module mem_ctrl ( 
    pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8,
    pi9, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17,
    pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26,
    pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35,
    pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44,
    pi45, pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53,
    pi54, pi55, pi56, pi57, pi58, pi59, pi60, pi61, pi62,
    pi63, pi64, pi65, pi66, pi67, pi68, pi69, pi70, pi71,
    pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79, pi80,
    pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88, pi89,
    pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97, pi98,
    pi99, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107,
    pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116,
    pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125,
    pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134,
    pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143,
    pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152,
    pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161,
    pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170,
    pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197,
    pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206,
    pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214, pi215,
    pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223, pi224,
    pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232, pi233,
    pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241, pi242,
    pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250, pi251,
    pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259, pi260,
    pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269,
    pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278,
    pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287,
    pi288, pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296,
    pi297, pi298, pi299, pi300, pi301, pi302, pi303, pi304, pi305,
    pi306, pi307, pi308, pi309, pi310, pi311, pi312, pi313, pi314,
    pi315, pi316, pi317, pi318, pi319, pi320, pi321, pi322, pi323,
    pi324, pi325, pi326, pi327, pi328, pi329, pi330, pi331, pi332,
    pi333, pi334, pi335, pi336, pi337, pi338, pi339, pi340, pi341,
    pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349, pi350,
    pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358, pi359,
    pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368,
    pi369, pi370, pi371, pi372, pi373, pi374, pi375, pi376, pi377,
    pi378, pi379, pi380, pi381, pi382, pi383, pi384, pi385, pi386,
    pi387, pi388, pi389, pi390, pi391, pi392, pi393, pi394, pi395,
    pi396, pi397, pi398, pi399, pi400, pi401, pi402, pi403, pi404,
    pi405, pi406, pi407, pi408, pi409, pi410, pi411, pi412, pi413,
    pi414, pi415, pi416, pi417, pi418, pi419, pi420, pi421, pi422,
    pi423, pi424, pi425, pi426, pi427, pi428, pi429, pi430, pi431,
    pi432, pi433, pi434, pi435, pi436, pi437, pi438, pi439, pi440,
    pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448, pi449,
    pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457, pi458,
    pi459, pi460, pi461, pi462, pi463, pi464, pi465, pi466, pi467,
    pi468, pi469, pi470, pi471, pi472, pi473, pi474, pi475, pi476,
    pi477, pi478, pi479, pi480, pi481, pi482, pi483, pi484, pi485,
    pi486, pi487, pi488, pi489, pi490, pi491, pi492, pi493, pi494,
    pi495, pi496, pi497, pi498, pi499, pi500, pi501, pi502, pi503,
    pi504, pi505, pi506, pi507, pi508, pi509, pi510, pi511, pi512,
    pi513, pi514, pi515, pi516, pi517, pi518, pi519, pi520, pi521,
    pi522, pi523, pi524, pi525, pi526, pi527, pi528, pi529, pi530,
    pi531, pi532, pi533, pi534, pi535, pi536, pi537, pi538, pi539,
    pi540, pi541, pi542, pi543, pi544, pi545, pi546, pi547, pi548,
    pi549, pi550, pi551, pi552, pi553, pi554, pi555, pi556, pi557,
    pi558, pi559, pi560, pi561, pi562, pi563, pi564, pi565, pi566,
    pi567, pi568, pi569, pi570, pi571, pi572, pi573, pi574, pi575,
    pi576, pi577, pi578, pi579, pi580, pi581, pi582, pi583, pi584,
    pi585, pi586, pi587, pi588, pi589, pi590, pi591, pi592, pi593,
    pi594, pi595, pi596, pi597, pi598, pi599, pi600, pi601, pi602,
    pi603, pi604, pi605, pi606, pi607, pi608, pi609, pi610, pi611,
    pi612, pi613, pi614, pi615, pi616, pi617, pi618, pi619, pi620,
    pi621, pi622, pi623, pi624, pi625, pi626, pi627, pi628, pi629,
    pi630, pi631, pi632, pi633, pi634, pi635, pi636, pi637, pi638,
    pi639, pi640, pi641, pi642, pi643, pi644, pi645, pi646, pi647,
    pi648, pi649, pi650, pi651, pi652, pi653, pi654, pi655, pi656,
    pi657, pi658, pi659, pi660, pi661, pi662, pi663, pi664, pi665,
    pi666, pi667, pi668, pi669, pi670, pi671, pi672, pi673, pi674,
    pi675, pi676, pi677, pi678, pi679, pi680, pi681, pi682, pi683,
    pi684, pi685, pi686, pi687, pi688, pi689, pi690, pi691, pi692,
    pi693, pi694, pi695, pi696, pi697, pi698, pi699, pi700, pi701,
    pi702, pi703, pi704, pi705, pi706, pi707, pi708, pi709, pi710,
    pi711, pi712, pi713, pi714, pi715, pi716, pi717, pi718, pi719,
    pi720, pi721, pi722, pi723, pi724, pi725, pi726, pi727, pi728,
    pi729, pi730, pi731, pi732, pi733, pi734, pi735, pi736, pi737,
    pi738, pi739, pi740, pi741, pi742, pi743, pi744, pi745, pi746,
    pi747, pi748, pi749, pi750, pi751, pi752, pi753, pi754, pi755,
    pi756, pi757, pi758, pi759, pi760, pi761, pi762, pi763, pi764,
    pi765, pi766, pi767, pi768, pi769, pi770, pi771, pi772, pi773,
    pi774, pi775, pi776, pi777, pi778, pi779, pi780, pi781, pi782,
    pi783, pi784, pi785, pi786, pi787, pi788, pi789, pi790, pi791,
    pi792, pi793, pi794, pi795, pi796, pi797, pi798, pi799, pi800,
    pi801, pi802, pi803, pi804, pi805, pi806, pi807, pi808, pi809,
    pi810, pi811, pi812, pi813, pi814, pi815, pi816, pi817, pi818,
    pi819, pi820, pi821, pi822, pi823, pi824, pi825, pi826, pi827,
    pi828, pi829, pi830, pi831, pi832, pi833, pi834, pi835, pi836,
    pi837, pi838, pi839, pi840, pi841, pi842, pi843, pi844, pi845,
    pi846, pi847, pi848, pi849, pi850, pi851, pi852, pi853, pi854,
    pi855, pi856, pi857, pi858, pi859, pi860, pi861, pi862, pi863,
    pi864, pi865, pi866, pi867, pi868, pi869, pi870, pi871, pi872,
    pi873, pi874, pi875, pi876, pi877, pi878, pi879, pi880, pi881,
    pi882, pi883, pi884, pi885, pi886, pi887, pi888, pi889, pi890,
    pi891, pi892, pi893, pi894, pi895, pi896, pi897, pi898, pi899,
    pi900, pi901, pi902, pi903, pi904, pi905, pi906, pi907, pi908,
    pi909, pi910, pi911, pi912, pi913, pi914, pi915, pi916, pi917,
    pi918, pi919, pi920, pi921, pi922, pi923, pi924, pi925, pi926,
    pi927, pi928, pi929, pi930, pi931, pi932, pi933, pi934, pi935,
    pi936, pi937, pi938, pi939, pi940, pi941, pi942, pi943, pi944,
    pi945, pi946, pi947, pi948, pi949, pi950, pi951, pi952, pi953,
    pi954, pi955, pi956, pi957, pi958, pi959, pi960, pi961, pi962,
    pi963, pi964, pi965, pi966, pi967, pi968, pi969, pi970, pi971,
    pi972, pi973, pi974, pi975, pi976, pi977, pi978, pi979, pi980,
    pi981, pi982, pi983, pi984, pi985, pi986, pi987, pi988, pi989,
    pi990, pi991, pi992, pi993, pi994, pi995, pi996, pi997, pi998,
    pi999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007,
    pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016,
    pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025,
    pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034,
    pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043,
    pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052,
    pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061,
    pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070,
    pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079,
    pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088,
    pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097,
    pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106,
    pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115,
    pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124,
    pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133,
    pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142,
    pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151,
    pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160,
    pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169,
    pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178,
    pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187,
    pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196,
    pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203,
    po0, po1, po2, po3, po4, po5, po6, po7, po8,
    po9, po10, po11, po12, po13, po14, po15, po16, po17,
    po18, po19, po20, po21, po22, po23, po24, po25, po26,
    po27, po28, po29, po30, po31, po32, po33, po34, po35,
    po36, po37, po38, po39, po40, po41, po42, po43, po44,
    po45, po46, po47, po48, po49, po50, po51, po52, po53,
    po54, po55, po56, po57, po58, po59, po60, po61, po62,
    po63, po64, po65, po66, po67, po68, po69, po70, po71,
    po72, po73, po74, po75, po76, po77, po78, po79, po80,
    po81, po82, po83, po84, po85, po86, po87, po88, po89,
    po90, po91, po92, po93, po94, po95, po96, po97, po98,
    po99, po100, po101, po102, po103, po104, po105, po106, po107,
    po108, po109, po110, po111, po112, po113, po114, po115, po116,
    po117, po118, po119, po120, po121, po122, po123, po124, po125,
    po126, po127, po128, po129, po130, po131, po132, po133, po134,
    po135, po136, po137, po138, po139, po140, po141, po142, po143,
    po144, po145, po146, po147, po148, po149, po150, po151, po152,
    po153, po154, po155, po156, po157, po158, po159, po160, po161,
    po162, po163, po164, po165, po166, po167, po168, po169, po170,
    po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188,
    po189, po190, po191, po192, po193, po194, po195, po196, po197,
    po198, po199, po200, po201, po202, po203, po204, po205, po206,
    po207, po208, po209, po210, po211, po212, po213, po214, po215,
    po216, po217, po218, po219, po220, po221, po222, po223, po224,
    po225, po226, po227, po228, po229, po230, po231, po232, po233,
    po234, po235, po236, po237, po238, po239, po240, po241, po242,
    po243, po244, po245, po246, po247, po248, po249, po250, po251,
    po252, po253, po254, po255, po256, po257, po258, po259, po260,
    po261, po262, po263, po264, po265, po266, po267, po268, po269,
    po270, po271, po272, po273, po274, po275, po276, po277, po278,
    po279, po280, po281, po282, po283, po284, po285, po286, po287,
    po288, po289, po290, po291, po292, po293, po294, po295, po296,
    po297, po298, po299, po300, po301, po302, po303, po304, po305,
    po306, po307, po308, po309, po310, po311, po312, po313, po314,
    po315, po316, po317, po318, po319, po320, po321, po322, po323,
    po324, po325, po326, po327, po328, po329, po330, po331, po332,
    po333, po334, po335, po336, po337, po338, po339, po340, po341,
    po342, po343, po344, po345, po346, po347, po348, po349, po350,
    po351, po352, po353, po354, po355, po356, po357, po358, po359,
    po360, po361, po362, po363, po364, po365, po366, po367, po368,
    po369, po370, po371, po372, po373, po374, po375, po376, po377,
    po378, po379, po380, po381, po382, po383, po384, po385, po386,
    po387, po388, po389, po390, po391, po392, po393, po394, po395,
    po396, po397, po398, po399, po400, po401, po402, po403, po404,
    po405, po406, po407, po408, po409, po410, po411, po412, po413,
    po414, po415, po416, po417, po418, po419, po420, po421, po422,
    po423, po424, po425, po426, po427, po428, po429, po430, po431,
    po432, po433, po434, po435, po436, po437, po438, po439, po440,
    po441, po442, po443, po444, po445, po446, po447, po448, po449,
    po450, po451, po452, po453, po454, po455, po456, po457, po458,
    po459, po460, po461, po462, po463, po464, po465, po466, po467,
    po468, po469, po470, po471, po472, po473, po474, po475, po476,
    po477, po478, po479, po480, po481, po482, po483, po484, po485,
    po486, po487, po488, po489, po490, po491, po492, po493, po494,
    po495, po496, po497, po498, po499, po500, po501, po502, po503,
    po504, po505, po506, po507, po508, po509, po510, po511, po512,
    po513, po514, po515, po516, po517, po518, po519, po520, po521,
    po522, po523, po524, po525, po526, po527, po528, po529, po530,
    po531, po532, po533, po534, po535, po536, po537, po538, po539,
    po540, po541, po542, po543, po544, po545, po546, po547, po548,
    po549, po550, po551, po552, po553, po554, po555, po556, po557,
    po558, po559, po560, po561, po562, po563, po564, po565, po566,
    po567, po568, po569, po570, po571, po572, po573, po574, po575,
    po576, po577, po578, po579, po580, po581, po582, po583, po584,
    po585, po586, po587, po588, po589, po590, po591, po592, po593,
    po594, po595, po596, po597, po598, po599, po600, po601, po602,
    po603, po604, po605, po606, po607, po608, po609, po610, po611,
    po612, po613, po614, po615, po616, po617, po618, po619, po620,
    po621, po622, po623, po624, po625, po626, po627, po628, po629,
    po630, po631, po632, po633, po634, po635, po636, po637, po638,
    po639, po640, po641, po642, po643, po644, po645, po646, po647,
    po648, po649, po650, po651, po652, po653, po654, po655, po656,
    po657, po658, po659, po660, po661, po662, po663, po664, po665,
    po666, po667, po668, po669, po670, po671, po672, po673, po674,
    po675, po676, po677, po678, po679, po680, po681, po682, po683,
    po684, po685, po686, po687, po688, po689, po690, po691, po692,
    po693, po694, po695, po696, po697, po698, po699, po700, po701,
    po702, po703, po704, po705, po706, po707, po708, po709, po710,
    po711, po712, po713, po714, po715, po716, po717, po718, po719,
    po720, po721, po722, po723, po724, po725, po726, po727, po728,
    po729, po730, po731, po732, po733, po734, po735, po736, po737,
    po738, po739, po740, po741, po742, po743, po744, po745, po746,
    po747, po748, po749, po750, po751, po752, po753, po754, po755,
    po756, po757, po758, po759, po760, po761, po762, po763, po764,
    po765, po766, po767, po768, po769, po770, po771, po772, po773,
    po774, po775, po776, po777, po778, po779, po780, po781, po782,
    po783, po784, po785, po786, po787, po788, po789, po790, po791,
    po792, po793, po794, po795, po796, po797, po798, po799, po800,
    po801, po802, po803, po804, po805, po806, po807, po808, po809,
    po810, po811, po812, po813, po814, po815, po816, po817, po818,
    po819, po820, po821, po822, po823, po824, po825, po826, po827,
    po828, po829, po830, po831, po832, po833, po834, po835, po836,
    po837, po838, po839, po840, po841, po842, po843, po844, po845,
    po846, po847, po848, po849, po850, po851, po852, po853, po854,
    po855, po856, po857, po858, po859, po860, po861, po862, po863,
    po864, po865, po866, po867, po868, po869, po870, po871, po872,
    po873, po874, po875, po876, po877, po878, po879, po880, po881,
    po882, po883, po884, po885, po886, po887, po888, po889, po890,
    po891, po892, po893, po894, po895, po896, po897, po898, po899,
    po900, po901, po902, po903, po904, po905, po906, po907, po908,
    po909, po910, po911, po912, po913, po914, po915, po916, po917,
    po918, po919, po920, po921, po922, po923, po924, po925, po926,
    po927, po928, po929, po930, po931, po932, po933, po934, po935,
    po936, po937, po938, po939, po940, po941, po942, po943, po944,
    po945, po946, po947, po948, po949, po950, po951, po952, po953,
    po954, po955, po956, po957, po958, po959, po960, po961, po962,
    po963, po964, po965, po966, po967, po968, po969, po970, po971,
    po972, po973, po974, po975, po976, po977, po978, po979, po980,
    po981, po982, po983, po984, po985, po986, po987, po988, po989,
    po990, po991, po992, po993, po994, po995, po996, po997, po998,
    po999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007,
    po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016,
    po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025,
    po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034,
    po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043,
    po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052,
    po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061,
    po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070,
    po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079,
    po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088,
    po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097,
    po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106,
    po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115,
    po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124,
    po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133,
    po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142,
    po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151,
    po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160,
    po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169,
    po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178,
    po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187,
    po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196,
    po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205,
    po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214,
    po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223,
    po1224, po1225, po1226, po1227, po1228, po1229, po1230  );
  input  pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7,
    pi8, pi9, pi10, pi11, pi12, pi13, pi14, pi15, pi16,
    pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25,
    pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34,
    pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43,
    pi44, pi45, pi46, pi47, pi48, pi49, pi50, pi51, pi52,
    pi53, pi54, pi55, pi56, pi57, pi58, pi59, pi60, pi61,
    pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69, pi70,
    pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79,
    pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88,
    pi89, pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97,
    pi98, pi99, pi100, pi101, pi102, pi103, pi104, pi105, pi106,
    pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115,
    pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124,
    pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133,
    pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142,
    pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151,
    pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160,
    pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187,
    pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196,
    pi197, pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205,
    pi206, pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214,
    pi215, pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223,
    pi224, pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232,
    pi233, pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241,
    pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250,
    pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259,
    pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268,
    pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277,
    pi278, pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286,
    pi287, pi288, pi289, pi290, pi291, pi292, pi293, pi294, pi295,
    pi296, pi297, pi298, pi299, pi300, pi301, pi302, pi303, pi304,
    pi305, pi306, pi307, pi308, pi309, pi310, pi311, pi312, pi313,
    pi314, pi315, pi316, pi317, pi318, pi319, pi320, pi321, pi322,
    pi323, pi324, pi325, pi326, pi327, pi328, pi329, pi330, pi331,
    pi332, pi333, pi334, pi335, pi336, pi337, pi338, pi339, pi340,
    pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349,
    pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358,
    pi359, pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367,
    pi368, pi369, pi370, pi371, pi372, pi373, pi374, pi375, pi376,
    pi377, pi378, pi379, pi380, pi381, pi382, pi383, pi384, pi385,
    pi386, pi387, pi388, pi389, pi390, pi391, pi392, pi393, pi394,
    pi395, pi396, pi397, pi398, pi399, pi400, pi401, pi402, pi403,
    pi404, pi405, pi406, pi407, pi408, pi409, pi410, pi411, pi412,
    pi413, pi414, pi415, pi416, pi417, pi418, pi419, pi420, pi421,
    pi422, pi423, pi424, pi425, pi426, pi427, pi428, pi429, pi430,
    pi431, pi432, pi433, pi434, pi435, pi436, pi437, pi438, pi439,
    pi440, pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448,
    pi449, pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457,
    pi458, pi459, pi460, pi461, pi462, pi463, pi464, pi465, pi466,
    pi467, pi468, pi469, pi470, pi471, pi472, pi473, pi474, pi475,
    pi476, pi477, pi478, pi479, pi480, pi481, pi482, pi483, pi484,
    pi485, pi486, pi487, pi488, pi489, pi490, pi491, pi492, pi493,
    pi494, pi495, pi496, pi497, pi498, pi499, pi500, pi501, pi502,
    pi503, pi504, pi505, pi506, pi507, pi508, pi509, pi510, pi511,
    pi512, pi513, pi514, pi515, pi516, pi517, pi518, pi519, pi520,
    pi521, pi522, pi523, pi524, pi525, pi526, pi527, pi528, pi529,
    pi530, pi531, pi532, pi533, pi534, pi535, pi536, pi537, pi538,
    pi539, pi540, pi541, pi542, pi543, pi544, pi545, pi546, pi547,
    pi548, pi549, pi550, pi551, pi552, pi553, pi554, pi555, pi556,
    pi557, pi558, pi559, pi560, pi561, pi562, pi563, pi564, pi565,
    pi566, pi567, pi568, pi569, pi570, pi571, pi572, pi573, pi574,
    pi575, pi576, pi577, pi578, pi579, pi580, pi581, pi582, pi583,
    pi584, pi585, pi586, pi587, pi588, pi589, pi590, pi591, pi592,
    pi593, pi594, pi595, pi596, pi597, pi598, pi599, pi600, pi601,
    pi602, pi603, pi604, pi605, pi606, pi607, pi608, pi609, pi610,
    pi611, pi612, pi613, pi614, pi615, pi616, pi617, pi618, pi619,
    pi620, pi621, pi622, pi623, pi624, pi625, pi626, pi627, pi628,
    pi629, pi630, pi631, pi632, pi633, pi634, pi635, pi636, pi637,
    pi638, pi639, pi640, pi641, pi642, pi643, pi644, pi645, pi646,
    pi647, pi648, pi649, pi650, pi651, pi652, pi653, pi654, pi655,
    pi656, pi657, pi658, pi659, pi660, pi661, pi662, pi663, pi664,
    pi665, pi666, pi667, pi668, pi669, pi670, pi671, pi672, pi673,
    pi674, pi675, pi676, pi677, pi678, pi679, pi680, pi681, pi682,
    pi683, pi684, pi685, pi686, pi687, pi688, pi689, pi690, pi691,
    pi692, pi693, pi694, pi695, pi696, pi697, pi698, pi699, pi700,
    pi701, pi702, pi703, pi704, pi705, pi706, pi707, pi708, pi709,
    pi710, pi711, pi712, pi713, pi714, pi715, pi716, pi717, pi718,
    pi719, pi720, pi721, pi722, pi723, pi724, pi725, pi726, pi727,
    pi728, pi729, pi730, pi731, pi732, pi733, pi734, pi735, pi736,
    pi737, pi738, pi739, pi740, pi741, pi742, pi743, pi744, pi745,
    pi746, pi747, pi748, pi749, pi750, pi751, pi752, pi753, pi754,
    pi755, pi756, pi757, pi758, pi759, pi760, pi761, pi762, pi763,
    pi764, pi765, pi766, pi767, pi768, pi769, pi770, pi771, pi772,
    pi773, pi774, pi775, pi776, pi777, pi778, pi779, pi780, pi781,
    pi782, pi783, pi784, pi785, pi786, pi787, pi788, pi789, pi790,
    pi791, pi792, pi793, pi794, pi795, pi796, pi797, pi798, pi799,
    pi800, pi801, pi802, pi803, pi804, pi805, pi806, pi807, pi808,
    pi809, pi810, pi811, pi812, pi813, pi814, pi815, pi816, pi817,
    pi818, pi819, pi820, pi821, pi822, pi823, pi824, pi825, pi826,
    pi827, pi828, pi829, pi830, pi831, pi832, pi833, pi834, pi835,
    pi836, pi837, pi838, pi839, pi840, pi841, pi842, pi843, pi844,
    pi845, pi846, pi847, pi848, pi849, pi850, pi851, pi852, pi853,
    pi854, pi855, pi856, pi857, pi858, pi859, pi860, pi861, pi862,
    pi863, pi864, pi865, pi866, pi867, pi868, pi869, pi870, pi871,
    pi872, pi873, pi874, pi875, pi876, pi877, pi878, pi879, pi880,
    pi881, pi882, pi883, pi884, pi885, pi886, pi887, pi888, pi889,
    pi890, pi891, pi892, pi893, pi894, pi895, pi896, pi897, pi898,
    pi899, pi900, pi901, pi902, pi903, pi904, pi905, pi906, pi907,
    pi908, pi909, pi910, pi911, pi912, pi913, pi914, pi915, pi916,
    pi917, pi918, pi919, pi920, pi921, pi922, pi923, pi924, pi925,
    pi926, pi927, pi928, pi929, pi930, pi931, pi932, pi933, pi934,
    pi935, pi936, pi937, pi938, pi939, pi940, pi941, pi942, pi943,
    pi944, pi945, pi946, pi947, pi948, pi949, pi950, pi951, pi952,
    pi953, pi954, pi955, pi956, pi957, pi958, pi959, pi960, pi961,
    pi962, pi963, pi964, pi965, pi966, pi967, pi968, pi969, pi970,
    pi971, pi972, pi973, pi974, pi975, pi976, pi977, pi978, pi979,
    pi980, pi981, pi982, pi983, pi984, pi985, pi986, pi987, pi988,
    pi989, pi990, pi991, pi992, pi993, pi994, pi995, pi996, pi997,
    pi998, pi999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006,
    pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015,
    pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024,
    pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033,
    pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042,
    pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051,
    pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060,
    pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069,
    pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078,
    pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087,
    pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096,
    pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105,
    pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114,
    pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123,
    pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132,
    pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141,
    pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150,
    pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159,
    pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168,
    pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177,
    pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186,
    pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195,
    pi1196, pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203;
  output po0, po1, po2, po3, po4, po5, po6, po7,
    po8, po9, po10, po11, po12, po13, po14, po15, po16,
    po17, po18, po19, po20, po21, po22, po23, po24, po25,
    po26, po27, po28, po29, po30, po31, po32, po33, po34,
    po35, po36, po37, po38, po39, po40, po41, po42, po43,
    po44, po45, po46, po47, po48, po49, po50, po51, po52,
    po53, po54, po55, po56, po57, po58, po59, po60, po61,
    po62, po63, po64, po65, po66, po67, po68, po69, po70,
    po71, po72, po73, po74, po75, po76, po77, po78, po79,
    po80, po81, po82, po83, po84, po85, po86, po87, po88,
    po89, po90, po91, po92, po93, po94, po95, po96, po97,
    po98, po99, po100, po101, po102, po103, po104, po105, po106,
    po107, po108, po109, po110, po111, po112, po113, po114, po115,
    po116, po117, po118, po119, po120, po121, po122, po123, po124,
    po125, po126, po127, po128, po129, po130, po131, po132, po133,
    po134, po135, po136, po137, po138, po139, po140, po141, po142,
    po143, po144, po145, po146, po147, po148, po149, po150, po151,
    po152, po153, po154, po155, po156, po157, po158, po159, po160,
    po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178,
    po179, po180, po181, po182, po183, po184, po185, po186, po187,
    po188, po189, po190, po191, po192, po193, po194, po195, po196,
    po197, po198, po199, po200, po201, po202, po203, po204, po205,
    po206, po207, po208, po209, po210, po211, po212, po213, po214,
    po215, po216, po217, po218, po219, po220, po221, po222, po223,
    po224, po225, po226, po227, po228, po229, po230, po231, po232,
    po233, po234, po235, po236, po237, po238, po239, po240, po241,
    po242, po243, po244, po245, po246, po247, po248, po249, po250,
    po251, po252, po253, po254, po255, po256, po257, po258, po259,
    po260, po261, po262, po263, po264, po265, po266, po267, po268,
    po269, po270, po271, po272, po273, po274, po275, po276, po277,
    po278, po279, po280, po281, po282, po283, po284, po285, po286,
    po287, po288, po289, po290, po291, po292, po293, po294, po295,
    po296, po297, po298, po299, po300, po301, po302, po303, po304,
    po305, po306, po307, po308, po309, po310, po311, po312, po313,
    po314, po315, po316, po317, po318, po319, po320, po321, po322,
    po323, po324, po325, po326, po327, po328, po329, po330, po331,
    po332, po333, po334, po335, po336, po337, po338, po339, po340,
    po341, po342, po343, po344, po345, po346, po347, po348, po349,
    po350, po351, po352, po353, po354, po355, po356, po357, po358,
    po359, po360, po361, po362, po363, po364, po365, po366, po367,
    po368, po369, po370, po371, po372, po373, po374, po375, po376,
    po377, po378, po379, po380, po381, po382, po383, po384, po385,
    po386, po387, po388, po389, po390, po391, po392, po393, po394,
    po395, po396, po397, po398, po399, po400, po401, po402, po403,
    po404, po405, po406, po407, po408, po409, po410, po411, po412,
    po413, po414, po415, po416, po417, po418, po419, po420, po421,
    po422, po423, po424, po425, po426, po427, po428, po429, po430,
    po431, po432, po433, po434, po435, po436, po437, po438, po439,
    po440, po441, po442, po443, po444, po445, po446, po447, po448,
    po449, po450, po451, po452, po453, po454, po455, po456, po457,
    po458, po459, po460, po461, po462, po463, po464, po465, po466,
    po467, po468, po469, po470, po471, po472, po473, po474, po475,
    po476, po477, po478, po479, po480, po481, po482, po483, po484,
    po485, po486, po487, po488, po489, po490, po491, po492, po493,
    po494, po495, po496, po497, po498, po499, po500, po501, po502,
    po503, po504, po505, po506, po507, po508, po509, po510, po511,
    po512, po513, po514, po515, po516, po517, po518, po519, po520,
    po521, po522, po523, po524, po525, po526, po527, po528, po529,
    po530, po531, po532, po533, po534, po535, po536, po537, po538,
    po539, po540, po541, po542, po543, po544, po545, po546, po547,
    po548, po549, po550, po551, po552, po553, po554, po555, po556,
    po557, po558, po559, po560, po561, po562, po563, po564, po565,
    po566, po567, po568, po569, po570, po571, po572, po573, po574,
    po575, po576, po577, po578, po579, po580, po581, po582, po583,
    po584, po585, po586, po587, po588, po589, po590, po591, po592,
    po593, po594, po595, po596, po597, po598, po599, po600, po601,
    po602, po603, po604, po605, po606, po607, po608, po609, po610,
    po611, po612, po613, po614, po615, po616, po617, po618, po619,
    po620, po621, po622, po623, po624, po625, po626, po627, po628,
    po629, po630, po631, po632, po633, po634, po635, po636, po637,
    po638, po639, po640, po641, po642, po643, po644, po645, po646,
    po647, po648, po649, po650, po651, po652, po653, po654, po655,
    po656, po657, po658, po659, po660, po661, po662, po663, po664,
    po665, po666, po667, po668, po669, po670, po671, po672, po673,
    po674, po675, po676, po677, po678, po679, po680, po681, po682,
    po683, po684, po685, po686, po687, po688, po689, po690, po691,
    po692, po693, po694, po695, po696, po697, po698, po699, po700,
    po701, po702, po703, po704, po705, po706, po707, po708, po709,
    po710, po711, po712, po713, po714, po715, po716, po717, po718,
    po719, po720, po721, po722, po723, po724, po725, po726, po727,
    po728, po729, po730, po731, po732, po733, po734, po735, po736,
    po737, po738, po739, po740, po741, po742, po743, po744, po745,
    po746, po747, po748, po749, po750, po751, po752, po753, po754,
    po755, po756, po757, po758, po759, po760, po761, po762, po763,
    po764, po765, po766, po767, po768, po769, po770, po771, po772,
    po773, po774, po775, po776, po777, po778, po779, po780, po781,
    po782, po783, po784, po785, po786, po787, po788, po789, po790,
    po791, po792, po793, po794, po795, po796, po797, po798, po799,
    po800, po801, po802, po803, po804, po805, po806, po807, po808,
    po809, po810, po811, po812, po813, po814, po815, po816, po817,
    po818, po819, po820, po821, po822, po823, po824, po825, po826,
    po827, po828, po829, po830, po831, po832, po833, po834, po835,
    po836, po837, po838, po839, po840, po841, po842, po843, po844,
    po845, po846, po847, po848, po849, po850, po851, po852, po853,
    po854, po855, po856, po857, po858, po859, po860, po861, po862,
    po863, po864, po865, po866, po867, po868, po869, po870, po871,
    po872, po873, po874, po875, po876, po877, po878, po879, po880,
    po881, po882, po883, po884, po885, po886, po887, po888, po889,
    po890, po891, po892, po893, po894, po895, po896, po897, po898,
    po899, po900, po901, po902, po903, po904, po905, po906, po907,
    po908, po909, po910, po911, po912, po913, po914, po915, po916,
    po917, po918, po919, po920, po921, po922, po923, po924, po925,
    po926, po927, po928, po929, po930, po931, po932, po933, po934,
    po935, po936, po937, po938, po939, po940, po941, po942, po943,
    po944, po945, po946, po947, po948, po949, po950, po951, po952,
    po953, po954, po955, po956, po957, po958, po959, po960, po961,
    po962, po963, po964, po965, po966, po967, po968, po969, po970,
    po971, po972, po973, po974, po975, po976, po977, po978, po979,
    po980, po981, po982, po983, po984, po985, po986, po987, po988,
    po989, po990, po991, po992, po993, po994, po995, po996, po997,
    po998, po999, po1000, po1001, po1002, po1003, po1004, po1005, po1006,
    po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015,
    po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024,
    po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033,
    po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042,
    po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051,
    po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060,
    po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069,
    po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078,
    po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087,
    po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096,
    po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105,
    po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114,
    po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123,
    po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132,
    po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141,
    po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150,
    po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159,
    po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168,
    po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177,
    po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186,
    po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195,
    po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204,
    po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213,
    po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222,
    po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230;
  wire n2437, n2438, n2439, n2440, n2441, n2442,
    n2443, n2444, n2445, n2446, n2447, n2448,
    n2449, n2450, n2451, n2452, n2453, n2454,
    n2455, n2456, n2457, n2458, n2459, n2460,
    n2461, n2462, n2463, n2464, n2465, n2466,
    n2467, n2468, n2469, n2470, n2471, n2472,
    n2473, n2474, n2475, n2476, n2477, n2478,
    n2479, n2480, n2481, n2482, n2483, n2484,
    n2485, n2486, n2487, n2488, n2489, n2490,
    n2491, n2492, n2493, n2494, n2495, n2496,
    n2497, n2498, n2499, n2500, n2501, n2502,
    n2503, n2504, n2505, n2506, n2507, n2508,
    n2509, n2510, n2511, n2512, n2513, n2514,
    n2515, n2516, n2517, n2518, n2519, n2520,
    n2521, n2522, n2523, n2524, n2525, n2526,
    n2527, n2528, n2529, n2530, n2531, n2532,
    n2533, n2534, n2535, n2536, n2537, n2538,
    n2539, n2540, n2541, n2542, n2543, n2544,
    n2545, n2546, n2547, n2548, n2549, n2550,
    n2551, n2552, n2553, n2554, n2555, n2556,
    n2557, n2558, n2559, n2560, n2561, n2562,
    n2563, n2564, n2565, n2566, n2567, n2568,
    n2569, n2570, n2571, n2572, n2573, n2574,
    n2575, n2576, n2577, n2578, n2579, n2580,
    n2581, n2582, n2583, n2584, n2585, n2586,
    n2587, n2588, n2589, n2590, n2591, n2592,
    n2593, n2594, n2595, n2596, n2597, n2598,
    n2599, n2600, n2601, n2602, n2603, n2604,
    n2605, n2606, n2607, n2608, n2609, n2610,
    n2611, n2612, n2613, n2614, n2615, n2616,
    n2617, n2618, n2619, n2620, n2621, n2622,
    n2623, n2624, n2625, n2626, n2627, n2628,
    n2629, n2630, n2631, n2632, n2633, n2634,
    n2635, n2636, n2637, n2638, n2639, n2640,
    n2641, n2642, n2643, n2644, n2645, n2646,
    n2647, n2648, n2649, n2650, n2651, n2652,
    n2653, n2654, n2655, n2656, n2657, n2658,
    n2659, n2660, n2661, n2662, n2663, n2664,
    n2665, n2666, n2667, n2668, n2669, n2670,
    n2671, n2672, n2673, n2674, n2675, n2676,
    n2677, n2678, n2679, n2680, n2681, n2682,
    n2683, n2684, n2685, n2686, n2687, n2688,
    n2689, n2690, n2691, n2692, n2693, n2694,
    n2695, n2696, n2697, n2698, n2699, n2700,
    n2701, n2702, n2703, n2704, n2705, n2706,
    n2707, n2708, n2709, n2710, n2711, n2712,
    n2713, n2714, n2715, n2716, n2717, n2718,
    n2719, n2720, n2721, n2722, n2723, n2724,
    n2725, n2726, n2727, n2728, n2729, n2730,
    n2731, n2732, n2733, n2734, n2735, n2736,
    n2737, n2738, n2739, n2740, n2741, n2742,
    n2743, n2744, n2745, n2746, n2747, n2748,
    n2749, n2750, n2751, n2752, n2753, n2754,
    n2755, n2756, n2757, n2758, n2759, n2760,
    n2761, n2762, n2763, n2764, n2765, n2766,
    n2767, n2768, n2769, n2770, n2771, n2772,
    n2773, n2774, n2775, n2776, n2777, n2778,
    n2779, n2780, n2781, n2782, n2783, n2784,
    n2785, n2786, n2787, n2788, n2789, n2790,
    n2791, n2792, n2793, n2794, n2795, n2796,
    n2797, n2798, n2799, n2800, n2801, n2802,
    n2803, n2804, n2805, n2806, n2807, n2808,
    n2809, n2810, n2811, n2812, n2813, n2814,
    n2815, n2816, n2817, n2818, n2819, n2820,
    n2821, n2822, n2823, n2824, n2825, n2826,
    n2827, n2828, n2829, n2830, n2831, n2832,
    n2833, n2834, n2835, n2836, n2837, n2838,
    n2839, n2840, n2841, n2842, n2843, n2844,
    n2845, n2846, n2847, n2848, n2849, n2850,
    n2851, n2852, n2853, n2854, n2855, n2856,
    n2857, n2858, n2859, n2860, n2861, n2862,
    n2863, n2864, n2865, n2866, n2867, n2868,
    n2869, n2870, n2871, n2872, n2873, n2874,
    n2875, n2876, n2877, n2878, n2879, n2880,
    n2881, n2882, n2883, n2884, n2885, n2886,
    n2887, n2888, n2889, n2890, n2891, n2892,
    n2893, n2894, n2895, n2896, n2897, n2898,
    n2899, n2900, n2901, n2902, n2903, n2904,
    n2905, n2906, n2907, n2908, n2909, n2910,
    n2911, n2912, n2913, n2914, n2915, n2916,
    n2917, n2918, n2919, n2920, n2921, n2922,
    n2923, n2924, n2925, n2926, n2927, n2928,
    n2929, n2930, n2931, n2932, n2933, n2934,
    n2935, n2936, n2937, n2938, n2939, n2940,
    n2941, n2942, n2943, n2944, n2945, n2946,
    n2947, n2948, n2949, n2950, n2951, n2952,
    n2953, n2954, n2955, n2956, n2957, n2958,
    n2959, n2960, n2961, n2962, n2963, n2964,
    n2965, n2966, n2967, n2968, n2969, n2970,
    n2971, n2972, n2973, n2974, n2975, n2976,
    n2977, n2978, n2979, n2980, n2981, n2982,
    n2983, n2984, n2985, n2986, n2987, n2988,
    n2989, n2990, n2991, n2992, n2993, n2994,
    n2995, n2996, n2997, n2998, n2999, n3000,
    n3001, n3002, n3003, n3004, n3005, n3006,
    n3007, n3008, n3009, n3010, n3011, n3012,
    n3013, n3014, n3015, n3016, n3017, n3018,
    n3019, n3020, n3021, n3022, n3023, n3024,
    n3025, n3026, n3027, n3028, n3029, n3030,
    n3031, n3032, n3033, n3034, n3035, n3036,
    n3037, n3038, n3039, n3040, n3041, n3042,
    n3043, n3044, n3045, n3046, n3047, n3048,
    n3049, n3050, n3051, n3052, n3053, n3054,
    n3055, n3056, n3057, n3058, n3059, n3060,
    n3061, n3062, n3063, n3064, n3065, n3066,
    n3067, n3068, n3069, n3070, n3071, n3072,
    n3073, n3074, n3075, n3076, n3077, n3078,
    n3079, n3080, n3081, n3082, n3083, n3084,
    n3085, n3086, n3087, n3088, n3089, n3090,
    n3091, n3092, n3093, n3094, n3095, n3096,
    n3097, n3098, n3099, n3100, n3101, n3102,
    n3103, n3104, n3105, n3106, n3107, n3108,
    n3109, n3110, n3111, n3112, n3113, n3114,
    n3115, n3116, n3117, n3118, n3119, n3120,
    n3121, n3122, n3123, n3124, n3125, n3126,
    n3127, n3128, n3129, n3130, n3131, n3132,
    n3133, n3134, n3135, n3136, n3137, n3138,
    n3139, n3140, n3141, n3142, n3143, n3144,
    n3145, n3146, n3147, n3148, n3149, n3150,
    n3151, n3152, n3153, n3154, n3155, n3156,
    n3157, n3158, n3159, n3160, n3161, n3162,
    n3163, n3164, n3165, n3166, n3167, n3168,
    n3169, n3170, n3171, n3172, n3173, n3174,
    n3175, n3176, n3177, n3178, n3179, n3180,
    n3181, n3182, n3183, n3184, n3185, n3186,
    n3187, n3188, n3189, n3190, n3191, n3192,
    n3193, n3194, n3195, n3196, n3197, n3198,
    n3199, n3200, n3201, n3202, n3203, n3204,
    n3205, n3206, n3207, n3208, n3209, n3210,
    n3211, n3212, n3213, n3214, n3215, n3216,
    n3217, n3218, n3219, n3220, n3221, n3222,
    n3223, n3224, n3225, n3226, n3227, n3228,
    n3229, n3230, n3231, n3232, n3233, n3234,
    n3235, n3236, n3237, n3238, n3239, n3240,
    n3241, n3242, n3243, n3244, n3245, n3246,
    n3247, n3248, n3249, n3250, n3251, n3252,
    n3253, n3254, n3255, n3256, n3257, n3258,
    n3259, n3260, n3261, n3262, n3263, n3264,
    n3265, n3266, n3267, n3268, n3269, n3270,
    n3271, n3272, n3273, n3274, n3275, n3276,
    n3277, n3278, n3279, n3280, n3281, n3282,
    n3283, n3284, n3285, n3286, n3287, n3288,
    n3289, n3290, n3291, n3292, n3293, n3294,
    n3295, n3296, n3297, n3298, n3299, n3300,
    n3301, n3302, n3303, n3305, n3306, n3307,
    n3308, n3309, n3310, n3311, n3312, n3313,
    n3314, n3315, n3316, n3317, n3318, n3319,
    n3320, n3321, n3322, n3323, n3324, n3325,
    n3326, n3327, n3328, n3329, n3330, n3331,
    n3332, n3333, n3334, n3335, n3336, n3337,
    n3338, n3339, n3340, n3341, n3342, n3343,
    n3344, n3345, n3346, n3347, n3348, n3349,
    n3350, n3351, n3352, n3353, n3354, n3355,
    n3356, n3357, n3358, n3359, n3360, n3361,
    n3362, n3363, n3364, n3365, n3366, n3367,
    n3368, n3369, n3370, n3371, n3372, n3373,
    n3374, n3375, n3376, n3377, n3378, n3379,
    n3380, n3381, n3382, n3383, n3384, n3385,
    n3386, n3387, n3388, n3389, n3390, n3391,
    n3392, n3393, n3394, n3395, n3396, n3397,
    n3398, n3399, n3400, n3401, n3402, n3403,
    n3404, n3405, n3406, n3407, n3408, n3409,
    n3410, n3411, n3412, n3413, n3414, n3415,
    n3416, n3417, n3418, n3419, n3420, n3421,
    n3422, n3423, n3424, n3425, n3426, n3427,
    n3428, n3429, n3430, n3431, n3432, n3433,
    n3434, n3435, n3436, n3437, n3438, n3439,
    n3440, n3441, n3442, n3443, n3444, n3445,
    n3446, n3447, n3448, n3449, n3450, n3451,
    n3452, n3453, n3454, n3455, n3456, n3457,
    n3458, n3459, n3460, n3461, n3462, n3463,
    n3464, n3465, n3466, n3467, n3468, n3469,
    n3470, n3471, n3472, n3473, n3474, n3475,
    n3476, n3477, n3478, n3479, n3480, n3481,
    n3482, n3483, n3484, n3485, n3486, n3487,
    n3488, n3489, n3490, n3491, n3492, n3493,
    n3494, n3495, n3496, n3497, n3498, n3499,
    n3500, n3501, n3502, n3503, n3504, n3505,
    n3506, n3507, n3508, n3509, n3510, n3511,
    n3512, n3513, n3514, n3515, n3516, n3517,
    n3518, n3519, n3520, n3521, n3522, n3523,
    n3524, n3525, n3526, n3527, n3528, n3529,
    n3530, n3531, n3532, n3533, n3534, n3535,
    n3537, n3538, n3539, n3540, n3541, n3542,
    n3543, n3544, n3545, n3546, n3547, n3548,
    n3549, n3550, n3551, n3552, n3553, n3554,
    n3555, n3556, n3557, n3558, n3559, n3560,
    n3561, n3562, n3563, n3564, n3565, n3566,
    n3567, n3568, n3569, n3570, n3571, n3572,
    n3573, n3574, n3575, n3576, n3577, n3578,
    n3579, n3580, n3581, n3582, n3583, n3584,
    n3585, n3586, n3587, n3588, n3589, n3590,
    n3591, n3592, n3593, n3594, n3595, n3596,
    n3597, n3598, n3599, n3600, n3601, n3602,
    n3603, n3604, n3605, n3606, n3607, n3608,
    n3609, n3610, n3611, n3612, n3613, n3614,
    n3615, n3616, n3617, n3618, n3619, n3620,
    n3621, n3622, n3623, n3624, n3625, n3626,
    n3627, n3628, n3629, n3630, n3631, n3632,
    n3633, n3634, n3635, n3636, n3637, n3638,
    n3639, n3640, n3641, n3642, n3643, n3644,
    n3645, n3646, n3647, n3648, n3649, n3650,
    n3651, n3652, n3653, n3654, n3655, n3656,
    n3657, n3658, n3659, n3660, n3661, n3662,
    n3663, n3664, n3665, n3666, n3667, n3668,
    n3669, n3670, n3671, n3672, n3673, n3674,
    n3675, n3676, n3677, n3678, n3679, n3680,
    n3681, n3682, n3683, n3684, n3685, n3686,
    n3687, n3688, n3689, n3690, n3691, n3692,
    n3693, n3694, n3695, n3696, n3697, n3698,
    n3699, n3700, n3701, n3702, n3703, n3704,
    n3705, n3706, n3708, n3709, n3710, n3711,
    n3712, n3713, n3714, n3715, n3716, n3717,
    n3718, n3719, n3720, n3721, n3722, n3723,
    n3724, n3725, n3726, n3727, n3728, n3729,
    n3730, n3731, n3732, n3733, n3734, n3735,
    n3736, n3737, n3738, n3739, n3740, n3741,
    n3742, n3743, n3744, n3745, n3746, n3747,
    n3748, n3749, n3750, n3751, n3752, n3753,
    n3754, n3755, n3756, n3757, n3758, n3759,
    n3760, n3761, n3762, n3763, n3764, n3765,
    n3766, n3767, n3768, n3769, n3770, n3771,
    n3772, n3773, n3774, n3775, n3776, n3777,
    n3778, n3779, n3780, n3781, n3782, n3783,
    n3784, n3785, n3786, n3787, n3788, n3789,
    n3790, n3791, n3792, n3793, n3794, n3795,
    n3796, n3797, n3798, n3799, n3800, n3801,
    n3802, n3803, n3804, n3805, n3806, n3807,
    n3808, n3809, n3810, n3811, n3812, n3813,
    n3814, n3815, n3816, n3817, n3818, n3819,
    n3820, n3821, n3822, n3823, n3824, n3825,
    n3826, n3827, n3828, n3829, n3830, n3831,
    n3832, n3833, n3834, n3835, n3836, n3837,
    n3838, n3839, n3840, n3841, n3842, n3843,
    n3844, n3845, n3846, n3847, n3848, n3849,
    n3850, n3851, n3852, n3853, n3854, n3855,
    n3856, n3857, n3858, n3859, n3860, n3861,
    n3862, n3863, n3864, n3865, n3866, n3867,
    n3868, n3869, n3870, n3871, n3872, n3873,
    n3874, n3875, n3876, n3877, n3878, n3879,
    n3880, n3881, n3882, n3883, n3884, n3885,
    n3886, n3887, n3888, n3889, n3890, n3891,
    n3892, n3893, n3894, n3895, n3896, n3897,
    n3898, n3899, n3900, n3901, n3902, n3903,
    n3904, n3905, n3906, n3907, n3908, n3909,
    n3910, n3911, n3912, n3913, n3914, n3915,
    n3916, n3917, n3918, n3919, n3920, n3921,
    n3922, n3923, n3924, n3925, n3926, n3927,
    n3928, n3929, n3930, n3931, n3932, n3933,
    n3934, n3935, n3936, n3938, n3939, n3940,
    n3941, n3942, n3943, n3944, n3945, n3946,
    n3947, n3948, n3949, n3950, n3951, n3952,
    n3953, n3954, n3955, n3956, n3957, n3958,
    n3959, n3960, n3961, n3962, n3963, n3964,
    n3965, n3966, n3967, n3968, n3969, n3970,
    n3971, n3972, n3973, n3974, n3975, n3976,
    n3977, n3978, n3979, n3980, n3981, n3982,
    n3983, n3984, n3985, n3986, n3987, n3988,
    n3989, n3990, n3991, n3992, n3993, n3994,
    n3995, n3996, n3997, n3998, n3999, n4000,
    n4001, n4002, n4003, n4004, n4005, n4006,
    n4007, n4008, n4009, n4010, n4011, n4012,
    n4013, n4014, n4015, n4016, n4017, n4018,
    n4019, n4020, n4021, n4022, n4023, n4024,
    n4025, n4026, n4027, n4028, n4029, n4030,
    n4031, n4032, n4033, n4034, n4035, n4036,
    n4037, n4038, n4039, n4040, n4041, n4042,
    n4043, n4044, n4045, n4046, n4047, n4048,
    n4049, n4050, n4051, n4052, n4053, n4054,
    n4055, n4056, n4057, n4058, n4059, n4060,
    n4061, n4062, n4063, n4064, n4065, n4066,
    n4067, n4068, n4069, n4070, n4071, n4072,
    n4073, n4074, n4075, n4076, n4077, n4078,
    n4079, n4080, n4081, n4082, n4083, n4084,
    n4085, n4086, n4087, n4088, n4089, n4090,
    n4091, n4092, n4093, n4094, n4095, n4096,
    n4097, n4098, n4099, n4100, n4101, n4102,
    n4103, n4104, n4105, n4106, n4107, n4108,
    n4109, n4110, n4111, n4112, n4113, n4114,
    n4115, n4116, n4117, n4118, n4119, n4120,
    n4121, n4122, n4123, n4124, n4125, n4126,
    n4127, n4128, n4129, n4130, n4131, n4132,
    n4133, n4134, n4135, n4136, n4137, n4138,
    n4139, n4140, n4141, n4142, n4143, n4144,
    n4145, n4146, n4147, n4148, n4149, n4150,
    n4151, n4152, n4153, n4154, n4155, n4156,
    n4157, n4158, n4159, n4160, n4161, n4162,
    n4163, n4165, n4166, n4167, n4168, n4169,
    n4170, n4171, n4172, n4173, n4174, n4175,
    n4176, n4177, n4178, n4179, n4180, n4181,
    n4182, n4183, n4184, n4185, n4186, n4187,
    n4188, n4189, n4190, n4191, n4192, n4193,
    n4194, n4195, n4196, n4197, n4198, n4199,
    n4200, n4201, n4202, n4203, n4204, n4205,
    n4206, n4207, n4208, n4209, n4210, n4211,
    n4212, n4213, n4214, n4215, n4216, n4217,
    n4218, n4219, n4220, n4221, n4222, n4223,
    n4224, n4225, n4226, n4227, n4228, n4229,
    n4230, n4231, n4232, n4233, n4234, n4235,
    n4236, n4237, n4238, n4239, n4240, n4241,
    n4242, n4243, n4244, n4245, n4246, n4247,
    n4248, n4249, n4250, n4251, n4252, n4253,
    n4254, n4255, n4256, n4257, n4258, n4259,
    n4260, n4261, n4262, n4263, n4264, n4265,
    n4266, n4267, n4268, n4269, n4270, n4271,
    n4272, n4273, n4274, n4275, n4276, n4277,
    n4278, n4279, n4280, n4281, n4282, n4283,
    n4284, n4285, n4286, n4287, n4288, n4289,
    n4290, n4291, n4292, n4293, n4294, n4295,
    n4296, n4297, n4298, n4299, n4300, n4301,
    n4302, n4303, n4304, n4305, n4306, n4307,
    n4308, n4309, n4310, n4311, n4312, n4313,
    n4314, n4315, n4316, n4317, n4318, n4319,
    n4320, n4321, n4322, n4323, n4324, n4325,
    n4326, n4327, n4328, n4329, n4330, n4331,
    n4332, n4333, n4334, n4335, n4336, n4337,
    n4338, n4339, n4340, n4341, n4342, n4343,
    n4344, n4345, n4346, n4347, n4348, n4349,
    n4350, n4351, n4352, n4353, n4354, n4355,
    n4356, n4357, n4358, n4359, n4360, n4361,
    n4362, n4363, n4364, n4365, n4366, n4367,
    n4368, n4369, n4370, n4371, n4372, n4373,
    n4374, n4375, n4376, n4377, n4378, n4379,
    n4380, n4381, n4382, n4383, n4384, n4385,
    n4387, n4388, n4389, n4390, n4391, n4392,
    n4393, n4394, n4395, n4396, n4397, n4398,
    n4399, n4400, n4401, n4402, n4403, n4404,
    n4405, n4406, n4407, n4408, n4409, n4410,
    n4411, n4412, n4413, n4414, n4415, n4416,
    n4417, n4418, n4419, n4420, n4421, n4422,
    n4423, n4424, n4425, n4426, n4427, n4428,
    n4429, n4430, n4431, n4432, n4433, n4434,
    n4435, n4436, n4437, n4438, n4439, n4440,
    n4441, n4442, n4443, n4444, n4445, n4446,
    n4447, n4448, n4449, n4450, n4451, n4452,
    n4453, n4454, n4455, n4456, n4457, n4458,
    n4459, n4460, n4461, n4462, n4463, n4464,
    n4465, n4466, n4467, n4468, n4469, n4470,
    n4471, n4472, n4473, n4474, n4475, n4476,
    n4477, n4478, n4479, n4480, n4481, n4482,
    n4483, n4484, n4485, n4486, n4487, n4488,
    n4489, n4490, n4491, n4492, n4493, n4494,
    n4495, n4496, n4497, n4498, n4499, n4500,
    n4501, n4502, n4503, n4504, n4505, n4506,
    n4507, n4508, n4509, n4510, n4511, n4512,
    n4513, n4514, n4515, n4516, n4517, n4518,
    n4519, n4520, n4521, n4522, n4523, n4524,
    n4525, n4526, n4527, n4528, n4529, n4530,
    n4531, n4532, n4533, n4534, n4535, n4536,
    n4537, n4538, n4539, n4540, n4541, n4542,
    n4543, n4544, n4545, n4546, n4547, n4548,
    n4549, n4550, n4551, n4552, n4553, n4554,
    n4555, n4556, n4557, n4558, n4559, n4560,
    n4561, n4562, n4563, n4564, n4565, n4566,
    n4567, n4568, n4569, n4570, n4571, n4572,
    n4573, n4574, n4575, n4576, n4577, n4578,
    n4579, n4580, n4581, n4582, n4583, n4584,
    n4585, n4586, n4587, n4588, n4589, n4590,
    n4591, n4592, n4593, n4594, n4595, n4596,
    n4597, n4598, n4599, n4600, n4601, n4602,
    n4603, n4604, n4605, n4606, n4607, n4609,
    n4610, n4611, n4612, n4613, n4614, n4615,
    n4616, n4617, n4618, n4619, n4620, n4621,
    n4622, n4623, n4624, n4625, n4626, n4627,
    n4628, n4629, n4630, n4631, n4632, n4633,
    n4634, n4635, n4636, n4637, n4638, n4639,
    n4640, n4641, n4642, n4643, n4644, n4645,
    n4646, n4647, n4648, n4649, n4650, n4651,
    n4652, n4653, n4654, n4655, n4656, n4657,
    n4658, n4659, n4660, n4661, n4662, n4663,
    n4664, n4665, n4666, n4667, n4668, n4669,
    n4670, n4671, n4672, n4673, n4674, n4675,
    n4676, n4677, n4678, n4679, n4680, n4681,
    n4682, n4683, n4684, n4685, n4686, n4687,
    n4688, n4689, n4690, n4691, n4692, n4693,
    n4694, n4695, n4696, n4697, n4698, n4699,
    n4700, n4701, n4702, n4703, n4704, n4705,
    n4706, n4707, n4708, n4709, n4710, n4711,
    n4712, n4713, n4714, n4715, n4716, n4717,
    n4718, n4719, n4720, n4721, n4722, n4723,
    n4724, n4725, n4726, n4727, n4728, n4729,
    n4730, n4731, n4732, n4733, n4734, n4735,
    n4736, n4737, n4738, n4739, n4740, n4741,
    n4742, n4743, n4744, n4745, n4746, n4747,
    n4748, n4749, n4750, n4751, n4752, n4753,
    n4754, n4755, n4756, n4757, n4758, n4759,
    n4760, n4761, n4762, n4763, n4764, n4765,
    n4766, n4767, n4768, n4769, n4770, n4771,
    n4772, n4773, n4774, n4775, n4776, n4777,
    n4778, n4779, n4780, n4781, n4782, n4783,
    n4784, n4785, n4786, n4787, n4788, n4789,
    n4790, n4791, n4792, n4793, n4794, n4795,
    n4796, n4797, n4798, n4799, n4800, n4801,
    n4802, n4803, n4804, n4805, n4806, n4807,
    n4808, n4809, n4810, n4811, n4812, n4813,
    n4814, n4815, n4816, n4817, n4818, n4819,
    n4820, n4821, n4822, n4823, n4824, n4825,
    n4826, n4827, n4828, n4829, n4830, n4831,
    n4832, n4833, n4834, n4835, n4836, n4837,
    n4839, n4840, n4841, n4842, n4843, n4844,
    n4845, n4846, n4847, n4848, n4849, n4850,
    n4851, n4852, n4853, n4854, n4855, n4856,
    n4857, n4858, n4859, n4860, n4861, n4862,
    n4863, n4864, n4865, n4866, n4867, n4868,
    n4869, n4870, n4871, n4872, n4873, n4874,
    n4875, n4876, n4877, n4878, n4879, n4880,
    n4881, n4882, n4883, n4884, n4885, n4886,
    n4887, n4888, n4889, n4890, n4891, n4892,
    n4893, n4894, n4895, n4896, n4897, n4898,
    n4899, n4900, n4901, n4902, n4903, n4904,
    n4905, n4906, n4907, n4908, n4909, n4910,
    n4911, n4912, n4913, n4914, n4915, n4916,
    n4917, n4918, n4919, n4920, n4921, n4922,
    n4923, n4924, n4925, n4926, n4927, n4928,
    n4929, n4930, n4931, n4932, n4933, n4934,
    n4935, n4936, n4937, n4938, n4939, n4940,
    n4941, n4942, n4943, n4944, n4945, n4946,
    n4947, n4948, n4949, n4950, n4951, n4952,
    n4953, n4954, n4955, n4956, n4957, n4958,
    n4959, n4960, n4961, n4962, n4963, n4964,
    n4965, n4966, n4967, n4968, n4969, n4970,
    n4971, n4972, n4973, n4974, n4975, n4976,
    n4977, n4978, n4979, n4980, n4981, n4982,
    n4983, n4984, n4985, n4986, n4987, n4988,
    n4989, n4990, n4991, n4992, n4993, n4994,
    n4995, n4996, n4997, n4998, n4999, n5000,
    n5001, n5002, n5003, n5004, n5005, n5006,
    n5007, n5008, n5009, n5010, n5011, n5012,
    n5013, n5014, n5015, n5016, n5017, n5018,
    n5019, n5020, n5021, n5022, n5023, n5024,
    n5025, n5026, n5027, n5028, n5029, n5030,
    n5031, n5032, n5033, n5034, n5035, n5036,
    n5037, n5038, n5039, n5040, n5041, n5042,
    n5043, n5044, n5045, n5046, n5047, n5048,
    n5049, n5050, n5051, n5052, n5053, n5054,
    n5055, n5056, n5057, n5058, n5060, n5061,
    n5062, n5063, n5064, n5065, n5066, n5067,
    n5068, n5069, n5070, n5071, n5072, n5073,
    n5074, n5075, n5076, n5077, n5078, n5079,
    n5080, n5081, n5082, n5083, n5084, n5085,
    n5086, n5087, n5088, n5089, n5090, n5091,
    n5092, n5093, n5094, n5095, n5096, n5097,
    n5098, n5099, n5100, n5101, n5102, n5103,
    n5104, n5105, n5106, n5107, n5108, n5109,
    n5110, n5111, n5112, n5113, n5114, n5115,
    n5116, n5117, n5118, n5119, n5120, n5121,
    n5122, n5123, n5124, n5125, n5126, n5127,
    n5128, n5129, n5130, n5131, n5132, n5133,
    n5134, n5135, n5136, n5137, n5138, n5139,
    n5140, n5141, n5142, n5143, n5144, n5145,
    n5146, n5147, n5148, n5149, n5150, n5151,
    n5152, n5153, n5154, n5155, n5156, n5157,
    n5158, n5159, n5160, n5161, n5162, n5163,
    n5164, n5165, n5166, n5167, n5168, n5169,
    n5170, n5171, n5172, n5173, n5174, n5175,
    n5176, n5177, n5178, n5179, n5180, n5181,
    n5182, n5183, n5184, n5185, n5186, n5187,
    n5188, n5189, n5190, n5191, n5192, n5193,
    n5194, n5195, n5196, n5197, n5198, n5199,
    n5200, n5201, n5202, n5203, n5204, n5205,
    n5206, n5207, n5208, n5209, n5210, n5211,
    n5212, n5213, n5214, n5215, n5216, n5217,
    n5218, n5219, n5220, n5221, n5222, n5223,
    n5224, n5225, n5226, n5227, n5228, n5229,
    n5230, n5231, n5232, n5233, n5234, n5235,
    n5236, n5237, n5238, n5239, n5240, n5241,
    n5242, n5243, n5244, n5245, n5246, n5247,
    n5248, n5249, n5250, n5251, n5252, n5253,
    n5254, n5255, n5256, n5257, n5258, n5259,
    n5260, n5261, n5262, n5263, n5264, n5265,
    n5266, n5267, n5268, n5269, n5270, n5271,
    n5272, n5273, n5274, n5275, n5276, n5277,
    n5278, n5279, n5281, n5282, n5283, n5284,
    n5285, n5286, n5287, n5288, n5289, n5290,
    n5291, n5292, n5293, n5294, n5295, n5296,
    n5297, n5298, n5299, n5300, n5301, n5302,
    n5303, n5304, n5305, n5306, n5307, n5308,
    n5309, n5310, n5311, n5312, n5313, n5314,
    n5315, n5316, n5317, n5318, n5319, n5320,
    n5321, n5322, n5323, n5324, n5325, n5326,
    n5327, n5328, n5329, n5330, n5331, n5332,
    n5333, n5334, n5335, n5336, n5337, n5338,
    n5339, n5340, n5341, n5342, n5343, n5344,
    n5345, n5346, n5347, n5348, n5349, n5350,
    n5351, n5352, n5353, n5354, n5355, n5356,
    n5357, n5358, n5359, n5360, n5361, n5362,
    n5363, n5364, n5365, n5366, n5367, n5368,
    n5369, n5370, n5371, n5372, n5373, n5374,
    n5375, n5376, n5377, n5378, n5379, n5380,
    n5381, n5382, n5383, n5384, n5385, n5386,
    n5387, n5388, n5389, n5390, n5391, n5392,
    n5393, n5394, n5395, n5396, n5397, n5398,
    n5399, n5400, n5401, n5402, n5403, n5404,
    n5405, n5406, n5407, n5408, n5409, n5410,
    n5411, n5412, n5413, n5414, n5415, n5416,
    n5417, n5418, n5419, n5420, n5421, n5422,
    n5423, n5424, n5425, n5426, n5427, n5428,
    n5429, n5430, n5431, n5432, n5433, n5434,
    n5435, n5436, n5437, n5438, n5439, n5440,
    n5441, n5442, n5443, n5444, n5445, n5446,
    n5447, n5448, n5449, n5450, n5451, n5452,
    n5453, n5454, n5455, n5456, n5457, n5458,
    n5459, n5460, n5461, n5462, n5463, n5464,
    n5465, n5466, n5467, n5468, n5469, n5470,
    n5471, n5472, n5473, n5474, n5475, n5476,
    n5477, n5478, n5479, n5480, n5481, n5482,
    n5483, n5484, n5485, n5486, n5487, n5488,
    n5489, n5490, n5491, n5492, n5493, n5494,
    n5495, n5496, n5497, n5498, n5499, n5500,
    n5501, n5502, n5503, n5504, n5505, n5506,
    n5507, n5508, n5509, n5510, n5511, n5512,
    n5513, n5514, n5516, n5517, n5518, n5519,
    n5520, n5521, n5522, n5523, n5524, n5525,
    n5526, n5527, n5528, n5529, n5530, n5531,
    n5532, n5533, n5534, n5535, n5536, n5537,
    n5538, n5539, n5540, n5541, n5542, n5543,
    n5544, n5545, n5546, n5547, n5548, n5549,
    n5550, n5551, n5552, n5553, n5554, n5555,
    n5556, n5557, n5558, n5559, n5560, n5561,
    n5562, n5563, n5564, n5565, n5566, n5567,
    n5568, n5569, n5570, n5571, n5572, n5573,
    n5574, n5575, n5576, n5577, n5578, n5579,
    n5580, n5581, n5582, n5583, n5584, n5585,
    n5586, n5587, n5588, n5589, n5590, n5591,
    n5592, n5593, n5594, n5595, n5596, n5597,
    n5598, n5599, n5600, n5601, n5602, n5603,
    n5604, n5605, n5606, n5607, n5608, n5609,
    n5610, n5611, n5612, n5613, n5614, n5615,
    n5616, n5617, n5618, n5619, n5620, n5621,
    n5622, n5623, n5624, n5625, n5626, n5627,
    n5628, n5629, n5630, n5631, n5632, n5633,
    n5634, n5635, n5636, n5637, n5638, n5639,
    n5640, n5641, n5642, n5643, n5644, n5645,
    n5646, n5647, n5648, n5649, n5650, n5651,
    n5652, n5653, n5654, n5655, n5656, n5657,
    n5658, n5659, n5660, n5661, n5662, n5663,
    n5664, n5665, n5666, n5667, n5668, n5669,
    n5670, n5671, n5672, n5673, n5674, n5675,
    n5676, n5677, n5678, n5679, n5680, n5681,
    n5682, n5683, n5684, n5685, n5686, n5687,
    n5688, n5689, n5690, n5691, n5692, n5693,
    n5694, n5695, n5696, n5697, n5698, n5699,
    n5700, n5701, n5702, n5703, n5704, n5705,
    n5706, n5707, n5708, n5709, n5710, n5711,
    n5712, n5713, n5714, n5715, n5716, n5717,
    n5718, n5719, n5720, n5721, n5722, n5723,
    n5724, n5725, n5726, n5727, n5728, n5729,
    n5730, n5731, n5732, n5733, n5734, n5735,
    n5736, n5737, n5738, n5739, n5740, n5741,
    n5742, n5743, n5744, n5745, n5746, n5747,
    n5748, n5749, n5751, n5752, n5753, n5754,
    n5755, n5756, n5757, n5758, n5759, n5760,
    n5761, n5762, n5763, n5764, n5765, n5766,
    n5767, n5768, n5769, n5770, n5771, n5772,
    n5773, n5774, n5775, n5776, n5777, n5778,
    n5779, n5780, n5781, n5782, n5783, n5784,
    n5785, n5786, n5787, n5788, n5789, n5790,
    n5791, n5792, n5793, n5794, n5795, n5796,
    n5797, n5798, n5799, n5800, n5801, n5802,
    n5803, n5804, n5805, n5806, n5807, n5808,
    n5809, n5810, n5811, n5812, n5813, n5814,
    n5815, n5816, n5817, n5818, n5819, n5820,
    n5821, n5822, n5823, n5824, n5825, n5826,
    n5827, n5828, n5829, n5830, n5831, n5832,
    n5833, n5834, n5835, n5836, n5837, n5838,
    n5839, n5840, n5841, n5842, n5843, n5844,
    n5845, n5846, n5847, n5848, n5849, n5850,
    n5851, n5852, n5853, n5854, n5855, n5856,
    n5857, n5858, n5859, n5860, n5861, n5862,
    n5863, n5864, n5865, n5866, n5867, n5868,
    n5869, n5870, n5871, n5872, n5873, n5874,
    n5875, n5876, n5877, n5878, n5879, n5880,
    n5881, n5882, n5883, n5884, n5885, n5886,
    n5887, n5888, n5889, n5890, n5891, n5892,
    n5893, n5894, n5895, n5896, n5897, n5898,
    n5899, n5900, n5901, n5902, n5903, n5904,
    n5905, n5906, n5907, n5908, n5909, n5910,
    n5911, n5912, n5913, n5914, n5915, n5916,
    n5917, n5918, n5919, n5920, n5921, n5922,
    n5923, n5924, n5925, n5926, n5927, n5928,
    n5929, n5930, n5931, n5932, n5933, n5934,
    n5935, n5936, n5937, n5938, n5939, n5940,
    n5941, n5942, n5943, n5944, n5945, n5946,
    n5947, n5948, n5949, n5950, n5951, n5952,
    n5953, n5954, n5955, n5956, n5957, n5958,
    n5959, n5960, n5961, n5962, n5963, n5964,
    n5965, n5966, n5967, n5968, n5969, n5970,
    n5971, n5972, n5973, n5974, n5975, n5976,
    n5977, n5978, n5979, n5980, n5981, n5982,
    n5983, n5984, n5985, n5986, n5987, n5988,
    n5989, n5990, n5991, n5992, n5993, n5994,
    n5995, n5996, n5997, n5998, n5999, n6000,
    n6001, n6002, n6003, n6004, n6005, n6006,
    n6007, n6008, n6009, n6010, n6011, n6012,
    n6013, n6014, n6015, n6016, n6017, n6018,
    n6019, n6020, n6021, n6022, n6023, n6024,
    n6025, n6026, n6027, n6028, n6029, n6030,
    n6031, n6032, n6033, n6034, n6035, n6036,
    n6037, n6038, n6039, n6040, n6041, n6042,
    n6043, n6044, n6045, n6046, n6047, n6048,
    n6049, n6050, n6051, n6052, n6053, n6054,
    n6055, n6056, n6057, n6058, n6059, n6060,
    n6061, n6062, n6063, n6064, n6065, n6066,
    n6067, n6068, n6069, n6070, n6071, n6072,
    n6073, n6074, n6075, n6076, n6077, n6078,
    n6079, n6080, n6081, n6082, n6083, n6084,
    n6085, n6086, n6087, n6088, n6089, n6090,
    n6091, n6092, n6093, n6094, n6095, n6096,
    n6097, n6098, n6099, n6100, n6101, n6102,
    n6103, n6105, n6106, n6107, n6108, n6109,
    n6110, n6111, n6112, n6113, n6114, n6115,
    n6116, n6117, n6118, n6119, n6120, n6121,
    n6122, n6123, n6124, n6125, n6126, n6127,
    n6128, n6129, n6130, n6131, n6132, n6133,
    n6134, n6135, n6136, n6137, n6138, n6139,
    n6140, n6141, n6142, n6143, n6144, n6145,
    n6146, n6147, n6148, n6149, n6150, n6151,
    n6152, n6153, n6154, n6155, n6156, n6157,
    n6158, n6159, n6160, n6161, n6162, n6163,
    n6164, n6165, n6166, n6167, n6168, n6170,
    n6171, n6172, n6173, n6174, n6175, n6176,
    n6177, n6178, n6179, n6180, n6181, n6182,
    n6183, n6184, n6185, n6186, n6187, n6188,
    n6189, n6190, n6191, n6192, n6193, n6194,
    n6195, n6196, n6197, n6198, n6199, n6200,
    n6201, n6202, n6203, n6204, n6205, n6206,
    n6207, n6208, n6209, n6210, n6211, n6212,
    n6213, n6214, n6215, n6216, n6217, n6218,
    n6219, n6220, n6221, n6222, n6223, n6224,
    n6225, n6226, n6227, n6228, n6229, n6230,
    n6231, n6232, n6233, n6234, n6235, n6236,
    n6237, n6238, n6239, n6240, n6241, n6242,
    n6243, n6244, n6245, n6246, n6247, n6248,
    n6249, n6250, n6251, n6252, n6253, n6254,
    n6255, n6256, n6257, n6258, n6259, n6260,
    n6261, n6263, n6264, n6265, n6266, n6268,
    n6269, n6270, n6271, n6272, n6273, n6274,
    n6275, n6276, n6277, n6278, n6279, n6280,
    n6281, n6282, n6283, n6284, n6285, n6286,
    n6287, n6288, n6289, n6290, n6291, n6293,
    n6294, n6295, n6296, n6297, n6298, n6299,
    n6300, n6301, n6302, n6303, n6304, n6305,
    n6306, n6307, n6308, n6309, n6310, n6311,
    n6312, n6313, n6314, n6315, n6316, n6317,
    n6318, n6319, n6320, n6321, n6322, n6323,
    n6324, n6325, n6326, n6328, n6329, n6330,
    n6331, n6332, n6333, n6334, n6335, n6336,
    n6337, n6338, n6339, n6340, n6341, n6342,
    n6343, n6344, n6345, n6346, n6347, n6348,
    n6349, n6350, n6351, n6352, n6353, n6354,
    n6355, n6356, n6357, n6358, n6359, n6360,
    n6361, n6362, n6363, n6364, n6365, n6366,
    n6367, n6368, n6369, n6370, n6371, n6372,
    n6373, n6374, n6375, n6376, n6377, n6378,
    n6379, n6380, n6381, n6382, n6383, n6384,
    n6385, n6386, n6387, n6388, n6389, n6390,
    n6391, n6392, n6393, n6394, n6395, n6396,
    n6397, n6398, n6399, n6400, n6401, n6402,
    n6403, n6404, n6405, n6406, n6407, n6408,
    n6409, n6410, n6411, n6412, n6413, n6414,
    n6415, n6416, n6417, n6418, n6419, n6420,
    n6421, n6422, n6423, n6424, n6425, n6426,
    n6427, n6428, n6429, n6430, n6431, n6432,
    n6433, n6434, n6435, n6436, n6437, n6438,
    n6439, n6440, n6441, n6442, n6443, n6444,
    n6445, n6446, n6447, n6448, n6449, n6450,
    n6451, n6452, n6453, n6454, n6455, n6456,
    n6457, n6458, n6459, n6460, n6461, n6462,
    n6463, n6464, n6465, n6466, n6467, n6468,
    n6469, n6470, n6471, n6472, n6473, n6474,
    n6475, n6476, n6477, n6478, n6479, n6480,
    n6481, n6482, n6483, n6484, n6485, n6486,
    n6487, n6488, n6489, n6490, n6491, n6492,
    n6493, n6494, n6495, n6496, n6497, n6498,
    n6499, n6500, n6501, n6502, n6503, n6504,
    n6505, n6506, n6507, n6508, n6509, n6510,
    n6511, n6512, n6513, n6514, n6515, n6516,
    n6517, n6518, n6519, n6520, n6521, n6522,
    n6523, n6524, n6525, n6526, n6527, n6528,
    n6529, n6530, n6531, n6532, n6533, n6534,
    n6535, n6536, n6537, n6538, n6539, n6540,
    n6541, n6542, n6543, n6544, n6545, n6546,
    n6547, n6548, n6549, n6550, n6551, n6552,
    n6553, n6554, n6555, n6556, n6557, n6558,
    n6559, n6560, n6562, n6563, n6564, n6565,
    n6566, n6567, n6568, n6569, n6570, n6571,
    n6572, n6573, n6574, n6575, n6576, n6577,
    n6578, n6579, n6580, n6581, n6582, n6583,
    n6584, n6585, n6586, n6587, n6588, n6589,
    n6590, n6591, n6592, n6593, n6594, n6595,
    n6596, n6597, n6598, n6599, n6600, n6601,
    n6602, n6603, n6604, n6605, n6606, n6607,
    n6608, n6609, n6610, n6611, n6612, n6613,
    n6614, n6615, n6616, n6617, n6618, n6619,
    n6620, n6621, n6622, n6623, n6624, n6625,
    n6626, n6627, n6628, n6629, n6630, n6631,
    n6632, n6633, n6634, n6635, n6636, n6637,
    n6638, n6639, n6640, n6641, n6642, n6643,
    n6644, n6645, n6646, n6647, n6648, n6649,
    n6650, n6651, n6652, n6653, n6654, n6655,
    n6656, n6657, n6658, n6659, n6660, n6661,
    n6662, n6663, n6664, n6665, n6666, n6667,
    n6668, n6669, n6670, n6671, n6672, n6673,
    n6674, n6675, n6676, n6677, n6678, n6679,
    n6680, n6681, n6682, n6683, n6685, n6686,
    n6687, n6688, n6689, n6690, n6691, n6692,
    n6693, n6694, n6695, n6696, n6697, n6698,
    n6699, n6700, n6701, n6702, n6703, n6704,
    n6705, n6706, n6707, n6708, n6709, n6710,
    n6711, n6712, n6713, n6714, n6715, n6716,
    n6717, n6718, n6719, n6720, n6721, n6722,
    n6723, n6724, n6725, n6726, n6727, n6728,
    n6729, n6730, n6731, n6732, n6733, n6734,
    n6735, n6736, n6737, n6738, n6739, n6740,
    n6741, n6742, n6743, n6744, n6745, n6746,
    n6747, n6748, n6749, n6750, n6751, n6752,
    n6753, n6754, n6755, n6756, n6757, n6758,
    n6759, n6760, n6761, n6762, n6763, n6764,
    n6765, n6766, n6767, n6768, n6769, n6770,
    n6771, n6772, n6773, n6774, n6775, n6776,
    n6777, n6778, n6779, n6780, n6781, n6782,
    n6783, n6784, n6785, n6786, n6787, n6788,
    n6789, n6790, n6791, n6792, n6793, n6794,
    n6795, n6796, n6797, n6798, n6799, n6800,
    n6801, n6802, n6803, n6804, n6805, n6806,
    n6807, n6808, n6809, n6810, n6811, n6812,
    n6813, n6815, n6816, n6817, n6818, n6819,
    n6820, n6821, n6822, n6823, n6824, n6825,
    n6826, n6827, n6828, n6829, n6830, n6831,
    n6832, n6833, n6834, n6835, n6836, n6837,
    n6838, n6839, n6840, n6841, n6842, n6843,
    n6844, n6845, n6846, n6847, n6848, n6849,
    n6850, n6851, n6852, n6853, n6854, n6855,
    n6856, n6857, n6858, n6859, n6860, n6861,
    n6862, n6863, n6864, n6865, n6866, n6867,
    n6868, n6869, n6870, n6871, n6872, n6873,
    n6874, n6875, n6876, n6877, n6878, n6879,
    n6880, n6881, n6882, n6883, n6884, n6885,
    n6886, n6887, n6888, n6889, n6890, n6891,
    n6892, n6893, n6894, n6895, n6896, n6897,
    n6898, n6899, n6900, n6901, n6902, n6903,
    n6904, n6905, n6906, n6907, n6908, n6909,
    n6911, n6912, n6913, n6914, n6915, n6916,
    n6917, n6918, n6919, n6920, n6921, n6922,
    n6923, n6924, n6925, n6926, n6927, n6928,
    n6929, n6930, n6931, n6932, n6933, n6934,
    n6935, n6936, n6937, n6938, n6939, n6940,
    n6941, n6942, n6943, n6944, n6945, n6946,
    n6947, n6948, n6949, n6950, n6951, n6952,
    n6953, n6954, n6955, n6956, n6957, n6958,
    n6959, n6960, n6961, n6962, n6963, n6964,
    n6965, n6966, n6967, n6968, n6969, n6970,
    n6971, n6972, n6973, n6974, n6975, n6976,
    n6977, n6978, n6979, n6980, n6981, n6982,
    n6983, n6984, n6985, n6986, n6987, n6988,
    n6989, n6990, n6991, n6992, n6993, n6994,
    n6995, n6996, n6997, n6998, n6999, n7000,
    n7001, n7002, n7003, n7004, n7005, n7007,
    n7008, n7009, n7010, n7011, n7012, n7013,
    n7014, n7015, n7016, n7017, n7018, n7019,
    n7020, n7021, n7022, n7023, n7024, n7025,
    n7026, n7027, n7028, n7029, n7030, n7031,
    n7032, n7033, n7034, n7035, n7036, n7037,
    n7038, n7039, n7040, n7041, n7042, n7043,
    n7044, n7045, n7046, n7047, n7048, n7049,
    n7050, n7051, n7052, n7053, n7054, n7055,
    n7056, n7057, n7058, n7059, n7060, n7061,
    n7062, n7063, n7064, n7065, n7066, n7067,
    n7068, n7069, n7070, n7071, n7072, n7073,
    n7074, n7075, n7076, n7077, n7078, n7079,
    n7080, n7081, n7082, n7083, n7084, n7085,
    n7086, n7087, n7088, n7089, n7090, n7091,
    n7092, n7093, n7094, n7095, n7096, n7097,
    n7098, n7099, n7100, n7101, n7103, n7104,
    n7105, n7106, n7107, n7108, n7109, n7110,
    n7111, n7112, n7113, n7114, n7115, n7116,
    n7117, n7118, n7119, n7120, n7121, n7122,
    n7123, n7124, n7125, n7126, n7127, n7128,
    n7129, n7130, n7131, n7132, n7133, n7134,
    n7135, n7136, n7137, n7138, n7139, n7140,
    n7141, n7142, n7143, n7144, n7145, n7146,
    n7147, n7148, n7149, n7150, n7151, n7152,
    n7153, n7154, n7155, n7156, n7157, n7158,
    n7159, n7160, n7161, n7162, n7163, n7164,
    n7165, n7166, n7167, n7168, n7169, n7170,
    n7171, n7172, n7173, n7174, n7175, n7176,
    n7177, n7178, n7179, n7180, n7181, n7182,
    n7183, n7184, n7185, n7186, n7187, n7188,
    n7189, n7190, n7191, n7192, n7193, n7194,
    n7195, n7196, n7197, n7199, n7200, n7201,
    n7202, n7203, n7204, n7205, n7206, n7207,
    n7208, n7209, n7210, n7211, n7212, n7213,
    n7214, n7215, n7216, n7217, n7218, n7219,
    n7220, n7221, n7222, n7223, n7224, n7225,
    n7226, n7227, n7228, n7229, n7230, n7231,
    n7232, n7233, n7234, n7235, n7236, n7237,
    n7238, n7239, n7240, n7241, n7242, n7243,
    n7244, n7245, n7246, n7247, n7248, n7249,
    n7250, n7251, n7252, n7253, n7254, n7255,
    n7256, n7257, n7258, n7259, n7260, n7261,
    n7262, n7263, n7264, n7265, n7266, n7267,
    n7268, n7269, n7270, n7271, n7272, n7273,
    n7274, n7275, n7276, n7277, n7278, n7279,
    n7280, n7281, n7282, n7283, n7284, n7285,
    n7286, n7287, n7288, n7289, n7291, n7292,
    n7293, n7294, n7295, n7296, n7297, n7298,
    n7299, n7300, n7301, n7302, n7303, n7304,
    n7305, n7306, n7307, n7308, n7309, n7310,
    n7311, n7312, n7313, n7314, n7315, n7316,
    n7317, n7318, n7319, n7320, n7321, n7322,
    n7323, n7324, n7325, n7326, n7327, n7328,
    n7329, n7330, n7331, n7332, n7333, n7334,
    n7335, n7336, n7337, n7338, n7339, n7340,
    n7341, n7343, n7344, n7346, n7347, n7348,
    n7349, n7350, n7351, n7352, n7353, n7354,
    n7355, n7356, n7357, n7358, n7359, n7360,
    n7361, n7362, n7363, n7364, n7365, n7366,
    n7367, n7368, n7369, n7370, n7371, n7372,
    n7373, n7374, n7375, n7376, n7377, n7378,
    n7379, n7380, n7381, n7382, n7383, n7384,
    n7385, n7386, n7387, n7388, n7389, n7390,
    n7391, n7392, n7393, n7394, n7396, n7397,
    n7398, n7399, n7401, n7403, n7405, n7407,
    n7408, n7409, n7410, n7411, n7412, n7413,
    n7414, n7415, n7416, n7417, n7418, n7419,
    n7420, n7421, n7422, n7423, n7424, n7425,
    n7426, n7427, n7428, n7429, n7430, n7431,
    n7432, n7433, n7434, n7435, n7436, n7437,
    n7438, n7439, n7440, n7441, n7442, n7443,
    n7444, n7445, n7446, n7447, n7448, n7449,
    n7450, n7451, n7452, n7453, n7454, n7455,
    n7456, n7457, n7458, n7459, n7460, n7461,
    n7462, n7463, n7464, n7465, n7466, n7467,
    n7468, n7469, n7470, n7471, n7472, n7473,
    n7474, n7475, n7476, n7477, n7478, n7479,
    n7480, n7481, n7482, n7483, n7484, n7485,
    n7486, n7487, n7488, n7489, n7490, n7491,
    n7492, n7493, n7494, n7495, n7496, n7497,
    n7498, n7499, n7500, n7501, n7502, n7503,
    n7504, n7505, n7506, n7507, n7508, n7509,
    n7510, n7511, n7512, n7513, n7514, n7515,
    n7516, n7517, n7518, n7519, n7520, n7521,
    n7522, n7523, n7524, n7525, n7526, n7527,
    n7528, n7529, n7530, n7531, n7532, n7533,
    n7534, n7535, n7536, n7537, n7538, n7539,
    n7540, n7541, n7542, n7543, n7544, n7545,
    n7546, n7547, n7548, n7549, n7550, n7551,
    n7552, n7553, n7554, n7555, n7556, n7557,
    n7558, n7559, n7560, n7561, n7562, n7563,
    n7564, n7565, n7566, n7567, n7568, n7569,
    n7570, n7571, n7572, n7573, n7574, n7575,
    n7576, n7577, n7578, n7579, n7580, n7581,
    n7582, n7583, n7584, n7585, n7586, n7587,
    n7588, n7589, n7590, n7591, n7592, n7593,
    n7594, n7595, n7596, n7597, n7598, n7599,
    n7600, n7601, n7602, n7603, n7604, n7605,
    n7606, n7607, n7608, n7609, n7610, n7611,
    n7612, n7613, n7614, n7615, n7616, n7617,
    n7618, n7619, n7620, n7621, n7622, n7623,
    n7624, n7625, n7626, n7627, n7628, n7629,
    n7630, n7631, n7632, n7633, n7634, n7635,
    n7636, n7637, n7638, n7639, n7640, n7641,
    n7642, n7643, n7644, n7645, n7646, n7647,
    n7648, n7649, n7650, n7651, n7652, n7653,
    n7654, n7655, n7656, n7657, n7658, n7659,
    n7660, n7661, n7662, n7663, n7664, n7665,
    n7666, n7667, n7668, n7669, n7670, n7671,
    n7672, n7673, n7674, n7675, n7676, n7677,
    n7678, n7679, n7680, n7681, n7682, n7683,
    n7684, n7685, n7686, n7687, n7688, n7689,
    n7690, n7691, n7692, n7693, n7694, n7695,
    n7696, n7697, n7698, n7699, n7700, n7701,
    n7702, n7703, n7704, n7705, n7706, n7707,
    n7708, n7709, n7710, n7711, n7712, n7713,
    n7714, n7715, n7716, n7717, n7718, n7719,
    n7720, n7721, n7722, n7723, n7724, n7725,
    n7726, n7727, n7728, n7729, n7730, n7731,
    n7732, n7733, n7734, n7735, n7736, n7737,
    n7738, n7739, n7740, n7741, n7742, n7743,
    n7744, n7745, n7746, n7747, n7748, n7749,
    n7750, n7751, n7752, n7753, n7754, n7755,
    n7756, n7757, n7758, n7759, n7760, n7761,
    n7762, n7763, n7764, n7765, n7766, n7767,
    n7768, n7769, n7770, n7771, n7772, n7773,
    n7774, n7775, n7776, n7777, n7778, n7779,
    n7780, n7781, n7782, n7783, n7784, n7785,
    n7786, n7787, n7788, n7789, n7790, n7791,
    n7792, n7793, n7794, n7795, n7796, n7797,
    n7798, n7799, n7800, n7801, n7802, n7803,
    n7804, n7805, n7806, n7807, n7808, n7809,
    n7810, n7811, n7812, n7813, n7814, n7815,
    n7816, n7817, n7818, n7819, n7820, n7821,
    n7822, n7823, n7824, n7825, n7826, n7827,
    n7828, n7829, n7830, n7831, n7832, n7833,
    n7834, n7835, n7836, n7837, n7838, n7839,
    n7840, n7841, n7842, n7843, n7844, n7845,
    n7846, n7847, n7848, n7849, n7850, n7851,
    n7852, n7853, n7854, n7855, n7856, n7857,
    n7858, n7859, n7860, n7861, n7862, n7863,
    n7864, n7865, n7866, n7867, n7868, n7869,
    n7870, n7871, n7872, n7873, n7874, n7875,
    n7876, n7877, n7878, n7879, n7880, n7881,
    n7882, n7883, n7884, n7885, n7886, n7887,
    n7888, n7889, n7890, n7891, n7892, n7893,
    n7894, n7895, n7896, n7897, n7898, n7899,
    n7900, n7901, n7902, n7903, n7904, n7905,
    n7906, n7907, n7908, n7909, n7910, n7911,
    n7912, n7913, n7914, n7915, n7916, n7917,
    n7918, n7919, n7920, n7921, n7922, n7923,
    n7924, n7925, n7926, n7927, n7928, n7929,
    n7930, n7931, n7932, n7933, n7934, n7935,
    n7936, n7937, n7938, n7939, n7940, n7941,
    n7942, n7943, n7944, n7945, n7946, n7947,
    n7948, n7949, n7950, n7951, n7952, n7953,
    n7954, n7955, n7956, n7957, n7958, n7959,
    n7960, n7961, n7962, n7963, n7964, n7965,
    n7966, n7967, n7968, n7969, n7970, n7971,
    n7972, n7973, n7974, n7975, n7976, n7977,
    n7978, n7979, n7980, n7981, n7982, n7983,
    n7984, n7985, n7986, n7987, n7988, n7989,
    n7990, n7991, n7992, n7993, n7994, n7995,
    n7996, n7997, n7998, n7999, n8000, n8001,
    n8002, n8003, n8004, n8005, n8006, n8007,
    n8008, n8009, n8010, n8011, n8012, n8013,
    n8014, n8015, n8016, n8017, n8018, n8019,
    n8020, n8021, n8022, n8023, n8024, n8025,
    n8026, n8027, n8028, n8029, n8030, n8031,
    n8032, n8033, n8034, n8035, n8036, n8037,
    n8038, n8039, n8040, n8041, n8042, n8043,
    n8044, n8045, n8046, n8047, n8048, n8049,
    n8050, n8051, n8052, n8053, n8054, n8055,
    n8056, n8057, n8058, n8059, n8060, n8061,
    n8062, n8063, n8064, n8065, n8066, n8067,
    n8068, n8069, n8070, n8071, n8072, n8073,
    n8074, n8075, n8076, n8077, n8078, n8079,
    n8080, n8081, n8082, n8083, n8084, n8085,
    n8086, n8087, n8088, n8089, n8090, n8091,
    n8092, n8093, n8094, n8095, n8096, n8097,
    n8098, n8099, n8100, n8101, n8102, n8103,
    n8104, n8105, n8106, n8107, n8108, n8109,
    n8110, n8111, n8112, n8113, n8114, n8115,
    n8116, n8117, n8118, n8119, n8120, n8121,
    n8122, n8123, n8124, n8125, n8126, n8127,
    n8128, n8129, n8130, n8131, n8132, n8133,
    n8134, n8135, n8136, n8137, n8138, n8139,
    n8140, n8141, n8142, n8143, n8144, n8145,
    n8146, n8147, n8148, n8149, n8150, n8151,
    n8152, n8153, n8154, n8155, n8156, n8157,
    n8158, n8159, n8160, n8161, n8162, n8163,
    n8164, n8165, n8166, n8167, n8168, n8169,
    n8170, n8171, n8172, n8173, n8174, n8175,
    n8176, n8177, n8178, n8179, n8180, n8181,
    n8182, n8183, n8184, n8185, n8186, n8187,
    n8188, n8189, n8190, n8191, n8192, n8193,
    n8194, n8195, n8196, n8197, n8198, n8199,
    n8200, n8201, n8202, n8203, n8204, n8205,
    n8206, n8207, n8208, n8209, n8210, n8211,
    n8212, n8213, n8214, n8215, n8216, n8217,
    n8218, n8219, n8220, n8221, n8222, n8223,
    n8224, n8225, n8226, n8227, n8228, n8229,
    n8230, n8231, n8232, n8233, n8234, n8235,
    n8236, n8237, n8238, n8239, n8240, n8241,
    n8242, n8243, n8244, n8245, n8246, n8247,
    n8248, n8249, n8250, n8251, n8252, n8253,
    n8254, n8255, n8256, n8257, n8258, n8259,
    n8260, n8261, n8262, n8263, n8264, n8265,
    n8266, n8267, n8268, n8269, n8270, n8271,
    n8272, n8273, n8274, n8275, n8276, n8277,
    n8278, n8279, n8280, n8281, n8282, n8283,
    n8284, n8285, n8286, n8287, n8288, n8289,
    n8290, n8291, n8292, n8293, n8294, n8295,
    n8296, n8297, n8298, n8299, n8300, n8301,
    n8302, n8303, n8304, n8305, n8306, n8307,
    n8308, n8309, n8310, n8311, n8312, n8313,
    n8314, n8315, n8316, n8317, n8318, n8319,
    n8320, n8321, n8322, n8323, n8324, n8325,
    n8326, n8327, n8328, n8329, n8330, n8331,
    n8332, n8333, n8334, n8335, n8336, n8337,
    n8338, n8339, n8340, n8341, n8342, n8343,
    n8344, n8345, n8346, n8347, n8348, n8349,
    n8350, n8351, n8352, n8353, n8354, n8355,
    n8356, n8357, n8358, n8359, n8360, n8361,
    n8362, n8363, n8364, n8365, n8366, n8367,
    n8368, n8369, n8370, n8371, n8372, n8373,
    n8374, n8375, n8376, n8377, n8378, n8379,
    n8380, n8381, n8382, n8383, n8384, n8385,
    n8386, n8387, n8388, n8389, n8390, n8391,
    n8392, n8393, n8394, n8395, n8396, n8397,
    n8398, n8399, n8400, n8401, n8402, n8403,
    n8404, n8405, n8406, n8407, n8408, n8409,
    n8410, n8411, n8412, n8413, n8414, n8415,
    n8416, n8417, n8418, n8419, n8420, n8421,
    n8422, n8423, n8424, n8425, n8426, n8427,
    n8428, n8429, n8430, n8431, n8432, n8433,
    n8434, n8435, n8436, n8437, n8438, n8439,
    n8440, n8441, n8442, n8443, n8444, n8445,
    n8446, n8448, n8449, n8450, n8451, n8452,
    n8453, n8454, n8455, n8456, n8457, n8458,
    n8459, n8460, n8461, n8462, n8463, n8464,
    n8465, n8466, n8467, n8468, n8469, n8470,
    n8471, n8472, n8473, n8474, n8475, n8476,
    n8477, n8478, n8479, n8480, n8481, n8482,
    n8483, n8484, n8485, n8486, n8487, n8488,
    n8489, n8490, n8491, n8492, n8493, n8494,
    n8495, n8496, n8497, n8498, n8499, n8500,
    n8501, n8502, n8503, n8504, n8505, n8506,
    n8507, n8508, n8509, n8510, n8511, n8512,
    n8513, n8514, n8515, n8516, n8517, n8518,
    n8519, n8520, n8521, n8522, n8523, n8524,
    n8525, n8526, n8527, n8528, n8529, n8530,
    n8531, n8532, n8533, n8534, n8535, n8536,
    n8537, n8538, n8539, n8540, n8541, n8542,
    n8543, n8544, n8545, n8546, n8547, n8548,
    n8549, n8550, n8551, n8552, n8553, n8554,
    n8555, n8556, n8557, n8558, n8559, n8560,
    n8561, n8562, n8563, n8564, n8565, n8566,
    n8567, n8568, n8569, n8570, n8571, n8572,
    n8573, n8574, n8575, n8576, n8577, n8578,
    n8579, n8580, n8581, n8582, n8583, n8584,
    n8585, n8586, n8587, n8588, n8589, n8590,
    n8591, n8592, n8593, n8594, n8595, n8596,
    n8597, n8598, n8599, n8600, n8601, n8602,
    n8603, n8604, n8605, n8606, n8607, n8608,
    n8609, n8610, n8611, n8612, n8613, n8614,
    n8615, n8616, n8617, n8618, n8619, n8620,
    n8621, n8622, n8623, n8624, n8625, n8626,
    n8627, n8628, n8629, n8630, n8631, n8632,
    n8633, n8634, n8635, n8636, n8637, n8638,
    n8639, n8640, n8641, n8642, n8643, n8644,
    n8645, n8646, n8647, n8648, n8649, n8650,
    n8651, n8652, n8653, n8654, n8655, n8656,
    n8657, n8658, n8659, n8660, n8661, n8662,
    n8663, n8664, n8665, n8666, n8667, n8668,
    n8669, n8670, n8671, n8672, n8673, n8674,
    n8675, n8676, n8677, n8678, n8679, n8680,
    n8681, n8682, n8683, n8684, n8685, n8686,
    n8687, n8688, n8689, n8690, n8691, n8692,
    n8693, n8694, n8695, n8696, n8697, n8698,
    n8699, n8700, n8701, n8702, n8703, n8704,
    n8705, n8706, n8707, n8708, n8709, n8710,
    n8711, n8712, n8713, n8714, n8715, n8716,
    n8717, n8718, n8719, n8720, n8721, n8722,
    n8723, n8724, n8725, n8726, n8727, n8728,
    n8729, n8730, n8731, n8732, n8733, n8734,
    n8735, n8736, n8737, n8738, n8739, n8740,
    n8741, n8742, n8743, n8744, n8745, n8746,
    n8747, n8748, n8749, n8750, n8751, n8752,
    n8753, n8754, n8755, n8756, n8757, n8758,
    n8759, n8760, n8761, n8762, n8763, n8764,
    n8765, n8766, n8767, n8768, n8769, n8770,
    n8771, n8772, n8773, n8774, n8775, n8776,
    n8777, n8778, n8779, n8780, n8781, n8782,
    n8783, n8784, n8785, n8786, n8787, n8788,
    n8789, n8790, n8791, n8792, n8793, n8794,
    n8795, n8796, n8797, n8798, n8799, n8800,
    n8801, n8802, n8803, n8804, n8805, n8806,
    n8807, n8808, n8809, n8810, n8811, n8812,
    n8813, n8814, n8815, n8816, n8817, n8818,
    n8819, n8820, n8821, n8822, n8823, n8824,
    n8825, n8826, n8827, n8828, n8829, n8830,
    n8831, n8832, n8833, n8834, n8835, n8836,
    n8837, n8838, n8839, n8840, n8841, n8842,
    n8843, n8844, n8845, n8846, n8847, n8848,
    n8849, n8850, n8851, n8852, n8853, n8854,
    n8855, n8856, n8857, n8858, n8859, n8860,
    n8861, n8862, n8864, n8865, n8866, n8867,
    n8868, n8869, n8870, n8871, n8872, n8873,
    n8874, n8875, n8876, n8877, n8878, n8879,
    n8880, n8881, n8882, n8883, n8884, n8885,
    n8886, n8887, n8888, n8889, n8890, n8892,
    n8893, n8894, n8895, n8896, n8897, n8898,
    n8899, n8900, n8901, n8902, n8903, n8904,
    n8905, n8906, n8907, n8908, n8909, n8910,
    n8911, n8912, n8913, n8914, n8915, n8916,
    n8917, n8918, n8919, n8920, n8921, n8922,
    n8923, n8924, n8925, n8926, n8927, n8928,
    n8929, n8930, n8931, n8932, n8933, n8934,
    n8935, n8936, n8937, n8938, n8939, n8940,
    n8941, n8942, n8943, n8944, n8945, n8946,
    n8947, n8948, n8949, n8950, n8951, n8952,
    n8953, n8954, n8955, n8956, n8957, n8958,
    n8960, n8961, n8962, n8963, n8964, n8965,
    n8966, n8967, n8968, n8969, n8970, n8971,
    n8972, n8973, n8974, n8975, n8976, n8977,
    n8978, n8979, n8980, n8981, n8982, n8983,
    n8984, n8985, n8986, n8987, n8988, n8989,
    n8990, n8991, n8992, n8993, n8994, n8995,
    n8996, n8997, n8998, n8999, n9000, n9001,
    n9002, n9003, n9004, n9005, n9006, n9007,
    n9008, n9009, n9010, n9011, n9012, n9013,
    n9014, n9015, n9016, n9017, n9018, n9019,
    n9020, n9021, n9022, n9023, n9024, n9025,
    n9026, n9027, n9028, n9029, n9030, n9031,
    n9032, n9033, n9034, n9035, n9036, n9037,
    n9038, n9039, n9040, n9041, n9042, n9043,
    n9044, n9045, n9046, n9047, n9048, n9049,
    n9050, n9051, n9052, n9053, n9054, n9055,
    n9056, n9057, n9058, n9059, n9060, n9061,
    n9062, n9063, n9064, n9065, n9066, n9067,
    n9068, n9069, n9070, n9071, n9072, n9073,
    n9074, n9075, n9076, n9077, n9078, n9079,
    n9080, n9081, n9082, n9083, n9084, n9085,
    n9086, n9087, n9088, n9089, n9090, n9091,
    n9092, n9093, n9094, n9095, n9096, n9097,
    n9098, n9099, n9100, n9101, n9102, n9103,
    n9104, n9105, n9106, n9107, n9108, n9109,
    n9110, n9111, n9112, n9113, n9114, n9115,
    n9116, n9117, n9118, n9119, n9120, n9121,
    n9122, n9123, n9124, n9125, n9126, n9127,
    n9128, n9129, n9130, n9131, n9132, n9133,
    n9134, n9135, n9136, n9137, n9138, n9139,
    n9140, n9141, n9142, n9143, n9144, n9145,
    n9146, n9147, n9148, n9149, n9150, n9151,
    n9152, n9153, n9154, n9155, n9156, n9157,
    n9158, n9159, n9160, n9161, n9162, n9163,
    n9164, n9165, n9166, n9167, n9168, n9169,
    n9170, n9171, n9172, n9173, n9174, n9175,
    n9176, n9177, n9178, n9179, n9180, n9181,
    n9182, n9183, n9184, n9185, n9186, n9187,
    n9188, n9189, n9190, n9191, n9192, n9193,
    n9194, n9195, n9196, n9197, n9198, n9199,
    n9200, n9201, n9202, n9203, n9204, n9205,
    n9206, n9207, n9208, n9209, n9210, n9211,
    n9212, n9213, n9214, n9215, n9216, n9217,
    n9218, n9219, n9220, n9221, n9222, n9223,
    n9224, n9225, n9226, n9227, n9228, n9229,
    n9230, n9231, n9232, n9233, n9234, n9235,
    n9236, n9237, n9238, n9239, n9240, n9241,
    n9242, n9243, n9244, n9245, n9246, n9247,
    n9248, n9249, n9250, n9251, n9252, n9253,
    n9254, n9255, n9256, n9257, n9258, n9259,
    n9260, n9261, n9262, n9263, n9264, n9265,
    n9266, n9267, n9268, n9269, n9270, n9271,
    n9272, n9273, n9274, n9275, n9276, n9277,
    n9278, n9279, n9280, n9281, n9282, n9283,
    n9284, n9285, n9286, n9287, n9288, n9289,
    n9290, n9291, n9292, n9293, n9294, n9295,
    n9296, n9297, n9298, n9299, n9300, n9301,
    n9302, n9303, n9304, n9305, n9306, n9307,
    n9308, n9309, n9310, n9311, n9312, n9313,
    n9314, n9315, n9316, n9317, n9318, n9319,
    n9320, n9321, n9322, n9323, n9324, n9325,
    n9326, n9327, n9328, n9329, n9330, n9331,
    n9332, n9333, n9334, n9335, n9336, n9337,
    n9338, n9339, n9340, n9341, n9342, n9343,
    n9344, n9345, n9346, n9347, n9348, n9349,
    n9350, n9351, n9352, n9353, n9354, n9355,
    n9356, n9357, n9358, n9359, n9360, n9361,
    n9362, n9363, n9364, n9365, n9366, n9367,
    n9368, n9369, n9370, n9371, n9372, n9373,
    n9374, n9375, n9376, n9377, n9378, n9379,
    n9380, n9381, n9382, n9383, n9384, n9385,
    n9386, n9387, n9388, n9389, n9390, n9391,
    n9392, n9393, n9394, n9395, n9396, n9397,
    n9398, n9399, n9400, n9401, n9402, n9403,
    n9404, n9405, n9406, n9407, n9408, n9409,
    n9410, n9411, n9412, n9413, n9414, n9415,
    n9416, n9417, n9418, n9419, n9420, n9421,
    n9422, n9423, n9424, n9425, n9426, n9427,
    n9428, n9429, n9430, n9431, n9432, n9433,
    n9434, n9435, n9436, n9437, n9438, n9439,
    n9440, n9441, n9442, n9443, n9444, n9445,
    n9446, n9447, n9448, n9449, n9450, n9451,
    n9452, n9453, n9454, n9455, n9456, n9457,
    n9458, n9459, n9460, n9461, n9462, n9463,
    n9464, n9465, n9466, n9467, n9468, n9469,
    n9470, n9471, n9472, n9473, n9474, n9475,
    n9476, n9477, n9478, n9479, n9480, n9481,
    n9482, n9483, n9484, n9485, n9486, n9487,
    n9488, n9489, n9490, n9491, n9492, n9493,
    n9494, n9495, n9496, n9497, n9498, n9499,
    n9500, n9501, n9502, n9503, n9504, n9505,
    n9506, n9507, n9508, n9509, n9510, n9511,
    n9512, n9513, n9514, n9515, n9516, n9517,
    n9518, n9519, n9520, n9521, n9522, n9523,
    n9524, n9525, n9526, n9527, n9528, n9529,
    n9530, n9531, n9532, n9533, n9534, n9535,
    n9536, n9537, n9538, n9539, n9540, n9541,
    n9542, n9543, n9544, n9545, n9546, n9547,
    n9548, n9549, n9550, n9551, n9552, n9553,
    n9554, n9555, n9556, n9557, n9558, n9559,
    n9560, n9561, n9562, n9563, n9564, n9565,
    n9566, n9567, n9568, n9569, n9570, n9571,
    n9572, n9573, n9574, n9575, n9576, n9577,
    n9578, n9579, n9580, n9581, n9582, n9583,
    n9584, n9585, n9586, n9587, n9588, n9589,
    n9590, n9591, n9592, n9593, n9594, n9595,
    n9596, n9597, n9598, n9599, n9600, n9601,
    n9602, n9603, n9604, n9605, n9606, n9607,
    n9608, n9609, n9610, n9611, n9612, n9613,
    n9614, n9615, n9616, n9617, n9618, n9619,
    n9620, n9621, n9622, n9623, n9624, n9625,
    n9626, n9627, n9628, n9629, n9630, n9631,
    n9632, n9633, n9634, n9635, n9636, n9637,
    n9638, n9639, n9640, n9641, n9642, n9643,
    n9644, n9645, n9646, n9647, n9648, n9649,
    n9650, n9651, n9652, n9653, n9654, n9655,
    n9656, n9657, n9658, n9659, n9660, n9661,
    n9662, n9663, n9664, n9665, n9666, n9667,
    n9668, n9669, n9670, n9671, n9672, n9673,
    n9674, n9676, n9677, n9678, n9679, n9680,
    n9681, n9682, n9683, n9684, n9685, n9686,
    n9687, n9688, n9689, n9690, n9691, n9692,
    n9693, n9694, n9695, n9696, n9697, n9698,
    n9699, n9700, n9701, n9702, n9703, n9704,
    n9705, n9706, n9707, n9708, n9709, n9710,
    n9711, n9712, n9713, n9714, n9715, n9716,
    n9717, n9718, n9719, n9720, n9721, n9722,
    n9723, n9724, n9725, n9726, n9727, n9728,
    n9729, n9730, n9731, n9732, n9733, n9734,
    n9735, n9736, n9737, n9738, n9739, n9740,
    n9741, n9742, n9743, n9744, n9745, n9746,
    n9747, n9748, n9749, n9750, n9751, n9752,
    n9753, n9754, n9755, n9756, n9757, n9758,
    n9759, n9760, n9761, n9762, n9763, n9764,
    n9765, n9766, n9767, n9768, n9769, n9770,
    n9771, n9772, n9773, n9774, n9775, n9776,
    n9777, n9778, n9779, n9780, n9781, n9782,
    n9783, n9784, n9785, n9786, n9787, n9788,
    n9789, n9790, n9791, n9792, n9793, n9794,
    n9795, n9796, n9797, n9798, n9799, n9800,
    n9801, n9802, n9803, n9804, n9805, n9806,
    n9807, n9808, n9809, n9810, n9811, n9812,
    n9813, n9814, n9815, n9816, n9817, n9818,
    n9819, n9820, n9821, n9822, n9823, n9824,
    n9825, n9826, n9827, n9828, n9829, n9830,
    n9831, n9832, n9833, n9834, n9835, n9836,
    n9837, n9838, n9839, n9840, n9841, n9842,
    n9843, n9844, n9845, n9846, n9847, n9848,
    n9849, n9850, n9851, n9852, n9853, n9854,
    n9855, n9856, n9857, n9858, n9859, n9860,
    n9861, n9862, n9863, n9864, n9865, n9866,
    n9867, n9868, n9869, n9870, n9871, n9872,
    n9873, n9874, n9875, n9876, n9877, n9878,
    n9879, n9880, n9881, n9882, n9883, n9884,
    n9885, n9886, n9887, n9888, n9889, n9890,
    n9891, n9892, n9893, n9894, n9895, n9896,
    n9897, n9898, n9899, n9900, n9901, n9902,
    n9903, n9904, n9905, n9906, n9907, n9908,
    n9909, n9910, n9911, n9912, n9913, n9914,
    n9915, n9916, n9917, n9918, n9919, n9920,
    n9921, n9922, n9923, n9924, n9925, n9926,
    n9927, n9928, n9929, n9930, n9931, n9932,
    n9933, n9934, n9935, n9936, n9937, n9938,
    n9939, n9940, n9941, n9942, n9943, n9944,
    n9945, n9946, n9947, n9948, n9949, n9950,
    n9951, n9952, n9953, n9954, n9955, n9956,
    n9957, n9958, n9959, n9960, n9961, n9962,
    n9963, n9964, n9965, n9966, n9967, n9968,
    n9969, n9970, n9971, n9972, n9973, n9974,
    n9975, n9976, n9977, n9978, n9979, n9980,
    n9981, n9982, n9983, n9984, n9985, n9986,
    n9987, n9988, n9989, n9990, n9991, n9992,
    n9993, n9994, n9995, n9996, n9997, n9998,
    n9999, n10000, n10001, n10002, n10003, n10004,
    n10005, n10006, n10007, n10008, n10009, n10010,
    n10011, n10012, n10013, n10014, n10015, n10016,
    n10017, n10018, n10019, n10020, n10021, n10022,
    n10023, n10024, n10025, n10026, n10027, n10028,
    n10029, n10030, n10031, n10032, n10033, n10034,
    n10035, n10036, n10037, n10038, n10039, n10040,
    n10041, n10042, n10043, n10044, n10045, n10046,
    n10047, n10048, n10049, n10050, n10052, n10053,
    n10054, n10055, n10056, n10057, n10058, n10059,
    n10060, n10061, n10062, n10063, n10064, n10065,
    n10066, n10067, n10068, n10069, n10070, n10071,
    n10072, n10073, n10074, n10075, n10076, n10077,
    n10078, n10079, n10080, n10081, n10082, n10083,
    n10084, n10085, n10086, n10087, n10088, n10089,
    n10090, n10091, n10092, n10093, n10094, n10095,
    n10096, n10097, n10098, n10099, n10100, n10101,
    n10102, n10103, n10104, n10105, n10106, n10107,
    n10108, n10109, n10110, n10111, n10112, n10113,
    n10114, n10115, n10116, n10117, n10118, n10119,
    n10120, n10121, n10122, n10123, n10124, n10125,
    n10126, n10128, n10129, n10130, n10131, n10132,
    n10133, n10134, n10135, n10136, n10137, n10138,
    n10139, n10140, n10141, n10142, n10143, n10144,
    n10145, n10146, n10147, n10148, n10150, n10151,
    n10152, n10153, n10154, n10155, n10156, n10157,
    n10158, n10159, n10160, n10161, n10162, n10163,
    n10164, n10165, n10166, n10167, n10168, n10169,
    n10170, n10171, n10172, n10173, n10174, n10175,
    n10176, n10177, n10178, n10179, n10181, n10182,
    n10183, n10184, n10185, n10186, n10187, n10188,
    n10189, n10190, n10191, n10192, n10193, n10194,
    n10195, n10196, n10197, n10198, n10199, n10200,
    n10201, n10202, n10203, n10204, n10205, n10206,
    n10207, n10208, n10209, n10210, n10211, n10212,
    n10213, n10214, n10215, n10216, n10217, n10218,
    n10219, n10220, n10221, n10222, n10223, n10224,
    n10225, n10226, n10227, n10228, n10229, n10230,
    n10231, n10232, n10233, n10234, n10235, n10236,
    n10237, n10238, n10239, n10240, n10241, n10242,
    n10243, n10244, n10245, n10246, n10247, n10248,
    n10249, n10250, n10251, n10252, n10253, n10254,
    n10255, n10256, n10257, n10258, n10259, n10260,
    n10262, n10263, n10264, n10265, n10266, n10267,
    n10268, n10269, n10270, n10271, n10272, n10273,
    n10275, n10276, n10277, n10278, n10279, n10280,
    n10281, n10282, n10283, n10284, n10285, n10286,
    n10287, n10288, n10289, n10290, n10291, n10292,
    n10293, n10294, n10295, n10296, n10297, n10298,
    n10299, n10300, n10301, n10302, n10303, n10304,
    n10305, n10306, n10307, n10308, n10309, n10310,
    n10311, n10312, n10313, n10314, n10315, n10316,
    n10317, n10318, n10319, n10320, n10321, n10322,
    n10323, n10324, n10325, n10326, n10327, n10328,
    n10329, n10330, n10331, n10332, n10333, n10334,
    n10335, n10336, n10337, n10338, n10339, n10340,
    n10341, n10342, n10343, n10344, n10345, n10346,
    n10347, n10348, n10349, n10350, n10351, n10352,
    n10353, n10354, n10355, n10356, n10357, n10358,
    n10359, n10360, n10361, n10362, n10363, n10364,
    n10365, n10366, n10367, n10368, n10369, n10370,
    n10371, n10372, n10373, n10374, n10375, n10376,
    n10377, n10378, n10379, n10380, n10381, n10382,
    n10383, n10384, n10385, n10386, n10387, n10388,
    n10389, n10390, n10391, n10392, n10393, n10394,
    n10395, n10396, n10397, n10398, n10399, n10400,
    n10401, n10402, n10403, n10404, n10405, n10406,
    n10407, n10408, n10409, n10410, n10411, n10412,
    n10413, n10414, n10415, n10416, n10417, n10418,
    n10419, n10420, n10421, n10422, n10423, n10424,
    n10425, n10426, n10427, n10428, n10429, n10430,
    n10431, n10432, n10433, n10434, n10435, n10436,
    n10437, n10438, n10439, n10440, n10441, n10442,
    n10443, n10444, n10445, n10446, n10447, n10448,
    n10449, n10450, n10451, n10452, n10453, n10454,
    n10455, n10456, n10457, n10458, n10459, n10460,
    n10461, n10463, n10464, n10465, n10466, n10467,
    n10468, n10469, n10470, n10471, n10472, n10473,
    n10474, n10475, n10476, n10477, n10478, n10479,
    n10480, n10481, n10482, n10483, n10484, n10485,
    n10486, n10487, n10488, n10489, n10490, n10491,
    n10492, n10493, n10494, n10495, n10496, n10497,
    n10498, n10499, n10500, n10501, n10502, n10503,
    n10504, n10505, n10506, n10507, n10508, n10509,
    n10510, n10511, n10512, n10513, n10514, n10515,
    n10516, n10517, n10518, n10519, n10520, n10521,
    n10522, n10523, n10524, n10525, n10526, n10527,
    n10528, n10529, n10530, n10531, n10532, n10533,
    n10534, n10535, n10536, n10537, n10538, n10539,
    n10540, n10541, n10542, n10543, n10544, n10545,
    n10546, n10547, n10548, n10549, n10550, n10551,
    n10552, n10553, n10554, n10555, n10556, n10557,
    n10558, n10559, n10560, n10561, n10562, n10563,
    n10564, n10565, n10566, n10567, n10568, n10569,
    n10570, n10571, n10572, n10573, n10574, n10575,
    n10576, n10577, n10578, n10579, n10580, n10581,
    n10582, n10583, n10584, n10585, n10586, n10587,
    n10588, n10589, n10590, n10591, n10592, n10593,
    n10594, n10595, n10596, n10597, n10598, n10599,
    n10600, n10601, n10602, n10603, n10604, n10605,
    n10606, n10607, n10608, n10609, n10610, n10611,
    n10612, n10613, n10614, n10615, n10616, n10617,
    n10618, n10619, n10620, n10621, n10622, n10623,
    n10624, n10625, n10626, n10627, n10628, n10629,
    n10630, n10631, n10632, n10633, n10634, n10635,
    n10636, n10637, n10638, n10639, n10640, n10641,
    n10642, n10643, n10644, n10645, n10646, n10647,
    n10648, n10649, n10650, n10651, n10652, n10653,
    n10654, n10655, n10656, n10657, n10658, n10659,
    n10660, n10661, n10662, n10663, n10664, n10665,
    n10666, n10667, n10668, n10669, n10670, n10671,
    n10672, n10673, n10674, n10675, n10676, n10677,
    n10678, n10679, n10680, n10681, n10682, n10683,
    n10684, n10685, n10686, n10687, n10688, n10689,
    n10690, n10691, n10692, n10693, n10694, n10695,
    n10696, n10697, n10698, n10699, n10700, n10701,
    n10702, n10703, n10704, n10705, n10706, n10708,
    n10709, n10710, n10711, n10712, n10713, n10714,
    n10715, n10716, n10717, n10718, n10719, n10720,
    n10721, n10722, n10723, n10724, n10725, n10726,
    n10727, n10728, n10729, n10730, n10731, n10732,
    n10733, n10734, n10735, n10736, n10737, n10738,
    n10739, n10740, n10741, n10742, n10743, n10744,
    n10745, n10746, n10747, n10748, n10749, n10750,
    n10751, n10752, n10753, n10754, n10755, n10756,
    n10757, n10758, n10759, n10760, n10761, n10762,
    n10763, n10764, n10765, n10766, n10767, n10768,
    n10769, n10770, n10771, n10772, n10773, n10774,
    n10775, n10776, n10777, n10778, n10779, n10780,
    n10781, n10782, n10783, n10784, n10785, n10786,
    n10787, n10788, n10789, n10790, n10791, n10792,
    n10793, n10794, n10795, n10796, n10797, n10798,
    n10799, n10800, n10801, n10802, n10803, n10804,
    n10805, n10806, n10807, n10808, n10809, n10810,
    n10811, n10812, n10813, n10814, n10815, n10816,
    n10817, n10818, n10819, n10820, n10821, n10822,
    n10823, n10824, n10825, n10826, n10827, n10828,
    n10829, n10830, n10831, n10832, n10833, n10834,
    n10835, n10836, n10837, n10838, n10839, n10840,
    n10841, n10842, n10843, n10844, n10845, n10846,
    n10847, n10848, n10849, n10850, n10851, n10852,
    n10853, n10854, n10855, n10856, n10857, n10858,
    n10859, n10860, n10861, n10862, n10863, n10864,
    n10865, n10866, n10867, n10868, n10869, n10870,
    n10871, n10872, n10873, n10874, n10875, n10876,
    n10877, n10878, n10879, n10880, n10881, n10882,
    n10883, n10884, n10886, n10887, n10888, n10889,
    n10890, n10891, n10892, n10893, n10894, n10895,
    n10896, n10897, n10898, n10899, n10900, n10901,
    n10902, n10903, n10904, n10905, n10906, n10907,
    n10908, n10909, n10910, n10911, n10912, n10913,
    n10914, n10915, n10916, n10917, n10918, n10919,
    n10920, n10921, n10922, n10923, n10924, n10925,
    n10926, n10927, n10928, n10929, n10930, n10931,
    n10932, n10933, n10934, n10935, n10936, n10937,
    n10938, n10939, n10940, n10941, n10942, n10943,
    n10944, n10945, n10946, n10947, n10948, n10949,
    n10950, n10951, n10952, n10953, n10954, n10955,
    n10956, n10957, n10959, n10960, n10961, n10963,
    n10964, n10965, n10966, n10967, n10968, n10969,
    n10970, n10971, n10972, n10973, n10974, n10975,
    n10976, n10977, n10978, n10979, n10980, n10981,
    n10983, n10984, n10985, n10986, n10987, n10988,
    n10989, n10990, n10991, n10992, n10993, n10994,
    n10995, n10996, n10997, n10998, n10999, n11000,
    n11001, n11002, n11003, n11004, n11005, n11006,
    n11007, n11008, n11009, n11010, n11011, n11012,
    n11013, n11014, n11015, n11016, n11017, n11018,
    n11019, n11020, n11021, n11022, n11023, n11024,
    n11025, n11026, n11028, n11029, n11030, n11031,
    n11032, n11034, n11035, n11036, n11037, n11038,
    n11039, n11040, n11041, n11042, n11043, n11044,
    n11045, n11046, n11047, n11048, n11049, n11050,
    n11051, n11053, n11054, n11055, n11056, n11057,
    n11058, n11059, n11060, n11061, n11062, n11063,
    n11064, n11065, n11066, n11067, n11068, n11069,
    n11070, n11071, n11072, n11073, n11074, n11075,
    n11076, n11077, n11079, n11080, n11081, n11082,
    n11083, n11084, n11085, n11087, n11088, n11089,
    n11090, n11091, n11092, n11093, n11094, n11095,
    n11096, n11097, n11098, n11099, n11100, n11101,
    n11102, n11103, n11104, n11105, n11106, n11107,
    n11108, n11109, n11110, n11111, n11112, n11113,
    n11114, n11115, n11116, n11117, n11118, n11119,
    n11120, n11121, n11122, n11123, n11124, n11125,
    n11126, n11127, n11128, n11129, n11130, n11131,
    n11132, n11133, n11134, n11135, n11136, n11137,
    n11138, n11139, n11140, n11141, n11142, n11143,
    n11144, n11145, n11146, n11147, n11148, n11149,
    n11150, n11151, n11152, n11153, n11154, n11155,
    n11156, n11157, n11158, n11159, n11160, n11161,
    n11162, n11163, n11164, n11165, n11166, n11167,
    n11168, n11169, n11170, n11171, n11172, n11173,
    n11174, n11175, n11176, n11177, n11178, n11179,
    n11180, n11181, n11182, n11183, n11184, n11185,
    n11186, n11187, n11188, n11189, n11190, n11191,
    n11192, n11193, n11194, n11195, n11196, n11197,
    n11198, n11199, n11200, n11201, n11202, n11203,
    n11204, n11205, n11206, n11207, n11208, n11209,
    n11210, n11211, n11212, n11213, n11214, n11215,
    n11216, n11217, n11218, n11219, n11220, n11221,
    n11222, n11223, n11224, n11225, n11226, n11227,
    n11228, n11229, n11230, n11231, n11232, n11233,
    n11234, n11235, n11236, n11238, n11239, n11240,
    n11241, n11242, n11243, n11244, n11245, n11246,
    n11247, n11248, n11250, n11251, n11252, n11253,
    n11254, n11255, n11256, n11257, n11258, n11259,
    n11260, n11261, n11262, n11263, n11264, n11265,
    n11266, n11267, n11268, n11270, n11271, n11272,
    n11273, n11274, n11275, n11276, n11277, n11278,
    n11279, n11280, n11281, n11282, n11284, n11285,
    n11286, n11287, n11288, n11289, n11290, n11292,
    n11293, n11294, n11295, n11296, n11297, n11298,
    n11299, n11300, n11302, n11303, n11305, n11306,
    n11307, n11308, n11309, n11311, n11312, n11313,
    n11314, n11315, n11316, n11317, n11318, n11320,
    n11321, n11322, n11323, n11325, n11326, n11327,
    n11328, n11330, n11331, n11332, n11333, n11334,
    n11336, n11337, n11338, n11339, n11340, n11341,
    n11342, n11344, n11345, n11346, n11348, n11349,
    n11350, n11351, n11352, n11353, n11354, n11355,
    n11356, n11357, n11358, n11359, n11360, n11361,
    n11362, n11363, n11365, n11366, n11367, n11368,
    n11370, n11371, n11372, n11373, n11374, n11375,
    n11376, n11378, n11379, n11380, n11381, n11382,
    n11383, n11384, n11385, n11386, n11387, n11388,
    n11389, n11391, n11392, n11393, n11394, n11395,
    n11396, n11397, n11398, n11399, n11400, n11401,
    n11402, n11403, n11404, n11405, n11406, n11407,
    n11408, n11409, n11411, n11412, n11413, n11414,
    n11415, n11416, n11417, n11418, n11419, n11420,
    n11421, n11422, n11423, n11424, n11425, n11426,
    n11427, n11428, n11429, n11430, n11431, n11433,
    n11434, n11435, n11436, n11437, n11438, n11439,
    n11440, n11441, n11442, n11443, n11444, n11445,
    n11446, n11448, n11449, n11450, n11451, n11452,
    n11453, n11454, n11455, n11456, n11457, n11458,
    n11460, n11461, n11462, n11463, n11464, n11465,
    n11466, n11467, n11468, n11469, n11470, n11471,
    n11472, n11473, n11475, n11476, n11477, n11478,
    n11479, n11480, n11481, n11482, n11483, n11484,
    n11486, n11487, n11488, n11489, n11490, n11491,
    n11492, n11493, n11494, n11495, n11496, n11497,
    n11498, n11499, n11500, n11501, n11502, n11503,
    n11504, n11505, n11506, n11507, n11508, n11509,
    n11510, n11511, n11512, n11513, n11514, n11515,
    n11516, n11517, n11518, n11519, n11520, n11521,
    n11522, n11523, n11524, n11525, n11526, n11527,
    n11528, n11529, n11530, n11531, n11532, n11533,
    n11534, n11535, n11536, n11537, n11538, n11539,
    n11540, n11541, n11542, n11543, n11544, n11545,
    n11546, n11547, n11548, n11549, n11550, n11551,
    n11552, n11553, n11554, n11555, n11556, n11557,
    n11558, n11559, n11560, n11561, n11562, n11563,
    n11564, n11565, n11566, n11567, n11568, n11569,
    n11570, n11571, n11572, n11573, n11574, n11575,
    n11576, n11577, n11578, n11579, n11580, n11581,
    n11582, n11583, n11584, n11585, n11586, n11587,
    n11588, n11589, n11590, n11591, n11592, n11593,
    n11594, n11595, n11596, n11597, n11598, n11599,
    n11600, n11601, n11602, n11603, n11604, n11605,
    n11606, n11607, n11608, n11609, n11610, n11611,
    n11612, n11613, n11614, n11615, n11616, n11617,
    n11618, n11619, n11620, n11621, n11622, n11623,
    n11624, n11625, n11626, n11627, n11628, n11629,
    n11630, n11631, n11632, n11633, n11634, n11635,
    n11636, n11637, n11639, n11640, n11641, n11642,
    n11643, n11644, n11645, n11646, n11647, n11649,
    n11651, n11652, n11653, n11654, n11655, n11656,
    n11657, n11658, n11659, n11660, n11661, n11662,
    n11663, n11664, n11665, n11666, n11667, n11668,
    n11669, n11670, n11671, n11672, n11673, n11674,
    n11675, n11676, n11677, n11678, n11679, n11680,
    n11681, n11682, n11683, n11684, n11685, n11686,
    n11687, n11688, n11689, n11690, n11691, n11692,
    n11693, n11694, n11695, n11696, n11697, n11698,
    n11699, n11700, n11701, n11702, n11703, n11704,
    n11705, n11706, n11707, n11708, n11709, n11710,
    n11711, n11712, n11713, n11714, n11715, n11716,
    n11717, n11718, n11719, n11720, n11721, n11722,
    n11723, n11724, n11725, n11726, n11727, n11728,
    n11729, n11730, n11731, n11732, n11733, n11734,
    n11735, n11736, n11737, n11738, n11739, n11740,
    n11741, n11742, n11743, n11744, n11745, n11746,
    n11747, n11748, n11749, n11750, n11751, n11752,
    n11753, n11754, n11755, n11756, n11757, n11758,
    n11759, n11760, n11761, n11762, n11763, n11764,
    n11765, n11766, n11767, n11768, n11769, n11770,
    n11771, n11772, n11773, n11774, n11775, n11776,
    n11777, n11778, n11779, n11780, n11781, n11782,
    n11783, n11784, n11785, n11786, n11787, n11788,
    n11789, n11790, n11791, n11792, n11793, n11794,
    n11795, n11796, n11797, n11798, n11799, n11800,
    n11801, n11802, n11803, n11804, n11805, n11806,
    n11807, n11808, n11809, n11810, n11811, n11812,
    n11813, n11814, n11815, n11816, n11817, n11818,
    n11819, n11820, n11821, n11822, n11823, n11824,
    n11825, n11826, n11827, n11828, n11829, n11830,
    n11831, n11832, n11833, n11834, n11835, n11836,
    n11837, n11838, n11839, n11840, n11841, n11842,
    n11843, n11844, n11845, n11846, n11847, n11848,
    n11849, n11850, n11851, n11852, n11853, n11854,
    n11855, n11856, n11857, n11858, n11859, n11860,
    n11861, n11862, n11863, n11864, n11865, n11866,
    n11867, n11868, n11869, n11870, n11871, n11872,
    n11873, n11874, n11875, n11876, n11877, n11878,
    n11879, n11880, n11881, n11882, n11883, n11884,
    n11885, n11886, n11887, n11888, n11889, n11890,
    n11891, n11892, n11893, n11894, n11895, n11896,
    n11897, n11898, n11899, n11900, n11901, n11902,
    n11903, n11904, n11905, n11906, n11907, n11908,
    n11909, n11910, n11911, n11912, n11913, n11914,
    n11915, n11916, n11917, n11918, n11919, n11920,
    n11921, n11922, n11923, n11924, n11925, n11926,
    n11927, n11928, n11929, n11930, n11931, n11932,
    n11933, n11934, n11935, n11936, n11937, n11938,
    n11939, n11940, n11941, n11942, n11943, n11944,
    n11945, n11946, n11947, n11948, n11949, n11950,
    n11951, n11952, n11953, n11954, n11955, n11956,
    n11957, n11958, n11959, n11960, n11961, n11962,
    n11963, n11964, n11965, n11966, n11967, n11968,
    n11969, n11970, n11971, n11972, n11973, n11974,
    n11975, n11976, n11977, n11978, n11979, n11980,
    n11981, n11982, n11983, n11984, n11985, n11986,
    n11987, n11988, n11989, n11990, n11991, n11992,
    n11993, n11994, n11995, n11996, n11997, n11998,
    n11999, n12000, n12001, n12002, n12003, n12004,
    n12005, n12006, n12007, n12008, n12009, n12010,
    n12011, n12012, n12013, n12014, n12015, n12016,
    n12017, n12018, n12019, n12020, n12021, n12022,
    n12023, n12024, n12025, n12026, n12027, n12028,
    n12029, n12030, n12031, n12032, n12033, n12034,
    n12035, n12036, n12037, n12038, n12039, n12040,
    n12041, n12042, n12043, n12044, n12045, n12046,
    n12047, n12048, n12049, n12050, n12051, n12052,
    n12053, n12054, n12055, n12056, n12057, n12058,
    n12059, n12060, n12061, n12062, n12063, n12064,
    n12065, n12066, n12067, n12068, n12069, n12070,
    n12071, n12072, n12073, n12074, n12075, n12076,
    n12077, n12078, n12079, n12080, n12081, n12082,
    n12083, n12084, n12085, n12086, n12087, n12088,
    n12089, n12090, n12091, n12092, n12093, n12094,
    n12095, n12096, n12097, n12098, n12099, n12100,
    n12101, n12102, n12103, n12104, n12105, n12106,
    n12107, n12108, n12109, n12110, n12111, n12112,
    n12113, n12114, n12115, n12116, n12117, n12118,
    n12119, n12120, n12121, n12122, n12123, n12124,
    n12125, n12126, n12127, n12128, n12129, n12130,
    n12131, n12132, n12133, n12134, n12135, n12136,
    n12137, n12138, n12139, n12140, n12141, n12142,
    n12143, n12144, n12145, n12146, n12147, n12148,
    n12149, n12150, n12151, n12152, n12154, n12155,
    n12156, n12157, n12158, n12159, n12160, n12161,
    n12162, n12163, n12164, n12165, n12166, n12167,
    n12168, n12169, n12170, n12171, n12172, n12173,
    n12174, n12175, n12176, n12177, n12178, n12179,
    n12180, n12181, n12182, n12183, n12184, n12185,
    n12186, n12187, n12188, n12189, n12190, n12191,
    n12192, n12193, n12194, n12195, n12196, n12197,
    n12198, n12199, n12200, n12201, n12202, n12203,
    n12204, n12205, n12206, n12207, n12208, n12209,
    n12210, n12211, n12212, n12213, n12214, n12215,
    n12216, n12217, n12218, n12219, n12220, n12221,
    n12222, n12223, n12224, n12225, n12226, n12227,
    n12228, n12229, n12230, n12231, n12232, n12233,
    n12234, n12235, n12236, n12237, n12238, n12239,
    n12240, n12241, n12242, n12243, n12244, n12245,
    n12246, n12247, n12248, n12249, n12250, n12251,
    n12252, n12253, n12254, n12255, n12256, n12257,
    n12258, n12259, n12260, n12261, n12262, n12263,
    n12264, n12265, n12266, n12267, n12268, n12269,
    n12270, n12271, n12272, n12273, n12274, n12275,
    n12276, n12277, n12278, n12279, n12280, n12281,
    n12282, n12283, n12284, n12285, n12286, n12287,
    n12288, n12289, n12290, n12291, n12292, n12293,
    n12294, n12295, n12296, n12297, n12298, n12299,
    n12300, n12301, n12302, n12303, n12304, n12305,
    n12306, n12307, n12308, n12309, n12310, n12311,
    n12312, n12313, n12314, n12315, n12316, n12317,
    n12318, n12319, n12320, n12321, n12322, n12323,
    n12324, n12325, n12326, n12327, n12328, n12329,
    n12330, n12331, n12332, n12333, n12334, n12335,
    n12336, n12337, n12338, n12339, n12340, n12341,
    n12342, n12343, n12344, n12345, n12346, n12347,
    n12348, n12349, n12350, n12351, n12352, n12353,
    n12354, n12355, n12356, n12357, n12358, n12359,
    n12360, n12361, n12362, n12363, n12364, n12365,
    n12366, n12367, n12368, n12369, n12370, n12371,
    n12372, n12373, n12374, n12375, n12376, n12377,
    n12378, n12379, n12380, n12381, n12382, n12383,
    n12384, n12385, n12386, n12387, n12388, n12389,
    n12390, n12391, n12392, n12393, n12394, n12395,
    n12396, n12397, n12398, n12399, n12400, n12401,
    n12402, n12403, n12404, n12405, n12406, n12407,
    n12408, n12409, n12410, n12411, n12412, n12413,
    n12414, n12415, n12416, n12417, n12418, n12419,
    n12420, n12421, n12422, n12423, n12424, n12425,
    n12426, n12427, n12428, n12429, n12430, n12431,
    n12432, n12433, n12434, n12435, n12436, n12437,
    n12438, n12439, n12440, n12441, n12442, n12443,
    n12444, n12445, n12446, n12447, n12448, n12449,
    n12450, n12451, n12452, n12453, n12454, n12455,
    n12456, n12457, n12458, n12459, n12460, n12461,
    n12462, n12463, n12464, n12465, n12466, n12467,
    n12468, n12469, n12470, n12471, n12472, n12473,
    n12474, n12475, n12476, n12477, n12478, n12479,
    n12480, n12481, n12482, n12483, n12484, n12485,
    n12486, n12487, n12488, n12489, n12490, n12491,
    n12492, n12493, n12494, n12495, n12496, n12497,
    n12498, n12499, n12500, n12501, n12502, n12503,
    n12504, n12505, n12506, n12507, n12508, n12509,
    n12510, n12511, n12512, n12513, n12514, n12515,
    n12516, n12517, n12518, n12519, n12520, n12521,
    n12522, n12523, n12524, n12525, n12526, n12527,
    n12528, n12529, n12530, n12531, n12532, n12533,
    n12534, n12535, n12536, n12537, n12538, n12539,
    n12540, n12541, n12542, n12543, n12544, n12545,
    n12546, n12547, n12548, n12549, n12550, n12551,
    n12552, n12553, n12554, n12555, n12556, n12557,
    n12558, n12559, n12560, n12561, n12562, n12563,
    n12564, n12565, n12566, n12567, n12568, n12569,
    n12570, n12571, n12572, n12573, n12574, n12575,
    n12576, n12577, n12578, n12579, n12580, n12581,
    n12582, n12583, n12584, n12585, n12586, n12587,
    n12588, n12589, n12590, n12591, n12592, n12593,
    n12594, n12595, n12596, n12597, n12598, n12599,
    n12600, n12601, n12602, n12603, n12604, n12605,
    n12606, n12607, n12608, n12609, n12610, n12611,
    n12612, n12613, n12614, n12615, n12616, n12617,
    n12618, n12619, n12620, n12621, n12622, n12623,
    n12624, n12625, n12626, n12627, n12628, n12629,
    n12630, n12631, n12632, n12633, n12634, n12635,
    n12636, n12637, n12638, n12639, n12640, n12641,
    n12642, n12643, n12644, n12645, n12646, n12647,
    n12648, n12649, n12650, n12651, n12652, n12653,
    n12654, n12655, n12656, n12657, n12658, n12659,
    n12660, n12661, n12662, n12663, n12664, n12665,
    n12666, n12667, n12668, n12669, n12670, n12671,
    n12672, n12673, n12674, n12675, n12676, n12677,
    n12678, n12679, n12680, n12681, n12682, n12683,
    n12684, n12685, n12686, n12687, n12688, n12689,
    n12690, n12691, n12692, n12693, n12694, n12695,
    n12696, n12697, n12698, n12699, n12700, n12701,
    n12702, n12703, n12704, n12705, n12706, n12707,
    n12708, n12709, n12710, n12711, n12712, n12713,
    n12714, n12715, n12716, n12717, n12718, n12719,
    n12720, n12721, n12722, n12723, n12724, n12725,
    n12726, n12727, n12728, n12729, n12730, n12731,
    n12732, n12733, n12734, n12735, n12736, n12737,
    n12738, n12739, n12740, n12741, n12742, n12743,
    n12744, n12745, n12746, n12747, n12748, n12749,
    n12750, n12751, n12752, n12753, n12754, n12755,
    n12756, n12757, n12758, n12759, n12760, n12761,
    n12762, n12763, n12764, n12765, n12766, n12767,
    n12768, n12769, n12770, n12771, n12772, n12773,
    n12774, n12775, n12776, n12777, n12778, n12779,
    n12780, n12781, n12782, n12783, n12784, n12785,
    n12786, n12787, n12788, n12789, n12790, n12791,
    n12792, n12793, n12794, n12795, n12796, n12797,
    n12798, n12799, n12800, n12801, n12802, n12803,
    n12804, n12805, n12806, n12807, n12808, n12809,
    n12810, n12811, n12812, n12813, n12814, n12815,
    n12816, n12817, n12818, n12819, n12820, n12821,
    n12822, n12823, n12824, n12825, n12826, n12827,
    n12828, n12829, n12830, n12831, n12832, n12833,
    n12834, n12835, n12836, n12837, n12838, n12839,
    n12840, n12841, n12842, n12843, n12844, n12845,
    n12846, n12847, n12848, n12849, n12850, n12851,
    n12852, n12853, n12854, n12855, n12856, n12857,
    n12858, n12859, n12860, n12861, n12862, n12863,
    n12864, n12865, n12866, n12867, n12868, n12869,
    n12870, n12871, n12872, n12873, n12874, n12875,
    n12876, n12877, n12878, n12879, n12880, n12881,
    n12882, n12883, n12884, n12885, n12886, n12887,
    n12888, n12889, n12890, n12891, n12892, n12893,
    n12894, n12895, n12896, n12897, n12898, n12899,
    n12900, n12901, n12902, n12903, n12904, n12905,
    n12906, n12907, n12908, n12909, n12910, n12911,
    n12912, n12913, n12914, n12915, n12916, n12917,
    n12918, n12919, n12920, n12921, n12922, n12923,
    n12924, n12925, n12926, n12927, n12928, n12929,
    n12930, n12931, n12932, n12933, n12934, n12935,
    n12936, n12937, n12938, n12939, n12940, n12941,
    n12942, n12943, n12944, n12945, n12946, n12947,
    n12948, n12949, n12950, n12951, n12952, n12953,
    n12954, n12955, n12956, n12957, n12958, n12959,
    n12960, n12961, n12962, n12963, n12964, n12965,
    n12966, n12967, n12968, n12969, n12970, n12971,
    n12972, n12973, n12974, n12975, n12976, n12977,
    n12978, n12979, n12980, n12981, n12982, n12983,
    n12984, n12985, n12986, n12987, n12988, n12989,
    n12990, n12991, n12993, n12994, n12995, n12996,
    n12997, n12998, n12999, n13000, n13001, n13003,
    n13004, n13005, n13006, n13007, n13008, n13009,
    n13011, n13012, n13013, n13014, n13015, n13016,
    n13017, n13018, n13019, n13020, n13021, n13022,
    n13023, n13025, n13026, n13027, n13028, n13029,
    n13031, n13032, n13033, n13034, n13036, n13037,
    n13038, n13040, n13041, n13042, n13044, n13045,
    n13046, n13047, n13048, n13049, n13050, n13051,
    n13052, n13053, n13054, n13055, n13056, n13057,
    n13058, n13059, n13060, n13061, n13062, n13064,
    n13065, n13066, n13067, n13068, n13069, n13070,
    n13071, n13072, n13074, n13075, n13076, n13077,
    n13079, n13080, n13081, n13082, n13083, n13084,
    n13085, n13086, n13087, n13088, n13089, n13091,
    n13092, n13093, n13094, n13095, n13096, n13097,
    n13098, n13099, n13100, n13101, n13103, n13104,
    n13105, n13106, n13107, n13108, n13110, n13111,
    n13112, n13113, n13114, n13115, n13116, n13117,
    n13118, n13119, n13120, n13121, n13122, n13123,
    n13124, n13125, n13126, n13128, n13129, n13130,
    n13131, n13132, n13133, n13134, n13135, n13136,
    n13137, n13138, n13139, n13140, n13141, n13142,
    n13144, n13145, n13146, n13147, n13148, n13149,
    n13150, n13151, n13152, n13153, n13155, n13156,
    n13157, n13158, n13159, n13160, n13161, n13162,
    n13163, n13165, n13166, n13167, n13168, n13170,
    n13171, n13172, n13173, n13174, n13175, n13176,
    n13177, n13178, n13179, n13180, n13181, n13182,
    n13183, n13184, n13185, n13186, n13187, n13188,
    n13189, n13190, n13191, n13192, n13193, n13194,
    n13195, n13196, n13197, n13198, n13199, n13200,
    n13201, n13202, n13203, n13204, n13205, n13206,
    n13207, n13208, n13209, n13210, n13211, n13212,
    n13213, n13214, n13215, n13216, n13217, n13218,
    n13219, n13220, n13221, n13222, n13223, n13224,
    n13225, n13226, n13227, n13228, n13229, n13230,
    n13231, n13232, n13233, n13234, n13235, n13236,
    n13237, n13238, n13239, n13240, n13241, n13242,
    n13243, n13244, n13245, n13247, n13248, n13249,
    n13250, n13251, n13252, n13253, n13254, n13255,
    n13256, n13257, n13258, n13259, n13260, n13261,
    n13262, n13264, n13265, n13266, n13267, n13268,
    n13269, n13270, n13271, n13272, n13273, n13274,
    n13275, n13276, n13277, n13278, n13279, n13280,
    n13281, n13282, n13283, n13284, n13285, n13286,
    n13287, n13288, n13289, n13290, n13291, n13292,
    n13293, n13294, n13295, n13296, n13297, n13298,
    n13299, n13300, n13301, n13302, n13303, n13304,
    n13305, n13306, n13307, n13308, n13309, n13310,
    n13311, n13312, n13313, n13314, n13315, n13316,
    n13317, n13318, n13319, n13320, n13321, n13322,
    n13323, n13324, n13325, n13326, n13327, n13328,
    n13329, n13330, n13331, n13332, n13333, n13334,
    n13335, n13336, n13337, n13338, n13339, n13340,
    n13341, n13342, n13343, n13345, n13347, n13348,
    n13349, n13350, n13351, n13352, n13353, n13355,
    n13356, n13357, n13358, n13359, n13360, n13361,
    n13362, n13363, n13364, n13365, n13366, n13367,
    n13368, n13369, n13370, n13371, n13373, n13374,
    n13375, n13376, n13377, n13378, n13379, n13380,
    n13381, n13383, n13385, n13386, n13387, n13388,
    n13389, n13390, n13391, n13392, n13393, n13394,
    n13395, n13396, n13397, n13398, n13399, n13400,
    n13401, n13403, n13405, n13406, n13407, n13408,
    n13409, n13410, n13411, n13412, n13413, n13414,
    n13416, n13417, n13418, n13419, n13420, n13423,
    n13424, n13425, n13426, n13427, n13428, n13429,
    n13430, n13431, n13432, n13433, n13434, n13435,
    n13436, n13437, n13438, n13439, n13440, n13441,
    n13442, n13443, n13444, n13445, n13446, n13447,
    n13448, n13449, n13450, n13451, n13452, n13453,
    n13454, n13455, n13456, n13457, n13458, n13459,
    n13460, n13461, n13462, n13463, n13464, n13465,
    n13466, n13467, n13468, n13469, n13470, n13471,
    n13472, n13474, n13475, n13476, n13477, n13478,
    n13479, n13480, n13481, n13482, n13483, n13484,
    n13485, n13486, n13487, n13488, n13489, n13490,
    n13491, n13492, n13493, n13494, n13495, n13496,
    n13497, n13498, n13499, n13500, n13501, n13502,
    n13503, n13504, n13505, n13506, n13507, n13508,
    n13509, n13510, n13511, n13512, n13513, n13514,
    n13515, n13517, n13518, n13519, n13520, n13521,
    n13522, n13523, n13524, n13525, n13526, n13527,
    n13528, n13529, n13530, n13531, n13532, n13533,
    n13534, n13535, n13536, n13537, n13538, n13539,
    n13540, n13541, n13542, n13543, n13544, n13545,
    n13546, n13547, n13548, n13549, n13550, n13551,
    n13552, n13553, n13554, n13555, n13556, n13557,
    n13559, n13560, n13561, n13562, n13563, n13564,
    n13565, n13566, n13567, n13568, n13569, n13570,
    n13571, n13572, n13573, n13574, n13575, n13576,
    n13577, n13578, n13579, n13580, n13581, n13582,
    n13583, n13584, n13585, n13586, n13587, n13588,
    n13589, n13590, n13591, n13592, n13593, n13594,
    n13595, n13596, n13597, n13598, n13599, n13600,
    n13601, n13602, n13603, n13604, n13605, n13606,
    n13607, n13608, n13610, n13611, n13612, n13613,
    n13614, n13615, n13616, n13617, n13618, n13619,
    n13620, n13621, n13622, n13623, n13624, n13626,
    n13627, n13628, n13629, n13630, n13631, n13632,
    n13633, n13634, n13635, n13636, n13637, n13638,
    n13639, n13640, n13641, n13642, n13643, n13644,
    n13645, n13646, n13647, n13648, n13649, n13650,
    n13651, n13652, n13653, n13654, n13655, n13656,
    n13657, n13658, n13659, n13660, n13661, n13662,
    n13663, n13664, n13665, n13666, n13667, n13668,
    n13669, n13670, n13671, n13672, n13673, n13674,
    n13675, n13676, n13677, n13678, n13679, n13680,
    n13681, n13682, n13683, n13684, n13685, n13686,
    n13687, n13688, n13689, n13690, n13691, n13692,
    n13693, n13694, n13695, n13696, n13697, n13698,
    n13699, n13700, n13701, n13702, n13703, n13704,
    n13705, n13706, n13707, n13708, n13709, n13710,
    n13711, n13712, n13713, n13714, n13715, n13716,
    n13717, n13718, n13719, n13720, n13721, n13722,
    n13723, n13724, n13725, n13726, n13727, n13728,
    n13729, n13730, n13731, n13732, n13733, n13734,
    n13735, n13736, n13737, n13738, n13739, n13740,
    n13741, n13742, n13743, n13744, n13745, n13746,
    n13747, n13748, n13749, n13750, n13751, n13752,
    n13753, n13754, n13755, n13756, n13757, n13758,
    n13759, n13760, n13761, n13762, n13763, n13764,
    n13765, n13766, n13767, n13768, n13769, n13770,
    n13771, n13772, n13773, n13774, n13775, n13776,
    n13777, n13778, n13779, n13780, n13781, n13782,
    n13783, n13784, n13785, n13786, n13787, n13788,
    n13789, n13790, n13791, n13792, n13793, n13794,
    n13795, n13796, n13797, n13798, n13799, n13800,
    n13801, n13802, n13803, n13804, n13805, n13806,
    n13807, n13808, n13809, n13810, n13811, n13812,
    n13813, n13814, n13815, n13816, n13817, n13818,
    n13819, n13820, n13821, n13822, n13823, n13824,
    n13825, n13826, n13827, n13828, n13829, n13830,
    n13831, n13832, n13833, n13834, n13835, n13836,
    n13837, n13838, n13839, n13840, n13841, n13842,
    n13843, n13844, n13845, n13846, n13847, n13848,
    n13849, n13850, n13851, n13852, n13853, n13854,
    n13855, n13856, n13857, n13858, n13859, n13860,
    n13861, n13862, n13863, n13864, n13865, n13866,
    n13867, n13868, n13869, n13870, n13871, n13872,
    n13873, n13874, n13875, n13876, n13877, n13878,
    n13879, n13880, n13881, n13882, n13883, n13884,
    n13885, n13886, n13887, n13888, n13889, n13890,
    n13891, n13892, n13893, n13894, n13895, n13896,
    n13897, n13898, n13899, n13900, n13901, n13902,
    n13903, n13904, n13905, n13906, n13907, n13908,
    n13909, n13910, n13911, n13912, n13913, n13914,
    n13915, n13916, n13917, n13918, n13919, n13920,
    n13921, n13922, n13923, n13924, n13925, n13926,
    n13927, n13928, n13930, n13931, n13932, n13933,
    n13934, n13935, n13936, n13937, n13938, n13939,
    n13940, n13941, n13942, n13943, n13944, n13945,
    n13946, n13947, n13948, n13949, n13950, n13951,
    n13952, n13953, n13954, n13955, n13956, n13957,
    n13958, n13959, n13960, n13961, n13962, n13963,
    n13964, n13965, n13966, n13967, n13968, n13969,
    n13970, n13971, n13972, n13973, n13974, n13975,
    n13976, n13977, n13978, n13979, n13980, n13981,
    n13982, n13983, n13985, n13986, n13987, n13988,
    n13989, n13990, n13991, n13992, n13993, n13994,
    n13995, n13996, n13997, n13998, n13999, n14000,
    n14001, n14002, n14003, n14004, n14005, n14006,
    n14007, n14008, n14009, n14010, n14011, n14012,
    n14013, n14014, n14015, n14016, n14017, n14018,
    n14019, n14020, n14021, n14022, n14023, n14024,
    n14025, n14026, n14027, n14028, n14029, n14030,
    n14031, n14032, n14033, n14034, n14035, n14036,
    n14037, n14038, n14039, n14040, n14041, n14042,
    n14043, n14044, n14045, n14046, n14047, n14048,
    n14049, n14050, n14051, n14052, n14053, n14054,
    n14055, n14056, n14057, n14058, n14059, n14060,
    n14061, n14062, n14063, n14064, n14065, n14066,
    n14067, n14068, n14069, n14070, n14071, n14072,
    n14073, n14074, n14075, n14076, n14077, n14078,
    n14079, n14080, n14081, n14082, n14083, n14084,
    n14085, n14086, n14087, n14088, n14089, n14090,
    n14091, n14092, n14093, n14094, n14095, n14096,
    n14097, n14098, n14099, n14100, n14101, n14102,
    n14103, n14104, n14105, n14106, n14107, n14108,
    n14109, n14110, n14111, n14112, n14113, n14114,
    n14115, n14116, n14117, n14118, n14119, n14120,
    n14121, n14122, n14123, n14124, n14125, n14126,
    n14127, n14128, n14129, n14130, n14131, n14132,
    n14133, n14134, n14135, n14136, n14137, n14138,
    n14139, n14140, n14141, n14142, n14143, n14144,
    n14145, n14146, n14147, n14148, n14149, n14150,
    n14151, n14152, n14153, n14154, n14155, n14156,
    n14157, n14158, n14159, n14160, n14161, n14162,
    n14163, n14164, n14165, n14166, n14167, n14168,
    n14169, n14170, n14171, n14172, n14173, n14174,
    n14175, n14176, n14177, n14178, n14179, n14180,
    n14181, n14182, n14183, n14184, n14185, n14186,
    n14187, n14188, n14189, n14190, n14191, n14192,
    n14193, n14194, n14195, n14196, n14197, n14198,
    n14199, n14200, n14201, n14202, n14203, n14204,
    n14205, n14206, n14207, n14208, n14209, n14210,
    n14211, n14212, n14213, n14214, n14215, n14216,
    n14217, n14218, n14219, n14220, n14221, n14222,
    n14223, n14224, n14225, n14226, n14227, n14228,
    n14229, n14230, n14231, n14232, n14233, n14234,
    n14235, n14236, n14237, n14238, n14239, n14240,
    n14241, n14242, n14243, n14244, n14245, n14246,
    n14247, n14248, n14249, n14250, n14251, n14252,
    n14253, n14254, n14255, n14256, n14257, n14258,
    n14259, n14260, n14261, n14262, n14263, n14264,
    n14265, n14266, n14267, n14268, n14269, n14270,
    n14271, n14272, n14273, n14274, n14275, n14276,
    n14277, n14278, n14279, n14280, n14281, n14282,
    n14283, n14284, n14285, n14286, n14287, n14288,
    n14289, n14290, n14291, n14292, n14293, n14294,
    n14295, n14296, n14297, n14298, n14299, n14300,
    n14301, n14302, n14303, n14304, n14305, n14306,
    n14307, n14308, n14309, n14310, n14311, n14312,
    n14313, n14314, n14315, n14316, n14317, n14318,
    n14319, n14320, n14321, n14322, n14323, n14324,
    n14325, n14326, n14327, n14328, n14329, n14330,
    n14331, n14332, n14333, n14334, n14335, n14336,
    n14337, n14338, n14339, n14340, n14341, n14342,
    n14343, n14344, n14345, n14346, n14347, n14348,
    n14349, n14350, n14351, n14352, n14353, n14354,
    n14355, n14356, n14357, n14358, n14359, n14360,
    n14361, n14362, n14363, n14364, n14365, n14366,
    n14367, n14368, n14369, n14370, n14371, n14372,
    n14373, n14374, n14375, n14376, n14377, n14378,
    n14379, n14380, n14382, n14383, n14384, n14385,
    n14386, n14387, n14388, n14389, n14390, n14391,
    n14392, n14393, n14394, n14395, n14396, n14397,
    n14398, n14399, n14400, n14401, n14402, n14403,
    n14404, n14405, n14406, n14407, n14408, n14409,
    n14410, n14411, n14412, n14413, n14414, n14415,
    n14416, n14417, n14418, n14419, n14420, n14421,
    n14422, n14423, n14424, n14425, n14426, n14427,
    n14428, n14429, n14430, n14431, n14432, n14433,
    n14434, n14435, n14436, n14437, n14438, n14439,
    n14440, n14441, n14442, n14443, n14444, n14445,
    n14446, n14447, n14448, n14449, n14450, n14451,
    n14452, n14453, n14454, n14455, n14456, n14457,
    n14458, n14459, n14460, n14461, n14462, n14463,
    n14464, n14465, n14466, n14467, n14468, n14469,
    n14470, n14471, n14472, n14473, n14474, n14475,
    n14476, n14477, n14478, n14479, n14480, n14481,
    n14482, n14483, n14484, n14485, n14486, n14487,
    n14488, n14489, n14490, n14491, n14492, n14493,
    n14494, n14495, n14496, n14497, n14498, n14499,
    n14500, n14501, n14502, n14503, n14504, n14505,
    n14506, n14507, n14508, n14509, n14510, n14511,
    n14512, n14513, n14514, n14515, n14516, n14517,
    n14518, n14519, n14520, n14521, n14522, n14523,
    n14524, n14525, n14526, n14527, n14528, n14529,
    n14530, n14531, n14532, n14533, n14534, n14535,
    n14536, n14537, n14538, n14539, n14540, n14541,
    n14542, n14543, n14544, n14545, n14546, n14547,
    n14548, n14549, n14550, n14551, n14552, n14553,
    n14554, n14555, n14556, n14557, n14558, n14559,
    n14560, n14561, n14562, n14563, n14564, n14565,
    n14566, n14567, n14568, n14569, n14570, n14571,
    n14572, n14573, n14574, n14575, n14576, n14577,
    n14578, n14579, n14580, n14581, n14582, n14583,
    n14584, n14585, n14586, n14587, n14588, n14589,
    n14590, n14591, n14592, n14593, n14594, n14595,
    n14596, n14597, n14598, n14599, n14600, n14601,
    n14602, n14603, n14604, n14605, n14606, n14607,
    n14608, n14609, n14610, n14611, n14612, n14613,
    n14614, n14615, n14616, n14617, n14618, n14619,
    n14620, n14621, n14622, n14623, n14624, n14625,
    n14626, n14627, n14628, n14629, n14630, n14631,
    n14632, n14633, n14634, n14635, n14636, n14637,
    n14638, n14639, n14640, n14641, n14642, n14643,
    n14644, n14645, n14646, n14647, n14648, n14649,
    n14650, n14651, n14652, n14653, n14654, n14655,
    n14656, n14657, n14658, n14659, n14660, n14661,
    n14662, n14663, n14664, n14665, n14666, n14667,
    n14668, n14669, n14670, n14671, n14672, n14673,
    n14674, n14675, n14676, n14677, n14678, n14679,
    n14680, n14681, n14682, n14683, n14684, n14685,
    n14686, n14687, n14688, n14689, n14690, n14691,
    n14692, n14693, n14694, n14695, n14696, n14697,
    n14698, n14699, n14700, n14701, n14702, n14703,
    n14704, n14705, n14706, n14707, n14708, n14709,
    n14710, n14711, n14712, n14713, n14714, n14715,
    n14716, n14717, n14718, n14719, n14720, n14721,
    n14722, n14723, n14724, n14725, n14726, n14727,
    n14728, n14729, n14730, n14731, n14732, n14733,
    n14734, n14735, n14736, n14737, n14738, n14739,
    n14740, n14741, n14742, n14743, n14744, n14745,
    n14746, n14747, n14748, n14749, n14750, n14751,
    n14752, n14753, n14754, n14755, n14756, n14757,
    n14758, n14759, n14760, n14761, n14762, n14763,
    n14764, n14765, n14766, n14767, n14768, n14769,
    n14770, n14771, n14772, n14773, n14774, n14775,
    n14776, n14777, n14778, n14779, n14780, n14781,
    n14782, n14783, n14784, n14785, n14786, n14787,
    n14788, n14789, n14790, n14791, n14792, n14793,
    n14794, n14795, n14796, n14797, n14798, n14799,
    n14801, n14802, n14803, n14804, n14805, n14806,
    n14807, n14809, n14810, n14811, n14812, n14813,
    n14814, n14815, n14816, n14817, n14818, n14819,
    n14820, n14821, n14822, n14823, n14824, n14825,
    n14826, n14827, n14828, n14829, n14830, n14831,
    n14832, n14833, n14834, n14835, n14836, n14837,
    n14838, n14839, n14840, n14841, n14842, n14843,
    n14844, n14845, n14846, n14847, n14848, n14849,
    n14850, n14851, n14852, n14853, n14854, n14855,
    n14856, n14857, n14858, n14859, n14860, n14861,
    n14863, n14864, n14865, n14866, n14867, n14868,
    n14869, n14870, n14871, n14872, n14873, n14874,
    n14875, n14876, n14877, n14878, n14879, n14880,
    n14881, n14882, n14883, n14884, n14885, n14886,
    n14887, n14888, n14889, n14890, n14891, n14892,
    n14893, n14894, n14895, n14896, n14897, n14898,
    n14899, n14900, n14901, n14902, n14903, n14904,
    n14905, n14906, n14907, n14908, n14909, n14910,
    n14911, n14912, n14913, n14914, n14915, n14916,
    n14917, n14918, n14919, n14920, n14921, n14922,
    n14923, n14924, n14925, n14926, n14927, n14928,
    n14929, n14930, n14931, n14932, n14933, n14934,
    n14935, n14936, n14937, n14938, n14939, n14940,
    n14941, n14942, n14943, n14944, n14945, n14946,
    n14947, n14948, n14949, n14950, n14951, n14952,
    n14953, n14954, n14955, n14956, n14957, n14958,
    n14959, n14960, n14961, n14962, n14963, n14964,
    n14965, n14966, n14967, n14968, n14969, n14970,
    n14971, n14972, n14973, n14974, n14975, n14976,
    n14977, n14978, n14979, n14980, n14981, n14982,
    n14983, n14984, n14985, n14986, n14987, n14988,
    n14989, n14990, n14991, n14992, n14993, n14994,
    n14995, n14996, n14997, n14998, n14999, n15000,
    n15001, n15002, n15003, n15004, n15005, n15006,
    n15007, n15008, n15009, n15010, n15011, n15012,
    n15013, n15014, n15015, n15016, n15017, n15018,
    n15019, n15020, n15021, n15022, n15023, n15024,
    n15025, n15026, n15027, n15028, n15029, n15030,
    n15031, n15032, n15033, n15034, n15035, n15036,
    n15037, n15038, n15039, n15040, n15041, n15042,
    n15043, n15044, n15045, n15046, n15047, n15048,
    n15049, n15050, n15051, n15052, n15053, n15054,
    n15055, n15056, n15057, n15058, n15059, n15060,
    n15061, n15062, n15063, n15064, n15065, n15066,
    n15067, n15068, n15069, n15070, n15071, n15072,
    n15073, n15074, n15075, n15076, n15077, n15078,
    n15079, n15080, n15081, n15082, n15083, n15084,
    n15085, n15086, n15087, n15088, n15089, n15090,
    n15091, n15092, n15093, n15094, n15095, n15096,
    n15097, n15098, n15099, n15100, n15101, n15102,
    n15103, n15104, n15105, n15106, n15107, n15108,
    n15109, n15110, n15111, n15112, n15113, n15114,
    n15115, n15116, n15117, n15118, n15119, n15120,
    n15121, n15122, n15123, n15124, n15125, n15126,
    n15127, n15128, n15129, n15130, n15131, n15132,
    n15133, n15134, n15135, n15136, n15137, n15138,
    n15139, n15140, n15141, n15142, n15143, n15144,
    n15145, n15146, n15147, n15148, n15149, n15150,
    n15151, n15152, n15153, n15154, n15155, n15156,
    n15157, n15158, n15159, n15160, n15161, n15162,
    n15163, n15164, n15165, n15166, n15167, n15168,
    n15169, n15170, n15171, n15172, n15173, n15174,
    n15175, n15176, n15177, n15178, n15179, n15180,
    n15181, n15182, n15183, n15184, n15185, n15186,
    n15187, n15188, n15189, n15190, n15191, n15192,
    n15193, n15194, n15195, n15196, n15197, n15198,
    n15199, n15200, n15201, n15202, n15203, n15204,
    n15205, n15206, n15207, n15208, n15209, n15210,
    n15211, n15212, n15213, n15214, n15215, n15216,
    n15217, n15218, n15219, n15220, n15221, n15222,
    n15223, n15224, n15225, n15226, n15227, n15228,
    n15229, n15230, n15231, n15232, n15233, n15234,
    n15235, n15236, n15237, n15238, n15239, n15240,
    n15241, n15242, n15243, n15244, n15245, n15246,
    n15247, n15248, n15249, n15250, n15251, n15252,
    n15253, n15254, n15255, n15256, n15257, n15258,
    n15259, n15260, n15261, n15262, n15263, n15264,
    n15265, n15267, n15268, n15269, n15270, n15271,
    n15272, n15273, n15274, n15275, n15276, n15277,
    n15278, n15279, n15280, n15281, n15282, n15283,
    n15284, n15285, n15286, n15287, n15288, n15289,
    n15290, n15291, n15292, n15293, n15294, n15295,
    n15296, n15297, n15298, n15299, n15300, n15301,
    n15302, n15303, n15304, n15305, n15306, n15307,
    n15308, n15309, n15310, n15311, n15312, n15313,
    n15314, n15315, n15316, n15317, n15318, n15319,
    n15320, n15321, n15322, n15323, n15324, n15325,
    n15326, n15327, n15328, n15329, n15330, n15331,
    n15332, n15333, n15334, n15335, n15336, n15337,
    n15338, n15339, n15340, n15341, n15342, n15343,
    n15344, n15345, n15346, n15347, n15348, n15349,
    n15350, n15351, n15352, n15353, n15354, n15355,
    n15356, n15357, n15358, n15359, n15360, n15361,
    n15362, n15363, n15364, n15365, n15366, n15367,
    n15368, n15369, n15370, n15371, n15372, n15373,
    n15374, n15375, n15376, n15377, n15378, n15379,
    n15380, n15381, n15382, n15383, n15384, n15385,
    n15386, n15387, n15388, n15389, n15390, n15391,
    n15392, n15393, n15394, n15395, n15396, n15397,
    n15398, n15399, n15400, n15401, n15402, n15403,
    n15404, n15405, n15406, n15407, n15408, n15409,
    n15410, n15411, n15412, n15413, n15414, n15415,
    n15416, n15417, n15418, n15419, n15420, n15421,
    n15422, n15423, n15424, n15425, n15426, n15427,
    n15428, n15429, n15430, n15431, n15432, n15433,
    n15434, n15435, n15436, n15437, n15438, n15439,
    n15440, n15441, n15442, n15443, n15444, n15445,
    n15446, n15447, n15448, n15449, n15450, n15451,
    n15452, n15453, n15454, n15455, n15456, n15457,
    n15458, n15459, n15460, n15461, n15462, n15463,
    n15464, n15465, n15466, n15467, n15468, n15469,
    n15470, n15471, n15472, n15473, n15474, n15475,
    n15476, n15477, n15478, n15479, n15480, n15481,
    n15482, n15483, n15484, n15485, n15486, n15487,
    n15488, n15489, n15490, n15491, n15492, n15493,
    n15494, n15495, n15496, n15497, n15498, n15499,
    n15500, n15501, n15502, n15503, n15504, n15505,
    n15506, n15507, n15508, n15509, n15510, n15511,
    n15512, n15513, n15514, n15515, n15516, n15517,
    n15518, n15519, n15520, n15521, n15522, n15523,
    n15524, n15525, n15526, n15527, n15528, n15529,
    n15530, n15531, n15532, n15533, n15534, n15535,
    n15536, n15537, n15538, n15539, n15540, n15541,
    n15542, n15543, n15544, n15545, n15546, n15547,
    n15548, n15549, n15550, n15551, n15552, n15553,
    n15554, n15555, n15556, n15557, n15558, n15559,
    n15560, n15561, n15562, n15563, n15564, n15565,
    n15566, n15567, n15569, n15570, n15571, n15572,
    n15573, n15574, n15575, n15576, n15577, n15578,
    n15579, n15580, n15581, n15582, n15583, n15584,
    n15585, n15586, n15587, n15588, n15589, n15590,
    n15591, n15592, n15593, n15594, n15595, n15596,
    n15597, n15598, n15599, n15600, n15601, n15602,
    n15603, n15604, n15605, n15606, n15607, n15608,
    n15609, n15610, n15611, n15612, n15613, n15614,
    n15615, n15616, n15617, n15618, n15619, n15620,
    n15621, n15622, n15623, n15624, n15625, n15626,
    n15627, n15628, n15629, n15630, n15631, n15632,
    n15633, n15634, n15635, n15636, n15637, n15638,
    n15639, n15640, n15641, n15642, n15643, n15644,
    n15645, n15646, n15647, n15648, n15649, n15650,
    n15651, n15652, n15653, n15654, n15655, n15656,
    n15657, n15658, n15659, n15660, n15661, n15663,
    n15664, n15665, n15666, n15667, n15668, n15669,
    n15670, n15671, n15672, n15673, n15674, n15675,
    n15676, n15677, n15678, n15679, n15680, n15681,
    n15682, n15683, n15684, n15685, n15686, n15688,
    n15689, n15690, n15691, n15692, n15693, n15694,
    n15695, n15696, n15697, n15698, n15699, n15700,
    n15701, n15702, n15703, n15704, n15705, n15706,
    n15707, n15708, n15709, n15710, n15711, n15712,
    n15713, n15714, n15715, n15716, n15717, n15718,
    n15719, n15720, n15721, n15722, n15723, n15724,
    n15725, n15726, n15727, n15728, n15729, n15730,
    n15731, n15732, n15733, n15734, n15735, n15736,
    n15737, n15738, n15739, n15740, n15741, n15742,
    n15743, n15744, n15745, n15746, n15747, n15748,
    n15749, n15750, n15751, n15752, n15753, n15754,
    n15755, n15756, n15757, n15758, n15759, n15760,
    n15761, n15762, n15763, n15764, n15765, n15766,
    n15767, n15768, n15769, n15770, n15771, n15772,
    n15773, n15774, n15775, n15776, n15777, n15778,
    n15779, n15780, n15781, n15782, n15783, n15784,
    n15785, n15786, n15787, n15788, n15789, n15790,
    n15791, n15792, n15793, n15794, n15795, n15796,
    n15797, n15798, n15799, n15800, n15801, n15802,
    n15803, n15804, n15805, n15806, n15807, n15808,
    n15809, n15810, n15811, n15812, n15813, n15814,
    n15815, n15816, n15817, n15818, n15819, n15820,
    n15821, n15823, n15824, n15825, n15826, n15827,
    n15828, n15829, n15831, n15832, n15833, n15834,
    n15835, n15836, n15837, n15838, n15839, n15840,
    n15841, n15842, n15843, n15844, n15845, n15846,
    n15847, n15848, n15849, n15850, n15851, n15852,
    n15853, n15854, n15855, n15856, n15857, n15858,
    n15859, n15860, n15861, n15862, n15863, n15864,
    n15865, n15866, n15867, n15868, n15869, n15870,
    n15871, n15872, n15873, n15874, n15875, n15876,
    n15877, n15878, n15879, n15880, n15881, n15882,
    n15883, n15884, n15885, n15886, n15887, n15888,
    n15889, n15890, n15891, n15892, n15893, n15894,
    n15895, n15896, n15897, n15898, n15899, n15900,
    n15901, n15902, n15903, n15904, n15905, n15906,
    n15907, n15908, n15909, n15910, n15911, n15912,
    n15913, n15914, n15915, n15916, n15917, n15918,
    n15919, n15920, n15921, n15922, n15923, n15924,
    n15925, n15926, n15927, n15928, n15929, n15930,
    n15931, n15932, n15933, n15934, n15935, n15936,
    n15937, n15938, n15939, n15940, n15941, n15942,
    n15943, n15944, n15945, n15946, n15947, n15948,
    n15949, n15950, n15951, n15952, n15953, n15954,
    n15955, n15956, n15957, n15958, n15959, n15960,
    n15961, n15962, n15963, n15964, n15965, n15966,
    n15967, n15968, n15969, n15970, n15971, n15972,
    n15973, n15974, n15975, n15976, n15977, n15978,
    n15979, n15980, n15981, n15982, n15983, n15984,
    n15985, n15986, n15987, n15988, n15989, n15990,
    n15991, n15992, n15993, n15994, n15995, n15996,
    n15997, n15998, n15999, n16000, n16001, n16002,
    n16003, n16004, n16005, n16006, n16007, n16008,
    n16009, n16010, n16011, n16012, n16013, n16014,
    n16015, n16016, n16017, n16018, n16019, n16020,
    n16021, n16022, n16023, n16024, n16025, n16026,
    n16027, n16028, n16029, n16030, n16031, n16032,
    n16033, n16034, n16035, n16036, n16037, n16038,
    n16039, n16040, n16041, n16042, n16043, n16044,
    n16045, n16047, n16048, n16049, n16050, n16051,
    n16052, n16053, n16054, n16055, n16056, n16057,
    n16058, n16059, n16060, n16061, n16062, n16063,
    n16064, n16065, n16066, n16067, n16068, n16069,
    n16070, n16071, n16072, n16073, n16074, n16075,
    n16076, n16077, n16078, n16079, n16080, n16081,
    n16082, n16083, n16084, n16085, n16086, n16087,
    n16088, n16089, n16090, n16091, n16092, n16093,
    n16094, n16095, n16096, n16097, n16098, n16099,
    n16100, n16101, n16102, n16103, n16104, n16105,
    n16107, n16108, n16109, n16110, n16111, n16112,
    n16113, n16114, n16115, n16116, n16117, n16118,
    n16119, n16120, n16121, n16122, n16123, n16124,
    n16125, n16126, n16127, n16128, n16129, n16130,
    n16131, n16132, n16133, n16134, n16135, n16136,
    n16137, n16138, n16139, n16140, n16141, n16142,
    n16143, n16144, n16145, n16146, n16147, n16148,
    n16149, n16150, n16151, n16152, n16153, n16154,
    n16155, n16156, n16157, n16158, n16159, n16160,
    n16161, n16162, n16163, n16164, n16165, n16166,
    n16167, n16168, n16169, n16170, n16171, n16172,
    n16173, n16174, n16175, n16176, n16177, n16178,
    n16179, n16180, n16181, n16182, n16183, n16184,
    n16185, n16186, n16187, n16188, n16189, n16190,
    n16191, n16192, n16193, n16194, n16195, n16196,
    n16197, n16198, n16199, n16200, n16201, n16202,
    n16203, n16204, n16205, n16206, n16207, n16208,
    n16209, n16210, n16211, n16212, n16213, n16214,
    n16215, n16216, n16217, n16218, n16219, n16221,
    n16222, n16223, n16224, n16225, n16226, n16227,
    n16228, n16229, n16230, n16231, n16232, n16233,
    n16234, n16235, n16236, n16237, n16238, n16239,
    n16240, n16241, n16242, n16243, n16244, n16245,
    n16246, n16247, n16248, n16249, n16250, n16251,
    n16252, n16253, n16254, n16255, n16256, n16257,
    n16258, n16259, n16260, n16261, n16262, n16263,
    n16264, n16265, n16266, n16267, n16268, n16269,
    n16270, n16271, n16272, n16273, n16274, n16275,
    n16276, n16277, n16278, n16279, n16280, n16281,
    n16282, n16283, n16284, n16285, n16286, n16287,
    n16288, n16289, n16290, n16291, n16292, n16293,
    n16294, n16295, n16296, n16297, n16298, n16299,
    n16300, n16301, n16302, n16303, n16304, n16305,
    n16306, n16307, n16308, n16309, n16310, n16311,
    n16312, n16313, n16314, n16315, n16316, n16317,
    n16318, n16319, n16320, n16321, n16322, n16323,
    n16324, n16325, n16326, n16327, n16328, n16329,
    n16330, n16331, n16332, n16333, n16334, n16335,
    n16336, n16337, n16338, n16340, n16341, n16342,
    n16343, n16344, n16345, n16346, n16347, n16348,
    n16349, n16350, n16351, n16352, n16353, n16354,
    n16355, n16356, n16357, n16358, n16359, n16360,
    n16361, n16362, n16363, n16364, n16365, n16366,
    n16367, n16368, n16369, n16370, n16371, n16372,
    n16373, n16374, n16375, n16376, n16377, n16378,
    n16379, n16380, n16381, n16382, n16383, n16384,
    n16385, n16386, n16387, n16388, n16389, n16390,
    n16391, n16392, n16393, n16394, n16395, n16396,
    n16397, n16398, n16399, n16400, n16401, n16402,
    n16403, n16404, n16405, n16406, n16407, n16408,
    n16409, n16410, n16411, n16412, n16413, n16414,
    n16415, n16416, n16417, n16418, n16419, n16420,
    n16421, n16422, n16423, n16424, n16426, n16427,
    n16428, n16429, n16430, n16431, n16432, n16433,
    n16434, n16435, n16436, n16437, n16439, n16440,
    n16441, n16442, n16443, n16444, n16445, n16446,
    n16447, n16448, n16449, n16450, n16451, n16452,
    n16453, n16454, n16455, n16456, n16457, n16458,
    n16459, n16460, n16461, n16462, n16463, n16464,
    n16465, n16466, n16467, n16468, n16469, n16470,
    n16471, n16472, n16473, n16474, n16475, n16476,
    n16477, n16478, n16479, n16480, n16481, n16482,
    n16483, n16484, n16485, n16486, n16487, n16488,
    n16489, n16490, n16491, n16492, n16493, n16494,
    n16495, n16496, n16497, n16498, n16499, n16500,
    n16501, n16502, n16503, n16504, n16505, n16506,
    n16507, n16508, n16509, n16510, n16511, n16512,
    n16513, n16514, n16515, n16516, n16517, n16518,
    n16519, n16520, n16521, n16522, n16524, n16525,
    n16526, n16527, n16528, n16529, n16530, n16531,
    n16532, n16533, n16534, n16535, n16536, n16537,
    n16538, n16539, n16540, n16541, n16542, n16543,
    n16544, n16545, n16546, n16547, n16548, n16549,
    n16550, n16551, n16552, n16553, n16554, n16555,
    n16556, n16557, n16558, n16559, n16560, n16561,
    n16562, n16563, n16564, n16565, n16566, n16567,
    n16568, n16569, n16570, n16571, n16572, n16573,
    n16574, n16575, n16576, n16578, n16579, n16580,
    n16581, n16582, n16583, n16584, n16585, n16586,
    n16587, n16588, n16589, n16590, n16591, n16592,
    n16593, n16594, n16595, n16596, n16597, n16598,
    n16599, n16600, n16601, n16602, n16603, n16604,
    n16605, n16606, n16607, n16608, n16609, n16610,
    n16611, n16612, n16613, n16614, n16615, n16616,
    n16617, n16618, n16619, n16620, n16621, n16622,
    n16624, n16625, n16626, n16627, n16628, n16629,
    n16630, n16631, n16632, n16633, n16634, n16635,
    n16636, n16637, n16638, n16639, n16640, n16641,
    n16642, n16643, n16644, n16645, n16646, n16647,
    n16648, n16649, n16650, n16651, n16652, n16653,
    n16654, n16655, n16656, n16657, n16658, n16659,
    n16660, n16661, n16662, n16663, n16664, n16665,
    n16666, n16667, n16668, n16669, n16670, n16671,
    n16672, n16673, n16674, n16675, n16676, n16677,
    n16678, n16679, n16680, n16681, n16682, n16683,
    n16684, n16685, n16686, n16687, n16688, n16689,
    n16690, n16691, n16692, n16693, n16694, n16695,
    n16696, n16697, n16698, n16699, n16700, n16701,
    n16702, n16703, n16704, n16705, n16706, n16707,
    n16708, n16709, n16710, n16711, n16712, n16713,
    n16714, n16715, n16716, n16717, n16718, n16719,
    n16720, n16721, n16722, n16723, n16724, n16725,
    n16726, n16727, n16728, n16729, n16730, n16731,
    n16732, n16733, n16734, n16735, n16736, n16737,
    n16738, n16739, n16740, n16741, n16742, n16743,
    n16744, n16745, n16746, n16747, n16748, n16749,
    n16750, n16751, n16752, n16753, n16754, n16755,
    n16756, n16757, n16758, n16759, n16760, n16761,
    n16762, n16763, n16764, n16765, n16766, n16767,
    n16768, n16769, n16770, n16771, n16772, n16773,
    n16774, n16775, n16776, n16777, n16778, n16779,
    n16780, n16781, n16782, n16783, n16784, n16785,
    n16786, n16787, n16788, n16789, n16790, n16791,
    n16792, n16793, n16794, n16795, n16796, n16797,
    n16798, n16799, n16800, n16801, n16802, n16803,
    n16804, n16805, n16806, n16807, n16808, n16809,
    n16810, n16811, n16812, n16813, n16814, n16815,
    n16816, n16817, n16818, n16819, n16820, n16821,
    n16822, n16823, n16824, n16825, n16826, n16827,
    n16828, n16829, n16830, n16831, n16832, n16833,
    n16834, n16835, n16836, n16837, n16838, n16839,
    n16840, n16841, n16842, n16843, n16844, n16845,
    n16846, n16847, n16848, n16849, n16850, n16851,
    n16852, n16853, n16854, n16855, n16856, n16857,
    n16858, n16859, n16860, n16861, n16862, n16863,
    n16864, n16865, n16866, n16867, n16868, n16869,
    n16870, n16871, n16872, n16873, n16874, n16875,
    n16876, n16877, n16878, n16879, n16880, n16881,
    n16882, n16883, n16884, n16885, n16886, n16887,
    n16888, n16889, n16890, n16891, n16892, n16893,
    n16894, n16895, n16896, n16897, n16898, n16899,
    n16900, n16901, n16902, n16903, n16904, n16905,
    n16906, n16907, n16908, n16909, n16910, n16911,
    n16912, n16913, n16914, n16915, n16916, n16917,
    n16918, n16919, n16920, n16921, n16922, n16923,
    n16924, n16925, n16926, n16927, n16928, n16929,
    n16930, n16931, n16932, n16933, n16934, n16935,
    n16936, n16937, n16938, n16939, n16940, n16941,
    n16942, n16943, n16944, n16945, n16946, n16947,
    n16948, n16949, n16950, n16951, n16952, n16953,
    n16954, n16955, n16956, n16957, n16958, n16959,
    n16960, n16961, n16962, n16963, n16964, n16965,
    n16966, n16967, n16968, n16969, n16970, n16971,
    n16972, n16973, n16974, n16975, n16976, n16977,
    n16978, n16979, n16980, n16981, n16982, n16983,
    n16984, n16985, n16986, n16987, n16988, n16989,
    n16990, n16991, n16992, n16993, n16994, n16995,
    n16996, n16997, n16998, n16999, n17000, n17001,
    n17002, n17003, n17004, n17005, n17006, n17007,
    n17008, n17009, n17010, n17011, n17012, n17013,
    n17014, n17015, n17016, n17017, n17018, n17019,
    n17020, n17021, n17022, n17023, n17024, n17025,
    n17026, n17027, n17028, n17029, n17030, n17031,
    n17032, n17033, n17034, n17035, n17036, n17037,
    n17038, n17039, n17040, n17041, n17042, n17043,
    n17044, n17045, n17046, n17047, n17048, n17049,
    n17050, n17051, n17052, n17053, n17054, n17055,
    n17056, n17057, n17058, n17059, n17060, n17061,
    n17062, n17063, n17064, n17065, n17066, n17067,
    n17068, n17069, n17070, n17071, n17072, n17073,
    n17074, n17075, n17076, n17077, n17078, n17079,
    n17080, n17081, n17082, n17083, n17084, n17085,
    n17086, n17087, n17088, n17089, n17090, n17091,
    n17092, n17093, n17094, n17095, n17096, n17097,
    n17098, n17099, n17100, n17101, n17102, n17103,
    n17104, n17105, n17106, n17107, n17108, n17109,
    n17110, n17111, n17112, n17113, n17114, n17115,
    n17116, n17117, n17118, n17119, n17120, n17121,
    n17122, n17123, n17124, n17125, n17126, n17127,
    n17128, n17129, n17130, n17131, n17132, n17133,
    n17134, n17135, n17136, n17137, n17138, n17139,
    n17140, n17141, n17142, n17143, n17144, n17145,
    n17146, n17147, n17148, n17149, n17150, n17151,
    n17152, n17153, n17154, n17155, n17156, n17157,
    n17158, n17159, n17160, n17161, n17162, n17163,
    n17164, n17165, n17166, n17167, n17168, n17169,
    n17170, n17171, n17172, n17173, n17174, n17175,
    n17176, n17177, n17178, n17179, n17180, n17181,
    n17182, n17183, n17184, n17185, n17186, n17187,
    n17188, n17189, n17190, n17191, n17192, n17193,
    n17194, n17195, n17196, n17197, n17198, n17199,
    n17200, n17201, n17202, n17203, n17204, n17205,
    n17206, n17207, n17208, n17209, n17210, n17211,
    n17212, n17213, n17214, n17215, n17216, n17217,
    n17218, n17219, n17220, n17221, n17222, n17223,
    n17224, n17225, n17226, n17227, n17228, n17229,
    n17230, n17231, n17232, n17233, n17234, n17235,
    n17236, n17237, n17238, n17239, n17240, n17241,
    n17242, n17243, n17244, n17245, n17246, n17247,
    n17248, n17249, n17250, n17251, n17252, n17253,
    n17254, n17255, n17256, n17257, n17258, n17259,
    n17260, n17261, n17262, n17263, n17264, n17265,
    n17266, n17267, n17268, n17269, n17270, n17271,
    n17272, n17273, n17274, n17275, n17276, n17277,
    n17278, n17279, n17280, n17281, n17282, n17283,
    n17284, n17285, n17286, n17287, n17288, n17289,
    n17290, n17291, n17292, n17293, n17294, n17295,
    n17296, n17297, n17298, n17299, n17300, n17301,
    n17302, n17303, n17304, n17305, n17306, n17307,
    n17308, n17309, n17310, n17311, n17312, n17313,
    n17314, n17315, n17316, n17317, n17318, n17319,
    n17320, n17321, n17322, n17323, n17324, n17325,
    n17326, n17327, n17328, n17329, n17330, n17331,
    n17332, n17333, n17334, n17335, n17336, n17337,
    n17338, n17339, n17340, n17341, n17342, n17343,
    n17344, n17345, n17346, n17347, n17348, n17349,
    n17350, n17351, n17352, n17353, n17354, n17355,
    n17356, n17357, n17358, n17359, n17360, n17361,
    n17362, n17363, n17364, n17365, n17366, n17367,
    n17368, n17369, n17370, n17371, n17372, n17373,
    n17374, n17375, n17376, n17377, n17378, n17379,
    n17380, n17381, n17382, n17383, n17384, n17385,
    n17386, n17387, n17388, n17389, n17390, n17391,
    n17392, n17393, n17394, n17395, n17396, n17397,
    n17398, n17399, n17400, n17401, n17402, n17403,
    n17404, n17405, n17406, n17407, n17408, n17409,
    n17410, n17411, n17412, n17413, n17414, n17415,
    n17416, n17417, n17418, n17419, n17420, n17421,
    n17422, n17423, n17424, n17425, n17426, n17427,
    n17428, n17429, n17430, n17431, n17432, n17433,
    n17434, n17435, n17436, n17437, n17438, n17439,
    n17440, n17441, n17442, n17443, n17444, n17445,
    n17446, n17447, n17448, n17449, n17450, n17451,
    n17452, n17453, n17454, n17455, n17456, n17457,
    n17458, n17459, n17460, n17461, n17462, n17463,
    n17464, n17465, n17466, n17467, n17468, n17469,
    n17470, n17471, n17472, n17473, n17474, n17475,
    n17476, n17477, n17478, n17479, n17480, n17481,
    n17482, n17483, n17484, n17485, n17486, n17487,
    n17488, n17489, n17490, n17491, n17492, n17493,
    n17494, n17495, n17496, n17497, n17498, n17499,
    n17500, n17501, n17502, n17503, n17504, n17505,
    n17506, n17507, n17508, n17509, n17510, n17511,
    n17512, n17513, n17514, n17515, n17516, n17517,
    n17518, n17519, n17520, n17521, n17522, n17523,
    n17524, n17525, n17526, n17527, n17528, n17529,
    n17530, n17531, n17532, n17533, n17534, n17535,
    n17536, n17537, n17538, n17539, n17540, n17541,
    n17542, n17543, n17544, n17545, n17546, n17547,
    n17548, n17549, n17550, n17551, n17552, n17553,
    n17554, n17555, n17556, n17557, n17558, n17559,
    n17560, n17561, n17562, n17563, n17564, n17565,
    n17566, n17567, n17568, n17569, n17570, n17571,
    n17572, n17573, n17574, n17575, n17576, n17577,
    n17578, n17579, n17580, n17581, n17582, n17583,
    n17584, n17585, n17586, n17587, n17588, n17589,
    n17590, n17591, n17592, n17593, n17594, n17595,
    n17596, n17597, n17598, n17599, n17600, n17601,
    n17602, n17603, n17604, n17605, n17606, n17607,
    n17608, n17609, n17610, n17611, n17612, n17613,
    n17614, n17615, n17616, n17617, n17618, n17619,
    n17620, n17621, n17622, n17623, n17624, n17625,
    n17626, n17627, n17628, n17629, n17630, n17631,
    n17632, n17633, n17634, n17635, n17636, n17637,
    n17638, n17639, n17640, n17641, n17642, n17643,
    n17644, n17645, n17646, n17647, n17648, n17649,
    n17650, n17651, n17652, n17653, n17654, n17655,
    n17656, n17657, n17658, n17659, n17660, n17661,
    n17662, n17663, n17664, n17665, n17666, n17667,
    n17668, n17669, n17670, n17671, n17672, n17673,
    n17674, n17675, n17676, n17677, n17678, n17679,
    n17680, n17681, n17682, n17683, n17684, n17685,
    n17686, n17687, n17688, n17689, n17690, n17691,
    n17692, n17693, n17694, n17695, n17696, n17697,
    n17698, n17699, n17700, n17701, n17702, n17703,
    n17704, n17705, n17706, n17707, n17708, n17709,
    n17710, n17711, n17712, n17713, n17714, n17715,
    n17716, n17717, n17718, n17719, n17720, n17721,
    n17722, n17723, n17724, n17725, n17726, n17727,
    n17728, n17729, n17730, n17731, n17732, n17733,
    n17734, n17735, n17736, n17737, n17738, n17739,
    n17740, n17741, n17742, n17743, n17744, n17745,
    n17746, n17747, n17748, n17749, n17750, n17751,
    n17752, n17753, n17754, n17755, n17756, n17757,
    n17758, n17759, n17760, n17761, n17762, n17763,
    n17764, n17765, n17766, n17767, n17768, n17769,
    n17770, n17771, n17772, n17773, n17774, n17775,
    n17776, n17777, n17778, n17779, n17780, n17781,
    n17782, n17783, n17784, n17785, n17786, n17787,
    n17788, n17789, n17790, n17791, n17792, n17793,
    n17794, n17795, n17796, n17797, n17798, n17799,
    n17800, n17801, n17802, n17803, n17804, n17805,
    n17806, n17807, n17808, n17809, n17810, n17811,
    n17812, n17813, n17814, n17815, n17816, n17817,
    n17818, n17819, n17820, n17821, n17822, n17823,
    n17824, n17825, n17826, n17827, n17828, n17829,
    n17830, n17831, n17832, n17833, n17834, n17835,
    n17836, n17837, n17838, n17839, n17840, n17841,
    n17842, n17843, n17844, n17845, n17846, n17847,
    n17848, n17849, n17850, n17851, n17852, n17853,
    n17854, n17855, n17856, n17857, n17858, n17859,
    n17860, n17861, n17862, n17863, n17864, n17865,
    n17866, n17867, n17868, n17869, n17870, n17871,
    n17872, n17873, n17874, n17875, n17876, n17877,
    n17878, n17879, n17880, n17881, n17882, n17883,
    n17884, n17885, n17886, n17887, n17888, n17889,
    n17890, n17891, n17892, n17893, n17894, n17895,
    n17896, n17897, n17898, n17899, n17900, n17901,
    n17902, n17903, n17904, n17905, n17906, n17907,
    n17908, n17909, n17910, n17911, n17912, n17913,
    n17914, n17915, n17916, n17917, n17918, n17919,
    n17920, n17921, n17922, n17923, n17924, n17925,
    n17926, n17927, n17928, n17929, n17930, n17931,
    n17932, n17933, n17934, n17935, n17936, n17937,
    n17938, n17939, n17940, n17941, n17942, n17943,
    n17944, n17945, n17946, n17947, n17948, n17949,
    n17950, n17951, n17952, n17953, n17954, n17955,
    n17956, n17957, n17958, n17959, n17960, n17961,
    n17962, n17963, n17964, n17965, n17966, n17967,
    n17968, n17969, n17970, n17971, n17972, n17973,
    n17974, n17975, n17976, n17977, n17978, n17979,
    n17980, n17981, n17982, n17983, n17984, n17985,
    n17986, n17987, n17988, n17989, n17990, n17991,
    n17992, n17993, n17994, n17995, n17996, n17997,
    n17998, n17999, n18000, n18002, n18003, n18004,
    n18005, n18006, n18007, n18008, n18009, n18010,
    n18011, n18012, n18013, n18014, n18015, n18016,
    n18017, n18018, n18019, n18020, n18021, n18022,
    n18023, n18024, n18025, n18026, n18027, n18028,
    n18029, n18030, n18031, n18032, n18033, n18034,
    n18035, n18036, n18037, n18038, n18039, n18040,
    n18041, n18042, n18043, n18044, n18045, n18046,
    n18047, n18048, n18049, n18050, n18051, n18052,
    n18053, n18054, n18055, n18056, n18057, n18058,
    n18059, n18060, n18061, n18062, n18063, n18064,
    n18065, n18066, n18067, n18068, n18069, n18070,
    n18071, n18072, n18073, n18074, n18075, n18076,
    n18077, n18078, n18079, n18080, n18081, n18082,
    n18083, n18084, n18085, n18086, n18087, n18088,
    n18089, n18090, n18091, n18092, n18093, n18094,
    n18095, n18096, n18097, n18098, n18099, n18100,
    n18101, n18102, n18103, n18104, n18105, n18106,
    n18107, n18108, n18109, n18110, n18111, n18112,
    n18113, n18114, n18115, n18116, n18117, n18118,
    n18119, n18120, n18121, n18122, n18123, n18124,
    n18125, n18126, n18127, n18128, n18129, n18130,
    n18131, n18132, n18133, n18134, n18135, n18136,
    n18137, n18138, n18139, n18140, n18141, n18142,
    n18143, n18144, n18145, n18146, n18147, n18148,
    n18149, n18150, n18151, n18152, n18153, n18154,
    n18155, n18156, n18157, n18158, n18159, n18160,
    n18161, n18162, n18163, n18164, n18165, n18166,
    n18167, n18168, n18169, n18170, n18171, n18172,
    n18173, n18174, n18175, n18176, n18177, n18178,
    n18179, n18180, n18181, n18182, n18183, n18184,
    n18185, n18186, n18187, n18188, n18189, n18190,
    n18191, n18192, n18193, n18194, n18195, n18196,
    n18197, n18198, n18199, n18200, n18201, n18202,
    n18203, n18204, n18205, n18206, n18207, n18208,
    n18209, n18210, n18211, n18212, n18213, n18214,
    n18215, n18216, n18217, n18218, n18219, n18220,
    n18221, n18222, n18223, n18224, n18225, n18226,
    n18227, n18228, n18229, n18230, n18231, n18232,
    n18233, n18234, n18235, n18236, n18237, n18238,
    n18239, n18240, n18241, n18242, n18243, n18244,
    n18245, n18246, n18247, n18248, n18249, n18250,
    n18251, n18252, n18253, n18254, n18255, n18256,
    n18257, n18258, n18259, n18260, n18261, n18262,
    n18263, n18264, n18265, n18266, n18267, n18268,
    n18269, n18270, n18271, n18272, n18273, n18274,
    n18275, n18276, n18277, n18278, n18279, n18280,
    n18281, n18282, n18283, n18284, n18285, n18286,
    n18287, n18288, n18289, n18290, n18291, n18292,
    n18293, n18294, n18295, n18296, n18297, n18298,
    n18299, n18300, n18301, n18302, n18303, n18304,
    n18305, n18306, n18307, n18308, n18309, n18310,
    n18311, n18312, n18313, n18314, n18315, n18316,
    n18317, n18318, n18319, n18320, n18321, n18322,
    n18323, n18324, n18325, n18326, n18327, n18328,
    n18329, n18330, n18331, n18332, n18333, n18334,
    n18335, n18336, n18337, n18338, n18339, n18340,
    n18341, n18342, n18343, n18344, n18345, n18346,
    n18347, n18348, n18349, n18350, n18351, n18352,
    n18353, n18354, n18355, n18356, n18357, n18358,
    n18359, n18360, n18361, n18362, n18363, n18364,
    n18365, n18366, n18367, n18368, n18369, n18370,
    n18371, n18372, n18373, n18374, n18375, n18376,
    n18377, n18378, n18379, n18380, n18381, n18382,
    n18383, n18384, n18385, n18386, n18387, n18388,
    n18389, n18390, n18391, n18392, n18393, n18394,
    n18395, n18396, n18397, n18398, n18399, n18400,
    n18401, n18402, n18403, n18404, n18405, n18406,
    n18407, n18408, n18409, n18410, n18411, n18412,
    n18413, n18414, n18415, n18416, n18417, n18418,
    n18419, n18420, n18421, n18422, n18423, n18424,
    n18425, n18426, n18427, n18428, n18429, n18430,
    n18431, n18432, n18433, n18434, n18435, n18436,
    n18437, n18438, n18439, n18440, n18441, n18442,
    n18443, n18444, n18445, n18446, n18447, n18448,
    n18449, n18450, n18451, n18452, n18453, n18454,
    n18455, n18456, n18457, n18458, n18459, n18460,
    n18461, n18462, n18463, n18464, n18465, n18466,
    n18467, n18468, n18469, n18470, n18471, n18472,
    n18473, n18474, n18475, n18476, n18477, n18478,
    n18479, n18480, n18481, n18482, n18483, n18484,
    n18485, n18486, n18487, n18488, n18489, n18490,
    n18491, n18492, n18493, n18494, n18495, n18496,
    n18497, n18498, n18499, n18500, n18501, n18502,
    n18503, n18504, n18505, n18506, n18507, n18508,
    n18509, n18510, n18511, n18512, n18513, n18514,
    n18515, n18516, n18517, n18518, n18519, n18520,
    n18521, n18522, n18523, n18524, n18525, n18527,
    n18528, n18529, n18530, n18531, n18532, n18533,
    n18534, n18535, n18536, n18537, n18538, n18539,
    n18540, n18541, n18542, n18543, n18544, n18545,
    n18546, n18547, n18548, n18549, n18550, n18551,
    n18552, n18553, n18554, n18555, n18556, n18557,
    n18558, n18559, n18560, n18561, n18562, n18563,
    n18564, n18565, n18566, n18567, n18568, n18569,
    n18570, n18571, n18572, n18573, n18574, n18575,
    n18576, n18577, n18578, n18579, n18580, n18581,
    n18582, n18583, n18584, n18585, n18586, n18587,
    n18588, n18589, n18590, n18591, n18592, n18593,
    n18594, n18595, n18596, n18597, n18598, n18599,
    n18600, n18601, n18602, n18603, n18604, n18605,
    n18606, n18607, n18608, n18609, n18610, n18611,
    n18612, n18613, n18614, n18615, n18616, n18617,
    n18618, n18619, n18620, n18621, n18622, n18623,
    n18624, n18625, n18626, n18627, n18628, n18629,
    n18630, n18631, n18632, n18633, n18634, n18635,
    n18636, n18637, n18638, n18639, n18640, n18641,
    n18642, n18643, n18644, n18645, n18646, n18647,
    n18648, n18649, n18650, n18651, n18652, n18653,
    n18654, n18655, n18656, n18657, n18658, n18659,
    n18660, n18661, n18662, n18663, n18664, n18665,
    n18666, n18667, n18668, n18669, n18670, n18671,
    n18672, n18673, n18674, n18675, n18676, n18677,
    n18678, n18679, n18680, n18681, n18682, n18683,
    n18684, n18685, n18686, n18687, n18688, n18689,
    n18690, n18691, n18692, n18693, n18694, n18695,
    n18696, n18697, n18698, n18699, n18700, n18701,
    n18702, n18703, n18704, n18705, n18706, n18707,
    n18708, n18709, n18710, n18711, n18712, n18713,
    n18714, n18715, n18716, n18717, n18718, n18719,
    n18720, n18721, n18722, n18723, n18724, n18725,
    n18726, n18727, n18728, n18729, n18730, n18731,
    n18732, n18733, n18734, n18735, n18736, n18737,
    n18738, n18739, n18740, n18741, n18742, n18743,
    n18744, n18745, n18746, n18747, n18748, n18749,
    n18750, n18751, n18752, n18753, n18754, n18755,
    n18756, n18757, n18758, n18759, n18760, n18761,
    n18762, n18763, n18764, n18765, n18766, n18767,
    n18768, n18769, n18770, n18771, n18772, n18773,
    n18774, n18775, n18776, n18777, n18778, n18779,
    n18780, n18781, n18782, n18783, n18784, n18785,
    n18786, n18787, n18788, n18789, n18790, n18791,
    n18792, n18793, n18794, n18795, n18796, n18797,
    n18798, n18799, n18800, n18801, n18802, n18803,
    n18804, n18805, n18806, n18807, n18808, n18809,
    n18810, n18811, n18812, n18813, n18814, n18815,
    n18816, n18817, n18818, n18819, n18820, n18821,
    n18822, n18823, n18824, n18825, n18826, n18827,
    n18828, n18829, n18830, n18831, n18832, n18833,
    n18834, n18835, n18836, n18837, n18838, n18839,
    n18840, n18841, n18842, n18843, n18844, n18845,
    n18846, n18847, n18848, n18849, n18850, n18851,
    n18852, n18853, n18854, n18855, n18856, n18857,
    n18858, n18859, n18860, n18861, n18862, n18863,
    n18864, n18865, n18866, n18867, n18868, n18869,
    n18870, n18871, n18872, n18873, n18874, n18875,
    n18876, n18877, n18878, n18879, n18880, n18881,
    n18882, n18883, n18884, n18885, n18886, n18887,
    n18888, n18889, n18890, n18891, n18892, n18893,
    n18894, n18895, n18896, n18897, n18898, n18899,
    n18900, n18901, n18902, n18903, n18904, n18905,
    n18906, n18907, n18908, n18909, n18910, n18911,
    n18912, n18913, n18914, n18915, n18916, n18917,
    n18918, n18919, n18920, n18921, n18922, n18923,
    n18924, n18925, n18926, n18927, n18928, n18929,
    n18930, n18931, n18932, n18933, n18934, n18935,
    n18936, n18937, n18938, n18939, n18940, n18941,
    n18942, n18943, n18944, n18945, n18946, n18947,
    n18948, n18949, n18950, n18951, n18952, n18953,
    n18954, n18955, n18956, n18957, n18958, n18959,
    n18960, n18961, n18962, n18963, n18964, n18965,
    n18966, n18967, n18968, n18969, n18970, n18971,
    n18972, n18973, n18974, n18975, n18976, n18977,
    n18978, n18979, n18980, n18981, n18982, n18983,
    n18984, n18985, n18986, n18987, n18988, n18989,
    n18990, n18991, n18992, n18993, n18994, n18995,
    n18996, n18997, n18998, n18999, n19000, n19001,
    n19002, n19003, n19004, n19005, n19006, n19007,
    n19008, n19009, n19010, n19011, n19012, n19013,
    n19014, n19015, n19016, n19017, n19018, n19019,
    n19020, n19021, n19022, n19023, n19024, n19025,
    n19026, n19027, n19028, n19029, n19030, n19031,
    n19032, n19033, n19034, n19035, n19036, n19037,
    n19038, n19039, n19040, n19041, n19042, n19043,
    n19044, n19045, n19046, n19047, n19048, n19049,
    n19050, n19051, n19052, n19053, n19054, n19055,
    n19056, n19057, n19058, n19059, n19060, n19061,
    n19062, n19063, n19064, n19065, n19066, n19067,
    n19068, n19069, n19070, n19071, n19072, n19073,
    n19074, n19075, n19076, n19077, n19078, n19079,
    n19080, n19081, n19082, n19083, n19084, n19085,
    n19086, n19087, n19088, n19089, n19090, n19091,
    n19092, n19093, n19094, n19095, n19096, n19097,
    n19098, n19099, n19100, n19101, n19102, n19103,
    n19104, n19105, n19106, n19107, n19108, n19109,
    n19110, n19111, n19112, n19113, n19114, n19115,
    n19116, n19117, n19118, n19119, n19120, n19121,
    n19122, n19123, n19124, n19125, n19126, n19127,
    n19128, n19129, n19130, n19131, n19132, n19133,
    n19134, n19135, n19136, n19137, n19138, n19139,
    n19140, n19141, n19142, n19143, n19144, n19145,
    n19146, n19147, n19148, n19149, n19150, n19151,
    n19152, n19153, n19154, n19155, n19156, n19157,
    n19158, n19159, n19160, n19161, n19162, n19163,
    n19164, n19165, n19166, n19167, n19168, n19169,
    n19170, n19171, n19172, n19173, n19174, n19175,
    n19176, n19177, n19178, n19179, n19180, n19181,
    n19182, n19183, n19184, n19185, n19186, n19187,
    n19188, n19189, n19190, n19191, n19192, n19193,
    n19194, n19195, n19196, n19197, n19198, n19199,
    n19200, n19201, n19202, n19203, n19204, n19205,
    n19206, n19207, n19208, n19209, n19210, n19211,
    n19212, n19213, n19214, n19215, n19216, n19217,
    n19218, n19219, n19220, n19221, n19222, n19223,
    n19224, n19225, n19226, n19227, n19228, n19229,
    n19230, n19231, n19232, n19233, n19234, n19235,
    n19236, n19237, n19238, n19239, n19240, n19241,
    n19242, n19243, n19244, n19245, n19246, n19247,
    n19248, n19249, n19250, n19251, n19252, n19253,
    n19254, n19255, n19256, n19257, n19258, n19259,
    n19260, n19261, n19262, n19263, n19264, n19265,
    n19266, n19267, n19268, n19269, n19270, n19271,
    n19272, n19273, n19274, n19275, n19276, n19277,
    n19278, n19279, n19280, n19281, n19282, n19283,
    n19284, n19285, n19286, n19287, n19288, n19289,
    n19290, n19291, n19292, n19293, n19294, n19295,
    n19296, n19297, n19298, n19299, n19300, n19302,
    n19303, n19304, n19305, n19306, n19307, n19308,
    n19309, n19310, n19311, n19312, n19313, n19314,
    n19315, n19316, n19317, n19318, n19319, n19320,
    n19321, n19322, n19323, n19324, n19325, n19326,
    n19327, n19328, n19329, n19330, n19331, n19332,
    n19333, n19334, n19335, n19336, n19337, n19338,
    n19339, n19340, n19341, n19342, n19343, n19344,
    n19345, n19346, n19347, n19348, n19349, n19350,
    n19351, n19352, n19353, n19354, n19355, n19356,
    n19357, n19358, n19359, n19360, n19361, n19362,
    n19363, n19364, n19365, n19366, n19367, n19368,
    n19369, n19370, n19371, n19372, n19373, n19374,
    n19375, n19376, n19377, n19378, n19379, n19380,
    n19381, n19382, n19383, n19384, n19385, n19386,
    n19387, n19388, n19389, n19390, n19391, n19392,
    n19393, n19394, n19395, n19396, n19397, n19398,
    n19399, n19400, n19401, n19402, n19403, n19404,
    n19405, n19406, n19407, n19408, n19409, n19410,
    n19411, n19412, n19413, n19414, n19415, n19416,
    n19417, n19418, n19419, n19420, n19421, n19422,
    n19423, n19424, n19425, n19426, n19427, n19428,
    n19429, n19430, n19431, n19432, n19433, n19434,
    n19435, n19436, n19437, n19438, n19439, n19440,
    n19441, n19442, n19443, n19444, n19445, n19446,
    n19447, n19448, n19449, n19450, n19451, n19452,
    n19453, n19454, n19455, n19456, n19457, n19458,
    n19459, n19460, n19461, n19462, n19463, n19464,
    n19465, n19466, n19467, n19468, n19469, n19470,
    n19471, n19472, n19473, n19474, n19475, n19476,
    n19477, n19478, n19479, n19480, n19481, n19482,
    n19483, n19484, n19485, n19486, n19487, n19488,
    n19489, n19490, n19491, n19492, n19493, n19494,
    n19495, n19496, n19497, n19498, n19499, n19500,
    n19501, n19502, n19503, n19504, n19505, n19506,
    n19507, n19508, n19509, n19510, n19511, n19512,
    n19513, n19514, n19515, n19516, n19517, n19518,
    n19519, n19520, n19521, n19522, n19523, n19524,
    n19525, n19526, n19527, n19528, n19529, n19530,
    n19531, n19532, n19533, n19534, n19535, n19536,
    n19537, n19538, n19539, n19540, n19541, n19542,
    n19543, n19544, n19545, n19546, n19547, n19548,
    n19549, n19550, n19551, n19552, n19553, n19554,
    n19555, n19556, n19557, n19558, n19559, n19560,
    n19561, n19562, n19563, n19564, n19565, n19566,
    n19567, n19568, n19569, n19570, n19571, n19572,
    n19573, n19574, n19575, n19576, n19577, n19578,
    n19579, n19580, n19581, n19582, n19583, n19584,
    n19585, n19586, n19587, n19588, n19589, n19590,
    n19591, n19592, n19593, n19594, n19595, n19596,
    n19597, n19598, n19599, n19600, n19601, n19602,
    n19603, n19604, n19605, n19606, n19607, n19608,
    n19609, n19610, n19611, n19612, n19613, n19614,
    n19615, n19616, n19617, n19618, n19619, n19620,
    n19621, n19622, n19623, n19624, n19625, n19626,
    n19627, n19628, n19629, n19630, n19631, n19632,
    n19633, n19634, n19635, n19636, n19637, n19638,
    n19639, n19640, n19641, n19642, n19643, n19644,
    n19645, n19646, n19647, n19648, n19649, n19650,
    n19651, n19652, n19653, n19654, n19655, n19656,
    n19657, n19658, n19659, n19660, n19661, n19662,
    n19663, n19664, n19665, n19666, n19667, n19668,
    n19669, n19670, n19671, n19672, n19673, n19674,
    n19675, n19676, n19677, n19678, n19679, n19680,
    n19681, n19682, n19683, n19684, n19685, n19686,
    n19687, n19688, n19689, n19690, n19691, n19692,
    n19693, n19694, n19695, n19696, n19697, n19698,
    n19699, n19700, n19701, n19702, n19703, n19704,
    n19705, n19706, n19707, n19708, n19709, n19710,
    n19711, n19712, n19713, n19714, n19715, n19716,
    n19717, n19718, n19719, n19720, n19721, n19722,
    n19723, n19724, n19725, n19726, n19727, n19728,
    n19729, n19730, n19731, n19732, n19733, n19734,
    n19735, n19736, n19737, n19738, n19739, n19740,
    n19741, n19742, n19743, n19744, n19745, n19746,
    n19747, n19748, n19749, n19750, n19751, n19752,
    n19753, n19754, n19755, n19756, n19757, n19758,
    n19759, n19760, n19761, n19762, n19763, n19764,
    n19765, n19766, n19767, n19768, n19769, n19770,
    n19771, n19772, n19773, n19774, n19775, n19776,
    n19777, n19778, n19779, n19780, n19781, n19782,
    n19783, n19784, n19785, n19786, n19787, n19788,
    n19789, n19790, n19791, n19792, n19793, n19794,
    n19795, n19796, n19797, n19798, n19799, n19800,
    n19801, n19802, n19803, n19804, n19805, n19806,
    n19807, n19808, n19809, n19810, n19811, n19812,
    n19813, n19814, n19815, n19816, n19817, n19818,
    n19819, n19820, n19821, n19822, n19823, n19824,
    n19825, n19826, n19828, n19829, n19830, n19831,
    n19832, n19833, n19834, n19835, n19836, n19837,
    n19838, n19839, n19840, n19841, n19842, n19843,
    n19844, n19845, n19846, n19847, n19848, n19849,
    n19850, n19851, n19852, n19853, n19854, n19855,
    n19856, n19857, n19858, n19859, n19860, n19861,
    n19862, n19863, n19864, n19865, n19866, n19867,
    n19868, n19869, n19870, n19871, n19872, n19873,
    n19874, n19875, n19876, n19877, n19878, n19879,
    n19880, n19881, n19882, n19883, n19884, n19885,
    n19886, n19887, n19888, n19889, n19890, n19891,
    n19892, n19893, n19894, n19895, n19896, n19897,
    n19898, n19899, n19900, n19901, n19902, n19903,
    n19904, n19905, n19906, n19907, n19908, n19909,
    n19910, n19911, n19912, n19913, n19914, n19915,
    n19916, n19917, n19918, n19919, n19920, n19921,
    n19922, n19923, n19924, n19925, n19926, n19927,
    n19928, n19929, n19930, n19931, n19932, n19933,
    n19934, n19935, n19936, n19937, n19938, n19939,
    n19940, n19941, n19942, n19943, n19944, n19945,
    n19946, n19947, n19948, n19949, n19950, n19951,
    n19952, n19953, n19954, n19955, n19956, n19957,
    n19958, n19959, n19960, n19961, n19962, n19963,
    n19964, n19965, n19966, n19967, n19968, n19969,
    n19970, n19971, n19972, n19973, n19974, n19975,
    n19976, n19977, n19978, n19979, n19980, n19981,
    n19982, n19983, n19984, n19985, n19986, n19987,
    n19988, n19989, n19990, n19991, n19992, n19993,
    n19994, n19995, n19996, n19997, n19998, n19999,
    n20000, n20001, n20002, n20003, n20004, n20005,
    n20006, n20007, n20008, n20009, n20010, n20011,
    n20012, n20013, n20014, n20015, n20016, n20017,
    n20018, n20019, n20020, n20021, n20022, n20023,
    n20024, n20025, n20026, n20027, n20028, n20029,
    n20030, n20031, n20032, n20033, n20034, n20035,
    n20036, n20037, n20038, n20039, n20040, n20041,
    n20042, n20043, n20044, n20045, n20046, n20047,
    n20048, n20049, n20050, n20051, n20052, n20053,
    n20054, n20055, n20056, n20057, n20058, n20059,
    n20060, n20061, n20062, n20063, n20064, n20065,
    n20066, n20067, n20068, n20069, n20070, n20071,
    n20072, n20073, n20074, n20075, n20076, n20077,
    n20078, n20079, n20080, n20081, n20082, n20083,
    n20084, n20085, n20086, n20087, n20088, n20089,
    n20090, n20091, n20092, n20093, n20094, n20095,
    n20096, n20097, n20098, n20099, n20100, n20101,
    n20102, n20103, n20104, n20105, n20106, n20107,
    n20108, n20109, n20110, n20111, n20112, n20113,
    n20114, n20115, n20116, n20117, n20118, n20119,
    n20120, n20121, n20122, n20123, n20124, n20125,
    n20126, n20127, n20128, n20129, n20130, n20131,
    n20132, n20133, n20134, n20135, n20136, n20137,
    n20138, n20139, n20140, n20141, n20142, n20143,
    n20144, n20145, n20146, n20147, n20148, n20149,
    n20150, n20151, n20152, n20153, n20154, n20155,
    n20156, n20157, n20158, n20159, n20160, n20161,
    n20162, n20163, n20164, n20165, n20166, n20167,
    n20168, n20169, n20170, n20171, n20172, n20173,
    n20174, n20175, n20176, n20177, n20178, n20179,
    n20180, n20181, n20182, n20183, n20184, n20185,
    n20186, n20187, n20188, n20189, n20190, n20191,
    n20192, n20193, n20194, n20195, n20196, n20197,
    n20198, n20199, n20200, n20201, n20202, n20203,
    n20204, n20205, n20206, n20207, n20208, n20209,
    n20210, n20211, n20212, n20213, n20214, n20215,
    n20216, n20217, n20218, n20219, n20220, n20221,
    n20222, n20223, n20224, n20225, n20226, n20227,
    n20228, n20229, n20230, n20231, n20232, n20233,
    n20234, n20235, n20236, n20237, n20238, n20239,
    n20240, n20241, n20242, n20243, n20244, n20245,
    n20246, n20247, n20248, n20249, n20250, n20251,
    n20252, n20253, n20254, n20255, n20256, n20257,
    n20258, n20259, n20260, n20261, n20262, n20263,
    n20264, n20265, n20266, n20267, n20268, n20269,
    n20270, n20271, n20272, n20273, n20274, n20275,
    n20276, n20277, n20278, n20279, n20280, n20281,
    n20282, n20283, n20284, n20285, n20286, n20287,
    n20288, n20289, n20290, n20291, n20292, n20293,
    n20294, n20295, n20296, n20297, n20298, n20299,
    n20300, n20301, n20302, n20303, n20304, n20305,
    n20306, n20307, n20308, n20309, n20310, n20311,
    n20312, n20313, n20314, n20315, n20316, n20317,
    n20318, n20319, n20320, n20321, n20322, n20323,
    n20324, n20325, n20326, n20327, n20328, n20329,
    n20330, n20331, n20332, n20333, n20334, n20335,
    n20336, n20337, n20338, n20339, n20340, n20341,
    n20342, n20343, n20344, n20346, n20347, n20348,
    n20349, n20350, n20351, n20352, n20353, n20354,
    n20355, n20356, n20357, n20358, n20359, n20360,
    n20361, n20362, n20363, n20364, n20365, n20366,
    n20367, n20368, n20369, n20370, n20371, n20372,
    n20373, n20374, n20375, n20376, n20377, n20378,
    n20379, n20380, n20381, n20382, n20383, n20384,
    n20385, n20386, n20387, n20388, n20389, n20390,
    n20391, n20392, n20393, n20394, n20395, n20396,
    n20397, n20398, n20399, n20400, n20401, n20402,
    n20403, n20404, n20405, n20406, n20407, n20408,
    n20409, n20410, n20411, n20412, n20413, n20414,
    n20415, n20416, n20417, n20418, n20419, n20420,
    n20421, n20422, n20423, n20424, n20425, n20426,
    n20427, n20428, n20429, n20430, n20431, n20432,
    n20433, n20434, n20435, n20436, n20437, n20438,
    n20439, n20440, n20441, n20442, n20443, n20444,
    n20445, n20446, n20447, n20448, n20449, n20450,
    n20451, n20452, n20453, n20454, n20455, n20456,
    n20457, n20458, n20459, n20460, n20461, n20462,
    n20463, n20464, n20465, n20466, n20467, n20468,
    n20469, n20470, n20471, n20472, n20473, n20474,
    n20475, n20476, n20477, n20478, n20479, n20480,
    n20481, n20482, n20483, n20484, n20485, n20486,
    n20487, n20488, n20489, n20490, n20491, n20492,
    n20493, n20494, n20495, n20496, n20497, n20498,
    n20499, n20500, n20501, n20502, n20503, n20504,
    n20505, n20506, n20507, n20508, n20509, n20510,
    n20511, n20512, n20513, n20514, n20515, n20516,
    n20517, n20518, n20519, n20520, n20521, n20522,
    n20523, n20524, n20525, n20526, n20527, n20528,
    n20529, n20530, n20531, n20532, n20533, n20534,
    n20535, n20536, n20537, n20538, n20539, n20540,
    n20541, n20542, n20543, n20544, n20545, n20546,
    n20547, n20548, n20549, n20550, n20551, n20552,
    n20553, n20554, n20555, n20556, n20557, n20558,
    n20559, n20560, n20561, n20562, n20563, n20564,
    n20565, n20566, n20567, n20568, n20569, n20570,
    n20571, n20572, n20573, n20574, n20575, n20576,
    n20577, n20578, n20579, n20580, n20581, n20582,
    n20583, n20584, n20585, n20586, n20587, n20588,
    n20589, n20590, n20591, n20592, n20593, n20594,
    n20595, n20596, n20597, n20598, n20599, n20600,
    n20601, n20602, n20603, n20604, n20605, n20606,
    n20607, n20608, n20609, n20610, n20611, n20612,
    n20613, n20614, n20615, n20616, n20617, n20618,
    n20619, n20620, n20621, n20622, n20623, n20624,
    n20625, n20626, n20627, n20628, n20629, n20630,
    n20631, n20632, n20633, n20634, n20635, n20636,
    n20637, n20638, n20639, n20640, n20641, n20642,
    n20643, n20644, n20645, n20646, n20647, n20648,
    n20649, n20650, n20651, n20652, n20653, n20654,
    n20655, n20656, n20657, n20658, n20659, n20660,
    n20661, n20662, n20663, n20664, n20665, n20666,
    n20667, n20668, n20669, n20670, n20671, n20672,
    n20673, n20674, n20675, n20676, n20677, n20678,
    n20679, n20680, n20681, n20682, n20683, n20684,
    n20685, n20686, n20687, n20688, n20689, n20690,
    n20691, n20692, n20693, n20694, n20695, n20696,
    n20697, n20698, n20699, n20700, n20701, n20702,
    n20703, n20704, n20705, n20706, n20707, n20708,
    n20709, n20710, n20711, n20712, n20713, n20714,
    n20715, n20716, n20717, n20718, n20719, n20720,
    n20721, n20722, n20723, n20724, n20725, n20726,
    n20727, n20728, n20729, n20730, n20731, n20732,
    n20733, n20734, n20735, n20736, n20737, n20738,
    n20739, n20740, n20741, n20742, n20743, n20744,
    n20745, n20746, n20747, n20748, n20749, n20750,
    n20751, n20752, n20753, n20754, n20755, n20756,
    n20757, n20758, n20759, n20760, n20761, n20762,
    n20763, n20764, n20765, n20766, n20767, n20768,
    n20769, n20770, n20771, n20772, n20773, n20774,
    n20775, n20776, n20777, n20778, n20779, n20780,
    n20781, n20782, n20783, n20784, n20785, n20786,
    n20787, n20788, n20789, n20790, n20791, n20792,
    n20793, n20794, n20795, n20796, n20797, n20798,
    n20799, n20800, n20801, n20802, n20803, n20804,
    n20805, n20806, n20807, n20808, n20809, n20810,
    n20811, n20812, n20813, n20814, n20815, n20816,
    n20817, n20818, n20819, n20820, n20821, n20822,
    n20823, n20824, n20825, n20826, n20827, n20828,
    n20829, n20830, n20832, n20833, n20834, n20835,
    n20836, n20837, n20838, n20839, n20840, n20841,
    n20842, n20843, n20844, n20845, n20846, n20847,
    n20848, n20849, n20850, n20851, n20852, n20853,
    n20854, n20855, n20856, n20857, n20858, n20859,
    n20860, n20861, n20862, n20863, n20864, n20865,
    n20866, n20867, n20868, n20869, n20870, n20871,
    n20872, n20873, n20874, n20875, n20876, n20877,
    n20878, n20879, n20880, n20881, n20882, n20883,
    n20884, n20885, n20886, n20887, n20888, n20889,
    n20890, n20891, n20892, n20893, n20894, n20895,
    n20896, n20897, n20898, n20899, n20900, n20901,
    n20902, n20903, n20904, n20905, n20906, n20907,
    n20908, n20909, n20910, n20911, n20913, n20914,
    n20915, n20916, n20917, n20918, n20919, n20920,
    n20921, n20922, n20923, n20924, n20925, n20926,
    n20927, n20928, n20929, n20930, n20931, n20932,
    n20933, n20934, n20935, n20936, n20937, n20938,
    n20939, n20940, n20941, n20942, n20943, n20944,
    n20945, n20946, n20947, n20948, n20949, n20950,
    n20951, n20952, n20953, n20954, n20955, n20956,
    n20957, n20958, n20959, n20960, n20961, n20962,
    n20963, n20964, n20965, n20966, n20967, n20968,
    n20969, n20970, n20971, n20972, n20973, n20974,
    n20975, n20976, n20977, n20978, n20979, n20980,
    n20981, n20982, n20983, n20984, n20985, n20986,
    n20987, n20988, n20989, n20990, n20991, n20992,
    n20993, n20994, n20995, n20996, n20997, n20998,
    n20999, n21000, n21001, n21002, n21003, n21004,
    n21005, n21006, n21007, n21008, n21009, n21010,
    n21011, n21012, n21013, n21014, n21015, n21016,
    n21017, n21018, n21019, n21020, n21021, n21022,
    n21023, n21024, n21025, n21026, n21027, n21028,
    n21029, n21030, n21031, n21032, n21033, n21034,
    n21035, n21036, n21037, n21038, n21039, n21040,
    n21041, n21042, n21043, n21044, n21045, n21046,
    n21047, n21048, n21049, n21050, n21051, n21052,
    n21053, n21054, n21055, n21056, n21057, n21058,
    n21059, n21061, n21062, n21063, n21064, n21065,
    n21066, n21067, n21068, n21069, n21070, n21071,
    n21072, n21073, n21074, n21075, n21076, n21077,
    n21078, n21079, n21080, n21081, n21082, n21083,
    n21084, n21085, n21086, n21087, n21088, n21089,
    n21090, n21091, n21092, n21093, n21094, n21095,
    n21096, n21097, n21098, n21099, n21100, n21101,
    n21102, n21103, n21104, n21105, n21106, n21107,
    n21108, n21109, n21110, n21111, n21112, n21113,
    n21114, n21115, n21116, n21117, n21118, n21119,
    n21120, n21121, n21122, n21123, n21125, n21126,
    n21127, n21128, n21129, n21130, n21131, n21132,
    n21133, n21134, n21135, n21136, n21137, n21138,
    n21139, n21140, n21141, n21142, n21143, n21144,
    n21145, n21146, n21147, n21148, n21149, n21150,
    n21151, n21152, n21153, n21154, n21155, n21156,
    n21157, n21158, n21159, n21160, n21161, n21162,
    n21163, n21164, n21165, n21166, n21167, n21168,
    n21169, n21170, n21171, n21172, n21173, n21174,
    n21175, n21176, n21177, n21178, n21179, n21180,
    n21181, n21182, n21184, n21185, n21186, n21187,
    n21188, n21189, n21190, n21191, n21192, n21193,
    n21194, n21195, n21196, n21197, n21198, n21199,
    n21200, n21201, n21202, n21203, n21204, n21205,
    n21206, n21207, n21208, n21209, n21210, n21211,
    n21212, n21213, n21214, n21215, n21216, n21217,
    n21218, n21219, n21220, n21221, n21222, n21223,
    n21224, n21225, n21226, n21227, n21228, n21229,
    n21230, n21231, n21232, n21233, n21234, n21235,
    n21236, n21237, n21238, n21240, n21241, n21242,
    n21243, n21244, n21245, n21246, n21247, n21248,
    n21249, n21250, n21251, n21252, n21253, n21254,
    n21255, n21256, n21257, n21258, n21259, n21260,
    n21261, n21262, n21263, n21264, n21265, n21266,
    n21267, n21268, n21269, n21270, n21271, n21272,
    n21273, n21274, n21275, n21276, n21277, n21278,
    n21279, n21280, n21281, n21282, n21283, n21284,
    n21285, n21286, n21287, n21288, n21289, n21290,
    n21291, n21292, n21293, n21294, n21295, n21296,
    n21297, n21298, n21299, n21300, n21301, n21302,
    n21303, n21304, n21305, n21306, n21307, n21308,
    n21309, n21310, n21311, n21312, n21313, n21314,
    n21315, n21316, n21318, n21319, n21320, n21321,
    n21322, n21323, n21324, n21325, n21326, n21327,
    n21328, n21329, n21330, n21331, n21332, n21333,
    n21334, n21335, n21336, n21337, n21338, n21339,
    n21340, n21341, n21342, n21343, n21344, n21345,
    n21346, n21347, n21348, n21349, n21350, n21351,
    n21352, n21353, n21354, n21355, n21356, n21357,
    n21358, n21359, n21360, n21361, n21362, n21363,
    n21364, n21365, n21366, n21367, n21368, n21369,
    n21370, n21371, n21372, n21373, n21374, n21375,
    n21376, n21377, n21378, n21379, n21380, n21381,
    n21382, n21383, n21384, n21385, n21386, n21387,
    n21388, n21389, n21390, n21391, n21392, n21393,
    n21394, n21395, n21396, n21397, n21398, n21399,
    n21400, n21401, n21402, n21403, n21404, n21405,
    n21406, n21407, n21408, n21409, n21410, n21411,
    n21412, n21413, n21414, n21415, n21416, n21417,
    n21418, n21419, n21421, n21422, n21423, n21424,
    n21425, n21426, n21427, n21428, n21429, n21430,
    n21431, n21432, n21433, n21434, n21435, n21436,
    n21437, n21438, n21439, n21440, n21441, n21442,
    n21443, n21444, n21445, n21446, n21447, n21448,
    n21449, n21450, n21451, n21452, n21453, n21454,
    n21455, n21456, n21457, n21458, n21459, n21460,
    n21461, n21462, n21463, n21464, n21465, n21466,
    n21467, n21468, n21469, n21470, n21471, n21472,
    n21473, n21474, n21475, n21476, n21477, n21478,
    n21479, n21480, n21481, n21482, n21483, n21484,
    n21485, n21486, n21487, n21488, n21489, n21490,
    n21491, n21492, n21493, n21494, n21495, n21496,
    n21497, n21498, n21499, n21500, n21502, n21503,
    n21504, n21505, n21506, n21507, n21508, n21509,
    n21510, n21511, n21512, n21513, n21514, n21515,
    n21516, n21517, n21518, n21519, n21520, n21521,
    n21522, n21523, n21524, n21525, n21526, n21527,
    n21528, n21529, n21530, n21531, n21532, n21533,
    n21534, n21535, n21536, n21537, n21538, n21539,
    n21540, n21541, n21542, n21543, n21544, n21545,
    n21546, n21547, n21548, n21549, n21550, n21551,
    n21552, n21554, n21555, n21556, n21557, n21558,
    n21559, n21560, n21561, n21562, n21563, n21564,
    n21565, n21566, n21567, n21568, n21569, n21570,
    n21571, n21572, n21573, n21574, n21575, n21576,
    n21577, n21578, n21579, n21580, n21581, n21582,
    n21583, n21584, n21585, n21586, n21587, n21588,
    n21589, n21590, n21591, n21592, n21594, n21595,
    n21596, n21597, n21598, n21599, n21600, n21601,
    n21602, n21603, n21604, n21605, n21606, n21607,
    n21608, n21609, n21610, n21611, n21612, n21613,
    n21614, n21615, n21616, n21617, n21618, n21619,
    n21620, n21621, n21622, n21624, n21625, n21626,
    n21627, n21628, n21629, n21630, n21631, n21632,
    n21633, n21634, n21635, n21636, n21637, n21638,
    n21639, n21640, n21641, n21642, n21643, n21644,
    n21645, n21646, n21647, n21648, n21649, n21650,
    n21651, n21652, n21653, n21654, n21655, n21656,
    n21657, n21658, n21659, n21660, n21661, n21662,
    n21663, n21664, n21665, n21666, n21667, n21668,
    n21669, n21670, n21671, n21672, n21673, n21674,
    n21675, n21676, n21677, n21678, n21679, n21681,
    n21682, n21683, n21684, n21685, n21686, n21687,
    n21688, n21689, n21690, n21691, n21692, n21693,
    n21694, n21695, n21696, n21697, n21698, n21699,
    n21700, n21701, n21702, n21703, n21704, n21705,
    n21706, n21707, n21708, n21709, n21710, n21711,
    n21712, n21713, n21714, n21715, n21716, n21717,
    n21718, n21719, n21720, n21721, n21722, n21723,
    n21724, n21725, n21726, n21727, n21728, n21729,
    n21730, n21731, n21732, n21733, n21734, n21735,
    n21737, n21738, n21739, n21740, n21741, n21742,
    n21743, n21744, n21745, n21746, n21747, n21748,
    n21749, n21750, n21751, n21752, n21753, n21754,
    n21755, n21756, n21757, n21758, n21759, n21760,
    n21761, n21762, n21763, n21764, n21765, n21766,
    n21767, n21768, n21769, n21770, n21771, n21772,
    n21773, n21774, n21775, n21776, n21777, n21778,
    n21779, n21780, n21781, n21782, n21783, n21784,
    n21785, n21786, n21787, n21788, n21789, n21790,
    n21791, n21793, n21794, n21795, n21796, n21797,
    n21798, n21799, n21800, n21801, n21802, n21803,
    n21804, n21805, n21806, n21807, n21808, n21809,
    n21810, n21811, n21812, n21813, n21814, n21815,
    n21816, n21817, n21818, n21819, n21820, n21821,
    n21822, n21823, n21824, n21825, n21826, n21827,
    n21828, n21829, n21830, n21831, n21832, n21833,
    n21834, n21835, n21836, n21837, n21838, n21839,
    n21840, n21841, n21842, n21843, n21844, n21845,
    n21846, n21847, n21848, n21849, n21850, n21852,
    n21853, n21854, n21855, n21856, n21857, n21858,
    n21859, n21860, n21861, n21862, n21863, n21864,
    n21865, n21866, n21867, n21868, n21869, n21870,
    n21871, n21872, n21873, n21874, n21875, n21876,
    n21877, n21878, n21879, n21880, n21881, n21882,
    n21883, n21884, n21885, n21886, n21887, n21888,
    n21889, n21890, n21891, n21892, n21893, n21894,
    n21895, n21896, n21897, n21898, n21899, n21900,
    n21901, n21902, n21903, n21904, n21905, n21906,
    n21907, n21908, n21909, n21910, n21911, n21912,
    n21913, n21914, n21915, n21916, n21917, n21918,
    n21919, n21920, n21921, n21922, n21923, n21924,
    n21925, n21926, n21927, n21928, n21929, n21930,
    n21931, n21932, n21933, n21934, n21935, n21936,
    n21937, n21938, n21939, n21940, n21941, n21942,
    n21943, n21944, n21946, n21947, n21948, n21949,
    n21950, n21951, n21952, n21953, n21954, n21955,
    n21956, n21957, n21958, n21959, n21960, n21961,
    n21962, n21963, n21964, n21965, n21966, n21967,
    n21968, n21969, n21970, n21971, n21972, n21973,
    n21974, n21975, n21976, n21977, n21978, n21979,
    n21980, n21981, n21982, n21983, n21984, n21985,
    n21986, n21987, n21988, n21989, n21990, n21991,
    n21992, n21993, n21994, n21995, n21996, n21997,
    n21998, n21999, n22001, n22002, n22003, n22004,
    n22005, n22006, n22007, n22008, n22009, n22010,
    n22011, n22012, n22013, n22014, n22015, n22016,
    n22017, n22018, n22019, n22020, n22021, n22022,
    n22023, n22024, n22025, n22026, n22027, n22028,
    n22029, n22030, n22031, n22032, n22033, n22034,
    n22035, n22036, n22037, n22038, n22039, n22040,
    n22041, n22042, n22043, n22044, n22045, n22046,
    n22047, n22048, n22049, n22050, n22051, n22052,
    n22053, n22054, n22055, n22056, n22057, n22059,
    n22060, n22061, n22062, n22063, n22064, n22065,
    n22066, n22067, n22068, n22069, n22070, n22071,
    n22072, n22073, n22074, n22075, n22076, n22077,
    n22078, n22079, n22080, n22081, n22082, n22083,
    n22084, n22085, n22086, n22087, n22088, n22089,
    n22090, n22091, n22092, n22093, n22094, n22095,
    n22096, n22097, n22099, n22100, n22101, n22102,
    n22103, n22104, n22105, n22106, n22107, n22108,
    n22109, n22110, n22111, n22112, n22113, n22114,
    n22115, n22116, n22117, n22118, n22119, n22120,
    n22121, n22122, n22123, n22124, n22125, n22126,
    n22127, n22128, n22129, n22130, n22131, n22132,
    n22133, n22134, n22135, n22136, n22137, n22139,
    n22140, n22141, n22142, n22143, n22144, n22145,
    n22146, n22147, n22148, n22149, n22150, n22151,
    n22152, n22153, n22154, n22155, n22156, n22157,
    n22158, n22159, n22160, n22161, n22162, n22163,
    n22164, n22165, n22166, n22167, n22168, n22169,
    n22170, n22171, n22172, n22173, n22174, n22175,
    n22176, n22177, n22178, n22179, n22180, n22181,
    n22182, n22183, n22184, n22185, n22186, n22187,
    n22188, n22189, n22190, n22191, n22192, n22193,
    n22194, n22195, n22196, n22197, n22198, n22199,
    n22200, n22201, n22202, n22203, n22204, n22205,
    n22206, n22207, n22208, n22209, n22210, n22211,
    n22212, n22213, n22214, n22215, n22216, n22217,
    n22218, n22219, n22220, n22221, n22222, n22223,
    n22224, n22225, n22226, n22227, n22228, n22229,
    n22230, n22231, n22232, n22233, n22234, n22236,
    n22237, n22238, n22239, n22240, n22241, n22242,
    n22243, n22244, n22245, n22246, n22247, n22248,
    n22249, n22250, n22251, n22252, n22253, n22254,
    n22255, n22256, n22257, n22258, n22259, n22260,
    n22261, n22262, n22263, n22264, n22265, n22266,
    n22267, n22268, n22269, n22270, n22271, n22272,
    n22273, n22274, n22275, n22276, n22277, n22279,
    n22280, n22281, n22282, n22283, n22284, n22285,
    n22286, n22287, n22288, n22289, n22290, n22291,
    n22292, n22293, n22294, n22295, n22296, n22297,
    n22298, n22299, n22300, n22301, n22302, n22303,
    n22304, n22305, n22306, n22307, n22308, n22309,
    n22310, n22311, n22312, n22313, n22314, n22315,
    n22316, n22317, n22318, n22319, n22320, n22321,
    n22322, n22323, n22324, n22325, n22326, n22327,
    n22328, n22329, n22330, n22331, n22332, n22333,
    n22334, n22335, n22336, n22337, n22338, n22339,
    n22340, n22341, n22342, n22343, n22344, n22345,
    n22346, n22347, n22348, n22349, n22350, n22351,
    n22352, n22353, n22354, n22355, n22356, n22357,
    n22358, n22360, n22361, n22362, n22363, n22364,
    n22365, n22366, n22367, n22368, n22369, n22370,
    n22371, n22372, n22373, n22374, n22375, n22376,
    n22377, n22378, n22379, n22380, n22381, n22382,
    n22383, n22384, n22385, n22386, n22387, n22388,
    n22389, n22390, n22391, n22392, n22393, n22394,
    n22395, n22396, n22397, n22398, n22399, n22400,
    n22401, n22402, n22403, n22404, n22405, n22406,
    n22407, n22408, n22409, n22410, n22411, n22412,
    n22413, n22414, n22415, n22416, n22417, n22418,
    n22419, n22420, n22421, n22422, n22423, n22424,
    n22425, n22426, n22427, n22428, n22429, n22430,
    n22431, n22432, n22433, n22434, n22435, n22436,
    n22437, n22438, n22439, n22441, n22442, n22443,
    n22444, n22445, n22446, n22447, n22448, n22449,
    n22450, n22451, n22452, n22453, n22454, n22455,
    n22456, n22457, n22458, n22459, n22460, n22461,
    n22462, n22463, n22464, n22465, n22466, n22467,
    n22468, n22469, n22470, n22471, n22472, n22473,
    n22474, n22475, n22476, n22477, n22478, n22479,
    n22480, n22481, n22482, n22483, n22484, n22485,
    n22486, n22487, n22488, n22489, n22490, n22491,
    n22492, n22493, n22494, n22495, n22496, n22497,
    n22498, n22499, n22500, n22501, n22502, n22503,
    n22504, n22505, n22506, n22507, n22508, n22509,
    n22510, n22511, n22512, n22513, n22514, n22515,
    n22516, n22517, n22518, n22519, n22521, n22522,
    n22523, n22524, n22525, n22526, n22527, n22528,
    n22529, n22530, n22531, n22532, n22533, n22534,
    n22535, n22536, n22537, n22538, n22539, n22540,
    n22541, n22542, n22543, n22544, n22545, n22546,
    n22547, n22548, n22549, n22550, n22551, n22552,
    n22553, n22554, n22555, n22556, n22557, n22558,
    n22559, n22560, n22561, n22562, n22563, n22564,
    n22565, n22566, n22567, n22568, n22569, n22570,
    n22571, n22572, n22573, n22574, n22575, n22576,
    n22577, n22578, n22579, n22580, n22581, n22582,
    n22583, n22584, n22585, n22586, n22587, n22588,
    n22589, n22590, n22591, n22592, n22593, n22594,
    n22595, n22596, n22597, n22598, n22599, n22600,
    n22602, n22603, n22604, n22605, n22606, n22607,
    n22608, n22609, n22610, n22611, n22612, n22613,
    n22614, n22615, n22616, n22617, n22618, n22619,
    n22620, n22621, n22622, n22623, n22624, n22625,
    n22626, n22627, n22628, n22629, n22630, n22631,
    n22632, n22633, n22634, n22635, n22636, n22637,
    n22638, n22639, n22640, n22641, n22642, n22643,
    n22644, n22645, n22646, n22647, n22648, n22649,
    n22650, n22651, n22652, n22653, n22654, n22655,
    n22656, n22657, n22658, n22659, n22660, n22661,
    n22662, n22663, n22664, n22665, n22666, n22667,
    n22668, n22669, n22670, n22671, n22672, n22673,
    n22674, n22675, n22676, n22677, n22678, n22679,
    n22680, n22681, n22683, n22684, n22685, n22686,
    n22687, n22688, n22689, n22690, n22691, n22692,
    n22693, n22694, n22695, n22696, n22697, n22698,
    n22699, n22700, n22701, n22702, n22703, n22704,
    n22705, n22706, n22707, n22708, n22709, n22710,
    n22711, n22712, n22713, n22714, n22715, n22716,
    n22717, n22718, n22719, n22720, n22721, n22722,
    n22723, n22724, n22725, n22726, n22727, n22728,
    n22729, n22730, n22731, n22732, n22733, n22734,
    n22735, n22736, n22737, n22738, n22739, n22740,
    n22741, n22742, n22743, n22744, n22745, n22746,
    n22747, n22748, n22749, n22750, n22751, n22752,
    n22753, n22754, n22755, n22756, n22757, n22758,
    n22759, n22760, n22761, n22762, n22763, n22764,
    n22765, n22766, n22767, n22768, n22769, n22770,
    n22771, n22772, n22773, n22774, n22775, n22776,
    n22777, n22778, n22779, n22780, n22781, n22782,
    n22783, n22784, n22785, n22786, n22787, n22788,
    n22789, n22790, n22791, n22792, n22793, n22794,
    n22795, n22796, n22797, n22798, n22799, n22800,
    n22801, n22802, n22803, n22804, n22805, n22806,
    n22807, n22808, n22809, n22810, n22811, n22812,
    n22813, n22814, n22815, n22816, n22817, n22818,
    n22819, n22820, n22821, n22822, n22823, n22824,
    n22825, n22826, n22827, n22828, n22829, n22830,
    n22831, n22832, n22833, n22834, n22835, n22836,
    n22837, n22838, n22839, n22840, n22841, n22842,
    n22843, n22844, n22845, n22846, n22847, n22848,
    n22849, n22850, n22851, n22852, n22853, n22854,
    n22855, n22856, n22857, n22858, n22859, n22860,
    n22861, n22862, n22863, n22864, n22865, n22866,
    n22867, n22868, n22869, n22870, n22871, n22872,
    n22873, n22874, n22875, n22876, n22877, n22878,
    n22879, n22880, n22881, n22882, n22883, n22884,
    n22885, n22886, n22887, n22888, n22889, n22890,
    n22891, n22892, n22893, n22894, n22895, n22896,
    n22897, n22898, n22899, n22900, n22901, n22902,
    n22903, n22904, n22905, n22906, n22907, n22908,
    n22909, n22910, n22911, n22912, n22913, n22914,
    n22915, n22916, n22917, n22918, n22919, n22920,
    n22921, n22922, n22923, n22924, n22925, n22926,
    n22927, n22928, n22929, n22930, n22931, n22932,
    n22933, n22934, n22935, n22936, n22937, n22938,
    n22939, n22940, n22941, n22942, n22943, n22944,
    n22945, n22946, n22947, n22948, n22949, n22950,
    n22951, n22952, n22953, n22954, n22955, n22956,
    n22957, n22958, n22959, n22960, n22961, n22962,
    n22963, n22964, n22965, n22966, n22967, n22968,
    n22969, n22970, n22971, n22972, n22973, n22974,
    n22975, n22976, n22977, n22978, n22979, n22980,
    n22981, n22982, n22983, n22984, n22985, n22986,
    n22987, n22988, n22989, n22990, n22991, n22992,
    n22993, n22994, n22995, n22996, n22997, n22998,
    n22999, n23000, n23001, n23002, n23003, n23004,
    n23005, n23006, n23007, n23008, n23009, n23010,
    n23011, n23012, n23013, n23014, n23015, n23016,
    n23017, n23018, n23019, n23020, n23021, n23022,
    n23023, n23024, n23025, n23026, n23027, n23028,
    n23029, n23030, n23031, n23032, n23033, n23034,
    n23035, n23036, n23037, n23038, n23039, n23040,
    n23041, n23042, n23043, n23044, n23045, n23046,
    n23047, n23048, n23049, n23050, n23051, n23052,
    n23053, n23054, n23055, n23056, n23057, n23058,
    n23059, n23060, n23061, n23062, n23063, n23064,
    n23065, n23066, n23067, n23068, n23069, n23070,
    n23071, n23072, n23073, n23074, n23075, n23076,
    n23077, n23078, n23079, n23080, n23081, n23082,
    n23083, n23084, n23085, n23086, n23087, n23088,
    n23089, n23090, n23091, n23092, n23093, n23094,
    n23095, n23096, n23097, n23098, n23099, n23100,
    n23101, n23102, n23103, n23104, n23105, n23106,
    n23107, n23108, n23109, n23110, n23111, n23112,
    n23113, n23114, n23115, n23116, n23117, n23118,
    n23119, n23120, n23121, n23122, n23123, n23124,
    n23125, n23126, n23127, n23128, n23129, n23130,
    n23131, n23132, n23133, n23134, n23135, n23136,
    n23137, n23138, n23139, n23140, n23141, n23142,
    n23143, n23144, n23145, n23146, n23147, n23148,
    n23149, n23150, n23151, n23152, n23153, n23154,
    n23156, n23157, n23158, n23159, n23160, n23161,
    n23162, n23163, n23164, n23165, n23166, n23167,
    n23168, n23169, n23170, n23171, n23172, n23173,
    n23174, n23175, n23176, n23177, n23178, n23179,
    n23180, n23181, n23182, n23183, n23184, n23185,
    n23186, n23187, n23188, n23189, n23190, n23191,
    n23192, n23193, n23194, n23195, n23196, n23197,
    n23198, n23199, n23200, n23201, n23202, n23203,
    n23204, n23205, n23206, n23207, n23208, n23209,
    n23210, n23211, n23212, n23213, n23214, n23215,
    n23216, n23217, n23218, n23219, n23220, n23221,
    n23222, n23223, n23224, n23225, n23226, n23227,
    n23228, n23229, n23230, n23231, n23232, n23233,
    n23234, n23235, n23236, n23237, n23238, n23239,
    n23240, n23241, n23242, n23243, n23244, n23245,
    n23246, n23247, n23248, n23249, n23250, n23251,
    n23252, n23253, n23254, n23255, n23256, n23257,
    n23258, n23259, n23260, n23261, n23262, n23263,
    n23264, n23265, n23266, n23267, n23268, n23269,
    n23270, n23271, n23272, n23273, n23274, n23275,
    n23276, n23277, n23278, n23279, n23280, n23281,
    n23282, n23283, n23284, n23285, n23286, n23287,
    n23288, n23289, n23290, n23291, n23292, n23293,
    n23294, n23295, n23296, n23297, n23298, n23299,
    n23300, n23301, n23302, n23303, n23304, n23305,
    n23306, n23307, n23308, n23309, n23310, n23311,
    n23312, n23313, n23314, n23315, n23316, n23317,
    n23318, n23319, n23320, n23321, n23322, n23323,
    n23324, n23325, n23326, n23327, n23328, n23329,
    n23330, n23331, n23332, n23333, n23334, n23335,
    n23336, n23337, n23338, n23339, n23340, n23341,
    n23342, n23343, n23344, n23345, n23346, n23347,
    n23348, n23349, n23350, n23351, n23352, n23353,
    n23354, n23355, n23356, n23357, n23358, n23359,
    n23360, n23361, n23362, n23363, n23364, n23365,
    n23366, n23367, n23368, n23369, n23370, n23371,
    n23372, n23373, n23374, n23375, n23376, n23377,
    n23378, n23379, n23380, n23381, n23382, n23383,
    n23384, n23385, n23386, n23387, n23388, n23389,
    n23390, n23391, n23392, n23393, n23394, n23395,
    n23396, n23397, n23398, n23399, n23400, n23401,
    n23402, n23403, n23404, n23405, n23406, n23407,
    n23408, n23409, n23410, n23411, n23412, n23413,
    n23414, n23415, n23416, n23417, n23418, n23419,
    n23420, n23421, n23422, n23423, n23424, n23425,
    n23426, n23427, n23428, n23429, n23430, n23431,
    n23432, n23433, n23434, n23435, n23436, n23437,
    n23438, n23439, n23440, n23441, n23442, n23443,
    n23444, n23445, n23446, n23447, n23448, n23449,
    n23450, n23451, n23452, n23453, n23454, n23455,
    n23456, n23457, n23458, n23459, n23460, n23461,
    n23462, n23463, n23464, n23465, n23466, n23467,
    n23468, n23469, n23470, n23471, n23472, n23473,
    n23474, n23475, n23476, n23477, n23478, n23479,
    n23480, n23481, n23482, n23483, n23484, n23485,
    n23486, n23487, n23488, n23489, n23490, n23491,
    n23492, n23493, n23494, n23495, n23496, n23497,
    n23498, n23499, n23500, n23501, n23502, n23503,
    n23504, n23505, n23506, n23507, n23508, n23509,
    n23510, n23511, n23512, n23513, n23514, n23515,
    n23516, n23517, n23518, n23519, n23520, n23521,
    n23522, n23523, n23524, n23525, n23526, n23527,
    n23528, n23529, n23530, n23531, n23532, n23533,
    n23534, n23535, n23536, n23537, n23538, n23539,
    n23540, n23541, n23542, n23543, n23544, n23545,
    n23546, n23547, n23548, n23549, n23550, n23551,
    n23552, n23553, n23554, n23555, n23556, n23557,
    n23558, n23559, n23560, n23561, n23562, n23563,
    n23564, n23565, n23566, n23567, n23568, n23569,
    n23570, n23571, n23572, n23573, n23574, n23575,
    n23576, n23577, n23578, n23579, n23580, n23581,
    n23582, n23583, n23584, n23585, n23586, n23587,
    n23588, n23589, n23590, n23591, n23592, n23593,
    n23594, n23595, n23596, n23597, n23598, n23599,
    n23600, n23601, n23602, n23603, n23604, n23605,
    n23606, n23607, n23608, n23609, n23610, n23611,
    n23612, n23613, n23614, n23615, n23616, n23617,
    n23618, n23619, n23620, n23621, n23622, n23623,
    n23624, n23625, n23626, n23627, n23628, n23629,
    n23630, n23631, n23632, n23633, n23634, n23635,
    n23636, n23637, n23638, n23640, n23641, n23642,
    n23643, n23644, n23645, n23646, n23647, n23648,
    n23649, n23650, n23651, n23652, n23653, n23654,
    n23655, n23656, n23657, n23658, n23659, n23660,
    n23661, n23662, n23663, n23664, n23665, n23666,
    n23667, n23668, n23669, n23670, n23671, n23672,
    n23673, n23674, n23675, n23676, n23677, n23678,
    n23679, n23680, n23681, n23682, n23683, n23684,
    n23685, n23686, n23687, n23688, n23689, n23690,
    n23691, n23692, n23693, n23694, n23695, n23696,
    n23697, n23698, n23699, n23700, n23701, n23702,
    n23703, n23704, n23705, n23706, n23707, n23708,
    n23709, n23710, n23711, n23712, n23713, n23714,
    n23715, n23716, n23717, n23718, n23719, n23720,
    n23721, n23722, n23723, n23724, n23725, n23726,
    n23727, n23728, n23729, n23730, n23731, n23732,
    n23733, n23734, n23735, n23736, n23737, n23738,
    n23739, n23740, n23741, n23742, n23743, n23744,
    n23745, n23746, n23747, n23748, n23749, n23750,
    n23751, n23752, n23753, n23754, n23755, n23756,
    n23757, n23758, n23759, n23760, n23761, n23762,
    n23763, n23764, n23765, n23766, n23767, n23768,
    n23769, n23770, n23771, n23772, n23773, n23774,
    n23775, n23776, n23777, n23778, n23779, n23780,
    n23781, n23782, n23783, n23784, n23785, n23786,
    n23787, n23788, n23789, n23790, n23791, n23792,
    n23793, n23794, n23795, n23796, n23797, n23798,
    n23799, n23800, n23801, n23802, n23803, n23804,
    n23805, n23806, n23807, n23808, n23809, n23810,
    n23811, n23812, n23813, n23814, n23815, n23816,
    n23817, n23818, n23819, n23820, n23821, n23822,
    n23823, n23824, n23825, n23826, n23827, n23828,
    n23829, n23830, n23831, n23832, n23833, n23834,
    n23835, n23836, n23837, n23838, n23839, n23840,
    n23841, n23842, n23843, n23844, n23845, n23846,
    n23847, n23848, n23849, n23850, n23851, n23852,
    n23853, n23854, n23855, n23856, n23857, n23858,
    n23859, n23860, n23861, n23862, n23863, n23864,
    n23865, n23866, n23867, n23868, n23869, n23870,
    n23871, n23872, n23873, n23874, n23875, n23876,
    n23877, n23878, n23879, n23880, n23881, n23882,
    n23883, n23884, n23885, n23886, n23887, n23888,
    n23889, n23890, n23891, n23892, n23893, n23894,
    n23895, n23896, n23897, n23898, n23899, n23900,
    n23901, n23902, n23903, n23904, n23905, n23906,
    n23907, n23908, n23909, n23910, n23911, n23912,
    n23913, n23914, n23915, n23916, n23917, n23918,
    n23919, n23920, n23921, n23922, n23923, n23924,
    n23925, n23926, n23927, n23928, n23929, n23930,
    n23931, n23932, n23933, n23934, n23935, n23936,
    n23937, n23938, n23939, n23940, n23941, n23942,
    n23943, n23944, n23945, n23946, n23947, n23948,
    n23949, n23950, n23951, n23952, n23953, n23954,
    n23955, n23956, n23957, n23958, n23959, n23960,
    n23961, n23962, n23963, n23964, n23965, n23966,
    n23967, n23968, n23969, n23970, n23971, n23972,
    n23973, n23974, n23975, n23976, n23977, n23978,
    n23979, n23980, n23981, n23982, n23983, n23984,
    n23985, n23986, n23987, n23988, n23989, n23990,
    n23991, n23992, n23993, n23994, n23995, n23996,
    n23997, n23998, n23999, n24000, n24001, n24002,
    n24003, n24004, n24005, n24006, n24007, n24008,
    n24009, n24010, n24011, n24012, n24013, n24014,
    n24015, n24016, n24017, n24018, n24019, n24020,
    n24021, n24022, n24023, n24024, n24025, n24026,
    n24027, n24028, n24029, n24030, n24031, n24032,
    n24033, n24034, n24035, n24036, n24037, n24038,
    n24039, n24040, n24041, n24042, n24043, n24044,
    n24045, n24046, n24047, n24048, n24049, n24050,
    n24051, n24052, n24053, n24054, n24055, n24056,
    n24057, n24058, n24059, n24060, n24061, n24062,
    n24063, n24064, n24065, n24066, n24067, n24068,
    n24069, n24070, n24071, n24072, n24073, n24074,
    n24075, n24076, n24077, n24078, n24079, n24080,
    n24081, n24082, n24083, n24084, n24085, n24086,
    n24087, n24088, n24089, n24090, n24091, n24092,
    n24093, n24094, n24095, n24096, n24097, n24098,
    n24099, n24100, n24101, n24102, n24103, n24104,
    n24105, n24106, n24107, n24108, n24109, n24110,
    n24111, n24112, n24113, n24114, n24116, n24117,
    n24118, n24119, n24120, n24121, n24122, n24123,
    n24124, n24125, n24126, n24127, n24128, n24129,
    n24130, n24131, n24132, n24133, n24134, n24135,
    n24136, n24137, n24138, n24139, n24140, n24141,
    n24142, n24143, n24144, n24145, n24146, n24147,
    n24148, n24149, n24150, n24151, n24152, n24153,
    n24154, n24155, n24156, n24157, n24158, n24159,
    n24160, n24161, n24162, n24163, n24164, n24165,
    n24166, n24167, n24168, n24169, n24170, n24171,
    n24172, n24173, n24174, n24175, n24176, n24177,
    n24178, n24179, n24180, n24181, n24182, n24183,
    n24184, n24185, n24186, n24187, n24188, n24189,
    n24190, n24191, n24192, n24193, n24194, n24195,
    n24196, n24197, n24198, n24199, n24200, n24201,
    n24202, n24203, n24204, n24205, n24206, n24207,
    n24208, n24209, n24210, n24211, n24212, n24213,
    n24214, n24215, n24216, n24217, n24218, n24219,
    n24220, n24221, n24222, n24223, n24224, n24225,
    n24226, n24227, n24228, n24229, n24230, n24231,
    n24232, n24233, n24234, n24235, n24236, n24237,
    n24238, n24239, n24240, n24241, n24242, n24243,
    n24244, n24245, n24246, n24247, n24248, n24249,
    n24250, n24251, n24252, n24253, n24254, n24255,
    n24256, n24257, n24258, n24259, n24260, n24261,
    n24262, n24263, n24264, n24265, n24266, n24267,
    n24268, n24269, n24270, n24271, n24272, n24273,
    n24274, n24275, n24276, n24277, n24278, n24279,
    n24280, n24281, n24282, n24283, n24284, n24285,
    n24286, n24287, n24288, n24289, n24290, n24291,
    n24292, n24293, n24294, n24295, n24296, n24297,
    n24298, n24299, n24300, n24301, n24302, n24303,
    n24304, n24305, n24306, n24307, n24308, n24309,
    n24310, n24311, n24312, n24313, n24314, n24315,
    n24316, n24317, n24318, n24319, n24320, n24321,
    n24322, n24323, n24324, n24325, n24326, n24327,
    n24328, n24329, n24330, n24331, n24332, n24333,
    n24334, n24335, n24336, n24337, n24338, n24339,
    n24340, n24341, n24342, n24343, n24344, n24345,
    n24346, n24347, n24348, n24349, n24350, n24351,
    n24352, n24353, n24354, n24355, n24356, n24357,
    n24358, n24359, n24360, n24361, n24362, n24363,
    n24364, n24365, n24366, n24367, n24368, n24369,
    n24370, n24371, n24372, n24373, n24374, n24375,
    n24376, n24377, n24378, n24379, n24380, n24381,
    n24382, n24383, n24384, n24385, n24386, n24387,
    n24388, n24389, n24390, n24391, n24392, n24393,
    n24394, n24395, n24396, n24397, n24398, n24399,
    n24400, n24401, n24402, n24403, n24404, n24405,
    n24406, n24407, n24408, n24409, n24410, n24411,
    n24412, n24413, n24414, n24415, n24416, n24417,
    n24418, n24419, n24420, n24421, n24422, n24423,
    n24424, n24425, n24426, n24427, n24428, n24429,
    n24430, n24431, n24432, n24433, n24434, n24435,
    n24436, n24437, n24438, n24439, n24440, n24441,
    n24442, n24443, n24444, n24445, n24446, n24447,
    n24448, n24449, n24450, n24451, n24452, n24453,
    n24454, n24455, n24456, n24457, n24458, n24459,
    n24460, n24461, n24462, n24463, n24464, n24465,
    n24466, n24467, n24468, n24469, n24470, n24471,
    n24472, n24473, n24474, n24475, n24476, n24477,
    n24478, n24479, n24480, n24481, n24482, n24483,
    n24484, n24485, n24486, n24487, n24488, n24489,
    n24490, n24491, n24492, n24493, n24494, n24495,
    n24496, n24497, n24498, n24499, n24500, n24501,
    n24502, n24503, n24504, n24505, n24506, n24507,
    n24508, n24509, n24510, n24511, n24512, n24513,
    n24514, n24515, n24516, n24517, n24518, n24519,
    n24520, n24521, n24522, n24523, n24524, n24525,
    n24526, n24527, n24528, n24529, n24530, n24531,
    n24532, n24533, n24534, n24535, n24536, n24537,
    n24538, n24539, n24540, n24541, n24542, n24543,
    n24544, n24545, n24546, n24547, n24548, n24549,
    n24550, n24551, n24552, n24553, n24554, n24555,
    n24556, n24557, n24558, n24559, n24560, n24561,
    n24562, n24564, n24565, n24566, n24567, n24568,
    n24569, n24570, n24571, n24572, n24573, n24574,
    n24575, n24576, n24577, n24578, n24579, n24580,
    n24581, n24582, n24583, n24584, n24585, n24586,
    n24587, n24588, n24589, n24590, n24591, n24592,
    n24593, n24594, n24595, n24596, n24597, n24598,
    n24599, n24600, n24601, n24602, n24603, n24604,
    n24605, n24606, n24607, n24608, n24609, n24610,
    n24611, n24612, n24613, n24614, n24615, n24616,
    n24617, n24618, n24619, n24620, n24621, n24622,
    n24623, n24624, n24625, n24626, n24627, n24628,
    n24629, n24630, n24631, n24632, n24633, n24634,
    n24635, n24636, n24637, n24638, n24639, n24640,
    n24641, n24642, n24643, n24644, n24645, n24646,
    n24647, n24648, n24649, n24650, n24651, n24652,
    n24653, n24654, n24655, n24656, n24657, n24658,
    n24659, n24660, n24661, n24662, n24663, n24664,
    n24665, n24666, n24667, n24668, n24669, n24670,
    n24671, n24672, n24673, n24674, n24675, n24676,
    n24677, n24678, n24679, n24680, n24681, n24682,
    n24683, n24684, n24685, n24686, n24687, n24688,
    n24689, n24690, n24691, n24692, n24693, n24694,
    n24695, n24696, n24697, n24698, n24699, n24700,
    n24701, n24702, n24703, n24704, n24705, n24706,
    n24707, n24708, n24709, n24710, n24711, n24712,
    n24713, n24714, n24715, n24716, n24717, n24718,
    n24719, n24720, n24721, n24722, n24723, n24724,
    n24725, n24726, n24727, n24728, n24729, n24730,
    n24731, n24732, n24733, n24734, n24735, n24736,
    n24737, n24738, n24739, n24740, n24741, n24742,
    n24743, n24744, n24745, n24746, n24747, n24748,
    n24749, n24750, n24751, n24752, n24753, n24754,
    n24755, n24756, n24757, n24758, n24759, n24760,
    n24761, n24762, n24763, n24764, n24765, n24766,
    n24767, n24768, n24769, n24770, n24771, n24772,
    n24773, n24774, n24775, n24776, n24777, n24778,
    n24779, n24780, n24781, n24782, n24783, n24784,
    n24785, n24786, n24787, n24788, n24789, n24790,
    n24791, n24792, n24793, n24794, n24795, n24796,
    n24797, n24798, n24799, n24800, n24801, n24802,
    n24803, n24804, n24805, n24806, n24807, n24808,
    n24809, n24810, n24811, n24812, n24813, n24814,
    n24815, n24816, n24817, n24818, n24819, n24820,
    n24821, n24822, n24823, n24824, n24825, n24826,
    n24827, n24828, n24829, n24830, n24831, n24832,
    n24833, n24834, n24835, n24836, n24837, n24838,
    n24839, n24840, n24841, n24842, n24843, n24844,
    n24845, n24846, n24847, n24848, n24849, n24850,
    n24851, n24852, n24853, n24854, n24855, n24856,
    n24857, n24858, n24859, n24860, n24861, n24862,
    n24863, n24864, n24865, n24866, n24867, n24868,
    n24869, n24870, n24871, n24872, n24873, n24874,
    n24875, n24876, n24877, n24878, n24879, n24880,
    n24881, n24882, n24883, n24884, n24885, n24886,
    n24887, n24888, n24889, n24890, n24891, n24892,
    n24893, n24894, n24895, n24896, n24897, n24898,
    n24899, n24900, n24901, n24902, n24903, n24904,
    n24905, n24906, n24907, n24908, n24909, n24910,
    n24911, n24912, n24913, n24914, n24915, n24916,
    n24917, n24918, n24919, n24920, n24921, n24922,
    n24923, n24924, n24925, n24926, n24927, n24928,
    n24929, n24930, n24931, n24932, n24933, n24934,
    n24935, n24936, n24937, n24938, n24939, n24940,
    n24941, n24942, n24943, n24944, n24945, n24946,
    n24947, n24948, n24949, n24950, n24951, n24952,
    n24953, n24954, n24955, n24956, n24957, n24958,
    n24959, n24960, n24961, n24962, n24963, n24964,
    n24965, n24966, n24967, n24968, n24969, n24970,
    n24971, n24972, n24973, n24974, n24975, n24976,
    n24977, n24978, n24979, n24980, n24981, n24982,
    n24983, n24984, n24985, n24986, n24987, n24988,
    n24989, n24990, n24991, n24992, n24993, n24994,
    n24995, n24996, n24997, n24998, n24999, n25000,
    n25001, n25002, n25003, n25004, n25005, n25006,
    n25007, n25008, n25009, n25010, n25011, n25012,
    n25013, n25014, n25015, n25016, n25017, n25018,
    n25019, n25020, n25021, n25022, n25023, n25024,
    n25025, n25026, n25027, n25028, n25029, n25030,
    n25031, n25032, n25033, n25034, n25035, n25036,
    n25037, n25038, n25039, n25040, n25041, n25042,
    n25043, n25044, n25046, n25047, n25048, n25049,
    n25050, n25051, n25052, n25053, n25054, n25055,
    n25056, n25057, n25058, n25059, n25060, n25061,
    n25062, n25063, n25064, n25065, n25066, n25067,
    n25068, n25069, n25070, n25071, n25072, n25073,
    n25074, n25075, n25076, n25077, n25078, n25079,
    n25080, n25081, n25082, n25083, n25084, n25085,
    n25086, n25087, n25088, n25089, n25090, n25091,
    n25092, n25093, n25094, n25095, n25096, n25097,
    n25098, n25099, n25100, n25101, n25102, n25103,
    n25104, n25105, n25106, n25107, n25108, n25109,
    n25110, n25111, n25112, n25113, n25114, n25115,
    n25116, n25117, n25118, n25119, n25120, n25121,
    n25122, n25123, n25124, n25125, n25126, n25127,
    n25128, n25129, n25130, n25131, n25132, n25133,
    n25134, n25135, n25136, n25137, n25138, n25139,
    n25140, n25141, n25142, n25143, n25144, n25145,
    n25146, n25147, n25148, n25149, n25150, n25151,
    n25152, n25153, n25154, n25155, n25156, n25157,
    n25158, n25159, n25160, n25161, n25162, n25163,
    n25164, n25165, n25166, n25167, n25168, n25169,
    n25170, n25171, n25172, n25173, n25174, n25175,
    n25176, n25177, n25178, n25179, n25180, n25181,
    n25182, n25183, n25184, n25185, n25186, n25187,
    n25188, n25189, n25190, n25191, n25192, n25193,
    n25194, n25195, n25196, n25197, n25198, n25199,
    n25200, n25201, n25202, n25203, n25204, n25205,
    n25206, n25207, n25208, n25209, n25210, n25211,
    n25212, n25213, n25214, n25215, n25216, n25217,
    n25218, n25219, n25220, n25221, n25222, n25223,
    n25224, n25225, n25226, n25227, n25228, n25229,
    n25230, n25231, n25232, n25233, n25234, n25235,
    n25236, n25237, n25238, n25239, n25240, n25241,
    n25242, n25243, n25244, n25245, n25246, n25247,
    n25248, n25249, n25250, n25251, n25252, n25253,
    n25254, n25255, n25256, n25257, n25258, n25259,
    n25260, n25261, n25262, n25263, n25264, n25265,
    n25266, n25267, n25268, n25269, n25270, n25271,
    n25272, n25273, n25274, n25275, n25276, n25277,
    n25278, n25279, n25280, n25281, n25282, n25283,
    n25284, n25285, n25286, n25287, n25288, n25289,
    n25290, n25291, n25292, n25293, n25294, n25295,
    n25296, n25297, n25298, n25299, n25300, n25301,
    n25302, n25303, n25304, n25305, n25306, n25307,
    n25308, n25309, n25310, n25311, n25312, n25313,
    n25314, n25315, n25316, n25317, n25318, n25319,
    n25320, n25321, n25322, n25323, n25324, n25325,
    n25326, n25327, n25328, n25329, n25330, n25331,
    n25332, n25333, n25334, n25335, n25336, n25337,
    n25338, n25339, n25340, n25341, n25342, n25343,
    n25344, n25345, n25346, n25347, n25348, n25349,
    n25350, n25351, n25352, n25353, n25354, n25355,
    n25356, n25357, n25358, n25359, n25360, n25361,
    n25362, n25363, n25364, n25365, n25366, n25367,
    n25368, n25369, n25370, n25371, n25372, n25373,
    n25374, n25375, n25376, n25377, n25378, n25379,
    n25380, n25381, n25382, n25383, n25384, n25385,
    n25386, n25387, n25388, n25389, n25390, n25391,
    n25392, n25393, n25394, n25395, n25396, n25397,
    n25398, n25399, n25400, n25401, n25402, n25403,
    n25404, n25405, n25406, n25407, n25408, n25409,
    n25410, n25411, n25412, n25413, n25414, n25415,
    n25416, n25417, n25418, n25419, n25420, n25421,
    n25422, n25423, n25424, n25425, n25426, n25427,
    n25428, n25429, n25430, n25431, n25432, n25433,
    n25434, n25435, n25436, n25437, n25438, n25439,
    n25440, n25441, n25442, n25443, n25444, n25445,
    n25446, n25447, n25448, n25449, n25450, n25451,
    n25452, n25453, n25454, n25455, n25456, n25457,
    n25458, n25459, n25460, n25461, n25462, n25463,
    n25464, n25465, n25466, n25467, n25468, n25469,
    n25470, n25471, n25472, n25473, n25474, n25475,
    n25476, n25477, n25478, n25479, n25480, n25481,
    n25482, n25483, n25484, n25485, n25486, n25487,
    n25488, n25489, n25490, n25491, n25492, n25493,
    n25494, n25495, n25496, n25497, n25498, n25499,
    n25500, n25501, n25502, n25503, n25504, n25505,
    n25506, n25507, n25508, n25509, n25510, n25511,
    n25512, n25513, n25515, n25516, n25517, n25518,
    n25519, n25520, n25521, n25522, n25523, n25524,
    n25525, n25526, n25527, n25528, n25529, n25530,
    n25531, n25532, n25533, n25534, n25535, n25536,
    n25537, n25538, n25539, n25540, n25541, n25542,
    n25543, n25544, n25545, n25546, n25547, n25548,
    n25549, n25550, n25551, n25552, n25553, n25554,
    n25555, n25556, n25557, n25558, n25559, n25560,
    n25561, n25562, n25563, n25564, n25565, n25566,
    n25567, n25568, n25569, n25570, n25571, n25572,
    n25573, n25574, n25575, n25576, n25577, n25578,
    n25579, n25580, n25581, n25582, n25583, n25584,
    n25585, n25586, n25587, n25588, n25589, n25590,
    n25591, n25592, n25593, n25594, n25595, n25596,
    n25597, n25598, n25599, n25600, n25601, n25602,
    n25603, n25604, n25605, n25606, n25607, n25608,
    n25609, n25610, n25611, n25612, n25613, n25614,
    n25615, n25616, n25617, n25618, n25619, n25620,
    n25621, n25622, n25623, n25624, n25625, n25626,
    n25627, n25628, n25629, n25630, n25631, n25632,
    n25633, n25634, n25635, n25636, n25637, n25638,
    n25639, n25640, n25641, n25642, n25643, n25644,
    n25645, n25646, n25647, n25648, n25649, n25650,
    n25651, n25652, n25653, n25654, n25655, n25656,
    n25657, n25658, n25659, n25660, n25661, n25662,
    n25663, n25664, n25665, n25666, n25667, n25668,
    n25669, n25670, n25671, n25672, n25673, n25674,
    n25675, n25676, n25677, n25678, n25679, n25680,
    n25681, n25682, n25683, n25684, n25685, n25686,
    n25687, n25688, n25689, n25690, n25691, n25692,
    n25693, n25694, n25695, n25696, n25697, n25698,
    n25699, n25700, n25701, n25702, n25703, n25704,
    n25705, n25706, n25707, n25708, n25709, n25710,
    n25711, n25712, n25713, n25714, n25715, n25716,
    n25717, n25718, n25719, n25720, n25721, n25722,
    n25723, n25724, n25725, n25726, n25727, n25728,
    n25729, n25730, n25731, n25732, n25733, n25734,
    n25735, n25736, n25737, n25738, n25739, n25740,
    n25741, n25742, n25743, n25744, n25745, n25746,
    n25747, n25748, n25749, n25750, n25751, n25752,
    n25753, n25754, n25755, n25756, n25757, n25758,
    n25759, n25760, n25761, n25762, n25763, n25764,
    n25765, n25766, n25767, n25768, n25769, n25770,
    n25771, n25772, n25773, n25774, n25775, n25776,
    n25777, n25778, n25779, n25780, n25781, n25782,
    n25783, n25784, n25785, n25786, n25787, n25788,
    n25789, n25790, n25791, n25792, n25793, n25794,
    n25795, n25796, n25797, n25798, n25799, n25800,
    n25801, n25802, n25803, n25804, n25805, n25806,
    n25807, n25808, n25809, n25810, n25811, n25812,
    n25813, n25814, n25815, n25816, n25817, n25818,
    n25819, n25820, n25821, n25822, n25823, n25824,
    n25825, n25826, n25827, n25828, n25829, n25830,
    n25831, n25832, n25833, n25834, n25835, n25836,
    n25837, n25838, n25839, n25840, n25841, n25842,
    n25843, n25844, n25845, n25846, n25847, n25848,
    n25849, n25850, n25851, n25852, n25853, n25854,
    n25855, n25856, n25857, n25858, n25859, n25860,
    n25861, n25862, n25863, n25864, n25865, n25866,
    n25867, n25868, n25869, n25870, n25871, n25872,
    n25873, n25874, n25875, n25876, n25877, n25878,
    n25879, n25880, n25881, n25882, n25883, n25884,
    n25885, n25886, n25887, n25888, n25889, n25890,
    n25891, n25892, n25893, n25894, n25895, n25896,
    n25897, n25898, n25899, n25900, n25901, n25902,
    n25903, n25904, n25905, n25906, n25907, n25908,
    n25909, n25910, n25911, n25912, n25913, n25914,
    n25915, n25916, n25917, n25918, n25919, n25920,
    n25921, n25922, n25923, n25924, n25925, n25926,
    n25927, n25928, n25929, n25930, n25931, n25932,
    n25933, n25934, n25935, n25936, n25937, n25938,
    n25939, n25940, n25941, n25942, n25943, n25944,
    n25945, n25946, n25947, n25948, n25949, n25950,
    n25951, n25952, n25953, n25954, n25955, n25956,
    n25957, n25958, n25959, n25960, n25961, n25962,
    n25963, n25964, n25965, n25966, n25967, n25968,
    n25969, n25970, n25971, n25972, n25973, n25974,
    n25975, n25976, n25977, n25978, n25979, n25980,
    n25981, n25982, n25983, n25984, n25985, n25986,
    n25987, n25988, n25989, n25990, n25991, n25992,
    n25994, n25995, n25996, n25997, n25998, n25999,
    n26000, n26001, n26002, n26003, n26004, n26005,
    n26006, n26007, n26008, n26009, n26010, n26011,
    n26012, n26013, n26014, n26015, n26016, n26017,
    n26018, n26019, n26020, n26021, n26022, n26023,
    n26024, n26025, n26026, n26027, n26028, n26029,
    n26030, n26031, n26032, n26033, n26034, n26035,
    n26036, n26037, n26038, n26039, n26040, n26041,
    n26042, n26043, n26044, n26045, n26046, n26047,
    n26048, n26049, n26050, n26051, n26052, n26053,
    n26054, n26055, n26056, n26057, n26058, n26059,
    n26060, n26061, n26062, n26063, n26064, n26065,
    n26066, n26067, n26068, n26069, n26070, n26071,
    n26072, n26073, n26074, n26075, n26076, n26077,
    n26078, n26079, n26080, n26081, n26082, n26083,
    n26084, n26085, n26086, n26087, n26088, n26089,
    n26090, n26091, n26092, n26093, n26094, n26095,
    n26096, n26097, n26098, n26099, n26100, n26101,
    n26102, n26103, n26104, n26105, n26106, n26107,
    n26108, n26109, n26110, n26111, n26112, n26113,
    n26114, n26115, n26116, n26117, n26118, n26119,
    n26120, n26121, n26122, n26123, n26124, n26125,
    n26126, n26127, n26128, n26129, n26130, n26131,
    n26132, n26133, n26134, n26135, n26136, n26137,
    n26138, n26139, n26140, n26141, n26142, n26143,
    n26144, n26145, n26146, n26147, n26148, n26149,
    n26150, n26151, n26152, n26153, n26154, n26155,
    n26156, n26157, n26158, n26159, n26160, n26161,
    n26162, n26163, n26164, n26165, n26166, n26167,
    n26168, n26169, n26170, n26171, n26172, n26173,
    n26174, n26175, n26176, n26177, n26178, n26179,
    n26180, n26181, n26182, n26183, n26184, n26185,
    n26186, n26187, n26188, n26189, n26190, n26191,
    n26192, n26193, n26194, n26195, n26196, n26197,
    n26198, n26199, n26200, n26201, n26202, n26203,
    n26204, n26205, n26206, n26207, n26208, n26209,
    n26210, n26211, n26212, n26213, n26214, n26215,
    n26216, n26217, n26218, n26219, n26220, n26221,
    n26222, n26223, n26224, n26225, n26226, n26227,
    n26228, n26229, n26230, n26231, n26232, n26233,
    n26234, n26235, n26236, n26237, n26238, n26239,
    n26240, n26241, n26242, n26243, n26244, n26245,
    n26246, n26247, n26248, n26249, n26250, n26251,
    n26252, n26253, n26254, n26255, n26256, n26257,
    n26258, n26259, n26260, n26261, n26262, n26263,
    n26264, n26265, n26266, n26267, n26268, n26269,
    n26270, n26271, n26272, n26273, n26274, n26275,
    n26276, n26277, n26278, n26279, n26280, n26281,
    n26282, n26283, n26284, n26285, n26286, n26287,
    n26288, n26289, n26290, n26291, n26292, n26293,
    n26294, n26295, n26296, n26297, n26298, n26299,
    n26300, n26301, n26302, n26303, n26304, n26305,
    n26306, n26307, n26308, n26309, n26310, n26311,
    n26312, n26313, n26314, n26315, n26316, n26317,
    n26318, n26319, n26320, n26321, n26322, n26323,
    n26324, n26325, n26326, n26327, n26328, n26329,
    n26330, n26331, n26332, n26333, n26334, n26335,
    n26336, n26337, n26338, n26339, n26340, n26341,
    n26342, n26343, n26344, n26345, n26346, n26347,
    n26348, n26349, n26350, n26351, n26352, n26353,
    n26354, n26355, n26356, n26357, n26358, n26359,
    n26360, n26361, n26362, n26363, n26364, n26365,
    n26366, n26367, n26368, n26369, n26370, n26371,
    n26372, n26373, n26374, n26375, n26376, n26377,
    n26378, n26379, n26380, n26381, n26382, n26383,
    n26384, n26385, n26386, n26387, n26388, n26389,
    n26390, n26391, n26392, n26393, n26394, n26395,
    n26396, n26397, n26398, n26399, n26400, n26401,
    n26402, n26403, n26404, n26405, n26406, n26407,
    n26408, n26409, n26410, n26411, n26412, n26413,
    n26414, n26415, n26416, n26417, n26418, n26419,
    n26420, n26421, n26422, n26423, n26424, n26425,
    n26426, n26427, n26428, n26429, n26430, n26431,
    n26432, n26433, n26434, n26435, n26436, n26437,
    n26438, n26439, n26440, n26441, n26442, n26443,
    n26444, n26445, n26446, n26447, n26448, n26449,
    n26450, n26451, n26452, n26453, n26454, n26455,
    n26456, n26457, n26458, n26459, n26460, n26461,
    n26462, n26463, n26464, n26465, n26466, n26467,
    n26469, n26470, n26471, n26472, n26473, n26474,
    n26475, n26476, n26477, n26478, n26479, n26480,
    n26481, n26482, n26483, n26484, n26485, n26486,
    n26487, n26488, n26489, n26490, n26491, n26492,
    n26493, n26494, n26495, n26496, n26497, n26498,
    n26499, n26500, n26501, n26502, n26503, n26504,
    n26505, n26506, n26507, n26508, n26509, n26510,
    n26511, n26512, n26513, n26514, n26515, n26516,
    n26517, n26518, n26519, n26520, n26521, n26522,
    n26523, n26524, n26525, n26526, n26527, n26528,
    n26529, n26530, n26531, n26532, n26533, n26534,
    n26535, n26536, n26537, n26538, n26539, n26540,
    n26541, n26542, n26543, n26544, n26545, n26546,
    n26547, n26548, n26549, n26550, n26551, n26552,
    n26553, n26554, n26555, n26556, n26557, n26558,
    n26559, n26560, n26561, n26562, n26563, n26564,
    n26565, n26566, n26567, n26568, n26569, n26570,
    n26571, n26572, n26573, n26574, n26575, n26576,
    n26577, n26578, n26579, n26580, n26581, n26582,
    n26583, n26584, n26585, n26586, n26587, n26588,
    n26589, n26590, n26591, n26592, n26593, n26594,
    n26595, n26596, n26597, n26598, n26599, n26600,
    n26601, n26602, n26603, n26604, n26605, n26606,
    n26607, n26608, n26609, n26610, n26611, n26612,
    n26613, n26614, n26615, n26616, n26617, n26618,
    n26619, n26620, n26621, n26622, n26623, n26624,
    n26625, n26626, n26627, n26628, n26629, n26630,
    n26631, n26632, n26633, n26634, n26635, n26636,
    n26637, n26638, n26639, n26640, n26641, n26642,
    n26643, n26644, n26645, n26646, n26647, n26648,
    n26649, n26650, n26651, n26652, n26653, n26654,
    n26655, n26656, n26657, n26658, n26659, n26660,
    n26661, n26662, n26663, n26664, n26665, n26666,
    n26667, n26668, n26669, n26670, n26671, n26672,
    n26673, n26674, n26675, n26676, n26677, n26678,
    n26679, n26680, n26681, n26682, n26683, n26684,
    n26685, n26686, n26687, n26688, n26689, n26690,
    n26691, n26692, n26693, n26694, n26695, n26696,
    n26697, n26698, n26699, n26700, n26701, n26702,
    n26703, n26704, n26705, n26706, n26707, n26708,
    n26709, n26710, n26711, n26712, n26713, n26714,
    n26715, n26716, n26717, n26718, n26719, n26720,
    n26721, n26722, n26723, n26724, n26725, n26726,
    n26727, n26728, n26729, n26730, n26731, n26732,
    n26733, n26734, n26735, n26736, n26737, n26738,
    n26739, n26740, n26741, n26742, n26743, n26744,
    n26745, n26746, n26747, n26748, n26749, n26750,
    n26751, n26752, n26753, n26754, n26755, n26756,
    n26757, n26758, n26759, n26760, n26761, n26762,
    n26763, n26764, n26765, n26766, n26767, n26768,
    n26769, n26770, n26771, n26772, n26773, n26774,
    n26775, n26776, n26777, n26778, n26779, n26780,
    n26781, n26782, n26783, n26784, n26785, n26786,
    n26787, n26788, n26789, n26790, n26791, n26792,
    n26793, n26794, n26795, n26796, n26797, n26798,
    n26799, n26800, n26801, n26802, n26803, n26804,
    n26805, n26806, n26807, n26808, n26809, n26810,
    n26811, n26812, n26813, n26814, n26815, n26816,
    n26817, n26818, n26819, n26820, n26821, n26822,
    n26823, n26824, n26825, n26826, n26827, n26828,
    n26829, n26830, n26831, n26832, n26833, n26834,
    n26835, n26836, n26837, n26838, n26839, n26840,
    n26841, n26842, n26843, n26844, n26845, n26846,
    n26847, n26848, n26849, n26850, n26851, n26852,
    n26853, n26854, n26855, n26856, n26857, n26858,
    n26859, n26860, n26861, n26862, n26863, n26864,
    n26865, n26866, n26867, n26868, n26869, n26870,
    n26871, n26872, n26873, n26874, n26875, n26876,
    n26877, n26878, n26879, n26880, n26881, n26882,
    n26883, n26884, n26885, n26886, n26887, n26888,
    n26889, n26890, n26891, n26892, n26893, n26894,
    n26895, n26896, n26897, n26898, n26899, n26900,
    n26901, n26902, n26903, n26904, n26905, n26906,
    n26907, n26908, n26909, n26910, n26911, n26912,
    n26913, n26914, n26915, n26916, n26917, n26918,
    n26919, n26920, n26921, n26922, n26923, n26924,
    n26925, n26926, n26927, n26928, n26929, n26930,
    n26931, n26932, n26933, n26934, n26935, n26936,
    n26937, n26938, n26939, n26940, n26941, n26942,
    n26944, n26945, n26946, n26947, n26948, n26949,
    n26950, n26951, n26952, n26953, n26954, n26955,
    n26956, n26957, n26958, n26959, n26960, n26961,
    n26962, n26963, n26964, n26965, n26966, n26967,
    n26968, n26969, n26970, n26971, n26972, n26973,
    n26974, n26975, n26976, n26977, n26978, n26979,
    n26980, n26981, n26982, n26983, n26984, n26985,
    n26986, n26987, n26988, n26989, n26990, n26991,
    n26992, n26993, n26994, n26995, n26996, n26997,
    n26998, n26999, n27000, n27001, n27002, n27003,
    n27004, n27005, n27006, n27007, n27008, n27009,
    n27010, n27011, n27012, n27013, n27014, n27015,
    n27016, n27017, n27018, n27019, n27020, n27021,
    n27022, n27023, n27024, n27025, n27026, n27027,
    n27028, n27029, n27030, n27031, n27032, n27033,
    n27034, n27035, n27036, n27037, n27038, n27039,
    n27040, n27041, n27042, n27043, n27044, n27045,
    n27046, n27047, n27048, n27049, n27050, n27051,
    n27052, n27053, n27054, n27055, n27056, n27057,
    n27058, n27059, n27060, n27061, n27062, n27063,
    n27064, n27065, n27066, n27067, n27068, n27069,
    n27070, n27071, n27072, n27073, n27074, n27075,
    n27076, n27077, n27078, n27079, n27080, n27081,
    n27082, n27083, n27084, n27085, n27086, n27087,
    n27088, n27089, n27090, n27091, n27092, n27093,
    n27094, n27095, n27096, n27097, n27098, n27099,
    n27100, n27101, n27102, n27103, n27104, n27105,
    n27106, n27107, n27108, n27109, n27110, n27111,
    n27112, n27113, n27114, n27115, n27116, n27117,
    n27118, n27119, n27120, n27121, n27122, n27123,
    n27124, n27125, n27126, n27127, n27128, n27129,
    n27130, n27131, n27132, n27133, n27134, n27135,
    n27136, n27137, n27138, n27139, n27140, n27141,
    n27142, n27143, n27144, n27145, n27146, n27147,
    n27148, n27149, n27150, n27151, n27152, n27153,
    n27154, n27155, n27156, n27157, n27158, n27159,
    n27160, n27161, n27162, n27163, n27164, n27165,
    n27166, n27167, n27168, n27169, n27170, n27171,
    n27172, n27173, n27174, n27175, n27176, n27177,
    n27178, n27179, n27180, n27181, n27182, n27183,
    n27184, n27185, n27186, n27187, n27188, n27189,
    n27190, n27191, n27192, n27193, n27194, n27195,
    n27196, n27197, n27198, n27199, n27200, n27201,
    n27202, n27203, n27204, n27205, n27206, n27207,
    n27208, n27209, n27210, n27211, n27212, n27213,
    n27214, n27215, n27216, n27217, n27218, n27219,
    n27220, n27221, n27222, n27223, n27224, n27225,
    n27226, n27227, n27228, n27229, n27230, n27231,
    n27232, n27233, n27234, n27235, n27236, n27237,
    n27238, n27239, n27240, n27241, n27242, n27243,
    n27244, n27245, n27246, n27247, n27248, n27249,
    n27250, n27251, n27252, n27253, n27254, n27255,
    n27256, n27257, n27258, n27259, n27260, n27261,
    n27262, n27263, n27264, n27265, n27266, n27267,
    n27268, n27269, n27270, n27271, n27272, n27273,
    n27274, n27275, n27276, n27277, n27278, n27279,
    n27280, n27281, n27282, n27283, n27284, n27285,
    n27286, n27287, n27288, n27289, n27290, n27291,
    n27292, n27293, n27294, n27295, n27296, n27297,
    n27298, n27299, n27300, n27301, n27302, n27303,
    n27304, n27305, n27306, n27307, n27308, n27309,
    n27310, n27311, n27312, n27313, n27314, n27315,
    n27316, n27317, n27318, n27319, n27320, n27321,
    n27322, n27323, n27324, n27325, n27326, n27327,
    n27328, n27329, n27330, n27331, n27332, n27333,
    n27334, n27335, n27336, n27337, n27338, n27339,
    n27340, n27341, n27342, n27343, n27344, n27345,
    n27346, n27347, n27348, n27349, n27350, n27351,
    n27352, n27353, n27354, n27355, n27356, n27357,
    n27358, n27359, n27360, n27361, n27362, n27363,
    n27364, n27365, n27366, n27367, n27368, n27369,
    n27370, n27371, n27372, n27373, n27374, n27375,
    n27376, n27377, n27378, n27379, n27380, n27381,
    n27382, n27383, n27384, n27385, n27386, n27387,
    n27388, n27389, n27390, n27391, n27392, n27393,
    n27394, n27395, n27396, n27397, n27398, n27399,
    n27400, n27401, n27402, n27403, n27404, n27405,
    n27406, n27407, n27408, n27409, n27410, n27411,
    n27413, n27414, n27415, n27416, n27417, n27418,
    n27419, n27420, n27421, n27422, n27423, n27424,
    n27425, n27426, n27427, n27428, n27429, n27430,
    n27431, n27432, n27433, n27434, n27435, n27436,
    n27437, n27438, n27439, n27440, n27441, n27442,
    n27443, n27444, n27445, n27446, n27447, n27448,
    n27449, n27450, n27451, n27452, n27453, n27454,
    n27455, n27456, n27457, n27458, n27459, n27460,
    n27461, n27462, n27463, n27464, n27465, n27466,
    n27467, n27468, n27469, n27470, n27471, n27472,
    n27473, n27474, n27475, n27476, n27477, n27478,
    n27479, n27480, n27481, n27482, n27483, n27484,
    n27485, n27486, n27487, n27488, n27489, n27490,
    n27491, n27492, n27493, n27494, n27495, n27496,
    n27497, n27498, n27499, n27500, n27501, n27502,
    n27503, n27504, n27505, n27506, n27507, n27508,
    n27509, n27510, n27511, n27512, n27513, n27514,
    n27515, n27516, n27517, n27518, n27519, n27520,
    n27521, n27522, n27523, n27524, n27525, n27526,
    n27527, n27528, n27529, n27530, n27531, n27532,
    n27533, n27534, n27535, n27536, n27537, n27538,
    n27539, n27540, n27541, n27542, n27543, n27544,
    n27545, n27546, n27547, n27548, n27549, n27550,
    n27551, n27552, n27553, n27554, n27555, n27556,
    n27557, n27558, n27559, n27560, n27561, n27562,
    n27563, n27564, n27565, n27566, n27567, n27568,
    n27569, n27570, n27571, n27572, n27573, n27574,
    n27575, n27576, n27577, n27578, n27579, n27580,
    n27581, n27582, n27583, n27584, n27585, n27586,
    n27587, n27588, n27589, n27590, n27591, n27592,
    n27593, n27594, n27595, n27596, n27597, n27598,
    n27599, n27600, n27601, n27602, n27603, n27604,
    n27605, n27606, n27607, n27608, n27609, n27610,
    n27611, n27612, n27613, n27614, n27615, n27616,
    n27617, n27618, n27619, n27620, n27621, n27622,
    n27623, n27624, n27625, n27626, n27627, n27628,
    n27629, n27630, n27631, n27632, n27633, n27634,
    n27635, n27636, n27637, n27638, n27639, n27640,
    n27641, n27642, n27643, n27644, n27645, n27646,
    n27647, n27648, n27649, n27650, n27651, n27652,
    n27653, n27654, n27655, n27656, n27657, n27658,
    n27659, n27660, n27661, n27662, n27663, n27664,
    n27665, n27666, n27667, n27668, n27669, n27670,
    n27671, n27672, n27673, n27674, n27675, n27676,
    n27677, n27678, n27679, n27680, n27681, n27682,
    n27683, n27684, n27685, n27686, n27687, n27688,
    n27689, n27690, n27691, n27692, n27693, n27694,
    n27695, n27696, n27697, n27698, n27699, n27700,
    n27701, n27702, n27703, n27704, n27705, n27706,
    n27707, n27708, n27709, n27710, n27711, n27712,
    n27713, n27714, n27715, n27716, n27717, n27718,
    n27719, n27720, n27721, n27722, n27723, n27724,
    n27725, n27726, n27727, n27728, n27729, n27730,
    n27731, n27732, n27733, n27734, n27735, n27736,
    n27737, n27738, n27739, n27740, n27741, n27742,
    n27743, n27744, n27745, n27746, n27747, n27748,
    n27749, n27750, n27751, n27752, n27753, n27754,
    n27755, n27756, n27757, n27758, n27759, n27760,
    n27761, n27762, n27763, n27764, n27765, n27766,
    n27767, n27768, n27769, n27770, n27771, n27772,
    n27773, n27774, n27775, n27776, n27777, n27778,
    n27779, n27780, n27781, n27782, n27783, n27784,
    n27785, n27786, n27787, n27788, n27789, n27790,
    n27791, n27792, n27793, n27794, n27795, n27796,
    n27797, n27798, n27799, n27800, n27801, n27802,
    n27803, n27804, n27805, n27806, n27807, n27808,
    n27809, n27810, n27811, n27812, n27813, n27814,
    n27815, n27816, n27817, n27818, n27819, n27820,
    n27821, n27822, n27823, n27824, n27825, n27826,
    n27827, n27828, n27829, n27830, n27831, n27832,
    n27833, n27834, n27835, n27836, n27837, n27838,
    n27839, n27840, n27841, n27842, n27843, n27844,
    n27845, n27846, n27847, n27848, n27849, n27850,
    n27851, n27852, n27853, n27854, n27855, n27856,
    n27857, n27858, n27859, n27860, n27861, n27862,
    n27863, n27864, n27865, n27866, n27867, n27868,
    n27869, n27870, n27871, n27872, n27873, n27874,
    n27875, n27876, n27877, n27878, n27879, n27880,
    n27882, n27883, n27884, n27885, n27886, n27887,
    n27888, n27889, n27890, n27891, n27892, n27893,
    n27894, n27895, n27896, n27897, n27898, n27899,
    n27900, n27901, n27902, n27903, n27904, n27905,
    n27906, n27907, n27908, n27909, n27910, n27911,
    n27912, n27913, n27914, n27915, n27916, n27917,
    n27918, n27919, n27920, n27921, n27922, n27923,
    n27924, n27925, n27926, n27927, n27928, n27929,
    n27930, n27931, n27932, n27933, n27934, n27935,
    n27936, n27937, n27938, n27939, n27940, n27941,
    n27942, n27943, n27944, n27945, n27946, n27947,
    n27948, n27949, n27950, n27951, n27952, n27953,
    n27954, n27955, n27956, n27957, n27958, n27959,
    n27960, n27961, n27962, n27963, n27964, n27965,
    n27966, n27967, n27968, n27969, n27970, n27971,
    n27972, n27973, n27974, n27975, n27976, n27977,
    n27978, n27979, n27980, n27981, n27982, n27983,
    n27984, n27985, n27986, n27987, n27988, n27989,
    n27990, n27991, n27992, n27993, n27994, n27995,
    n27996, n27997, n27998, n27999, n28000, n28001,
    n28002, n28003, n28004, n28005, n28006, n28007,
    n28008, n28009, n28010, n28011, n28012, n28013,
    n28014, n28015, n28016, n28017, n28018, n28019,
    n28020, n28021, n28022, n28023, n28024, n28025,
    n28026, n28027, n28028, n28029, n28030, n28031,
    n28032, n28033, n28034, n28035, n28036, n28037,
    n28038, n28039, n28040, n28041, n28042, n28043,
    n28044, n28045, n28046, n28047, n28048, n28049,
    n28050, n28051, n28052, n28053, n28054, n28055,
    n28056, n28057, n28058, n28059, n28060, n28061,
    n28062, n28063, n28064, n28065, n28066, n28067,
    n28068, n28069, n28070, n28071, n28072, n28073,
    n28074, n28075, n28076, n28077, n28078, n28079,
    n28080, n28081, n28082, n28083, n28084, n28085,
    n28086, n28087, n28088, n28089, n28090, n28091,
    n28092, n28093, n28094, n28095, n28096, n28097,
    n28098, n28099, n28100, n28101, n28102, n28103,
    n28104, n28105, n28106, n28107, n28108, n28109,
    n28110, n28111, n28112, n28113, n28114, n28115,
    n28116, n28117, n28118, n28119, n28120, n28121,
    n28122, n28123, n28124, n28125, n28126, n28127,
    n28128, n28129, n28130, n28131, n28132, n28133,
    n28134, n28135, n28136, n28137, n28138, n28139,
    n28140, n28141, n28142, n28143, n28144, n28145,
    n28146, n28147, n28148, n28149, n28150, n28151,
    n28152, n28153, n28154, n28155, n28156, n28157,
    n28158, n28159, n28160, n28161, n28162, n28163,
    n28164, n28165, n28166, n28167, n28168, n28169,
    n28170, n28171, n28172, n28173, n28174, n28175,
    n28176, n28177, n28178, n28179, n28180, n28181,
    n28182, n28183, n28184, n28185, n28186, n28187,
    n28188, n28189, n28190, n28191, n28192, n28193,
    n28194, n28195, n28196, n28197, n28198, n28199,
    n28200, n28201, n28202, n28203, n28204, n28205,
    n28206, n28207, n28208, n28209, n28210, n28211,
    n28212, n28213, n28214, n28215, n28216, n28217,
    n28218, n28219, n28220, n28221, n28222, n28223,
    n28224, n28225, n28226, n28227, n28228, n28229,
    n28230, n28231, n28232, n28233, n28234, n28235,
    n28236, n28237, n28238, n28239, n28240, n28241,
    n28242, n28243, n28244, n28245, n28246, n28247,
    n28248, n28249, n28250, n28251, n28252, n28253,
    n28254, n28255, n28256, n28257, n28258, n28259,
    n28260, n28261, n28262, n28263, n28264, n28265,
    n28266, n28267, n28268, n28269, n28270, n28271,
    n28272, n28273, n28274, n28275, n28276, n28277,
    n28278, n28279, n28280, n28281, n28282, n28283,
    n28284, n28285, n28286, n28287, n28288, n28289,
    n28290, n28291, n28292, n28293, n28294, n28295,
    n28296, n28297, n28298, n28299, n28300, n28301,
    n28302, n28303, n28304, n28305, n28306, n28307,
    n28308, n28309, n28310, n28311, n28312, n28313,
    n28314, n28315, n28316, n28317, n28318, n28319,
    n28320, n28321, n28322, n28323, n28324, n28325,
    n28326, n28327, n28328, n28329, n28330, n28331,
    n28332, n28333, n28334, n28335, n28336, n28337,
    n28338, n28339, n28340, n28341, n28342, n28343,
    n28344, n28345, n28346, n28347, n28348, n28349,
    n28351, n28352, n28353, n28354, n28355, n28356,
    n28357, n28358, n28359, n28360, n28361, n28362,
    n28363, n28364, n28365, n28366, n28367, n28368,
    n28369, n28370, n28371, n28372, n28373, n28374,
    n28375, n28376, n28377, n28378, n28379, n28380,
    n28381, n28382, n28383, n28384, n28385, n28386,
    n28387, n28388, n28389, n28390, n28391, n28392,
    n28393, n28394, n28395, n28396, n28397, n28398,
    n28399, n28400, n28401, n28402, n28403, n28404,
    n28405, n28406, n28407, n28408, n28409, n28410,
    n28411, n28412, n28413, n28414, n28415, n28416,
    n28417, n28418, n28419, n28420, n28421, n28422,
    n28423, n28424, n28425, n28426, n28427, n28428,
    n28429, n28430, n28431, n28432, n28433, n28434,
    n28435, n28436, n28437, n28438, n28439, n28440,
    n28441, n28442, n28443, n28444, n28445, n28446,
    n28447, n28448, n28449, n28450, n28451, n28452,
    n28453, n28454, n28455, n28456, n28457, n28458,
    n28459, n28460, n28461, n28462, n28463, n28464,
    n28465, n28466, n28467, n28468, n28469, n28470,
    n28471, n28472, n28473, n28474, n28475, n28476,
    n28477, n28478, n28479, n28480, n28481, n28482,
    n28483, n28484, n28485, n28486, n28487, n28488,
    n28489, n28490, n28491, n28492, n28493, n28494,
    n28495, n28496, n28497, n28498, n28499, n28500,
    n28501, n28502, n28503, n28504, n28505, n28506,
    n28507, n28508, n28509, n28510, n28511, n28512,
    n28513, n28514, n28515, n28516, n28517, n28518,
    n28519, n28520, n28521, n28522, n28523, n28524,
    n28525, n28526, n28527, n28528, n28529, n28530,
    n28531, n28532, n28533, n28534, n28535, n28536,
    n28537, n28538, n28539, n28540, n28541, n28542,
    n28543, n28544, n28545, n28546, n28547, n28548,
    n28549, n28550, n28551, n28552, n28553, n28554,
    n28555, n28556, n28557, n28558, n28559, n28560,
    n28561, n28562, n28563, n28564, n28565, n28566,
    n28567, n28568, n28569, n28570, n28571, n28572,
    n28573, n28574, n28575, n28576, n28577, n28578,
    n28579, n28580, n28581, n28582, n28583, n28584,
    n28585, n28586, n28587, n28588, n28589, n28590,
    n28591, n28592, n28593, n28594, n28595, n28596,
    n28597, n28598, n28599, n28600, n28601, n28602,
    n28603, n28604, n28605, n28606, n28607, n28608,
    n28609, n28610, n28611, n28612, n28613, n28614,
    n28615, n28616, n28617, n28618, n28619, n28620,
    n28621, n28622, n28623, n28624, n28625, n28626,
    n28627, n28628, n28629, n28630, n28631, n28632,
    n28633, n28634, n28635, n28636, n28637, n28638,
    n28639, n28640, n28641, n28642, n28643, n28644,
    n28645, n28646, n28647, n28648, n28649, n28650,
    n28651, n28652, n28653, n28654, n28655, n28656,
    n28657, n28658, n28659, n28660, n28661, n28662,
    n28663, n28664, n28665, n28666, n28667, n28668,
    n28669, n28670, n28671, n28672, n28673, n28674,
    n28675, n28676, n28677, n28678, n28679, n28680,
    n28681, n28682, n28683, n28684, n28685, n28686,
    n28687, n28688, n28689, n28690, n28691, n28692,
    n28693, n28694, n28695, n28696, n28697, n28698,
    n28699, n28700, n28701, n28702, n28703, n28704,
    n28705, n28706, n28707, n28708, n28709, n28710,
    n28711, n28712, n28713, n28714, n28715, n28716,
    n28717, n28718, n28719, n28720, n28721, n28722,
    n28723, n28724, n28725, n28726, n28727, n28728,
    n28729, n28730, n28731, n28732, n28733, n28734,
    n28735, n28736, n28737, n28738, n28739, n28740,
    n28741, n28742, n28743, n28744, n28745, n28746,
    n28747, n28748, n28749, n28750, n28751, n28752,
    n28753, n28754, n28755, n28756, n28757, n28758,
    n28759, n28760, n28761, n28762, n28763, n28764,
    n28765, n28766, n28767, n28768, n28769, n28770,
    n28771, n28772, n28773, n28774, n28775, n28776,
    n28777, n28778, n28779, n28780, n28781, n28782,
    n28783, n28784, n28785, n28786, n28787, n28788,
    n28789, n28790, n28791, n28792, n28793, n28794,
    n28795, n28796, n28797, n28798, n28799, n28800,
    n28801, n28802, n28803, n28804, n28805, n28806,
    n28807, n28808, n28809, n28810, n28811, n28812,
    n28813, n28814, n28815, n28816, n28817, n28818,
    n28819, n28820, n28821, n28822, n28823, n28824,
    n28826, n28827, n28828, n28829, n28830, n28831,
    n28832, n28833, n28834, n28835, n28836, n28837,
    n28838, n28839, n28840, n28841, n28842, n28843,
    n28844, n28845, n28846, n28847, n28848, n28849,
    n28850, n28851, n28852, n28853, n28854, n28855,
    n28856, n28857, n28858, n28859, n28860, n28861,
    n28862, n28863, n28864, n28865, n28866, n28867,
    n28868, n28869, n28870, n28871, n28872, n28873,
    n28874, n28875, n28876, n28877, n28878, n28879,
    n28880, n28881, n28882, n28883, n28884, n28885,
    n28886, n28887, n28888, n28889, n28890, n28891,
    n28892, n28893, n28894, n28895, n28896, n28897,
    n28898, n28899, n28900, n28901, n28902, n28903,
    n28904, n28905, n28906, n28907, n28908, n28909,
    n28910, n28911, n28912, n28913, n28914, n28915,
    n28916, n28917, n28918, n28919, n28920, n28921,
    n28922, n28923, n28924, n28925, n28926, n28927,
    n28928, n28929, n28930, n28931, n28932, n28933,
    n28934, n28935, n28936, n28937, n28938, n28939,
    n28940, n28941, n28942, n28943, n28944, n28945,
    n28946, n28947, n28948, n28949, n28950, n28951,
    n28952, n28953, n28954, n28955, n28956, n28957,
    n28958, n28959, n28960, n28961, n28962, n28963,
    n28964, n28965, n28966, n28967, n28968, n28969,
    n28970, n28971, n28972, n28973, n28974, n28975,
    n28976, n28977, n28978, n28979, n28980, n28981,
    n28982, n28983, n28984, n28985, n28986, n28987,
    n28988, n28989, n28990, n28991, n28992, n28993,
    n28994, n28995, n28996, n28997, n28998, n28999,
    n29000, n29001, n29002, n29003, n29004, n29005,
    n29006, n29007, n29008, n29009, n29010, n29011,
    n29012, n29013, n29014, n29015, n29016, n29017,
    n29018, n29019, n29020, n29021, n29022, n29023,
    n29024, n29025, n29026, n29027, n29028, n29029,
    n29030, n29031, n29032, n29033, n29034, n29035,
    n29036, n29037, n29038, n29039, n29040, n29041,
    n29042, n29043, n29044, n29045, n29046, n29047,
    n29048, n29049, n29050, n29051, n29052, n29053,
    n29054, n29055, n29056, n29057, n29058, n29059,
    n29060, n29061, n29062, n29063, n29064, n29065,
    n29066, n29067, n29068, n29069, n29070, n29071,
    n29072, n29073, n29074, n29075, n29076, n29077,
    n29078, n29079, n29080, n29081, n29082, n29083,
    n29084, n29085, n29086, n29087, n29088, n29089,
    n29090, n29091, n29092, n29093, n29094, n29095,
    n29096, n29097, n29098, n29099, n29100, n29101,
    n29102, n29103, n29104, n29105, n29106, n29107,
    n29108, n29109, n29110, n29111, n29112, n29113,
    n29114, n29115, n29116, n29117, n29118, n29119,
    n29120, n29121, n29122, n29123, n29124, n29125,
    n29126, n29127, n29128, n29129, n29130, n29131,
    n29132, n29133, n29134, n29135, n29136, n29137,
    n29138, n29139, n29140, n29141, n29142, n29143,
    n29144, n29145, n29146, n29147, n29148, n29149,
    n29150, n29151, n29152, n29153, n29154, n29155,
    n29156, n29157, n29158, n29159, n29160, n29161,
    n29162, n29163, n29164, n29165, n29166, n29167,
    n29168, n29169, n29170, n29171, n29172, n29173,
    n29174, n29175, n29176, n29177, n29178, n29179,
    n29180, n29181, n29182, n29183, n29184, n29185,
    n29186, n29187, n29188, n29189, n29190, n29191,
    n29192, n29193, n29194, n29195, n29196, n29197,
    n29198, n29199, n29200, n29201, n29202, n29203,
    n29204, n29205, n29206, n29207, n29208, n29209,
    n29210, n29211, n29212, n29213, n29214, n29215,
    n29216, n29217, n29218, n29219, n29220, n29221,
    n29222, n29223, n29224, n29225, n29226, n29227,
    n29228, n29229, n29230, n29231, n29232, n29233,
    n29234, n29235, n29236, n29237, n29238, n29239,
    n29240, n29241, n29242, n29243, n29244, n29245,
    n29246, n29247, n29248, n29249, n29250, n29251,
    n29252, n29253, n29254, n29255, n29256, n29257,
    n29258, n29259, n29260, n29261, n29262, n29263,
    n29264, n29265, n29266, n29267, n29268, n29269,
    n29270, n29271, n29272, n29273, n29274, n29275,
    n29276, n29277, n29278, n29279, n29280, n29281,
    n29282, n29283, n29284, n29285, n29286, n29287,
    n29288, n29289, n29290, n29291, n29292, n29293,
    n29294, n29295, n29296, n29297, n29299, n29300,
    n29301, n29302, n29303, n29304, n29305, n29306,
    n29307, n29308, n29309, n29310, n29311, n29312,
    n29313, n29314, n29315, n29316, n29317, n29318,
    n29319, n29320, n29321, n29322, n29323, n29324,
    n29325, n29326, n29327, n29328, n29329, n29330,
    n29331, n29332, n29333, n29334, n29335, n29336,
    n29337, n29338, n29339, n29340, n29341, n29342,
    n29343, n29344, n29345, n29346, n29347, n29348,
    n29349, n29350, n29351, n29352, n29353, n29354,
    n29355, n29356, n29357, n29358, n29359, n29360,
    n29361, n29362, n29363, n29364, n29365, n29366,
    n29367, n29368, n29369, n29370, n29371, n29372,
    n29373, n29374, n29375, n29376, n29377, n29378,
    n29379, n29380, n29381, n29382, n29383, n29384,
    n29385, n29386, n29387, n29388, n29389, n29390,
    n29391, n29392, n29393, n29394, n29395, n29396,
    n29397, n29398, n29399, n29400, n29401, n29402,
    n29403, n29404, n29405, n29406, n29407, n29408,
    n29409, n29410, n29411, n29412, n29413, n29414,
    n29415, n29416, n29417, n29418, n29419, n29420,
    n29421, n29422, n29423, n29424, n29425, n29426,
    n29427, n29428, n29429, n29430, n29431, n29432,
    n29433, n29434, n29435, n29436, n29437, n29438,
    n29439, n29440, n29441, n29442, n29443, n29444,
    n29445, n29446, n29447, n29448, n29449, n29450,
    n29451, n29452, n29453, n29454, n29455, n29456,
    n29457, n29458, n29459, n29460, n29461, n29462,
    n29463, n29464, n29465, n29466, n29467, n29468,
    n29469, n29470, n29471, n29472, n29473, n29474,
    n29475, n29476, n29477, n29478, n29479, n29480,
    n29481, n29482, n29483, n29484, n29485, n29486,
    n29487, n29488, n29489, n29490, n29491, n29492,
    n29493, n29494, n29495, n29496, n29497, n29498,
    n29499, n29500, n29501, n29502, n29503, n29504,
    n29505, n29506, n29507, n29508, n29509, n29510,
    n29511, n29512, n29513, n29514, n29515, n29516,
    n29517, n29518, n29519, n29520, n29521, n29522,
    n29523, n29524, n29525, n29526, n29527, n29528,
    n29529, n29530, n29531, n29532, n29533, n29534,
    n29535, n29536, n29537, n29538, n29539, n29540,
    n29541, n29542, n29543, n29544, n29545, n29546,
    n29547, n29548, n29549, n29550, n29551, n29552,
    n29553, n29554, n29555, n29556, n29557, n29558,
    n29559, n29560, n29561, n29562, n29563, n29564,
    n29565, n29566, n29567, n29568, n29569, n29570,
    n29571, n29572, n29573, n29574, n29575, n29576,
    n29577, n29578, n29579, n29580, n29581, n29582,
    n29583, n29584, n29585, n29586, n29587, n29588,
    n29589, n29590, n29591, n29592, n29593, n29594,
    n29595, n29596, n29597, n29598, n29599, n29600,
    n29601, n29602, n29603, n29604, n29605, n29606,
    n29607, n29608, n29609, n29610, n29611, n29612,
    n29613, n29614, n29615, n29616, n29617, n29618,
    n29619, n29620, n29621, n29622, n29623, n29624,
    n29625, n29626, n29627, n29628, n29629, n29630,
    n29631, n29632, n29633, n29634, n29635, n29636,
    n29637, n29638, n29639, n29640, n29641, n29642,
    n29643, n29644, n29645, n29646, n29647, n29648,
    n29649, n29650, n29651, n29652, n29653, n29654,
    n29655, n29656, n29657, n29658, n29659, n29660,
    n29661, n29662, n29663, n29664, n29665, n29666,
    n29667, n29668, n29669, n29670, n29671, n29672,
    n29673, n29674, n29675, n29676, n29677, n29678,
    n29679, n29680, n29681, n29682, n29683, n29684,
    n29685, n29686, n29687, n29688, n29689, n29690,
    n29691, n29692, n29693, n29694, n29695, n29696,
    n29697, n29698, n29699, n29700, n29701, n29702,
    n29703, n29704, n29705, n29706, n29707, n29708,
    n29709, n29710, n29711, n29712, n29713, n29714,
    n29715, n29716, n29717, n29718, n29719, n29720,
    n29721, n29722, n29723, n29724, n29725, n29726,
    n29727, n29728, n29729, n29730, n29731, n29732,
    n29733, n29734, n29735, n29736, n29737, n29738,
    n29739, n29740, n29741, n29742, n29743, n29744,
    n29745, n29746, n29747, n29748, n29749, n29750,
    n29751, n29752, n29753, n29754, n29755, n29756,
    n29757, n29758, n29759, n29760, n29761, n29762,
    n29763, n29764, n29765, n29766, n29767, n29768,
    n29769, n29770, n29772, n29773, n29774, n29775,
    n29776, n29777, n29778, n29779, n29780, n29781,
    n29782, n29783, n29784, n29785, n29786, n29787,
    n29788, n29789, n29790, n29791, n29792, n29793,
    n29794, n29795, n29796, n29797, n29798, n29799,
    n29800, n29801, n29802, n29803, n29804, n29805,
    n29806, n29807, n29808, n29809, n29810, n29811,
    n29812, n29813, n29814, n29815, n29816, n29817,
    n29818, n29819, n29820, n29821, n29822, n29823,
    n29824, n29825, n29826, n29827, n29828, n29829,
    n29830, n29831, n29832, n29833, n29834, n29835,
    n29836, n29837, n29838, n29839, n29840, n29841,
    n29842, n29843, n29844, n29845, n29846, n29847,
    n29848, n29849, n29850, n29851, n29852, n29853,
    n29854, n29855, n29856, n29857, n29858, n29859,
    n29860, n29861, n29862, n29863, n29864, n29865,
    n29866, n29867, n29868, n29869, n29870, n29871,
    n29872, n29873, n29874, n29875, n29876, n29877,
    n29878, n29879, n29880, n29881, n29882, n29883,
    n29884, n29885, n29886, n29887, n29888, n29889,
    n29890, n29891, n29892, n29893, n29894, n29895,
    n29896, n29897, n29898, n29899, n29900, n29901,
    n29902, n29903, n29904, n29905, n29906, n29907,
    n29908, n29909, n29910, n29911, n29912, n29913,
    n29914, n29915, n29916, n29917, n29918, n29919,
    n29920, n29921, n29922, n29923, n29924, n29925,
    n29926, n29927, n29928, n29929, n29930, n29931,
    n29932, n29933, n29934, n29935, n29936, n29937,
    n29938, n29939, n29940, n29941, n29942, n29943,
    n29944, n29945, n29946, n29947, n29948, n29949,
    n29950, n29951, n29952, n29953, n29954, n29955,
    n29956, n29957, n29958, n29959, n29960, n29961,
    n29962, n29963, n29964, n29965, n29966, n29967,
    n29968, n29969, n29970, n29971, n29972, n29973,
    n29974, n29975, n29976, n29977, n29978, n29979,
    n29980, n29981, n29982, n29983, n29984, n29985,
    n29986, n29987, n29988, n29989, n29990, n29991,
    n29992, n29993, n29994, n29995, n29996, n29997,
    n29998, n29999, n30000, n30001, n30002, n30003,
    n30004, n30005, n30006, n30007, n30008, n30009,
    n30010, n30011, n30012, n30013, n30014, n30015,
    n30016, n30017, n30018, n30019, n30020, n30021,
    n30022, n30023, n30024, n30025, n30026, n30027,
    n30028, n30029, n30030, n30031, n30032, n30033,
    n30034, n30035, n30036, n30037, n30038, n30039,
    n30040, n30041, n30042, n30043, n30044, n30045,
    n30046, n30047, n30048, n30049, n30050, n30051,
    n30052, n30053, n30054, n30055, n30056, n30057,
    n30058, n30059, n30060, n30061, n30062, n30063,
    n30064, n30065, n30066, n30067, n30068, n30069,
    n30070, n30071, n30072, n30073, n30074, n30075,
    n30076, n30077, n30078, n30079, n30080, n30081,
    n30082, n30083, n30084, n30085, n30086, n30087,
    n30088, n30089, n30090, n30091, n30092, n30093,
    n30094, n30095, n30096, n30097, n30098, n30099,
    n30100, n30101, n30102, n30103, n30104, n30105,
    n30106, n30107, n30108, n30109, n30110, n30111,
    n30112, n30113, n30114, n30115, n30116, n30117,
    n30118, n30119, n30120, n30121, n30122, n30123,
    n30124, n30125, n30126, n30127, n30128, n30129,
    n30130, n30131, n30132, n30133, n30134, n30135,
    n30136, n30137, n30138, n30139, n30140, n30141,
    n30142, n30143, n30144, n30145, n30146, n30147,
    n30148, n30149, n30150, n30151, n30152, n30153,
    n30154, n30155, n30156, n30157, n30158, n30159,
    n30160, n30161, n30162, n30163, n30164, n30165,
    n30166, n30167, n30168, n30169, n30170, n30171,
    n30172, n30173, n30174, n30175, n30176, n30177,
    n30178, n30179, n30180, n30181, n30182, n30183,
    n30184, n30185, n30186, n30187, n30188, n30189,
    n30190, n30191, n30192, n30193, n30194, n30195,
    n30196, n30197, n30198, n30199, n30200, n30201,
    n30202, n30203, n30204, n30205, n30206, n30207,
    n30208, n30209, n30210, n30211, n30212, n30213,
    n30214, n30215, n30216, n30217, n30218, n30219,
    n30220, n30221, n30222, n30223, n30224, n30225,
    n30226, n30227, n30228, n30229, n30230, n30231,
    n30232, n30233, n30234, n30235, n30236, n30237,
    n30238, n30239, n30240, n30241, n30242, n30243,
    n30245, n30246, n30247, n30248, n30249, n30250,
    n30251, n30252, n30253, n30254, n30255, n30256,
    n30257, n30258, n30259, n30260, n30261, n30262,
    n30263, n30264, n30265, n30266, n30267, n30268,
    n30269, n30270, n30271, n30272, n30273, n30274,
    n30275, n30276, n30277, n30278, n30279, n30280,
    n30281, n30282, n30283, n30284, n30285, n30286,
    n30287, n30288, n30289, n30290, n30291, n30292,
    n30293, n30294, n30295, n30296, n30297, n30298,
    n30299, n30300, n30301, n30302, n30303, n30304,
    n30305, n30306, n30307, n30308, n30309, n30310,
    n30311, n30312, n30313, n30314, n30315, n30316,
    n30317, n30318, n30319, n30320, n30321, n30322,
    n30323, n30324, n30325, n30326, n30327, n30328,
    n30329, n30330, n30331, n30332, n30333, n30334,
    n30335, n30336, n30337, n30338, n30339, n30340,
    n30341, n30342, n30343, n30344, n30345, n30346,
    n30347, n30348, n30349, n30350, n30351, n30352,
    n30353, n30354, n30355, n30356, n30357, n30358,
    n30359, n30360, n30361, n30362, n30363, n30364,
    n30365, n30366, n30367, n30368, n30369, n30370,
    n30371, n30372, n30373, n30374, n30375, n30376,
    n30377, n30378, n30379, n30380, n30381, n30382,
    n30383, n30384, n30385, n30386, n30387, n30388,
    n30389, n30390, n30391, n30392, n30393, n30394,
    n30395, n30396, n30397, n30398, n30399, n30400,
    n30401, n30402, n30403, n30404, n30405, n30406,
    n30407, n30408, n30409, n30410, n30411, n30412,
    n30413, n30414, n30415, n30416, n30417, n30418,
    n30419, n30420, n30421, n30422, n30423, n30424,
    n30425, n30426, n30427, n30428, n30429, n30430,
    n30431, n30432, n30433, n30434, n30435, n30436,
    n30437, n30438, n30439, n30440, n30441, n30442,
    n30443, n30444, n30445, n30446, n30447, n30448,
    n30449, n30450, n30451, n30452, n30453, n30454,
    n30455, n30456, n30457, n30458, n30459, n30460,
    n30461, n30462, n30463, n30464, n30465, n30466,
    n30467, n30468, n30469, n30470, n30471, n30472,
    n30473, n30474, n30475, n30476, n30477, n30478,
    n30479, n30480, n30481, n30482, n30483, n30484,
    n30485, n30486, n30487, n30488, n30489, n30490,
    n30491, n30492, n30493, n30494, n30495, n30496,
    n30497, n30498, n30499, n30500, n30501, n30502,
    n30503, n30504, n30505, n30506, n30507, n30508,
    n30509, n30510, n30511, n30512, n30513, n30514,
    n30515, n30516, n30517, n30518, n30519, n30520,
    n30521, n30522, n30523, n30524, n30525, n30526,
    n30527, n30528, n30529, n30530, n30531, n30532,
    n30533, n30534, n30535, n30536, n30537, n30538,
    n30539, n30540, n30541, n30542, n30543, n30544,
    n30545, n30546, n30547, n30548, n30549, n30550,
    n30551, n30552, n30553, n30554, n30555, n30556,
    n30557, n30558, n30559, n30560, n30561, n30562,
    n30563, n30564, n30565, n30566, n30567, n30568,
    n30569, n30570, n30571, n30572, n30573, n30574,
    n30575, n30576, n30577, n30578, n30579, n30580,
    n30581, n30582, n30583, n30584, n30585, n30586,
    n30587, n30588, n30589, n30590, n30591, n30592,
    n30593, n30594, n30595, n30596, n30597, n30598,
    n30599, n30600, n30601, n30602, n30603, n30604,
    n30605, n30606, n30607, n30608, n30609, n30610,
    n30611, n30612, n30613, n30614, n30615, n30616,
    n30617, n30618, n30619, n30620, n30621, n30622,
    n30623, n30624, n30625, n30626, n30627, n30628,
    n30629, n30630, n30631, n30632, n30633, n30634,
    n30635, n30636, n30637, n30638, n30639, n30640,
    n30641, n30642, n30643, n30644, n30645, n30646,
    n30647, n30648, n30649, n30650, n30651, n30652,
    n30653, n30654, n30655, n30656, n30657, n30658,
    n30659, n30660, n30661, n30662, n30663, n30664,
    n30665, n30666, n30667, n30668, n30669, n30670,
    n30671, n30672, n30673, n30674, n30675, n30676,
    n30677, n30678, n30679, n30680, n30681, n30682,
    n30683, n30684, n30685, n30686, n30687, n30688,
    n30689, n30690, n30691, n30692, n30693, n30694,
    n30695, n30696, n30697, n30698, n30699, n30700,
    n30701, n30702, n30703, n30704, n30705, n30706,
    n30707, n30708, n30709, n30710, n30711, n30712,
    n30713, n30714, n30715, n30716, n30717, n30718,
    n30719, n30720, n30721, n30722, n30724, n30725,
    n30726, n30727, n30728, n30729, n30730, n30731,
    n30732, n30733, n30734, n30735, n30736, n30737,
    n30738, n30739, n30740, n30741, n30742, n30743,
    n30744, n30745, n30746, n30747, n30748, n30749,
    n30750, n30751, n30752, n30753, n30754, n30755,
    n30756, n30757, n30758, n30759, n30760, n30761,
    n30762, n30763, n30764, n30765, n30766, n30767,
    n30768, n30769, n30770, n30771, n30772, n30773,
    n30774, n30775, n30776, n30777, n30778, n30779,
    n30780, n30781, n30782, n30783, n30784, n30785,
    n30786, n30787, n30788, n30789, n30790, n30791,
    n30792, n30793, n30794, n30795, n30796, n30797,
    n30798, n30799, n30800, n30801, n30802, n30803,
    n30804, n30805, n30806, n30807, n30808, n30809,
    n30810, n30811, n30812, n30813, n30814, n30815,
    n30816, n30817, n30818, n30819, n30820, n30821,
    n30822, n30823, n30824, n30825, n30826, n30827,
    n30828, n30829, n30830, n30831, n30832, n30833,
    n30834, n30835, n30836, n30837, n30838, n30839,
    n30840, n30841, n30842, n30843, n30844, n30845,
    n30846, n30847, n30848, n30849, n30850, n30851,
    n30852, n30853, n30854, n30855, n30856, n30857,
    n30858, n30859, n30860, n30861, n30862, n30863,
    n30864, n30865, n30866, n30867, n30868, n30869,
    n30870, n30871, n30872, n30873, n30874, n30875,
    n30876, n30877, n30878, n30879, n30880, n30881,
    n30882, n30883, n30884, n30885, n30886, n30887,
    n30888, n30889, n30890, n30891, n30892, n30893,
    n30894, n30895, n30896, n30897, n30898, n30899,
    n30900, n30901, n30902, n30903, n30904, n30905,
    n30906, n30907, n30908, n30909, n30910, n30911,
    n30912, n30913, n30914, n30915, n30916, n30917,
    n30918, n30919, n30920, n30921, n30922, n30923,
    n30924, n30925, n30926, n30927, n30928, n30929,
    n30930, n30931, n30932, n30933, n30934, n30935,
    n30936, n30937, n30938, n30939, n30940, n30941,
    n30942, n30943, n30944, n30945, n30946, n30947,
    n30948, n30949, n30950, n30951, n30952, n30953,
    n30954, n30955, n30956, n30957, n30958, n30959,
    n30960, n30961, n30962, n30963, n30964, n30965,
    n30966, n30967, n30968, n30969, n30970, n30971,
    n30972, n30973, n30974, n30975, n30976, n30977,
    n30978, n30979, n30980, n30981, n30982, n30983,
    n30984, n30985, n30986, n30987, n30988, n30989,
    n30990, n30991, n30992, n30993, n30994, n30995,
    n30996, n30997, n30998, n30999, n31000, n31001,
    n31002, n31003, n31004, n31005, n31006, n31007,
    n31008, n31009, n31010, n31011, n31012, n31013,
    n31014, n31015, n31016, n31017, n31018, n31019,
    n31020, n31021, n31022, n31023, n31024, n31025,
    n31026, n31027, n31028, n31029, n31030, n31031,
    n31032, n31033, n31034, n31035, n31036, n31037,
    n31038, n31039, n31040, n31041, n31042, n31043,
    n31044, n31045, n31046, n31047, n31048, n31049,
    n31050, n31051, n31052, n31053, n31054, n31055,
    n31056, n31057, n31058, n31059, n31060, n31061,
    n31062, n31063, n31064, n31065, n31066, n31067,
    n31068, n31069, n31070, n31071, n31072, n31073,
    n31074, n31075, n31076, n31077, n31078, n31079,
    n31080, n31081, n31082, n31083, n31084, n31085,
    n31086, n31087, n31088, n31089, n31090, n31091,
    n31092, n31093, n31094, n31095, n31096, n31097,
    n31098, n31099, n31100, n31101, n31102, n31103,
    n31104, n31105, n31106, n31107, n31108, n31109,
    n31110, n31111, n31112, n31113, n31114, n31115,
    n31116, n31117, n31118, n31119, n31120, n31121,
    n31122, n31123, n31124, n31125, n31126, n31127,
    n31128, n31129, n31130, n31131, n31132, n31133,
    n31134, n31135, n31136, n31137, n31138, n31139,
    n31140, n31141, n31142, n31143, n31144, n31145,
    n31146, n31147, n31148, n31149, n31150, n31151,
    n31152, n31153, n31154, n31155, n31156, n31157,
    n31158, n31159, n31160, n31161, n31162, n31163,
    n31164, n31165, n31166, n31167, n31168, n31169,
    n31170, n31171, n31172, n31173, n31174, n31175,
    n31176, n31177, n31178, n31179, n31180, n31181,
    n31182, n31183, n31184, n31185, n31186, n31187,
    n31188, n31189, n31190, n31191, n31192, n31193,
    n31194, n31195, n31196, n31197, n31199, n31200,
    n31201, n31202, n31203, n31204, n31205, n31206,
    n31207, n31208, n31209, n31210, n31211, n31212,
    n31213, n31214, n31215, n31216, n31217, n31218,
    n31219, n31220, n31221, n31222, n31223, n31224,
    n31225, n31226, n31227, n31228, n31229, n31230,
    n31231, n31232, n31233, n31234, n31235, n31236,
    n31237, n31238, n31239, n31240, n31241, n31242,
    n31243, n31244, n31245, n31246, n31247, n31248,
    n31249, n31250, n31251, n31252, n31253, n31254,
    n31255, n31256, n31257, n31258, n31259, n31260,
    n31261, n31262, n31263, n31264, n31265, n31266,
    n31267, n31268, n31269, n31270, n31271, n31272,
    n31273, n31274, n31275, n31276, n31277, n31278,
    n31279, n31280, n31281, n31282, n31283, n31284,
    n31285, n31286, n31287, n31288, n31289, n31290,
    n31291, n31292, n31293, n31294, n31295, n31296,
    n31297, n31298, n31299, n31300, n31301, n31302,
    n31303, n31304, n31305, n31306, n31307, n31308,
    n31309, n31310, n31311, n31312, n31313, n31314,
    n31315, n31316, n31317, n31318, n31319, n31320,
    n31321, n31322, n31323, n31324, n31325, n31326,
    n31327, n31328, n31329, n31330, n31331, n31332,
    n31333, n31334, n31335, n31336, n31337, n31338,
    n31339, n31340, n31341, n31342, n31343, n31344,
    n31345, n31346, n31347, n31348, n31349, n31350,
    n31351, n31352, n31353, n31354, n31355, n31356,
    n31357, n31358, n31359, n31360, n31361, n31362,
    n31363, n31364, n31365, n31366, n31367, n31368,
    n31369, n31370, n31371, n31372, n31373, n31374,
    n31375, n31376, n31377, n31378, n31379, n31380,
    n31381, n31382, n31383, n31384, n31385, n31386,
    n31387, n31388, n31389, n31390, n31391, n31392,
    n31393, n31394, n31395, n31396, n31397, n31398,
    n31399, n31400, n31401, n31402, n31403, n31404,
    n31405, n31406, n31407, n31408, n31409, n31410,
    n31411, n31412, n31413, n31414, n31415, n31416,
    n31417, n31418, n31419, n31420, n31421, n31422,
    n31423, n31424, n31425, n31426, n31427, n31428,
    n31429, n31430, n31431, n31432, n31433, n31434,
    n31435, n31436, n31437, n31438, n31439, n31440,
    n31441, n31442, n31443, n31444, n31445, n31446,
    n31447, n31448, n31449, n31450, n31451, n31452,
    n31453, n31454, n31455, n31456, n31457, n31458,
    n31459, n31460, n31461, n31462, n31463, n31464,
    n31465, n31466, n31467, n31468, n31469, n31470,
    n31471, n31472, n31473, n31474, n31475, n31476,
    n31477, n31478, n31479, n31480, n31481, n31482,
    n31483, n31484, n31485, n31486, n31487, n31488,
    n31489, n31490, n31491, n31492, n31493, n31494,
    n31495, n31496, n31497, n31498, n31499, n31500,
    n31501, n31502, n31503, n31504, n31505, n31506,
    n31507, n31508, n31509, n31510, n31511, n31512,
    n31513, n31514, n31515, n31516, n31517, n31518,
    n31519, n31520, n31521, n31522, n31523, n31524,
    n31525, n31526, n31527, n31528, n31529, n31530,
    n31531, n31532, n31533, n31534, n31535, n31536,
    n31537, n31538, n31539, n31540, n31541, n31542,
    n31543, n31544, n31545, n31546, n31547, n31548,
    n31549, n31550, n31551, n31552, n31553, n31554,
    n31555, n31556, n31557, n31558, n31559, n31560,
    n31561, n31562, n31563, n31564, n31565, n31566,
    n31567, n31568, n31569, n31570, n31571, n31572,
    n31573, n31574, n31575, n31576, n31577, n31578,
    n31579, n31580, n31581, n31582, n31583, n31584,
    n31585, n31586, n31587, n31588, n31589, n31590,
    n31591, n31592, n31593, n31594, n31595, n31596,
    n31597, n31598, n31599, n31600, n31601, n31602,
    n31603, n31604, n31605, n31606, n31607, n31608,
    n31609, n31610, n31611, n31612, n31613, n31614,
    n31615, n31616, n31617, n31618, n31619, n31620,
    n31621, n31622, n31623, n31624, n31625, n31626,
    n31627, n31628, n31629, n31630, n31631, n31632,
    n31633, n31634, n31635, n31636, n31637, n31638,
    n31639, n31640, n31641, n31642, n31643, n31644,
    n31645, n31646, n31647, n31648, n31649, n31650,
    n31651, n31652, n31653, n31654, n31655, n31656,
    n31657, n31658, n31659, n31660, n31661, n31662,
    n31663, n31664, n31665, n31666, n31667, n31668,
    n31669, n31670, n31671, n31672, n31674, n31675,
    n31676, n31677, n31678, n31679, n31680, n31681,
    n31682, n31683, n31684, n31685, n31686, n31687,
    n31688, n31689, n31690, n31691, n31692, n31693,
    n31694, n31695, n31696, n31697, n31698, n31699,
    n31700, n31701, n31702, n31703, n31704, n31705,
    n31706, n31707, n31708, n31709, n31710, n31711,
    n31712, n31713, n31714, n31715, n31716, n31717,
    n31718, n31719, n31720, n31721, n31722, n31723,
    n31724, n31725, n31726, n31727, n31728, n31729,
    n31730, n31731, n31732, n31733, n31734, n31735,
    n31736, n31737, n31738, n31739, n31740, n31741,
    n31742, n31743, n31744, n31745, n31746, n31747,
    n31748, n31749, n31750, n31751, n31752, n31753,
    n31754, n31755, n31756, n31757, n31758, n31759,
    n31760, n31761, n31762, n31763, n31764, n31765,
    n31766, n31767, n31768, n31769, n31770, n31771,
    n31772, n31773, n31774, n31775, n31776, n31777,
    n31778, n31779, n31780, n31781, n31782, n31783,
    n31784, n31785, n31786, n31787, n31788, n31789,
    n31790, n31791, n31792, n31793, n31794, n31795,
    n31796, n31797, n31798, n31799, n31800, n31801,
    n31802, n31803, n31804, n31805, n31806, n31807,
    n31808, n31809, n31810, n31811, n31812, n31813,
    n31814, n31815, n31816, n31817, n31818, n31819,
    n31820, n31821, n31822, n31823, n31824, n31825,
    n31826, n31827, n31828, n31829, n31830, n31831,
    n31832, n31833, n31834, n31835, n31836, n31837,
    n31838, n31839, n31840, n31841, n31842, n31843,
    n31844, n31845, n31846, n31847, n31848, n31849,
    n31850, n31851, n31852, n31853, n31854, n31855,
    n31856, n31857, n31858, n31859, n31860, n31861,
    n31862, n31863, n31864, n31865, n31866, n31867,
    n31868, n31869, n31870, n31871, n31872, n31873,
    n31874, n31875, n31876, n31877, n31878, n31879,
    n31880, n31881, n31882, n31883, n31884, n31885,
    n31886, n31887, n31888, n31889, n31890, n31891,
    n31892, n31893, n31894, n31895, n31896, n31897,
    n31898, n31899, n31900, n31901, n31902, n31903,
    n31904, n31905, n31906, n31907, n31908, n31909,
    n31910, n31911, n31912, n31913, n31914, n31915,
    n31916, n31917, n31918, n31919, n31920, n31921,
    n31922, n31923, n31924, n31925, n31926, n31927,
    n31928, n31929, n31930, n31931, n31932, n31933,
    n31934, n31935, n31936, n31937, n31938, n31939,
    n31940, n31941, n31942, n31943, n31944, n31945,
    n31946, n31947, n31948, n31949, n31950, n31951,
    n31952, n31953, n31954, n31955, n31956, n31957,
    n31958, n31959, n31960, n31961, n31962, n31963,
    n31964, n31965, n31966, n31967, n31968, n31969,
    n31970, n31971, n31972, n31973, n31974, n31975,
    n31976, n31977, n31978, n31979, n31980, n31981,
    n31982, n31983, n31984, n31985, n31986, n31987,
    n31988, n31989, n31990, n31991, n31992, n31993,
    n31994, n31995, n31996, n31997, n31998, n31999,
    n32000, n32001, n32002, n32003, n32004, n32005,
    n32006, n32007, n32008, n32009, n32010, n32011,
    n32012, n32013, n32014, n32015, n32016, n32017,
    n32018, n32019, n32020, n32021, n32022, n32023,
    n32024, n32025, n32026, n32027, n32028, n32029,
    n32030, n32031, n32032, n32033, n32034, n32035,
    n32036, n32037, n32038, n32039, n32040, n32041,
    n32042, n32043, n32044, n32045, n32046, n32047,
    n32048, n32049, n32050, n32051, n32052, n32053,
    n32054, n32055, n32056, n32057, n32058, n32059,
    n32060, n32061, n32062, n32063, n32064, n32065,
    n32066, n32067, n32068, n32069, n32070, n32071,
    n32072, n32073, n32074, n32075, n32076, n32077,
    n32078, n32079, n32080, n32081, n32082, n32083,
    n32084, n32085, n32086, n32087, n32088, n32089,
    n32090, n32091, n32092, n32093, n32094, n32095,
    n32096, n32097, n32098, n32099, n32100, n32101,
    n32102, n32103, n32104, n32105, n32106, n32107,
    n32108, n32109, n32110, n32111, n32112, n32113,
    n32114, n32115, n32116, n32117, n32118, n32119,
    n32120, n32121, n32122, n32123, n32124, n32125,
    n32126, n32127, n32128, n32129, n32130, n32131,
    n32132, n32133, n32134, n32135, n32136, n32137,
    n32138, n32139, n32140, n32141, n32142, n32143,
    n32144, n32145, n32146, n32147, n32149, n32150,
    n32151, n32152, n32153, n32154, n32155, n32156,
    n32157, n32158, n32159, n32160, n32161, n32162,
    n32163, n32164, n32165, n32166, n32167, n32168,
    n32169, n32170, n32171, n32172, n32173, n32174,
    n32175, n32176, n32177, n32178, n32179, n32180,
    n32181, n32182, n32183, n32184, n32185, n32186,
    n32187, n32188, n32189, n32190, n32191, n32192,
    n32193, n32194, n32195, n32196, n32197, n32198,
    n32199, n32200, n32201, n32202, n32203, n32204,
    n32205, n32206, n32207, n32208, n32209, n32210,
    n32211, n32212, n32213, n32214, n32215, n32216,
    n32217, n32218, n32219, n32220, n32221, n32222,
    n32223, n32224, n32225, n32226, n32227, n32228,
    n32229, n32230, n32231, n32232, n32233, n32234,
    n32235, n32236, n32237, n32238, n32239, n32240,
    n32241, n32242, n32243, n32244, n32245, n32246,
    n32247, n32248, n32249, n32250, n32251, n32252,
    n32253, n32254, n32255, n32256, n32257, n32258,
    n32259, n32260, n32261, n32262, n32263, n32264,
    n32265, n32266, n32267, n32268, n32269, n32270,
    n32271, n32272, n32273, n32274, n32275, n32276,
    n32277, n32278, n32279, n32280, n32281, n32282,
    n32283, n32284, n32285, n32286, n32287, n32288,
    n32289, n32290, n32291, n32292, n32293, n32294,
    n32295, n32296, n32297, n32298, n32299, n32300,
    n32301, n32302, n32303, n32304, n32305, n32306,
    n32307, n32308, n32309, n32310, n32311, n32312,
    n32313, n32314, n32315, n32316, n32317, n32318,
    n32319, n32320, n32321, n32322, n32323, n32324,
    n32325, n32326, n32327, n32328, n32329, n32330,
    n32331, n32332, n32333, n32334, n32335, n32336,
    n32337, n32338, n32339, n32340, n32341, n32342,
    n32343, n32344, n32345, n32346, n32347, n32348,
    n32349, n32350, n32351, n32352, n32353, n32354,
    n32355, n32356, n32357, n32358, n32359, n32360,
    n32361, n32362, n32363, n32364, n32365, n32366,
    n32367, n32368, n32369, n32370, n32371, n32372,
    n32373, n32374, n32375, n32376, n32377, n32378,
    n32379, n32380, n32381, n32382, n32383, n32384,
    n32385, n32386, n32387, n32388, n32389, n32390,
    n32391, n32392, n32393, n32394, n32395, n32396,
    n32397, n32398, n32399, n32400, n32401, n32402,
    n32403, n32404, n32405, n32406, n32407, n32408,
    n32409, n32410, n32411, n32412, n32413, n32414,
    n32415, n32416, n32417, n32418, n32419, n32420,
    n32421, n32422, n32423, n32424, n32425, n32426,
    n32427, n32428, n32429, n32430, n32431, n32432,
    n32433, n32434, n32435, n32436, n32437, n32438,
    n32439, n32440, n32441, n32442, n32443, n32444,
    n32445, n32446, n32447, n32448, n32449, n32450,
    n32451, n32452, n32453, n32454, n32455, n32456,
    n32457, n32458, n32459, n32460, n32461, n32462,
    n32463, n32464, n32465, n32466, n32467, n32468,
    n32469, n32470, n32471, n32472, n32473, n32474,
    n32475, n32476, n32477, n32478, n32479, n32480,
    n32481, n32482, n32483, n32484, n32485, n32486,
    n32487, n32488, n32489, n32490, n32491, n32492,
    n32493, n32494, n32495, n32496, n32497, n32498,
    n32499, n32500, n32501, n32502, n32503, n32504,
    n32505, n32506, n32507, n32508, n32509, n32510,
    n32511, n32512, n32513, n32514, n32515, n32516,
    n32517, n32518, n32519, n32520, n32521, n32522,
    n32523, n32524, n32525, n32526, n32527, n32528,
    n32529, n32530, n32531, n32532, n32533, n32534,
    n32535, n32536, n32537, n32538, n32539, n32540,
    n32541, n32542, n32543, n32544, n32545, n32546,
    n32547, n32548, n32549, n32550, n32551, n32552,
    n32553, n32554, n32555, n32556, n32557, n32558,
    n32559, n32560, n32561, n32562, n32563, n32564,
    n32565, n32566, n32567, n32568, n32569, n32570,
    n32571, n32572, n32573, n32574, n32575, n32576,
    n32577, n32578, n32579, n32580, n32581, n32582,
    n32583, n32584, n32585, n32586, n32587, n32588,
    n32589, n32590, n32591, n32592, n32593, n32594,
    n32595, n32596, n32597, n32598, n32599, n32600,
    n32601, n32602, n32603, n32604, n32605, n32606,
    n32607, n32608, n32609, n32610, n32611, n32612,
    n32613, n32614, n32615, n32616, n32617, n32619,
    n32620, n32621, n32622, n32623, n32624, n32625,
    n32626, n32627, n32628, n32629, n32630, n32631,
    n32632, n32633, n32634, n32635, n32636, n32637,
    n32638, n32639, n32640, n32641, n32642, n32643,
    n32644, n32645, n32646, n32647, n32648, n32649,
    n32650, n32651, n32652, n32653, n32654, n32655,
    n32656, n32657, n32658, n32659, n32660, n32661,
    n32662, n32663, n32664, n32665, n32666, n32667,
    n32668, n32669, n32670, n32671, n32672, n32673,
    n32674, n32675, n32676, n32677, n32678, n32679,
    n32680, n32681, n32682, n32683, n32684, n32685,
    n32686, n32687, n32688, n32689, n32690, n32691,
    n32692, n32693, n32694, n32695, n32696, n32697,
    n32698, n32699, n32700, n32701, n32702, n32703,
    n32704, n32705, n32706, n32707, n32708, n32709,
    n32710, n32711, n32712, n32713, n32714, n32715,
    n32716, n32717, n32718, n32719, n32720, n32721,
    n32722, n32723, n32724, n32725, n32726, n32727,
    n32728, n32729, n32730, n32731, n32732, n32733,
    n32734, n32735, n32736, n32737, n32738, n32739,
    n32740, n32741, n32742, n32743, n32744, n32745,
    n32746, n32747, n32748, n32749, n32750, n32751,
    n32752, n32753, n32754, n32755, n32756, n32757,
    n32758, n32759, n32760, n32761, n32762, n32763,
    n32764, n32765, n32766, n32767, n32768, n32769,
    n32770, n32771, n32772, n32773, n32774, n32775,
    n32776, n32777, n32778, n32779, n32780, n32781,
    n32782, n32783, n32784, n32785, n32786, n32787,
    n32788, n32789, n32790, n32791, n32792, n32793,
    n32794, n32795, n32796, n32797, n32798, n32799,
    n32800, n32801, n32802, n32803, n32804, n32805,
    n32806, n32807, n32808, n32809, n32810, n32811,
    n32812, n32813, n32814, n32815, n32816, n32817,
    n32818, n32819, n32820, n32821, n32822, n32823,
    n32824, n32825, n32826, n32827, n32828, n32829,
    n32830, n32831, n32832, n32833, n32834, n32835,
    n32836, n32837, n32838, n32839, n32840, n32841,
    n32842, n32843, n32844, n32845, n32846, n32847,
    n32848, n32849, n32850, n32851, n32852, n32853,
    n32854, n32855, n32856, n32857, n32858, n32859,
    n32860, n32861, n32862, n32863, n32864, n32865,
    n32866, n32867, n32868, n32869, n32870, n32871,
    n32872, n32873, n32874, n32875, n32876, n32877,
    n32878, n32879, n32880, n32881, n32882, n32883,
    n32884, n32885, n32886, n32887, n32888, n32889,
    n32890, n32891, n32892, n32893, n32894, n32895,
    n32896, n32897, n32898, n32899, n32900, n32901,
    n32902, n32903, n32904, n32905, n32906, n32907,
    n32908, n32909, n32910, n32911, n32912, n32913,
    n32914, n32915, n32916, n32917, n32918, n32919,
    n32920, n32921, n32922, n32923, n32924, n32925,
    n32926, n32927, n32928, n32929, n32930, n32931,
    n32932, n32933, n32934, n32935, n32936, n32937,
    n32938, n32939, n32940, n32941, n32942, n32943,
    n32944, n32945, n32946, n32947, n32948, n32949,
    n32950, n32951, n32952, n32953, n32954, n32955,
    n32956, n32957, n32958, n32959, n32960, n32961,
    n32962, n32963, n32964, n32965, n32966, n32967,
    n32968, n32969, n32970, n32971, n32972, n32973,
    n32974, n32975, n32976, n32977, n32978, n32979,
    n32980, n32981, n32982, n32983, n32984, n32985,
    n32986, n32987, n32988, n32989, n32990, n32991,
    n32992, n32993, n32994, n32995, n32996, n32997,
    n32998, n32999, n33000, n33001, n33002, n33003,
    n33004, n33005, n33006, n33007, n33008, n33009,
    n33010, n33011, n33012, n33013, n33014, n33015,
    n33016, n33017, n33018, n33019, n33020, n33021,
    n33022, n33023, n33024, n33025, n33026, n33027,
    n33028, n33029, n33030, n33031, n33032, n33033,
    n33034, n33035, n33036, n33037, n33038, n33039,
    n33040, n33041, n33042, n33043, n33044, n33045,
    n33046, n33047, n33048, n33049, n33050, n33051,
    n33052, n33053, n33054, n33055, n33056, n33057,
    n33058, n33059, n33060, n33061, n33062, n33063,
    n33064, n33065, n33066, n33067, n33068, n33069,
    n33070, n33071, n33072, n33073, n33074, n33075,
    n33076, n33077, n33078, n33079, n33080, n33081,
    n33082, n33083, n33085, n33086, n33087, n33088,
    n33089, n33090, n33091, n33092, n33093, n33094,
    n33095, n33096, n33097, n33098, n33099, n33100,
    n33101, n33102, n33103, n33104, n33105, n33106,
    n33107, n33108, n33109, n33110, n33111, n33112,
    n33113, n33114, n33115, n33116, n33117, n33118,
    n33119, n33120, n33121, n33122, n33123, n33124,
    n33125, n33126, n33127, n33128, n33129, n33130,
    n33131, n33132, n33133, n33135, n33136, n33137,
    n33138, n33139, n33140, n33141, n33142, n33143,
    n33144, n33145, n33146, n33147, n33148, n33149,
    n33150, n33151, n33152, n33153, n33154, n33155,
    n33156, n33157, n33158, n33159, n33160, n33161,
    n33162, n33163, n33164, n33165, n33166, n33167,
    n33168, n33169, n33170, n33171, n33172, n33173,
    n33174, n33175, n33176, n33177, n33178, n33179,
    n33180, n33181, n33182, n33183, n33184, n33185,
    n33186, n33187, n33188, n33189, n33190, n33191,
    n33192, n33193, n33194, n33195, n33196, n33197,
    n33198, n33199, n33200, n33201, n33202, n33204,
    n33205, n33206, n33207, n33208, n33209, n33210,
    n33211, n33212, n33213, n33214, n33215, n33216,
    n33217, n33218, n33219, n33220, n33221, n33222,
    n33223, n33224, n33225, n33226, n33227, n33228,
    n33229, n33230, n33231, n33232, n33233, n33234,
    n33235, n33236, n33237, n33238, n33239, n33240,
    n33241, n33242, n33243, n33244, n33245, n33246,
    n33247, n33248, n33249, n33250, n33251, n33252,
    n33253, n33254, n33255, n33256, n33257, n33258,
    n33259, n33260, n33261, n33262, n33263, n33265,
    n33266, n33267, n33268, n33269, n33270, n33271,
    n33272, n33273, n33274, n33275, n33276, n33277,
    n33278, n33279, n33280, n33281, n33282, n33283,
    n33284, n33285, n33286, n33287, n33288, n33289,
    n33290, n33291, n33292, n33293, n33294, n33295,
    n33296, n33297, n33298, n33299, n33300, n33301,
    n33302, n33303, n33304, n33305, n33306, n33307,
    n33308, n33309, n33310, n33311, n33312, n33313,
    n33314, n33315, n33316, n33317, n33318, n33319,
    n33320, n33321, n33322, n33323, n33324, n33325,
    n33326, n33327, n33328, n33329, n33330, n33331,
    n33332, n33333, n33334, n33335, n33336, n33337,
    n33338, n33339, n33340, n33341, n33342, n33343,
    n33344, n33345, n33346, n33347, n33348, n33349,
    n33350, n33351, n33352, n33353, n33354, n33355,
    n33356, n33357, n33358, n33359, n33360, n33361,
    n33362, n33363, n33364, n33365, n33366, n33367,
    n33368, n33369, n33370, n33371, n33372, n33373,
    n33374, n33375, n33376, n33377, n33378, n33379,
    n33380, n33381, n33382, n33383, n33384, n33385,
    n33386, n33387, n33388, n33389, n33390, n33391,
    n33392, n33393, n33394, n33395, n33396, n33397,
    n33398, n33399, n33400, n33401, n33402, n33403,
    n33404, n33405, n33406, n33407, n33408, n33409,
    n33410, n33411, n33412, n33413, n33414, n33415,
    n33416, n33417, n33418, n33419, n33420, n33421,
    n33422, n33423, n33424, n33425, n33426, n33427,
    n33428, n33429, n33430, n33431, n33432, n33433,
    n33434, n33435, n33436, n33437, n33438, n33439,
    n33440, n33441, n33442, n33443, n33444, n33445,
    n33446, n33447, n33448, n33449, n33450, n33451,
    n33452, n33453, n33454, n33455, n33456, n33457,
    n33458, n33459, n33460, n33461, n33462, n33463,
    n33464, n33465, n33466, n33467, n33468, n33469,
    n33470, n33471, n33472, n33473, n33474, n33475,
    n33476, n33477, n33478, n33479, n33480, n33481,
    n33482, n33483, n33484, n33485, n33486, n33487,
    n33488, n33489, n33490, n33491, n33492, n33493,
    n33494, n33495, n33496, n33497, n33498, n33499,
    n33500, n33501, n33502, n33503, n33504, n33505,
    n33506, n33507, n33508, n33509, n33510, n33511,
    n33512, n33513, n33514, n33515, n33516, n33517,
    n33518, n33519, n33520, n33521, n33522, n33523,
    n33524, n33525, n33526, n33527, n33528, n33529,
    n33530, n33531, n33532, n33533, n33534, n33535,
    n33536, n33537, n33538, n33539, n33540, n33541,
    n33542, n33543, n33544, n33545, n33546, n33547,
    n33548, n33549, n33550, n33551, n33552, n33553,
    n33554, n33555, n33556, n33557, n33558, n33559,
    n33560, n33561, n33562, n33563, n33564, n33565,
    n33566, n33567, n33568, n33569, n33570, n33571,
    n33572, n33573, n33574, n33575, n33576, n33577,
    n33578, n33579, n33580, n33581, n33582, n33583,
    n33584, n33585, n33586, n33587, n33588, n33589,
    n33590, n33591, n33592, n33593, n33594, n33595,
    n33596, n33597, n33598, n33599, n33600, n33601,
    n33602, n33603, n33604, n33605, n33606, n33607,
    n33608, n33609, n33610, n33611, n33612, n33613,
    n33614, n33615, n33616, n33617, n33618, n33619,
    n33620, n33621, n33622, n33623, n33624, n33625,
    n33626, n33627, n33628, n33629, n33630, n33631,
    n33632, n33633, n33634, n33635, n33636, n33637,
    n33638, n33639, n33640, n33641, n33642, n33643,
    n33644, n33645, n33646, n33647, n33648, n33649,
    n33650, n33651, n33652, n33653, n33654, n33655,
    n33656, n33657, n33658, n33659, n33660, n33661,
    n33662, n33663, n33664, n33665, n33666, n33667,
    n33668, n33669, n33670, n33671, n33672, n33673,
    n33674, n33675, n33676, n33677, n33678, n33679,
    n33680, n33681, n33682, n33683, n33684, n33685,
    n33686, n33687, n33688, n33689, n33690, n33691,
    n33692, n33693, n33694, n33695, n33696, n33697,
    n33698, n33699, n33700, n33701, n33702, n33703,
    n33704, n33705, n33706, n33707, n33708, n33709,
    n33710, n33711, n33712, n33713, n33714, n33715,
    n33716, n33717, n33718, n33719, n33720, n33721,
    n33722, n33723, n33724, n33725, n33726, n33727,
    n33728, n33729, n33730, n33731, n33732, n33733,
    n33734, n33735, n33736, n33737, n33738, n33739,
    n33740, n33741, n33742, n33743, n33744, n33745,
    n33746, n33747, n33748, n33749, n33750, n33751,
    n33752, n33753, n33754, n33755, n33756, n33757,
    n33758, n33759, n33760, n33761, n33762, n33763,
    n33764, n33765, n33766, n33767, n33768, n33769,
    n33770, n33771, n33772, n33773, n33774, n33775,
    n33776, n33777, n33778, n33779, n33780, n33781,
    n33782, n33783, n33784, n33785, n33786, n33787,
    n33788, n33789, n33790, n33791, n33792, n33793,
    n33794, n33795, n33796, n33797, n33798, n33799,
    n33800, n33801, n33802, n33803, n33804, n33805,
    n33806, n33807, n33808, n33809, n33810, n33811,
    n33812, n33813, n33814, n33815, n33816, n33817,
    n33818, n33819, n33820, n33821, n33822, n33823,
    n33824, n33825, n33826, n33827, n33828, n33829,
    n33830, n33831, n33832, n33833, n33834, n33835,
    n33836, n33837, n33838, n33839, n33840, n33841,
    n33842, n33843, n33844, n33845, n33846, n33847,
    n33848, n33849, n33850, n33851, n33852, n33853,
    n33854, n33855, n33856, n33857, n33858, n33859,
    n33860, n33861, n33862, n33863, n33864, n33865,
    n33866, n33867, n33868, n33869, n33870, n33871,
    n33872, n33873, n33874, n33875, n33876, n33877,
    n33878, n33879, n33880, n33881, n33882, n33883,
    n33884, n33885, n33886, n33887, n33888, n33889,
    n33890, n33891, n33892, n33893, n33894, n33895,
    n33896, n33897, n33899, n33900, n33901, n33902,
    n33903, n33904, n33905, n33906, n33907, n33908,
    n33909, n33910, n33911, n33912, n33913, n33914,
    n33915, n33916, n33917, n33918, n33919, n33920,
    n33921, n33922, n33923, n33924, n33925, n33926,
    n33927, n33928, n33929, n33930, n33931, n33932,
    n33933, n33934, n33935, n33936, n33937, n33938,
    n33939, n33940, n33941, n33942, n33943, n33944,
    n33945, n33946, n33947, n33948, n33949, n33950,
    n33951, n33952, n33953, n33954, n33955, n33956,
    n33957, n33958, n33959, n33960, n33961, n33962,
    n33963, n33964, n33965, n33966, n33967, n33968,
    n33969, n33970, n33971, n33972, n33973, n33974,
    n33975, n33976, n33977, n33978, n33979, n33980,
    n33981, n33982, n33983, n33984, n33985, n33986,
    n33987, n33988, n33989, n33990, n33991, n33992,
    n33993, n33994, n33995, n33996, n33997, n33998,
    n33999, n34000, n34001, n34002, n34003, n34004,
    n34005, n34006, n34007, n34008, n34009, n34010,
    n34011, n34012, n34013, n34014, n34015, n34016,
    n34017, n34018, n34019, n34020, n34021, n34022,
    n34023, n34024, n34025, n34026, n34027, n34028,
    n34029, n34030, n34031, n34032, n34033, n34034,
    n34035, n34036, n34037, n34038, n34039, n34040,
    n34041, n34042, n34043, n34044, n34045, n34046,
    n34047, n34048, n34049, n34050, n34051, n34052,
    n34053, n34054, n34055, n34056, n34057, n34058,
    n34059, n34060, n34061, n34062, n34063, n34064,
    n34065, n34066, n34067, n34068, n34069, n34070,
    n34071, n34072, n34073, n34074, n34075, n34076,
    n34077, n34078, n34079, n34080, n34081, n34082,
    n34083, n34084, n34085, n34086, n34087, n34088,
    n34089, n34090, n34091, n34092, n34093, n34094,
    n34095, n34096, n34097, n34098, n34099, n34100,
    n34101, n34102, n34103, n34104, n34105, n34106,
    n34107, n34108, n34109, n34110, n34111, n34112,
    n34113, n34114, n34115, n34116, n34117, n34118,
    n34119, n34120, n34121, n34122, n34123, n34124,
    n34125, n34126, n34127, n34128, n34129, n34130,
    n34131, n34132, n34133, n34134, n34135, n34136,
    n34137, n34138, n34139, n34140, n34141, n34142,
    n34143, n34144, n34145, n34146, n34147, n34148,
    n34149, n34150, n34151, n34152, n34153, n34154,
    n34155, n34156, n34157, n34158, n34159, n34160,
    n34161, n34162, n34163, n34164, n34165, n34166,
    n34167, n34168, n34169, n34170, n34171, n34172,
    n34173, n34174, n34175, n34176, n34177, n34178,
    n34179, n34180, n34181, n34182, n34183, n34184,
    n34185, n34186, n34187, n34188, n34190, n34191,
    n34192, n34193, n34194, n34195, n34196, n34197,
    n34198, n34199, n34200, n34201, n34202, n34203,
    n34204, n34205, n34206, n34207, n34208, n34209,
    n34210, n34211, n34212, n34213, n34214, n34215,
    n34216, n34217, n34218, n34219, n34220, n34221,
    n34222, n34223, n34224, n34225, n34226, n34227,
    n34228, n34229, n34230, n34231, n34232, n34233,
    n34234, n34235, n34236, n34237, n34238, n34239,
    n34240, n34241, n34242, n34243, n34244, n34245,
    n34246, n34247, n34248, n34249, n34250, n34251,
    n34252, n34253, n34254, n34255, n34256, n34257,
    n34258, n34259, n34260, n34261, n34262, n34263,
    n34264, n34265, n34266, n34267, n34268, n34269,
    n34270, n34271, n34272, n34273, n34274, n34275,
    n34276, n34277, n34278, n34279, n34280, n34281,
    n34282, n34283, n34284, n34285, n34286, n34287,
    n34288, n34289, n34290, n34291, n34292, n34293,
    n34294, n34295, n34296, n34297, n34298, n34299,
    n34300, n34301, n34302, n34303, n34304, n34305,
    n34306, n34307, n34308, n34309, n34310, n34311,
    n34312, n34313, n34314, n34315, n34316, n34317,
    n34318, n34319, n34320, n34321, n34322, n34323,
    n34324, n34325, n34326, n34327, n34328, n34329,
    n34330, n34331, n34332, n34333, n34334, n34335,
    n34336, n34337, n34338, n34339, n34340, n34341,
    n34342, n34343, n34344, n34345, n34346, n34347,
    n34348, n34349, n34350, n34351, n34352, n34353,
    n34354, n34355, n34356, n34357, n34358, n34359,
    n34360, n34361, n34362, n34363, n34364, n34365,
    n34366, n34367, n34368, n34369, n34370, n34371,
    n34372, n34373, n34374, n34375, n34376, n34377,
    n34378, n34379, n34380, n34381, n34382, n34383,
    n34384, n34385, n34386, n34387, n34388, n34389,
    n34390, n34391, n34392, n34393, n34394, n34395,
    n34396, n34397, n34398, n34399, n34400, n34401,
    n34402, n34403, n34404, n34405, n34406, n34407,
    n34408, n34409, n34410, n34411, n34412, n34413,
    n34414, n34415, n34416, n34417, n34418, n34419,
    n34420, n34421, n34422, n34423, n34424, n34425,
    n34426, n34427, n34428, n34429, n34430, n34431,
    n34432, n34433, n34434, n34435, n34436, n34437,
    n34438, n34439, n34440, n34441, n34442, n34443,
    n34444, n34445, n34446, n34447, n34448, n34449,
    n34450, n34451, n34452, n34453, n34454, n34455,
    n34456, n34457, n34458, n34459, n34460, n34461,
    n34462, n34463, n34464, n34465, n34466, n34468,
    n34469, n34470, n34471, n34472, n34473, n34474,
    n34475, n34476, n34477, n34478, n34479, n34480,
    n34481, n34482, n34483, n34484, n34485, n34486,
    n34487, n34488, n34489, n34490, n34491, n34492,
    n34493, n34494, n34495, n34496, n34497, n34498,
    n34499, n34500, n34501, n34502, n34503, n34504,
    n34505, n34506, n34507, n34508, n34509, n34510,
    n34511, n34512, n34513, n34514, n34515, n34516,
    n34517, n34518, n34519, n34520, n34521, n34522,
    n34523, n34524, n34525, n34526, n34527, n34528,
    n34529, n34530, n34531, n34532, n34533, n34534,
    n34535, n34536, n34537, n34538, n34539, n34540,
    n34541, n34542, n34543, n34544, n34545, n34546,
    n34547, n34548, n34549, n34550, n34551, n34552,
    n34553, n34554, n34555, n34556, n34557, n34558,
    n34559, n34560, n34561, n34562, n34563, n34564,
    n34565, n34566, n34567, n34568, n34569, n34570,
    n34571, n34572, n34573, n34574, n34575, n34576,
    n34577, n34578, n34579, n34580, n34581, n34582,
    n34583, n34584, n34585, n34586, n34587, n34588,
    n34589, n34590, n34591, n34592, n34593, n34594,
    n34595, n34596, n34597, n34598, n34599, n34600,
    n34601, n34602, n34603, n34604, n34605, n34606,
    n34607, n34608, n34609, n34610, n34611, n34612,
    n34613, n34614, n34615, n34616, n34617, n34618,
    n34619, n34620, n34621, n34622, n34623, n34624,
    n34625, n34626, n34627, n34628, n34629, n34630,
    n34631, n34632, n34633, n34634, n34635, n34636,
    n34637, n34638, n34639, n34640, n34641, n34642,
    n34643, n34644, n34645, n34646, n34647, n34648,
    n34649, n34650, n34651, n34652, n34653, n34654,
    n34655, n34656, n34657, n34658, n34659, n34660,
    n34661, n34663, n34664, n34665, n34666, n34667,
    n34668, n34669, n34671, n34672, n34673, n34674,
    n34675, n34676, n34677, n34679, n34680, n34681,
    n34682, n34683, n34684, n34685, n34686, n34687,
    n34688, n34689, n34690, n34691, n34692, n34693,
    n34694, n34695, n34696, n34697, n34698, n34699,
    n34700, n34701, n34702, n34703, n34704, n34705,
    n34706, n34707, n34708, n34709, n34710, n34711,
    n34712, n34713, n34714, n34715, n34716, n34717,
    n34718, n34719, n34720, n34721, n34722, n34723,
    n34724, n34725, n34726, n34727, n34728, n34729,
    n34730, n34731, n34732, n34733, n34734, n34735,
    n34736, n34737, n34738, n34739, n34740, n34741,
    n34742, n34743, n34744, n34745, n34746, n34747,
    n34748, n34749, n34750, n34751, n34752, n34753,
    n34754, n34755, n34756, n34757, n34758, n34759,
    n34760, n34761, n34762, n34763, n34764, n34765,
    n34766, n34767, n34768, n34769, n34770, n34771,
    n34772, n34773, n34774, n34775, n34776, n34777,
    n34778, n34779, n34780, n34781, n34782, n34783,
    n34784, n34785, n34786, n34788, n34789, n34790,
    n34791, n34792, n34793, n34795, n34796, n34797,
    n34798, n34799, n34800, n34801, n34803, n34804,
    n34805, n34806, n34807, n34808, n34809, n34810,
    n34811, n34812, n34813, n34814, n34815, n34816,
    n34817, n34818, n34819, n34820, n34821, n34822,
    n34823, n34824, n34825, n34826, n34827, n34828,
    n34829, n34830, n34831, n34832, n34833, n34834,
    n34835, n34836, n34837, n34838, n34839, n34840,
    n34841, n34842, n34843, n34844, n34845, n34846,
    n34847, n34848, n34849, n34850, n34851, n34852,
    n34853, n34854, n34855, n34856, n34857, n34858,
    n34859, n34860, n34861, n34862, n34863, n34864,
    n34865, n34866, n34867, n34868, n34869, n34870,
    n34871, n34872, n34873, n34874, n34875, n34876,
    n34877, n34878, n34879, n34880, n34881, n34882,
    n34883, n34884, n34885, n34886, n34887, n34888,
    n34889, n34890, n34891, n34892, n34893, n34894,
    n34895, n34896, n34897, n34898, n34899, n34900,
    n34901, n34902, n34903, n34904, n34905, n34906,
    n34907, n34908, n34909, n34910, n34911, n34912,
    n34913, n34914, n34915, n34916, n34917, n34918,
    n34919, n34920, n34921, n34922, n34923, n34924,
    n34925, n34926, n34927, n34928, n34929, n34930,
    n34931, n34932, n34933, n34934, n34935, n34936,
    n34937, n34938, n34939, n34940, n34941, n34942,
    n34943, n34944, n34945, n34946, n34947, n34948,
    n34949, n34950, n34951, n34952, n34953, n34954,
    n34955, n34956, n34957, n34958, n34959, n34960,
    n34961, n34962, n34963, n34964, n34965, n34966,
    n34967, n34968, n34969, n34970, n34971, n34972,
    n34973, n34974, n34975, n34976, n34977, n34978,
    n34979, n34980, n34981, n34982, n34983, n34984,
    n34985, n34986, n34987, n34988, n34989, n34990,
    n34991, n34992, n34993, n34994, n34995, n34996,
    n34997, n34998, n34999, n35000, n35001, n35002,
    n35003, n35004, n35005, n35006, n35007, n35008,
    n35009, n35010, n35011, n35012, n35013, n35014,
    n35015, n35016, n35017, n35018, n35019, n35020,
    n35021, n35022, n35023, n35024, n35025, n35026,
    n35027, n35028, n35029, n35030, n35031, n35032,
    n35033, n35034, n35035, n35036, n35037, n35038,
    n35039, n35040, n35041, n35042, n35043, n35044,
    n35045, n35046, n35047, n35048, n35049, n35050,
    n35051, n35052, n35053, n35054, n35055, n35056,
    n35057, n35058, n35059, n35060, n35061, n35062,
    n35063, n35064, n35065, n35066, n35067, n35068,
    n35069, n35070, n35071, n35072, n35073, n35074,
    n35075, n35076, n35077, n35078, n35079, n35080,
    n35081, n35082, n35083, n35084, n35085, n35086,
    n35087, n35088, n35089, n35090, n35091, n35092,
    n35093, n35094, n35095, n35096, n35097, n35098,
    n35099, n35100, n35101, n35102, n35103, n35104,
    n35105, n35106, n35107, n35108, n35109, n35110,
    n35111, n35112, n35113, n35114, n35115, n35116,
    n35117, n35118, n35119, n35120, n35121, n35122,
    n35123, n35124, n35125, n35126, n35127, n35128,
    n35129, n35130, n35131, n35132, n35133, n35134,
    n35135, n35136, n35137, n35138, n35139, n35140,
    n35141, n35142, n35143, n35144, n35145, n35146,
    n35147, n35148, n35149, n35150, n35151, n35152,
    n35153, n35154, n35155, n35156, n35157, n35158,
    n35159, n35160, n35161, n35162, n35163, n35164,
    n35165, n35166, n35167, n35168, n35169, n35170,
    n35171, n35172, n35173, n35174, n35175, n35176,
    n35177, n35178, n35179, n35180, n35181, n35182,
    n35183, n35184, n35185, n35186, n35187, n35188,
    n35189, n35190, n35191, n35192, n35193, n35194,
    n35195, n35196, n35197, n35198, n35199, n35200,
    n35201, n35202, n35203, n35204, n35205, n35206,
    n35207, n35208, n35209, n35210, n35211, n35212,
    n35213, n35214, n35215, n35216, n35217, n35218,
    n35219, n35220, n35221, n35222, n35223, n35224,
    n35225, n35226, n35227, n35228, n35229, n35230,
    n35231, n35232, n35233, n35234, n35235, n35236,
    n35237, n35238, n35239, n35240, n35241, n35242,
    n35243, n35244, n35245, n35246, n35247, n35248,
    n35249, n35250, n35251, n35252, n35253, n35254,
    n35255, n35256, n35257, n35258, n35259, n35260,
    n35261, n35262, n35263, n35264, n35265, n35266,
    n35267, n35268, n35269, n35270, n35271, n35272,
    n35273, n35274, n35275, n35276, n35277, n35278,
    n35279, n35280, n35281, n35282, n35283, n35284,
    n35285, n35286, n35287, n35288, n35289, n35290,
    n35291, n35292, n35293, n35295, n35296, n35297,
    n35298, n35299, n35300, n35301, n35302, n35303,
    n35304, n35305, n35306, n35307, n35308, n35309,
    n35310, n35311, n35312, n35313, n35314, n35315,
    n35316, n35317, n35318, n35319, n35320, n35321,
    n35322, n35323, n35324, n35325, n35326, n35327,
    n35328, n35329, n35330, n35331, n35332, n35333,
    n35334, n35335, n35336, n35337, n35338, n35339,
    n35340, n35341, n35342, n35343, n35344, n35345,
    n35346, n35347, n35348, n35349, n35350, n35351,
    n35352, n35353, n35354, n35355, n35356, n35357,
    n35358, n35359, n35360, n35361, n35362, n35363,
    n35364, n35365, n35366, n35367, n35368, n35370,
    n35371, n35372, n35373, n35374, n35375, n35376,
    n35377, n35378, n35379, n35380, n35381, n35382,
    n35383, n35384, n35385, n35386, n35387, n35388,
    n35389, n35390, n35391, n35392, n35393, n35394,
    n35395, n35396, n35397, n35398, n35399, n35400,
    n35401, n35402, n35403, n35404, n35405, n35406,
    n35407, n35408, n35409, n35410, n35411, n35412,
    n35413, n35414, n35415, n35416, n35417, n35418,
    n35419, n35420, n35421, n35422, n35423, n35424,
    n35425, n35426, n35427, n35428, n35429, n35430,
    n35431, n35432, n35433, n35434, n35435, n35436,
    n35437, n35438, n35439, n35440, n35441, n35442,
    n35443, n35444, n35445, n35446, n35447, n35448,
    n35449, n35450, n35451, n35452, n35453, n35454,
    n35455, n35456, n35457, n35458, n35459, n35460,
    n35461, n35462, n35463, n35464, n35465, n35466,
    n35467, n35468, n35469, n35470, n35471, n35472,
    n35473, n35474, n35475, n35476, n35477, n35478,
    n35479, n35480, n35481, n35482, n35483, n35484,
    n35485, n35486, n35487, n35488, n35489, n35490,
    n35491, n35492, n35493, n35494, n35495, n35496,
    n35497, n35498, n35499, n35500, n35501, n35502,
    n35503, n35504, n35505, n35506, n35507, n35508,
    n35509, n35510, n35511, n35512, n35513, n35514,
    n35515, n35516, n35517, n35518, n35519, n35520,
    n35521, n35522, n35523, n35524, n35525, n35526,
    n35527, n35529, n35530, n35531, n35532, n35533,
    n35534, n35535, n35536, n35537, n35538, n35539,
    n35540, n35541, n35542, n35543, n35544, n35545,
    n35546, n35547, n35548, n35549, n35550, n35551,
    n35552, n35553, n35554, n35555, n35556, n35557,
    n35558, n35559, n35560, n35561, n35562, n35563,
    n35564, n35565, n35566, n35567, n35568, n35569,
    n35570, n35571, n35572, n35573, n35574, n35575,
    n35576, n35577, n35578, n35579, n35580, n35581,
    n35582, n35583, n35584, n35585, n35586, n35587,
    n35588, n35589, n35590, n35591, n35592, n35593,
    n35594, n35595, n35596, n35597, n35598, n35599,
    n35600, n35601, n35602, n35603, n35604, n35605,
    n35606, n35607, n35608, n35609, n35610, n35611,
    n35612, n35613, n35614, n35615, n35616, n35617,
    n35618, n35619, n35620, n35621, n35622, n35623,
    n35624, n35625, n35626, n35627, n35628, n35629,
    n35630, n35631, n35632, n35633, n35634, n35635,
    n35636, n35637, n35638, n35639, n35640, n35641,
    n35642, n35643, n35644, n35645, n35646, n35647,
    n35648, n35649, n35650, n35651, n35652, n35653,
    n35655, n35656, n35657, n35658, n35659, n35660,
    n35661, n35662, n35663, n35664, n35665, n35666,
    n35667, n35668, n35669, n35670, n35671, n35672,
    n35673, n35674, n35675, n35676, n35677, n35678,
    n35679, n35680, n35682, n35683, n35684, n35685,
    n35686, n35687, n35688, n35689, n35690, n35691,
    n35692, n35693, n35694, n35695, n35696, n35697,
    n35698, n35699, n35700, n35701, n35703, n35704,
    n35705, n35706, n35707, n35708, n35709, n35710,
    n35711, n35712, n35713, n35714, n35715, n35716,
    n35717, n35718, n35719, n35720, n35721, n35722,
    n35724, n35725, n35726, n35727, n35728, n35729,
    n35730, n35731, n35732, n35733, n35734, n35735,
    n35736, n35737, n35738, n35739, n35740, n35741,
    n35742, n35743, n35745, n35746, n35747, n35748,
    n35749, n35750, n35751, n35752, n35753, n35754,
    n35755, n35756, n35757, n35758, n35759, n35760,
    n35761, n35762, n35763, n35764, n35765, n35766,
    n35767, n35768, n35769, n35770, n35771, n35772,
    n35773, n35774, n35775, n35776, n35777, n35778,
    n35779, n35780, n35781, n35782, n35783, n35784,
    n35785, n35786, n35787, n35788, n35789, n35790,
    n35791, n35792, n35793, n35794, n35795, n35796,
    n35797, n35798, n35799, n35800, n35801, n35802,
    n35803, n35804, n35805, n35806, n35807, n35808,
    n35809, n35810, n35811, n35812, n35813, n35814,
    n35815, n35816, n35817, n35818, n35819, n35820,
    n35821, n35822, n35823, n35824, n35825, n35826,
    n35827, n35828, n35829, n35830, n35831, n35832,
    n35833, n35834, n35835, n35836, n35837, n35838,
    n35839, n35840, n35841, n35842, n35843, n35844,
    n35845, n35846, n35847, n35848, n35849, n35850,
    n35851, n35852, n35853, n35854, n35855, n35856,
    n35857, n35858, n35859, n35861, n35862, n35863,
    n35864, n35865, n35866, n35867, n35868, n35869,
    n35870, n35871, n35872, n35873, n35874, n35875,
    n35876, n35877, n35878, n35879, n35880, n35881,
    n35882, n35883, n35884, n35885, n35886, n35887,
    n35888, n35889, n35890, n35891, n35892, n35893,
    n35894, n35895, n35896, n35897, n35898, n35899,
    n35900, n35901, n35902, n35903, n35904, n35905,
    n35906, n35907, n35908, n35909, n35910, n35911,
    n35912, n35913, n35914, n35915, n35916, n35917,
    n35918, n35919, n35920, n35921, n35922, n35923,
    n35924, n35925, n35926, n35927, n35928, n35929,
    n35930, n35931, n35932, n35933, n35934, n35935,
    n35936, n35937, n35938, n35939, n35940, n35941,
    n35942, n35943, n35944, n35945, n35946, n35947,
    n35948, n35949, n35950, n35951, n35952, n35953,
    n35954, n35955, n35956, n35957, n35958, n35959,
    n35960, n35961, n35962, n35963, n35964, n35965,
    n35966, n35967, n35968, n35969, n35970, n35972,
    n35973, n35974, n35975, n35976, n35977, n35978,
    n35979, n35980, n35981, n35982, n35983, n35984,
    n35985, n35986, n35987, n35988, n35989, n35991,
    n35992, n35993, n35994, n35995, n35996, n35998,
    n35999, n36000, n36001, n36002, n36003, n36004,
    n36005, n36006, n36007, n36008, n36009, n36010,
    n36011, n36012, n36013, n36014, n36015, n36016,
    n36017, n36019, n36020, n36021, n36022, n36023,
    n36024, n36026, n36027, n36028, n36029, n36030,
    n36031, n36032, n36033, n36034, n36035, n36036,
    n36037, n36038, n36039, n36040, n36041, n36042,
    n36043, n36044, n36045, n36046, n36047, n36048,
    n36049, n36050, n36051, n36052, n36053, n36054,
    n36055, n36056, n36057, n36058, n36059, n36060,
    n36061, n36062, n36063, n36064, n36065, n36066,
    n36067, n36068, n36069, n36070, n36071, n36072,
    n36073, n36074, n36075, n36076, n36077, n36078,
    n36079, n36080, n36081, n36082, n36083, n36084,
    n36085, n36086, n36087, n36088, n36089, n36090,
    n36091, n36092, n36093, n36094, n36095, n36096,
    n36097, n36098, n36099, n36100, n36101, n36102,
    n36103, n36104, n36105, n36106, n36107, n36108,
    n36109, n36110, n36111, n36112, n36113, n36114,
    n36115, n36116, n36117, n36118, n36119, n36120,
    n36121, n36122, n36123, n36124, n36125, n36126,
    n36127, n36128, n36129, n36130, n36131, n36132,
    n36133, n36135, n36136, n36137, n36138, n36139,
    n36140, n36141, n36142, n36143, n36144, n36145,
    n36146, n36147, n36148, n36149, n36150, n36151,
    n36152, n36153, n36154, n36155, n36156, n36157,
    n36158, n36159, n36160, n36161, n36162, n36163,
    n36164, n36165, n36166, n36167, n36168, n36169,
    n36170, n36171, n36172, n36173, n36174, n36175,
    n36176, n36177, n36178, n36179, n36180, n36181,
    n36182, n36183, n36184, n36185, n36186, n36187,
    n36188, n36189, n36190, n36191, n36192, n36193,
    n36194, n36195, n36196, n36197, n36198, n36199,
    n36200, n36201, n36202, n36203, n36204, n36205,
    n36206, n36207, n36208, n36209, n36210, n36211,
    n36212, n36213, n36214, n36215, n36216, n36217,
    n36218, n36219, n36220, n36221, n36222, n36223,
    n36224, n36225, n36226, n36227, n36228, n36229,
    n36230, n36231, n36232, n36233, n36234, n36235,
    n36236, n36237, n36238, n36239, n36240, n36241,
    n36242, n36243, n36244, n36245, n36246, n36247,
    n36248, n36249, n36250, n36251, n36252, n36253,
    n36254, n36255, n36256, n36257, n36258, n36259,
    n36260, n36261, n36262, n36263, n36264, n36265,
    n36266, n36267, n36268, n36269, n36270, n36271,
    n36272, n36273, n36274, n36275, n36276, n36277,
    n36278, n36279, n36280, n36281, n36282, n36283,
    n36284, n36285, n36286, n36287, n36288, n36289,
    n36290, n36291, n36292, n36293, n36294, n36295,
    n36296, n36297, n36298, n36299, n36300, n36301,
    n36302, n36303, n36304, n36305, n36306, n36307,
    n36308, n36309, n36310, n36311, n36312, n36313,
    n36314, n36315, n36316, n36317, n36318, n36319,
    n36320, n36321, n36322, n36323, n36324, n36325,
    n36326, n36327, n36328, n36329, n36330, n36331,
    n36332, n36333, n36334, n36335, n36336, n36337,
    n36338, n36339, n36340, n36341, n36342, n36343,
    n36344, n36345, n36346, n36347, n36348, n36349,
    n36350, n36351, n36352, n36353, n36354, n36355,
    n36356, n36357, n36358, n36359, n36360, n36361,
    n36362, n36363, n36364, n36365, n36366, n36367,
    n36368, n36369, n36370, n36371, n36372, n36373,
    n36374, n36375, n36376, n36377, n36378, n36379,
    n36380, n36381, n36382, n36383, n36384, n36385,
    n36386, n36387, n36388, n36389, n36390, n36391,
    n36392, n36393, n36394, n36395, n36396, n36397,
    n36398, n36399, n36400, n36401, n36402, n36403,
    n36404, n36405, n36406, n36407, n36408, n36409,
    n36410, n36411, n36412, n36413, n36414, n36415,
    n36416, n36417, n36418, n36419, n36420, n36421,
    n36422, n36423, n36424, n36425, n36426, n36427,
    n36428, n36429, n36430, n36431, n36432, n36433,
    n36434, n36435, n36436, n36437, n36438, n36439,
    n36440, n36441, n36442, n36443, n36444, n36445,
    n36446, n36447, n36448, n36449, n36450, n36451,
    n36452, n36453, n36454, n36455, n36456, n36457,
    n36458, n36459, n36460, n36461, n36462, n36463,
    n36464, n36465, n36466, n36467, n36468, n36469,
    n36470, n36471, n36472, n36473, n36474, n36475,
    n36476, n36477, n36478, n36479, n36480, n36481,
    n36482, n36483, n36484, n36485, n36486, n36487,
    n36488, n36489, n36490, n36491, n36492, n36493,
    n36494, n36495, n36496, n36497, n36498, n36499,
    n36500, n36501, n36502, n36503, n36504, n36505,
    n36506, n36507, n36508, n36509, n36510, n36511,
    n36512, n36513, n36514, n36515, n36516, n36517,
    n36518, n36519, n36520, n36521, n36522, n36523,
    n36524, n36525, n36526, n36527, n36528, n36529,
    n36530, n36531, n36532, n36533, n36534, n36535,
    n36536, n36537, n36538, n36539, n36540, n36541,
    n36542, n36543, n36544, n36545, n36546, n36547,
    n36548, n36549, n36550, n36551, n36552, n36553,
    n36554, n36555, n36556, n36557, n36558, n36559,
    n36560, n36561, n36562, n36563, n36564, n36565,
    n36566, n36567, n36568, n36569, n36570, n36571,
    n36572, n36573, n36574, n36575, n36576, n36577,
    n36578, n36579, n36580, n36581, n36582, n36583,
    n36584, n36585, n36586, n36587, n36588, n36589,
    n36590, n36591, n36592, n36593, n36594, n36595,
    n36596, n36597, n36598, n36599, n36600, n36601,
    n36602, n36603, n36604, n36605, n36606, n36607,
    n36608, n36609, n36610, n36611, n36612, n36613,
    n36614, n36615, n36616, n36617, n36618, n36619,
    n36620, n36621, n36622, n36623, n36624, n36625,
    n36626, n36627, n36628, n36629, n36630, n36631,
    n36632, n36633, n36634, n36635, n36636, n36637,
    n36638, n36639, n36640, n36641, n36642, n36643,
    n36644, n36645, n36646, n36647, n36648, n36649,
    n36650, n36651, n36652, n36653, n36654, n36655,
    n36656, n36657, n36658, n36659, n36660, n36661,
    n36662, n36663, n36664, n36665, n36666, n36667,
    n36668, n36669, n36670, n36671, n36672, n36673,
    n36674, n36675, n36676, n36677, n36678, n36679,
    n36680, n36681, n36682, n36683, n36684, n36685,
    n36686, n36687, n36688, n36689, n36690, n36691,
    n36692, n36693, n36694, n36695, n36696, n36697,
    n36698, n36699, n36700, n36701, n36702, n36703,
    n36704, n36705, n36706, n36707, n36708, n36709,
    n36710, n36711, n36712, n36713, n36714, n36715,
    n36716, n36717, n36718, n36719, n36720, n36721,
    n36722, n36723, n36724, n36725, n36726, n36727,
    n36728, n36729, n36730, n36731, n36732, n36733,
    n36734, n36735, n36736, n36737, n36738, n36739,
    n36740, n36741, n36742, n36743, n36744, n36745,
    n36746, n36747, n36748, n36749, n36750, n36751,
    n36752, n36753, n36754, n36755, n36757, n36758,
    n36759, n36760, n36761, n36762, n36763, n36764,
    n36765, n36766, n36767, n36768, n36769, n36770,
    n36771, n36772, n36773, n36774, n36775, n36776,
    n36777, n36778, n36779, n36780, n36781, n36782,
    n36783, n36784, n36785, n36786, n36787, n36788,
    n36789, n36790, n36791, n36792, n36793, n36794,
    n36795, n36796, n36797, n36798, n36799, n36800,
    n36801, n36802, n36803, n36804, n36805, n36806,
    n36807, n36808, n36809, n36810, n36811, n36812,
    n36813, n36814, n36815, n36816, n36817, n36818,
    n36819, n36820, n36821, n36822, n36823, n36824,
    n36825, n36826, n36827, n36828, n36829, n36830,
    n36831, n36832, n36833, n36834, n36835, n36836,
    n36837, n36838, n36839, n36840, n36841, n36842,
    n36843, n36844, n36845, n36846, n36847, n36848,
    n36849, n36850, n36851, n36852, n36853, n36854,
    n36855, n36856, n36857, n36858, n36859, n36860,
    n36861, n36862, n36863, n36864, n36865, n36866,
    n36867, n36868, n36869, n36870, n36871, n36872,
    n36873, n36874, n36875, n36876, n36877, n36878,
    n36879, n36880, n36881, n36882, n36883, n36884,
    n36885, n36886, n36887, n36888, n36889, n36890,
    n36891, n36892, n36893, n36894, n36895, n36896,
    n36897, n36898, n36899, n36900, n36901, n36902,
    n36903, n36904, n36905, n36906, n36907, n36908,
    n36909, n36910, n36911, n36912, n36913, n36914,
    n36915, n36916, n36917, n36918, n36919, n36920,
    n36921, n36922, n36923, n36924, n36925, n36926,
    n36927, n36928, n36929, n36930, n36931, n36932,
    n36933, n36934, n36935, n36936, n36937, n36938,
    n36939, n36940, n36941, n36942, n36943, n36944,
    n36945, n36946, n36947, n36948, n36949, n36950,
    n36951, n36952, n36953, n36954, n36955, n36956,
    n36957, n36958, n36959, n36960, n36961, n36962,
    n36963, n36964, n36965, n36966, n36967, n36968,
    n36969, n36970, n36971, n36972, n36973, n36974,
    n36975, n36976, n36977, n36978, n36979, n36980,
    n36981, n36982, n36983, n36984, n36985, n36986,
    n36987, n36988, n36989, n36990, n36991, n36992,
    n36993, n36994, n36995, n36996, n36997, n36998,
    n36999, n37000, n37001, n37002, n37003, n37004,
    n37005, n37006, n37007, n37008, n37009, n37010,
    n37011, n37012, n37013, n37014, n37015, n37016,
    n37017, n37018, n37019, n37020, n37021, n37022,
    n37023, n37024, n37025, n37026, n37027, n37028,
    n37029, n37030, n37031, n37032, n37033, n37034,
    n37035, n37036, n37037, n37038, n37039, n37040,
    n37041, n37042, n37043, n37044, n37045, n37046,
    n37047, n37048, n37049, n37050, n37051, n37052,
    n37053, n37054, n37055, n37056, n37057, n37058,
    n37059, n37060, n37061, n37062, n37063, n37064,
    n37065, n37066, n37067, n37068, n37069, n37070,
    n37071, n37072, n37073, n37074, n37075, n37076,
    n37077, n37078, n37079, n37080, n37081, n37082,
    n37083, n37084, n37085, n37086, n37087, n37088,
    n37089, n37090, n37091, n37092, n37093, n37094,
    n37095, n37096, n37097, n37098, n37099, n37100,
    n37101, n37102, n37103, n37104, n37105, n37106,
    n37107, n37108, n37109, n37110, n37111, n37112,
    n37113, n37114, n37115, n37116, n37117, n37118,
    n37119, n37120, n37121, n37122, n37123, n37124,
    n37125, n37126, n37127, n37128, n37129, n37130,
    n37131, n37132, n37133, n37134, n37135, n37136,
    n37137, n37138, n37139, n37140, n37141, n37142,
    n37143, n37144, n37145, n37146, n37147, n37148,
    n37149, n37150, n37151, n37152, n37153, n37154,
    n37155, n37156, n37157, n37158, n37159, n37160,
    n37161, n37162, n37163, n37164, n37165, n37166,
    n37167, n37168, n37169, n37170, n37171, n37172,
    n37173, n37174, n37175, n37176, n37177, n37178,
    n37179, n37180, n37181, n37182, n37183, n37184,
    n37185, n37186, n37187, n37188, n37189, n37190,
    n37191, n37192, n37193, n37194, n37195, n37196,
    n37197, n37198, n37199, n37200, n37201, n37202,
    n37203, n37204, n37205, n37206, n37207, n37208,
    n37209, n37210, n37211, n37212, n37213, n37214,
    n37215, n37216, n37217, n37218, n37219, n37220,
    n37221, n37222, n37223, n37224, n37225, n37226,
    n37227, n37228, n37229, n37230, n37231, n37232,
    n37233, n37234, n37235, n37236, n37237, n37238,
    n37239, n37240, n37241, n37242, n37243, n37244,
    n37245, n37246, n37247, n37248, n37249, n37250,
    n37251, n37252, n37253, n37254, n37255, n37256,
    n37257, n37258, n37259, n37260, n37261, n37262,
    n37263, n37264, n37265, n37266, n37267, n37268,
    n37269, n37270, n37271, n37272, n37273, n37274,
    n37275, n37276, n37277, n37278, n37279, n37280,
    n37281, n37282, n37283, n37284, n37285, n37286,
    n37287, n37288, n37289, n37290, n37291, n37292,
    n37293, n37294, n37295, n37296, n37297, n37298,
    n37299, n37300, n37301, n37302, n37303, n37304,
    n37305, n37306, n37307, n37308, n37309, n37310,
    n37311, n37312, n37313, n37314, n37315, n37316,
    n37317, n37318, n37319, n37320, n37321, n37322,
    n37323, n37324, n37325, n37326, n37327, n37328,
    n37329, n37330, n37331, n37332, n37333, n37334,
    n37335, n37336, n37338, n37339, n37340, n37341,
    n37342, n37343, n37344, n37345, n37346, n37347,
    n37348, n37349, n37350, n37351, n37352, n37353,
    n37354, n37355, n37356, n37357, n37358, n37359,
    n37360, n37361, n37362, n37363, n37364, n37365,
    n37366, n37367, n37368, n37369, n37370, n37371,
    n37372, n37373, n37374, n37375, n37376, n37377,
    n37378, n37379, n37380, n37381, n37382, n37383,
    n37384, n37385, n37386, n37387, n37388, n37389,
    n37390, n37391, n37392, n37393, n37394, n37395,
    n37396, n37397, n37398, n37399, n37400, n37401,
    n37402, n37403, n37404, n37405, n37406, n37407,
    n37408, n37409, n37410, n37411, n37412, n37413,
    n37414, n37415, n37416, n37417, n37418, n37419,
    n37420, n37421, n37422, n37423, n37424, n37425,
    n37426, n37427, n37428, n37429, n37430, n37431,
    n37432, n37433, n37434, n37435, n37436, n37437,
    n37438, n37439, n37440, n37441, n37442, n37443,
    n37444, n37445, n37446, n37447, n37448, n37449,
    n37450, n37451, n37452, n37453, n37454, n37455,
    n37456, n37457, n37458, n37459, n37460, n37461,
    n37462, n37463, n37464, n37465, n37466, n37467,
    n37468, n37469, n37470, n37471, n37472, n37473,
    n37474, n37475, n37476, n37477, n37478, n37479,
    n37480, n37481, n37482, n37483, n37484, n37485,
    n37486, n37487, n37488, n37489, n37490, n37491,
    n37492, n37493, n37494, n37495, n37496, n37497,
    n37498, n37499, n37500, n37501, n37502, n37503,
    n37504, n37505, n37506, n37507, n37508, n37509,
    n37510, n37511, n37512, n37513, n37514, n37515,
    n37516, n37517, n37518, n37519, n37520, n37521,
    n37522, n37523, n37524, n37525, n37526, n37527,
    n37528, n37529, n37530, n37531, n37532, n37533,
    n37534, n37535, n37536, n37537, n37538, n37539,
    n37540, n37541, n37542, n37543, n37544, n37545,
    n37546, n37547, n37548, n37549, n37550, n37551,
    n37552, n37553, n37554, n37555, n37556, n37557,
    n37558, n37559, n37560, n37561, n37562, n37563,
    n37564, n37565, n37566, n37567, n37568, n37569,
    n37570, n37571, n37572, n37573, n37574, n37575,
    n37576, n37577, n37578, n37579, n37580, n37581,
    n37582, n37583, n37584, n37585, n37586, n37587,
    n37588, n37589, n37590, n37591, n37592, n37593,
    n37594, n37595, n37596, n37597, n37598, n37599,
    n37600, n37601, n37602, n37603, n37604, n37605,
    n37606, n37607, n37608, n37609, n37610, n37611,
    n37612, n37613, n37614, n37615, n37616, n37617,
    n37618, n37619, n37620, n37621, n37622, n37623,
    n37624, n37625, n37626, n37627, n37628, n37629,
    n37630, n37631, n37632, n37633, n37634, n37635,
    n37636, n37637, n37638, n37639, n37640, n37641,
    n37642, n37643, n37644, n37645, n37646, n37647,
    n37648, n37649, n37650, n37651, n37652, n37653,
    n37654, n37655, n37656, n37657, n37658, n37659,
    n37660, n37661, n37662, n37663, n37664, n37665,
    n37666, n37667, n37668, n37669, n37670, n37671,
    n37672, n37673, n37674, n37675, n37676, n37677,
    n37678, n37679, n37680, n37681, n37682, n37683,
    n37684, n37685, n37686, n37687, n37688, n37689,
    n37690, n37691, n37692, n37693, n37694, n37695,
    n37696, n37697, n37698, n37699, n37700, n37701,
    n37702, n37703, n37704, n37705, n37706, n37707,
    n37708, n37709, n37710, n37711, n37712, n37713,
    n37714, n37715, n37716, n37717, n37718, n37719,
    n37720, n37721, n37722, n37723, n37724, n37725,
    n37726, n37727, n37728, n37729, n37730, n37731,
    n37732, n37733, n37734, n37735, n37736, n37737,
    n37738, n37739, n37740, n37741, n37742, n37743,
    n37744, n37745, n37746, n37747, n37748, n37749,
    n37750, n37751, n37752, n37753, n37754, n37755,
    n37756, n37757, n37758, n37759, n37760, n37761,
    n37762, n37763, n37764, n37765, n37766, n37767,
    n37768, n37769, n37770, n37771, n37772, n37773,
    n37774, n37775, n37776, n37777, n37778, n37779,
    n37780, n37781, n37782, n37783, n37784, n37785,
    n37786, n37787, n37788, n37789, n37790, n37791,
    n37792, n37793, n37794, n37795, n37796, n37797,
    n37798, n37799, n37800, n37801, n37802, n37803,
    n37804, n37805, n37806, n37807, n37808, n37809,
    n37810, n37811, n37812, n37813, n37814, n37815,
    n37816, n37817, n37818, n37819, n37820, n37821,
    n37822, n37823, n37824, n37825, n37826, n37827,
    n37828, n37829, n37830, n37831, n37832, n37833,
    n37834, n37835, n37836, n37837, n37838, n37839,
    n37840, n37841, n37842, n37843, n37844, n37845,
    n37846, n37847, n37848, n37849, n37850, n37851,
    n37852, n37853, n37854, n37855, n37856, n37857,
    n37858, n37859, n37860, n37861, n37862, n37863,
    n37864, n37865, n37866, n37867, n37868, n37869,
    n37870, n37871, n37872, n37873, n37874, n37875,
    n37876, n37877, n37878, n37879, n37880, n37881,
    n37882, n37883, n37884, n37885, n37886, n37887,
    n37888, n37889, n37890, n37891, n37892, n37893,
    n37894, n37895, n37896, n37897, n37898, n37899,
    n37900, n37901, n37902, n37903, n37904, n37905,
    n37906, n37907, n37908, n37909, n37910, n37911,
    n37912, n37913, n37914, n37915, n37916, n37917,
    n37918, n37919, n37920, n37921, n37922, n37923,
    n37925, n37926, n37927, n37928, n37929, n37930,
    n37931, n37932, n37933, n37934, n37935, n37936,
    n37937, n37938, n37939, n37940, n37941, n37942,
    n37943, n37944, n37945, n37946, n37947, n37948,
    n37949, n37950, n37951, n37952, n37953, n37954,
    n37955, n37956, n37957, n37958, n37959, n37960,
    n37961, n37962, n37963, n37964, n37965, n37966,
    n37967, n37968, n37969, n37970, n37971, n37972,
    n37973, n37974, n37975, n37976, n37977, n37978,
    n37979, n37980, n37981, n37982, n37983, n37984,
    n37985, n37986, n37987, n37988, n37989, n37990,
    n37991, n37992, n37993, n37994, n37995, n37996,
    n37997, n37998, n37999, n38000, n38001, n38002,
    n38003, n38004, n38005, n38006, n38007, n38008,
    n38009, n38010, n38011, n38012, n38013, n38014,
    n38015, n38016, n38017, n38018, n38019, n38020,
    n38021, n38022, n38023, n38024, n38025, n38026,
    n38027, n38028, n38029, n38030, n38031, n38032,
    n38033, n38034, n38035, n38036, n38037, n38038,
    n38039, n38040, n38041, n38042, n38043, n38044,
    n38045, n38046, n38047, n38048, n38050, n38051,
    n38052, n38053, n38054, n38055, n38056, n38057,
    n38058, n38059, n38060, n38061, n38062, n38063,
    n38064, n38065, n38066, n38067, n38068, n38069,
    n38070, n38071, n38072, n38073, n38074, n38075,
    n38076, n38077, n38078, n38079, n38080, n38081,
    n38082, n38083, n38084, n38085, n38086, n38087,
    n38088, n38089, n38090, n38091, n38092, n38093,
    n38094, n38095, n38096, n38097, n38098, n38099,
    n38100, n38101, n38103, n38104, n38105, n38106,
    n38107, n38108, n38109, n38110, n38111, n38112,
    n38113, n38114, n38115, n38116, n38117, n38118,
    n38119, n38120, n38121, n38122, n38123, n38124,
    n38125, n38126, n38127, n38128, n38129, n38130,
    n38131, n38132, n38134, n38135, n38136, n38137,
    n38138, n38139, n38140, n38141, n38142, n38143,
    n38144, n38146, n38147, n38148, n38149, n38150,
    n38151, n38152, n38153, n38154, n38155, n38156,
    n38157, n38158, n38159, n38160, n38161, n38162,
    n38163, n38164, n38165, n38166, n38167, n38168,
    n38169, n38170, n38171, n38172, n38173, n38174,
    n38175, n38176, n38177, n38178, n38179, n38180,
    n38181, n38182, n38183, n38184, n38185, n38186,
    n38187, n38188, n38189, n38190, n38191, n38192,
    n38193, n38194, n38195, n38196, n38197, n38198,
    n38199, n38200, n38201, n38202, n38203, n38204,
    n38205, n38206, n38207, n38208, n38209, n38210,
    n38211, n38212, n38213, n38214, n38215, n38216,
    n38217, n38218, n38219, n38220, n38221, n38222,
    n38223, n38224, n38225, n38226, n38227, n38229,
    n38230, n38231, n38232, n38233, n38234, n38235,
    n38236, n38237, n38238, n38239, n38240, n38241,
    n38242, n38243, n38244, n38245, n38246, n38247,
    n38248, n38249, n38250, n38251, n38252, n38253,
    n38254, n38255, n38256, n38257, n38258, n38259,
    n38260, n38261, n38262, n38263, n38264, n38266,
    n38267, n38268, n38269, n38270, n38271, n38272,
    n38273, n38274, n38275, n38276, n38277, n38278,
    n38279, n38280, n38281, n38282, n38283, n38284,
    n38285, n38286, n38287, n38289, n38290, n38291,
    n38292, n38293, n38294, n38295, n38296, n38297,
    n38298, n38299, n38300, n38301, n38302, n38303,
    n38304, n38305, n38306, n38307, n38308, n38309,
    n38310, n38311, n38312, n38313, n38314, n38315,
    n38316, n38317, n38318, n38319, n38320, n38321,
    n38322, n38323, n38324, n38325, n38326, n38327,
    n38328, n38329, n38330, n38331, n38332, n38333,
    n38334, n38335, n38336, n38337, n38338, n38339,
    n38340, n38341, n38342, n38343, n38344, n38345,
    n38346, n38347, n38348, n38349, n38350, n38351,
    n38352, n38353, n38354, n38355, n38356, n38357,
    n38358, n38359, n38360, n38361, n38362, n38363,
    n38364, n38365, n38366, n38367, n38368, n38369,
    n38370, n38371, n38372, n38373, n38374, n38375,
    n38376, n38377, n38378, n38379, n38380, n38381,
    n38382, n38383, n38384, n38385, n38386, n38387,
    n38388, n38389, n38390, n38391, n38392, n38393,
    n38394, n38395, n38396, n38397, n38398, n38399,
    n38400, n38401, n38402, n38403, n38404, n38405,
    n38406, n38407, n38408, n38409, n38410, n38411,
    n38412, n38413, n38414, n38415, n38416, n38417,
    n38418, n38419, n38420, n38421, n38422, n38423,
    n38424, n38425, n38426, n38427, n38428, n38429,
    n38430, n38431, n38432, n38433, n38434, n38435,
    n38436, n38437, n38438, n38439, n38440, n38441,
    n38442, n38443, n38444, n38445, n38446, n38447,
    n38448, n38449, n38450, n38451, n38452, n38453,
    n38454, n38455, n38456, n38457, n38458, n38459,
    n38460, n38461, n38462, n38463, n38464, n38465,
    n38466, n38467, n38468, n38469, n38470, n38471,
    n38472, n38473, n38474, n38475, n38476, n38477,
    n38478, n38479, n38480, n38481, n38482, n38483,
    n38484, n38485, n38486, n38487, n38488, n38489,
    n38490, n38491, n38492, n38493, n38494, n38495,
    n38496, n38497, n38498, n38499, n38500, n38501,
    n38502, n38503, n38504, n38505, n38506, n38507,
    n38508, n38509, n38510, n38511, n38512, n38513,
    n38514, n38515, n38516, n38517, n38518, n38519,
    n38520, n38521, n38522, n38523, n38524, n38525,
    n38526, n38527, n38528, n38529, n38530, n38531,
    n38532, n38533, n38534, n38535, n38536, n38537,
    n38538, n38539, n38540, n38541, n38542, n38543,
    n38544, n38545, n38546, n38547, n38548, n38549,
    n38550, n38551, n38552, n38553, n38554, n38555,
    n38556, n38557, n38558, n38559, n38560, n38561,
    n38562, n38563, n38564, n38565, n38566, n38567,
    n38568, n38569, n38570, n38571, n38572, n38573,
    n38574, n38575, n38576, n38577, n38578, n38579,
    n38580, n38581, n38582, n38583, n38584, n38585,
    n38586, n38587, n38588, n38589, n38590, n38591,
    n38592, n38593, n38594, n38595, n38596, n38597,
    n38598, n38599, n38600, n38601, n38602, n38603,
    n38604, n38605, n38606, n38607, n38608, n38609,
    n38610, n38611, n38612, n38613, n38614, n38615,
    n38616, n38617, n38618, n38619, n38620, n38621,
    n38622, n38623, n38624, n38625, n38626, n38627,
    n38628, n38629, n38630, n38631, n38632, n38633,
    n38634, n38635, n38636, n38637, n38638, n38639,
    n38640, n38641, n38642, n38643, n38644, n38645,
    n38646, n38647, n38648, n38649, n38650, n38651,
    n38652, n38653, n38654, n38655, n38656, n38657,
    n38658, n38659, n38660, n38661, n38662, n38663,
    n38664, n38665, n38666, n38667, n38668, n38669,
    n38670, n38671, n38672, n38673, n38674, n38675,
    n38676, n38677, n38678, n38679, n38680, n38681,
    n38682, n38683, n38684, n38685, n38686, n38687,
    n38688, n38689, n38690, n38691, n38692, n38693,
    n38694, n38695, n38696, n38697, n38699, n38700,
    n38701, n38702, n38703, n38704, n38705, n38706,
    n38707, n38708, n38709, n38710, n38711, n38712,
    n38713, n38714, n38715, n38716, n38717, n38718,
    n38719, n38720, n38721, n38722, n38723, n38724,
    n38725, n38726, n38727, n38728, n38729, n38730,
    n38731, n38732, n38733, n38734, n38735, n38736,
    n38737, n38738, n38739, n38740, n38741, n38742,
    n38743, n38744, n38745, n38746, n38747, n38748,
    n38749, n38750, n38751, n38752, n38753, n38754,
    n38755, n38756, n38757, n38758, n38759, n38760,
    n38761, n38762, n38763, n38764, n38765, n38766,
    n38767, n38768, n38769, n38770, n38771, n38772,
    n38773, n38774, n38775, n38776, n38777, n38778,
    n38779, n38780, n38781, n38782, n38783, n38784,
    n38785, n38786, n38787, n38788, n38789, n38790,
    n38791, n38792, n38793, n38794, n38795, n38796,
    n38797, n38798, n38799, n38800, n38801, n38802,
    n38803, n38804, n38805, n38806, n38807, n38808,
    n38809, n38810, n38811, n38812, n38813, n38814,
    n38815, n38816, n38817, n38818, n38819, n38820,
    n38821, n38822, n38823, n38824, n38825, n38826,
    n38827, n38828, n38829, n38830, n38831, n38832,
    n38833, n38834, n38835, n38836, n38837, n38838,
    n38839, n38840, n38841, n38842, n38843, n38844,
    n38845, n38846, n38847, n38848, n38849, n38850,
    n38851, n38852, n38853, n38854, n38855, n38856,
    n38857, n38858, n38859, n38860, n38861, n38862,
    n38863, n38864, n38865, n38866, n38867, n38868,
    n38869, n38870, n38871, n38872, n38873, n38874,
    n38875, n38876, n38877, n38878, n38879, n38880,
    n38881, n38882, n38883, n38884, n38885, n38886,
    n38887, n38888, n38889, n38890, n38891, n38892,
    n38893, n38894, n38895, n38896, n38897, n38898,
    n38899, n38900, n38901, n38902, n38903, n38904,
    n38905, n38906, n38907, n38908, n38909, n38910,
    n38911, n38912, n38913, n38914, n38915, n38916,
    n38917, n38918, n38919, n38920, n38921, n38922,
    n38923, n38924, n38925, n38926, n38927, n38928,
    n38929, n38930, n38931, n38932, n38933, n38934,
    n38935, n38936, n38937, n38938, n38939, n38940,
    n38941, n38942, n38943, n38944, n38945, n38946,
    n38947, n38948, n38949, n38950, n38951, n38952,
    n38953, n38954, n38955, n38956, n38957, n38958,
    n38959, n38960, n38961, n38962, n38963, n38964,
    n38965, n38966, n38967, n38968, n38969, n38970,
    n38971, n38972, n38973, n38974, n38975, n38976,
    n38977, n38978, n38979, n38980, n38981, n38982,
    n38983, n38984, n38985, n38986, n38987, n38988,
    n38989, n38990, n38991, n38992, n38993, n38994,
    n38995, n38996, n38997, n38998, n38999, n39000,
    n39001, n39002, n39003, n39004, n39005, n39006,
    n39007, n39008, n39009, n39010, n39011, n39012,
    n39013, n39014, n39015, n39016, n39017, n39018,
    n39019, n39020, n39021, n39022, n39023, n39025,
    n39026, n39027, n39028, n39029, n39030, n39031,
    n39032, n39033, n39034, n39035, n39036, n39037,
    n39038, n39039, n39040, n39041, n39042, n39043,
    n39044, n39045, n39046, n39047, n39048, n39049,
    n39050, n39051, n39052, n39053, n39054, n39055,
    n39056, n39057, n39058, n39059, n39060, n39061,
    n39062, n39063, n39064, n39065, n39066, n39067,
    n39068, n39069, n39070, n39071, n39072, n39073,
    n39074, n39075, n39076, n39077, n39078, n39079,
    n39080, n39081, n39082, n39083, n39084, n39085,
    n39086, n39087, n39088, n39089, n39090, n39091,
    n39092, n39093, n39094, n39095, n39096, n39097,
    n39098, n39099, n39100, n39101, n39102, n39103,
    n39104, n39105, n39106, n39107, n39108, n39109,
    n39110, n39111, n39112, n39113, n39114, n39115,
    n39116, n39117, n39118, n39119, n39120, n39121,
    n39122, n39123, n39124, n39125, n39126, n39127,
    n39128, n39129, n39130, n39131, n39132, n39133,
    n39134, n39135, n39136, n39137, n39138, n39139,
    n39140, n39141, n39142, n39143, n39144, n39145,
    n39146, n39147, n39148, n39149, n39150, n39151,
    n39152, n39153, n39154, n39155, n39156, n39157,
    n39158, n39159, n39160, n39161, n39162, n39163,
    n39164, n39165, n39166, n39167, n39168, n39169,
    n39170, n39171, n39172, n39173, n39174, n39175,
    n39176, n39177, n39178, n39179, n39180, n39181,
    n39182, n39183, n39184, n39185, n39186, n39187,
    n39188, n39189, n39190, n39191, n39192, n39193,
    n39194, n39195, n39196, n39197, n39198, n39199,
    n39200, n39201, n39202, n39203, n39204, n39205,
    n39206, n39207, n39208, n39209, n39210, n39211,
    n39212, n39213, n39214, n39215, n39216, n39217,
    n39218, n39219, n39220, n39222, n39223, n39224,
    n39225, n39226, n39227, n39228, n39229, n39230,
    n39231, n39232, n39233, n39235, n39236, n39237,
    n39238, n39239, n39240, n39241, n39242, n39243,
    n39244, n39245, n39246, n39247, n39248, n39249,
    n39250, n39251, n39252, n39253, n39254, n39255,
    n39256, n39257, n39258, n39259, n39260, n39261,
    n39262, n39263, n39264, n39265, n39266, n39267,
    n39268, n39269, n39270, n39271, n39272, n39273,
    n39274, n39275, n39276, n39277, n39278, n39279,
    n39280, n39281, n39282, n39283, n39284, n39285,
    n39286, n39287, n39288, n39289, n39290, n39291,
    n39292, n39293, n39294, n39295, n39296, n39297,
    n39298, n39299, n39300, n39301, n39302, n39303,
    n39304, n39305, n39306, n39307, n39308, n39309,
    n39310, n39311, n39312, n39313, n39314, n39315,
    n39316, n39317, n39318, n39319, n39320, n39321,
    n39322, n39323, n39324, n39325, n39326, n39327,
    n39328, n39329, n39330, n39331, n39332, n39333,
    n39334, n39335, n39336, n39337, n39338, n39339,
    n39340, n39341, n39342, n39343, n39344, n39345,
    n39346, n39347, n39348, n39349, n39350, n39351,
    n39352, n39353, n39354, n39355, n39356, n39357,
    n39358, n39359, n39360, n39361, n39362, n39363,
    n39364, n39365, n39366, n39367, n39368, n39369,
    n39370, n39371, n39372, n39373, n39374, n39375,
    n39376, n39377, n39378, n39379, n39380, n39381,
    n39382, n39383, n39384, n39385, n39386, n39387,
    n39388, n39389, n39390, n39391, n39392, n39393,
    n39394, n39395, n39396, n39397, n39398, n39399,
    n39400, n39401, n39402, n39403, n39404, n39405,
    n39406, n39407, n39408, n39409, n39410, n39411,
    n39412, n39413, n39414, n39415, n39416, n39417,
    n39418, n39419, n39420, n39421, n39422, n39423,
    n39424, n39425, n39426, n39427, n39428, n39429,
    n39430, n39431, n39432, n39433, n39434, n39435,
    n39436, n39437, n39438, n39439, n39440, n39441,
    n39442, n39443, n39444, n39445, n39446, n39447,
    n39448, n39449, n39450, n39451, n39452, n39453,
    n39454, n39455, n39456, n39457, n39458, n39459,
    n39460, n39461, n39462, n39463, n39464, n39465,
    n39466, n39467, n39468, n39469, n39470, n39471,
    n39472, n39473, n39474, n39475, n39476, n39477,
    n39478, n39479, n39480, n39481, n39482, n39483,
    n39484, n39485, n39486, n39487, n39488, n39489,
    n39490, n39491, n39492, n39493, n39494, n39495,
    n39496, n39498, n39499, n39500, n39501, n39502,
    n39503, n39504, n39505, n39506, n39507, n39508,
    n39509, n39510, n39511, n39512, n39513, n39514,
    n39515, n39516, n39517, n39518, n39519, n39520,
    n39521, n39522, n39523, n39524, n39525, n39526,
    n39527, n39528, n39529, n39530, n39531, n39532,
    n39533, n39534, n39535, n39536, n39537, n39538,
    n39539, n39540, n39541, n39542, n39543, n39544,
    n39545, n39546, n39547, n39548, n39549, n39550,
    n39551, n39552, n39553, n39554, n39555, n39556,
    n39557, n39558, n39559, n39560, n39561, n39562,
    n39563, n39564, n39565, n39566, n39567, n39568,
    n39569, n39570, n39571, n39572, n39573, n39574,
    n39575, n39576, n39577, n39578, n39579, n39580,
    n39581, n39582, n39583, n39584, n39585, n39586,
    n39587, n39588, n39589, n39590, n39591, n39592,
    n39593, n39594, n39595, n39596, n39597, n39598,
    n39599, n39600, n39601, n39602, n39603, n39604,
    n39605, n39606, n39607, n39608, n39609, n39610,
    n39611, n39612, n39613, n39614, n39615, n39616,
    n39617, n39618, n39619, n39620, n39621, n39622,
    n39623, n39624, n39625, n39626, n39627, n39628,
    n39629, n39630, n39631, n39632, n39633, n39634,
    n39635, n39636, n39637, n39638, n39639, n39640,
    n39641, n39642, n39643, n39644, n39645, n39646,
    n39647, n39648, n39649, n39650, n39651, n39652,
    n39653, n39654, n39655, n39656, n39657, n39658,
    n39659, n39660, n39661, n39662, n39663, n39664,
    n39665, n39666, n39667, n39668, n39669, n39670,
    n39671, n39672, n39673, n39674, n39675, n39676,
    n39677, n39678, n39679, n39680, n39681, n39682,
    n39683, n39684, n39685, n39686, n39687, n39688,
    n39689, n39690, n39691, n39692, n39693, n39694,
    n39695, n39696, n39697, n39698, n39699, n39700,
    n39701, n39702, n39703, n39704, n39705, n39706,
    n39707, n39708, n39709, n39710, n39711, n39712,
    n39713, n39714, n39715, n39716, n39717, n39718,
    n39719, n39720, n39721, n39722, n39723, n39724,
    n39725, n39726, n39727, n39728, n39729, n39730,
    n39731, n39732, n39733, n39734, n39735, n39736,
    n39737, n39738, n39739, n39740, n39741, n39742,
    n39743, n39744, n39745, n39746, n39747, n39748,
    n39749, n39750, n39751, n39752, n39753, n39754,
    n39755, n39756, n39757, n39758, n39759, n39760,
    n39761, n39762, n39763, n39764, n39765, n39766,
    n39767, n39768, n39769, n39770, n39771, n39772,
    n39773, n39774, n39775, n39776, n39777, n39778,
    n39779, n39780, n39781, n39782, n39783, n39784,
    n39785, n39786, n39787, n39788, n39789, n39790,
    n39791, n39792, n39793, n39794, n39795, n39796,
    n39797, n39798, n39799, n39800, n39801, n39802,
    n39803, n39804, n39805, n39806, n39807, n39808,
    n39809, n39810, n39811, n39812, n39813, n39814,
    n39815, n39816, n39817, n39818, n39819, n39820,
    n39821, n39822, n39823, n39824, n39825, n39827,
    n39828, n39829, n39830, n39831, n39832, n39833,
    n39834, n39835, n39836, n39837, n39838, n39839,
    n39840, n39841, n39842, n39843, n39844, n39845,
    n39846, n39847, n39848, n39849, n39850, n39851,
    n39852, n39853, n39854, n39855, n39856, n39857,
    n39858, n39859, n39860, n39861, n39862, n39863,
    n39864, n39865, n39866, n39867, n39868, n39869,
    n39870, n39871, n39872, n39873, n39874, n39875,
    n39876, n39877, n39878, n39879, n39880, n39881,
    n39882, n39883, n39884, n39885, n39886, n39887,
    n39888, n39889, n39890, n39891, n39892, n39893,
    n39894, n39895, n39896, n39897, n39898, n39899,
    n39900, n39901, n39902, n39903, n39904, n39905,
    n39906, n39907, n39908, n39909, n39910, n39911,
    n39912, n39913, n39914, n39915, n39916, n39918,
    n39919, n39920, n39921, n39922, n39923, n39924,
    n39925, n39926, n39927, n39928, n39929, n39930,
    n39931, n39932, n39933, n39934, n39935, n39936,
    n39937, n39938, n39939, n39940, n39941, n39942,
    n39943, n39944, n39945, n39946, n39947, n39948,
    n39949, n39950, n39951, n39952, n39953, n39954,
    n39955, n39956, n39957, n39958, n39959, n39960,
    n39961, n39962, n39963, n39964, n39965, n39966,
    n39967, n39968, n39969, n39970, n39971, n39972,
    n39973, n39974, n39975, n39976, n39977, n39978,
    n39979, n39980, n39981, n39982, n39983, n39984,
    n39985, n39986, n39987, n39988, n39989, n39990,
    n39991, n39992, n39993, n39994, n39995, n39996,
    n39997, n39998, n39999, n40000, n40001, n40002,
    n40003, n40004, n40005, n40006, n40007, n40008,
    n40009, n40010, n40011, n40012, n40013, n40014,
    n40015, n40016, n40017, n40018, n40019, n40020,
    n40021, n40022, n40023, n40024, n40025, n40026,
    n40027, n40028, n40029, n40030, n40031, n40032,
    n40033, n40034, n40035, n40036, n40037, n40038,
    n40039, n40040, n40041, n40042, n40043, n40044,
    n40045, n40046, n40047, n40048, n40049, n40050,
    n40051, n40052, n40053, n40054, n40055, n40056,
    n40057, n40058, n40059, n40060, n40061, n40062,
    n40063, n40064, n40065, n40066, n40067, n40068,
    n40069, n40070, n40071, n40072, n40073, n40074,
    n40075, n40076, n40077, n40078, n40079, n40080,
    n40081, n40082, n40083, n40084, n40085, n40086,
    n40087, n40088, n40089, n40090, n40091, n40092,
    n40093, n40094, n40095, n40096, n40097, n40098,
    n40099, n40100, n40101, n40102, n40103, n40104,
    n40105, n40106, n40107, n40108, n40109, n40110,
    n40111, n40112, n40113, n40114, n40115, n40116,
    n40117, n40118, n40119, n40120, n40121, n40122,
    n40123, n40124, n40125, n40126, n40127, n40128,
    n40129, n40130, n40131, n40132, n40133, n40134,
    n40135, n40136, n40137, n40138, n40139, n40140,
    n40141, n40142, n40143, n40144, n40145, n40146,
    n40147, n40148, n40149, n40150, n40151, n40152,
    n40153, n40154, n40155, n40156, n40157, n40158,
    n40159, n40160, n40161, n40162, n40163, n40164,
    n40165, n40166, n40167, n40168, n40169, n40170,
    n40171, n40172, n40173, n40174, n40175, n40176,
    n40177, n40178, n40179, n40180, n40181, n40182,
    n40183, n40184, n40185, n40186, n40187, n40188,
    n40189, n40190, n40191, n40192, n40193, n40194,
    n40195, n40196, n40197, n40198, n40199, n40200,
    n40201, n40202, n40203, n40204, n40205, n40206,
    n40207, n40208, n40209, n40210, n40211, n40212,
    n40213, n40214, n40215, n40216, n40217, n40218,
    n40219, n40220, n40221, n40222, n40223, n40224,
    n40225, n40226, n40227, n40228, n40229, n40230,
    n40231, n40232, n40233, n40234, n40235, n40236,
    n40237, n40238, n40239, n40240, n40241, n40242,
    n40243, n40244, n40245, n40246, n40247, n40248,
    n40249, n40250, n40251, n40252, n40253, n40254,
    n40255, n40256, n40257, n40258, n40259, n40260,
    n40261, n40262, n40263, n40264, n40265, n40266,
    n40267, n40268, n40269, n40270, n40271, n40272,
    n40273, n40274, n40275, n40276, n40277, n40278,
    n40279, n40280, n40281, n40282, n40283, n40284,
    n40285, n40286, n40287, n40288, n40289, n40290,
    n40291, n40292, n40293, n40294, n40295, n40296,
    n40297, n40298, n40299, n40300, n40301, n40302,
    n40303, n40304, n40305, n40306, n40307, n40308,
    n40309, n40310, n40311, n40312, n40313, n40314,
    n40315, n40316, n40317, n40318, n40319, n40320,
    n40321, n40322, n40323, n40324, n40325, n40326,
    n40327, n40328, n40329, n40331, n40332, n40333,
    n40334, n40335, n40336, n40337, n40338, n40339,
    n40340, n40341, n40342, n40343, n40344, n40345,
    n40346, n40347, n40348, n40349, n40350, n40351,
    n40352, n40353, n40354, n40355, n40356, n40357,
    n40358, n40359, n40360, n40361, n40362, n40363,
    n40364, n40365, n40366, n40367, n40368, n40369,
    n40370, n40371, n40372, n40373, n40374, n40375,
    n40376, n40377, n40378, n40379, n40380, n40381,
    n40382, n40383, n40384, n40385, n40386, n40387,
    n40388, n40389, n40390, n40391, n40392, n40393,
    n40394, n40395, n40396, n40397, n40398, n40399,
    n40400, n40401, n40402, n40403, n40404, n40405,
    n40406, n40407, n40408, n40409, n40410, n40411,
    n40412, n40413, n40414, n40415, n40416, n40417,
    n40418, n40419, n40420, n40421, n40422, n40423,
    n40424, n40425, n40426, n40427, n40428, n40429,
    n40430, n40431, n40432, n40433, n40434, n40435,
    n40436, n40437, n40438, n40439, n40440, n40441,
    n40442, n40443, n40444, n40445, n40446, n40447,
    n40448, n40449, n40450, n40451, n40452, n40453,
    n40454, n40455, n40456, n40457, n40458, n40459,
    n40460, n40461, n40462, n40463, n40464, n40465,
    n40466, n40467, n40468, n40469, n40470, n40471,
    n40472, n40473, n40474, n40475, n40476, n40477,
    n40478, n40479, n40480, n40481, n40482, n40483,
    n40484, n40485, n40486, n40487, n40488, n40489,
    n40490, n40491, n40492, n40493, n40494, n40495,
    n40496, n40497, n40498, n40499, n40500, n40501,
    n40502, n40503, n40504, n40505, n40506, n40507,
    n40508, n40509, n40510, n40511, n40512, n40513,
    n40514, n40515, n40516, n40517, n40518, n40519,
    n40520, n40521, n40522, n40523, n40524, n40525,
    n40526, n40527, n40528, n40529, n40530, n40531,
    n40532, n40533, n40534, n40535, n40536, n40537,
    n40538, n40539, n40540, n40541, n40542, n40543,
    n40544, n40545, n40546, n40547, n40548, n40549,
    n40550, n40551, n40552, n40553, n40554, n40555,
    n40556, n40557, n40558, n40559, n40560, n40561,
    n40562, n40563, n40564, n40565, n40566, n40567,
    n40568, n40569, n40570, n40571, n40572, n40573,
    n40574, n40575, n40576, n40577, n40578, n40579,
    n40580, n40581, n40582, n40583, n40584, n40585,
    n40586, n40587, n40588, n40589, n40590, n40591,
    n40592, n40593, n40594, n40595, n40596, n40597,
    n40598, n40599, n40600, n40601, n40602, n40603,
    n40604, n40605, n40606, n40607, n40608, n40609,
    n40610, n40611, n40612, n40613, n40614, n40615,
    n40616, n40617, n40618, n40620, n40621, n40622,
    n40623, n40624, n40625, n40626, n40627, n40628,
    n40629, n40630, n40631, n40632, n40633, n40634,
    n40635, n40636, n40637, n40638, n40639, n40640,
    n40641, n40642, n40643, n40644, n40645, n40646,
    n40647, n40648, n40649, n40650, n40651, n40652,
    n40653, n40654, n40655, n40656, n40657, n40658,
    n40659, n40660, n40661, n40662, n40663, n40664,
    n40665, n40666, n40667, n40668, n40669, n40670,
    n40671, n40672, n40673, n40674, n40675, n40676,
    n40677, n40678, n40679, n40680, n40681, n40682,
    n40683, n40684, n40685, n40686, n40687, n40688,
    n40689, n40690, n40691, n40692, n40693, n40694,
    n40695, n40696, n40697, n40698, n40699, n40700,
    n40701, n40702, n40704, n40705, n40706, n40707,
    n40708, n40709, n40710, n40711, n40712, n40713,
    n40714, n40715, n40716, n40717, n40718, n40719,
    n40720, n40721, n40722, n40723, n40724, n40725,
    n40726, n40727, n40728, n40729, n40730, n40731,
    n40732, n40733, n40734, n40735, n40736, n40737,
    n40738, n40739, n40740, n40741, n40742, n40743,
    n40744, n40745, n40746, n40747, n40748, n40749,
    n40750, n40751, n40752, n40753, n40754, n40755,
    n40756, n40757, n40758, n40759, n40760, n40761,
    n40762, n40763, n40764, n40765, n40766, n40767,
    n40768, n40769, n40770, n40771, n40772, n40773,
    n40774, n40775, n40776, n40777, n40778, n40779,
    n40780, n40781, n40782, n40783, n40784, n40785,
    n40786, n40787, n40788, n40789, n40790, n40791,
    n40792, n40793, n40794, n40795, n40796, n40797,
    n40798, n40799, n40800, n40801, n40802, n40803,
    n40804, n40805, n40806, n40807, n40808, n40809,
    n40810, n40811, n40812, n40813, n40814, n40815,
    n40816, n40817, n40818, n40819, n40820, n40821,
    n40822, n40823, n40824, n40825, n40826, n40827,
    n40828, n40829, n40830, n40831, n40832, n40833,
    n40834, n40835, n40836, n40837, n40838, n40839,
    n40840, n40841, n40842, n40843, n40844, n40845,
    n40846, n40847, n40848, n40849, n40850, n40851,
    n40852, n40853, n40854, n40855, n40856, n40857,
    n40858, n40859, n40860, n40861, n40862, n40863,
    n40864, n40865, n40866, n40867, n40868, n40869,
    n40870, n40871, n40872, n40873, n40874, n40875,
    n40876, n40877, n40878, n40879, n40880, n40881,
    n40882, n40883, n40884, n40885, n40886, n40887,
    n40888, n40889, n40890, n40891, n40892, n40893,
    n40894, n40895, n40896, n40897, n40898, n40899,
    n40900, n40901, n40902, n40903, n40904, n40905,
    n40906, n40907, n40908, n40909, n40910, n40911,
    n40912, n40913, n40914, n40915, n40916, n40917,
    n40918, n40919, n40920, n40921, n40922, n40923,
    n40924, n40925, n40926, n40927, n40928, n40929,
    n40930, n40931, n40932, n40933, n40934, n40935,
    n40936, n40937, n40938, n40939, n40940, n40941,
    n40942, n40943, n40944, n40945, n40946, n40947,
    n40948, n40949, n40950, n40951, n40952, n40953,
    n40954, n40955, n40956, n40957, n40958, n40959,
    n40960, n40961, n40962, n40963, n40964, n40965,
    n40966, n40967, n40968, n40969, n40970, n40971,
    n40972, n40973, n40974, n40975, n40976, n40977,
    n40978, n40979, n40980, n40981, n40982, n40983,
    n40984, n40985, n40986, n40987, n40988, n40989,
    n40990, n40991, n40992, n40993, n40994, n40995,
    n40996, n40997, n40998, n40999, n41000, n41001,
    n41002, n41003, n41004, n41005, n41006, n41007,
    n41008, n41009, n41010, n41011, n41012, n41014,
    n41015, n41016, n41017, n41018, n41019, n41020,
    n41021, n41022, n41023, n41024, n41025, n41026,
    n41027, n41028, n41029, n41030, n41031, n41032,
    n41033, n41034, n41035, n41036, n41037, n41038,
    n41039, n41040, n41041, n41042, n41043, n41044,
    n41045, n41046, n41047, n41048, n41049, n41050,
    n41051, n41052, n41053, n41054, n41055, n41056,
    n41057, n41058, n41059, n41060, n41061, n41062,
    n41063, n41064, n41065, n41067, n41068, n41069,
    n41070, n41071, n41072, n41073, n41074, n41075,
    n41076, n41077, n41078, n41079, n41080, n41081,
    n41082, n41083, n41084, n41085, n41086, n41087,
    n41088, n41089, n41090, n41091, n41092, n41093,
    n41094, n41095, n41096, n41097, n41098, n41099,
    n41100, n41101, n41102, n41103, n41104, n41105,
    n41106, n41107, n41108, n41109, n41110, n41111,
    n41112, n41113, n41114, n41115, n41116, n41117,
    n41118, n41119, n41120, n41121, n41122, n41123,
    n41124, n41125, n41126, n41127, n41128, n41129,
    n41130, n41131, n41132, n41133, n41134, n41135,
    n41136, n41137, n41138, n41139, n41140, n41141,
    n41142, n41143, n41144, n41145, n41146, n41147,
    n41148, n41149, n41150, n41151, n41152, n41153,
    n41154, n41155, n41156, n41157, n41158, n41159,
    n41160, n41161, n41162, n41163, n41164, n41165,
    n41166, n41167, n41168, n41169, n41170, n41171,
    n41172, n41173, n41174, n41175, n41176, n41177,
    n41178, n41179, n41180, n41181, n41182, n41183,
    n41184, n41185, n41186, n41187, n41188, n41189,
    n41190, n41191, n41192, n41193, n41194, n41195,
    n41196, n41197, n41198, n41199, n41200, n41201,
    n41202, n41203, n41204, n41205, n41206, n41207,
    n41208, n41209, n41210, n41211, n41212, n41213,
    n41214, n41215, n41216, n41217, n41218, n41219,
    n41220, n41221, n41222, n41223, n41224, n41225,
    n41226, n41227, n41228, n41229, n41230, n41231,
    n41232, n41233, n41234, n41235, n41236, n41237,
    n41238, n41239, n41240, n41241, n41242, n41243,
    n41244, n41245, n41246, n41247, n41248, n41249,
    n41250, n41251, n41252, n41253, n41254, n41255,
    n41256, n41257, n41258, n41259, n41260, n41261,
    n41262, n41263, n41264, n41265, n41266, n41267,
    n41268, n41269, n41270, n41271, n41272, n41273,
    n41274, n41275, n41276, n41277, n41278, n41279,
    n41280, n41281, n41282, n41283, n41284, n41285,
    n41286, n41287, n41288, n41289, n41290, n41291,
    n41292, n41293, n41294, n41295, n41296, n41297,
    n41298, n41299, n41300, n41301, n41302, n41303,
    n41304, n41305, n41307, n41308, n41309, n41310,
    n41311, n41312, n41313, n41314, n41315, n41316,
    n41317, n41318, n41319, n41320, n41321, n41322,
    n41323, n41324, n41325, n41326, n41327, n41328,
    n41329, n41330, n41331, n41332, n41333, n41334,
    n41335, n41336, n41337, n41338, n41339, n41340,
    n41341, n41342, n41343, n41344, n41345, n41346,
    n41347, n41348, n41349, n41350, n41351, n41352,
    n41353, n41354, n41355, n41356, n41357, n41358,
    n41359, n41360, n41361, n41362, n41363, n41364,
    n41365, n41366, n41367, n41368, n41369, n41370,
    n41371, n41372, n41373, n41374, n41375, n41376,
    n41377, n41378, n41379, n41380, n41381, n41382,
    n41383, n41384, n41385, n41386, n41387, n41388,
    n41389, n41390, n41391, n41392, n41393, n41394,
    n41395, n41396, n41397, n41398, n41399, n41400,
    n41401, n41402, n41403, n41404, n41405, n41406,
    n41407, n41408, n41409, n41410, n41411, n41412,
    n41413, n41414, n41415, n41416, n41417, n41418,
    n41419, n41420, n41421, n41422, n41423, n41424,
    n41425, n41426, n41427, n41428, n41429, n41430,
    n41431, n41432, n41433, n41434, n41435, n41436,
    n41437, n41438, n41439, n41440, n41441, n41442,
    n41443, n41444, n41445, n41446, n41447, n41448,
    n41449, n41450, n41451, n41452, n41453, n41454,
    n41455, n41456, n41457, n41458, n41459, n41460,
    n41461, n41462, n41463, n41464, n41465, n41466,
    n41467, n41468, n41469, n41470, n41471, n41472,
    n41473, n41474, n41475, n41476, n41477, n41478,
    n41479, n41480, n41481, n41482, n41483, n41484,
    n41485, n41486, n41487, n41488, n41489, n41490,
    n41491, n41492, n41493, n41494, n41495, n41496,
    n41497, n41498, n41499, n41500, n41501, n41502,
    n41503, n41504, n41505, n41506, n41507, n41508,
    n41509, n41510, n41511, n41512, n41513, n41514,
    n41515, n41516, n41517, n41518, n41519, n41520,
    n41521, n41522, n41523, n41524, n41525, n41526,
    n41527, n41528, n41529, n41530, n41531, n41532,
    n41533, n41534, n41535, n41536, n41537, n41538,
    n41539, n41540, n41541, n41542, n41543, n41544,
    n41545, n41546, n41547, n41548, n41549, n41550,
    n41551, n41552, n41553, n41554, n41555, n41556,
    n41557, n41558, n41559, n41560, n41561, n41562,
    n41563, n41564, n41565, n41566, n41567, n41568,
    n41569, n41570, n41571, n41572, n41573, n41574,
    n41575, n41576, n41577, n41578, n41580, n41581,
    n41582, n41583, n41584, n41585, n41586, n41587,
    n41588, n41589, n41590, n41591, n41592, n41593,
    n41594, n41595, n41596, n41597, n41598, n41599,
    n41600, n41601, n41602, n41603, n41604, n41605,
    n41606, n41607, n41608, n41609, n41610, n41611,
    n41612, n41613, n41614, n41615, n41616, n41617,
    n41618, n41619, n41620, n41621, n41622, n41623,
    n41624, n41625, n41626, n41627, n41628, n41629,
    n41630, n41631, n41632, n41633, n41634, n41635,
    n41636, n41637, n41638, n41639, n41640, n41641,
    n41642, n41643, n41644, n41645, n41646, n41647,
    n41648, n41649, n41650, n41651, n41652, n41653,
    n41654, n41655, n41656, n41657, n41658, n41659,
    n41660, n41661, n41662, n41663, n41664, n41665,
    n41666, n41667, n41668, n41669, n41670, n41671,
    n41672, n41673, n41674, n41675, n41676, n41677,
    n41678, n41679, n41680, n41681, n41682, n41683,
    n41684, n41685, n41686, n41687, n41688, n41689,
    n41690, n41691, n41692, n41693, n41694, n41695,
    n41696, n41697, n41698, n41699, n41700, n41701,
    n41702, n41703, n41704, n41705, n41706, n41707,
    n41708, n41709, n41710, n41711, n41712, n41713,
    n41714, n41715, n41716, n41717, n41718, n41719,
    n41720, n41721, n41722, n41723, n41724, n41725,
    n41726, n41727, n41728, n41729, n41730, n41731,
    n41732, n41733, n41734, n41735, n41736, n41737,
    n41738, n41739, n41740, n41741, n41742, n41743,
    n41744, n41745, n41746, n41747, n41748, n41749,
    n41750, n41751, n41752, n41753, n41754, n41755,
    n41756, n41757, n41758, n41759, n41760, n41761,
    n41762, n41763, n41764, n41765, n41766, n41767,
    n41768, n41769, n41770, n41771, n41772, n41773,
    n41774, n41775, n41776, n41777, n41778, n41779,
    n41780, n41781, n41782, n41783, n41784, n41785,
    n41786, n41787, n41788, n41789, n41790, n41791,
    n41792, n41793, n41794, n41795, n41796, n41797,
    n41798, n41799, n41800, n41801, n41802, n41803,
    n41804, n41805, n41806, n41807, n41808, n41810,
    n41811, n41812, n41813, n41814, n41815, n41816,
    n41817, n41818, n41819, n41820, n41821, n41822,
    n41823, n41824, n41825, n41826, n41827, n41828,
    n41829, n41830, n41831, n41832, n41833, n41834,
    n41835, n41836, n41837, n41838, n41839, n41840,
    n41841, n41842, n41843, n41844, n41845, n41846,
    n41847, n41848, n41849, n41850, n41851, n41852,
    n41853, n41854, n41855, n41856, n41857, n41858,
    n41859, n41860, n41861, n41862, n41863, n41864,
    n41865, n41866, n41867, n41868, n41869, n41870,
    n41871, n41872, n41873, n41874, n41875, n41876,
    n41877, n41878, n41879, n41880, n41881, n41882,
    n41883, n41884, n41885, n41886, n41887, n41888,
    n41889, n41890, n41891, n41892, n41893, n41894,
    n41895, n41896, n41897, n41898, n41899, n41900,
    n41901, n41902, n41903, n41904, n41905, n41906,
    n41907, n41908, n41909, n41910, n41911, n41912,
    n41913, n41914, n41915, n41916, n41917, n41918,
    n41919, n41920, n41921, n41922, n41923, n41924,
    n41925, n41926, n41927, n41928, n41929, n41930,
    n41931, n41932, n41933, n41934, n41935, n41936,
    n41937, n41938, n41939, n41940, n41941, n41942,
    n41943, n41944, n41945, n41946, n41947, n41948,
    n41949, n41950, n41951, n41952, n41953, n41954,
    n41955, n41956, n41957, n41958, n41959, n41960,
    n41961, n41962, n41963, n41964, n41965, n41966,
    n41967, n41968, n41969, n41970, n41971, n41973,
    n41974, n41975, n41976, n41977, n41978, n41979,
    n41980, n41981, n41982, n41983, n41984, n41985,
    n41986, n41987, n41988, n41989, n41990, n41991,
    n41992, n41993, n41994, n41995, n41996, n41997,
    n41998, n41999, n42000, n42001, n42002, n42003,
    n42004, n42005, n42006, n42007, n42008, n42009,
    n42010, n42011, n42012, n42013, n42014, n42015,
    n42016, n42017, n42018, n42019, n42020, n42021,
    n42022, n42023, n42024, n42025, n42026, n42027,
    n42028, n42029, n42030, n42031, n42032, n42033,
    n42034, n42035, n42036, n42037, n42038, n42039,
    n42040, n42041, n42042, n42043, n42044, n42045,
    n42046, n42047, n42048, n42049, n42050, n42051,
    n42052, n42053, n42054, n42055, n42056, n42057,
    n42058, n42059, n42060, n42061, n42062, n42063,
    n42064, n42065, n42066, n42067, n42068, n42069,
    n42070, n42071, n42072, n42073, n42074, n42075,
    n42076, n42077, n42078, n42079, n42080, n42081,
    n42082, n42083, n42084, n42085, n42086, n42087,
    n42088, n42089, n42090, n42091, n42092, n42093,
    n42094, n42095, n42096, n42097, n42098, n42099,
    n42100, n42101, n42102, n42103, n42104, n42105,
    n42106, n42107, n42108, n42109, n42110, n42111,
    n42112, n42113, n42114, n42115, n42116, n42117,
    n42118, n42119, n42120, n42121, n42122, n42123,
    n42124, n42125, n42126, n42127, n42128, n42129,
    n42130, n42131, n42132, n42133, n42134, n42135,
    n42136, n42137, n42138, n42139, n42140, n42141,
    n42142, n42143, n42144, n42145, n42146, n42147,
    n42148, n42149, n42150, n42151, n42152, n42153,
    n42154, n42155, n42156, n42157, n42158, n42159,
    n42161, n42162, n42163, n42164, n42165, n42166,
    n42167, n42169, n42170, n42171, n42172, n42173,
    n42174, n42175, n42176, n42177, n42179, n42180,
    n42181, n42182, n42183, n42184, n42185, n42186,
    n42187, n42188, n42189, n42190, n42191, n42192,
    n42193, n42194, n42195, n42196, n42197, n42198,
    n42199, n42200, n42201, n42202, n42203, n42204,
    n42205, n42206, n42207, n42208, n42209, n42210,
    n42211, n42212, n42213, n42214, n42215, n42216,
    n42217, n42218, n42219, n42221, n42222, n42223,
    n42224, n42225, n42226, n42227, n42228, n42229,
    n42230, n42231, n42232, n42233, n42234, n42235,
    n42236, n42237, n42238, n42239, n42240, n42241,
    n42242, n42243, n42244, n42245, n42246, n42247,
    n42248, n42249, n42250, n42251, n42252, n42253,
    n42254, n42255, n42256, n42257, n42258, n42259,
    n42260, n42261, n42262, n42263, n42264, n42265,
    n42266, n42267, n42268, n42269, n42270, n42271,
    n42272, n42273, n42274, n42275, n42276, n42277,
    n42278, n42279, n42280, n42281, n42282, n42283,
    n42284, n42285, n42286, n42287, n42288, n42289,
    n42290, n42291, n42292, n42293, n42294, n42295,
    n42296, n42297, n42298, n42299, n42300, n42301,
    n42302, n42303, n42304, n42305, n42306, n42307,
    n42308, n42309, n42310, n42311, n42312, n42313,
    n42314, n42315, n42316, n42317, n42318, n42319,
    n42320, n42321, n42322, n42323, n42324, n42325,
    n42326, n42327, n42328, n42329, n42330, n42331,
    n42332, n42333, n42334, n42335, n42336, n42337,
    n42338, n42339, n42340, n42341, n42342, n42343,
    n42344, n42345, n42346, n42347, n42348, n42349,
    n42350, n42351, n42352, n42353, n42354, n42355,
    n42356, n42357, n42358, n42359, n42360, n42361,
    n42362, n42363, n42364, n42365, n42366, n42367,
    n42368, n42369, n42370, n42371, n42372, n42373,
    n42374, n42375, n42376, n42377, n42378, n42379,
    n42380, n42381, n42382, n42383, n42384, n42385,
    n42386, n42387, n42388, n42389, n42390, n42391,
    n42392, n42393, n42394, n42395, n42396, n42397,
    n42398, n42399, n42400, n42401, n42402, n42403,
    n42404, n42405, n42406, n42407, n42408, n42409,
    n42410, n42411, n42412, n42413, n42414, n42415,
    n42416, n42417, n42418, n42419, n42420, n42421,
    n42422, n42423, n42424, n42425, n42426, n42427,
    n42428, n42429, n42430, n42431, n42432, n42433,
    n42434, n42435, n42436, n42437, n42438, n42439,
    n42440, n42441, n42442, n42443, n42444, n42445,
    n42446, n42447, n42448, n42449, n42450, n42451,
    n42452, n42453, n42454, n42455, n42457, n42458,
    n42459, n42460, n42461, n42462, n42463, n42464,
    n42465, n42466, n42467, n42468, n42469, n42470,
    n42471, n42472, n42473, n42474, n42475, n42476,
    n42477, n42478, n42479, n42480, n42481, n42482,
    n42483, n42484, n42485, n42486, n42487, n42488,
    n42489, n42490, n42491, n42492, n42493, n42494,
    n42495, n42496, n42497, n42498, n42499, n42500,
    n42501, n42502, n42503, n42504, n42505, n42506,
    n42507, n42508, n42509, n42510, n42511, n42512,
    n42513, n42514, n42515, n42516, n42517, n42518,
    n42519, n42520, n42521, n42522, n42523, n42524,
    n42525, n42526, n42527, n42528, n42529, n42530,
    n42531, n42532, n42533, n42534, n42535, n42536,
    n42537, n42538, n42539, n42540, n42541, n42542,
    n42543, n42544, n42545, n42546, n42547, n42548,
    n42549, n42550, n42551, n42552, n42553, n42554,
    n42555, n42556, n42557, n42558, n42559, n42560,
    n42561, n42562, n42563, n42564, n42565, n42566,
    n42567, n42568, n42569, n42570, n42571, n42572,
    n42573, n42574, n42575, n42576, n42577, n42578,
    n42579, n42580, n42581, n42582, n42583, n42584,
    n42585, n42586, n42587, n42588, n42589, n42590,
    n42591, n42592, n42593, n42594, n42595, n42596,
    n42597, n42598, n42599, n42600, n42601, n42602,
    n42603, n42604, n42605, n42606, n42607, n42608,
    n42609, n42610, n42611, n42612, n42613, n42614,
    n42615, n42616, n42617, n42618, n42619, n42620,
    n42621, n42622, n42623, n42624, n42625, n42626,
    n42627, n42628, n42629, n42630, n42631, n42632,
    n42633, n42634, n42635, n42636, n42637, n42638,
    n42639, n42640, n42641, n42642, n42643, n42644,
    n42645, n42646, n42647, n42648, n42649, n42650,
    n42651, n42652, n42653, n42654, n42655, n42656,
    n42657, n42658, n42659, n42660, n42661, n42662,
    n42663, n42664, n42665, n42666, n42667, n42668,
    n42669, n42670, n42671, n42672, n42673, n42674,
    n42675, n42676, n42677, n42678, n42679, n42681,
    n42682, n42683, n42684, n42685, n42687, n42688,
    n42689, n42690, n42691, n42693, n42694, n42695,
    n42696, n42697, n42699, n42700, n42701, n42702,
    n42703, n42705, n42706, n42707, n42708, n42709,
    n42711, n42712, n42713, n42714, n42715, n42716,
    n42718, n42719, n42720, n42721, n42722, n42723,
    n42725, n42726, n42727, n42728, n42729, n42730,
    n42731, n42732, n42733, n42734, n42735, n42736,
    n42737, n42738, n42739, n42740, n42741, n42742,
    n42743, n42744, n42745, n42746, n42747, n42748,
    n42749, n42750, n42751, n42752, n42753, n42754,
    n42755, n42756, n42757, n42759, n42760, n42761,
    n42762, n42763, n42764, n42765, n42766, n42767,
    n42768, n42769, n42770, n42771, n42772, n42773,
    n42774, n42775, n42776, n42777, n42778, n42779,
    n42780, n42781, n42782, n42783, n42784, n42785,
    n42786, n42787, n42788, n42789, n42790, n42791,
    n42792, n42793, n42794, n42795, n42796, n42797,
    n42798, n42799, n42800, n42801, n42802, n42803,
    n42804, n42805, n42806, n42807, n42808, n42809,
    n42810, n42811, n42812, n42813, n42814, n42815,
    n42816, n42817, n42818, n42819, n42820, n42821,
    n42822, n42823, n42824, n42825, n42826, n42827,
    n42828, n42829, n42830, n42831, n42832, n42833,
    n42834, n42835, n42836, n42837, n42838, n42839,
    n42840, n42841, n42842, n42843, n42844, n42845,
    n42846, n42847, n42848, n42849, n42850, n42851,
    n42852, n42853, n42854, n42855, n42856, n42857,
    n42858, n42859, n42860, n42861, n42862, n42863,
    n42864, n42865, n42866, n42867, n42868, n42869,
    n42870, n42871, n42872, n42873, n42874, n42875,
    n42876, n42877, n42878, n42879, n42880, n42881,
    n42882, n42883, n42884, n42885, n42886, n42887,
    n42888, n42889, n42890, n42891, n42892, n42893,
    n42894, n42895, n42896, n42897, n42898, n42899,
    n42900, n42901, n42902, n42903, n42904, n42905,
    n42906, n42907, n42908, n42909, n42910, n42911,
    n42912, n42913, n42914, n42915, n42916, n42917,
    n42918, n42919, n42920, n42921, n42922, n42923,
    n42924, n42925, n42926, n42927, n42928, n42929,
    n42930, n42931, n42932, n42933, n42934, n42935,
    n42936, n42937, n42938, n42939, n42940, n42941,
    n42942, n42943, n42944, n42945, n42946, n42947,
    n42948, n42949, n42950, n42951, n42952, n42953,
    n42954, n42955, n42956, n42957, n42958, n42959,
    n42960, n42961, n42962, n42963, n42964, n42965,
    n42966, n42967, n42969, n42970, n42971, n42972,
    n42973, n42974, n42975, n42976, n42977, n42978,
    n42979, n42980, n42981, n42982, n42983, n42984,
    n42985, n42986, n42987, n42988, n42989, n42990,
    n42991, n42992, n42993, n42994, n42995, n42996,
    n42997, n42998, n42999, n43000, n43001, n43002,
    n43003, n43004, n43005, n43006, n43007, n43008,
    n43009, n43010, n43011, n43012, n43014, n43015,
    n43016, n43017, n43018, n43019, n43020, n43021,
    n43022, n43023, n43024, n43025, n43026, n43027,
    n43028, n43029, n43030, n43031, n43032, n43033,
    n43034, n43035, n43036, n43037, n43038, n43039,
    n43040, n43041, n43042, n43043, n43044, n43045,
    n43046, n43047, n43048, n43049, n43050, n43051,
    n43052, n43053, n43055, n43056, n43057, n43058,
    n43059, n43060, n43061, n43062, n43063, n43064,
    n43065, n43066, n43067, n43068, n43069, n43070,
    n43071, n43072, n43073, n43074, n43075, n43076,
    n43077, n43078, n43079, n43080, n43081, n43082,
    n43083, n43084, n43085, n43086, n43087, n43088,
    n43089, n43090, n43091, n43092, n43093, n43094,
    n43095, n43096, n43097, n43098, n43099, n43100,
    n43101, n43102, n43103, n43104, n43105, n43106,
    n43107, n43108, n43109, n43110, n43111, n43112,
    n43113, n43114, n43115, n43116, n43117, n43118,
    n43119, n43120, n43122, n43123, n43124, n43125,
    n43126, n43127, n43128, n43129, n43130, n43131,
    n43132, n43133, n43134, n43135, n43136, n43137,
    n43138, n43139, n43140, n43141, n43142, n43143,
    n43144, n43145, n43146, n43147, n43148, n43149,
    n43150, n43151, n43152, n43153, n43154, n43155,
    n43156, n43157, n43158, n43159, n43160, n43161,
    n43162, n43163, n43164, n43165, n43166, n43167,
    n43168, n43169, n43170, n43171, n43172, n43173,
    n43174, n43175, n43176, n43177, n43178, n43179,
    n43180, n43181, n43182, n43183, n43184, n43185,
    n43186, n43187, n43188, n43189, n43190, n43191,
    n43192, n43193, n43194, n43195, n43196, n43197,
    n43198, n43199, n43200, n43201, n43202, n43203,
    n43204, n43205, n43206, n43207, n43208, n43209,
    n43210, n43211, n43212, n43213, n43214, n43215,
    n43216, n43217, n43218, n43219, n43220, n43221,
    n43222, n43223, n43224, n43225, n43226, n43227,
    n43228, n43229, n43230, n43231, n43232, n43233,
    n43234, n43235, n43236, n43237, n43238, n43239,
    n43240, n43241, n43242, n43243, n43244, n43245,
    n43246, n43247, n43248, n43249, n43250, n43251,
    n43252, n43253, n43254, n43255, n43256, n43257,
    n43258, n43259, n43260, n43261, n43262, n43263,
    n43264, n43265, n43266, n43267, n43268, n43269,
    n43270, n43271, n43272, n43273, n43274, n43275,
    n43276, n43277, n43278, n43279, n43280, n43281,
    n43282, n43283, n43284, n43285, n43286, n43287,
    n43288, n43289, n43290, n43291, n43292, n43293,
    n43294, n43295, n43296, n43297, n43298, n43299,
    n43300, n43301, n43302, n43303, n43304, n43305,
    n43306, n43307, n43308, n43309, n43310, n43311,
    n43312, n43313, n43314, n43315, n43316, n43317,
    n43318, n43319, n43320, n43321, n43322, n43323,
    n43324, n43325, n43326, n43327, n43329, n43330,
    n43331, n43332, n43333, n43334, n43335, n43336,
    n43337, n43338, n43339, n43340, n43341, n43342,
    n43343, n43344, n43345, n43346, n43347, n43348,
    n43349, n43350, n43351, n43352, n43353, n43354,
    n43355, n43356, n43357, n43358, n43359, n43360,
    n43361, n43362, n43363, n43364, n43365, n43366,
    n43367, n43368, n43369, n43370, n43371, n43372,
    n43373, n43374, n43375, n43376, n43377, n43378,
    n43379, n43380, n43381, n43382, n43383, n43384,
    n43385, n43386, n43387, n43388, n43389, n43390,
    n43391, n43392, n43393, n43394, n43395, n43396,
    n43397, n43398, n43399, n43400, n43401, n43402,
    n43403, n43404, n43405, n43406, n43407, n43408,
    n43409, n43410, n43411, n43412, n43413, n43414,
    n43415, n43416, n43417, n43418, n43419, n43420,
    n43421, n43422, n43423, n43424, n43425, n43426,
    n43427, n43428, n43429, n43430, n43431, n43432,
    n43433, n43434, n43435, n43436, n43437, n43438,
    n43439, n43440, n43441, n43442, n43443, n43444,
    n43445, n43446, n43447, n43448, n43449, n43450,
    n43451, n43452, n43453, n43454, n43455, n43456,
    n43457, n43458, n43459, n43460, n43461, n43462,
    n43463, n43464, n43465, n43466, n43467, n43468,
    n43469, n43470, n43471, n43472, n43473, n43474,
    n43475, n43476, n43477, n43478, n43479, n43480,
    n43481, n43482, n43483, n43484, n43486, n43487,
    n43488, n43489, n43490, n43491, n43492, n43493,
    n43494, n43495, n43496, n43497, n43498, n43499,
    n43500, n43501, n43502, n43503, n43504, n43505,
    n43506, n43507, n43508, n43509, n43510, n43511,
    n43512, n43513, n43514, n43515, n43516, n43517,
    n43518, n43519, n43520, n43521, n43522, n43523,
    n43524, n43525, n43526, n43527, n43528, n43529,
    n43531, n43532, n43533, n43534, n43535, n43536,
    n43537, n43538, n43539, n43540, n43541, n43542,
    n43543, n43544, n43545, n43546, n43547, n43548,
    n43549, n43550, n43551, n43552, n43553, n43554,
    n43555, n43556, n43557, n43558, n43559, n43560,
    n43561, n43562, n43563, n43564, n43565, n43566,
    n43567, n43568, n43569, n43570, n43571, n43572,
    n43573, n43575, n43576, n43577, n43578, n43579,
    n43580, n43581, n43582, n43583, n43584, n43585,
    n43586, n43587, n43588, n43589, n43590, n43591,
    n43592, n43593, n43594, n43595, n43596, n43597,
    n43598, n43599, n43600, n43601, n43602, n43603,
    n43604, n43605, n43606, n43607, n43608, n43609,
    n43610, n43611, n43612, n43613, n43614, n43615,
    n43616, n43617, n43618, n43619, n43620, n43621,
    n43622, n43624, n43625, n43626, n43627, n43628,
    n43629, n43630, n43631, n43632, n43633, n43634,
    n43635, n43636, n43637, n43638, n43639, n43640,
    n43641, n43642, n43643, n43644, n43645, n43646,
    n43647, n43648, n43649, n43650, n43651, n43652,
    n43653, n43654, n43655, n43656, n43657, n43658,
    n43659, n43660, n43661, n43662, n43663, n43664,
    n43665, n43666, n43667, n43668, n43669, n43670,
    n43671, n43672, n43673, n43674, n43675, n43676,
    n43677, n43678, n43679, n43680, n43681, n43682,
    n43683, n43684, n43685, n43686, n43687, n43688,
    n43689, n43690, n43691, n43692, n43693, n43694,
    n43695, n43696, n43697, n43698, n43699, n43700,
    n43701, n43702, n43703, n43704, n43705, n43706,
    n43707, n43708, n43709, n43710, n43711, n43712,
    n43713, n43714, n43715, n43717, n43718, n43719,
    n43720, n43721, n43722, n43723, n43724, n43725,
    n43726, n43727, n43728, n43729, n43730, n43731,
    n43732, n43733, n43734, n43735, n43736, n43737,
    n43738, n43739, n43740, n43741, n43742, n43743,
    n43744, n43745, n43746, n43747, n43748, n43749,
    n43750, n43751, n43752, n43753, n43754, n43755,
    n43756, n43757, n43758, n43759, n43760, n43761,
    n43762, n43763, n43764, n43765, n43766, n43767,
    n43768, n43769, n43770, n43771, n43772, n43773,
    n43774, n43775, n43776, n43777, n43778, n43780,
    n43781, n43782, n43783, n43784, n43785, n43786,
    n43787, n43788, n43789, n43790, n43791, n43792,
    n43793, n43794, n43795, n43796, n43797, n43798,
    n43799, n43800, n43801, n43802, n43803, n43804,
    n43805, n43806, n43807, n43808, n43809, n43810,
    n43811, n43812, n43813, n43814, n43815, n43816,
    n43817, n43818, n43819, n43821, n43822, n43823,
    n43824, n43825, n43826, n43827, n43828, n43829,
    n43830, n43831, n43832, n43833, n43834, n43835,
    n43836, n43837, n43838, n43839, n43840, n43841,
    n43842, n43843, n43844, n43845, n43846, n43847,
    n43848, n43849, n43850, n43851, n43852, n43853,
    n43854, n43855, n43856, n43857, n43858, n43859,
    n43860, n43861, n43862, n43863, n43864, n43865,
    n43866, n43867, n43868, n43869, n43870, n43871,
    n43872, n43873, n43874, n43875, n43876, n43877,
    n43878, n43879, n43880, n43881, n43882, n43883,
    n43884, n43885, n43886, n43887, n43888, n43889,
    n43890, n43891, n43892, n43893, n43894, n43896,
    n43897, n43898, n43899, n43900, n43901, n43902,
    n43903, n43904, n43905, n43906, n43907, n43908,
    n43909, n43910, n43911, n43912, n43913, n43914,
    n43915, n43916, n43917, n43918, n43919, n43920,
    n43921, n43922, n43923, n43925, n43926, n43927,
    n43928, n43929, n43930, n43931, n43932, n43933,
    n43934, n43935, n43936, n43937, n43938, n43939,
    n43940, n43941, n43942, n43943, n43944, n43945,
    n43946, n43947, n43948, n43949, n43950, n43951,
    n43952, n43953, n43954, n43955, n43956, n43957,
    n43958, n43959, n43960, n43961, n43962, n43963,
    n43964, n43965, n43966, n43968, n43969, n43970,
    n43971, n43972, n43973, n43974, n43975, n43976,
    n43977, n43978, n43979, n43980, n43981, n43982,
    n43983, n43984, n43985, n43986, n43987, n43988,
    n43989, n43990, n43991, n43992, n43993, n43994,
    n43995, n43996, n43997, n43998, n43999, n44000,
    n44001, n44002, n44003, n44004, n44005, n44006,
    n44007, n44008, n44009, n44010, n44011, n44012,
    n44013, n44014, n44015, n44016, n44017, n44018,
    n44019, n44020, n44021, n44022, n44023, n44024,
    n44025, n44026, n44027, n44028, n44029, n44030,
    n44031, n44032, n44033, n44035, n44036, n44037,
    n44038, n44039, n44040, n44041, n44042, n44043,
    n44044, n44045, n44046, n44047, n44048, n44049,
    n44050, n44051, n44052, n44053, n44054, n44055,
    n44056, n44057, n44058, n44059, n44060, n44061,
    n44062, n44063, n44064, n44065, n44066, n44067,
    n44068, n44069, n44070, n44071, n44072, n44073,
    n44074, n44075, n44076, n44077, n44078, n44079,
    n44080, n44081, n44082, n44083, n44084, n44085,
    n44086, n44087, n44088, n44089, n44090, n44091,
    n44092, n44094, n44095, n44096, n44097, n44098,
    n44099, n44100, n44101, n44102, n44103, n44104,
    n44105, n44106, n44107, n44108, n44109, n44110,
    n44111, n44112, n44113, n44114, n44115, n44116,
    n44117, n44118, n44119, n44120, n44121, n44122,
    n44123, n44124, n44125, n44126, n44127, n44128,
    n44129, n44130, n44131, n44132, n44133, n44134,
    n44135, n44136, n44138, n44139, n44140, n44141,
    n44142, n44143, n44144, n44145, n44146, n44147,
    n44148, n44149, n44150, n44151, n44152, n44153,
    n44154, n44155, n44156, n44157, n44158, n44159,
    n44160, n44161, n44162, n44163, n44164, n44165,
    n44166, n44167, n44168, n44169, n44170, n44171,
    n44172, n44173, n44174, n44175, n44177, n44178,
    n44179, n44180, n44181, n44182, n44183, n44184,
    n44185, n44186, n44187, n44188, n44189, n44190,
    n44191, n44192, n44193, n44194, n44195, n44196,
    n44197, n44198, n44199, n44200, n44201, n44202,
    n44203, n44204, n44205, n44206, n44207, n44208,
    n44209, n44210, n44211, n44212, n44213, n44214,
    n44216, n44217, n44218, n44219, n44220, n44221,
    n44222, n44223, n44224, n44225, n44226, n44227,
    n44228, n44229, n44230, n44231, n44232, n44233,
    n44234, n44235, n44236, n44237, n44238, n44239,
    n44240, n44241, n44242, n44243, n44244, n44245,
    n44246, n44247, n44248, n44249, n44250, n44251,
    n44252, n44253, n44254, n44255, n44256, n44257,
    n44258, n44259, n44260, n44261, n44262, n44263,
    n44264, n44265, n44266, n44267, n44268, n44269,
    n44270, n44271, n44272, n44273, n44275, n44276,
    n44277, n44279, n44280, n44281, n44282, n44283,
    n44284, n44285, n44286, n44287, n44288, n44289,
    n44290, n44291, n44292, n44293, n44294, n44295,
    n44296, n44298, n44299, n44300, n44301, n44302,
    n44303, n44304, n44305, n44306, n44307, n44308,
    n44309, n44310, n44311, n44312, n44313, n44314,
    n44316, n44318, n44319, n44321, n44322, n44323,
    n44325, n44326, n44327, n44328, n44329, n44330,
    n44331, n44332, n44333, n44334, n44335, n44336,
    n44338, n44339, n44341, n44342, n44344, n44345,
    n44347, n44348, n44350, n44351, n44353, n44354,
    n44356, n44357, n44359, n44360, n44362, n44363,
    n44365, n44366, n44367, n44368, n44369, n44370,
    n44371, n44373, n44374, n44375, n44376, n44377,
    n44378, n44380, n44381, n44382, n44384, n44385,
    n44386, n44387, n44388, n44389, n44390, n44391,
    n44392, n44393, n44394, n44395, n44396, n44397,
    n44398, n44399, n44400, n44401, n44402, n44403,
    n44404, n44406, n44407, n44409, n44410, n44412,
    n44413, n44415, n44416, n44418, n44419, n44421,
    n44422, n44424, n44425, n44427, n44428, n44429,
    n44430, n44431, n44432, n44433, n44434, n44435,
    n44436, n44437, n44438, n44439, n44440, n44441,
    n44442, n44443, n44444, n44445, n44446, n44447,
    n44448, n44449, n44450, n44451, n44452, n44454,
    n44455, n44456, n44458, n44459, n44461, n44462,
    n44463, n44465, n44466, n44468, n44469, n44470,
    n44471, n44472, n44473, n44474, n44475, n44476,
    n44477, n44478, n44480, n44481, n44482, n44483,
    n44485, n44486, n44488, n44489, n44490, n44492,
    n44493, n44494, n44495, n44497, n44498, n44500,
    n44501, n44503, n44504, n44506, n44507, n44509,
    n44510, n44512, n44513, n44515, n44516, n44518,
    n44519, n44521, n44522, n44524, n44525, n44527,
    n44528, n44530, n44531, n44532, n44533, n44534,
    n44535, n44536, n44538, n44539, n44540, n44541,
    n44543, n44544, n44545, n44546, n44547, n44548,
    n44549, n44550, n44551, n44552, n44553, n44555,
    n44556, n44558, n44559, n44561, n44562, n44564,
    n44565, n44567, n44568, n44570, n44571, n44573,
    n44574, n44576, n44577, n44578, n44579, n44580,
    n44582, n44583, n44585, n44586, n44588, n44589,
    n44591, n44592, n44594, n44595, n44597, n44598,
    n44600, n44601, n44603, n44604, n44606, n44607,
    n44609, n44610, n44612, n44613, n44615, n44616,
    n44618, n44619, n44621, n44622, n44624, n44625,
    n44627, n44628, n44630, n44631, n44633, n44634,
    n44636, n44637, n44639, n44640, n44642, n44643,
    n44645, n44646, n44648, n44649, n44651, n44652,
    n44654, n44655, n44657, n44658, n44660, n44661,
    n44663, n44664, n44666, n44667, n44669, n44670,
    n44672, n44673, n44675, n44676, n44678, n44679,
    n44681, n44682, n44684, n44685, n44687, n44688,
    n44690, n44691, n44693, n44694, n44696, n44697,
    n44699, n44700, n44702, n44703, n44705, n44706,
    n44708, n44709, n44711, n44712, n44714, n44715,
    n44717, n44718, n44720, n44721, n44723, n44724,
    n44726, n44727, n44729, n44730, n44732, n44733,
    n44735, n44736, n44738, n44739, n44741, n44742,
    n44744, n44745, n44747, n44748, n44750, n44751,
    n44753, n44754, n44756, n44757, n44759, n44760,
    n44762, n44763, n44765, n44766, n44768, n44769,
    n44771, n44772, n44774, n44775, n44777, n44778,
    n44780, n44781, n44783, n44784, n44786, n44787,
    n44789, n44790, n44792, n44793, n44795, n44796,
    n44798, n44799, n44801, n44802, n44803, n44805,
    n44806, n44808, n44809, n44811, n44812, n44814,
    n44815, n44817, n44818, n44820, n44821, n44823,
    n44824, n44826, n44827, n44829, n44830, n44832,
    n44833, n44835, n44836, n44838, n44839, n44841,
    n44842, n44844, n44845, n44847, n44848, n44850,
    n44851, n44853, n44854, n44856, n44857, n44859,
    n44860, n44862, n44863, n44865, n44866, n44868,
    n44869, n44871, n44872, n44874, n44875, n44877,
    n44878, n44880, n44881, n44883, n44884, n44886,
    n44887, n44889, n44890, n44892, n44893, n44895,
    n44896, n44898, n44899, n44901, n44902, n44904,
    n44905, n44907, n44908, n44910, n44911, n44913,
    n44914, n44916, n44917, n44919, n44920, n44922,
    n44923, n44925, n44926, n44928, n44929, n44931,
    n44932, n44933, n44934, n44935, n44936, n44937,
    n44938, n44939, n44940, n44941, n44942, n44943,
    n44944, n44945, n44946, n44947, n44948, n44949,
    n44950, n44951, n44952, n44953, n44955, n44956,
    n44958, n44959, n44961, n44962, n44964, n44965,
    n44967, n44968, n44970, n44971, n44973, n44974,
    n44976, n44977, n44978, n44979, n44980, n44981,
    n44982, n44983, n44984, n44985, n44986, n44987,
    n44988, n44989, n44990, n44991, n44992, n44993,
    n44994, n44995, n44996, n44997, n44998, n44999,
    n45001, n45002, n45003, n45004, n45005, n45006,
    n45007, n45008, n45009, n45010, n45011, n45012,
    n45013, n45014, n45015, n45016, n45017, n45019,
    n45020, n45021, n45022, n45023, n45024, n45025,
    n45026, n45027, n45028, n45029, n45030, n45031,
    n45032, n45033, n45034, n45035, n45036, n45037,
    n45038, n45039, n45040, n45041, n45042, n45043,
    n45044, n45045, n45046, n45047, n45049, n45050,
    n45051, n45052, n45053, n45055, n45056, n45057,
    n45058, n45059, n45060, n45061, n45062, n45063,
    n45064, n45065, n45066, n45067, n45068, n45069,
    n45070, n45071, n45072, n45073, n45075, n45076,
    n45077, n45078, n45079, n45080, n45081, n45082,
    n45083, n45084, n45085, n45086, n45087, n45088,
    n45089, n45090, n45091, n45092, n45093, n45095,
    n45096, n45097, n45098, n45099, n45100, n45101,
    n45102, n45103, n45104, n45105, n45106, n45107,
    n45108, n45109, n45110, n45111, n45112, n45113,
    n45115, n45116, n45117, n45118, n45119, n45120,
    n45121, n45122, n45123, n45124, n45125, n45126,
    n45127, n45128, n45129, n45130, n45131, n45132,
    n45133, n45135, n45136, n45137, n45138, n45139,
    n45140, n45141, n45142, n45143, n45144, n45146,
    n45147, n45148, n45149, n45150, n45151, n45152,
    n45153, n45154, n45155, n45157, n45158, n45159,
    n45160, n45161, n45162, n45163, n45164, n45165,
    n45166, n45168, n45169, n45170, n45171, n45172,
    n45173, n45174, n45175, n45176, n45177, n45178,
    n45181, n45182, n45184, n45185, n45187, n45188,
    n45190, n45191, n45193, n45194, n45196, n45197,
    n45199, n45200, n45202, n45203, n45205, n45206,
    n45208, n45209, n45211, n45212, n45214, n45215,
    n45217, n45218, n45220, n45221, n45223, n45224,
    n45226, n45227, n45229, n45230, n45232, n45233,
    n45235, n45236, n45238, n45239, n45241, n45242,
    n45244, n45245, n45247, n45248, n45250, n45251,
    n45253, n45254, n45255, n45256, n45257, n45258,
    n45259, n45260, n45262, n45263, n45265, n45266,
    n45268, n45269, n45271, n45272, n45274, n45275,
    n45277, n45278, n45279, n45280, n45281, n45283,
    n45284, n45286, n45287, n45289, n45290, n45292,
    n45293, n45295, n45296, n45298, n45299, n45301,
    n45302, n45303, n45304, n45305, n45307, n45308,
    n45310, n45311, n45313, n45314, n45316, n45317,
    n45319, n45320, n45321, n45322, n45324, n45325,
    n45327, n45328, n45330, n45331, n45333, n45334,
    n45336, n45337, n45339, n45340, n45342, n45343,
    n45345, n45346, n45348, n45349, n45351, n45352,
    n45354, n45355, n45357, n45358, n45360, n45361,
    n45363, n45364, n45366, n45367, n45369, n45370,
    n45372, n45373, n45375, n45376, n45378, n45379,
    n45381, n45382, n45384, n45385, n45386, n45387,
    n45389, n45390, n45392, n45393, n45395, n45396,
    n45398, n45399, n45401, n45402, n45404, n45405,
    n45407, n45408, n45410, n45411, n45413, n45414,
    n45416, n45417, n45419, n45420, n45422, n45423,
    n45425, n45426, n45427, n45428, n45430, n45431,
    n45433, n45434, n45436, n45437, n45439, n45440,
    n45442, n45443, n45445, n45446, n45448, n45449,
    n45451, n45452, n45454, n45455, n45457, n45458,
    n45459, n45460, n45461, n45462, n45463, n45464,
    n45465, n45466, n45467, n45468, n45469, n45470,
    n45471, n45472, n45473, n45474, n45475, n45476,
    n45477, n45478, n45479, n45480, n45481, n45482,
    n45483, n45484, n45485, n45486, n45487, n45488,
    n45489, n45490, n45491, n45492, n45493, n45494,
    n45495, n45496, n45497, n45498, n45499, n45500,
    n45501, n45502, n45503, n45504, n45505, n45506,
    n45507, n45508, n45509, n45510, n45511, n45512,
    n45513, n45514, n45515, n45516, n45517, n45518,
    n45519, n45520, n45521, n45522, n45523, n45524,
    n45525, n45526, n45527, n45528, n45529, n45530,
    n45531, n45532, n45533, n45534, n45535, n45536,
    n45537, n45538, n45539, n45540, n45541, n45542,
    n45543, n45544, n45545, n45546, n45547, n45548,
    n45549, n45550, n45551, n45552, n45553, n45554,
    n45555, n45556, n45557, n45558, n45559, n45560,
    n45561, n45562, n45563, n45564, n45565, n45567,
    n45568, n45570, n45571, n45573, n45574, n45575,
    n45576, n45578, n45579, n45581, n45582, n45584,
    n45585, n45587, n45588, n45590, n45591, n45593,
    n45594, n45596, n45597, n45599, n45600, n45602,
    n45603, n45605, n45606, n45608, n45609, n45611,
    n45612, n45614, n45615, n45617, n45618, n45620,
    n45621, n45623, n45624, n45625, n45626, n45627,
    n45628, n45630, n45631, n45632, n45633, n45635,
    n45636, n45637, n45638, n45639, n45640, n45641,
    n45642, n45643, n45644, n45645, n45646, n45647,
    n45648, n45649, n45650, n45651, n45652, n45653,
    n45654, n45656, n45657, n45658, n45660, n45661,
    n45662, n45664, n45665, n45666, n45668, n45669,
    n45670, n45671, n45672, n45673, n45674, n45675,
    n45676, n45677, n45678, n45679, n45680, n45681,
    n45682, n45683, n45684, n45685, n45686, n45687,
    n45688, n45689, n45690, n45691, n45692, n45693,
    n45694, n45695, n45696, n45697, n45698, n45699,
    n45700, n45701, n45702, n45703, n45704, n45705,
    n45706, n45707, n45708, n45709, n45710, n45711,
    n45712, n45713, n45714, n45715, n45716, n45717,
    n45718, n45719, n45720, n45721, n45722, n45723,
    n45724, n45725, n45726, n45727, n45728, n45729,
    n45730, n45731, n45732, n45733, n45734, n45735,
    n45736, n45737, n45738, n45739, n45740, n45741,
    n45742, n45743, n45744, n45745, n45746, n45747,
    n45748, n45749, n45750, n45751, n45752, n45753,
    n45754, n45755, n45756, n45757, n45758, n45759,
    n45760, n45761, n45762, n45763, n45764, n45765,
    n45766, n45767, n45768, n45769, n45770, n45771,
    n45772, n45773, n45774, n45775, n45776, n45777,
    n45778, n45779, n45780, n45781, n45782, n45783,
    n45784, n45785, n45786, n45787, n45788, n45789,
    n45790, n45791, n45792, n45793, n45794, n45795,
    n45796, n45797, n45798, n45799, n45800, n45801,
    n45802, n45803, n45804, n45805, n45806, n45807,
    n45808, n45809, n45810, n45811, n45812, n45813,
    n45814, n45815, n45816, n45817, n45818, n45819,
    n45820, n45821, n45822, n45823, n45824, n45825,
    n45826, n45827, n45828, n45829, n45830, n45831,
    n45832, n45833, n45834, n45835, n45836, n45837,
    n45838, n45839, n45840, n45841, n45842, n45843,
    n45844, n45845, n45846, n45847, n45848, n45849,
    n45850, n45851, n45852, n45853, n45854, n45855,
    n45856, n45857, n45858, n45859, n45860, n45861,
    n45862, n45863, n45864, n45865, n45866, n45867,
    n45868, n45869, n45870, n45871, n45872, n45873,
    n45874, n45875, n45876, n45877, n45878, n45879,
    n45880, n45881, n45882, n45883, n45884, n45885,
    n45886, n45887, n45888, n45889, n45890, n45891,
    n45892, n45893, n45894, n45895, n45896, n45897,
    n45898, n45899, n45900, n45901, n45902, n45903,
    n45904, n45905, n45906, n45907, n45908, n45909,
    n45910, n45911, n45912, n45913, n45914, n45915,
    n45916, n45917, n45918, n45919, n45920, n45921,
    n45922, n45923, n45924, n45925, n45926, n45927,
    n45928, n45929, n45930, n45931, n45932, n45933,
    n45934, n45935, n45936, n45937, n45938, n45939,
    n45940, n45941, n45942, n45943, n45944, n45945,
    n45946, n45947, n45948, n45949, n45950, n45951,
    n45952, n45953, n45954, n45955, n45956, n45957,
    n45958, n45959, n45960, n45961, n45962, n45963,
    n45964, n45965, n45966, n45967, n45968, n45969,
    n45970, n45971, n45972, n45973, n45974, n45975,
    n45976, n45977, n45978, n45979, n45980, n45981,
    n45982, n45983, n45984, n45985, n45986, n45987,
    n45988, n45989, n45990, n45991, n45992, n45993,
    n45994, n45995, n45996, n45997, n45998, n45999,
    n46000, n46001, n46002, n46003, n46004, n46005,
    n46006, n46007, n46008, n46009, n46010, n46011,
    n46012, n46013, n46014, n46015, n46016, n46017,
    n46018, n46019, n46020, n46021, n46022, n46023,
    n46024, n46025, n46026, n46027, n46028, n46029,
    n46030, n46031, n46032, n46033, n46034, n46035,
    n46036, n46037, n46038, n46039, n46040, n46041,
    n46042, n46043, n46044, n46045, n46046, n46047,
    n46048, n46049, n46050, n46051, n46052, n46053,
    n46054, n46055, n46056, n46057, n46058, n46059,
    n46060, n46061, n46062, n46063, n46064, n46065,
    n46066, n46067, n46068, n46069, n46070, n46071,
    n46072, n46073, n46074, n46075, n46076, n46077,
    n46078, n46079, n46080, n46081, n46082, n46083,
    n46084, n46085, n46086, n46087, n46088, n46089,
    n46090, n46091, n46092, n46093, n46094, n46095,
    n46096, n46097, n46098, n46099, n46100, n46101,
    n46102, n46103, n46104, n46105, n46106, n46107,
    n46108, n46109, n46110, n46111, n46112, n46113,
    n46114, n46115, n46116, n46117, n46118, n46119,
    n46120, n46121, n46122, n46123, n46124, n46125,
    n46126, n46127, n46128, n46129, n46130, n46131,
    n46132, n46133, n46134, n46135, n46136, n46137,
    n46138, n46139, n46140, n46141, n46142, n46143,
    n46144, n46145, n46146, n46147, n46148, n46149,
    n46150, n46151, n46152, n46153, n46154, n46155,
    n46156, n46157, n46158, n46159, n46160, n46161,
    n46162, n46163, n46164, n46165, n46166, n46167,
    n46168, n46169, n46170, n46171, n46172, n46173,
    n46174, n46175, n46176, n46177, n46178, n46179,
    n46180, n46181, n46182, n46183, n46184, n46185,
    n46186, n46187, n46188, n46189, n46190, n46191,
    n46192, n46193, n46194, n46195, n46196, n46197,
    n46198, n46199, n46200, n46201, n46202, n46203,
    n46204, n46205, n46206, n46207, n46208, n46209,
    n46210, n46211, n46212, n46213, n46214, n46215,
    n46216, n46217, n46218, n46219, n46220, n46221,
    n46222, n46223, n46224, n46225, n46226, n46227,
    n46228, n46229, n46230, n46231, n46232, n46233,
    n46234, n46235, n46236, n46237, n46238, n46239,
    n46240, n46241, n46242, n46243, n46244, n46245,
    n46246, n46247, n46248, n46249, n46250, n46251,
    n46252, n46253, n46254, n46255, n46256, n46257,
    n46258, n46259, n46260, n46261, n46262, n46263,
    n46264, n46265, n46266, n46267, n46268, n46269,
    n46270, n46271, n46272, n46273, n46274, n46275,
    n46276, n46277, n46278, n46279, n46280, n46281,
    n46282, n46283, n46284, n46285, n46286, n46287,
    n46288, n46289, n46290, n46291, n46292, n46293,
    n46294, n46295, n46296, n46297, n46298, n46299,
    n46300, n46301, n46302, n46303, n46304, n46305,
    n46306, n46307, n46308, n46309, n46310, n46311,
    n46312, n46313, n46314, n46315, n46316, n46317,
    n46318, n46319, n46320, n46321, n46322, n46323,
    n46324, n46325, n46326, n46327, n46328, n46329,
    n46330, n46331, n46332, n46333, n46334, n46335,
    n46336, n46337, n46338, n46339, n46340, n46341,
    n46342, n46343, n46344, n46345, n46346, n46347,
    n46348, n46349, n46350, n46351, n46352, n46353,
    n46354, n46355, n46356, n46357, n46358, n46359,
    n46360, n46361, n46362, n46363, n46364, n46365,
    n46366, n46367, n46368, n46369, n46370, n46371,
    n46372, n46373, n46374, n46375, n46376, n46377,
    n46378, n46379, n46380, n46382, n46383, n46384,
    n46385, n46386, n46387, n46389, n46390, n46391,
    n46392, n46393, n46395, n46396, n46397, n46398,
    n46399, n46401, n46402, n46403, n46405, n46406,
    n46407, n46408, n46409, n46411, n46412, n46413,
    n46415, n46416, n46418, n46419, n46420, n46422,
    n46423, n46424, n46425, n46426, n46427, n46428,
    n46429, n46430, n46431, n46432, n46434, n46435,
    n46436, n46437, n46439, n46440, n46441, n46442,
    n46443, n46444, n46445, n46446, n46448, n46449,
    n46450, n46451, n46452, n46453, n46455, n46456,
    n46458, n46459, n46460, n46461, n46462, n46464,
    n46465, n46466, n46468, n46469, n46470, n46472,
    n46473, n46474, n46476, n46477, n46478, n46480,
    n46481, n46482, n46484, n46485, n46486, n46488,
    n46489, n46490, n46492, n46493, n46494, n46495,
    n46497, n46498, n46499, n46500, n46502, n46503,
    n46504, n46505, n46507, n46508, n46509, n46510,
    n46511, n46513, n46514, n46515, n46517, n46518,
    n46519, n46521, n46522, n46523, n46525, n46526,
    n46527, n46529, n46530, n46531, n46533, n46534,
    n46535, n46537, n46538, n46539, n46540, n46541,
    n46543, n46544, n46545, n46546, n46548, n46549,
    n46550, n46552, n46553, n46554, n46556, n46557,
    n46558, n46560, n46561, n46562, n46564, n46565,
    n46566, n46568, n46569, n46570, n46572, n46573,
    n46574, n46576, n46577, n46578, n46580, n46581,
    n46582, n46584, n46585, n46586, n46588, n46589,
    n46590, n46592, n46593, n46594, n46596, n46597,
    n46598, n46600, n46601, n46602, n46604, n46605,
    n46606, n46608, n46609, n46610, n46612, n46613,
    n46614, n46616, n46617, n46618, n46620, n46621,
    n46622, n46624, n46625, n46626, n46628, n46629,
    n46630, n46632, n46633, n46634, n46636, n46637,
    n46638, n46640, n46641, n46642, n46644, n46645,
    n46646, n46648, n46649, n46650, n46652, n46653,
    n46654, n46656, n46657, n46658, n46660, n46661,
    n46662, n46664, n46665, n46666, n46668, n46669,
    n46670, n46672, n46673, n46674, n46676, n46677,
    n46678, n46680, n46681, n46682, n46684, n46685,
    n46686, n46687, n46688, n46689, n46690, n46691,
    n46692, n46694, n46696, n46697, n46698, n46700,
    n46701, n46702, n46704, n46705, n46706, n46708,
    n46709, n46710, n46711, n46712, n46713, n46714,
    n46715, n46716, n46717, n46718, n46719, n46720,
    n46721, n46722, n46723, n46724, n46725, n46726,
    n46727, n46728, n46729, n46730, n46731, n46732,
    n46733, n46734, n46735, n46736, n46737, n46738,
    n46739, n46740, n46741, n46742, n46743, n46744,
    n46745, n46746, n46747, n46748, n46749, n46750,
    n46751, n46752, n46753, n46754, n46755, n46757,
    n46758, n46759, n46760, n46761, n46762, n46763,
    n46764, n46765, n46766, n46767, n46768, n46769,
    n46770, n46771, n46772, n46773, n46774, n46775,
    n46776, n46777, n46778, n46779, n46780, n46781,
    n46782, n46783, n46784, n46785, n46786, n46787,
    n46788, n46789, n46790, n46791, n46792, n46793,
    n46794, n46795, n46796, n46797, n46799, n46800,
    n46801, n46803, n46804, n46805, n46806, n46807,
    n46808, n46809, n46810, n46811, n46812, n46813,
    n46814, n46815, n46816, n46817, n46818, n46819,
    n46820, n46821, n46822, n46823, n46824, n46825,
    n46826, n46827, n46828, n46829, n46830, n46831,
    n46832, n46833, n46834, n46835, n46836, n46837,
    n46839, n46840, n46841, n46842, n46843, n46844,
    n46845, n46846, n46847, n46848, n46849, n46850,
    n46851, n46852, n46853, n46854, n46855, n46856,
    n46857, n46858, n46859, n46860, n46861, n46862,
    n46863, n46864, n46865, n46866, n46867, n46868,
    n46869, n46870, n46871, n46872, n46873, n46874,
    n46876, n46877, n46878, n46879, n46880, n46881,
    n46882, n46883, n46884, n46885, n46886, n46887,
    n46888, n46889, n46890, n46891, n46892, n46893,
    n46894, n46895, n46896, n46897, n46898, n46899,
    n46900, n46901, n46902, n46903, n46904, n46905,
    n46906, n46907, n46908, n46909, n46910, n46912,
    n46913, n46914, n46916, n46917, n46918, n46919,
    n46920, n46921, n46922, n46923, n46924, n46925,
    n46926, n46927, n46928, n46929, n46930, n46931,
    n46932, n46933, n46934, n46935, n46936, n46937,
    n46938, n46939, n46940, n46941, n46942, n46943,
    n46944, n46945, n46946, n46947, n46949, n46950,
    n46951, n46952, n46953, n46954, n46955, n46956,
    n46957, n46958, n46959, n46960, n46961, n46962,
    n46963, n46964, n46965, n46966, n46967, n46968,
    n46969, n46970, n46971, n46972, n46973, n46974,
    n46975, n46976, n46977, n46978, n46979, n46981,
    n46982, n46983, n46984, n46985, n46986, n46987,
    n46988, n46989, n46990, n46991, n46992, n46993,
    n46994, n46995, n46996, n46997, n46998, n46999,
    n47000, n47001, n47002, n47003, n47004, n47005,
    n47006, n47007, n47008, n47009, n47010, n47011,
    n47012, n47013, n47014, n47015, n47017, n47018,
    n47019, n47020, n47021, n47022, n47023, n47024,
    n47025, n47026, n47027, n47028, n47029, n47030,
    n47031, n47032, n47033, n47034, n47035, n47036,
    n47037, n47038, n47039, n47040, n47041, n47042,
    n47043, n47044, n47045, n47046, n47047, n47048,
    n47049, n47050, n47051, n47053, n47054, n47055,
    n47056, n47057, n47058, n47059, n47060, n47061,
    n47062, n47063, n47064, n47065, n47066, n47067,
    n47068, n47069, n47070, n47071, n47072, n47073,
    n47074, n47075, n47076, n47077, n47078, n47079,
    n47080, n47081, n47082, n47083, n47084, n47085,
    n47086, n47087, n47088, n47089, n47091, n47092,
    n47093, n47094, n47095, n47096, n47097, n47098,
    n47099, n47100, n47101, n47102, n47103, n47104,
    n47105, n47106, n47107, n47108, n47109, n47110,
    n47111, n47112, n47113, n47114, n47115, n47116,
    n47117, n47118, n47119, n47120, n47121, n47122,
    n47123, n47124, n47125, n47127, n47128, n47129,
    n47130, n47131, n47132, n47133, n47134, n47135,
    n47136, n47137, n47138, n47139, n47140, n47141,
    n47142, n47143, n47144, n47145, n47146, n47147,
    n47148, n47149, n47150, n47151, n47152, n47153,
    n47154, n47155, n47156, n47157, n47158, n47159,
    n47160, n47161, n47163, n47164, n47165, n47166,
    n47167, n47168, n47169, n47170, n47171, n47172,
    n47173, n47174, n47175, n47176, n47177, n47178,
    n47179, n47180, n47181, n47182, n47183, n47184,
    n47185, n47186, n47187, n47188, n47189, n47190,
    n47191, n47192, n47193, n47195, n47196, n47197,
    n47198, n47199, n47200, n47201, n47202, n47203,
    n47204, n47205, n47206, n47207, n47208, n47209,
    n47210, n47211, n47212, n47213, n47214, n47215,
    n47216, n47217, n47218, n47219, n47220, n47221,
    n47222, n47223, n47224, n47225, n47227, n47228,
    n47229, n47230, n47231, n47232, n47233, n47234,
    n47235, n47236, n47237, n47238, n47239, n47240,
    n47241, n47242, n47243, n47244, n47245, n47246,
    n47247, n47248, n47249, n47250, n47251, n47252,
    n47253, n47254, n47255, n47256, n47257, n47258,
    n47259, n47260, n47261, n47262, n47264, n47265,
    n47266, n47268, n47269, n47270, n47272, n47273,
    n47274, n47275, n47276, n47277, n47278, n47279,
    n47280, n47281, n47282, n47283, n47284, n47285,
    n47286, n47287, n47288, n47289, n47290, n47291,
    n47292, n47293, n47294, n47295, n47296, n47297,
    n47298, n47299, n47300, n47301, n47302, n47305,
    n47306, n47307, n47309, n47310, n47311, n47312,
    n47313, n47314, n47315, n47316, n47317, n47318,
    n47319, n47320, n47321, n47322, n47323, n47324,
    n47325, n47326, n47327, n47328, n47329, n47330,
    n47331, n47332, n47333, n47334, n47335, n47336,
    n47337, n47338, n47339, n47340, n47341, n47342,
    n47343, n47344, n47345, n47346, n47348, n47349,
    n47350, n47352, n47353, n47354, n47356, n47357,
    n47358, n47360, n47361, n47362, n47363, n47364,
    n47365, n47366, n47367, n47368, n47369, n47370,
    n47371, n47372, n47373, n47374, n47375, n47376,
    n47377, n47378, n47379, n47380, n47381, n47382,
    n47383, n47384, n47385, n47386, n47387, n47388,
    n47389, n47390, n47391, n47392, n47394, n47395,
    n47396, n47398, n47399, n47400, n47402, n47403,
    n47404, n47405, n47406, n47407, n47408, n47409,
    n47410, n47411, n47412, n47413, n47414, n47415,
    n47416, n47417, n47418, n47419, n47420, n47421,
    n47422, n47423, n47424, n47425, n47426, n47427,
    n47428, n47429, n47430, n47431, n47432, n47433,
    n47434, n47435, n47437, n47438, n47439, n47441,
    n47442, n47443, n47445, n47446, n47447, n47449,
    n47450, n47451, n47453, n47454, n47455, n47457,
    n47458, n47459, n47461, n47462, n47463, n47465,
    n47466, n47467, n47469, n47470, n47471, n47473,
    n47474, n47475, n47477, n47478, n47479, n47481,
    n47482, n47483, n47485, n47486, n47487, n47489,
    n47490, n47491, n47493, n47494, n47495, n47496,
    n47497, n47498, n47499, n47500, n47501, n47502,
    n47503, n47504, n47505, n47506, n47507, n47508,
    n47509, n47510, n47511, n47512, n47513, n47514,
    n47515, n47516, n47517, n47518, n47519, n47520,
    n47521, n47522, n47523, n47524, n47525, n47526,
    n47527, n47529, n47530, n47531, n47532, n47533,
    n47534, n47535, n47536, n47537, n47538, n47539,
    n47540, n47541, n47542, n47543, n47544, n47545,
    n47546, n47547, n47548, n47549, n47550, n47551,
    n47552, n47553, n47554, n47555, n47556, n47557,
    n47558, n47559, n47560, n47561, n47562, n47563,
    n47564, n47565, n47566, n47567, n47569, n47570,
    n47571, n47573, n47574, n47575, n47577, n47578,
    n47579, n47580, n47581, n47582, n47583, n47584,
    n47585, n47586, n47587, n47588, n47589, n47590,
    n47591, n47592, n47593, n47594, n47595, n47596,
    n47597, n47598, n47599, n47600, n47601, n47602,
    n47603, n47604, n47605, n47606, n47607, n47608,
    n47609, n47611, n47612, n47613, n47614, n47615,
    n47616, n47617, n47618, n47619, n47620, n47621,
    n47622, n47623, n47624, n47625, n47626, n47627,
    n47628, n47629, n47630, n47631, n47632, n47633,
    n47634, n47635, n47636, n47637, n47638, n47639,
    n47640, n47641, n47642, n47643, n47644, n47646,
    n47647, n47648, n47649, n47650, n47651, n47652,
    n47653, n47654, n47655, n47656, n47657, n47658,
    n47659, n47660, n47661, n47662, n47663, n47664,
    n47665, n47666, n47667, n47668, n47669, n47670,
    n47671, n47672, n47673, n47674, n47675, n47676,
    n47677, n47678, n47680, n47681, n47682, n47683,
    n47684, n47685, n47686, n47687, n47688, n47689,
    n47690, n47691, n47692, n47693, n47694, n47695,
    n47696, n47697, n47698, n47699, n47700, n47701,
    n47702, n47703, n47704, n47705, n47706, n47707,
    n47708, n47709, n47710, n47711, n47712, n47713,
    n47715, n47716, n47717, n47719, n47720, n47721,
    n47722, n47723, n47724, n47725, n47726, n47727,
    n47728, n47729, n47730, n47731, n47732, n47733,
    n47734, n47735, n47736, n47737, n47738, n47739,
    n47740, n47741, n47742, n47743, n47744, n47745,
    n47746, n47747, n47748, n47749, n47750, n47751,
    n47752, n47753, n47755, n47756, n47757, n47758,
    n47759, n47760, n47761, n47762, n47763, n47764,
    n47765, n47766, n47767, n47768, n47769, n47770,
    n47771, n47772, n47773, n47774, n47775, n47776,
    n47777, n47778, n47779, n47780, n47781, n47782,
    n47783, n47784, n47785, n47786, n47787, n47789,
    n47790, n47791, n47792, n47793, n47794, n47795,
    n47796, n47797, n47798, n47799, n47800, n47801,
    n47802, n47803, n47804, n47805, n47806, n47807,
    n47808, n47809, n47810, n47811, n47812, n47813,
    n47814, n47815, n47816, n47817, n47818, n47819,
    n47820, n47821, n47822, n47823, n47825, n47826,
    n47827, n47828, n47829, n47830, n47831, n47832,
    n47833, n47834, n47835, n47836, n47837, n47838,
    n47839, n47840, n47841, n47842, n47843, n47844,
    n47845, n47846, n47847, n47848, n47849, n47850,
    n47851, n47852, n47853, n47854, n47855, n47856,
    n47857, n47859, n47860, n47861, n47862, n47863,
    n47864, n47865, n47866, n47867, n47868, n47869,
    n47870, n47871, n47872, n47873, n47874, n47875,
    n47876, n47877, n47878, n47879, n47880, n47881,
    n47882, n47883, n47884, n47885, n47886, n47887,
    n47888, n47889, n47890, n47891, n47892, n47894,
    n47895, n47896, n47897, n47898, n47899, n47900,
    n47901, n47902, n47903, n47904, n47905, n47906,
    n47907, n47908, n47909, n47910, n47911, n47912,
    n47913, n47914, n47915, n47916, n47917, n47918,
    n47919, n47920, n47921, n47922, n47923, n47924,
    n47925, n47926, n47927, n47928, n47929, n47930,
    n47931, n47932, n47933, n47934, n47935, n47936,
    n47937, n47938, n47939, n47940, n47941, n47942,
    n47943, n47944, n47945, n47946, n47947, n47948,
    n47950, n47951, n47952, n47953, n47954, n47955,
    n47956, n47957, n47958, n47959, n47960, n47961,
    n47962, n47963, n47964, n47965, n47966, n47967,
    n47968, n47969, n47970, n47971, n47972, n47973,
    n47974, n47975, n47976, n47977, n47978, n47979,
    n47980, n47981, n47982, n47983, n47985, n47986,
    n47987, n47989, n47990, n47991, n47993, n47994,
    n47995, n47997, n47998, n47999, n48001, n48002,
    n48003, n48005, n48006, n48007, n48009, n48010,
    n48011, n48013, n48014, n48015, n48017, n48018,
    n48019, n48020, n48021, n48022, n48023, n48024,
    n48025, n48026, n48027, n48028, n48029, n48030,
    n48031, n48032, n48034, n48035, n48036, n48038,
    n48039, n48040, n48041, n48042, n48043, n48044,
    n48045, n48046, n48047, n48048, n48049, n48050,
    n48051, n48052, n48053, n48054, n48055, n48056,
    n48057, n48058, n48059, n48060, n48061, n48062,
    n48063, n48064, n48065, n48066, n48067, n48068,
    n48069, n48070, n48071, n48072, n48074, n48075,
    n48076, n48078, n48079, n48080, n48082, n48083,
    n48084, n48086, n48087, n48088, n48090, n48091,
    n48092, n48094, n48095, n48097, n48098, n48099,
    n48101, n48102, n48103, n48105, n48106, n48107,
    n48109, n48110, n48111, n48113, n48114, n48115,
    n48117, n48118, n48119, n48121, n48122, n48123,
    n48125, n48126, n48127, n48128, n48129, n48130,
    n48131, n48132, n48133, n48134, n48135, n48136,
    n48138, n48139, n48140, n48142, n48143, n48144,
    n48146, n48147, n48148, n48150, n48151, n48152,
    n48154, n48155, n48156, n48158, n48159, n48160,
    n48162, n48163, n48164, n48166, n48167, n48168,
    n48170, n48171, n48172, n48174, n48175, n48176,
    n48178, n48179, n48180, n48182, n48183, n48184,
    n48186, n48187, n48188, n48190, n48191, n48192,
    n48194, n48195, n48196, n48198, n48199, n48200,
    n48202, n48203, n48204, n48207, n48208, n48209,
    n48210, n48211, n48212, n48213, n48214, n48215,
    n48216, n48217, n48218, n48219, n48220, n48222,
    n48223, n48225, n48226, n48227, n48229, n48230,
    n48231, n48233, n48234, n48235, n48237, n48238,
    n48239, n48240, n48241, n48242, n48243, n48244,
    n48245, n48246, n48247, n48248, n48249, n48250,
    n48251, n48252, n48253, n48255, n48256, n48257,
    n48259, n48260, n48261, n48262, n48264, n48265,
    n48266, n48268, n48269, n48270, n48271, n48272,
    n48273, n48274, n48276, n48277, n48278, n48280,
    n48281, n48282, n48283, n48284, n48285, n48286,
    n48287, n48288, n48289, n48290, n48291, n48292,
    n48293, n48294, n48295, n48297, n48298, n48299,
    n48301, n48302, n48303, n48305, n48306, n48307,
    n48308, n48309, n48310, n48311, n48315, n48316,
    n48318, n48320, n48321, n48323, n48324, n48326,
    n48327, n48329, n48330, n48332, n48333, n48335,
    n48336, n48338, n48339, n48341, n48342, n48344,
    n48345, n48347, n48348, n48350, n48351, n48352,
    n48354, n48355, n48357, n48358, n48359, n48360,
    n48361, n48362, n48363, n48364, n48366, n48367,
    n48369, n48370, n48372, n48373, n48375, n48376,
    n48378, n48379, n48381, n48382, n48384, n48385,
    n48386, n48388, n48389, n48391, n48392, n48394,
    n48395, n48397, n48398, n48400, n48401, n48403,
    n48404, n48406, n48407, n48409, n48410, n48412,
    n48413, n48415, n48416, n48418, n48420, n48422,
    n48424, n48427, n48428, n48429, n48431, n48432,
    n48433, n48434, n48435, n48436, n48437, n48438,
    n48439, n48440, n48441, n48442, n48443, n48444,
    n48445, n48446, n48447, n48448, n48449, n48450,
    n48451, n48452, n48453, n48454, n48455, n48456,
    n48457, n48458, n48460, n48461, n48462, n48463,
    n48464, n48465, n48466, n48467, n48468, n48469,
    n48470, n48471, n48472, n48473, n48474, n48475,
    n48476, n48477, n48478, n48479, n48480, n48481,
    n48482, n48483, n48484, n48485, n48486, n48488,
    n48489, n48490, n48491, n48492, n48493, n48494,
    n48495, n48496, n48497, n48498, n48499, n48500,
    n48501, n48502, n48503, n48504, n48505, n48506,
    n48507, n48508, n48509, n48510, n48511, n48512,
    n48513, n48514, n48516, n48517, n48518, n48519,
    n48520, n48521, n48522, n48523, n48524, n48525,
    n48526, n48527, n48528, n48529, n48530, n48531,
    n48532, n48533, n48534, n48535, n48536, n48537,
    n48538, n48539, n48540, n48541, n48542, n48544,
    n48545, n48547, n48549, n48550, n48552, n48555,
    n48557, n48558, n48560, n48561, n48563, n48564,
    n48566, n48567, n48570, n48571, n48573, n48574,
    n48576, n48577, n48579, n48580, n48582, n48583,
    n48585, n48586, n48588, n48589, n48591, n48592,
    n48594, n48595, n48597, n48598, n48600, n48601,
    n48603, n48604, n48606, n48607, n48609, n48610,
    n48612, n48613, n48615, n48616, n48618, n48619,
    n48621, n48622, n48624, n48625, n48627, n48628,
    n48629, n48630, n48631, n48632, n48633, n48634,
    n48636, n48637, n48639, n48640, n48642, n48643,
    n48645, n48646, n48648, n48649, n48651, n48652,
    n48654, n48655, n48657, n48658, n48659, n48660,
    n48661, n48662, n48663, n48664, n48666, n48667,
    n48669, n48670, n48672, n48673, n48675, n48676,
    n48678, n48679, n48681, n48682, n48683, n48684,
    n48685, n48686, n48687, n48688, n48690, n48691,
    n48693, n48694, n48695, n48696, n48697, n48698,
    n48699, n48700, n48702, n48703, n48704, n48705,
    n48706, n48707, n48708, n48709, n48711, n48712,
    n48713, n48714, n48715, n48716, n48717, n48718,
    n48720, n48721, n48723, n48724, n48726, n48728,
    n48729, n48731, n48732, n48734, n48735, n48737,
    n48739, n48740, n48742, n48743, n48745, n48746,
    n48748, n48749, n48751, n48752, n48754, n48755,
    n48757, n48758, n48760, n48761, n48763, n48764,
    n48766, n48768, n48769, n48771, n48772, n48774,
    n48775, n48777, n48779, n48781, n48782, n48784,
    n48785, n48786, n48787, n48788, n48789, n48790,
    n48791, n48792, n48793, n48795, n48797, n48798,
    n48800, n48801, n48803, n48804, n48806, n48808,
    n48809, n48811, n48813, n48814, n48816, n48818,
    n48819, n48821, n48822, n48824, n48825, n48827,
    n48828, n48830, n48832, n48833, n48835, n48836,
    n48838, n48839, n48841, n48842, n48844, n48845,
    n48847, n48848, n48850, n48852, n48853, n48855,
    n48856, n48858, n48859, n48861, n48863, n48865,
    n48866, n48868, n48870, n48871, n48873, n48874,
    n48876, n48878, n48879, n48881, n48883, n48884,
    n48886, n48887, n48889, n48890, n48892, n48893,
    n48896, n48898, n48900, n48901, n48904;
  assign n2437 = ~pi216 & pi833;
  assign n2438 = pi1144 & ~n2437;
  assign n2439 = pi929 & n2437;
  assign n2440 = ~pi332 & ~n2438;
  assign n2441 = ~n2439 & n2440;
  assign n2442 = pi221 & ~n2441;
  assign n2443 = pi265 & ~pi332;
  assign n2444 = pi216 & ~n2443;
  assign n2445 = pi153 & ~pi332;
  assign n2446 = ~pi105 & ~n2445;
  assign n2447 = ~pi152 & ~pi161;
  assign n2448 = ~pi166 & n2447;
  assign n2449 = pi95 & ~pi479;
  assign n2450 = ~pi40 & ~pi72;
  assign n2451 = ~pi88 & ~pi98;
  assign n2452 = ~pi77 & n2451;
  assign n2453 = ~pi50 & n2452;
  assign n2454 = ~pi102 & n2453;
  assign n2455 = ~pi65 & ~pi71;
  assign n2456 = ~pi83 & ~pi103;
  assign n2457 = ~pi67 & ~pi69;
  assign n2458 = ~pi66 & ~pi73;
  assign n2459 = ~pi61 & ~pi76;
  assign n2460 = ~pi85 & ~pi106;
  assign n2461 = n2459 & n2460;
  assign n2462 = ~pi48 & n2461;
  assign n2463 = ~pi89 & n2462;
  assign n2464 = ~pi49 & n2463;
  assign n2465 = ~pi104 & n2464;
  assign n2466 = ~pi45 & n2465;
  assign n2467 = ~pi68 & ~pi84;
  assign n2468 = ~pi82 & ~pi111;
  assign n2469 = ~pi36 & n2468;
  assign n2470 = n2467 & n2469;
  assign n2471 = n2466 & n2470;
  assign n2472 = n2458 & n2471;
  assign n2473 = n2457 & n2472;
  assign n2474 = n2456 & n2473;
  assign n2475 = n2455 & n2474;
  assign n2476 = ~pi63 & ~pi107;
  assign n2477 = n2475 & n2476;
  assign n2478 = ~pi64 & n2477;
  assign n2479 = ~pi81 & n2478;
  assign n2480 = n2454 & n2479;
  assign n2481 = ~pi53 & ~pi60;
  assign n2482 = ~pi86 & n2481;
  assign n2483 = ~pi97 & ~pi108;
  assign n2484 = ~pi94 & n2483;
  assign n2485 = ~pi46 & n2482;
  assign n2486 = n2484 & n2485;
  assign n2487 = n2480 & n2486;
  assign n2488 = ~pi109 & ~pi110;
  assign n2489 = ~pi58 & ~pi91;
  assign n2490 = ~pi47 & n2489;
  assign n2491 = n2488 & n2490;
  assign n2492 = n2487 & n2491;
  assign n2493 = ~pi90 & ~pi93;
  assign n2494 = ~pi70 & ~pi96;
  assign n2495 = ~pi35 & ~pi51;
  assign n2496 = n2494 & n2495;
  assign n2497 = n2493 & n2496;
  assign n2498 = n2492 & n2497;
  assign n2499 = n2450 & n2498;
  assign n2500 = pi225 & n2499;
  assign n2501 = pi32 & ~n2500;
  assign n2502 = ~pi95 & ~n2501;
  assign n2503 = pi60 & n2480;
  assign n2504 = ~pi53 & ~n2503;
  assign n2505 = ~pi86 & ~pi94;
  assign n2506 = ~pi60 & n2480;
  assign n2507 = pi53 & ~n2506;
  assign n2508 = n2505 & ~n2507;
  assign n2509 = ~n2504 & n2508;
  assign n2510 = ~pi46 & n2488;
  assign n2511 = ~pi47 & ~pi91;
  assign n2512 = n2483 & n2511;
  assign n2513 = n2510 & n2512;
  assign n2514 = ~pi58 & n2513;
  assign n2515 = n2493 & n2514;
  assign n2516 = n2509 & n2515;
  assign n2517 = ~pi35 & ~n2516;
  assign n2518 = ~pi58 & ~pi90;
  assign n2519 = n2486 & n2488;
  assign n2520 = n2511 & n2519;
  assign n2521 = n2480 & n2520;
  assign n2522 = n2518 & n2521;
  assign n2523 = ~pi93 & n2522;
  assign n2524 = pi35 & ~n2523;
  assign n2525 = pi35 & n2523;
  assign n2526 = ~pi225 & n2525;
  assign n2527 = ~pi70 & ~n2526;
  assign n2528 = ~pi51 & n2527;
  assign n2529 = ~n2524 & n2528;
  assign n2530 = ~n2517 & n2529;
  assign n2531 = ~pi96 & ~n2530;
  assign n2532 = ~pi47 & n2519;
  assign n2533 = n2480 & n2532;
  assign n2534 = ~pi93 & n2518;
  assign n2535 = ~pi35 & ~pi70;
  assign n2536 = ~pi51 & n2535;
  assign n2537 = ~pi91 & n2534;
  assign n2538 = n2536 & n2537;
  assign n2539 = n2533 & n2538;
  assign n2540 = pi96 & ~n2539;
  assign n2541 = n2450 & ~n2540;
  assign n2542 = ~n2531 & n2541;
  assign n2543 = ~pi32 & ~n2542;
  assign n2544 = n2502 & ~n2543;
  assign n2545 = ~n2449 & ~n2544;
  assign n2546 = ~pi137 & n2545;
  assign n2547 = ~pi35 & ~pi93;
  assign n2548 = n2522 & n2547;
  assign n2549 = ~pi72 & ~pi96;
  assign n2550 = ~pi51 & ~pi70;
  assign n2551 = n2549 & n2550;
  assign n2552 = n2548 & n2551;
  assign n2553 = pi40 & n2552;
  assign n2554 = ~pi32 & ~n2553;
  assign n2555 = pi72 & ~n2498;
  assign n2556 = ~pi40 & ~n2555;
  assign n2557 = ~pi70 & n2548;
  assign n2558 = pi51 & ~n2557;
  assign n2559 = ~pi96 & ~n2558;
  assign n2560 = ~pi51 & pi70;
  assign n2561 = n2559 & ~n2560;
  assign n2562 = ~n2524 & ~n2526;
  assign n2563 = pi93 & n2522;
  assign n2564 = ~pi35 & ~n2563;
  assign n2565 = pi91 & n2533;
  assign n2566 = n2518 & ~n2565;
  assign n2567 = ~pi109 & n2487;
  assign n2568 = pi110 & ~n2567;
  assign n2569 = pi47 & n2480;
  assign n2570 = n2519 & n2569;
  assign n2571 = pi47 & ~n2570;
  assign n2572 = ~pi91 & ~n2571;
  assign n2573 = ~n2568 & n2572;
  assign n2574 = ~pi47 & ~pi110;
  assign n2575 = pi109 & ~n2487;
  assign n2576 = ~pi102 & n2479;
  assign n2577 = n2451 & n2576;
  assign n2578 = ~pi50 & n2481;
  assign n2579 = ~pi77 & n2578;
  assign n2580 = n2505 & n2579;
  assign n2581 = n2577 & n2580;
  assign n2582 = ~pi97 & n2581;
  assign n2583 = pi108 & ~n2582;
  assign n2584 = ~pi46 & ~n2583;
  assign n2585 = pi97 & ~n2581;
  assign n2586 = n2452 & n2576;
  assign n2587 = n2578 & n2586;
  assign n2588 = ~pi86 & pi94;
  assign n2589 = n2587 & n2588;
  assign n2590 = ~pi97 & ~n2589;
  assign n2591 = pi86 & ~n2587;
  assign n2592 = ~pi94 & ~n2591;
  assign n2593 = pi77 & n2577;
  assign n2594 = ~pi50 & ~n2593;
  assign n2595 = pi81 & ~n2478;
  assign n2596 = pi102 & ~n2479;
  assign n2597 = ~n2595 & ~n2596;
  assign n2598 = pi64 & ~n2477;
  assign n2599 = pi71 & ~n2474;
  assign n2600 = ~pi65 & ~n2599;
  assign n2601 = ~pi67 & n2472;
  assign n2602 = pi69 & ~n2601;
  assign n2603 = pi83 & ~n2473;
  assign n2604 = ~pi103 & ~n2603;
  assign n2605 = ~n2602 & n2604;
  assign n2606 = ~pi69 & ~pi83;
  assign n2607 = ~pi68 & ~pi111;
  assign n2608 = n2458 & n2466;
  assign n2609 = pi84 & ~n2608;
  assign n2610 = pi85 & pi106;
  assign n2611 = n2459 & ~n2610;
  assign n2612 = pi61 & pi76;
  assign n2613 = n2460 & ~n2612;
  assign n2614 = ~n2611 & ~n2613;
  assign n2615 = ~pi48 & ~n2614;
  assign n2616 = ~n2461 & ~n2615;
  assign n2617 = pi89 & ~n2462;
  assign n2618 = ~pi49 & ~n2617;
  assign n2619 = ~n2616 & n2618;
  assign n2620 = ~n2463 & ~n2619;
  assign n2621 = pi104 & ~n2464;
  assign n2622 = ~pi45 & ~n2621;
  assign n2623 = ~n2620 & n2622;
  assign n2624 = ~n2465 & ~n2623;
  assign n2625 = ~n2466 & ~n2624;
  assign n2626 = n2458 & ~n2625;
  assign n2627 = pi66 & pi73;
  assign n2628 = ~n2458 & ~n2466;
  assign n2629 = ~n2627 & ~n2628;
  assign n2630 = ~n2626 & n2629;
  assign n2631 = ~pi84 & ~n2630;
  assign n2632 = ~n2609 & ~n2631;
  assign n2633 = n2607 & ~n2632;
  assign n2634 = ~pi84 & n2608;
  assign n2635 = ~pi68 & n2634;
  assign n2636 = pi111 & ~n2635;
  assign n2637 = ~pi82 & ~n2636;
  assign n2638 = pi68 & ~n2634;
  assign n2639 = n2637 & ~n2638;
  assign n2640 = ~n2633 & n2639;
  assign n2641 = ~pi36 & ~pi67;
  assign n2642 = pi82 & n2607;
  assign n2643 = n2634 & n2642;
  assign n2644 = n2641 & ~n2643;
  assign n2645 = ~n2640 & n2644;
  assign n2646 = pi67 & ~n2472;
  assign n2647 = n2468 & n2635;
  assign n2648 = pi36 & ~n2647;
  assign n2649 = ~n2646 & ~n2648;
  assign n2650 = ~n2645 & n2649;
  assign n2651 = n2606 & ~n2650;
  assign n2652 = n2605 & ~n2651;
  assign n2653 = pi103 & n2606;
  assign n2654 = n2601 & n2653;
  assign n2655 = ~pi71 & ~n2654;
  assign n2656 = ~n2652 & n2655;
  assign n2657 = n2600 & ~n2656;
  assign n2658 = ~pi107 & ~n2657;
  assign n2659 = pi65 & ~pi71;
  assign n2660 = n2474 & n2659;
  assign n2661 = n2658 & ~n2660;
  assign n2662 = ~pi63 & pi107;
  assign n2663 = n2475 & n2662;
  assign n2664 = ~n2476 & ~n2663;
  assign n2665 = ~n2661 & ~n2664;
  assign n2666 = ~pi64 & ~n2665;
  assign n2667 = ~n2598 & ~n2666;
  assign n2668 = ~pi81 & ~pi102;
  assign n2669 = ~n2667 & n2668;
  assign n2670 = ~n2658 & ~n2664;
  assign n2671 = pi63 & ~pi107;
  assign n2672 = n2475 & n2671;
  assign n2673 = ~pi64 & ~n2672;
  assign n2674 = ~n2670 & n2673;
  assign n2675 = ~n2598 & ~n2674;
  assign n2676 = n2669 & ~n2675;
  assign n2677 = n2597 & ~n2676;
  assign n2678 = n2451 & ~n2677;
  assign n2679 = ~pi98 & n2576;
  assign n2680 = pi88 & ~n2679;
  assign n2681 = pi98 & ~n2576;
  assign n2682 = ~pi77 & ~n2681;
  assign n2683 = ~n2680 & n2682;
  assign n2684 = ~n2678 & n2683;
  assign n2685 = n2594 & ~n2684;
  assign n2686 = pi50 & ~n2586;
  assign n2687 = ~pi60 & ~n2686;
  assign n2688 = ~n2685 & n2687;
  assign n2689 = n2504 & ~n2688;
  assign n2690 = ~n2507 & ~n2689;
  assign n2691 = ~pi86 & ~n2690;
  assign n2692 = n2592 & ~n2691;
  assign n2693 = n2590 & ~n2692;
  assign n2694 = ~n2585 & ~n2693;
  assign n2695 = ~pi108 & ~n2694;
  assign n2696 = n2584 & ~n2695;
  assign n2697 = pi46 & n2483;
  assign n2698 = n2581 & n2697;
  assign n2699 = ~pi109 & ~n2698;
  assign n2700 = ~n2696 & n2699;
  assign n2701 = ~n2575 & ~n2700;
  assign n2702 = n2574 & ~n2701;
  assign n2703 = n2573 & ~n2702;
  assign n2704 = n2566 & ~n2703;
  assign n2705 = pi58 & ~n2521;
  assign n2706 = pi90 & ~n2492;
  assign n2707 = ~pi93 & ~n2706;
  assign n2708 = ~n2705 & n2707;
  assign n2709 = ~n2704 & n2708;
  assign n2710 = n2564 & ~n2709;
  assign n2711 = n2562 & ~n2710;
  assign n2712 = ~pi51 & ~n2711;
  assign n2713 = n2561 & ~n2712;
  assign n2714 = ~pi72 & ~n2713;
  assign n2715 = n2556 & ~n2714;
  assign n2716 = n2554 & ~n2715;
  assign n2717 = pi96 & n2539;
  assign n2718 = ~pi51 & ~pi72;
  assign n2719 = ~pi40 & n2718;
  assign n2720 = n2548 & n2719;
  assign n2721 = n2717 & n2720;
  assign n2722 = n2716 & ~n2721;
  assign n2723 = ~n2501 & ~n2722;
  assign n2724 = ~pi95 & ~n2723;
  assign n2725 = ~pi32 & ~pi40;
  assign n2726 = n2552 & n2725;
  assign n2727 = pi95 & ~n2726;
  assign n2728 = pi479 & n2727;
  assign n2729 = ~n2724 & ~n2728;
  assign n2730 = pi137 & ~n2729;
  assign n2731 = ~n2546 & ~n2730;
  assign n2732 = pi210 & ~n2731;
  assign n2733 = ~pi833 & pi957;
  assign n2734 = pi1091 & ~n2733;
  assign n2735 = pi841 & n2522;
  assign n2736 = ~pi93 & n2735;
  assign n2737 = n2718 & n2736;
  assign n2738 = ~pi35 & ~pi40;
  assign n2739 = pi225 & n2738;
  assign n2740 = n2494 & n2739;
  assign n2741 = n2737 & n2740;
  assign n2742 = pi32 & ~n2741;
  assign n2743 = ~n2722 & ~n2742;
  assign n2744 = ~pi95 & ~n2743;
  assign n2745 = ~n2728 & ~n2744;
  assign n2746 = pi137 & ~n2745;
  assign n2747 = pi95 & pi479;
  assign n2748 = ~n2543 & ~n2742;
  assign n2749 = ~pi95 & ~n2748;
  assign n2750 = ~n2747 & ~n2749;
  assign n2751 = ~pi137 & ~n2750;
  assign n2752 = ~n2746 & ~n2751;
  assign n2753 = ~n2734 & n2752;
  assign n2754 = pi829 & pi950;
  assign n2755 = pi1092 & pi1093;
  assign n2756 = n2754 & n2755;
  assign n2757 = n2750 & ~n2756;
  assign n2758 = ~pi108 & ~n2585;
  assign n2759 = ~pi110 & n2758;
  assign n2760 = ~pi97 & ~n2509;
  assign n2761 = ~pi46 & ~pi109;
  assign n2762 = n2511 & n2761;
  assign n2763 = n2534 & n2762;
  assign n2764 = n2759 & n2763;
  assign n2765 = ~n2760 & n2764;
  assign n2766 = ~pi35 & ~n2765;
  assign n2767 = n2529 & ~n2766;
  assign n2768 = ~pi96 & ~n2767;
  assign n2769 = n2541 & ~n2768;
  assign n2770 = ~pi32 & ~n2769;
  assign n2771 = ~n2742 & ~n2770;
  assign n2772 = ~pi95 & ~n2771;
  assign n2773 = ~n2747 & n2756;
  assign n2774 = ~n2772 & n2773;
  assign n2775 = ~pi137 & ~n2774;
  assign n2776 = ~n2757 & n2775;
  assign n2777 = n2734 & ~n2776;
  assign n2778 = ~n2746 & n2777;
  assign n2779 = ~n2753 & ~n2778;
  assign n2780 = ~pi210 & n2779;
  assign n2781 = ~n2732 & ~n2780;
  assign n2782 = pi234 & n2781;
  assign n2783 = ~pi40 & n2549;
  assign n2784 = n2530 & n2783;
  assign n2785 = ~pi32 & ~n2784;
  assign n2786 = n2502 & ~n2785;
  assign n2787 = ~pi137 & ~n2786;
  assign n2788 = ~n2449 & ~n2727;
  assign n2789 = ~n2501 & ~n2716;
  assign n2790 = ~pi95 & ~n2789;
  assign n2791 = n2788 & ~n2790;
  assign n2792 = pi137 & ~n2791;
  assign n2793 = ~n2787 & ~n2792;
  assign n2794 = pi210 & ~n2793;
  assign n2795 = ~pi95 & ~n2742;
  assign n2796 = n2734 & n2756;
  assign n2797 = ~n2517 & ~n2796;
  assign n2798 = ~n2766 & n2796;
  assign n2799 = ~n2797 & ~n2798;
  assign n2800 = n2529 & n2783;
  assign n2801 = ~n2799 & n2800;
  assign n2802 = ~pi32 & ~n2801;
  assign n2803 = n2795 & ~n2802;
  assign n2804 = ~pi137 & ~n2803;
  assign n2805 = ~n2716 & ~n2742;
  assign n2806 = ~pi95 & ~n2805;
  assign n2807 = n2788 & ~n2806;
  assign n2808 = pi137 & ~n2807;
  assign n2809 = ~n2804 & ~n2808;
  assign n2810 = ~pi210 & ~n2809;
  assign n2811 = ~n2794 & ~n2810;
  assign n2812 = ~pi234 & n2811;
  assign n2813 = ~pi332 & ~n2812;
  assign n2814 = ~n2782 & n2813;
  assign n2815 = n2448 & ~n2814;
  assign n2816 = pi146 & n2781;
  assign n2817 = pi234 & ~pi332;
  assign n2818 = ~pi210 & ~n2752;
  assign n2819 = ~pi146 & ~n2732;
  assign n2820 = ~n2818 & n2819;
  assign n2821 = n2817 & ~n2820;
  assign n2822 = ~n2816 & n2821;
  assign n2823 = pi146 & n2811;
  assign n2824 = ~n2785 & n2795;
  assign n2825 = ~pi137 & ~n2824;
  assign n2826 = ~n2808 & ~n2825;
  assign n2827 = ~pi210 & ~n2826;
  assign n2828 = ~pi146 & ~n2794;
  assign n2829 = ~n2827 & n2828;
  assign n2830 = ~pi234 & ~pi332;
  assign n2831 = ~n2823 & n2830;
  assign n2832 = ~n2829 & n2831;
  assign n2833 = ~n2448 & ~n2832;
  assign n2834 = ~n2822 & n2833;
  assign n2835 = ~n2815 & ~n2834;
  assign n2836 = pi105 & ~n2835;
  assign n2837 = ~n2446 & ~n2836;
  assign n2838 = pi228 & ~n2837;
  assign n2839 = ~pi109 & ~n2696;
  assign n2840 = ~n2575 & ~n2839;
  assign n2841 = n2574 & ~n2840;
  assign n2842 = n2573 & ~n2841;
  assign n2843 = n2566 & ~n2842;
  assign n2844 = n2708 & ~n2843;
  assign n2845 = n2564 & ~n2844;
  assign n2846 = n2562 & ~n2845;
  assign n2847 = ~pi51 & ~n2846;
  assign n2848 = n2561 & ~n2847;
  assign n2849 = ~pi72 & ~n2848;
  assign n2850 = n2556 & ~n2849;
  assign n2851 = n2554 & ~n2850;
  assign n2852 = ~n2721 & n2851;
  assign n2853 = ~n2742 & ~n2852;
  assign n2854 = ~pi95 & ~n2853;
  assign n2855 = ~n2727 & ~n2854;
  assign n2856 = pi137 & ~n2855;
  assign n2857 = ~pi146 & ~n2448;
  assign n2858 = n2734 & ~n2857;
  assign n2859 = ~n2757 & n2858;
  assign n2860 = ~n2727 & n2750;
  assign n2861 = ~n2859 & n2860;
  assign n2862 = ~n2727 & n2858;
  assign n2863 = n2774 & n2862;
  assign n2864 = ~pi137 & ~n2863;
  assign n2865 = ~n2861 & n2864;
  assign n2866 = ~n2856 & ~n2865;
  assign n2867 = ~pi210 & ~n2866;
  assign n2868 = pi234 & ~n2867;
  assign n2869 = ~n2742 & ~n2851;
  assign n2870 = ~pi95 & ~n2869;
  assign n2871 = n2788 & ~n2870;
  assign n2872 = pi137 & ~n2871;
  assign n2873 = n2804 & ~n2857;
  assign n2874 = n2825 & n2857;
  assign n2875 = ~pi210 & ~pi234;
  assign n2876 = ~n2874 & n2875;
  assign n2877 = ~n2873 & n2876;
  assign n2878 = ~n2872 & n2877;
  assign n2879 = ~n2501 & ~n2851;
  assign n2880 = ~pi95 & ~n2879;
  assign n2881 = n2788 & ~n2880;
  assign n2882 = pi137 & ~n2881;
  assign n2883 = pi210 & ~n2787;
  assign n2884 = ~n2882 & n2883;
  assign n2885 = ~n2878 & ~n2884;
  assign n2886 = ~n2868 & n2885;
  assign n2887 = ~n2501 & ~n2852;
  assign n2888 = ~pi95 & ~n2887;
  assign n2889 = pi137 & ~n2727;
  assign n2890 = ~n2888 & n2889;
  assign n2891 = ~pi137 & ~n2727;
  assign n2892 = ~n2545 & n2891;
  assign n2893 = pi210 & pi234;
  assign n2894 = ~n2892 & n2893;
  assign n2895 = ~n2890 & n2894;
  assign n2896 = ~n2886 & ~n2895;
  assign n2897 = n2445 & ~n2896;
  assign n2898 = pi93 & ~n2522;
  assign n2899 = ~pi35 & ~n2898;
  assign n2900 = ~n2705 & ~n2706;
  assign n2901 = ~pi53 & n2688;
  assign n2902 = ~pi86 & ~n2901;
  assign n2903 = n2592 & ~n2902;
  assign n2904 = n2590 & ~n2903;
  assign n2905 = ~n2585 & ~n2904;
  assign n2906 = ~pi108 & ~n2905;
  assign n2907 = n2584 & ~n2906;
  assign n2908 = ~pi109 & ~n2907;
  assign n2909 = ~n2575 & ~n2908;
  assign n2910 = n2574 & ~n2909;
  assign n2911 = n2573 & ~n2910;
  assign n2912 = n2566 & ~n2911;
  assign n2913 = n2900 & ~n2912;
  assign n2914 = ~pi93 & ~n2913;
  assign n2915 = n2899 & ~n2914;
  assign n2916 = n2528 & ~n2915;
  assign n2917 = pi70 & ~n2548;
  assign n2918 = n2559 & ~n2917;
  assign n2919 = ~n2916 & n2918;
  assign n2920 = ~pi72 & ~n2717;
  assign n2921 = ~n2919 & n2920;
  assign n2922 = n2556 & ~n2921;
  assign n2923 = n2554 & ~n2922;
  assign n2924 = ~n2796 & n2923;
  assign n2925 = pi225 & pi841;
  assign n2926 = n2499 & ~n2925;
  assign n2927 = pi32 & ~n2926;
  assign n2928 = n2554 & n2796;
  assign n2929 = ~pi97 & ~n2904;
  assign n2930 = ~pi108 & ~n2929;
  assign n2931 = n2584 & ~n2930;
  assign n2932 = ~pi109 & ~n2931;
  assign n2933 = ~n2575 & ~n2932;
  assign n2934 = n2574 & ~n2933;
  assign n2935 = n2573 & ~n2934;
  assign n2936 = n2566 & ~n2935;
  assign n2937 = n2900 & ~n2936;
  assign n2938 = ~pi93 & ~n2937;
  assign n2939 = n2899 & ~n2938;
  assign n2940 = n2528 & ~n2939;
  assign n2941 = n2918 & ~n2940;
  assign n2942 = n2920 & ~n2941;
  assign n2943 = n2556 & ~n2942;
  assign n2944 = n2928 & ~n2943;
  assign n2945 = ~n2927 & ~n2944;
  assign n2946 = ~n2924 & n2945;
  assign n2947 = ~pi95 & ~n2946;
  assign n2948 = ~n2727 & ~n2947;
  assign n2949 = ~pi137 & ~n2948;
  assign n2950 = ~pi95 & ~n2927;
  assign n2951 = ~pi51 & ~pi96;
  assign n2952 = ~n2917 & n2951;
  assign n2953 = n2450 & n2952;
  assign n2954 = ~n2527 & n2953;
  assign n2955 = ~pi32 & ~n2954;
  assign n2956 = ~pi72 & n2725;
  assign n2957 = n2717 & n2956;
  assign n2958 = n2955 & ~n2957;
  assign n2959 = n2950 & ~n2958;
  assign n2960 = n2449 & n2726;
  assign n2961 = pi137 & ~n2960;
  assign n2962 = ~n2959 & n2961;
  assign n2963 = ~n2949 & ~n2962;
  assign n2964 = ~pi210 & ~n2963;
  assign n2965 = pi146 & n2964;
  assign n2966 = ~pi225 & n2499;
  assign n2967 = pi32 & ~n2966;
  assign n2968 = ~n2923 & ~n2967;
  assign n2969 = ~pi95 & ~n2968;
  assign n2970 = n2891 & ~n2969;
  assign n2971 = ~pi95 & ~n2967;
  assign n2972 = ~n2958 & n2971;
  assign n2973 = ~n2960 & ~n2972;
  assign n2974 = pi137 & ~n2973;
  assign n2975 = pi210 & ~n2974;
  assign n2976 = ~n2970 & n2975;
  assign n2977 = n2830 & ~n2976;
  assign n2978 = ~pi146 & ~pi210;
  assign n2979 = ~n2923 & ~n2927;
  assign n2980 = ~pi95 & ~n2979;
  assign n2981 = ~n2727 & ~n2980;
  assign n2982 = ~pi137 & ~n2981;
  assign n2983 = ~n2962 & ~n2982;
  assign n2984 = n2978 & ~n2983;
  assign n2985 = n2977 & ~n2984;
  assign n2986 = ~n2965 & n2985;
  assign n2987 = n2950 & ~n2955;
  assign n2988 = pi137 & ~n2987;
  assign n2989 = ~pi72 & ~n2919;
  assign n2990 = n2556 & ~n2989;
  assign n2991 = n2554 & ~n2990;
  assign n2992 = ~n2796 & n2991;
  assign n2993 = ~pi72 & ~n2941;
  assign n2994 = n2556 & ~n2993;
  assign n2995 = n2928 & ~n2994;
  assign n2996 = ~n2927 & ~n2995;
  assign n2997 = ~n2992 & n2996;
  assign n2998 = ~pi95 & ~n2997;
  assign n2999 = n2788 & ~n2998;
  assign n3000 = ~pi137 & ~n2999;
  assign n3001 = ~n2988 & ~n3000;
  assign n3002 = ~pi210 & ~n3001;
  assign n3003 = pi146 & n3002;
  assign n3004 = ~n2967 & ~n2991;
  assign n3005 = ~pi95 & ~n3004;
  assign n3006 = ~pi137 & n2788;
  assign n3007 = ~n3005 & n3006;
  assign n3008 = pi137 & n2971;
  assign n3009 = ~n2955 & n3008;
  assign n3010 = pi210 & ~n3009;
  assign n3011 = ~n3007 & n3010;
  assign n3012 = n2817 & ~n3011;
  assign n3013 = ~n2927 & ~n2991;
  assign n3014 = ~pi95 & ~n3013;
  assign n3015 = n2788 & ~n3014;
  assign n3016 = ~pi137 & ~n3015;
  assign n3017 = ~n2988 & ~n3016;
  assign n3018 = n2978 & ~n3017;
  assign n3019 = n3012 & ~n3018;
  assign n3020 = ~n3003 & n3019;
  assign n3021 = ~n2448 & ~n2986;
  assign n3022 = ~n3020 & n3021;
  assign n3023 = ~n3002 & n3012;
  assign n3024 = ~n2964 & n2977;
  assign n3025 = n2448 & ~n3023;
  assign n3026 = ~n3024 & n3025;
  assign n3027 = ~pi153 & ~n3026;
  assign n3028 = ~n3022 & n3027;
  assign n3029 = ~pi228 & ~n2897;
  assign n3030 = ~n3028 & n3029;
  assign n3031 = ~n2838 & ~n3030;
  assign n3032 = ~pi216 & ~n3031;
  assign n3033 = ~n2444 & ~n3032;
  assign n3034 = ~pi221 & ~n3033;
  assign n3035 = ~n2442 & ~n3034;
  assign n3036 = ~pi215 & ~n3035;
  assign n3037 = ~pi332 & ~pi1144;
  assign n3038 = pi215 & ~n3037;
  assign n3039 = pi299 & ~n3038;
  assign n3040 = ~n3036 & n3039;
  assign n3041 = ~pi224 & pi833;
  assign n3042 = pi222 & ~n3041;
  assign n3043 = ~pi223 & ~n3042;
  assign n3044 = n3037 & ~n3043;
  assign n3045 = pi224 & ~n2443;
  assign n3046 = ~pi222 & ~n3045;
  assign n3047 = ~pi332 & ~pi929;
  assign n3048 = n3041 & n3047;
  assign n3049 = ~n3046 & ~n3048;
  assign n3050 = ~pi223 & ~n3049;
  assign n3051 = ~n3044 & ~n3050;
  assign n3052 = ~pi299 & ~n3051;
  assign n3053 = ~pi222 & ~pi224;
  assign n3054 = pi198 & ~n2731;
  assign n3055 = ~pi198 & n2779;
  assign n3056 = ~n3054 & ~n3055;
  assign n3057 = pi142 & n3056;
  assign n3058 = ~pi198 & ~n2752;
  assign n3059 = ~pi142 & ~n3054;
  assign n3060 = ~n3058 & n3059;
  assign n3061 = n2817 & ~n3060;
  assign n3062 = ~n3057 & n3061;
  assign n3063 = ~pi144 & ~pi174;
  assign n3064 = ~pi189 & n3063;
  assign n3065 = ~pi223 & ~n3064;
  assign n3066 = pi198 & ~n2793;
  assign n3067 = ~pi198 & ~n2809;
  assign n3068 = ~n3066 & ~n3067;
  assign n3069 = pi142 & n3068;
  assign n3070 = ~pi198 & ~n2826;
  assign n3071 = ~pi142 & ~n3066;
  assign n3072 = ~n3070 & n3071;
  assign n3073 = n2830 & ~n3069;
  assign n3074 = ~n3072 & n3073;
  assign n3075 = n3065 & ~n3074;
  assign n3076 = ~n3062 & n3075;
  assign n3077 = ~pi223 & n3064;
  assign n3078 = pi234 & n3056;
  assign n3079 = ~pi234 & n3068;
  assign n3080 = ~pi332 & ~n3079;
  assign n3081 = ~n3078 & n3080;
  assign n3082 = n3077 & ~n3081;
  assign n3083 = ~n3076 & ~n3082;
  assign n3084 = n3053 & ~n3083;
  assign n3085 = n3052 & ~n3084;
  assign n3086 = ~pi39 & ~n3085;
  assign n3087 = ~n3040 & n3086;
  assign n3088 = pi234 & n2449;
  assign n3089 = ~pi332 & ~n3088;
  assign n3090 = ~pi95 & n2726;
  assign n3091 = ~n2449 & ~n3090;
  assign n3092 = pi234 & ~n3091;
  assign n3093 = ~pi32 & ~pi95;
  assign n3094 = n2450 & n3093;
  assign n3095 = n2951 & n3094;
  assign n3096 = n2557 & n3095;
  assign n3097 = ~pi234 & n3096;
  assign n3098 = ~n3092 & ~n3097;
  assign n3099 = pi137 & ~n3098;
  assign n3100 = n3089 & ~n3099;
  assign n3101 = ~pi223 & n3053;
  assign n3102 = ~n3100 & n3101;
  assign n3103 = ~n3051 & ~n3102;
  assign n3104 = ~pi299 & ~n3103;
  assign n3105 = pi105 & ~n3100;
  assign n3106 = ~n2446 & ~n3105;
  assign n3107 = pi228 & ~n3106;
  assign n3108 = ~pi332 & n3090;
  assign n3109 = ~pi137 & ~pi153;
  assign n3110 = n3108 & n3109;
  assign n3111 = pi137 & n3096;
  assign n3112 = n2445 & ~n3111;
  assign n3113 = ~pi228 & ~n3112;
  assign n3114 = ~n3110 & n3113;
  assign n3115 = ~n3107 & ~n3114;
  assign n3116 = ~pi216 & ~n3115;
  assign n3117 = ~n2444 & ~n3116;
  assign n3118 = ~pi221 & ~n3117;
  assign n3119 = ~n2442 & ~n3118;
  assign n3120 = ~pi215 & ~n3119;
  assign n3121 = ~n3038 & ~n3120;
  assign n3122 = pi299 & ~n3121;
  assign n3123 = ~n3104 & ~n3122;
  assign n3124 = pi39 & ~n3123;
  assign n3125 = ~pi38 & ~n3124;
  assign n3126 = ~n3087 & n3125;
  assign n3127 = pi105 & pi228;
  assign n3128 = n3089 & n3127;
  assign n3129 = n2445 & ~n3127;
  assign n3130 = ~pi216 & ~n3129;
  assign n3131 = ~n3128 & n3130;
  assign n3132 = ~n2444 & ~n3131;
  assign n3133 = ~pi221 & ~n3132;
  assign n3134 = ~n2442 & ~n3133;
  assign n3135 = ~pi215 & ~n3134;
  assign n3136 = ~n3038 & ~n3135;
  assign n3137 = ~pi215 & ~pi221;
  assign n3138 = n3130 & n3137;
  assign n3139 = ~n3100 & n3138;
  assign n3140 = n3136 & ~n3139;
  assign n3141 = pi299 & ~n3140;
  assign n3142 = ~n3104 & ~n3141;
  assign n3143 = ~pi39 & ~n3142;
  assign n3144 = pi299 & n3136;
  assign n3145 = ~n3089 & n3101;
  assign n3146 = n3052 & ~n3145;
  assign n3147 = ~n3144 & ~n3146;
  assign n3148 = pi39 & n3147;
  assign n3149 = pi38 & ~n3148;
  assign n3150 = ~n3143 & n3149;
  assign n3151 = ~pi100 & ~n3150;
  assign n3152 = ~n3126 & n3151;
  assign n3153 = pi228 & ~n2446;
  assign n3154 = ~pi210 & ~n2857;
  assign n3155 = pi95 & pi234;
  assign n3156 = ~pi137 & ~n3155;
  assign n3157 = ~n3154 & n3156;
  assign n3158 = ~n3098 & ~n3157;
  assign n3159 = ~pi332 & ~n3158;
  assign n3160 = pi105 & ~n3159;
  assign n3161 = n3153 & ~n3160;
  assign n3162 = ~pi137 & pi210;
  assign n3163 = ~pi252 & ~n3162;
  assign n3164 = ~n2857 & n3163;
  assign n3165 = n3108 & n3164;
  assign n3166 = n2857 & n3111;
  assign n3167 = n2445 & ~n3166;
  assign n3168 = ~n3165 & n3167;
  assign n3169 = pi252 & ~n2857;
  assign n3170 = ~n3154 & ~n3169;
  assign n3171 = n3110 & n3170;
  assign n3172 = ~n3168 & ~n3171;
  assign n3173 = ~pi228 & ~n3172;
  assign n3174 = ~pi216 & ~n3173;
  assign n3175 = ~n3161 & n3174;
  assign n3176 = ~n2444 & ~n3175;
  assign n3177 = ~pi221 & ~n3176;
  assign n3178 = ~n2442 & ~n3177;
  assign n3179 = ~pi215 & ~n3178;
  assign n3180 = ~n3038 & ~n3179;
  assign n3181 = pi299 & ~n3180;
  assign n3182 = ~pi38 & ~pi39;
  assign n3183 = pi142 & ~pi198;
  assign n3184 = ~pi137 & ~n3183;
  assign n3185 = ~n3098 & ~n3184;
  assign n3186 = n3089 & ~n3185;
  assign n3187 = n3065 & ~n3186;
  assign n3188 = ~pi137 & pi198;
  assign n3189 = ~pi95 & n3188;
  assign n3190 = ~n3091 & ~n3189;
  assign n3191 = n2817 & ~n3190;
  assign n3192 = n3096 & ~n3188;
  assign n3193 = n2830 & ~n3192;
  assign n3194 = n3077 & ~n3193;
  assign n3195 = ~n3191 & n3194;
  assign n3196 = ~n3187 & ~n3195;
  assign n3197 = n3053 & ~n3196;
  assign n3198 = ~n3051 & ~n3197;
  assign n3199 = ~pi299 & ~n3198;
  assign n3200 = n3182 & ~n3199;
  assign n3201 = ~n3181 & n3200;
  assign n3202 = ~n3147 & ~n3182;
  assign n3203 = pi100 & ~n3202;
  assign n3204 = ~n3201 & n3203;
  assign n3205 = ~pi87 & ~n3204;
  assign n3206 = ~n3152 & n3205;
  assign n3207 = ~pi38 & ~pi100;
  assign n3208 = ~pi39 & n3207;
  assign n3209 = ~n3147 & ~n3208;
  assign n3210 = n3123 & n3208;
  assign n3211 = ~n3209 & ~n3210;
  assign n3212 = pi87 & ~n3211;
  assign n3213 = ~pi75 & ~n3212;
  assign n3214 = ~n3206 & n3213;
  assign n3215 = n3130 & ~n3161;
  assign n3216 = ~n2444 & ~n3215;
  assign n3217 = ~pi221 & ~n3216;
  assign n3218 = ~n2442 & ~n3217;
  assign n3219 = ~pi215 & ~n3218;
  assign n3220 = ~n3038 & ~n3219;
  assign n3221 = pi299 & ~n3220;
  assign n3222 = ~pi39 & ~pi87;
  assign n3223 = n3207 & n3222;
  assign n3224 = ~n3199 & n3223;
  assign n3225 = ~n3221 & n3224;
  assign n3226 = ~n3147 & ~n3223;
  assign n3227 = pi75 & ~n3226;
  assign n3228 = ~n3225 & n3227;
  assign n3229 = ~n3214 & ~n3228;
  assign n3230 = ~pi92 & ~n3229;
  assign n3231 = ~pi75 & ~pi87;
  assign n3232 = ~n3211 & n3231;
  assign n3233 = ~n3147 & ~n3231;
  assign n3234 = pi92 & ~n3233;
  assign n3235 = ~n3232 & n3234;
  assign n3236 = ~pi54 & ~n3235;
  assign n3237 = ~n3230 & n3236;
  assign n3238 = ~pi75 & ~pi92;
  assign n3239 = n3223 & n3238;
  assign n3240 = n3147 & ~n3239;
  assign n3241 = ~pi87 & ~pi100;
  assign n3242 = ~pi38 & n3241;
  assign n3243 = n3238 & n3242;
  assign n3244 = n3143 & n3243;
  assign n3245 = ~n3240 & ~n3244;
  assign n3246 = pi54 & n3245;
  assign n3247 = ~pi74 & ~n3246;
  assign n3248 = ~n3237 & n3247;
  assign n3249 = ~pi54 & n3245;
  assign n3250 = pi54 & ~n3147;
  assign n3251 = pi74 & ~n3250;
  assign n3252 = ~n3249 & n3251;
  assign n3253 = ~n3248 & ~n3252;
  assign n3254 = ~pi55 & ~n3253;
  assign n3255 = ~pi332 & n3098;
  assign n3256 = pi105 & ~n3255;
  assign n3257 = n3153 & ~n3256;
  assign n3258 = ~pi228 & n2445;
  assign n3259 = ~n3096 & n3258;
  assign n3260 = ~pi216 & ~n3259;
  assign n3261 = ~n3257 & n3260;
  assign n3262 = ~n2444 & ~n3261;
  assign n3263 = ~pi221 & ~n3262;
  assign n3264 = ~n2442 & ~n3263;
  assign n3265 = ~pi215 & ~n3264;
  assign n3266 = ~pi54 & ~pi74;
  assign n3267 = n3238 & n3266;
  assign n3268 = n3241 & n3267;
  assign n3269 = n3182 & n3268;
  assign n3270 = ~n3038 & n3269;
  assign n3271 = ~n3265 & n3270;
  assign n3272 = n3136 & ~n3269;
  assign n3273 = pi55 & ~n3272;
  assign n3274 = ~n3271 & n3273;
  assign n3275 = ~pi56 & ~n3274;
  assign n3276 = ~n3254 & n3275;
  assign n3277 = ~pi100 & n3182;
  assign n3278 = ~pi92 & n3231;
  assign n3279 = n3266 & n3278;
  assign n3280 = ~pi55 & n3279;
  assign n3281 = n3277 & n3280;
  assign n3282 = n3136 & ~n3281;
  assign n3283 = n3121 & n3281;
  assign n3284 = ~n3282 & ~n3283;
  assign n3285 = pi56 & ~n3284;
  assign n3286 = ~pi62 & ~n3285;
  assign n3287 = ~n3276 & n3286;
  assign n3288 = ~pi56 & ~n3284;
  assign n3289 = pi56 & n3136;
  assign n3290 = pi62 & ~n3289;
  assign n3291 = ~n3288 & n3290;
  assign n3292 = ~pi59 & ~n3291;
  assign n3293 = ~n3287 & n3292;
  assign n3294 = ~pi56 & ~pi62;
  assign n3295 = n3281 & n3294;
  assign n3296 = n3139 & n3295;
  assign n3297 = pi59 & n3136;
  assign n3298 = ~n3296 & n3297;
  assign n3299 = ~pi57 & ~n3298;
  assign n3300 = ~n3293 & n3299;
  assign n3301 = ~pi59 & n3296;
  assign n3302 = n3136 & ~n3301;
  assign n3303 = pi57 & ~n3302;
  assign po153 = n3300 | n3303;
  assign n3305 = ~pi222 & pi224;
  assign n3306 = pi276 & n3305;
  assign n3307 = ~pi1146 & ~n3041;
  assign n3308 = ~pi939 & n3041;
  assign n3309 = pi222 & ~n3307;
  assign n3310 = ~n3308 & n3309;
  assign n3311 = ~pi223 & ~n3310;
  assign n3312 = ~n3306 & n3311;
  assign n3313 = pi223 & ~pi1146;
  assign n3314 = ~pi299 & ~n3313;
  assign n3315 = ~n3312 & n3314;
  assign n3316 = pi215 & pi1146;
  assign n3317 = ~pi1146 & ~n2437;
  assign n3318 = ~pi939 & n2437;
  assign n3319 = pi221 & ~n3317;
  assign n3320 = ~n3318 & n3319;
  assign n3321 = ~n3316 & ~n3320;
  assign n3322 = ~pi228 & n3096;
  assign n3323 = ~pi216 & n3322;
  assign n3324 = n3321 & n3323;
  assign n3325 = pi216 & ~pi221;
  assign n3326 = pi276 & n3325;
  assign n3327 = ~pi216 & ~n3127;
  assign n3328 = ~n3326 & ~n3327;
  assign n3329 = ~pi221 & ~n3328;
  assign n3330 = ~n3320 & ~n3329;
  assign n3331 = ~pi215 & ~n3330;
  assign n3332 = ~n3316 & ~n3331;
  assign n3333 = pi299 & ~n3332;
  assign n3334 = ~n3324 & n3333;
  assign n3335 = ~n3315 & ~n3334;
  assign n3336 = ~pi154 & ~n3335;
  assign n3337 = ~n3320 & ~n3326;
  assign n3338 = ~pi215 & ~n3337;
  assign n3339 = ~n3316 & ~n3338;
  assign n3340 = pi299 & ~n3339;
  assign n3341 = ~n3315 & ~n3340;
  assign n3342 = pi154 & ~n3341;
  assign n3343 = n3208 & ~n3342;
  assign n3344 = ~n3336 & n3343;
  assign n3345 = pi154 & ~n3339;
  assign n3346 = ~pi154 & ~n3332;
  assign n3347 = ~n3345 & ~n3346;
  assign n3348 = pi299 & ~n3347;
  assign n3349 = ~n3315 & ~n3348;
  assign n3350 = ~n3208 & n3349;
  assign n3351 = ~n3344 & ~n3350;
  assign n3352 = pi87 & ~n3351;
  assign n3353 = pi39 & ~n3096;
  assign n3354 = ~pi70 & n2845;
  assign n3355 = ~n2524 & ~n2917;
  assign n3356 = ~n3354 & n3355;
  assign n3357 = ~pi51 & ~n3356;
  assign n3358 = n2559 & ~n3357;
  assign n3359 = n2920 & ~n3358;
  assign n3360 = ~n2555 & ~n3359;
  assign n3361 = n2725 & ~n3360;
  assign n3362 = pi40 & ~n2552;
  assign n3363 = pi32 & ~n2499;
  assign n3364 = ~n3362 & ~n3363;
  assign n3365 = ~n3361 & n3364;
  assign n3366 = ~pi95 & ~n3365;
  assign n3367 = ~n2727 & ~n3366;
  assign n3368 = ~pi39 & ~n3367;
  assign n3369 = ~n3353 & ~n3368;
  assign n3370 = ~pi216 & ~pi228;
  assign n3371 = n3321 & n3370;
  assign n3372 = n3369 & n3371;
  assign n3373 = n3333 & ~n3372;
  assign n3374 = ~n3315 & ~n3373;
  assign n3375 = ~pi154 & ~n3374;
  assign n3376 = ~pi38 & ~n3342;
  assign n3377 = ~n3375 & n3376;
  assign n3378 = pi38 & n3349;
  assign n3379 = ~pi100 & ~n3378;
  assign n3380 = ~n3377 & n3379;
  assign n3381 = ~pi146 & ~n3096;
  assign n3382 = ~pi252 & n3096;
  assign n3383 = pi146 & ~n3382;
  assign n3384 = ~n3381 & ~n3383;
  assign n3385 = pi152 & ~n3384;
  assign n3386 = ~pi161 & ~pi166;
  assign n3387 = n3384 & ~n3386;
  assign n3388 = n3382 & n3386;
  assign n3389 = ~pi152 & ~n3388;
  assign n3390 = ~n3387 & n3389;
  assign n3391 = ~n3385 & ~n3390;
  assign n3392 = ~pi38 & ~pi216;
  assign n3393 = ~pi228 & n3392;
  assign n3394 = ~pi154 & pi299;
  assign n3395 = ~pi39 & n3394;
  assign n3396 = n3393 & n3395;
  assign n3397 = n3321 & n3396;
  assign n3398 = n3391 & n3397;
  assign n3399 = pi100 & ~n3349;
  assign n3400 = ~n3398 & n3399;
  assign n3401 = ~pi87 & ~n3400;
  assign n3402 = ~n3380 & n3401;
  assign n3403 = ~n3352 & ~n3402;
  assign n3404 = ~pi75 & ~n3403;
  assign n3405 = pi75 & n3349;
  assign n3406 = ~pi92 & ~n3405;
  assign n3407 = ~n3404 & n3406;
  assign n3408 = n3231 & n3344;
  assign n3409 = n3231 & n3277;
  assign n3410 = n3349 & ~n3409;
  assign n3411 = pi92 & ~n3410;
  assign n3412 = ~n3408 & n3411;
  assign n3413 = n3266 & ~n3412;
  assign n3414 = ~n3407 & n3413;
  assign n3415 = ~n3266 & n3349;
  assign n3416 = ~pi55 & ~n3415;
  assign n3417 = ~n3414 & n3416;
  assign n3418 = n3324 & ~n3345;
  assign n3419 = n3269 & n3418;
  assign n3420 = pi55 & ~n3347;
  assign n3421 = ~n3419 & n3420;
  assign n3422 = ~pi56 & ~n3421;
  assign n3423 = ~n3417 & n3422;
  assign n3424 = ~pi55 & n3269;
  assign n3425 = ~n3347 & n3424;
  assign n3426 = ~n3418 & n3425;
  assign n3427 = ~n3281 & ~n3347;
  assign n3428 = pi56 & ~n3427;
  assign n3429 = ~n3426 & n3428;
  assign n3430 = ~pi62 & ~n3429;
  assign n3431 = ~n3423 & n3430;
  assign n3432 = ~pi57 & ~pi59;
  assign n3433 = ~pi56 & n3280;
  assign n3434 = n3277 & n3433;
  assign n3435 = ~n3347 & ~n3434;
  assign n3436 = ~n3426 & ~n3435;
  assign n3437 = pi62 & ~n3436;
  assign n3438 = n3432 & ~n3437;
  assign n3439 = ~n3431 & n3438;
  assign n3440 = n3347 & ~n3432;
  assign n3441 = ~pi239 & ~n3440;
  assign n3442 = ~n3439 & n3441;
  assign n3443 = n2717 & n3094;
  assign n3444 = ~n2449 & ~n3443;
  assign n3445 = ~pi224 & n3444;
  assign n3446 = ~n3053 & ~n3306;
  assign n3447 = ~n3445 & ~n3446;
  assign n3448 = n3311 & ~n3447;
  assign n3449 = ~n3313 & ~n3448;
  assign n3450 = ~pi299 & ~n3449;
  assign n3451 = ~pi72 & ~n3358;
  assign n3452 = ~n2555 & ~n3451;
  assign n3453 = n2725 & ~n3452;
  assign n3454 = n3364 & ~n3453;
  assign n3455 = ~pi95 & ~n3454;
  assign n3456 = n2788 & ~n3455;
  assign n3457 = ~pi228 & n3456;
  assign n3458 = n3127 & n3444;
  assign n3459 = ~n3457 & ~n3458;
  assign n3460 = ~pi154 & ~n3459;
  assign n3461 = ~pi216 & ~pi221;
  assign n3462 = ~pi215 & n3461;
  assign n3463 = pi105 & ~n3444;
  assign n3464 = pi228 & ~n3463;
  assign n3465 = ~n2727 & ~n3444;
  assign n3466 = ~pi228 & ~n3465;
  assign n3467 = ~n3464 & ~n3466;
  assign n3468 = pi154 & ~n3467;
  assign n3469 = n3462 & ~n3468;
  assign n3470 = ~n3460 & n3469;
  assign n3471 = pi299 & n3339;
  assign n3472 = ~n3470 & n3471;
  assign n3473 = ~n3450 & ~n3472;
  assign n3474 = ~pi39 & ~n3473;
  assign n3475 = n2449 & n3127;
  assign n3476 = n3462 & n3475;
  assign n3477 = n3339 & ~n3476;
  assign n3478 = ~pi215 & ~n3477;
  assign n3479 = pi154 & ~n3477;
  assign n3480 = ~n3346 & ~n3478;
  assign n3481 = ~n3479 & n3480;
  assign n3482 = pi299 & ~n3481;
  assign n3483 = ~pi223 & ~pi299;
  assign n3484 = n3053 & n3483;
  assign n3485 = n2449 & n3484;
  assign n3486 = ~n3315 & ~n3485;
  assign n3487 = ~n3482 & n3486;
  assign n3488 = n3324 & ~n3479;
  assign n3489 = ~n3481 & ~n3488;
  assign n3490 = pi299 & ~n3489;
  assign n3491 = ~n3487 & ~n3490;
  assign n3492 = pi39 & ~n3491;
  assign n3493 = n3207 & ~n3492;
  assign n3494 = ~n3474 & n3493;
  assign n3495 = pi100 & n3398;
  assign n3496 = ~n3207 & ~n3487;
  assign n3497 = ~n3495 & n3496;
  assign n3498 = ~n3494 & ~n3497;
  assign n3499 = ~pi87 & ~n3498;
  assign n3500 = n3208 & n3490;
  assign n3501 = pi87 & ~n3487;
  assign n3502 = ~n3500 & n3501;
  assign n3503 = ~pi75 & ~n3502;
  assign n3504 = ~n3499 & n3503;
  assign n3505 = pi75 & n3487;
  assign n3506 = ~pi92 & ~n3505;
  assign n3507 = ~n3504 & n3506;
  assign n3508 = n3409 & n3490;
  assign n3509 = pi92 & ~n3487;
  assign n3510 = ~n3508 & n3509;
  assign n3511 = n3266 & ~n3510;
  assign n3512 = ~n3507 & n3511;
  assign n3513 = ~n3266 & n3487;
  assign n3514 = ~pi55 & ~n3513;
  assign n3515 = ~n3512 & n3514;
  assign n3516 = n3269 & n3488;
  assign n3517 = pi55 & ~n3481;
  assign n3518 = ~n3516 & n3517;
  assign n3519 = ~pi56 & ~n3518;
  assign n3520 = ~n3515 & n3519;
  assign n3521 = n3424 & n3489;
  assign n3522 = ~n3281 & ~n3481;
  assign n3523 = pi56 & ~n3522;
  assign n3524 = ~n3521 & n3523;
  assign n3525 = ~pi62 & ~n3524;
  assign n3526 = ~n3520 & n3525;
  assign n3527 = ~n3434 & ~n3481;
  assign n3528 = ~pi56 & n3521;
  assign n3529 = ~n3527 & ~n3528;
  assign n3530 = pi62 & ~n3529;
  assign n3531 = n3432 & ~n3530;
  assign n3532 = ~n3526 & n3531;
  assign n3533 = ~n3432 & n3481;
  assign n3534 = pi239 & ~n3533;
  assign n3535 = ~n3532 & n3534;
  assign po154 = n3442 | n3535;
  assign n3537 = ~pi1145 & ~n2437;
  assign n3538 = ~pi927 & n2437;
  assign n3539 = pi221 & ~n3537;
  assign n3540 = ~n3538 & n3539;
  assign n3541 = pi216 & pi274;
  assign n3542 = ~pi221 & ~n3541;
  assign n3543 = ~pi151 & n3459;
  assign n3544 = pi151 & n3467;
  assign n3545 = ~pi216 & ~n3544;
  assign n3546 = ~n3543 & n3545;
  assign n3547 = n3542 & ~n3546;
  assign n3548 = ~n3540 & ~n3547;
  assign n3549 = ~pi215 & ~n3548;
  assign n3550 = pi215 & pi1145;
  assign n3551 = pi299 & ~n3550;
  assign n3552 = ~n3549 & n3551;
  assign n3553 = ~pi1145 & ~n3041;
  assign n3554 = ~pi927 & n3041;
  assign n3555 = pi222 & ~n3553;
  assign n3556 = ~n3554 & n3555;
  assign n3557 = pi224 & pi274;
  assign n3558 = ~pi222 & ~n3557;
  assign n3559 = ~n3445 & n3558;
  assign n3560 = ~n3556 & ~n3559;
  assign n3561 = ~pi223 & ~n3560;
  assign n3562 = pi223 & pi1145;
  assign n3563 = ~pi299 & ~n3562;
  assign n3564 = ~n3561 & n3563;
  assign n3565 = ~pi39 & ~n3564;
  assign n3566 = ~n3552 & n3565;
  assign n3567 = n3305 & ~n3557;
  assign n3568 = ~n3556 & ~n3567;
  assign n3569 = ~pi223 & ~n3568;
  assign n3570 = ~n3562 & ~n3569;
  assign n3571 = ~pi299 & ~n3570;
  assign n3572 = ~n3485 & ~n3571;
  assign n3573 = ~pi151 & ~n3127;
  assign n3574 = ~n3475 & ~n3573;
  assign n3575 = ~pi151 & n3322;
  assign n3576 = ~n3574 & ~n3575;
  assign n3577 = ~pi216 & ~n3576;
  assign n3578 = n3542 & ~n3577;
  assign n3579 = ~n3540 & ~n3578;
  assign n3580 = ~pi215 & ~n3579;
  assign n3581 = ~n3550 & ~n3580;
  assign n3582 = pi299 & ~n3581;
  assign n3583 = n3572 & ~n3582;
  assign n3584 = pi39 & ~n3583;
  assign n3585 = ~pi38 & ~n3584;
  assign n3586 = ~n3566 & n3585;
  assign n3587 = ~pi216 & ~n3573;
  assign n3588 = n3542 & ~n3587;
  assign n3589 = ~n3540 & ~n3588;
  assign n3590 = ~pi215 & ~n3589;
  assign n3591 = ~n3550 & ~n3590;
  assign n3592 = n3137 & n3475;
  assign n3593 = ~n3541 & n3592;
  assign n3594 = n3591 & ~n3593;
  assign n3595 = pi299 & ~n3594;
  assign n3596 = n3572 & ~n3595;
  assign n3597 = pi38 & n3596;
  assign n3598 = ~pi100 & ~n3597;
  assign n3599 = ~n3586 & n3598;
  assign n3600 = ~pi228 & n3391;
  assign n3601 = ~n2449 & n3127;
  assign n3602 = ~n3600 & ~n3601;
  assign n3603 = ~pi151 & n3602;
  assign n3604 = n3577 & ~n3603;
  assign n3605 = n3542 & ~n3604;
  assign n3606 = ~n3540 & ~n3605;
  assign n3607 = ~pi215 & ~n3606;
  assign n3608 = ~n3550 & ~n3607;
  assign n3609 = pi299 & ~n3608;
  assign n3610 = n3182 & n3572;
  assign n3611 = ~n3609 & n3610;
  assign n3612 = ~n3182 & n3596;
  assign n3613 = pi100 & ~n3612;
  assign n3614 = ~n3611 & n3613;
  assign n3615 = ~n3599 & ~n3614;
  assign n3616 = ~pi87 & ~n3615;
  assign n3617 = ~n3208 & n3596;
  assign n3618 = n3208 & n3583;
  assign n3619 = ~n3617 & ~n3618;
  assign n3620 = pi87 & n3619;
  assign n3621 = ~pi75 & ~n3620;
  assign n3622 = ~n3616 & n3621;
  assign n3623 = pi75 & n3596;
  assign n3624 = ~pi92 & ~n3623;
  assign n3625 = ~n3622 & n3624;
  assign n3626 = n3231 & ~n3619;
  assign n3627 = ~n3231 & n3596;
  assign n3628 = pi92 & ~n3627;
  assign n3629 = ~n3626 & n3628;
  assign n3630 = n3266 & ~n3629;
  assign n3631 = ~n3625 & n3630;
  assign n3632 = ~n3266 & n3596;
  assign n3633 = ~pi55 & ~n3632;
  assign n3634 = ~n3631 & n3633;
  assign n3635 = n3269 & n3581;
  assign n3636 = ~n3269 & n3594;
  assign n3637 = pi55 & ~n3636;
  assign n3638 = ~n3635 & n3637;
  assign n3639 = ~pi56 & ~n3638;
  assign n3640 = ~n3634 & n3639;
  assign n3641 = n3281 & ~n3581;
  assign n3642 = ~n3281 & ~n3594;
  assign n3643 = pi56 & ~n3642;
  assign n3644 = ~n3641 & n3643;
  assign n3645 = ~pi62 & ~n3644;
  assign n3646 = ~n3640 & n3645;
  assign n3647 = n3434 & n3581;
  assign n3648 = ~n3434 & n3594;
  assign n3649 = pi62 & ~n3648;
  assign n3650 = ~n3647 & n3649;
  assign n3651 = pi235 & n3432;
  assign n3652 = ~n3650 & n3651;
  assign n3653 = ~n3646 & n3652;
  assign n3654 = ~n3540 & ~n3550;
  assign n3655 = n3323 & n3654;
  assign n3656 = pi299 & ~n3591;
  assign n3657 = ~n3655 & n3656;
  assign n3658 = n3277 & ~n3571;
  assign n3659 = ~n3657 & n3658;
  assign n3660 = ~n3571 & ~n3656;
  assign n3661 = ~n3208 & n3660;
  assign n3662 = ~n3659 & ~n3661;
  assign n3663 = pi87 & ~n3662;
  assign n3664 = ~pi100 & n3369;
  assign n3665 = ~pi39 & pi100;
  assign n3666 = n3391 & n3665;
  assign n3667 = ~n3664 & ~n3666;
  assign n3668 = n3393 & n3654;
  assign n3669 = ~n3667 & n3668;
  assign n3670 = n3656 & ~n3669;
  assign n3671 = ~pi87 & ~n3571;
  assign n3672 = ~n3670 & n3671;
  assign n3673 = ~n3663 & ~n3672;
  assign n3674 = ~pi75 & ~n3673;
  assign n3675 = pi75 & n3660;
  assign n3676 = ~pi92 & ~n3675;
  assign n3677 = ~n3674 & n3676;
  assign n3678 = n3231 & n3659;
  assign n3679 = ~n3409 & n3660;
  assign n3680 = pi92 & ~n3679;
  assign n3681 = ~n3678 & n3680;
  assign n3682 = n3266 & ~n3681;
  assign n3683 = ~n3677 & n3682;
  assign n3684 = ~n3266 & n3660;
  assign n3685 = ~pi55 & ~n3684;
  assign n3686 = ~n3683 & n3685;
  assign n3687 = n3269 & n3655;
  assign n3688 = pi55 & ~n3591;
  assign n3689 = ~n3687 & n3688;
  assign n3690 = ~pi56 & ~n3689;
  assign n3691 = ~n3686 & n3690;
  assign n3692 = n3281 & n3655;
  assign n3693 = ~n3591 & ~n3692;
  assign n3694 = pi56 & ~n3693;
  assign n3695 = ~pi62 & ~n3694;
  assign n3696 = ~n3691 & n3695;
  assign n3697 = ~pi56 & n3692;
  assign n3698 = pi62 & ~n3591;
  assign n3699 = ~n3697 & n3698;
  assign n3700 = ~pi235 & n3432;
  assign n3701 = ~n3699 & n3700;
  assign n3702 = ~n3696 & n3701;
  assign n3703 = pi235 & n3593;
  assign n3704 = ~n3432 & ~n3703;
  assign n3705 = n3591 & n3704;
  assign n3706 = ~n3702 & ~n3705;
  assign po155 = ~n3653 & n3706;
  assign n3708 = pi215 & pi1143;
  assign n3709 = pi299 & ~n3708;
  assign n3710 = ~pi1143 & ~n2437;
  assign n3711 = ~pi944 & n2437;
  assign n3712 = pi221 & ~n3710;
  assign n3713 = ~n3711 & n3712;
  assign n3714 = pi216 & pi264;
  assign n3715 = ~pi221 & ~n3714;
  assign n3716 = ~pi146 & ~n3456;
  assign n3717 = pi146 & n3465;
  assign n3718 = ~pi284 & ~n3717;
  assign n3719 = pi146 & pi284;
  assign n3720 = ~n3367 & n3719;
  assign n3721 = ~n3718 & ~n3720;
  assign n3722 = ~n3716 & ~n3721;
  assign n3723 = ~pi228 & ~n3722;
  assign n3724 = pi284 & ~n2449;
  assign n3725 = pi105 & ~n3724;
  assign n3726 = ~pi105 & pi146;
  assign n3727 = pi228 & ~n3726;
  assign n3728 = ~n3725 & n3727;
  assign n3729 = n3127 & ~n3444;
  assign n3730 = ~n3728 & ~n3729;
  assign n3731 = ~n3723 & n3730;
  assign n3732 = ~pi216 & ~n3731;
  assign n3733 = n3715 & ~n3732;
  assign n3734 = ~n3713 & ~n3733;
  assign n3735 = ~pi215 & ~n3734;
  assign n3736 = n3709 & ~n3735;
  assign n3737 = pi223 & pi1143;
  assign n3738 = ~pi299 & ~n3737;
  assign n3739 = ~pi1143 & ~n3041;
  assign n3740 = ~pi944 & n3041;
  assign n3741 = pi222 & ~n3739;
  assign n3742 = ~n3740 & n3741;
  assign n3743 = pi224 & pi264;
  assign n3744 = ~pi222 & ~n3743;
  assign n3745 = ~pi284 & n3444;
  assign n3746 = ~pi224 & ~n3745;
  assign n3747 = n3744 & ~n3746;
  assign n3748 = ~n3742 & ~n3747;
  assign n3749 = ~n3444 & n3744;
  assign n3750 = n3748 & ~n3749;
  assign n3751 = ~pi223 & ~n3750;
  assign n3752 = n3738 & ~n3751;
  assign n3753 = ~pi39 & ~n3752;
  assign n3754 = n3738 & n3748;
  assign n3755 = n3753 & ~n3754;
  assign n3756 = ~n3736 & n3755;
  assign n3757 = ~pi224 & n3724;
  assign n3758 = n3744 & ~n3757;
  assign n3759 = ~n3742 & ~n3758;
  assign n3760 = ~pi223 & ~n3759;
  assign n3761 = ~n3737 & ~n3760;
  assign n3762 = ~pi299 & ~n3761;
  assign n3763 = n2449 & n3101;
  assign n3764 = n3762 & ~n3763;
  assign n3765 = pi284 & n3096;
  assign n3766 = ~n3381 & ~n3765;
  assign n3767 = ~pi228 & ~n3766;
  assign n3768 = ~n3475 & ~n3728;
  assign n3769 = ~n3767 & n3768;
  assign n3770 = ~pi216 & ~n3769;
  assign n3771 = n3715 & ~n3770;
  assign n3772 = ~n3713 & ~n3771;
  assign n3773 = ~pi215 & ~n3772;
  assign n3774 = ~n3708 & ~n3773;
  assign n3775 = pi299 & ~n3774;
  assign n3776 = ~n3764 & ~n3775;
  assign n3777 = pi39 & ~n3776;
  assign n3778 = ~pi38 & ~n3777;
  assign n3779 = ~n3756 & n3778;
  assign n3780 = ~pi146 & ~pi228;
  assign n3781 = n3768 & ~n3780;
  assign n3782 = ~pi216 & ~n3781;
  assign n3783 = n3715 & ~n3782;
  assign n3784 = ~n3713 & ~n3783;
  assign n3785 = ~pi215 & ~n3784;
  assign n3786 = ~n3708 & ~n3785;
  assign n3787 = pi299 & ~n3786;
  assign n3788 = ~n3764 & ~n3787;
  assign n3789 = pi38 & n3788;
  assign n3790 = ~pi100 & ~n3789;
  assign n3791 = ~n3779 & n3790;
  assign n3792 = pi252 & n2448;
  assign n3793 = ~pi284 & ~n3792;
  assign n3794 = n3096 & n3793;
  assign n3795 = ~pi228 & ~n3794;
  assign n3796 = ~n3383 & n3795;
  assign n3797 = n3768 & ~n3796;
  assign n3798 = ~pi216 & ~n3797;
  assign n3799 = n3715 & ~n3798;
  assign n3800 = ~n3713 & ~n3799;
  assign n3801 = ~pi215 & ~n3800;
  assign n3802 = ~n3708 & ~n3801;
  assign n3803 = pi299 & ~n3802;
  assign n3804 = n3182 & ~n3764;
  assign n3805 = ~n3803 & n3804;
  assign n3806 = ~n3182 & n3788;
  assign n3807 = pi100 & ~n3806;
  assign n3808 = ~n3805 & n3807;
  assign n3809 = ~n3791 & ~n3808;
  assign n3810 = ~pi87 & ~n3809;
  assign n3811 = ~n3208 & n3788;
  assign n3812 = n3208 & n3776;
  assign n3813 = ~n3811 & ~n3812;
  assign n3814 = pi87 & n3813;
  assign n3815 = ~pi75 & ~n3814;
  assign n3816 = ~n3810 & n3815;
  assign n3817 = pi75 & n3788;
  assign n3818 = ~pi92 & ~n3817;
  assign n3819 = ~n3816 & n3818;
  assign n3820 = n3231 & ~n3813;
  assign n3821 = ~n3231 & n3788;
  assign n3822 = pi92 & ~n3821;
  assign n3823 = ~n3820 & n3822;
  assign n3824 = n3266 & ~n3823;
  assign n3825 = ~n3819 & n3824;
  assign n3826 = ~n3266 & n3788;
  assign n3827 = ~pi55 & ~n3826;
  assign n3828 = ~n3825 & n3827;
  assign n3829 = n3269 & n3774;
  assign n3830 = ~n3269 & n3786;
  assign n3831 = pi55 & ~n3830;
  assign n3832 = ~n3829 & n3831;
  assign n3833 = ~pi56 & ~n3832;
  assign n3834 = ~n3828 & n3833;
  assign n3835 = n3281 & ~n3774;
  assign n3836 = ~n3281 & ~n3786;
  assign n3837 = pi56 & ~n3836;
  assign n3838 = ~n3835 & n3837;
  assign n3839 = ~pi62 & ~n3838;
  assign n3840 = ~n3834 & n3839;
  assign n3841 = n3434 & n3774;
  assign n3842 = ~n3434 & n3786;
  assign n3843 = pi62 & ~n3842;
  assign n3844 = ~n3841 & n3843;
  assign n3845 = ~pi238 & n3432;
  assign n3846 = ~n3844 & n3845;
  assign n3847 = ~n3840 & n3846;
  assign n3848 = ~n3463 & n3728;
  assign n3849 = pi146 & ~n3456;
  assign n3850 = ~pi146 & n3465;
  assign n3851 = pi284 & ~n3850;
  assign n3852 = ~n3849 & n3851;
  assign n3853 = ~pi146 & ~pi284;
  assign n3854 = ~n3367 & n3853;
  assign n3855 = ~n3852 & ~n3854;
  assign n3856 = ~pi228 & ~n3855;
  assign n3857 = ~n3848 & ~n3856;
  assign n3858 = ~pi216 & ~n3857;
  assign n3859 = n3715 & ~n3858;
  assign n3860 = ~n3713 & ~n3859;
  assign n3861 = ~pi215 & ~n3860;
  assign n3862 = n3709 & ~n3861;
  assign n3863 = n3753 & ~n3862;
  assign n3864 = ~n3728 & ~n3767;
  assign n3865 = ~pi216 & ~n3864;
  assign n3866 = n3715 & ~n3865;
  assign n3867 = ~n3713 & ~n3866;
  assign n3868 = ~pi215 & ~n3867;
  assign n3869 = ~n3708 & ~n3868;
  assign n3870 = pi299 & ~n3869;
  assign n3871 = ~n3762 & ~n3870;
  assign n3872 = pi39 & ~n3871;
  assign n3873 = ~pi38 & ~n3872;
  assign n3874 = ~n3863 & n3873;
  assign n3875 = n3592 & ~n3714;
  assign n3876 = n3786 & ~n3875;
  assign n3877 = pi299 & ~n3876;
  assign n3878 = ~n3762 & ~n3877;
  assign n3879 = pi38 & n3878;
  assign n3880 = ~pi100 & ~n3879;
  assign n3881 = ~n3874 & n3880;
  assign n3882 = ~n3728 & ~n3796;
  assign n3883 = ~pi216 & ~n3882;
  assign n3884 = n3715 & ~n3883;
  assign n3885 = ~n3713 & ~n3884;
  assign n3886 = ~pi215 & ~n3885;
  assign n3887 = ~n3708 & ~n3886;
  assign n3888 = pi299 & ~n3887;
  assign n3889 = n3182 & ~n3762;
  assign n3890 = ~n3888 & n3889;
  assign n3891 = ~n3182 & n3878;
  assign n3892 = pi100 & ~n3891;
  assign n3893 = ~n3890 & n3892;
  assign n3894 = ~n3881 & ~n3893;
  assign n3895 = ~pi87 & ~n3894;
  assign n3896 = ~n3208 & n3878;
  assign n3897 = n3208 & n3871;
  assign n3898 = ~n3896 & ~n3897;
  assign n3899 = pi87 & n3898;
  assign n3900 = ~pi75 & ~n3899;
  assign n3901 = ~n3895 & n3900;
  assign n3902 = pi75 & n3878;
  assign n3903 = ~pi92 & ~n3902;
  assign n3904 = ~n3901 & n3903;
  assign n3905 = n3231 & ~n3898;
  assign n3906 = ~n3231 & n3878;
  assign n3907 = pi92 & ~n3906;
  assign n3908 = ~n3905 & n3907;
  assign n3909 = n3266 & ~n3908;
  assign n3910 = ~n3904 & n3909;
  assign n3911 = ~n3266 & n3878;
  assign n3912 = ~pi55 & ~n3911;
  assign n3913 = ~n3910 & n3912;
  assign n3914 = n3269 & n3869;
  assign n3915 = ~n3269 & n3876;
  assign n3916 = pi55 & ~n3915;
  assign n3917 = ~n3914 & n3916;
  assign n3918 = ~pi56 & ~n3917;
  assign n3919 = ~n3913 & n3918;
  assign n3920 = n3281 & ~n3869;
  assign n3921 = ~n3281 & ~n3876;
  assign n3922 = pi56 & ~n3921;
  assign n3923 = ~n3920 & n3922;
  assign n3924 = ~pi62 & ~n3923;
  assign n3925 = ~n3919 & n3924;
  assign n3926 = n3434 & n3869;
  assign n3927 = ~n3434 & n3876;
  assign n3928 = pi62 & ~n3927;
  assign n3929 = ~n3926 & n3928;
  assign n3930 = pi238 & n3432;
  assign n3931 = ~n3929 & n3930;
  assign n3932 = ~n3925 & n3931;
  assign n3933 = pi238 & n3875;
  assign n3934 = ~n3432 & ~n3933;
  assign n3935 = n3786 & n3934;
  assign n3936 = ~n3847 & ~n3935;
  assign po156 = ~n3932 & n3936;
  assign n3938 = pi215 & pi1142;
  assign n3939 = pi299 & ~n3938;
  assign n3940 = ~pi1142 & ~n2437;
  assign n3941 = ~pi932 & n2437;
  assign n3942 = pi221 & ~n3940;
  assign n3943 = ~n3941 & n3942;
  assign n3944 = pi216 & pi277;
  assign n3945 = ~pi221 & ~n3944;
  assign n3946 = ~pi262 & n3465;
  assign n3947 = ~pi172 & ~n3946;
  assign n3948 = pi172 & ~pi262;
  assign n3949 = n3456 & n3948;
  assign n3950 = ~n3947 & ~n3949;
  assign n3951 = pi262 & n3367;
  assign n3952 = ~pi228 & ~n3951;
  assign n3953 = ~n3950 & n3952;
  assign n3954 = pi262 & ~n2449;
  assign n3955 = pi105 & n3954;
  assign n3956 = ~n3443 & n3955;
  assign n3957 = ~pi105 & pi172;
  assign n3958 = pi228 & ~n3957;
  assign n3959 = ~n3956 & n3958;
  assign n3960 = ~n3463 & n3959;
  assign n3961 = ~pi216 & ~n3960;
  assign n3962 = ~n3953 & n3961;
  assign n3963 = n3945 & ~n3962;
  assign n3964 = ~n3943 & ~n3963;
  assign n3965 = ~pi215 & ~n3964;
  assign n3966 = n3939 & ~n3965;
  assign n3967 = pi223 & pi1142;
  assign n3968 = ~pi299 & ~n3967;
  assign n3969 = ~pi1142 & ~n3041;
  assign n3970 = ~pi932 & n3041;
  assign n3971 = pi222 & ~n3969;
  assign n3972 = ~n3970 & n3971;
  assign n3973 = pi224 & pi277;
  assign n3974 = ~pi222 & ~n3973;
  assign n3975 = ~pi262 & n3444;
  assign n3976 = ~pi224 & ~n3975;
  assign n3977 = n3974 & ~n3976;
  assign n3978 = ~n3972 & ~n3977;
  assign n3979 = n3968 & n3978;
  assign n3980 = ~n3444 & n3974;
  assign n3981 = n3978 & ~n3980;
  assign n3982 = ~pi223 & ~n3981;
  assign n3983 = n3968 & ~n3982;
  assign n3984 = ~pi39 & ~n3983;
  assign n3985 = ~n3979 & n3984;
  assign n3986 = ~n3966 & n3985;
  assign n3987 = ~pi224 & n3954;
  assign n3988 = n3974 & ~n3987;
  assign n3989 = ~n3972 & ~n3988;
  assign n3990 = ~pi223 & ~n3989;
  assign n3991 = ~n3967 & ~n3990;
  assign n3992 = ~pi299 & ~n3991;
  assign n3993 = ~n3763 & n3992;
  assign n3994 = ~pi262 & n3096;
  assign n3995 = pi172 & ~pi228;
  assign n3996 = ~n3322 & ~n3995;
  assign n3997 = ~n3994 & ~n3996;
  assign n3998 = ~n3955 & ~n3957;
  assign n3999 = pi228 & ~n3998;
  assign n4000 = ~n3475 & ~n3999;
  assign n4001 = ~n3997 & n4000;
  assign n4002 = ~pi216 & ~n4001;
  assign n4003 = n3945 & ~n4002;
  assign n4004 = ~n3943 & ~n4003;
  assign n4005 = ~pi215 & ~n4004;
  assign n4006 = ~n3938 & ~n4005;
  assign n4007 = pi299 & ~n4006;
  assign n4008 = ~n3993 & ~n4007;
  assign n4009 = pi39 & ~n4008;
  assign n4010 = ~pi38 & ~n4009;
  assign n4011 = ~n3986 & n4010;
  assign n4012 = ~n3995 & ~n3999;
  assign n4013 = ~pi216 & ~n4012;
  assign n4014 = n3945 & ~n4013;
  assign n4015 = ~n3943 & ~n4014;
  assign n4016 = ~pi215 & ~n4015;
  assign n4017 = ~n3938 & ~n4016;
  assign n4018 = ~n3476 & ~n4017;
  assign n4019 = pi299 & n4018;
  assign n4020 = ~n3993 & ~n4019;
  assign n4021 = pi38 & n4020;
  assign n4022 = ~pi100 & ~n4021;
  assign n4023 = ~n4011 & n4022;
  assign n4024 = ~pi262 & n3391;
  assign n4025 = ~n3600 & ~n3995;
  assign n4026 = ~n4024 & ~n4025;
  assign n4027 = n4000 & ~n4026;
  assign n4028 = ~pi216 & ~n4027;
  assign n4029 = n3945 & ~n4028;
  assign n4030 = ~n3943 & ~n4029;
  assign n4031 = ~pi215 & ~n4030;
  assign n4032 = ~n3938 & ~n4031;
  assign n4033 = pi299 & ~n4032;
  assign n4034 = n3182 & ~n3993;
  assign n4035 = ~n4033 & n4034;
  assign n4036 = ~n3182 & n4020;
  assign n4037 = pi100 & ~n4036;
  assign n4038 = ~n4035 & n4037;
  assign n4039 = ~n4023 & ~n4038;
  assign n4040 = ~pi87 & ~n4039;
  assign n4041 = ~n3208 & n4020;
  assign n4042 = n3208 & n4008;
  assign n4043 = ~n4041 & ~n4042;
  assign n4044 = pi87 & n4043;
  assign n4045 = ~pi75 & ~n4044;
  assign n4046 = ~n4040 & n4045;
  assign n4047 = pi75 & n4020;
  assign n4048 = ~pi92 & ~n4047;
  assign n4049 = ~n4046 & n4048;
  assign n4050 = n3231 & ~n4043;
  assign n4051 = ~n3231 & n4020;
  assign n4052 = pi92 & ~n4051;
  assign n4053 = ~n4050 & n4052;
  assign n4054 = n3266 & ~n4053;
  assign n4055 = ~n4049 & n4054;
  assign n4056 = ~n3266 & n4020;
  assign n4057 = ~pi55 & ~n4056;
  assign n4058 = ~n4055 & n4057;
  assign n4059 = n3269 & n4006;
  assign n4060 = ~n3269 & ~n4018;
  assign n4061 = pi55 & ~n4060;
  assign n4062 = ~n4059 & n4061;
  assign n4063 = ~pi56 & ~n4062;
  assign n4064 = ~n4058 & n4063;
  assign n4065 = n3281 & ~n4006;
  assign n4066 = ~n3281 & n4018;
  assign n4067 = pi56 & ~n4066;
  assign n4068 = ~n4065 & n4067;
  assign n4069 = ~pi62 & ~n4068;
  assign n4070 = ~n4064 & n4069;
  assign n4071 = n3434 & n4006;
  assign n4072 = ~n3434 & ~n4018;
  assign n4073 = pi62 & ~n4072;
  assign n4074 = ~n4071 & n4073;
  assign n4075 = n3432 & ~n4074;
  assign n4076 = ~n4070 & n4075;
  assign n4077 = ~n3432 & ~n4018;
  assign n4078 = ~pi249 & ~n4077;
  assign n4079 = ~n4076 & n4078;
  assign n4080 = pi262 & n3456;
  assign n4081 = ~pi172 & ~n4080;
  assign n4082 = ~pi262 & ~n3367;
  assign n4083 = pi262 & ~n3465;
  assign n4084 = pi172 & ~n4083;
  assign n4085 = ~n4082 & n4084;
  assign n4086 = ~n4081 & ~n4085;
  assign n4087 = ~pi228 & ~n4086;
  assign n4088 = ~pi216 & ~n3959;
  assign n4089 = ~n4087 & n4088;
  assign n4090 = n3945 & ~n4089;
  assign n4091 = ~n3943 & ~n4090;
  assign n4092 = ~pi215 & ~n4091;
  assign n4093 = n3939 & ~n4092;
  assign n4094 = n3984 & ~n4093;
  assign n4095 = ~n3997 & ~n3999;
  assign n4096 = ~pi216 & ~n4095;
  assign n4097 = n3945 & ~n4096;
  assign n4098 = ~n3943 & ~n4097;
  assign n4099 = ~pi215 & ~n4098;
  assign n4100 = ~n3938 & ~n4099;
  assign n4101 = pi299 & ~n4100;
  assign n4102 = ~n3992 & ~n4101;
  assign n4103 = pi39 & ~n4102;
  assign n4104 = ~pi38 & ~n4103;
  assign n4105 = ~n4094 & n4104;
  assign n4106 = pi299 & ~n4017;
  assign n4107 = ~n3992 & ~n4106;
  assign n4108 = pi38 & n4107;
  assign n4109 = ~pi100 & ~n4108;
  assign n4110 = ~n4105 & n4109;
  assign n4111 = ~n3999 & ~n4026;
  assign n4112 = ~pi216 & ~n4111;
  assign n4113 = n3945 & ~n4112;
  assign n4114 = ~n3943 & ~n4113;
  assign n4115 = ~pi215 & ~n4114;
  assign n4116 = ~n3938 & ~n4115;
  assign n4117 = pi299 & ~n4116;
  assign n4118 = n3182 & ~n3992;
  assign n4119 = ~n4117 & n4118;
  assign n4120 = ~n3182 & n4107;
  assign n4121 = pi100 & ~n4120;
  assign n4122 = ~n4119 & n4121;
  assign n4123 = ~n4110 & ~n4122;
  assign n4124 = ~pi87 & ~n4123;
  assign n4125 = ~n3208 & n4107;
  assign n4126 = n3208 & n4102;
  assign n4127 = ~n4125 & ~n4126;
  assign n4128 = pi87 & n4127;
  assign n4129 = ~pi75 & ~n4128;
  assign n4130 = ~n4124 & n4129;
  assign n4131 = pi75 & n4107;
  assign n4132 = ~pi92 & ~n4131;
  assign n4133 = ~n4130 & n4132;
  assign n4134 = n3231 & ~n4127;
  assign n4135 = ~n3231 & n4107;
  assign n4136 = pi92 & ~n4135;
  assign n4137 = ~n4134 & n4136;
  assign n4138 = n3266 & ~n4137;
  assign n4139 = ~n4133 & n4138;
  assign n4140 = ~n3266 & n4107;
  assign n4141 = ~pi55 & ~n4140;
  assign n4142 = ~n4139 & n4141;
  assign n4143 = n3269 & n4100;
  assign n4144 = ~n3269 & n4017;
  assign n4145 = pi55 & ~n4144;
  assign n4146 = ~n4143 & n4145;
  assign n4147 = ~pi56 & ~n4146;
  assign n4148 = ~n4142 & n4147;
  assign n4149 = n3281 & ~n4100;
  assign n4150 = ~n3281 & ~n4017;
  assign n4151 = pi56 & ~n4150;
  assign n4152 = ~n4149 & n4151;
  assign n4153 = ~pi62 & ~n4152;
  assign n4154 = ~n4148 & n4153;
  assign n4155 = n3434 & n4100;
  assign n4156 = ~n3434 & n4017;
  assign n4157 = pi62 & ~n4156;
  assign n4158 = ~n4155 & n4157;
  assign n4159 = n3432 & ~n4158;
  assign n4160 = ~n4154 & n4159;
  assign n4161 = ~n3432 & n4017;
  assign n4162 = pi249 & ~n4161;
  assign n4163 = ~n4160 & n4162;
  assign po157 = n4079 | n4163;
  assign n4165 = pi215 & pi1141;
  assign n4166 = pi299 & ~n4165;
  assign n4167 = ~pi1141 & ~n2437;
  assign n4168 = ~pi935 & n2437;
  assign n4169 = pi221 & ~n4167;
  assign n4170 = ~n4168 & n4169;
  assign n4171 = pi216 & pi270;
  assign n4172 = ~pi221 & ~n4171;
  assign n4173 = pi861 & n3465;
  assign n4174 = ~pi171 & ~n4173;
  assign n4175 = pi171 & n3456;
  assign n4176 = ~n4174 & ~n4175;
  assign n4177 = pi861 & ~n4176;
  assign n4178 = ~n3367 & n4174;
  assign n4179 = ~n4177 & ~n4178;
  assign n4180 = ~pi228 & ~n4179;
  assign n4181 = pi861 & ~n2449;
  assign n4182 = pi105 & ~n4181;
  assign n4183 = ~pi105 & pi171;
  assign n4184 = pi228 & ~n4183;
  assign n4185 = ~n4182 & n4184;
  assign n4186 = ~n3463 & n4185;
  assign n4187 = ~pi216 & ~n4186;
  assign n4188 = ~n4180 & n4187;
  assign n4189 = n4172 & ~n4188;
  assign n4190 = ~n4170 & ~n4189;
  assign n4191 = ~pi215 & ~n4190;
  assign n4192 = n4166 & ~n4191;
  assign n4193 = pi223 & pi1141;
  assign n4194 = ~pi299 & ~n4193;
  assign n4195 = ~pi1141 & ~n3041;
  assign n4196 = ~pi935 & n3041;
  assign n4197 = pi222 & ~n4195;
  assign n4198 = ~n4196 & n4197;
  assign n4199 = pi224 & pi270;
  assign n4200 = ~pi222 & ~n4199;
  assign n4201 = pi861 & n3444;
  assign n4202 = ~pi224 & ~n4201;
  assign n4203 = n4200 & ~n4202;
  assign n4204 = ~n4198 & ~n4203;
  assign n4205 = n4194 & n4204;
  assign n4206 = ~n3444 & n4200;
  assign n4207 = n4204 & ~n4206;
  assign n4208 = ~pi223 & ~n4207;
  assign n4209 = n4194 & ~n4208;
  assign n4210 = ~pi39 & ~n4209;
  assign n4211 = ~n4205 & n4210;
  assign n4212 = ~n4192 & n4211;
  assign n4213 = ~pi224 & ~n4181;
  assign n4214 = n4200 & ~n4213;
  assign n4215 = ~n4198 & ~n4214;
  assign n4216 = ~pi223 & ~n4215;
  assign n4217 = ~n4193 & ~n4216;
  assign n4218 = ~pi299 & ~n4217;
  assign n4219 = ~pi216 & ~n4185;
  assign n4220 = ~pi861 & n3096;
  assign n4221 = pi171 & ~n3096;
  assign n4222 = ~pi228 & ~n4220;
  assign n4223 = ~n4221 & n4222;
  assign n4224 = n4219 & ~n4223;
  assign n4225 = n4172 & ~n4224;
  assign n4226 = ~n4170 & ~n4225;
  assign n4227 = ~pi215 & ~n4226;
  assign n4228 = ~n4165 & ~n4227;
  assign n4229 = pi299 & ~n4228;
  assign n4230 = ~n4218 & ~n4229;
  assign n4231 = pi39 & ~n4230;
  assign n4232 = ~pi38 & ~n4231;
  assign n4233 = ~n4212 & n4232;
  assign n4234 = ~pi171 & ~pi228;
  assign n4235 = n4219 & ~n4234;
  assign n4236 = n4172 & ~n4235;
  assign n4237 = ~n4170 & ~n4236;
  assign n4238 = ~pi215 & ~n4237;
  assign n4239 = ~n4165 & ~n4238;
  assign n4240 = pi299 & ~n4239;
  assign n4241 = ~n4218 & ~n4240;
  assign n4242 = pi38 & n4241;
  assign n4243 = ~pi100 & ~n4242;
  assign n4244 = ~n4233 & n4243;
  assign n4245 = ~pi861 & n3391;
  assign n4246 = ~n3600 & ~n4234;
  assign n4247 = ~n4245 & ~n4246;
  assign n4248 = n4219 & ~n4247;
  assign n4249 = n4172 & ~n4248;
  assign n4250 = ~n4170 & ~n4249;
  assign n4251 = ~pi215 & ~n4250;
  assign n4252 = ~n4165 & ~n4251;
  assign n4253 = pi299 & ~n4252;
  assign n4254 = n3182 & ~n4218;
  assign n4255 = ~n4253 & n4254;
  assign n4256 = ~n3182 & n4241;
  assign n4257 = pi100 & ~n4256;
  assign n4258 = ~n4255 & n4257;
  assign n4259 = ~n4244 & ~n4258;
  assign n4260 = ~pi87 & ~n4259;
  assign n4261 = ~n3208 & n4241;
  assign n4262 = n3208 & n4230;
  assign n4263 = ~n4261 & ~n4262;
  assign n4264 = pi87 & n4263;
  assign n4265 = ~pi75 & ~n4264;
  assign n4266 = ~n4260 & n4265;
  assign n4267 = pi75 & n4241;
  assign n4268 = ~pi92 & ~n4267;
  assign n4269 = ~n4266 & n4268;
  assign n4270 = n3231 & ~n4263;
  assign n4271 = ~n3231 & n4241;
  assign n4272 = pi92 & ~n4271;
  assign n4273 = ~n4270 & n4272;
  assign n4274 = n3266 & ~n4273;
  assign n4275 = ~n4269 & n4274;
  assign n4276 = ~n3266 & n4241;
  assign n4277 = ~pi55 & ~n4276;
  assign n4278 = ~n4275 & n4277;
  assign n4279 = n3269 & n4228;
  assign n4280 = ~n3269 & n4239;
  assign n4281 = pi55 & ~n4280;
  assign n4282 = ~n4279 & n4281;
  assign n4283 = ~pi56 & ~n4282;
  assign n4284 = ~n4278 & n4283;
  assign n4285 = n3281 & ~n4228;
  assign n4286 = ~n3281 & ~n4239;
  assign n4287 = pi56 & ~n4286;
  assign n4288 = ~n4285 & n4287;
  assign n4289 = ~pi62 & ~n4288;
  assign n4290 = ~n4284 & n4289;
  assign n4291 = n3434 & n4228;
  assign n4292 = ~n3434 & n4239;
  assign n4293 = pi62 & ~n4292;
  assign n4294 = ~n4291 & n4293;
  assign n4295 = ~pi241 & n3432;
  assign n4296 = ~n4294 & n4295;
  assign n4297 = ~n4290 & n4296;
  assign n4298 = ~pi861 & n3456;
  assign n4299 = ~pi171 & ~n4298;
  assign n4300 = pi861 & ~n3367;
  assign n4301 = ~pi861 & ~n3465;
  assign n4302 = pi171 & ~n4301;
  assign n4303 = ~n4300 & n4302;
  assign n4304 = ~n4299 & ~n4303;
  assign n4305 = ~pi228 & ~n4304;
  assign n4306 = ~n3729 & n4219;
  assign n4307 = ~n4305 & n4306;
  assign n4308 = n4172 & ~n4307;
  assign n4309 = ~n4170 & ~n4308;
  assign n4310 = ~pi215 & ~n4309;
  assign n4311 = n4166 & ~n4310;
  assign n4312 = n4210 & ~n4311;
  assign n4313 = ~n3485 & ~n4218;
  assign n4314 = ~n3475 & n4219;
  assign n4315 = ~n4223 & n4314;
  assign n4316 = n4172 & ~n4315;
  assign n4317 = ~n4170 & ~n4316;
  assign n4318 = ~pi215 & ~n4317;
  assign n4319 = ~n4165 & ~n4318;
  assign n4320 = pi299 & ~n4319;
  assign n4321 = n4313 & ~n4320;
  assign n4322 = pi39 & ~n4321;
  assign n4323 = ~pi38 & ~n4322;
  assign n4324 = ~n4312 & n4323;
  assign n4325 = n3592 & ~n4171;
  assign n4326 = n4239 & ~n4325;
  assign n4327 = pi299 & ~n4326;
  assign n4328 = n4313 & ~n4327;
  assign n4329 = pi38 & n4328;
  assign n4330 = ~pi100 & ~n4329;
  assign n4331 = ~n4324 & n4330;
  assign n4332 = ~n4247 & n4314;
  assign n4333 = n4172 & ~n4332;
  assign n4334 = ~n4170 & ~n4333;
  assign n4335 = ~pi215 & ~n4334;
  assign n4336 = ~n4165 & ~n4335;
  assign n4337 = pi299 & ~n4336;
  assign n4338 = n3182 & n4313;
  assign n4339 = ~n4337 & n4338;
  assign n4340 = ~n3182 & n4328;
  assign n4341 = pi100 & ~n4340;
  assign n4342 = ~n4339 & n4341;
  assign n4343 = ~n4331 & ~n4342;
  assign n4344 = ~pi87 & ~n4343;
  assign n4345 = ~n3208 & n4328;
  assign n4346 = n3208 & n4321;
  assign n4347 = ~n4345 & ~n4346;
  assign n4348 = pi87 & n4347;
  assign n4349 = ~pi75 & ~n4348;
  assign n4350 = ~n4344 & n4349;
  assign n4351 = pi75 & n4328;
  assign n4352 = ~pi92 & ~n4351;
  assign n4353 = ~n4350 & n4352;
  assign n4354 = n3231 & ~n4347;
  assign n4355 = ~n3231 & n4328;
  assign n4356 = pi92 & ~n4355;
  assign n4357 = ~n4354 & n4356;
  assign n4358 = n3266 & ~n4357;
  assign n4359 = ~n4353 & n4358;
  assign n4360 = ~n3266 & n4328;
  assign n4361 = ~pi55 & ~n4360;
  assign n4362 = ~n4359 & n4361;
  assign n4363 = n3269 & n4319;
  assign n4364 = ~n3269 & n4326;
  assign n4365 = pi55 & ~n4364;
  assign n4366 = ~n4363 & n4365;
  assign n4367 = ~pi56 & ~n4366;
  assign n4368 = ~n4362 & n4367;
  assign n4369 = n3281 & ~n4319;
  assign n4370 = ~n3281 & ~n4326;
  assign n4371 = pi56 & ~n4370;
  assign n4372 = ~n4369 & n4371;
  assign n4373 = ~pi62 & ~n4372;
  assign n4374 = ~n4368 & n4373;
  assign n4375 = n3434 & n4319;
  assign n4376 = ~n3434 & n4326;
  assign n4377 = pi62 & ~n4376;
  assign n4378 = ~n4375 & n4377;
  assign n4379 = pi241 & n3432;
  assign n4380 = ~n4378 & n4379;
  assign n4381 = ~n4374 & n4380;
  assign n4382 = pi241 & n4325;
  assign n4383 = ~n3432 & ~n4382;
  assign n4384 = n4239 & n4383;
  assign n4385 = ~n4381 & ~n4384;
  assign po158 = ~n4297 & n4385;
  assign n4387 = pi215 & pi1140;
  assign n4388 = pi299 & ~n4387;
  assign n4389 = ~pi1140 & ~n2437;
  assign n4390 = ~pi921 & n2437;
  assign n4391 = pi221 & ~n4389;
  assign n4392 = ~n4390 & n4391;
  assign n4393 = pi216 & pi282;
  assign n4394 = ~pi221 & ~n4393;
  assign n4395 = pi869 & n3465;
  assign n4396 = ~pi170 & ~n4395;
  assign n4397 = pi170 & n3456;
  assign n4398 = ~n4396 & ~n4397;
  assign n4399 = pi869 & ~n4398;
  assign n4400 = ~n3367 & n4396;
  assign n4401 = ~n4399 & ~n4400;
  assign n4402 = ~pi228 & ~n4401;
  assign n4403 = pi869 & ~n2449;
  assign n4404 = pi105 & ~n4403;
  assign n4405 = ~pi105 & pi170;
  assign n4406 = pi228 & ~n4405;
  assign n4407 = ~n4404 & n4406;
  assign n4408 = ~n3463 & n4407;
  assign n4409 = ~pi216 & ~n4408;
  assign n4410 = ~n4402 & n4409;
  assign n4411 = n4394 & ~n4410;
  assign n4412 = ~n4392 & ~n4411;
  assign n4413 = ~pi215 & ~n4412;
  assign n4414 = n4388 & ~n4413;
  assign n4415 = pi223 & pi1140;
  assign n4416 = ~pi299 & ~n4415;
  assign n4417 = ~pi1140 & ~n3041;
  assign n4418 = ~pi921 & n3041;
  assign n4419 = pi222 & ~n4417;
  assign n4420 = ~n4418 & n4419;
  assign n4421 = pi224 & pi282;
  assign n4422 = ~pi222 & ~n4421;
  assign n4423 = pi869 & n3444;
  assign n4424 = ~pi224 & ~n4423;
  assign n4425 = n4422 & ~n4424;
  assign n4426 = ~n4420 & ~n4425;
  assign n4427 = n4416 & n4426;
  assign n4428 = ~n3444 & n4422;
  assign n4429 = n4426 & ~n4428;
  assign n4430 = ~pi223 & ~n4429;
  assign n4431 = n4416 & ~n4430;
  assign n4432 = ~pi39 & ~n4431;
  assign n4433 = ~n4427 & n4432;
  assign n4434 = ~n4414 & n4433;
  assign n4435 = ~pi224 & ~n4403;
  assign n4436 = n4422 & ~n4435;
  assign n4437 = ~n4420 & ~n4436;
  assign n4438 = ~pi223 & ~n4437;
  assign n4439 = ~n4415 & ~n4438;
  assign n4440 = ~pi299 & ~n4439;
  assign n4441 = ~pi216 & ~n4407;
  assign n4442 = ~pi869 & n3096;
  assign n4443 = pi170 & ~n3096;
  assign n4444 = ~pi228 & ~n4442;
  assign n4445 = ~n4443 & n4444;
  assign n4446 = n4441 & ~n4445;
  assign n4447 = n4394 & ~n4446;
  assign n4448 = ~n4392 & ~n4447;
  assign n4449 = ~pi215 & ~n4448;
  assign n4450 = ~n4387 & ~n4449;
  assign n4451 = pi299 & ~n4450;
  assign n4452 = ~n4440 & ~n4451;
  assign n4453 = pi39 & ~n4452;
  assign n4454 = ~pi38 & ~n4453;
  assign n4455 = ~n4434 & n4454;
  assign n4456 = ~pi170 & ~pi228;
  assign n4457 = n4441 & ~n4456;
  assign n4458 = n4394 & ~n4457;
  assign n4459 = ~n4392 & ~n4458;
  assign n4460 = ~pi215 & ~n4459;
  assign n4461 = ~n4387 & ~n4460;
  assign n4462 = pi299 & ~n4461;
  assign n4463 = ~n4440 & ~n4462;
  assign n4464 = pi38 & n4463;
  assign n4465 = ~pi100 & ~n4464;
  assign n4466 = ~n4455 & n4465;
  assign n4467 = ~pi869 & n3391;
  assign n4468 = ~n3600 & ~n4456;
  assign n4469 = ~n4467 & ~n4468;
  assign n4470 = n4441 & ~n4469;
  assign n4471 = n4394 & ~n4470;
  assign n4472 = ~n4392 & ~n4471;
  assign n4473 = ~pi215 & ~n4472;
  assign n4474 = ~n4387 & ~n4473;
  assign n4475 = pi299 & ~n4474;
  assign n4476 = n3182 & ~n4440;
  assign n4477 = ~n4475 & n4476;
  assign n4478 = ~n3182 & n4463;
  assign n4479 = pi100 & ~n4478;
  assign n4480 = ~n4477 & n4479;
  assign n4481 = ~n4466 & ~n4480;
  assign n4482 = ~pi87 & ~n4481;
  assign n4483 = ~n3208 & n4463;
  assign n4484 = n3208 & n4452;
  assign n4485 = ~n4483 & ~n4484;
  assign n4486 = pi87 & n4485;
  assign n4487 = ~pi75 & ~n4486;
  assign n4488 = ~n4482 & n4487;
  assign n4489 = pi75 & n4463;
  assign n4490 = ~pi92 & ~n4489;
  assign n4491 = ~n4488 & n4490;
  assign n4492 = n3231 & ~n4485;
  assign n4493 = ~n3231 & n4463;
  assign n4494 = pi92 & ~n4493;
  assign n4495 = ~n4492 & n4494;
  assign n4496 = n3266 & ~n4495;
  assign n4497 = ~n4491 & n4496;
  assign n4498 = ~n3266 & n4463;
  assign n4499 = ~pi55 & ~n4498;
  assign n4500 = ~n4497 & n4499;
  assign n4501 = n3269 & n4450;
  assign n4502 = ~n3269 & n4461;
  assign n4503 = pi55 & ~n4502;
  assign n4504 = ~n4501 & n4503;
  assign n4505 = ~pi56 & ~n4504;
  assign n4506 = ~n4500 & n4505;
  assign n4507 = n3281 & ~n4450;
  assign n4508 = ~n3281 & ~n4461;
  assign n4509 = pi56 & ~n4508;
  assign n4510 = ~n4507 & n4509;
  assign n4511 = ~pi62 & ~n4510;
  assign n4512 = ~n4506 & n4511;
  assign n4513 = n3434 & n4450;
  assign n4514 = ~n3434 & n4461;
  assign n4515 = pi62 & ~n4514;
  assign n4516 = ~n4513 & n4515;
  assign n4517 = ~pi248 & n3432;
  assign n4518 = ~n4516 & n4517;
  assign n4519 = ~n4512 & n4518;
  assign n4520 = ~pi869 & n3456;
  assign n4521 = ~pi170 & ~n4520;
  assign n4522 = pi869 & ~n3367;
  assign n4523 = ~pi869 & ~n3465;
  assign n4524 = pi170 & ~n4523;
  assign n4525 = ~n4522 & n4524;
  assign n4526 = ~n4521 & ~n4525;
  assign n4527 = ~pi228 & ~n4526;
  assign n4528 = ~n3729 & n4441;
  assign n4529 = ~n4527 & n4528;
  assign n4530 = n4394 & ~n4529;
  assign n4531 = ~n4392 & ~n4530;
  assign n4532 = ~pi215 & ~n4531;
  assign n4533 = n4388 & ~n4532;
  assign n4534 = n4432 & ~n4533;
  assign n4535 = ~n3485 & ~n4440;
  assign n4536 = ~n3475 & n4441;
  assign n4537 = ~n4445 & n4536;
  assign n4538 = n4394 & ~n4537;
  assign n4539 = ~n4392 & ~n4538;
  assign n4540 = ~pi215 & ~n4539;
  assign n4541 = ~n4387 & ~n4540;
  assign n4542 = pi299 & ~n4541;
  assign n4543 = n4535 & ~n4542;
  assign n4544 = pi39 & ~n4543;
  assign n4545 = ~pi38 & ~n4544;
  assign n4546 = ~n4534 & n4545;
  assign n4547 = n3592 & ~n4393;
  assign n4548 = n4461 & ~n4547;
  assign n4549 = pi299 & ~n4548;
  assign n4550 = n4535 & ~n4549;
  assign n4551 = pi38 & n4550;
  assign n4552 = ~pi100 & ~n4551;
  assign n4553 = ~n4546 & n4552;
  assign n4554 = ~n4469 & n4536;
  assign n4555 = n4394 & ~n4554;
  assign n4556 = ~n4392 & ~n4555;
  assign n4557 = ~pi215 & ~n4556;
  assign n4558 = ~n4387 & ~n4557;
  assign n4559 = pi299 & ~n4558;
  assign n4560 = n3182 & n4535;
  assign n4561 = ~n4559 & n4560;
  assign n4562 = ~n3182 & n4550;
  assign n4563 = pi100 & ~n4562;
  assign n4564 = ~n4561 & n4563;
  assign n4565 = ~n4553 & ~n4564;
  assign n4566 = ~pi87 & ~n4565;
  assign n4567 = ~n3208 & n4550;
  assign n4568 = n3208 & n4543;
  assign n4569 = ~n4567 & ~n4568;
  assign n4570 = pi87 & n4569;
  assign n4571 = ~pi75 & ~n4570;
  assign n4572 = ~n4566 & n4571;
  assign n4573 = pi75 & n4550;
  assign n4574 = ~pi92 & ~n4573;
  assign n4575 = ~n4572 & n4574;
  assign n4576 = n3231 & ~n4569;
  assign n4577 = ~n3231 & n4550;
  assign n4578 = pi92 & ~n4577;
  assign n4579 = ~n4576 & n4578;
  assign n4580 = n3266 & ~n4579;
  assign n4581 = ~n4575 & n4580;
  assign n4582 = ~n3266 & n4550;
  assign n4583 = ~pi55 & ~n4582;
  assign n4584 = ~n4581 & n4583;
  assign n4585 = n3269 & n4541;
  assign n4586 = ~n3269 & n4548;
  assign n4587 = pi55 & ~n4586;
  assign n4588 = ~n4585 & n4587;
  assign n4589 = ~pi56 & ~n4588;
  assign n4590 = ~n4584 & n4589;
  assign n4591 = n3281 & ~n4541;
  assign n4592 = ~n3281 & ~n4548;
  assign n4593 = pi56 & ~n4592;
  assign n4594 = ~n4591 & n4593;
  assign n4595 = ~pi62 & ~n4594;
  assign n4596 = ~n4590 & n4595;
  assign n4597 = n3434 & n4541;
  assign n4598 = ~n3434 & n4548;
  assign n4599 = pi62 & ~n4598;
  assign n4600 = ~n4597 & n4599;
  assign n4601 = pi248 & n3432;
  assign n4602 = ~n4600 & n4601;
  assign n4603 = ~n4596 & n4602;
  assign n4604 = pi248 & n4547;
  assign n4605 = ~n3432 & ~n4604;
  assign n4606 = n4461 & n4605;
  assign n4607 = ~n4603 & ~n4606;
  assign po159 = ~n4519 & n4607;
  assign n4609 = ~pi148 & ~pi215;
  assign n4610 = pi833 & pi920;
  assign n4611 = ~pi833 & pi1139;
  assign n4612 = ~pi216 & ~n4610;
  assign n4613 = ~n4611 & n4612;
  assign n4614 = pi216 & ~pi1139;
  assign n4615 = pi221 & ~n4614;
  assign n4616 = ~n4613 & n4615;
  assign n4617 = pi216 & pi281;
  assign n4618 = ~pi221 & ~n4617;
  assign n4619 = ~n3127 & ~n3322;
  assign n4620 = pi862 & ~n3475;
  assign n4621 = ~pi216 & ~n4620;
  assign n4622 = ~n4619 & n4621;
  assign n4623 = n4618 & ~n4622;
  assign n4624 = ~n4616 & ~n4623;
  assign n4625 = ~n3127 & ~n3600;
  assign n4626 = n4618 & n4625;
  assign n4627 = n4624 & ~n4626;
  assign n4628 = n4609 & ~n4627;
  assign n4629 = ~pi216 & ~pi862;
  assign n4630 = ~n3322 & ~n3601;
  assign n4631 = n4629 & ~n4630;
  assign n4632 = n4618 & ~n4631;
  assign n4633 = ~n4616 & ~n4632;
  assign n4634 = n3602 & n4618;
  assign n4635 = n4633 & ~n4634;
  assign n4636 = pi148 & ~pi215;
  assign n4637 = ~pi216 & ~n4616;
  assign n4638 = n3602 & n4637;
  assign n4639 = n4636 & ~n4638;
  assign n4640 = ~n4635 & n4639;
  assign n4641 = pi215 & pi1139;
  assign n4642 = ~n4628 & ~n4641;
  assign n4643 = ~n4640 & n4642;
  assign n4644 = pi299 & ~n4643;
  assign n4645 = ~pi1139 & ~n3041;
  assign n4646 = ~pi920 & n3041;
  assign n4647 = pi222 & ~n4645;
  assign n4648 = ~n4646 & n4647;
  assign n4649 = pi223 & pi1139;
  assign n4650 = ~pi224 & ~n4649;
  assign n4651 = ~n4648 & n4650;
  assign n4652 = n2449 & n4651;
  assign n4653 = ~pi862 & n4651;
  assign n4654 = pi224 & pi281;
  assign n4655 = ~pi222 & ~n4654;
  assign n4656 = ~n4648 & ~n4655;
  assign n4657 = ~pi223 & ~n4656;
  assign n4658 = ~n4649 & ~n4657;
  assign n4659 = ~pi299 & ~n4658;
  assign n4660 = ~n4653 & n4659;
  assign n4661 = ~n4652 & n4660;
  assign n4662 = n3182 & ~n4661;
  assign n4663 = ~n4644 & n4662;
  assign n4664 = n3601 & n4629;
  assign n4665 = n4618 & ~n4664;
  assign n4666 = ~n4616 & ~n4665;
  assign n4667 = pi148 & ~n3127;
  assign n4668 = n4637 & n4667;
  assign n4669 = ~pi215 & ~n4668;
  assign n4670 = ~n4666 & n4669;
  assign n4671 = ~n4641 & ~n4670;
  assign n4672 = ~n3476 & ~n4671;
  assign n4673 = pi299 & n4672;
  assign n4674 = ~n4661 & ~n4673;
  assign n4675 = ~n3182 & n4674;
  assign n4676 = pi100 & ~n4675;
  assign n4677 = ~n4663 & n4676;
  assign n4678 = ~pi228 & n3367;
  assign n4679 = ~n3127 & ~n4678;
  assign n4680 = ~pi862 & n4679;
  assign n4681 = pi862 & ~n3467;
  assign n4682 = ~pi216 & ~n4681;
  assign n4683 = ~n4680 & n4682;
  assign n4684 = n4618 & ~n4683;
  assign n4685 = ~n4616 & ~n4684;
  assign n4686 = n4609 & ~n4685;
  assign n4687 = ~n3459 & n4629;
  assign n4688 = n4618 & ~n4687;
  assign n4689 = ~n4616 & ~n4688;
  assign n4690 = n3459 & n4637;
  assign n4691 = n4636 & ~n4690;
  assign n4692 = ~n4689 & n4691;
  assign n4693 = pi299 & ~n4641;
  assign n4694 = ~n4692 & n4693;
  assign n4695 = ~n4686 & n4694;
  assign n4696 = ~n3444 & n4651;
  assign n4697 = ~n4653 & ~n4658;
  assign n4698 = ~n4696 & n4697;
  assign n4699 = ~pi299 & ~n4698;
  assign n4700 = ~pi39 & ~n4699;
  assign n4701 = ~n4695 & n4700;
  assign n4702 = n4609 & ~n4624;
  assign n4703 = n4630 & n4637;
  assign n4704 = n4636 & ~n4703;
  assign n4705 = ~n4633 & n4704;
  assign n4706 = ~n4641 & ~n4705;
  assign n4707 = ~n4702 & n4706;
  assign n4708 = pi299 & ~n4707;
  assign n4709 = ~n4661 & ~n4708;
  assign n4710 = pi39 & ~n4709;
  assign n4711 = ~pi38 & ~n4710;
  assign n4712 = ~n4701 & n4711;
  assign n4713 = pi38 & n4674;
  assign n4714 = ~pi100 & ~n4713;
  assign n4715 = ~n4712 & n4714;
  assign n4716 = ~n4677 & ~n4715;
  assign n4717 = ~pi87 & ~n4716;
  assign n4718 = ~n3208 & n4674;
  assign n4719 = n3208 & n4709;
  assign n4720 = ~n4718 & ~n4719;
  assign n4721 = pi87 & n4720;
  assign n4722 = ~pi75 & ~n4721;
  assign n4723 = ~n4717 & n4722;
  assign n4724 = pi75 & n4674;
  assign n4725 = ~pi92 & ~n4724;
  assign n4726 = ~n4723 & n4725;
  assign n4727 = n3231 & ~n4720;
  assign n4728 = ~n3231 & n4674;
  assign n4729 = pi92 & ~n4728;
  assign n4730 = ~n4727 & n4729;
  assign n4731 = n3266 & ~n4730;
  assign n4732 = ~n4726 & n4731;
  assign n4733 = ~n3266 & n4674;
  assign n4734 = ~pi55 & ~n4733;
  assign n4735 = ~n4732 & n4734;
  assign n4736 = n3269 & n4707;
  assign n4737 = ~n3269 & ~n4672;
  assign n4738 = pi55 & ~n4737;
  assign n4739 = ~n4736 & n4738;
  assign n4740 = ~pi56 & ~n4739;
  assign n4741 = ~n4735 & n4740;
  assign n4742 = n3281 & ~n4707;
  assign n4743 = ~n3281 & n4672;
  assign n4744 = pi56 & ~n4743;
  assign n4745 = ~n4742 & n4744;
  assign n4746 = ~pi62 & ~n4745;
  assign n4747 = ~n4741 & n4746;
  assign n4748 = n3434 & n4707;
  assign n4749 = ~n3434 & ~n4672;
  assign n4750 = pi62 & ~n4749;
  assign n4751 = ~n4748 & n4750;
  assign n4752 = n3432 & ~n4751;
  assign n4753 = ~n4747 & n4752;
  assign n4754 = ~n3432 & ~n4672;
  assign n4755 = ~pi247 & ~n4754;
  assign n4756 = ~n4753 & n4755;
  assign n4757 = n4609 & ~n4635;
  assign n4758 = n4625 & n4637;
  assign n4759 = ~n4633 & n4636;
  assign n4760 = ~n4758 & n4759;
  assign n4761 = ~n4641 & ~n4760;
  assign n4762 = ~n4757 & n4761;
  assign n4763 = pi299 & ~n4762;
  assign n4764 = ~n3485 & ~n4660;
  assign n4765 = n3182 & n4764;
  assign n4766 = ~n4763 & n4765;
  assign n4767 = pi299 & ~n4671;
  assign n4768 = n4764 & ~n4767;
  assign n4769 = ~n3182 & n4768;
  assign n4770 = pi100 & ~n4769;
  assign n4771 = ~n4766 & n4770;
  assign n4772 = n3444 & n4653;
  assign n4773 = n4659 & ~n4772;
  assign n4774 = pi862 & ~n4679;
  assign n4775 = ~pi862 & n3467;
  assign n4776 = ~pi216 & ~n4775;
  assign n4777 = ~n4774 & n4776;
  assign n4778 = n4618 & ~n4777;
  assign n4779 = ~n4616 & ~n4778;
  assign n4780 = n4636 & ~n4779;
  assign n4781 = n4609 & ~n4689;
  assign n4782 = ~n4641 & ~n4781;
  assign n4783 = ~n4780 & n4782;
  assign n4784 = pi299 & ~n4783;
  assign n4785 = ~n4773 & ~n4784;
  assign n4786 = ~pi39 & ~n4785;
  assign n4787 = ~n4633 & n4669;
  assign n4788 = n4706 & ~n4787;
  assign n4789 = pi299 & ~n4788;
  assign n4790 = n4764 & ~n4789;
  assign n4791 = pi39 & ~n4790;
  assign n4792 = ~pi38 & ~n4791;
  assign n4793 = ~n4786 & n4792;
  assign n4794 = pi38 & n4768;
  assign n4795 = ~pi100 & ~n4794;
  assign n4796 = ~n4793 & n4795;
  assign n4797 = ~n4771 & ~n4796;
  assign n4798 = ~pi87 & ~n4797;
  assign n4799 = ~n3208 & n4768;
  assign n4800 = n3208 & n4790;
  assign n4801 = ~n4799 & ~n4800;
  assign n4802 = pi87 & n4801;
  assign n4803 = ~pi75 & ~n4802;
  assign n4804 = ~n4798 & n4803;
  assign n4805 = pi75 & n4768;
  assign n4806 = ~pi92 & ~n4805;
  assign n4807 = ~n4804 & n4806;
  assign n4808 = n3231 & ~n4801;
  assign n4809 = ~n3231 & n4768;
  assign n4810 = pi92 & ~n4809;
  assign n4811 = ~n4808 & n4810;
  assign n4812 = n3266 & ~n4811;
  assign n4813 = ~n4807 & n4812;
  assign n4814 = ~n3266 & n4768;
  assign n4815 = ~pi55 & ~n4814;
  assign n4816 = ~n4813 & n4815;
  assign n4817 = n3269 & n4788;
  assign n4818 = ~n3269 & n4671;
  assign n4819 = pi55 & ~n4818;
  assign n4820 = ~n4817 & n4819;
  assign n4821 = ~pi56 & ~n4820;
  assign n4822 = ~n4816 & n4821;
  assign n4823 = n3281 & ~n4788;
  assign n4824 = ~n3281 & ~n4671;
  assign n4825 = pi56 & ~n4824;
  assign n4826 = ~n4823 & n4825;
  assign n4827 = ~pi62 & ~n4826;
  assign n4828 = ~n4822 & n4827;
  assign n4829 = n3434 & n4788;
  assign n4830 = ~n3434 & n4671;
  assign n4831 = pi62 & ~n4830;
  assign n4832 = ~n4829 & n4831;
  assign n4833 = n3432 & ~n4832;
  assign n4834 = ~n4828 & n4833;
  assign n4835 = ~n3432 & n4671;
  assign n4836 = pi247 & ~n4835;
  assign n4837 = ~n4834 & n4836;
  assign po160 = n4756 | n4837;
  assign n4839 = pi215 & pi1138;
  assign n4840 = pi299 & ~n4839;
  assign n4841 = ~pi1138 & ~n2437;
  assign n4842 = ~pi940 & n2437;
  assign n4843 = pi221 & ~n4841;
  assign n4844 = ~n4842 & n4843;
  assign n4845 = pi216 & pi269;
  assign n4846 = ~pi221 & ~n4845;
  assign n4847 = pi877 & n3465;
  assign n4848 = ~pi169 & ~n4847;
  assign n4849 = pi169 & n3456;
  assign n4850 = ~n4848 & ~n4849;
  assign n4851 = pi877 & ~n4850;
  assign n4852 = ~n3367 & n4848;
  assign n4853 = ~n4851 & ~n4852;
  assign n4854 = ~pi228 & ~n4853;
  assign n4855 = pi877 & ~n2449;
  assign n4856 = pi105 & ~n4855;
  assign n4857 = ~pi105 & pi169;
  assign n4858 = pi228 & ~n4857;
  assign n4859 = ~n4856 & n4858;
  assign n4860 = ~n3463 & n4859;
  assign n4861 = ~pi216 & ~n4860;
  assign n4862 = ~n4854 & n4861;
  assign n4863 = n4846 & ~n4862;
  assign n4864 = ~n4844 & ~n4863;
  assign n4865 = ~pi215 & ~n4864;
  assign n4866 = n4840 & ~n4865;
  assign n4867 = pi223 & pi1138;
  assign n4868 = ~pi299 & ~n4867;
  assign n4869 = ~pi1138 & ~n3041;
  assign n4870 = ~pi940 & n3041;
  assign n4871 = pi222 & ~n4869;
  assign n4872 = ~n4870 & n4871;
  assign n4873 = pi224 & pi269;
  assign n4874 = ~pi222 & ~n4873;
  assign n4875 = pi877 & n3444;
  assign n4876 = ~pi224 & ~n4875;
  assign n4877 = n4874 & ~n4876;
  assign n4878 = ~n4872 & ~n4877;
  assign n4879 = n4868 & n4878;
  assign n4880 = ~n3444 & n4874;
  assign n4881 = n4878 & ~n4880;
  assign n4882 = ~pi223 & ~n4881;
  assign n4883 = n4868 & ~n4882;
  assign n4884 = ~pi39 & ~n4883;
  assign n4885 = ~n4879 & n4884;
  assign n4886 = ~n4866 & n4885;
  assign n4887 = ~pi224 & ~n4855;
  assign n4888 = n4874 & ~n4887;
  assign n4889 = ~n4872 & ~n4888;
  assign n4890 = ~pi223 & ~n4889;
  assign n4891 = ~n4867 & ~n4890;
  assign n4892 = ~pi299 & ~n4891;
  assign n4893 = ~pi216 & ~n4859;
  assign n4894 = ~pi877 & n3096;
  assign n4895 = ~pi169 & ~pi228;
  assign n4896 = ~n3322 & ~n4895;
  assign n4897 = ~n4894 & ~n4896;
  assign n4898 = n4893 & ~n4897;
  assign n4899 = n4846 & ~n4898;
  assign n4900 = ~n4844 & ~n4899;
  assign n4901 = ~pi215 & ~n4900;
  assign n4902 = ~n4839 & ~n4901;
  assign n4903 = pi299 & ~n4902;
  assign n4904 = ~n4892 & ~n4903;
  assign n4905 = pi39 & ~n4904;
  assign n4906 = ~pi38 & ~n4905;
  assign n4907 = ~n4886 & n4906;
  assign n4908 = n4893 & ~n4895;
  assign n4909 = n4846 & ~n4908;
  assign n4910 = ~n4844 & ~n4909;
  assign n4911 = ~pi215 & ~n4910;
  assign n4912 = ~n4839 & ~n4911;
  assign n4913 = pi299 & ~n4912;
  assign n4914 = ~n4892 & ~n4913;
  assign n4915 = pi38 & n4914;
  assign n4916 = ~pi100 & ~n4915;
  assign n4917 = ~n4907 & n4916;
  assign n4918 = ~pi877 & n3391;
  assign n4919 = ~n3600 & ~n4895;
  assign n4920 = ~n4918 & ~n4919;
  assign n4921 = n4893 & ~n4920;
  assign n4922 = n4846 & ~n4921;
  assign n4923 = ~n4844 & ~n4922;
  assign n4924 = ~pi215 & ~n4923;
  assign n4925 = ~n4839 & ~n4924;
  assign n4926 = pi299 & ~n4925;
  assign n4927 = n3182 & ~n4892;
  assign n4928 = ~n4926 & n4927;
  assign n4929 = ~n3182 & n4914;
  assign n4930 = pi100 & ~n4929;
  assign n4931 = ~n4928 & n4930;
  assign n4932 = ~n4917 & ~n4931;
  assign n4933 = ~pi87 & ~n4932;
  assign n4934 = ~n3208 & n4914;
  assign n4935 = n3208 & n4904;
  assign n4936 = ~n4934 & ~n4935;
  assign n4937 = pi87 & n4936;
  assign n4938 = ~pi75 & ~n4937;
  assign n4939 = ~n4933 & n4938;
  assign n4940 = pi75 & n4914;
  assign n4941 = ~pi92 & ~n4940;
  assign n4942 = ~n4939 & n4941;
  assign n4943 = n3231 & ~n4936;
  assign n4944 = ~n3231 & n4914;
  assign n4945 = pi92 & ~n4944;
  assign n4946 = ~n4943 & n4945;
  assign n4947 = n3266 & ~n4946;
  assign n4948 = ~n4942 & n4947;
  assign n4949 = ~n3266 & n4914;
  assign n4950 = ~pi55 & ~n4949;
  assign n4951 = ~n4948 & n4950;
  assign n4952 = n3269 & n4902;
  assign n4953 = ~n3269 & n4912;
  assign n4954 = pi55 & ~n4953;
  assign n4955 = ~n4952 & n4954;
  assign n4956 = ~pi56 & ~n4955;
  assign n4957 = ~n4951 & n4956;
  assign n4958 = n3281 & ~n4902;
  assign n4959 = ~n3281 & ~n4912;
  assign n4960 = pi56 & ~n4959;
  assign n4961 = ~n4958 & n4960;
  assign n4962 = ~pi62 & ~n4961;
  assign n4963 = ~n4957 & n4962;
  assign n4964 = n3434 & n4902;
  assign n4965 = ~n3434 & n4912;
  assign n4966 = pi62 & ~n4965;
  assign n4967 = ~n4964 & n4966;
  assign n4968 = ~pi246 & n3432;
  assign n4969 = ~n4967 & n4968;
  assign n4970 = ~n4963 & n4969;
  assign n4971 = ~pi877 & n3456;
  assign n4972 = ~pi169 & ~n4971;
  assign n4973 = pi877 & ~n3367;
  assign n4974 = ~pi877 & ~n3465;
  assign n4975 = pi169 & ~n4974;
  assign n4976 = ~n4973 & n4975;
  assign n4977 = ~n4972 & ~n4976;
  assign n4978 = ~pi228 & ~n4977;
  assign n4979 = ~n3729 & n4893;
  assign n4980 = ~n4978 & n4979;
  assign n4981 = n4846 & ~n4980;
  assign n4982 = ~n4844 & ~n4981;
  assign n4983 = ~pi215 & ~n4982;
  assign n4984 = n4840 & ~n4983;
  assign n4985 = n4884 & ~n4984;
  assign n4986 = ~n3485 & ~n4892;
  assign n4987 = ~n3475 & n4893;
  assign n4988 = ~n4897 & n4987;
  assign n4989 = n4846 & ~n4988;
  assign n4990 = ~n4844 & ~n4989;
  assign n4991 = ~pi215 & ~n4990;
  assign n4992 = ~n4839 & ~n4991;
  assign n4993 = pi299 & ~n4992;
  assign n4994 = n4986 & ~n4993;
  assign n4995 = pi39 & ~n4994;
  assign n4996 = ~pi38 & ~n4995;
  assign n4997 = ~n4985 & n4996;
  assign n4998 = n3592 & ~n4845;
  assign n4999 = n4912 & ~n4998;
  assign n5000 = pi299 & ~n4999;
  assign n5001 = n4986 & ~n5000;
  assign n5002 = pi38 & n5001;
  assign n5003 = ~pi100 & ~n5002;
  assign n5004 = ~n4997 & n5003;
  assign n5005 = ~n4920 & n4987;
  assign n5006 = n4846 & ~n5005;
  assign n5007 = ~n4844 & ~n5006;
  assign n5008 = ~pi215 & ~n5007;
  assign n5009 = ~n4839 & ~n5008;
  assign n5010 = pi299 & ~n5009;
  assign n5011 = n3182 & n4986;
  assign n5012 = ~n5010 & n5011;
  assign n5013 = ~n3182 & n5001;
  assign n5014 = pi100 & ~n5013;
  assign n5015 = ~n5012 & n5014;
  assign n5016 = ~n5004 & ~n5015;
  assign n5017 = ~pi87 & ~n5016;
  assign n5018 = ~n3208 & n5001;
  assign n5019 = n3208 & n4994;
  assign n5020 = ~n5018 & ~n5019;
  assign n5021 = pi87 & n5020;
  assign n5022 = ~pi75 & ~n5021;
  assign n5023 = ~n5017 & n5022;
  assign n5024 = pi75 & n5001;
  assign n5025 = ~pi92 & ~n5024;
  assign n5026 = ~n5023 & n5025;
  assign n5027 = n3231 & ~n5020;
  assign n5028 = ~n3231 & n5001;
  assign n5029 = pi92 & ~n5028;
  assign n5030 = ~n5027 & n5029;
  assign n5031 = n3266 & ~n5030;
  assign n5032 = ~n5026 & n5031;
  assign n5033 = ~n3266 & n5001;
  assign n5034 = ~pi55 & ~n5033;
  assign n5035 = ~n5032 & n5034;
  assign n5036 = n3269 & n4992;
  assign n5037 = ~n3269 & n4999;
  assign n5038 = pi55 & ~n5037;
  assign n5039 = ~n5036 & n5038;
  assign n5040 = ~pi56 & ~n5039;
  assign n5041 = ~n5035 & n5040;
  assign n5042 = n3281 & ~n4992;
  assign n5043 = ~n3281 & ~n4999;
  assign n5044 = pi56 & ~n5043;
  assign n5045 = ~n5042 & n5044;
  assign n5046 = ~pi62 & ~n5045;
  assign n5047 = ~n5041 & n5046;
  assign n5048 = n3434 & n4992;
  assign n5049 = ~n3434 & n4999;
  assign n5050 = pi62 & ~n5049;
  assign n5051 = ~n5048 & n5050;
  assign n5052 = pi246 & n3432;
  assign n5053 = ~n5051 & n5052;
  assign n5054 = ~n5047 & n5053;
  assign n5055 = pi246 & n4998;
  assign n5056 = ~n3432 & ~n5055;
  assign n5057 = n4912 & n5056;
  assign n5058 = ~n5054 & ~n5057;
  assign po161 = ~n4970 & n5058;
  assign n5060 = pi215 & pi1137;
  assign n5061 = pi299 & ~n5060;
  assign n5062 = ~pi1137 & ~n2437;
  assign n5063 = ~pi933 & n2437;
  assign n5064 = pi221 & ~n5062;
  assign n5065 = ~n5063 & n5064;
  assign n5066 = pi216 & pi280;
  assign n5067 = ~pi221 & ~n5066;
  assign n5068 = pi878 & n3465;
  assign n5069 = ~pi168 & ~n5068;
  assign n5070 = pi168 & n3456;
  assign n5071 = ~n5069 & ~n5070;
  assign n5072 = pi878 & ~n5071;
  assign n5073 = ~n3367 & n5069;
  assign n5074 = ~n5072 & ~n5073;
  assign n5075 = ~pi228 & ~n5074;
  assign n5076 = pi878 & ~n2449;
  assign n5077 = pi105 & ~n5076;
  assign n5078 = ~pi105 & pi168;
  assign n5079 = pi228 & ~n5078;
  assign n5080 = ~n5077 & n5079;
  assign n5081 = ~n3463 & n5080;
  assign n5082 = ~pi216 & ~n5081;
  assign n5083 = ~n5075 & n5082;
  assign n5084 = n5067 & ~n5083;
  assign n5085 = ~n5065 & ~n5084;
  assign n5086 = ~pi215 & ~n5085;
  assign n5087 = n5061 & ~n5086;
  assign n5088 = pi223 & pi1137;
  assign n5089 = ~pi299 & ~n5088;
  assign n5090 = ~pi1137 & ~n3041;
  assign n5091 = ~pi933 & n3041;
  assign n5092 = pi222 & ~n5090;
  assign n5093 = ~n5091 & n5092;
  assign n5094 = pi224 & pi280;
  assign n5095 = ~pi222 & ~n5094;
  assign n5096 = pi878 & n3444;
  assign n5097 = ~pi224 & ~n5096;
  assign n5098 = n5095 & ~n5097;
  assign n5099 = ~n5093 & ~n5098;
  assign n5100 = n5089 & n5099;
  assign n5101 = ~n3444 & n5095;
  assign n5102 = n5099 & ~n5101;
  assign n5103 = ~pi223 & ~n5102;
  assign n5104 = n5089 & ~n5103;
  assign n5105 = ~pi39 & ~n5104;
  assign n5106 = ~n5100 & n5105;
  assign n5107 = ~n5087 & n5106;
  assign n5108 = ~pi224 & ~n5076;
  assign n5109 = n5095 & ~n5108;
  assign n5110 = ~n5093 & ~n5109;
  assign n5111 = ~pi223 & ~n5110;
  assign n5112 = ~n5088 & ~n5111;
  assign n5113 = ~pi299 & ~n5112;
  assign n5114 = ~pi216 & ~n5080;
  assign n5115 = ~pi878 & n3096;
  assign n5116 = ~pi168 & ~pi228;
  assign n5117 = ~n3322 & ~n5116;
  assign n5118 = ~n5115 & ~n5117;
  assign n5119 = n5114 & ~n5118;
  assign n5120 = n5067 & ~n5119;
  assign n5121 = ~n5065 & ~n5120;
  assign n5122 = ~pi215 & ~n5121;
  assign n5123 = ~n5060 & ~n5122;
  assign n5124 = pi299 & ~n5123;
  assign n5125 = ~n5113 & ~n5124;
  assign n5126 = pi39 & ~n5125;
  assign n5127 = ~pi38 & ~n5126;
  assign n5128 = ~n5107 & n5127;
  assign n5129 = n5114 & ~n5116;
  assign n5130 = n5067 & ~n5129;
  assign n5131 = ~n5065 & ~n5130;
  assign n5132 = ~pi215 & ~n5131;
  assign n5133 = ~n5060 & ~n5132;
  assign n5134 = pi299 & ~n5133;
  assign n5135 = ~n5113 & ~n5134;
  assign n5136 = pi38 & n5135;
  assign n5137 = ~pi100 & ~n5136;
  assign n5138 = ~n5128 & n5137;
  assign n5139 = ~pi878 & n3391;
  assign n5140 = ~n3600 & ~n5116;
  assign n5141 = ~n5139 & ~n5140;
  assign n5142 = n5114 & ~n5141;
  assign n5143 = n5067 & ~n5142;
  assign n5144 = ~n5065 & ~n5143;
  assign n5145 = ~pi215 & ~n5144;
  assign n5146 = ~n5060 & ~n5145;
  assign n5147 = pi299 & ~n5146;
  assign n5148 = n3182 & ~n5113;
  assign n5149 = ~n5147 & n5148;
  assign n5150 = ~n3182 & n5135;
  assign n5151 = pi100 & ~n5150;
  assign n5152 = ~n5149 & n5151;
  assign n5153 = ~n5138 & ~n5152;
  assign n5154 = ~pi87 & ~n5153;
  assign n5155 = ~n3208 & n5135;
  assign n5156 = n3208 & n5125;
  assign n5157 = ~n5155 & ~n5156;
  assign n5158 = pi87 & n5157;
  assign n5159 = ~pi75 & ~n5158;
  assign n5160 = ~n5154 & n5159;
  assign n5161 = pi75 & n5135;
  assign n5162 = ~pi92 & ~n5161;
  assign n5163 = ~n5160 & n5162;
  assign n5164 = n3231 & ~n5157;
  assign n5165 = ~n3231 & n5135;
  assign n5166 = pi92 & ~n5165;
  assign n5167 = ~n5164 & n5166;
  assign n5168 = n3266 & ~n5167;
  assign n5169 = ~n5163 & n5168;
  assign n5170 = ~n3266 & n5135;
  assign n5171 = ~pi55 & ~n5170;
  assign n5172 = ~n5169 & n5171;
  assign n5173 = n3269 & n5123;
  assign n5174 = ~n3269 & n5133;
  assign n5175 = pi55 & ~n5174;
  assign n5176 = ~n5173 & n5175;
  assign n5177 = ~pi56 & ~n5176;
  assign n5178 = ~n5172 & n5177;
  assign n5179 = n3281 & ~n5123;
  assign n5180 = ~n3281 & ~n5133;
  assign n5181 = pi56 & ~n5180;
  assign n5182 = ~n5179 & n5181;
  assign n5183 = ~pi62 & ~n5182;
  assign n5184 = ~n5178 & n5183;
  assign n5185 = n3434 & n5123;
  assign n5186 = ~n3434 & n5133;
  assign n5187 = pi62 & ~n5186;
  assign n5188 = ~n5185 & n5187;
  assign n5189 = ~pi240 & n3432;
  assign n5190 = ~n5188 & n5189;
  assign n5191 = ~n5184 & n5190;
  assign n5192 = ~pi878 & n3456;
  assign n5193 = ~pi168 & ~n5192;
  assign n5194 = pi878 & ~n3367;
  assign n5195 = ~pi878 & ~n3465;
  assign n5196 = pi168 & ~n5195;
  assign n5197 = ~n5194 & n5196;
  assign n5198 = ~n5193 & ~n5197;
  assign n5199 = ~pi228 & ~n5198;
  assign n5200 = ~n3729 & n5114;
  assign n5201 = ~n5199 & n5200;
  assign n5202 = n5067 & ~n5201;
  assign n5203 = ~n5065 & ~n5202;
  assign n5204 = ~pi215 & ~n5203;
  assign n5205 = n5061 & ~n5204;
  assign n5206 = n5105 & ~n5205;
  assign n5207 = ~n3485 & ~n5113;
  assign n5208 = ~n3475 & n5114;
  assign n5209 = ~n5118 & n5208;
  assign n5210 = n5067 & ~n5209;
  assign n5211 = ~n5065 & ~n5210;
  assign n5212 = ~pi215 & ~n5211;
  assign n5213 = ~n5060 & ~n5212;
  assign n5214 = pi299 & ~n5213;
  assign n5215 = n5207 & ~n5214;
  assign n5216 = pi39 & ~n5215;
  assign n5217 = ~pi38 & ~n5216;
  assign n5218 = ~n5206 & n5217;
  assign n5219 = n3592 & ~n5066;
  assign n5220 = n5133 & ~n5219;
  assign n5221 = pi299 & ~n5220;
  assign n5222 = n5207 & ~n5221;
  assign n5223 = pi38 & n5222;
  assign n5224 = ~pi100 & ~n5223;
  assign n5225 = ~n5218 & n5224;
  assign n5226 = ~n5141 & n5208;
  assign n5227 = n5067 & ~n5226;
  assign n5228 = ~n5065 & ~n5227;
  assign n5229 = ~pi215 & ~n5228;
  assign n5230 = ~n5060 & ~n5229;
  assign n5231 = pi299 & ~n5230;
  assign n5232 = n3182 & n5207;
  assign n5233 = ~n5231 & n5232;
  assign n5234 = ~n3182 & n5222;
  assign n5235 = pi100 & ~n5234;
  assign n5236 = ~n5233 & n5235;
  assign n5237 = ~n5225 & ~n5236;
  assign n5238 = ~pi87 & ~n5237;
  assign n5239 = ~n3208 & n5222;
  assign n5240 = n3208 & n5215;
  assign n5241 = ~n5239 & ~n5240;
  assign n5242 = pi87 & n5241;
  assign n5243 = ~pi75 & ~n5242;
  assign n5244 = ~n5238 & n5243;
  assign n5245 = pi75 & n5222;
  assign n5246 = ~pi92 & ~n5245;
  assign n5247 = ~n5244 & n5246;
  assign n5248 = n3231 & ~n5241;
  assign n5249 = ~n3231 & n5222;
  assign n5250 = pi92 & ~n5249;
  assign n5251 = ~n5248 & n5250;
  assign n5252 = n3266 & ~n5251;
  assign n5253 = ~n5247 & n5252;
  assign n5254 = ~n3266 & n5222;
  assign n5255 = ~pi55 & ~n5254;
  assign n5256 = ~n5253 & n5255;
  assign n5257 = n3269 & n5213;
  assign n5258 = ~n3269 & n5220;
  assign n5259 = pi55 & ~n5258;
  assign n5260 = ~n5257 & n5259;
  assign n5261 = ~pi56 & ~n5260;
  assign n5262 = ~n5256 & n5261;
  assign n5263 = n3281 & ~n5213;
  assign n5264 = ~n3281 & ~n5220;
  assign n5265 = pi56 & ~n5264;
  assign n5266 = ~n5263 & n5265;
  assign n5267 = ~pi62 & ~n5266;
  assign n5268 = ~n5262 & n5267;
  assign n5269 = n3434 & n5213;
  assign n5270 = ~n3434 & n5220;
  assign n5271 = pi62 & ~n5270;
  assign n5272 = ~n5269 & n5271;
  assign n5273 = pi240 & n3432;
  assign n5274 = ~n5272 & n5273;
  assign n5275 = ~n5268 & n5274;
  assign n5276 = pi240 & n5219;
  assign n5277 = ~n3432 & ~n5276;
  assign n5278 = n5133 & n5277;
  assign n5279 = ~n5275 & ~n5278;
  assign po162 = ~n5191 & n5279;
  assign n5281 = ~pi1136 & ~n2437;
  assign n5282 = ~pi928 & n2437;
  assign n5283 = pi221 & ~n5281;
  assign n5284 = ~n5282 & n5283;
  assign n5285 = pi216 & pi266;
  assign n5286 = pi875 & ~n2449;
  assign n5287 = pi105 & ~n5286;
  assign n5288 = ~pi105 & ~pi166;
  assign n5289 = ~n5287 & ~n5288;
  assign n5290 = n3464 & ~n5289;
  assign n5291 = ~pi216 & ~n5290;
  assign n5292 = ~pi166 & ~n3456;
  assign n5293 = pi166 & n3465;
  assign n5294 = pi875 & ~n5293;
  assign n5295 = ~n5292 & n5294;
  assign n5296 = pi166 & ~pi875;
  assign n5297 = ~n3367 & n5296;
  assign n5298 = ~n5295 & ~n5297;
  assign n5299 = ~pi228 & ~n5298;
  assign n5300 = ~n3464 & ~n5299;
  assign n5301 = n5291 & ~n5300;
  assign n5302 = ~n5285 & ~n5301;
  assign n5303 = ~pi221 & ~n5302;
  assign n5304 = ~n5284 & ~n5303;
  assign n5305 = ~pi215 & ~n5304;
  assign n5306 = pi215 & pi1136;
  assign n5307 = pi299 & ~n5306;
  assign n5308 = ~n5305 & n5307;
  assign n5309 = ~pi224 & ~pi875;
  assign n5310 = ~n2449 & n5309;
  assign n5311 = pi224 & ~pi266;
  assign n5312 = ~pi222 & ~n5311;
  assign n5313 = ~n5310 & n5312;
  assign n5314 = n3053 & ~n3444;
  assign n5315 = n5313 & ~n5314;
  assign n5316 = ~pi1136 & ~n3041;
  assign n5317 = ~pi928 & n3041;
  assign n5318 = pi222 & ~n5316;
  assign n5319 = ~n5317 & n5318;
  assign n5320 = pi223 & pi1136;
  assign n5321 = ~pi299 & ~n5320;
  assign n5322 = ~n5319 & n5321;
  assign n5323 = ~n5315 & n5322;
  assign n5324 = ~n5313 & ~n5319;
  assign n5325 = ~n5314 & n5324;
  assign n5326 = ~pi223 & ~n5325;
  assign n5327 = n5321 & ~n5326;
  assign n5328 = ~pi39 & ~n5327;
  assign n5329 = ~n5323 & n5328;
  assign n5330 = ~n5308 & n5329;
  assign n5331 = ~pi223 & ~n5324;
  assign n5332 = ~n5320 & ~n5331;
  assign n5333 = ~pi299 & ~n5332;
  assign n5334 = n3101 & ~n5286;
  assign n5335 = n5333 & ~n5334;
  assign n5336 = pi228 & n5289;
  assign n5337 = ~pi875 & n3096;
  assign n5338 = pi166 & ~pi228;
  assign n5339 = ~n3322 & ~n5338;
  assign n5340 = ~n5337 & ~n5339;
  assign n5341 = ~n5336 & ~n5340;
  assign n5342 = ~pi216 & ~n5341;
  assign n5343 = ~n5285 & ~n5342;
  assign n5344 = ~pi221 & ~n5343;
  assign n5345 = ~n5284 & ~n5344;
  assign n5346 = ~pi215 & ~n5345;
  assign n5347 = ~n5306 & ~n5346;
  assign n5348 = pi299 & ~n5347;
  assign n5349 = ~n5335 & ~n5348;
  assign n5350 = pi39 & ~n5349;
  assign n5351 = ~pi38 & ~n5350;
  assign n5352 = ~n5330 & n5351;
  assign n5353 = ~n5336 & ~n5338;
  assign n5354 = ~pi216 & ~n5353;
  assign n5355 = ~n5285 & ~n5354;
  assign n5356 = ~pi221 & ~n5355;
  assign n5357 = ~n5284 & ~n5356;
  assign n5358 = ~pi215 & ~n5357;
  assign n5359 = ~n5306 & ~n5358;
  assign n5360 = pi299 & ~n5359;
  assign n5361 = ~n5335 & ~n5360;
  assign n5362 = pi38 & n5361;
  assign n5363 = ~pi100 & ~n5362;
  assign n5364 = ~n5352 & n5363;
  assign n5365 = ~pi875 & n3384;
  assign n5366 = pi166 & ~n5365;
  assign n5367 = ~n2447 & ~n3384;
  assign n5368 = n2447 & ~n3382;
  assign n5369 = pi875 & ~n5368;
  assign n5370 = ~n5367 & n5369;
  assign n5371 = ~n5366 & ~n5370;
  assign n5372 = ~pi228 & ~n5371;
  assign n5373 = ~n5336 & ~n5372;
  assign n5374 = ~pi216 & ~n5373;
  assign n5375 = ~n5285 & ~n5374;
  assign n5376 = ~pi221 & ~n5375;
  assign n5377 = ~n5284 & ~n5376;
  assign n5378 = ~pi215 & ~n5377;
  assign n5379 = ~n5306 & ~n5378;
  assign n5380 = pi299 & ~n5379;
  assign n5381 = n3182 & ~n5335;
  assign n5382 = ~n5380 & n5381;
  assign n5383 = ~n3182 & n5361;
  assign n5384 = pi100 & ~n5383;
  assign n5385 = ~n5382 & n5384;
  assign n5386 = ~n5364 & ~n5385;
  assign n5387 = ~pi87 & ~n5386;
  assign n5388 = ~n3208 & n5361;
  assign n5389 = n3208 & n5349;
  assign n5390 = ~n5388 & ~n5389;
  assign n5391 = pi87 & n5390;
  assign n5392 = ~pi75 & ~n5391;
  assign n5393 = ~n5387 & n5392;
  assign n5394 = pi75 & n5361;
  assign n5395 = ~pi92 & ~n5394;
  assign n5396 = ~n5393 & n5395;
  assign n5397 = n3231 & ~n5390;
  assign n5398 = ~n3231 & n5361;
  assign n5399 = pi92 & ~n5398;
  assign n5400 = ~n5397 & n5399;
  assign n5401 = n3266 & ~n5400;
  assign n5402 = ~n5396 & n5401;
  assign n5403 = ~n3266 & n5361;
  assign n5404 = ~pi55 & ~n5403;
  assign n5405 = ~n5402 & n5404;
  assign n5406 = n3269 & n5347;
  assign n5407 = ~n3269 & n5359;
  assign n5408 = pi55 & ~n5407;
  assign n5409 = ~n5406 & n5408;
  assign n5410 = ~pi56 & ~n5409;
  assign n5411 = ~n5405 & n5410;
  assign n5412 = n3281 & ~n5347;
  assign n5413 = ~n3281 & ~n5359;
  assign n5414 = pi56 & ~n5413;
  assign n5415 = ~n5412 & n5414;
  assign n5416 = ~pi62 & ~n5415;
  assign n5417 = ~n5411 & n5416;
  assign n5418 = n3434 & n5347;
  assign n5419 = ~n3434 & n5359;
  assign n5420 = pi62 & ~n5419;
  assign n5421 = ~n5418 & n5420;
  assign n5422 = n3432 & ~n5421;
  assign n5423 = ~n5417 & n5422;
  assign n5424 = ~n3432 & n5359;
  assign n5425 = ~pi245 & ~n5424;
  assign n5426 = ~n5423 & n5425;
  assign n5427 = pi166 & n3456;
  assign n5428 = ~pi166 & ~n3465;
  assign n5429 = ~pi875 & ~n5428;
  assign n5430 = ~n5427 & n5429;
  assign n5431 = ~pi166 & ~n3367;
  assign n5432 = pi875 & ~n5431;
  assign n5433 = ~pi228 & ~n5430;
  assign n5434 = ~n5432 & n5433;
  assign n5435 = n5291 & ~n5434;
  assign n5436 = ~n5285 & ~n5435;
  assign n5437 = ~pi221 & ~n5436;
  assign n5438 = ~n5284 & ~n5437;
  assign n5439 = ~pi215 & ~n5438;
  assign n5440 = n5307 & ~n5439;
  assign n5441 = n5328 & ~n5440;
  assign n5442 = ~n3475 & ~n5336;
  assign n5443 = ~n5340 & n5442;
  assign n5444 = ~pi216 & ~n5443;
  assign n5445 = ~n5285 & ~n5444;
  assign n5446 = ~pi221 & ~n5445;
  assign n5447 = ~n5284 & ~n5446;
  assign n5448 = ~pi215 & ~n5447;
  assign n5449 = ~n5306 & ~n5448;
  assign n5450 = pi299 & ~n5449;
  assign n5451 = ~n5333 & ~n5450;
  assign n5452 = pi39 & ~n5451;
  assign n5453 = ~pi38 & ~n5452;
  assign n5454 = ~n5441 & n5453;
  assign n5455 = ~n3476 & n5359;
  assign n5456 = pi299 & ~n5455;
  assign n5457 = ~n5333 & ~n5456;
  assign n5458 = pi38 & n5457;
  assign n5459 = ~pi100 & ~n5458;
  assign n5460 = ~n5454 & n5459;
  assign n5461 = ~n5372 & n5442;
  assign n5462 = ~pi216 & ~n5461;
  assign n5463 = ~n5285 & ~n5462;
  assign n5464 = ~pi221 & ~n5463;
  assign n5465 = ~n5284 & ~n5464;
  assign n5466 = ~pi215 & ~n5465;
  assign n5467 = ~n5306 & ~n5466;
  assign n5468 = pi299 & ~n5467;
  assign n5469 = n3182 & ~n5333;
  assign n5470 = ~n5468 & n5469;
  assign n5471 = ~n3182 & n5457;
  assign n5472 = pi100 & ~n5471;
  assign n5473 = ~n5470 & n5472;
  assign n5474 = ~n5460 & ~n5473;
  assign n5475 = ~pi87 & ~n5474;
  assign n5476 = ~n3208 & n5457;
  assign n5477 = n3208 & n5451;
  assign n5478 = ~n5476 & ~n5477;
  assign n5479 = pi87 & n5478;
  assign n5480 = ~pi75 & ~n5479;
  assign n5481 = ~n5475 & n5480;
  assign n5482 = pi75 & n5457;
  assign n5483 = ~pi92 & ~n5482;
  assign n5484 = ~n5481 & n5483;
  assign n5485 = n3231 & ~n5478;
  assign n5486 = ~n3231 & n5457;
  assign n5487 = pi92 & ~n5486;
  assign n5488 = ~n5485 & n5487;
  assign n5489 = n3266 & ~n5488;
  assign n5490 = ~n5484 & n5489;
  assign n5491 = ~n3266 & n5457;
  assign n5492 = ~pi55 & ~n5491;
  assign n5493 = ~n5490 & n5492;
  assign n5494 = n3269 & n5449;
  assign n5495 = ~n3269 & n5455;
  assign n5496 = pi55 & ~n5495;
  assign n5497 = ~n5494 & n5496;
  assign n5498 = ~pi56 & ~n5497;
  assign n5499 = ~n5493 & n5498;
  assign n5500 = n3281 & ~n5449;
  assign n5501 = ~n3281 & ~n5455;
  assign n5502 = pi56 & ~n5501;
  assign n5503 = ~n5500 & n5502;
  assign n5504 = ~pi62 & ~n5503;
  assign n5505 = ~n5499 & n5504;
  assign n5506 = n3434 & n5449;
  assign n5507 = ~n3434 & n5455;
  assign n5508 = pi62 & ~n5507;
  assign n5509 = ~n5506 & n5508;
  assign n5510 = n3432 & ~n5509;
  assign n5511 = ~n5505 & n5510;
  assign n5512 = ~n3432 & n5455;
  assign n5513 = pi245 & ~n5512;
  assign n5514 = ~n5511 & n5513;
  assign po163 = n5426 | n5514;
  assign n5516 = ~pi1135 & ~n2437;
  assign n5517 = ~pi938 & n2437;
  assign n5518 = pi221 & ~n5516;
  assign n5519 = ~n5517 & n5518;
  assign n5520 = pi216 & pi279;
  assign n5521 = pi879 & ~n2449;
  assign n5522 = pi105 & ~n5521;
  assign n5523 = ~pi105 & ~pi161;
  assign n5524 = ~n5522 & ~n5523;
  assign n5525 = n3464 & ~n5524;
  assign n5526 = ~pi216 & ~n5525;
  assign n5527 = ~pi161 & ~n3456;
  assign n5528 = pi161 & n3465;
  assign n5529 = pi879 & ~n5528;
  assign n5530 = ~n5527 & n5529;
  assign n5531 = pi161 & ~pi879;
  assign n5532 = ~n3367 & n5531;
  assign n5533 = ~n5530 & ~n5532;
  assign n5534 = ~pi228 & ~n5533;
  assign n5535 = ~n3464 & ~n5534;
  assign n5536 = n5526 & ~n5535;
  assign n5537 = ~n5520 & ~n5536;
  assign n5538 = ~pi221 & ~n5537;
  assign n5539 = ~n5519 & ~n5538;
  assign n5540 = ~pi215 & ~n5539;
  assign n5541 = pi215 & pi1135;
  assign n5542 = pi299 & ~n5541;
  assign n5543 = ~n5540 & n5542;
  assign n5544 = pi223 & pi1135;
  assign n5545 = ~pi299 & ~n5544;
  assign n5546 = ~pi1135 & ~n3041;
  assign n5547 = ~pi938 & n3041;
  assign n5548 = pi222 & ~n5546;
  assign n5549 = ~n5547 & n5548;
  assign n5550 = ~pi224 & ~pi879;
  assign n5551 = ~n2449 & n5550;
  assign n5552 = pi224 & ~pi279;
  assign n5553 = ~pi222 & ~n5552;
  assign n5554 = ~n5551 & n5553;
  assign n5555 = ~n5549 & ~n5554;
  assign n5556 = ~pi223 & ~n5555;
  assign n5557 = n5314 & ~n5549;
  assign n5558 = n5556 & ~n5557;
  assign n5559 = n5545 & ~n5558;
  assign n5560 = ~pi39 & ~n5559;
  assign n5561 = ~n5543 & n5560;
  assign n5562 = ~n5544 & ~n5556;
  assign n5563 = ~pi299 & ~n5562;
  assign n5564 = n3101 & ~n5521;
  assign n5565 = n5563 & ~n5564;
  assign n5566 = pi228 & n5524;
  assign n5567 = ~pi879 & n3096;
  assign n5568 = pi161 & ~pi228;
  assign n5569 = ~n3322 & ~n5568;
  assign n5570 = ~n5567 & ~n5569;
  assign n5571 = ~n5566 & ~n5570;
  assign n5572 = ~pi216 & ~n5571;
  assign n5573 = ~n5520 & ~n5572;
  assign n5574 = ~pi221 & ~n5573;
  assign n5575 = ~n5519 & ~n5574;
  assign n5576 = ~pi215 & ~n5575;
  assign n5577 = ~n5541 & ~n5576;
  assign n5578 = pi299 & ~n5577;
  assign n5579 = ~n5565 & ~n5578;
  assign n5580 = pi39 & ~n5579;
  assign n5581 = ~pi38 & ~n5580;
  assign n5582 = ~n5561 & n5581;
  assign n5583 = ~n5566 & ~n5568;
  assign n5584 = ~pi216 & ~n5583;
  assign n5585 = ~n5520 & ~n5584;
  assign n5586 = ~pi221 & ~n5585;
  assign n5587 = ~n5519 & ~n5586;
  assign n5588 = ~pi215 & ~n5587;
  assign n5589 = ~n5541 & ~n5588;
  assign n5590 = pi299 & ~n5589;
  assign n5591 = ~n5565 & ~n5590;
  assign n5592 = pi38 & n5591;
  assign n5593 = ~pi100 & ~n5592;
  assign n5594 = ~n5582 & n5593;
  assign n5595 = ~pi879 & n3384;
  assign n5596 = pi161 & ~n5595;
  assign n5597 = ~pi152 & ~pi166;
  assign n5598 = ~n3384 & ~n5597;
  assign n5599 = ~n3382 & n5597;
  assign n5600 = pi879 & ~n5599;
  assign n5601 = ~n5598 & n5600;
  assign n5602 = ~n5596 & ~n5601;
  assign n5603 = ~pi228 & ~n5602;
  assign n5604 = ~n5566 & ~n5603;
  assign n5605 = ~pi216 & ~n5604;
  assign n5606 = ~n5520 & ~n5605;
  assign n5607 = ~pi221 & ~n5606;
  assign n5608 = ~n5519 & ~n5607;
  assign n5609 = ~pi215 & ~n5608;
  assign n5610 = ~n5541 & ~n5609;
  assign n5611 = pi299 & ~n5610;
  assign n5612 = n3182 & ~n5565;
  assign n5613 = ~n5611 & n5612;
  assign n5614 = ~n3182 & n5591;
  assign n5615 = pi100 & ~n5614;
  assign n5616 = ~n5613 & n5615;
  assign n5617 = ~n5594 & ~n5616;
  assign n5618 = ~pi87 & ~n5617;
  assign n5619 = ~n3208 & n5591;
  assign n5620 = n3208 & n5579;
  assign n5621 = ~n5619 & ~n5620;
  assign n5622 = pi87 & n5621;
  assign n5623 = ~pi75 & ~n5622;
  assign n5624 = ~n5618 & n5623;
  assign n5625 = pi75 & n5591;
  assign n5626 = ~pi92 & ~n5625;
  assign n5627 = ~n5624 & n5626;
  assign n5628 = n3231 & ~n5621;
  assign n5629 = ~n3231 & n5591;
  assign n5630 = pi92 & ~n5629;
  assign n5631 = ~n5628 & n5630;
  assign n5632 = n3266 & ~n5631;
  assign n5633 = ~n5627 & n5632;
  assign n5634 = ~n3266 & n5591;
  assign n5635 = ~pi55 & ~n5634;
  assign n5636 = ~n5633 & n5635;
  assign n5637 = n3269 & n5577;
  assign n5638 = ~n3269 & n5589;
  assign n5639 = pi55 & ~n5638;
  assign n5640 = ~n5637 & n5639;
  assign n5641 = ~pi56 & ~n5640;
  assign n5642 = ~n5636 & n5641;
  assign n5643 = n3281 & ~n5577;
  assign n5644 = ~n3281 & ~n5589;
  assign n5645 = pi56 & ~n5644;
  assign n5646 = ~n5643 & n5645;
  assign n5647 = ~pi62 & ~n5646;
  assign n5648 = ~n5642 & n5647;
  assign n5649 = n3434 & n5577;
  assign n5650 = ~n3434 & n5589;
  assign n5651 = pi62 & ~n5650;
  assign n5652 = ~n5649 & n5651;
  assign n5653 = n3432 & ~n5652;
  assign n5654 = ~n5648 & n5653;
  assign n5655 = ~n3432 & n5589;
  assign n5656 = ~pi244 & ~n5655;
  assign n5657 = ~n5654 & n5656;
  assign n5658 = pi161 & n3456;
  assign n5659 = ~pi161 & ~n3465;
  assign n5660 = ~pi879 & ~n5659;
  assign n5661 = ~n5658 & n5660;
  assign n5662 = ~pi161 & ~n3367;
  assign n5663 = pi879 & ~n5662;
  assign n5664 = ~pi228 & ~n5661;
  assign n5665 = ~n5663 & n5664;
  assign n5666 = n5526 & ~n5665;
  assign n5667 = ~n5520 & ~n5666;
  assign n5668 = ~pi221 & ~n5667;
  assign n5669 = ~n5519 & ~n5668;
  assign n5670 = ~pi215 & ~n5669;
  assign n5671 = n5542 & ~n5670;
  assign n5672 = ~n5314 & n5555;
  assign n5673 = ~pi223 & ~n5672;
  assign n5674 = n5545 & ~n5673;
  assign n5675 = ~pi39 & ~n5674;
  assign n5676 = ~n5671 & n5675;
  assign n5677 = ~n3475 & ~n5566;
  assign n5678 = ~n5570 & n5677;
  assign n5679 = ~pi216 & ~n5678;
  assign n5680 = ~n5520 & ~n5679;
  assign n5681 = ~pi221 & ~n5680;
  assign n5682 = ~n5519 & ~n5681;
  assign n5683 = ~pi215 & ~n5682;
  assign n5684 = ~n5541 & ~n5683;
  assign n5685 = pi299 & ~n5684;
  assign n5686 = ~n5563 & ~n5685;
  assign n5687 = pi39 & ~n5686;
  assign n5688 = ~pi38 & ~n5687;
  assign n5689 = ~n5676 & n5688;
  assign n5690 = ~n3476 & n5589;
  assign n5691 = pi299 & ~n5690;
  assign n5692 = ~n5563 & ~n5691;
  assign n5693 = pi38 & n5692;
  assign n5694 = ~pi100 & ~n5693;
  assign n5695 = ~n5689 & n5694;
  assign n5696 = ~n5603 & n5677;
  assign n5697 = ~pi216 & ~n5696;
  assign n5698 = ~n5520 & ~n5697;
  assign n5699 = ~pi221 & ~n5698;
  assign n5700 = ~n5519 & ~n5699;
  assign n5701 = ~pi215 & ~n5700;
  assign n5702 = ~n5541 & ~n5701;
  assign n5703 = pi299 & ~n5702;
  assign n5704 = n3182 & ~n5563;
  assign n5705 = ~n5703 & n5704;
  assign n5706 = ~n3182 & n5692;
  assign n5707 = pi100 & ~n5706;
  assign n5708 = ~n5705 & n5707;
  assign n5709 = ~n5695 & ~n5708;
  assign n5710 = ~pi87 & ~n5709;
  assign n5711 = ~n3208 & n5692;
  assign n5712 = n3208 & n5686;
  assign n5713 = ~n5711 & ~n5712;
  assign n5714 = pi87 & n5713;
  assign n5715 = ~pi75 & ~n5714;
  assign n5716 = ~n5710 & n5715;
  assign n5717 = pi75 & n5692;
  assign n5718 = ~pi92 & ~n5717;
  assign n5719 = ~n5716 & n5718;
  assign n5720 = n3231 & ~n5713;
  assign n5721 = ~n3231 & n5692;
  assign n5722 = pi92 & ~n5721;
  assign n5723 = ~n5720 & n5722;
  assign n5724 = n3266 & ~n5723;
  assign n5725 = ~n5719 & n5724;
  assign n5726 = ~n3266 & n5692;
  assign n5727 = ~pi55 & ~n5726;
  assign n5728 = ~n5725 & n5727;
  assign n5729 = n3269 & n5684;
  assign n5730 = ~n3269 & n5690;
  assign n5731 = pi55 & ~n5730;
  assign n5732 = ~n5729 & n5731;
  assign n5733 = ~pi56 & ~n5732;
  assign n5734 = ~n5728 & n5733;
  assign n5735 = n3281 & ~n5684;
  assign n5736 = ~n3281 & ~n5690;
  assign n5737 = pi56 & ~n5736;
  assign n5738 = ~n5735 & n5737;
  assign n5739 = ~pi62 & ~n5738;
  assign n5740 = ~n5734 & n5739;
  assign n5741 = n3434 & n5684;
  assign n5742 = ~n3434 & n5690;
  assign n5743 = pi62 & ~n5742;
  assign n5744 = ~n5741 & n5743;
  assign n5745 = n3432 & ~n5744;
  assign n5746 = ~n5740 & n5745;
  assign n5747 = ~n3432 & n5690;
  assign n5748 = pi244 & ~n5747;
  assign n5749 = ~n5746 & n5748;
  assign po164 = n5657 | n5749;
  assign n5751 = pi833 & ~pi930;
  assign n5752 = ~pi216 & pi221;
  assign n5753 = n5751 & n5752;
  assign n5754 = pi216 & pi278;
  assign n5755 = ~pi221 & ~n5754;
  assign n5756 = ~pi105 & pi152;
  assign n5757 = pi228 & ~n5756;
  assign n5758 = ~pi846 & n3444;
  assign n5759 = pi105 & ~n5758;
  assign n5760 = n5757 & ~n5759;
  assign n5761 = ~pi216 & ~n5760;
  assign n5762 = pi152 & ~n3456;
  assign n5763 = ~pi152 & n3465;
  assign n5764 = ~pi846 & ~n5763;
  assign n5765 = ~n5762 & n5764;
  assign n5766 = ~pi152 & pi846;
  assign n5767 = ~n3367 & n5766;
  assign n5768 = ~n5765 & ~n5767;
  assign n5769 = ~pi228 & ~n5768;
  assign n5770 = n5761 & ~n5769;
  assign n5771 = n5755 & ~n5770;
  assign n5772 = ~n5753 & ~n5771;
  assign n5773 = pi221 & ~n2437;
  assign n5774 = ~pi215 & pi299;
  assign n5775 = ~n5773 & n5774;
  assign n5776 = n5772 & n5775;
  assign n5777 = pi222 & ~pi224;
  assign n5778 = n5751 & n5777;
  assign n5779 = pi224 & pi278;
  assign n5780 = ~pi222 & ~n5779;
  assign n5781 = ~pi224 & ~n5758;
  assign n5782 = n5780 & ~n5781;
  assign n5783 = ~n5778 & ~n5782;
  assign n5784 = ~n3042 & n3483;
  assign n5785 = n5783 & n5784;
  assign n5786 = ~pi39 & ~n5785;
  assign n5787 = ~n5776 & n5786;
  assign n5788 = pi846 & ~n2449;
  assign n5789 = ~pi224 & n5788;
  assign n5790 = n5780 & ~n5789;
  assign n5791 = n3043 & ~n5778;
  assign n5792 = ~n5790 & n5791;
  assign n5793 = ~pi299 & ~n5792;
  assign n5794 = ~n3763 & n5793;
  assign n5795 = ~pi215 & ~n5773;
  assign n5796 = ~n5753 & n5795;
  assign n5797 = pi105 & n5788;
  assign n5798 = ~n5756 & ~n5797;
  assign n5799 = pi228 & ~n5798;
  assign n5800 = ~n3475 & ~n5799;
  assign n5801 = ~pi846 & n3096;
  assign n5802 = pi152 & ~pi228;
  assign n5803 = ~n3322 & ~n5802;
  assign n5804 = ~n5801 & ~n5803;
  assign n5805 = n5800 & ~n5804;
  assign n5806 = ~pi216 & ~n5805;
  assign n5807 = n5755 & ~n5806;
  assign n5808 = n5796 & ~n5807;
  assign n5809 = pi299 & ~n5808;
  assign n5810 = ~n5794 & ~n5809;
  assign n5811 = pi39 & ~n5810;
  assign n5812 = ~pi38 & ~n5811;
  assign n5813 = ~n5787 & n5812;
  assign n5814 = ~n5799 & ~n5802;
  assign n5815 = ~pi216 & ~n5814;
  assign n5816 = n5755 & ~n5815;
  assign n5817 = n5796 & ~n5816;
  assign n5818 = ~n3476 & ~n5817;
  assign n5819 = pi299 & n5818;
  assign n5820 = ~n5794 & ~n5819;
  assign n5821 = pi38 & n5820;
  assign n5822 = ~pi100 & ~n5821;
  assign n5823 = ~n5813 & n5822;
  assign n5824 = pi846 & ~n3390;
  assign n5825 = ~n3385 & ~n5824;
  assign n5826 = ~pi228 & ~n5825;
  assign n5827 = n5800 & ~n5826;
  assign n5828 = ~pi216 & ~n5827;
  assign n5829 = n5755 & ~n5828;
  assign n5830 = n5796 & ~n5829;
  assign n5831 = pi299 & ~n5830;
  assign n5832 = n3182 & ~n5794;
  assign n5833 = ~n5831 & n5832;
  assign n5834 = ~n3182 & n5820;
  assign n5835 = pi100 & ~n5834;
  assign n5836 = ~n5833 & n5835;
  assign n5837 = ~n5823 & ~n5836;
  assign n5838 = ~pi87 & ~n5837;
  assign n5839 = ~n3208 & n5820;
  assign n5840 = n3208 & n5810;
  assign n5841 = ~n5839 & ~n5840;
  assign n5842 = pi87 & n5841;
  assign n5843 = ~pi75 & ~n5842;
  assign n5844 = ~n5838 & n5843;
  assign n5845 = pi75 & n5820;
  assign n5846 = ~pi92 & ~n5845;
  assign n5847 = ~n5844 & n5846;
  assign n5848 = n3231 & ~n5841;
  assign n5849 = ~n3231 & n5820;
  assign n5850 = pi92 & ~n5849;
  assign n5851 = ~n5848 & n5850;
  assign n5852 = n3266 & ~n5851;
  assign n5853 = ~n5847 & n5852;
  assign n5854 = ~n3266 & n5820;
  assign n5855 = ~pi55 & ~n5854;
  assign n5856 = ~n5853 & n5855;
  assign n5857 = n3269 & n5808;
  assign n5858 = ~n3269 & ~n5818;
  assign n5859 = pi55 & ~n5858;
  assign n5860 = ~n5857 & n5859;
  assign n5861 = ~pi56 & ~n5860;
  assign n5862 = ~n5856 & n5861;
  assign n5863 = n3281 & ~n5808;
  assign n5864 = ~n3281 & n5818;
  assign n5865 = pi56 & ~n5864;
  assign n5866 = ~n5863 & n5865;
  assign n5867 = ~pi62 & ~n5866;
  assign n5868 = ~n5862 & n5867;
  assign n5869 = n3434 & n5808;
  assign n5870 = ~n3434 & ~n5818;
  assign n5871 = pi62 & ~n5870;
  assign n5872 = ~n5869 & n5871;
  assign n5873 = n3432 & ~n5872;
  assign n5874 = ~n5868 & n5873;
  assign n5875 = ~n3432 & ~n5818;
  assign n5876 = pi242 & ~n5875;
  assign n5877 = ~n5874 & n5876;
  assign n5878 = ~pi152 & ~n3456;
  assign n5879 = pi152 & n3465;
  assign n5880 = pi846 & ~n5879;
  assign n5881 = ~n5878 & n5880;
  assign n5882 = pi152 & ~pi846;
  assign n5883 = ~n3367 & n5882;
  assign n5884 = ~pi228 & ~n5883;
  assign n5885 = ~n5881 & n5884;
  assign n5886 = ~n3444 & n5757;
  assign n5887 = n5761 & ~n5886;
  assign n5888 = ~n5885 & n5887;
  assign n5889 = n5755 & ~n5888;
  assign n5890 = ~n5753 & ~n5889;
  assign n5891 = n5775 & n5890;
  assign n5892 = ~n3443 & n5789;
  assign n5893 = n5780 & ~n5892;
  assign n5894 = ~n5778 & n5784;
  assign n5895 = ~n5893 & n5894;
  assign n5896 = ~pi39 & ~n5895;
  assign n5897 = ~n5891 & n5896;
  assign n5898 = ~n5799 & ~n5804;
  assign n5899 = ~pi216 & ~n5898;
  assign n5900 = n5755 & ~n5899;
  assign n5901 = n5796 & ~n5900;
  assign n5902 = pi299 & ~n5901;
  assign n5903 = ~n5793 & ~n5902;
  assign n5904 = pi39 & ~n5903;
  assign n5905 = ~pi38 & ~n5904;
  assign n5906 = ~n5897 & n5905;
  assign n5907 = pi299 & ~n5817;
  assign n5908 = ~n5793 & ~n5907;
  assign n5909 = pi38 & n5908;
  assign n5910 = ~pi100 & ~n5909;
  assign n5911 = ~n5906 & n5910;
  assign n5912 = ~n5799 & ~n5826;
  assign n5913 = ~pi216 & ~n5912;
  assign n5914 = n5755 & ~n5913;
  assign n5915 = n5796 & ~n5914;
  assign n5916 = pi299 & ~n5915;
  assign n5917 = n3182 & ~n5793;
  assign n5918 = ~n5916 & n5917;
  assign n5919 = ~n3182 & n5908;
  assign n5920 = pi100 & ~n5919;
  assign n5921 = ~n5918 & n5920;
  assign n5922 = ~n5911 & ~n5921;
  assign n5923 = ~pi87 & ~n5922;
  assign n5924 = ~n3208 & n5908;
  assign n5925 = n3208 & n5903;
  assign n5926 = ~n5924 & ~n5925;
  assign n5927 = pi87 & n5926;
  assign n5928 = ~pi75 & ~n5927;
  assign n5929 = ~n5923 & n5928;
  assign n5930 = pi75 & n5908;
  assign n5931 = ~pi92 & ~n5930;
  assign n5932 = ~n5929 & n5931;
  assign n5933 = n3231 & ~n5926;
  assign n5934 = ~n3231 & n5908;
  assign n5935 = pi92 & ~n5934;
  assign n5936 = ~n5933 & n5935;
  assign n5937 = n3266 & ~n5936;
  assign n5938 = ~n5932 & n5937;
  assign n5939 = ~n3266 & n5908;
  assign n5940 = ~pi55 & ~n5939;
  assign n5941 = ~n5938 & n5940;
  assign n5942 = n3269 & n5901;
  assign n5943 = ~n3269 & n5817;
  assign n5944 = pi55 & ~n5943;
  assign n5945 = ~n5942 & n5944;
  assign n5946 = ~pi56 & ~n5945;
  assign n5947 = ~n5941 & n5946;
  assign n5948 = n3281 & ~n5901;
  assign n5949 = ~n3281 & ~n5817;
  assign n5950 = pi56 & ~n5949;
  assign n5951 = ~n5948 & n5950;
  assign n5952 = ~pi62 & ~n5951;
  assign n5953 = ~n5947 & n5952;
  assign n5954 = n3434 & n5901;
  assign n5955 = ~n3434 & n5817;
  assign n5956 = pi62 & ~n5955;
  assign n5957 = ~n5954 & n5956;
  assign n5958 = n3432 & ~n5957;
  assign n5959 = ~n5953 & n5958;
  assign n5960 = ~n3432 & n5817;
  assign n5961 = ~pi242 & ~n5960;
  assign n5962 = ~n5959 & n5961;
  assign n5963 = ~n5877 & ~n5962;
  assign n5964 = ~pi1134 & ~n5963;
  assign n5965 = n3483 & ~n5783;
  assign n5966 = ~pi39 & ~n5965;
  assign n5967 = ~n5772 & n5774;
  assign n5968 = n5966 & ~n5967;
  assign n5969 = n3043 & n5794;
  assign n5970 = ~pi299 & ~n5969;
  assign n5971 = ~n5753 & ~n5807;
  assign n5972 = ~pi215 & ~n5971;
  assign n5973 = pi299 & ~n5972;
  assign n5974 = ~n5970 & ~n5973;
  assign n5975 = pi39 & ~n5974;
  assign n5976 = ~pi38 & ~n5975;
  assign n5977 = ~n5968 & n5976;
  assign n5978 = ~n5753 & ~n5816;
  assign n5979 = ~pi215 & ~n5978;
  assign n5980 = ~n3476 & n5979;
  assign n5981 = pi299 & ~n5980;
  assign n5982 = ~n5970 & ~n5981;
  assign n5983 = pi38 & n5982;
  assign n5984 = ~pi100 & ~n5983;
  assign n5985 = ~n5977 & n5984;
  assign n5986 = ~n5753 & ~n5829;
  assign n5987 = ~pi215 & ~n5986;
  assign n5988 = pi299 & ~n5987;
  assign n5989 = n3182 & ~n5970;
  assign n5990 = ~n5988 & n5989;
  assign n5991 = ~n3182 & n5982;
  assign n5992 = pi100 & ~n5991;
  assign n5993 = ~n5990 & n5992;
  assign n5994 = ~n5985 & ~n5993;
  assign n5995 = ~pi87 & ~n5994;
  assign n5996 = ~n3208 & n5982;
  assign n5997 = n3208 & n5974;
  assign n5998 = ~n5996 & ~n5997;
  assign n5999 = pi87 & n5998;
  assign n6000 = ~pi75 & ~n5999;
  assign n6001 = ~n5995 & n6000;
  assign n6002 = pi75 & n5982;
  assign n6003 = ~pi92 & ~n6002;
  assign n6004 = ~n6001 & n6003;
  assign n6005 = n3231 & ~n5998;
  assign n6006 = ~n3231 & n5982;
  assign n6007 = pi92 & ~n6006;
  assign n6008 = ~n6005 & n6007;
  assign n6009 = n3266 & ~n6008;
  assign n6010 = ~n6004 & n6009;
  assign n6011 = ~n3266 & n5982;
  assign n6012 = ~pi55 & ~n6011;
  assign n6013 = ~n6010 & n6012;
  assign n6014 = n3269 & n5972;
  assign n6015 = ~n3269 & n5980;
  assign n6016 = pi55 & ~n6015;
  assign n6017 = ~n6014 & n6016;
  assign n6018 = ~pi56 & ~n6017;
  assign n6019 = ~n6013 & n6018;
  assign n6020 = n3281 & ~n5972;
  assign n6021 = ~n3281 & ~n5980;
  assign n6022 = pi56 & ~n6021;
  assign n6023 = ~n6020 & n6022;
  assign n6024 = ~pi62 & ~n6023;
  assign n6025 = ~n6019 & n6024;
  assign n6026 = n3434 & n5972;
  assign n6027 = ~n3434 & n5980;
  assign n6028 = pi62 & ~n6027;
  assign n6029 = ~n6026 & n6028;
  assign n6030 = n3432 & ~n6029;
  assign n6031 = ~n6025 & n6030;
  assign n6032 = ~n3432 & n5980;
  assign n6033 = pi242 & ~n6032;
  assign n6034 = ~n6031 & n6033;
  assign n6035 = n5774 & ~n5890;
  assign n6036 = n3483 & n5893;
  assign n6037 = n5966 & ~n6036;
  assign n6038 = ~n6035 & n6037;
  assign n6039 = ~pi223 & n5790;
  assign n6040 = n5970 & ~n6039;
  assign n6041 = ~n5753 & ~n5900;
  assign n6042 = ~pi215 & ~n6041;
  assign n6043 = pi299 & ~n6042;
  assign n6044 = ~n6040 & ~n6043;
  assign n6045 = pi39 & ~n6044;
  assign n6046 = ~pi38 & ~n6045;
  assign n6047 = ~n6038 & n6046;
  assign n6048 = pi299 & ~n5979;
  assign n6049 = ~n6040 & ~n6048;
  assign n6050 = pi38 & n6049;
  assign n6051 = ~pi100 & ~n6050;
  assign n6052 = ~n6047 & n6051;
  assign n6053 = ~n5753 & ~n5914;
  assign n6054 = ~pi215 & ~n6053;
  assign n6055 = pi299 & ~n6054;
  assign n6056 = n3182 & ~n6040;
  assign n6057 = ~n6055 & n6056;
  assign n6058 = ~n3182 & n6049;
  assign n6059 = pi100 & ~n6058;
  assign n6060 = ~n6057 & n6059;
  assign n6061 = ~n6052 & ~n6060;
  assign n6062 = ~pi87 & ~n6061;
  assign n6063 = ~n3208 & n6049;
  assign n6064 = n3208 & n6044;
  assign n6065 = ~n6063 & ~n6064;
  assign n6066 = pi87 & n6065;
  assign n6067 = ~pi75 & ~n6066;
  assign n6068 = ~n6062 & n6067;
  assign n6069 = pi75 & n6049;
  assign n6070 = ~pi92 & ~n6069;
  assign n6071 = ~n6068 & n6070;
  assign n6072 = n3231 & ~n6065;
  assign n6073 = ~n3231 & n6049;
  assign n6074 = pi92 & ~n6073;
  assign n6075 = ~n6072 & n6074;
  assign n6076 = n3266 & ~n6075;
  assign n6077 = ~n6071 & n6076;
  assign n6078 = ~n3266 & n6049;
  assign n6079 = ~pi55 & ~n6078;
  assign n6080 = ~n6077 & n6079;
  assign n6081 = n3269 & n6042;
  assign n6082 = ~n3269 & n5979;
  assign n6083 = pi55 & ~n6082;
  assign n6084 = ~n6081 & n6083;
  assign n6085 = ~pi56 & ~n6084;
  assign n6086 = ~n6080 & n6085;
  assign n6087 = n3281 & ~n6042;
  assign n6088 = ~n3281 & ~n5979;
  assign n6089 = pi56 & ~n6088;
  assign n6090 = ~n6087 & n6089;
  assign n6091 = ~pi62 & ~n6090;
  assign n6092 = ~n6086 & n6091;
  assign n6093 = n3434 & n6042;
  assign n6094 = ~n3434 & n5979;
  assign n6095 = pi62 & ~n6094;
  assign n6096 = ~n6093 & n6095;
  assign n6097 = n3432 & ~n6096;
  assign n6098 = ~n6092 & n6097;
  assign n6099 = ~n3432 & n5979;
  assign n6100 = ~pi242 & ~n6099;
  assign n6101 = ~n6098 & n6100;
  assign n6102 = pi1134 & ~n6101;
  assign n6103 = ~n6034 & n6102;
  assign po165 = ~n5964 & ~n6103;
  assign n6105 = pi57 & pi59;
  assign n6106 = n3096 & n3295;
  assign n6107 = ~n3432 & ~n6106;
  assign n6108 = ~n6105 & ~n6107;
  assign n6109 = pi57 & ~n6108;
  assign n6110 = n3090 & n3208;
  assign n6111 = n3280 & n6110;
  assign n6112 = pi56 & ~n6111;
  assign n6113 = ~pi54 & n3278;
  assign n6114 = n6110 & n6113;
  assign n6115 = pi74 & ~n6114;
  assign n6116 = ~pi55 & ~n6115;
  assign n6117 = ~pi39 & n3090;
  assign n6118 = pi38 & ~n6117;
  assign n6119 = ~pi100 & ~n6118;
  assign n6120 = pi58 & n2521;
  assign n6121 = ~pi90 & ~n6120;
  assign n6122 = n2505 & n2578;
  assign n6123 = n2684 & n6122;
  assign n6124 = n2590 & ~n6123;
  assign n6125 = ~n2585 & ~n6124;
  assign n6126 = ~pi108 & ~n6125;
  assign n6127 = n2584 & ~n6126;
  assign n6128 = ~pi110 & n2699;
  assign n6129 = ~n6127 & n6128;
  assign n6130 = ~n2568 & ~n2575;
  assign n6131 = ~n6129 & n6130;
  assign n6132 = ~pi47 & ~n6131;
  assign n6133 = n2489 & ~n2571;
  assign n6134 = ~n6132 & n6133;
  assign n6135 = n6121 & ~n6134;
  assign n6136 = ~n2706 & ~n6135;
  assign n6137 = ~pi93 & ~n6136;
  assign n6138 = ~pi841 & n2522;
  assign n6139 = pi93 & ~n6138;
  assign n6140 = ~n6137 & ~n6139;
  assign n6141 = ~pi35 & ~n6140;
  assign n6142 = ~pi70 & ~n2524;
  assign n6143 = ~n6141 & n6142;
  assign n6144 = ~pi51 & ~n6143;
  assign n6145 = n2559 & ~n6144;
  assign n6146 = n2920 & ~n6145;
  assign n6147 = n2556 & ~n6146;
  assign n6148 = n2554 & ~n6147;
  assign n6149 = ~pi198 & ~pi299;
  assign n6150 = ~pi210 & pi299;
  assign n6151 = ~n6149 & ~n6150;
  assign n6152 = ~pi35 & n2551;
  assign n6153 = ~pi40 & n6152;
  assign n6154 = n2736 & n6153;
  assign n6155 = pi32 & ~n6154;
  assign n6156 = ~n6151 & ~n6155;
  assign n6157 = ~n3363 & n6151;
  assign n6158 = ~n6156 & ~n6157;
  assign n6159 = ~n6148 & ~n6158;
  assign n6160 = ~pi95 & ~n6159;
  assign n6161 = ~n2727 & ~n6160;
  assign n6162 = ~pi39 & ~n6161;
  assign n6163 = pi603 & ~pi642;
  assign n6164 = ~pi614 & ~pi616;
  assign n6165 = n6163 & n6164;
  assign n6166 = ~pi662 & pi680;
  assign n6167 = ~pi661 & n6166;
  assign n6168 = ~pi681 & n6167;
  assign po1101 = n6165 | n6168;
  assign n6170 = ~pi332 & ~pi468;
  assign n6171 = pi835 & pi984;
  assign n6172 = ~pi252 & ~pi1001;
  assign n6173 = ~pi979 & ~n6172;
  assign n6174 = ~n6171 & n6173;
  assign n6175 = ~pi287 & n6174;
  assign n6176 = pi835 & pi950;
  assign n6177 = n6175 & n6176;
  assign n6178 = pi1092 & n6177;
  assign n6179 = ~pi824 & ~pi829;
  assign n6180 = pi824 & ~pi1091;
  assign n6181 = pi1093 & ~n2734;
  assign n6182 = ~n6180 & n6181;
  assign n6183 = ~n6179 & ~n6182;
  assign n6184 = n6178 & n6183;
  assign n6185 = ~n6170 & ~n6184;
  assign n6186 = po1101 & ~n6185;
  assign n6187 = n3096 & ~n6186;
  assign n6188 = n3090 & n6170;
  assign n6189 = po1101 & n6188;
  assign n6190 = ~n6187 & ~n6189;
  assign n6191 = ~pi587 & ~pi602;
  assign n6192 = ~pi961 & ~pi967;
  assign n6193 = ~pi969 & ~pi971;
  assign n6194 = ~pi974 & ~pi977;
  assign n6195 = n6193 & n6194;
  assign n6196 = n6191 & n6192;
  assign n6197 = n6195 & n6196;
  assign n6198 = ~n6190 & n6197;
  assign n6199 = ~n6165 & ~n6170;
  assign n6200 = ~n6168 & n6199;
  assign n6201 = n6184 & ~n6200;
  assign n6202 = n3096 & ~n6201;
  assign n6203 = ~n6197 & n6202;
  assign n6204 = pi223 & ~n6203;
  assign n6205 = ~n6198 & n6204;
  assign n6206 = po1101 & ~n6170;
  assign n6207 = n6170 & ~n6197;
  assign n6208 = ~n6206 & ~n6207;
  assign n6209 = n2796 & n6177;
  assign n6210 = pi222 & pi224;
  assign n6211 = ~n6208 & n6210;
  assign n6212 = n6209 & n6211;
  assign n6213 = n3096 & ~n6212;
  assign n6214 = ~pi223 & ~n6213;
  assign n6215 = ~pi299 & ~n6214;
  assign n6216 = ~n6205 & n6215;
  assign n6217 = ~pi907 & ~pi947;
  assign n6218 = ~pi960 & ~pi963;
  assign n6219 = ~pi970 & ~pi972;
  assign n6220 = ~pi975 & ~pi978;
  assign n6221 = n6219 & n6220;
  assign n6222 = n6218 & n6221;
  assign n6223 = n6217 & n6222;
  assign n6224 = ~n6190 & n6223;
  assign n6225 = n6202 & ~n6223;
  assign n6226 = pi215 & ~n6225;
  assign n6227 = ~n6224 & n6226;
  assign n6228 = n6170 & ~n6223;
  assign n6229 = ~n6206 & ~n6228;
  assign n6230 = pi216 & pi221;
  assign n6231 = n6209 & n6230;
  assign n6232 = ~n6229 & n6231;
  assign n6233 = n3096 & ~n6232;
  assign n6234 = ~pi215 & ~n6233;
  assign n6235 = pi299 & ~n6234;
  assign n6236 = ~n6227 & n6235;
  assign n6237 = pi39 & ~n6216;
  assign n6238 = ~n6236 & n6237;
  assign n6239 = ~n6162 & ~n6238;
  assign n6240 = ~pi38 & ~n6239;
  assign n6241 = n6119 & ~n6240;
  assign n6242 = ~pi299 & ~n3064;
  assign n6243 = pi299 & ~n2448;
  assign n6244 = ~n6242 & ~n6243;
  assign n6245 = pi146 & n6243;
  assign n6246 = pi142 & n6242;
  assign n6247 = ~n6245 & ~n6246;
  assign n6248 = ~n6244 & n6247;
  assign n6249 = ~n3382 & ~n6248;
  assign n6250 = ~pi39 & n3096;
  assign n6251 = ~pi38 & pi100;
  assign n6252 = n6250 & n6251;
  assign n6253 = ~pi41 & ~pi99;
  assign n6254 = ~pi101 & n6253;
  assign n6255 = ~pi42 & ~pi43;
  assign n6256 = ~pi52 & n6255;
  assign n6257 = ~pi113 & ~pi116;
  assign n6258 = ~pi114 & ~pi115;
  assign n6259 = n6257 & n6258;
  assign n6260 = n6256 & n6259;
  assign n6261 = n6254 & n6260;
  assign po1057 = pi44 | ~n6261;
  assign n6263 = ~pi683 & po1057;
  assign n6264 = pi129 & pi250;
  assign n6265 = pi950 & pi1092;
  assign n6266 = ~n6179 & n6265;
  assign po740 = ~pi1093 & n6266;
  assign n6268 = ~pi250 & ~po740;
  assign n6269 = ~n6264 & ~n6268;
  assign n6270 = ~n6263 & ~n6269;
  assign n6271 = n6248 & po1057;
  assign n6272 = n6270 & n6271;
  assign n6273 = ~n6249 & ~n6272;
  assign n6274 = n6252 & n6273;
  assign n6275 = ~pi87 & ~n6274;
  assign n6276 = ~n6241 & n6275;
  assign n6277 = pi87 & ~n6110;
  assign n6278 = ~pi75 & ~n6277;
  assign n6279 = ~pi54 & ~pi92;
  assign n6280 = n6278 & n6279;
  assign n6281 = ~n6276 & n6280;
  assign n6282 = ~pi74 & ~n6281;
  assign n6283 = n6116 & ~n6282;
  assign n6284 = ~pi56 & ~n6283;
  assign n6285 = ~n6112 & ~n6284;
  assign n6286 = ~pi62 & ~n6285;
  assign n6287 = n3433 & n6110;
  assign n6288 = pi62 & ~n6287;
  assign n6289 = ~pi59 & ~n6288;
  assign n6290 = ~n6286 & n6289;
  assign n6291 = ~pi57 & ~n6290;
  assign po167 = ~n6109 & ~n6291;
  assign n6293 = ~pi55 & n3294;
  assign n6294 = ~pi59 & n6293;
  assign n6295 = ~pi228 & ~n6294;
  assign n6296 = pi57 & ~n6295;
  assign n6297 = ~n6168 & ~n6170;
  assign n6298 = ~pi907 & n6170;
  assign n6299 = ~n6297 & ~n6298;
  assign n6300 = ~pi228 & ~n3269;
  assign n6301 = pi30 & pi228;
  assign n6302 = ~n3322 & ~n6301;
  assign n6303 = ~n6300 & ~n6302;
  assign n6304 = n6299 & n6303;
  assign n6305 = n6296 & n6304;
  assign n6306 = n6299 & n6301;
  assign n6307 = pi299 & ~n6306;
  assign n6308 = pi158 & pi159;
  assign n6309 = pi160 & pi197;
  assign n6310 = n6308 & n6309;
  assign n6311 = ~pi91 & ~pi314;
  assign n6312 = n2574 & ~n2575;
  assign n6313 = pi85 & n2625;
  assign n6314 = n2458 & ~n6313;
  assign n6315 = n2629 & ~n6314;
  assign n6316 = n2467 & ~n6315;
  assign n6317 = ~n2609 & ~n2638;
  assign n6318 = ~n6316 & n6317;
  assign n6319 = n2468 & n6318;
  assign n6320 = ~n2643 & ~n6319;
  assign n6321 = n2641 & ~n6320;
  assign n6322 = pi67 & n2472;
  assign n6323 = n2606 & ~n6322;
  assign n6324 = ~n6321 & n6323;
  assign n6325 = n2605 & ~n6324;
  assign n6326 = ~pi71 & ~n6325;
  assign po1049 = pi64 | ~n2476;
  assign n6328 = n2600 & ~po1049;
  assign n6329 = ~n6326 & n6328;
  assign n6330 = ~pi81 & ~n6329;
  assign n6331 = n2654 & n6328;
  assign n6332 = n6330 & ~n6331;
  assign n6333 = ~pi102 & ~n2595;
  assign n6334 = n2452 & n6333;
  assign n6335 = ~n6332 & n6334;
  assign n6336 = n2594 & ~n6335;
  assign n6337 = n2687 & ~n6336;
  assign n6338 = n2504 & ~n6337;
  assign n6339 = ~n2507 & ~n6338;
  assign n6340 = ~pi86 & ~n6339;
  assign n6341 = ~pi46 & n2483;
  assign n6342 = n2592 & n6341;
  assign n6343 = ~n6340 & n6342;
  assign n6344 = n2699 & ~n6343;
  assign n6345 = n6312 & ~n6344;
  assign n6346 = n6311 & ~n6345;
  assign n6347 = pi91 & ~n2533;
  assign n6348 = ~pi58 & ~n6347;
  assign n6349 = ~pi91 & pi314;
  assign n6350 = ~n6330 & n6334;
  assign n6351 = n2594 & ~n6350;
  assign n6352 = n2687 & ~n6351;
  assign n6353 = n2504 & ~n6352;
  assign n6354 = ~n2507 & ~n6353;
  assign n6355 = ~pi86 & ~n6354;
  assign n6356 = n6342 & ~n6355;
  assign n6357 = n2699 & ~n6356;
  assign n6358 = n6312 & ~n6357;
  assign n6359 = n6349 & ~n6358;
  assign n6360 = n6348 & ~n6359;
  assign n6361 = ~n6346 & n6360;
  assign n6362 = ~pi90 & ~n6361;
  assign n6363 = ~n2706 & ~n6362;
  assign n6364 = ~pi93 & ~n6363;
  assign n6365 = pi93 & ~n2735;
  assign n6366 = ~pi35 & ~n6365;
  assign n6367 = ~n6364 & n6366;
  assign n6368 = ~pi70 & ~n6367;
  assign n6369 = n2952 & ~n6368;
  assign n6370 = ~pi72 & ~n6369;
  assign n6371 = ~pi95 & n2725;
  assign n6372 = ~n2555 & n6371;
  assign n6373 = ~n6370 & n6372;
  assign n6374 = ~n2960 & ~n6373;
  assign n6375 = ~pi841 & n2523;
  assign n6376 = n2536 & n6375;
  assign n6377 = n2783 & n6376;
  assign n6378 = pi32 & n6377;
  assign n6379 = ~pi95 & n6378;
  assign n6380 = ~pi210 & n6379;
  assign n6381 = n6374 & ~n6380;
  assign n6382 = ~n6170 & ~n6381;
  assign n6383 = ~pi47 & n2488;
  assign n6384 = ~n2698 & ~n6343;
  assign n6385 = n6383 & ~n6384;
  assign n6386 = n6311 & ~n6385;
  assign n6387 = ~n2698 & ~n6356;
  assign n6388 = n6383 & ~n6387;
  assign n6389 = n6349 & ~n6388;
  assign n6390 = n6348 & ~n6389;
  assign n6391 = ~n6386 & n6390;
  assign n6392 = ~pi90 & ~n6391;
  assign n6393 = ~n2706 & ~n6392;
  assign n6394 = ~pi93 & ~n6393;
  assign n6395 = n6366 & ~n6394;
  assign n6396 = ~pi70 & ~n6395;
  assign n6397 = n2952 & ~n6396;
  assign n6398 = ~pi72 & ~n6397;
  assign n6399 = n6372 & ~n6398;
  assign n6400 = ~n2960 & ~n6399;
  assign n6401 = ~n6380 & n6400;
  assign n6402 = n6170 & ~n6401;
  assign n6403 = ~n6382 & ~n6402;
  assign n6404 = n6299 & ~n6403;
  assign n6405 = n6310 & ~n6404;
  assign n6406 = n6299 & ~n6381;
  assign n6407 = ~n6310 & ~n6406;
  assign n6408 = ~pi228 & ~n6407;
  assign n6409 = ~n6405 & n6408;
  assign n6410 = n6307 & ~n6409;
  assign n6411 = ~pi602 & n6170;
  assign n6412 = ~n6297 & ~n6411;
  assign n6413 = ~pi198 & n6379;
  assign n6414 = n6374 & ~n6413;
  assign n6415 = ~pi228 & ~n6414;
  assign n6416 = ~n6301 & ~n6415;
  assign n6417 = n6412 & ~n6416;
  assign n6418 = ~pi299 & ~n6417;
  assign n6419 = pi145 & pi180;
  assign n6420 = pi181 & pi182;
  assign n6421 = n6419 & n6420;
  assign n6422 = ~pi299 & n6421;
  assign n6423 = ~n6418 & ~n6422;
  assign n6424 = n6301 & n6412;
  assign n6425 = ~n6170 & ~n6414;
  assign n6426 = n6400 & ~n6413;
  assign n6427 = n6170 & ~n6426;
  assign n6428 = ~n6425 & ~n6427;
  assign n6429 = ~pi228 & n6412;
  assign n6430 = ~n6428 & n6429;
  assign n6431 = ~n6424 & ~n6430;
  assign n6432 = n6421 & ~n6431;
  assign n6433 = ~n6423 & ~n6432;
  assign n6434 = pi232 & ~n6410;
  assign n6435 = ~n6433 & n6434;
  assign n6436 = ~pi228 & n6406;
  assign n6437 = n6307 & ~n6436;
  assign n6438 = ~pi232 & ~n6437;
  assign n6439 = ~n6418 & n6438;
  assign n6440 = ~n6435 & ~n6439;
  assign n6441 = ~pi39 & ~n6440;
  assign n6442 = ~pi215 & pi221;
  assign n6443 = ~pi287 & n3096;
  assign n6444 = pi835 & n6174;
  assign n6445 = n6443 & n6444;
  assign n6446 = pi824 & pi1093;
  assign n6447 = n6265 & n6446;
  assign n6448 = n6445 & n6447;
  assign n6449 = ~pi1091 & n6448;
  assign n6450 = pi1091 & n2733;
  assign n6451 = n6447 & ~n6450;
  assign n6452 = ~n2796 & ~n6451;
  assign n6453 = pi1091 & ~n6452;
  assign n6454 = n6445 & n6453;
  assign n6455 = ~n6449 & ~n6454;
  assign n6456 = pi216 & ~n6455;
  assign n6457 = ~pi829 & ~n2733;
  assign n6458 = pi1091 & ~n6457;
  assign n6459 = n6448 & ~n6458;
  assign n6460 = ~pi216 & n6459;
  assign n6461 = ~n6456 & ~n6460;
  assign n6462 = ~pi228 & ~n6461;
  assign n6463 = ~n6301 & ~n6462;
  assign n6464 = n6442 & ~n6463;
  assign n6465 = ~n6301 & ~n6464;
  assign n6466 = n6299 & ~n6465;
  assign n6467 = pi299 & ~n6466;
  assign n6468 = pi224 & n6455;
  assign n6469 = pi222 & ~pi223;
  assign n6470 = ~pi224 & ~n6459;
  assign n6471 = n6469 & ~n6470;
  assign n6472 = ~n6468 & n6471;
  assign n6473 = ~pi228 & n6472;
  assign n6474 = ~n6301 & ~n6473;
  assign n6475 = n6412 & ~n6474;
  assign n6476 = ~pi299 & ~n6475;
  assign n6477 = pi39 & ~n6476;
  assign n6478 = ~n6467 & n6477;
  assign n6479 = ~pi38 & ~n6478;
  assign n6480 = ~n6441 & n6479;
  assign n6481 = pi299 & n6299;
  assign n6482 = ~pi299 & n6412;
  assign n6483 = ~n6481 & ~n6482;
  assign n6484 = ~pi39 & ~n6302;
  assign n6485 = ~n6483 & n6484;
  assign n6486 = n6301 & ~n6483;
  assign n6487 = pi38 & ~n6486;
  assign n6488 = ~n6485 & n6487;
  assign n6489 = ~n6480 & ~n6488;
  assign n6490 = ~pi100 & ~n6489;
  assign n6491 = ~pi142 & ~n3064;
  assign n6492 = n3096 & ~n6269;
  assign n6493 = pi683 & po1057;
  assign n6494 = n6492 & n6493;
  assign n6495 = ~n6297 & n6494;
  assign n6496 = n6491 & n6495;
  assign n6497 = pi252 & ~n6491;
  assign n6498 = pi252 & n6188;
  assign n6499 = ~n6168 & n6498;
  assign n6500 = pi252 & n3096;
  assign n6501 = n6168 & n6500;
  assign n6502 = ~n6499 & ~n6501;
  assign n6503 = n6497 & ~n6502;
  assign n6504 = ~n6496 & ~n6503;
  assign n6505 = ~pi228 & ~n6411;
  assign n6506 = ~n6504 & n6505;
  assign n6507 = ~pi299 & ~n6424;
  assign n6508 = ~n6506 & n6507;
  assign n6509 = ~n2857 & n6502;
  assign n6510 = n2857 & ~n6495;
  assign n6511 = ~pi228 & ~n6298;
  assign n6512 = ~n6510 & n6511;
  assign n6513 = ~n6509 & n6512;
  assign n6514 = n6307 & ~n6513;
  assign n6515 = n3182 & ~n6514;
  assign n6516 = ~n6508 & n6515;
  assign n6517 = ~n3182 & n6486;
  assign n6518 = pi100 & ~n6517;
  assign n6519 = ~n6516 & n6518;
  assign n6520 = ~pi87 & ~n6519;
  assign n6521 = ~n6490 & n6520;
  assign n6522 = pi87 & n6486;
  assign n6523 = ~pi75 & ~n6522;
  assign n6524 = ~n6521 & n6523;
  assign n6525 = ~n3223 & n6486;
  assign n6526 = n3242 & n6485;
  assign n6527 = ~n6525 & ~n6526;
  assign n6528 = pi75 & n6527;
  assign n6529 = ~pi92 & ~n6528;
  assign n6530 = ~n6524 & n6529;
  assign n6531 = ~pi75 & n6527;
  assign n6532 = pi75 & ~n6486;
  assign n6533 = pi92 & ~n6532;
  assign n6534 = ~n6531 & n6533;
  assign n6535 = ~pi54 & ~n6534;
  assign n6536 = ~n6530 & n6535;
  assign n6537 = n3238 & n6527;
  assign n6538 = ~n3238 & ~n6486;
  assign n6539 = ~n6537 & ~n6538;
  assign n6540 = pi54 & ~n6539;
  assign n6541 = ~pi74 & ~n6540;
  assign n6542 = ~n6536 & n6541;
  assign n6543 = ~pi54 & n6537;
  assign n6544 = ~pi54 & n3238;
  assign n6545 = ~n6486 & ~n6544;
  assign n6546 = pi74 & ~n6545;
  assign n6547 = ~n6543 & n6546;
  assign n6548 = ~pi55 & ~n6547;
  assign n6549 = ~n6542 & n6548;
  assign n6550 = pi55 & ~n6304;
  assign n6551 = n3294 & ~n6550;
  assign n6552 = ~n6549 & n6551;
  assign n6553 = ~n3294 & n6306;
  assign n6554 = ~pi59 & ~n6553;
  assign n6555 = ~n6552 & n6554;
  assign n6556 = ~pi228 & ~n6293;
  assign n6557 = n6304 & ~n6556;
  assign n6558 = pi59 & ~n6557;
  assign n6559 = ~pi57 & ~n6558;
  assign n6560 = ~n6555 & n6559;
  assign po171 = ~n6305 & ~n6560;
  assign n6562 = ~pi947 & n6170;
  assign n6563 = ~n6199 & ~n6562;
  assign n6564 = n6303 & n6563;
  assign n6565 = n6296 & n6564;
  assign n6566 = n6301 & n6563;
  assign n6567 = pi299 & ~n6566;
  assign n6568 = ~n6403 & n6563;
  assign n6569 = n6310 & ~n6568;
  assign n6570 = ~n6381 & n6563;
  assign n6571 = ~n6310 & ~n6570;
  assign n6572 = ~pi228 & ~n6571;
  assign n6573 = ~n6569 & n6572;
  assign n6574 = n6567 & ~n6573;
  assign n6575 = ~pi587 & n6170;
  assign n6576 = ~n6199 & ~n6575;
  assign n6577 = n6301 & n6576;
  assign n6578 = ~pi228 & n6576;
  assign n6579 = ~n6428 & n6578;
  assign n6580 = ~n6577 & ~n6579;
  assign n6581 = n6421 & ~n6580;
  assign n6582 = ~n6416 & n6576;
  assign n6583 = ~n6421 & n6582;
  assign n6584 = ~pi299 & ~n6583;
  assign n6585 = ~n6581 & n6584;
  assign n6586 = pi232 & ~n6574;
  assign n6587 = ~n6585 & n6586;
  assign n6588 = ~pi299 & ~n6582;
  assign n6589 = ~pi228 & n6570;
  assign n6590 = n6567 & ~n6589;
  assign n6591 = ~pi232 & ~n6590;
  assign n6592 = ~n6588 & n6591;
  assign n6593 = ~n6587 & ~n6592;
  assign n6594 = ~pi39 & ~n6593;
  assign n6595 = pi299 & n6442;
  assign n6596 = ~n6567 & ~n6595;
  assign n6597 = n6464 & n6563;
  assign n6598 = ~n6596 & ~n6597;
  assign n6599 = ~n6474 & n6576;
  assign n6600 = ~pi299 & ~n6599;
  assign n6601 = pi39 & ~n6600;
  assign n6602 = ~n6598 & n6601;
  assign n6603 = ~pi38 & ~n6602;
  assign n6604 = ~n6594 & n6603;
  assign n6605 = pi299 & ~n6563;
  assign n6606 = ~pi299 & ~n6576;
  assign n6607 = ~n6605 & ~n6606;
  assign n6608 = n6484 & n6607;
  assign n6609 = n6301 & n6607;
  assign n6610 = pi38 & ~n6609;
  assign n6611 = ~n6608 & n6610;
  assign n6612 = ~n6604 & ~n6611;
  assign n6613 = ~pi100 & ~n6612;
  assign n6614 = ~pi228 & n3064;
  assign n6615 = ~n6165 & ~n6498;
  assign n6616 = n6165 & ~n6500;
  assign n6617 = ~n6615 & ~n6616;
  assign n6618 = ~n6575 & n6617;
  assign n6619 = n6614 & ~n6618;
  assign n6620 = pi142 & ~n6617;
  assign n6621 = ~n6199 & n6494;
  assign n6622 = ~pi142 & ~n6621;
  assign n6623 = n6165 & ~n6170;
  assign n6624 = ~pi587 & ~n6623;
  assign n6625 = ~pi228 & ~n6624;
  assign n6626 = ~n6622 & n6625;
  assign n6627 = ~n6620 & n6626;
  assign n6628 = ~n6577 & ~n6614;
  assign n6629 = ~n6627 & n6628;
  assign n6630 = ~n6619 & ~n6629;
  assign n6631 = ~pi299 & ~n6630;
  assign n6632 = n2857 & ~n6562;
  assign n6633 = n6621 & n6632;
  assign n6634 = ~pi947 & ~n6623;
  assign n6635 = ~n2857 & ~n6634;
  assign n6636 = n6617 & n6635;
  assign n6637 = ~n6633 & ~n6636;
  assign n6638 = ~pi228 & ~n6637;
  assign n6639 = n6567 & ~n6638;
  assign n6640 = n3182 & ~n6639;
  assign n6641 = ~n6631 & n6640;
  assign n6642 = ~n3182 & n6609;
  assign n6643 = pi100 & ~n6642;
  assign n6644 = ~n6641 & n6643;
  assign n6645 = ~pi87 & ~n6644;
  assign n6646 = ~n6613 & n6645;
  assign n6647 = pi87 & n6609;
  assign n6648 = ~pi75 & ~n6647;
  assign n6649 = ~n6646 & n6648;
  assign n6650 = ~n3223 & n6609;
  assign n6651 = n3242 & n6608;
  assign n6652 = ~n6650 & ~n6651;
  assign n6653 = pi75 & n6652;
  assign n6654 = ~pi92 & ~n6653;
  assign n6655 = ~n6649 & n6654;
  assign n6656 = ~pi75 & n6652;
  assign n6657 = pi75 & ~n6609;
  assign n6658 = pi92 & ~n6657;
  assign n6659 = ~n6656 & n6658;
  assign n6660 = ~pi54 & ~n6659;
  assign n6661 = ~n6655 & n6660;
  assign n6662 = n3238 & n6652;
  assign n6663 = ~n3238 & ~n6609;
  assign n6664 = ~n6662 & ~n6663;
  assign n6665 = pi54 & ~n6664;
  assign n6666 = ~pi74 & ~n6665;
  assign n6667 = ~n6661 & n6666;
  assign n6668 = ~pi54 & n6662;
  assign n6669 = ~n6544 & ~n6609;
  assign n6670 = pi74 & ~n6669;
  assign n6671 = ~n6668 & n6670;
  assign n6672 = ~pi55 & ~n6671;
  assign n6673 = ~n6667 & n6672;
  assign n6674 = pi55 & ~n6564;
  assign n6675 = n3294 & ~n6674;
  assign n6676 = ~n6673 & n6675;
  assign n6677 = ~n3294 & n6566;
  assign n6678 = ~pi59 & ~n6677;
  assign n6679 = ~n6676 & n6678;
  assign n6680 = ~n6556 & n6564;
  assign n6681 = pi59 & ~n6680;
  assign n6682 = ~pi57 & ~n6681;
  assign n6683 = ~n6679 & n6682;
  assign po172 = ~n6565 & ~n6683;
  assign n6685 = pi30 & n6170;
  assign n6686 = pi228 & n6685;
  assign n6687 = pi970 & n6686;
  assign n6688 = ~pi228 & pi970;
  assign n6689 = n6188 & n6688;
  assign n6690 = n3269 & n6689;
  assign n6691 = n6294 & n6690;
  assign n6692 = ~n6687 & ~n6691;
  assign n6693 = pi57 & ~n6692;
  assign n6694 = pi299 & ~n6687;
  assign n6695 = n6170 & ~n6381;
  assign n6696 = n6688 & n6695;
  assign n6697 = n6694 & ~n6696;
  assign n6698 = pi299 & n6308;
  assign n6699 = ~n6697 & ~n6698;
  assign n6700 = n6309 & ~n6402;
  assign n6701 = ~n6309 & n6381;
  assign n6702 = ~n6700 & ~n6701;
  assign n6703 = n6170 & n6702;
  assign n6704 = n6688 & n6703;
  assign n6705 = ~n6687 & ~n6704;
  assign n6706 = n6308 & ~n6705;
  assign n6707 = ~n6699 & ~n6706;
  assign n6708 = n6170 & ~n6416;
  assign n6709 = ~n6421 & ~n6708;
  assign n6710 = ~pi228 & n6427;
  assign n6711 = ~n6414 & ~n6421;
  assign n6712 = ~n6686 & ~n6711;
  assign n6713 = ~n6710 & n6712;
  assign n6714 = ~n6709 & ~n6713;
  assign n6715 = pi967 & n6714;
  assign n6716 = ~pi299 & ~n6715;
  assign n6717 = pi232 & ~n6716;
  assign n6718 = ~n6707 & n6717;
  assign n6719 = pi967 & n6708;
  assign n6720 = ~pi299 & ~n6719;
  assign n6721 = ~pi232 & ~n6697;
  assign n6722 = ~n6720 & n6721;
  assign n6723 = ~n6718 & ~n6722;
  assign n6724 = ~pi39 & ~n6723;
  assign n6725 = pi299 & pi970;
  assign n6726 = n6442 & ~n6461;
  assign n6727 = n6170 & n6726;
  assign n6728 = ~pi228 & ~n6727;
  assign n6729 = n6725 & ~n6728;
  assign n6730 = ~pi299 & pi967;
  assign n6731 = n6170 & n6472;
  assign n6732 = ~pi228 & ~n6731;
  assign n6733 = n6730 & ~n6732;
  assign n6734 = ~n6729 & ~n6733;
  assign n6735 = pi228 & ~n6685;
  assign n6736 = pi39 & ~n6735;
  assign n6737 = ~n6734 & n6736;
  assign n6738 = ~pi38 & ~n6737;
  assign n6739 = ~n6724 & n6738;
  assign n6740 = ~pi228 & ~n6188;
  assign n6741 = ~n6735 & ~n6740;
  assign n6742 = pi967 & n6741;
  assign n6743 = ~pi299 & ~n6742;
  assign n6744 = ~n6689 & n6694;
  assign n6745 = ~pi39 & ~n6744;
  assign n6746 = ~n6743 & n6745;
  assign n6747 = ~n6725 & ~n6730;
  assign n6748 = n6686 & ~n6747;
  assign n6749 = pi39 & n6748;
  assign n6750 = pi38 & ~n6749;
  assign n6751 = ~n6746 & n6750;
  assign n6752 = ~n6739 & ~n6751;
  assign n6753 = ~pi100 & ~n6752;
  assign n6754 = ~n6491 & n6498;
  assign n6755 = n6170 & n6494;
  assign n6756 = n6491 & n6755;
  assign n6757 = ~pi228 & ~n6754;
  assign n6758 = ~n6756 & n6757;
  assign n6759 = ~n6735 & ~n6758;
  assign n6760 = pi967 & n6759;
  assign n6761 = ~pi299 & ~n6760;
  assign n6762 = ~n2857 & ~n6498;
  assign n6763 = n2857 & ~n6755;
  assign n6764 = ~pi228 & ~n6762;
  assign n6765 = ~n6763 & n6764;
  assign n6766 = pi970 & n6765;
  assign n6767 = n6694 & ~n6766;
  assign n6768 = n3182 & ~n6767;
  assign n6769 = ~n6761 & n6768;
  assign n6770 = ~n3182 & n6748;
  assign n6771 = pi100 & ~n6770;
  assign n6772 = ~n6769 & n6771;
  assign n6773 = ~pi87 & ~n6772;
  assign n6774 = ~n6753 & n6773;
  assign n6775 = pi87 & n6748;
  assign n6776 = ~pi75 & ~n6775;
  assign n6777 = ~n6774 & n6776;
  assign n6778 = ~n3223 & n6748;
  assign n6779 = n3242 & n6746;
  assign n6780 = ~n6778 & ~n6779;
  assign n6781 = pi75 & n6780;
  assign n6782 = ~pi92 & ~n6781;
  assign n6783 = ~n6777 & n6782;
  assign n6784 = ~pi75 & n6780;
  assign n6785 = pi75 & ~n6748;
  assign n6786 = pi92 & ~n6785;
  assign n6787 = ~n6784 & n6786;
  assign n6788 = ~pi54 & ~n6787;
  assign n6789 = ~n6783 & n6788;
  assign n6790 = n3238 & n6780;
  assign n6791 = ~n3238 & ~n6748;
  assign n6792 = ~n6790 & ~n6791;
  assign n6793 = pi54 & ~n6792;
  assign n6794 = ~pi74 & ~n6793;
  assign n6795 = ~n6789 & n6794;
  assign n6796 = ~pi54 & n6790;
  assign n6797 = ~n6544 & ~n6748;
  assign n6798 = pi74 & ~n6797;
  assign n6799 = ~n6796 & n6798;
  assign n6800 = ~pi55 & ~n6799;
  assign n6801 = ~n6795 & n6800;
  assign n6802 = pi55 & ~n6687;
  assign n6803 = ~n6690 & n6802;
  assign n6804 = n3294 & ~n6803;
  assign n6805 = ~n6801 & n6804;
  assign n6806 = ~n3294 & n6687;
  assign n6807 = ~pi59 & ~n6806;
  assign n6808 = ~n6805 & n6807;
  assign n6809 = n6293 & n6690;
  assign n6810 = pi59 & ~n6687;
  assign n6811 = ~n6809 & n6810;
  assign n6812 = ~pi57 & ~n6811;
  assign n6813 = ~n6808 & n6812;
  assign po173 = ~n6693 & ~n6813;
  assign n6815 = pi972 & n6686;
  assign n6816 = ~pi228 & pi972;
  assign n6817 = n6188 & n6816;
  assign n6818 = n3269 & n6817;
  assign n6819 = n6294 & n6818;
  assign n6820 = ~n6815 & ~n6819;
  assign n6821 = pi57 & ~n6820;
  assign n6822 = pi299 & ~n6815;
  assign n6823 = n6695 & n6816;
  assign n6824 = n6822 & ~n6823;
  assign n6825 = ~n6698 & ~n6824;
  assign n6826 = n6703 & n6816;
  assign n6827 = ~n6815 & ~n6826;
  assign n6828 = n6308 & ~n6827;
  assign n6829 = ~n6825 & ~n6828;
  assign n6830 = pi961 & n6714;
  assign n6831 = ~pi299 & ~n6830;
  assign n6832 = pi232 & ~n6831;
  assign n6833 = ~n6829 & n6832;
  assign n6834 = pi961 & n6708;
  assign n6835 = ~pi299 & ~n6834;
  assign n6836 = ~pi232 & ~n6824;
  assign n6837 = ~n6835 & n6836;
  assign n6838 = ~n6833 & ~n6837;
  assign n6839 = ~pi39 & ~n6838;
  assign n6840 = ~pi299 & pi961;
  assign n6841 = ~n6732 & n6840;
  assign n6842 = pi299 & pi972;
  assign n6843 = ~n6728 & n6842;
  assign n6844 = ~n6841 & ~n6843;
  assign n6845 = n6736 & ~n6844;
  assign n6846 = ~pi38 & ~n6845;
  assign n6847 = ~n6839 & n6846;
  assign n6848 = pi961 & n6741;
  assign n6849 = ~pi299 & ~n6848;
  assign n6850 = ~n6817 & n6822;
  assign n6851 = ~pi39 & ~n6850;
  assign n6852 = ~n6849 & n6851;
  assign n6853 = ~n6840 & ~n6842;
  assign n6854 = n6686 & ~n6853;
  assign n6855 = pi39 & n6854;
  assign n6856 = pi38 & ~n6855;
  assign n6857 = ~n6852 & n6856;
  assign n6858 = ~n6847 & ~n6857;
  assign n6859 = ~pi100 & ~n6858;
  assign n6860 = pi961 & n6759;
  assign n6861 = ~pi299 & ~n6860;
  assign n6862 = pi972 & n6765;
  assign n6863 = n6822 & ~n6862;
  assign n6864 = n3182 & ~n6863;
  assign n6865 = ~n6861 & n6864;
  assign n6866 = ~n3182 & n6854;
  assign n6867 = pi100 & ~n6866;
  assign n6868 = ~n6865 & n6867;
  assign n6869 = ~pi87 & ~n6868;
  assign n6870 = ~n6859 & n6869;
  assign n6871 = pi87 & n6854;
  assign n6872 = ~pi75 & ~n6871;
  assign n6873 = ~n6870 & n6872;
  assign n6874 = ~n3223 & n6854;
  assign n6875 = n3242 & n6852;
  assign n6876 = ~n6874 & ~n6875;
  assign n6877 = pi75 & n6876;
  assign n6878 = ~pi92 & ~n6877;
  assign n6879 = ~n6873 & n6878;
  assign n6880 = ~pi75 & n6876;
  assign n6881 = pi75 & ~n6854;
  assign n6882 = pi92 & ~n6881;
  assign n6883 = ~n6880 & n6882;
  assign n6884 = ~pi54 & ~n6883;
  assign n6885 = ~n6879 & n6884;
  assign n6886 = n3238 & n6876;
  assign n6887 = ~n3238 & ~n6854;
  assign n6888 = ~n6886 & ~n6887;
  assign n6889 = pi54 & ~n6888;
  assign n6890 = ~pi74 & ~n6889;
  assign n6891 = ~n6885 & n6890;
  assign n6892 = ~pi54 & n6886;
  assign n6893 = ~n6544 & ~n6854;
  assign n6894 = pi74 & ~n6893;
  assign n6895 = ~n6892 & n6894;
  assign n6896 = ~pi55 & ~n6895;
  assign n6897 = ~n6891 & n6896;
  assign n6898 = pi55 & ~n6815;
  assign n6899 = ~n6818 & n6898;
  assign n6900 = n3294 & ~n6899;
  assign n6901 = ~n6897 & n6900;
  assign n6902 = ~n3294 & n6815;
  assign n6903 = ~pi59 & ~n6902;
  assign n6904 = ~n6901 & n6903;
  assign n6905 = n6293 & n6818;
  assign n6906 = pi59 & ~n6815;
  assign n6907 = ~n6905 & n6906;
  assign n6908 = ~pi57 & ~n6907;
  assign n6909 = ~n6904 & n6908;
  assign po174 = ~n6821 & ~n6909;
  assign n6911 = pi960 & n6686;
  assign n6912 = ~pi228 & pi960;
  assign n6913 = n6188 & n6912;
  assign n6914 = n3269 & n6913;
  assign n6915 = n6294 & n6914;
  assign n6916 = ~n6911 & ~n6915;
  assign n6917 = pi57 & ~n6916;
  assign n6918 = pi299 & ~n6911;
  assign n6919 = n6695 & n6912;
  assign n6920 = n6918 & ~n6919;
  assign n6921 = ~n6698 & ~n6920;
  assign n6922 = n6703 & n6912;
  assign n6923 = ~n6911 & ~n6922;
  assign n6924 = n6308 & ~n6923;
  assign n6925 = ~n6921 & ~n6924;
  assign n6926 = pi977 & n6714;
  assign n6927 = ~pi299 & ~n6926;
  assign n6928 = pi232 & ~n6927;
  assign n6929 = ~n6925 & n6928;
  assign n6930 = pi977 & n6708;
  assign n6931 = ~pi299 & ~n6930;
  assign n6932 = ~pi232 & ~n6920;
  assign n6933 = ~n6931 & n6932;
  assign n6934 = ~n6929 & ~n6933;
  assign n6935 = ~pi39 & ~n6934;
  assign n6936 = ~pi299 & pi977;
  assign n6937 = ~n6732 & n6936;
  assign n6938 = pi299 & pi960;
  assign n6939 = ~n6728 & n6938;
  assign n6940 = ~n6937 & ~n6939;
  assign n6941 = n6736 & ~n6940;
  assign n6942 = ~pi38 & ~n6941;
  assign n6943 = ~n6935 & n6942;
  assign n6944 = pi977 & n6741;
  assign n6945 = ~pi299 & ~n6944;
  assign n6946 = ~n6913 & n6918;
  assign n6947 = ~pi39 & ~n6946;
  assign n6948 = ~n6945 & n6947;
  assign n6949 = ~n6936 & ~n6938;
  assign n6950 = n6686 & ~n6949;
  assign n6951 = pi39 & n6950;
  assign n6952 = pi38 & ~n6951;
  assign n6953 = ~n6948 & n6952;
  assign n6954 = ~n6943 & ~n6953;
  assign n6955 = ~pi100 & ~n6954;
  assign n6956 = pi977 & n6759;
  assign n6957 = ~pi299 & ~n6956;
  assign n6958 = pi960 & n6765;
  assign n6959 = n6918 & ~n6958;
  assign n6960 = n3182 & ~n6959;
  assign n6961 = ~n6957 & n6960;
  assign n6962 = ~n3182 & n6950;
  assign n6963 = pi100 & ~n6962;
  assign n6964 = ~n6961 & n6963;
  assign n6965 = ~pi87 & ~n6964;
  assign n6966 = ~n6955 & n6965;
  assign n6967 = pi87 & n6950;
  assign n6968 = ~pi75 & ~n6967;
  assign n6969 = ~n6966 & n6968;
  assign n6970 = ~n3223 & n6950;
  assign n6971 = n3242 & n6948;
  assign n6972 = ~n6970 & ~n6971;
  assign n6973 = pi75 & n6972;
  assign n6974 = ~pi92 & ~n6973;
  assign n6975 = ~n6969 & n6974;
  assign n6976 = ~pi75 & n6972;
  assign n6977 = pi75 & ~n6950;
  assign n6978 = pi92 & ~n6977;
  assign n6979 = ~n6976 & n6978;
  assign n6980 = ~pi54 & ~n6979;
  assign n6981 = ~n6975 & n6980;
  assign n6982 = n3238 & n6972;
  assign n6983 = ~n3238 & ~n6950;
  assign n6984 = ~n6982 & ~n6983;
  assign n6985 = pi54 & ~n6984;
  assign n6986 = ~pi74 & ~n6985;
  assign n6987 = ~n6981 & n6986;
  assign n6988 = ~pi54 & n6982;
  assign n6989 = ~n6544 & ~n6950;
  assign n6990 = pi74 & ~n6989;
  assign n6991 = ~n6988 & n6990;
  assign n6992 = ~pi55 & ~n6991;
  assign n6993 = ~n6987 & n6992;
  assign n6994 = pi55 & ~n6911;
  assign n6995 = ~n6914 & n6994;
  assign n6996 = n3294 & ~n6995;
  assign n6997 = ~n6993 & n6996;
  assign n6998 = ~n3294 & n6911;
  assign n6999 = ~pi59 & ~n6998;
  assign n7000 = ~n6997 & n6999;
  assign n7001 = n6293 & n6914;
  assign n7002 = pi59 & ~n6911;
  assign n7003 = ~n7001 & n7002;
  assign n7004 = ~pi57 & ~n7003;
  assign n7005 = ~n7000 & n7004;
  assign po175 = ~n6917 & ~n7005;
  assign n7007 = pi963 & n6686;
  assign n7008 = ~pi228 & pi963;
  assign n7009 = n6188 & n7008;
  assign n7010 = n3269 & n7009;
  assign n7011 = n6294 & n7010;
  assign n7012 = ~n7007 & ~n7011;
  assign n7013 = pi57 & ~n7012;
  assign n7014 = pi299 & ~n7007;
  assign n7015 = n6695 & n7008;
  assign n7016 = n7014 & ~n7015;
  assign n7017 = ~n6698 & ~n7016;
  assign n7018 = n6703 & n7008;
  assign n7019 = ~n7007 & ~n7018;
  assign n7020 = n6308 & ~n7019;
  assign n7021 = ~n7017 & ~n7020;
  assign n7022 = pi969 & n6714;
  assign n7023 = ~pi299 & ~n7022;
  assign n7024 = pi232 & ~n7023;
  assign n7025 = ~n7021 & n7024;
  assign n7026 = pi969 & n6708;
  assign n7027 = ~pi299 & ~n7026;
  assign n7028 = ~pi232 & ~n7016;
  assign n7029 = ~n7027 & n7028;
  assign n7030 = ~n7025 & ~n7029;
  assign n7031 = ~pi39 & ~n7030;
  assign n7032 = ~pi299 & pi969;
  assign n7033 = ~n6732 & n7032;
  assign n7034 = pi299 & pi963;
  assign n7035 = ~n6728 & n7034;
  assign n7036 = ~n7033 & ~n7035;
  assign n7037 = n6736 & ~n7036;
  assign n7038 = ~pi38 & ~n7037;
  assign n7039 = ~n7031 & n7038;
  assign n7040 = pi969 & n6741;
  assign n7041 = ~pi299 & ~n7040;
  assign n7042 = ~n7009 & n7014;
  assign n7043 = ~pi39 & ~n7042;
  assign n7044 = ~n7041 & n7043;
  assign n7045 = ~n7032 & ~n7034;
  assign n7046 = n6686 & ~n7045;
  assign n7047 = pi39 & n7046;
  assign n7048 = pi38 & ~n7047;
  assign n7049 = ~n7044 & n7048;
  assign n7050 = ~n7039 & ~n7049;
  assign n7051 = ~pi100 & ~n7050;
  assign n7052 = pi969 & n6759;
  assign n7053 = ~pi299 & ~n7052;
  assign n7054 = pi963 & n6765;
  assign n7055 = n7014 & ~n7054;
  assign n7056 = n3182 & ~n7055;
  assign n7057 = ~n7053 & n7056;
  assign n7058 = ~n3182 & n7046;
  assign n7059 = pi100 & ~n7058;
  assign n7060 = ~n7057 & n7059;
  assign n7061 = ~pi87 & ~n7060;
  assign n7062 = ~n7051 & n7061;
  assign n7063 = pi87 & n7046;
  assign n7064 = ~pi75 & ~n7063;
  assign n7065 = ~n7062 & n7064;
  assign n7066 = ~n3223 & n7046;
  assign n7067 = n3242 & n7044;
  assign n7068 = ~n7066 & ~n7067;
  assign n7069 = pi75 & n7068;
  assign n7070 = ~pi92 & ~n7069;
  assign n7071 = ~n7065 & n7070;
  assign n7072 = ~pi75 & n7068;
  assign n7073 = pi75 & ~n7046;
  assign n7074 = pi92 & ~n7073;
  assign n7075 = ~n7072 & n7074;
  assign n7076 = ~pi54 & ~n7075;
  assign n7077 = ~n7071 & n7076;
  assign n7078 = n3238 & n7068;
  assign n7079 = ~n3238 & ~n7046;
  assign n7080 = ~n7078 & ~n7079;
  assign n7081 = pi54 & ~n7080;
  assign n7082 = ~pi74 & ~n7081;
  assign n7083 = ~n7077 & n7082;
  assign n7084 = ~pi54 & n7078;
  assign n7085 = ~n6544 & ~n7046;
  assign n7086 = pi74 & ~n7085;
  assign n7087 = ~n7084 & n7086;
  assign n7088 = ~pi55 & ~n7087;
  assign n7089 = ~n7083 & n7088;
  assign n7090 = pi55 & ~n7007;
  assign n7091 = ~n7010 & n7090;
  assign n7092 = n3294 & ~n7091;
  assign n7093 = ~n7089 & n7092;
  assign n7094 = ~n3294 & n7007;
  assign n7095 = ~pi59 & ~n7094;
  assign n7096 = ~n7093 & n7095;
  assign n7097 = n6293 & n7010;
  assign n7098 = pi59 & ~n7007;
  assign n7099 = ~n7097 & n7098;
  assign n7100 = ~pi57 & ~n7099;
  assign n7101 = ~n7096 & n7100;
  assign po176 = ~n7013 & ~n7101;
  assign n7103 = pi975 & n6686;
  assign n7104 = ~pi228 & pi975;
  assign n7105 = n6188 & n7104;
  assign n7106 = n3269 & n7105;
  assign n7107 = n6294 & n7106;
  assign n7108 = ~n7103 & ~n7107;
  assign n7109 = pi57 & ~n7108;
  assign n7110 = pi299 & ~n7103;
  assign n7111 = n6695 & n7104;
  assign n7112 = n7110 & ~n7111;
  assign n7113 = ~n6698 & ~n7112;
  assign n7114 = n6703 & n7104;
  assign n7115 = ~n7103 & ~n7114;
  assign n7116 = n6308 & ~n7115;
  assign n7117 = ~n7113 & ~n7116;
  assign n7118 = pi971 & n6714;
  assign n7119 = ~pi299 & ~n7118;
  assign n7120 = pi232 & ~n7119;
  assign n7121 = ~n7117 & n7120;
  assign n7122 = pi971 & n6708;
  assign n7123 = ~pi299 & ~n7122;
  assign n7124 = ~pi232 & ~n7112;
  assign n7125 = ~n7123 & n7124;
  assign n7126 = ~n7121 & ~n7125;
  assign n7127 = ~pi39 & ~n7126;
  assign n7128 = ~pi299 & pi971;
  assign n7129 = ~n6732 & n7128;
  assign n7130 = pi299 & pi975;
  assign n7131 = ~n6728 & n7130;
  assign n7132 = ~n7129 & ~n7131;
  assign n7133 = n6736 & ~n7132;
  assign n7134 = ~pi38 & ~n7133;
  assign n7135 = ~n7127 & n7134;
  assign n7136 = pi971 & n6741;
  assign n7137 = ~pi299 & ~n7136;
  assign n7138 = ~n7105 & n7110;
  assign n7139 = ~pi39 & ~n7138;
  assign n7140 = ~n7137 & n7139;
  assign n7141 = ~n7128 & ~n7130;
  assign n7142 = n6686 & ~n7141;
  assign n7143 = pi39 & n7142;
  assign n7144 = pi38 & ~n7143;
  assign n7145 = ~n7140 & n7144;
  assign n7146 = ~n7135 & ~n7145;
  assign n7147 = ~pi100 & ~n7146;
  assign n7148 = pi971 & n6759;
  assign n7149 = ~pi299 & ~n7148;
  assign n7150 = pi975 & n6765;
  assign n7151 = n7110 & ~n7150;
  assign n7152 = n3182 & ~n7151;
  assign n7153 = ~n7149 & n7152;
  assign n7154 = ~n3182 & n7142;
  assign n7155 = pi100 & ~n7154;
  assign n7156 = ~n7153 & n7155;
  assign n7157 = ~pi87 & ~n7156;
  assign n7158 = ~n7147 & n7157;
  assign n7159 = pi87 & n7142;
  assign n7160 = ~pi75 & ~n7159;
  assign n7161 = ~n7158 & n7160;
  assign n7162 = ~n3223 & n7142;
  assign n7163 = n3242 & n7140;
  assign n7164 = ~n7162 & ~n7163;
  assign n7165 = pi75 & n7164;
  assign n7166 = ~pi92 & ~n7165;
  assign n7167 = ~n7161 & n7166;
  assign n7168 = ~pi75 & n7164;
  assign n7169 = pi75 & ~n7142;
  assign n7170 = pi92 & ~n7169;
  assign n7171 = ~n7168 & n7170;
  assign n7172 = ~pi54 & ~n7171;
  assign n7173 = ~n7167 & n7172;
  assign n7174 = n3238 & n7164;
  assign n7175 = ~n3238 & ~n7142;
  assign n7176 = ~n7174 & ~n7175;
  assign n7177 = pi54 & ~n7176;
  assign n7178 = ~pi74 & ~n7177;
  assign n7179 = ~n7173 & n7178;
  assign n7180 = ~pi54 & n7174;
  assign n7181 = ~n6544 & ~n7142;
  assign n7182 = pi74 & ~n7181;
  assign n7183 = ~n7180 & n7182;
  assign n7184 = ~pi55 & ~n7183;
  assign n7185 = ~n7179 & n7184;
  assign n7186 = pi55 & ~n7103;
  assign n7187 = ~n7106 & n7186;
  assign n7188 = n3294 & ~n7187;
  assign n7189 = ~n7185 & n7188;
  assign n7190 = ~n3294 & n7103;
  assign n7191 = ~pi59 & ~n7190;
  assign n7192 = ~n7189 & n7191;
  assign n7193 = n6293 & n7106;
  assign n7194 = pi59 & ~n7103;
  assign n7195 = ~n7193 & n7194;
  assign n7196 = ~pi57 & ~n7195;
  assign n7197 = ~n7192 & n7196;
  assign po177 = ~n7109 & ~n7197;
  assign n7199 = pi978 & n6686;
  assign n7200 = ~pi228 & pi978;
  assign n7201 = n3269 & n7200;
  assign n7202 = n6188 & n7201;
  assign n7203 = n6294 & n7202;
  assign n7204 = ~n7199 & ~n7203;
  assign n7205 = pi57 & ~n7204;
  assign n7206 = ~pi299 & pi974;
  assign n7207 = pi299 & pi978;
  assign n7208 = ~n7206 & ~n7207;
  assign n7209 = n6741 & ~n7208;
  assign n7210 = ~pi39 & n7209;
  assign n7211 = n6686 & ~n7208;
  assign n7212 = pi39 & n7211;
  assign n7213 = pi38 & ~n7212;
  assign n7214 = ~n7210 & n7213;
  assign n7215 = pi299 & ~n7199;
  assign n7216 = n6695 & n7200;
  assign n7217 = n7215 & ~n7216;
  assign n7218 = ~n6698 & ~n7217;
  assign n7219 = n6703 & n7200;
  assign n7220 = ~n7199 & ~n7219;
  assign n7221 = n6308 & ~n7220;
  assign n7222 = ~n7218 & ~n7221;
  assign n7223 = pi974 & n6714;
  assign n7224 = ~pi299 & ~n7223;
  assign n7225 = pi232 & ~n7224;
  assign n7226 = ~n7222 & n7225;
  assign n7227 = pi974 & n6708;
  assign n7228 = ~pi299 & ~n7227;
  assign n7229 = ~pi232 & ~n7217;
  assign n7230 = ~n7228 & n7229;
  assign n7231 = ~n7226 & ~n7230;
  assign n7232 = ~pi39 & ~n7231;
  assign n7233 = ~n6732 & n7206;
  assign n7234 = ~n6728 & n7207;
  assign n7235 = ~n7233 & ~n7234;
  assign n7236 = n6736 & ~n7235;
  assign n7237 = ~pi38 & ~n7236;
  assign n7238 = ~n7232 & n7237;
  assign n7239 = ~n7214 & ~n7238;
  assign n7240 = ~pi100 & ~n7239;
  assign n7241 = pi974 & n6759;
  assign n7242 = ~pi299 & ~n7241;
  assign n7243 = pi978 & n6765;
  assign n7244 = n7215 & ~n7243;
  assign n7245 = n3182 & ~n7244;
  assign n7246 = ~n7242 & n7245;
  assign n7247 = ~n3182 & n7211;
  assign n7248 = pi100 & ~n7247;
  assign n7249 = ~n7246 & n7248;
  assign n7250 = ~pi87 & ~n7249;
  assign n7251 = ~n7240 & n7250;
  assign n7252 = pi87 & n7211;
  assign n7253 = ~pi75 & ~n7252;
  assign n7254 = ~n7251 & n7253;
  assign n7255 = ~pi228 & ~n3223;
  assign n7256 = n7209 & ~n7255;
  assign n7257 = pi75 & ~n7256;
  assign n7258 = ~pi92 & ~n7257;
  assign n7259 = ~n7254 & n7258;
  assign n7260 = ~pi75 & ~n7256;
  assign n7261 = pi75 & ~n7211;
  assign n7262 = pi92 & ~n7261;
  assign n7263 = ~n7260 & n7262;
  assign n7264 = ~pi54 & ~n7263;
  assign n7265 = ~n7259 & n7264;
  assign n7266 = n3238 & ~n7256;
  assign n7267 = ~n3238 & ~n7211;
  assign n7268 = ~n7266 & ~n7267;
  assign n7269 = pi54 & ~n7268;
  assign n7270 = ~pi74 & ~n7269;
  assign n7271 = ~n7265 & n7270;
  assign n7272 = ~pi54 & n7266;
  assign n7273 = ~n6544 & ~n7211;
  assign n7274 = pi74 & ~n7273;
  assign n7275 = ~n7272 & n7274;
  assign n7276 = ~pi55 & ~n7275;
  assign n7277 = ~n7271 & n7276;
  assign n7278 = pi55 & ~n7199;
  assign n7279 = ~n7202 & n7278;
  assign n7280 = n3294 & ~n7279;
  assign n7281 = ~n7277 & n7280;
  assign n7282 = ~n3294 & n7199;
  assign n7283 = ~pi59 & ~n7282;
  assign n7284 = ~n7281 & n7283;
  assign n7285 = n6293 & n7202;
  assign n7286 = pi59 & ~n7199;
  assign n7287 = ~n7285 & n7286;
  assign n7288 = ~pi57 & ~n7287;
  assign n7289 = ~n7284 & n7288;
  assign po178 = ~n7205 & ~n7289;
  assign n7291 = n3242 & n6250;
  assign n7292 = pi75 & ~n7291;
  assign n7293 = n3207 & n3231;
  assign n7294 = n6250 & n7293;
  assign n7295 = pi92 & ~n7294;
  assign n7296 = ~n7292 & ~n7295;
  assign n7297 = pi299 & ~n6229;
  assign n7298 = n6726 & n7297;
  assign n7299 = ~pi299 & ~n6208;
  assign n7300 = n6472 & n7299;
  assign n7301 = pi39 & ~n7300;
  assign n7302 = ~n7298 & n7301;
  assign n7303 = n6421 & n6427;
  assign n7304 = ~pi299 & ~n6425;
  assign n7305 = ~n6711 & n7304;
  assign n7306 = ~n7303 & n7305;
  assign n7307 = ~n6382 & n6698;
  assign n7308 = ~n6702 & n7307;
  assign n7309 = pi299 & n6381;
  assign n7310 = ~n6308 & n7309;
  assign n7311 = pi232 & ~n7310;
  assign n7312 = ~n7306 & n7311;
  assign n7313 = ~n7308 & n7312;
  assign n7314 = ~pi299 & n6414;
  assign n7315 = ~pi232 & ~n7309;
  assign n7316 = ~n7314 & n7315;
  assign n7317 = ~pi39 & ~n7316;
  assign n7318 = ~n7313 & n7317;
  assign n7319 = ~n7302 & ~n7318;
  assign n7320 = ~pi38 & ~n7319;
  assign n7321 = ~n6118 & ~n7320;
  assign n7322 = ~pi100 & ~n7321;
  assign n7323 = ~pi38 & n6250;
  assign n7324 = pi100 & ~n7323;
  assign n7325 = n6275 & ~n7324;
  assign n7326 = ~n7322 & n7325;
  assign n7327 = n3238 & ~n7326;
  assign n7328 = n7296 & ~n7327;
  assign n7329 = ~pi54 & ~n7328;
  assign n7330 = ~pi92 & n7294;
  assign n7331 = pi54 & ~n7330;
  assign n7332 = ~n7329 & ~n7331;
  assign n7333 = ~pi74 & ~n7332;
  assign n7334 = ~n6115 & ~n7333;
  assign n7335 = ~pi55 & ~n7334;
  assign n7336 = n3279 & n6110;
  assign n7337 = pi55 & ~n7336;
  assign n7338 = ~pi56 & ~n7337;
  assign n7339 = ~pi62 & n7338;
  assign n7340 = ~n7335 & n7339;
  assign n7341 = n3432 & ~n7340;
  assign po195 = n6108 & ~n7341;
  assign n7343 = ~pi954 & ~po195;
  assign n7344 = pi24 & pi954;
  assign po182 = ~n7343 & ~n7344;
  assign n7346 = n3277 & n3322;
  assign n7347 = n3433 & n7346;
  assign n7348 = ~n3127 & ~n7347;
  assign n7349 = pi62 & ~n7348;
  assign n7350 = ~pi100 & n4678;
  assign n7351 = n3096 & ~n6497;
  assign n7352 = ~pi299 & ~n7351;
  assign n7353 = pi299 & ~n3391;
  assign n7354 = ~n7352 & ~n7353;
  assign n7355 = pi100 & n3322;
  assign n7356 = n7354 & n7355;
  assign n7357 = ~pi39 & ~n7356;
  assign n7358 = ~n7350 & n7357;
  assign n7359 = ~pi100 & n3322;
  assign n7360 = pi39 & ~n7359;
  assign n7361 = ~pi38 & ~n7360;
  assign n7362 = ~n7358 & n7361;
  assign n7363 = ~n3127 & ~n7362;
  assign n7364 = ~pi87 & ~n7363;
  assign n7365 = ~n3127 & ~n7346;
  assign n7366 = pi87 & ~n7365;
  assign n7367 = ~pi75 & ~n7366;
  assign n7368 = ~n7364 & n7367;
  assign n7369 = pi75 & ~n3127;
  assign n7370 = ~pi92 & ~n7369;
  assign n7371 = ~n7368 & n7370;
  assign n7372 = n3322 & n3409;
  assign n7373 = ~n3127 & ~n7372;
  assign n7374 = pi92 & ~n7373;
  assign n7375 = n3266 & ~n7374;
  assign n7376 = ~n7371 & n7375;
  assign n7377 = ~n3127 & ~n3266;
  assign n7378 = ~pi55 & ~n7377;
  assign n7379 = ~n7376 & n7378;
  assign n7380 = n3277 & n6113;
  assign n7381 = n3322 & n7380;
  assign n7382 = ~pi74 & n7381;
  assign n7383 = ~n3127 & ~n7382;
  assign n7384 = pi55 & ~n7383;
  assign n7385 = ~pi56 & ~n7384;
  assign n7386 = ~n7379 & n7385;
  assign n7387 = n3281 & n3322;
  assign n7388 = pi56 & ~n3127;
  assign n7389 = ~n7387 & n7388;
  assign n7390 = ~pi62 & ~n7389;
  assign n7391 = ~n7386 & n7390;
  assign n7392 = ~n7349 & ~n7391;
  assign n7393 = n3432 & ~n7392;
  assign n7394 = n3127 & ~n3432;
  assign po183 = n7393 | n7394;
  assign n7396 = pi119 & pi1056;
  assign n7397 = ~pi228 & pi252;
  assign n7398 = ~pi119 & ~n7397;
  assign n7399 = ~pi468 & ~n7398;
  assign po184 = n7396 | ~n7399;
  assign n7401 = pi119 & pi1077;
  assign po185 = ~n7399 | n7401;
  assign n7403 = pi119 & pi1073;
  assign po186 = ~n7399 | n7403;
  assign n7405 = pi119 & pi1041;
  assign po187 = ~n7399 | n7405;
  assign n7407 = pi360 & ~pi462;
  assign n7408 = ~pi360 & pi462;
  assign n7409 = ~n7407 & ~n7408;
  assign n7410 = pi352 & ~pi353;
  assign n7411 = ~pi352 & pi353;
  assign n7412 = ~n7410 & ~n7411;
  assign n7413 = n7409 & n7412;
  assign n7414 = ~n7409 & ~n7412;
  assign n7415 = ~n7413 & ~n7414;
  assign n7416 = pi354 & ~n7415;
  assign n7417 = ~pi354 & n7415;
  assign n7418 = ~n7416 & ~n7417;
  assign n7419 = pi345 & ~pi346;
  assign n7420 = ~pi345 & pi346;
  assign n7421 = ~n7419 & ~n7420;
  assign n7422 = pi323 & ~n7421;
  assign n7423 = ~pi323 & n7421;
  assign n7424 = ~n7422 & ~n7423;
  assign n7425 = pi358 & ~pi450;
  assign n7426 = ~pi358 & pi450;
  assign n7427 = ~n7425 & ~n7426;
  assign n7428 = n7424 & ~n7427;
  assign n7429 = ~n7424 & n7427;
  assign n7430 = ~n7428 & ~n7429;
  assign n7431 = ~pi327 & ~pi362;
  assign n7432 = pi327 & pi362;
  assign n7433 = ~n7431 & ~n7432;
  assign n7434 = pi343 & ~pi344;
  assign n7435 = ~pi343 & pi344;
  assign n7436 = ~n7434 & ~n7435;
  assign n7437 = n7433 & ~n7436;
  assign n7438 = ~n7433 & n7436;
  assign n7439 = ~n7437 & ~n7438;
  assign n7440 = n7430 & n7439;
  assign n7441 = ~n7430 & ~n7439;
  assign n7442 = pi1197 & ~n7440;
  assign n7443 = ~n7441 & n7442;
  assign n7444 = ~pi74 & n6279;
  assign n7445 = n2535 & ~n6139;
  assign n7446 = ~pi841 & n2492;
  assign n7447 = pi90 & n7446;
  assign n7448 = ~pi93 & ~n7447;
  assign n7449 = n7445 & ~n7448;
  assign n7450 = ~pi51 & ~n7449;
  assign n7451 = ~pi50 & ~pi77;
  assign n7452 = ~pi94 & n7451;
  assign n7453 = n2576 & n7452;
  assign n7454 = ~pi88 & pi98;
  assign n7455 = n2482 & n7454;
  assign n7456 = n7453 & n7455;
  assign n7457 = ~pi97 & ~n7456;
  assign n7458 = n2514 & ~n7457;
  assign n7459 = ~pi35 & n2493;
  assign n7460 = ~pi70 & n7459;
  assign n7461 = n7458 & n7460;
  assign n7462 = n7450 & ~n7461;
  assign n7463 = ~n2558 & ~n7462;
  assign n7464 = ~pi96 & n3094;
  assign n7465 = n7463 & n7464;
  assign n7466 = n6266 & n7465;
  assign n7467 = ~pi96 & ~n7463;
  assign n7468 = pi96 & ~n6376;
  assign n7469 = n3094 & ~n7468;
  assign n7470 = ~pi122 & pi829;
  assign n7471 = n6265 & n7470;
  assign n7472 = n7469 & n7471;
  assign n7473 = ~n7467 & n7472;
  assign n7474 = ~n7466 & ~n7473;
  assign n7475 = ~pi1093 & ~n7474;
  assign n7476 = ~pi87 & ~n7475;
  assign n7477 = n3096 & po740;
  assign n7478 = pi87 & ~n7477;
  assign n7479 = ~pi75 & n3277;
  assign n7480 = ~n7478 & n7479;
  assign n7481 = ~n7476 & n7480;
  assign n7482 = ~pi567 & ~n7481;
  assign n7483 = n7444 & ~n7482;
  assign n7484 = pi232 & n6170;
  assign n7485 = n6244 & n7484;
  assign n7486 = n3223 & ~n7485;
  assign n7487 = ~pi24 & n6500;
  assign n7488 = ~n2733 & po1057;
  assign n7489 = pi1091 & n7488;
  assign n7490 = n7471 & n7489;
  assign n7491 = n7487 & n7490;
  assign n7492 = pi1093 & n7491;
  assign n7493 = n7486 & n7492;
  assign n7494 = pi75 & ~n7493;
  assign n7495 = pi1093 & ~n2733;
  assign n7496 = pi824 & n6265;
  assign n7497 = ~n2558 & n7464;
  assign n7498 = ~n7450 & n7497;
  assign n7499 = n7496 & n7498;
  assign n7500 = ~pi829 & n7499;
  assign n7501 = ~pi24 & n2565;
  assign n7502 = ~pi46 & pi97;
  assign n7503 = ~pi108 & n7502;
  assign n7504 = n6383 & n7503;
  assign n7505 = n2581 & n7504;
  assign n7506 = ~pi91 & n7505;
  assign n7507 = ~n7501 & ~n7506;
  assign n7508 = n2518 & n7445;
  assign n7509 = ~n7507 & n7508;
  assign n7510 = n7450 & ~n7509;
  assign n7511 = ~n2558 & ~n7510;
  assign n7512 = ~pi96 & ~n7511;
  assign n7513 = pi829 & n6265;
  assign n7514 = n7469 & n7513;
  assign n7515 = ~n7512 & n7514;
  assign n7516 = ~n7500 & ~n7515;
  assign n7517 = ~pi122 & ~n7516;
  assign n7518 = pi122 & n6266;
  assign n7519 = n7498 & n7518;
  assign n7520 = ~n7517 & ~n7519;
  assign n7521 = n7495 & ~n7520;
  assign n7522 = pi1091 & ~n7521;
  assign n7523 = ~n7475 & n7522;
  assign n7524 = ~pi1091 & ~n7475;
  assign n7525 = ~n7523 & ~n7524;
  assign n7526 = ~pi39 & ~n7525;
  assign n7527 = ~n2733 & n2754;
  assign n7528 = n6445 & n7527;
  assign n7529 = n2755 & n7528;
  assign n7530 = pi1091 & n7529;
  assign n7531 = ~n6229 & n7530;
  assign n7532 = ~pi216 & n6595;
  assign n7533 = n7531 & n7532;
  assign n7534 = ~n6208 & n7530;
  assign n7535 = ~pi299 & n6469;
  assign n7536 = ~pi224 & n7535;
  assign n7537 = n7534 & n7536;
  assign n7538 = pi39 & ~n7533;
  assign n7539 = ~n7537 & n7538;
  assign n7540 = ~pi38 & ~n7539;
  assign n7541 = ~n7526 & n7540;
  assign n7542 = ~pi100 & ~n7541;
  assign n7543 = n6447 & n7498;
  assign n7544 = n7540 & n7543;
  assign n7545 = ~n7522 & n7544;
  assign n7546 = n7542 & ~n7545;
  assign n7547 = pi1093 & n7471;
  assign n7548 = n7488 & n7547;
  assign n7549 = n3096 & n7548;
  assign n7550 = pi1091 & n7549;
  assign n7551 = pi228 & n7550;
  assign n7552 = n3182 & ~n7485;
  assign n7553 = n7551 & n7552;
  assign n7554 = pi100 & ~n7553;
  assign n7555 = ~n7546 & ~n7554;
  assign n7556 = ~pi87 & ~n7555;
  assign n7557 = n3096 & n7496;
  assign n7558 = ~pi1091 & pi1093;
  assign n7559 = ~n7557 & n7558;
  assign n7560 = pi1093 & n2733;
  assign n7561 = n6266 & ~n7560;
  assign n7562 = n3096 & n7561;
  assign n7563 = ~n7558 & ~n7562;
  assign n7564 = n3208 & ~n7563;
  assign n7565 = ~n7559 & n7564;
  assign n7566 = pi87 & ~n7565;
  assign n7567 = ~n7556 & ~n7566;
  assign n7568 = ~pi75 & ~n7567;
  assign n7569 = ~n7494 & ~n7568;
  assign n7570 = pi567 & ~n7569;
  assign n7571 = n7483 & ~n7570;
  assign n7572 = ~pi350 & ~pi592;
  assign n7573 = ~n7571 & ~n7572;
  assign n7574 = pi321 & ~pi347;
  assign n7575 = ~pi321 & pi347;
  assign n7576 = ~n7574 & ~n7575;
  assign n7577 = pi316 & ~pi349;
  assign n7578 = ~pi316 & pi349;
  assign n7579 = ~n7577 & ~n7578;
  assign n7580 = pi348 & n7579;
  assign n7581 = ~pi348 & ~n7579;
  assign n7582 = ~n7580 & ~n7581;
  assign n7583 = pi315 & ~pi359;
  assign n7584 = ~pi315 & pi359;
  assign n7585 = ~n7583 & ~n7584;
  assign n7586 = pi322 & n7585;
  assign n7587 = ~pi322 & ~n7585;
  assign n7588 = ~n7586 & ~n7587;
  assign n7589 = n7582 & ~n7588;
  assign n7590 = ~n7582 & n7588;
  assign n7591 = ~n7589 & ~n7590;
  assign n7592 = n7576 & n7591;
  assign n7593 = ~n7576 & ~n7591;
  assign n7594 = ~n7592 & ~n7593;
  assign n7595 = ~pi87 & ~n7554;
  assign n7596 = ~n7542 & n7595;
  assign n7597 = pi1091 & ~n7562;
  assign n7598 = ~pi1091 & ~n7477;
  assign n7599 = pi87 & ~pi100;
  assign n7600 = n3182 & n7599;
  assign n7601 = ~n7597 & n7600;
  assign n7602 = ~n7598 & n7601;
  assign n7603 = ~pi75 & ~n7602;
  assign n7604 = ~n7596 & n7603;
  assign n7605 = ~n7494 & ~n7604;
  assign n7606 = pi567 & ~n7605;
  assign n7607 = n7483 & ~n7606;
  assign n7608 = n7572 & ~n7607;
  assign n7609 = n7594 & ~n7608;
  assign n7610 = ~n7573 & n7609;
  assign n7611 = pi350 & ~pi592;
  assign n7612 = ~n7571 & ~n7611;
  assign n7613 = ~n7607 & n7611;
  assign n7614 = ~n7594 & ~n7613;
  assign n7615 = ~n7612 & n7614;
  assign n7616 = pi452 & ~pi455;
  assign n7617 = ~pi452 & pi455;
  assign n7618 = ~n7616 & ~n7617;
  assign n7619 = pi355 & n7618;
  assign n7620 = ~pi355 & ~n7618;
  assign n7621 = ~n7619 & ~n7620;
  assign n7622 = pi320 & ~pi460;
  assign n7623 = ~pi320 & pi460;
  assign n7624 = ~n7622 & ~n7623;
  assign n7625 = pi342 & ~n7624;
  assign n7626 = ~pi342 & n7624;
  assign n7627 = ~n7625 & ~n7626;
  assign n7628 = pi361 & ~pi441;
  assign n7629 = ~pi361 & pi441;
  assign n7630 = ~n7628 & ~n7629;
  assign n7631 = n7627 & n7630;
  assign n7632 = ~n7627 & ~n7630;
  assign n7633 = ~n7631 & ~n7632;
  assign n7634 = pi458 & n7633;
  assign n7635 = ~pi458 & ~n7633;
  assign n7636 = ~n7634 & ~n7635;
  assign n7637 = n7621 & n7636;
  assign n7638 = ~n7621 & ~n7636;
  assign n7639 = ~n7637 & ~n7638;
  assign n7640 = pi1196 & n7639;
  assign n7641 = ~n7610 & ~n7640;
  assign n7642 = ~n7615 & n7641;
  assign n7643 = ~pi592 & ~n7607;
  assign n7644 = pi592 & ~n7571;
  assign n7645 = ~n7643 & ~n7644;
  assign n7646 = n7640 & ~n7645;
  assign n7647 = pi1198 & ~n7646;
  assign n7648 = ~n7642 & n7647;
  assign n7649 = ~pi455 & ~n7645;
  assign n7650 = pi455 & ~n7571;
  assign n7651 = ~n7649 & ~n7650;
  assign n7652 = ~pi452 & ~n7651;
  assign n7653 = pi455 & ~n7645;
  assign n7654 = ~pi455 & ~n7571;
  assign n7655 = ~n7653 & ~n7654;
  assign n7656 = pi452 & ~n7655;
  assign n7657 = ~n7652 & ~n7656;
  assign n7658 = ~pi355 & ~n7657;
  assign n7659 = ~pi452 & ~n7655;
  assign n7660 = pi452 & ~n7651;
  assign n7661 = ~n7659 & ~n7660;
  assign n7662 = pi355 & ~n7661;
  assign n7663 = ~n7658 & ~n7662;
  assign n7664 = pi458 & ~n7663;
  assign n7665 = ~pi355 & ~n7661;
  assign n7666 = pi355 & ~n7657;
  assign n7667 = ~n7665 & ~n7666;
  assign n7668 = ~pi458 & ~n7667;
  assign n7669 = n7633 & ~n7664;
  assign n7670 = ~n7668 & n7669;
  assign n7671 = pi458 & ~n7667;
  assign n7672 = ~pi458 & ~n7663;
  assign n7673 = ~n7633 & ~n7671;
  assign n7674 = ~n7672 & n7673;
  assign n7675 = pi1196 & ~n7670;
  assign n7676 = ~n7674 & n7675;
  assign n7677 = ~pi1196 & ~n7571;
  assign n7678 = ~pi1198 & ~n7677;
  assign n7679 = ~n7676 & n7678;
  assign n7680 = ~n7648 & ~n7679;
  assign n7681 = ~n7443 & ~n7680;
  assign n7682 = n7443 & n7645;
  assign n7683 = ~n7681 & ~n7682;
  assign n7684 = ~pi351 & pi1199;
  assign n7685 = n7683 & ~n7684;
  assign n7686 = pi1199 & ~n7645;
  assign n7687 = ~pi351 & n7686;
  assign n7688 = ~n7685 & ~n7687;
  assign n7689 = ~pi461 & ~n7688;
  assign n7690 = pi351 & pi1199;
  assign n7691 = n7683 & ~n7690;
  assign n7692 = pi351 & n7686;
  assign n7693 = ~n7691 & ~n7692;
  assign n7694 = pi461 & ~n7693;
  assign n7695 = ~n7689 & ~n7694;
  assign n7696 = ~pi357 & ~n7695;
  assign n7697 = ~pi461 & ~n7693;
  assign n7698 = pi461 & ~n7688;
  assign n7699 = ~n7697 & ~n7698;
  assign n7700 = pi357 & ~n7699;
  assign n7701 = ~n7696 & ~n7700;
  assign n7702 = ~pi356 & ~n7701;
  assign n7703 = ~pi357 & ~n7699;
  assign n7704 = pi357 & ~n7695;
  assign n7705 = ~n7703 & ~n7704;
  assign n7706 = pi356 & ~n7705;
  assign n7707 = ~n7702 & ~n7706;
  assign n7708 = ~n7418 & ~n7707;
  assign n7709 = ~pi356 & ~n7705;
  assign n7710 = pi356 & ~n7701;
  assign n7711 = ~n7709 & ~n7710;
  assign n7712 = n7418 & ~n7711;
  assign n7713 = ~pi591 & ~n7708;
  assign n7714 = ~n7712 & n7713;
  assign n7715 = pi591 & n7571;
  assign n7716 = pi590 & ~n7715;
  assign n7717 = ~n7714 & n7716;
  assign n7718 = ~pi285 & ~pi286;
  assign n7719 = ~pi289 & n7718;
  assign n7720 = ~pi288 & n7719;
  assign n7721 = ~pi363 & ~pi372;
  assign n7722 = pi363 & pi372;
  assign n7723 = ~n7721 & ~n7722;
  assign n7724 = pi386 & ~n7723;
  assign n7725 = ~pi386 & n7723;
  assign n7726 = ~n7724 & ~n7725;
  assign n7727 = pi338 & ~pi388;
  assign n7728 = ~pi338 & pi388;
  assign n7729 = ~n7727 & ~n7728;
  assign n7730 = pi337 & ~pi339;
  assign n7731 = ~pi337 & pi339;
  assign n7732 = ~n7730 & ~n7731;
  assign n7733 = pi387 & n7732;
  assign n7734 = ~pi387 & ~n7732;
  assign n7735 = ~n7733 & ~n7734;
  assign n7736 = pi380 & ~n7735;
  assign n7737 = ~pi380 & n7735;
  assign n7738 = ~n7736 & ~n7737;
  assign n7739 = n7729 & ~n7738;
  assign n7740 = ~n7729 & n7738;
  assign n7741 = ~n7739 & ~n7740;
  assign n7742 = n7726 & n7741;
  assign n7743 = ~n7726 & ~n7741;
  assign n7744 = ~n7742 & ~n7743;
  assign n7745 = pi1196 & ~n7744;
  assign n7746 = ~pi368 & ~pi389;
  assign n7747 = pi368 & pi389;
  assign n7748 = ~n7746 & ~n7747;
  assign n7749 = pi365 & ~pi447;
  assign n7750 = ~pi365 & pi447;
  assign n7751 = ~n7749 & ~n7750;
  assign n7752 = pi336 & ~pi383;
  assign n7753 = ~pi336 & pi383;
  assign n7754 = ~n7752 & ~n7753;
  assign n7755 = pi364 & ~pi366;
  assign n7756 = ~pi364 & pi366;
  assign n7757 = ~n7755 & ~n7756;
  assign n7758 = n7754 & n7757;
  assign n7759 = ~n7754 & ~n7757;
  assign n7760 = ~n7758 & ~n7759;
  assign n7761 = n7751 & n7760;
  assign n7762 = ~n7751 & ~n7760;
  assign n7763 = ~n7761 & ~n7762;
  assign n7764 = n7748 & n7763;
  assign n7765 = ~n7748 & ~n7763;
  assign n7766 = ~n7764 & ~n7765;
  assign n7767 = pi367 & ~n7766;
  assign n7768 = ~pi367 & n7766;
  assign n7769 = ~n7767 & ~n7768;
  assign n7770 = pi1197 & n7769;
  assign n7771 = ~n7745 & ~n7770;
  assign n7772 = pi377 & pi592;
  assign n7773 = ~n7571 & ~n7772;
  assign n7774 = pi379 & ~pi382;
  assign n7775 = ~pi379 & pi382;
  assign n7776 = ~n7774 & ~n7775;
  assign n7777 = pi376 & ~pi439;
  assign n7778 = ~pi376 & pi439;
  assign n7779 = ~n7777 & ~n7778;
  assign n7780 = pi381 & n7779;
  assign n7781 = ~pi381 & ~n7779;
  assign n7782 = ~n7780 & ~n7781;
  assign n7783 = pi317 & ~pi385;
  assign n7784 = ~pi317 & pi385;
  assign n7785 = ~n7783 & ~n7784;
  assign n7786 = pi378 & n7785;
  assign n7787 = ~pi378 & ~n7785;
  assign n7788 = ~n7786 & ~n7787;
  assign n7789 = n7782 & ~n7788;
  assign n7790 = ~n7782 & n7788;
  assign n7791 = ~n7789 & ~n7790;
  assign n7792 = n7776 & n7791;
  assign n7793 = ~n7776 & ~n7791;
  assign n7794 = ~n7792 & ~n7793;
  assign n7795 = ~n7607 & n7772;
  assign n7796 = ~n7794 & ~n7795;
  assign n7797 = ~n7773 & n7796;
  assign n7798 = ~pi377 & pi592;
  assign n7799 = ~n7571 & ~n7798;
  assign n7800 = ~n7607 & n7798;
  assign n7801 = n7794 & ~n7800;
  assign n7802 = ~n7799 & n7801;
  assign n7803 = ~n7797 & ~n7802;
  assign n7804 = n7771 & ~n7803;
  assign n7805 = pi592 & ~n7607;
  assign n7806 = ~pi592 & ~n7571;
  assign n7807 = ~n7805 & ~n7806;
  assign n7808 = ~n7771 & n7807;
  assign n7809 = ~n7804 & ~n7808;
  assign n7810 = pi1199 & n7809;
  assign n7811 = n7571 & ~n7770;
  assign n7812 = n7770 & n7807;
  assign n7813 = ~n7811 & ~n7812;
  assign n7814 = n7744 & ~n7813;
  assign n7815 = ~pi1196 & ~n7770;
  assign n7816 = n7807 & ~n7815;
  assign n7817 = ~pi1196 & n7811;
  assign n7818 = ~n7816 & ~n7817;
  assign n7819 = ~n7744 & ~n7818;
  assign n7820 = ~pi1199 & ~n7814;
  assign n7821 = ~n7819 & n7820;
  assign n7822 = ~n7810 & ~n7821;
  assign n7823 = ~pi374 & ~n7822;
  assign n7824 = ~pi1198 & n7821;
  assign n7825 = ~pi1198 & pi1199;
  assign n7826 = n7809 & n7825;
  assign n7827 = pi1198 & ~n7807;
  assign n7828 = ~n7826 & ~n7827;
  assign n7829 = ~n7824 & n7828;
  assign n7830 = pi374 & ~n7829;
  assign n7831 = ~n7823 & ~n7830;
  assign n7832 = pi369 & ~n7831;
  assign n7833 = ~pi374 & ~n7829;
  assign n7834 = pi374 & ~n7822;
  assign n7835 = ~n7833 & ~n7834;
  assign n7836 = ~pi369 & ~n7835;
  assign n7837 = ~n7832 & ~n7836;
  assign n7838 = ~pi370 & ~n7837;
  assign n7839 = ~pi369 & ~n7831;
  assign n7840 = pi369 & ~n7835;
  assign n7841 = ~n7839 & ~n7840;
  assign n7842 = pi370 & ~n7841;
  assign n7843 = ~n7838 & ~n7842;
  assign n7844 = ~pi371 & ~n7843;
  assign n7845 = ~pi370 & ~n7841;
  assign n7846 = pi370 & ~n7837;
  assign n7847 = ~n7845 & ~n7846;
  assign n7848 = pi371 & ~n7847;
  assign n7849 = ~n7844 & ~n7848;
  assign n7850 = ~pi373 & ~n7849;
  assign n7851 = ~pi371 & ~n7847;
  assign n7852 = pi371 & ~n7843;
  assign n7853 = ~n7851 & ~n7852;
  assign n7854 = pi373 & ~n7853;
  assign n7855 = ~n7850 & ~n7854;
  assign n7856 = ~pi375 & n7855;
  assign n7857 = pi384 & ~pi442;
  assign n7858 = ~pi384 & pi442;
  assign n7859 = ~n7857 & ~n7858;
  assign n7860 = pi440 & ~n7859;
  assign n7861 = ~pi440 & n7859;
  assign n7862 = ~n7860 & ~n7861;
  assign n7863 = ~pi373 & ~n7853;
  assign n7864 = pi373 & ~n7849;
  assign n7865 = ~n7863 & ~n7864;
  assign n7866 = pi375 & n7865;
  assign n7867 = ~n7856 & n7862;
  assign n7868 = ~n7866 & n7867;
  assign n7869 = pi375 & n7855;
  assign n7870 = ~pi375 & n7865;
  assign n7871 = ~n7862 & ~n7869;
  assign n7872 = ~n7870 & n7871;
  assign n7873 = ~pi591 & ~n7868;
  assign n7874 = ~n7872 & n7873;
  assign n7875 = pi1197 & ~n7645;
  assign n7876 = pi328 & ~pi408;
  assign n7877 = ~pi328 & pi408;
  assign n7878 = ~n7876 & ~n7877;
  assign n7879 = ~pi394 & ~pi396;
  assign n7880 = pi394 & pi396;
  assign n7881 = ~n7879 & ~n7880;
  assign n7882 = n7878 & ~n7881;
  assign n7883 = ~n7878 & n7881;
  assign n7884 = ~n7882 & ~n7883;
  assign n7885 = pi398 & ~pi399;
  assign n7886 = ~pi398 & pi399;
  assign n7887 = ~n7885 & ~n7886;
  assign n7888 = pi395 & n7887;
  assign n7889 = ~pi395 & ~n7887;
  assign n7890 = ~n7888 & ~n7889;
  assign n7891 = pi329 & ~n7890;
  assign n7892 = ~pi329 & n7890;
  assign n7893 = ~n7891 & ~n7892;
  assign n7894 = pi400 & ~n7893;
  assign n7895 = ~pi400 & n7893;
  assign n7896 = ~n7894 & ~n7895;
  assign n7897 = n7884 & n7896;
  assign n7898 = ~n7884 & ~n7896;
  assign n7899 = ~n7897 & ~n7898;
  assign n7900 = pi1198 & ~n7899;
  assign n7901 = n7645 & n7900;
  assign n7902 = pi390 & ~pi410;
  assign n7903 = ~pi390 & pi410;
  assign n7904 = ~n7902 & ~n7903;
  assign n7905 = pi397 & ~pi412;
  assign n7906 = ~pi397 & pi412;
  assign n7907 = ~n7905 & ~n7906;
  assign n7908 = pi404 & n7907;
  assign n7909 = ~pi404 & ~n7907;
  assign n7910 = ~n7908 & ~n7909;
  assign n7911 = pi319 & ~pi324;
  assign n7912 = ~pi319 & pi324;
  assign n7913 = ~n7911 & ~n7912;
  assign n7914 = pi456 & ~n7913;
  assign n7915 = ~pi456 & n7913;
  assign n7916 = ~n7914 & ~n7915;
  assign n7917 = n7910 & ~n7916;
  assign n7918 = ~n7910 & n7916;
  assign n7919 = ~n7917 & ~n7918;
  assign n7920 = n7904 & n7919;
  assign n7921 = ~n7904 & ~n7919;
  assign n7922 = ~n7920 & ~n7921;
  assign n7923 = pi411 & n7922;
  assign n7924 = ~pi411 & ~n7922;
  assign n7925 = ~n7923 & ~n7924;
  assign n7926 = n7545 & n7925;
  assign n7927 = n7542 & ~n7926;
  assign n7928 = n7595 & ~n7927;
  assign n7929 = ~n7563 & n7600;
  assign n7930 = n7557 & n7925;
  assign n7931 = n7558 & ~n7930;
  assign n7932 = n7929 & ~n7931;
  assign n7933 = ~pi75 & ~pi592;
  assign n7934 = pi1196 & n7933;
  assign n7935 = ~n7932 & n7934;
  assign n7936 = ~n7928 & n7935;
  assign n7937 = ~pi1196 & n7568;
  assign n7938 = ~n7936 & ~n7937;
  assign n7939 = ~pi1199 & ~n7938;
  assign n7940 = pi318 & ~pi409;
  assign n7941 = ~pi318 & pi409;
  assign n7942 = ~n7940 & ~n7941;
  assign n7943 = pi401 & ~pi402;
  assign n7944 = ~pi401 & pi402;
  assign n7945 = ~n7943 & ~n7944;
  assign n7946 = pi406 & n7945;
  assign n7947 = ~pi406 & ~n7945;
  assign n7948 = ~n7946 & ~n7947;
  assign n7949 = ~pi403 & ~pi405;
  assign n7950 = pi403 & pi405;
  assign n7951 = ~n7949 & ~n7950;
  assign n7952 = pi325 & ~pi326;
  assign n7953 = ~pi325 & pi326;
  assign n7954 = ~n7952 & ~n7953;
  assign n7955 = n7951 & n7954;
  assign n7956 = ~n7951 & ~n7954;
  assign n7957 = ~n7955 & ~n7956;
  assign n7958 = n7948 & ~n7957;
  assign n7959 = ~n7948 & n7957;
  assign n7960 = ~n7958 & ~n7959;
  assign n7961 = n7942 & n7960;
  assign n7962 = ~n7942 & ~n7960;
  assign n7963 = ~n7961 & ~n7962;
  assign n7964 = pi1196 & ~n7925;
  assign n7965 = ~pi75 & n7964;
  assign n7966 = ~n7963 & ~n7965;
  assign n7967 = n7545 & n7966;
  assign n7968 = n7542 & ~n7967;
  assign n7969 = n7595 & ~n7968;
  assign n7970 = n7557 & ~n7963;
  assign n7971 = n7558 & ~n7970;
  assign n7972 = n7929 & ~n7971;
  assign n7973 = ~pi1196 & n7972;
  assign n7974 = ~n7931 & n7972;
  assign n7975 = pi1199 & n7933;
  assign n7976 = ~n7973 & n7975;
  assign n7977 = ~n7974 & n7976;
  assign n7978 = ~n7969 & n7977;
  assign n7979 = ~n7569 & ~n7933;
  assign n7980 = ~n7978 & ~n7979;
  assign n7981 = ~n7939 & n7980;
  assign n7982 = pi567 & ~n7981;
  assign n7983 = n7483 & ~n7900;
  assign n7984 = ~n7982 & n7983;
  assign n7985 = ~n7901 & ~n7984;
  assign n7986 = ~pi1197 & n7985;
  assign n7987 = ~n7875 & ~n7986;
  assign n7988 = pi333 & ~n7987;
  assign n7989 = ~pi333 & n7985;
  assign n7990 = ~n7988 & ~n7989;
  assign n7991 = pi391 & ~n7990;
  assign n7992 = pi333 & ~n7985;
  assign n7993 = ~pi333 & n7987;
  assign n7994 = ~n7992 & ~n7993;
  assign n7995 = ~pi391 & n7994;
  assign n7996 = ~n7991 & ~n7995;
  assign n7997 = ~pi392 & ~n7996;
  assign n7998 = ~pi391 & ~n7990;
  assign n7999 = pi391 & n7994;
  assign n8000 = ~n7998 & ~n7999;
  assign n8001 = pi392 & ~n8000;
  assign n8002 = ~n7997 & ~n8001;
  assign n8003 = ~pi393 & ~n8002;
  assign n8004 = ~pi392 & ~n8000;
  assign n8005 = pi392 & ~n7996;
  assign n8006 = ~n8004 & ~n8005;
  assign n8007 = pi393 & ~n8006;
  assign n8008 = ~n8003 & ~n8007;
  assign n8009 = ~pi334 & n8008;
  assign n8010 = pi407 & ~pi463;
  assign n8011 = ~pi407 & pi463;
  assign n8012 = ~n8010 & ~n8011;
  assign n8013 = pi335 & ~pi413;
  assign n8014 = ~pi335 & pi413;
  assign n8015 = ~n8013 & ~n8014;
  assign n8016 = n8012 & n8015;
  assign n8017 = ~n8012 & ~n8015;
  assign n8018 = ~n8016 & ~n8017;
  assign n8019 = ~pi393 & ~n8006;
  assign n8020 = pi393 & ~n8002;
  assign n8021 = ~n8019 & ~n8020;
  assign n8022 = pi334 & n8021;
  assign n8023 = ~n8009 & n8018;
  assign n8024 = ~n8022 & n8023;
  assign n8025 = ~pi334 & n8021;
  assign n8026 = pi334 & n8008;
  assign n8027 = ~n8018 & ~n8025;
  assign n8028 = ~n8026 & n8027;
  assign n8029 = pi591 & ~n8024;
  assign n8030 = ~n8028 & n8029;
  assign n8031 = ~pi590 & ~n8030;
  assign n8032 = ~n7874 & n8031;
  assign n8033 = n7720 & ~n8032;
  assign n8034 = ~n7717 & n8033;
  assign n8035 = n7487 & n7548;
  assign n8036 = pi1091 & ~n8035;
  assign n8037 = n7486 & ~n8036;
  assign n8038 = ~pi122 & pi1093;
  assign n8039 = ~pi98 & n7496;
  assign n8040 = n8038 & n8039;
  assign n8041 = ~pi1091 & ~n8040;
  assign n8042 = n8037 & ~n8041;
  assign n8043 = n7496 & n8038;
  assign n8044 = ~pi1091 & n8043;
  assign n8045 = ~pi98 & n8044;
  assign n8046 = ~n7486 & n8045;
  assign n8047 = pi75 & ~n8046;
  assign n8048 = ~n8042 & n8047;
  assign n8049 = ~pi39 & ~n7523;
  assign n8050 = ~pi122 & n8039;
  assign n8051 = pi122 & n7499;
  assign n8052 = ~n8050 & ~n8051;
  assign n8053 = pi1093 & ~n8052;
  assign n8054 = n7524 & ~n8053;
  assign n8055 = n8049 & ~n8054;
  assign n8056 = pi1091 & ~n7529;
  assign n8057 = ~n8041 & ~n8056;
  assign n8058 = n6206 & n8057;
  assign n8059 = ~n6206 & n8045;
  assign n8060 = ~n8058 & ~n8059;
  assign n8061 = n6197 & n8060;
  assign n8062 = ~n6200 & n8057;
  assign n8063 = n6200 & n8045;
  assign n8064 = ~n8062 & ~n8063;
  assign n8065 = ~n6197 & n8064;
  assign n8066 = ~pi223 & n5777;
  assign n8067 = ~n8061 & n8066;
  assign n8068 = ~n8065 & n8067;
  assign n8069 = n8045 & ~n8066;
  assign n8070 = ~pi299 & ~n8069;
  assign n8071 = ~n8068 & n8070;
  assign n8072 = n6223 & n8060;
  assign n8073 = ~n6223 & n8064;
  assign n8074 = ~pi216 & n6442;
  assign n8075 = ~n8072 & n8074;
  assign n8076 = ~n8073 & n8075;
  assign n8077 = n8045 & ~n8074;
  assign n8078 = pi299 & ~n8077;
  assign n8079 = ~n8076 & n8078;
  assign n8080 = pi39 & ~n8071;
  assign n8081 = ~n8079 & n8080;
  assign n8082 = ~n8055 & ~n8081;
  assign n8083 = ~pi38 & ~n8082;
  assign n8084 = pi38 & n8045;
  assign n8085 = ~pi100 & ~n8084;
  assign n8086 = ~n8083 & n8085;
  assign n8087 = pi228 & ~n7485;
  assign n8088 = pi1091 & ~n7549;
  assign n8089 = ~n8041 & ~n8088;
  assign n8090 = n8087 & ~n8089;
  assign n8091 = ~n8045 & ~n8087;
  assign n8092 = n3182 & ~n8091;
  assign n8093 = ~n8090 & n8092;
  assign n8094 = ~n3182 & n8045;
  assign n8095 = pi100 & ~n8094;
  assign n8096 = ~n8093 & n8095;
  assign n8097 = ~pi87 & ~n8096;
  assign n8098 = ~n8086 & n8097;
  assign n8099 = pi122 & n7557;
  assign n8100 = ~n8050 & ~n8099;
  assign n8101 = pi1093 & ~n8100;
  assign n8102 = n7598 & ~n8101;
  assign n8103 = n3208 & ~n7597;
  assign n8104 = ~n8102 & n8103;
  assign n8105 = ~n8045 & ~n8104;
  assign n8106 = pi87 & ~n8105;
  assign n8107 = ~pi75 & ~n8106;
  assign n8108 = ~n8098 & n8107;
  assign n8109 = ~n8048 & ~n8108;
  assign n8110 = pi567 & ~n8109;
  assign n8111 = n7483 & ~n8110;
  assign n8112 = pi567 & n8045;
  assign n8113 = ~n7444 & n8112;
  assign n8114 = ~n8111 & ~n8113;
  assign n8115 = pi592 & n8114;
  assign n8116 = ~n7643 & ~n8115;
  assign n8117 = n7443 & ~n8116;
  assign n8118 = pi455 & ~n8116;
  assign n8119 = ~pi455 & n8114;
  assign n8120 = ~n8118 & ~n8119;
  assign n8121 = ~pi452 & ~n8120;
  assign n8122 = pi355 & ~n7636;
  assign n8123 = ~pi355 & n7636;
  assign n8124 = ~n8122 & ~n8123;
  assign n8125 = ~pi455 & ~n8116;
  assign n8126 = pi455 & n8114;
  assign n8127 = ~n8125 & ~n8126;
  assign n8128 = pi452 & ~n8127;
  assign n8129 = ~n8121 & ~n8124;
  assign n8130 = ~n8128 & n8129;
  assign n8131 = ~pi452 & ~n8127;
  assign n8132 = pi452 & ~n8120;
  assign n8133 = n8124 & ~n8131;
  assign n8134 = ~n8132 & n8133;
  assign n8135 = pi1196 & ~n8130;
  assign n8136 = ~n8134 & n8135;
  assign n8137 = ~pi1196 & n8114;
  assign n8138 = ~pi1198 & ~n8137;
  assign n8139 = ~n8136 & n8138;
  assign n8140 = ~n7611 & n8114;
  assign n8141 = n7614 & ~n8140;
  assign n8142 = ~n7572 & n8114;
  assign n8143 = n7609 & ~n8142;
  assign n8144 = ~n7640 & ~n8141;
  assign n8145 = ~n8143 & n8144;
  assign n8146 = n7640 & ~n8116;
  assign n8147 = pi1198 & ~n8146;
  assign n8148 = ~n8145 & n8147;
  assign n8149 = ~n7443 & ~n8148;
  assign n8150 = ~n8139 & n8149;
  assign n8151 = ~n8117 & ~n8150;
  assign n8152 = ~n7684 & ~n8151;
  assign n8153 = pi1199 & ~n8116;
  assign n8154 = ~pi351 & n8153;
  assign n8155 = ~n8152 & ~n8154;
  assign n8156 = ~pi461 & ~n8155;
  assign n8157 = ~n7690 & ~n8151;
  assign n8158 = pi351 & n8153;
  assign n8159 = ~n8157 & ~n8158;
  assign n8160 = pi461 & ~n8159;
  assign n8161 = ~n8156 & ~n8160;
  assign n8162 = ~pi357 & ~n8161;
  assign n8163 = ~pi461 & ~n8159;
  assign n8164 = pi461 & ~n8155;
  assign n8165 = ~n8163 & ~n8164;
  assign n8166 = pi357 & ~n8165;
  assign n8167 = ~n8162 & ~n8166;
  assign n8168 = ~pi356 & ~n8167;
  assign n8169 = ~pi357 & ~n8165;
  assign n8170 = pi357 & ~n8161;
  assign n8171 = ~n8169 & ~n8170;
  assign n8172 = pi356 & ~n8171;
  assign n8173 = ~n8168 & ~n8172;
  assign n8174 = ~n7418 & ~n8173;
  assign n8175 = ~pi356 & ~n8171;
  assign n8176 = pi356 & ~n8167;
  assign n8177 = ~n8175 & ~n8176;
  assign n8178 = n7418 & ~n8177;
  assign n8179 = ~pi591 & ~n8174;
  assign n8180 = ~n8178 & n8179;
  assign n8181 = pi591 & ~n8114;
  assign n8182 = pi590 & ~n8181;
  assign n8183 = ~n8180 & n8182;
  assign n8184 = pi375 & n7862;
  assign n8185 = ~pi375 & ~n7862;
  assign n8186 = ~n8184 & ~n8185;
  assign n8187 = pi373 & ~n8186;
  assign n8188 = ~pi373 & n8186;
  assign n8189 = ~n8187 & ~n8188;
  assign n8190 = ~pi592 & n8114;
  assign n8191 = ~n7805 & ~n8190;
  assign n8192 = ~n7771 & n8191;
  assign n8193 = n7771 & ~n8114;
  assign n8194 = ~pi1199 & ~n8193;
  assign n8195 = ~n8192 & n8194;
  assign n8196 = ~n7798 & n8114;
  assign n8197 = n7801 & ~n8196;
  assign n8198 = ~n7772 & n8114;
  assign n8199 = n7796 & ~n8198;
  assign n8200 = ~n8197 & ~n8199;
  assign n8201 = n7771 & ~n8200;
  assign n8202 = pi1199 & ~n8192;
  assign n8203 = ~n8201 & n8202;
  assign n8204 = ~n8195 & ~n8203;
  assign n8205 = ~pi374 & ~n8204;
  assign n8206 = ~pi1198 & ~n8204;
  assign n8207 = pi1198 & ~n8191;
  assign n8208 = ~n8206 & ~n8207;
  assign n8209 = pi374 & ~n8208;
  assign n8210 = ~n8205 & ~n8209;
  assign n8211 = pi369 & ~n8210;
  assign n8212 = ~pi374 & ~n8208;
  assign n8213 = pi374 & ~n8204;
  assign n8214 = ~n8212 & ~n8213;
  assign n8215 = ~pi369 & ~n8214;
  assign n8216 = ~n8211 & ~n8215;
  assign n8217 = ~pi370 & ~n8216;
  assign n8218 = ~pi369 & ~n8210;
  assign n8219 = pi369 & ~n8214;
  assign n8220 = ~n8218 & ~n8219;
  assign n8221 = pi370 & ~n8220;
  assign n8222 = ~n8217 & ~n8221;
  assign n8223 = ~pi371 & ~n8222;
  assign n8224 = ~pi370 & ~n8220;
  assign n8225 = pi370 & ~n8216;
  assign n8226 = ~n8224 & ~n8225;
  assign n8227 = pi371 & ~n8226;
  assign n8228 = ~n8223 & ~n8227;
  assign n8229 = ~n8189 & ~n8228;
  assign n8230 = ~pi371 & ~n8226;
  assign n8231 = pi371 & ~n8222;
  assign n8232 = ~n8230 & ~n8231;
  assign n8233 = n8189 & ~n8232;
  assign n8234 = ~pi591 & ~n8229;
  assign n8235 = ~n8233 & n8234;
  assign n8236 = pi334 & ~n8018;
  assign n8237 = ~pi334 & n8018;
  assign n8238 = ~n8236 & ~n8237;
  assign n8239 = pi393 & n8238;
  assign n8240 = ~pi393 & ~n8238;
  assign n8241 = ~n8239 & ~n8240;
  assign n8242 = ~pi592 & pi1196;
  assign n8243 = n7925 & n8040;
  assign n8244 = ~pi1091 & n8243;
  assign n8245 = pi567 & n8244;
  assign n8246 = ~n7444 & n8245;
  assign n8247 = ~n7963 & n8039;
  assign n8248 = n8246 & n8247;
  assign n8249 = n8242 & ~n8248;
  assign n8250 = ~n8074 & n8244;
  assign n8251 = pi299 & ~n8250;
  assign n8252 = ~n7963 & n8040;
  assign n8253 = ~pi1091 & n8252;
  assign n8254 = ~n8074 & n8253;
  assign n8255 = pi299 & ~n8254;
  assign n8256 = ~n8251 & ~n8255;
  assign n8257 = ~n7963 & n8244;
  assign n8258 = n6206 & n7530;
  assign n8259 = ~n8257 & ~n8258;
  assign n8260 = n6223 & n8259;
  assign n8261 = ~n6200 & n7530;
  assign n8262 = ~n8257 & ~n8261;
  assign n8263 = ~n6223 & n8262;
  assign n8264 = n8074 & ~n8260;
  assign n8265 = ~n8263 & n8264;
  assign n8266 = ~n8256 & ~n8265;
  assign n8267 = ~n8066 & n8244;
  assign n8268 = ~pi299 & ~n8267;
  assign n8269 = ~n8066 & n8253;
  assign n8270 = ~pi299 & ~n8269;
  assign n8271 = ~n8268 & ~n8270;
  assign n8272 = n6197 & n8259;
  assign n8273 = ~n6197 & n8262;
  assign n8274 = n8066 & ~n8272;
  assign n8275 = ~n8273 & n8274;
  assign n8276 = ~n8271 & ~n8275;
  assign n8277 = pi39 & ~n8266;
  assign n8278 = ~n8276 & n8277;
  assign n8279 = n7524 & ~n7925;
  assign n8280 = n8055 & ~n8279;
  assign n8281 = n7499 & ~n7963;
  assign n8282 = pi122 & ~n8281;
  assign n8283 = ~pi122 & ~n8247;
  assign n8284 = pi1093 & ~n8283;
  assign n8285 = ~n8282 & n8284;
  assign n8286 = n7524 & ~n8285;
  assign n8287 = n8280 & ~n8286;
  assign n8288 = ~n8278 & ~n8287;
  assign n8289 = ~pi38 & ~n8288;
  assign n8290 = pi38 & n8244;
  assign n8291 = ~pi100 & ~n8290;
  assign n8292 = pi38 & n8253;
  assign n8293 = ~pi100 & ~n8292;
  assign n8294 = ~n8291 & ~n8293;
  assign n8295 = ~n8289 & ~n8294;
  assign n8296 = n6242 & n7550;
  assign n8297 = n6170 & ~n6243;
  assign n8298 = ~n6242 & ~n8297;
  assign n8299 = ~pi1091 & ~n8257;
  assign n8300 = n8298 & ~n8299;
  assign n8301 = ~n8088 & n8300;
  assign n8302 = ~n8296 & ~n8301;
  assign n8303 = pi228 & ~n8302;
  assign n8304 = pi228 & n8298;
  assign n8305 = n8257 & ~n8304;
  assign n8306 = pi232 & ~n8305;
  assign n8307 = ~n8303 & n8306;
  assign n8308 = ~pi232 & ~n8257;
  assign n8309 = ~n7551 & n8308;
  assign n8310 = n3182 & ~n8309;
  assign n8311 = ~n8307 & n8310;
  assign n8312 = ~n3182 & n8257;
  assign n8313 = pi100 & ~n8312;
  assign n8314 = ~n8311 & n8313;
  assign n8315 = ~n8295 & ~n8314;
  assign n8316 = ~pi87 & ~n8315;
  assign n8317 = ~n3208 & n8244;
  assign n8318 = pi87 & ~n8317;
  assign n8319 = ~n3208 & n8253;
  assign n8320 = pi87 & ~n8319;
  assign n8321 = ~n8318 & ~n8320;
  assign n8322 = n7598 & ~n7925;
  assign n8323 = n7598 & n7963;
  assign n8324 = n8104 & ~n8323;
  assign n8325 = ~n8322 & n8324;
  assign n8326 = ~n8321 & ~n8325;
  assign n8327 = ~n8316 & ~n8326;
  assign n8328 = ~pi75 & ~n8327;
  assign n8329 = ~n7486 & n8244;
  assign n8330 = pi75 & ~n8329;
  assign n8331 = ~n7486 & n8253;
  assign n8332 = pi75 & ~n8331;
  assign n8333 = ~n8330 & ~n8332;
  assign n8334 = n8037 & ~n8299;
  assign n8335 = ~n8333 & ~n8334;
  assign n8336 = ~n8328 & ~n8335;
  assign n8337 = n8249 & ~n8336;
  assign n8338 = pi567 & n8253;
  assign n8339 = ~n7444 & n8338;
  assign n8340 = ~pi592 & ~pi1196;
  assign n8341 = ~n8339 & n8340;
  assign n8342 = n8320 & ~n8324;
  assign n8343 = n7554 & ~n8253;
  assign n8344 = n8049 & ~n8286;
  assign n8345 = ~n8253 & ~n8261;
  assign n8346 = ~n6223 & n8345;
  assign n8347 = ~n8253 & ~n8258;
  assign n8348 = n6223 & n8347;
  assign n8349 = n8074 & ~n8346;
  assign n8350 = ~n8348 & n8349;
  assign n8351 = n8255 & ~n8350;
  assign n8352 = ~n6197 & n8345;
  assign n8353 = n6197 & n8347;
  assign n8354 = n8066 & ~n8352;
  assign n8355 = ~n8353 & n8354;
  assign n8356 = n8270 & ~n8355;
  assign n8357 = pi39 & ~n8351;
  assign n8358 = ~n8356 & n8357;
  assign n8359 = ~n8344 & ~n8358;
  assign n8360 = ~pi38 & ~n8359;
  assign n8361 = n8293 & ~n8360;
  assign n8362 = ~n8343 & ~n8361;
  assign n8363 = ~pi87 & ~n8362;
  assign n8364 = ~n8342 & ~n8363;
  assign n8365 = ~pi75 & ~n8364;
  assign n8366 = ~pi1091 & ~n8252;
  assign n8367 = n8037 & ~n8366;
  assign n8368 = n8332 & ~n8367;
  assign n8369 = ~n8365 & ~n8368;
  assign n8370 = n8341 & ~n8369;
  assign n8371 = ~n8337 & ~n8370;
  assign n8372 = pi567 & ~n8371;
  assign n8373 = ~n8249 & ~n8341;
  assign n8374 = ~n7483 & ~n8373;
  assign n8375 = pi1199 & ~n8374;
  assign n8376 = ~n8372 & n8375;
  assign n8377 = ~n8244 & ~n8261;
  assign n8378 = ~n6223 & n8377;
  assign n8379 = ~n8244 & ~n8258;
  assign n8380 = n6223 & n8379;
  assign n8381 = n8074 & ~n8378;
  assign n8382 = ~n8380 & n8381;
  assign n8383 = n8251 & ~n8382;
  assign n8384 = ~n6197 & n8377;
  assign n8385 = n6197 & n8379;
  assign n8386 = n8066 & ~n8384;
  assign n8387 = ~n8385 & n8386;
  assign n8388 = n8268 & ~n8387;
  assign n8389 = pi39 & ~n8383;
  assign n8390 = ~n8388 & n8389;
  assign n8391 = ~n8280 & ~n8390;
  assign n8392 = ~pi38 & ~n8391;
  assign n8393 = n8291 & ~n8392;
  assign n8394 = n7554 & ~n8244;
  assign n8395 = ~n8393 & ~n8394;
  assign n8396 = ~pi87 & ~n8395;
  assign n8397 = n8104 & ~n8322;
  assign n8398 = n8318 & ~n8397;
  assign n8399 = ~n8396 & ~n8398;
  assign n8400 = ~pi75 & ~n8399;
  assign n8401 = ~pi1091 & ~n8243;
  assign n8402 = n8037 & ~n8401;
  assign n8403 = n8330 & ~n8402;
  assign n8404 = ~n8400 & ~n8403;
  assign n8405 = pi567 & ~n8404;
  assign n8406 = n7483 & ~n8405;
  assign n8407 = n8242 & ~n8246;
  assign n8408 = ~n8406 & n8407;
  assign n8409 = ~pi1199 & ~n8137;
  assign n8410 = ~n8408 & n8409;
  assign n8411 = ~n7900 & ~n8410;
  assign n8412 = ~n8376 & n8411;
  assign n8413 = n7643 & n7900;
  assign n8414 = ~n8115 & ~n8413;
  assign n8415 = ~n8412 & n8414;
  assign n8416 = ~pi1197 & ~n8415;
  assign n8417 = pi1197 & ~n8116;
  assign n8418 = ~n8416 & ~n8417;
  assign n8419 = ~pi333 & ~n8418;
  assign n8420 = pi333 & ~n8415;
  assign n8421 = ~n8419 & ~n8420;
  assign n8422 = ~pi391 & ~n8421;
  assign n8423 = ~pi333 & ~n8415;
  assign n8424 = pi333 & ~n8418;
  assign n8425 = ~n8423 & ~n8424;
  assign n8426 = pi391 & ~n8425;
  assign n8427 = ~n8422 & ~n8426;
  assign n8428 = ~pi392 & ~n8427;
  assign n8429 = ~pi391 & ~n8425;
  assign n8430 = pi391 & ~n8421;
  assign n8431 = ~n8429 & ~n8430;
  assign n8432 = pi392 & ~n8431;
  assign n8433 = ~n8428 & ~n8432;
  assign n8434 = ~n8241 & ~n8433;
  assign n8435 = ~pi392 & ~n8431;
  assign n8436 = pi392 & ~n8427;
  assign n8437 = ~n8435 & ~n8436;
  assign n8438 = n8241 & ~n8437;
  assign n8439 = pi591 & ~n8434;
  assign n8440 = ~n8438 & n8439;
  assign n8441 = ~pi590 & ~n8440;
  assign n8442 = ~n8235 & n8441;
  assign n8443 = ~n7720 & ~n8442;
  assign n8444 = ~n8183 & n8443;
  assign n8445 = ~pi588 & ~n8444;
  assign n8446 = ~n8034 & n8445;
  assign po1038 = pi57 | ~n6294;
  assign n8448 = pi433 & ~pi451;
  assign n8449 = ~pi433 & pi451;
  assign n8450 = ~n8448 & ~n8449;
  assign n8451 = pi449 & n8450;
  assign n8452 = ~pi449 & ~n8450;
  assign n8453 = ~n8451 & ~n8452;
  assign n8454 = pi448 & ~n8453;
  assign n8455 = ~pi448 & n8453;
  assign n8456 = ~n8454 & ~n8455;
  assign n8457 = ~pi417 & ~pi418;
  assign n8458 = pi417 & pi418;
  assign n8459 = ~n8457 & ~n8458;
  assign n8460 = pi437 & n8459;
  assign n8461 = ~pi437 & ~n8459;
  assign n8462 = ~n8460 & ~n8461;
  assign n8463 = pi453 & ~pi464;
  assign n8464 = ~pi453 & pi464;
  assign n8465 = ~n8463 & ~n8464;
  assign n8466 = n8462 & n8465;
  assign n8467 = ~n8462 & ~n8465;
  assign n8468 = ~n8466 & ~n8467;
  assign n8469 = pi415 & ~pi431;
  assign n8470 = ~pi415 & pi431;
  assign n8471 = ~n8469 & ~n8470;
  assign n8472 = pi416 & ~pi438;
  assign n8473 = ~pi416 & pi438;
  assign n8474 = ~n8472 & ~n8473;
  assign n8475 = n8471 & n8474;
  assign n8476 = ~n8471 & ~n8474;
  assign n8477 = ~n8475 & ~n8476;
  assign n8478 = n8468 & ~n8477;
  assign n8479 = ~n8468 & n8477;
  assign n8480 = pi1197 & ~n8478;
  assign n8481 = ~n8479 & n8480;
  assign n8482 = pi421 & ~pi454;
  assign n8483 = ~pi421 & pi454;
  assign n8484 = ~n8482 & ~n8483;
  assign n8485 = pi432 & ~pi459;
  assign n8486 = ~pi432 & pi459;
  assign n8487 = ~n8485 & ~n8486;
  assign n8488 = n8484 & ~n8487;
  assign n8489 = ~n8484 & n8487;
  assign n8490 = ~n8488 & ~n8489;
  assign n8491 = ~pi419 & ~pi420;
  assign n8492 = pi419 & pi420;
  assign n8493 = ~n8491 & ~n8492;
  assign n8494 = pi423 & ~pi424;
  assign n8495 = ~pi423 & pi424;
  assign n8496 = ~n8494 & ~n8495;
  assign n8497 = n8493 & ~n8496;
  assign n8498 = ~n8493 & n8496;
  assign n8499 = ~n8497 & ~n8498;
  assign n8500 = n8490 & n8499;
  assign n8501 = ~n8490 & ~n8499;
  assign n8502 = ~n8500 & ~n8501;
  assign n8503 = pi425 & ~n8502;
  assign n8504 = ~pi425 & n8502;
  assign n8505 = pi1198 & ~n8503;
  assign n8506 = ~n8504 & n8505;
  assign n8507 = ~n8481 & ~n8506;
  assign n8508 = n7645 & ~n8507;
  assign n8509 = ~pi443 & ~pi592;
  assign n8510 = ~n7571 & ~n8509;
  assign n8511 = ~n7607 & n8509;
  assign n8512 = ~n8510 & ~n8511;
  assign n8513 = ~pi444 & ~n8512;
  assign n8514 = pi443 & ~pi592;
  assign n8515 = ~n7571 & ~n8514;
  assign n8516 = ~n7607 & n8514;
  assign n8517 = ~n8515 & ~n8516;
  assign n8518 = pi444 & ~n8517;
  assign n8519 = ~n8513 & ~n8518;
  assign n8520 = ~pi436 & ~n8519;
  assign n8521 = ~pi429 & ~pi435;
  assign n8522 = pi429 & pi435;
  assign n8523 = ~n8521 & ~n8522;
  assign n8524 = pi434 & ~pi446;
  assign n8525 = ~pi434 & pi446;
  assign n8526 = ~n8524 & ~n8525;
  assign n8527 = pi414 & ~pi422;
  assign n8528 = ~pi414 & pi422;
  assign n8529 = ~n8527 & ~n8528;
  assign n8530 = n8526 & n8529;
  assign n8531 = ~n8526 & ~n8529;
  assign n8532 = ~n8530 & ~n8531;
  assign n8533 = n8523 & n8532;
  assign n8534 = ~n8523 & ~n8532;
  assign n8535 = ~n8533 & ~n8534;
  assign n8536 = ~pi444 & ~n8517;
  assign n8537 = pi444 & ~n8512;
  assign n8538 = ~n8536 & ~n8537;
  assign n8539 = pi436 & ~n8538;
  assign n8540 = ~n8520 & n8535;
  assign n8541 = ~n8539 & n8540;
  assign n8542 = ~pi436 & ~n8538;
  assign n8543 = pi436 & ~n8519;
  assign n8544 = ~n8535 & ~n8542;
  assign n8545 = ~n8543 & n8544;
  assign n8546 = pi1196 & ~n8541;
  assign n8547 = ~n8545 & n8546;
  assign n8548 = ~n7677 & n8507;
  assign n8549 = ~n8547 & n8548;
  assign n8550 = ~n8508 & ~n8549;
  assign n8551 = pi428 & ~n8550;
  assign n8552 = ~pi428 & n7645;
  assign n8553 = ~n8551 & ~n8552;
  assign n8554 = ~pi427 & ~n8553;
  assign n8555 = ~pi428 & ~n8550;
  assign n8556 = pi428 & n7645;
  assign n8557 = ~n8555 & ~n8556;
  assign n8558 = pi427 & ~n8557;
  assign n8559 = ~n8554 & ~n8558;
  assign n8560 = pi430 & ~n8559;
  assign n8561 = ~pi427 & ~n8557;
  assign n8562 = pi427 & ~n8553;
  assign n8563 = ~n8561 & ~n8562;
  assign n8564 = ~pi430 & ~n8563;
  assign n8565 = ~n8560 & ~n8564;
  assign n8566 = pi426 & ~n8565;
  assign n8567 = pi430 & ~n8563;
  assign n8568 = ~pi430 & ~n8559;
  assign n8569 = ~n8567 & ~n8568;
  assign n8570 = ~pi426 & ~n8569;
  assign n8571 = ~n8566 & ~n8570;
  assign n8572 = pi445 & ~n8571;
  assign n8573 = pi426 & ~n8569;
  assign n8574 = ~pi426 & ~n8565;
  assign n8575 = ~n8573 & ~n8574;
  assign n8576 = ~pi445 & ~n8575;
  assign n8577 = ~n8572 & ~n8576;
  assign n8578 = ~n8456 & ~n8577;
  assign n8579 = pi445 & ~n8575;
  assign n8580 = ~pi445 & ~n8571;
  assign n8581 = ~n8579 & ~n8580;
  assign n8582 = n8456 & ~n8581;
  assign n8583 = pi1199 & ~n8578;
  assign n8584 = ~n8582 & n8583;
  assign n8585 = ~pi590 & ~pi591;
  assign n8586 = ~pi1199 & n8550;
  assign n8587 = n8585 & ~n8586;
  assign n8588 = ~n8584 & n8587;
  assign n8589 = n7571 & ~n8585;
  assign n8590 = n7720 & ~n8589;
  assign n8591 = ~n8588 & n8590;
  assign n8592 = n8114 & ~n8509;
  assign n8593 = ~pi436 & pi444;
  assign n8594 = pi436 & ~pi444;
  assign n8595 = ~n8593 & ~n8594;
  assign n8596 = n8535 & ~n8595;
  assign n8597 = ~n8535 & n8595;
  assign n8598 = ~n8596 & ~n8597;
  assign n8599 = ~n8511 & n8598;
  assign n8600 = ~n8592 & n8599;
  assign n8601 = n8114 & ~n8514;
  assign n8602 = ~n8516 & ~n8598;
  assign n8603 = ~n8601 & n8602;
  assign n8604 = pi1196 & ~n8600;
  assign n8605 = ~n8603 & n8604;
  assign n8606 = ~n8137 & ~n8605;
  assign n8607 = n8507 & ~n8606;
  assign n8608 = ~n8116 & ~n8507;
  assign n8609 = ~n8607 & ~n8608;
  assign n8610 = pi428 & n8609;
  assign n8611 = ~pi428 & n8116;
  assign n8612 = pi427 & ~n8611;
  assign n8613 = ~n8610 & n8612;
  assign n8614 = ~pi428 & n8609;
  assign n8615 = pi428 & n8116;
  assign n8616 = ~pi427 & ~n8615;
  assign n8617 = ~n8614 & n8616;
  assign n8618 = ~n8613 & ~n8617;
  assign n8619 = ~pi430 & ~n8618;
  assign n8620 = ~pi427 & pi428;
  assign n8621 = pi427 & ~pi428;
  assign n8622 = ~n8620 & ~n8621;
  assign n8623 = n8116 & n8622;
  assign n8624 = n8609 & ~n8622;
  assign n8625 = ~n8623 & ~n8624;
  assign n8626 = pi430 & n8625;
  assign n8627 = ~n8619 & ~n8626;
  assign n8628 = ~pi426 & ~n8627;
  assign n8629 = pi430 & ~n8618;
  assign n8630 = ~pi430 & n8625;
  assign n8631 = ~n8629 & ~n8630;
  assign n8632 = pi426 & ~n8631;
  assign n8633 = ~n8628 & ~n8632;
  assign n8634 = ~pi445 & ~n8633;
  assign n8635 = ~pi426 & ~n8631;
  assign n8636 = pi426 & ~n8627;
  assign n8637 = ~n8635 & ~n8636;
  assign n8638 = pi445 & ~n8637;
  assign n8639 = ~n8634 & ~n8638;
  assign n8640 = pi448 & n8639;
  assign n8641 = ~pi445 & ~n8637;
  assign n8642 = pi445 & ~n8633;
  assign n8643 = ~n8641 & ~n8642;
  assign n8644 = ~pi448 & n8643;
  assign n8645 = ~n8453 & ~n8640;
  assign n8646 = ~n8644 & n8645;
  assign n8647 = ~pi448 & n8639;
  assign n8648 = pi448 & n8643;
  assign n8649 = n8453 & ~n8647;
  assign n8650 = ~n8648 & n8649;
  assign n8651 = ~n8646 & ~n8650;
  assign n8652 = pi1199 & ~n8651;
  assign n8653 = ~pi1199 & ~n8609;
  assign n8654 = n8585 & ~n8653;
  assign n8655 = ~n8652 & n8654;
  assign n8656 = ~n8114 & ~n8585;
  assign n8657 = ~n7720 & ~n8656;
  assign n8658 = ~n8655 & n8657;
  assign n8659 = ~n8591 & ~n8658;
  assign n8660 = pi588 & ~n8659;
  assign n8661 = ~po1038 & ~n8660;
  assign n8662 = ~n8446 & n8661;
  assign n8663 = ~pi592 & n7639;
  assign n8664 = ~n7627 & n8112;
  assign n8665 = ~n8663 & n8664;
  assign n8666 = pi361 & ~pi458;
  assign n8667 = ~pi361 & pi458;
  assign n8668 = ~n8666 & ~n8667;
  assign n8669 = n7621 & n8668;
  assign n8670 = ~n7621 & ~n8668;
  assign n8671 = ~n8669 & ~n8670;
  assign n8672 = ~pi441 & n8671;
  assign n8673 = pi441 & ~n8671;
  assign n8674 = ~pi592 & ~n8672;
  assign n8675 = ~n8673 & n8674;
  assign n8676 = n7627 & n8112;
  assign n8677 = ~n8675 & n8676;
  assign n8678 = pi1196 & ~n8677;
  assign n8679 = ~n8665 & n8678;
  assign n8680 = ~pi1198 & ~n8679;
  assign n8681 = pi350 & ~n7594;
  assign n8682 = ~pi350 & n7594;
  assign n8683 = ~n8681 & ~n8682;
  assign n8684 = ~n7640 & n8683;
  assign n8685 = ~pi592 & n8112;
  assign n8686 = pi1198 & n8685;
  assign n8687 = n8684 & n8686;
  assign n8688 = ~n8680 & ~n8687;
  assign n8689 = ~n7443 & ~n8688;
  assign n8690 = ~pi592 & ~n8689;
  assign n8691 = n8112 & ~n8690;
  assign n8692 = ~n7690 & ~n8691;
  assign n8693 = pi592 & n8112;
  assign n8694 = pi1199 & ~n8693;
  assign n8695 = pi351 & n8694;
  assign n8696 = ~n8692 & ~n8695;
  assign n8697 = ~pi461 & ~n8696;
  assign n8698 = ~n7684 & ~n8691;
  assign n8699 = ~pi351 & n8694;
  assign n8700 = ~n8698 & ~n8699;
  assign n8701 = pi461 & ~n8700;
  assign n8702 = ~n8697 & ~n8701;
  assign n8703 = ~pi357 & ~n8702;
  assign n8704 = ~pi461 & ~n8700;
  assign n8705 = pi461 & ~n8696;
  assign n8706 = ~n8704 & ~n8705;
  assign n8707 = pi357 & ~n8706;
  assign n8708 = ~n8703 & ~n8707;
  assign n8709 = ~pi356 & ~n8708;
  assign n8710 = ~pi357 & ~n8706;
  assign n8711 = pi357 & ~n8702;
  assign n8712 = ~n8710 & ~n8711;
  assign n8713 = pi356 & ~n8712;
  assign n8714 = n7418 & ~n8709;
  assign n8715 = ~n8713 & n8714;
  assign n8716 = ~pi356 & ~n8712;
  assign n8717 = pi356 & ~n8708;
  assign n8718 = ~n7418 & ~n8716;
  assign n8719 = ~n8717 & n8718;
  assign n8720 = ~n8715 & ~n8719;
  assign n8721 = pi590 & ~n8720;
  assign n8722 = ~pi377 & ~n7794;
  assign n8723 = pi377 & n7794;
  assign n8724 = ~n8722 & ~n8723;
  assign n8725 = n7771 & ~n8724;
  assign n8726 = pi592 & ~n8725;
  assign n8727 = n8112 & ~n8726;
  assign n8728 = pi1199 & ~n8727;
  assign n8729 = n7771 & n8693;
  assign n8730 = ~n8728 & n8729;
  assign n8731 = ~pi1198 & n8730;
  assign n8732 = ~pi369 & ~pi374;
  assign n8733 = pi369 & pi374;
  assign n8734 = ~n8732 & ~n8733;
  assign n8735 = ~pi370 & ~n8734;
  assign n8736 = pi370 & n8734;
  assign n8737 = ~n8735 & ~n8736;
  assign n8738 = ~pi371 & ~n8737;
  assign n8739 = pi371 & n8737;
  assign n8740 = ~n8738 & ~n8739;
  assign n8741 = ~pi373 & ~n8740;
  assign n8742 = pi373 & n8740;
  assign n8743 = ~n8741 & ~n8742;
  assign n8744 = pi375 & ~n8743;
  assign n8745 = ~pi375 & n8743;
  assign n8746 = ~n8744 & ~n8745;
  assign n8747 = ~n7862 & ~n8746;
  assign n8748 = n7862 & n8746;
  assign n8749 = ~n8747 & ~n8748;
  assign n8750 = n8730 & n8749;
  assign n8751 = ~n8685 & ~n8731;
  assign n8752 = ~n8750 & n8751;
  assign n8753 = ~pi590 & ~n8752;
  assign n8754 = ~pi591 & ~n8753;
  assign n8755 = ~n8721 & n8754;
  assign n8756 = pi1197 & ~n8693;
  assign n8757 = ~pi592 & ~n7964;
  assign n8758 = n8338 & n8757;
  assign n8759 = n8694 & ~n8758;
  assign n8760 = n8242 & n8245;
  assign n8761 = n8112 & ~n8242;
  assign n8762 = ~pi1199 & ~n8761;
  assign n8763 = ~n8760 & n8762;
  assign n8764 = ~n8759 & ~n8763;
  assign n8765 = ~pi1197 & ~n8764;
  assign n8766 = ~n8756 & ~n8765;
  assign n8767 = pi333 & ~n8766;
  assign n8768 = pi1198 & ~n8693;
  assign n8769 = n8764 & ~n8768;
  assign n8770 = ~n7899 & ~n8769;
  assign n8771 = ~pi333 & ~n8764;
  assign n8772 = ~n8770 & ~n8771;
  assign n8773 = ~n8767 & n8772;
  assign n8774 = ~pi391 & ~n8773;
  assign n8775 = ~pi333 & ~n8766;
  assign n8776 = n8764 & ~n8770;
  assign n8777 = ~n8775 & n8776;
  assign n8778 = pi391 & ~n8777;
  assign n8779 = ~n8774 & ~n8778;
  assign n8780 = ~pi392 & ~n8779;
  assign n8781 = ~pi391 & ~n8777;
  assign n8782 = pi391 & ~n8773;
  assign n8783 = ~n8781 & ~n8782;
  assign n8784 = pi392 & ~n8783;
  assign n8785 = ~n8780 & ~n8784;
  assign n8786 = ~pi393 & ~n8785;
  assign n8787 = ~pi392 & ~n8783;
  assign n8788 = pi392 & ~n8779;
  assign n8789 = ~n8787 & ~n8788;
  assign n8790 = pi393 & ~n8789;
  assign n8791 = n8238 & ~n8786;
  assign n8792 = ~n8790 & n8791;
  assign n8793 = ~pi393 & ~n8789;
  assign n8794 = pi393 & ~n8785;
  assign n8795 = ~n8238 & ~n8793;
  assign n8796 = ~n8794 & n8795;
  assign n8797 = ~n8792 & ~n8796;
  assign n8798 = ~pi590 & ~n8797;
  assign n8799 = pi590 & n8112;
  assign n8800 = pi591 & ~n8799;
  assign n8801 = ~n8798 & n8800;
  assign n8802 = ~n8755 & ~n8801;
  assign n8803 = ~pi588 & ~n8802;
  assign n8804 = ~n7720 & po1038;
  assign n8805 = pi436 & ~pi443;
  assign n8806 = ~pi436 & pi443;
  assign n8807 = ~n8805 & ~n8806;
  assign n8808 = ~pi444 & n8807;
  assign n8809 = pi444 & ~n8807;
  assign n8810 = ~n8808 & ~n8809;
  assign n8811 = ~n8535 & ~n8810;
  assign n8812 = n8535 & n8810;
  assign n8813 = n8242 & ~n8811;
  assign n8814 = ~n8812 & n8813;
  assign n8815 = n8507 & ~n8814;
  assign n8816 = n8685 & n8815;
  assign n8817 = pi430 & ~n8622;
  assign n8818 = ~pi430 & n8622;
  assign n8819 = ~n8817 & ~n8818;
  assign n8820 = ~pi426 & ~n8819;
  assign n8821 = pi426 & n8819;
  assign n8822 = ~n8820 & ~n8821;
  assign n8823 = ~pi445 & ~n8822;
  assign n8824 = pi445 & n8822;
  assign n8825 = ~n8823 & ~n8824;
  assign n8826 = ~pi448 & ~n8825;
  assign n8827 = pi448 & n8825;
  assign n8828 = ~n8826 & ~n8827;
  assign n8829 = n8816 & ~n8828;
  assign n8830 = ~n8693 & ~n8829;
  assign n8831 = n8453 & ~n8830;
  assign n8832 = n8816 & n8828;
  assign n8833 = ~n8693 & ~n8832;
  assign n8834 = ~n8453 & ~n8833;
  assign n8835 = pi1199 & ~n8831;
  assign n8836 = ~n8834 & n8835;
  assign n8837 = ~pi1199 & ~n8693;
  assign n8838 = ~n8816 & n8837;
  assign n8839 = n8585 & ~n8838;
  assign n8840 = ~n8836 & n8839;
  assign n8841 = n8112 & ~n8585;
  assign n8842 = pi588 & ~n8841;
  assign n8843 = ~n8840 & n8842;
  assign n8844 = n8804 & ~n8843;
  assign n8845 = ~n8803 & n8844;
  assign n8846 = ~pi217 & ~n8845;
  assign n8847 = ~n8662 & n8846;
  assign n8848 = ~n7571 & n7720;
  assign n8849 = ~n7720 & n8114;
  assign n8850 = ~po1038 & ~n8849;
  assign n8851 = ~n8848 & n8850;
  assign n8852 = n8112 & n8804;
  assign n8853 = pi217 & ~n8852;
  assign n8854 = ~n8851 & n8853;
  assign n8855 = ~pi1161 & ~pi1162;
  assign n8856 = ~pi1163 & n8855;
  assign n8857 = ~n8854 & n8856;
  assign n8858 = ~n8847 & n8857;
  assign n8859 = pi1161 & ~pi1163;
  assign n8860 = n2755 & n8859;
  assign n8861 = ~pi31 & pi1162;
  assign n8862 = n8860 & n8861;
  assign po189 = n8858 | n8862;
  assign n8864 = n3294 & n3432;
  assign n8865 = ~pi55 & ~pi74;
  assign n8866 = n8864 & n8865;
  assign n8867 = n6279 & n8866;
  assign n8868 = pi100 & n3182;
  assign n8869 = n6248 & ~po1057;
  assign n8870 = n6492 & n8869;
  assign n8871 = ~pi137 & n8870;
  assign n8872 = pi129 & n3096;
  assign n8873 = ~pi137 & pi252;
  assign n8874 = po1057 & ~n7485;
  assign n8875 = ~n6248 & ~n8874;
  assign n8876 = n8873 & n8875;
  assign n8877 = n8872 & n8876;
  assign n8878 = ~n8871 & ~n8877;
  assign n8879 = n8868 & ~n8878;
  assign n8880 = ~pi24 & ~pi90;
  assign n8881 = n6153 & n8880;
  assign n8882 = pi50 & n2586;
  assign n8883 = n2482 & n8882;
  assign n8884 = n2484 & n2510;
  assign n8885 = n2490 & n8884;
  assign n8886 = ~pi93 & n8885;
  assign n8887 = n8883 & n8886;
  assign n8888 = n8881 & n8887;
  assign n8889 = pi829 & ~pi1093;
  assign n8890 = n6265 & n8889;
  assign po840 = n2796 | n8890;
  assign n8892 = ~n7720 & ~po840;
  assign n8893 = ~pi137 & ~n8892;
  assign n8894 = n8888 & ~n8893;
  assign n8895 = ~pi68 & ~pi73;
  assign n8896 = ~pi49 & ~pi66;
  assign n8897 = ~pi89 & ~pi102;
  assign n8898 = n7451 & n8897;
  assign n8899 = ~pi64 & ~pi81;
  assign n8900 = n2476 & n8899;
  assign n8901 = n2451 & n2641;
  assign n8902 = ~pi103 & n2460;
  assign n8903 = n8901 & n8902;
  assign n8904 = n2455 & n2606;
  assign n8905 = ~pi45 & ~pi48;
  assign n8906 = ~pi61 & ~pi104;
  assign n8907 = n8905 & n8906;
  assign n8908 = n8904 & n8907;
  assign n8909 = pi76 & ~pi84;
  assign n8910 = n2468 & n8909;
  assign n8911 = n8895 & n8896;
  assign n8912 = n8910 & n8911;
  assign n8913 = n8898 & n8900;
  assign n8914 = n8912 & n8913;
  assign n8915 = n8903 & n8908;
  assign n8916 = n8914 & n8915;
  assign n8917 = ~n8882 & ~n8916;
  assign n8918 = n2486 & n2491;
  assign n8919 = ~n8917 & n8918;
  assign n8920 = ~pi24 & ~n8919;
  assign n8921 = n2482 & n8916;
  assign n8922 = n8885 & n8921;
  assign n8923 = pi24 & ~n8922;
  assign n8924 = n2550 & n2783;
  assign n8925 = ~pi137 & n7459;
  assign n8926 = n8924 & n8925;
  assign n8927 = ~n8892 & n8926;
  assign n8928 = ~n8923 & n8927;
  assign n8929 = ~n8920 & n8928;
  assign n8930 = ~n8894 & ~n8929;
  assign n8931 = ~pi32 & ~n8930;
  assign n8932 = ~pi24 & ~pi841;
  assign n8933 = pi32 & ~n8932;
  assign n8934 = n2499 & n8933;
  assign n8935 = ~n8931 & ~n8934;
  assign n8936 = ~n6151 & ~n8935;
  assign n8937 = ~pi32 & ~n8888;
  assign n8938 = n6151 & ~n6155;
  assign n8939 = ~n8937 & n8938;
  assign n8940 = ~n8936 & ~n8939;
  assign n8941 = ~pi95 & n3277;
  assign n8942 = ~n8940 & n8941;
  assign n8943 = ~n8879 & ~n8942;
  assign n8944 = n3231 & ~n8943;
  assign n8945 = ~pi24 & n2548;
  assign n8946 = n2494 & n3094;
  assign n8947 = ~pi51 & n8946;
  assign n8948 = n8945 & n8947;
  assign n8949 = ~po840 & n8948;
  assign n8950 = pi252 & ~n8874;
  assign n8951 = ~pi87 & n3182;
  assign n8952 = pi75 & ~pi100;
  assign n8953 = n8951 & n8952;
  assign n8954 = ~pi137 & n8953;
  assign n8955 = ~n6271 & n8954;
  assign n8956 = ~n8950 & n8955;
  assign n8957 = n8949 & n8956;
  assign n8958 = ~n8944 & ~n8957;
  assign po190 = n8867 & ~n8958;
  assign n8960 = ~pi195 & ~pi196;
  assign n8961 = ~pi138 & n8960;
  assign n8962 = ~pi139 & n8961;
  assign n8963 = ~pi118 & n8962;
  assign n8964 = ~pi79 & n8963;
  assign n8965 = ~pi34 & n8964;
  assign n8966 = ~pi33 & ~n8965;
  assign n8967 = pi149 & pi157;
  assign n8968 = ~pi149 & ~pi157;
  assign n8969 = n6170 & ~n8968;
  assign n8970 = ~n8967 & n8969;
  assign n8971 = pi232 & n8970;
  assign n8972 = pi75 & ~n8971;
  assign n8973 = pi100 & ~n8971;
  assign n8974 = ~n8972 & ~n8973;
  assign n8975 = ~pi75 & ~pi100;
  assign n8976 = n7484 & n8975;
  assign n8977 = pi164 & n8976;
  assign n8978 = n8974 & ~n8977;
  assign n8979 = ~pi74 & ~n8978;
  assign n8980 = pi169 & n8976;
  assign n8981 = n8974 & ~n8980;
  assign n8982 = pi74 & ~n8981;
  assign n8983 = ~n3432 & ~n8979;
  assign n8984 = ~n8982 & n8983;
  assign n8985 = pi299 & ~n8970;
  assign n8986 = pi178 & pi183;
  assign n8987 = ~pi178 & ~pi183;
  assign n8988 = n6170 & ~n8987;
  assign n8989 = ~n8986 & n8988;
  assign n8990 = ~pi299 & ~n8989;
  assign n8991 = pi232 & ~n8985;
  assign n8992 = ~n8990 & n8991;
  assign n8993 = pi100 & ~n8992;
  assign n8994 = pi75 & ~n8992;
  assign n8995 = ~n8993 & ~n8994;
  assign n8996 = pi191 & ~pi299;
  assign n8997 = pi169 & pi299;
  assign n8998 = ~n8996 & ~n8997;
  assign n8999 = n8976 & ~n8998;
  assign n9000 = n8995 & ~n8999;
  assign n9001 = pi74 & ~n9000;
  assign n9002 = ~pi55 & ~n9001;
  assign n9003 = ~pi186 & ~pi299;
  assign n9004 = ~pi164 & pi299;
  assign n9005 = ~n9003 & ~n9004;
  assign n9006 = n7484 & n9005;
  assign n9007 = n8975 & n9006;
  assign n9008 = n8995 & ~n9007;
  assign n9009 = pi54 & ~n9008;
  assign n9010 = pi299 & n7484;
  assign n9011 = ~n6117 & n9010;
  assign n9012 = ~pi186 & ~n9011;
  assign n9013 = ~n6250 & n7484;
  assign n9014 = pi186 & ~n9013;
  assign n9015 = pi164 & ~n9014;
  assign n9016 = ~n9012 & n9015;
  assign n9017 = ~pi299 & n7484;
  assign n9018 = ~n6117 & n9017;
  assign n9019 = ~pi164 & pi186;
  assign n9020 = n9018 & n9019;
  assign n9021 = ~n9016 & ~n9020;
  assign n9022 = pi38 & ~n9021;
  assign n9023 = ~pi176 & pi232;
  assign n9024 = ~pi40 & n2476;
  assign n9025 = ~pi102 & n8899;
  assign n9026 = n2455 & n9025;
  assign n9027 = n2453 & n9026;
  assign n9028 = n2474 & n9027;
  assign n9029 = ~pi60 & n9028;
  assign n9030 = n2505 & n2513;
  assign n9031 = ~pi53 & n9030;
  assign n9032 = n9029 & n9031;
  assign n9033 = ~pi58 & n9032;
  assign n9034 = n7459 & n9033;
  assign n9035 = ~pi32 & n2551;
  assign n9036 = n9034 & n9035;
  assign n9037 = ~pi95 & n9036;
  assign n9038 = n6446 & ~n6458;
  assign n9039 = n6178 & n9038;
  assign n9040 = ~n6209 & ~n9039;
  assign n9041 = n9037 & ~n9040;
  assign n9042 = n6206 & n9041;
  assign n9043 = n9024 & ~n9042;
  assign n9044 = pi224 & n6469;
  assign n9045 = n9024 & ~n9044;
  assign n9046 = ~n9043 & ~n9045;
  assign n9047 = n9037 & n9039;
  assign n9048 = n6170 & n9047;
  assign n9049 = n9024 & ~n9048;
  assign n9050 = ~n6197 & ~n9049;
  assign n9051 = ~n9045 & n9050;
  assign n9052 = pi174 & n9051;
  assign n9053 = ~n9046 & ~n9052;
  assign n9054 = ~pi299 & ~n9053;
  assign n9055 = pi216 & n6442;
  assign n9056 = n9024 & ~n9055;
  assign n9057 = pi299 & ~n9056;
  assign n9058 = n6170 & n9041;
  assign n9059 = n9024 & ~n9058;
  assign n9060 = ~n6223 & ~n9059;
  assign n9061 = n9043 & ~n9060;
  assign n9062 = n6209 & n9037;
  assign n9063 = ~n6200 & n9062;
  assign n9064 = n9024 & ~n9063;
  assign n9065 = n6170 & n9064;
  assign n9066 = ~pi152 & n9065;
  assign n9067 = ~pi154 & ~n9061;
  assign n9068 = ~n9066 & n9067;
  assign n9069 = n9024 & ~n9047;
  assign n9070 = n6228 & ~n9069;
  assign n9071 = pi152 & n9070;
  assign n9072 = n9043 & ~n9071;
  assign n9073 = pi154 & ~n9072;
  assign n9074 = n9055 & ~n9073;
  assign n9075 = ~n9068 & n9074;
  assign n9076 = n9057 & ~n9075;
  assign n9077 = ~n9054 & ~n9076;
  assign n9078 = n6207 & n9062;
  assign n9079 = n9024 & n9044;
  assign n9080 = ~n9078 & n9079;
  assign n9081 = ~n9045 & ~n9080;
  assign n9082 = ~pi299 & n9081;
  assign n9083 = n9077 & ~n9082;
  assign n9084 = n9023 & ~n9083;
  assign n9085 = pi176 & pi232;
  assign n9086 = ~n9077 & n9085;
  assign n9087 = n9057 & ~n9061;
  assign n9088 = ~n6197 & ~n9059;
  assign n9089 = ~n9045 & n9088;
  assign n9090 = ~n9046 & ~n9089;
  assign n9091 = ~pi299 & ~n9090;
  assign n9092 = ~n9087 & ~n9091;
  assign n9093 = ~pi232 & ~n9092;
  assign n9094 = pi39 & ~n9093;
  assign n9095 = ~n9086 & n9094;
  assign n9096 = ~n9084 & n9095;
  assign n9097 = pi95 & ~n9024;
  assign n9098 = ~n2449 & ~n9097;
  assign n9099 = ~pi40 & ~pi479;
  assign n9100 = n2476 & ~n9036;
  assign n9101 = n9099 & n9100;
  assign n9102 = ~n9098 & ~n9101;
  assign n9103 = pi32 & ~n9024;
  assign n9104 = n2476 & ~n2549;
  assign n9105 = n2476 & ~n9034;
  assign n9106 = pi70 & ~n9105;
  assign n9107 = n2476 & ~n9032;
  assign n9108 = pi58 & ~n9107;
  assign n9109 = pi53 & ~n9029;
  assign n9110 = ~pi60 & n8882;
  assign n9111 = n2504 & ~n9110;
  assign n9112 = ~n9109 & ~n9111;
  assign n9113 = ~pi68 & n2457;
  assign n9114 = ~pi111 & n2456;
  assign n9115 = ~pi36 & n9113;
  assign n9116 = n9114 & n9115;
  assign n9117 = ~pi66 & ~pi84;
  assign n9118 = pi73 & ~pi82;
  assign n9119 = n9117 & n9118;
  assign n9120 = n9027 & n9119;
  assign n9121 = n9116 & n9120;
  assign n9122 = n2466 & n9121;
  assign n9123 = n2481 & n9122;
  assign n9124 = n2476 & ~n9123;
  assign n9125 = ~n9112 & n9124;
  assign n9126 = n2505 & ~n9125;
  assign n9127 = ~n2476 & ~n2505;
  assign n9128 = n2513 & ~n9127;
  assign n9129 = ~n9126 & n9128;
  assign n9130 = n2476 & ~n2513;
  assign n9131 = ~pi58 & ~n9130;
  assign n9132 = ~n9129 & n9131;
  assign n9133 = ~n9108 & ~n9132;
  assign n9134 = ~pi90 & ~n9133;
  assign n9135 = ~pi841 & n9033;
  assign n9136 = n2476 & ~n9135;
  assign n9137 = pi90 & ~n9136;
  assign n9138 = n2547 & ~n9137;
  assign n9139 = ~n9134 & n9138;
  assign n9140 = n2476 & ~n2547;
  assign n9141 = ~pi70 & ~n9140;
  assign n9142 = ~n9139 & n9141;
  assign n9143 = ~n9106 & ~n9142;
  assign n9144 = ~pi51 & ~n9143;
  assign n9145 = pi51 & ~n2476;
  assign n9146 = n2549 & ~n9145;
  assign n9147 = ~n9144 & n9146;
  assign n9148 = ~n9104 & ~n9147;
  assign n9149 = ~pi40 & ~n9148;
  assign n9150 = ~pi32 & ~n9149;
  assign n9151 = ~n9103 & ~n9150;
  assign n9152 = ~pi95 & ~n9151;
  assign n9153 = ~n9102 & ~n9152;
  assign n9154 = n2493 & n6152;
  assign n9155 = n9135 & n9154;
  assign n9156 = n9024 & ~n9155;
  assign n9157 = pi32 & ~n9156;
  assign n9158 = ~n9150 & ~n9157;
  assign n9159 = ~pi95 & ~n9158;
  assign n9160 = ~pi198 & n9159;
  assign n9161 = n9153 & ~n9160;
  assign n9162 = ~n6170 & n9161;
  assign n9163 = n9030 & n9112;
  assign n9164 = n2476 & ~n9163;
  assign n9165 = ~pi58 & ~n9164;
  assign n9166 = ~n9108 & ~n9165;
  assign n9167 = ~pi90 & ~n9166;
  assign n9168 = n9138 & ~n9167;
  assign n9169 = n9141 & ~n9168;
  assign n9170 = ~n9106 & ~n9169;
  assign n9171 = ~pi51 & ~n9170;
  assign n9172 = n9146 & ~n9171;
  assign n9173 = ~n9104 & ~n9172;
  assign n9174 = ~pi40 & ~n9173;
  assign n9175 = ~pi32 & ~n9174;
  assign n9176 = ~n9157 & ~n9175;
  assign n9177 = ~pi95 & ~n9176;
  assign n9178 = ~pi198 & n9177;
  assign n9179 = n6170 & ~n9097;
  assign n9180 = ~n9103 & ~n9175;
  assign n9181 = ~pi95 & ~n9180;
  assign n9182 = n9179 & ~n9181;
  assign n9183 = ~n9178 & n9182;
  assign n9184 = ~n9162 & ~n9183;
  assign n9185 = ~pi183 & ~n9184;
  assign n9186 = ~pi40 & ~n9103;
  assign n9187 = n2476 & ~n6152;
  assign n9188 = ~pi32 & ~n9187;
  assign n9189 = pi93 & ~n2476;
  assign n9190 = n6152 & ~n9189;
  assign n9191 = n2476 & ~n9108;
  assign n9192 = ~pi90 & ~n9191;
  assign n9193 = ~n9137 & ~n9192;
  assign n9194 = ~pi93 & ~n9193;
  assign n9195 = n9190 & ~n9194;
  assign n9196 = n9188 & ~n9195;
  assign n9197 = n9186 & ~n9196;
  assign n9198 = ~pi95 & ~n9197;
  assign n9199 = n9179 & ~n9198;
  assign n9200 = ~n9162 & ~n9199;
  assign n9201 = pi183 & ~n9200;
  assign n9202 = ~n9185 & ~n9201;
  assign n9203 = ~pi95 & n9202;
  assign n9204 = ~pi174 & ~n9102;
  assign n9205 = ~n9203 & n9204;
  assign n9206 = pi183 & n6170;
  assign n9207 = ~n9161 & ~n9206;
  assign n9208 = n8918 & n9122;
  assign n9209 = ~pi90 & n9208;
  assign n9210 = n9193 & ~n9209;
  assign n9211 = ~pi93 & ~n9210;
  assign n9212 = n9190 & ~n9211;
  assign n9213 = n9188 & ~n9212;
  assign n9214 = n9186 & ~n9213;
  assign n9215 = ~pi95 & ~n9214;
  assign n9216 = ~n9102 & ~n9215;
  assign n9217 = n6170 & ~n9216;
  assign n9218 = pi183 & n9217;
  assign n9219 = pi174 & ~n9218;
  assign n9220 = ~n9207 & n9219;
  assign n9221 = ~pi180 & ~n9220;
  assign n9222 = ~n9205 & n9221;
  assign n9223 = ~pi174 & ~n9202;
  assign n9224 = n9179 & ~n9215;
  assign n9225 = ~n9162 & ~n9224;
  assign n9226 = pi183 & ~n9225;
  assign n9227 = ~pi40 & n6170;
  assign n9228 = ~n9097 & ~n9152;
  assign n9229 = ~n9160 & n9228;
  assign n9230 = n9227 & n9229;
  assign n9231 = ~n9162 & ~n9230;
  assign n9232 = ~pi183 & ~n9231;
  assign n9233 = ~n9226 & ~n9232;
  assign n9234 = pi174 & ~n9233;
  assign n9235 = pi180 & ~n9223;
  assign n9236 = ~n9234 & n9235;
  assign n9237 = ~n9222 & ~n9236;
  assign n9238 = ~pi193 & ~n9237;
  assign n9239 = ~pi40 & ~n2476;
  assign n9240 = pi32 & ~n9239;
  assign n9241 = n2518 & n2547;
  assign n9242 = ~n2476 & ~n9241;
  assign n9243 = n7459 & n9132;
  assign n9244 = ~n9242 & ~n9243;
  assign n9245 = ~pi70 & ~n9244;
  assign n9246 = ~n9106 & ~n9245;
  assign n9247 = ~pi51 & ~n9246;
  assign n9248 = n9146 & ~n9247;
  assign n9249 = ~pi40 & ~n9104;
  assign n9250 = ~n9248 & n9249;
  assign n9251 = ~pi32 & ~n9250;
  assign n9252 = ~n9240 & ~n9251;
  assign n9253 = ~n2783 & ~n9024;
  assign n9254 = ~n9252 & ~n9253;
  assign n9255 = ~pi95 & ~n9254;
  assign n9256 = ~n9102 & ~n9255;
  assign n9257 = n6170 & ~n9024;
  assign n9258 = ~n9097 & ~n9255;
  assign n9259 = pi95 & ~n9239;
  assign n9260 = ~pi40 & ~n9156;
  assign n9261 = pi32 & ~n9260;
  assign n9262 = ~n9251 & ~n9261;
  assign n9263 = ~pi95 & ~n9262;
  assign n9264 = ~n9259 & ~n9263;
  assign n9265 = n9258 & ~n9264;
  assign n9266 = ~pi198 & ~n9265;
  assign n9267 = n6170 & ~n9266;
  assign n9268 = ~n9257 & ~n9267;
  assign n9269 = n9256 & ~n9268;
  assign n9270 = ~n9162 & ~n9269;
  assign n9271 = ~pi183 & ~n9270;
  assign n9272 = n8918 & n9154;
  assign n9273 = ~pi32 & n9272;
  assign n9274 = n9122 & n9273;
  assign n9275 = n9024 & ~n9274;
  assign n9276 = ~pi95 & ~n9275;
  assign n9277 = n6170 & ~n9276;
  assign n9278 = ~n9102 & n9277;
  assign n9279 = ~n9162 & ~n9278;
  assign n9280 = pi183 & ~n9279;
  assign n9281 = pi174 & ~n9280;
  assign n9282 = ~n9271 & n9281;
  assign n9283 = ~n6170 & ~n9161;
  assign n9284 = n7459 & n9165;
  assign n9285 = ~n9242 & ~n9284;
  assign n9286 = ~pi70 & ~n9285;
  assign n9287 = ~n9106 & ~n9286;
  assign n9288 = ~pi51 & ~n9287;
  assign n9289 = n9146 & ~n9288;
  assign n9290 = ~n9104 & ~n9289;
  assign n9291 = ~pi40 & ~n9290;
  assign n9292 = ~pi32 & ~n9291;
  assign n9293 = ~n9103 & ~n9292;
  assign n9294 = ~pi95 & ~n9293;
  assign n9295 = ~n9102 & ~n9294;
  assign n9296 = ~n9157 & ~n9292;
  assign n9297 = ~pi95 & ~n9296;
  assign n9298 = ~pi198 & n9297;
  assign n9299 = n9295 & ~n9298;
  assign n9300 = n6170 & ~n9299;
  assign n9301 = ~n9283 & ~n9300;
  assign n9302 = ~pi183 & n9301;
  assign n9303 = ~pi95 & ~n9024;
  assign n9304 = ~n9102 & ~n9303;
  assign n9305 = n6170 & n9304;
  assign n9306 = ~n9162 & ~n9305;
  assign n9307 = pi183 & ~n9306;
  assign n9308 = ~pi174 & ~n9302;
  assign n9309 = ~n9307 & n9308;
  assign n9310 = ~pi180 & ~n9309;
  assign n9311 = ~n9282 & n9310;
  assign n9312 = n9258 & n9267;
  assign n9313 = ~n9162 & ~n9312;
  assign n9314 = ~pi183 & ~n9313;
  assign n9315 = n9179 & ~n9276;
  assign n9316 = ~n9162 & ~n9315;
  assign n9317 = pi183 & ~n9316;
  assign n9318 = pi174 & ~n9317;
  assign n9319 = ~n9314 & n9318;
  assign n9320 = ~n9257 & ~n9283;
  assign n9321 = pi183 & n9320;
  assign n9322 = ~pi40 & n9290;
  assign n9323 = ~pi32 & ~n9322;
  assign n9324 = ~n9240 & ~n9323;
  assign n9325 = ~pi95 & ~n9324;
  assign n9326 = ~n9259 & ~n9325;
  assign n9327 = pi198 & ~n9326;
  assign n9328 = ~n9261 & ~n9323;
  assign n9329 = ~pi95 & ~n9328;
  assign n9330 = ~n9259 & ~n9329;
  assign n9331 = ~pi198 & ~n9330;
  assign n9332 = ~n9327 & ~n9331;
  assign n9333 = n9227 & ~n9332;
  assign n9334 = ~n9162 & ~n9333;
  assign n9335 = ~pi183 & ~n9334;
  assign n9336 = ~pi174 & ~n9321;
  assign n9337 = ~n9335 & n9336;
  assign n9338 = pi180 & ~n9319;
  assign n9339 = ~n9337 & n9338;
  assign n9340 = pi193 & ~n9311;
  assign n9341 = ~n9339 & n9340;
  assign n9342 = ~n9238 & ~n9341;
  assign n9343 = ~pi299 & ~n9342;
  assign n9344 = pi158 & pi299;
  assign n9345 = ~pi210 & n9159;
  assign n9346 = n9153 & ~n9345;
  assign n9347 = ~n6170 & n9346;
  assign n9348 = ~pi210 & n9177;
  assign n9349 = n9182 & ~n9348;
  assign n9350 = ~n9347 & ~n9349;
  assign n9351 = ~pi152 & ~n9350;
  assign n9352 = ~n6170 & ~n9346;
  assign n9353 = n9228 & ~n9345;
  assign n9354 = n6170 & ~n9353;
  assign n9355 = ~n9352 & ~n9354;
  assign n9356 = pi152 & n9355;
  assign n9357 = ~pi172 & ~n9351;
  assign n9358 = ~n9356 & n9357;
  assign n9359 = ~pi210 & ~n9265;
  assign n9360 = n6170 & ~n9359;
  assign n9361 = n9258 & n9360;
  assign n9362 = ~n9347 & ~n9361;
  assign n9363 = pi152 & ~n9362;
  assign n9364 = ~n9097 & ~n9297;
  assign n9365 = ~pi210 & ~n9364;
  assign n9366 = n6170 & ~n9365;
  assign n9367 = ~n9097 & ~n9294;
  assign n9368 = n9366 & n9367;
  assign n9369 = ~n9347 & ~n9368;
  assign n9370 = ~pi152 & ~n9369;
  assign n9371 = pi172 & ~n9370;
  assign n9372 = ~n9363 & n9371;
  assign n9373 = ~n9358 & ~n9372;
  assign n9374 = n9344 & ~n9373;
  assign n9375 = ~n9257 & ~n9360;
  assign n9376 = n9256 & ~n9375;
  assign n9377 = pi152 & ~n9376;
  assign n9378 = ~n9257 & ~n9366;
  assign n9379 = n9295 & ~n9378;
  assign n9380 = ~pi152 & ~n9379;
  assign n9381 = pi172 & ~n9380;
  assign n9382 = ~n9377 & n9381;
  assign n9383 = ~n9102 & ~n9181;
  assign n9384 = ~n9348 & n9383;
  assign n9385 = n6170 & n9384;
  assign n9386 = ~pi152 & ~n9385;
  assign n9387 = pi152 & ~n9346;
  assign n9388 = ~pi172 & ~n9386;
  assign n9389 = ~n9387 & n9388;
  assign n9390 = ~pi158 & pi299;
  assign n9391 = ~n9347 & n9390;
  assign n9392 = ~n9389 & n9391;
  assign n9393 = ~n9382 & n9392;
  assign n9394 = ~pi149 & ~n9393;
  assign n9395 = ~n9374 & n9394;
  assign n9396 = ~n9224 & ~n9347;
  assign n9397 = pi152 & ~n9396;
  assign n9398 = ~n9199 & ~n9347;
  assign n9399 = ~pi152 & ~n9398;
  assign n9400 = ~pi172 & ~n9397;
  assign n9401 = ~n9399 & n9400;
  assign n9402 = ~n9315 & ~n9347;
  assign n9403 = pi152 & ~n9402;
  assign n9404 = ~n9257 & ~n9352;
  assign n9405 = ~pi152 & n9404;
  assign n9406 = pi172 & ~n9403;
  assign n9407 = ~n9405 & n9406;
  assign n9408 = ~n9401 & ~n9407;
  assign n9409 = n9344 & ~n9408;
  assign n9410 = ~n9278 & ~n9347;
  assign n9411 = pi152 & ~n9410;
  assign n9412 = ~n9305 & ~n9347;
  assign n9413 = ~pi152 & ~n9412;
  assign n9414 = pi172 & ~n9411;
  assign n9415 = ~n9413 & n9414;
  assign n9416 = ~n9102 & ~n9198;
  assign n9417 = n6170 & ~n9416;
  assign n9418 = ~n9352 & ~n9417;
  assign n9419 = ~pi152 & n9418;
  assign n9420 = ~n9217 & ~n9352;
  assign n9421 = pi152 & n9420;
  assign n9422 = ~pi172 & ~n9419;
  assign n9423 = ~n9421 & n9422;
  assign n9424 = ~n9415 & ~n9423;
  assign n9425 = n9390 & ~n9424;
  assign n9426 = pi149 & ~n9409;
  assign n9427 = ~n9425 & n9426;
  assign n9428 = ~n9395 & ~n9427;
  assign n9429 = ~n9343 & ~n9428;
  assign n9430 = pi232 & ~n9429;
  assign n9431 = ~n6151 & n9159;
  assign n9432 = n9153 & ~n9431;
  assign n9433 = ~pi232 & ~n9432;
  assign n9434 = ~pi39 & ~n9433;
  assign n9435 = ~n9430 & n9434;
  assign n9436 = ~n9096 & ~n9435;
  assign n9437 = ~pi38 & ~n9436;
  assign n9438 = ~n9022 & ~n9437;
  assign n9439 = ~pi100 & ~n9438;
  assign n9440 = ~pi87 & ~n8993;
  assign n9441 = ~n9439 & n9440;
  assign n9442 = pi38 & n9006;
  assign n9443 = ~pi100 & n9442;
  assign n9444 = ~n8993 & ~n9443;
  assign n9445 = n3207 & n9024;
  assign n9446 = pi87 & ~n9445;
  assign n9447 = n9444 & n9446;
  assign n9448 = n3238 & ~n9447;
  assign n9449 = ~n9441 & n9448;
  assign n9450 = ~pi75 & pi92;
  assign n9451 = pi232 & ~n3394;
  assign n9452 = ~pi176 & ~pi299;
  assign n9453 = n6170 & ~n9452;
  assign n9454 = n9451 & n9453;
  assign n9455 = n3222 & n9037;
  assign n9456 = ~n9454 & n9455;
  assign n9457 = n9445 & ~n9456;
  assign n9458 = n9444 & ~n9457;
  assign n9459 = n9450 & ~n9458;
  assign n9460 = ~n8994 & ~n9459;
  assign n9461 = ~n9449 & n9460;
  assign n9462 = ~pi54 & ~n9461;
  assign n9463 = ~n9009 & ~n9462;
  assign n9464 = ~pi74 & ~n9463;
  assign n9465 = n9002 & ~n9464;
  assign n9466 = pi55 & ~n8982;
  assign n9467 = pi54 & ~n8978;
  assign n9468 = ~pi92 & ~n8972;
  assign n9469 = pi164 & n7484;
  assign n9470 = pi38 & ~n9469;
  assign n9471 = n3241 & ~n9470;
  assign n9472 = pi149 & n7484;
  assign n9473 = ~pi39 & ~n9472;
  assign n9474 = n9037 & n9473;
  assign n9475 = n9024 & ~n9474;
  assign n9476 = ~pi38 & ~n9475;
  assign n9477 = n9471 & ~n9476;
  assign n9478 = ~pi38 & ~n9024;
  assign n9479 = ~pi100 & ~n9478;
  assign n9480 = ~n9470 & n9479;
  assign n9481 = pi87 & n9480;
  assign n9482 = ~n8973 & ~n9481;
  assign n9483 = ~n9477 & n9482;
  assign n9484 = ~pi75 & ~n9483;
  assign n9485 = n9468 & ~n9484;
  assign n9486 = ~pi75 & n9480;
  assign n9487 = pi92 & n8974;
  assign n9488 = ~n9486 & n9487;
  assign n9489 = ~pi54 & ~n9488;
  assign n9490 = ~n9485 & n9489;
  assign n9491 = ~n9467 & ~n9490;
  assign n9492 = ~pi74 & ~n9491;
  assign n9493 = n9466 & ~n9492;
  assign n9494 = n3294 & ~n9493;
  assign n9495 = ~n9465 & n9494;
  assign n9496 = pi38 & n9469;
  assign n9497 = n8975 & n9496;
  assign n9498 = n8974 & ~n9497;
  assign n9499 = ~n9467 & n9498;
  assign n9500 = ~pi74 & ~n9499;
  assign n9501 = ~n8982 & ~n9500;
  assign n9502 = ~n3294 & ~n9501;
  assign n9503 = n3432 & ~n9502;
  assign n9504 = ~pi38 & n9024;
  assign n9505 = n8975 & n9504;
  assign n9506 = n3266 & n9505;
  assign n9507 = ~n3294 & n9506;
  assign n9508 = n9503 & ~n9507;
  assign n9509 = ~n9495 & n9508;
  assign n9510 = ~n8984 & ~n9509;
  assign n9511 = ~n8966 & ~n9510;
  assign n9512 = n6228 & ~n6455;
  assign n9513 = pi154 & ~n9512;
  assign n9514 = n6228 & n6459;
  assign n9515 = ~pi154 & ~n9514;
  assign n9516 = ~pi152 & ~n9515;
  assign n9517 = ~n9513 & n9516;
  assign n9518 = n6170 & n7530;
  assign n9519 = ~n6223 & n9518;
  assign n9520 = pi152 & pi154;
  assign n9521 = n9519 & n9520;
  assign n9522 = ~n9517 & ~n9521;
  assign n9523 = n9055 & ~n9522;
  assign n9524 = pi299 & ~n9523;
  assign n9525 = n6207 & n6459;
  assign n9526 = n9044 & n9525;
  assign n9527 = ~pi174 & n9526;
  assign n9528 = ~pi299 & ~n9527;
  assign n9529 = n9023 & ~n9528;
  assign n9530 = ~n6455 & n9044;
  assign n9531 = n6207 & n9530;
  assign n9532 = ~pi174 & n9531;
  assign n9533 = n6207 & n9044;
  assign n9534 = n7530 & n9533;
  assign n9535 = pi174 & n9534;
  assign n9536 = ~pi299 & ~n9535;
  assign n9537 = ~n9532 & n9536;
  assign n9538 = n9085 & ~n9537;
  assign n9539 = ~n9529 & ~n9538;
  assign n9540 = pi39 & ~n9524;
  assign n9541 = ~n9539 & n9540;
  assign n9542 = pi90 & ~n7446;
  assign n9543 = n2547 & ~n6121;
  assign n9544 = ~n9542 & n9543;
  assign n9545 = ~pi90 & n2514;
  assign n9546 = n2547 & n9545;
  assign n9547 = n2508 & n9546;
  assign n9548 = n2476 & n9547;
  assign n9549 = n9126 & n9548;
  assign n9550 = ~pi70 & ~n9549;
  assign n9551 = ~n9544 & n9550;
  assign n9552 = n2952 & n3094;
  assign n9553 = ~n9551 & n9552;
  assign n9554 = ~n9550 & n9552;
  assign n9555 = ~n6379 & ~n9554;
  assign n9556 = ~pi198 & ~n9555;
  assign n9557 = ~n9553 & ~n9556;
  assign n9558 = n9206 & ~n9557;
  assign n9559 = ~pi72 & ~pi93;
  assign n9560 = n2496 & n9559;
  assign n9561 = ~n9542 & n9560;
  assign n9562 = n2476 & n9208;
  assign n9563 = n6121 & ~n9562;
  assign n9564 = n9561 & ~n9563;
  assign n9565 = n3093 & n6170;
  assign n9566 = ~pi40 & n9565;
  assign n9567 = n9564 & n9566;
  assign n9568 = ~pi183 & n9567;
  assign n9569 = ~pi174 & ~n9568;
  assign n9570 = ~n9558 & n9569;
  assign n9571 = ~n9111 & n9547;
  assign n9572 = ~pi70 & ~n9571;
  assign n9573 = ~n9544 & n9572;
  assign n9574 = n9552 & ~n9573;
  assign n9575 = ~n6413 & ~n9574;
  assign n9576 = n6170 & ~n9575;
  assign n9577 = pi183 & n9576;
  assign n9578 = ~n6121 & n9561;
  assign n9579 = n9566 & n9578;
  assign n9580 = ~pi183 & n9579;
  assign n9581 = pi174 & ~n9580;
  assign n9582 = ~n9577 & n9581;
  assign n9583 = ~n9570 & ~n9582;
  assign n9584 = pi193 & ~n9583;
  assign n9585 = ~n6413 & ~n9554;
  assign n9586 = ~pi174 & n9585;
  assign n9587 = n9552 & ~n9572;
  assign n9588 = ~n6413 & ~n9587;
  assign n9589 = pi174 & n9588;
  assign n9590 = n9206 & ~n9589;
  assign n9591 = ~n9586 & n9590;
  assign n9592 = n9154 & n9562;
  assign n9593 = n3093 & n9592;
  assign n9594 = n9227 & n9593;
  assign n9595 = ~pi174 & ~pi183;
  assign n9596 = n9594 & n9595;
  assign n9597 = ~pi193 & ~n9596;
  assign n9598 = ~n9591 & n9597;
  assign n9599 = ~n9584 & ~n9598;
  assign n9600 = n2960 & n6170;
  assign n9601 = pi180 & n9600;
  assign n9602 = ~pi299 & ~n9601;
  assign n9603 = ~n9599 & n9602;
  assign n9604 = ~pi39 & pi232;
  assign n9605 = pi172 & n9553;
  assign n9606 = ~n6380 & ~n9554;
  assign n9607 = ~pi152 & n9606;
  assign n9608 = ~n9605 & n9607;
  assign n9609 = ~n6380 & ~n9587;
  assign n9610 = pi172 & n9574;
  assign n9611 = pi152 & ~n9610;
  assign n9612 = n9609 & n9611;
  assign n9613 = pi149 & n6170;
  assign n9614 = ~n9612 & n9613;
  assign n9615 = ~n9608 & n9614;
  assign n9616 = ~pi152 & n9567;
  assign n9617 = ~n9579 & ~n9616;
  assign n9618 = pi172 & ~n9617;
  assign n9619 = ~pi152 & ~pi172;
  assign n9620 = n9594 & n9619;
  assign n9621 = ~n9618 & ~n9620;
  assign n9622 = ~pi149 & ~n9621;
  assign n9623 = pi158 & n9600;
  assign n9624 = pi299 & ~n9623;
  assign n9625 = ~n9622 & n9624;
  assign n9626 = ~n9615 & n9625;
  assign n9627 = n9604 & ~n9626;
  assign n9628 = ~n9603 & n9627;
  assign n9629 = ~n9541 & ~n9628;
  assign n9630 = ~pi38 & ~n9629;
  assign n9631 = ~pi87 & ~n9022;
  assign n9632 = ~n9630 & n9631;
  assign n9633 = pi87 & ~n9442;
  assign n9634 = ~pi100 & ~n9633;
  assign n9635 = ~n9632 & n9634;
  assign n9636 = ~n8993 & ~n9635;
  assign n9637 = n3238 & ~n9636;
  assign n9638 = ~pi38 & ~pi87;
  assign n9639 = ~pi100 & n9638;
  assign n9640 = n9454 & n9639;
  assign n9641 = n6117 & n9640;
  assign n9642 = n9444 & ~n9641;
  assign n9643 = n9450 & ~n9642;
  assign n9644 = ~n8994 & ~n9643;
  assign n9645 = ~n9637 & n9644;
  assign n9646 = ~pi54 & ~n9645;
  assign n9647 = ~n9009 & ~n9646;
  assign n9648 = ~pi74 & ~n9647;
  assign n9649 = n9002 & ~n9648;
  assign n9650 = n6117 & n9472;
  assign n9651 = ~pi38 & ~n9650;
  assign n9652 = n9471 & ~n9651;
  assign n9653 = n7599 & n9496;
  assign n9654 = ~n8973 & ~n9653;
  assign n9655 = ~n9652 & n9654;
  assign n9656 = ~pi75 & ~n9655;
  assign n9657 = n9468 & ~n9656;
  assign n9658 = pi92 & n9498;
  assign n9659 = ~pi54 & ~n9658;
  assign n9660 = ~n9657 & n9659;
  assign n9661 = ~n9467 & ~n9660;
  assign n9662 = ~pi74 & ~n9661;
  assign n9663 = n9466 & ~n9662;
  assign n9664 = n3294 & ~n9663;
  assign n9665 = ~n9649 & n9664;
  assign n9666 = n9503 & ~n9665;
  assign n9667 = ~n8984 & ~n9666;
  assign n9668 = n8966 & ~n9667;
  assign n9669 = ~pi954 & ~n9668;
  assign n9670 = ~n9511 & n9669;
  assign n9671 = ~pi33 & ~n9510;
  assign n9672 = pi33 & ~n9667;
  assign n9673 = pi954 & ~n9672;
  assign n9674 = ~n9671 & n9673;
  assign po191 = ~n9670 & ~n9674;
  assign n9676 = pi197 & n8968;
  assign n9677 = ~pi197 & ~n8968;
  assign n9678 = ~n9676 & ~n9677;
  assign n9679 = pi162 & n6170;
  assign n9680 = n9678 & ~n9679;
  assign n9681 = n9676 & n9679;
  assign n9682 = ~pi162 & ~pi197;
  assign n9683 = n8969 & ~n9682;
  assign n9684 = n6170 & ~n9683;
  assign n9685 = ~n9681 & n9684;
  assign n9686 = ~n9678 & ~n9685;
  assign n9687 = ~n9680 & ~n9686;
  assign n9688 = pi232 & n9687;
  assign n9689 = ~n8975 & n9688;
  assign n9690 = pi167 & n7484;
  assign n9691 = n8975 & n9690;
  assign n9692 = ~n9689 & ~n9691;
  assign n9693 = ~pi74 & n9692;
  assign n9694 = pi148 & n8976;
  assign n9695 = pi74 & ~n9694;
  assign n9696 = ~n9689 & n9695;
  assign n9697 = ~n9693 & ~n9696;
  assign n9698 = ~n3432 & n9697;
  assign n9699 = ~pi54 & ~n9689;
  assign n9700 = pi38 & n9691;
  assign n9701 = n9699 & ~n9700;
  assign n9702 = ~pi74 & n9701;
  assign n9703 = n9697 & ~n9702;
  assign n9704 = ~n3294 & ~n9703;
  assign n9705 = n3432 & ~n9704;
  assign n9706 = ~n3294 & ~n9506;
  assign n9707 = n3432 & ~n9706;
  assign n9708 = ~n9705 & ~n9707;
  assign n9709 = pi299 & ~n9687;
  assign n9710 = pi140 & pi145;
  assign n9711 = n8987 & ~n9710;
  assign n9712 = ~pi140 & ~pi145;
  assign n9713 = n6170 & ~n9712;
  assign n9714 = n9711 & n9713;
  assign n9715 = ~n9710 & ~n9712;
  assign n9716 = n8988 & ~n9715;
  assign n9717 = ~pi299 & ~n9714;
  assign n9718 = ~n9716 & n9717;
  assign n9719 = pi232 & ~n9718;
  assign n9720 = ~n9709 & n9719;
  assign n9721 = pi100 & ~n9720;
  assign n9722 = pi75 & ~n9720;
  assign n9723 = ~n9721 & ~n9722;
  assign n9724 = pi141 & ~pi299;
  assign n9725 = pi148 & pi299;
  assign n9726 = ~n9724 & ~n9725;
  assign n9727 = n7484 & ~n9726;
  assign n9728 = n8975 & ~n9727;
  assign n9729 = n9723 & ~n9728;
  assign n9730 = pi74 & ~n9729;
  assign n9731 = ~pi55 & ~n9730;
  assign n9732 = pi188 & ~pi299;
  assign n9733 = pi167 & pi299;
  assign n9734 = ~n9732 & ~n9733;
  assign n9735 = n7484 & ~n9734;
  assign n9736 = ~pi100 & ~n9735;
  assign n9737 = ~pi75 & n9736;
  assign n9738 = n9723 & ~n9737;
  assign n9739 = pi54 & ~n9738;
  assign n9740 = ~pi142 & ~n9270;
  assign n9741 = pi142 & n9161;
  assign n9742 = ~pi140 & ~n9741;
  assign n9743 = ~n9740 & n9742;
  assign n9744 = ~pi142 & ~n9279;
  assign n9745 = pi142 & ~n9217;
  assign n9746 = ~n9283 & n9745;
  assign n9747 = pi140 & ~n9746;
  assign n9748 = ~n9744 & n9747;
  assign n9749 = ~n9743 & ~n9748;
  assign n9750 = ~pi181 & ~n9749;
  assign n9751 = ~pi142 & ~n9313;
  assign n9752 = pi142 & ~n9231;
  assign n9753 = ~pi140 & ~n9752;
  assign n9754 = ~n9751 & n9753;
  assign n9755 = pi142 & ~n9225;
  assign n9756 = ~pi142 & ~n9316;
  assign n9757 = pi140 & ~n9755;
  assign n9758 = ~n9756 & n9757;
  assign n9759 = ~n9754 & ~n9758;
  assign n9760 = pi181 & ~n9759;
  assign n9761 = pi144 & ~n9760;
  assign n9762 = ~n9750 & n9761;
  assign n9763 = pi142 & ~n9184;
  assign n9764 = ~pi142 & ~n9334;
  assign n9765 = ~pi140 & ~n9763;
  assign n9766 = ~n9764 & n9765;
  assign n9767 = ~pi142 & n9320;
  assign n9768 = pi142 & ~n9200;
  assign n9769 = pi140 & ~n9767;
  assign n9770 = ~n9768 & n9769;
  assign n9771 = ~n9766 & ~n9770;
  assign n9772 = pi181 & ~n9771;
  assign n9773 = ~pi142 & n9301;
  assign n9774 = ~n9178 & n9383;
  assign n9775 = n6170 & ~n9774;
  assign n9776 = pi142 & ~n9775;
  assign n9777 = ~n9283 & n9776;
  assign n9778 = ~pi140 & ~n9777;
  assign n9779 = ~n9773 & n9778;
  assign n9780 = ~pi142 & ~n9306;
  assign n9781 = pi142 & ~n9417;
  assign n9782 = ~n9283 & n9781;
  assign n9783 = pi140 & ~n9782;
  assign n9784 = ~n9780 & n9783;
  assign n9785 = ~n9779 & ~n9784;
  assign n9786 = ~pi181 & ~n9785;
  assign n9787 = ~pi144 & ~n9786;
  assign n9788 = ~n9772 & n9787;
  assign n9789 = ~pi299 & ~n9788;
  assign n9790 = ~n9762 & n9789;
  assign n9791 = ~pi159 & pi299;
  assign n9792 = pi146 & n9418;
  assign n9793 = ~pi146 & ~n9412;
  assign n9794 = ~pi161 & ~n9792;
  assign n9795 = ~n9793 & n9794;
  assign n9796 = pi146 & n9420;
  assign n9797 = ~pi146 & ~n9410;
  assign n9798 = pi161 & ~n9796;
  assign n9799 = ~n9797 & n9798;
  assign n9800 = ~n9795 & ~n9799;
  assign n9801 = pi162 & ~n9800;
  assign n9802 = pi161 & ~n9376;
  assign n9803 = ~pi161 & ~n9379;
  assign n9804 = ~pi146 & ~n9803;
  assign n9805 = ~n9802 & n9804;
  assign n9806 = ~pi161 & ~n9385;
  assign n9807 = pi161 & ~n9346;
  assign n9808 = pi146 & ~n9806;
  assign n9809 = ~n9807 & n9808;
  assign n9810 = ~pi162 & ~n9347;
  assign n9811 = ~n9809 & n9810;
  assign n9812 = ~n9805 & n9811;
  assign n9813 = ~n9801 & ~n9812;
  assign n9814 = n9791 & ~n9813;
  assign n9815 = ~pi146 & ~n9362;
  assign n9816 = pi146 & n9355;
  assign n9817 = pi161 & ~n9816;
  assign n9818 = ~n9815 & n9817;
  assign n9819 = pi146 & ~n9350;
  assign n9820 = ~pi146 & ~n9369;
  assign n9821 = ~pi161 & ~n9819;
  assign n9822 = ~n9820 & n9821;
  assign n9823 = ~pi162 & ~n9818;
  assign n9824 = ~n9822 & n9823;
  assign n9825 = ~pi146 & n9404;
  assign n9826 = pi146 & ~n9398;
  assign n9827 = ~pi161 & ~n9825;
  assign n9828 = ~n9826 & n9827;
  assign n9829 = pi146 & ~n9396;
  assign n9830 = ~pi146 & ~n9402;
  assign n9831 = pi161 & ~n9829;
  assign n9832 = ~n9830 & n9831;
  assign n9833 = pi162 & ~n9828;
  assign n9834 = ~n9832 & n9833;
  assign n9835 = pi159 & pi299;
  assign n9836 = ~n9824 & n9835;
  assign n9837 = ~n9834 & n9836;
  assign n9838 = ~n9814 & ~n9837;
  assign n9839 = ~n9790 & n9838;
  assign n9840 = pi232 & ~n9839;
  assign n9841 = ~n9433 & ~n9840;
  assign n9842 = n3182 & ~n9841;
  assign n9843 = pi144 & n9090;
  assign n9844 = ~pi177 & ~pi299;
  assign n9845 = ~pi144 & ~n9046;
  assign n9846 = ~n9081 & n9845;
  assign n9847 = n9844 & ~n9846;
  assign n9848 = ~n9843 & n9847;
  assign n9849 = ~n9046 & ~n9051;
  assign n9850 = pi177 & ~pi299;
  assign n9851 = ~n9845 & n9850;
  assign n9852 = ~n9849 & n9851;
  assign n9853 = ~n9848 & ~n9852;
  assign n9854 = pi232 & ~n9853;
  assign n9855 = ~n9093 & ~n9854;
  assign n9856 = ~pi38 & ~n9855;
  assign n9857 = ~pi161 & n9065;
  assign n9858 = ~n9061 & ~n9857;
  assign n9859 = n9055 & ~n9858;
  assign n9860 = ~pi38 & ~pi155;
  assign n9861 = n9057 & n9860;
  assign n9862 = ~n9859 & n9861;
  assign n9863 = pi161 & n9070;
  assign n9864 = n9043 & n9055;
  assign n9865 = ~n9863 & n9864;
  assign n9866 = ~pi38 & pi155;
  assign n9867 = n9057 & n9866;
  assign n9868 = ~n9865 & n9867;
  assign n9869 = ~n9862 & ~n9868;
  assign n9870 = pi232 & ~n9869;
  assign n9871 = ~n9856 & ~n9870;
  assign n9872 = pi39 & ~n9871;
  assign n9873 = pi188 & n9018;
  assign n9874 = ~pi167 & ~n9873;
  assign n9875 = ~pi188 & ~n9011;
  assign n9876 = pi167 & pi188;
  assign n9877 = ~n9013 & n9876;
  assign n9878 = ~n9875 & ~n9877;
  assign n9879 = ~n9874 & n9878;
  assign n9880 = pi38 & ~n9879;
  assign n9881 = ~pi87 & ~n9880;
  assign n9882 = ~n9872 & n9881;
  assign n9883 = ~n9842 & n9882;
  assign n9884 = pi38 & ~n9735;
  assign n9885 = ~n9478 & ~n9884;
  assign n9886 = pi87 & n9885;
  assign n9887 = ~pi100 & ~n9886;
  assign n9888 = ~n9883 & n9887;
  assign n9889 = ~n9721 & ~n9888;
  assign n9890 = n3238 & ~n9889;
  assign n9891 = pi155 & pi299;
  assign n9892 = ~n9850 & ~n9891;
  assign n9893 = ~pi38 & n9892;
  assign n9894 = n7484 & ~n9893;
  assign n9895 = n9455 & ~n9894;
  assign n9896 = n9885 & ~n9895;
  assign n9897 = ~pi100 & ~n9896;
  assign n9898 = ~n9721 & ~n9897;
  assign n9899 = n9450 & ~n9898;
  assign n9900 = ~n9722 & ~n9899;
  assign n9901 = ~n9890 & n9900;
  assign n9902 = ~pi54 & ~n9901;
  assign n9903 = ~n9739 & ~n9902;
  assign n9904 = ~pi74 & ~n9903;
  assign n9905 = n9731 & ~n9904;
  assign n9906 = pi55 & ~n9696;
  assign n9907 = pi54 & n9692;
  assign n9908 = ~n9505 & n9701;
  assign n9909 = ~n6279 & ~n9908;
  assign n9910 = pi100 & ~n9688;
  assign n9911 = pi38 & n9690;
  assign n9912 = n9455 & ~n9679;
  assign n9913 = n9504 & ~n9912;
  assign n9914 = ~pi100 & ~n9913;
  assign n9915 = ~pi232 & n9455;
  assign n9916 = ~n9914 & ~n9915;
  assign n9917 = ~n9911 & ~n9916;
  assign n9918 = ~n9910 & ~n9917;
  assign n9919 = ~pi75 & ~n9918;
  assign n9920 = pi75 & ~n9688;
  assign n9921 = ~pi92 & ~n9920;
  assign n9922 = ~n9919 & n9921;
  assign n9923 = ~n9909 & ~n9922;
  assign n9924 = ~n9907 & ~n9923;
  assign n9925 = ~pi74 & ~n9924;
  assign n9926 = n9906 & ~n9925;
  assign n9927 = n3294 & ~n9926;
  assign n9928 = ~n9905 & n9927;
  assign n9929 = ~n9708 & ~n9928;
  assign n9930 = ~n9698 & ~n9929;
  assign n9931 = ~pi34 & n9930;
  assign n9932 = ~pi146 & ~n9567;
  assign n9933 = pi146 & ~n9594;
  assign n9934 = ~pi161 & ~n9933;
  assign n9935 = ~n9932 & n9934;
  assign n9936 = ~pi146 & pi161;
  assign n9937 = n9579 & n9936;
  assign n9938 = ~n9935 & ~n9937;
  assign n9939 = ~pi162 & ~n9938;
  assign n9940 = ~pi162 & n9600;
  assign n9941 = n9835 & ~n9940;
  assign n9942 = ~n9791 & ~n9941;
  assign n9943 = ~n9679 & ~n9942;
  assign n9944 = ~pi146 & n9553;
  assign n9945 = n9606 & ~n9944;
  assign n9946 = ~pi161 & ~n9945;
  assign n9947 = ~pi146 & n9574;
  assign n9948 = n9609 & ~n9947;
  assign n9949 = pi161 & ~n9948;
  assign n9950 = pi159 & n2960;
  assign n9951 = pi299 & ~n9950;
  assign n9952 = ~n9949 & n9951;
  assign n9953 = ~n9946 & n9952;
  assign n9954 = ~n9943 & ~n9953;
  assign n9955 = ~n9939 & ~n9954;
  assign n9956 = ~pi142 & n9567;
  assign n9957 = pi142 & n9594;
  assign n9958 = ~pi140 & ~n9957;
  assign n9959 = ~n9956 & n9958;
  assign n9960 = ~pi142 & n9553;
  assign n9961 = pi140 & n9585;
  assign n9962 = ~n9960 & n9961;
  assign n9963 = ~n9959 & ~n9962;
  assign n9964 = ~pi144 & ~n9963;
  assign n9965 = pi140 & ~n6170;
  assign n9966 = ~pi142 & n9579;
  assign n9967 = ~pi140 & ~n9966;
  assign n9968 = ~pi142 & n9574;
  assign n9969 = pi140 & ~n9968;
  assign n9970 = n9588 & n9969;
  assign n9971 = ~n9967 & ~n9970;
  assign n9972 = pi144 & ~n9971;
  assign n9973 = ~n9965 & ~n9972;
  assign n9974 = ~n9964 & n9973;
  assign n9975 = pi181 & n9600;
  assign n9976 = ~pi299 & ~n9975;
  assign n9977 = ~n9974 & n9976;
  assign n9978 = pi232 & ~n9955;
  assign n9979 = ~n9977 & n9978;
  assign n9980 = n3182 & ~n9979;
  assign n9981 = pi161 & ~n9519;
  assign n9982 = ~pi161 & ~n9512;
  assign n9983 = n9055 & ~n9982;
  assign n9984 = ~n9981 & n9983;
  assign n9985 = n9866 & ~n9984;
  assign n9986 = ~pi161 & n9055;
  assign n9987 = n9514 & n9986;
  assign n9988 = n9860 & ~n9987;
  assign n9989 = ~n9985 & ~n9988;
  assign n9990 = pi299 & ~n9989;
  assign n9991 = ~pi144 & n9531;
  assign n9992 = pi144 & n9534;
  assign n9993 = n9850 & ~n9992;
  assign n9994 = ~n9991 & n9993;
  assign n9995 = ~pi144 & n9526;
  assign n9996 = n9844 & ~n9995;
  assign n9997 = pi232 & ~n9996;
  assign n9998 = ~n9994 & n9997;
  assign n9999 = ~pi38 & ~n9998;
  assign n10000 = ~n9990 & ~n9999;
  assign n10001 = pi39 & ~n10000;
  assign n10002 = ~n9880 & ~n10001;
  assign n10003 = ~n9980 & n10002;
  assign n10004 = ~pi100 & ~n10003;
  assign n10005 = ~n9721 & ~n10004;
  assign n10006 = ~pi87 & ~n10005;
  assign n10007 = ~n3207 & ~n9736;
  assign n10008 = ~n9721 & n10007;
  assign n10009 = pi87 & ~n10008;
  assign n10010 = ~n10006 & ~n10009;
  assign n10011 = n3238 & ~n10010;
  assign n10012 = pi38 & ~n9734;
  assign n10013 = n3182 & ~n9892;
  assign n10014 = n3090 & n10013;
  assign n10015 = ~n10012 & ~n10014;
  assign n10016 = n7484 & ~n10015;
  assign n10017 = ~pi100 & ~n10016;
  assign n10018 = ~n9721 & ~n10017;
  assign n10019 = ~pi87 & ~n10018;
  assign n10020 = ~n10009 & ~n10019;
  assign n10021 = n9450 & ~n10020;
  assign n10022 = ~n9722 & ~n10021;
  assign n10023 = ~n10011 & n10022;
  assign n10024 = ~pi54 & ~n10023;
  assign n10025 = ~n9739 & ~n10024;
  assign n10026 = ~pi74 & ~n10025;
  assign n10027 = n9731 & ~n10026;
  assign n10028 = ~pi92 & pi162;
  assign n10029 = n9604 & n10028;
  assign n10030 = n9638 & n10029;
  assign n10031 = n6188 & n10030;
  assign n10032 = ~n9911 & ~n10031;
  assign n10033 = n8975 & ~n10032;
  assign n10034 = n9699 & ~n10033;
  assign n10035 = ~n9907 & ~n10034;
  assign n10036 = ~pi74 & ~n10035;
  assign n10037 = n9906 & ~n10036;
  assign n10038 = n3294 & ~n10037;
  assign n10039 = ~n10027 & n10038;
  assign n10040 = n9705 & ~n10039;
  assign n10041 = ~n9698 & ~n10040;
  assign n10042 = pi34 & n10041;
  assign n10043 = ~pi33 & ~pi954;
  assign n10044 = ~n10042 & ~n10043;
  assign n10045 = ~n9931 & n10044;
  assign n10046 = ~pi34 & ~n8964;
  assign n10047 = n9930 & ~n10046;
  assign n10048 = n10041 & n10046;
  assign n10049 = n10043 & ~n10048;
  assign n10050 = ~n10047 & n10049;
  assign po192 = ~n10045 & ~n10050;
  assign n10052 = pi137 & n8870;
  assign n10053 = pi1091 & pi1093;
  assign n10054 = n2733 & n10053;
  assign n10055 = n7496 & ~n10054;
  assign n10056 = pi683 & n10055;
  assign n10057 = pi252 & po1057;
  assign n10058 = ~n10056 & n10057;
  assign n10059 = ~n6248 & ~n8875;
  assign n10060 = ~n10058 & n10059;
  assign n10061 = ~n8875 & ~n10060;
  assign n10062 = ~n8873 & ~n10061;
  assign n10063 = ~n10060 & ~n10062;
  assign n10064 = n8872 & ~n10063;
  assign n10065 = ~n10052 & ~n10064;
  assign n10066 = n8868 & ~n10065;
  assign n10067 = ~pi90 & n6120;
  assign n10068 = ~pi93 & ~n10067;
  assign n10069 = ~n6139 & ~n10068;
  assign n10070 = ~pi35 & ~n10069;
  assign n10071 = pi35 & ~n2736;
  assign n10072 = n8924 & ~n10071;
  assign n10073 = ~n10070 & n10072;
  assign n10074 = ~pi32 & n10073;
  assign n10075 = pi32 & ~pi93;
  assign n10076 = n8881 & n10075;
  assign n10077 = n7446 & n10076;
  assign n10078 = ~n10074 & ~n10077;
  assign n10079 = ~pi95 & ~n6151;
  assign n10080 = ~n10078 & n10079;
  assign n10081 = n6151 & ~n10070;
  assign n10082 = n2734 & n7547;
  assign n10083 = ~pi137 & ~n6151;
  assign n10084 = ~n7720 & ~n10083;
  assign n10085 = n10082 & n10084;
  assign n10086 = ~pi122 & ~po740;
  assign n10087 = n7720 & ~n10083;
  assign n10088 = n10086 & n10087;
  assign n10089 = ~n10085 & ~n10088;
  assign n10090 = ~n10081 & n10089;
  assign n10091 = n2493 & n8922;
  assign n10092 = n10070 & ~n10091;
  assign n10093 = n3093 & n10072;
  assign n10094 = ~n10092 & n10093;
  assign n10095 = ~n10090 & n10094;
  assign n10096 = ~n2553 & ~n10073;
  assign n10097 = pi1082 & n3093;
  assign n10098 = ~n10096 & n10097;
  assign n10099 = ~pi38 & ~n10095;
  assign n10100 = ~n10098 & n10099;
  assign n10101 = ~n10080 & n10100;
  assign n10102 = pi38 & ~n8948;
  assign n10103 = ~pi39 & ~pi100;
  assign n10104 = ~n10102 & n10103;
  assign n10105 = ~n10101 & n10104;
  assign n10106 = ~n10066 & ~n10105;
  assign n10107 = n3231 & ~n10106;
  assign n10108 = pi137 & ~po840;
  assign n10109 = ~n6271 & n10108;
  assign n10110 = ~n8950 & ~n10109;
  assign n10111 = n8953 & ~n10110;
  assign n10112 = n8948 & n10111;
  assign n10113 = ~n10107 & ~n10112;
  assign n10114 = ~pi92 & ~n10113;
  assign n10115 = ~pi54 & ~n10114;
  assign n10116 = ~pi24 & n7330;
  assign n10117 = pi54 & ~n10116;
  assign n10118 = n3294 & n8865;
  assign n10119 = ~n10117 & n10118;
  assign n10120 = ~n10115 & n10119;
  assign n10121 = ~pi59 & ~n10120;
  assign n10122 = n3269 & n3294;
  assign n10123 = n8948 & n10122;
  assign n10124 = ~pi55 & n10123;
  assign n10125 = pi59 & ~n10124;
  assign n10126 = ~pi57 & ~n10125;
  assign po193 = ~n10121 & n10126;
  assign n10128 = n2514 & n2580;
  assign n10129 = ~pi83 & n2647;
  assign n10130 = ~pi65 & n2451;
  assign n10131 = n2476 & n10130;
  assign n10132 = n9025 & n10131;
  assign n10133 = ~pi69 & n10132;
  assign n10134 = ~pi67 & ~pi71;
  assign n10135 = pi36 & ~pi103;
  assign n10136 = n10134 & n10135;
  assign n10137 = n10133 & n10136;
  assign n10138 = n10129 & n10137;
  assign n10139 = n10128 & n10138;
  assign n10140 = ~pi58 & n7501;
  assign n10141 = ~n10139 & ~n10140;
  assign n10142 = n2493 & n6371;
  assign n10143 = n6152 & n10142;
  assign n10144 = n3266 & ~po1038;
  assign n10145 = n3409 & n10144;
  assign n10146 = ~pi92 & n10145;
  assign n10147 = n10143 & n10146;
  assign n10148 = po740 & n10147;
  assign po194 = ~n10141 & n10148;
  assign n10150 = ~pi39 & n3094;
  assign n10151 = pi24 & n10150;
  assign n10152 = n2498 & n10151;
  assign n10153 = pi38 & ~n10152;
  assign n10154 = ~pi81 & ~n2598;
  assign n10155 = ~pi71 & n2476;
  assign n10156 = ~pi104 & n2461;
  assign n10157 = n10155 & n10156;
  assign n10158 = ~pi45 & ~pi73;
  assign n10159 = n8896 & n10158;
  assign n10160 = ~pi48 & ~pi65;
  assign n10161 = ~pi82 & ~pi84;
  assign n10162 = pi89 & n10161;
  assign n10163 = n10160 & n10162;
  assign n10164 = n10159 & n10163;
  assign n10165 = n9116 & n10164;
  assign n10166 = n10157 & n10165;
  assign n10167 = pi332 & n10166;
  assign n10168 = ~pi64 & ~n10167;
  assign n10169 = n6371 & n9241;
  assign n10170 = n2520 & n10169;
  assign n10171 = n2551 & n10170;
  assign n10172 = ~pi39 & ~pi841;
  assign n10173 = n2454 & n10172;
  assign n10174 = ~n10168 & n10173;
  assign n10175 = n10171 & n10174;
  assign n10176 = n10154 & n10175;
  assign n10177 = ~pi38 & ~n10176;
  assign n10178 = n3268 & ~po1038;
  assign n10179 = ~n10177 & n10178;
  assign po196 = ~n10153 & n10179;
  assign n10181 = ~pi38 & n10178;
  assign n10182 = ~pi984 & ~n6265;
  assign n10183 = pi835 & ~n10182;
  assign n10184 = n6173 & ~n10183;
  assign n10185 = n6183 & ~n10184;
  assign n10186 = pi1093 & n10185;
  assign n10187 = n6174 & n6443;
  assign n10188 = ~n10186 & n10187;
  assign n10189 = ~pi223 & n10188;
  assign n10190 = n6206 & n10185;
  assign n10191 = n10187 & ~n10190;
  assign n10192 = n6197 & n10191;
  assign n10193 = ~n6200 & n10185;
  assign n10194 = n10187 & ~n10193;
  assign n10195 = ~n6197 & n10194;
  assign n10196 = ~pi299 & ~n10192;
  assign n10197 = ~n10195 & n10196;
  assign n10198 = ~n10189 & n10197;
  assign n10199 = ~pi215 & n10188;
  assign n10200 = n6223 & n10191;
  assign n10201 = ~n6223 & n10194;
  assign n10202 = pi299 & ~n10200;
  assign n10203 = ~n10201 & n10202;
  assign n10204 = ~n10199 & n10203;
  assign n10205 = pi786 & ~pi1082;
  assign n10206 = ~n10198 & ~n10205;
  assign n10207 = ~n10204 & n10206;
  assign n10208 = n5774 & ~n6229;
  assign n10209 = n3483 & ~n6208;
  assign n10210 = ~n10208 & ~n10209;
  assign n10211 = po740 & n10205;
  assign n10212 = ~n10210 & n10211;
  assign n10213 = n6445 & n10212;
  assign n10214 = ~n10207 & ~n10213;
  assign n10215 = pi39 & ~n10214;
  assign n10216 = ~pi39 & ~pi95;
  assign n10217 = n6151 & n6378;
  assign n10218 = n2510 & ~n2583;
  assign n10219 = n8899 & n9117;
  assign n10220 = ~pi65 & ~pi69;
  assign n10221 = n10219 & n10220;
  assign n10222 = pi48 & ~pi49;
  assign n10223 = ~pi68 & ~pi82;
  assign n10224 = n10222 & n10223;
  assign n10225 = n10158 & n10224;
  assign n10226 = n8898 & n8901;
  assign n10227 = n9114 & n10226;
  assign n10228 = n10221 & n10225;
  assign n10229 = n10227 & n10228;
  assign n10230 = n10157 & n10229;
  assign n10231 = ~pi841 & n2481;
  assign n10232 = n2505 & n10231;
  assign n10233 = ~pi97 & n10232;
  assign n10234 = n10230 & n10233;
  assign n10235 = n10218 & n10234;
  assign n10236 = pi108 & n2510;
  assign n10237 = n2582 & n10236;
  assign n10238 = ~pi47 & ~n10237;
  assign n10239 = ~n10235 & n10238;
  assign n10240 = ~pi986 & ~po740;
  assign n10241 = pi252 & ~n10240;
  assign n10242 = pi314 & ~n10241;
  assign n10243 = n6133 & n10242;
  assign n10244 = ~n10239 & n10243;
  assign n10245 = ~pi47 & ~pi841;
  assign n10246 = n10230 & n10245;
  assign n10247 = ~n2569 & ~n10246;
  assign n10248 = n2489 & n2519;
  assign n10249 = ~n10242 & n10248;
  assign n10250 = ~n10247 & n10249;
  assign n10251 = ~n10244 & ~n10250;
  assign n10252 = n2493 & ~n10251;
  assign n10253 = ~pi35 & ~n10252;
  assign n10254 = pi35 & ~n6375;
  assign n10255 = n2551 & ~n10254;
  assign n10256 = n2725 & n10255;
  assign n10257 = ~n10253 & n10256;
  assign n10258 = ~n10217 & ~n10257;
  assign n10259 = n10216 & ~n10258;
  assign n10260 = ~n10215 & ~n10259;
  assign po197 = n10181 & ~n10260;
  assign n10262 = n3093 & ~n3362;
  assign n10263 = pi102 & n2534;
  assign n10264 = n2453 & n10263;
  assign n10265 = n6152 & n10264;
  assign n10266 = n2520 & n10265;
  assign n10267 = n2479 & n10266;
  assign n10268 = ~pi40 & ~n10267;
  assign n10269 = n10262 & ~n10268;
  assign n10270 = ~pi1082 & ~n10269;
  assign n10271 = n6371 & n10267;
  assign n10272 = pi1082 & ~n10271;
  assign n10273 = n10146 & ~n10272;
  assign po198 = ~n10270 & n10273;
  assign n10275 = ~pi41 & ~pi72;
  assign n10276 = ~n8087 & ~n10275;
  assign n10277 = ~n2734 & n10275;
  assign n10278 = n8087 & ~n10277;
  assign n10279 = ~pi44 & n3096;
  assign n10280 = ~pi101 & n10279;
  assign n10281 = n7547 & n10280;
  assign n10282 = n7487 & n10281;
  assign n10283 = pi41 & ~n10282;
  assign n10284 = ~pi41 & pi72;
  assign n10285 = n2734 & ~n10284;
  assign n10286 = ~pi99 & n6260;
  assign n10287 = ~pi72 & pi101;
  assign n10288 = ~pi41 & ~n10287;
  assign n10289 = ~pi24 & n2498;
  assign n10290 = pi252 & n6371;
  assign n10291 = n7547 & n10290;
  assign n10292 = n10289 & n10291;
  assign n10293 = ~pi44 & n10292;
  assign n10294 = n10288 & n10293;
  assign n10295 = ~n10286 & n10294;
  assign n10296 = n10285 & ~n10295;
  assign n10297 = ~n10283 & n10296;
  assign n10298 = n10278 & ~n10297;
  assign n10299 = ~n10276 & ~n10298;
  assign n10300 = ~pi39 & ~n10299;
  assign n10301 = ~pi189 & n6170;
  assign n10302 = pi144 & n10301;
  assign n10303 = ~pi174 & n10302;
  assign n10304 = ~pi299 & ~n10303;
  assign n10305 = ~pi166 & n6170;
  assign n10306 = pi161 & n10305;
  assign n10307 = ~pi152 & n10306;
  assign n10308 = ~n6242 & ~n10307;
  assign n10309 = pi232 & ~n10304;
  assign n10310 = ~n10308 & n10309;
  assign n10311 = ~pi72 & ~n10310;
  assign n10312 = pi39 & ~n10311;
  assign n10313 = n3242 & ~n10312;
  assign n10314 = ~n10300 & n10313;
  assign n10315 = ~pi39 & ~n10275;
  assign n10316 = ~n10312 & ~n10315;
  assign n10317 = ~n3242 & n10316;
  assign n10318 = pi75 & ~n10317;
  assign n10319 = ~n10314 & n10318;
  assign n10320 = n7465 & ~n7471;
  assign n10321 = ~pi1093 & ~n7473;
  assign n10322 = ~n10320 & n10321;
  assign n10323 = ~pi44 & ~n10322;
  assign n10324 = n2762 & ~n7457;
  assign n10325 = n2759 & n10324;
  assign n10326 = ~n7501 & ~n10325;
  assign n10327 = n2518 & ~n10326;
  assign n10328 = n7448 & ~n10327;
  assign n10329 = n7445 & ~n10328;
  assign n10330 = ~pi51 & ~n10329;
  assign n10331 = ~n2558 & ~n10330;
  assign n10332 = ~pi96 & ~n10331;
  assign n10333 = n6371 & ~n7468;
  assign n10334 = ~pi72 & n7471;
  assign n10335 = n10333 & n10334;
  assign n10336 = ~n10332 & n10335;
  assign n10337 = ~n10320 & ~n10336;
  assign n10338 = pi1093 & n10337;
  assign n10339 = n10323 & ~n10338;
  assign n10340 = ~pi101 & n10339;
  assign n10341 = pi41 & ~n10340;
  assign n10342 = pi44 & pi72;
  assign n10343 = ~pi72 & ~n7465;
  assign n10344 = ~n7471 & n10343;
  assign n10345 = ~n7467 & n10333;
  assign n10346 = n10334 & ~n10345;
  assign n10347 = ~pi1093 & ~n10344;
  assign n10348 = ~n10346 & n10347;
  assign n10349 = ~pi72 & n10337;
  assign n10350 = pi1093 & ~n10349;
  assign n10351 = ~n10348 & ~n10350;
  assign n10352 = ~pi44 & ~n10351;
  assign n10353 = ~n10342 & ~n10352;
  assign n10354 = ~pi101 & n10353;
  assign n10355 = n10288 & ~n10354;
  assign n10356 = n2734 & ~n10355;
  assign n10357 = ~n10341 & n10356;
  assign n10358 = pi1093 & ~n7465;
  assign n10359 = n10323 & ~n10358;
  assign n10360 = ~pi101 & n10359;
  assign n10361 = pi41 & ~n10360;
  assign n10362 = n10343 & ~n10348;
  assign n10363 = pi44 & ~pi72;
  assign n10364 = ~n10362 & ~n10363;
  assign n10365 = ~pi101 & ~n10364;
  assign n10366 = n10288 & ~n10365;
  assign n10367 = ~n2734 & ~n10366;
  assign n10368 = ~n10361 & n10367;
  assign n10369 = pi228 & ~n10368;
  assign n10370 = ~n10357 & n10369;
  assign n10371 = ~pi480 & pi949;
  assign n10372 = n2514 & n2589;
  assign n10373 = n2497 & n10372;
  assign n10374 = ~n10371 & n10373;
  assign n10375 = ~pi109 & n6341;
  assign n10376 = n2589 & n10375;
  assign n10377 = ~pi110 & ~n10376;
  assign n10378 = n2489 & ~n2568;
  assign n10379 = n2497 & n10371;
  assign n10380 = ~pi47 & n10379;
  assign n10381 = n10378 & n10380;
  assign n10382 = ~n10377 & n10381;
  assign n10383 = pi901 & ~pi959;
  assign n10384 = ~n10374 & n10383;
  assign n10385 = ~n10382 & n10384;
  assign n10386 = n2490 & n2567;
  assign n10387 = pi110 & n10386;
  assign n10388 = n10379 & n10387;
  assign n10389 = ~n10383 & ~n10388;
  assign n10390 = ~pi250 & pi252;
  assign n10391 = n6371 & n10390;
  assign n10392 = ~n10389 & n10391;
  assign n10393 = ~n10385 & n10392;
  assign n10394 = ~pi72 & n10393;
  assign n10395 = n10143 & n10387;
  assign n10396 = n10371 & ~n10390;
  assign n10397 = n10395 & n10396;
  assign n10398 = ~n10394 & ~n10397;
  assign n10399 = ~pi44 & ~n10398;
  assign n10400 = ~pi101 & n10399;
  assign n10401 = pi41 & ~n10400;
  assign n10402 = n6371 & ~n10390;
  assign n10403 = n10388 & n10402;
  assign n10404 = ~pi72 & ~n10403;
  assign n10405 = ~n10393 & n10404;
  assign n10406 = ~n10363 & ~n10405;
  assign n10407 = ~pi101 & ~n10406;
  assign n10408 = n10288 & ~n10407;
  assign n10409 = ~n10401 & ~n10408;
  assign n10410 = ~pi228 & ~n10409;
  assign n10411 = ~pi39 & ~n10410;
  assign n10412 = ~n10370 & n10411;
  assign n10413 = pi287 & n3096;
  assign n10414 = n10310 & n10413;
  assign n10415 = ~n10311 & ~n10414;
  assign n10416 = pi39 & ~n10415;
  assign n10417 = n3207 & ~n10416;
  assign n10418 = ~n10412 & n10417;
  assign n10419 = pi41 & ~n10281;
  assign n10420 = n2498 & n6371;
  assign n10421 = ~pi44 & n10420;
  assign n10422 = n10288 & n10421;
  assign n10423 = ~n10284 & ~n10422;
  assign n10424 = ~pi72 & ~n7547;
  assign n10425 = ~n10423 & ~n10424;
  assign n10426 = ~n10286 & n10425;
  assign n10427 = n2734 & ~n10286;
  assign n10428 = ~n10285 & ~n10427;
  assign n10429 = ~n10419 & ~n10428;
  assign n10430 = ~n10426 & n10429;
  assign n10431 = n10278 & ~n10430;
  assign n10432 = ~n10276 & ~n10431;
  assign n10433 = ~pi39 & ~n10432;
  assign n10434 = ~n10312 & ~n10433;
  assign n10435 = n6251 & ~n10434;
  assign n10436 = pi38 & ~n10316;
  assign n10437 = ~pi87 & ~n10436;
  assign n10438 = ~n10435 & n10437;
  assign n10439 = ~n10418 & n10438;
  assign n10440 = pi41 & ~n10280;
  assign n10441 = pi228 & n10423;
  assign n10442 = ~n10440 & n10441;
  assign n10443 = ~pi228 & n10275;
  assign n10444 = n3208 & ~n10443;
  assign n10445 = ~n10442 & n10444;
  assign n10446 = ~n3207 & n10315;
  assign n10447 = pi87 & ~n10446;
  assign n10448 = ~n10312 & n10447;
  assign n10449 = ~n10445 & n10448;
  assign n10450 = ~pi75 & ~n10449;
  assign n10451 = ~n10439 & n10450;
  assign n10452 = ~n10319 & ~n10451;
  assign n10453 = n7444 & ~n10452;
  assign n10454 = ~n7444 & ~n10316;
  assign n10455 = ~po1038 & ~n10454;
  assign n10456 = ~n10453 & n10455;
  assign n10457 = pi39 & pi232;
  assign n10458 = n10307 & n10457;
  assign n10459 = ~pi72 & ~n10315;
  assign n10460 = po1038 & n10459;
  assign n10461 = ~n10458 & n10460;
  assign po199 = ~n10456 & ~n10461;
  assign n10463 = pi207 & pi208;
  assign n10464 = ~pi115 & n2734;
  assign n10465 = pi42 & ~pi114;
  assign n10466 = pi72 & pi116;
  assign n10467 = pi72 & pi113;
  assign n10468 = pi72 & ~n6253;
  assign n10469 = ~pi99 & n10355;
  assign n10470 = ~n10468 & ~n10469;
  assign n10471 = ~pi113 & ~n10470;
  assign n10472 = ~n10467 & ~n10471;
  assign n10473 = ~pi116 & ~n10472;
  assign n10474 = ~n10466 & ~n10473;
  assign n10475 = n10465 & ~n10474;
  assign n10476 = pi42 & ~pi72;
  assign n10477 = pi114 & ~n10476;
  assign n10478 = n6253 & n10340;
  assign n10479 = n6257 & n10478;
  assign n10480 = ~pi42 & ~n10479;
  assign n10481 = ~n10477 & ~n10480;
  assign n10482 = ~n10475 & n10481;
  assign n10483 = n10464 & ~n10482;
  assign n10484 = ~pi115 & ~n2734;
  assign n10485 = ~pi99 & n10366;
  assign n10486 = ~n10468 & ~n10485;
  assign n10487 = ~pi113 & ~n10486;
  assign n10488 = ~n10467 & ~n10487;
  assign n10489 = ~pi116 & ~n10488;
  assign n10490 = ~n10466 & ~n10489;
  assign n10491 = pi42 & n10490;
  assign n10492 = n6253 & n10360;
  assign n10493 = n6257 & n10492;
  assign n10494 = ~pi42 & n10493;
  assign n10495 = ~pi114 & ~n10494;
  assign n10496 = ~n10491 & n10495;
  assign n10497 = ~n10477 & ~n10496;
  assign n10498 = n10484 & ~n10497;
  assign n10499 = pi115 & ~n10476;
  assign n10500 = pi228 & ~n10499;
  assign n10501 = ~n10498 & n10500;
  assign n10502 = ~n10483 & n10501;
  assign n10503 = ~pi99 & n10408;
  assign n10504 = ~n10468 & ~n10503;
  assign n10505 = ~pi72 & pi113;
  assign n10506 = ~n10504 & ~n10505;
  assign n10507 = ~pi116 & n10506;
  assign n10508 = ~n10466 & ~n10507;
  assign n10509 = n10465 & ~n10508;
  assign n10510 = n6253 & n10400;
  assign n10511 = ~pi113 & n10510;
  assign n10512 = ~pi116 & n10511;
  assign n10513 = ~pi42 & ~n10512;
  assign n10514 = ~n10477 & ~n10513;
  assign n10515 = ~n10509 & n10514;
  assign n10516 = ~pi115 & ~n10515;
  assign n10517 = ~pi228 & ~n10499;
  assign n10518 = ~n10516 & n10517;
  assign n10519 = ~pi39 & ~n10518;
  assign n10520 = ~n10502 & n10519;
  assign n10521 = ~pi72 & ~n10301;
  assign n10522 = n6170 & n10413;
  assign n10523 = ~pi189 & n10522;
  assign n10524 = ~n10521 & ~n10523;
  assign n10525 = pi199 & ~n10524;
  assign n10526 = pi232 & ~pi299;
  assign n10527 = ~n10525 & n10526;
  assign n10528 = n10305 & n10413;
  assign n10529 = ~pi166 & n7484;
  assign n10530 = ~pi72 & ~n10529;
  assign n10531 = pi232 & pi299;
  assign n10532 = ~n10530 & n10531;
  assign n10533 = ~n10528 & n10532;
  assign n10534 = ~pi72 & pi199;
  assign n10535 = ~pi232 & ~n10534;
  assign n10536 = pi72 & ~pi232;
  assign n10537 = pi299 & ~n10536;
  assign n10538 = n10535 & ~n10537;
  assign n10539 = ~n10533 & ~n10538;
  assign n10540 = ~n10527 & n10539;
  assign n10541 = pi39 & ~n10540;
  assign n10542 = ~n10520 & ~n10541;
  assign n10543 = n3207 & ~n10542;
  assign n10544 = ~n8087 & ~n10476;
  assign n10545 = ~n10464 & n10476;
  assign n10546 = n8087 & ~n10545;
  assign n10547 = n10464 & ~n10477;
  assign n10548 = n6253 & n10280;
  assign n10549 = n6257 & n10548;
  assign n10550 = n7547 & n10549;
  assign n10551 = ~pi114 & ~n6256;
  assign n10552 = n10550 & n10551;
  assign n10553 = ~pi42 & n10552;
  assign n10554 = n6254 & n10421;
  assign n10555 = n6257 & n10554;
  assign n10556 = ~pi72 & ~n10555;
  assign n10557 = ~n10424 & ~n10556;
  assign n10558 = pi42 & ~n10557;
  assign n10559 = ~pi114 & ~n10558;
  assign n10560 = ~n10553 & n10559;
  assign n10561 = n10547 & ~n10560;
  assign n10562 = n10546 & ~n10561;
  assign n10563 = ~n10544 & ~n10562;
  assign n10564 = ~pi39 & ~n10563;
  assign n10565 = ~pi299 & ~n10535;
  assign n10566 = pi199 & n10521;
  assign n10567 = pi232 & ~n10566;
  assign n10568 = n10565 & ~n10567;
  assign n10569 = pi299 & n10530;
  assign n10570 = pi39 & ~n10569;
  assign n10571 = ~n10568 & n10570;
  assign n10572 = ~n10564 & ~n10571;
  assign n10573 = n6251 & ~n10572;
  assign n10574 = ~pi39 & ~n10476;
  assign n10575 = ~n10571 & ~n10574;
  assign n10576 = pi38 & ~n10575;
  assign n10577 = ~pi87 & ~n10576;
  assign n10578 = ~n10573 & n10577;
  assign n10579 = ~n10543 & n10578;
  assign n10580 = pi228 & n10549;
  assign n10581 = ~pi115 & n10580;
  assign n10582 = ~pi114 & n10581;
  assign n10583 = ~pi42 & n10582;
  assign n10584 = pi228 & n10554;
  assign n10585 = n6259 & n10584;
  assign n10586 = n10476 & ~n10585;
  assign n10587 = n3208 & ~n10586;
  assign n10588 = ~n10583 & n10587;
  assign n10589 = ~n3207 & n10574;
  assign n10590 = pi87 & ~n10589;
  assign n10591 = ~n10588 & n10590;
  assign n10592 = ~n10571 & n10591;
  assign n10593 = ~pi75 & ~n10592;
  assign n10594 = ~n10579 & n10593;
  assign n10595 = n7487 & n10552;
  assign n10596 = ~pi42 & n10595;
  assign n10597 = n6254 & n10293;
  assign n10598 = ~pi113 & n10597;
  assign n10599 = ~pi116 & n10598;
  assign n10600 = n10476 & ~n10599;
  assign n10601 = ~pi114 & ~n10600;
  assign n10602 = ~n10596 & n10601;
  assign n10603 = n10547 & ~n10602;
  assign n10604 = n10546 & ~n10603;
  assign n10605 = n3242 & ~n10544;
  assign n10606 = ~n10604 & n10605;
  assign n10607 = ~n3242 & n10476;
  assign n10608 = ~pi39 & ~n10607;
  assign n10609 = ~n10606 & n10608;
  assign n10610 = ~n10571 & ~n10609;
  assign n10611 = pi75 & ~n10610;
  assign n10612 = n7444 & ~n10611;
  assign n10613 = ~n10594 & n10612;
  assign n10614 = ~n10463 & ~n10613;
  assign n10615 = ~pi72 & pi200;
  assign n10616 = ~pi232 & ~n10615;
  assign n10617 = ~pi299 & ~n10616;
  assign n10618 = pi200 & n10521;
  assign n10619 = pi232 & ~n10618;
  assign n10620 = n10617 & ~n10619;
  assign n10621 = pi39 & ~n10620;
  assign n10622 = ~n10568 & n10621;
  assign n10623 = ~n10574 & ~n10622;
  assign n10624 = ~n7444 & n10623;
  assign n10625 = n10463 & ~n10624;
  assign n10626 = pi232 & ~n10525;
  assign n10627 = pi200 & ~n10524;
  assign n10628 = n10626 & ~n10627;
  assign n10629 = ~pi299 & n10628;
  assign n10630 = n10538 & ~n10615;
  assign n10631 = ~n10533 & ~n10630;
  assign n10632 = ~n10629 & n10631;
  assign n10633 = pi39 & ~n10632;
  assign n10634 = ~n10520 & ~n10633;
  assign n10635 = n3207 & ~n10634;
  assign n10636 = n10571 & n10621;
  assign n10637 = ~n10564 & ~n10636;
  assign n10638 = n6251 & ~n10637;
  assign n10639 = pi38 & ~n10623;
  assign n10640 = ~pi87 & ~n10639;
  assign n10641 = ~n10577 & ~n10640;
  assign n10642 = ~n10638 & ~n10641;
  assign n10643 = ~n10635 & n10642;
  assign n10644 = n10590 & ~n10636;
  assign n10645 = ~n10588 & n10644;
  assign n10646 = ~pi75 & ~n10645;
  assign n10647 = ~n10643 & n10646;
  assign n10648 = ~n10609 & ~n10636;
  assign n10649 = pi75 & ~n10648;
  assign n10650 = n7444 & ~n10649;
  assign n10651 = ~n10647 & n10650;
  assign n10652 = n10625 & ~n10651;
  assign n10653 = ~n10614 & ~n10652;
  assign n10654 = pi211 & pi214;
  assign n10655 = pi212 & n10654;
  assign n10656 = ~pi219 & ~n10655;
  assign n10657 = ~n7444 & n10575;
  assign n10658 = ~n10656 & ~n10657;
  assign n10659 = ~n10653 & n10658;
  assign n10660 = n10565 & ~n10626;
  assign n10661 = pi39 & ~n10660;
  assign n10662 = ~n10520 & ~n10661;
  assign n10663 = n3207 & ~n10662;
  assign n10664 = pi39 & ~n10568;
  assign n10665 = ~n10564 & ~n10664;
  assign n10666 = n6251 & ~n10665;
  assign n10667 = ~n10574 & ~n10664;
  assign n10668 = pi38 & ~n10667;
  assign n10669 = ~pi87 & ~n10668;
  assign n10670 = ~n10666 & n10669;
  assign n10671 = ~n10663 & n10670;
  assign n10672 = n10591 & ~n10664;
  assign n10673 = ~pi75 & ~n10672;
  assign n10674 = ~n10671 & n10673;
  assign n10675 = ~n10609 & ~n10664;
  assign n10676 = pi75 & ~n10675;
  assign n10677 = n7444 & ~n10676;
  assign n10678 = ~n10674 & n10677;
  assign n10679 = ~n7444 & n10667;
  assign n10680 = ~n10463 & ~n10679;
  assign n10681 = ~n10678 & n10680;
  assign n10682 = ~n10565 & ~n10617;
  assign n10683 = ~n10628 & ~n10682;
  assign n10684 = pi39 & ~n10683;
  assign n10685 = ~n10520 & ~n10684;
  assign n10686 = n3207 & ~n10685;
  assign n10687 = ~n10564 & ~n10622;
  assign n10688 = n6251 & ~n10687;
  assign n10689 = n10640 & ~n10688;
  assign n10690 = ~n10686 & n10689;
  assign n10691 = n10591 & ~n10622;
  assign n10692 = ~pi75 & ~n10691;
  assign n10693 = ~n10690 & n10692;
  assign n10694 = ~n10609 & ~n10622;
  assign n10695 = pi75 & ~n10694;
  assign n10696 = n7444 & ~n10695;
  assign n10697 = ~n10693 & n10696;
  assign n10698 = n10625 & ~n10697;
  assign n10699 = ~n10681 & ~n10698;
  assign n10700 = n10656 & ~n10699;
  assign n10701 = ~po1038 & ~n10659;
  assign n10702 = ~n10700 & n10701;
  assign n10703 = n10530 & ~n10656;
  assign n10704 = pi39 & ~n10703;
  assign n10705 = po1038 & ~n10574;
  assign n10706 = ~n10704 & n10705;
  assign po200 = n10702 | n10706;
  assign n10708 = pi212 & pi214;
  assign n10709 = ~pi211 & ~pi219;
  assign n10710 = n10708 & ~n10709;
  assign n10711 = ~pi211 & ~n10708;
  assign n10712 = ~n10710 & ~n10711;
  assign n10713 = ~n2734 & ~n10490;
  assign n10714 = n2734 & ~n10474;
  assign n10715 = ~n10713 & ~n10714;
  assign n10716 = pi228 & ~n10715;
  assign n10717 = ~pi228 & ~n10508;
  assign n10718 = ~n10716 & ~n10717;
  assign n10719 = ~pi42 & n6258;
  assign n10720 = pi43 & n10719;
  assign n10721 = ~n10718 & n10720;
  assign n10722 = ~pi228 & ~n10512;
  assign n10723 = ~n2734 & ~n10492;
  assign n10724 = n2734 & ~n10478;
  assign n10725 = ~n10723 & ~n10724;
  assign n10726 = n6257 & n10725;
  assign n10727 = pi228 & ~n10726;
  assign n10728 = ~n10722 & ~n10727;
  assign n10729 = ~pi43 & ~n10728;
  assign n10730 = pi43 & ~pi72;
  assign n10731 = ~n10719 & ~n10730;
  assign n10732 = ~n10729 & ~n10731;
  assign n10733 = ~n10721 & n10732;
  assign n10734 = ~pi39 & ~n10733;
  assign n10735 = pi232 & ~n10627;
  assign n10736 = n10617 & ~n10735;
  assign n10737 = pi39 & ~n10736;
  assign n10738 = ~n10734 & ~n10737;
  assign n10739 = n3207 & ~n10738;
  assign n10740 = ~n8087 & ~n10730;
  assign n10741 = n2734 & n10719;
  assign n10742 = n10730 & ~n10741;
  assign n10743 = n8087 & ~n10742;
  assign n10744 = ~pi43 & pi52;
  assign n10745 = n10550 & n10744;
  assign n10746 = pi43 & ~n10557;
  assign n10747 = ~n10745 & ~n10746;
  assign n10748 = n10741 & ~n10747;
  assign n10749 = n10743 & ~n10748;
  assign n10750 = ~n10740 & ~n10749;
  assign n10751 = ~pi39 & ~n10750;
  assign n10752 = ~n10621 & ~n10751;
  assign n10753 = n6251 & ~n10752;
  assign n10754 = ~pi39 & ~n10730;
  assign n10755 = ~n10621 & ~n10754;
  assign n10756 = pi38 & ~n10755;
  assign n10757 = ~pi87 & ~n10756;
  assign n10758 = ~n10753 & n10757;
  assign n10759 = ~n10739 & n10758;
  assign n10760 = ~pi43 & ~n10549;
  assign n10761 = pi43 & ~n10556;
  assign n10762 = pi228 & n10719;
  assign n10763 = ~n10761 & n10762;
  assign n10764 = ~n10760 & n10763;
  assign n10765 = n10730 & ~n10762;
  assign n10766 = n3208 & ~n10765;
  assign n10767 = ~n10764 & n10766;
  assign n10768 = ~n3207 & n10754;
  assign n10769 = pi87 & ~n10768;
  assign n10770 = ~n10767 & n10769;
  assign n10771 = ~n10621 & n10770;
  assign n10772 = ~pi75 & ~n10771;
  assign n10773 = ~n10759 & n10772;
  assign n10774 = ~pi72 & ~n10599;
  assign n10775 = pi43 & n10774;
  assign n10776 = n7487 & n10550;
  assign n10777 = n10744 & n10776;
  assign n10778 = ~n10775 & ~n10777;
  assign n10779 = n10741 & ~n10778;
  assign n10780 = n10743 & ~n10779;
  assign n10781 = ~n10740 & ~n10780;
  assign n10782 = ~pi39 & ~n10781;
  assign n10783 = n3242 & ~n10782;
  assign n10784 = ~n3242 & ~n10754;
  assign n10785 = ~n10783 & ~n10784;
  assign n10786 = ~n10621 & ~n10785;
  assign n10787 = pi75 & ~n10786;
  assign n10788 = n7444 & ~n10787;
  assign n10789 = ~n10773 & n10788;
  assign n10790 = ~n7444 & n10755;
  assign n10791 = ~n10463 & ~n10790;
  assign n10792 = ~n10789 & n10791;
  assign n10793 = ~pi199 & ~pi200;
  assign n10794 = ~pi299 & ~n10793;
  assign n10795 = ~pi72 & ~n10794;
  assign n10796 = ~pi232 & ~n10795;
  assign n10797 = ~pi299 & ~n10796;
  assign n10798 = ~n10524 & n10793;
  assign n10799 = pi232 & ~n10798;
  assign n10800 = n10797 & ~n10799;
  assign n10801 = pi39 & ~n10800;
  assign n10802 = ~n10734 & ~n10801;
  assign n10803 = n3207 & ~n10802;
  assign n10804 = n10521 & n10793;
  assign n10805 = pi232 & ~n10804;
  assign n10806 = n10797 & ~n10805;
  assign n10807 = pi39 & ~n10806;
  assign n10808 = ~n10751 & ~n10807;
  assign n10809 = n6251 & ~n10808;
  assign n10810 = ~n10754 & ~n10807;
  assign n10811 = pi38 & ~n10810;
  assign n10812 = ~pi87 & ~n10811;
  assign n10813 = ~n10809 & n10812;
  assign n10814 = ~n10803 & n10813;
  assign n10815 = ~n3277 & ~n10810;
  assign n10816 = n10770 & ~n10815;
  assign n10817 = ~pi75 & ~n10816;
  assign n10818 = ~n10814 & n10817;
  assign n10819 = ~n10785 & ~n10807;
  assign n10820 = pi75 & ~n10819;
  assign n10821 = n7444 & ~n10820;
  assign n10822 = ~n10818 & n10821;
  assign n10823 = ~n7444 & n10810;
  assign n10824 = n10463 & ~n10823;
  assign n10825 = ~n10822 & n10824;
  assign n10826 = ~n10792 & ~n10825;
  assign n10827 = ~n10712 & ~n10826;
  assign n10828 = n10526 & ~n10627;
  assign n10829 = ~n10537 & n10616;
  assign n10830 = ~n10533 & ~n10829;
  assign n10831 = ~n10828 & n10830;
  assign n10832 = pi39 & ~n10831;
  assign n10833 = ~n10734 & ~n10832;
  assign n10834 = n3207 & ~n10833;
  assign n10835 = n10570 & ~n10620;
  assign n10836 = ~n10751 & ~n10835;
  assign n10837 = n6251 & ~n10836;
  assign n10838 = ~n10754 & ~n10835;
  assign n10839 = pi38 & ~n10838;
  assign n10840 = ~pi87 & ~n10839;
  assign n10841 = ~n10837 & n10840;
  assign n10842 = ~n10834 & n10841;
  assign n10843 = n10770 & ~n10835;
  assign n10844 = ~pi75 & ~n10843;
  assign n10845 = ~n10842 & n10844;
  assign n10846 = ~n10785 & ~n10835;
  assign n10847 = pi75 & ~n10846;
  assign n10848 = n7444 & ~n10847;
  assign n10849 = ~n10845 & n10848;
  assign n10850 = ~n7444 & n10838;
  assign n10851 = ~n10463 & ~n10850;
  assign n10852 = ~n10849 & n10851;
  assign n10853 = n10526 & ~n10798;
  assign n10854 = ~n10533 & ~n10796;
  assign n10855 = ~n10853 & n10854;
  assign n10856 = pi39 & ~n10855;
  assign n10857 = ~n10734 & ~n10856;
  assign n10858 = n3207 & ~n10857;
  assign n10859 = ~n10569 & n10807;
  assign n10860 = ~n10751 & ~n10859;
  assign n10861 = n6251 & ~n10860;
  assign n10862 = ~n10754 & ~n10859;
  assign n10863 = pi38 & ~n10862;
  assign n10864 = ~pi87 & ~n10863;
  assign n10865 = ~n10861 & n10864;
  assign n10866 = ~n10858 & n10865;
  assign n10867 = n10770 & ~n10859;
  assign n10868 = ~pi75 & ~n10867;
  assign n10869 = ~n10866 & n10868;
  assign n10870 = ~n10785 & ~n10859;
  assign n10871 = pi75 & ~n10870;
  assign n10872 = n7444 & ~n10871;
  assign n10873 = ~n10869 & n10872;
  assign n10874 = ~n7444 & n10862;
  assign n10875 = n10463 & ~n10874;
  assign n10876 = ~n10873 & n10875;
  assign n10877 = ~n10852 & ~n10876;
  assign n10878 = n10712 & ~n10877;
  assign n10879 = ~po1038 & ~n10827;
  assign n10880 = ~n10878 & n10879;
  assign n10881 = n10530 & n10712;
  assign n10882 = pi39 & ~n10881;
  assign n10883 = po1038 & ~n10754;
  assign n10884 = ~n10882 & n10883;
  assign po201 = n10880 | n10884;
  assign n10886 = ~n8087 & ~n10363;
  assign n10887 = ~pi39 & ~n10886;
  assign n10888 = ~n2734 & n10363;
  assign n10889 = n8087 & ~n10888;
  assign n10890 = n7489 & ~n10342;
  assign n10891 = n7547 & n10279;
  assign n10892 = n7487 & n10891;
  assign n10893 = pi44 & ~n10292;
  assign n10894 = ~n10892 & ~n10893;
  assign n10895 = n10890 & ~n10894;
  assign n10896 = n10889 & ~n10895;
  assign n10897 = n10887 & ~n10896;
  assign n10898 = pi39 & n7485;
  assign n10899 = ~pi72 & n10898;
  assign n10900 = ~n10897 & ~n10899;
  assign n10901 = n3242 & ~n10900;
  assign n10902 = ~pi39 & ~n10363;
  assign n10903 = pi39 & ~n10899;
  assign n10904 = ~n10902 & ~n10903;
  assign n10905 = ~n3242 & n10904;
  assign n10906 = pi75 & ~n10905;
  assign n10907 = ~n10901 & n10906;
  assign n10908 = pi44 & n10351;
  assign n10909 = n2734 & ~n10339;
  assign n10910 = ~n10908 & n10909;
  assign n10911 = pi44 & n10362;
  assign n10912 = ~n2734 & ~n10359;
  assign n10913 = ~n10911 & n10912;
  assign n10914 = ~n10910 & ~n10913;
  assign n10915 = pi228 & ~n10914;
  assign n10916 = pi44 & n10405;
  assign n10917 = ~pi228 & ~n10916;
  assign n10918 = ~n10399 & n10917;
  assign n10919 = ~pi39 & ~n10918;
  assign n10920 = ~n10915 & n10919;
  assign n10921 = pi287 & n10420;
  assign n10922 = ~pi72 & ~n10921;
  assign n10923 = n10898 & n10922;
  assign n10924 = n3207 & ~n10923;
  assign n10925 = ~n10920 & n10924;
  assign n10926 = n7547 & n10420;
  assign n10927 = pi44 & ~n10926;
  assign n10928 = ~n10891 & ~n10927;
  assign n10929 = n10890 & ~n10928;
  assign n10930 = n10889 & ~n10929;
  assign n10931 = n10887 & ~n10930;
  assign n10932 = n6251 & ~n10899;
  assign n10933 = ~n10931 & n10932;
  assign n10934 = pi38 & ~n10904;
  assign n10935 = ~pi87 & ~n10934;
  assign n10936 = ~n10933 & n10935;
  assign n10937 = ~n10925 & n10936;
  assign n10938 = pi228 & n3207;
  assign n10939 = n10279 & n10938;
  assign n10940 = n10420 & n10938;
  assign n10941 = n10363 & ~n10940;
  assign n10942 = ~pi39 & ~n10941;
  assign n10943 = ~n10939 & n10942;
  assign n10944 = pi87 & ~n10903;
  assign n10945 = ~n10943 & n10944;
  assign n10946 = ~pi75 & ~n10945;
  assign n10947 = ~n10937 & n10946;
  assign n10948 = ~n10907 & ~n10947;
  assign n10949 = n7444 & ~n10948;
  assign n10950 = ~n7444 & ~n10904;
  assign n10951 = ~po1038 & ~n10950;
  assign n10952 = ~n10949 & n10951;
  assign n10953 = n2448 & n7484;
  assign n10954 = ~pi72 & n10953;
  assign n10955 = pi39 & ~n10954;
  assign n10956 = po1038 & ~n10902;
  assign n10957 = ~n10955 & n10956;
  assign po202 = n10952 | n10957;
  assign n10959 = ~pi38 & pi39;
  assign n10960 = n10178 & n10959;
  assign n10961 = pi979 & n10960;
  assign po203 = n6443 & n10961;
  assign n10963 = ~pi102 & ~pi104;
  assign n10964 = ~pi111 & n10963;
  assign n10965 = ~pi49 & ~pi76;
  assign n10966 = n8895 & n10965;
  assign n10967 = pi61 & ~pi82;
  assign n10968 = ~pi83 & ~pi89;
  assign n10969 = n10967 & n10968;
  assign n10970 = n7451 & n8905;
  assign n10971 = n10969 & n10970;
  assign n10972 = n10155 & n10964;
  assign n10973 = n10966 & n10972;
  assign n10974 = n8903 & n10971;
  assign n10975 = n10221 & n10974;
  assign n10976 = n10973 & n10975;
  assign n10977 = n8918 & n10976;
  assign n10978 = ~pi841 & n10977;
  assign n10979 = n2491 & n2698;
  assign n10980 = pi24 & n10979;
  assign n10981 = ~n10978 & ~n10980;
  assign po204 = n10147 & ~n10981;
  assign n10983 = ~n2680 & n7451;
  assign n10984 = ~pi82 & n2463;
  assign n10985 = ~pi84 & pi104;
  assign n10986 = n2607 & n10985;
  assign n10987 = n10159 & n10986;
  assign n10988 = n10984 & n10987;
  assign n10989 = ~pi36 & ~n10988;
  assign n10990 = n8904 & n9025;
  assign n10991 = ~pi67 & ~pi103;
  assign n10992 = n2476 & n10991;
  assign n10993 = ~pi98 & n10992;
  assign n10994 = n10990 & n10993;
  assign n10995 = ~n10989 & n10994;
  assign n10996 = ~n2648 & n10995;
  assign n10997 = ~pi88 & ~n10996;
  assign n10998 = n2532 & ~n10997;
  assign n10999 = n10983 & n10998;
  assign n11000 = n2489 & n10999;
  assign n11001 = ~n10140 & ~n11000;
  assign n11002 = n10143 & ~n11001;
  assign n11003 = n7560 & ~n11002;
  assign n11004 = ~n6265 & n11002;
  assign n11005 = ~pi36 & n10995;
  assign n11006 = ~pi88 & ~n11005;
  assign n11007 = n10983 & ~n11006;
  assign n11008 = n10171 & n11007;
  assign n11009 = ~pi824 & n6265;
  assign n11010 = n11008 & n11009;
  assign n11011 = pi829 & ~n11010;
  assign n11012 = ~n11004 & n11011;
  assign n11013 = ~n2733 & n11012;
  assign n11014 = ~n11003 & ~n11013;
  assign n11015 = pi1091 & ~n11014;
  assign n11016 = ~n7496 & n11002;
  assign n11017 = ~pi829 & ~n11016;
  assign n11018 = ~n11012 & ~n11017;
  assign n11019 = ~pi1093 & ~n11018;
  assign n11020 = n7496 & n10143;
  assign n11021 = ~n10141 & n11020;
  assign n11022 = ~n6457 & ~n7558;
  assign n11023 = ~n11021 & ~n11022;
  assign n11024 = ~n11016 & n11023;
  assign n11025 = n10146 & ~n11024;
  assign n11026 = ~n11019 & n11025;
  assign po205 = ~n11015 & n11026;
  assign n11028 = ~pi72 & pi841;
  assign n11029 = n2494 & n11028;
  assign n11030 = ~pi51 & n11029;
  assign n11031 = n10230 & n11030;
  assign n11032 = n10146 & n11031;
  assign po206 = n10170 & n11032;
  assign n11034 = pi74 & ~n8948;
  assign n11035 = n2453 & n2476;
  assign n11036 = ~pi103 & n2641;
  assign n11037 = n10219 & n11036;
  assign n11038 = n8895 & n8904;
  assign n11039 = n11037 & n11038;
  assign n11040 = ~pi45 & pi49;
  assign n11041 = n10964 & n11040;
  assign n11042 = n11035 & n11041;
  assign n11043 = n11039 & n11042;
  assign n11044 = n10984 & n11043;
  assign n11045 = n2495 & n8918;
  assign n11046 = n11044 & n11045;
  assign n11047 = n10142 & n11029;
  assign n11048 = n11046 & n11047;
  assign n11049 = ~pi74 & ~n11048;
  assign n11050 = n7380 & ~po1038;
  assign n11051 = ~n11049 & n11050;
  assign po207 = ~n11034 & n11051;
  assign n11053 = pi24 & n8885;
  assign n11054 = ~n10372 & ~n11053;
  assign n11055 = pi24 & ~pi94;
  assign n11056 = ~n8883 & n11055;
  assign n11057 = ~pi252 & ~n8874;
  assign n11058 = pi252 & ~po840;
  assign n11059 = ~n11057 & ~n11058;
  assign n11060 = n10143 & n11059;
  assign n11061 = ~n11056 & n11060;
  assign n11062 = ~n11054 & n11061;
  assign n11063 = n2536 & n7464;
  assign n11064 = pi24 & ~pi90;
  assign n11065 = n11063 & n11064;
  assign n11066 = ~n11059 & n11065;
  assign n11067 = n8887 & n11066;
  assign n11068 = ~n11062 & ~n11067;
  assign n11069 = ~pi100 & ~n11068;
  assign n11070 = pi100 & n6248;
  assign n11071 = n6494 & n11070;
  assign n11072 = ~n11069 & ~n11071;
  assign n11073 = n3182 & n3231;
  assign n11074 = ~n11072 & n11073;
  assign n11075 = n6271 & n8953;
  assign n11076 = n8949 & n11075;
  assign n11077 = ~n11074 & ~n11076;
  assign po208 = n8867 & ~n11077;
  assign n11079 = n2489 & n10147;
  assign n11080 = n2532 & n11079;
  assign n11081 = n9026 & n11035;
  assign n11082 = n2456 & n11081;
  assign n11083 = ~pi69 & n11082;
  assign n11084 = n2641 & n11083;
  assign n11085 = n2643 & n11084;
  assign po209 = n11080 & n11085;
  assign n11087 = ~pi219 & n10711;
  assign n11088 = pi52 & ~pi72;
  assign n11089 = ~pi39 & n11088;
  assign n11090 = pi38 & ~n11089;
  assign n11091 = n6255 & n6258;
  assign n11092 = pi228 & n11091;
  assign n11093 = ~pi52 & n10549;
  assign n11094 = pi52 & n10556;
  assign n11095 = ~n11093 & ~n11094;
  assign n11096 = n11092 & ~n11095;
  assign n11097 = n11088 & ~n11092;
  assign n11098 = ~n11096 & ~n11097;
  assign n11099 = ~pi38 & n11098;
  assign n11100 = ~n11090 & ~n11099;
  assign n11101 = ~pi100 & ~n11100;
  assign n11102 = pi100 & ~n11089;
  assign n11103 = ~pi100 & n10959;
  assign n11104 = pi87 & ~n11103;
  assign n11105 = ~n11102 & n11104;
  assign n11106 = ~n11101 & n11105;
  assign n11107 = ~pi114 & n6255;
  assign n11108 = pi52 & n10474;
  assign n11109 = ~pi52 & n10479;
  assign n11110 = n10464 & ~n11109;
  assign n11111 = ~n11108 & n11110;
  assign n11112 = pi52 & n10490;
  assign n11113 = ~pi52 & n10493;
  assign n11114 = n10484 & ~n11113;
  assign n11115 = ~n11112 & n11114;
  assign n11116 = ~n11111 & ~n11115;
  assign n11117 = n11107 & ~n11116;
  assign n11118 = ~n11088 & ~n11091;
  assign n11119 = pi228 & ~n11118;
  assign n11120 = ~n11117 & n11119;
  assign n11121 = pi52 & n10508;
  assign n11122 = ~pi52 & n10512;
  assign n11123 = n11091 & ~n11122;
  assign n11124 = ~n11121 & n11123;
  assign n11125 = ~pi228 & ~n11118;
  assign n11126 = ~n11124 & n11125;
  assign n11127 = ~pi39 & ~n11126;
  assign n11128 = ~n11120 & n11127;
  assign n11129 = ~pi100 & n11128;
  assign n11130 = n8087 & n10464;
  assign n11131 = n11107 & n11130;
  assign n11132 = n7547 & n11131;
  assign n11133 = n10555 & n11132;
  assign n11134 = n11088 & ~n11133;
  assign n11135 = pi100 & ~n11134;
  assign n11136 = ~pi39 & ~n11135;
  assign n11137 = ~n11129 & n11136;
  assign n11138 = ~pi38 & ~n11137;
  assign n11139 = ~pi87 & ~n11090;
  assign n11140 = ~n11138 & n11139;
  assign n11141 = ~n11106 & ~n11140;
  assign n11142 = ~pi75 & ~n11141;
  assign n11143 = n10599 & n11131;
  assign n11144 = n3242 & n11143;
  assign n11145 = n11089 & ~n11144;
  assign n11146 = pi75 & n11145;
  assign n11147 = n7444 & ~n11146;
  assign n11148 = ~n11142 & n11147;
  assign n11149 = ~n7444 & ~n11089;
  assign n11150 = n10463 & ~n11149;
  assign n11151 = ~n11148 & n11150;
  assign n11152 = ~n10801 & ~n11128;
  assign n11153 = n3207 & ~n11152;
  assign n11154 = ~pi39 & ~n11134;
  assign n11155 = ~n10807 & ~n11154;
  assign n11156 = n6251 & ~n11155;
  assign n11157 = ~pi39 & ~n11088;
  assign n11158 = ~n10807 & ~n11157;
  assign n11159 = pi38 & ~n11158;
  assign n11160 = ~pi87 & ~n11159;
  assign n11161 = ~n11156 & n11160;
  assign n11162 = ~n11153 & n11161;
  assign n11163 = ~n3207 & n11158;
  assign n11164 = ~pi39 & n11098;
  assign n11165 = n3207 & ~n10807;
  assign n11166 = ~n11164 & n11165;
  assign n11167 = ~n11163 & ~n11166;
  assign n11168 = pi87 & ~n11167;
  assign n11169 = ~pi75 & ~n11168;
  assign n11170 = ~n11162 & n11169;
  assign n11171 = n11088 & ~n11143;
  assign n11172 = ~pi39 & ~n11171;
  assign n11173 = n3242 & ~n10807;
  assign n11174 = ~n11172 & n11173;
  assign n11175 = ~n3242 & n11158;
  assign n11176 = pi75 & ~n11175;
  assign n11177 = ~n11174 & n11176;
  assign n11178 = n7444 & ~n10463;
  assign n11179 = ~n11177 & n11178;
  assign n11180 = ~n11170 & n11179;
  assign n11181 = ~n11151 & ~n11180;
  assign n11182 = ~n11087 & ~n11181;
  assign n11183 = ~n10533 & n10537;
  assign n11184 = pi39 & ~n11183;
  assign n11185 = ~n11128 & ~n11184;
  assign n11186 = n3207 & ~n11185;
  assign n11187 = ~n10570 & ~n11157;
  assign n11188 = pi38 & ~n11187;
  assign n11189 = ~n10570 & ~n11154;
  assign n11190 = n6251 & ~n11189;
  assign n11191 = ~n11188 & ~n11190;
  assign n11192 = ~n11186 & n11191;
  assign n11193 = ~pi87 & ~n11192;
  assign n11194 = ~n3207 & n11187;
  assign n11195 = pi87 & ~n11194;
  assign n11196 = n3207 & ~n10570;
  assign n11197 = ~n11164 & n11196;
  assign n11198 = n11195 & ~n11197;
  assign n11199 = n10463 & ~n11198;
  assign n11200 = ~n11193 & n11199;
  assign n11201 = ~n10856 & ~n11128;
  assign n11202 = n3207 & ~n11201;
  assign n11203 = ~n10859 & ~n11154;
  assign n11204 = n6251 & ~n11203;
  assign n11205 = n11159 & ~n11187;
  assign n11206 = ~n11204 & ~n11205;
  assign n11207 = ~n11202 & n11206;
  assign n11208 = ~pi87 & ~n11207;
  assign n11209 = n3207 & ~n10859;
  assign n11210 = ~n11164 & n11209;
  assign n11211 = ~n11163 & n11195;
  assign n11212 = ~n11210 & n11211;
  assign n11213 = ~n10463 & ~n11212;
  assign n11214 = ~n11208 & n11213;
  assign n11215 = ~n11200 & ~n11214;
  assign n11216 = ~pi75 & ~n11215;
  assign n11217 = ~pi39 & ~n11145;
  assign n11218 = ~n10463 & n10859;
  assign n11219 = n10463 & n10570;
  assign n11220 = pi75 & ~n11219;
  assign n11221 = ~n11218 & n11220;
  assign n11222 = ~n11217 & n11221;
  assign n11223 = n7444 & ~n11222;
  assign n11224 = ~n11216 & n11223;
  assign n11225 = ~n7444 & ~n11187;
  assign n11226 = n11087 & ~n11225;
  assign n11227 = ~n11224 & n11226;
  assign n11228 = ~n7444 & ~n10463;
  assign n11229 = n11158 & n11228;
  assign n11230 = ~po1038 & ~n11229;
  assign n11231 = ~n11227 & n11230;
  assign n11232 = ~n11182 & n11231;
  assign n11233 = pi39 & n11087;
  assign n11234 = n10530 & n11233;
  assign n11235 = po1038 & ~n11089;
  assign n11236 = ~n11234 & n11235;
  assign po210 = ~n11232 & ~n11236;
  assign n11238 = pi24 & n10143;
  assign n11239 = pi53 & n2505;
  assign n11240 = n2514 & n11239;
  assign n11241 = n2506 & n11240;
  assign n11242 = n11238 & n11241;
  assign n11243 = ~pi39 & ~n11242;
  assign n11244 = ~pi287 & ~pi979;
  assign n11245 = n6171 & n11244;
  assign n11246 = pi39 & ~n11245;
  assign n11247 = n10181 & ~n11246;
  assign n11248 = ~n11243 & n11247;
  assign po211 = ~n3353 & n11248;
  assign n11250 = n3243 & n10152;
  assign n11251 = pi54 & ~n11250;
  assign n11252 = n8885 & n9031;
  assign n11253 = ~pi60 & ~pi85;
  assign n11254 = pi106 & n11253;
  assign n11255 = n2468 & n8897;
  assign n11256 = n11254 & n11255;
  assign n11257 = n10966 & n11256;
  assign n11258 = n8908 & n11037;
  assign n11259 = n11257 & n11258;
  assign n11260 = n11035 & n11259;
  assign n11261 = n11252 & n11260;
  assign n11262 = ~pi841 & n2493;
  assign n11263 = n8946 & n11262;
  assign n11264 = n2495 & n3239;
  assign n11265 = n11263 & n11264;
  assign n11266 = n11261 & n11265;
  assign n11267 = ~pi54 & ~n11266;
  assign n11268 = n8866 & ~n11267;
  assign po212 = ~n11251 & n11268;
  assign n11270 = ~pi54 & n11250;
  assign n11271 = ~pi74 & n11270;
  assign n11272 = pi55 & ~n11271;
  assign n11273 = pi45 & n2468;
  assign n11274 = n2476 & n11273;
  assign n11275 = n11039 & n11274;
  assign n11276 = n2465 & n11275;
  assign n11277 = n6371 & n9272;
  assign n11278 = n2454 & n3269;
  assign n11279 = n11277 & n11278;
  assign n11280 = n11276 & n11279;
  assign n11281 = ~pi55 & ~n11280;
  assign n11282 = n8864 & ~n11281;
  assign po213 = ~n11272 & n11282;
  assign n11284 = pi56 & ~pi62;
  assign n11285 = pi55 & n10123;
  assign n11286 = ~n11284 & ~n11285;
  assign n11287 = n3093 & n3281;
  assign n11288 = n6154 & n11287;
  assign n11289 = pi56 & ~n11288;
  assign n11290 = n3432 & ~n11289;
  assign po214 = ~n11286 & n11290;
  assign n11292 = n6293 & n11271;
  assign n11293 = pi57 & ~n11292;
  assign n11294 = n6377 & n11287;
  assign n11295 = ~pi56 & pi62;
  assign n11296 = ~pi924 & n11295;
  assign n11297 = ~n11284 & ~n11296;
  assign n11298 = n11294 & ~n11297;
  assign n11299 = ~pi57 & ~n11298;
  assign n11300 = ~pi59 & ~n11293;
  assign po215 = ~n11299 & n11300;
  assign n11302 = ~pi93 & n11063;
  assign n11303 = n10146 & n11302;
  assign po216 = n7447 & n11303;
  assign n11305 = pi59 & ~n11292;
  assign n11306 = pi924 & n11295;
  assign n11307 = n11294 & n11306;
  assign n11308 = ~pi59 & ~n11307;
  assign n11309 = ~pi57 & ~n11305;
  assign po217 = ~n11308 & n11309;
  assign n11311 = pi39 & ~pi979;
  assign n11312 = ~n6171 & n11311;
  assign n11313 = n6172 & n11312;
  assign n11314 = n6443 & n11313;
  assign n11315 = ~pi39 & n11238;
  assign n11316 = n11252 & n11315;
  assign n11317 = n2503 & n11316;
  assign n11318 = ~n11314 & ~n11317;
  assign po218 = n10181 & ~n11318;
  assign n11320 = pi841 & n10977;
  assign n11321 = ~pi24 & n11252;
  assign n11322 = n2503 & n11321;
  assign n11323 = ~n11320 & ~n11322;
  assign po219 = n10147 & ~n11323;
  assign n11325 = pi57 & ~n10124;
  assign n11326 = n11288 & n11295;
  assign n11327 = ~pi57 & ~n11326;
  assign n11328 = ~pi59 & ~n11325;
  assign po220 = ~n11327 & n11328;
  assign n11330 = n2671 & n8918;
  assign n11331 = n9028 & n11330;
  assign n11332 = pi999 & n11331;
  assign n11333 = ~pi24 & n10979;
  assign n11334 = ~n11332 & ~n11333;
  assign po221 = n10147 & ~n11334;
  assign n11336 = ~pi64 & ~n2663;
  assign n11337 = n2454 & ~n11336;
  assign n11338 = n10154 & n11337;
  assign n11339 = pi841 & ~n11338;
  assign n11340 = n2662 & n9028;
  assign n11341 = ~pi841 & ~n11340;
  assign n11342 = n11080 & ~n11341;
  assign po222 = ~n11339 & n11342;
  assign n11344 = pi39 & n10205;
  assign n11345 = n10181 & n11344;
  assign n11346 = ~n10197 & n11345;
  assign po223 = ~n10203 & n11346;
  assign n11348 = ~pi199 & ~pi299;
  assign n11349 = pi314 & n2453;
  assign n11350 = n11277 & n11349;
  assign n11351 = pi81 & ~pi102;
  assign n11352 = n11350 & n11351;
  assign n11353 = n2478 & n11352;
  assign n11354 = n3269 & n11353;
  assign n11355 = ~n11348 & n11354;
  assign n11356 = pi219 & ~n11355;
  assign n11357 = n3207 & n3267;
  assign n11358 = pi199 & ~pi299;
  assign n11359 = n3222 & n11358;
  assign n11360 = n11357 & n11359;
  assign n11361 = n11353 & n11360;
  assign n11362 = ~pi219 & ~n11361;
  assign n11363 = ~po1038 & ~n11362;
  assign po224 = ~n11356 & n11363;
  assign n11365 = pi83 & ~pi103;
  assign n11366 = n11081 & n11365;
  assign n11367 = n10146 & n11366;
  assign n11368 = n11350 & n11367;
  assign po225 = n2473 & n11368;
  assign n11370 = ~n6229 & n6459;
  assign n11371 = n3325 & n5774;
  assign n11372 = n11370 & n11371;
  assign n11373 = ~n6208 & n6459;
  assign n11374 = n3305 & n3483;
  assign n11375 = n11373 & n11374;
  assign n11376 = ~n11372 & ~n11375;
  assign po226 = n10960 & ~n11376;
  assign n11378 = pi69 & n11036;
  assign n11379 = n10129 & n11378;
  assign n11380 = ~pi71 & ~n11379;
  assign n11381 = ~pi81 & ~pi314;
  assign n11382 = n2454 & n11381;
  assign n11383 = n6328 & n11382;
  assign n11384 = ~n11380 & n11383;
  assign n11385 = pi71 & pi314;
  assign n11386 = n7451 & n11385;
  assign n11387 = n10132 & n11386;
  assign n11388 = n2474 & n11387;
  assign n11389 = ~n11384 & ~n11388;
  assign po227 = n11080 & ~n11389;
  assign n11391 = n2548 & n2560;
  assign n11392 = ~pi96 & n11391;
  assign n11393 = n10151 & n11392;
  assign n11394 = pi198 & pi589;
  assign n11395 = n3484 & ~n6208;
  assign n11396 = n11394 & n11395;
  assign n11397 = pi210 & pi589;
  assign n11398 = ~pi221 & n5774;
  assign n11399 = ~pi216 & n11398;
  assign n11400 = ~n6229 & n11399;
  assign n11401 = n11397 & n11400;
  assign n11402 = ~n11396 & ~n11401;
  assign n11403 = ~pi593 & n6444;
  assign n11404 = ~n6452 & n11403;
  assign n11405 = ~n11402 & n11404;
  assign n11406 = ~pi287 & ~n11405;
  assign n11407 = pi39 & ~n11406;
  assign n11408 = n3096 & n11407;
  assign n11409 = ~n11393 & ~n11408;
  assign po228 = n10181 & ~n11409;
  assign n11411 = ~pi50 & n8918;
  assign n11412 = n6334 & n11411;
  assign n11413 = n2458 & n2470;
  assign n11414 = n6313 & n11413;
  assign n11415 = n10992 & n11414;
  assign n11416 = ~pi64 & n8904;
  assign n11417 = n11415 & n11416;
  assign n11418 = ~pi81 & ~n11417;
  assign n11419 = ~pi199 & pi200;
  assign n11420 = ~pi299 & n11419;
  assign n11421 = pi211 & ~pi219;
  assign n11422 = pi299 & n11421;
  assign n11423 = ~n11420 & ~n11422;
  assign n11424 = pi314 & ~n11423;
  assign n11425 = n10143 & n11424;
  assign n11426 = ~n11418 & n11425;
  assign n11427 = n11412 & n11426;
  assign n11428 = n10990 & n11423;
  assign n11429 = n11350 & n11428;
  assign n11430 = n11415 & n11429;
  assign n11431 = ~n11427 & ~n11430;
  assign po229 = n10146 & ~n11431;
  assign n11433 = pi24 & n2498;
  assign n11434 = pi72 & n11433;
  assign n11435 = pi88 & n10128;
  assign n11436 = n6451 & n9154;
  assign n11437 = n11435 & n11436;
  assign n11438 = n2679 & n11437;
  assign n11439 = ~n11434 & ~n11438;
  assign n11440 = n6371 & ~n11439;
  assign n11441 = ~pi39 & ~n11440;
  assign n11442 = n7532 & n11370;
  assign n11443 = n7536 & n11373;
  assign n11444 = pi39 & ~n11442;
  assign n11445 = ~n11443 & n11444;
  assign n11446 = n10181 & ~n11445;
  assign po230 = ~n11441 & n11446;
  assign n11448 = n9044 & n11373;
  assign n11449 = ~pi299 & ~n11448;
  assign n11450 = n9055 & n11370;
  assign n11451 = pi299 & ~n11450;
  assign n11452 = ~n11449 & ~n11451;
  assign n11453 = pi39 & ~n11452;
  assign n11454 = ~pi314 & pi1050;
  assign n11455 = n9562 & n10143;
  assign n11456 = n11454 & n11455;
  assign n11457 = ~pi39 & ~n11456;
  assign n11458 = n10181 & ~n11457;
  assign po231 = ~n11453 & n11458;
  assign n11460 = pi74 & n11270;
  assign n11461 = n2538 & n7505;
  assign n11462 = ~pi96 & ~n11461;
  assign n11463 = ~pi96 & ~pi1093;
  assign n11464 = n7496 & n11463;
  assign n11465 = ~pi96 & ~n6151;
  assign n11466 = pi479 & ~n11465;
  assign n11467 = n3409 & n7444;
  assign n11468 = ~n11464 & n11467;
  assign n11469 = ~po840 & ~n11466;
  assign n11470 = n11468 & n11469;
  assign n11471 = ~n11462 & n11470;
  assign n11472 = n7469 & n11471;
  assign n11473 = ~n11460 & ~n11472;
  assign po232 = ~po1038 & ~n11473;
  assign n11475 = pi96 & ~pi1093;
  assign n11476 = ~n2733 & n10053;
  assign n11477 = ~n11462 & n11476;
  assign n11478 = ~n11475 & ~n11477;
  assign n11479 = n3223 & ~n11478;
  assign n11480 = n7514 & n11479;
  assign n11481 = ~pi75 & ~n11480;
  assign n11482 = n3242 & n10152;
  assign n11483 = pi75 & ~n11482;
  assign n11484 = n8867 & ~n11483;
  assign po233 = ~n11481 & n11484;
  assign n11486 = n3094 & n10373;
  assign n11487 = pi252 & n7513;
  assign n11488 = n11486 & ~n11487;
  assign n11489 = ~pi137 & n11488;
  assign n11490 = ~pi137 & n2734;
  assign n11491 = ~n8885 & ~n10372;
  assign n11492 = ~pi94 & ~n8921;
  assign n11493 = n10143 & ~n11492;
  assign n11494 = ~n11491 & n11493;
  assign n11495 = ~n7513 & ~n11494;
  assign n11496 = ~pi252 & n11494;
  assign n11497 = n8916 & n10171;
  assign n11498 = pi252 & n11497;
  assign n11499 = n7513 & ~n11498;
  assign n11500 = ~n11496 & n11499;
  assign n11501 = ~n11495 & ~n11500;
  assign n11502 = pi122 & ~n11501;
  assign n11503 = n7496 & n11495;
  assign n11504 = ~n6266 & ~n11486;
  assign n11505 = ~n11500 & ~n11504;
  assign n11506 = ~n11503 & n11505;
  assign n11507 = ~pi122 & ~n11506;
  assign n11508 = ~n11502 & ~n11507;
  assign n11509 = ~pi1093 & ~n11508;
  assign n11510 = ~pi122 & ~n11488;
  assign n11511 = ~n11502 & ~n11510;
  assign n11512 = pi1093 & ~n11511;
  assign n11513 = ~n11509 & ~n11512;
  assign n11514 = n2734 & ~n11513;
  assign n11515 = ~n11490 & ~n11514;
  assign n11516 = ~n11489 & ~n11515;
  assign n11517 = ~pi122 & n11486;
  assign n11518 = pi1093 & ~n11494;
  assign n11519 = ~n8038 & ~n11518;
  assign n11520 = ~n11517 & ~n11519;
  assign n11521 = ~n11509 & ~n11520;
  assign n11522 = ~n2734 & ~n11521;
  assign n11523 = ~pi137 & ~n2734;
  assign n11524 = ~n11522 & ~n11523;
  assign n11525 = pi252 & pi1092;
  assign n11526 = ~pi1093 & n11525;
  assign n11527 = n2754 & n11526;
  assign n11528 = ~pi137 & ~n11527;
  assign n11529 = n11486 & n11528;
  assign n11530 = ~n11524 & ~n11529;
  assign n11531 = ~n11516 & ~n11530;
  assign n11532 = ~po1057 & ~n11531;
  assign n11533 = ~n10086 & n11497;
  assign n11534 = po1057 & ~n11533;
  assign n11535 = ~pi137 & po1057;
  assign n11536 = ~n11534 & ~n11535;
  assign n11537 = ~n11532 & n11536;
  assign n11538 = ~pi210 & ~n11537;
  assign n11539 = ~n11514 & ~n11522;
  assign n11540 = ~po1057 & ~n11539;
  assign n11541 = ~n11534 & ~n11540;
  assign n11542 = pi210 & ~n11541;
  assign n11543 = ~n11538 & ~n11542;
  assign n11544 = n2447 & n10305;
  assign n11545 = ~n11543 & ~n11544;
  assign n11546 = ~pi210 & ~n11531;
  assign n11547 = pi210 & ~n11539;
  assign n11548 = ~n11546 & ~n11547;
  assign n11549 = n11544 & ~n11548;
  assign n11550 = pi299 & ~n11549;
  assign n11551 = ~n11545 & n11550;
  assign n11552 = ~pi198 & ~n11537;
  assign n11553 = pi198 & ~n11541;
  assign n11554 = ~n11552 & ~n11553;
  assign n11555 = n3064 & n6170;
  assign n11556 = ~n11554 & ~n11555;
  assign n11557 = pi198 & ~n11539;
  assign n11558 = ~pi198 & ~n11531;
  assign n11559 = ~n11557 & ~n11558;
  assign n11560 = n11555 & ~n11559;
  assign n11561 = ~pi299 & ~n11560;
  assign n11562 = ~n11556 & n11561;
  assign n11563 = ~n11551 & ~n11562;
  assign n11564 = pi232 & ~n11563;
  assign n11565 = pi299 & ~n11543;
  assign n11566 = ~pi299 & ~n11554;
  assign n11567 = ~pi232 & ~n11565;
  assign n11568 = ~n11566 & n11567;
  assign n11569 = ~n11564 & ~n11568;
  assign n11570 = n7720 & ~n11569;
  assign n11571 = n7513 & ~n11486;
  assign n11572 = ~n11487 & ~n11495;
  assign n11573 = ~n11571 & n11572;
  assign n11574 = n8038 & ~n11573;
  assign n11575 = ~n11502 & ~n11574;
  assign n11576 = n2734 & ~n11575;
  assign n11577 = ~n2734 & n11518;
  assign n11578 = ~pi1093 & ~n11501;
  assign n11579 = ~n11577 & ~n11578;
  assign n11580 = ~n11576 & n11579;
  assign n11581 = ~po1057 & n11580;
  assign n11582 = po1057 & n11497;
  assign n11583 = ~n10082 & n11582;
  assign n11584 = ~n11581 & ~n11583;
  assign n11585 = pi210 & ~n11584;
  assign n11586 = pi137 & n11578;
  assign n11587 = ~pi137 & ~n11573;
  assign n11588 = ~pi1093 & n11587;
  assign n11589 = ~n11518 & ~n11586;
  assign n11590 = ~n11588 & n11589;
  assign n11591 = ~po1057 & n11590;
  assign n11592 = ~n11582 & ~n11591;
  assign n11593 = n8890 & n11535;
  assign n11594 = ~n2734 & ~n11593;
  assign n11595 = ~n11592 & n11594;
  assign n11596 = pi137 & ~n11575;
  assign n11597 = ~n11586 & ~n11587;
  assign n11598 = ~n11596 & n11597;
  assign n11599 = ~po1057 & ~n11598;
  assign n11600 = pi137 & ~n8038;
  assign n11601 = n7513 & ~n11600;
  assign n11602 = n11497 & ~n11601;
  assign n11603 = po1057 & ~n11602;
  assign n11604 = n2734 & ~n11603;
  assign n11605 = ~n11599 & n11604;
  assign n11606 = ~n11595 & ~n11605;
  assign n11607 = ~pi210 & ~n11606;
  assign n11608 = ~n11585 & ~n11607;
  assign n11609 = ~n11544 & ~n11608;
  assign n11610 = ~n2734 & n11590;
  assign n11611 = n2734 & n11598;
  assign n11612 = ~n11610 & ~n11611;
  assign n11613 = ~pi210 & n11612;
  assign n11614 = pi210 & ~n11580;
  assign n11615 = n11544 & ~n11614;
  assign n11616 = ~n11613 & n11615;
  assign n11617 = pi299 & ~n11616;
  assign n11618 = ~n11609 & n11617;
  assign n11619 = pi198 & ~n11584;
  assign n11620 = ~pi198 & ~n11606;
  assign n11621 = ~n11619 & ~n11620;
  assign n11622 = ~n11555 & ~n11621;
  assign n11623 = ~pi198 & ~n11612;
  assign n11624 = pi198 & n11580;
  assign n11625 = ~n11623 & ~n11624;
  assign n11626 = n11555 & ~n11625;
  assign n11627 = ~pi299 & ~n11626;
  assign n11628 = ~n11622 & n11627;
  assign n11629 = ~n11618 & ~n11628;
  assign n11630 = pi232 & ~n11629;
  assign n11631 = ~pi299 & ~n11621;
  assign n11632 = pi299 & ~n11608;
  assign n11633 = ~pi232 & ~n11631;
  assign n11634 = ~n11632 & n11633;
  assign n11635 = ~n7720 & ~n11634;
  assign n11636 = ~n11630 & n11635;
  assign n11637 = ~n11570 & ~n11636;
  assign po234 = n10146 & ~n11637;
  assign n11639 = n2578 & n2593;
  assign n11640 = ~pi86 & ~n11639;
  assign n11641 = n6342 & ~n11640;
  assign n11642 = n2491 & n11641;
  assign n11643 = ~pi314 & ~n11642;
  assign n11644 = pi86 & n8885;
  assign n11645 = n2587 & n11644;
  assign n11646 = pi314 & ~n11645;
  assign n11647 = n10147 & ~n11646;
  assign po235 = ~n11643 & n11647;
  assign n11649 = pi119 & pi232;
  assign po236 = ~pi468 & n11649;
  assign n11651 = pi163 & ~n9685;
  assign n11652 = ~pi163 & ~n9681;
  assign n11653 = ~n9683 & n11652;
  assign n11654 = ~n11651 & ~n11653;
  assign n11655 = pi232 & n11654;
  assign n11656 = pi75 & ~n11655;
  assign n11657 = pi100 & ~n11655;
  assign n11658 = ~n11656 & ~n11657;
  assign n11659 = pi147 & n7484;
  assign n11660 = n8975 & n11659;
  assign n11661 = n11658 & ~n11660;
  assign n11662 = ~n8975 & n11655;
  assign n11663 = pi74 & ~n11662;
  assign n11664 = ~n3432 & ~n11663;
  assign n11665 = n11661 & n11664;
  assign n11666 = pi299 & ~n11654;
  assign n11667 = ~n9711 & n9713;
  assign n11668 = ~pi184 & n11667;
  assign n11669 = pi184 & n6170;
  assign n11670 = ~n11667 & n11669;
  assign n11671 = ~pi299 & ~n11668;
  assign n11672 = ~n11670 & n11671;
  assign n11673 = pi232 & ~n11672;
  assign n11674 = ~n11666 & n11673;
  assign n11675 = ~n8975 & n11674;
  assign n11676 = pi74 & ~n11675;
  assign n11677 = ~pi55 & ~n11676;
  assign n11678 = ~pi187 & ~pi299;
  assign n11679 = ~pi147 & pi299;
  assign n11680 = ~n11678 & ~n11679;
  assign n11681 = n7484 & n11680;
  assign n11682 = n8975 & ~n11681;
  assign n11683 = pi54 & ~n11682;
  assign n11684 = ~n11675 & n11683;
  assign n11685 = ~pi187 & ~n9011;
  assign n11686 = pi187 & ~n9013;
  assign n11687 = pi147 & ~n11686;
  assign n11688 = ~n11685 & n11687;
  assign n11689 = ~pi147 & pi187;
  assign n11690 = n9018 & n11689;
  assign n11691 = ~n11688 & ~n11690;
  assign n11692 = pi38 & ~n11691;
  assign n11693 = ~pi40 & ~n9197;
  assign n11694 = ~pi95 & ~n11693;
  assign n11695 = ~pi40 & ~n9214;
  assign n11696 = pi166 & n11695;
  assign n11697 = n11694 & ~n11696;
  assign n11698 = n6170 & ~n9259;
  assign n11699 = ~n11697 & n11698;
  assign n11700 = ~pi153 & ~n11699;
  assign n11701 = ~pi40 & ~n9275;
  assign n11702 = ~pi95 & ~n11701;
  assign n11703 = pi166 & ~n11702;
  assign n11704 = n11698 & n11703;
  assign n11705 = n9239 & n10305;
  assign n11706 = pi153 & ~n11705;
  assign n11707 = ~n11704 & n11706;
  assign n11708 = pi160 & ~n11707;
  assign n11709 = ~n11700 & n11708;
  assign n11710 = ~pi153 & n11697;
  assign n11711 = ~n2449 & ~n9259;
  assign n11712 = n9099 & ~n9100;
  assign n11713 = ~n11711 & ~n11712;
  assign n11714 = ~n11455 & ~n11702;
  assign n11715 = pi153 & ~n11703;
  assign n11716 = ~n11714 & n11715;
  assign n11717 = ~pi160 & n6170;
  assign n11718 = ~n11716 & n11717;
  assign n11719 = ~n11713 & n11718;
  assign n11720 = ~n11710 & n11719;
  assign n11721 = pi163 & ~n11720;
  assign n11722 = ~n11709 & n11721;
  assign n11723 = ~pi40 & ~n9353;
  assign n11724 = ~pi95 & ~n11723;
  assign n11725 = ~n11713 & ~n11724;
  assign n11726 = pi166 & n11725;
  assign n11727 = ~pi40 & n9173;
  assign n11728 = ~pi32 & ~n11727;
  assign n11729 = ~n9240 & ~n11728;
  assign n11730 = ~pi95 & ~n11729;
  assign n11731 = ~n11713 & ~n11730;
  assign n11732 = pi210 & ~n11731;
  assign n11733 = ~n9261 & ~n11728;
  assign n11734 = ~pi95 & ~n11733;
  assign n11735 = ~n11713 & ~n11734;
  assign n11736 = ~pi210 & ~n11735;
  assign n11737 = n10305 & ~n11732;
  assign n11738 = ~n11736 & n11737;
  assign n11739 = ~pi153 & ~n11738;
  assign n11740 = ~n11726 & n11739;
  assign n11741 = ~pi95 & ~n9252;
  assign n11742 = ~n11713 & ~n11741;
  assign n11743 = pi210 & ~n11742;
  assign n11744 = ~n9263 & ~n11713;
  assign n11745 = ~pi210 & ~n11744;
  assign n11746 = pi166 & n6170;
  assign n11747 = ~n11743 & n11746;
  assign n11748 = ~n11745 & n11747;
  assign n11749 = ~n9329 & ~n11713;
  assign n11750 = ~pi210 & ~n11749;
  assign n11751 = ~n9325 & ~n11713;
  assign n11752 = pi210 & ~n11751;
  assign n11753 = n10305 & ~n11750;
  assign n11754 = ~n11752 & n11753;
  assign n11755 = pi153 & ~n11748;
  assign n11756 = ~n11754 & n11755;
  assign n11757 = ~pi160 & ~n11756;
  assign n11758 = ~n11740 & n11757;
  assign n11759 = n11723 & n11746;
  assign n11760 = ~n9259 & ~n11734;
  assign n11761 = ~pi210 & ~n11760;
  assign n11762 = ~n9259 & ~n11730;
  assign n11763 = pi210 & ~n11762;
  assign n11764 = n10305 & ~n11761;
  assign n11765 = ~n11763 & n11764;
  assign n11766 = ~pi153 & ~n11765;
  assign n11767 = ~n11759 & n11766;
  assign n11768 = pi210 & ~n9326;
  assign n11769 = ~pi210 & ~n9330;
  assign n11770 = n10305 & ~n11768;
  assign n11771 = ~n11769 & n11770;
  assign n11772 = ~pi210 & ~n9264;
  assign n11773 = ~n9259 & ~n11741;
  assign n11774 = pi210 & ~n11773;
  assign n11775 = n11746 & ~n11772;
  assign n11776 = ~n11774 & n11775;
  assign n11777 = pi153 & ~n11771;
  assign n11778 = ~n11776 & n11777;
  assign n11779 = pi160 & ~n11778;
  assign n11780 = ~n11767 & n11779;
  assign n11781 = ~pi163 & ~n11780;
  assign n11782 = ~n11758 & n11781;
  assign n11783 = ~n11722 & ~n11782;
  assign n11784 = ~n6170 & n11725;
  assign n11785 = pi299 & ~n11784;
  assign n11786 = ~n11783 & n11785;
  assign n11787 = ~pi40 & ~n9229;
  assign n11788 = ~pi95 & ~n11787;
  assign n11789 = ~n11713 & ~n11788;
  assign n11790 = ~n6170 & n11789;
  assign n11791 = ~pi175 & ~pi299;
  assign n11792 = pi189 & n11695;
  assign n11793 = n11694 & ~n11792;
  assign n11794 = ~pi182 & n11713;
  assign n11795 = pi182 & n9259;
  assign n11796 = n6170 & ~n11795;
  assign n11797 = ~n11794 & n11796;
  assign n11798 = ~n11793 & n11797;
  assign n11799 = pi184 & ~n11798;
  assign n11800 = pi189 & n6170;
  assign n11801 = n11787 & n11800;
  assign n11802 = ~pi198 & ~n11760;
  assign n11803 = pi198 & ~n11762;
  assign n11804 = n10301 & ~n11802;
  assign n11805 = ~n11803 & n11804;
  assign n11806 = pi182 & ~pi184;
  assign n11807 = ~n11805 & n11806;
  assign n11808 = ~n11801 & n11807;
  assign n11809 = ~n11799 & ~n11808;
  assign n11810 = n11791 & ~n11809;
  assign n11811 = n9332 & n10301;
  assign n11812 = ~pi198 & ~n9264;
  assign n11813 = pi198 & ~n11773;
  assign n11814 = n11800 & ~n11812;
  assign n11815 = ~n11813 & n11814;
  assign n11816 = pi182 & ~n11811;
  assign n11817 = ~n11815 & n11816;
  assign n11818 = ~pi198 & ~n11744;
  assign n11819 = pi198 & ~n11742;
  assign n11820 = n11800 & ~n11818;
  assign n11821 = ~n11819 & n11820;
  assign n11822 = ~pi182 & ~n11821;
  assign n11823 = ~n11817 & ~n11822;
  assign n11824 = pi95 & ~pi182;
  assign n11825 = ~n9332 & ~n11824;
  assign n11826 = n10301 & ~n11713;
  assign n11827 = ~n11825 & n11826;
  assign n11828 = ~n11823 & ~n11827;
  assign n11829 = ~pi184 & ~n11828;
  assign n11830 = pi175 & ~pi299;
  assign n11831 = ~pi95 & pi189;
  assign n11832 = n2476 & ~n11831;
  assign n11833 = n11701 & ~n11832;
  assign n11834 = ~n11824 & ~n11833;
  assign n11835 = n11669 & ~n11834;
  assign n11836 = ~n11794 & n11835;
  assign n11837 = n11830 & ~n11836;
  assign n11838 = ~n11829 & n11837;
  assign n11839 = ~n11810 & ~n11838;
  assign n11840 = ~n11790 & ~n11839;
  assign n11841 = ~n10301 & n11789;
  assign n11842 = pi198 & ~n11731;
  assign n11843 = ~pi198 & ~n11735;
  assign n11844 = n10301 & ~n11842;
  assign n11845 = ~n11843 & n11844;
  assign n11846 = ~pi182 & ~pi184;
  assign n11847 = n11791 & n11846;
  assign n11848 = ~n11845 & n11847;
  assign n11849 = ~n11841 & n11848;
  assign n11850 = ~n11840 & ~n11849;
  assign n11851 = ~n11786 & n11850;
  assign n11852 = pi232 & ~n11851;
  assign n11853 = ~pi299 & n11789;
  assign n11854 = pi299 & n11725;
  assign n11855 = ~pi232 & ~n11853;
  assign n11856 = ~n11854 & n11855;
  assign n11857 = ~pi39 & ~n11856;
  assign n11858 = ~n11852 & n11857;
  assign n11859 = ~n9044 & ~n9239;
  assign n11860 = ~pi40 & ~n9043;
  assign n11861 = ~pi189 & ~n11860;
  assign n11862 = n2476 & ~n9047;
  assign n11863 = n9227 & ~n11862;
  assign n11864 = n6200 & n9239;
  assign n11865 = n2476 & ~n9041;
  assign n11866 = ~pi40 & ~n11865;
  assign n11867 = n6206 & n11866;
  assign n11868 = ~n11864 & ~n11867;
  assign n11869 = ~n11863 & n11868;
  assign n11870 = pi189 & ~n6197;
  assign n11871 = n11869 & n11870;
  assign n11872 = ~n11861 & ~n11871;
  assign n11873 = pi179 & ~n11872;
  assign n11874 = n6197 & ~n11860;
  assign n11875 = n9062 & n9227;
  assign n11876 = ~n2476 & n9227;
  assign n11877 = ~n11875 & ~n11876;
  assign n11878 = n11868 & n11877;
  assign n11879 = ~pi189 & ~n11878;
  assign n11880 = ~n6200 & n11866;
  assign n11881 = ~n11864 & ~n11880;
  assign n11882 = pi189 & ~n11881;
  assign n11883 = ~pi179 & ~n6197;
  assign n11884 = ~n11882 & n11883;
  assign n11885 = ~n11879 & n11884;
  assign n11886 = ~n11874 & ~n11885;
  assign n11887 = ~n11873 & n11886;
  assign n11888 = n9044 & ~n11887;
  assign n11889 = ~n11859 & ~n11888;
  assign n11890 = ~pi299 & ~n11889;
  assign n11891 = ~n9055 & n9239;
  assign n11892 = pi299 & ~n11891;
  assign n11893 = n6223 & ~n11860;
  assign n11894 = ~n6223 & n11881;
  assign n11895 = ~n11893 & ~n11894;
  assign n11896 = ~pi166 & ~n6223;
  assign n11897 = ~n11895 & ~n11896;
  assign n11898 = n11878 & n11896;
  assign n11899 = n9055 & ~n11898;
  assign n11900 = ~n11897 & n11899;
  assign n11901 = n11892 & ~n11900;
  assign n11902 = ~n11890 & ~n11901;
  assign n11903 = ~pi156 & pi232;
  assign n11904 = ~n11902 & n11903;
  assign n11905 = pi166 & ~n6223;
  assign n11906 = n11869 & n11905;
  assign n11907 = ~n11860 & ~n11905;
  assign n11908 = n9055 & ~n11907;
  assign n11909 = ~n11906 & n11908;
  assign n11910 = n11892 & ~n11909;
  assign n11911 = ~n11890 & ~n11910;
  assign n11912 = pi156 & pi232;
  assign n11913 = ~n11911 & n11912;
  assign n11914 = ~n6197 & n11881;
  assign n11915 = ~n11874 & ~n11914;
  assign n11916 = n9044 & ~n11915;
  assign n11917 = ~pi299 & ~n11859;
  assign n11918 = ~n11916 & n11917;
  assign n11919 = n9057 & n11895;
  assign n11920 = ~pi232 & ~n11919;
  assign n11921 = ~n11918 & n11920;
  assign n11922 = pi39 & ~n11921;
  assign n11923 = ~n11904 & n11922;
  assign n11924 = ~n11913 & n11923;
  assign n11925 = ~pi38 & ~n11924;
  assign n11926 = ~n11858 & n11925;
  assign n11927 = ~n11692 & ~n11926;
  assign n11928 = n3241 & ~n11927;
  assign n11929 = pi100 & ~n11674;
  assign n11930 = pi38 & ~n11681;
  assign n11931 = ~pi100 & ~n11930;
  assign n11932 = ~pi38 & ~pi40;
  assign n11933 = pi87 & ~n2476;
  assign n11934 = n11932 & n11933;
  assign n11935 = n11931 & ~n11934;
  assign n11936 = pi87 & n11935;
  assign n11937 = ~n11929 & ~n11936;
  assign n11938 = ~n11928 & n11937;
  assign n11939 = n3238 & ~n11938;
  assign n11940 = pi75 & ~n11674;
  assign n11941 = pi39 & ~n9239;
  assign n11942 = n9638 & ~n11941;
  assign n11943 = n2476 & ~n9037;
  assign n11944 = ~pi40 & ~n11943;
  assign n11945 = ~pi179 & ~pi299;
  assign n11946 = ~pi156 & pi299;
  assign n11947 = ~n11945 & ~n11946;
  assign n11948 = n7484 & n11947;
  assign n11949 = n2476 & n11948;
  assign n11950 = n11944 & ~n11949;
  assign n11951 = ~pi39 & ~n11950;
  assign n11952 = n11942 & ~n11951;
  assign n11953 = n11935 & ~n11952;
  assign n11954 = ~n11929 & ~n11953;
  assign n11955 = n9450 & ~n11954;
  assign n11956 = ~n11940 & ~n11955;
  assign n11957 = ~n11939 & n11956;
  assign n11958 = ~pi54 & ~n11957;
  assign n11959 = ~n11684 & ~n11958;
  assign n11960 = ~pi74 & ~n11959;
  assign n11961 = n11677 & ~n11960;
  assign n11962 = pi55 & ~n11663;
  assign n11963 = pi54 & ~n11661;
  assign n11964 = pi163 & pi232;
  assign n11965 = ~n6170 & n9037;
  assign n11966 = n9024 & ~n11965;
  assign n11967 = n11964 & n11966;
  assign n11968 = n11944 & ~n11967;
  assign n11969 = ~pi39 & ~n11968;
  assign n11970 = n11942 & ~n11969;
  assign n11971 = pi38 & ~n11659;
  assign n11972 = ~pi100 & ~n11971;
  assign n11973 = ~n11934 & n11972;
  assign n11974 = ~n11970 & n11973;
  assign n11975 = ~n11657 & ~n11974;
  assign n11976 = n3238 & ~n11975;
  assign n11977 = ~n11932 & n11972;
  assign n11978 = ~n11657 & ~n11977;
  assign n11979 = ~n9445 & n11978;
  assign n11980 = n9450 & ~n11979;
  assign n11981 = ~n11656 & ~n11980;
  assign n11982 = ~n11976 & n11981;
  assign n11983 = ~pi54 & ~n11982;
  assign n11984 = ~n11963 & ~n11983;
  assign n11985 = ~pi74 & ~n11984;
  assign n11986 = n11962 & ~n11985;
  assign n11987 = n3294 & ~n11986;
  assign n11988 = ~n11961 & n11987;
  assign n11989 = ~pi75 & ~n11978;
  assign n11990 = ~n11656 & ~n11989;
  assign n11991 = ~pi54 & ~n11990;
  assign n11992 = ~n11963 & ~n11991;
  assign n11993 = ~pi74 & ~n11992;
  assign n11994 = ~n11663 & ~n11993;
  assign n11995 = ~n3294 & ~n11994;
  assign n11996 = n3432 & ~n11995;
  assign n11997 = ~n9507 & n11996;
  assign n11998 = ~n11988 & n11997;
  assign n11999 = ~n11665 & ~n11998;
  assign n12000 = ~pi79 & n11999;
  assign n12001 = ~pi32 & pi95;
  assign n12002 = ~pi479 & n12001;
  assign n12003 = n2552 & n12002;
  assign n12004 = ~pi40 & ~n12003;
  assign n12005 = n9606 & n12004;
  assign n12006 = n10305 & ~n12005;
  assign n12007 = n9609 & n12004;
  assign n12008 = n11746 & ~n12007;
  assign n12009 = ~pi153 & ~n12008;
  assign n12010 = ~n12006 & n12009;
  assign n12011 = ~pi210 & ~n9555;
  assign n12012 = ~n9553 & n12004;
  assign n12013 = ~n12011 & n12012;
  assign n12014 = n10305 & ~n12013;
  assign n12015 = ~n9574 & n12007;
  assign n12016 = n11746 & ~n12015;
  assign n12017 = pi153 & ~n12016;
  assign n12018 = ~n12014 & n12017;
  assign n12019 = ~n12010 & ~n12018;
  assign n12020 = pi40 & ~n6170;
  assign n12021 = pi163 & ~n12020;
  assign n12022 = ~n12019 & n12021;
  assign n12023 = pi160 & ~n12022;
  assign n12024 = pi153 & n9553;
  assign n12025 = n9606 & ~n12024;
  assign n12026 = n10305 & ~n12025;
  assign n12027 = pi153 & n9574;
  assign n12028 = n9609 & ~n12027;
  assign n12029 = n11746 & ~n12028;
  assign n12030 = ~pi40 & pi163;
  assign n12031 = ~n12029 & n12030;
  assign n12032 = ~n12026 & n12031;
  assign n12033 = pi153 & n9565;
  assign n12034 = n9578 & n12033;
  assign n12035 = n9593 & n10305;
  assign n12036 = ~pi40 & ~pi163;
  assign n12037 = ~n12035 & n12036;
  assign n12038 = ~n12034 & n12037;
  assign n12039 = ~pi160 & ~n12038;
  assign n12040 = ~n12032 & n12039;
  assign n12041 = ~n12023 & ~n12040;
  assign n12042 = n6170 & n12003;
  assign n12043 = n12038 & ~n12042;
  assign n12044 = pi299 & ~n12043;
  assign n12045 = ~n12041 & n12044;
  assign n12046 = pi184 & n9585;
  assign n12047 = ~pi184 & ~n9593;
  assign n12048 = ~pi189 & ~n12047;
  assign n12049 = ~n12046 & n12048;
  assign n12050 = pi182 & n12003;
  assign n12051 = pi184 & pi189;
  assign n12052 = ~n9588 & n12051;
  assign n12053 = ~n12050 & ~n12052;
  assign n12054 = ~n12049 & n12053;
  assign n12055 = n6170 & ~n12054;
  assign n12056 = ~pi40 & ~n12055;
  assign n12057 = n11791 & ~n12056;
  assign n12058 = pi189 & ~n9578;
  assign n12059 = ~pi189 & ~n9564;
  assign n12060 = n3093 & ~n12058;
  assign n12061 = ~n12059 & n12060;
  assign n12062 = ~n12050 & ~n12061;
  assign n12063 = n6170 & ~n12062;
  assign n12064 = ~pi184 & ~n12063;
  assign n12065 = ~n9557 & n10301;
  assign n12066 = pi189 & n9576;
  assign n12067 = ~pi182 & pi184;
  assign n12068 = ~n12066 & n12067;
  assign n12069 = ~n12065 & n12068;
  assign n12070 = ~n12064 & ~n12069;
  assign n12071 = ~pi40 & ~n12070;
  assign n12072 = ~n9556 & n12012;
  assign n12073 = n10301 & ~n12072;
  assign n12074 = n9575 & n12004;
  assign n12075 = n11800 & ~n12074;
  assign n12076 = pi182 & pi184;
  assign n12077 = ~n12020 & n12076;
  assign n12078 = ~n12075 & n12077;
  assign n12079 = ~n12073 & n12078;
  assign n12080 = n11830 & ~n12079;
  assign n12081 = ~n12071 & n12080;
  assign n12082 = ~n12057 & ~n12081;
  assign n12083 = ~n12045 & n12082;
  assign n12084 = ~pi39 & ~n12083;
  assign n12085 = n2552 & n9565;
  assign n12086 = ~n6223 & n9055;
  assign n12087 = pi156 & n6209;
  assign n12088 = ~pi166 & n9039;
  assign n12089 = ~n12087 & ~n12088;
  assign n12090 = n12086 & ~n12089;
  assign n12091 = n12085 & n12090;
  assign n12092 = ~pi40 & pi299;
  assign n12093 = ~n12091 & n12092;
  assign n12094 = ~pi189 & n9039;
  assign n12095 = pi179 & n6209;
  assign n12096 = ~n12094 & ~n12095;
  assign n12097 = ~n6197 & n9044;
  assign n12098 = ~n12096 & n12097;
  assign n12099 = n12085 & n12098;
  assign n12100 = ~pi40 & ~pi299;
  assign n12101 = ~n12099 & n12100;
  assign n12102 = pi39 & ~n12093;
  assign n12103 = ~n12101 & n12102;
  assign n12104 = pi232 & ~n12103;
  assign n12105 = ~n12084 & n12104;
  assign n12106 = ~pi40 & ~pi232;
  assign n12107 = ~pi38 & ~n12106;
  assign n12108 = ~n12105 & n12107;
  assign n12109 = ~n11692 & ~n12108;
  assign n12110 = n3241 & ~n12109;
  assign n12111 = pi87 & ~n11932;
  assign n12112 = n11931 & n12111;
  assign n12113 = ~n11929 & ~n12112;
  assign n12114 = ~n12110 & n12113;
  assign n12115 = n3238 & ~n12114;
  assign n12116 = n3093 & n3222;
  assign n12117 = n11948 & n12116;
  assign n12118 = n2552 & n12117;
  assign n12119 = n11932 & ~n12118;
  assign n12120 = n11931 & ~n12119;
  assign n12121 = ~n11929 & ~n12120;
  assign n12122 = n9450 & ~n12121;
  assign n12123 = ~n11940 & ~n12122;
  assign n12124 = ~n12115 & n12123;
  assign n12125 = ~pi54 & ~n12124;
  assign n12126 = ~n11684 & ~n12125;
  assign n12127 = ~pi74 & ~n12126;
  assign n12128 = n11677 & ~n12127;
  assign n12129 = ~pi92 & n3222;
  assign n12130 = n11964 & n12129;
  assign n12131 = n12085 & n12130;
  assign n12132 = n11932 & ~n12131;
  assign n12133 = ~pi75 & n11972;
  assign n12134 = ~n12132 & n12133;
  assign n12135 = n11658 & ~n12134;
  assign n12136 = ~pi54 & ~n12135;
  assign n12137 = ~n11963 & ~n12136;
  assign n12138 = ~pi74 & ~n12137;
  assign n12139 = n11962 & ~n12138;
  assign n12140 = n3294 & ~n12139;
  assign n12141 = ~n12128 & n12140;
  assign n12142 = n11996 & ~n12141;
  assign n12143 = ~n11665 & ~n12142;
  assign n12144 = pi79 & n12143;
  assign n12145 = ~pi34 & n10043;
  assign n12146 = ~n12144 & ~n12145;
  assign n12147 = ~n12000 & n12146;
  assign n12148 = ~pi79 & ~n8963;
  assign n12149 = n11999 & ~n12148;
  assign n12150 = n12143 & n12148;
  assign n12151 = n12145 & ~n12150;
  assign n12152 = ~n12149 & n12151;
  assign po237 = n12147 | n12152;
  assign n12154 = pi98 & pi1092;
  assign n12155 = pi1093 & n12154;
  assign n12156 = ~pi567 & n2755;
  assign n12157 = ~n12155 & ~n12156;
  assign n12158 = ~n8585 & n12157;
  assign n12159 = pi588 & ~n12158;
  assign n12160 = pi592 & ~n12157;
  assign n12161 = ~n7444 & n12157;
  assign n12162 = n7444 & ~n12156;
  assign n12163 = pi75 & n12155;
  assign n12164 = pi1091 & n12155;
  assign n12165 = ~pi110 & n2490;
  assign n12166 = ~pi88 & n2482;
  assign n12167 = n10375 & n12166;
  assign n12168 = n12165 & n12167;
  assign n12169 = n7453 & n12168;
  assign n12170 = n7460 & n12169;
  assign n12171 = pi51 & n12170;
  assign n12172 = pi90 & pi93;
  assign n12173 = ~pi841 & ~n2493;
  assign n12174 = ~n12172 & n12173;
  assign n12175 = n2536 & n12174;
  assign n12176 = n12169 & n12175;
  assign n12177 = ~n12171 & ~n12176;
  assign n12178 = pi824 & pi950;
  assign n12179 = n7464 & n12178;
  assign n12180 = ~n12177 & n12179;
  assign n12181 = ~pi98 & ~n12180;
  assign n12182 = pi1092 & ~n12181;
  assign n12183 = ~n12164 & ~n12182;
  assign n12184 = ~n7558 & ~n12164;
  assign n12185 = n3223 & ~n12184;
  assign n12186 = ~n12183 & n12185;
  assign n12187 = n3095 & n12178;
  assign n12188 = n12170 & n12187;
  assign n12189 = ~pi98 & ~n12188;
  assign n12190 = pi1092 & ~n12189;
  assign n12191 = ~n12164 & ~n12190;
  assign n12192 = n7600 & ~n12184;
  assign n12193 = ~n12191 & n12192;
  assign n12194 = ~n3208 & n12155;
  assign n12195 = ~n12193 & ~n12194;
  assign n12196 = ~n12186 & n12195;
  assign n12197 = ~pi75 & ~n12196;
  assign n12198 = ~n12163 & ~n12197;
  assign n12199 = pi567 & ~n12198;
  assign n12200 = n12162 & ~n12199;
  assign n12201 = ~n12161 & ~n12200;
  assign n12202 = ~pi592 & n12201;
  assign n12203 = ~n12160 & ~n12202;
  assign n12204 = ~n8507 & n12203;
  assign n12205 = ~pi1196 & ~n12157;
  assign n12206 = n8507 & ~n12205;
  assign n12207 = ~pi443 & ~n12157;
  assign n12208 = pi443 & ~n12203;
  assign n12209 = ~n12207 & ~n12208;
  assign n12210 = n8595 & n12209;
  assign n12211 = pi443 & ~n12157;
  assign n12212 = ~pi443 & ~n12203;
  assign n12213 = ~n12211 & ~n12212;
  assign n12214 = ~n8595 & n12213;
  assign n12215 = ~n12210 & ~n12214;
  assign n12216 = pi435 & ~n12215;
  assign n12217 = ~pi444 & n12213;
  assign n12218 = pi444 & n12209;
  assign n12219 = ~pi436 & ~n12217;
  assign n12220 = ~n12218 & n12219;
  assign n12221 = ~pi444 & n12209;
  assign n12222 = pi444 & n12213;
  assign n12223 = pi436 & ~n12221;
  assign n12224 = ~n12222 & n12223;
  assign n12225 = ~n12220 & ~n12224;
  assign n12226 = ~pi435 & n12225;
  assign n12227 = ~n12216 & ~n12226;
  assign n12228 = ~pi429 & n12227;
  assign n12229 = ~pi435 & ~n12215;
  assign n12230 = pi435 & n12225;
  assign n12231 = ~n12229 & ~n12230;
  assign n12232 = pi429 & n12231;
  assign n12233 = n8532 & ~n12228;
  assign n12234 = ~n12232 & n12233;
  assign n12235 = ~pi429 & n12231;
  assign n12236 = pi429 & n12227;
  assign n12237 = ~n8532 & ~n12235;
  assign n12238 = ~n12236 & n12237;
  assign n12239 = pi1196 & ~n12234;
  assign n12240 = ~n12238 & n12239;
  assign n12241 = n12206 & ~n12240;
  assign n12242 = ~n12204 & ~n12241;
  assign n12243 = ~pi428 & ~n12242;
  assign n12244 = pi428 & n12203;
  assign n12245 = ~n12243 & ~n12244;
  assign n12246 = ~pi427 & ~n12245;
  assign n12247 = pi428 & ~n12242;
  assign n12248 = ~pi428 & n12203;
  assign n12249 = ~n12247 & ~n12248;
  assign n12250 = pi427 & ~n12249;
  assign n12251 = ~n12246 & ~n12250;
  assign n12252 = pi430 & ~n12251;
  assign n12253 = ~pi427 & ~n12249;
  assign n12254 = pi427 & ~n12245;
  assign n12255 = ~n12253 & ~n12254;
  assign n12256 = ~pi430 & ~n12255;
  assign n12257 = ~n12252 & ~n12256;
  assign n12258 = pi426 & ~n12257;
  assign n12259 = pi430 & ~n12255;
  assign n12260 = ~pi430 & ~n12251;
  assign n12261 = ~n12259 & ~n12260;
  assign n12262 = ~pi426 & ~n12261;
  assign n12263 = ~n12258 & ~n12262;
  assign n12264 = pi445 & ~n12263;
  assign n12265 = pi426 & ~n12261;
  assign n12266 = ~pi426 & ~n12257;
  assign n12267 = ~n12265 & ~n12266;
  assign n12268 = ~pi445 & ~n12267;
  assign n12269 = ~n12264 & ~n12268;
  assign n12270 = pi448 & n12269;
  assign n12271 = pi445 & ~n12267;
  assign n12272 = ~pi445 & ~n12263;
  assign n12273 = ~n12271 & ~n12272;
  assign n12274 = ~pi448 & n12273;
  assign n12275 = n8453 & ~n12270;
  assign n12276 = ~n12274 & n12275;
  assign n12277 = pi448 & n12273;
  assign n12278 = ~pi448 & n12269;
  assign n12279 = ~n8453 & ~n12277;
  assign n12280 = ~n12278 & n12279;
  assign n12281 = pi1199 & ~n12276;
  assign n12282 = ~n12280 & n12281;
  assign n12283 = ~pi1199 & n12242;
  assign n12284 = n8585 & ~n12283;
  assign n12285 = ~n12282 & n12284;
  assign n12286 = n12159 & ~n12285;
  assign n12287 = pi591 & ~n12157;
  assign n12288 = pi590 & ~n12287;
  assign n12289 = n8684 & n12157;
  assign n12290 = ~n8684 & n12203;
  assign n12291 = ~n12289 & ~n12290;
  assign n12292 = pi1198 & ~n12291;
  assign n12293 = ~pi1198 & ~n12205;
  assign n12294 = n7618 & n12157;
  assign n12295 = ~n7618 & n12203;
  assign n12296 = ~n12294 & ~n12295;
  assign n12297 = pi355 & ~n12296;
  assign n12298 = pi455 & ~n12157;
  assign n12299 = ~pi455 & ~n12203;
  assign n12300 = ~n12298 & ~n12299;
  assign n12301 = ~pi452 & ~n12300;
  assign n12302 = ~pi455 & ~n12157;
  assign n12303 = pi455 & ~n12203;
  assign n12304 = ~n12302 & ~n12303;
  assign n12305 = pi452 & ~n12304;
  assign n12306 = ~n12301 & ~n12305;
  assign n12307 = ~pi355 & n12306;
  assign n12308 = ~n12297 & ~n12307;
  assign n12309 = ~pi458 & n12308;
  assign n12310 = ~pi355 & ~n12296;
  assign n12311 = pi355 & n12306;
  assign n12312 = ~n12310 & ~n12311;
  assign n12313 = pi458 & n12312;
  assign n12314 = ~n7633 & ~n12309;
  assign n12315 = ~n12313 & n12314;
  assign n12316 = ~pi458 & n12312;
  assign n12317 = pi458 & n12308;
  assign n12318 = n7633 & ~n12316;
  assign n12319 = ~n12317 & n12318;
  assign n12320 = pi1196 & ~n12315;
  assign n12321 = ~n12319 & n12320;
  assign n12322 = n12293 & ~n12321;
  assign n12323 = ~n12292 & ~n12322;
  assign n12324 = ~n7443 & ~n12323;
  assign n12325 = n7443 & n12203;
  assign n12326 = ~n12324 & ~n12325;
  assign n12327 = ~n7690 & n12326;
  assign n12328 = pi1199 & ~n12203;
  assign n12329 = pi351 & n12328;
  assign n12330 = ~n12327 & ~n12329;
  assign n12331 = ~pi461 & ~n12330;
  assign n12332 = ~n7684 & n12326;
  assign n12333 = ~pi351 & n12328;
  assign n12334 = ~n12332 & ~n12333;
  assign n12335 = pi461 & ~n12334;
  assign n12336 = ~n12331 & ~n12335;
  assign n12337 = ~pi357 & ~n12336;
  assign n12338 = ~pi461 & ~n12334;
  assign n12339 = pi461 & ~n12330;
  assign n12340 = ~n12338 & ~n12339;
  assign n12341 = pi357 & ~n12340;
  assign n12342 = ~n12337 & ~n12341;
  assign n12343 = ~pi356 & ~n12342;
  assign n12344 = ~pi357 & ~n12340;
  assign n12345 = pi357 & ~n12336;
  assign n12346 = ~n12344 & ~n12345;
  assign n12347 = pi356 & ~n12346;
  assign n12348 = ~n12343 & ~n12347;
  assign n12349 = ~pi354 & ~n12348;
  assign n12350 = ~pi356 & ~n12346;
  assign n12351 = pi356 & ~n12342;
  assign n12352 = ~n12350 & ~n12351;
  assign n12353 = pi354 & ~n12352;
  assign n12354 = ~n7415 & ~n12349;
  assign n12355 = ~n12353 & n12354;
  assign n12356 = ~pi354 & ~n12352;
  assign n12357 = pi354 & ~n12348;
  assign n12358 = n7415 & ~n12356;
  assign n12359 = ~n12357 & n12358;
  assign n12360 = ~pi591 & ~n12355;
  assign n12361 = ~n12359 & n12360;
  assign n12362 = n12288 & ~n12361;
  assign n12363 = ~pi1197 & ~n7900;
  assign n12364 = ~n12203 & ~n12363;
  assign n12365 = n8242 & ~n12161;
  assign n12366 = ~pi411 & n12154;
  assign n12367 = n7922 & ~n12366;
  assign n12368 = pi411 & n12182;
  assign n12369 = n12367 & ~n12368;
  assign n12370 = ~n7922 & ~n12154;
  assign n12371 = ~n7924 & ~n12370;
  assign n12372 = ~pi411 & n12182;
  assign n12373 = ~n12371 & ~n12372;
  assign n12374 = ~n12369 & ~n12373;
  assign n12375 = ~n12164 & ~n12374;
  assign n12376 = n12185 & ~n12375;
  assign n12377 = pi411 & n12190;
  assign n12378 = n12367 & ~n12377;
  assign n12379 = ~pi411 & n12190;
  assign n12380 = ~n12371 & ~n12379;
  assign n12381 = ~n12378 & ~n12380;
  assign n12382 = ~n12164 & ~n12381;
  assign n12383 = n12192 & ~n12382;
  assign n12384 = ~n12194 & ~n12383;
  assign n12385 = ~n12376 & n12384;
  assign n12386 = ~pi75 & ~n12385;
  assign n12387 = ~n12163 & ~n12386;
  assign n12388 = pi567 & ~n12387;
  assign n12389 = n12162 & ~n12388;
  assign n12390 = n12365 & ~n12389;
  assign n12391 = ~n12160 & ~n12205;
  assign n12392 = ~pi1199 & n12391;
  assign n12393 = ~n12390 & n12392;
  assign n12394 = n7963 & n12193;
  assign n12395 = n7963 & n12182;
  assign n12396 = ~n7963 & n12154;
  assign n12397 = ~n12395 & ~n12396;
  assign n12398 = n12186 & ~n12397;
  assign n12399 = ~n12394 & ~n12398;
  assign n12400 = n12385 & n12399;
  assign n12401 = n12365 & ~n12400;
  assign n12402 = n7963 & n12190;
  assign n12403 = ~n12396 & ~n12402;
  assign n12404 = n12193 & ~n12403;
  assign n12405 = ~n12194 & ~n12404;
  assign n12406 = ~n12398 & n12405;
  assign n12407 = n8340 & ~n12161;
  assign n12408 = ~n12406 & n12407;
  assign n12409 = ~n12401 & ~n12408;
  assign n12410 = ~pi75 & pi567;
  assign n12411 = ~n12409 & n12410;
  assign n12412 = n7933 & n12162;
  assign n12413 = ~n12157 & ~n12412;
  assign n12414 = pi1199 & ~n12413;
  assign n12415 = ~n12411 & n12414;
  assign n12416 = ~n7900 & ~n12415;
  assign n12417 = ~n12393 & n12416;
  assign n12418 = ~pi1197 & n12417;
  assign n12419 = ~n12364 & ~n12418;
  assign n12420 = ~pi333 & ~n12419;
  assign n12421 = n7900 & ~n12203;
  assign n12422 = ~n12417 & ~n12421;
  assign n12423 = pi333 & ~n12422;
  assign n12424 = ~n12420 & ~n12423;
  assign n12425 = ~pi391 & ~n12424;
  assign n12426 = pi333 & ~n12419;
  assign n12427 = ~pi333 & ~n12422;
  assign n12428 = ~n12426 & ~n12427;
  assign n12429 = pi391 & ~n12428;
  assign n12430 = ~n12425 & ~n12429;
  assign n12431 = ~pi392 & ~n12430;
  assign n12432 = ~pi391 & ~n12428;
  assign n12433 = pi391 & ~n12424;
  assign n12434 = ~n12432 & ~n12433;
  assign n12435 = pi392 & ~n12434;
  assign n12436 = ~n12431 & ~n12435;
  assign n12437 = ~pi393 & ~n12436;
  assign n12438 = ~pi392 & ~n12434;
  assign n12439 = pi392 & ~n12430;
  assign n12440 = ~n12438 & ~n12439;
  assign n12441 = pi393 & ~n12440;
  assign n12442 = ~n8238 & ~n12437;
  assign n12443 = ~n12441 & n12442;
  assign n12444 = ~pi393 & ~n12440;
  assign n12445 = pi393 & ~n12436;
  assign n12446 = n8238 & ~n12444;
  assign n12447 = ~n12445 & n12446;
  assign n12448 = pi591 & ~n12443;
  assign n12449 = ~n12447 & n12448;
  assign n12450 = ~pi592 & ~n12157;
  assign n12451 = pi592 & n12201;
  assign n12452 = ~n12450 & ~n12451;
  assign n12453 = ~n8725 & n12452;
  assign n12454 = n8725 & n12157;
  assign n12455 = pi1199 & ~n12454;
  assign n12456 = ~n12453 & n12455;
  assign n12457 = ~pi1197 & ~n12157;
  assign n12458 = ~n7745 & ~n12457;
  assign n12459 = n7769 & n12452;
  assign n12460 = ~n7769 & n12157;
  assign n12461 = pi1197 & ~n12460;
  assign n12462 = ~n12459 & n12461;
  assign n12463 = n12458 & ~n12462;
  assign n12464 = n7745 & n12452;
  assign n12465 = ~pi1199 & ~n12464;
  assign n12466 = ~n12463 & n12465;
  assign n12467 = ~n12456 & ~n12466;
  assign n12468 = ~pi374 & ~n12467;
  assign n12469 = ~pi1198 & ~n12467;
  assign n12470 = pi1198 & ~n12452;
  assign n12471 = ~n12469 & ~n12470;
  assign n12472 = pi374 & ~n12471;
  assign n12473 = ~n12468 & ~n12472;
  assign n12474 = ~pi369 & ~n12473;
  assign n12475 = pi371 & n8189;
  assign n12476 = ~pi371 & ~n8189;
  assign n12477 = ~n12475 & ~n12476;
  assign n12478 = pi370 & ~n12477;
  assign n12479 = ~pi370 & n12477;
  assign n12480 = ~n12478 & ~n12479;
  assign n12481 = ~pi374 & ~n12471;
  assign n12482 = pi374 & ~n12467;
  assign n12483 = ~n12481 & ~n12482;
  assign n12484 = pi369 & ~n12483;
  assign n12485 = ~n12474 & ~n12480;
  assign n12486 = ~n12484 & n12485;
  assign n12487 = pi369 & ~n12473;
  assign n12488 = ~pi369 & ~n12483;
  assign n12489 = n12480 & ~n12487;
  assign n12490 = ~n12488 & n12489;
  assign n12491 = ~pi591 & ~n12486;
  assign n12492 = ~n12490 & n12491;
  assign n12493 = ~pi590 & ~n12492;
  assign n12494 = ~n12449 & n12493;
  assign n12495 = ~pi588 & ~n12494;
  assign n12496 = ~n12362 & n12495;
  assign n12497 = n7720 & ~n12496;
  assign n12498 = ~n12286 & n12497;
  assign n12499 = ~n8044 & ~n12155;
  assign n12500 = ~pi122 & n12499;
  assign n12501 = n7558 & ~n12500;
  assign n12502 = n3208 & ~n12164;
  assign n12503 = ~n12501 & n12502;
  assign n12504 = ~pi87 & n12502;
  assign n12505 = ~n12182 & n12504;
  assign n12506 = pi87 & n12502;
  assign n12507 = ~n12190 & n12506;
  assign n12508 = ~n12505 & ~n12507;
  assign n12509 = pi122 & ~n12508;
  assign n12510 = ~n12503 & ~n12509;
  assign n12511 = ~pi75 & ~n12510;
  assign n12512 = pi567 & n7444;
  assign n12513 = ~n7479 & n12499;
  assign n12514 = n12512 & ~n12513;
  assign n12515 = ~n12511 & n12514;
  assign n12516 = ~n7444 & ~n12499;
  assign n12517 = ~n12156 & ~n12516;
  assign n12518 = ~n12515 & n12517;
  assign n12519 = ~pi592 & ~n12518;
  assign n12520 = ~n12160 & ~n12519;
  assign n12521 = ~n8507 & n12520;
  assign n12522 = pi443 & ~n12520;
  assign n12523 = ~n12207 & ~n12522;
  assign n12524 = n8595 & n12523;
  assign n12525 = ~pi443 & ~n12520;
  assign n12526 = ~n12211 & ~n12525;
  assign n12527 = ~n8595 & n12526;
  assign n12528 = ~n12524 & ~n12527;
  assign n12529 = pi435 & ~n12528;
  assign n12530 = ~pi444 & n12526;
  assign n12531 = pi444 & n12523;
  assign n12532 = ~pi436 & ~n12530;
  assign n12533 = ~n12531 & n12532;
  assign n12534 = ~pi444 & n12523;
  assign n12535 = pi444 & n12526;
  assign n12536 = pi436 & ~n12534;
  assign n12537 = ~n12535 & n12536;
  assign n12538 = ~n12533 & ~n12537;
  assign n12539 = ~pi435 & n12538;
  assign n12540 = ~n12529 & ~n12539;
  assign n12541 = ~pi429 & n12540;
  assign n12542 = ~pi435 & ~n12528;
  assign n12543 = pi435 & n12538;
  assign n12544 = ~n12542 & ~n12543;
  assign n12545 = pi429 & n12544;
  assign n12546 = n8532 & ~n12541;
  assign n12547 = ~n12545 & n12546;
  assign n12548 = ~pi429 & n12544;
  assign n12549 = pi429 & n12540;
  assign n12550 = ~n8532 & ~n12548;
  assign n12551 = ~n12549 & n12550;
  assign n12552 = pi1196 & ~n12547;
  assign n12553 = ~n12551 & n12552;
  assign n12554 = n12206 & ~n12553;
  assign n12555 = ~n12521 & ~n12554;
  assign n12556 = pi428 & ~n12555;
  assign n12557 = ~pi428 & n12520;
  assign n12558 = ~n12556 & ~n12557;
  assign n12559 = ~pi427 & ~n12558;
  assign n12560 = ~pi428 & ~n12555;
  assign n12561 = pi428 & n12520;
  assign n12562 = ~n12560 & ~n12561;
  assign n12563 = pi427 & ~n12562;
  assign n12564 = ~n12559 & ~n12563;
  assign n12565 = pi430 & ~n12564;
  assign n12566 = ~pi427 & ~n12562;
  assign n12567 = pi427 & ~n12558;
  assign n12568 = ~n12566 & ~n12567;
  assign n12569 = ~pi430 & ~n12568;
  assign n12570 = ~n12565 & ~n12569;
  assign n12571 = pi426 & ~n12570;
  assign n12572 = pi430 & ~n12568;
  assign n12573 = ~pi430 & ~n12564;
  assign n12574 = ~n12572 & ~n12573;
  assign n12575 = ~pi426 & ~n12574;
  assign n12576 = ~n12571 & ~n12575;
  assign n12577 = pi445 & ~n12576;
  assign n12578 = pi426 & ~n12574;
  assign n12579 = ~pi426 & ~n12570;
  assign n12580 = ~n12578 & ~n12579;
  assign n12581 = ~pi445 & ~n12580;
  assign n12582 = ~n12577 & ~n12581;
  assign n12583 = pi448 & n12582;
  assign n12584 = pi445 & ~n12580;
  assign n12585 = ~pi445 & ~n12576;
  assign n12586 = ~n12584 & ~n12585;
  assign n12587 = ~pi448 & n12586;
  assign n12588 = ~n8453 & ~n12583;
  assign n12589 = ~n12587 & n12588;
  assign n12590 = ~pi448 & n12582;
  assign n12591 = pi448 & n12586;
  assign n12592 = n8453 & ~n12590;
  assign n12593 = ~n12591 & n12592;
  assign n12594 = pi1199 & ~n12589;
  assign n12595 = ~n12593 & n12594;
  assign n12596 = ~pi1199 & n12555;
  assign n12597 = n8585 & ~n12596;
  assign n12598 = ~n12595 & n12597;
  assign n12599 = n12159 & ~n12598;
  assign n12600 = ~n8684 & n12520;
  assign n12601 = ~n12289 & ~n12600;
  assign n12602 = pi1198 & ~n12601;
  assign n12603 = ~n7618 & n12520;
  assign n12604 = ~n12294 & ~n12603;
  assign n12605 = ~pi355 & ~n12604;
  assign n12606 = ~pi455 & ~n12520;
  assign n12607 = ~n12298 & ~n12606;
  assign n12608 = ~pi452 & ~n12607;
  assign n12609 = pi455 & ~n12520;
  assign n12610 = ~n12302 & ~n12609;
  assign n12611 = pi452 & ~n12610;
  assign n12612 = ~n12608 & ~n12611;
  assign n12613 = pi355 & n12612;
  assign n12614 = ~n12605 & ~n12613;
  assign n12615 = ~pi458 & n12614;
  assign n12616 = pi355 & ~n12604;
  assign n12617 = ~pi355 & n12612;
  assign n12618 = ~n12616 & ~n12617;
  assign n12619 = pi458 & n12618;
  assign n12620 = n7633 & ~n12615;
  assign n12621 = ~n12619 & n12620;
  assign n12622 = ~pi458 & n12618;
  assign n12623 = pi458 & n12614;
  assign n12624 = ~n7633 & ~n12622;
  assign n12625 = ~n12623 & n12624;
  assign n12626 = pi1196 & ~n12621;
  assign n12627 = ~n12625 & n12626;
  assign n12628 = n12293 & ~n12627;
  assign n12629 = ~n12602 & ~n12628;
  assign n12630 = ~n7443 & ~n12629;
  assign n12631 = n7443 & n12520;
  assign n12632 = ~n12630 & ~n12631;
  assign n12633 = ~n7690 & n12632;
  assign n12634 = pi1199 & ~n12520;
  assign n12635 = pi351 & n12634;
  assign n12636 = ~n12633 & ~n12635;
  assign n12637 = ~pi461 & ~n12636;
  assign n12638 = ~n7684 & n12632;
  assign n12639 = ~pi351 & n12634;
  assign n12640 = ~n12638 & ~n12639;
  assign n12641 = pi461 & ~n12640;
  assign n12642 = ~n12637 & ~n12641;
  assign n12643 = ~pi357 & ~n12642;
  assign n12644 = ~pi461 & ~n12640;
  assign n12645 = pi461 & ~n12636;
  assign n12646 = ~n12644 & ~n12645;
  assign n12647 = pi357 & ~n12646;
  assign n12648 = ~n12643 & ~n12647;
  assign n12649 = ~pi356 & ~n12648;
  assign n12650 = ~pi357 & ~n12646;
  assign n12651 = pi357 & ~n12642;
  assign n12652 = ~n12650 & ~n12651;
  assign n12653 = pi356 & ~n12652;
  assign n12654 = ~n12649 & ~n12653;
  assign n12655 = ~pi354 & ~n12654;
  assign n12656 = ~pi356 & ~n12652;
  assign n12657 = pi356 & ~n12648;
  assign n12658 = ~n12656 & ~n12657;
  assign n12659 = pi354 & ~n12658;
  assign n12660 = ~n7415 & ~n12655;
  assign n12661 = ~n12659 & n12660;
  assign n12662 = ~pi354 & ~n12658;
  assign n12663 = pi354 & ~n12654;
  assign n12664 = n7415 & ~n12662;
  assign n12665 = ~n12663 & n12664;
  assign n12666 = ~pi591 & ~n12661;
  assign n12667 = ~n12665 & n12666;
  assign n12668 = n12288 & ~n12667;
  assign n12669 = pi367 & ~n12157;
  assign n12670 = pi592 & ~n12518;
  assign n12671 = ~n12450 & ~n12670;
  assign n12672 = ~pi367 & ~n12671;
  assign n12673 = ~n12669 & ~n12672;
  assign n12674 = n7748 & ~n12673;
  assign n12675 = ~pi367 & ~n12157;
  assign n12676 = pi367 & ~n12671;
  assign n12677 = ~n12675 & ~n12676;
  assign n12678 = ~n7748 & ~n12677;
  assign n12679 = ~n12674 & ~n12678;
  assign n12680 = n7751 & ~n12679;
  assign n12681 = ~n7748 & n12673;
  assign n12682 = n7748 & n12677;
  assign n12683 = ~n12681 & ~n12682;
  assign n12684 = ~n7751 & n12683;
  assign n12685 = ~n7760 & ~n12680;
  assign n12686 = ~n12684 & n12685;
  assign n12687 = ~n7751 & ~n12679;
  assign n12688 = n7751 & n12683;
  assign n12689 = n7760 & ~n12687;
  assign n12690 = ~n12688 & n12689;
  assign n12691 = pi1197 & ~n12686;
  assign n12692 = ~n12690 & n12691;
  assign n12693 = n12458 & ~n12692;
  assign n12694 = n7745 & n12671;
  assign n12695 = ~pi1199 & ~n12694;
  assign n12696 = ~n12693 & n12695;
  assign n12697 = ~n8725 & n12671;
  assign n12698 = ~n12454 & ~n12697;
  assign n12699 = pi1199 & n12698;
  assign n12700 = ~n12696 & ~n12699;
  assign n12701 = ~pi374 & ~n12700;
  assign n12702 = ~pi1198 & n12696;
  assign n12703 = n7825 & n12698;
  assign n12704 = pi1198 & ~n12671;
  assign n12705 = ~n12703 & ~n12704;
  assign n12706 = ~n12702 & n12705;
  assign n12707 = pi374 & ~n12706;
  assign n12708 = ~n12701 & ~n12707;
  assign n12709 = pi369 & ~n12708;
  assign n12710 = ~pi374 & ~n12706;
  assign n12711 = pi374 & ~n12700;
  assign n12712 = ~n12710 & ~n12711;
  assign n12713 = ~pi369 & ~n12712;
  assign n12714 = n12480 & ~n12709;
  assign n12715 = ~n12713 & n12714;
  assign n12716 = ~pi369 & ~n12708;
  assign n12717 = pi369 & ~n12712;
  assign n12718 = ~n12480 & ~n12716;
  assign n12719 = ~n12717 & n12718;
  assign n12720 = ~pi591 & ~n12715;
  assign n12721 = ~n12719 & n12720;
  assign n12722 = ~n12363 & n12520;
  assign n12723 = pi397 & ~pi404;
  assign n12724 = ~pi397 & pi404;
  assign n12725 = ~n12723 & ~n12724;
  assign n12726 = pi411 & ~n12725;
  assign n12727 = ~pi411 & n12725;
  assign n12728 = ~n12726 & ~n12727;
  assign n12729 = ~n7904 & n12728;
  assign n12730 = n7904 & ~n12728;
  assign n12731 = ~n12729 & ~n12730;
  assign n12732 = n7496 & ~n12731;
  assign n12733 = ~n12154 & ~n12732;
  assign n12734 = ~pi412 & ~n12733;
  assign n12735 = n7496 & n12731;
  assign n12736 = ~n12154 & ~n12735;
  assign n12737 = pi412 & ~n12736;
  assign n12738 = n7916 & ~n12734;
  assign n12739 = ~n12737 & n12738;
  assign n12740 = pi412 & ~n12733;
  assign n12741 = ~pi412 & ~n12736;
  assign n12742 = ~n7916 & ~n12740;
  assign n12743 = ~n12741 & n12742;
  assign n12744 = ~pi122 & ~n12739;
  assign n12745 = ~n12743 & n12744;
  assign n12746 = ~n12154 & ~n12745;
  assign n12747 = n7558 & ~n12746;
  assign n12748 = ~n12164 & ~n12747;
  assign n12749 = pi567 & ~n12748;
  assign n12750 = ~n12156 & ~n12749;
  assign n12751 = ~n12162 & ~n12750;
  assign n12752 = pi122 & n12374;
  assign n12753 = ~n12745 & ~n12752;
  assign n12754 = n7558 & ~n12753;
  assign n12755 = n12504 & ~n12754;
  assign n12756 = pi122 & n12381;
  assign n12757 = ~n12745 & ~n12756;
  assign n12758 = n7558 & ~n12757;
  assign n12759 = n12506 & ~n12758;
  assign n12760 = ~n3208 & n12748;
  assign n12761 = ~n12759 & ~n12760;
  assign n12762 = ~n12755 & n12761;
  assign n12763 = ~pi75 & ~n12762;
  assign n12764 = pi75 & n12748;
  assign n12765 = n12512 & ~n12764;
  assign n12766 = ~n12763 & n12765;
  assign n12767 = ~n12751 & ~n12766;
  assign n12768 = n8242 & ~n12767;
  assign n12769 = ~n12205 & ~n12768;
  assign n12770 = ~pi1199 & ~n12769;
  assign n12771 = ~pi122 & n7496;
  assign n12772 = ~n12154 & ~n12771;
  assign n12773 = n7496 & n7963;
  assign n12774 = ~pi122 & ~n12154;
  assign n12775 = ~n12773 & n12774;
  assign n12776 = ~n12184 & ~n12775;
  assign n12777 = ~n12772 & n12776;
  assign n12778 = pi567 & n12777;
  assign n12779 = ~n12156 & ~n12778;
  assign n12780 = ~n12749 & n12779;
  assign n12781 = ~n12162 & ~n12780;
  assign n12782 = n3208 & ~n12776;
  assign n12783 = ~n12747 & n12782;
  assign n12784 = ~n12402 & n12506;
  assign n12785 = ~n12381 & n12784;
  assign n12786 = n12397 & n12504;
  assign n12787 = ~n12374 & n12786;
  assign n12788 = ~n12785 & ~n12787;
  assign n12789 = ~pi122 & n12773;
  assign n12790 = ~n12745 & ~n12789;
  assign n12791 = ~n12788 & n12790;
  assign n12792 = ~n12783 & ~n12791;
  assign n12793 = ~pi75 & ~n12792;
  assign n12794 = ~n7479 & ~n12777;
  assign n12795 = ~n12747 & n12794;
  assign n12796 = n12512 & ~n12795;
  assign n12797 = ~n12793 & n12796;
  assign n12798 = ~n12781 & ~n12797;
  assign n12799 = n8242 & ~n12798;
  assign n12800 = ~n12162 & ~n12779;
  assign n12801 = n12403 & n12506;
  assign n12802 = ~n12786 & ~n12801;
  assign n12803 = pi122 & ~n12802;
  assign n12804 = ~n12782 & ~n12803;
  assign n12805 = ~pi75 & ~n12804;
  assign n12806 = n12512 & ~n12794;
  assign n12807 = ~n12805 & n12806;
  assign n12808 = ~n12800 & ~n12807;
  assign n12809 = n8340 & ~n12808;
  assign n12810 = ~n12799 & ~n12809;
  assign n12811 = pi1199 & ~n12810;
  assign n12812 = ~n12160 & ~n12811;
  assign n12813 = ~n12770 & n12812;
  assign n12814 = n12363 & n12813;
  assign n12815 = ~n12722 & ~n12814;
  assign n12816 = pi333 & ~n12815;
  assign n12817 = n7900 & ~n12520;
  assign n12818 = ~n7900 & ~n12813;
  assign n12819 = ~n12817 & ~n12818;
  assign n12820 = ~pi333 & n12819;
  assign n12821 = ~n12816 & ~n12820;
  assign n12822 = pi391 & ~n12821;
  assign n12823 = pi333 & ~n12819;
  assign n12824 = ~pi333 & n12815;
  assign n12825 = ~n12823 & ~n12824;
  assign n12826 = ~pi391 & n12825;
  assign n12827 = ~n12822 & ~n12826;
  assign n12828 = pi392 & ~n12827;
  assign n12829 = ~pi391 & n12821;
  assign n12830 = pi391 & ~n12825;
  assign n12831 = ~n12829 & ~n12830;
  assign n12832 = ~pi392 & n12831;
  assign n12833 = ~n12828 & ~n12832;
  assign n12834 = pi393 & ~n12833;
  assign n12835 = ~pi392 & ~n12827;
  assign n12836 = pi392 & n12831;
  assign n12837 = ~n12835 & ~n12836;
  assign n12838 = ~pi393 & ~n12837;
  assign n12839 = ~n12834 & ~n12838;
  assign n12840 = ~n8238 & ~n12839;
  assign n12841 = pi393 & ~n12837;
  assign n12842 = ~pi393 & ~n12833;
  assign n12843 = ~n12841 & ~n12842;
  assign n12844 = n8238 & ~n12843;
  assign n12845 = pi591 & ~n12840;
  assign n12846 = ~n12844 & n12845;
  assign n12847 = ~pi590 & ~n12846;
  assign n12848 = ~n12721 & n12847;
  assign n12849 = ~pi588 & ~n12848;
  assign n12850 = ~n12668 & n12849;
  assign n12851 = ~n7720 & ~n12850;
  assign n12852 = ~n12599 & n12851;
  assign n12853 = ~pi80 & ~po1038;
  assign n12854 = ~n12852 & n12853;
  assign n12855 = ~n12498 & n12854;
  assign n12856 = ~n8685 & n12157;
  assign n12857 = ~n12363 & ~n12856;
  assign n12858 = n8242 & ~n12750;
  assign n12859 = n12391 & ~n12858;
  assign n12860 = ~pi1199 & ~n12859;
  assign n12861 = n8242 & ~n12780;
  assign n12862 = n8340 & ~n12779;
  assign n12863 = ~n12160 & ~n12862;
  assign n12864 = ~n12861 & n12863;
  assign n12865 = pi1199 & ~n12864;
  assign n12866 = ~n12860 & ~n12865;
  assign n12867 = n12363 & ~n12866;
  assign n12868 = ~n12857 & ~n12867;
  assign n12869 = pi333 & ~n12868;
  assign n12870 = n7900 & ~n12856;
  assign n12871 = ~n7900 & ~n12866;
  assign n12872 = ~n12870 & ~n12871;
  assign n12873 = ~pi333 & ~n12872;
  assign n12874 = ~n12869 & ~n12873;
  assign n12875 = pi391 & ~n12874;
  assign n12876 = pi392 & n8241;
  assign n12877 = ~pi392 & ~n8241;
  assign n12878 = ~n12876 & ~n12877;
  assign n12879 = ~pi333 & ~n12868;
  assign n12880 = pi333 & ~n12872;
  assign n12881 = ~n12879 & ~n12880;
  assign n12882 = ~pi391 & ~n12881;
  assign n12883 = ~n12875 & ~n12878;
  assign n12884 = ~n12882 & n12883;
  assign n12885 = pi391 & ~n12881;
  assign n12886 = ~pi391 & ~n12874;
  assign n12887 = n12878 & ~n12885;
  assign n12888 = ~n12886 & n12887;
  assign n12889 = pi591 & ~n12884;
  assign n12890 = ~n12888 & n12889;
  assign n12891 = n8112 & n8752;
  assign n12892 = n12157 & ~n12891;
  assign n12893 = ~pi591 & ~n12892;
  assign n12894 = ~pi590 & ~n12893;
  assign n12895 = ~n12890 & n12894;
  assign n12896 = ~n8693 & n12157;
  assign n12897 = n8689 & n12896;
  assign n12898 = ~n7690 & n12897;
  assign n12899 = ~n12856 & ~n12898;
  assign n12900 = pi461 & ~n12899;
  assign n12901 = ~n7684 & n12897;
  assign n12902 = ~n12856 & ~n12901;
  assign n12903 = ~pi461 & ~n12902;
  assign n12904 = ~n12900 & ~n12903;
  assign n12905 = pi357 & ~n12904;
  assign n12906 = pi461 & ~n12902;
  assign n12907 = ~pi461 & ~n12899;
  assign n12908 = ~n12906 & ~n12907;
  assign n12909 = ~pi357 & ~n12908;
  assign n12910 = ~n12905 & ~n12909;
  assign n12911 = pi356 & ~n12910;
  assign n12912 = pi357 & ~n12908;
  assign n12913 = ~pi357 & ~n12904;
  assign n12914 = ~n12912 & ~n12913;
  assign n12915 = ~pi356 & ~n12914;
  assign n12916 = ~n12911 & ~n12915;
  assign n12917 = pi354 & n12916;
  assign n12918 = pi356 & ~n12914;
  assign n12919 = ~pi356 & ~n12910;
  assign n12920 = ~n12918 & ~n12919;
  assign n12921 = ~pi354 & n12920;
  assign n12922 = ~n7415 & ~n12917;
  assign n12923 = ~n12921 & n12922;
  assign n12924 = pi354 & n12920;
  assign n12925 = ~pi354 & n12916;
  assign n12926 = n7415 & ~n12924;
  assign n12927 = ~n12925 & n12926;
  assign n12928 = ~pi591 & ~n12923;
  assign n12929 = ~n12927 & n12928;
  assign n12930 = n12288 & ~n12929;
  assign n12931 = ~pi588 & ~n12930;
  assign n12932 = ~n12895 & n12931;
  assign n12933 = pi592 & ~n8507;
  assign n12934 = n8112 & ~n8815;
  assign n12935 = ~n12933 & n12934;
  assign n12936 = n12157 & ~n12935;
  assign n12937 = pi428 & ~n12936;
  assign n12938 = ~pi428 & ~n12856;
  assign n12939 = ~n12937 & ~n12938;
  assign n12940 = ~pi427 & ~n12939;
  assign n12941 = ~pi428 & ~n12936;
  assign n12942 = pi428 & ~n12856;
  assign n12943 = ~n12941 & ~n12942;
  assign n12944 = pi427 & ~n12943;
  assign n12945 = ~n12940 & ~n12944;
  assign n12946 = ~pi430 & ~n12945;
  assign n12947 = ~pi427 & ~n12943;
  assign n12948 = pi427 & ~n12939;
  assign n12949 = ~n12947 & ~n12948;
  assign n12950 = pi430 & ~n12949;
  assign n12951 = ~n12946 & ~n12950;
  assign n12952 = ~pi426 & ~n12951;
  assign n12953 = ~pi430 & ~n12949;
  assign n12954 = pi430 & ~n12945;
  assign n12955 = ~n12953 & ~n12954;
  assign n12956 = pi426 & ~n12955;
  assign n12957 = ~n12952 & ~n12956;
  assign n12958 = ~pi445 & ~n12957;
  assign n12959 = ~pi426 & ~n12955;
  assign n12960 = pi426 & ~n12951;
  assign n12961 = ~n12959 & ~n12960;
  assign n12962 = pi445 & ~n12961;
  assign n12963 = ~n12958 & ~n12962;
  assign n12964 = pi448 & ~n12963;
  assign n12965 = ~pi445 & ~n12961;
  assign n12966 = pi445 & ~n12957;
  assign n12967 = ~n12965 & ~n12966;
  assign n12968 = ~pi448 & ~n12967;
  assign n12969 = n8453 & ~n12964;
  assign n12970 = ~n12968 & n12969;
  assign n12971 = ~pi448 & ~n12963;
  assign n12972 = pi448 & ~n12967;
  assign n12973 = ~n8453 & ~n12971;
  assign n12974 = ~n12972 & n12973;
  assign n12975 = pi1199 & ~n12970;
  assign n12976 = ~n12974 & n12975;
  assign n12977 = ~pi1199 & ~n12936;
  assign n12978 = n8585 & ~n12977;
  assign n12979 = ~n12976 & n12978;
  assign n12980 = n12159 & ~n12979;
  assign n12981 = ~n7720 & ~n12980;
  assign n12982 = ~n12932 & n12981;
  assign n12983 = n7720 & n12157;
  assign n12984 = ~pi80 & po1038;
  assign n12985 = ~n12983 & n12984;
  assign n12986 = ~n12982 & n12985;
  assign n12987 = ~pi217 & ~n12986;
  assign n12988 = ~n12855 & n12987;
  assign n12989 = ~pi80 & ~n12157;
  assign n12990 = pi217 & ~n12989;
  assign n12991 = n8856 & ~n12990;
  assign po238 = ~n12988 & n12991;
  assign n12993 = ~po1038 & n11279;
  assign n12994 = pi81 & ~pi314;
  assign n12995 = n2478 & n12994;
  assign n12996 = pi68 & ~pi81;
  assign n12997 = n2469 & n12996;
  assign n12998 = n10992 & n12997;
  assign n12999 = n11416 & n12998;
  assign n13000 = n2634 & n12999;
  assign n13001 = ~n12995 & ~n13000;
  assign po239 = n12993 & ~n13001;
  assign n13003 = pi69 & pi314;
  assign n13004 = n2601 & n13003;
  assign n13005 = pi66 & ~pi73;
  assign n13006 = n2457 & n13005;
  assign n13007 = n2471 & n13006;
  assign n13008 = ~n13004 & ~n13007;
  assign n13009 = n11080 & n11082;
  assign po240 = ~n13008 & n13009;
  assign n13011 = n2486 & n11081;
  assign n13012 = n2491 & n13011;
  assign n13013 = n2469 & n2608;
  assign n13014 = pi84 & n9113;
  assign n13015 = n13013 & n13014;
  assign n13016 = ~pi83 & ~n13015;
  assign n13017 = n13012 & ~n13016;
  assign n13018 = n2604 & n13017;
  assign n13019 = ~pi314 & ~n13018;
  assign n13020 = n2456 & n13015;
  assign n13021 = n13012 & n13020;
  assign n13022 = pi314 & ~n13021;
  assign n13023 = n10147 & ~n13022;
  assign po241 = ~n13019 & n13023;
  assign n13025 = pi211 & pi299;
  assign n13026 = pi219 & pi299;
  assign n13027 = ~n13025 & ~n13026;
  assign n13028 = ~n10794 & n13027;
  assign n13029 = ~po1038 & n13028;
  assign po242 = n11354 & n13029;
  assign n13031 = n6322 & n11083;
  assign n13032 = ~pi314 & n11084;
  assign n13033 = n11414 & n13032;
  assign n13034 = ~n13031 & ~n13033;
  assign po243 = n11080 & ~n13034;
  assign n13036 = n7531 & n11371;
  assign n13037 = n7534 & n11374;
  assign n13038 = ~n13036 & ~n13037;
  assign po244 = n10960 & ~n13038;
  assign n13040 = n2654 & n13011;
  assign n13041 = pi314 & n10147;
  assign n13042 = n2491 & n13041;
  assign po245 = n13040 & n13042;
  assign n13044 = n7496 & n11008;
  assign n13045 = ~pi1093 & ~n13044;
  assign n13046 = n7452 & n12167;
  assign n13047 = n11005 & n13046;
  assign n13048 = n11020 & n12165;
  assign n13049 = n13047 & n13048;
  assign n13050 = pi1093 & ~n13049;
  assign n13051 = n3269 & ~n10054;
  assign n13052 = ~n13050 & n13051;
  assign n13053 = ~n13045 & n13052;
  assign n13054 = n7720 & ~n13053;
  assign n13055 = n2497 & n7496;
  assign n13056 = ~pi1093 & n3094;
  assign n13057 = n3269 & n13056;
  assign n13058 = n13055 & n13057;
  assign n13059 = n11435 & n13058;
  assign n13060 = n2679 & n13059;
  assign n13061 = ~n7720 & ~n13060;
  assign n13062 = ~po1038 & ~n13061;
  assign po246 = ~n13054 & n13062;
  assign n13064 = pi70 & ~n8945;
  assign n13065 = n2454 & n8899;
  assign n13066 = n8918 & n13065;
  assign n13067 = n10166 & n13066;
  assign n13068 = pi841 & n7459;
  assign n13069 = n13067 & n13068;
  assign n13070 = ~pi70 & ~n13069;
  assign n13071 = n3095 & n10146;
  assign n13072 = ~n13070 & n13071;
  assign po247 = ~n13064 & n13072;
  assign n13074 = ~pi1050 & n9562;
  assign n13075 = ~pi90 & ~n13074;
  assign n13076 = n11303 & ~n13075;
  assign n13077 = ~n2706 & n13076;
  assign po248 = ~n7447 & n13077;
  assign n13079 = ~pi58 & n2565;
  assign n13080 = ~n10139 & ~n13079;
  assign n13081 = n2796 & n10143;
  assign n13082 = ~n13080 & n13081;
  assign n13083 = pi24 & n2534;
  assign n13084 = ~n2796 & n13083;
  assign n13085 = n11063 & n13084;
  assign n13086 = n2565 & n13085;
  assign n13087 = ~pi39 & ~n13086;
  assign n13088 = ~n13082 & n13087;
  assign n13089 = n10178 & ~n13088;
  assign po249 = n7540 & n13089;
  assign n13091 = pi92 & n3096;
  assign n13092 = n3409 & n11454;
  assign n13093 = n13091 & n13092;
  assign n13094 = n5774 & n6230;
  assign n13095 = n7531 & n13094;
  assign n13096 = n3483 & n6210;
  assign n13097 = n7534 & n13096;
  assign n13098 = ~n13095 & ~n13097;
  assign n13099 = n3278 & n11103;
  assign n13100 = ~n13098 & n13099;
  assign n13101 = ~n13093 & ~n13100;
  assign po250 = n10144 & ~n13101;
  assign n13103 = ~pi1050 & n3096;
  assign n13104 = pi92 & ~n13103;
  assign n13105 = pi93 & n11063;
  assign n13106 = n2735 & n13105;
  assign n13107 = ~pi92 & ~n13106;
  assign n13108 = n10145 & ~n13107;
  assign po251 = ~n13104 & n13108;
  assign n13110 = n11046 & n11263;
  assign n13111 = n2734 & n13110;
  assign n13112 = pi1093 & ~n13111;
  assign n13113 = n7513 & ~n13112;
  assign n13114 = n10232 & n11044;
  assign n13115 = ~n2589 & ~n13114;
  assign n13116 = n2514 & n10143;
  assign n13117 = pi252 & n13116;
  assign n13118 = ~n13115 & n13117;
  assign n13119 = ~n13113 & ~n13118;
  assign n13120 = ~po840 & ~n13119;
  assign n13121 = ~n13110 & ~n13120;
  assign n13122 = pi252 & n13119;
  assign n13123 = ~n13121 & ~n13122;
  assign n13124 = n8874 & ~n13123;
  assign n13125 = ~n8874 & ~n13110;
  assign n13126 = n10146 & ~n13125;
  assign po252 = ~n13124 & n13126;
  assign n13128 = ~n6208 & ~n6455;
  assign n13129 = n3484 & ~n11394;
  assign n13130 = n13128 & n13129;
  assign n13131 = ~n11397 & n11400;
  assign n13132 = ~n6455 & n13131;
  assign n13133 = pi39 & ~n13132;
  assign n13134 = ~n13130 & n13133;
  assign n13135 = n2450 & n12001;
  assign n13136 = n11433 & n13135;
  assign n13137 = ~pi332 & n10143;
  assign n13138 = n11262 & n13137;
  assign n13139 = n13067 & n13138;
  assign n13140 = ~pi39 & ~n13139;
  assign n13141 = ~n13136 & n13140;
  assign n13142 = n10181 & ~n13141;
  assign po253 = ~n13134 & n13142;
  assign n13144 = n10289 & n13135;
  assign n13145 = pi479 & ~po840;
  assign n13146 = n2957 & n13145;
  assign n13147 = pi96 & n2535;
  assign n13148 = n2725 & n13147;
  assign n13149 = ~n13145 & n13148;
  assign n13150 = n2737 & n13149;
  assign n13151 = ~n13146 & ~n13150;
  assign n13152 = ~pi95 & ~n13151;
  assign n13153 = ~n13144 & ~n13152;
  assign po254 = n10146 & ~n13153;
  assign n13155 = pi39 & pi593;
  assign n13156 = ~n11402 & n13155;
  assign n13157 = ~n6455 & n13156;
  assign n13158 = n6151 & n13145;
  assign n13159 = ~po740 & ~n13158;
  assign n13160 = ~pi96 & n10150;
  assign n13161 = ~n13159 & n13160;
  assign n13162 = n11461 & n13161;
  assign n13163 = ~n13157 & ~n13162;
  assign po255 = n10181 & ~n13163;
  assign n13165 = ~pi92 & n11455;
  assign n13166 = ~n13091 & ~n13165;
  assign n13167 = pi314 & pi1050;
  assign n13168 = n10145 & n13167;
  assign po256 = ~n13166 & n13168;
  assign n13170 = ~pi72 & pi99;
  assign n13171 = ~n8087 & ~n13170;
  assign n13172 = ~n2734 & n13170;
  assign n13173 = n8087 & ~n13172;
  assign n13174 = ~n10294 & n13170;
  assign n13175 = n6254 & n10892;
  assign n13176 = ~n13174 & ~n13175;
  assign n13177 = n10427 & ~n13176;
  assign n13178 = n13173 & ~n13177;
  assign n13179 = ~n13171 & ~n13178;
  assign n13180 = ~pi39 & ~n13179;
  assign n13181 = ~pi72 & pi152;
  assign n13182 = n10306 & n13181;
  assign n13183 = pi299 & n13182;
  assign n13184 = ~pi72 & pi174;
  assign n13185 = ~pi299 & n13184;
  assign n13186 = n10302 & n13185;
  assign n13187 = ~n13183 & ~n13186;
  assign n13188 = pi232 & ~n13187;
  assign n13189 = pi39 & ~n13188;
  assign n13190 = n3242 & ~n13189;
  assign n13191 = ~n13180 & n13190;
  assign n13192 = ~pi39 & ~n13170;
  assign n13193 = ~n13189 & ~n13192;
  assign n13194 = ~n3242 & n13193;
  assign n13195 = pi75 & ~n13194;
  assign n13196 = ~n13191 & n13195;
  assign n13197 = pi41 & pi72;
  assign n13198 = pi99 & ~n13197;
  assign n13199 = ~n10355 & n13198;
  assign n13200 = n10724 & ~n13199;
  assign n13201 = ~n10366 & n13198;
  assign n13202 = n10723 & ~n13201;
  assign n13203 = ~n13200 & ~n13202;
  assign n13204 = pi228 & ~n13203;
  assign n13205 = ~n10408 & n13198;
  assign n13206 = ~pi228 & ~n10510;
  assign n13207 = ~n13205 & n13206;
  assign n13208 = ~pi39 & ~n13207;
  assign n13209 = ~n13204 & n13208;
  assign n13210 = n10457 & ~n13187;
  assign n13211 = ~n10921 & n13210;
  assign n13212 = n3207 & ~n13211;
  assign n13213 = ~n13209 & n13212;
  assign n13214 = ~n10425 & n13170;
  assign n13215 = n6253 & n10281;
  assign n13216 = ~n13214 & ~n13215;
  assign n13217 = n10427 & ~n13216;
  assign n13218 = n13173 & ~n13217;
  assign n13219 = ~n13171 & ~n13218;
  assign n13220 = ~pi39 & ~n13219;
  assign n13221 = ~n13189 & ~n13220;
  assign n13222 = n6251 & ~n13221;
  assign n13223 = pi38 & ~n13193;
  assign n13224 = ~pi87 & ~n13223;
  assign n13225 = ~n13222 & n13224;
  assign n13226 = ~n13213 & n13225;
  assign n13227 = pi228 & n10548;
  assign n13228 = pi228 & n10422;
  assign n13229 = n13170 & ~n13228;
  assign n13230 = n3277 & ~n13229;
  assign n13231 = ~n13227 & n13230;
  assign n13232 = ~n3277 & ~n13193;
  assign n13233 = pi87 & ~n13232;
  assign n13234 = ~n13231 & n13233;
  assign n13235 = ~pi75 & ~n13234;
  assign n13236 = ~n13226 & n13235;
  assign n13237 = ~n13196 & ~n13236;
  assign n13238 = n7444 & ~n13237;
  assign n13239 = ~n7444 & ~n13193;
  assign n13240 = ~po1038 & ~n13239;
  assign n13241 = ~n13238 & n13240;
  assign n13242 = pi232 & n13182;
  assign n13243 = pi39 & ~n13242;
  assign n13244 = po1038 & ~n13192;
  assign n13245 = ~n13243 & n13244;
  assign po257 = n13241 | n13245;
  assign n13247 = ~n7484 & n10058;
  assign n13248 = pi129 & ~n13247;
  assign n13249 = n6244 & ~n13248;
  assign n13250 = n6248 & ~n6270;
  assign n13251 = pi129 & ~n10058;
  assign n13252 = ~n6247 & ~n13251;
  assign n13253 = ~n13250 & ~n13252;
  assign n13254 = ~n13249 & n13253;
  assign n13255 = ~pi75 & n3222;
  assign n13256 = n6251 & n13255;
  assign n13257 = ~n13254 & n13256;
  assign n13258 = ~pi24 & n8953;
  assign n13259 = po840 & n13258;
  assign n13260 = ~n8950 & n13259;
  assign n13261 = ~n13257 & ~n13260;
  assign n13262 = n8867 & ~n13261;
  assign po258 = n3096 & n13262;
  assign n13264 = ~n8087 & ~n10287;
  assign n13265 = ~n2734 & n10287;
  assign n13266 = n8087 & ~n13265;
  assign n13267 = n2734 & ~n6261;
  assign n13268 = n10287 & ~n10293;
  assign n13269 = ~n10282 & ~n13268;
  assign n13270 = n13267 & ~n13269;
  assign n13271 = n13266 & ~n13270;
  assign n13272 = ~n13264 & ~n13271;
  assign n13273 = ~pi39 & ~n13272;
  assign n13274 = pi152 & n3386;
  assign n13275 = n6170 & n13274;
  assign n13276 = ~pi72 & n13275;
  assign n13277 = pi299 & ~n13276;
  assign n13278 = ~pi144 & pi174;
  assign n13279 = n10301 & n13278;
  assign n13280 = ~pi72 & n13279;
  assign n13281 = ~pi299 & ~n13280;
  assign n13282 = pi232 & ~n13277;
  assign n13283 = ~n13281 & n13282;
  assign n13284 = pi39 & ~n13283;
  assign n13285 = n3242 & ~n13284;
  assign n13286 = ~n13273 & n13285;
  assign n13287 = ~pi39 & ~n10287;
  assign n13288 = ~n13284 & ~n13287;
  assign n13289 = ~n3242 & n13288;
  assign n13290 = pi75 & ~n13289;
  assign n13291 = ~n13286 & n13290;
  assign n13292 = pi101 & n10353;
  assign n13293 = n2734 & ~n10340;
  assign n13294 = ~n13292 & n13293;
  assign n13295 = pi101 & ~n10364;
  assign n13296 = ~n2734 & ~n10360;
  assign n13297 = ~n13295 & n13296;
  assign n13298 = ~n13294 & ~n13297;
  assign n13299 = pi228 & ~n13298;
  assign n13300 = pi101 & ~n10406;
  assign n13301 = ~pi228 & ~n13300;
  assign n13302 = ~n10400 & n13301;
  assign n13303 = ~pi39 & ~n13302;
  assign n13304 = ~n13299 & n13303;
  assign n13305 = n10922 & n13275;
  assign n13306 = pi299 & ~n13305;
  assign n13307 = n10922 & n13279;
  assign n13308 = ~pi299 & ~n13307;
  assign n13309 = n10457 & ~n13306;
  assign n13310 = ~n13308 & n13309;
  assign n13311 = n3207 & ~n13310;
  assign n13312 = ~n13304 & n13311;
  assign n13313 = ~pi44 & n10926;
  assign n13314 = n10287 & ~n13313;
  assign n13315 = ~n10281 & ~n13314;
  assign n13316 = n13267 & ~n13315;
  assign n13317 = n13266 & ~n13316;
  assign n13318 = ~n13264 & ~n13317;
  assign n13319 = ~pi39 & ~n13318;
  assign n13320 = ~n13284 & ~n13319;
  assign n13321 = n6251 & ~n13320;
  assign n13322 = pi38 & ~n13288;
  assign n13323 = ~pi87 & ~n13322;
  assign n13324 = ~n13321 & n13323;
  assign n13325 = ~n13312 & n13324;
  assign n13326 = ~pi101 & n10939;
  assign n13327 = n10421 & n10938;
  assign n13328 = n10287 & ~n13327;
  assign n13329 = ~pi39 & ~n13328;
  assign n13330 = ~n13326 & n13329;
  assign n13331 = pi87 & ~n13284;
  assign n13332 = ~n13330 & n13331;
  assign n13333 = ~pi75 & ~n13332;
  assign n13334 = ~n13325 & n13333;
  assign n13335 = ~n13291 & ~n13334;
  assign n13336 = n7444 & ~n13335;
  assign n13337 = ~n7444 & ~n13288;
  assign n13338 = ~po1038 & ~n13337;
  assign n13339 = ~n13336 & n13338;
  assign n13340 = pi232 & n13276;
  assign n13341 = pi39 & ~n13340;
  assign n13342 = po1038 & ~n13287;
  assign n13343 = ~n13341 & n13342;
  assign po259 = n13339 | n13343;
  assign n13345 = n2660 & n8900;
  assign po260 = n12993 & n13345;
  assign n13347 = ~pi109 & ~n13040;
  assign n13348 = n6312 & ~n13347;
  assign n13349 = ~pi314 & ~n13348;
  assign n13350 = pi109 & n2574;
  assign n13351 = n2487 & n13350;
  assign n13352 = pi314 & ~n13351;
  assign n13353 = n11079 & ~n13352;
  assign po261 = ~n13349 & n13353;
  assign n13355 = n7720 & ~n8874;
  assign n13356 = n10055 & ~n13355;
  assign n13357 = n10395 & ~n13356;
  assign n13358 = ~pi110 & ~n13047;
  assign n13359 = ~pi47 & n11020;
  assign n13360 = ~n13358 & n13359;
  assign n13361 = n10378 & n13360;
  assign n13362 = ~po1057 & ~n13361;
  assign n13363 = po1057 & ~n13049;
  assign n13364 = ~n7485 & ~n10054;
  assign n13365 = ~n13363 & n13364;
  assign n13366 = ~n13362 & n13365;
  assign n13367 = n7485 & ~n10054;
  assign n13368 = n13361 & n13367;
  assign n13369 = ~n13366 & ~n13368;
  assign n13370 = ~n7720 & ~n13369;
  assign n13371 = ~n13357 & ~n13370;
  assign po262 = n10146 & ~n13371;
  assign n13373 = pi24 & n11261;
  assign n13374 = ~pi53 & ~n11260;
  assign n13375 = n2508 & ~n13374;
  assign n13376 = ~pi24 & n2514;
  assign n13377 = n13375 & n13376;
  assign n13378 = ~n13373 & ~n13377;
  assign n13379 = pi841 & ~n13378;
  assign n13380 = n8932 & n11241;
  assign n13381 = ~n13379 & ~n13380;
  assign po264 = n10147 & ~n13381;
  assign n13383 = ~pi999 & n10147;
  assign po265 = n11331 & n13383;
  assign n13385 = ~pi97 & n7456;
  assign n13386 = ~pi108 & ~n13385;
  assign n13387 = n2490 & ~n13386;
  assign n13388 = n10218 & n13387;
  assign n13389 = ~pi314 & ~n13388;
  assign n13390 = pi314 & ~n7458;
  assign n13391 = n7460 & ~n10241;
  assign n13392 = ~n13390 & n13391;
  assign n13393 = ~n13389 & n13392;
  assign n13394 = n7460 & n10241;
  assign n13395 = n13388 & n13394;
  assign n13396 = ~pi51 & ~n13395;
  assign n13397 = ~n13393 & n13396;
  assign n13398 = n3208 & n7497;
  assign n13399 = ~n13397 & n13398;
  assign n13400 = ~pi87 & ~n13399;
  assign n13401 = n6278 & n8867;
  assign po266 = ~n13400 & n13401;
  assign n13403 = n2593 & n11411;
  assign po267 = n13041 & n13403;
  assign n13405 = ~pi82 & ~pi109;
  assign n13406 = pi111 & n13405;
  assign n13407 = n12165 & n13406;
  assign n13408 = n2486 & n13407;
  assign n13409 = n11084 & n13408;
  assign n13410 = n2635 & n13409;
  assign n13411 = pi314 & n13410;
  assign n13412 = n8874 & n10055;
  assign n13413 = n10387 & n13412;
  assign n13414 = ~n13411 & ~n13413;
  assign po268 = n10147 & ~n13414;
  assign n13416 = pi72 & n10289;
  assign n13417 = ~pi314 & n13410;
  assign n13418 = n9154 & n13417;
  assign n13419 = ~n13416 & ~n13418;
  assign n13420 = n6371 & n10146;
  assign po269 = ~n13419 & n13420;
  assign po270 = ~pi124 | pi468;
  assign n13423 = ~pi99 & ~n10367;
  assign n13424 = ~n10356 & n13423;
  assign n13425 = pi113 & ~n10468;
  assign n13426 = ~n13424 & n13425;
  assign n13427 = ~pi113 & n10725;
  assign n13428 = pi228 & ~n13427;
  assign n13429 = ~n13426 & n13428;
  assign n13430 = pi113 & n10504;
  assign n13431 = ~pi228 & ~n10511;
  assign n13432 = ~n13430 & n13431;
  assign n13433 = ~pi39 & ~n13432;
  assign n13434 = ~n13429 & n13433;
  assign n13435 = n3207 & ~n13434;
  assign n13436 = ~pi39 & n10505;
  assign n13437 = pi38 & ~n13436;
  assign n13438 = n2734 & n8087;
  assign n13439 = n7547 & n10554;
  assign n13440 = ~n6260 & ~n13439;
  assign n13441 = n13438 & ~n13440;
  assign n13442 = n10505 & ~n13441;
  assign n13443 = ~n6260 & n13438;
  assign n13444 = ~pi113 & n13443;
  assign n13445 = n13215 & n13444;
  assign n13446 = ~n13442 & ~n13445;
  assign n13447 = ~pi39 & ~n13446;
  assign n13448 = n6251 & ~n13447;
  assign n13449 = ~n13437 & ~n13448;
  assign n13450 = ~n13435 & n13449;
  assign n13451 = ~pi87 & ~n13450;
  assign n13452 = n10505 & ~n10584;
  assign n13453 = ~pi113 & n13227;
  assign n13454 = ~n13452 & ~n13453;
  assign n13455 = n3277 & ~n13454;
  assign n13456 = ~n3207 & n13436;
  assign n13457 = pi87 & ~n13456;
  assign n13458 = ~n13455 & n13457;
  assign n13459 = ~n13451 & ~n13458;
  assign n13460 = ~pi75 & ~n13459;
  assign n13461 = n7487 & n13445;
  assign n13462 = ~n6260 & ~n10597;
  assign n13463 = n13438 & ~n13462;
  assign n13464 = n10505 & ~n13463;
  assign n13465 = ~n13461 & ~n13464;
  assign n13466 = n3223 & ~n13465;
  assign n13467 = ~n3242 & n13436;
  assign n13468 = pi75 & ~n13467;
  assign n13469 = ~n13466 & n13468;
  assign n13470 = ~n13460 & ~n13469;
  assign n13471 = n8867 & ~n13470;
  assign n13472 = ~n8867 & ~n13436;
  assign po271 = ~n13471 & ~n13472;
  assign n13474 = pi114 & n10774;
  assign n13475 = n11130 & ~n13474;
  assign n13476 = ~n10595 & n13475;
  assign n13477 = ~pi72 & pi114;
  assign n13478 = ~n11130 & ~n13477;
  assign n13479 = n3223 & ~n13478;
  assign n13480 = ~n13476 & n13479;
  assign n13481 = ~pi39 & n13477;
  assign n13482 = ~n3242 & n13481;
  assign n13483 = pi75 & ~n13482;
  assign n13484 = ~n13480 & n13483;
  assign n13485 = ~pi114 & ~n10728;
  assign n13486 = pi114 & ~n10718;
  assign n13487 = ~n13485 & ~n13486;
  assign n13488 = ~pi115 & ~n13487;
  assign n13489 = pi115 & ~n13477;
  assign n13490 = ~pi39 & ~n13489;
  assign n13491 = ~n13488 & n13490;
  assign n13492 = n3207 & ~n13491;
  assign n13493 = pi114 & ~n10557;
  assign n13494 = n11130 & ~n13493;
  assign n13495 = ~n10552 & n13494;
  assign n13496 = ~pi39 & ~n13478;
  assign n13497 = ~n13495 & n13496;
  assign n13498 = n6251 & ~n13497;
  assign n13499 = pi38 & ~n13481;
  assign n13500 = ~pi87 & ~n13499;
  assign n13501 = ~n13498 & n13500;
  assign n13502 = ~n13492 & n13501;
  assign n13503 = pi228 & n10555;
  assign n13504 = ~pi115 & n13503;
  assign n13505 = n13477 & ~n13504;
  assign n13506 = n3207 & ~n13505;
  assign n13507 = ~n10582 & n13506;
  assign n13508 = ~n3207 & ~n13481;
  assign n13509 = n11104 & ~n13508;
  assign n13510 = ~n13507 & n13509;
  assign n13511 = ~pi75 & ~n13510;
  assign n13512 = ~n13502 & n13511;
  assign n13513 = ~n13484 & ~n13512;
  assign n13514 = n8867 & ~n13513;
  assign n13515 = ~n8867 & ~n13481;
  assign po272 = ~n13514 & ~n13515;
  assign n13517 = ~pi52 & n11107;
  assign n13518 = ~pi115 & ~n13517;
  assign n13519 = n10550 & n13518;
  assign n13520 = n7487 & n13519;
  assign n13521 = pi115 & n10774;
  assign n13522 = n13438 & ~n13521;
  assign n13523 = ~n13520 & n13522;
  assign n13524 = ~pi72 & pi115;
  assign n13525 = ~n13438 & ~n13524;
  assign n13526 = n3223 & ~n13525;
  assign n13527 = ~n13523 & n13526;
  assign n13528 = ~pi39 & n13524;
  assign n13529 = ~n3242 & n13528;
  assign n13530 = pi75 & ~n13529;
  assign n13531 = ~n13527 & n13530;
  assign n13532 = pi115 & ~n10718;
  assign n13533 = ~pi115 & ~n10728;
  assign n13534 = ~pi39 & ~n13533;
  assign n13535 = ~n13532 & n13534;
  assign n13536 = n3207 & ~n13535;
  assign n13537 = pi115 & ~n10557;
  assign n13538 = n13438 & ~n13537;
  assign n13539 = ~n13519 & n13538;
  assign n13540 = ~pi39 & ~n13525;
  assign n13541 = ~n13539 & n13540;
  assign n13542 = n6251 & ~n13541;
  assign n13543 = pi38 & ~n13528;
  assign n13544 = ~pi87 & ~n13543;
  assign n13545 = ~n13542 & n13544;
  assign n13546 = ~n13536 & n13545;
  assign n13547 = ~n13503 & n13524;
  assign n13548 = n3207 & ~n13547;
  assign n13549 = ~n10581 & n13548;
  assign n13550 = ~n3207 & ~n13528;
  assign n13551 = n11104 & ~n13550;
  assign n13552 = ~n13549 & n13551;
  assign n13553 = ~pi75 & ~n13552;
  assign n13554 = ~n13546 & n13553;
  assign n13555 = ~n13531 & ~n13554;
  assign n13556 = n8867 & ~n13555;
  assign n13557 = ~n8867 & ~n13528;
  assign po273 = ~n13556 & ~n13557;
  assign n13559 = pi116 & n10488;
  assign n13560 = ~n2734 & ~n13559;
  assign n13561 = n2734 & ~n10472;
  assign n13562 = pi116 & ~n13561;
  assign n13563 = ~n10479 & ~n13562;
  assign n13564 = ~n13560 & ~n13563;
  assign n13565 = ~n2734 & n10493;
  assign n13566 = pi228 & ~n13565;
  assign n13567 = ~n13564 & n13566;
  assign n13568 = pi116 & ~n10506;
  assign n13569 = n10722 & ~n13568;
  assign n13570 = ~pi39 & ~n13569;
  assign n13571 = ~n13567 & n13570;
  assign n13572 = n3207 & ~n13571;
  assign n13573 = ~pi72 & pi116;
  assign n13574 = ~n13438 & n13573;
  assign n13575 = ~pi113 & n13439;
  assign n13576 = n13573 & ~n13575;
  assign n13577 = ~n10550 & ~n13576;
  assign n13578 = n13443 & ~n13577;
  assign n13579 = ~n13574 & ~n13578;
  assign n13580 = ~pi39 & ~n13579;
  assign n13581 = n6251 & ~n13580;
  assign n13582 = ~pi39 & n13573;
  assign n13583 = pi38 & ~n13582;
  assign n13584 = ~pi87 & ~n13583;
  assign n13585 = ~n13581 & n13584;
  assign n13586 = ~n13572 & n13585;
  assign n13587 = ~pi113 & n10584;
  assign n13588 = n13573 & ~n13587;
  assign n13589 = ~pi38 & ~n13588;
  assign n13590 = ~n10580 & n13589;
  assign n13591 = ~n13583 & ~n13590;
  assign n13592 = ~pi100 & ~n13591;
  assign n13593 = pi100 & ~n13582;
  assign n13594 = n11104 & ~n13593;
  assign n13595 = ~n13592 & n13594;
  assign n13596 = ~pi75 & ~n13595;
  assign n13597 = ~n13586 & n13596;
  assign n13598 = ~n10598 & n13573;
  assign n13599 = ~n10776 & ~n13598;
  assign n13600 = n13443 & ~n13599;
  assign n13601 = ~n13574 & ~n13600;
  assign n13602 = n3223 & ~n13601;
  assign n13603 = ~n3242 & n13582;
  assign n13604 = pi75 & ~n13603;
  assign n13605 = ~n13602 & n13604;
  assign n13606 = ~n13597 & ~n13605;
  assign n13607 = n8867 & ~n13606;
  assign n13608 = ~n8867 & ~n13582;
  assign po274 = ~n13607 & ~n13608;
  assign n13610 = n3665 & n7354;
  assign n13611 = ~n3664 & ~n13610;
  assign n13612 = ~pi38 & ~n13611;
  assign n13613 = ~pi87 & ~n13612;
  assign n13614 = n6278 & ~n13613;
  assign n13615 = ~pi92 & ~n13614;
  assign n13616 = ~pi54 & ~n7295;
  assign n13617 = ~pi74 & n13616;
  assign n13618 = ~n13615 & n13617;
  assign n13619 = ~pi55 & ~n13618;
  assign n13620 = ~n7337 & ~n13619;
  assign n13621 = ~pi56 & ~n13620;
  assign n13622 = ~n6112 & ~n13621;
  assign n13623 = ~pi62 & ~n13622;
  assign n13624 = ~pi57 & n6289;
  assign po275 = ~n13623 & n13624;
  assign n13626 = pi163 & n6170;
  assign n13627 = ~n11654 & ~n13626;
  assign n13628 = ~pi150 & ~n13627;
  assign n13629 = pi150 & n9684;
  assign n13630 = n11652 & n13629;
  assign n13631 = ~n13628 & ~n13630;
  assign n13632 = pi232 & ~n13631;
  assign n13633 = ~n8975 & n13632;
  assign n13634 = pi74 & ~n13633;
  assign n13635 = pi165 & n7484;
  assign n13636 = ~pi38 & ~pi54;
  assign n13637 = ~n13635 & ~n13636;
  assign n13638 = n8975 & n13637;
  assign n13639 = ~pi74 & ~n13633;
  assign n13640 = ~n13638 & n13639;
  assign n13641 = ~n13634 & ~n13640;
  assign n13642 = ~n3294 & ~n13641;
  assign n13643 = n3432 & ~n13642;
  assign n13644 = ~n9707 & ~n13643;
  assign n13645 = pi299 & n13631;
  assign n13646 = ~pi184 & ~n11667;
  assign n13647 = pi185 & ~n13646;
  assign n13648 = ~pi185 & n13646;
  assign n13649 = n6170 & ~n13647;
  assign n13650 = ~n13648 & n13649;
  assign n13651 = ~pi299 & ~n13650;
  assign n13652 = pi232 & ~n13651;
  assign n13653 = ~n13645 & n13652;
  assign n13654 = ~n8975 & n13653;
  assign n13655 = pi74 & ~n13654;
  assign n13656 = ~pi55 & ~n13655;
  assign n13657 = ~pi143 & ~pi299;
  assign n13658 = ~pi165 & pi299;
  assign n13659 = ~n13657 & ~n13658;
  assign n13660 = n7484 & n13659;
  assign n13661 = n8975 & ~n13660;
  assign n13662 = pi54 & ~n13661;
  assign n13663 = ~n13654 & n13662;
  assign n13664 = ~pi143 & ~n9011;
  assign n13665 = pi143 & ~n9013;
  assign n13666 = pi165 & ~n13665;
  assign n13667 = ~n13664 & n13666;
  assign n13668 = pi143 & ~pi165;
  assign n13669 = n9018 & n13668;
  assign n13670 = pi38 & ~n13669;
  assign n13671 = ~n13667 & n13670;
  assign n13672 = n3241 & ~n13671;
  assign n13673 = ~n6170 & n9304;
  assign n13674 = pi151 & ~pi168;
  assign n13675 = ~n9385 & n13674;
  assign n13676 = pi168 & n9376;
  assign n13677 = ~pi168 & n9379;
  assign n13678 = ~pi151 & ~n13677;
  assign n13679 = ~n13676 & n13678;
  assign n13680 = ~n13675 & ~n13679;
  assign n13681 = ~n13673 & ~n13680;
  assign n13682 = ~n6170 & ~n9304;
  assign n13683 = n6170 & ~n9346;
  assign n13684 = ~n13682 & ~n13683;
  assign n13685 = pi151 & pi168;
  assign n13686 = ~n13684 & n13685;
  assign n13687 = pi150 & ~n13686;
  assign n13688 = ~n13681 & n13687;
  assign n13689 = ~n9217 & ~n13682;
  assign n13690 = pi168 & n13689;
  assign n13691 = ~n9417 & ~n13682;
  assign n13692 = ~pi168 & n13691;
  assign n13693 = pi151 & ~n13692;
  assign n13694 = ~n13690 & n13693;
  assign n13695 = pi168 & n6170;
  assign n13696 = n9304 & ~n13695;
  assign n13697 = pi168 & n9278;
  assign n13698 = ~pi151 & ~n13696;
  assign n13699 = ~n13697 & n13698;
  assign n13700 = ~pi150 & ~n13699;
  assign n13701 = ~n13694 & n13700;
  assign n13702 = pi299 & ~n13701;
  assign n13703 = ~n13688 & n13702;
  assign n13704 = ~n9269 & ~n13673;
  assign n13705 = ~pi173 & ~n13704;
  assign n13706 = n6170 & ~n9161;
  assign n13707 = pi173 & ~n13682;
  assign n13708 = ~n13706 & n13707;
  assign n13709 = pi185 & ~n13708;
  assign n13710 = ~n13705 & n13709;
  assign n13711 = pi173 & n13689;
  assign n13712 = ~n9278 & ~n13673;
  assign n13713 = ~pi173 & ~n13712;
  assign n13714 = ~pi185 & ~n13713;
  assign n13715 = ~n13711 & n13714;
  assign n13716 = pi190 & ~n13715;
  assign n13717 = ~n13710 & n13716;
  assign n13718 = pi173 & ~n9774;
  assign n13719 = ~pi173 & ~n9299;
  assign n13720 = n6170 & ~n13719;
  assign n13721 = ~n13718 & n13720;
  assign n13722 = pi185 & ~n13673;
  assign n13723 = ~n13721 & n13722;
  assign n13724 = pi173 & n13691;
  assign n13725 = ~pi173 & n9304;
  assign n13726 = ~pi185 & ~n13725;
  assign n13727 = ~n13724 & n13726;
  assign n13728 = ~pi190 & ~n13727;
  assign n13729 = ~n13723 & n13728;
  assign n13730 = ~pi299 & ~n13729;
  assign n13731 = ~n13717 & n13730;
  assign n13732 = pi232 & ~n13731;
  assign n13733 = ~n13703 & n13732;
  assign n13734 = ~pi232 & n9304;
  assign n13735 = ~pi39 & ~n13734;
  assign n13736 = ~n13733 & n13735;
  assign n13737 = ~pi178 & ~pi299;
  assign n13738 = pi168 & n9047;
  assign n13739 = pi157 & n9062;
  assign n13740 = ~n13738 & ~n13739;
  assign n13741 = n6170 & n12086;
  assign n13742 = ~n13740 & n13741;
  assign n13743 = pi299 & ~n13742;
  assign n13744 = ~n13737 & ~n13743;
  assign n13745 = n9024 & ~n13744;
  assign n13746 = pi178 & ~n9081;
  assign n13747 = ~pi190 & ~n13746;
  assign n13748 = ~pi299 & ~n13747;
  assign n13749 = ~n13745 & ~n13748;
  assign n13750 = ~n9079 & ~n12097;
  assign n13751 = ~pi178 & ~n13750;
  assign n13752 = ~n9050 & n13751;
  assign n13753 = pi178 & ~n13750;
  assign n13754 = ~n9088 & n13753;
  assign n13755 = ~pi299 & ~n9045;
  assign n13756 = pi190 & n13755;
  assign n13757 = ~n13752 & n13756;
  assign n13758 = ~n13754 & n13757;
  assign n13759 = pi232 & ~n13758;
  assign n13760 = ~n13749 & n13759;
  assign n13761 = ~pi232 & n9024;
  assign n13762 = pi39 & ~n13761;
  assign n13763 = ~n13760 & n13762;
  assign n13764 = ~pi38 & ~n13763;
  assign n13765 = ~n13736 & n13764;
  assign n13766 = n13672 & ~n13765;
  assign n13767 = pi100 & ~n13653;
  assign n13768 = pi38 & ~n13660;
  assign n13769 = n7599 & ~n13768;
  assign n13770 = ~n9504 & n13769;
  assign n13771 = ~n13767 & ~n13770;
  assign n13772 = ~n13766 & n13771;
  assign n13773 = n3238 & ~n13772;
  assign n13774 = pi75 & ~n13653;
  assign n13775 = ~pi100 & ~n13768;
  assign n13776 = ~pi157 & pi299;
  assign n13777 = ~n13737 & ~n13776;
  assign n13778 = n7484 & n13777;
  assign n13779 = n9455 & n13778;
  assign n13780 = n9504 & ~n13779;
  assign n13781 = n13775 & ~n13780;
  assign n13782 = ~n13767 & ~n13781;
  assign n13783 = n9450 & ~n13782;
  assign n13784 = ~n13774 & ~n13783;
  assign n13785 = ~n13773 & n13784;
  assign n13786 = ~pi54 & ~n13785;
  assign n13787 = ~n13663 & ~n13786;
  assign n13788 = ~pi74 & ~n13787;
  assign n13789 = n13656 & ~n13788;
  assign n13790 = pi55 & ~n13634;
  assign n13791 = pi150 & n7484;
  assign n13792 = ~pi92 & n9455;
  assign n13793 = n13791 & n13792;
  assign n13794 = n9024 & n13636;
  assign n13795 = ~n13793 & n13794;
  assign n13796 = ~n13637 & ~n13795;
  assign n13797 = n8975 & ~n13796;
  assign n13798 = n13639 & ~n13797;
  assign n13799 = n13790 & ~n13798;
  assign n13800 = n3294 & ~n13799;
  assign n13801 = ~n13789 & n13800;
  assign n13802 = ~n13644 & ~n13801;
  assign n13803 = ~n8975 & ~n13632;
  assign n13804 = n8975 & n13635;
  assign n13805 = ~n3432 & ~n13804;
  assign n13806 = ~n13803 & n13805;
  assign n13807 = ~n13634 & n13806;
  assign n13808 = ~n13802 & ~n13807;
  assign n13809 = pi118 & n13808;
  assign n13810 = ~pi79 & n12145;
  assign n13811 = n6206 & ~n6455;
  assign n13812 = ~pi157 & n9519;
  assign n13813 = pi168 & ~n13812;
  assign n13814 = pi157 & ~n9514;
  assign n13815 = ~pi157 & ~pi168;
  assign n13816 = ~n9512 & n13815;
  assign n13817 = ~n13814 & ~n13816;
  assign n13818 = ~n13813 & n13817;
  assign n13819 = ~n13811 & ~n13818;
  assign n13820 = n13094 & ~n13819;
  assign n13821 = ~pi178 & ~n6197;
  assign n13822 = n9518 & n13821;
  assign n13823 = ~n13811 & ~n13822;
  assign n13824 = pi190 & ~n13823;
  assign n13825 = pi178 & ~n9525;
  assign n13826 = ~n13811 & n13825;
  assign n13827 = ~pi178 & ~n13128;
  assign n13828 = ~pi190 & ~n13826;
  assign n13829 = ~n13827 & n13828;
  assign n13830 = ~n13824 & ~n13829;
  assign n13831 = n13096 & ~n13830;
  assign n13832 = pi232 & ~n13831;
  assign n13833 = ~n13820 & n13832;
  assign n13834 = n7299 & n9530;
  assign n13835 = ~n6229 & n13094;
  assign n13836 = ~n6455 & n13835;
  assign n13837 = ~pi232 & ~n13836;
  assign n13838 = ~n13834 & n13837;
  assign n13839 = pi39 & ~n13838;
  assign n13840 = ~n13833 & n13839;
  assign n13841 = n9592 & n13674;
  assign n13842 = pi168 & ~n9578;
  assign n13843 = ~pi168 & ~n9564;
  assign n13844 = ~pi151 & ~n13842;
  assign n13845 = ~n13843 & n13844;
  assign n13846 = ~n13841 & ~n13845;
  assign n13847 = n9566 & ~n13846;
  assign n13848 = pi150 & ~n13847;
  assign n13849 = ~pi151 & n9553;
  assign n13850 = n9606 & ~n13849;
  assign n13851 = ~pi168 & ~n13850;
  assign n13852 = ~pi151 & n9574;
  assign n13853 = n9609 & ~n13852;
  assign n13854 = n13695 & ~n13853;
  assign n13855 = ~pi150 & ~n13854;
  assign n13856 = ~n13851 & n13855;
  assign n13857 = ~n13848 & ~n13856;
  assign n13858 = ~n9553 & ~n12011;
  assign n13859 = ~n6170 & ~n13858;
  assign n13860 = pi299 & ~n13859;
  assign n13861 = ~n13857 & n13860;
  assign n13862 = n6371 & n9592;
  assign n13863 = pi173 & n13862;
  assign n13864 = ~pi173 & n6371;
  assign n13865 = n9564 & n13864;
  assign n13866 = ~n13863 & ~n13865;
  assign n13867 = ~pi190 & n6170;
  assign n13868 = ~n13866 & n13867;
  assign n13869 = ~pi173 & pi190;
  assign n13870 = n9579 & n13869;
  assign n13871 = pi185 & ~n13870;
  assign n13872 = ~n13868 & n13871;
  assign n13873 = ~pi173 & n9553;
  assign n13874 = n9585 & ~n13873;
  assign n13875 = ~pi190 & ~n13874;
  assign n13876 = pi173 & n9588;
  assign n13877 = pi190 & n9576;
  assign n13878 = ~n13876 & n13877;
  assign n13879 = ~pi185 & ~n13878;
  assign n13880 = ~n13875 & n13879;
  assign n13881 = ~n13872 & ~n13880;
  assign n13882 = ~n6170 & ~n9557;
  assign n13883 = ~pi299 & ~n13882;
  assign n13884 = ~n13881 & n13883;
  assign n13885 = ~n13861 & ~n13884;
  assign n13886 = pi232 & ~n13885;
  assign n13887 = ~n6151 & ~n9555;
  assign n13888 = ~pi232 & ~n9553;
  assign n13889 = ~n13887 & n13888;
  assign n13890 = ~pi39 & ~n13889;
  assign n13891 = ~n13886 & n13890;
  assign n13892 = ~n13840 & ~n13891;
  assign n13893 = ~pi38 & ~n13892;
  assign n13894 = n13672 & ~n13893;
  assign n13895 = ~n13767 & ~n13769;
  assign n13896 = ~n13894 & n13895;
  assign n13897 = n3238 & ~n13896;
  assign n13898 = n8951 & ~n13778;
  assign n13899 = n3096 & n13898;
  assign n13900 = n13775 & ~n13899;
  assign n13901 = ~n13767 & ~n13900;
  assign n13902 = n9450 & ~n13901;
  assign n13903 = ~n13774 & ~n13902;
  assign n13904 = ~n13897 & n13903;
  assign n13905 = ~pi54 & ~n13904;
  assign n13906 = ~n13663 & ~n13905;
  assign n13907 = ~pi74 & ~n13906;
  assign n13908 = n13656 & ~n13907;
  assign n13909 = pi54 & n13635;
  assign n13910 = ~pi92 & n8975;
  assign n13911 = n8951 & n13910;
  assign n13912 = ~n13791 & n13911;
  assign n13913 = ~n13909 & n13912;
  assign n13914 = n3096 & n13913;
  assign n13915 = n13640 & ~n13914;
  assign n13916 = n13790 & ~n13915;
  assign n13917 = n3294 & ~n13916;
  assign n13918 = ~n13908 & n13917;
  assign n13919 = n13643 & ~n13918;
  assign n13920 = ~n13807 & ~n13919;
  assign n13921 = ~pi118 & n13920;
  assign n13922 = ~n13810 & ~n13921;
  assign n13923 = ~n13809 & n13922;
  assign n13924 = ~pi118 & ~n8962;
  assign n13925 = n13808 & n13924;
  assign n13926 = n13920 & ~n13924;
  assign n13927 = n13810 & ~n13926;
  assign n13928 = ~n13925 & n13927;
  assign po276 = n13923 | n13928;
  assign n13930 = pi128 & pi228;
  assign n13931 = ~n10144 & n13930;
  assign n13932 = ~n3053 & n3483;
  assign n13933 = n7534 & n13932;
  assign n13934 = ~n3461 & n5774;
  assign n13935 = n7531 & n13934;
  assign n13936 = ~n13933 & ~n13935;
  assign n13937 = pi39 & ~n13936;
  assign n13938 = n2579 & n10138;
  assign n13939 = n11640 & ~n13938;
  assign n13940 = n2592 & ~n13939;
  assign n13941 = ~pi97 & ~n13940;
  assign n13942 = ~pi46 & n2796;
  assign n13943 = n2758 & n13942;
  assign n13944 = ~n13941 & n13943;
  assign n13945 = pi299 & n6310;
  assign n13946 = ~n6422 & ~n13945;
  assign n13947 = n7484 & ~n13946;
  assign n13948 = pi109 & ~n13947;
  assign n13949 = ~n2796 & n11641;
  assign n13950 = ~n13948 & ~n13949;
  assign n13951 = ~n13944 & n13950;
  assign n13952 = ~n6312 & ~n13947;
  assign n13953 = ~n6383 & n13947;
  assign n13954 = ~n13952 & ~n13953;
  assign n13955 = ~n13951 & n13954;
  assign n13956 = ~pi91 & ~n13955;
  assign n13957 = n2534 & ~n6347;
  assign n13958 = ~n13956 & n13957;
  assign n13959 = ~n2563 & ~n13958;
  assign n13960 = ~pi39 & n11063;
  assign n13961 = ~n13959 & n13960;
  assign n13962 = ~n13937 & ~n13961;
  assign n13963 = ~pi38 & ~n13962;
  assign n13964 = ~pi228 & n13963;
  assign n13965 = ~n13930 & ~n13964;
  assign n13966 = ~pi100 & ~n13965;
  assign n13967 = n3182 & n3322;
  assign n13968 = ~n13930 & ~n13967;
  assign n13969 = pi100 & ~n13968;
  assign n13970 = ~pi87 & ~n13969;
  assign n13971 = ~n13966 & n13970;
  assign n13972 = pi87 & ~n13930;
  assign n13973 = ~pi75 & ~n13972;
  assign n13974 = ~n13971 & n13973;
  assign n13975 = n7359 & n8951;
  assign n13976 = ~n13930 & ~n13975;
  assign n13977 = pi75 & ~n13976;
  assign n13978 = ~pi92 & ~n13977;
  assign n13979 = ~n13974 & n13978;
  assign n13980 = pi92 & ~n13930;
  assign n13981 = ~n7372 & n13980;
  assign n13982 = n10144 & ~n13981;
  assign n13983 = ~n13979 & n13982;
  assign po277 = n13931 | n13983;
  assign n13985 = ~pi31 & ~pi80;
  assign n13986 = pi818 & n13985;
  assign n13987 = ~n7444 & n8044;
  assign n13988 = ~n7720 & ~n13987;
  assign n13989 = ~pi120 & ~n7444;
  assign n13990 = ~pi1093 & n13989;
  assign n13991 = n13988 & ~n13990;
  assign n13992 = n3096 & n7490;
  assign n13993 = pi120 & ~n8044;
  assign n13994 = ~n7550 & n13993;
  assign n13995 = n13992 & ~n13994;
  assign n13996 = ~pi120 & pi1093;
  assign n13997 = n7550 & ~n13996;
  assign n13998 = ~n13995 & ~n13997;
  assign n13999 = n3182 & n8087;
  assign n14000 = ~n13998 & n13999;
  assign n14001 = ~n8044 & n13996;
  assign n14002 = ~n13993 & ~n14001;
  assign n14003 = pi100 & ~n14002;
  assign n14004 = ~n14000 & n14003;
  assign n14005 = ~pi1093 & n7474;
  assign n14006 = pi120 & n14005;
  assign n14007 = ~pi39 & ~n14006;
  assign n14008 = n7514 & ~n10332;
  assign n14009 = n7465 & n7496;
  assign n14010 = ~pi829 & n14009;
  assign n14011 = ~pi122 & ~n14010;
  assign n14012 = ~n14008 & n14011;
  assign n14013 = pi122 & ~n7466;
  assign n14014 = ~n2733 & ~n14013;
  assign n14015 = ~n14012 & n14014;
  assign n14016 = n10053 & ~n14015;
  assign n14017 = n7558 & ~n14009;
  assign n14018 = ~n12771 & n14017;
  assign n14019 = ~n14016 & ~n14018;
  assign n14020 = n14007 & n14019;
  assign n14021 = ~n6206 & n14002;
  assign n14022 = ~n7530 & n13993;
  assign n14023 = pi1091 & pi1092;
  assign n14024 = n7528 & n14023;
  assign n14025 = n14001 & ~n14024;
  assign n14026 = ~n14022 & ~n14025;
  assign n14027 = n6206 & n14026;
  assign n14028 = ~n14021 & ~n14027;
  assign n14029 = n6223 & n14028;
  assign n14030 = n6200 & ~n14002;
  assign n14031 = ~n6200 & ~n14026;
  assign n14032 = ~n14030 & ~n14031;
  assign n14033 = ~n6223 & ~n14032;
  assign n14034 = n8074 & ~n14029;
  assign n14035 = ~n14033 & n14034;
  assign n14036 = ~n8074 & n14002;
  assign n14037 = pi299 & ~n14036;
  assign n14038 = ~n14035 & n14037;
  assign n14039 = n6197 & n14028;
  assign n14040 = ~n6197 & ~n14032;
  assign n14041 = n8066 & ~n14039;
  assign n14042 = ~n14040 & n14041;
  assign n14043 = ~n8066 & n14002;
  assign n14044 = ~pi299 & ~n14043;
  assign n14045 = ~n14042 & n14044;
  assign n14046 = pi39 & ~n14038;
  assign n14047 = ~n14045 & n14046;
  assign n14048 = ~n14020 & ~n14047;
  assign n14049 = ~pi38 & ~n14048;
  assign n14050 = pi38 & n8044;
  assign n14051 = ~pi120 & ~pi1093;
  assign n14052 = pi38 & n14051;
  assign n14053 = ~pi100 & ~n14052;
  assign n14054 = ~n14050 & n14053;
  assign n14055 = ~n14049 & n14054;
  assign n14056 = ~n14004 & ~n14055;
  assign n14057 = ~pi87 & ~n14056;
  assign n14058 = n7566 & ~n14051;
  assign n14059 = n7558 & ~n12771;
  assign n14060 = ~n8099 & n14059;
  assign n14061 = n7564 & ~n14060;
  assign n14062 = ~n3208 & n8044;
  assign n14063 = pi87 & ~n14062;
  assign n14064 = ~n14061 & n14063;
  assign n14065 = n14058 & n14064;
  assign n14066 = ~n14057 & ~n14065;
  assign n14067 = ~pi75 & ~n14066;
  assign n14068 = n7485 & n14002;
  assign n14069 = ~n7491 & n14001;
  assign n14070 = ~pi1091 & ~n8043;
  assign n14071 = ~n8036 & ~n14070;
  assign n14072 = pi120 & ~n14071;
  assign n14073 = ~n7485 & ~n14072;
  assign n14074 = ~n14069 & n14073;
  assign n14075 = ~n14068 & ~n14074;
  assign n14076 = n3223 & ~n14075;
  assign n14077 = ~n3223 & n14002;
  assign n14078 = pi75 & ~n14077;
  assign n14079 = ~n14076 & n14078;
  assign n14080 = n7444 & ~n14079;
  assign n14081 = ~n14067 & n14080;
  assign n14082 = n13991 & ~n14081;
  assign n14083 = ~n14016 & ~n14017;
  assign n14084 = n14007 & n14083;
  assign n14085 = pi1093 & ~n6206;
  assign n14086 = n6223 & n14085;
  assign n14087 = n6200 & ~n6223;
  assign n14088 = n8074 & ~n14087;
  assign n14089 = ~n14086 & n14088;
  assign n14090 = n7530 & n14089;
  assign n14091 = pi299 & ~n14051;
  assign n14092 = ~n14090 & n14091;
  assign n14093 = n6197 & n14085;
  assign n14094 = ~n6197 & n6200;
  assign n14095 = n8066 & ~n14094;
  assign n14096 = ~n14093 & n14095;
  assign n14097 = n7530 & n14096;
  assign n14098 = ~pi299 & ~n14051;
  assign n14099 = ~n14097 & n14098;
  assign n14100 = pi39 & ~n14092;
  assign n14101 = ~n14099 & n14100;
  assign n14102 = ~n14084 & ~n14101;
  assign n14103 = ~pi38 & ~n14102;
  assign n14104 = n14053 & ~n14103;
  assign n14105 = pi120 & n7550;
  assign n14106 = ~pi120 & n13992;
  assign n14107 = ~n14105 & ~n14106;
  assign n14108 = n13999 & ~n14107;
  assign n14109 = pi100 & ~n14051;
  assign n14110 = ~n14108 & n14109;
  assign n14111 = ~n14104 & ~n14110;
  assign n14112 = ~pi87 & ~n14111;
  assign n14113 = ~n14058 & ~n14112;
  assign n14114 = ~pi75 & ~n14113;
  assign n14115 = n7494 & ~n14051;
  assign n14116 = n7444 & ~n14115;
  assign n14117 = ~n14114 & n14116;
  assign n14118 = n7720 & ~n13990;
  assign n14119 = ~n14117 & n14118;
  assign n14120 = ~n14082 & ~n14119;
  assign n14121 = n13986 & ~n14120;
  assign n14122 = ~po1038 & ~n14121;
  assign n14123 = ~n7720 & n14002;
  assign n14124 = pi120 & ~n14123;
  assign n14125 = n13986 & ~n14051;
  assign n14126 = ~n14123 & n14125;
  assign n14127 = po1038 & ~n14126;
  assign n14128 = ~n14124 & n14127;
  assign n14129 = ~n8856 & ~n14128;
  assign n14130 = pi951 & pi982;
  assign n14131 = pi1092 & n14130;
  assign n14132 = pi1093 & n14131;
  assign n14133 = ~pi120 & ~n14132;
  assign n14134 = ~n14123 & ~n14133;
  assign n14135 = n14127 & ~n14134;
  assign n14136 = n8856 & ~n14135;
  assign n14137 = ~n14129 & ~n14136;
  assign n14138 = ~n14122 & ~n14137;
  assign n14139 = pi120 & n7492;
  assign n14140 = ~pi1091 & n14132;
  assign n14141 = ~pi120 & ~n14140;
  assign n14142 = n10053 & n14131;
  assign n14143 = ~pi93 & ~pi122;
  assign n14144 = n2549 & n14143;
  assign n14145 = n2754 & n8880;
  assign n14146 = n14144 & n14145;
  assign n14147 = n2536 & n14146;
  assign n14148 = n10290 & n14147;
  assign n14149 = n7488 & n14148;
  assign n14150 = n2492 & n14149;
  assign n14151 = n14142 & ~n14150;
  assign n14152 = n14141 & ~n14151;
  assign n14153 = ~n14139 & ~n14152;
  assign n14154 = ~n7485 & ~n14153;
  assign n14155 = n7485 & n14133;
  assign n14156 = n3223 & ~n14155;
  assign n14157 = ~n14154 & n14156;
  assign n14158 = ~n3223 & ~n14133;
  assign n14159 = pi75 & ~n14158;
  assign n14160 = ~n14157 & n14159;
  assign n14161 = pi950 & n3096;
  assign n14162 = n7470 & n7488;
  assign n14163 = n14161 & n14162;
  assign n14164 = n14142 & ~n14163;
  assign n14165 = n14141 & ~n14164;
  assign n14166 = ~n14105 & ~n14165;
  assign n14167 = ~pi39 & n8087;
  assign n14168 = ~n14166 & n14167;
  assign n14169 = pi100 & ~n14168;
  assign n14170 = ~pi38 & ~n14169;
  assign n14171 = ~n13999 & n14133;
  assign n14172 = ~n14170 & ~n14171;
  assign n14173 = ~n8066 & n14133;
  assign n14174 = ~pi299 & ~n14173;
  assign n14175 = ~n8261 & ~n14133;
  assign n14176 = ~n6197 & n14175;
  assign n14177 = ~n8258 & ~n14133;
  assign n14178 = n6197 & n14177;
  assign n14179 = n8066 & ~n14176;
  assign n14180 = ~n14178 & n14179;
  assign n14181 = n14174 & ~n14180;
  assign n14182 = ~n8074 & n14133;
  assign n14183 = pi299 & ~n14182;
  assign n14184 = ~n6223 & n14175;
  assign n14185 = n6223 & n14177;
  assign n14186 = n8074 & ~n14184;
  assign n14187 = ~n14185 & n14186;
  assign n14188 = n14183 & ~n14187;
  assign n14189 = ~n14181 & ~n14188;
  assign n14190 = pi39 & ~n14189;
  assign n14191 = n2580 & n7454;
  assign n14192 = n2576 & n14191;
  assign n14193 = ~pi97 & ~n14192;
  assign n14194 = n2762 & ~n14193;
  assign n14195 = n2759 & n14194;
  assign n14196 = ~n7501 & ~n14195;
  assign n14197 = n2518 & ~n14196;
  assign n14198 = n7448 & ~n14197;
  assign n14199 = n7445 & ~n14198;
  assign n14200 = ~pi51 & ~n14199;
  assign n14201 = ~n2558 & ~n14200;
  assign n14202 = ~pi96 & ~n14201;
  assign n14203 = ~pi72 & pi950;
  assign n14204 = n10333 & n14203;
  assign n14205 = ~n14202 & n14204;
  assign n14206 = n7470 & n14131;
  assign n14207 = ~n14205 & n14206;
  assign n14208 = n9545 & n14192;
  assign n14209 = n7445 & n14208;
  assign n14210 = n7450 & ~n14209;
  assign n14211 = pi950 & n7497;
  assign n14212 = ~n14210 & n14211;
  assign n14213 = pi824 & n14212;
  assign n14214 = n14131 & ~n14213;
  assign n14215 = ~pi829 & n14214;
  assign n14216 = pi829 & pi1092;
  assign n14217 = pi122 & n14130;
  assign n14218 = n14216 & n14217;
  assign n14219 = ~n14212 & n14218;
  assign n14220 = ~n14215 & ~n14219;
  assign n14221 = ~n14207 & n14220;
  assign n14222 = n7495 & ~n14221;
  assign n14223 = n2733 & n14132;
  assign n14224 = ~n14222 & ~n14223;
  assign n14225 = pi1091 & ~n14224;
  assign n14226 = n14140 & ~n14213;
  assign n14227 = ~pi120 & ~n14226;
  assign n14228 = ~n14225 & n14227;
  assign n14229 = ~n14005 & n14083;
  assign n14230 = pi120 & n14229;
  assign n14231 = ~pi39 & ~n14228;
  assign n14232 = ~n14230 & n14231;
  assign n14233 = ~n14190 & ~n14232;
  assign n14234 = n3207 & ~n14233;
  assign n14235 = ~n14172 & ~n14234;
  assign n14236 = ~pi87 & ~n14235;
  assign n14237 = ~n3208 & n14133;
  assign n14238 = pi87 & ~n14237;
  assign n14239 = ~n2733 & ~n6179;
  assign n14240 = n14161 & n14239;
  assign n14241 = n14142 & ~n14240;
  assign n14242 = pi824 & n14161;
  assign n14243 = n14140 & ~n14242;
  assign n14244 = ~n14241 & ~n14243;
  assign n14245 = ~pi120 & ~n14244;
  assign n14246 = ~n7559 & ~n7563;
  assign n14247 = pi120 & ~n14246;
  assign n14248 = n3208 & ~n14247;
  assign n14249 = ~n14245 & n14248;
  assign n14250 = n14238 & ~n14249;
  assign n14251 = ~pi75 & ~n14250;
  assign n14252 = ~n14236 & n14251;
  assign n14253 = ~n14160 & ~n14252;
  assign n14254 = n7444 & ~n14253;
  assign n14255 = n7720 & ~n14254;
  assign n14256 = ~n12771 & n14140;
  assign n14257 = ~n14164 & ~n14256;
  assign n14258 = ~pi120 & ~n14257;
  assign n14259 = ~n13994 & ~n14258;
  assign n14260 = n8087 & ~n14259;
  assign n14261 = ~n14002 & ~n14133;
  assign n14262 = ~n8087 & n14261;
  assign n14263 = n3182 & ~n14262;
  assign n14264 = ~n14260 & n14263;
  assign n14265 = ~n3182 & ~n14261;
  assign n14266 = pi100 & ~n14265;
  assign n14267 = ~n14264 & n14266;
  assign n14268 = ~n14005 & n14019;
  assign n14269 = pi120 & n14268;
  assign n14270 = n14059 & n14214;
  assign n14271 = ~pi120 & ~n14270;
  assign n14272 = ~n14225 & n14271;
  assign n14273 = ~n14269 & ~n14272;
  assign n14274 = ~pi39 & ~n14273;
  assign n14275 = ~n7528 & n14142;
  assign n14276 = ~n14256 & ~n14275;
  assign n14277 = ~pi120 & ~n14276;
  assign n14278 = ~n14022 & ~n14277;
  assign n14279 = n6206 & ~n14278;
  assign n14280 = ~n6206 & n14261;
  assign n14281 = ~n14279 & ~n14280;
  assign n14282 = n6197 & ~n14281;
  assign n14283 = ~n6200 & ~n14278;
  assign n14284 = n6200 & n14261;
  assign n14285 = ~n14283 & ~n14284;
  assign n14286 = ~n6197 & ~n14285;
  assign n14287 = n8066 & ~n14282;
  assign n14288 = ~n14286 & n14287;
  assign n14289 = ~n14043 & n14174;
  assign n14290 = ~n14288 & n14289;
  assign n14291 = n6223 & ~n14281;
  assign n14292 = ~n6223 & ~n14285;
  assign n14293 = n8074 & ~n14291;
  assign n14294 = ~n14292 & n14293;
  assign n14295 = n8044 & ~n8074;
  assign n14296 = n14183 & ~n14295;
  assign n14297 = ~n14294 & n14296;
  assign n14298 = pi39 & ~n14290;
  assign n14299 = ~n14297 & n14298;
  assign n14300 = ~n14274 & ~n14299;
  assign n14301 = ~pi38 & ~n14300;
  assign n14302 = pi38 & ~n14261;
  assign n14303 = ~pi100 & ~n14302;
  assign n14304 = ~n14301 & n14303;
  assign n14305 = ~n14267 & ~n14304;
  assign n14306 = ~pi87 & ~n14305;
  assign n14307 = ~n14061 & ~n14248;
  assign n14308 = ~n14241 & ~n14256;
  assign n14309 = n14245 & ~n14308;
  assign n14310 = ~n14307 & ~n14309;
  assign n14311 = ~n14062 & n14238;
  assign n14312 = ~n14310 & n14311;
  assign n14313 = ~n14306 & ~n14312;
  assign n14314 = ~pi75 & ~n14313;
  assign n14315 = n7485 & ~n14261;
  assign n14316 = ~n14151 & ~n14256;
  assign n14317 = ~pi120 & ~n14316;
  assign n14318 = n14073 & ~n14317;
  assign n14319 = ~n14315 & ~n14318;
  assign n14320 = n3223 & ~n14319;
  assign n14321 = ~n3223 & ~n14261;
  assign n14322 = pi75 & ~n14321;
  assign n14323 = ~n14320 & n14322;
  assign n14324 = n7444 & ~n14323;
  assign n14325 = ~n14314 & n14324;
  assign n14326 = n13991 & ~n14325;
  assign n14327 = ~n14255 & ~n14326;
  assign n14328 = n13989 & ~n14132;
  assign n14329 = n14136 & ~n14328;
  assign n14330 = ~n14327 & n14329;
  assign n14331 = n7554 & ~n8044;
  assign n14332 = ~pi39 & ~n14268;
  assign n14333 = ~n8044 & ~n8258;
  assign n14334 = n6197 & n14333;
  assign n14335 = ~n8044 & ~n8261;
  assign n14336 = ~n6197 & n14335;
  assign n14337 = n8066 & ~n14334;
  assign n14338 = ~n14336 & n14337;
  assign n14339 = n8044 & ~n8066;
  assign n14340 = ~pi299 & ~n14339;
  assign n14341 = ~n14338 & n14340;
  assign n14342 = n6223 & n14333;
  assign n14343 = ~n6223 & n14335;
  assign n14344 = n8074 & ~n14342;
  assign n14345 = ~n14343 & n14344;
  assign n14346 = pi299 & ~n14295;
  assign n14347 = ~n14345 & n14346;
  assign n14348 = ~n14341 & ~n14347;
  assign n14349 = pi39 & ~n14348;
  assign n14350 = ~pi38 & ~n14349;
  assign n14351 = ~n14332 & n14350;
  assign n14352 = ~pi100 & ~n14050;
  assign n14353 = ~n14351 & n14352;
  assign n14354 = ~n14331 & ~n14353;
  assign n14355 = ~pi87 & ~n14354;
  assign n14356 = ~n14064 & ~n14355;
  assign n14357 = ~pi75 & ~n14356;
  assign n14358 = n7486 & n14071;
  assign n14359 = ~n7486 & n8044;
  assign n14360 = pi75 & ~n14359;
  assign n14361 = ~n14358 & n14360;
  assign n14362 = ~n14357 & ~n14361;
  assign n14363 = n13988 & ~n14362;
  assign n14364 = ~pi39 & ~n14229;
  assign n14365 = n7540 & ~n14364;
  assign n14366 = ~pi100 & ~n14365;
  assign n14367 = ~n7554 & ~n14366;
  assign n14368 = ~pi87 & ~n14367;
  assign n14369 = ~n7566 & ~n14368;
  assign n14370 = ~pi75 & ~n14369;
  assign n14371 = ~n7494 & ~n14370;
  assign n14372 = n7720 & ~n13989;
  assign n14373 = ~n14371 & n14372;
  assign n14374 = ~n7444 & ~n14123;
  assign n14375 = ~n14363 & ~n14374;
  assign n14376 = ~n14373 & n14375;
  assign n14377 = pi120 & n14129;
  assign n14378 = ~n14376 & n14377;
  assign n14379 = ~n14330 & ~n14378;
  assign n14380 = ~n13986 & ~n14379;
  assign po278 = n14138 | n14380;
  assign n14382 = ~pi134 & ~pi135;
  assign n14383 = ~pi136 & n14382;
  assign n14384 = ~pi130 & n14383;
  assign n14385 = ~pi132 & n14384;
  assign n14386 = ~pi126 & n14385;
  assign n14387 = ~pi121 & n14386;
  assign n14388 = ~pi125 & ~pi133;
  assign n14389 = pi121 & ~n14388;
  assign n14390 = ~pi121 & n14388;
  assign n14391 = ~n14389 & ~n14390;
  assign n14392 = ~n14387 & ~n14391;
  assign n14393 = n2467 & n10134;
  assign n14394 = ~pi51 & n14393;
  assign n14395 = ~pi87 & n14394;
  assign n14396 = ~n14392 & n14395;
  assign n14397 = pi51 & n6170;
  assign n14398 = ~pi146 & n14397;
  assign n14399 = pi161 & ~n14398;
  assign n14400 = n6170 & ~n14394;
  assign n14401 = pi51 & pi146;
  assign n14402 = ~n14399 & ~n14401;
  assign n14403 = n14400 & n14402;
  assign n14404 = ~pi87 & ~n14403;
  assign n14405 = pi87 & ~n13626;
  assign n14406 = pi232 & ~n14405;
  assign n14407 = ~n14404 & n14406;
  assign n14408 = po1038 & ~n14396;
  assign n14409 = ~n14407 & n14408;
  assign n14410 = ~pi142 & n14397;
  assign n14411 = pi144 & ~n14410;
  assign n14412 = pi51 & pi142;
  assign n14413 = n14400 & ~n14412;
  assign n14414 = ~n14411 & n14413;
  assign n14415 = ~pi299 & ~n14414;
  assign n14416 = pi299 & ~n14403;
  assign n14417 = pi232 & ~n14415;
  assign n14418 = ~n14416 & n14417;
  assign n14419 = pi38 & ~n14418;
  assign n14420 = ~pi100 & ~n14419;
  assign n14421 = pi38 & ~n14394;
  assign n14422 = ~pi100 & ~n14421;
  assign n14423 = ~n14420 & ~n14422;
  assign n14424 = n2456 & n10133;
  assign n14425 = n13013 & n14424;
  assign n14426 = n2579 & n14425;
  assign n14427 = n2494 & n7459;
  assign n14428 = ~pi58 & n14427;
  assign n14429 = n9030 & n14428;
  assign n14430 = n14426 & n14429;
  assign n14431 = pi72 & n6371;
  assign n14432 = n14430 & n14431;
  assign n14433 = ~pi50 & pi77;
  assign n14434 = n2482 & n14433;
  assign n14435 = n14425 & n14434;
  assign n14436 = pi86 & n14426;
  assign n14437 = ~n14435 & ~n14436;
  assign n14438 = n11053 & ~n14437;
  assign n14439 = ~pi24 & n11644;
  assign n14440 = n14426 & n14439;
  assign n14441 = n14393 & ~n14440;
  assign n14442 = ~n14438 & n14441;
  assign n14443 = ~pi51 & ~n14393;
  assign n14444 = ~n2497 & ~n14443;
  assign n14445 = ~n14442 & ~n14444;
  assign n14446 = n3094 & n14445;
  assign n14447 = ~pi24 & pi314;
  assign n14448 = n14427 & n14447;
  assign n14449 = n8885 & n14448;
  assign n14450 = n14435 & n14449;
  assign n14451 = n3094 & n14450;
  assign n14452 = n14394 & ~n14451;
  assign n14453 = ~n14446 & n14452;
  assign n14454 = ~n6170 & ~n14453;
  assign n14455 = ~n14400 & ~n14454;
  assign n14456 = ~n14432 & n14455;
  assign n14457 = pi144 & ~n14456;
  assign n14458 = n14394 & ~n14446;
  assign n14459 = ~n14432 & n14458;
  assign n14460 = ~n14451 & n14459;
  assign n14461 = ~n6170 & ~n14460;
  assign n14462 = pi72 & n10420;
  assign n14463 = ~n14397 & ~n14462;
  assign n14464 = n6170 & ~n14463;
  assign n14465 = ~n14461 & ~n14464;
  assign n14466 = ~pi144 & ~n14465;
  assign n14467 = ~n14457 & ~n14466;
  assign n14468 = ~n14410 & ~n14467;
  assign n14469 = pi180 & ~n14468;
  assign n14470 = ~pi51 & n14448;
  assign n14471 = n13403 & n14470;
  assign n14472 = n3094 & n6170;
  assign n14473 = n14471 & n14472;
  assign n14474 = n14465 & ~n14473;
  assign n14475 = pi142 & n14474;
  assign n14476 = ~n6170 & n14460;
  assign n14477 = ~pi72 & ~n14471;
  assign n14478 = n6372 & ~n14477;
  assign n14479 = n6170 & ~n14478;
  assign n14480 = ~n14476 & ~n14479;
  assign n14481 = ~pi142 & ~n14480;
  assign n14482 = ~pi144 & ~n14481;
  assign n14483 = ~n14475 & n14482;
  assign n14484 = ~n14451 & n14456;
  assign n14485 = n14411 & ~n14484;
  assign n14486 = ~pi180 & ~n14485;
  assign n14487 = ~n14483 & n14486;
  assign n14488 = pi179 & ~n14469;
  assign n14489 = ~n14487 & n14488;
  assign n14490 = ~pi24 & ~n11645;
  assign n14491 = pi24 & ~n11642;
  assign n14492 = ~n14490 & ~n14491;
  assign n14493 = ~pi314 & ~n14492;
  assign n14494 = pi314 & ~n11642;
  assign n14495 = ~n14493 & ~n14494;
  assign n14496 = n7459 & n8946;
  assign n14497 = n14495 & n14496;
  assign n14498 = ~pi51 & ~n14497;
  assign n14499 = ~n14462 & n14498;
  assign n14500 = n6170 & ~n14499;
  assign n14501 = ~n14461 & ~n14500;
  assign n14502 = pi142 & n14501;
  assign n14503 = n2497 & n14495;
  assign n14504 = ~pi72 & ~n14503;
  assign n14505 = n6372 & ~n14504;
  assign n14506 = n6170 & ~n14505;
  assign n14507 = ~n14476 & ~n14506;
  assign n14508 = ~pi142 & ~n14507;
  assign n14509 = ~pi144 & ~n14502;
  assign n14510 = ~n14508 & n14509;
  assign n14511 = n14411 & ~n14460;
  assign n14512 = ~pi180 & ~n14511;
  assign n14513 = ~n14510 & n14512;
  assign n14514 = n2497 & n14492;
  assign n14515 = ~pi72 & ~n14514;
  assign n14516 = n6372 & ~n14515;
  assign n14517 = n6170 & ~n14516;
  assign n14518 = ~n14476 & ~n14517;
  assign n14519 = ~pi142 & ~n14518;
  assign n14520 = n14472 & n14514;
  assign n14521 = ~n14464 & ~n14520;
  assign n14522 = ~n14461 & n14521;
  assign n14523 = pi142 & n14522;
  assign n14524 = ~pi144 & ~n14523;
  assign n14525 = ~n14519 & n14524;
  assign n14526 = ~pi51 & n6170;
  assign n14527 = ~n14459 & n14526;
  assign n14528 = ~n14461 & ~n14527;
  assign n14529 = n6170 & ~n14458;
  assign n14530 = ~pi142 & ~n14529;
  assign n14531 = n6170 & n14443;
  assign n14532 = ~n14472 & ~n14531;
  assign n14533 = n3094 & ~n14445;
  assign n14534 = ~n14532 & ~n14533;
  assign n14535 = pi142 & ~n14534;
  assign n14536 = ~n14530 & ~n14535;
  assign n14537 = ~n14455 & ~n14536;
  assign n14538 = n14528 & ~n14537;
  assign n14539 = pi144 & ~n14538;
  assign n14540 = pi180 & ~n14539;
  assign n14541 = ~n14525 & n14540;
  assign n14542 = ~pi179 & ~n14541;
  assign n14543 = ~n14513 & n14542;
  assign n14544 = ~n14489 & ~n14543;
  assign n14545 = ~pi299 & ~n14544;
  assign n14546 = ~pi161 & ~n14398;
  assign n14547 = ~n14465 & n14546;
  assign n14548 = pi146 & n14456;
  assign n14549 = n14393 & ~n14432;
  assign n14550 = n14526 & ~n14549;
  assign n14551 = ~pi146 & ~n14550;
  assign n14552 = ~n14461 & n14551;
  assign n14553 = pi161 & ~n14548;
  assign n14554 = ~n14552 & n14553;
  assign n14555 = ~n14547 & ~n14554;
  assign n14556 = n9344 & ~n14555;
  assign n14557 = pi146 & n14474;
  assign n14558 = ~pi146 & ~n14480;
  assign n14559 = ~pi161 & ~n14558;
  assign n14560 = ~n14557 & n14559;
  assign n14561 = n14526 & n14549;
  assign n14562 = ~n14451 & n14561;
  assign n14563 = ~n14397 & ~n14562;
  assign n14564 = pi146 & ~n14394;
  assign n14565 = ~n14563 & ~n14564;
  assign n14566 = pi161 & ~n14565;
  assign n14567 = ~n14476 & n14566;
  assign n14568 = ~n14560 & ~n14567;
  assign n14569 = n9390 & ~n14568;
  assign n14570 = ~n14556 & ~n14569;
  assign n14571 = pi156 & ~n14570;
  assign n14572 = ~pi146 & ~n14507;
  assign n14573 = pi146 & n14501;
  assign n14574 = n9390 & ~n14572;
  assign n14575 = ~n14573 & n14574;
  assign n14576 = ~pi146 & ~n14518;
  assign n14577 = pi146 & n14522;
  assign n14578 = n9344 & ~n14577;
  assign n14579 = ~n14576 & n14578;
  assign n14580 = ~pi161 & ~n14579;
  assign n14581 = ~n14575 & n14580;
  assign n14582 = ~pi146 & ~n14529;
  assign n14583 = pi146 & ~n14534;
  assign n14584 = ~n14582 & ~n14583;
  assign n14585 = ~n14455 & ~n14584;
  assign n14586 = n14528 & ~n14585;
  assign n14587 = n9344 & ~n14586;
  assign n14588 = n9390 & ~n14398;
  assign n14589 = ~n14460 & n14588;
  assign n14590 = pi161 & ~n14589;
  assign n14591 = ~n14587 & n14590;
  assign n14592 = ~pi156 & ~n14591;
  assign n14593 = ~n14581 & n14592;
  assign n14594 = ~n14571 & ~n14593;
  assign n14595 = ~n14545 & n14594;
  assign n14596 = n9604 & ~n14595;
  assign n14597 = n3094 & n14430;
  assign n14598 = n14394 & ~n14597;
  assign n14599 = ~n6170 & ~n14598;
  assign n14600 = ~n6188 & ~n14599;
  assign n14601 = ~pi142 & ~n14600;
  assign n14602 = n2557 & n7464;
  assign n14603 = ~pi51 & ~n14602;
  assign n14604 = n6170 & ~n14603;
  assign n14605 = ~n14599 & ~n14604;
  assign n14606 = pi142 & ~n14605;
  assign n14607 = n6469 & ~n14601;
  assign n14608 = ~n14606 & n14607;
  assign n14609 = ~n9044 & ~n14608;
  assign n14610 = ~pi287 & n6170;
  assign n14611 = ~pi51 & n14610;
  assign n14612 = ~n14605 & ~n14611;
  assign n14613 = pi224 & ~n14410;
  assign n14614 = n14612 & n14613;
  assign n14615 = ~n14609 & ~n14614;
  assign n14616 = ~n14394 & ~n14410;
  assign n14617 = ~n6469 & ~n14616;
  assign n14618 = pi144 & ~n14617;
  assign n14619 = ~n6469 & n14531;
  assign n14620 = ~n14617 & ~n14619;
  assign n14621 = ~n14618 & n14620;
  assign n14622 = ~n14615 & n14621;
  assign n14623 = ~pi51 & ~n14598;
  assign n14624 = ~pi287 & ~n14623;
  assign n14625 = ~n14531 & ~n14610;
  assign n14626 = ~n14624 & ~n14625;
  assign n14627 = ~n14413 & ~n14626;
  assign n14628 = n9044 & ~n14627;
  assign n14629 = n14393 & n14628;
  assign n14630 = pi51 & ~n6170;
  assign n14631 = ~n14623 & ~n14630;
  assign n14632 = n6469 & ~n14412;
  assign n14633 = n14631 & n14632;
  assign n14634 = n14618 & ~n14633;
  assign n14635 = ~n14629 & n14634;
  assign n14636 = pi181 & ~n14635;
  assign n14637 = ~n14622 & n14636;
  assign n14638 = ~n14608 & n14621;
  assign n14639 = ~pi181 & ~n14634;
  assign n14640 = ~n14638 & n14639;
  assign n14641 = ~pi299 & ~n14640;
  assign n14642 = ~n14637 & n14641;
  assign n14643 = ~n14398 & ~n14598;
  assign n14644 = pi161 & ~n14643;
  assign n14645 = ~pi146 & ~n14600;
  assign n14646 = pi146 & ~n14605;
  assign n14647 = ~pi161 & ~n14645;
  assign n14648 = ~n14646 & n14647;
  assign n14649 = ~n14644 & ~n14648;
  assign n14650 = n6442 & ~n14649;
  assign n14651 = ~n9055 & ~n14650;
  assign n14652 = n14546 & n14612;
  assign n14653 = n14597 & ~n14610;
  assign n14654 = n14394 & ~n14653;
  assign n14655 = n14399 & ~n14654;
  assign n14656 = ~n14652 & ~n14655;
  assign n14657 = pi216 & ~n14656;
  assign n14658 = ~n14651 & ~n14657;
  assign n14659 = ~n14394 & ~n14403;
  assign n14660 = ~n6442 & ~n14659;
  assign n14661 = n9835 & ~n14660;
  assign n14662 = ~n14658 & n14661;
  assign n14663 = n9791 & ~n14660;
  assign n14664 = ~n14650 & n14663;
  assign n14665 = pi232 & ~n14664;
  assign n14666 = ~n14642 & n14665;
  assign n14667 = ~n14662 & n14666;
  assign n14668 = ~n6595 & ~n7535;
  assign n14669 = n14597 & ~n14668;
  assign n14670 = ~pi232 & n14394;
  assign n14671 = ~n14669 & n14670;
  assign n14672 = pi39 & ~n14671;
  assign n14673 = ~n14667 & n14672;
  assign n14674 = ~pi39 & ~pi232;
  assign n14675 = ~n14460 & n14674;
  assign n14676 = ~n14673 & ~n14675;
  assign n14677 = ~n14596 & n14676;
  assign n14678 = ~pi38 & ~n14677;
  assign n14679 = ~n14423 & ~n14678;
  assign n14680 = pi100 & n14394;
  assign n14681 = n3279 & ~n14680;
  assign n14682 = pi100 & n14418;
  assign n14683 = n14681 & ~n14682;
  assign n14684 = ~n14679 & n14683;
  assign n14685 = ~pi87 & ~n3267;
  assign n14686 = ~n14394 & n14685;
  assign n14687 = ~n14418 & n14686;
  assign n14688 = ~pi184 & ~pi299;
  assign n14689 = ~pi163 & pi299;
  assign n14690 = ~n14688 & ~n14689;
  assign n14691 = n7484 & n14690;
  assign n14692 = pi87 & ~n14691;
  assign n14693 = ~n14392 & ~n14692;
  assign n14694 = ~n14687 & n14693;
  assign n14695 = ~n14684 & n14694;
  assign n14696 = n6170 & ~n14498;
  assign n14697 = ~n14401 & n14696;
  assign n14698 = pi161 & ~n14697;
  assign n14699 = n6170 & ~n14453;
  assign n14700 = ~pi146 & n14699;
  assign n14701 = n14393 & ~n14450;
  assign n14702 = n14427 & n14701;
  assign n14703 = n14442 & n14702;
  assign n14704 = ~n14444 & ~n14703;
  assign n14705 = n3094 & ~n14704;
  assign n14706 = ~n14532 & ~n14705;
  assign n14707 = pi146 & n14706;
  assign n14708 = ~pi161 & ~n14700;
  assign n14709 = ~n14707 & n14708;
  assign n14710 = ~n14698 & ~n14709;
  assign n14711 = n9344 & ~n14710;
  assign n14712 = n14399 & ~n14520;
  assign n14713 = ~pi161 & ~n14584;
  assign n14714 = ~n14712 & ~n14713;
  assign n14715 = n9390 & ~n14714;
  assign n14716 = pi232 & ~n14715;
  assign n14717 = ~n14711 & n14716;
  assign n14718 = pi156 & ~n14717;
  assign n14719 = ~n14412 & n14696;
  assign n14720 = pi144 & ~n14719;
  assign n14721 = ~pi142 & n14699;
  assign n14722 = pi142 & n14706;
  assign n14723 = ~pi144 & ~n14721;
  assign n14724 = ~n14722 & n14723;
  assign n14725 = pi180 & ~n14724;
  assign n14726 = ~n14720 & n14725;
  assign n14727 = n14411 & ~n14520;
  assign n14728 = ~pi144 & ~n14536;
  assign n14729 = ~pi180 & ~n14728;
  assign n14730 = ~n14727 & n14729;
  assign n14731 = pi179 & ~n14730;
  assign n14732 = ~n14726 & n14731;
  assign n14733 = n14411 & ~n14473;
  assign n14734 = ~pi51 & ~n14701;
  assign n14735 = n3094 & ~n14734;
  assign n14736 = ~n14532 & ~n14735;
  assign n14737 = pi142 & n14736;
  assign n14738 = n6170 & ~n14452;
  assign n14739 = ~pi142 & n14738;
  assign n14740 = ~pi144 & ~n14739;
  assign n14741 = ~n14737 & n14740;
  assign n14742 = pi180 & ~n14741;
  assign n14743 = ~n14733 & n14742;
  assign n14744 = ~pi180 & n14414;
  assign n14745 = ~pi179 & ~n14744;
  assign n14746 = ~n14743 & n14745;
  assign n14747 = ~n14732 & ~n14746;
  assign n14748 = ~pi299 & ~n14747;
  assign n14749 = ~pi39 & ~n14718;
  assign n14750 = ~n14748 & n14749;
  assign n14751 = pi142 & ~n3096;
  assign n14752 = ~pi142 & ~n14602;
  assign n14753 = n9044 & n14610;
  assign n14754 = ~n14751 & n14753;
  assign n14755 = ~n14752 & n14754;
  assign n14756 = n14411 & ~n14755;
  assign n14757 = ~pi144 & ~n14413;
  assign n14758 = ~n14628 & n14757;
  assign n14759 = pi181 & ~n14758;
  assign n14760 = ~n14756 & n14759;
  assign n14761 = ~pi181 & n14414;
  assign n14762 = ~pi299 & ~n14761;
  assign n14763 = ~n14760 & n14762;
  assign n14764 = n6170 & n6443;
  assign n14765 = n14399 & ~n14764;
  assign n14766 = n14546 & ~n14626;
  assign n14767 = n9055 & ~n14766;
  assign n14768 = ~n14765 & n14767;
  assign n14769 = ~n9055 & n14403;
  assign n14770 = n9835 & ~n14769;
  assign n14771 = ~n14768 & n14770;
  assign n14772 = ~pi159 & n14416;
  assign n14773 = n10457 & ~n14772;
  assign n14774 = ~n14771 & n14773;
  assign n14775 = ~n14763 & n14774;
  assign n14776 = ~pi38 & ~n14775;
  assign n14777 = ~n14750 & n14776;
  assign n14778 = n14399 & ~n14473;
  assign n14779 = pi146 & n14736;
  assign n14780 = ~pi146 & n14738;
  assign n14781 = ~pi161 & ~n14780;
  assign n14782 = ~n14779 & n14781;
  assign n14783 = ~n14778 & ~n14782;
  assign n14784 = n9344 & ~n14783;
  assign n14785 = ~pi158 & n14416;
  assign n14786 = pi232 & ~n14785;
  assign n14787 = ~n14784 & n14786;
  assign n14788 = ~pi156 & n3182;
  assign n14789 = ~n14787 & n14788;
  assign n14790 = n14420 & ~n14789;
  assign n14791 = ~n14777 & n14790;
  assign n14792 = n3279 & ~n14682;
  assign n14793 = ~n14791 & n14792;
  assign n14794 = ~n14418 & n14685;
  assign n14795 = n14392 & ~n14692;
  assign n14796 = ~n14794 & n14795;
  assign n14797 = ~n14793 & n14796;
  assign n14798 = ~po1038 & ~n14797;
  assign n14799 = ~n14695 & n14798;
  assign po279 = n14409 | n14799;
  assign n14801 = n8044 & n8804;
  assign n14802 = n7444 & n14362;
  assign n14803 = n13988 & ~n14802;
  assign n14804 = n7444 & n14371;
  assign n14805 = n7720 & ~n14804;
  assign n14806 = ~po1038 & ~n14803;
  assign n14807 = ~n14805 & n14806;
  assign po280 = n14801 | n14807;
  assign n14809 = ~pi110 & n9039;
  assign n14810 = ~n6229 & n6442;
  assign n14811 = n14809 & n14810;
  assign n14812 = pi39 & ~n14811;
  assign n14813 = pi110 & n10055;
  assign n14814 = ~n10953 & n14813;
  assign n14815 = po1057 & n14814;
  assign n14816 = ~pi39 & ~n14815;
  assign n14817 = po1038 & ~n14816;
  assign n14818 = ~n14812 & n14817;
  assign n14819 = ~pi38 & n3268;
  assign n14820 = pi299 & n14811;
  assign n14821 = ~n6208 & n7535;
  assign n14822 = n14809 & n14821;
  assign n14823 = pi39 & ~n14822;
  assign n14824 = ~n14820 & n14823;
  assign n14825 = ~pi111 & ~n6318;
  assign n14826 = ~pi36 & n2637;
  assign n14827 = ~n14825 & n14826;
  assign n14828 = n2457 & ~n14827;
  assign n14829 = ~n2602 & ~n2646;
  assign n14830 = ~n14828 & n14829;
  assign n14831 = ~pi83 & ~n14830;
  assign n14832 = n2604 & ~n14831;
  assign n14833 = ~pi71 & ~n14832;
  assign n14834 = n6328 & ~n14833;
  assign n14835 = ~pi81 & ~n14834;
  assign n14836 = n11412 & ~n14835;
  assign n14837 = ~pi90 & ~n14836;
  assign n14838 = n2496 & ~n14837;
  assign n14839 = pi90 & ~n10386;
  assign n14840 = n9559 & ~n14839;
  assign n14841 = n14838 & n14840;
  assign n14842 = pi72 & n2497;
  assign n14843 = n10386 & n14842;
  assign n14844 = ~n14841 & ~n14843;
  assign n14845 = n6371 & ~n14844;
  assign n14846 = ~pi110 & ~n14845;
  assign n14847 = n13412 & ~n14846;
  assign n14848 = n2707 & n14838;
  assign n14849 = ~pi72 & ~n14848;
  assign n14850 = n6372 & ~n13412;
  assign n14851 = ~n14849 & n14850;
  assign n14852 = ~pi39 & ~n14851;
  assign n14853 = ~n14847 & n14852;
  assign n14854 = ~n14824 & ~n14853;
  assign n14855 = n14819 & ~n14854;
  assign n14856 = pi110 & n13412;
  assign n14857 = ~pi39 & ~n14856;
  assign n14858 = ~n14824 & ~n14857;
  assign n14859 = ~n14819 & ~n14858;
  assign n14860 = ~po1038 & ~n14859;
  assign n14861 = ~n14855 & n14860;
  assign po281 = ~n14818 & ~n14861;
  assign n14863 = ~pi125 & n14387;
  assign n14864 = pi125 & pi133;
  assign n14865 = ~n14388 & ~n14864;
  assign n14866 = ~n14863 & ~n14865;
  assign n14867 = n14394 & ~n14866;
  assign n14868 = pi172 & n14397;
  assign n14869 = ~pi152 & n14531;
  assign n14870 = ~n14868 & ~n14869;
  assign n14871 = pi232 & ~n14870;
  assign n14872 = ~n14867 & ~n14871;
  assign n14873 = ~pi87 & ~n14872;
  assign n14874 = pi87 & n7484;
  assign n14875 = pi162 & n14874;
  assign n14876 = po1038 & ~n14875;
  assign n14877 = ~n14873 & n14876;
  assign n14878 = ~pi152 & n6170;
  assign n14879 = n14462 & ~n14878;
  assign n14880 = ~pi152 & n14550;
  assign n14881 = ~pi197 & ~n14880;
  assign n14882 = ~n14879 & n14881;
  assign n14883 = ~n6170 & n14462;
  assign n14884 = ~n14526 & ~n14883;
  assign n14885 = ~n14562 & ~n14884;
  assign n14886 = ~pi152 & pi197;
  assign n14887 = ~n14885 & n14886;
  assign n14888 = ~n14882 & ~n14887;
  assign n14889 = ~n14868 & ~n14888;
  assign n14890 = ~n6170 & ~n14462;
  assign n14891 = ~n14479 & ~n14890;
  assign n14892 = ~pi172 & n14891;
  assign n14893 = ~n14397 & ~n14473;
  assign n14894 = ~n14462 & n14893;
  assign n14895 = pi172 & ~n14894;
  assign n14896 = pi152 & pi197;
  assign n14897 = ~n14895 & n14896;
  assign n14898 = ~n14892 & n14897;
  assign n14899 = ~n14889 & ~n14898;
  assign n14900 = n9860 & ~n14899;
  assign n14901 = ~n14506 & ~n14890;
  assign n14902 = ~pi172 & n14901;
  assign n14903 = ~n14499 & ~n14890;
  assign n14904 = pi172 & n14903;
  assign n14905 = pi152 & ~n14904;
  assign n14906 = ~n14902 & n14905;
  assign n14907 = n6170 & n14460;
  assign n14908 = ~n14884 & ~n14907;
  assign n14909 = ~pi152 & ~n14868;
  assign n14910 = ~n14908 & n14909;
  assign n14911 = pi197 & ~n14910;
  assign n14912 = ~n14906 & n14911;
  assign n14913 = ~n14517 & ~n14890;
  assign n14914 = pi152 & n14913;
  assign n14915 = ~n14527 & ~n14883;
  assign n14916 = ~pi152 & ~n14915;
  assign n14917 = ~pi172 & ~n14916;
  assign n14918 = ~n14914 & n14917;
  assign n14919 = n14463 & ~n14520;
  assign n14920 = pi152 & ~n14919;
  assign n14921 = n14459 & n14561;
  assign n14922 = ~n14890 & ~n14921;
  assign n14923 = ~pi152 & n14922;
  assign n14924 = pi172 & ~n14923;
  assign n14925 = ~n14920 & n14924;
  assign n14926 = ~pi197 & ~n14925;
  assign n14927 = ~n14918 & n14926;
  assign n14928 = n9866 & ~n14927;
  assign n14929 = ~n14912 & n14928;
  assign n14930 = ~n14900 & ~n14929;
  assign n14931 = pi299 & ~n14930;
  assign n14932 = pi145 & n14891;
  assign n14933 = ~pi145 & n14462;
  assign n14934 = pi174 & ~n14933;
  assign n14935 = ~n14932 & n14934;
  assign n14936 = pi145 & n14885;
  assign n14937 = ~n14550 & ~n14883;
  assign n14938 = ~pi145 & ~n14937;
  assign n14939 = ~pi174 & ~n14938;
  assign n14940 = ~n14936 & n14939;
  assign n14941 = ~n14935 & ~n14940;
  assign n14942 = ~pi193 & ~n14941;
  assign n14943 = ~pi145 & n14473;
  assign n14944 = ~n14893 & ~n14943;
  assign n14945 = ~n14462 & ~n14944;
  assign n14946 = pi174 & ~n14945;
  assign n14947 = ~n14397 & ~n14451;
  assign n14948 = pi145 & ~n14947;
  assign n14949 = n14561 & ~n14948;
  assign n14950 = ~pi174 & ~n14949;
  assign n14951 = ~n14890 & n14950;
  assign n14952 = pi193 & ~n14951;
  assign n14953 = ~n14946 & n14952;
  assign n14954 = ~n14942 & ~n14953;
  assign n14955 = n9844 & ~n14954;
  assign n14956 = pi145 & n14901;
  assign n14957 = ~pi145 & n14913;
  assign n14958 = ~pi193 & ~n14957;
  assign n14959 = ~n14956 & n14958;
  assign n14960 = pi145 & n14903;
  assign n14961 = ~pi145 & ~n14919;
  assign n14962 = pi193 & ~n14961;
  assign n14963 = ~n14960 & n14962;
  assign n14964 = pi174 & ~n14963;
  assign n14965 = ~n14959 & n14964;
  assign n14966 = pi193 & n14922;
  assign n14967 = ~pi193 & ~n14915;
  assign n14968 = ~pi145 & ~n14966;
  assign n14969 = ~n14967 & n14968;
  assign n14970 = pi193 & n14397;
  assign n14971 = pi145 & ~n14970;
  assign n14972 = ~n14908 & n14971;
  assign n14973 = ~pi174 & ~n14972;
  assign n14974 = ~n14969 & n14973;
  assign n14975 = n9850 & ~n14974;
  assign n14976 = ~n14965 & n14975;
  assign n14977 = ~n14955 & ~n14976;
  assign n14978 = ~pi38 & ~n14977;
  assign n14979 = ~n14931 & ~n14978;
  assign n14980 = n9604 & ~n14979;
  assign n14981 = ~n7532 & ~n7536;
  assign n14982 = n3096 & ~n14981;
  assign n14983 = ~pi232 & ~n14982;
  assign n14984 = pi39 & ~n14983;
  assign n14985 = ~n8074 & n14870;
  assign n14986 = n3096 & ~n6170;
  assign n14987 = n6170 & ~n14598;
  assign n14988 = ~n14986 & ~n14987;
  assign n14989 = ~pi152 & ~n14988;
  assign n14990 = ~n14604 & ~n14986;
  assign n14991 = pi152 & ~n14990;
  assign n14992 = ~n14989 & ~n14991;
  assign n14993 = pi51 & ~pi172;
  assign n14994 = ~n14992 & ~n14993;
  assign n14995 = ~pi216 & ~n14994;
  assign n14996 = n6442 & n14995;
  assign n14997 = ~n14985 & ~n14996;
  assign n14998 = n9390 & ~n14997;
  assign n14999 = n14602 & n14610;
  assign n15000 = ~n14397 & ~n14999;
  assign n15001 = pi224 & n15000;
  assign n15002 = n6469 & ~n15001;
  assign n15003 = n8066 & n14990;
  assign n15004 = n15002 & ~n15003;
  assign n15005 = ~n14397 & ~n15004;
  assign n15006 = pi174 & ~n15005;
  assign n15007 = n8066 & n14988;
  assign n15008 = n14597 & n14610;
  assign n15009 = pi224 & ~n15008;
  assign n15010 = n6469 & ~n15009;
  assign n15011 = ~n14400 & ~n15010;
  assign n15012 = ~n15007 & ~n15011;
  assign n15013 = ~pi174 & n15012;
  assign n15014 = pi193 & ~n15013;
  assign n15015 = ~n15006 & n15014;
  assign n15016 = n6170 & n14623;
  assign n15017 = ~n14986 & ~n15016;
  assign n15018 = ~pi224 & n15017;
  assign n15019 = pi224 & ~n14626;
  assign n15020 = n6469 & ~n15019;
  assign n15021 = ~n15018 & n15020;
  assign n15022 = ~n14619 & ~n15021;
  assign n15023 = ~pi174 & ~n15022;
  assign n15024 = ~n8066 & ~n14753;
  assign n15025 = n3096 & ~n15024;
  assign n15026 = pi174 & n15025;
  assign n15027 = ~pi193 & ~n15026;
  assign n15028 = ~n15023 & n15027;
  assign n15029 = pi180 & ~n15028;
  assign n15030 = ~n15015 & n15029;
  assign n15031 = ~n8066 & ~n14400;
  assign n15032 = ~n15017 & ~n15031;
  assign n15033 = ~pi174 & n15032;
  assign n15034 = n3096 & n8066;
  assign n15035 = pi174 & n15034;
  assign n15036 = ~n14970 & ~n15035;
  assign n15037 = ~n15033 & n15036;
  assign n15038 = ~pi180 & ~n15037;
  assign n15039 = ~pi299 & ~n15038;
  assign n15040 = ~n15030 & n15039;
  assign n15041 = pi152 & n15000;
  assign n15042 = ~n14400 & ~n15008;
  assign n15043 = ~pi152 & n15042;
  assign n15044 = pi172 & ~n15043;
  assign n15045 = ~n15041 & n15044;
  assign n15046 = pi152 & ~n14764;
  assign n15047 = ~pi152 & ~n14626;
  assign n15048 = ~pi172 & ~n15047;
  assign n15049 = ~n15046 & n15048;
  assign n15050 = pi216 & ~n15045;
  assign n15051 = ~n15049 & n15050;
  assign n15052 = n6442 & ~n15051;
  assign n15053 = ~n14995 & n15052;
  assign n15054 = ~n6442 & ~n14870;
  assign n15055 = n9344 & ~n15054;
  assign n15056 = ~n15053 & n15055;
  assign n15057 = ~n14998 & ~n15056;
  assign n15058 = ~n15040 & n15057;
  assign n15059 = pi232 & ~n15058;
  assign n15060 = n14984 & ~n15059;
  assign n15061 = ~pi232 & ~n14462;
  assign n15062 = ~pi39 & ~n15061;
  assign n15063 = ~pi38 & ~n15062;
  assign n15064 = ~n15060 & n15063;
  assign n15065 = pi299 & n14870;
  assign n15066 = ~pi174 & n14531;
  assign n15067 = ~pi299 & ~n14970;
  assign n15068 = ~n15066 & n15067;
  assign n15069 = pi232 & ~n15068;
  assign n15070 = ~n15065 & n15069;
  assign n15071 = pi38 & ~n15070;
  assign n15072 = ~pi100 & ~n15071;
  assign n15073 = ~n15064 & n15072;
  assign n15074 = ~n14980 & n15073;
  assign n15075 = pi100 & n15070;
  assign n15076 = n3279 & ~n15075;
  assign n15077 = ~n15074 & n15076;
  assign n15078 = n14685 & ~n15070;
  assign n15079 = pi140 & ~pi299;
  assign n15080 = pi162 & pi299;
  assign n15081 = ~n15079 & ~n15080;
  assign n15082 = n7484 & ~n15081;
  assign n15083 = pi87 & ~n15082;
  assign n15084 = n14866 & ~n15083;
  assign n15085 = ~n15078 & n15084;
  assign n15086 = ~n15077 & n15085;
  assign n15087 = n14472 & n14503;
  assign n15088 = ~n14454 & ~n15087;
  assign n15089 = ~pi145 & n15088;
  assign n15090 = ~n14454 & ~n14520;
  assign n15091 = pi145 & n15090;
  assign n15092 = ~pi174 & ~n15091;
  assign n15093 = ~n15089 & n15092;
  assign n15094 = ~n14454 & ~n14706;
  assign n15095 = ~pi145 & ~n14452;
  assign n15096 = ~n6170 & ~n14452;
  assign n15097 = ~n14400 & ~n15096;
  assign n15098 = ~n14446 & n15097;
  assign n15099 = ~n15095 & n15098;
  assign n15100 = n3094 & n15099;
  assign n15101 = pi174 & ~n15094;
  assign n15102 = ~n15100 & n15101;
  assign n15103 = pi193 & ~n15102;
  assign n15104 = ~n15093 & n15103;
  assign n15105 = ~pi145 & ~n14454;
  assign n15106 = ~n14696 & n15105;
  assign n15107 = ~pi51 & n15091;
  assign n15108 = ~pi174 & ~n15107;
  assign n15109 = ~n15106 & n15108;
  assign n15110 = pi174 & ~n15099;
  assign n15111 = ~pi193 & ~n15110;
  assign n15112 = ~n15109 & n15111;
  assign n15113 = n9844 & ~n15104;
  assign n15114 = ~n15112 & n15113;
  assign n15115 = ~n14397 & ~n14454;
  assign n15116 = ~pi174 & ~n14943;
  assign n15117 = pi145 & n14393;
  assign n15118 = ~n15116 & ~n15117;
  assign n15119 = n15115 & ~n15118;
  assign n15120 = ~n14454 & ~n14738;
  assign n15121 = pi174 & n15120;
  assign n15122 = ~n15119 & ~n15121;
  assign n15123 = ~pi193 & ~n15122;
  assign n15124 = pi145 & ~n14531;
  assign n15125 = ~pi145 & pi174;
  assign n15126 = ~n14736 & n15125;
  assign n15127 = ~n15124 & ~n15126;
  assign n15128 = ~n15116 & n15127;
  assign n15129 = pi193 & ~n14454;
  assign n15130 = ~n15128 & n15129;
  assign n15131 = n9850 & ~n15130;
  assign n15132 = ~n15123 & n15131;
  assign n15133 = ~n15114 & ~n15132;
  assign n15134 = ~pi38 & ~n15133;
  assign n15135 = ~pi152 & ~n15088;
  assign n15136 = pi152 & ~n15094;
  assign n15137 = pi172 & ~n15136;
  assign n15138 = ~n15135 & n15137;
  assign n15139 = ~pi152 & n14696;
  assign n15140 = ~n14453 & ~n14878;
  assign n15141 = ~pi172 & ~n15140;
  assign n15142 = ~n15139 & n15141;
  assign n15143 = ~n15138 & ~n15142;
  assign n15144 = ~pi197 & ~n15143;
  assign n15145 = ~pi152 & ~n15090;
  assign n15146 = ~n14454 & ~n14534;
  assign n15147 = pi172 & n15146;
  assign n15148 = ~pi172 & n15098;
  assign n15149 = pi152 & ~n15148;
  assign n15150 = ~n15147 & n15149;
  assign n15151 = ~pi172 & n14397;
  assign n15152 = pi197 & ~n15151;
  assign n15153 = ~n15150 & n15152;
  assign n15154 = ~n15145 & n15153;
  assign n15155 = pi299 & n9860;
  assign n15156 = ~n15154 & n15155;
  assign n15157 = ~n15144 & n15156;
  assign n15158 = ~n14454 & ~n14473;
  assign n15159 = ~pi152 & n15158;
  assign n15160 = ~n14397 & n15159;
  assign n15161 = pi152 & n15120;
  assign n15162 = ~pi172 & ~n15161;
  assign n15163 = ~n15160 & n15162;
  assign n15164 = ~n14454 & ~n14736;
  assign n15165 = pi152 & n15164;
  assign n15166 = pi172 & ~n15165;
  assign n15167 = ~n15159 & n15166;
  assign n15168 = ~pi197 & ~n15167;
  assign n15169 = ~n15163 & n15168;
  assign n15170 = pi152 & n14531;
  assign n15171 = ~n14454 & ~n15170;
  assign n15172 = pi172 & ~n15171;
  assign n15173 = ~pi172 & ~n14869;
  assign n15174 = ~n14455 & n15173;
  assign n15175 = pi197 & ~n15172;
  assign n15176 = ~n15174 & n15175;
  assign n15177 = pi299 & n9866;
  assign n15178 = ~n15176 & n15177;
  assign n15179 = ~n15169 & n15178;
  assign n15180 = ~n15157 & ~n15179;
  assign n15181 = ~n15134 & n15180;
  assign n15182 = n9604 & ~n15181;
  assign n15183 = ~n14422 & ~n15072;
  assign n15184 = ~n14394 & n14870;
  assign n15185 = ~n9055 & ~n15184;
  assign n15186 = ~n14598 & ~n14878;
  assign n15187 = ~pi152 & n14604;
  assign n15188 = ~n15186 & ~n15187;
  assign n15189 = ~pi172 & ~n15188;
  assign n15190 = ~pi152 & n14600;
  assign n15191 = pi152 & n14631;
  assign n15192 = pi172 & ~n15191;
  assign n15193 = ~n15190 & n15192;
  assign n15194 = n9055 & ~n15189;
  assign n15195 = ~n15193 & n15194;
  assign n15196 = n9390 & ~n15195;
  assign n15197 = n14612 & n14909;
  assign n15198 = pi152 & ~n14868;
  assign n15199 = ~n14654 & n15198;
  assign n15200 = n9055 & ~n15199;
  assign n15201 = ~n15197 & n15200;
  assign n15202 = n9344 & ~n15201;
  assign n15203 = ~n15196 & ~n15202;
  assign n15204 = ~n15185 & ~n15203;
  assign n15205 = ~n6170 & ~n14393;
  assign n15206 = ~n9044 & ~n15205;
  assign n15207 = ~n14630 & n15206;
  assign n15208 = n9044 & n14600;
  assign n15209 = ~n15207 & ~n15208;
  assign n15210 = ~pi174 & ~n15209;
  assign n15211 = n9044 & n14597;
  assign n15212 = n14394 & ~n15211;
  assign n15213 = ~n14397 & ~n15212;
  assign n15214 = pi174 & ~n15213;
  assign n15215 = ~pi180 & ~n15214;
  assign n15216 = ~n15210 & n15215;
  assign n15217 = n9044 & ~n14599;
  assign n15218 = ~n10522 & n15217;
  assign n15219 = ~n15207 & ~n15218;
  assign n15220 = ~pi174 & ~n15219;
  assign n15221 = ~pi51 & ~n14654;
  assign n15222 = n6170 & ~n15221;
  assign n15223 = ~n15212 & ~n15222;
  assign n15224 = pi174 & ~n15223;
  assign n15225 = pi180 & ~n15224;
  assign n15226 = ~n15220 & n15225;
  assign n15227 = pi193 & ~n15226;
  assign n15228 = ~n15216 & n15227;
  assign n15229 = n9044 & n14605;
  assign n15230 = ~pi51 & n15206;
  assign n15231 = ~n15229 & ~n15230;
  assign n15232 = pi180 & n14611;
  assign n15233 = ~pi174 & ~n15232;
  assign n15234 = n15231 & n15233;
  assign n15235 = pi180 & n14654;
  assign n15236 = pi174 & ~n15212;
  assign n15237 = ~n15235 & n15236;
  assign n15238 = ~pi193 & ~n15237;
  assign n15239 = ~n15234 & n15238;
  assign n15240 = ~pi299 & ~n15239;
  assign n15241 = ~n15228 & n15240;
  assign n15242 = ~n15204 & ~n15241;
  assign n15243 = pi232 & ~n15242;
  assign n15244 = ~pi299 & ~n15212;
  assign n15245 = n9055 & n14597;
  assign n15246 = n14394 & ~n15245;
  assign n15247 = pi299 & ~n15246;
  assign n15248 = ~n15244 & ~n15247;
  assign n15249 = ~pi232 & ~n15248;
  assign n15250 = pi39 & ~n15249;
  assign n15251 = ~n15243 & n15250;
  assign n15252 = ~pi232 & ~n14453;
  assign n15253 = ~pi39 & ~n15252;
  assign n15254 = ~pi38 & ~n15253;
  assign n15255 = ~n15251 & n15254;
  assign n15256 = ~n15183 & ~n15255;
  assign n15257 = ~n15182 & n15256;
  assign n15258 = n14681 & ~n15075;
  assign n15259 = ~n15257 & n15258;
  assign n15260 = n14686 & ~n15070;
  assign n15261 = ~n14866 & ~n15083;
  assign n15262 = ~n15260 & n15261;
  assign n15263 = ~n15259 & n15262;
  assign n15264 = ~po1038 & ~n15263;
  assign n15265 = ~n15086 & n15264;
  assign po282 = n14877 | n15265;
  assign n15267 = ~pi153 & n14901;
  assign n15268 = pi153 & n14903;
  assign n15269 = pi157 & ~n15268;
  assign n15270 = ~n15267 & n15269;
  assign n15271 = ~pi153 & n14891;
  assign n15272 = pi153 & ~n14894;
  assign n15273 = ~pi157 & ~n15272;
  assign n15274 = ~n15271 & n15273;
  assign n15275 = ~n15270 & ~n15274;
  assign n15276 = pi166 & ~n15275;
  assign n15277 = pi157 & n14908;
  assign n15278 = ~pi157 & n14885;
  assign n15279 = pi153 & n14397;
  assign n15280 = ~pi166 & ~n15279;
  assign n15281 = ~n15277 & n15280;
  assign n15282 = ~n15278 & n15281;
  assign n15283 = ~n15276 & ~n15282;
  assign n15284 = n9835 & ~n15283;
  assign n15285 = ~pi189 & n14908;
  assign n15286 = pi189 & n14901;
  assign n15287 = ~n15285 & ~n15286;
  assign n15288 = pi178 & ~n15287;
  assign n15289 = ~pi189 & ~n14885;
  assign n15290 = pi189 & ~n14891;
  assign n15291 = ~pi178 & ~n15289;
  assign n15292 = ~n15290 & n15291;
  assign n15293 = ~n15288 & ~n15292;
  assign n15294 = pi181 & ~n15293;
  assign n15295 = pi189 & n14913;
  assign n15296 = ~pi189 & ~n14915;
  assign n15297 = pi178 & ~n15296;
  assign n15298 = ~n15295 & n15297;
  assign n15299 = ~pi189 & ~n14937;
  assign n15300 = pi189 & n14462;
  assign n15301 = ~pi178 & ~n15300;
  assign n15302 = ~n14397 & n15301;
  assign n15303 = ~n15299 & n15302;
  assign n15304 = ~pi181 & ~n15303;
  assign n15305 = n14937 & n15301;
  assign n15306 = n15304 & ~n15305;
  assign n15307 = ~n15298 & n15306;
  assign n15308 = n11791 & ~n15307;
  assign n15309 = ~n15294 & n15308;
  assign n15310 = pi166 & ~n14919;
  assign n15311 = ~pi166 & n14922;
  assign n15312 = pi153 & ~n15311;
  assign n15313 = ~n15310 & n15312;
  assign n15314 = pi166 & n14913;
  assign n15315 = ~pi166 & ~n14915;
  assign n15316 = ~pi153 & ~n15315;
  assign n15317 = ~n15314 & n15316;
  assign n15318 = ~n15313 & ~n15317;
  assign n15319 = pi157 & ~n15318;
  assign n15320 = ~pi166 & ~n14937;
  assign n15321 = pi166 & n14462;
  assign n15322 = ~pi157 & ~n15279;
  assign n15323 = ~n15321 & n15322;
  assign n15324 = ~n15320 & n15323;
  assign n15325 = ~n15319 & ~n15324;
  assign n15326 = n9791 & ~n15325;
  assign n15327 = ~pi189 & n15115;
  assign n15328 = n14903 & ~n15327;
  assign n15329 = pi178 & ~n15285;
  assign n15330 = ~n15328 & n15329;
  assign n15331 = pi189 & n14894;
  assign n15332 = ~n14397 & n15289;
  assign n15333 = ~n15331 & ~n15332;
  assign n15334 = ~pi178 & ~n15333;
  assign n15335 = pi181 & ~n15334;
  assign n15336 = ~n15330 & n15335;
  assign n15337 = pi189 & ~n14919;
  assign n15338 = ~pi189 & n14922;
  assign n15339 = pi178 & ~n15338;
  assign n15340 = ~n15337 & n15339;
  assign n15341 = n15304 & ~n15340;
  assign n15342 = n11830 & ~n15341;
  assign n15343 = ~n15336 & n15342;
  assign n15344 = ~n15326 & ~n15343;
  assign n15345 = ~n15284 & n15344;
  assign n15346 = ~n15309 & n15345;
  assign n15347 = pi232 & ~n15346;
  assign n15348 = n15062 & ~n15347;
  assign n15349 = ~pi126 & n14390;
  assign n15350 = pi126 & ~n14390;
  assign n15351 = ~n15349 & ~n15350;
  assign n15352 = ~n14386 & ~n15351;
  assign n15353 = ~pi189 & n15032;
  assign n15354 = pi189 & n15034;
  assign n15355 = ~pi182 & ~n15354;
  assign n15356 = ~n15353 & n15355;
  assign n15357 = ~n14397 & n15356;
  assign n15358 = pi189 & ~n15005;
  assign n15359 = ~pi189 & n15012;
  assign n15360 = pi182 & ~n15359;
  assign n15361 = ~n15358 & n15360;
  assign n15362 = ~n15357 & ~n15361;
  assign n15363 = n11830 & ~n15362;
  assign n15364 = pi166 & n14764;
  assign n15365 = ~pi166 & n14626;
  assign n15366 = ~pi153 & ~n15365;
  assign n15367 = ~n15364 & n15366;
  assign n15368 = pi166 & ~n15000;
  assign n15369 = ~pi166 & ~n15042;
  assign n15370 = pi153 & ~n15369;
  assign n15371 = ~n15368 & n15370;
  assign n15372 = pi160 & ~n15367;
  assign n15373 = ~n15371 & n15372;
  assign n15374 = pi216 & ~n15373;
  assign n15375 = ~pi166 & ~n14988;
  assign n15376 = pi166 & ~n14990;
  assign n15377 = ~n15375 & ~n15376;
  assign n15378 = pi51 & ~pi153;
  assign n15379 = ~n15377 & ~n15378;
  assign n15380 = ~pi216 & ~n15379;
  assign n15381 = n6442 & ~n15374;
  assign n15382 = ~n15380 & n15381;
  assign n15383 = ~pi51 & ~n14531;
  assign n15384 = ~n10305 & ~n14393;
  assign n15385 = ~pi51 & ~n15384;
  assign n15386 = ~n15279 & ~n15385;
  assign n15387 = ~n15383 & ~n15386;
  assign n15388 = ~pi160 & pi216;
  assign n15389 = n6442 & ~n15388;
  assign n15390 = n15387 & ~n15389;
  assign n15391 = pi299 & ~n15390;
  assign n15392 = ~n15382 & n15391;
  assign n15393 = ~pi189 & ~n15022;
  assign n15394 = pi189 & n15025;
  assign n15395 = pi182 & ~n15394;
  assign n15396 = ~n15393 & n15395;
  assign n15397 = ~n15356 & ~n15396;
  assign n15398 = n11791 & ~n15397;
  assign n15399 = ~n15363 & ~n15398;
  assign n15400 = ~n15392 & n15399;
  assign n15401 = pi232 & ~n15400;
  assign n15402 = n14984 & ~n15401;
  assign n15403 = n15352 & ~n15402;
  assign n15404 = ~n15348 & n15403;
  assign n15405 = ~n10301 & ~n14453;
  assign n15406 = ~pi189 & n14696;
  assign n15407 = ~n15405 & ~n15406;
  assign n15408 = ~pi178 & ~n15407;
  assign n15409 = pi189 & n15120;
  assign n15410 = pi178 & ~n15327;
  assign n15411 = ~pi189 & n15158;
  assign n15412 = pi178 & ~n15411;
  assign n15413 = ~n15410 & ~n15412;
  assign n15414 = ~n15409 & ~n15413;
  assign n15415 = ~pi181 & ~n15414;
  assign n15416 = ~n15408 & n15415;
  assign n15417 = ~n14520 & n15327;
  assign n15418 = pi189 & n15098;
  assign n15419 = ~pi178 & ~n15418;
  assign n15420 = ~n15417 & n15419;
  assign n15421 = ~n14455 & n15410;
  assign n15422 = pi181 & ~n15421;
  assign n15423 = ~n15420 & n15422;
  assign n15424 = n11791 & ~n15423;
  assign n15425 = ~n15416 & n15424;
  assign n15426 = ~pi166 & ~n15088;
  assign n15427 = pi166 & ~n15094;
  assign n15428 = pi153 & ~n15427;
  assign n15429 = ~n15426 & n15428;
  assign n15430 = ~pi166 & n14696;
  assign n15431 = ~n10305 & ~n14453;
  assign n15432 = ~pi153 & ~n15431;
  assign n15433 = ~n15430 & n15432;
  assign n15434 = ~n15429 & ~n15433;
  assign n15435 = ~pi157 & ~n15434;
  assign n15436 = ~pi166 & ~n15158;
  assign n15437 = pi51 & n10305;
  assign n15438 = pi166 & ~n15120;
  assign n15439 = ~n15437 & ~n15438;
  assign n15440 = ~pi153 & ~n15439;
  assign n15441 = pi153 & pi166;
  assign n15442 = ~n15164 & n15441;
  assign n15443 = pi157 & ~n15442;
  assign n15444 = ~n15436 & n15443;
  assign n15445 = ~n15440 & n15444;
  assign n15446 = n9791 & ~n15445;
  assign n15447 = ~n15435 & n15446;
  assign n15448 = ~pi189 & n15088;
  assign n15449 = pi189 & n15094;
  assign n15450 = ~pi178 & ~n15449;
  assign n15451 = ~n15448 & n15450;
  assign n15452 = pi189 & n15164;
  assign n15453 = n15412 & ~n15452;
  assign n15454 = ~pi181 & ~n15453;
  assign n15455 = ~n15451 & n15454;
  assign n15456 = ~pi189 & ~n14520;
  assign n15457 = pi189 & ~n14534;
  assign n15458 = ~pi178 & ~n15457;
  assign n15459 = ~n15456 & n15458;
  assign n15460 = pi178 & n11800;
  assign n15461 = n14443 & n15460;
  assign n15462 = pi181 & ~n15461;
  assign n15463 = ~n14454 & n15462;
  assign n15464 = ~n15459 & n15463;
  assign n15465 = n11830 & ~n15464;
  assign n15466 = ~n15455 & n15465;
  assign n15467 = ~pi166 & ~n15090;
  assign n15468 = ~n15146 & n15441;
  assign n15469 = pi166 & ~n15098;
  assign n15470 = ~n15437 & ~n15469;
  assign n15471 = ~pi153 & ~n15470;
  assign n15472 = ~pi157 & ~n15468;
  assign n15473 = ~n15471 & n15472;
  assign n15474 = ~n15467 & n15473;
  assign n15475 = pi166 & n14531;
  assign n15476 = ~n14454 & ~n15475;
  assign n15477 = pi153 & ~n15476;
  assign n15478 = ~pi153 & ~n15387;
  assign n15479 = ~n14455 & n15478;
  assign n15480 = pi157 & ~n15477;
  assign n15481 = ~n15479 & n15480;
  assign n15482 = n9835 & ~n15481;
  assign n15483 = ~n15474 & n15482;
  assign n15484 = ~n15466 & ~n15483;
  assign n15485 = ~n15425 & n15484;
  assign n15486 = ~n15447 & n15485;
  assign n15487 = pi232 & ~n15486;
  assign n15488 = n15253 & ~n15487;
  assign n15489 = ~pi166 & n14612;
  assign n15490 = pi166 & ~n14654;
  assign n15491 = ~n15489 & ~n15490;
  assign n15492 = pi160 & ~n15279;
  assign n15493 = ~n15491 & n15492;
  assign n15494 = ~n10305 & ~n14598;
  assign n15495 = ~pi166 & n14604;
  assign n15496 = ~n15494 & ~n15495;
  assign n15497 = ~pi153 & ~n15496;
  assign n15498 = ~pi166 & n14600;
  assign n15499 = pi166 & n14631;
  assign n15500 = pi153 & ~n15499;
  assign n15501 = ~n15498 & n15500;
  assign n15502 = ~n15497 & ~n15501;
  assign n15503 = ~pi160 & ~n15502;
  assign n15504 = n9055 & ~n15493;
  assign n15505 = ~n15503 & n15504;
  assign n15506 = ~n9055 & ~n15386;
  assign n15507 = pi299 & ~n15506;
  assign n15508 = ~n15505 & n15507;
  assign n15509 = pi182 & n14654;
  assign n15510 = pi189 & ~n15212;
  assign n15511 = ~n15509 & n15510;
  assign n15512 = pi182 & n14611;
  assign n15513 = ~pi189 & ~n15512;
  assign n15514 = n15231 & n15513;
  assign n15515 = ~n15511 & ~n15514;
  assign n15516 = n11791 & ~n15515;
  assign n15517 = ~pi189 & ~n15209;
  assign n15518 = pi189 & ~n15213;
  assign n15519 = ~pi182 & ~n15518;
  assign n15520 = ~n15517 & n15519;
  assign n15521 = ~pi189 & ~n15219;
  assign n15522 = pi189 & ~n15223;
  assign n15523 = pi182 & ~n15522;
  assign n15524 = ~n15521 & n15523;
  assign n15525 = ~n15520 & ~n15524;
  assign n15526 = n11830 & ~n15525;
  assign n15527 = ~n15516 & ~n15526;
  assign n15528 = ~n15508 & n15527;
  assign n15529 = pi232 & ~n15528;
  assign n15530 = n15250 & ~n15529;
  assign n15531 = ~n15352 & ~n15530;
  assign n15532 = ~n15488 & n15531;
  assign n15533 = n3207 & ~n15532;
  assign n15534 = ~n15404 & n15533;
  assign n15535 = pi299 & ~n15387;
  assign n15536 = ~pi189 & n14531;
  assign n15537 = pi175 & n14397;
  assign n15538 = ~pi299 & ~n15537;
  assign n15539 = ~n15536 & n15538;
  assign n15540 = pi232 & ~n15539;
  assign n15541 = ~n15535 & n15540;
  assign n15542 = ~n3207 & n15541;
  assign n15543 = ~n3207 & n14394;
  assign n15544 = ~n15352 & n15543;
  assign n15545 = n3279 & ~n15544;
  assign n15546 = ~n15542 & n15545;
  assign n15547 = ~n15534 & n15546;
  assign n15548 = n14685 & ~n15541;
  assign n15549 = ~pi150 & pi299;
  assign n15550 = ~pi185 & ~pi299;
  assign n15551 = ~n15549 & ~n15550;
  assign n15552 = n7484 & n15551;
  assign n15553 = pi87 & ~n15552;
  assign n15554 = ~n15548 & ~n15553;
  assign n15555 = n14395 & ~n15352;
  assign n15556 = ~n15554 & ~n15555;
  assign n15557 = ~po1038 & ~n15556;
  assign n15558 = ~n15547 & n15557;
  assign n15559 = pi232 & ~n15383;
  assign n15560 = n15352 & ~n15559;
  assign n15561 = ~pi232 & ~n14394;
  assign n15562 = ~n15386 & ~n15561;
  assign n15563 = ~n15560 & n15562;
  assign n15564 = ~pi87 & ~n15563;
  assign n15565 = pi87 & ~n13791;
  assign n15566 = po1038 & ~n15565;
  assign n15567 = ~n15564 & n15566;
  assign po283 = ~n15558 & ~n15567;
  assign n15569 = n3281 & n8872;
  assign n15570 = ~n3294 & ~n15569;
  assign n15571 = pi129 & n6117;
  assign n15572 = pi38 & ~n15571;
  assign n15573 = ~n2524 & ~n2898;
  assign n15574 = n2597 & ~n2669;
  assign n15575 = n2451 & ~n15574;
  assign n15576 = n2683 & ~n15575;
  assign n15577 = n2594 & ~n15576;
  assign n15578 = n2687 & ~n15577;
  assign n15579 = n2504 & ~n15578;
  assign n15580 = ~n2507 & ~n15579;
  assign n15581 = ~pi86 & ~n15580;
  assign n15582 = n2592 & ~n15581;
  assign n15583 = ~pi97 & ~n15582;
  assign n15584 = ~n2585 & ~n15583;
  assign n15585 = ~pi108 & ~n15584;
  assign n15586 = n2584 & ~n15585;
  assign n15587 = n2699 & ~n15586;
  assign n15588 = ~n2575 & ~n15587;
  assign n15589 = n2574 & ~n15588;
  assign n15590 = n2573 & ~n15589;
  assign n15591 = po740 & n15590;
  assign n15592 = n2590 & ~n15582;
  assign n15593 = ~n2585 & ~n15592;
  assign n15594 = ~pi108 & ~n15593;
  assign n15595 = n2584 & ~n15594;
  assign n15596 = n2699 & ~n15595;
  assign n15597 = ~n2575 & ~n15596;
  assign n15598 = n2574 & ~n15597;
  assign n15599 = n2573 & ~n15598;
  assign n15600 = ~po740 & n15599;
  assign n15601 = pi250 & ~n7485;
  assign n15602 = n10057 & n15601;
  assign n15603 = ~n15591 & n15602;
  assign n15604 = ~n15600 & n15603;
  assign n15605 = ~pi127 & n15590;
  assign n15606 = pi127 & n15599;
  assign n15607 = ~n15602 & ~n15605;
  assign n15608 = ~n15606 & n15607;
  assign n15609 = ~n15604 & ~n15608;
  assign n15610 = n2566 & ~n15609;
  assign n15611 = n2900 & ~n15610;
  assign n15612 = n2547 & ~n15611;
  assign n15613 = n15573 & ~n15612;
  assign n15614 = ~pi70 & ~n15613;
  assign n15615 = ~n2917 & ~n15614;
  assign n15616 = ~pi51 & ~n15615;
  assign n15617 = n2559 & ~n15616;
  assign n15618 = n2920 & ~n15617;
  assign n15619 = ~n2555 & ~n15618;
  assign n15620 = n2725 & ~n15619;
  assign n15621 = n3364 & ~n15620;
  assign n15622 = ~pi95 & ~n15621;
  assign n15623 = ~pi39 & pi129;
  assign n15624 = ~n2727 & n15623;
  assign n15625 = ~n15622 & n15624;
  assign n15626 = pi39 & n8872;
  assign n15627 = ~pi38 & ~n15626;
  assign n15628 = ~n15625 & n15627;
  assign n15629 = ~n15572 & ~n15628;
  assign n15630 = n3241 & ~n15629;
  assign n15631 = ~n3208 & ~n8951;
  assign n15632 = n8872 & ~n15631;
  assign n15633 = ~n3241 & ~n15632;
  assign n15634 = ~pi75 & ~n15633;
  assign n15635 = ~n15630 & n15634;
  assign n15636 = pi129 & n7291;
  assign n15637 = pi75 & n15636;
  assign n15638 = ~pi92 & ~n15637;
  assign n15639 = ~n15635 & n15638;
  assign n15640 = pi92 & ~pi129;
  assign n15641 = n13616 & ~n15640;
  assign n15642 = ~n15639 & n15641;
  assign n15643 = pi54 & n3239;
  assign n15644 = n8872 & n15643;
  assign n15645 = ~pi74 & ~n15644;
  assign n15646 = ~n15642 & n15645;
  assign n15647 = n6544 & n15636;
  assign n15648 = pi74 & ~n15647;
  assign n15649 = ~pi55 & ~n15648;
  assign n15650 = ~n15646 & n15649;
  assign n15651 = pi55 & n3267;
  assign n15652 = n15636 & n15651;
  assign n15653 = ~n15650 & ~n15652;
  assign n15654 = ~pi56 & ~n15653;
  assign n15655 = ~n11284 & ~n11295;
  assign n15656 = ~n15654 & n15655;
  assign n15657 = ~n15570 & ~n15656;
  assign n15658 = n3432 & ~n15657;
  assign n15659 = n3294 & n15569;
  assign n15660 = ~n3432 & ~n15659;
  assign n15661 = ~n6105 & ~n15660;
  assign po284 = ~n15658 & n15661;
  assign n15663 = ~n6115 & ~n7337;
  assign n15664 = ~pi38 & ~n3369;
  assign n15665 = n6119 & ~n15664;
  assign n15666 = n6252 & ~n6269;
  assign n15667 = ~pi87 & ~n15666;
  assign n15668 = ~n15665 & n15667;
  assign n15669 = n6278 & ~n15668;
  assign n15670 = n8874 & n10390;
  assign n15671 = po740 & n15670;
  assign n15672 = ~pi129 & ~n15670;
  assign n15673 = n8953 & ~n15671;
  assign n15674 = ~n15672 & n15673;
  assign n15675 = n3096 & n15674;
  assign n15676 = n6279 & ~n15675;
  assign n15677 = ~n15669 & n15676;
  assign n15678 = ~n7295 & ~n7331;
  assign n15679 = ~n15677 & n15678;
  assign n15680 = n8865 & ~n15679;
  assign n15681 = n15663 & ~n15680;
  assign n15682 = ~pi56 & ~n15681;
  assign n15683 = ~n6112 & ~n15682;
  assign n15684 = ~pi62 & ~n15683;
  assign n15685 = ~n6288 & ~n15684;
  assign n15686 = n3432 & ~n15685;
  assign po286 = n6108 & ~n15686;
  assign n15688 = ~pi51 & ~n15248;
  assign n15689 = ~pi232 & ~n15688;
  assign n15690 = n10959 & ~n15689;
  assign n15691 = ~pi51 & n15231;
  assign n15692 = pi140 & n14610;
  assign n15693 = n15691 & ~n15692;
  assign n15694 = n8996 & ~n15693;
  assign n15695 = ~pi51 & ~n14605;
  assign n15696 = ~n14610 & n15695;
  assign n15697 = pi169 & ~n15696;
  assign n15698 = pi162 & n9055;
  assign n15699 = ~pi169 & ~n15221;
  assign n15700 = n15698 & ~n15699;
  assign n15701 = ~n15697 & n15700;
  assign n15702 = pi169 & n6170;
  assign n15703 = ~n3096 & n15702;
  assign n15704 = ~n14623 & ~n15702;
  assign n15705 = ~pi162 & n9055;
  assign n15706 = ~n15704 & n15705;
  assign n15707 = ~n15703 & n15706;
  assign n15708 = ~n9055 & n14443;
  assign n15709 = ~n15702 & n15708;
  assign n15710 = pi299 & ~n15709;
  assign n15711 = ~n15707 & n15710;
  assign n15712 = ~n15701 & n15711;
  assign n15713 = ~pi191 & ~pi299;
  assign n15714 = ~pi51 & ~n15212;
  assign n15715 = pi140 & n15222;
  assign n15716 = n15714 & ~n15715;
  assign n15717 = n15713 & ~n15716;
  assign n15718 = ~n15694 & ~n15717;
  assign n15719 = ~n15712 & n15718;
  assign n15720 = pi232 & ~n15719;
  assign n15721 = n15690 & ~n15720;
  assign n15722 = n7484 & ~n8998;
  assign n15723 = n14443 & ~n15722;
  assign n15724 = ~n10959 & n15723;
  assign n15725 = ~pi100 & ~n15724;
  assign n15726 = ~n15721 & n15725;
  assign n15727 = ~n15383 & ~n15723;
  assign n15728 = pi100 & n15727;
  assign n15729 = n3279 & ~n15728;
  assign n15730 = ~n14680 & n15729;
  assign n15731 = ~n15726 & n15730;
  assign n15732 = pi87 & ~n9735;
  assign n15733 = n14685 & ~n15727;
  assign n15734 = ~n15732 & ~n15733;
  assign n15735 = ~n14395 & ~n15734;
  assign n15736 = ~pi132 & n15349;
  assign n15737 = pi130 & ~n15736;
  assign n15738 = ~pi130 & n15736;
  assign n15739 = ~n15737 & ~n15738;
  assign n15740 = ~n14384 & ~n15739;
  assign n15741 = ~n15735 & ~n15740;
  assign n15742 = ~n15731 & n15741;
  assign n15743 = ~n14630 & n15042;
  assign n15744 = pi224 & ~n15743;
  assign n15745 = ~n6170 & ~n14603;
  assign n15746 = ~n14987 & ~n15745;
  assign n15747 = ~pi224 & ~n15746;
  assign n15748 = ~n15744 & ~n15747;
  assign n15749 = n6469 & ~n15748;
  assign n15750 = ~n6469 & ~n15383;
  assign n15751 = ~n15749 & ~n15750;
  assign n15752 = pi140 & n15751;
  assign n15753 = n8066 & ~n15746;
  assign n15754 = ~n8066 & ~n15383;
  assign n15755 = ~n15753 & ~n15754;
  assign n15756 = ~pi140 & n15755;
  assign n15757 = n8996 & ~n15756;
  assign n15758 = ~n15752 & n15757;
  assign n15759 = ~n14603 & ~n15702;
  assign n15760 = pi169 & n14987;
  assign n15761 = ~n15759 & ~n15760;
  assign n15762 = ~pi216 & ~n15761;
  assign n15763 = ~pi51 & ~n14999;
  assign n15764 = ~pi169 & n15763;
  assign n15765 = pi169 & n15743;
  assign n15766 = pi162 & pi216;
  assign n15767 = ~n15765 & n15766;
  assign n15768 = ~n15764 & n15767;
  assign n15769 = ~n15762 & ~n15768;
  assign n15770 = n6442 & ~n15769;
  assign n15771 = pi169 & n14531;
  assign n15772 = ~pi51 & ~n15771;
  assign n15773 = ~n8074 & ~n15698;
  assign n15774 = ~n15772 & n15773;
  assign n15775 = ~n15770 & ~n15774;
  assign n15776 = pi299 & ~n15775;
  assign n15777 = n14602 & n15002;
  assign n15778 = ~pi51 & ~n15777;
  assign n15779 = pi140 & n15778;
  assign n15780 = n8066 & n14602;
  assign n15781 = ~pi51 & ~n15780;
  assign n15782 = ~pi140 & n15781;
  assign n15783 = n15713 & ~n15782;
  assign n15784 = ~n15779 & n15783;
  assign n15785 = ~n15776 & ~n15784;
  assign n15786 = ~n15758 & n15785;
  assign n15787 = pi232 & ~n15786;
  assign n15788 = n14602 & ~n14981;
  assign n15789 = ~pi51 & ~n15788;
  assign n15790 = ~pi232 & ~n15789;
  assign n15791 = pi39 & ~n15790;
  assign n15792 = ~n15787 & n15791;
  assign n15793 = ~pi232 & ~n14499;
  assign n15794 = ~pi39 & ~n15793;
  assign n15795 = ~n6170 & n14499;
  assign n15796 = ~n14907 & ~n15795;
  assign n15797 = ~n8998 & ~n15796;
  assign n15798 = n8998 & n14499;
  assign n15799 = pi232 & ~n15798;
  assign n15800 = ~n15797 & n15799;
  assign n15801 = n15794 & ~n15800;
  assign n15802 = ~n15792 & ~n15801;
  assign n15803 = ~pi38 & ~n15802;
  assign n15804 = pi38 & ~n15727;
  assign n15805 = ~pi100 & ~n15804;
  assign n15806 = ~n15803 & n15805;
  assign n15807 = n15729 & ~n15806;
  assign n15808 = n15734 & n15740;
  assign n15809 = ~n15807 & n15808;
  assign n15810 = ~n15742 & ~n15809;
  assign n15811 = ~po1038 & ~n15810;
  assign n15812 = ~pi51 & ~pi87;
  assign n15813 = ~n15771 & n15812;
  assign n15814 = n15740 & n15813;
  assign n15815 = pi169 & n7484;
  assign n15816 = ~pi87 & n14443;
  assign n15817 = ~n15815 & n15816;
  assign n15818 = pi87 & ~n9690;
  assign n15819 = po1038 & ~n15818;
  assign n15820 = ~n15817 & n15819;
  assign n15821 = ~n15814 & n15820;
  assign po287 = ~n15811 & ~n15821;
  assign n15823 = ~pi100 & ~n13963;
  assign n15824 = ~pi87 & ~n7324;
  assign n15825 = ~n15823 & n15824;
  assign n15826 = ~pi75 & ~n15825;
  assign n15827 = ~n7292 & ~n15826;
  assign n15828 = ~pi92 & ~n15827;
  assign n15829 = n8866 & n13616;
  assign po288 = ~n15828 & n15829;
  assign n15831 = pi51 & ~pi151;
  assign n15832 = ~n13695 & ~n14397;
  assign n15833 = ~n15831 & ~n15832;
  assign n15834 = n14400 & n15833;
  assign n15835 = pi232 & n15834;
  assign n15836 = pi132 & ~n15349;
  assign n15837 = ~n15736 & ~n15836;
  assign n15838 = ~n14385 & ~n15837;
  assign n15839 = n14394 & ~n15838;
  assign n15840 = ~n15835 & ~n15839;
  assign n15841 = ~pi87 & ~n15840;
  assign n15842 = pi164 & n14874;
  assign n15843 = po1038 & ~n15842;
  assign n15844 = ~n15841 & n15843;
  assign n15845 = pi151 & n14499;
  assign n15846 = ~pi151 & ~n14505;
  assign n15847 = ~pi168 & ~n15845;
  assign n15848 = ~n15846 & n15847;
  assign n15849 = pi168 & ~n15831;
  assign n15850 = ~n14460 & n15849;
  assign n15851 = n6170 & ~n15850;
  assign n15852 = ~n15848 & n15851;
  assign n15853 = ~n6170 & ~n14516;
  assign n15854 = pi160 & ~n15853;
  assign n15855 = ~n15852 & n15854;
  assign n15856 = ~n6170 & n14516;
  assign n15857 = n14521 & ~n15856;
  assign n15858 = ~pi168 & ~n15857;
  assign n15859 = pi168 & ~n14921;
  assign n15860 = ~n15853 & n15859;
  assign n15861 = pi151 & ~n15860;
  assign n15862 = ~n15858 & n15861;
  assign n15863 = ~n13695 & n14516;
  assign n15864 = pi168 & n14527;
  assign n15865 = ~pi151 & ~n15864;
  assign n15866 = ~n15863 & n15865;
  assign n15867 = ~pi160 & ~n15866;
  assign n15868 = ~n15862 & n15867;
  assign n15869 = pi299 & ~n15868;
  assign n15870 = ~n15855 & n15869;
  assign n15871 = ~pi190 & ~pi299;
  assign n15872 = pi182 & ~n15853;
  assign n15873 = ~n14506 & n15872;
  assign n15874 = ~pi182 & n14516;
  assign n15875 = ~pi173 & ~n15874;
  assign n15876 = ~n15873 & n15875;
  assign n15877 = ~n14500 & ~n15856;
  assign n15878 = pi182 & ~n15877;
  assign n15879 = ~pi182 & ~n15857;
  assign n15880 = pi173 & ~n15879;
  assign n15881 = ~n15878 & n15880;
  assign n15882 = ~n15876 & ~n15881;
  assign n15883 = n15871 & ~n15882;
  assign n15884 = pi190 & ~pi299;
  assign n15885 = pi182 & n14451;
  assign n15886 = n14459 & ~n15885;
  assign n15887 = pi51 & ~pi173;
  assign n15888 = n6170 & ~n15887;
  assign n15889 = ~n15886 & n15888;
  assign n15890 = n15884 & ~n15889;
  assign n15891 = ~n15856 & n15890;
  assign n15892 = pi232 & ~n15891;
  assign n15893 = ~n15870 & n15892;
  assign n15894 = ~n15883 & n15893;
  assign n15895 = ~pi232 & n14516;
  assign n15896 = ~n15894 & ~n15895;
  assign n15897 = ~pi39 & ~n15896;
  assign n15898 = ~pi168 & n14764;
  assign n15899 = pi168 & n14626;
  assign n15900 = ~pi151 & ~n15899;
  assign n15901 = ~n15898 & n15900;
  assign n15902 = ~pi168 & ~n15000;
  assign n15903 = pi168 & ~n15042;
  assign n15904 = pi151 & ~n15903;
  assign n15905 = ~n15902 & n15904;
  assign n15906 = pi149 & ~n15901;
  assign n15907 = ~n15905 & n15906;
  assign n15908 = pi216 & ~n15907;
  assign n15909 = pi168 & ~n14988;
  assign n15910 = ~pi168 & ~n14990;
  assign n15911 = ~n15909 & ~n15910;
  assign n15912 = ~n15831 & ~n15911;
  assign n15913 = ~pi216 & ~n15912;
  assign n15914 = n6442 & ~n15908;
  assign n15915 = ~n15913 & n15914;
  assign n15916 = ~pi149 & pi216;
  assign n15917 = n6442 & ~n15916;
  assign n15918 = n15834 & ~n15917;
  assign n15919 = pi299 & ~n15918;
  assign n15920 = ~n15915 & n15919;
  assign n15921 = pi183 & ~n15022;
  assign n15922 = ~pi183 & ~n15017;
  assign n15923 = ~pi173 & ~n15922;
  assign n15924 = ~n15921 & n15923;
  assign n15925 = ~pi183 & n15031;
  assign n15926 = ~pi183 & ~n15007;
  assign n15927 = pi173 & ~n15012;
  assign n15928 = ~n15926 & n15927;
  assign n15929 = ~n15925 & ~n15928;
  assign n15930 = ~n15924 & n15929;
  assign n15931 = n15884 & ~n15930;
  assign n15932 = pi183 & n15005;
  assign n15933 = ~pi183 & ~n14397;
  assign n15934 = ~n15034 & n15933;
  assign n15935 = pi173 & ~n15934;
  assign n15936 = ~n15932 & n15935;
  assign n15937 = ~pi183 & ~n8066;
  assign n15938 = ~pi173 & ~n15937;
  assign n15939 = n15025 & n15938;
  assign n15940 = n15871 & ~n15939;
  assign n15941 = ~n15936 & n15940;
  assign n15942 = ~n15931 & ~n15941;
  assign n15943 = ~n15920 & n15942;
  assign n15944 = pi232 & ~n15943;
  assign n15945 = n14984 & ~n15944;
  assign n15946 = ~n15897 & ~n15945;
  assign n15947 = n3207 & ~n15946;
  assign n15948 = pi190 & n14531;
  assign n15949 = pi173 & n14397;
  assign n15950 = ~pi299 & ~n15949;
  assign n15951 = ~n15948 & n15950;
  assign n15952 = pi299 & ~n15834;
  assign n15953 = pi232 & ~n15951;
  assign n15954 = ~n15952 & n15953;
  assign n15955 = ~n3207 & n15954;
  assign n15956 = n3279 & ~n15955;
  assign n15957 = ~n15947 & n15956;
  assign n15958 = n14685 & ~n15954;
  assign n15959 = pi87 & ~n9006;
  assign n15960 = n15838 & ~n15959;
  assign n15961 = ~n15958 & n15960;
  assign n15962 = ~n15957 & n15961;
  assign n15963 = ~n14394 & n15952;
  assign n15964 = ~n13094 & ~n15963;
  assign n15965 = pi168 & ~n14600;
  assign n15966 = ~pi168 & ~n14631;
  assign n15967 = pi151 & ~n15966;
  assign n15968 = ~n15965 & n15967;
  assign n15969 = pi168 & n14604;
  assign n15970 = ~n13695 & ~n14598;
  assign n15971 = ~pi151 & ~n15970;
  assign n15972 = ~n15969 & n15971;
  assign n15973 = ~pi149 & ~n15972;
  assign n15974 = ~n15968 & n15973;
  assign n15975 = ~n15000 & ~n15831;
  assign n15976 = ~n14605 & ~n15975;
  assign n15977 = pi168 & ~n15976;
  assign n15978 = ~n14654 & ~n15833;
  assign n15979 = ~pi168 & ~n15978;
  assign n15980 = pi149 & ~n15979;
  assign n15981 = ~n15977 & n15980;
  assign n15982 = n9055 & ~n15974;
  assign n15983 = ~n15981 & n15982;
  assign n15984 = ~n15964 & ~n15983;
  assign n15985 = ~pi183 & ~n15209;
  assign n15986 = pi183 & ~n15219;
  assign n15987 = pi173 & ~n15986;
  assign n15988 = ~n15985 & n15987;
  assign n15989 = pi183 & n14611;
  assign n15990 = ~pi173 & ~n15989;
  assign n15991 = n15231 & n15990;
  assign n15992 = ~n15988 & ~n15991;
  assign n15993 = n15884 & ~n15992;
  assign n15994 = pi183 & n14654;
  assign n15995 = n15871 & ~n15949;
  assign n15996 = ~n15212 & n15995;
  assign n15997 = ~n15994 & n15996;
  assign n15998 = ~n15984 & ~n15997;
  assign n15999 = ~n15993 & n15998;
  assign n16000 = pi232 & ~n15999;
  assign n16001 = ~n15249 & ~n16000;
  assign n16002 = pi39 & ~n16001;
  assign n16003 = pi151 & n14736;
  assign n16004 = ~pi151 & ~n14452;
  assign n16005 = ~pi168 & ~n16004;
  assign n16006 = ~n16003 & n16005;
  assign n16007 = ~pi151 & n14397;
  assign n16008 = pi168 & ~n16007;
  assign n16009 = ~n14473 & n16008;
  assign n16010 = ~n16006 & ~n16009;
  assign n16011 = ~pi160 & ~n15096;
  assign n16012 = ~n16010 & n16011;
  assign n16013 = ~pi168 & n14531;
  assign n16014 = ~n15096 & ~n16013;
  assign n16015 = pi151 & ~n16014;
  assign n16016 = ~pi151 & ~n15834;
  assign n16017 = ~n15097 & n16016;
  assign n16018 = pi160 & ~n16015;
  assign n16019 = ~n16017 & n16018;
  assign n16020 = pi299 & ~n16019;
  assign n16021 = ~n16012 & n16020;
  assign n16022 = ~pi182 & n14473;
  assign n16023 = ~n15096 & ~n15887;
  assign n16024 = ~n16022 & n16023;
  assign n16025 = n15884 & ~n16024;
  assign n16026 = pi182 & n15097;
  assign n16027 = ~n14452 & n15995;
  assign n16028 = ~n16026 & n16027;
  assign n16029 = pi232 & ~n16028;
  assign n16030 = ~n16025 & n16029;
  assign n16031 = ~n16021 & n16030;
  assign n16032 = ~pi232 & n14452;
  assign n16033 = ~pi39 & ~n16032;
  assign n16034 = ~n16031 & n16033;
  assign n16035 = n3207 & ~n16034;
  assign n16036 = ~n16002 & n16035;
  assign n16037 = n3279 & ~n15543;
  assign n16038 = ~n15955 & n16037;
  assign n16039 = ~n16036 & n16038;
  assign n16040 = n14686 & ~n15954;
  assign n16041 = ~n15838 & ~n15959;
  assign n16042 = ~n16040 & n16041;
  assign n16043 = ~n16039 & n16042;
  assign n16044 = ~po1038 & ~n16043;
  assign n16045 = ~n15962 & n16044;
  assign po289 = n15844 | n16045;
  assign n16047 = ~n6170 & ~n14478;
  assign n16048 = ~n14506 & ~n16047;
  assign n16049 = n9451 & n16048;
  assign n16050 = ~n9451 & n14478;
  assign n16051 = ~pi39 & pi176;
  assign n16052 = ~n16050 & n16051;
  assign n16053 = ~n16049 & n16052;
  assign n16054 = pi299 & n9451;
  assign n16055 = n16048 & n16054;
  assign n16056 = n14478 & ~n16054;
  assign n16057 = ~pi39 & ~pi176;
  assign n16058 = ~n16056 & n16057;
  assign n16059 = ~n16055 & n16058;
  assign n16060 = pi197 & n14610;
  assign n16061 = ~n5752 & ~n16060;
  assign n16062 = n6595 & ~n16061;
  assign n16063 = ~pi145 & ~n8066;
  assign n16064 = ~pi299 & ~n16063;
  assign n16065 = ~n15024 & n16064;
  assign n16066 = ~n16062 & ~n16065;
  assign n16067 = n3096 & ~n16066;
  assign n16068 = pi232 & ~n16067;
  assign n16069 = ~n14983 & ~n16068;
  assign n16070 = pi39 & ~n16069;
  assign n16071 = n11357 & ~n16070;
  assign n16072 = ~n16053 & n16071;
  assign n16073 = ~n16059 & n16072;
  assign n16074 = ~pi133 & ~n14863;
  assign n16075 = ~pi87 & n16074;
  assign n16076 = ~n16073 & n16075;
  assign n16077 = pi145 & n14654;
  assign n16078 = n15244 & ~n16077;
  assign n16079 = n15245 & ~n16060;
  assign n16080 = n14394 & ~n16079;
  assign n16081 = pi299 & ~n16080;
  assign n16082 = ~n16078 & ~n16081;
  assign n16083 = pi232 & ~n16082;
  assign n16084 = n15250 & ~n16083;
  assign n16085 = ~n9454 & n14446;
  assign n16086 = ~pi39 & n14394;
  assign n16087 = ~n16085 & n16086;
  assign n16088 = ~pi38 & ~n16087;
  assign n16089 = ~n16084 & n16088;
  assign n16090 = n14422 & ~n16089;
  assign n16091 = n14681 & ~n16090;
  assign n16092 = ~n14686 & ~n16091;
  assign n16093 = ~n16074 & ~n16092;
  assign n16094 = ~pi183 & ~pi299;
  assign n16095 = ~pi149 & pi299;
  assign n16096 = ~n16094 & ~n16095;
  assign n16097 = n7484 & n16096;
  assign n16098 = pi87 & ~n16097;
  assign n16099 = ~n16093 & ~n16098;
  assign n16100 = ~n16076 & n16099;
  assign n16101 = ~po1038 & ~n16100;
  assign n16102 = n14395 & ~n16074;
  assign n16103 = pi149 & n14874;
  assign n16104 = po1038 & ~n16103;
  assign n16105 = ~n16102 & n16104;
  assign po290 = n16101 | n16105;
  assign n16107 = ~pi136 & n15738;
  assign n16108 = ~pi135 & n16107;
  assign n16109 = pi134 & ~n16108;
  assign n16110 = n14393 & ~n16109;
  assign n16111 = po1038 & n15812;
  assign n16112 = pi171 & n6170;
  assign n16113 = ~n14393 & n16112;
  assign n16114 = pi232 & n16113;
  assign n16115 = n16111 & ~n16114;
  assign n16116 = ~n16110 & n16115;
  assign n16117 = pi39 & pi186;
  assign n16118 = pi192 & ~pi299;
  assign n16119 = ~n14610 & n15691;
  assign n16120 = n16118 & ~n16119;
  assign n16121 = ~pi192 & ~pi299;
  assign n16122 = ~n15222 & n15714;
  assign n16123 = n16121 & ~n16122;
  assign n16124 = ~n16120 & ~n16123;
  assign n16125 = n15708 & ~n16112;
  assign n16126 = pi299 & ~n16125;
  assign n16127 = n4221 & n6170;
  assign n16128 = ~n14623 & ~n16112;
  assign n16129 = n9055 & ~n16128;
  assign n16130 = ~n16127 & n16129;
  assign n16131 = n16126 & ~n16130;
  assign n16132 = n16124 & ~n16131;
  assign n16133 = pi232 & ~n16132;
  assign n16134 = ~n15689 & ~n16133;
  assign n16135 = n16117 & ~n16134;
  assign n16136 = pi39 & ~pi186;
  assign n16137 = ~n15691 & n16118;
  assign n16138 = ~n15714 & n16121;
  assign n16139 = ~n16137 & ~n16138;
  assign n16140 = ~n16131 & n16139;
  assign n16141 = pi232 & ~n16140;
  assign n16142 = ~n15689 & ~n16141;
  assign n16143 = n16136 & ~n16142;
  assign n16144 = pi171 & pi299;
  assign n16145 = ~n16118 & ~n16144;
  assign n16146 = n7484 & ~n16145;
  assign n16147 = n14443 & ~n16146;
  assign n16148 = ~pi39 & ~n16147;
  assign n16149 = ~pi164 & ~n16148;
  assign n16150 = ~n16143 & n16149;
  assign n16151 = ~n16135 & n16150;
  assign n16152 = pi171 & ~n15696;
  assign n16153 = ~pi171 & ~n15221;
  assign n16154 = n9055 & ~n16153;
  assign n16155 = ~n16152 & n16154;
  assign n16156 = n16126 & ~n16155;
  assign n16157 = n16124 & ~n16156;
  assign n16158 = pi232 & ~n16157;
  assign n16159 = ~n15689 & ~n16158;
  assign n16160 = n16117 & ~n16159;
  assign n16161 = n16139 & ~n16156;
  assign n16162 = pi232 & ~n16161;
  assign n16163 = ~n15689 & ~n16162;
  assign n16164 = n16136 & ~n16163;
  assign n16165 = pi164 & ~n16148;
  assign n16166 = ~n16164 & n16165;
  assign n16167 = ~n16160 & n16166;
  assign n16168 = n3207 & ~n16151;
  assign n16169 = ~n16167 & n16168;
  assign n16170 = ~n15383 & ~n16147;
  assign n16171 = ~n3207 & n16170;
  assign n16172 = n3279 & ~n16171;
  assign n16173 = ~n15543 & n16172;
  assign n16174 = ~n16169 & n16173;
  assign n16175 = n14685 & n16147;
  assign n16176 = ~n16109 & ~n16175;
  assign n16177 = ~n16174 & n16176;
  assign n16178 = ~pi51 & ~n16113;
  assign n16179 = ~pi164 & pi216;
  assign n16180 = n6442 & ~n16179;
  assign n16181 = ~n16178 & ~n16180;
  assign n16182 = ~n14603 & ~n16112;
  assign n16183 = pi171 & n14987;
  assign n16184 = ~n16182 & ~n16183;
  assign n16185 = ~pi216 & ~n16184;
  assign n16186 = ~pi171 & n15763;
  assign n16187 = pi171 & n15743;
  assign n16188 = pi164 & pi216;
  assign n16189 = ~n16187 & n16188;
  assign n16190 = ~n16186 & n16189;
  assign n16191 = ~n16185 & ~n16190;
  assign n16192 = n6442 & ~n16191;
  assign n16193 = ~n16181 & ~n16192;
  assign n16194 = pi299 & ~n16193;
  assign n16195 = ~n15755 & n16118;
  assign n16196 = ~n15781 & n16121;
  assign n16197 = ~n16117 & ~n16196;
  assign n16198 = ~n16195 & n16197;
  assign n16199 = ~n15751 & n16118;
  assign n16200 = ~n15778 & n16121;
  assign n16201 = pi186 & ~n16200;
  assign n16202 = ~n16199 & n16201;
  assign n16203 = ~n16198 & ~n16202;
  assign n16204 = ~n16194 & ~n16203;
  assign n16205 = pi232 & ~n16204;
  assign n16206 = n15791 & ~n16205;
  assign n16207 = pi232 & ~n16145;
  assign n16208 = n15796 & n16207;
  assign n16209 = ~n14499 & ~n16207;
  assign n16210 = ~pi39 & ~n16209;
  assign n16211 = ~n16208 & n16210;
  assign n16212 = n3207 & ~n16206;
  assign n16213 = ~n16211 & n16212;
  assign n16214 = n16172 & ~n16213;
  assign n16215 = n14685 & ~n16170;
  assign n16216 = n16109 & ~n16215;
  assign n16217 = ~n16214 & n16216;
  assign n16218 = ~po1038 & ~n16217;
  assign n16219 = ~n16177 & n16218;
  assign po291 = n16116 | n16219;
  assign n16221 = pi170 & n6170;
  assign n16222 = n10531 & n16221;
  assign n16223 = n14443 & ~n16222;
  assign n16224 = pi194 & n9017;
  assign n16225 = n16223 & ~n16224;
  assign n16226 = ~n15383 & ~n16225;
  assign n16227 = pi100 & n16226;
  assign n16228 = n3279 & ~n16227;
  assign n16229 = ~n14603 & ~n16221;
  assign n16230 = pi170 & n14987;
  assign n16231 = n8074 & ~n16230;
  assign n16232 = ~n16229 & n16231;
  assign n16233 = ~n9055 & ~n16232;
  assign n16234 = ~pi170 & n15763;
  assign n16235 = pi170 & n15743;
  assign n16236 = pi216 & ~n16235;
  assign n16237 = ~n16234 & n16236;
  assign n16238 = ~n16233 & ~n16237;
  assign n16239 = pi150 & pi299;
  assign n16240 = ~n14393 & n16221;
  assign n16241 = ~pi51 & ~n16240;
  assign n16242 = ~n6442 & n16241;
  assign n16243 = n16239 & ~n16242;
  assign n16244 = ~n16238 & n16243;
  assign n16245 = ~n8074 & n16241;
  assign n16246 = n15549 & ~n16245;
  assign n16247 = ~n16232 & n16246;
  assign n16248 = ~n16244 & ~n16247;
  assign n16249 = pi185 & n15778;
  assign n16250 = ~pi185 & n15781;
  assign n16251 = ~pi299 & ~n16250;
  assign n16252 = ~n16249 & n16251;
  assign n16253 = n16248 & ~n16252;
  assign n16254 = pi232 & ~n16253;
  assign n16255 = n15791 & ~n16254;
  assign n16256 = ~pi299 & ~n14499;
  assign n16257 = pi170 & ~n15796;
  assign n16258 = ~pi170 & n14499;
  assign n16259 = n10531 & ~n16258;
  assign n16260 = ~n16257 & n16259;
  assign n16261 = n15794 & ~n16260;
  assign n16262 = ~n16256 & n16261;
  assign n16263 = ~n16255 & ~n16262;
  assign n16264 = ~pi38 & ~n16263;
  assign n16265 = ~n15383 & ~n16223;
  assign n16266 = pi38 & ~n16265;
  assign n16267 = ~pi194 & ~n16266;
  assign n16268 = ~n16264 & n16267;
  assign n16269 = pi185 & n15751;
  assign n16270 = ~pi185 & n15755;
  assign n16271 = ~pi299 & ~n16270;
  assign n16272 = ~n16269 & n16271;
  assign n16273 = n16248 & ~n16272;
  assign n16274 = pi232 & ~n16273;
  assign n16275 = n15791 & ~n16274;
  assign n16276 = n10526 & n15796;
  assign n16277 = n16261 & ~n16276;
  assign n16278 = ~n16275 & ~n16277;
  assign n16279 = ~pi38 & ~n16278;
  assign n16280 = pi170 & n7484;
  assign n16281 = ~n9017 & ~n16280;
  assign n16282 = n14443 & n16281;
  assign n16283 = ~n15383 & ~n16282;
  assign n16284 = pi38 & ~n16283;
  assign n16285 = pi194 & ~n16284;
  assign n16286 = ~n16279 & n16285;
  assign n16287 = ~n16268 & ~n16286;
  assign n16288 = ~pi100 & ~n16287;
  assign n16289 = n16228 & ~n16288;
  assign n16290 = pi135 & ~n16107;
  assign n16291 = pi134 & n16108;
  assign n16292 = ~n16290 & ~n16291;
  assign n16293 = n14685 & ~n16226;
  assign n16294 = ~n16292 & ~n16293;
  assign n16295 = ~n16289 & n16294;
  assign n16296 = pi185 & n15222;
  assign n16297 = n15714 & ~n16296;
  assign n16298 = ~n10959 & n16223;
  assign n16299 = ~pi194 & ~n16298;
  assign n16300 = ~n16297 & n16299;
  assign n16301 = ~pi185 & n15691;
  assign n16302 = ~n10959 & n16282;
  assign n16303 = pi194 & ~n16302;
  assign n16304 = ~n16119 & n16303;
  assign n16305 = ~n16301 & n16304;
  assign n16306 = ~n16300 & ~n16305;
  assign n16307 = ~pi299 & ~n16306;
  assign n16308 = pi170 & ~n15696;
  assign n16309 = ~pi170 & ~n15221;
  assign n16310 = n9055 & ~n16309;
  assign n16311 = ~n16308 & n16310;
  assign n16312 = n16239 & ~n16311;
  assign n16313 = n4443 & n6170;
  assign n16314 = ~n14623 & ~n16221;
  assign n16315 = n9055 & ~n16314;
  assign n16316 = ~n16313 & n16315;
  assign n16317 = n15549 & ~n16316;
  assign n16318 = ~n16312 & ~n16317;
  assign n16319 = n15708 & ~n16221;
  assign n16320 = ~n16299 & ~n16303;
  assign n16321 = ~n16319 & ~n16320;
  assign n16322 = ~n16318 & n16321;
  assign n16323 = ~n16307 & ~n16322;
  assign n16324 = pi232 & ~n16323;
  assign n16325 = ~n15690 & ~n16320;
  assign n16326 = ~n16324 & ~n16325;
  assign n16327 = ~pi100 & ~n16326;
  assign n16328 = ~n14680 & n16228;
  assign n16329 = ~n16327 & n16328;
  assign n16330 = n14685 & n16225;
  assign n16331 = n16292 & ~n16330;
  assign n16332 = ~n16329 & n16331;
  assign n16333 = ~po1038 & ~n16332;
  assign n16334 = ~n16295 & n16333;
  assign n16335 = n14393 & n16292;
  assign n16336 = ~n14393 & n16280;
  assign n16337 = n16111 & ~n16336;
  assign n16338 = ~n16335 & n16337;
  assign po292 = n16334 | n16338;
  assign n16340 = pi136 & ~n15738;
  assign n16341 = ~n16107 & ~n16340;
  assign n16342 = ~n14383 & ~n16341;
  assign n16343 = ~n14443 & n16342;
  assign n16344 = pi148 & n7484;
  assign n16345 = ~n14393 & ~n16344;
  assign n16346 = ~n16343 & ~n16345;
  assign n16347 = n16111 & ~n16346;
  assign n16348 = ~n9726 & ~n15796;
  assign n16349 = n9726 & n14499;
  assign n16350 = pi232 & ~n16349;
  assign n16351 = ~n16348 & n16350;
  assign n16352 = n15794 & ~n16351;
  assign n16353 = pi184 & n15751;
  assign n16354 = ~pi184 & n15755;
  assign n16355 = n9724 & ~n16354;
  assign n16356 = ~n16353 & n16355;
  assign n16357 = pi184 & n15778;
  assign n16358 = ~pi141 & ~pi299;
  assign n16359 = ~pi184 & n15781;
  assign n16360 = n16358 & ~n16359;
  assign n16361 = ~n16357 & n16360;
  assign n16362 = n8074 & ~n15746;
  assign n16363 = pi163 & n6442;
  assign n16364 = n15743 & n16363;
  assign n16365 = ~n6442 & n15383;
  assign n16366 = ~n8074 & ~n15383;
  assign n16367 = ~pi163 & ~n16366;
  assign n16368 = ~n16365 & ~n16367;
  assign n16369 = ~n16364 & n16368;
  assign n16370 = pi148 & ~n16369;
  assign n16371 = ~n16362 & n16370;
  assign n16372 = ~pi287 & n13626;
  assign n16373 = pi216 & ~n16372;
  assign n16374 = n6442 & ~n16373;
  assign n16375 = n14602 & n16374;
  assign n16376 = ~pi51 & ~pi148;
  assign n16377 = ~n16375 & n16376;
  assign n16378 = pi299 & ~n16377;
  assign n16379 = ~n16371 & n16378;
  assign n16380 = ~n16361 & ~n16379;
  assign n16381 = ~n16356 & n16380;
  assign n16382 = pi232 & ~n16381;
  assign n16383 = n15791 & ~n16382;
  assign n16384 = n3207 & ~n16383;
  assign n16385 = ~n16352 & n16384;
  assign n16386 = n9727 & ~n14393;
  assign n16387 = ~pi51 & ~n16386;
  assign n16388 = ~n3207 & ~n16387;
  assign n16389 = n3279 & ~n16388;
  assign n16390 = ~n16385 & n16389;
  assign n16391 = n14685 & n16387;
  assign n16392 = n16342 & ~n16391;
  assign n16393 = ~n16390 & n16392;
  assign n16394 = ~n11103 & ~n14393;
  assign n16395 = n16387 & n16394;
  assign n16396 = pi184 & n14610;
  assign n16397 = n15691 & ~n16396;
  assign n16398 = n9724 & ~n16397;
  assign n16399 = n9055 & n15695;
  assign n16400 = ~n6170 & n15708;
  assign n16401 = pi148 & ~n16400;
  assign n16402 = ~n16399 & n16401;
  assign n16403 = ~pi51 & n15245;
  assign n16404 = ~pi148 & ~n16403;
  assign n16405 = ~n16372 & ~n16404;
  assign n16406 = ~pi148 & n14443;
  assign n16407 = ~n16405 & ~n16406;
  assign n16408 = ~n16402 & ~n16407;
  assign n16409 = pi299 & ~n16408;
  assign n16410 = pi184 & n15222;
  assign n16411 = n15714 & ~n16410;
  assign n16412 = n16358 & ~n16411;
  assign n16413 = ~n16398 & ~n16412;
  assign n16414 = ~n16409 & n16413;
  assign n16415 = pi232 & ~n16414;
  assign n16416 = ~pi100 & n15690;
  assign n16417 = ~n16415 & n16416;
  assign n16418 = ~n16395 & ~n16417;
  assign n16419 = n3279 & ~n16418;
  assign n16420 = ~n14393 & n16391;
  assign n16421 = ~n16342 & ~n16420;
  assign n16422 = ~n16419 & n16421;
  assign n16423 = ~po1038 & ~n16422;
  assign n16424 = ~n16393 & n16423;
  assign po293 = n16347 | n16424;
  assign n16426 = ~pi39 & pi137;
  assign n16427 = n10413 & n14819;
  assign n16428 = n6150 & n11544;
  assign n16429 = ~pi299 & ~po1038;
  assign n16430 = ~pi198 & n11555;
  assign n16431 = n16429 & n16430;
  assign n16432 = ~n16428 & ~n16431;
  assign n16433 = ~n16427 & ~n16432;
  assign n16434 = ~pi210 & n11544;
  assign n16435 = po1038 & n16434;
  assign n16436 = ~n16433 & ~n16435;
  assign n16437 = n10457 & ~n16436;
  assign po294 = n16426 | n16437;
  assign n16439 = ~n9455 & n9505;
  assign n16440 = pi92 & ~n16439;
  assign n16441 = n3266 & ~n16440;
  assign n16442 = ~pi75 & ~n9446;
  assign n16443 = pi299 & ~n9384;
  assign n16444 = ~pi299 & ~n9774;
  assign n16445 = ~pi232 & ~n16443;
  assign n16446 = ~n16444 & n16445;
  assign n16447 = ~pi39 & ~n16446;
  assign n16448 = ~n6170 & ~n9774;
  assign n16449 = ~n13706 & ~n16448;
  assign n16450 = ~pi299 & ~n16449;
  assign n16451 = pi141 & n16450;
  assign n16452 = pi148 & n6170;
  assign n16453 = ~n9384 & ~n16452;
  assign n16454 = pi148 & n13683;
  assign n16455 = ~n16453 & ~n16454;
  assign n16456 = pi299 & ~n16455;
  assign n16457 = ~pi141 & n16444;
  assign n16458 = pi232 & ~n16457;
  assign n16459 = ~n16451 & n16458;
  assign n16460 = ~n16456 & n16459;
  assign n16461 = n16447 & ~n16460;
  assign n16462 = ~n9064 & ~n11966;
  assign n16463 = n9080 & ~n16462;
  assign n16464 = n13755 & ~n16463;
  assign n16465 = ~n6223 & ~n9064;
  assign n16466 = n9055 & ~n16462;
  assign n16467 = ~n16465 & n16466;
  assign n16468 = n9057 & ~n16467;
  assign n16469 = ~n16464 & ~n16468;
  assign n16470 = ~pi232 & ~n16469;
  assign n16471 = ~n9060 & ~n16462;
  assign n16472 = ~n9056 & ~n16471;
  assign n16473 = pi148 & ~n16472;
  assign n16474 = ~n9725 & ~n16468;
  assign n16475 = ~n16473 & ~n16474;
  assign n16476 = ~pi141 & n16464;
  assign n16477 = ~n9088 & n16463;
  assign n16478 = n13755 & ~n16477;
  assign n16479 = pi141 & n16478;
  assign n16480 = ~n16476 & ~n16479;
  assign n16481 = ~n16475 & n16480;
  assign n16482 = pi232 & ~n16481;
  assign n16483 = ~n16470 & ~n16482;
  assign n16484 = pi39 & ~n16483;
  assign n16485 = n3207 & ~n16484;
  assign n16486 = ~n16461 & n16485;
  assign n16487 = ~pi87 & ~n16486;
  assign n16488 = n16442 & ~n16487;
  assign n16489 = ~pi92 & ~n16488;
  assign n16490 = n16441 & ~n16489;
  assign n16491 = ~pi55 & ~n16490;
  assign n16492 = n9506 & ~n13792;
  assign n16493 = pi55 & ~n16492;
  assign n16494 = ~n16491 & ~n16493;
  assign n16495 = n3294 & ~n16494;
  assign n16496 = n9707 & ~n16495;
  assign n16497 = pi138 & n16496;
  assign n16498 = ~pi232 & ~n11452;
  assign n16499 = ~n9724 & ~n11452;
  assign n16500 = n6206 & n6459;
  assign n16501 = n9044 & n16500;
  assign n16502 = n9724 & ~n16501;
  assign n16503 = ~n6206 & n9725;
  assign n16504 = ~n16502 & ~n16503;
  assign n16505 = ~n16499 & n16504;
  assign n16506 = pi232 & ~n16505;
  assign n16507 = ~n16498 & ~n16506;
  assign n16508 = pi39 & ~n16507;
  assign n16509 = ~n9727 & n13862;
  assign n16510 = ~pi39 & ~n16509;
  assign n16511 = n10181 & ~n16510;
  assign n16512 = ~n16508 & n16511;
  assign n16513 = ~pi138 & n16512;
  assign n16514 = ~pi118 & n13810;
  assign n16515 = ~pi139 & n16514;
  assign n16516 = ~n16513 & ~n16515;
  assign n16517 = ~n16497 & n16516;
  assign n16518 = ~pi138 & ~n8960;
  assign n16519 = n16496 & n16518;
  assign n16520 = n16512 & ~n16518;
  assign n16521 = n16515 & ~n16520;
  assign n16522 = ~n16519 & n16521;
  assign po295 = ~n16517 & ~n16522;
  assign n16524 = pi191 & n16450;
  assign n16525 = ~n9384 & ~n15702;
  assign n16526 = pi169 & n13683;
  assign n16527 = ~n16525 & ~n16526;
  assign n16528 = pi299 & ~n16527;
  assign n16529 = ~pi191 & n16444;
  assign n16530 = pi232 & ~n16529;
  assign n16531 = ~n16524 & n16530;
  assign n16532 = ~n16528 & n16531;
  assign n16533 = n16447 & ~n16532;
  assign n16534 = ~pi169 & n9064;
  assign n16535 = ~n16471 & ~n16534;
  assign n16536 = n9055 & ~n16535;
  assign n16537 = n9057 & ~n16536;
  assign n16538 = pi191 & n16478;
  assign n16539 = ~pi191 & n16464;
  assign n16540 = ~n16537 & ~n16539;
  assign n16541 = ~n16538 & n16540;
  assign n16542 = pi232 & ~n16541;
  assign n16543 = ~n16470 & ~n16542;
  assign n16544 = pi39 & ~n16543;
  assign n16545 = n3207 & ~n16544;
  assign n16546 = ~n16533 & n16545;
  assign n16547 = ~pi87 & ~n16546;
  assign n16548 = n16442 & ~n16547;
  assign n16549 = ~pi92 & ~n16548;
  assign n16550 = n16441 & ~n16549;
  assign n16551 = ~pi55 & ~n16550;
  assign n16552 = ~n16493 & ~n16551;
  assign n16553 = n3294 & ~n16552;
  assign n16554 = n9707 & ~n16553;
  assign n16555 = pi139 & n16554;
  assign n16556 = ~n6206 & n8997;
  assign n16557 = ~n11448 & n15713;
  assign n16558 = n8996 & ~n16501;
  assign n16559 = ~n11451 & ~n16556;
  assign n16560 = ~n16557 & ~n16558;
  assign n16561 = n16559 & n16560;
  assign n16562 = pi232 & ~n16561;
  assign n16563 = ~n16498 & ~n16562;
  assign n16564 = pi39 & ~n16563;
  assign n16565 = n13862 & ~n15722;
  assign n16566 = ~pi39 & ~n16565;
  assign n16567 = n10181 & ~n16566;
  assign n16568 = ~n16564 & n16567;
  assign n16569 = ~pi139 & n16568;
  assign n16570 = ~n16514 & ~n16569;
  assign n16571 = ~n16555 & n16570;
  assign n16572 = ~pi139 & ~n8961;
  assign n16573 = n16554 & n16572;
  assign n16574 = n16568 & ~n16572;
  assign n16575 = n16514 & ~n16574;
  assign n16576 = ~n16573 & n16575;
  assign po296 = ~n16571 & ~n16576;
  assign n16578 = pi140 & ~n3268;
  assign n16579 = ~pi102 & ~n11276;
  assign n16580 = ~pi98 & ~n2596;
  assign n16581 = ~n16579 & n16580;
  assign n16582 = n7451 & n12166;
  assign n16583 = n16581 & n16582;
  assign n16584 = n8885 & n9154;
  assign n16585 = n16583 & n16584;
  assign n16586 = ~pi40 & ~n16585;
  assign n16587 = n10262 & ~n16586;
  assign n16588 = ~pi252 & ~n16587;
  assign n16589 = n2534 & n2572;
  assign n16590 = n8884 & n16583;
  assign n16591 = ~pi47 & ~n16590;
  assign n16592 = pi314 & n10237;
  assign n16593 = n16591 & ~n16592;
  assign n16594 = n16589 & ~n16593;
  assign n16595 = ~pi35 & ~n16594;
  assign n16596 = ~pi40 & n10255;
  assign n16597 = ~n16595 & n16596;
  assign n16598 = pi252 & ~n2553;
  assign n16599 = ~n16597 & n16598;
  assign n16600 = ~n16588 & ~n16599;
  assign n16601 = n3093 & n16600;
  assign n16602 = pi1092 & ~n12178;
  assign n16603 = n16601 & n16602;
  assign n16604 = ~pi88 & ~n16581;
  assign n16605 = n10983 & ~n16604;
  assign n16606 = n2519 & n16605;
  assign n16607 = ~pi47 & ~n16592;
  assign n16608 = ~n16606 & n16607;
  assign n16609 = n16589 & ~n16608;
  assign n16610 = ~pi35 & ~n16609;
  assign n16611 = pi252 & n10255;
  assign n16612 = ~n16610 & n16611;
  assign n16613 = ~pi252 & n9272;
  assign n16614 = n16605 & n16613;
  assign n16615 = ~pi40 & ~n16614;
  assign n16616 = ~n16612 & n16615;
  assign n16617 = n7496 & n10262;
  assign n16618 = ~n16616 & n16617;
  assign n16619 = ~n16603 & ~n16618;
  assign n16620 = pi1093 & ~n16619;
  assign n16621 = ~n2733 & ~n16620;
  assign n16622 = pi1092 & n10053;
  assign po1106 = n2733 & n16622;
  assign n16624 = n16601 & po1106;
  assign n16625 = ~n2734 & ~n16624;
  assign n16626 = ~n16621 & ~n16625;
  assign n16627 = ~pi1091 & n16620;
  assign n16628 = ~n16626 & ~n16627;
  assign n16629 = ~pi210 & n16628;
  assign n16630 = ~n3362 & ~n16616;
  assign n16631 = ~pi32 & ~n16630;
  assign n16632 = pi32 & ~n6377;
  assign n16633 = ~pi95 & n6265;
  assign n16634 = ~n16632 & n16633;
  assign n16635 = ~n16631 & n16634;
  assign n16636 = pi824 & n16635;
  assign n16637 = ~n16603 & ~n16636;
  assign n16638 = n7558 & ~n16637;
  assign n16639 = ~pi32 & ~n16600;
  assign n16640 = n16634 & ~n16639;
  assign n16641 = ~pi824 & pi829;
  assign n16642 = n16640 & n16641;
  assign n16643 = n16637 & ~n16642;
  assign n16644 = pi1093 & ~n16643;
  assign n16645 = ~n2733 & ~n16644;
  assign n16646 = ~n16625 & ~n16645;
  assign n16647 = ~n16638 & ~n16646;
  assign n16648 = pi210 & n16647;
  assign n16649 = ~n16629 & ~n16648;
  assign n16650 = pi299 & ~n16649;
  assign n16651 = ~pi198 & n16628;
  assign n16652 = pi198 & n16647;
  assign n16653 = ~n16651 & ~n16652;
  assign n16654 = ~pi299 & ~n16653;
  assign n16655 = ~n16650 & ~n16654;
  assign n16656 = ~pi39 & ~n16655;
  assign n16657 = ~n6174 & n6443;
  assign n16658 = ~pi120 & ~n16657;
  assign n16659 = pi120 & ~n3096;
  assign n16660 = ~n16658 & ~n16659;
  assign n16661 = n2755 & n16660;
  assign n16662 = ~n6170 & n16661;
  assign n16663 = n2755 & n16657;
  assign n16664 = ~pi120 & ~n16663;
  assign n16665 = n2755 & n3096;
  assign n16666 = n6177 & n14239;
  assign n16667 = n16665 & ~n16666;
  assign n16668 = pi120 & ~n16667;
  assign n16669 = pi1091 & ~n16668;
  assign n16670 = ~n16664 & n16669;
  assign n16671 = pi120 & ~n16665;
  assign n16672 = ~pi1091 & ~n16671;
  assign n16673 = pi120 & pi824;
  assign n16674 = n6177 & n16673;
  assign n16675 = n16672 & ~n16674;
  assign n16676 = ~n16664 & n16675;
  assign n16677 = ~n16670 & ~n16676;
  assign n16678 = n6170 & ~n16677;
  assign n16679 = ~n16662 & ~n16678;
  assign n16680 = ~n6163 & ~n16661;
  assign n16681 = ~n6170 & n16677;
  assign n16682 = n6170 & ~n16661;
  assign n16683 = ~n16681 & ~n16682;
  assign n16684 = n6163 & ~n16683;
  assign n16685 = ~n16680 & ~n16684;
  assign n16686 = ~pi614 & ~n16685;
  assign n16687 = ~pi616 & n16686;
  assign n16688 = ~n16679 & ~n16687;
  assign n16689 = pi681 & ~n16688;
  assign n16690 = pi616 & ~n16661;
  assign n16691 = pi614 & ~n16661;
  assign n16692 = ~n16686 & ~n16691;
  assign n16693 = ~pi616 & ~n16692;
  assign n16694 = ~n16690 & ~n16693;
  assign n16695 = ~n6166 & ~n16694;
  assign n16696 = n6166 & n16677;
  assign n16697 = ~n6170 & ~n16696;
  assign n16698 = ~n16695 & n16697;
  assign n16699 = ~n16678 & ~n16698;
  assign n16700 = ~pi661 & ~n16699;
  assign n16701 = pi661 & n16688;
  assign n16702 = ~pi681 & ~n16701;
  assign n16703 = ~n16700 & n16702;
  assign n16704 = ~n16689 & ~n16703;
  assign n16705 = ~n6197 & ~n16704;
  assign n16706 = pi681 & ~n16694;
  assign n16707 = ~pi661 & ~pi681;
  assign n16708 = ~pi662 & n16707;
  assign n16709 = ~pi616 & ~n16708;
  assign n16710 = n16692 & n16709;
  assign n16711 = ~pi680 & n16693;
  assign n16712 = pi680 & ~n16683;
  assign n16713 = ~pi616 & n16708;
  assign n16714 = ~n16712 & n16713;
  assign n16715 = ~n16711 & n16714;
  assign n16716 = ~n16710 & ~n16715;
  assign n16717 = ~pi680 & ~n16661;
  assign n16718 = pi616 & n16708;
  assign n16719 = ~n16717 & n16718;
  assign n16720 = ~n16712 & n16719;
  assign n16721 = pi616 & n16661;
  assign n16722 = ~n16708 & n16721;
  assign n16723 = ~n16720 & ~n16722;
  assign n16724 = ~pi681 & n16723;
  assign n16725 = n16716 & n16724;
  assign n16726 = ~n16706 & ~n16725;
  assign n16727 = n6197 & ~n16726;
  assign n16728 = ~n16705 & ~n16727;
  assign n16729 = pi223 & ~n16728;
  assign n16730 = ~pi603 & ~n16661;
  assign n16731 = ~pi824 & ~n16657;
  assign n16732 = n6443 & ~n10184;
  assign n16733 = pi1092 & n16732;
  assign n16734 = ~n11009 & ~n16733;
  assign n16735 = ~n16731 & ~n16734;
  assign n16736 = pi1093 & n16735;
  assign n16737 = ~pi120 & ~n16736;
  assign n16738 = n16672 & ~n16737;
  assign n16739 = n2733 & n16663;
  assign n16740 = ~pi829 & ~n16735;
  assign n16741 = pi829 & ~n16733;
  assign n16742 = n7495 & ~n16741;
  assign n16743 = ~n16740 & n16742;
  assign n16744 = ~n16739 & ~n16743;
  assign n16745 = pi1091 & ~n16744;
  assign n16746 = ~pi120 & ~n16745;
  assign n16747 = ~n16671 & ~n16746;
  assign n16748 = ~n16738 & ~n16747;
  assign n16749 = ~n6170 & n16748;
  assign n16750 = ~n16682 & ~n16749;
  assign n16751 = pi603 & ~n16750;
  assign n16752 = ~n16730 & ~n16751;
  assign n16753 = ~pi642 & ~n16752;
  assign n16754 = ~n16680 & ~n16753;
  assign n16755 = ~pi614 & ~n16754;
  assign n16756 = ~n16691 & ~n16755;
  assign n16757 = ~pi616 & ~n16756;
  assign n16758 = ~n16690 & ~n16757;
  assign n16759 = pi681 & ~n16758;
  assign n16760 = ~pi616 & ~n16754;
  assign n16761 = ~pi614 & ~n6168;
  assign n16762 = ~n16690 & n16761;
  assign n16763 = ~n16760 & n16762;
  assign n16764 = ~pi614 & n6168;
  assign n16765 = n16750 & n16764;
  assign n16766 = ~n16763 & ~n16765;
  assign n16767 = pi680 & ~n16750;
  assign n16768 = pi614 & n16708;
  assign n16769 = ~n16717 & n16768;
  assign n16770 = ~n16767 & n16769;
  assign n16771 = pi614 & n16661;
  assign n16772 = ~n16708 & n16771;
  assign n16773 = ~n16770 & ~n16772;
  assign n16774 = ~pi681 & n16773;
  assign n16775 = n16766 & n16774;
  assign n16776 = ~n16759 & ~n16775;
  assign n16777 = n6197 & ~n16776;
  assign n16778 = n6170 & ~n16748;
  assign n16779 = ~n16662 & ~n16778;
  assign n16780 = ~n6165 & n16779;
  assign n16781 = n6165 & n16748;
  assign n16782 = ~n16780 & ~n16781;
  assign n16783 = ~n6168 & ~n16782;
  assign n16784 = n6168 & n16748;
  assign n16785 = ~n16783 & ~n16784;
  assign n16786 = ~n6197 & ~n16785;
  assign n16787 = ~n16777 & ~n16786;
  assign n16788 = ~n3053 & n16787;
  assign n16789 = n3053 & n16661;
  assign n16790 = ~pi223 & ~n16789;
  assign n16791 = ~n16788 & n16790;
  assign n16792 = ~n16729 & ~n16791;
  assign n16793 = ~pi299 & ~n16792;
  assign n16794 = n6222 & ~n16776;
  assign n16795 = ~n6222 & ~n16785;
  assign n16796 = n6217 & ~n16795;
  assign n16797 = ~n16794 & n16796;
  assign n16798 = ~n3461 & n16797;
  assign n16799 = n3461 & n16661;
  assign n16800 = ~pi215 & ~n16799;
  assign n16801 = ~n6217 & n16785;
  assign n16802 = ~n3461 & n16801;
  assign n16803 = n16800 & ~n16802;
  assign n16804 = ~n16798 & n16803;
  assign n16805 = ~n6217 & n16704;
  assign n16806 = ~n6222 & ~n16704;
  assign n16807 = n6222 & ~n16726;
  assign n16808 = n6217 & ~n16807;
  assign n16809 = ~n16806 & n16808;
  assign n16810 = ~n16805 & ~n16809;
  assign n16811 = pi215 & n16810;
  assign n16812 = ~n16804 & ~n16811;
  assign n16813 = pi299 & ~n16812;
  assign n16814 = ~n16793 & ~n16813;
  assign n16815 = pi39 & ~n16814;
  assign n16816 = ~n16656 & ~n16815;
  assign n16817 = pi761 & n16816;
  assign n16818 = pi621 & n16626;
  assign n16819 = ~pi210 & ~n16818;
  assign n16820 = pi621 & n16646;
  assign n16821 = pi210 & ~n16820;
  assign n16822 = ~n16819 & ~n16821;
  assign n16823 = pi603 & ~n16822;
  assign n16824 = n16649 & ~n16823;
  assign n16825 = pi299 & ~n16824;
  assign n16826 = ~pi198 & ~n16818;
  assign n16827 = pi198 & ~n16820;
  assign n16828 = ~n16826 & ~n16827;
  assign n16829 = pi621 & ~n16627;
  assign n16830 = ~n16628 & ~n16829;
  assign n16831 = ~pi198 & n16830;
  assign n16832 = pi621 & ~n16638;
  assign n16833 = ~n16647 & ~n16832;
  assign n16834 = pi198 & n16833;
  assign n16835 = ~n16831 & ~n16834;
  assign n16836 = ~pi603 & ~n16835;
  assign n16837 = ~n16828 & ~n16836;
  assign n16838 = ~pi299 & n16837;
  assign n16839 = ~n16825 & ~n16838;
  assign n16840 = ~pi39 & ~n16839;
  assign n16841 = pi621 & pi1091;
  assign n16842 = pi603 & ~n16841;
  assign n16843 = n16785 & ~n16842;
  assign n16844 = ~n6223 & ~n16843;
  assign n16845 = n16661 & n16841;
  assign n16846 = n6170 & ~n16845;
  assign n16847 = n16747 & n16841;
  assign n16848 = ~n6170 & ~n16847;
  assign n16849 = ~n16846 & ~n16848;
  assign n16850 = pi603 & ~n16849;
  assign n16851 = n16750 & ~n16850;
  assign n16852 = n6168 & ~n16851;
  assign n16853 = ~pi614 & ~pi642;
  assign n16854 = ~pi616 & n16853;
  assign n16855 = n16661 & ~n16842;
  assign n16856 = ~n16854 & n16855;
  assign n16857 = ~n16730 & n16854;
  assign n16858 = ~n16850 & n16857;
  assign n16859 = ~n16856 & ~n16858;
  assign n16860 = ~n6168 & n16859;
  assign n16861 = ~n16852 & ~n16860;
  assign n16862 = n6223 & ~n16861;
  assign n16863 = ~n3461 & ~n16844;
  assign n16864 = ~n16862 & n16863;
  assign n16865 = n3461 & n16855;
  assign n16866 = ~n16864 & ~n16865;
  assign n16867 = ~pi215 & ~n16866;
  assign n16868 = pi621 & n16670;
  assign n16869 = ~n6170 & ~n16868;
  assign n16870 = ~n16846 & ~n16869;
  assign n16871 = pi603 & ~n16870;
  assign n16872 = n6168 & n16683;
  assign n16873 = ~n16871 & n16872;
  assign n16874 = n16857 & ~n16871;
  assign n16875 = ~n16856 & ~n16874;
  assign n16876 = ~n6168 & ~n16875;
  assign n16877 = ~n16873 & ~n16876;
  assign n16878 = n6223 & n16877;
  assign n16879 = n2755 & ~n16842;
  assign n16880 = ~n16679 & n16879;
  assign n16881 = n6165 & ~n16670;
  assign n16882 = n16880 & ~n16881;
  assign n16883 = ~n6168 & ~n16882;
  assign n16884 = ~n16677 & n16879;
  assign n16885 = n6168 & ~n16884;
  assign n16886 = ~n16883 & ~n16885;
  assign n16887 = ~n6223 & ~n16886;
  assign n16888 = pi215 & ~n16887;
  assign n16889 = ~n16878 & n16888;
  assign n16890 = ~n16867 & ~n16889;
  assign n16891 = pi299 & ~n16890;
  assign n16892 = ~n6197 & ~n16843;
  assign n16893 = n6197 & ~n16861;
  assign n16894 = ~n3053 & ~n16892;
  assign n16895 = ~n16893 & n16894;
  assign n16896 = n3053 & n16855;
  assign n16897 = ~n16895 & ~n16896;
  assign n16898 = ~pi223 & ~n16897;
  assign n16899 = n6197 & n16877;
  assign n16900 = ~n6197 & ~n16886;
  assign n16901 = pi223 & ~n16900;
  assign n16902 = ~n16899 & n16901;
  assign n16903 = ~n16898 & ~n16902;
  assign n16904 = ~pi299 & ~n16903;
  assign n16905 = ~n16891 & ~n16904;
  assign n16906 = pi39 & n16905;
  assign n16907 = ~n16840 & ~n16906;
  assign n16908 = ~pi761 & n16907;
  assign n16909 = ~pi140 & ~n16908;
  assign n16910 = ~n16817 & n16909;
  assign n16911 = pi603 & ~n16835;
  assign n16912 = ~pi299 & ~n16911;
  assign n16913 = ~pi210 & ~n16830;
  assign n16914 = pi210 & ~n16833;
  assign n16915 = ~n16913 & ~n16914;
  assign n16916 = pi603 & n16915;
  assign n16917 = pi299 & ~n16916;
  assign n16918 = ~n16912 & ~n16917;
  assign n16919 = ~pi39 & ~n16918;
  assign n16920 = n16750 & n16842;
  assign n16921 = n6168 & n16920;
  assign n16922 = n16661 & n16842;
  assign n16923 = ~n16854 & n16922;
  assign n16924 = n16854 & n16920;
  assign n16925 = ~n16923 & ~n16924;
  assign n16926 = ~n6168 & ~n16925;
  assign n16927 = ~n16921 & ~n16926;
  assign n16928 = n6223 & n16927;
  assign n16929 = n16785 & n16842;
  assign n16930 = ~n6223 & ~n16929;
  assign n16931 = ~n3461 & ~n16928;
  assign n16932 = ~n16930 & n16931;
  assign n16933 = n2755 & n16842;
  assign n16934 = n3461 & n16660;
  assign n16935 = n16933 & n16934;
  assign n16936 = ~pi215 & ~n16935;
  assign n16937 = ~n16932 & n16936;
  assign n16938 = ~n16681 & n16922;
  assign n16939 = ~n16679 & n16922;
  assign n16940 = n16681 & n16854;
  assign n16941 = n16939 & ~n16940;
  assign n16942 = ~n6168 & n16941;
  assign n16943 = ~n16938 & ~n16942;
  assign n16944 = ~n6223 & n16679;
  assign n16945 = ~n16943 & ~n16944;
  assign n16946 = pi215 & ~n16945;
  assign n16947 = pi299 & ~n16946;
  assign n16948 = ~n16937 & n16947;
  assign n16949 = n16789 & n16842;
  assign n16950 = ~pi223 & ~n16949;
  assign n16951 = n6197 & n16927;
  assign n16952 = ~n6197 & ~n16929;
  assign n16953 = ~n3053 & ~n16951;
  assign n16954 = ~n16952 & n16953;
  assign n16955 = n16950 & ~n16954;
  assign n16956 = ~n6197 & n16679;
  assign n16957 = ~n16943 & ~n16956;
  assign n16958 = pi223 & ~n16957;
  assign n16959 = ~pi299 & ~n16958;
  assign n16960 = ~n16955 & n16959;
  assign n16961 = ~n16948 & ~n16960;
  assign n16962 = pi39 & n16961;
  assign n16963 = ~n16919 & ~n16962;
  assign n16964 = pi140 & ~pi761;
  assign n16965 = n16963 & n16964;
  assign n16966 = ~n16910 & ~n16965;
  assign n16967 = ~pi38 & ~n16966;
  assign n16968 = n2755 & n6250;
  assign n16969 = ~pi140 & ~n16968;
  assign n16970 = n6250 & n16933;
  assign n16971 = ~pi761 & n16970;
  assign n16972 = ~n16969 & ~n16971;
  assign n16973 = pi38 & ~n16972;
  assign n16974 = ~n16967 & ~n16973;
  assign n16975 = pi738 & ~n16974;
  assign n16976 = pi680 & ~n16708;
  assign n16977 = pi665 & pi1091;
  assign n16978 = ~n16842 & ~n16977;
  assign n16979 = n16661 & ~n16978;
  assign n16980 = pi616 & ~n16979;
  assign n16981 = pi614 & ~n16979;
  assign n16982 = pi642 & ~n16979;
  assign n16983 = pi665 & n16670;
  assign n16984 = ~n16677 & n16922;
  assign n16985 = ~n16983 & ~n16984;
  assign n16986 = n16662 & n16977;
  assign n16987 = ~pi603 & n16986;
  assign n16988 = n16985 & ~n16987;
  assign n16989 = n16661 & n16977;
  assign n16990 = n6170 & ~n16989;
  assign n16991 = ~n6170 & ~n16983;
  assign n16992 = ~n16990 & ~n16991;
  assign n16993 = ~pi642 & ~n16938;
  assign n16994 = ~n16992 & n16993;
  assign n16995 = n16988 & n16994;
  assign n16996 = ~n16982 & ~n16995;
  assign n16997 = ~pi614 & ~n16996;
  assign n16998 = ~n16981 & ~n16997;
  assign n16999 = ~pi616 & ~n16998;
  assign n17000 = ~n16980 & ~n16999;
  assign n17001 = n16976 & ~n17000;
  assign n17002 = ~pi680 & ~n16694;
  assign n17003 = n6168 & ~n16992;
  assign n17004 = ~n16938 & n17003;
  assign n17005 = ~n17002 & ~n17004;
  assign n17006 = ~n17001 & n17005;
  assign n17007 = n6197 & ~n17006;
  assign n17008 = ~pi680 & ~n16688;
  assign n17009 = n6168 & n16985;
  assign n17010 = ~n16983 & ~n16986;
  assign n17011 = ~n16939 & n17010;
  assign n17012 = n16854 & n16988;
  assign n17013 = ~n17011 & ~n17012;
  assign n17014 = n16976 & ~n17013;
  assign n17015 = ~n17009 & ~n17014;
  assign n17016 = ~n17008 & n17015;
  assign n17017 = ~n6197 & ~n17016;
  assign n17018 = pi223 & ~n17017;
  assign n17019 = ~n17007 & n17018;
  assign n17020 = n16752 & ~n16978;
  assign n17021 = ~pi642 & ~n17020;
  assign n17022 = ~n16982 & ~n17021;
  assign n17023 = ~pi614 & ~n17022;
  assign n17024 = ~n16981 & ~n17023;
  assign n17025 = ~pi616 & ~n17024;
  assign n17026 = ~n16980 & ~n17025;
  assign n17027 = n16976 & ~n17026;
  assign n17028 = ~pi680 & ~n16758;
  assign n17029 = n16747 & n16977;
  assign n17030 = ~n6170 & ~n17029;
  assign n17031 = ~n16990 & ~n17030;
  assign n17032 = ~pi603 & ~n17031;
  assign n17033 = pi603 & n16978;
  assign n17034 = ~n16751 & ~n17033;
  assign n17035 = ~n17032 & n17034;
  assign n17036 = n6168 & ~n17035;
  assign n17037 = ~n17028 & ~n17036;
  assign n17038 = ~n17027 & n17037;
  assign n17039 = n6197 & n17038;
  assign n17040 = n16782 & ~n16978;
  assign n17041 = n16976 & ~n17040;
  assign n17042 = ~pi680 & ~n16782;
  assign n17043 = ~n16748 & ~n16841;
  assign n17044 = pi603 & n17043;
  assign n17045 = pi603 & ~pi621;
  assign n17046 = n17029 & ~n17045;
  assign n17047 = n6168 & ~n17046;
  assign n17048 = ~n17044 & n17047;
  assign n17049 = ~n17042 & ~n17048;
  assign n17050 = ~n17041 & n17049;
  assign n17051 = ~n6197 & n17050;
  assign n17052 = ~n3053 & ~n17051;
  assign n17053 = ~n17039 & n17052;
  assign n17054 = pi680 & n16978;
  assign n17055 = n16661 & ~n17054;
  assign n17056 = n3053 & ~n17055;
  assign n17057 = ~pi223 & ~n17056;
  assign n17058 = ~n17053 & n17057;
  assign n17059 = ~n17019 & ~n17058;
  assign n17060 = ~pi299 & ~n17059;
  assign n17061 = ~n6223 & ~n17050;
  assign n17062 = n6223 & ~n17038;
  assign n17063 = ~n17061 & ~n17062;
  assign n17064 = ~n3461 & ~n17063;
  assign n17065 = n3461 & ~n17055;
  assign n17066 = ~pi215 & ~n17065;
  assign n17067 = ~n17064 & n17066;
  assign n17068 = n6223 & ~n17006;
  assign n17069 = ~n6223 & ~n17016;
  assign n17070 = pi215 & ~n17069;
  assign n17071 = ~n17068 & n17070;
  assign n17072 = ~n17067 & ~n17071;
  assign n17073 = pi299 & ~n17072;
  assign n17074 = ~n17060 & ~n17073;
  assign n17075 = ~pi140 & n17074;
  assign n17076 = n16661 & ~n16977;
  assign n17077 = ~n16748 & ~n16977;
  assign n17078 = ~n17076 & ~n17077;
  assign n17079 = ~pi603 & n16779;
  assign n17080 = n6170 & n16847;
  assign n17081 = n16662 & n16841;
  assign n17082 = pi603 & ~n17081;
  assign n17083 = ~n17080 & n17082;
  assign n17084 = ~n17079 & ~n17083;
  assign n17085 = ~n17078 & n17084;
  assign n17086 = pi616 & ~n17085;
  assign n17087 = ~pi665 & n16847;
  assign n17088 = pi603 & ~n17087;
  assign n17089 = ~n16779 & ~n17078;
  assign n17090 = ~pi603 & ~n17089;
  assign n17091 = ~n17088 & ~n17090;
  assign n17092 = n16854 & ~n17091;
  assign n17093 = n17085 & ~n17092;
  assign n17094 = n16853 & n17091;
  assign n17095 = ~pi616 & ~n17094;
  assign n17096 = ~n17093 & n17095;
  assign n17097 = ~n17086 & ~n17096;
  assign n17098 = ~n16708 & ~n17097;
  assign n17099 = n6168 & n17077;
  assign n17100 = ~n17088 & n17099;
  assign n17101 = ~n16976 & ~n17100;
  assign n17102 = ~n17098 & ~n17101;
  assign n17103 = ~n6223 & ~n17102;
  assign n17104 = n16855 & ~n16977;
  assign n17105 = pi616 & ~n17104;
  assign n17106 = n16976 & ~n17105;
  assign n17107 = pi603 & pi665;
  assign n17108 = ~pi603 & ~n17076;
  assign n17109 = ~n17107 & ~n17108;
  assign n17110 = ~n16850 & n17109;
  assign n17111 = n16853 & n17110;
  assign n17112 = ~n16853 & n17104;
  assign n17113 = ~pi616 & ~n17112;
  assign n17114 = ~n17111 & n17113;
  assign n17115 = n17106 & ~n17114;
  assign n17116 = n16750 & n17036;
  assign n17117 = ~n17115 & ~n17116;
  assign n17118 = n6223 & n17117;
  assign n17119 = ~n3461 & ~n17118;
  assign n17120 = ~n17103 & n17119;
  assign n17121 = ~n16800 & ~n17066;
  assign n17122 = ~n17120 & ~n17121;
  assign n17123 = n16880 & n17109;
  assign n17124 = pi616 & ~n17123;
  assign n17125 = pi614 & ~pi616;
  assign n17126 = ~n17123 & n17125;
  assign n17127 = ~n16871 & n17109;
  assign n17128 = ~pi642 & ~n17127;
  assign n17129 = n17123 & ~n17128;
  assign n17130 = n6164 & ~n17129;
  assign n17131 = ~n17126 & ~n17130;
  assign n17132 = ~n17124 & n17131;
  assign n17133 = ~n16708 & ~n17132;
  assign n17134 = ~n16677 & n17054;
  assign n17135 = ~n16976 & ~n17134;
  assign n17136 = ~n17133 & ~n17135;
  assign n17137 = ~n6223 & n17136;
  assign n17138 = ~n16875 & ~n16977;
  assign n17139 = ~pi616 & ~n17138;
  assign n17140 = n17106 & ~n17139;
  assign n17141 = n16873 & n17109;
  assign n17142 = ~n17140 & ~n17141;
  assign n17143 = n6223 & ~n17142;
  assign n17144 = pi215 & ~n17143;
  assign n17145 = ~n17137 & n17144;
  assign n17146 = ~n17122 & ~n17145;
  assign n17147 = pi299 & ~n17146;
  assign n17148 = ~n6197 & n17102;
  assign n17149 = n6197 & ~n17117;
  assign n17150 = ~n3053 & ~n17149;
  assign n17151 = ~n17148 & n17150;
  assign n17152 = pi680 & ~n16977;
  assign n17153 = n2755 & n17152;
  assign n17154 = ~n16842 & n17153;
  assign n17155 = ~n16933 & ~n17154;
  assign n17156 = n16661 & ~n17155;
  assign n17157 = n3053 & ~n17156;
  assign n17158 = n16950 & ~n17157;
  assign n17159 = ~n17151 & n17158;
  assign n17160 = ~n6197 & ~n17136;
  assign n17161 = n6197 & n17142;
  assign n17162 = pi223 & ~n17161;
  assign n17163 = ~n17160 & n17162;
  assign n17164 = ~pi299 & ~n17163;
  assign n17165 = ~n17159 & n17164;
  assign n17166 = ~n17147 & ~n17165;
  assign n17167 = pi140 & n17166;
  assign n17168 = pi761 & ~n17167;
  assign n17169 = ~n17075 & n17168;
  assign n17170 = ~n17044 & ~n17091;
  assign n17171 = n16854 & ~n17170;
  assign n17172 = ~n16779 & n16842;
  assign n17173 = ~n17089 & ~n17172;
  assign n17174 = ~n16854 & ~n17173;
  assign n17175 = n16976 & ~n17174;
  assign n17176 = ~n17171 & n17175;
  assign n17177 = ~n16976 & ~n17099;
  assign n17178 = ~n16929 & n17177;
  assign n17179 = ~n17176 & ~n17178;
  assign n17180 = ~n6197 & n17179;
  assign n17181 = n16977 & ~n17045;
  assign n17182 = n16661 & ~n17181;
  assign n17183 = ~n16854 & n17182;
  assign n17184 = n16976 & ~n17183;
  assign n17185 = ~n16920 & ~n17110;
  assign n17186 = n16854 & ~n17185;
  assign n17187 = n17184 & ~n17186;
  assign n17188 = ~pi680 & n16925;
  assign n17189 = n16750 & ~n17078;
  assign n17190 = n6168 & ~n16920;
  assign n17191 = ~n17189 & n17190;
  assign n17192 = ~n17188 & ~n17191;
  assign n17193 = ~n17187 & n17192;
  assign n17194 = n6197 & n17193;
  assign n17195 = ~n3053 & ~n17194;
  assign n17196 = ~n17180 & n17195;
  assign n17197 = ~pi223 & ~n17157;
  assign n17198 = ~n17196 & n17197;
  assign n17199 = ~n6165 & n17076;
  assign n17200 = ~n16681 & n17076;
  assign n17201 = ~n17199 & ~n17200;
  assign n17202 = ~n16938 & n17201;
  assign n17203 = n16854 & ~n17202;
  assign n17204 = n17184 & ~n17203;
  assign n17205 = n16708 & ~n17200;
  assign n17206 = pi680 & ~n17205;
  assign n17207 = n16943 & ~n17206;
  assign n17208 = ~n17204 & ~n17207;
  assign n17209 = n6197 & ~n17208;
  assign n17210 = ~n16942 & ~n16984;
  assign n17211 = ~n16679 & n17076;
  assign n17212 = ~n17201 & n17206;
  assign n17213 = n17211 & n17212;
  assign n17214 = n17210 & ~n17213;
  assign n17215 = ~n6197 & n17214;
  assign n17216 = pi223 & ~n17215;
  assign n17217 = ~n17209 & n17216;
  assign n17218 = ~pi299 & ~n17217;
  assign n17219 = ~n17198 & n17218;
  assign n17220 = ~n6223 & n17179;
  assign n17221 = n6223 & n17193;
  assign n17222 = ~n17220 & ~n17221;
  assign n17223 = ~n3461 & ~n17222;
  assign n17224 = n3461 & n17156;
  assign n17225 = ~pi215 & ~n17224;
  assign n17226 = ~n17223 & n17225;
  assign n17227 = n6223 & n17208;
  assign n17228 = ~n6223 & ~n17214;
  assign n17229 = pi215 & ~n17228;
  assign n17230 = ~n17227 & n17229;
  assign n17231 = ~n17226 & ~n17230;
  assign n17232 = pi299 & ~n17231;
  assign n17233 = ~n17219 & ~n17232;
  assign n17234 = pi140 & n17233;
  assign n17235 = n16782 & ~n16842;
  assign n17236 = ~pi680 & ~n17235;
  assign n17237 = ~n6199 & n17029;
  assign n17238 = ~n6165 & n16986;
  assign n17239 = ~n17237 & ~n17238;
  assign n17240 = n17181 & ~n17239;
  assign n17241 = n16976 & ~n17240;
  assign n17242 = ~n17047 & ~n17241;
  assign n17243 = ~n17236 & n17242;
  assign n17244 = ~n6197 & n17243;
  assign n17245 = ~pi680 & n16859;
  assign n17246 = n16858 & n16977;
  assign n17247 = n16989 & ~n17045;
  assign n17248 = ~n16854 & n17247;
  assign n17249 = n16976 & ~n17248;
  assign n17250 = ~n17246 & n17249;
  assign n17251 = n17031 & n17181;
  assign n17252 = n6168 & ~n17251;
  assign n17253 = ~n17245 & ~n17252;
  assign n17254 = ~n17250 & n17253;
  assign n17255 = n6197 & n17254;
  assign n17256 = ~n17244 & ~n17255;
  assign n17257 = ~n3053 & ~n17256;
  assign n17258 = ~n16842 & ~n17152;
  assign n17259 = n16665 & n17258;
  assign n17260 = ~n16658 & n17259;
  assign n17261 = n3053 & n17260;
  assign n17262 = ~pi223 & ~n17261;
  assign n17263 = ~n17257 & n17262;
  assign n17264 = n16876 & ~n17152;
  assign n17265 = n6168 & ~n17045;
  assign n17266 = n16992 & n17265;
  assign n17267 = ~n17264 & ~n17266;
  assign n17268 = n6197 & ~n17267;
  assign n17269 = ~n16875 & ~n17010;
  assign n17270 = n16976 & ~n17269;
  assign n17271 = ~pi680 & ~n16882;
  assign n17272 = pi680 & ~n16983;
  assign n17273 = ~n17045 & ~n17272;
  assign n17274 = n6168 & ~n17273;
  assign n17275 = ~n17271 & ~n17274;
  assign n17276 = ~n17270 & n17275;
  assign n17277 = ~n6197 & n17276;
  assign n17278 = pi223 & ~n17268;
  assign n17279 = ~n17277 & n17278;
  assign n17280 = ~n17263 & ~n17279;
  assign n17281 = ~pi299 & ~n17280;
  assign n17282 = ~n6223 & n17243;
  assign n17283 = n6223 & n17254;
  assign n17284 = ~n17282 & ~n17283;
  assign n17285 = ~n3461 & ~n17284;
  assign n17286 = n3461 & n17260;
  assign n17287 = ~pi215 & ~n17286;
  assign n17288 = ~n17285 & n17287;
  assign n17289 = n6223 & ~n17267;
  assign n17290 = ~n6223 & n17276;
  assign n17291 = pi215 & ~n17289;
  assign n17292 = ~n17290 & n17291;
  assign n17293 = ~n17288 & ~n17292;
  assign n17294 = pi299 & ~n17293;
  assign n17295 = ~n17281 & ~n17294;
  assign n17296 = ~pi140 & ~n17295;
  assign n17297 = ~pi761 & ~n17296;
  assign n17298 = ~n17234 & n17297;
  assign n17299 = ~n17169 & ~n17298;
  assign n17300 = pi39 & ~n17299;
  assign n17301 = pi665 & n16646;
  assign n17302 = pi198 & ~n17301;
  assign n17303 = pi665 & n16626;
  assign n17304 = ~pi198 & ~n17303;
  assign n17305 = ~n17302 & ~n17304;
  assign n17306 = pi680 & ~n17305;
  assign n17307 = n16653 & ~n17306;
  assign n17308 = ~pi299 & ~n17307;
  assign n17309 = ~pi210 & ~n17303;
  assign n17310 = pi210 & ~n17301;
  assign n17311 = ~n17309 & ~n17310;
  assign n17312 = pi680 & ~n17311;
  assign n17313 = n16649 & ~n17312;
  assign n17314 = pi299 & ~n17313;
  assign n17315 = ~n17308 & ~n17314;
  assign n17316 = pi680 & n16918;
  assign n17317 = ~n17315 & ~n17316;
  assign n17318 = ~pi140 & ~n17317;
  assign n17319 = pi665 & ~n16627;
  assign n17320 = ~n16628 & ~n17319;
  assign n17321 = ~pi198 & ~n17320;
  assign n17322 = pi665 & ~n16638;
  assign n17323 = ~n16647 & ~n17322;
  assign n17324 = pi198 & ~n17323;
  assign n17325 = ~n17321 & ~n17324;
  assign n17326 = ~pi603 & ~n17325;
  assign n17327 = pi603 & ~n16828;
  assign n17328 = ~n17107 & ~n17327;
  assign n17329 = ~n17326 & n17328;
  assign n17330 = pi680 & n17329;
  assign n17331 = ~pi299 & ~n17330;
  assign n17332 = pi210 & ~n17323;
  assign n17333 = ~pi210 & ~n17320;
  assign n17334 = ~n17332 & ~n17333;
  assign n17335 = ~pi603 & ~n17334;
  assign n17336 = ~n16823 & ~n17107;
  assign n17337 = ~n17335 & n17336;
  assign n17338 = pi680 & n17337;
  assign n17339 = pi299 & ~n17338;
  assign n17340 = ~n17331 & ~n17339;
  assign n17341 = pi140 & ~n17340;
  assign n17342 = pi761 & ~n17318;
  assign n17343 = ~n17341 & n17342;
  assign n17344 = n16839 & n17315;
  assign n17345 = ~pi140 & n17344;
  assign n17346 = pi680 & n17325;
  assign n17347 = ~pi299 & ~n17346;
  assign n17348 = pi680 & n17334;
  assign n17349 = pi299 & ~n17348;
  assign n17350 = ~n17347 & ~n17349;
  assign n17351 = ~n16918 & ~n17350;
  assign n17352 = pi140 & n17351;
  assign n17353 = ~pi761 & ~n17352;
  assign n17354 = ~n17345 & n17353;
  assign n17355 = ~pi39 & ~n17354;
  assign n17356 = ~n17343 & n17355;
  assign n17357 = ~pi38 & ~n17356;
  assign n17358 = ~n17300 & n17357;
  assign n17359 = ~pi140 & ~n17259;
  assign n17360 = pi140 & ~n17155;
  assign n17361 = n3096 & n17360;
  assign n17362 = ~pi761 & ~n17361;
  assign n17363 = ~n17359 & n17362;
  assign n17364 = ~pi140 & ~n16665;
  assign n17365 = n16665 & n17054;
  assign n17366 = pi761 & ~n17364;
  assign n17367 = ~n17365 & n17366;
  assign n17368 = ~n17363 & ~n17367;
  assign n17369 = ~pi39 & ~n17368;
  assign n17370 = pi39 & pi140;
  assign n17371 = pi38 & ~n17370;
  assign n17372 = ~n17369 & n17371;
  assign n17373 = ~n17358 & ~n17372;
  assign n17374 = ~pi738 & ~n17373;
  assign n17375 = n3268 & ~n16975;
  assign n17376 = ~n17374 & n17375;
  assign n17377 = ~n16578 & ~n17376;
  assign n17378 = ~pi625 & n17377;
  assign n17379 = n3268 & n16974;
  assign n17380 = ~n16578 & ~n17379;
  assign n17381 = pi625 & n17380;
  assign n17382 = ~pi1153 & ~n17381;
  assign n17383 = ~n17378 & n17382;
  assign n17384 = n16789 & n17152;
  assign n17385 = n6165 & n17189;
  assign n17386 = ~n17199 & ~n17385;
  assign n17387 = ~n16708 & n17386;
  assign n17388 = n16708 & ~n17189;
  assign n17389 = pi680 & ~n17388;
  assign n17390 = ~n17387 & n17389;
  assign n17391 = n6197 & ~n17390;
  assign n17392 = n16782 & n17152;
  assign n17393 = ~n16708 & n17392;
  assign n17394 = ~n17099 & ~n17393;
  assign n17395 = ~n6197 & n17394;
  assign n17396 = ~n3053 & ~n17391;
  assign n17397 = ~n17395 & n17396;
  assign n17398 = ~n17384 & ~n17397;
  assign n17399 = ~pi223 & ~n17398;
  assign n17400 = pi680 & ~n17201;
  assign n17401 = ~n16956 & n17400;
  assign n17402 = pi223 & ~n17205;
  assign n17403 = n17401 & n17402;
  assign n17404 = ~n17399 & ~n17403;
  assign n17405 = ~pi299 & ~n17404;
  assign n17406 = ~n6223 & n17394;
  assign n17407 = n6223 & ~n17390;
  assign n17408 = ~n3461 & ~n17406;
  assign n17409 = ~n17407 & n17408;
  assign n17410 = n16661 & n17152;
  assign n17411 = n3461 & n17410;
  assign n17412 = ~n17409 & ~n17411;
  assign n17413 = ~pi215 & ~n17412;
  assign n17414 = ~n16944 & n17400;
  assign n17415 = pi215 & ~n17205;
  assign n17416 = n17414 & n17415;
  assign n17417 = ~n17413 & ~n17416;
  assign n17418 = pi299 & ~n17417;
  assign n17419 = ~n17405 & ~n17418;
  assign n17420 = pi140 & ~n17419;
  assign n17421 = n6165 & n17031;
  assign n17422 = ~n6165 & n16989;
  assign n17423 = pi680 & ~n17422;
  assign n17424 = ~n17421 & n17423;
  assign n17425 = ~n17028 & ~n17424;
  assign n17426 = ~n16708 & n17425;
  assign n17427 = pi680 & ~n17031;
  assign n17428 = n16708 & ~n17427;
  assign n17429 = ~n17028 & n17428;
  assign n17430 = ~n17426 & ~n17429;
  assign n17431 = n6197 & n17430;
  assign n17432 = ~n16708 & ~n17239;
  assign n17433 = n16708 & n17029;
  assign n17434 = pi680 & ~n17433;
  assign n17435 = ~n17432 & n17434;
  assign n17436 = ~n17042 & ~n17435;
  assign n17437 = ~n6197 & ~n17436;
  assign n17438 = ~n3053 & ~n17437;
  assign n17439 = ~n17431 & n17438;
  assign n17440 = n16789 & ~n17152;
  assign n17441 = ~pi223 & ~n17440;
  assign n17442 = ~n17439 & n17441;
  assign n17443 = ~n16992 & n17423;
  assign n17444 = ~n17003 & ~n17443;
  assign n17445 = ~n17002 & n17444;
  assign n17446 = n6197 & n17445;
  assign n17447 = ~n17238 & n17272;
  assign n17448 = ~n17008 & ~n17447;
  assign n17449 = n17444 & n17448;
  assign n17450 = ~n6197 & n17449;
  assign n17451 = pi223 & ~n17446;
  assign n17452 = ~n17450 & n17451;
  assign n17453 = ~n17442 & ~n17452;
  assign n17454 = ~pi299 & ~n17453;
  assign n17455 = n6223 & n17430;
  assign n17456 = ~n6223 & ~n17436;
  assign n17457 = ~n3461 & ~n17456;
  assign n17458 = ~n17455 & n17457;
  assign n17459 = n2755 & ~n17152;
  assign n17460 = n16934 & n17459;
  assign n17461 = ~pi215 & ~n17460;
  assign n17462 = ~n17458 & n17461;
  assign n17463 = n6223 & n17445;
  assign n17464 = ~n6223 & n17449;
  assign n17465 = pi215 & ~n17463;
  assign n17466 = ~n17464 & n17465;
  assign n17467 = ~n17462 & ~n17466;
  assign n17468 = pi299 & ~n17467;
  assign n17469 = ~n17454 & ~n17468;
  assign n17470 = pi39 & n17469;
  assign n17471 = ~n17370 & ~n17470;
  assign n17472 = ~n17420 & ~n17471;
  assign n17473 = pi140 & n17350;
  assign n17474 = ~pi140 & ~n17315;
  assign n17475 = ~pi39 & ~n17473;
  assign n17476 = ~n17474 & n17475;
  assign n17477 = ~n17472 & ~n17476;
  assign n17478 = ~pi38 & ~n17477;
  assign n17479 = n6250 & n17153;
  assign n17480 = pi38 & ~n17479;
  assign n17481 = ~n16969 & n17480;
  assign n17482 = ~pi738 & ~n17481;
  assign n17483 = ~n17478 & n17482;
  assign n17484 = ~pi38 & ~n16816;
  assign n17485 = n2755 & n6117;
  assign n17486 = pi38 & ~n17485;
  assign n17487 = ~n17484 & ~n17486;
  assign n17488 = ~pi140 & pi738;
  assign n17489 = ~n17487 & n17488;
  assign n17490 = n3268 & ~n17489;
  assign n17491 = ~n17483 & n17490;
  assign n17492 = ~n16578 & ~n17491;
  assign n17493 = pi625 & n17492;
  assign n17494 = n3268 & n17487;
  assign n17495 = ~pi140 & ~n17494;
  assign n17496 = ~pi625 & n17495;
  assign n17497 = pi1153 & ~n17496;
  assign n17498 = ~n17493 & n17497;
  assign n17499 = ~pi608 & ~n17498;
  assign n17500 = ~n17383 & n17499;
  assign n17501 = pi625 & n17377;
  assign n17502 = ~pi625 & n17380;
  assign n17503 = pi1153 & ~n17502;
  assign n17504 = ~n17501 & n17503;
  assign n17505 = ~pi625 & n17492;
  assign n17506 = pi625 & n17495;
  assign n17507 = ~pi1153 & ~n17506;
  assign n17508 = ~n17505 & n17507;
  assign n17509 = pi608 & ~n17508;
  assign n17510 = ~n17504 & n17509;
  assign n17511 = ~n17500 & ~n17510;
  assign n17512 = pi778 & ~n17511;
  assign n17513 = ~pi778 & n17377;
  assign n17514 = ~n17512 & ~n17513;
  assign n17515 = ~pi609 & ~n17514;
  assign n17516 = ~pi778 & ~n17492;
  assign n17517 = ~n17498 & ~n17508;
  assign n17518 = pi778 & ~n17517;
  assign n17519 = ~n17516 & ~n17518;
  assign n17520 = pi609 & n17519;
  assign n17521 = ~pi1155 & ~n17520;
  assign n17522 = ~n17515 & n17521;
  assign n17523 = ~pi608 & pi1153;
  assign n17524 = pi608 & ~pi1153;
  assign n17525 = ~n17523 & ~n17524;
  assign n17526 = pi778 & ~n17525;
  assign n17527 = pi609 & ~n17526;
  assign n17528 = ~n17495 & ~n17527;
  assign n17529 = ~n17380 & ~n17526;
  assign n17530 = pi609 & n17529;
  assign n17531 = ~n17528 & ~n17530;
  assign n17532 = pi1155 & ~n17531;
  assign n17533 = ~pi660 & ~n17532;
  assign n17534 = ~n17522 & n17533;
  assign n17535 = pi609 & ~n17514;
  assign n17536 = ~pi609 & n17519;
  assign n17537 = pi1155 & ~n17536;
  assign n17538 = ~n17535 & n17537;
  assign n17539 = ~pi609 & ~n17526;
  assign n17540 = ~n17495 & ~n17539;
  assign n17541 = ~pi609 & n17529;
  assign n17542 = ~n17540 & ~n17541;
  assign n17543 = ~pi1155 & ~n17542;
  assign n17544 = pi660 & ~n17543;
  assign n17545 = ~n17538 & n17544;
  assign n17546 = ~n17534 & ~n17545;
  assign n17547 = pi785 & ~n17546;
  assign n17548 = ~pi785 & ~n17514;
  assign n17549 = ~n17547 & ~n17548;
  assign n17550 = ~pi618 & ~n17549;
  assign n17551 = pi660 & pi1155;
  assign n17552 = ~pi660 & ~pi1155;
  assign n17553 = pi785 & ~n17551;
  assign n17554 = ~n17552 & n17553;
  assign n17555 = ~n17519 & ~n17554;
  assign n17556 = ~n17495 & n17554;
  assign n17557 = ~n17555 & ~n17556;
  assign n17558 = pi618 & n17557;
  assign n17559 = ~pi1154 & ~n17558;
  assign n17560 = ~n17550 & n17559;
  assign n17561 = ~n17495 & n17526;
  assign n17562 = ~n17529 & ~n17561;
  assign n17563 = ~pi785 & ~n17562;
  assign n17564 = ~n17532 & ~n17543;
  assign n17565 = pi785 & ~n17564;
  assign n17566 = ~n17563 & ~n17565;
  assign n17567 = pi618 & n17566;
  assign n17568 = ~pi618 & n17495;
  assign n17569 = pi1154 & ~n17568;
  assign n17570 = ~n17567 & n17569;
  assign n17571 = ~pi627 & ~n17570;
  assign n17572 = ~n17560 & n17571;
  assign n17573 = pi618 & ~n17549;
  assign n17574 = ~pi618 & n17557;
  assign n17575 = pi1154 & ~n17574;
  assign n17576 = ~n17573 & n17575;
  assign n17577 = ~pi618 & n17566;
  assign n17578 = pi618 & n17495;
  assign n17579 = ~pi1154 & ~n17578;
  assign n17580 = ~n17577 & n17579;
  assign n17581 = pi627 & ~n17580;
  assign n17582 = ~n17576 & n17581;
  assign n17583 = ~n17572 & ~n17582;
  assign n17584 = pi781 & ~n17583;
  assign n17585 = ~pi781 & ~n17549;
  assign n17586 = ~n17584 & ~n17585;
  assign n17587 = ~pi619 & ~n17586;
  assign n17588 = pi627 & pi1154;
  assign n17589 = ~pi627 & ~pi1154;
  assign n17590 = pi781 & ~n17588;
  assign n17591 = ~n17589 & n17590;
  assign n17592 = n17557 & ~n17591;
  assign n17593 = n17495 & n17591;
  assign n17594 = ~n17592 & ~n17593;
  assign n17595 = pi619 & ~n17594;
  assign n17596 = ~pi1159 & ~n17595;
  assign n17597 = ~n17587 & n17596;
  assign n17598 = ~pi781 & ~n17566;
  assign n17599 = ~n17570 & ~n17580;
  assign n17600 = pi781 & ~n17599;
  assign n17601 = ~n17598 & ~n17600;
  assign n17602 = pi619 & n17601;
  assign n17603 = ~pi619 & n17495;
  assign n17604 = pi1159 & ~n17603;
  assign n17605 = ~n17602 & n17604;
  assign n17606 = ~pi648 & ~n17605;
  assign n17607 = ~n17597 & n17606;
  assign n17608 = pi619 & ~n17586;
  assign n17609 = ~pi619 & ~n17594;
  assign n17610 = pi1159 & ~n17609;
  assign n17611 = ~n17608 & n17610;
  assign n17612 = ~pi619 & n17601;
  assign n17613 = pi619 & n17495;
  assign n17614 = ~pi1159 & ~n17613;
  assign n17615 = ~n17612 & n17614;
  assign n17616 = pi648 & ~n17615;
  assign n17617 = ~n17611 & n17616;
  assign n17618 = ~n17607 & ~n17617;
  assign n17619 = pi789 & ~n17618;
  assign n17620 = ~pi789 & ~n17586;
  assign n17621 = ~n17619 & ~n17620;
  assign n17622 = ~pi788 & n17621;
  assign n17623 = ~pi626 & n17621;
  assign n17624 = ~pi648 & pi1159;
  assign n17625 = pi648 & ~pi1159;
  assign n17626 = ~n17624 & ~n17625;
  assign n17627 = pi789 & ~n17626;
  assign n17628 = n17594 & ~n17627;
  assign n17629 = ~n17495 & n17627;
  assign n17630 = ~n17628 & ~n17629;
  assign n17631 = pi626 & ~n17630;
  assign n17632 = ~pi641 & ~n17631;
  assign n17633 = ~n17623 & n17632;
  assign n17634 = ~pi641 & ~pi1158;
  assign n17635 = ~pi789 & ~n17601;
  assign n17636 = ~n17605 & ~n17615;
  assign n17637 = pi789 & ~n17636;
  assign n17638 = ~n17635 & ~n17637;
  assign n17639 = ~pi626 & n17638;
  assign n17640 = pi626 & n17495;
  assign n17641 = ~pi1158 & ~n17640;
  assign n17642 = ~n17639 & n17641;
  assign n17643 = ~n17634 & ~n17642;
  assign n17644 = ~n17633 & ~n17643;
  assign n17645 = pi626 & n17621;
  assign n17646 = ~pi626 & ~n17630;
  assign n17647 = pi641 & ~n17646;
  assign n17648 = ~n17645 & n17647;
  assign n17649 = pi641 & pi1158;
  assign n17650 = pi626 & n17638;
  assign n17651 = ~pi626 & n17495;
  assign n17652 = pi1158 & ~n17651;
  assign n17653 = ~n17650 & n17652;
  assign n17654 = ~n17649 & ~n17653;
  assign n17655 = ~n17648 & ~n17654;
  assign n17656 = ~n17644 & ~n17655;
  assign n17657 = pi788 & ~n17656;
  assign n17658 = ~n17622 & ~n17657;
  assign n17659 = ~pi628 & n17658;
  assign n17660 = ~n17642 & ~n17653;
  assign n17661 = pi788 & ~n17660;
  assign n17662 = ~pi788 & ~n17638;
  assign n17663 = ~n17661 & ~n17662;
  assign n17664 = pi628 & n17663;
  assign n17665 = ~pi1156 & ~n17664;
  assign n17666 = ~n17659 & n17665;
  assign n17667 = ~pi641 & pi1158;
  assign n17668 = pi641 & ~pi1158;
  assign n17669 = ~n17667 & ~n17668;
  assign n17670 = pi788 & ~n17669;
  assign n17671 = n17630 & ~n17670;
  assign n17672 = n17495 & n17670;
  assign n17673 = ~n17671 & ~n17672;
  assign n17674 = pi628 & ~n17673;
  assign n17675 = ~pi628 & n17495;
  assign n17676 = pi1156 & ~n17675;
  assign n17677 = ~n17674 & n17676;
  assign n17678 = ~pi629 & ~n17677;
  assign n17679 = ~n17666 & n17678;
  assign n17680 = pi628 & n17658;
  assign n17681 = ~pi628 & n17663;
  assign n17682 = pi1156 & ~n17681;
  assign n17683 = ~n17680 & n17682;
  assign n17684 = ~pi628 & ~n17673;
  assign n17685 = pi628 & n17495;
  assign n17686 = ~pi1156 & ~n17685;
  assign n17687 = ~n17684 & n17686;
  assign n17688 = pi629 & ~n17687;
  assign n17689 = ~n17683 & n17688;
  assign n17690 = ~n17679 & ~n17689;
  assign n17691 = pi792 & ~n17690;
  assign n17692 = ~pi792 & n17658;
  assign n17693 = ~n17691 & ~n17692;
  assign n17694 = ~pi647 & ~n17693;
  assign n17695 = ~pi629 & pi1156;
  assign n17696 = pi629 & ~pi1156;
  assign n17697 = ~n17695 & ~n17696;
  assign n17698 = pi792 & ~n17697;
  assign n17699 = n17663 & ~n17698;
  assign n17700 = n17495 & n17698;
  assign n17701 = ~n17699 & ~n17700;
  assign n17702 = pi647 & ~n17701;
  assign n17703 = ~pi1157 & ~n17702;
  assign n17704 = ~n17694 & n17703;
  assign n17705 = ~pi792 & n17673;
  assign n17706 = ~n17677 & ~n17687;
  assign n17707 = pi792 & ~n17706;
  assign n17708 = ~n17705 & ~n17707;
  assign n17709 = pi647 & n17708;
  assign n17710 = ~pi647 & n17495;
  assign n17711 = pi1157 & ~n17710;
  assign n17712 = ~n17709 & n17711;
  assign n17713 = ~pi630 & ~n17712;
  assign n17714 = ~n17704 & n17713;
  assign n17715 = pi647 & ~n17693;
  assign n17716 = ~pi647 & ~n17701;
  assign n17717 = pi1157 & ~n17716;
  assign n17718 = ~n17715 & n17717;
  assign n17719 = ~pi647 & n17708;
  assign n17720 = pi647 & n17495;
  assign n17721 = ~pi1157 & ~n17720;
  assign n17722 = ~n17719 & n17721;
  assign n17723 = pi630 & ~n17722;
  assign n17724 = ~n17718 & n17723;
  assign n17725 = ~n17714 & ~n17724;
  assign n17726 = pi787 & ~n17725;
  assign n17727 = ~pi787 & ~n17693;
  assign n17728 = ~n17726 & ~n17727;
  assign n17729 = pi644 & ~n17728;
  assign n17730 = ~pi787 & ~n17708;
  assign n17731 = ~n17712 & ~n17722;
  assign n17732 = pi787 & ~n17731;
  assign n17733 = ~n17730 & ~n17732;
  assign n17734 = ~pi644 & n17733;
  assign n17735 = pi715 & ~n17734;
  assign n17736 = ~n17729 & n17735;
  assign n17737 = ~pi630 & pi1157;
  assign n17738 = pi630 & ~pi1157;
  assign n17739 = ~n17737 & ~n17738;
  assign n17740 = pi787 & ~n17739;
  assign n17741 = n17701 & ~n17740;
  assign n17742 = ~n17495 & n17740;
  assign n17743 = ~n17741 & ~n17742;
  assign n17744 = pi644 & n17743;
  assign n17745 = ~pi644 & n17495;
  assign n17746 = ~pi715 & ~n17745;
  assign n17747 = ~n17744 & n17746;
  assign n17748 = pi1160 & ~n17747;
  assign n17749 = ~n17736 & n17748;
  assign n17750 = ~pi644 & ~n17728;
  assign n17751 = pi644 & n17733;
  assign n17752 = ~pi715 & ~n17751;
  assign n17753 = ~n17750 & n17752;
  assign n17754 = ~pi644 & n17743;
  assign n17755 = pi644 & n17495;
  assign n17756 = pi715 & ~n17755;
  assign n17757 = ~n17754 & n17756;
  assign n17758 = ~pi1160 & ~n17757;
  assign n17759 = ~n17753 & n17758;
  assign n17760 = pi790 & ~n17749;
  assign n17761 = ~n17759 & n17760;
  assign n17762 = ~pi790 & n17728;
  assign n17763 = ~po1038 & ~n17762;
  assign n17764 = ~n17761 & n17763;
  assign n17765 = ~pi140 & po1038;
  assign n17766 = ~pi832 & ~n17765;
  assign n17767 = ~n17764 & n17766;
  assign n17768 = ~pi140 & ~n2755;
  assign n17769 = ~pi738 & n17153;
  assign n17770 = ~n17768 & ~n17769;
  assign n17771 = ~pi778 & n17770;
  assign n17772 = ~pi625 & n17769;
  assign n17773 = ~n17770 & ~n17772;
  assign n17774 = pi1153 & ~n17773;
  assign n17775 = ~pi1153 & ~n17768;
  assign n17776 = ~n17772 & n17775;
  assign n17777 = ~n17774 & ~n17776;
  assign n17778 = pi778 & ~n17777;
  assign n17779 = ~n17771 & ~n17778;
  assign n17780 = n2755 & n17554;
  assign n17781 = n17779 & ~n17780;
  assign n17782 = n2755 & n17591;
  assign n17783 = n17781 & ~n17782;
  assign n17784 = n2755 & n17627;
  assign n17785 = n17783 & ~n17784;
  assign n17786 = ~pi626 & pi1158;
  assign n17787 = pi626 & ~pi1158;
  assign n17788 = ~n17786 & ~n17787;
  assign n17789 = ~pi626 & pi641;
  assign n17790 = pi626 & ~pi641;
  assign n17791 = ~n17789 & ~n17790;
  assign n17792 = ~n17788 & ~n17791;
  assign n17793 = n17785 & n17792;
  assign n17794 = n2755 & n17526;
  assign n17795 = ~pi761 & n16933;
  assign n17796 = ~n17768 & ~n17795;
  assign n17797 = ~n17794 & ~n17796;
  assign n17798 = ~pi785 & ~n17797;
  assign n17799 = n2755 & ~n17527;
  assign n17800 = ~n17796 & ~n17799;
  assign n17801 = pi1155 & ~n17800;
  assign n17802 = pi609 & n2755;
  assign n17803 = n17797 & ~n17802;
  assign n17804 = ~pi1155 & ~n17803;
  assign n17805 = ~n17801 & ~n17804;
  assign n17806 = pi785 & ~n17805;
  assign n17807 = ~n17798 & ~n17806;
  assign n17808 = ~pi781 & ~n17807;
  assign n17809 = ~pi618 & n2755;
  assign n17810 = n17807 & ~n17809;
  assign n17811 = pi1154 & ~n17810;
  assign n17812 = pi618 & n2755;
  assign n17813 = n17807 & ~n17812;
  assign n17814 = ~pi1154 & ~n17813;
  assign n17815 = ~n17811 & ~n17814;
  assign n17816 = pi781 & ~n17815;
  assign n17817 = ~n17808 & ~n17816;
  assign n17818 = ~pi789 & ~n17817;
  assign n17819 = pi619 & n17817;
  assign n17820 = ~pi619 & n17768;
  assign n17821 = pi1159 & ~n17820;
  assign n17822 = ~n17819 & n17821;
  assign n17823 = ~pi619 & n17817;
  assign n17824 = pi619 & n17768;
  assign n17825 = ~pi1159 & ~n17824;
  assign n17826 = ~n17823 & n17825;
  assign n17827 = ~n17822 & ~n17826;
  assign n17828 = pi789 & ~n17827;
  assign n17829 = ~n17818 & ~n17828;
  assign n17830 = pi626 & n17829;
  assign n17831 = ~pi626 & n17768;
  assign n17832 = pi1158 & ~n17831;
  assign n17833 = ~n17830 & n17832;
  assign n17834 = ~pi626 & n17829;
  assign n17835 = pi626 & n17768;
  assign n17836 = ~pi1158 & ~n17835;
  assign n17837 = ~n17834 & n17836;
  assign n17838 = ~n17833 & ~n17837;
  assign n17839 = ~n17669 & n17838;
  assign n17840 = ~n17793 & ~n17839;
  assign n17841 = pi788 & ~n17840;
  assign n17842 = ~n16842 & ~n17770;
  assign n17843 = pi625 & n17842;
  assign n17844 = n17796 & ~n17842;
  assign n17845 = ~n17843 & ~n17844;
  assign n17846 = n17775 & ~n17845;
  assign n17847 = ~pi608 & ~n17774;
  assign n17848 = ~n17846 & n17847;
  assign n17849 = pi1153 & n17796;
  assign n17850 = ~n17843 & n17849;
  assign n17851 = pi608 & ~n17776;
  assign n17852 = ~n17850 & n17851;
  assign n17853 = ~n17848 & ~n17852;
  assign n17854 = pi778 & ~n17853;
  assign n17855 = ~pi778 & ~n17844;
  assign n17856 = ~n17854 & ~n17855;
  assign n17857 = ~pi609 & ~n17856;
  assign n17858 = pi609 & n17779;
  assign n17859 = ~pi1155 & ~n17858;
  assign n17860 = ~n17857 & n17859;
  assign n17861 = ~pi660 & ~n17801;
  assign n17862 = ~n17860 & n17861;
  assign n17863 = pi609 & ~n17856;
  assign n17864 = ~pi609 & n17779;
  assign n17865 = pi1155 & ~n17864;
  assign n17866 = ~n17863 & n17865;
  assign n17867 = pi660 & ~n17804;
  assign n17868 = ~n17866 & n17867;
  assign n17869 = ~n17862 & ~n17868;
  assign n17870 = pi785 & ~n17869;
  assign n17871 = ~pi785 & ~n17856;
  assign n17872 = ~n17870 & ~n17871;
  assign n17873 = ~pi618 & ~n17872;
  assign n17874 = pi618 & n17781;
  assign n17875 = ~pi1154 & ~n17874;
  assign n17876 = ~n17873 & n17875;
  assign n17877 = ~pi627 & ~n17811;
  assign n17878 = ~n17876 & n17877;
  assign n17879 = pi618 & ~n17872;
  assign n17880 = ~pi618 & n17781;
  assign n17881 = pi1154 & ~n17880;
  assign n17882 = ~n17879 & n17881;
  assign n17883 = pi627 & ~n17814;
  assign n17884 = ~n17882 & n17883;
  assign n17885 = ~n17878 & ~n17884;
  assign n17886 = pi781 & ~n17885;
  assign n17887 = ~pi781 & ~n17872;
  assign n17888 = ~n17886 & ~n17887;
  assign n17889 = ~pi619 & ~n17888;
  assign n17890 = pi619 & n17783;
  assign n17891 = ~pi1159 & ~n17890;
  assign n17892 = ~n17889 & n17891;
  assign n17893 = ~pi648 & ~n17822;
  assign n17894 = ~n17892 & n17893;
  assign n17895 = pi619 & ~n17888;
  assign n17896 = ~pi619 & n17783;
  assign n17897 = pi1159 & ~n17896;
  assign n17898 = ~n17895 & n17897;
  assign n17899 = pi648 & ~n17826;
  assign n17900 = ~n17898 & n17899;
  assign n17901 = pi789 & ~n17894;
  assign n17902 = ~n17900 & n17901;
  assign n17903 = ~pi789 & n17888;
  assign n17904 = pi788 & ~n17788;
  assign n17905 = ~n17670 & ~n17904;
  assign n17906 = ~n17903 & n17905;
  assign n17907 = ~n17902 & n17906;
  assign n17908 = ~n17841 & ~n17907;
  assign n17909 = ~pi628 & ~n17908;
  assign n17910 = ~pi788 & ~n17829;
  assign n17911 = pi788 & ~n17838;
  assign n17912 = ~n17910 & ~n17911;
  assign n17913 = pi628 & n17912;
  assign n17914 = ~pi1156 & ~n17913;
  assign n17915 = ~n17909 & n17914;
  assign n17916 = n2755 & n17670;
  assign n17917 = n17785 & ~n17916;
  assign n17918 = ~pi628 & n2755;
  assign n17919 = n17917 & ~n17918;
  assign n17920 = pi1156 & ~n17919;
  assign n17921 = ~pi629 & ~n17920;
  assign n17922 = ~n17915 & n17921;
  assign n17923 = pi628 & ~n17908;
  assign n17924 = ~pi628 & n17912;
  assign n17925 = pi1156 & ~n17924;
  assign n17926 = ~n17923 & n17925;
  assign n17927 = pi628 & n2755;
  assign n17928 = n17917 & ~n17927;
  assign n17929 = ~pi1156 & ~n17928;
  assign n17930 = pi629 & ~n17929;
  assign n17931 = ~n17926 & n17930;
  assign n17932 = ~n17922 & ~n17931;
  assign n17933 = pi792 & ~n17932;
  assign n17934 = ~pi792 & ~n17908;
  assign n17935 = ~n17933 & ~n17934;
  assign n17936 = ~pi647 & ~n17935;
  assign n17937 = ~n17698 & n17912;
  assign n17938 = n17698 & n17768;
  assign n17939 = ~n17937 & ~n17938;
  assign n17940 = pi647 & ~n17939;
  assign n17941 = ~pi1157 & ~n17940;
  assign n17942 = ~n17936 & n17941;
  assign n17943 = ~pi628 & pi1156;
  assign n17944 = pi628 & ~pi1156;
  assign n17945 = ~n17943 & ~n17944;
  assign n17946 = pi792 & ~n17945;
  assign n17947 = n2755 & n17946;
  assign n17948 = n17917 & ~n17947;
  assign n17949 = pi647 & n17948;
  assign n17950 = ~pi647 & n17768;
  assign n17951 = pi1157 & ~n17950;
  assign n17952 = ~n17949 & n17951;
  assign n17953 = ~pi630 & ~n17952;
  assign n17954 = ~n17942 & n17953;
  assign n17955 = pi647 & ~n17935;
  assign n17956 = ~pi647 & ~n17939;
  assign n17957 = pi1157 & ~n17956;
  assign n17958 = ~n17955 & n17957;
  assign n17959 = ~pi647 & n17948;
  assign n17960 = pi647 & n17768;
  assign n17961 = ~pi1157 & ~n17960;
  assign n17962 = ~n17959 & n17961;
  assign n17963 = pi630 & ~n17962;
  assign n17964 = ~n17958 & n17963;
  assign n17965 = ~n17954 & ~n17964;
  assign n17966 = pi787 & ~n17965;
  assign n17967 = ~pi787 & ~n17935;
  assign n17968 = ~n17966 & ~n17967;
  assign n17969 = pi644 & ~n17968;
  assign n17970 = ~pi787 & ~n17948;
  assign n17971 = ~n17952 & ~n17962;
  assign n17972 = pi787 & ~n17971;
  assign n17973 = ~n17970 & ~n17972;
  assign n17974 = ~pi644 & n17973;
  assign n17975 = pi715 & ~n17974;
  assign n17976 = ~n17969 & n17975;
  assign n17977 = n17740 & ~n17768;
  assign n17978 = ~n17740 & n17939;
  assign n17979 = ~n17977 & ~n17978;
  assign n17980 = pi644 & n17979;
  assign n17981 = ~pi644 & n17768;
  assign n17982 = ~pi715 & ~n17981;
  assign n17983 = ~n17980 & n17982;
  assign n17984 = pi1160 & ~n17983;
  assign n17985 = ~n17976 & n17984;
  assign n17986 = ~pi644 & ~n17968;
  assign n17987 = pi644 & n17973;
  assign n17988 = ~pi715 & ~n17987;
  assign n17989 = ~n17986 & n17988;
  assign n17990 = ~pi644 & n17979;
  assign n17991 = pi644 & n17768;
  assign n17992 = pi715 & ~n17991;
  assign n17993 = ~n17990 & n17992;
  assign n17994 = ~pi1160 & ~n17993;
  assign n17995 = ~n17989 & n17994;
  assign n17996 = ~n17985 & ~n17995;
  assign n17997 = pi790 & ~n17996;
  assign n17998 = ~pi790 & ~n17968;
  assign n17999 = pi832 & ~n17998;
  assign n18000 = ~n17997 & n17999;
  assign po297 = ~n17767 & ~n18000;
  assign n18002 = pi141 & ~n3268;
  assign n18003 = ~pi141 & ~n16968;
  assign n18004 = pi749 & n16970;
  assign n18005 = ~n18003 & ~n18004;
  assign n18006 = pi38 & ~n18005;
  assign n18007 = ~pi749 & n16814;
  assign n18008 = pi141 & n16961;
  assign n18009 = ~n18007 & ~n18008;
  assign n18010 = pi39 & ~n18009;
  assign n18011 = ~pi141 & n16907;
  assign n18012 = pi141 & n16919;
  assign n18013 = pi749 & ~n18012;
  assign n18014 = ~n18011 & n18013;
  assign n18015 = ~pi39 & n16655;
  assign n18016 = ~pi141 & ~pi749;
  assign n18017 = ~n18015 & n18016;
  assign n18018 = ~n18014 & ~n18017;
  assign n18019 = ~pi38 & ~n18018;
  assign n18020 = ~n18010 & n18019;
  assign n18021 = ~n18006 & ~n18020;
  assign n18022 = ~pi706 & ~n18021;
  assign n18023 = ~pi141 & n17074;
  assign n18024 = pi141 & n17166;
  assign n18025 = ~pi749 & ~n18024;
  assign n18026 = ~n18023 & n18025;
  assign n18027 = pi141 & n17233;
  assign n18028 = ~pi141 & ~n17295;
  assign n18029 = pi749 & ~n18028;
  assign n18030 = ~n18027 & n18029;
  assign n18031 = pi39 & ~n18030;
  assign n18032 = ~n18026 & n18031;
  assign n18033 = ~pi141 & n17317;
  assign n18034 = pi141 & n17340;
  assign n18035 = ~pi749 & ~n18033;
  assign n18036 = ~n18034 & n18035;
  assign n18037 = ~pi141 & ~n17344;
  assign n18038 = pi141 & ~n17351;
  assign n18039 = pi749 & ~n18038;
  assign n18040 = ~n18037 & n18039;
  assign n18041 = ~pi39 & ~n18040;
  assign n18042 = ~n18036 & n18041;
  assign n18043 = ~pi38 & ~n18042;
  assign n18044 = ~n18032 & n18043;
  assign n18045 = ~pi39 & n17365;
  assign n18046 = pi38 & ~n18045;
  assign n18047 = n18005 & n18046;
  assign n18048 = pi706 & ~n18047;
  assign n18049 = ~n18044 & n18048;
  assign n18050 = n3268 & ~n18022;
  assign n18051 = ~n18049 & n18050;
  assign n18052 = ~n18002 & ~n18051;
  assign n18053 = ~pi625 & n18052;
  assign n18054 = n3268 & n18021;
  assign n18055 = ~n18002 & ~n18054;
  assign n18056 = pi625 & n18055;
  assign n18057 = ~pi1153 & ~n18056;
  assign n18058 = ~n18053 & n18057;
  assign n18059 = ~pi39 & n17315;
  assign n18060 = ~n17470 & ~n18059;
  assign n18061 = ~pi141 & n18060;
  assign n18062 = pi39 & ~n17419;
  assign n18063 = ~pi39 & n17350;
  assign n18064 = ~n18062 & ~n18063;
  assign n18065 = pi141 & ~n18064;
  assign n18066 = ~pi38 & ~n18065;
  assign n18067 = ~n18061 & n18066;
  assign n18068 = n17480 & ~n18003;
  assign n18069 = pi706 & ~n18068;
  assign n18070 = ~n18067 & n18069;
  assign n18071 = ~pi141 & ~pi706;
  assign n18072 = ~n17487 & n18071;
  assign n18073 = n3268 & ~n18072;
  assign n18074 = ~n18070 & n18073;
  assign n18075 = ~n18002 & ~n18074;
  assign n18076 = pi625 & n18075;
  assign n18077 = ~pi141 & ~n17494;
  assign n18078 = ~pi625 & n18077;
  assign n18079 = pi1153 & ~n18078;
  assign n18080 = ~n18076 & n18079;
  assign n18081 = ~pi608 & ~n18080;
  assign n18082 = ~n18058 & n18081;
  assign n18083 = pi625 & n18052;
  assign n18084 = ~pi625 & n18055;
  assign n18085 = pi1153 & ~n18084;
  assign n18086 = ~n18083 & n18085;
  assign n18087 = ~pi625 & n18075;
  assign n18088 = pi625 & n18077;
  assign n18089 = ~pi1153 & ~n18088;
  assign n18090 = ~n18087 & n18089;
  assign n18091 = pi608 & ~n18090;
  assign n18092 = ~n18086 & n18091;
  assign n18093 = ~n18082 & ~n18092;
  assign n18094 = pi778 & ~n18093;
  assign n18095 = ~pi778 & n18052;
  assign n18096 = ~n18094 & ~n18095;
  assign n18097 = ~pi609 & ~n18096;
  assign n18098 = ~pi778 & ~n18075;
  assign n18099 = ~n18080 & ~n18090;
  assign n18100 = pi778 & ~n18099;
  assign n18101 = ~n18098 & ~n18100;
  assign n18102 = pi609 & n18101;
  assign n18103 = ~pi1155 & ~n18102;
  assign n18104 = ~n18097 & n18103;
  assign n18105 = ~n17527 & ~n18077;
  assign n18106 = ~n17526 & ~n18055;
  assign n18107 = pi609 & n18106;
  assign n18108 = ~n18105 & ~n18107;
  assign n18109 = pi1155 & ~n18108;
  assign n18110 = ~pi660 & ~n18109;
  assign n18111 = ~n18104 & n18110;
  assign n18112 = pi609 & ~n18096;
  assign n18113 = ~pi609 & n18101;
  assign n18114 = pi1155 & ~n18113;
  assign n18115 = ~n18112 & n18114;
  assign n18116 = ~n17539 & ~n18077;
  assign n18117 = ~pi609 & n18106;
  assign n18118 = ~n18116 & ~n18117;
  assign n18119 = ~pi1155 & ~n18118;
  assign n18120 = pi660 & ~n18119;
  assign n18121 = ~n18115 & n18120;
  assign n18122 = ~n18111 & ~n18121;
  assign n18123 = pi785 & ~n18122;
  assign n18124 = ~pi785 & ~n18096;
  assign n18125 = ~n18123 & ~n18124;
  assign n18126 = ~pi618 & ~n18125;
  assign n18127 = ~n17554 & ~n18101;
  assign n18128 = n17554 & ~n18077;
  assign n18129 = ~n18127 & ~n18128;
  assign n18130 = pi618 & n18129;
  assign n18131 = ~pi1154 & ~n18130;
  assign n18132 = ~n18126 & n18131;
  assign n18133 = n17526 & ~n18077;
  assign n18134 = ~n18106 & ~n18133;
  assign n18135 = ~pi785 & ~n18134;
  assign n18136 = ~n18109 & ~n18119;
  assign n18137 = pi785 & ~n18136;
  assign n18138 = ~n18135 & ~n18137;
  assign n18139 = pi618 & n18138;
  assign n18140 = ~pi618 & n18077;
  assign n18141 = pi1154 & ~n18140;
  assign n18142 = ~n18139 & n18141;
  assign n18143 = ~pi627 & ~n18142;
  assign n18144 = ~n18132 & n18143;
  assign n18145 = pi618 & ~n18125;
  assign n18146 = ~pi618 & n18129;
  assign n18147 = pi1154 & ~n18146;
  assign n18148 = ~n18145 & n18147;
  assign n18149 = ~pi618 & n18138;
  assign n18150 = pi618 & n18077;
  assign n18151 = ~pi1154 & ~n18150;
  assign n18152 = ~n18149 & n18151;
  assign n18153 = pi627 & ~n18152;
  assign n18154 = ~n18148 & n18153;
  assign n18155 = ~n18144 & ~n18154;
  assign n18156 = pi781 & ~n18155;
  assign n18157 = ~pi781 & ~n18125;
  assign n18158 = ~n18156 & ~n18157;
  assign n18159 = ~pi619 & ~n18158;
  assign n18160 = ~n17591 & n18129;
  assign n18161 = n17591 & n18077;
  assign n18162 = ~n18160 & ~n18161;
  assign n18163 = pi619 & ~n18162;
  assign n18164 = ~pi1159 & ~n18163;
  assign n18165 = ~n18159 & n18164;
  assign n18166 = ~pi781 & ~n18138;
  assign n18167 = ~n18142 & ~n18152;
  assign n18168 = pi781 & ~n18167;
  assign n18169 = ~n18166 & ~n18168;
  assign n18170 = pi619 & n18169;
  assign n18171 = ~pi619 & n18077;
  assign n18172 = pi1159 & ~n18171;
  assign n18173 = ~n18170 & n18172;
  assign n18174 = ~pi648 & ~n18173;
  assign n18175 = ~n18165 & n18174;
  assign n18176 = pi619 & ~n18158;
  assign n18177 = ~pi619 & ~n18162;
  assign n18178 = pi1159 & ~n18177;
  assign n18179 = ~n18176 & n18178;
  assign n18180 = ~pi619 & n18169;
  assign n18181 = pi619 & n18077;
  assign n18182 = ~pi1159 & ~n18181;
  assign n18183 = ~n18180 & n18182;
  assign n18184 = pi648 & ~n18183;
  assign n18185 = ~n18179 & n18184;
  assign n18186 = ~n18175 & ~n18185;
  assign n18187 = pi789 & ~n18186;
  assign n18188 = ~pi789 & ~n18158;
  assign n18189 = ~n18187 & ~n18188;
  assign n18190 = ~pi788 & n18189;
  assign n18191 = ~pi626 & n18189;
  assign n18192 = n17627 & ~n18077;
  assign n18193 = ~n17627 & n18162;
  assign n18194 = ~n18192 & ~n18193;
  assign n18195 = pi626 & ~n18194;
  assign n18196 = ~pi641 & ~n18195;
  assign n18197 = ~n18191 & n18196;
  assign n18198 = ~pi789 & ~n18169;
  assign n18199 = ~n18173 & ~n18183;
  assign n18200 = pi789 & ~n18199;
  assign n18201 = ~n18198 & ~n18200;
  assign n18202 = ~pi626 & n18201;
  assign n18203 = pi626 & n18077;
  assign n18204 = ~pi1158 & ~n18203;
  assign n18205 = ~n18202 & n18204;
  assign n18206 = ~n17634 & ~n18205;
  assign n18207 = ~n18197 & ~n18206;
  assign n18208 = pi626 & n18189;
  assign n18209 = ~pi626 & ~n18194;
  assign n18210 = pi641 & ~n18209;
  assign n18211 = ~n18208 & n18210;
  assign n18212 = pi626 & n18201;
  assign n18213 = ~pi626 & n18077;
  assign n18214 = pi1158 & ~n18213;
  assign n18215 = ~n18212 & n18214;
  assign n18216 = ~n17649 & ~n18215;
  assign n18217 = ~n18211 & ~n18216;
  assign n18218 = ~n18207 & ~n18217;
  assign n18219 = pi788 & ~n18218;
  assign n18220 = ~n18190 & ~n18219;
  assign n18221 = ~pi628 & n18220;
  assign n18222 = ~n18205 & ~n18215;
  assign n18223 = pi788 & ~n18222;
  assign n18224 = ~pi788 & ~n18201;
  assign n18225 = ~n18223 & ~n18224;
  assign n18226 = pi628 & n18225;
  assign n18227 = ~pi1156 & ~n18226;
  assign n18228 = ~n18221 & n18227;
  assign n18229 = ~n17670 & n18194;
  assign n18230 = n17670 & n18077;
  assign n18231 = ~n18229 & ~n18230;
  assign n18232 = pi628 & ~n18231;
  assign n18233 = ~pi628 & n18077;
  assign n18234 = pi1156 & ~n18233;
  assign n18235 = ~n18232 & n18234;
  assign n18236 = ~pi629 & ~n18235;
  assign n18237 = ~n18228 & n18236;
  assign n18238 = pi628 & n18220;
  assign n18239 = ~pi628 & n18225;
  assign n18240 = pi1156 & ~n18239;
  assign n18241 = ~n18238 & n18240;
  assign n18242 = ~pi628 & ~n18231;
  assign n18243 = pi628 & n18077;
  assign n18244 = ~pi1156 & ~n18243;
  assign n18245 = ~n18242 & n18244;
  assign n18246 = pi629 & ~n18245;
  assign n18247 = ~n18241 & n18246;
  assign n18248 = ~n18237 & ~n18247;
  assign n18249 = pi792 & ~n18248;
  assign n18250 = ~pi792 & n18220;
  assign n18251 = ~n18249 & ~n18250;
  assign n18252 = ~pi647 & ~n18251;
  assign n18253 = ~n17698 & n18225;
  assign n18254 = n17698 & n18077;
  assign n18255 = ~n18253 & ~n18254;
  assign n18256 = pi647 & ~n18255;
  assign n18257 = ~pi1157 & ~n18256;
  assign n18258 = ~n18252 & n18257;
  assign n18259 = ~pi792 & n18231;
  assign n18260 = ~n18235 & ~n18245;
  assign n18261 = pi792 & ~n18260;
  assign n18262 = ~n18259 & ~n18261;
  assign n18263 = pi647 & n18262;
  assign n18264 = ~pi647 & n18077;
  assign n18265 = pi1157 & ~n18264;
  assign n18266 = ~n18263 & n18265;
  assign n18267 = ~pi630 & ~n18266;
  assign n18268 = ~n18258 & n18267;
  assign n18269 = pi647 & ~n18251;
  assign n18270 = ~pi647 & ~n18255;
  assign n18271 = pi1157 & ~n18270;
  assign n18272 = ~n18269 & n18271;
  assign n18273 = ~pi647 & n18262;
  assign n18274 = pi647 & n18077;
  assign n18275 = ~pi1157 & ~n18274;
  assign n18276 = ~n18273 & n18275;
  assign n18277 = pi630 & ~n18276;
  assign n18278 = ~n18272 & n18277;
  assign n18279 = ~n18268 & ~n18278;
  assign n18280 = pi787 & ~n18279;
  assign n18281 = ~pi787 & ~n18251;
  assign n18282 = ~n18280 & ~n18281;
  assign n18283 = pi644 & ~n18282;
  assign n18284 = ~pi787 & ~n18262;
  assign n18285 = ~n18266 & ~n18276;
  assign n18286 = pi787 & ~n18285;
  assign n18287 = ~n18284 & ~n18286;
  assign n18288 = ~pi644 & n18287;
  assign n18289 = pi715 & ~n18288;
  assign n18290 = ~n18283 & n18289;
  assign n18291 = n17740 & ~n18077;
  assign n18292 = ~n17740 & n18255;
  assign n18293 = ~n18291 & ~n18292;
  assign n18294 = pi644 & n18293;
  assign n18295 = ~pi644 & n18077;
  assign n18296 = ~pi715 & ~n18295;
  assign n18297 = ~n18294 & n18296;
  assign n18298 = pi1160 & ~n18297;
  assign n18299 = ~n18290 & n18298;
  assign n18300 = ~pi644 & ~n18282;
  assign n18301 = pi644 & n18287;
  assign n18302 = ~pi715 & ~n18301;
  assign n18303 = ~n18300 & n18302;
  assign n18304 = ~pi644 & n18293;
  assign n18305 = pi644 & n18077;
  assign n18306 = pi715 & ~n18305;
  assign n18307 = ~n18304 & n18306;
  assign n18308 = ~pi1160 & ~n18307;
  assign n18309 = ~n18303 & n18308;
  assign n18310 = pi790 & ~n18299;
  assign n18311 = ~n18309 & n18310;
  assign n18312 = ~pi790 & n18282;
  assign n18313 = ~po1038 & ~n18312;
  assign n18314 = ~n18311 & n18313;
  assign n18315 = ~pi141 & po1038;
  assign n18316 = ~pi832 & ~n18315;
  assign n18317 = ~n18314 & n18316;
  assign n18318 = ~pi141 & ~n2755;
  assign n18319 = pi706 & n17153;
  assign n18320 = ~n18318 & ~n18319;
  assign n18321 = ~pi778 & n18320;
  assign n18322 = ~pi625 & n18319;
  assign n18323 = ~n18320 & ~n18322;
  assign n18324 = pi1153 & ~n18323;
  assign n18325 = ~pi1153 & ~n18318;
  assign n18326 = ~n18322 & n18325;
  assign n18327 = ~n18324 & ~n18326;
  assign n18328 = pi778 & ~n18327;
  assign n18329 = ~n18321 & ~n18328;
  assign n18330 = ~n17780 & n18329;
  assign n18331 = ~n17782 & n18330;
  assign n18332 = ~n17784 & n18331;
  assign n18333 = n17792 & n18332;
  assign n18334 = pi749 & n16933;
  assign n18335 = ~n18318 & ~n18334;
  assign n18336 = ~n17794 & ~n18335;
  assign n18337 = ~pi785 & ~n18336;
  assign n18338 = ~n17799 & ~n18335;
  assign n18339 = pi1155 & ~n18338;
  assign n18340 = ~n17802 & n18336;
  assign n18341 = ~pi1155 & ~n18340;
  assign n18342 = ~n18339 & ~n18341;
  assign n18343 = pi785 & ~n18342;
  assign n18344 = ~n18337 & ~n18343;
  assign n18345 = ~pi781 & ~n18344;
  assign n18346 = ~n17809 & n18344;
  assign n18347 = pi1154 & ~n18346;
  assign n18348 = ~n17812 & n18344;
  assign n18349 = ~pi1154 & ~n18348;
  assign n18350 = ~n18347 & ~n18349;
  assign n18351 = pi781 & ~n18350;
  assign n18352 = ~n18345 & ~n18351;
  assign n18353 = ~pi789 & ~n18352;
  assign n18354 = pi619 & n18352;
  assign n18355 = ~pi619 & n18318;
  assign n18356 = pi1159 & ~n18355;
  assign n18357 = ~n18354 & n18356;
  assign n18358 = ~pi619 & n18352;
  assign n18359 = pi619 & n18318;
  assign n18360 = ~pi1159 & ~n18359;
  assign n18361 = ~n18358 & n18360;
  assign n18362 = ~n18357 & ~n18361;
  assign n18363 = pi789 & ~n18362;
  assign n18364 = ~n18353 & ~n18363;
  assign n18365 = pi626 & n18364;
  assign n18366 = ~pi626 & n18318;
  assign n18367 = pi1158 & ~n18366;
  assign n18368 = ~n18365 & n18367;
  assign n18369 = ~pi626 & n18364;
  assign n18370 = pi626 & n18318;
  assign n18371 = ~pi1158 & ~n18370;
  assign n18372 = ~n18369 & n18371;
  assign n18373 = ~n18368 & ~n18372;
  assign n18374 = ~n17669 & n18373;
  assign n18375 = ~n18333 & ~n18374;
  assign n18376 = pi788 & ~n18375;
  assign n18377 = ~n16842 & ~n18320;
  assign n18378 = pi625 & n18377;
  assign n18379 = n18335 & ~n18377;
  assign n18380 = ~n18378 & ~n18379;
  assign n18381 = n18325 & ~n18380;
  assign n18382 = ~pi608 & ~n18324;
  assign n18383 = ~n18381 & n18382;
  assign n18384 = pi1153 & n18335;
  assign n18385 = ~n18378 & n18384;
  assign n18386 = pi608 & ~n18326;
  assign n18387 = ~n18385 & n18386;
  assign n18388 = ~n18383 & ~n18387;
  assign n18389 = pi778 & ~n18388;
  assign n18390 = ~pi778 & ~n18379;
  assign n18391 = ~n18389 & ~n18390;
  assign n18392 = ~pi609 & ~n18391;
  assign n18393 = pi609 & n18329;
  assign n18394 = ~pi1155 & ~n18393;
  assign n18395 = ~n18392 & n18394;
  assign n18396 = ~pi660 & ~n18339;
  assign n18397 = ~n18395 & n18396;
  assign n18398 = pi609 & ~n18391;
  assign n18399 = ~pi609 & n18329;
  assign n18400 = pi1155 & ~n18399;
  assign n18401 = ~n18398 & n18400;
  assign n18402 = pi660 & ~n18341;
  assign n18403 = ~n18401 & n18402;
  assign n18404 = ~n18397 & ~n18403;
  assign n18405 = pi785 & ~n18404;
  assign n18406 = ~pi785 & ~n18391;
  assign n18407 = ~n18405 & ~n18406;
  assign n18408 = ~pi618 & ~n18407;
  assign n18409 = pi618 & n18330;
  assign n18410 = ~pi1154 & ~n18409;
  assign n18411 = ~n18408 & n18410;
  assign n18412 = ~pi627 & ~n18347;
  assign n18413 = ~n18411 & n18412;
  assign n18414 = pi618 & ~n18407;
  assign n18415 = ~pi618 & n18330;
  assign n18416 = pi1154 & ~n18415;
  assign n18417 = ~n18414 & n18416;
  assign n18418 = pi627 & ~n18349;
  assign n18419 = ~n18417 & n18418;
  assign n18420 = ~n18413 & ~n18419;
  assign n18421 = pi781 & ~n18420;
  assign n18422 = ~pi781 & ~n18407;
  assign n18423 = ~n18421 & ~n18422;
  assign n18424 = ~pi619 & ~n18423;
  assign n18425 = pi619 & n18331;
  assign n18426 = ~pi1159 & ~n18425;
  assign n18427 = ~n18424 & n18426;
  assign n18428 = ~pi648 & ~n18357;
  assign n18429 = ~n18427 & n18428;
  assign n18430 = pi619 & ~n18423;
  assign n18431 = ~pi619 & n18331;
  assign n18432 = pi1159 & ~n18431;
  assign n18433 = ~n18430 & n18432;
  assign n18434 = pi648 & ~n18361;
  assign n18435 = ~n18433 & n18434;
  assign n18436 = pi789 & ~n18429;
  assign n18437 = ~n18435 & n18436;
  assign n18438 = ~pi789 & n18423;
  assign n18439 = n17905 & ~n18438;
  assign n18440 = ~n18437 & n18439;
  assign n18441 = ~n18376 & ~n18440;
  assign n18442 = ~pi628 & ~n18441;
  assign n18443 = ~pi788 & ~n18364;
  assign n18444 = pi788 & ~n18373;
  assign n18445 = ~n18443 & ~n18444;
  assign n18446 = pi628 & n18445;
  assign n18447 = ~pi1156 & ~n18446;
  assign n18448 = ~n18442 & n18447;
  assign n18449 = ~n17916 & n18332;
  assign n18450 = ~n17918 & n18449;
  assign n18451 = pi1156 & ~n18450;
  assign n18452 = ~pi629 & ~n18451;
  assign n18453 = ~n18448 & n18452;
  assign n18454 = pi628 & ~n18441;
  assign n18455 = ~pi628 & n18445;
  assign n18456 = pi1156 & ~n18455;
  assign n18457 = ~n18454 & n18456;
  assign n18458 = ~n17927 & n18449;
  assign n18459 = ~pi1156 & ~n18458;
  assign n18460 = pi629 & ~n18459;
  assign n18461 = ~n18457 & n18460;
  assign n18462 = ~n18453 & ~n18461;
  assign n18463 = pi792 & ~n18462;
  assign n18464 = ~pi792 & ~n18441;
  assign n18465 = ~n18463 & ~n18464;
  assign n18466 = ~pi647 & ~n18465;
  assign n18467 = ~n17698 & n18445;
  assign n18468 = n17698 & n18318;
  assign n18469 = ~n18467 & ~n18468;
  assign n18470 = pi647 & ~n18469;
  assign n18471 = ~pi1157 & ~n18470;
  assign n18472 = ~n18466 & n18471;
  assign n18473 = ~n17947 & n18449;
  assign n18474 = pi647 & n18473;
  assign n18475 = ~pi647 & n18318;
  assign n18476 = pi1157 & ~n18475;
  assign n18477 = ~n18474 & n18476;
  assign n18478 = ~pi630 & ~n18477;
  assign n18479 = ~n18472 & n18478;
  assign n18480 = pi647 & ~n18465;
  assign n18481 = ~pi647 & ~n18469;
  assign n18482 = pi1157 & ~n18481;
  assign n18483 = ~n18480 & n18482;
  assign n18484 = ~pi647 & n18473;
  assign n18485 = pi647 & n18318;
  assign n18486 = ~pi1157 & ~n18485;
  assign n18487 = ~n18484 & n18486;
  assign n18488 = pi630 & ~n18487;
  assign n18489 = ~n18483 & n18488;
  assign n18490 = ~n18479 & ~n18489;
  assign n18491 = pi787 & ~n18490;
  assign n18492 = ~pi787 & ~n18465;
  assign n18493 = ~n18491 & ~n18492;
  assign n18494 = pi644 & ~n18493;
  assign n18495 = ~pi787 & ~n18473;
  assign n18496 = ~n18477 & ~n18487;
  assign n18497 = pi787 & ~n18496;
  assign n18498 = ~n18495 & ~n18497;
  assign n18499 = ~pi644 & n18498;
  assign n18500 = pi715 & ~n18499;
  assign n18501 = ~n18494 & n18500;
  assign n18502 = n17740 & ~n18318;
  assign n18503 = ~n17740 & n18469;
  assign n18504 = ~n18502 & ~n18503;
  assign n18505 = pi644 & n18504;
  assign n18506 = ~pi644 & n18318;
  assign n18507 = ~pi715 & ~n18506;
  assign n18508 = ~n18505 & n18507;
  assign n18509 = pi1160 & ~n18508;
  assign n18510 = ~n18501 & n18509;
  assign n18511 = ~pi644 & ~n18493;
  assign n18512 = pi644 & n18498;
  assign n18513 = ~pi715 & ~n18512;
  assign n18514 = ~n18511 & n18513;
  assign n18515 = ~pi644 & n18504;
  assign n18516 = pi644 & n18318;
  assign n18517 = pi715 & ~n18516;
  assign n18518 = ~n18515 & n18517;
  assign n18519 = ~pi1160 & ~n18518;
  assign n18520 = ~n18514 & n18519;
  assign n18521 = ~n18510 & ~n18520;
  assign n18522 = pi790 & ~n18521;
  assign n18523 = ~pi790 & ~n18493;
  assign n18524 = pi832 & ~n18523;
  assign n18525 = ~n18522 & n18524;
  assign po298 = ~n18317 & ~n18525;
  assign n18527 = pi142 & ~n3268;
  assign n18528 = pi142 & ~n16837;
  assign n18529 = n17307 & n18528;
  assign n18530 = ~pi142 & ~n16911;
  assign n18531 = ~n17346 & n18530;
  assign n18532 = ~n18529 & ~n18531;
  assign n18533 = pi743 & ~n18532;
  assign n18534 = ~pi142 & n17330;
  assign n18535 = pi142 & ~n16911;
  assign n18536 = ~n17307 & n18535;
  assign n18537 = ~pi743 & ~n18536;
  assign n18538 = ~n18534 & n18537;
  assign n18539 = ~pi299 & ~n18538;
  assign n18540 = ~n18533 & n18539;
  assign n18541 = ~pi142 & ~n16916;
  assign n18542 = ~n17348 & n18541;
  assign n18543 = pi142 & n16824;
  assign n18544 = ~n17312 & n18543;
  assign n18545 = ~n18542 & ~n18544;
  assign n18546 = pi743 & ~n18545;
  assign n18547 = ~pi142 & n17338;
  assign n18548 = pi142 & ~n16916;
  assign n18549 = ~n17313 & n18548;
  assign n18550 = ~pi743 & ~n18549;
  assign n18551 = ~n18547 & n18550;
  assign n18552 = pi299 & ~n18546;
  assign n18553 = ~n18551 & n18552;
  assign n18554 = ~n18540 & ~n18553;
  assign n18555 = pi735 & ~n18554;
  assign n18556 = pi743 & ~n18530;
  assign n18557 = ~n18528 & n18556;
  assign n18558 = pi142 & ~pi743;
  assign n18559 = ~n16653 & n18558;
  assign n18560 = ~pi299 & ~n18559;
  assign n18561 = ~n18557 & n18560;
  assign n18562 = pi142 & ~n16649;
  assign n18563 = ~pi743 & ~n18562;
  assign n18564 = ~n18541 & ~n18563;
  assign n18565 = ~n18543 & n18564;
  assign n18566 = pi299 & ~n18565;
  assign n18567 = ~n18561 & ~n18566;
  assign n18568 = ~pi735 & n18567;
  assign n18569 = ~pi39 & ~n18568;
  assign n18570 = ~n18555 & n18569;
  assign n18571 = pi142 & n17276;
  assign n18572 = ~pi142 & n17214;
  assign n18573 = pi743 & ~n18572;
  assign n18574 = ~n18571 & n18573;
  assign n18575 = ~pi142 & ~n17136;
  assign n18576 = pi142 & n17016;
  assign n18577 = ~pi743 & ~n18576;
  assign n18578 = ~n18575 & n18577;
  assign n18579 = ~n18574 & ~n18578;
  assign n18580 = pi735 & ~n18579;
  assign n18581 = pi142 & ~n16704;
  assign n18582 = ~pi743 & ~n18581;
  assign n18583 = pi142 & ~n16886;
  assign n18584 = pi743 & n17210;
  assign n18585 = ~n18583 & n18584;
  assign n18586 = ~n18582 & ~n18585;
  assign n18587 = ~pi735 & n18586;
  assign n18588 = ~n18580 & ~n18587;
  assign n18589 = ~n6197 & n18588;
  assign n18590 = ~pi142 & ~n17208;
  assign n18591 = pi142 & ~n17267;
  assign n18592 = pi743 & ~n18590;
  assign n18593 = ~n18591 & n18592;
  assign n18594 = pi142 & n17006;
  assign n18595 = ~pi142 & n17142;
  assign n18596 = ~pi743 & ~n18595;
  assign n18597 = ~n18594 & n18596;
  assign n18598 = ~n18593 & ~n18597;
  assign n18599 = pi735 & ~n18598;
  assign n18600 = pi142 & ~n16726;
  assign n18601 = ~pi743 & ~n18600;
  assign n18602 = pi142 & n16877;
  assign n18603 = pi743 & n16943;
  assign n18604 = ~n18602 & n18603;
  assign n18605 = ~n18601 & ~n18604;
  assign n18606 = ~pi735 & n18605;
  assign n18607 = ~n18599 & ~n18606;
  assign n18608 = n6197 & n18607;
  assign n18609 = pi223 & ~n18608;
  assign n18610 = ~n18589 & n18609;
  assign n18611 = pi142 & n17254;
  assign n18612 = ~pi142 & ~n17193;
  assign n18613 = pi743 & ~n18611;
  assign n18614 = ~n18612 & n18613;
  assign n18615 = pi142 & n17038;
  assign n18616 = ~pi142 & n17117;
  assign n18617 = ~pi743 & ~n18616;
  assign n18618 = ~n18615 & n18617;
  assign n18619 = ~n18614 & ~n18618;
  assign n18620 = pi735 & ~n18619;
  assign n18621 = ~pi142 & n16927;
  assign n18622 = pi142 & n16861;
  assign n18623 = ~n18621 & ~n18622;
  assign n18624 = pi743 & ~n18623;
  assign n18625 = pi142 & ~n16776;
  assign n18626 = ~pi743 & ~n18625;
  assign n18627 = ~n18624 & ~n18626;
  assign n18628 = ~pi735 & n18627;
  assign n18629 = ~n18620 & ~n18628;
  assign n18630 = n6197 & ~n18629;
  assign n18631 = ~pi142 & ~n17179;
  assign n18632 = pi142 & n17243;
  assign n18633 = pi743 & ~n18632;
  assign n18634 = ~n18631 & n18633;
  assign n18635 = ~pi142 & ~n17102;
  assign n18636 = pi142 & n17050;
  assign n18637 = ~pi743 & ~n18636;
  assign n18638 = ~n18635 & n18637;
  assign n18639 = ~n18634 & ~n18638;
  assign n18640 = pi735 & ~n18639;
  assign n18641 = pi142 & ~n16785;
  assign n18642 = ~pi743 & ~n18641;
  assign n18643 = pi142 & ~n16843;
  assign n18644 = pi743 & ~n16929;
  assign n18645 = ~n18643 & n18644;
  assign n18646 = ~n18642 & ~n18645;
  assign n18647 = ~pi735 & n18646;
  assign n18648 = ~n18640 & ~n18647;
  assign n18649 = ~n6197 & ~n18648;
  assign n18650 = ~n3053 & ~n18649;
  assign n18651 = ~n18630 & n18650;
  assign n18652 = pi142 & ~n16661;
  assign n18653 = pi743 & n16922;
  assign n18654 = ~n18652 & ~n18653;
  assign n18655 = ~pi735 & n18654;
  assign n18656 = pi142 & ~n16665;
  assign n18657 = pi743 & n16933;
  assign n18658 = n3096 & n18657;
  assign n18659 = ~n18656 & ~n18658;
  assign n18660 = ~n17365 & n18659;
  assign n18661 = ~n16658 & ~n18660;
  assign n18662 = pi735 & ~n18661;
  assign n18663 = ~n18652 & n18662;
  assign n18664 = ~n18655 & ~n18663;
  assign n18665 = n3053 & ~n18664;
  assign n18666 = ~pi223 & ~n18665;
  assign n18667 = ~n18651 & n18666;
  assign n18668 = ~n18610 & ~n18667;
  assign n18669 = ~pi299 & ~n18668;
  assign n18670 = ~n6223 & n18588;
  assign n18671 = n6223 & n18607;
  assign n18672 = pi215 & ~n18671;
  assign n18673 = ~n18670 & n18672;
  assign n18674 = n6223 & ~n18629;
  assign n18675 = ~n6223 & ~n18648;
  assign n18676 = ~n3461 & ~n18675;
  assign n18677 = ~n18674 & n18676;
  assign n18678 = n3461 & ~n18664;
  assign n18679 = ~pi215 & ~n18678;
  assign n18680 = ~n18677 & n18679;
  assign n18681 = ~n18673 & ~n18680;
  assign n18682 = pi299 & ~n18681;
  assign n18683 = pi39 & ~n18669;
  assign n18684 = ~n18682 & n18683;
  assign n18685 = ~n18570 & ~n18684;
  assign n18686 = ~pi38 & ~n18685;
  assign n18687 = pi39 & pi142;
  assign n18688 = pi38 & ~n18687;
  assign n18689 = pi735 & n17365;
  assign n18690 = n18659 & ~n18689;
  assign n18691 = ~pi39 & ~n18690;
  assign n18692 = n18688 & ~n18691;
  assign n18693 = n3268 & ~n18692;
  assign n18694 = ~n18686 & n18693;
  assign n18695 = ~n18527 & ~n18694;
  assign n18696 = pi625 & n18695;
  assign n18697 = ~n6223 & n18646;
  assign n18698 = n6223 & n18627;
  assign n18699 = ~n18697 & ~n18698;
  assign n18700 = ~n3461 & ~n18699;
  assign n18701 = n3461 & ~n18654;
  assign n18702 = ~pi215 & ~n18701;
  assign n18703 = ~n18700 & n18702;
  assign n18704 = ~n6223 & n18586;
  assign n18705 = n6223 & n18605;
  assign n18706 = pi215 & ~n18705;
  assign n18707 = ~n18704 & n18706;
  assign n18708 = ~n18703 & ~n18707;
  assign n18709 = pi299 & ~n18708;
  assign n18710 = n6197 & n18627;
  assign n18711 = ~n6197 & n18646;
  assign n18712 = ~n3053 & ~n18711;
  assign n18713 = ~n18710 & n18712;
  assign n18714 = n3053 & n18654;
  assign n18715 = ~pi223 & ~n18714;
  assign n18716 = ~n18713 & n18715;
  assign n18717 = ~n6197 & ~n18586;
  assign n18718 = n6197 & ~n18605;
  assign n18719 = pi223 & ~n18718;
  assign n18720 = ~n18717 & n18719;
  assign n18721 = ~pi299 & ~n18720;
  assign n18722 = ~n18716 & n18721;
  assign n18723 = pi39 & ~n18722;
  assign n18724 = ~n18709 & n18723;
  assign n18725 = ~pi39 & n18567;
  assign n18726 = ~pi38 & ~n18725;
  assign n18727 = ~n18724 & n18726;
  assign n18728 = ~pi39 & ~n18659;
  assign n18729 = n18688 & ~n18728;
  assign n18730 = n3268 & ~n18729;
  assign n18731 = ~n18727 & n18730;
  assign n18732 = ~n18527 & ~n18731;
  assign n18733 = ~pi625 & n18732;
  assign n18734 = pi1153 & ~n18733;
  assign n18735 = ~n18696 & n18734;
  assign n18736 = ~pi142 & ~n17390;
  assign n18737 = pi142 & ~n17430;
  assign n18738 = ~n18736 & ~n18737;
  assign n18739 = pi735 & ~n18738;
  assign n18740 = ~pi735 & ~n18625;
  assign n18741 = ~n18739 & ~n18740;
  assign n18742 = n6223 & n18741;
  assign n18743 = ~pi142 & n17394;
  assign n18744 = pi142 & n17436;
  assign n18745 = ~n18743 & ~n18744;
  assign n18746 = pi735 & ~n18745;
  assign n18747 = ~pi735 & ~n18641;
  assign n18748 = ~n18746 & ~n18747;
  assign n18749 = ~n6223 & n18748;
  assign n18750 = ~n3461 & ~n18749;
  assign n18751 = ~n18742 & n18750;
  assign n18752 = pi735 & n17153;
  assign n18753 = n16660 & n18752;
  assign n18754 = ~n18652 & ~n18753;
  assign n18755 = n3461 & n18754;
  assign n18756 = ~pi215 & ~n18755;
  assign n18757 = ~n18751 & n18756;
  assign n18758 = ~pi735 & ~n18581;
  assign n18759 = pi142 & ~n17449;
  assign n18760 = ~pi142 & n17212;
  assign n18761 = n17211 & n18760;
  assign n18762 = pi735 & ~n18761;
  assign n18763 = ~n18759 & n18762;
  assign n18764 = ~n18758 & ~n18763;
  assign n18765 = ~n6223 & ~n18764;
  assign n18766 = ~pi735 & ~n18600;
  assign n18767 = pi142 & ~n17445;
  assign n18768 = pi735 & ~n18760;
  assign n18769 = ~n18767 & n18768;
  assign n18770 = ~n18766 & ~n18769;
  assign n18771 = n6223 & ~n18770;
  assign n18772 = pi215 & ~n18771;
  assign n18773 = ~n18765 & n18772;
  assign n18774 = pi299 & ~n18773;
  assign n18775 = ~n18757 & n18774;
  assign n18776 = n6197 & n18741;
  assign n18777 = ~n6197 & n18748;
  assign n18778 = ~n3053 & ~n18777;
  assign n18779 = ~n18776 & n18778;
  assign n18780 = n3053 & n18754;
  assign n18781 = ~pi223 & ~n18780;
  assign n18782 = ~n18779 & n18781;
  assign n18783 = ~n6197 & ~n18764;
  assign n18784 = n6197 & ~n18770;
  assign n18785 = pi223 & ~n18784;
  assign n18786 = ~n18783 & n18785;
  assign n18787 = ~pi299 & ~n18786;
  assign n18788 = ~n18782 & n18787;
  assign n18789 = pi39 & ~n18775;
  assign n18790 = ~n18788 & n18789;
  assign n18791 = ~pi142 & ~n17350;
  assign n18792 = pi142 & n17315;
  assign n18793 = pi735 & ~n18791;
  assign n18794 = ~n18792 & n18793;
  assign n18795 = pi142 & ~pi735;
  assign n18796 = ~n16655 & n18795;
  assign n18797 = ~n18794 & ~n18796;
  assign n18798 = ~pi39 & ~n18797;
  assign n18799 = ~pi38 & ~n18798;
  assign n18800 = ~n18790 & n18799;
  assign n18801 = n3096 & n18752;
  assign n18802 = ~n18656 & ~n18801;
  assign n18803 = ~pi39 & ~n18802;
  assign n18804 = n18688 & ~n18803;
  assign n18805 = n3268 & ~n18804;
  assign n18806 = ~n18800 & n18805;
  assign n18807 = ~n18527 & ~n18806;
  assign n18808 = ~pi625 & n18807;
  assign n18809 = n3268 & ~n17486;
  assign n18810 = pi142 & ~n18809;
  assign n18811 = pi39 & ~n16793;
  assign n18812 = pi142 & ~n18015;
  assign n18813 = ~n18811 & n18812;
  assign n18814 = ~n6223 & ~n18581;
  assign n18815 = n6223 & ~n18600;
  assign n18816 = pi215 & ~n18815;
  assign n18817 = ~n18814 & n18816;
  assign n18818 = ~n6223 & ~n18641;
  assign n18819 = n6223 & ~n18625;
  assign n18820 = ~n18818 & ~n18819;
  assign n18821 = ~n3461 & ~n18820;
  assign n18822 = n3461 & ~n18652;
  assign n18823 = ~pi215 & ~n18822;
  assign n18824 = ~n18821 & n18823;
  assign n18825 = ~n18817 & ~n18824;
  assign n18826 = pi39 & pi299;
  assign n18827 = ~n18825 & n18826;
  assign n18828 = ~n18813 & ~n18827;
  assign n18829 = n14819 & ~n18828;
  assign n18830 = ~n18810 & ~n18829;
  assign n18831 = pi625 & n18830;
  assign n18832 = ~pi1153 & ~n18831;
  assign n18833 = ~n18808 & n18832;
  assign n18834 = pi608 & ~n18833;
  assign n18835 = ~n18735 & n18834;
  assign n18836 = ~pi625 & n18695;
  assign n18837 = pi625 & n18732;
  assign n18838 = ~pi1153 & ~n18837;
  assign n18839 = ~n18836 & n18838;
  assign n18840 = pi625 & n18807;
  assign n18841 = ~pi625 & n18830;
  assign n18842 = pi1153 & ~n18841;
  assign n18843 = ~n18840 & n18842;
  assign n18844 = ~pi608 & ~n18843;
  assign n18845 = ~n18839 & n18844;
  assign n18846 = ~n18835 & ~n18845;
  assign n18847 = pi778 & ~n18846;
  assign n18848 = ~pi778 & n18695;
  assign n18849 = ~n18847 & ~n18848;
  assign n18850 = ~pi609 & ~n18849;
  assign n18851 = ~pi778 & ~n18807;
  assign n18852 = ~n18833 & ~n18843;
  assign n18853 = pi778 & ~n18852;
  assign n18854 = ~n18851 & ~n18853;
  assign n18855 = pi609 & n18854;
  assign n18856 = ~pi1155 & ~n18855;
  assign n18857 = ~n18850 & n18856;
  assign n18858 = ~n17527 & ~n18830;
  assign n18859 = ~n17526 & ~n18732;
  assign n18860 = pi609 & n18859;
  assign n18861 = ~n18858 & ~n18860;
  assign n18862 = pi1155 & ~n18861;
  assign n18863 = ~pi660 & ~n18862;
  assign n18864 = ~n18857 & n18863;
  assign n18865 = pi609 & ~n18849;
  assign n18866 = ~pi609 & n18854;
  assign n18867 = pi1155 & ~n18866;
  assign n18868 = ~n18865 & n18867;
  assign n18869 = ~n17539 & ~n18830;
  assign n18870 = ~pi609 & n18859;
  assign n18871 = ~n18869 & ~n18870;
  assign n18872 = ~pi1155 & ~n18871;
  assign n18873 = pi660 & ~n18872;
  assign n18874 = ~n18868 & n18873;
  assign n18875 = ~n18864 & ~n18874;
  assign n18876 = pi785 & ~n18875;
  assign n18877 = ~pi785 & ~n18849;
  assign n18878 = ~n18876 & ~n18877;
  assign n18879 = ~pi618 & ~n18878;
  assign n18880 = ~n17554 & n18854;
  assign n18881 = n17554 & n18830;
  assign n18882 = ~n18880 & ~n18881;
  assign n18883 = pi618 & ~n18882;
  assign n18884 = ~pi1154 & ~n18883;
  assign n18885 = ~n18879 & n18884;
  assign n18886 = n17526 & ~n18830;
  assign n18887 = ~n18859 & ~n18886;
  assign n18888 = ~pi785 & ~n18887;
  assign n18889 = ~n18862 & ~n18872;
  assign n18890 = pi785 & ~n18889;
  assign n18891 = ~n18888 & ~n18890;
  assign n18892 = pi618 & n18891;
  assign n18893 = ~pi618 & n18830;
  assign n18894 = pi1154 & ~n18893;
  assign n18895 = ~n18892 & n18894;
  assign n18896 = ~pi627 & ~n18895;
  assign n18897 = ~n18885 & n18896;
  assign n18898 = pi618 & ~n18878;
  assign n18899 = ~pi618 & ~n18882;
  assign n18900 = pi1154 & ~n18899;
  assign n18901 = ~n18898 & n18900;
  assign n18902 = ~pi618 & n18891;
  assign n18903 = pi618 & n18830;
  assign n18904 = ~pi1154 & ~n18903;
  assign n18905 = ~n18902 & n18904;
  assign n18906 = pi627 & ~n18905;
  assign n18907 = ~n18901 & n18906;
  assign n18908 = ~n18897 & ~n18907;
  assign n18909 = pi781 & ~n18908;
  assign n18910 = ~pi781 & ~n18878;
  assign n18911 = ~n18909 & ~n18910;
  assign n18912 = ~pi619 & ~n18911;
  assign n18913 = n17591 & ~n18830;
  assign n18914 = ~n17591 & n18882;
  assign n18915 = ~n18913 & ~n18914;
  assign n18916 = pi619 & n18915;
  assign n18917 = ~pi1159 & ~n18916;
  assign n18918 = ~n18912 & n18917;
  assign n18919 = ~pi781 & ~n18891;
  assign n18920 = ~n18895 & ~n18905;
  assign n18921 = pi781 & ~n18920;
  assign n18922 = ~n18919 & ~n18921;
  assign n18923 = pi619 & n18922;
  assign n18924 = ~pi619 & n18830;
  assign n18925 = pi1159 & ~n18924;
  assign n18926 = ~n18923 & n18925;
  assign n18927 = ~pi648 & ~n18926;
  assign n18928 = ~n18918 & n18927;
  assign n18929 = pi619 & ~n18911;
  assign n18930 = ~pi619 & n18915;
  assign n18931 = pi1159 & ~n18930;
  assign n18932 = ~n18929 & n18931;
  assign n18933 = ~pi619 & n18922;
  assign n18934 = pi619 & n18830;
  assign n18935 = ~pi1159 & ~n18934;
  assign n18936 = ~n18933 & n18935;
  assign n18937 = pi648 & ~n18936;
  assign n18938 = ~n18932 & n18937;
  assign n18939 = ~n18928 & ~n18938;
  assign n18940 = pi789 & ~n18939;
  assign n18941 = ~pi789 & ~n18911;
  assign n18942 = ~n18940 & ~n18941;
  assign n18943 = ~pi788 & n18942;
  assign n18944 = ~pi626 & n18942;
  assign n18945 = ~n17627 & n18915;
  assign n18946 = n17627 & n18830;
  assign n18947 = ~n18945 & ~n18946;
  assign n18948 = pi626 & n18947;
  assign n18949 = ~pi641 & ~n18948;
  assign n18950 = ~n18944 & n18949;
  assign n18951 = ~pi789 & ~n18922;
  assign n18952 = ~n18926 & ~n18936;
  assign n18953 = pi789 & ~n18952;
  assign n18954 = ~n18951 & ~n18953;
  assign n18955 = ~pi626 & n18954;
  assign n18956 = pi626 & n18830;
  assign n18957 = ~pi1158 & ~n18956;
  assign n18958 = ~n18955 & n18957;
  assign n18959 = ~n17634 & ~n18958;
  assign n18960 = ~n18950 & ~n18959;
  assign n18961 = pi626 & n18942;
  assign n18962 = ~pi626 & n18947;
  assign n18963 = pi641 & ~n18962;
  assign n18964 = ~n18961 & n18963;
  assign n18965 = pi626 & n18954;
  assign n18966 = ~pi626 & n18830;
  assign n18967 = pi1158 & ~n18966;
  assign n18968 = ~n18965 & n18967;
  assign n18969 = ~n17649 & ~n18968;
  assign n18970 = ~n18964 & ~n18969;
  assign n18971 = ~n18960 & ~n18970;
  assign n18972 = pi788 & ~n18971;
  assign n18973 = ~n18943 & ~n18972;
  assign n18974 = ~pi628 & n18973;
  assign n18975 = ~n18958 & ~n18968;
  assign n18976 = pi788 & ~n18975;
  assign n18977 = ~pi788 & ~n18954;
  assign n18978 = ~n18976 & ~n18977;
  assign n18979 = pi628 & n18978;
  assign n18980 = ~pi1156 & ~n18979;
  assign n18981 = ~n18974 & n18980;
  assign n18982 = ~n17670 & ~n18947;
  assign n18983 = n17670 & n18830;
  assign n18984 = ~n18982 & ~n18983;
  assign n18985 = pi628 & ~n18984;
  assign n18986 = ~pi628 & n18830;
  assign n18987 = pi1156 & ~n18986;
  assign n18988 = ~n18985 & n18987;
  assign n18989 = ~pi629 & ~n18988;
  assign n18990 = ~n18981 & n18989;
  assign n18991 = pi628 & n18973;
  assign n18992 = ~pi628 & n18978;
  assign n18993 = pi1156 & ~n18992;
  assign n18994 = ~n18991 & n18993;
  assign n18995 = ~pi628 & ~n18984;
  assign n18996 = pi628 & n18830;
  assign n18997 = ~pi1156 & ~n18996;
  assign n18998 = ~n18995 & n18997;
  assign n18999 = pi629 & ~n18998;
  assign n19000 = ~n18994 & n18999;
  assign n19001 = ~n18990 & ~n19000;
  assign n19002 = pi792 & ~n19001;
  assign n19003 = ~pi792 & n18973;
  assign n19004 = ~n19002 & ~n19003;
  assign n19005 = ~pi647 & ~n19004;
  assign n19006 = ~n17698 & n18978;
  assign n19007 = n17698 & n18830;
  assign n19008 = ~n19006 & ~n19007;
  assign n19009 = pi647 & ~n19008;
  assign n19010 = ~pi1157 & ~n19009;
  assign n19011 = ~n19005 & n19010;
  assign n19012 = ~pi792 & n18984;
  assign n19013 = ~n18988 & ~n18998;
  assign n19014 = pi792 & ~n19013;
  assign n19015 = ~n19012 & ~n19014;
  assign n19016 = pi647 & n19015;
  assign n19017 = ~pi647 & n18830;
  assign n19018 = pi1157 & ~n19017;
  assign n19019 = ~n19016 & n19018;
  assign n19020 = ~pi630 & ~n19019;
  assign n19021 = ~n19011 & n19020;
  assign n19022 = pi647 & ~n19004;
  assign n19023 = ~pi647 & ~n19008;
  assign n19024 = pi1157 & ~n19023;
  assign n19025 = ~n19022 & n19024;
  assign n19026 = ~pi647 & n19015;
  assign n19027 = pi647 & n18830;
  assign n19028 = ~pi1157 & ~n19027;
  assign n19029 = ~n19026 & n19028;
  assign n19030 = pi630 & ~n19029;
  assign n19031 = ~n19025 & n19030;
  assign n19032 = ~n19021 & ~n19031;
  assign n19033 = pi787 & ~n19032;
  assign n19034 = ~pi787 & ~n19004;
  assign n19035 = ~n19033 & ~n19034;
  assign n19036 = pi644 & ~n19035;
  assign n19037 = ~pi787 & ~n19015;
  assign n19038 = ~n19019 & ~n19029;
  assign n19039 = pi787 & ~n19038;
  assign n19040 = ~n19037 & ~n19039;
  assign n19041 = ~pi644 & n19040;
  assign n19042 = pi715 & ~n19041;
  assign n19043 = ~n19036 & n19042;
  assign n19044 = n17740 & ~n18830;
  assign n19045 = ~n17740 & n19008;
  assign n19046 = ~n19044 & ~n19045;
  assign n19047 = pi644 & n19046;
  assign n19048 = ~pi644 & n18830;
  assign n19049 = ~pi715 & ~n19048;
  assign n19050 = ~n19047 & n19049;
  assign n19051 = pi1160 & ~n19050;
  assign n19052 = ~n19043 & n19051;
  assign n19053 = ~pi644 & ~n19035;
  assign n19054 = pi644 & n19040;
  assign n19055 = ~pi715 & ~n19054;
  assign n19056 = ~n19053 & n19055;
  assign n19057 = ~pi644 & n19046;
  assign n19058 = pi644 & n18830;
  assign n19059 = pi715 & ~n19058;
  assign n19060 = ~n19057 & n19059;
  assign n19061 = ~pi1160 & ~n19060;
  assign n19062 = ~n19056 & n19061;
  assign n19063 = pi790 & ~n19052;
  assign n19064 = ~n19062 & n19063;
  assign n19065 = ~pi790 & n19035;
  assign n19066 = n6294 & ~n19065;
  assign n19067 = ~n19064 & n19066;
  assign n19068 = ~pi142 & ~n6294;
  assign n19069 = ~pi57 & ~n19068;
  assign n19070 = ~n19067 & n19069;
  assign n19071 = pi57 & pi142;
  assign n19072 = ~pi832 & ~n19071;
  assign n19073 = ~n19070 & n19072;
  assign n19074 = ~n17526 & n18657;
  assign n19075 = pi609 & n19074;
  assign n19076 = pi142 & ~n2755;
  assign n19077 = pi1155 & ~n19076;
  assign n19078 = ~n19075 & n19077;
  assign n19079 = ~pi609 & n19074;
  assign n19080 = ~pi1155 & ~n19076;
  assign n19081 = ~n19079 & n19080;
  assign n19082 = ~n19078 & ~n19081;
  assign n19083 = pi785 & ~n19082;
  assign n19084 = ~pi785 & ~n19076;
  assign n19085 = ~n19074 & n19084;
  assign n19086 = ~n19083 & ~n19085;
  assign n19087 = ~pi781 & ~n19086;
  assign n19088 = pi618 & n19086;
  assign n19089 = ~pi618 & n19076;
  assign n19090 = pi1154 & ~n19089;
  assign n19091 = ~n19088 & n19090;
  assign n19092 = ~pi618 & n19086;
  assign n19093 = pi618 & n19076;
  assign n19094 = ~pi1154 & ~n19093;
  assign n19095 = ~n19092 & n19094;
  assign n19096 = ~n19091 & ~n19095;
  assign n19097 = pi781 & ~n19096;
  assign n19098 = ~n19087 & ~n19097;
  assign n19099 = ~pi789 & ~n19098;
  assign n19100 = pi619 & n19098;
  assign n19101 = ~pi619 & n19076;
  assign n19102 = pi1159 & ~n19101;
  assign n19103 = ~n19100 & n19102;
  assign n19104 = ~pi619 & n19098;
  assign n19105 = pi619 & n19076;
  assign n19106 = ~pi1159 & ~n19105;
  assign n19107 = ~n19104 & n19106;
  assign n19108 = ~n19103 & ~n19107;
  assign n19109 = pi789 & ~n19108;
  assign n19110 = ~n19099 & ~n19109;
  assign n19111 = pi626 & n19110;
  assign n19112 = ~pi626 & n19076;
  assign n19113 = pi1158 & ~n19112;
  assign n19114 = ~n19111 & n19113;
  assign n19115 = ~pi626 & n19110;
  assign n19116 = pi626 & n19076;
  assign n19117 = ~pi1158 & ~n19116;
  assign n19118 = ~n19115 & n19117;
  assign n19119 = ~n19114 & ~n19118;
  assign n19120 = ~n17669 & n19119;
  assign n19121 = ~pi625 & pi1153;
  assign n19122 = pi625 & ~pi1153;
  assign n19123 = ~n19121 & ~n19122;
  assign n19124 = pi778 & ~n19123;
  assign n19125 = n18752 & ~n19124;
  assign n19126 = ~n19076 & ~n19125;
  assign n19127 = ~n17554 & ~n19126;
  assign n19128 = ~n17591 & n19127;
  assign n19129 = ~n19076 & ~n19128;
  assign n19130 = n17627 & ~n19076;
  assign n19131 = n17792 & ~n19130;
  assign n19132 = ~n19129 & n19131;
  assign n19133 = ~n19120 & ~n19132;
  assign n19134 = pi788 & ~n19133;
  assign n19135 = pi735 & n17154;
  assign n19136 = pi625 & n19135;
  assign n19137 = ~n18657 & ~n19076;
  assign n19138 = ~n19135 & n19137;
  assign n19139 = ~n19136 & ~n19138;
  assign n19140 = ~pi1153 & ~n19139;
  assign n19141 = pi625 & n18752;
  assign n19142 = pi1153 & ~n19076;
  assign n19143 = ~n19141 & n19142;
  assign n19144 = ~pi608 & ~n19143;
  assign n19145 = ~n19140 & n19144;
  assign n19146 = ~n18657 & ~n19136;
  assign n19147 = pi1153 & ~n19146;
  assign n19148 = ~pi625 & ~pi1153;
  assign n19149 = n18752 & n19148;
  assign n19150 = ~n19076 & ~n19149;
  assign n19151 = ~n19147 & n19150;
  assign n19152 = pi608 & ~n19151;
  assign n19153 = ~n19145 & ~n19152;
  assign n19154 = pi778 & ~n19153;
  assign n19155 = ~pi778 & ~n19138;
  assign n19156 = ~n19154 & ~n19155;
  assign n19157 = ~pi609 & ~n19156;
  assign n19158 = pi609 & ~n19126;
  assign n19159 = ~pi1155 & ~n19158;
  assign n19160 = ~n19157 & n19159;
  assign n19161 = ~pi660 & ~n19078;
  assign n19162 = ~n19160 & n19161;
  assign n19163 = pi609 & ~n19156;
  assign n19164 = ~pi609 & ~n19126;
  assign n19165 = pi1155 & ~n19164;
  assign n19166 = ~n19163 & n19165;
  assign n19167 = pi660 & ~n19081;
  assign n19168 = ~n19166 & n19167;
  assign n19169 = ~n19162 & ~n19168;
  assign n19170 = pi785 & ~n19169;
  assign n19171 = ~pi785 & ~n19156;
  assign n19172 = ~n19170 & ~n19171;
  assign n19173 = ~pi618 & ~n19172;
  assign n19174 = ~n19076 & ~n19127;
  assign n19175 = pi618 & ~n19174;
  assign n19176 = ~pi1154 & ~n19175;
  assign n19177 = ~n19173 & n19176;
  assign n19178 = ~pi627 & ~n19091;
  assign n19179 = ~n19177 & n19178;
  assign n19180 = pi618 & ~n19172;
  assign n19181 = ~pi618 & ~n19174;
  assign n19182 = pi1154 & ~n19181;
  assign n19183 = ~n19180 & n19182;
  assign n19184 = pi627 & ~n19095;
  assign n19185 = ~n19183 & n19184;
  assign n19186 = ~n19179 & ~n19185;
  assign n19187 = pi781 & ~n19186;
  assign n19188 = ~pi781 & ~n19172;
  assign n19189 = ~n19187 & ~n19188;
  assign n19190 = ~pi619 & ~n19189;
  assign n19191 = pi619 & ~n19129;
  assign n19192 = ~pi1159 & ~n19191;
  assign n19193 = ~n19190 & n19192;
  assign n19194 = ~pi648 & ~n19103;
  assign n19195 = ~n19193 & n19194;
  assign n19196 = pi619 & ~n19189;
  assign n19197 = ~pi619 & ~n19129;
  assign n19198 = pi1159 & ~n19197;
  assign n19199 = ~n19196 & n19198;
  assign n19200 = pi648 & ~n19107;
  assign n19201 = ~n19199 & n19200;
  assign n19202 = pi789 & ~n19195;
  assign n19203 = ~n19201 & n19202;
  assign n19204 = ~pi789 & n19189;
  assign n19205 = n17905 & ~n19204;
  assign n19206 = ~n19203 & n19205;
  assign n19207 = ~n19134 & ~n19206;
  assign n19208 = ~pi628 & n19207;
  assign n19209 = ~pi788 & ~n19110;
  assign n19210 = pi788 & ~n19119;
  assign n19211 = ~n19209 & ~n19210;
  assign n19212 = pi628 & ~n19211;
  assign n19213 = ~pi1156 & ~n19212;
  assign n19214 = ~n19208 & n19213;
  assign n19215 = ~n17627 & ~n17670;
  assign n19216 = ~n17554 & ~n17591;
  assign n19217 = n19215 & n19216;
  assign n19218 = ~n19126 & n19217;
  assign n19219 = pi628 & n19218;
  assign n19220 = ~n19076 & ~n19219;
  assign n19221 = pi1156 & ~n19220;
  assign n19222 = ~pi629 & ~n19221;
  assign n19223 = ~n19214 & n19222;
  assign n19224 = pi628 & n19207;
  assign n19225 = ~pi628 & ~n19211;
  assign n19226 = pi1156 & ~n19225;
  assign n19227 = ~n19224 & n19226;
  assign n19228 = ~pi628 & n19218;
  assign n19229 = ~n19076 & ~n19228;
  assign n19230 = ~pi1156 & ~n19229;
  assign n19231 = pi629 & ~n19230;
  assign n19232 = ~n19227 & n19231;
  assign n19233 = ~n19223 & ~n19232;
  assign n19234 = pi792 & ~n19233;
  assign n19235 = ~pi792 & n19207;
  assign n19236 = ~n19234 & ~n19235;
  assign n19237 = ~pi647 & n19236;
  assign n19238 = ~n17698 & n19211;
  assign n19239 = n17698 & n19076;
  assign n19240 = ~n19238 & ~n19239;
  assign n19241 = pi647 & ~n19240;
  assign n19242 = ~pi1157 & ~n19241;
  assign n19243 = ~n19237 & n19242;
  assign n19244 = pi628 & pi1156;
  assign n19245 = ~pi628 & ~pi1156;
  assign n19246 = pi792 & ~n19244;
  assign n19247 = ~n19245 & n19246;
  assign n19248 = n19218 & ~n19247;
  assign n19249 = pi647 & n19248;
  assign n19250 = pi1157 & ~n19076;
  assign n19251 = ~n19249 & n19250;
  assign n19252 = ~pi630 & ~n19251;
  assign n19253 = ~n19243 & n19252;
  assign n19254 = pi647 & n19236;
  assign n19255 = ~pi647 & ~n19240;
  assign n19256 = pi1157 & ~n19255;
  assign n19257 = ~n19254 & n19256;
  assign n19258 = ~pi647 & n19248;
  assign n19259 = ~pi1157 & ~n19076;
  assign n19260 = ~n19258 & n19259;
  assign n19261 = pi630 & ~n19260;
  assign n19262 = ~n19257 & n19261;
  assign n19263 = ~n19253 & ~n19262;
  assign n19264 = pi787 & ~n19263;
  assign n19265 = ~pi787 & n19236;
  assign n19266 = ~n19264 & ~n19265;
  assign n19267 = pi644 & ~n19266;
  assign n19268 = ~pi647 & pi1157;
  assign n19269 = pi647 & ~pi1157;
  assign n19270 = ~n19268 & ~n19269;
  assign n19271 = pi787 & ~n19270;
  assign n19272 = n19248 & ~n19271;
  assign n19273 = ~n19076 & ~n19272;
  assign n19274 = ~pi644 & ~n19273;
  assign n19275 = pi715 & ~n19274;
  assign n19276 = ~n19267 & n19275;
  assign n19277 = n17740 & ~n19076;
  assign n19278 = ~n17740 & n19240;
  assign n19279 = ~n19277 & ~n19278;
  assign n19280 = pi644 & n19279;
  assign n19281 = ~pi644 & n19076;
  assign n19282 = ~pi715 & ~n19281;
  assign n19283 = ~n19280 & n19282;
  assign n19284 = pi1160 & ~n19283;
  assign n19285 = ~n19276 & n19284;
  assign n19286 = ~pi644 & ~n19266;
  assign n19287 = pi644 & ~n19273;
  assign n19288 = ~pi715 & ~n19287;
  assign n19289 = ~n19286 & n19288;
  assign n19290 = ~pi644 & n19279;
  assign n19291 = pi644 & n19076;
  assign n19292 = pi715 & ~n19291;
  assign n19293 = ~n19290 & n19292;
  assign n19294 = ~pi1160 & ~n19293;
  assign n19295 = ~n19289 & n19294;
  assign n19296 = ~n19285 & ~n19295;
  assign n19297 = pi790 & ~n19296;
  assign n19298 = ~pi790 & ~n19266;
  assign n19299 = pi832 & ~n19298;
  assign n19300 = ~n19297 & n19299;
  assign po299 = ~n19073 & ~n19300;
  assign n19302 = pi143 & ~n3268;
  assign n19303 = n16968 & ~n17054;
  assign n19304 = pi38 & n19303;
  assign n19305 = pi39 & ~n17074;
  assign n19306 = ~pi39 & ~n17317;
  assign n19307 = ~n19305 & ~n19306;
  assign n19308 = ~pi38 & ~n19307;
  assign n19309 = ~n19304 & ~n19308;
  assign n19310 = ~pi143 & n19309;
  assign n19311 = ~pi39 & ~n17340;
  assign n19312 = pi39 & ~n17166;
  assign n19313 = ~n19311 & ~n19312;
  assign n19314 = ~pi38 & n19313;
  assign n19315 = pi143 & n19314;
  assign n19316 = pi38 & n18045;
  assign n19317 = pi774 & ~n19316;
  assign n19318 = ~n19315 & n19317;
  assign n19319 = ~n19310 & n19318;
  assign n19320 = n6250 & ~n17155;
  assign n19321 = pi38 & ~n19320;
  assign n19322 = pi39 & ~n17233;
  assign n19323 = n16919 & ~n17350;
  assign n19324 = ~n19322 & ~n19323;
  assign n19325 = ~pi38 & ~n19324;
  assign n19326 = ~n19321 & ~n19325;
  assign n19327 = pi143 & n19326;
  assign n19328 = pi39 & ~n17295;
  assign n19329 = ~pi39 & ~n17344;
  assign n19330 = ~pi38 & n19329;
  assign n19331 = ~pi39 & n17259;
  assign n19332 = pi38 & ~n19331;
  assign n19333 = ~n19330 & ~n19332;
  assign n19334 = ~n19328 & n19333;
  assign n19335 = ~pi143 & ~n19334;
  assign n19336 = ~pi774 & ~n19335;
  assign n19337 = ~n19327 & n19336;
  assign n19338 = pi687 & ~n19337;
  assign n19339 = ~n19319 & n19338;
  assign n19340 = ~pi143 & ~n17487;
  assign n19341 = pi774 & ~n19340;
  assign n19342 = n6117 & n16933;
  assign n19343 = pi38 & n19342;
  assign n19344 = ~pi38 & n16963;
  assign n19345 = pi143 & ~n19344;
  assign n19346 = ~pi38 & ~n16907;
  assign n19347 = n6250 & n16879;
  assign n19348 = pi38 & ~n19347;
  assign n19349 = ~n19346 & ~n19348;
  assign n19350 = ~pi143 & ~pi774;
  assign n19351 = n19349 & n19350;
  assign n19352 = ~n19345 & ~n19351;
  assign n19353 = ~n19343 & ~n19352;
  assign n19354 = ~n19341 & ~n19353;
  assign n19355 = ~pi687 & n19354;
  assign n19356 = n3268 & ~n19339;
  assign n19357 = ~n19355 & n19356;
  assign n19358 = ~n19302 & ~n19357;
  assign n19359 = ~pi625 & n19358;
  assign n19360 = n3268 & ~n19354;
  assign n19361 = ~n19302 & ~n19360;
  assign n19362 = pi625 & n19361;
  assign n19363 = ~pi1153 & ~n19362;
  assign n19364 = ~n19359 & n19363;
  assign n19365 = ~pi687 & n19340;
  assign n19366 = ~pi143 & n18060;
  assign n19367 = pi143 & ~n18064;
  assign n19368 = ~pi38 & ~n19367;
  assign n19369 = ~n19366 & n19368;
  assign n19370 = ~pi143 & ~n16968;
  assign n19371 = n17480 & ~n19370;
  assign n19372 = pi687 & ~n19371;
  assign n19373 = ~n19369 & n19372;
  assign n19374 = n3268 & ~n19365;
  assign n19375 = ~n19373 & n19374;
  assign n19376 = ~n19302 & ~n19375;
  assign n19377 = pi625 & n19376;
  assign n19378 = ~pi143 & ~n17494;
  assign n19379 = ~pi625 & n19378;
  assign n19380 = pi1153 & ~n19379;
  assign n19381 = ~n19377 & n19380;
  assign n19382 = ~pi608 & ~n19381;
  assign n19383 = ~n19364 & n19382;
  assign n19384 = pi625 & n19358;
  assign n19385 = ~pi625 & n19361;
  assign n19386 = pi1153 & ~n19385;
  assign n19387 = ~n19384 & n19386;
  assign n19388 = ~pi625 & n19376;
  assign n19389 = pi625 & n19378;
  assign n19390 = ~pi1153 & ~n19389;
  assign n19391 = ~n19388 & n19390;
  assign n19392 = pi608 & ~n19391;
  assign n19393 = ~n19387 & n19392;
  assign n19394 = ~n19383 & ~n19393;
  assign n19395 = pi778 & ~n19394;
  assign n19396 = ~pi778 & n19358;
  assign n19397 = ~n19395 & ~n19396;
  assign n19398 = ~pi609 & ~n19397;
  assign n19399 = ~pi778 & ~n19376;
  assign n19400 = ~n19381 & ~n19391;
  assign n19401 = pi778 & ~n19400;
  assign n19402 = ~n19399 & ~n19401;
  assign n19403 = pi609 & n19402;
  assign n19404 = ~pi1155 & ~n19403;
  assign n19405 = ~n19398 & n19404;
  assign n19406 = ~n17527 & ~n19378;
  assign n19407 = ~n17526 & ~n19361;
  assign n19408 = pi609 & n19407;
  assign n19409 = ~n19406 & ~n19408;
  assign n19410 = pi1155 & ~n19409;
  assign n19411 = ~pi660 & ~n19410;
  assign n19412 = ~n19405 & n19411;
  assign n19413 = pi609 & ~n19397;
  assign n19414 = ~pi609 & n19402;
  assign n19415 = pi1155 & ~n19414;
  assign n19416 = ~n19413 & n19415;
  assign n19417 = ~n17539 & ~n19378;
  assign n19418 = ~pi609 & n19407;
  assign n19419 = ~n19417 & ~n19418;
  assign n19420 = ~pi1155 & ~n19419;
  assign n19421 = pi660 & ~n19420;
  assign n19422 = ~n19416 & n19421;
  assign n19423 = ~n19412 & ~n19422;
  assign n19424 = pi785 & ~n19423;
  assign n19425 = ~pi785 & ~n19397;
  assign n19426 = ~n19424 & ~n19425;
  assign n19427 = ~pi618 & ~n19426;
  assign n19428 = ~n17554 & ~n19402;
  assign n19429 = n17554 & ~n19378;
  assign n19430 = ~n19428 & ~n19429;
  assign n19431 = pi618 & n19430;
  assign n19432 = ~pi1154 & ~n19431;
  assign n19433 = ~n19427 & n19432;
  assign n19434 = n17526 & ~n19378;
  assign n19435 = ~n19407 & ~n19434;
  assign n19436 = ~pi785 & ~n19435;
  assign n19437 = ~n19410 & ~n19420;
  assign n19438 = pi785 & ~n19437;
  assign n19439 = ~n19436 & ~n19438;
  assign n19440 = pi618 & n19439;
  assign n19441 = ~pi618 & n19378;
  assign n19442 = pi1154 & ~n19441;
  assign n19443 = ~n19440 & n19442;
  assign n19444 = ~pi627 & ~n19443;
  assign n19445 = ~n19433 & n19444;
  assign n19446 = pi618 & ~n19426;
  assign n19447 = ~pi618 & n19430;
  assign n19448 = pi1154 & ~n19447;
  assign n19449 = ~n19446 & n19448;
  assign n19450 = ~pi618 & n19439;
  assign n19451 = pi618 & n19378;
  assign n19452 = ~pi1154 & ~n19451;
  assign n19453 = ~n19450 & n19452;
  assign n19454 = pi627 & ~n19453;
  assign n19455 = ~n19449 & n19454;
  assign n19456 = ~n19445 & ~n19455;
  assign n19457 = pi781 & ~n19456;
  assign n19458 = ~pi781 & ~n19426;
  assign n19459 = ~n19457 & ~n19458;
  assign n19460 = ~pi619 & ~n19459;
  assign n19461 = ~n17591 & n19430;
  assign n19462 = n17591 & n19378;
  assign n19463 = ~n19461 & ~n19462;
  assign n19464 = pi619 & ~n19463;
  assign n19465 = ~pi1159 & ~n19464;
  assign n19466 = ~n19460 & n19465;
  assign n19467 = ~pi781 & ~n19439;
  assign n19468 = ~n19443 & ~n19453;
  assign n19469 = pi781 & ~n19468;
  assign n19470 = ~n19467 & ~n19469;
  assign n19471 = pi619 & n19470;
  assign n19472 = ~pi619 & n19378;
  assign n19473 = pi1159 & ~n19472;
  assign n19474 = ~n19471 & n19473;
  assign n19475 = ~pi648 & ~n19474;
  assign n19476 = ~n19466 & n19475;
  assign n19477 = pi619 & ~n19459;
  assign n19478 = ~pi619 & ~n19463;
  assign n19479 = pi1159 & ~n19478;
  assign n19480 = ~n19477 & n19479;
  assign n19481 = ~pi619 & n19470;
  assign n19482 = pi619 & n19378;
  assign n19483 = ~pi1159 & ~n19482;
  assign n19484 = ~n19481 & n19483;
  assign n19485 = pi648 & ~n19484;
  assign n19486 = ~n19480 & n19485;
  assign n19487 = ~n19476 & ~n19486;
  assign n19488 = pi789 & ~n19487;
  assign n19489 = ~pi789 & ~n19459;
  assign n19490 = ~n19488 & ~n19489;
  assign n19491 = ~pi788 & n19490;
  assign n19492 = ~pi626 & n19490;
  assign n19493 = n17627 & ~n19378;
  assign n19494 = ~n17627 & n19463;
  assign n19495 = ~n19493 & ~n19494;
  assign n19496 = pi626 & ~n19495;
  assign n19497 = ~pi641 & ~n19496;
  assign n19498 = ~n19492 & n19497;
  assign n19499 = ~pi789 & ~n19470;
  assign n19500 = ~n19474 & ~n19484;
  assign n19501 = pi789 & ~n19500;
  assign n19502 = ~n19499 & ~n19501;
  assign n19503 = ~pi626 & n19502;
  assign n19504 = pi626 & n19378;
  assign n19505 = ~pi1158 & ~n19504;
  assign n19506 = ~n19503 & n19505;
  assign n19507 = ~n17634 & ~n19506;
  assign n19508 = ~n19498 & ~n19507;
  assign n19509 = pi626 & n19490;
  assign n19510 = ~pi626 & ~n19495;
  assign n19511 = pi641 & ~n19510;
  assign n19512 = ~n19509 & n19511;
  assign n19513 = pi626 & n19502;
  assign n19514 = ~pi626 & n19378;
  assign n19515 = pi1158 & ~n19514;
  assign n19516 = ~n19513 & n19515;
  assign n19517 = ~n17649 & ~n19516;
  assign n19518 = ~n19512 & ~n19517;
  assign n19519 = ~n19508 & ~n19518;
  assign n19520 = pi788 & ~n19519;
  assign n19521 = ~n19491 & ~n19520;
  assign n19522 = ~pi628 & n19521;
  assign n19523 = ~n19506 & ~n19516;
  assign n19524 = pi788 & ~n19523;
  assign n19525 = ~pi788 & ~n19502;
  assign n19526 = ~n19524 & ~n19525;
  assign n19527 = pi628 & n19526;
  assign n19528 = ~pi1156 & ~n19527;
  assign n19529 = ~n19522 & n19528;
  assign n19530 = ~n17670 & n19495;
  assign n19531 = n17670 & n19378;
  assign n19532 = ~n19530 & ~n19531;
  assign n19533 = pi628 & ~n19532;
  assign n19534 = ~pi628 & n19378;
  assign n19535 = pi1156 & ~n19534;
  assign n19536 = ~n19533 & n19535;
  assign n19537 = ~pi629 & ~n19536;
  assign n19538 = ~n19529 & n19537;
  assign n19539 = pi628 & n19521;
  assign n19540 = ~pi628 & n19526;
  assign n19541 = pi1156 & ~n19540;
  assign n19542 = ~n19539 & n19541;
  assign n19543 = ~pi628 & ~n19532;
  assign n19544 = pi628 & n19378;
  assign n19545 = ~pi1156 & ~n19544;
  assign n19546 = ~n19543 & n19545;
  assign n19547 = pi629 & ~n19546;
  assign n19548 = ~n19542 & n19547;
  assign n19549 = ~n19538 & ~n19548;
  assign n19550 = pi792 & ~n19549;
  assign n19551 = ~pi792 & n19521;
  assign n19552 = ~n19550 & ~n19551;
  assign n19553 = ~pi647 & ~n19552;
  assign n19554 = ~n17698 & n19526;
  assign n19555 = n17698 & n19378;
  assign n19556 = ~n19554 & ~n19555;
  assign n19557 = pi647 & ~n19556;
  assign n19558 = ~pi1157 & ~n19557;
  assign n19559 = ~n19553 & n19558;
  assign n19560 = ~pi792 & n19532;
  assign n19561 = ~n19536 & ~n19546;
  assign n19562 = pi792 & ~n19561;
  assign n19563 = ~n19560 & ~n19562;
  assign n19564 = pi647 & n19563;
  assign n19565 = ~pi647 & n19378;
  assign n19566 = pi1157 & ~n19565;
  assign n19567 = ~n19564 & n19566;
  assign n19568 = ~pi630 & ~n19567;
  assign n19569 = ~n19559 & n19568;
  assign n19570 = pi647 & ~n19552;
  assign n19571 = ~pi647 & ~n19556;
  assign n19572 = pi1157 & ~n19571;
  assign n19573 = ~n19570 & n19572;
  assign n19574 = ~pi647 & n19563;
  assign n19575 = pi647 & n19378;
  assign n19576 = ~pi1157 & ~n19575;
  assign n19577 = ~n19574 & n19576;
  assign n19578 = pi630 & ~n19577;
  assign n19579 = ~n19573 & n19578;
  assign n19580 = ~n19569 & ~n19579;
  assign n19581 = pi787 & ~n19580;
  assign n19582 = ~pi787 & ~n19552;
  assign n19583 = ~n19581 & ~n19582;
  assign n19584 = pi644 & ~n19583;
  assign n19585 = ~pi787 & ~n19563;
  assign n19586 = ~n19567 & ~n19577;
  assign n19587 = pi787 & ~n19586;
  assign n19588 = ~n19585 & ~n19587;
  assign n19589 = ~pi644 & n19588;
  assign n19590 = pi715 & ~n19589;
  assign n19591 = ~n19584 & n19590;
  assign n19592 = n17740 & ~n19378;
  assign n19593 = ~n17740 & n19556;
  assign n19594 = ~n19592 & ~n19593;
  assign n19595 = pi644 & n19594;
  assign n19596 = ~pi644 & n19378;
  assign n19597 = ~pi715 & ~n19596;
  assign n19598 = ~n19595 & n19597;
  assign n19599 = pi1160 & ~n19598;
  assign n19600 = ~n19591 & n19599;
  assign n19601 = ~pi644 & ~n19583;
  assign n19602 = pi644 & n19588;
  assign n19603 = ~pi715 & ~n19602;
  assign n19604 = ~n19601 & n19603;
  assign n19605 = ~pi644 & n19594;
  assign n19606 = pi644 & n19378;
  assign n19607 = pi715 & ~n19606;
  assign n19608 = ~n19605 & n19607;
  assign n19609 = ~pi1160 & ~n19608;
  assign n19610 = ~n19604 & n19609;
  assign n19611 = pi790 & ~n19600;
  assign n19612 = ~n19610 & n19611;
  assign n19613 = ~pi790 & n19583;
  assign n19614 = ~po1038 & ~n19613;
  assign n19615 = ~n19612 & n19614;
  assign n19616 = ~pi143 & po1038;
  assign n19617 = ~pi832 & ~n19616;
  assign n19618 = ~n19615 & n19617;
  assign n19619 = ~pi143 & ~n2755;
  assign n19620 = pi687 & n17153;
  assign n19621 = ~n19619 & ~n19620;
  assign n19622 = ~pi778 & n19621;
  assign n19623 = ~pi625 & n19620;
  assign n19624 = ~n19621 & ~n19623;
  assign n19625 = pi1153 & ~n19624;
  assign n19626 = ~pi1153 & ~n19619;
  assign n19627 = ~n19623 & n19626;
  assign n19628 = ~n19625 & ~n19627;
  assign n19629 = pi778 & ~n19628;
  assign n19630 = ~n19622 & ~n19629;
  assign n19631 = ~n17780 & n19630;
  assign n19632 = ~n17782 & n19631;
  assign n19633 = ~n17784 & n19632;
  assign n19634 = n17792 & n19633;
  assign n19635 = ~pi774 & n16933;
  assign n19636 = ~n19619 & ~n19635;
  assign n19637 = ~n17794 & ~n19636;
  assign n19638 = ~pi785 & ~n19637;
  assign n19639 = ~n17799 & ~n19636;
  assign n19640 = pi1155 & ~n19639;
  assign n19641 = ~n17802 & n19637;
  assign n19642 = ~pi1155 & ~n19641;
  assign n19643 = ~n19640 & ~n19642;
  assign n19644 = pi785 & ~n19643;
  assign n19645 = ~n19638 & ~n19644;
  assign n19646 = ~pi781 & ~n19645;
  assign n19647 = ~n17809 & n19645;
  assign n19648 = pi1154 & ~n19647;
  assign n19649 = ~n17812 & n19645;
  assign n19650 = ~pi1154 & ~n19649;
  assign n19651 = ~n19648 & ~n19650;
  assign n19652 = pi781 & ~n19651;
  assign n19653 = ~n19646 & ~n19652;
  assign n19654 = ~pi789 & ~n19653;
  assign n19655 = pi619 & n19653;
  assign n19656 = ~pi619 & n19619;
  assign n19657 = pi1159 & ~n19656;
  assign n19658 = ~n19655 & n19657;
  assign n19659 = ~pi619 & n19653;
  assign n19660 = pi619 & n19619;
  assign n19661 = ~pi1159 & ~n19660;
  assign n19662 = ~n19659 & n19661;
  assign n19663 = ~n19658 & ~n19662;
  assign n19664 = pi789 & ~n19663;
  assign n19665 = ~n19654 & ~n19664;
  assign n19666 = pi626 & n19665;
  assign n19667 = ~pi626 & n19619;
  assign n19668 = pi1158 & ~n19667;
  assign n19669 = ~n19666 & n19668;
  assign n19670 = ~pi626 & n19665;
  assign n19671 = pi626 & n19619;
  assign n19672 = ~pi1158 & ~n19671;
  assign n19673 = ~n19670 & n19672;
  assign n19674 = ~n19669 & ~n19673;
  assign n19675 = ~n17669 & n19674;
  assign n19676 = ~n19634 & ~n19675;
  assign n19677 = pi788 & ~n19676;
  assign n19678 = ~n16842 & ~n19621;
  assign n19679 = pi625 & n19678;
  assign n19680 = n19636 & ~n19678;
  assign n19681 = ~n19679 & ~n19680;
  assign n19682 = n19626 & ~n19681;
  assign n19683 = ~pi608 & ~n19625;
  assign n19684 = ~n19682 & n19683;
  assign n19685 = pi1153 & n19636;
  assign n19686 = ~n19679 & n19685;
  assign n19687 = pi608 & ~n19627;
  assign n19688 = ~n19686 & n19687;
  assign n19689 = ~n19684 & ~n19688;
  assign n19690 = pi778 & ~n19689;
  assign n19691 = ~pi778 & ~n19680;
  assign n19692 = ~n19690 & ~n19691;
  assign n19693 = ~pi609 & ~n19692;
  assign n19694 = pi609 & n19630;
  assign n19695 = ~pi1155 & ~n19694;
  assign n19696 = ~n19693 & n19695;
  assign n19697 = ~pi660 & ~n19640;
  assign n19698 = ~n19696 & n19697;
  assign n19699 = pi609 & ~n19692;
  assign n19700 = ~pi609 & n19630;
  assign n19701 = pi1155 & ~n19700;
  assign n19702 = ~n19699 & n19701;
  assign n19703 = pi660 & ~n19642;
  assign n19704 = ~n19702 & n19703;
  assign n19705 = ~n19698 & ~n19704;
  assign n19706 = pi785 & ~n19705;
  assign n19707 = ~pi785 & ~n19692;
  assign n19708 = ~n19706 & ~n19707;
  assign n19709 = ~pi618 & ~n19708;
  assign n19710 = pi618 & n19631;
  assign n19711 = ~pi1154 & ~n19710;
  assign n19712 = ~n19709 & n19711;
  assign n19713 = ~pi627 & ~n19648;
  assign n19714 = ~n19712 & n19713;
  assign n19715 = pi618 & ~n19708;
  assign n19716 = ~pi618 & n19631;
  assign n19717 = pi1154 & ~n19716;
  assign n19718 = ~n19715 & n19717;
  assign n19719 = pi627 & ~n19650;
  assign n19720 = ~n19718 & n19719;
  assign n19721 = ~n19714 & ~n19720;
  assign n19722 = pi781 & ~n19721;
  assign n19723 = ~pi781 & ~n19708;
  assign n19724 = ~n19722 & ~n19723;
  assign n19725 = ~pi619 & ~n19724;
  assign n19726 = pi619 & n19632;
  assign n19727 = ~pi1159 & ~n19726;
  assign n19728 = ~n19725 & n19727;
  assign n19729 = ~pi648 & ~n19658;
  assign n19730 = ~n19728 & n19729;
  assign n19731 = pi619 & ~n19724;
  assign n19732 = ~pi619 & n19632;
  assign n19733 = pi1159 & ~n19732;
  assign n19734 = ~n19731 & n19733;
  assign n19735 = pi648 & ~n19662;
  assign n19736 = ~n19734 & n19735;
  assign n19737 = pi789 & ~n19730;
  assign n19738 = ~n19736 & n19737;
  assign n19739 = ~pi789 & n19724;
  assign n19740 = n17905 & ~n19739;
  assign n19741 = ~n19738 & n19740;
  assign n19742 = ~n19677 & ~n19741;
  assign n19743 = ~pi628 & ~n19742;
  assign n19744 = ~pi788 & ~n19665;
  assign n19745 = pi788 & ~n19674;
  assign n19746 = ~n19744 & ~n19745;
  assign n19747 = pi628 & n19746;
  assign n19748 = ~pi1156 & ~n19747;
  assign n19749 = ~n19743 & n19748;
  assign n19750 = ~n17916 & n19633;
  assign n19751 = ~n17918 & n19750;
  assign n19752 = pi1156 & ~n19751;
  assign n19753 = ~pi629 & ~n19752;
  assign n19754 = ~n19749 & n19753;
  assign n19755 = pi628 & ~n19742;
  assign n19756 = ~pi628 & n19746;
  assign n19757 = pi1156 & ~n19756;
  assign n19758 = ~n19755 & n19757;
  assign n19759 = ~n17927 & n19750;
  assign n19760 = ~pi1156 & ~n19759;
  assign n19761 = pi629 & ~n19760;
  assign n19762 = ~n19758 & n19761;
  assign n19763 = ~n19754 & ~n19762;
  assign n19764 = pi792 & ~n19763;
  assign n19765 = ~pi792 & ~n19742;
  assign n19766 = ~n19764 & ~n19765;
  assign n19767 = ~pi647 & ~n19766;
  assign n19768 = ~n17698 & n19746;
  assign n19769 = n17698 & n19619;
  assign n19770 = ~n19768 & ~n19769;
  assign n19771 = pi647 & ~n19770;
  assign n19772 = ~pi1157 & ~n19771;
  assign n19773 = ~n19767 & n19772;
  assign n19774 = ~n17947 & n19750;
  assign n19775 = pi647 & n19774;
  assign n19776 = ~pi647 & n19619;
  assign n19777 = pi1157 & ~n19776;
  assign n19778 = ~n19775 & n19777;
  assign n19779 = ~pi630 & ~n19778;
  assign n19780 = ~n19773 & n19779;
  assign n19781 = pi647 & ~n19766;
  assign n19782 = ~pi647 & ~n19770;
  assign n19783 = pi1157 & ~n19782;
  assign n19784 = ~n19781 & n19783;
  assign n19785 = ~pi647 & n19774;
  assign n19786 = pi647 & n19619;
  assign n19787 = ~pi1157 & ~n19786;
  assign n19788 = ~n19785 & n19787;
  assign n19789 = pi630 & ~n19788;
  assign n19790 = ~n19784 & n19789;
  assign n19791 = ~n19780 & ~n19790;
  assign n19792 = pi787 & ~n19791;
  assign n19793 = ~pi787 & ~n19766;
  assign n19794 = ~n19792 & ~n19793;
  assign n19795 = pi644 & ~n19794;
  assign n19796 = ~pi787 & ~n19774;
  assign n19797 = ~n19778 & ~n19788;
  assign n19798 = pi787 & ~n19797;
  assign n19799 = ~n19796 & ~n19798;
  assign n19800 = ~pi644 & n19799;
  assign n19801 = pi715 & ~n19800;
  assign n19802 = ~n19795 & n19801;
  assign n19803 = n17740 & ~n19619;
  assign n19804 = ~n17740 & n19770;
  assign n19805 = ~n19803 & ~n19804;
  assign n19806 = pi644 & n19805;
  assign n19807 = ~pi644 & n19619;
  assign n19808 = ~pi715 & ~n19807;
  assign n19809 = ~n19806 & n19808;
  assign n19810 = pi1160 & ~n19809;
  assign n19811 = ~n19802 & n19810;
  assign n19812 = ~pi644 & ~n19794;
  assign n19813 = pi644 & n19799;
  assign n19814 = ~pi715 & ~n19813;
  assign n19815 = ~n19812 & n19814;
  assign n19816 = ~pi644 & n19805;
  assign n19817 = pi644 & n19619;
  assign n19818 = pi715 & ~n19817;
  assign n19819 = ~n19816 & n19818;
  assign n19820 = ~pi1160 & ~n19819;
  assign n19821 = ~n19815 & n19820;
  assign n19822 = ~n19811 & ~n19821;
  assign n19823 = pi790 & ~n19822;
  assign n19824 = ~pi790 & ~n19794;
  assign n19825 = pi832 & ~n19824;
  assign n19826 = ~n19823 & n19825;
  assign po300 = ~n19618 & ~n19826;
  assign n19828 = pi144 & ~n3268;
  assign n19829 = ~pi758 & ~n16814;
  assign n19830 = pi758 & n16905;
  assign n19831 = ~n19829 & ~n19830;
  assign n19832 = pi39 & ~n19831;
  assign n19833 = pi758 & n16839;
  assign n19834 = ~pi758 & n16655;
  assign n19835 = ~pi39 & ~n19834;
  assign n19836 = ~n19833 & n19835;
  assign n19837 = ~n19832 & ~n19836;
  assign n19838 = pi144 & ~n19837;
  assign n19839 = ~pi144 & pi758;
  assign n19840 = n16963 & n19839;
  assign n19841 = ~n19838 & ~n19840;
  assign n19842 = ~pi38 & ~n19841;
  assign n19843 = ~pi144 & ~n16968;
  assign n19844 = pi758 & n16842;
  assign n19845 = n16968 & ~n19844;
  assign n19846 = pi38 & ~n19843;
  assign n19847 = ~n19845 & n19846;
  assign n19848 = ~n19842 & ~n19847;
  assign n19849 = ~pi736 & n19848;
  assign n19850 = pi144 & ~n17074;
  assign n19851 = ~pi144 & ~n17166;
  assign n19852 = ~pi758 & ~n19851;
  assign n19853 = ~n19850 & n19852;
  assign n19854 = ~pi144 & ~n17233;
  assign n19855 = pi144 & n17295;
  assign n19856 = pi758 & ~n19855;
  assign n19857 = ~n19854 & n19856;
  assign n19858 = pi39 & ~n19857;
  assign n19859 = ~n19853 & n19858;
  assign n19860 = ~pi144 & ~n17340;
  assign n19861 = pi144 & ~n17317;
  assign n19862 = ~pi758 & ~n19860;
  assign n19863 = ~n19861 & n19862;
  assign n19864 = pi144 & n17344;
  assign n19865 = ~pi144 & n17351;
  assign n19866 = pi758 & ~n19865;
  assign n19867 = ~n19864 & n19866;
  assign n19868 = ~pi39 & ~n19867;
  assign n19869 = ~n19863 & n19868;
  assign n19870 = ~pi38 & ~n19869;
  assign n19871 = ~n19859 & n19870;
  assign n19872 = pi736 & ~n19316;
  assign n19873 = ~n19847 & n19872;
  assign n19874 = ~n19871 & n19873;
  assign n19875 = n3268 & ~n19874;
  assign n19876 = ~n19849 & n19875;
  assign n19877 = ~n19828 & ~n19876;
  assign n19878 = ~pi625 & n19877;
  assign n19879 = n3268 & ~n19848;
  assign n19880 = ~n19828 & ~n19879;
  assign n19881 = pi625 & n19880;
  assign n19882 = ~pi1153 & ~n19881;
  assign n19883 = ~n19878 & n19882;
  assign n19884 = pi144 & ~n17494;
  assign n19885 = pi736 & n3268;
  assign n19886 = ~n19884 & ~n19885;
  assign n19887 = pi144 & ~n18060;
  assign n19888 = ~pi144 & n18064;
  assign n19889 = ~pi38 & ~n19888;
  assign n19890 = ~n19887 & n19889;
  assign n19891 = n16968 & ~n17152;
  assign n19892 = pi38 & ~n19891;
  assign n19893 = ~n19843 & n19892;
  assign n19894 = n19885 & ~n19893;
  assign n19895 = ~n19890 & n19894;
  assign n19896 = ~n19886 & ~n19895;
  assign n19897 = pi625 & ~n19896;
  assign n19898 = ~pi625 & ~n19884;
  assign n19899 = pi1153 & ~n19898;
  assign n19900 = ~n19897 & n19899;
  assign n19901 = ~pi608 & ~n19900;
  assign n19902 = ~n19883 & n19901;
  assign n19903 = pi625 & n19877;
  assign n19904 = ~pi625 & n19880;
  assign n19905 = pi1153 & ~n19904;
  assign n19906 = ~n19903 & n19905;
  assign n19907 = ~pi625 & ~n19896;
  assign n19908 = pi625 & ~n19884;
  assign n19909 = ~pi1153 & ~n19908;
  assign n19910 = ~n19907 & n19909;
  assign n19911 = pi608 & ~n19910;
  assign n19912 = ~n19906 & n19911;
  assign n19913 = ~n19902 & ~n19912;
  assign n19914 = pi778 & ~n19913;
  assign n19915 = ~pi778 & n19877;
  assign n19916 = ~n19914 & ~n19915;
  assign n19917 = ~pi609 & ~n19916;
  assign n19918 = ~pi778 & n19896;
  assign n19919 = ~n19900 & ~n19910;
  assign n19920 = pi778 & ~n19919;
  assign n19921 = ~n19918 & ~n19920;
  assign n19922 = pi609 & n19921;
  assign n19923 = ~pi1155 & ~n19922;
  assign n19924 = ~n19917 & n19923;
  assign n19925 = n17526 & ~n19884;
  assign n19926 = ~n17526 & n19880;
  assign n19927 = ~n19925 & ~n19926;
  assign n19928 = pi609 & ~n19927;
  assign n19929 = ~pi609 & ~n19884;
  assign n19930 = pi1155 & ~n19929;
  assign n19931 = ~n19928 & n19930;
  assign n19932 = ~pi660 & ~n19931;
  assign n19933 = ~n19924 & n19932;
  assign n19934 = pi609 & ~n19916;
  assign n19935 = ~pi609 & n19921;
  assign n19936 = pi1155 & ~n19935;
  assign n19937 = ~n19934 & n19936;
  assign n19938 = ~pi609 & ~n19927;
  assign n19939 = pi609 & ~n19884;
  assign n19940 = ~pi1155 & ~n19939;
  assign n19941 = ~n19938 & n19940;
  assign n19942 = pi660 & ~n19941;
  assign n19943 = ~n19937 & n19942;
  assign n19944 = ~n19933 & ~n19943;
  assign n19945 = pi785 & ~n19944;
  assign n19946 = ~pi785 & ~n19916;
  assign n19947 = ~n19945 & ~n19946;
  assign n19948 = ~pi618 & ~n19947;
  assign n19949 = n17554 & ~n19884;
  assign n19950 = ~n17554 & n19921;
  assign n19951 = ~n19949 & ~n19950;
  assign n19952 = pi618 & ~n19951;
  assign n19953 = ~pi1154 & ~n19952;
  assign n19954 = ~n19948 & n19953;
  assign n19955 = ~pi785 & n19927;
  assign n19956 = ~n19931 & ~n19941;
  assign n19957 = pi785 & ~n19956;
  assign n19958 = ~n19955 & ~n19957;
  assign n19959 = pi618 & n19958;
  assign n19960 = ~pi618 & ~n19884;
  assign n19961 = pi1154 & ~n19960;
  assign n19962 = ~n19959 & n19961;
  assign n19963 = ~pi627 & ~n19962;
  assign n19964 = ~n19954 & n19963;
  assign n19965 = pi618 & ~n19947;
  assign n19966 = ~pi618 & ~n19951;
  assign n19967 = pi1154 & ~n19966;
  assign n19968 = ~n19965 & n19967;
  assign n19969 = ~pi618 & n19958;
  assign n19970 = pi618 & ~n19884;
  assign n19971 = ~pi1154 & ~n19970;
  assign n19972 = ~n19969 & n19971;
  assign n19973 = pi627 & ~n19972;
  assign n19974 = ~n19968 & n19973;
  assign n19975 = ~n19964 & ~n19974;
  assign n19976 = pi781 & ~n19975;
  assign n19977 = ~pi781 & ~n19947;
  assign n19978 = ~n19976 & ~n19977;
  assign n19979 = ~pi619 & ~n19978;
  assign n19980 = ~n17591 & n19951;
  assign n19981 = n17591 & n19884;
  assign n19982 = ~n19980 & ~n19981;
  assign n19983 = pi619 & n19982;
  assign n19984 = ~pi1159 & ~n19983;
  assign n19985 = ~n19979 & n19984;
  assign n19986 = ~pi781 & ~n19958;
  assign n19987 = ~n19962 & ~n19972;
  assign n19988 = pi781 & ~n19987;
  assign n19989 = ~n19986 & ~n19988;
  assign n19990 = pi619 & n19989;
  assign n19991 = ~pi619 & ~n19884;
  assign n19992 = pi1159 & ~n19991;
  assign n19993 = ~n19990 & n19992;
  assign n19994 = ~pi648 & ~n19993;
  assign n19995 = ~n19985 & n19994;
  assign n19996 = pi619 & ~n19978;
  assign n19997 = ~pi619 & n19982;
  assign n19998 = pi1159 & ~n19997;
  assign n19999 = ~n19996 & n19998;
  assign n20000 = ~pi619 & n19989;
  assign n20001 = pi619 & ~n19884;
  assign n20002 = ~pi1159 & ~n20001;
  assign n20003 = ~n20000 & n20002;
  assign n20004 = pi648 & ~n20003;
  assign n20005 = ~n19999 & n20004;
  assign n20006 = ~n19995 & ~n20005;
  assign n20007 = pi789 & ~n20006;
  assign n20008 = ~pi789 & ~n19978;
  assign n20009 = ~n20007 & ~n20008;
  assign n20010 = ~pi788 & n20009;
  assign n20011 = ~pi626 & n20009;
  assign n20012 = n17627 & ~n19884;
  assign n20013 = ~n17627 & n19982;
  assign n20014 = ~n20012 & ~n20013;
  assign n20015 = pi626 & n20014;
  assign n20016 = ~pi641 & ~n20015;
  assign n20017 = ~n20011 & n20016;
  assign n20018 = ~pi789 & ~n19989;
  assign n20019 = ~n19993 & ~n20003;
  assign n20020 = pi789 & ~n20019;
  assign n20021 = ~n20018 & ~n20020;
  assign n20022 = ~pi626 & n20021;
  assign n20023 = pi626 & ~n19884;
  assign n20024 = ~pi1158 & ~n20023;
  assign n20025 = ~n20022 & n20024;
  assign n20026 = ~n17634 & ~n20025;
  assign n20027 = ~n20017 & ~n20026;
  assign n20028 = pi626 & n20009;
  assign n20029 = ~pi626 & n20014;
  assign n20030 = pi641 & ~n20029;
  assign n20031 = ~n20028 & n20030;
  assign n20032 = pi626 & n20021;
  assign n20033 = ~pi626 & ~n19884;
  assign n20034 = pi1158 & ~n20033;
  assign n20035 = ~n20032 & n20034;
  assign n20036 = ~n17649 & ~n20035;
  assign n20037 = ~n20031 & ~n20036;
  assign n20038 = ~n20027 & ~n20037;
  assign n20039 = pi788 & ~n20038;
  assign n20040 = ~n20010 & ~n20039;
  assign n20041 = ~pi628 & n20040;
  assign n20042 = ~n20025 & ~n20035;
  assign n20043 = pi788 & ~n20042;
  assign n20044 = ~pi788 & ~n20021;
  assign n20045 = ~n20043 & ~n20044;
  assign n20046 = pi628 & n20045;
  assign n20047 = ~pi1156 & ~n20046;
  assign n20048 = ~n20041 & n20047;
  assign n20049 = ~n17670 & n20014;
  assign n20050 = n17670 & n19884;
  assign n20051 = ~n20049 & ~n20050;
  assign n20052 = pi628 & n20051;
  assign n20053 = ~pi628 & ~n19884;
  assign n20054 = pi1156 & ~n20053;
  assign n20055 = ~n20052 & n20054;
  assign n20056 = ~pi629 & ~n20055;
  assign n20057 = ~n20048 & n20056;
  assign n20058 = pi628 & n20040;
  assign n20059 = ~pi628 & n20045;
  assign n20060 = pi1156 & ~n20059;
  assign n20061 = ~n20058 & n20060;
  assign n20062 = ~pi628 & n20051;
  assign n20063 = pi628 & ~n19884;
  assign n20064 = ~pi1156 & ~n20063;
  assign n20065 = ~n20062 & n20064;
  assign n20066 = pi629 & ~n20065;
  assign n20067 = ~n20061 & n20066;
  assign n20068 = ~n20057 & ~n20067;
  assign n20069 = pi792 & ~n20068;
  assign n20070 = ~pi792 & n20040;
  assign n20071 = ~n20069 & ~n20070;
  assign n20072 = ~pi647 & ~n20071;
  assign n20073 = ~n17698 & ~n20045;
  assign n20074 = n17698 & n19884;
  assign n20075 = ~n20073 & ~n20074;
  assign n20076 = pi647 & n20075;
  assign n20077 = ~pi1157 & ~n20076;
  assign n20078 = ~n20072 & n20077;
  assign n20079 = ~pi792 & ~n20051;
  assign n20080 = ~n20055 & ~n20065;
  assign n20081 = pi792 & ~n20080;
  assign n20082 = ~n20079 & ~n20081;
  assign n20083 = pi647 & n20082;
  assign n20084 = ~pi647 & ~n19884;
  assign n20085 = pi1157 & ~n20084;
  assign n20086 = ~n20083 & n20085;
  assign n20087 = ~pi630 & ~n20086;
  assign n20088 = ~n20078 & n20087;
  assign n20089 = pi647 & ~n20071;
  assign n20090 = ~pi647 & n20075;
  assign n20091 = pi1157 & ~n20090;
  assign n20092 = ~n20089 & n20091;
  assign n20093 = ~pi647 & n20082;
  assign n20094 = pi647 & ~n19884;
  assign n20095 = ~pi1157 & ~n20094;
  assign n20096 = ~n20093 & n20095;
  assign n20097 = pi630 & ~n20096;
  assign n20098 = ~n20092 & n20097;
  assign n20099 = ~n20088 & ~n20098;
  assign n20100 = pi787 & ~n20099;
  assign n20101 = ~pi787 & ~n20071;
  assign n20102 = ~n20100 & ~n20101;
  assign n20103 = pi644 & ~n20102;
  assign n20104 = ~pi787 & ~n20082;
  assign n20105 = ~n20086 & ~n20096;
  assign n20106 = pi787 & ~n20105;
  assign n20107 = ~n20104 & ~n20106;
  assign n20108 = ~pi644 & n20107;
  assign n20109 = pi715 & ~n20108;
  assign n20110 = ~n20103 & n20109;
  assign n20111 = n17740 & ~n19884;
  assign n20112 = ~n17740 & n20075;
  assign n20113 = ~n20111 & ~n20112;
  assign n20114 = pi644 & ~n20113;
  assign n20115 = ~pi644 & ~n19884;
  assign n20116 = ~pi715 & ~n20115;
  assign n20117 = ~n20114 & n20116;
  assign n20118 = pi1160 & ~n20117;
  assign n20119 = ~n20110 & n20118;
  assign n20120 = ~pi644 & ~n20102;
  assign n20121 = pi644 & n20107;
  assign n20122 = ~pi715 & ~n20121;
  assign n20123 = ~n20120 & n20122;
  assign n20124 = ~pi644 & ~n20113;
  assign n20125 = pi644 & ~n19884;
  assign n20126 = pi715 & ~n20125;
  assign n20127 = ~n20124 & n20126;
  assign n20128 = ~pi1160 & ~n20127;
  assign n20129 = ~n20123 & n20128;
  assign n20130 = pi790 & ~n20119;
  assign n20131 = ~n20129 & n20130;
  assign n20132 = ~pi790 & n20102;
  assign n20133 = n6294 & ~n20132;
  assign n20134 = ~n20131 & n20133;
  assign n20135 = ~pi144 & ~n6294;
  assign n20136 = ~pi57 & ~n20135;
  assign n20137 = ~n20134 & n20136;
  assign n20138 = pi57 & pi144;
  assign n20139 = ~pi832 & ~n20138;
  assign n20140 = ~n20137 & n20139;
  assign n20141 = pi144 & ~n2755;
  assign n20142 = pi736 & n17153;
  assign n20143 = ~n20141 & ~n20142;
  assign n20144 = ~pi778 & n20143;
  assign n20145 = pi625 & n20142;
  assign n20146 = ~n20143 & ~n20145;
  assign n20147 = ~pi1153 & ~n20146;
  assign n20148 = pi1153 & ~n20141;
  assign n20149 = ~n20145 & n20148;
  assign n20150 = ~n20147 & ~n20149;
  assign n20151 = pi778 & ~n20150;
  assign n20152 = ~n20144 & ~n20151;
  assign n20153 = n19217 & n20152;
  assign n20154 = ~pi628 & n20153;
  assign n20155 = pi629 & ~n20154;
  assign n20156 = ~pi609 & ~pi1155;
  assign n20157 = pi609 & pi1155;
  assign n20158 = pi785 & ~n20156;
  assign n20159 = ~n20157 & n20158;
  assign n20160 = pi758 & n16933;
  assign n20161 = ~n20159 & n20160;
  assign n20162 = ~pi619 & pi1159;
  assign n20163 = pi619 & ~pi1159;
  assign n20164 = ~n20162 & ~n20163;
  assign n20165 = pi789 & ~n20164;
  assign n20166 = ~pi618 & ~pi1154;
  assign n20167 = pi618 & pi1154;
  assign n20168 = pi781 & ~n20166;
  assign n20169 = ~n20167 & n20168;
  assign n20170 = ~n17526 & ~n20169;
  assign n20171 = ~n20165 & n20170;
  assign n20172 = n20161 & n20171;
  assign n20173 = ~n17904 & n20172;
  assign n20174 = pi628 & ~n20173;
  assign n20175 = ~n20155 & ~n20174;
  assign n20176 = ~pi1156 & ~n20175;
  assign n20177 = pi628 & n20153;
  assign n20178 = ~pi628 & ~n20173;
  assign n20179 = pi629 & ~n20178;
  assign n20180 = pi1156 & ~n20179;
  assign n20181 = ~n20177 & n20180;
  assign n20182 = ~n20176 & ~n20181;
  assign n20183 = ~n20141 & ~n20182;
  assign n20184 = pi792 & n20183;
  assign n20185 = n17627 & ~n20141;
  assign n20186 = ~n17554 & n20152;
  assign n20187 = ~n17591 & n20186;
  assign n20188 = ~n20141 & ~n20187;
  assign n20189 = ~n20185 & ~n20188;
  assign n20190 = n17786 & n20189;
  assign n20191 = ~pi626 & n20172;
  assign n20192 = ~n20141 & ~n20191;
  assign n20193 = ~pi1158 & ~n20192;
  assign n20194 = pi641 & ~n20193;
  assign n20195 = ~n20190 & n20194;
  assign n20196 = n17787 & n20189;
  assign n20197 = pi626 & n20172;
  assign n20198 = ~n20141 & ~n20197;
  assign n20199 = pi1158 & ~n20198;
  assign n20200 = ~pi641 & ~n20199;
  assign n20201 = ~n20196 & n20200;
  assign n20202 = pi788 & ~n20195;
  assign n20203 = ~n20201 & n20202;
  assign n20204 = ~n20141 & ~n20160;
  assign n20205 = pi736 & n17154;
  assign n20206 = n20204 & ~n20205;
  assign n20207 = pi625 & n20205;
  assign n20208 = ~n20206 & ~n20207;
  assign n20209 = ~pi1153 & ~n20208;
  assign n20210 = ~pi608 & ~n20149;
  assign n20211 = ~n20209 & n20210;
  assign n20212 = pi1153 & n20204;
  assign n20213 = ~n20207 & n20212;
  assign n20214 = pi608 & ~n20147;
  assign n20215 = ~n20213 & n20214;
  assign n20216 = ~n20211 & ~n20215;
  assign n20217 = pi778 & ~n20216;
  assign n20218 = ~pi778 & ~n20206;
  assign n20219 = ~n20217 & ~n20218;
  assign n20220 = ~pi609 & ~n20219;
  assign n20221 = pi609 & n20152;
  assign n20222 = ~pi1155 & ~n20221;
  assign n20223 = ~n20220 & n20222;
  assign n20224 = n17527 & n20160;
  assign n20225 = pi1155 & ~n20141;
  assign n20226 = ~n20224 & n20225;
  assign n20227 = ~pi660 & ~n20226;
  assign n20228 = ~n20223 & n20227;
  assign n20229 = pi609 & ~n20219;
  assign n20230 = ~pi609 & n20152;
  assign n20231 = pi1155 & ~n20230;
  assign n20232 = ~n20229 & n20231;
  assign n20233 = n17539 & n20160;
  assign n20234 = ~pi1155 & ~n20141;
  assign n20235 = ~n20233 & n20234;
  assign n20236 = pi660 & ~n20235;
  assign n20237 = ~n20232 & n20236;
  assign n20238 = ~n20228 & ~n20237;
  assign n20239 = pi785 & ~n20238;
  assign n20240 = ~pi785 & ~n20219;
  assign n20241 = ~n20239 & ~n20240;
  assign n20242 = ~pi618 & ~n20241;
  assign n20243 = ~n20141 & ~n20186;
  assign n20244 = pi618 & ~n20243;
  assign n20245 = ~pi1154 & ~n20244;
  assign n20246 = ~n20242 & n20245;
  assign n20247 = pi618 & ~n17526;
  assign n20248 = n20161 & n20247;
  assign n20249 = pi1154 & ~n20141;
  assign n20250 = ~n20248 & n20249;
  assign n20251 = ~pi627 & ~n20250;
  assign n20252 = ~n20246 & n20251;
  assign n20253 = pi618 & ~n20241;
  assign n20254 = ~pi618 & ~n20243;
  assign n20255 = pi1154 & ~n20254;
  assign n20256 = ~n20253 & n20255;
  assign n20257 = ~pi618 & ~n17526;
  assign n20258 = n20161 & n20257;
  assign n20259 = ~pi1154 & ~n20141;
  assign n20260 = ~n20258 & n20259;
  assign n20261 = pi627 & ~n20260;
  assign n20262 = ~n20256 & n20261;
  assign n20263 = ~n20252 & ~n20262;
  assign n20264 = pi781 & ~n20263;
  assign n20265 = ~pi781 & ~n20241;
  assign n20266 = ~n20264 & ~n20265;
  assign n20267 = ~pi619 & ~n20266;
  assign n20268 = pi619 & ~n20188;
  assign n20269 = ~pi1159 & ~n20268;
  assign n20270 = ~n20267 & n20269;
  assign n20271 = n20161 & ~n20169;
  assign n20272 = pi619 & ~n17526;
  assign n20273 = n20271 & n20272;
  assign n20274 = pi1159 & ~n20141;
  assign n20275 = ~n20273 & n20274;
  assign n20276 = ~pi648 & ~n20275;
  assign n20277 = ~n20270 & n20276;
  assign n20278 = pi619 & ~n20266;
  assign n20279 = ~pi619 & ~n20188;
  assign n20280 = pi1159 & ~n20279;
  assign n20281 = ~n20278 & n20280;
  assign n20282 = ~pi619 & ~n17526;
  assign n20283 = n20271 & n20282;
  assign n20284 = ~pi1159 & ~n20141;
  assign n20285 = ~n20283 & n20284;
  assign n20286 = pi648 & ~n20285;
  assign n20287 = ~n20281 & n20286;
  assign n20288 = pi789 & ~n20277;
  assign n20289 = ~n20287 & n20288;
  assign n20290 = ~pi789 & n20266;
  assign n20291 = n17905 & ~n20290;
  assign n20292 = ~n20289 & n20291;
  assign n20293 = ~n20203 & ~n20292;
  assign n20294 = ~n20184 & ~n20293;
  assign n20295 = pi629 & n19244;
  assign n20296 = ~pi629 & n19245;
  assign n20297 = pi792 & ~n20295;
  assign n20298 = ~n20296 & n20297;
  assign n20299 = ~n20183 & n20298;
  assign n20300 = ~n17740 & ~n19271;
  assign n20301 = ~n20299 & n20300;
  assign n20302 = ~n20294 & n20301;
  assign n20303 = ~n17698 & n20173;
  assign n20304 = ~pi630 & n20303;
  assign n20305 = pi647 & ~n20304;
  assign n20306 = ~n19247 & n20153;
  assign n20307 = pi630 & ~n20306;
  assign n20308 = ~n20305 & ~n20307;
  assign n20309 = ~pi1157 & ~n20308;
  assign n20310 = ~pi630 & ~n20306;
  assign n20311 = pi647 & ~n20310;
  assign n20312 = pi630 & n20303;
  assign n20313 = pi1157 & ~n20312;
  assign n20314 = ~n20311 & n20313;
  assign n20315 = ~n20309 & ~n20314;
  assign n20316 = pi787 & ~n20141;
  assign n20317 = ~n20315 & n20316;
  assign n20318 = ~n20302 & ~n20317;
  assign n20319 = pi644 & n20318;
  assign n20320 = ~n19271 & n20306;
  assign n20321 = ~n20141 & ~n20320;
  assign n20322 = ~pi644 & ~n20321;
  assign n20323 = pi715 & ~n20322;
  assign n20324 = ~n20319 & n20323;
  assign n20325 = ~n17740 & n20303;
  assign n20326 = pi644 & n20325;
  assign n20327 = ~pi715 & ~n20141;
  assign n20328 = ~n20326 & n20327;
  assign n20329 = pi1160 & ~n20328;
  assign n20330 = ~n20324 & n20329;
  assign n20331 = ~pi644 & n20318;
  assign n20332 = pi644 & ~n20321;
  assign n20333 = ~pi715 & ~n20332;
  assign n20334 = ~n20331 & n20333;
  assign n20335 = ~pi644 & n20325;
  assign n20336 = pi715 & ~n20141;
  assign n20337 = ~n20335 & n20336;
  assign n20338 = ~pi1160 & ~n20337;
  assign n20339 = ~n20334 & n20338;
  assign n20340 = ~n20330 & ~n20339;
  assign n20341 = pi790 & ~n20340;
  assign n20342 = ~pi790 & n20318;
  assign n20343 = pi832 & ~n20342;
  assign n20344 = ~n20341 & n20343;
  assign po301 = ~n20140 & ~n20344;
  assign n20346 = ~pi145 & ~n17494;
  assign n20347 = n17627 & ~n20346;
  assign n20348 = ~pi698 & n3268;
  assign n20349 = n20346 & ~n20348;
  assign n20350 = pi145 & ~n18064;
  assign n20351 = ~pi38 & ~n20350;
  assign n20352 = n3268 & ~n20351;
  assign n20353 = ~pi145 & n18060;
  assign n20354 = ~n20352 & ~n20353;
  assign n20355 = ~pi145 & ~n16968;
  assign n20356 = n17480 & ~n20355;
  assign n20357 = ~pi698 & ~n20356;
  assign n20358 = ~n20354 & n20357;
  assign n20359 = ~n20349 & ~n20358;
  assign n20360 = ~pi778 & n20359;
  assign n20361 = pi625 & ~n20359;
  assign n20362 = ~pi625 & n20346;
  assign n20363 = pi1153 & ~n20362;
  assign n20364 = ~n20361 & n20363;
  assign n20365 = ~pi625 & ~n20359;
  assign n20366 = pi625 & n20346;
  assign n20367 = ~pi1153 & ~n20366;
  assign n20368 = ~n20365 & n20367;
  assign n20369 = ~n20364 & ~n20368;
  assign n20370 = pi778 & ~n20369;
  assign n20371 = ~n20360 & ~n20370;
  assign n20372 = ~n17554 & ~n20371;
  assign n20373 = n17554 & ~n20346;
  assign n20374 = ~n20372 & ~n20373;
  assign n20375 = ~n17591 & n20374;
  assign n20376 = n17591 & n20346;
  assign n20377 = ~n20375 & ~n20376;
  assign n20378 = ~n17627 & n20377;
  assign n20379 = ~n20347 & ~n20378;
  assign n20380 = ~n17670 & n20379;
  assign n20381 = n17670 & n20346;
  assign n20382 = ~n20380 & ~n20381;
  assign n20383 = ~pi792 & n20382;
  assign n20384 = pi628 & ~n20382;
  assign n20385 = ~pi628 & n20346;
  assign n20386 = pi1156 & ~n20385;
  assign n20387 = ~n20384 & n20386;
  assign n20388 = ~pi628 & ~n20382;
  assign n20389 = pi628 & n20346;
  assign n20390 = ~pi1156 & ~n20389;
  assign n20391 = ~n20388 & n20390;
  assign n20392 = ~n20387 & ~n20391;
  assign n20393 = pi792 & ~n20392;
  assign n20394 = ~n20383 & ~n20393;
  assign n20395 = ~pi647 & ~n20394;
  assign n20396 = pi647 & ~n20346;
  assign n20397 = ~n20395 & ~n20396;
  assign n20398 = ~pi1157 & n20397;
  assign n20399 = pi647 & ~n20394;
  assign n20400 = ~pi647 & ~n20346;
  assign n20401 = ~n20399 & ~n20400;
  assign n20402 = pi1157 & n20401;
  assign n20403 = ~n20398 & ~n20402;
  assign n20404 = pi787 & ~n20403;
  assign n20405 = ~pi787 & n20394;
  assign n20406 = ~n20404 & ~n20405;
  assign n20407 = ~pi644 & ~n20406;
  assign n20408 = pi715 & ~n20407;
  assign n20409 = pi145 & ~n3268;
  assign n20410 = ~pi145 & ~n16816;
  assign n20411 = pi767 & ~n20410;
  assign n20412 = pi145 & ~n16963;
  assign n20413 = ~pi145 & ~pi767;
  assign n20414 = n16907 & n20413;
  assign n20415 = ~n20412 & ~n20414;
  assign n20416 = ~n20411 & n20415;
  assign n20417 = ~pi38 & ~n20416;
  assign n20418 = ~pi767 & n16970;
  assign n20419 = pi38 & ~n20355;
  assign n20420 = ~n20418 & n20419;
  assign n20421 = ~n20417 & ~n20420;
  assign n20422 = n3268 & ~n20421;
  assign n20423 = ~n20409 & ~n20422;
  assign n20424 = ~n17526 & ~n20423;
  assign n20425 = n17526 & ~n20346;
  assign n20426 = ~n20424 & ~n20425;
  assign n20427 = ~pi785 & ~n20426;
  assign n20428 = ~n17527 & ~n20346;
  assign n20429 = pi609 & n20424;
  assign n20430 = ~n20428 & ~n20429;
  assign n20431 = pi1155 & ~n20430;
  assign n20432 = ~n17539 & ~n20346;
  assign n20433 = ~pi609 & n20424;
  assign n20434 = ~n20432 & ~n20433;
  assign n20435 = ~pi1155 & ~n20434;
  assign n20436 = ~n20431 & ~n20435;
  assign n20437 = pi785 & ~n20436;
  assign n20438 = ~n20427 & ~n20437;
  assign n20439 = ~pi781 & ~n20438;
  assign n20440 = pi618 & n20438;
  assign n20441 = ~pi618 & n20346;
  assign n20442 = pi1154 & ~n20441;
  assign n20443 = ~n20440 & n20442;
  assign n20444 = ~pi618 & n20438;
  assign n20445 = pi618 & n20346;
  assign n20446 = ~pi1154 & ~n20445;
  assign n20447 = ~n20444 & n20446;
  assign n20448 = ~n20443 & ~n20447;
  assign n20449 = pi781 & ~n20448;
  assign n20450 = ~n20439 & ~n20449;
  assign n20451 = ~pi789 & ~n20450;
  assign n20452 = pi619 & n20450;
  assign n20453 = ~pi619 & n20346;
  assign n20454 = pi1159 & ~n20453;
  assign n20455 = ~n20452 & n20454;
  assign n20456 = ~pi619 & n20450;
  assign n20457 = pi619 & n20346;
  assign n20458 = ~pi1159 & ~n20457;
  assign n20459 = ~n20456 & n20458;
  assign n20460 = ~n20455 & ~n20459;
  assign n20461 = pi789 & ~n20460;
  assign n20462 = ~n20451 & ~n20461;
  assign n20463 = ~pi788 & ~n20462;
  assign n20464 = pi626 & n20462;
  assign n20465 = ~pi626 & n20346;
  assign n20466 = pi1158 & ~n20465;
  assign n20467 = ~n20464 & n20466;
  assign n20468 = ~pi626 & n20462;
  assign n20469 = pi626 & n20346;
  assign n20470 = ~pi1158 & ~n20469;
  assign n20471 = ~n20468 & n20470;
  assign n20472 = ~n20467 & ~n20471;
  assign n20473 = pi788 & ~n20472;
  assign n20474 = ~n20463 & ~n20473;
  assign n20475 = ~n17698 & n20474;
  assign n20476 = n17698 & n20346;
  assign n20477 = ~n20475 & ~n20476;
  assign n20478 = ~n17740 & ~n20477;
  assign n20479 = n17740 & n20346;
  assign n20480 = ~n20478 & ~n20479;
  assign n20481 = pi644 & ~n20480;
  assign n20482 = ~pi644 & n20346;
  assign n20483 = ~pi715 & ~n20482;
  assign n20484 = ~n20481 & n20483;
  assign n20485 = pi1160 & ~n20484;
  assign n20486 = ~n20408 & n20485;
  assign n20487 = pi630 & ~pi647;
  assign n20488 = pi1157 & n20487;
  assign n20489 = ~pi630 & pi647;
  assign n20490 = ~pi1157 & n20489;
  assign n20491 = ~n20488 & ~n20490;
  assign n20492 = n20477 & ~n20491;
  assign n20493 = n17738 & ~n20397;
  assign n20494 = n17737 & ~n20401;
  assign n20495 = ~n20493 & ~n20494;
  assign n20496 = ~n20492 & n20495;
  assign n20497 = pi787 & ~n20496;
  assign n20498 = ~pi628 & pi629;
  assign n20499 = pi1156 & n20498;
  assign n20500 = pi628 & ~pi629;
  assign n20501 = ~pi1156 & n20500;
  assign n20502 = ~n20499 & ~n20501;
  assign n20503 = ~n20474 & ~n20502;
  assign n20504 = ~pi629 & n20387;
  assign n20505 = pi629 & n20391;
  assign n20506 = ~n20504 & ~n20505;
  assign n20507 = ~n20503 & n20506;
  assign n20508 = pi792 & ~n20507;
  assign n20509 = pi698 & n20421;
  assign n20510 = ~pi145 & n17074;
  assign n20511 = pi145 & n17166;
  assign n20512 = pi767 & ~n20511;
  assign n20513 = ~n20510 & n20512;
  assign n20514 = pi145 & n17233;
  assign n20515 = ~pi145 & ~n17295;
  assign n20516 = ~pi767 & ~n20515;
  assign n20517 = ~n20514 & n20516;
  assign n20518 = pi39 & ~n20517;
  assign n20519 = ~n20513 & n20518;
  assign n20520 = pi145 & ~n17340;
  assign n20521 = ~pi145 & ~n17317;
  assign n20522 = pi767 & ~n20520;
  assign n20523 = ~n20521 & n20522;
  assign n20524 = ~pi145 & n17344;
  assign n20525 = pi145 & n17351;
  assign n20526 = ~pi767 & ~n20525;
  assign n20527 = ~n20524 & n20526;
  assign n20528 = ~n20523 & ~n20527;
  assign n20529 = ~pi39 & ~n20528;
  assign n20530 = ~pi38 & ~n20529;
  assign n20531 = ~n20519 & n20530;
  assign n20532 = ~pi767 & ~n17259;
  assign n20533 = n19303 & ~n20532;
  assign n20534 = ~pi145 & ~n20533;
  assign n20535 = ~pi767 & n16933;
  assign n20536 = ~n17154 & ~n20535;
  assign n20537 = pi145 & ~n20536;
  assign n20538 = n6250 & n20537;
  assign n20539 = pi38 & ~n20538;
  assign n20540 = ~n20534 & n20539;
  assign n20541 = ~pi698 & ~n20540;
  assign n20542 = ~n20531 & n20541;
  assign n20543 = n3268 & ~n20542;
  assign n20544 = ~n20509 & n20543;
  assign n20545 = ~n20409 & ~n20544;
  assign n20546 = ~pi625 & n20545;
  assign n20547 = pi625 & n20423;
  assign n20548 = ~pi1153 & ~n20547;
  assign n20549 = ~n20546 & n20548;
  assign n20550 = ~pi608 & ~n20364;
  assign n20551 = ~n20549 & n20550;
  assign n20552 = pi625 & n20545;
  assign n20553 = ~pi625 & n20423;
  assign n20554 = pi1153 & ~n20553;
  assign n20555 = ~n20552 & n20554;
  assign n20556 = pi608 & ~n20368;
  assign n20557 = ~n20555 & n20556;
  assign n20558 = ~n20551 & ~n20557;
  assign n20559 = pi778 & ~n20558;
  assign n20560 = ~pi778 & n20545;
  assign n20561 = ~n20559 & ~n20560;
  assign n20562 = ~pi609 & ~n20561;
  assign n20563 = pi609 & n20371;
  assign n20564 = ~pi1155 & ~n20563;
  assign n20565 = ~n20562 & n20564;
  assign n20566 = ~pi660 & ~n20431;
  assign n20567 = ~n20565 & n20566;
  assign n20568 = pi609 & ~n20561;
  assign n20569 = ~pi609 & n20371;
  assign n20570 = pi1155 & ~n20569;
  assign n20571 = ~n20568 & n20570;
  assign n20572 = pi660 & ~n20435;
  assign n20573 = ~n20571 & n20572;
  assign n20574 = ~n20567 & ~n20573;
  assign n20575 = pi785 & ~n20574;
  assign n20576 = ~pi785 & ~n20561;
  assign n20577 = ~n20575 & ~n20576;
  assign n20578 = ~pi618 & ~n20577;
  assign n20579 = pi618 & n20374;
  assign n20580 = ~pi1154 & ~n20579;
  assign n20581 = ~n20578 & n20580;
  assign n20582 = ~pi627 & ~n20443;
  assign n20583 = ~n20581 & n20582;
  assign n20584 = pi618 & ~n20577;
  assign n20585 = ~pi618 & n20374;
  assign n20586 = pi1154 & ~n20585;
  assign n20587 = ~n20584 & n20586;
  assign n20588 = pi627 & ~n20447;
  assign n20589 = ~n20587 & n20588;
  assign n20590 = ~n20583 & ~n20589;
  assign n20591 = pi781 & ~n20590;
  assign n20592 = ~pi781 & ~n20577;
  assign n20593 = ~n20591 & ~n20592;
  assign n20594 = ~pi619 & ~n20593;
  assign n20595 = pi619 & ~n20377;
  assign n20596 = ~pi1159 & ~n20595;
  assign n20597 = ~n20594 & n20596;
  assign n20598 = ~pi648 & ~n20455;
  assign n20599 = ~n20597 & n20598;
  assign n20600 = pi619 & ~n20593;
  assign n20601 = ~pi619 & ~n20377;
  assign n20602 = pi1159 & ~n20601;
  assign n20603 = ~n20600 & n20602;
  assign n20604 = pi648 & ~n20459;
  assign n20605 = ~n20603 & n20604;
  assign n20606 = pi789 & ~n20599;
  assign n20607 = ~n20605 & n20606;
  assign n20608 = ~pi789 & n20593;
  assign n20609 = n17905 & ~n20608;
  assign n20610 = ~n20607 & n20609;
  assign n20611 = n17792 & n20379;
  assign n20612 = ~n17669 & n20472;
  assign n20613 = ~n20611 & ~n20612;
  assign n20614 = pi788 & ~n20613;
  assign n20615 = ~n20298 & ~n20614;
  assign n20616 = ~n20610 & n20615;
  assign n20617 = ~n20508 & ~n20616;
  assign n20618 = n20300 & ~n20617;
  assign n20619 = ~n20497 & ~n20618;
  assign n20620 = ~pi644 & n20619;
  assign n20621 = pi644 & ~n20406;
  assign n20622 = ~pi715 & ~n20621;
  assign n20623 = ~n20620 & n20622;
  assign n20624 = ~pi644 & ~n20480;
  assign n20625 = pi644 & n20346;
  assign n20626 = pi715 & ~n20625;
  assign n20627 = ~n20624 & n20626;
  assign n20628 = ~pi1160 & ~n20627;
  assign n20629 = ~n20623 & n20628;
  assign n20630 = ~n20486 & ~n20629;
  assign n20631 = pi790 & ~n20630;
  assign n20632 = pi644 & n20485;
  assign n20633 = pi790 & ~n20632;
  assign n20634 = n20619 & ~n20633;
  assign n20635 = ~n20631 & ~n20634;
  assign n20636 = ~po1038 & ~n20635;
  assign n20637 = ~pi145 & po1038;
  assign n20638 = ~pi832 & ~n20637;
  assign n20639 = ~n20636 & n20638;
  assign n20640 = ~pi145 & ~n2755;
  assign n20641 = ~n20535 & ~n20640;
  assign n20642 = ~n17794 & ~n20641;
  assign n20643 = ~pi785 & ~n20642;
  assign n20644 = ~n17799 & ~n20641;
  assign n20645 = pi1155 & ~n20644;
  assign n20646 = ~n17802 & n20642;
  assign n20647 = ~pi1155 & ~n20646;
  assign n20648 = ~n20645 & ~n20647;
  assign n20649 = pi785 & ~n20648;
  assign n20650 = ~n20643 & ~n20649;
  assign n20651 = ~pi781 & ~n20650;
  assign n20652 = ~n17809 & n20650;
  assign n20653 = pi1154 & ~n20652;
  assign n20654 = ~n17812 & n20650;
  assign n20655 = ~pi1154 & ~n20654;
  assign n20656 = ~n20653 & ~n20655;
  assign n20657 = pi781 & ~n20656;
  assign n20658 = ~n20651 & ~n20657;
  assign n20659 = ~pi789 & ~n20658;
  assign n20660 = pi619 & n20658;
  assign n20661 = ~pi619 & n20640;
  assign n20662 = pi1159 & ~n20661;
  assign n20663 = ~n20660 & n20662;
  assign n20664 = ~pi619 & n20658;
  assign n20665 = pi619 & n20640;
  assign n20666 = ~pi1159 & ~n20665;
  assign n20667 = ~n20664 & n20666;
  assign n20668 = ~n20663 & ~n20667;
  assign n20669 = pi789 & ~n20668;
  assign n20670 = ~n20659 & ~n20669;
  assign n20671 = ~pi788 & ~n20670;
  assign n20672 = pi626 & n20670;
  assign n20673 = ~pi626 & n20640;
  assign n20674 = pi1158 & ~n20673;
  assign n20675 = ~n20672 & n20674;
  assign n20676 = ~pi626 & n20670;
  assign n20677 = pi626 & n20640;
  assign n20678 = ~pi1158 & ~n20677;
  assign n20679 = ~n20676 & n20678;
  assign n20680 = ~n20675 & ~n20679;
  assign n20681 = pi788 & ~n20680;
  assign n20682 = ~n20671 & ~n20681;
  assign n20683 = ~n17698 & n20682;
  assign n20684 = n17698 & n20640;
  assign n20685 = ~n20683 & ~n20684;
  assign n20686 = ~n20491 & n20685;
  assign n20687 = ~pi698 & n17153;
  assign n20688 = ~n20640 & ~n20687;
  assign n20689 = ~pi778 & n20688;
  assign n20690 = ~pi625 & n20687;
  assign n20691 = ~n20688 & ~n20690;
  assign n20692 = pi1153 & ~n20691;
  assign n20693 = ~pi1153 & ~n20640;
  assign n20694 = ~n20690 & n20693;
  assign n20695 = ~n20692 & ~n20694;
  assign n20696 = pi778 & ~n20695;
  assign n20697 = ~n20689 & ~n20696;
  assign n20698 = ~n17780 & n20697;
  assign n20699 = ~n17782 & n20698;
  assign n20700 = ~n17784 & n20699;
  assign n20701 = ~n17916 & n20700;
  assign n20702 = ~n17947 & n20701;
  assign n20703 = ~pi647 & n20702;
  assign n20704 = pi647 & n20640;
  assign n20705 = ~pi1157 & ~n20704;
  assign n20706 = ~n20703 & n20705;
  assign n20707 = pi647 & ~n20702;
  assign n20708 = ~pi647 & ~n20640;
  assign n20709 = ~n20707 & ~n20708;
  assign n20710 = pi1157 & ~n20709;
  assign n20711 = ~n20706 & ~n20710;
  assign n20712 = ~n17739 & ~n20711;
  assign n20713 = ~n20686 & ~n20712;
  assign n20714 = pi787 & ~n20713;
  assign n20715 = n17792 & n20700;
  assign n20716 = ~n17669 & n20680;
  assign n20717 = ~n20715 & ~n20716;
  assign n20718 = pi788 & ~n20717;
  assign n20719 = ~n16842 & ~n20688;
  assign n20720 = pi625 & n20719;
  assign n20721 = n20641 & ~n20719;
  assign n20722 = ~n20720 & ~n20721;
  assign n20723 = n20693 & ~n20722;
  assign n20724 = ~pi608 & ~n20692;
  assign n20725 = ~n20723 & n20724;
  assign n20726 = pi1153 & n20641;
  assign n20727 = ~n20720 & n20726;
  assign n20728 = pi608 & ~n20694;
  assign n20729 = ~n20727 & n20728;
  assign n20730 = ~n20725 & ~n20729;
  assign n20731 = pi778 & ~n20730;
  assign n20732 = ~pi778 & ~n20721;
  assign n20733 = ~n20731 & ~n20732;
  assign n20734 = ~pi609 & ~n20733;
  assign n20735 = pi609 & n20697;
  assign n20736 = ~pi1155 & ~n20735;
  assign n20737 = ~n20734 & n20736;
  assign n20738 = ~pi660 & ~n20645;
  assign n20739 = ~n20737 & n20738;
  assign n20740 = pi609 & ~n20733;
  assign n20741 = ~pi609 & n20697;
  assign n20742 = pi1155 & ~n20741;
  assign n20743 = ~n20740 & n20742;
  assign n20744 = pi660 & ~n20647;
  assign n20745 = ~n20743 & n20744;
  assign n20746 = ~n20739 & ~n20745;
  assign n20747 = pi785 & ~n20746;
  assign n20748 = ~pi785 & ~n20733;
  assign n20749 = ~n20747 & ~n20748;
  assign n20750 = ~pi618 & ~n20749;
  assign n20751 = pi618 & n20698;
  assign n20752 = ~pi1154 & ~n20751;
  assign n20753 = ~n20750 & n20752;
  assign n20754 = ~pi627 & ~n20653;
  assign n20755 = ~n20753 & n20754;
  assign n20756 = pi618 & ~n20749;
  assign n20757 = ~pi618 & n20698;
  assign n20758 = pi1154 & ~n20757;
  assign n20759 = ~n20756 & n20758;
  assign n20760 = pi627 & ~n20655;
  assign n20761 = ~n20759 & n20760;
  assign n20762 = ~n20755 & ~n20761;
  assign n20763 = pi781 & ~n20762;
  assign n20764 = ~pi781 & ~n20749;
  assign n20765 = ~n20763 & ~n20764;
  assign n20766 = ~pi619 & ~n20765;
  assign n20767 = pi619 & n20699;
  assign n20768 = ~pi1159 & ~n20767;
  assign n20769 = ~n20766 & n20768;
  assign n20770 = ~pi648 & ~n20663;
  assign n20771 = ~n20769 & n20770;
  assign n20772 = pi619 & ~n20765;
  assign n20773 = ~pi619 & n20699;
  assign n20774 = pi1159 & ~n20773;
  assign n20775 = ~n20772 & n20774;
  assign n20776 = pi648 & ~n20667;
  assign n20777 = ~n20775 & n20776;
  assign n20778 = pi789 & ~n20771;
  assign n20779 = ~n20777 & n20778;
  assign n20780 = ~pi789 & n20765;
  assign n20781 = n17905 & ~n20780;
  assign n20782 = ~n20779 & n20781;
  assign n20783 = ~n20718 & ~n20782;
  assign n20784 = ~n20298 & ~n20783;
  assign n20785 = n17944 & n20682;
  assign n20786 = pi1156 & ~n17918;
  assign n20787 = n20701 & n20786;
  assign n20788 = ~n20785 & ~n20787;
  assign n20789 = ~pi629 & ~n20788;
  assign n20790 = ~pi1156 & ~n17927;
  assign n20791 = n20701 & n20790;
  assign n20792 = n17943 & n20682;
  assign n20793 = ~n20791 & ~n20792;
  assign n20794 = pi629 & ~n20793;
  assign n20795 = ~n20789 & ~n20794;
  assign n20796 = pi792 & ~n20795;
  assign n20797 = n20300 & ~n20796;
  assign n20798 = ~n20784 & n20797;
  assign n20799 = ~n20714 & ~n20798;
  assign n20800 = pi644 & n20799;
  assign n20801 = ~pi787 & ~n20702;
  assign n20802 = pi787 & ~n20711;
  assign n20803 = ~n20801 & ~n20802;
  assign n20804 = ~pi644 & n20803;
  assign n20805 = pi715 & ~n20804;
  assign n20806 = ~n20800 & n20805;
  assign n20807 = ~n17740 & ~n20685;
  assign n20808 = n17740 & n20640;
  assign n20809 = ~n20807 & ~n20808;
  assign n20810 = pi644 & ~n20809;
  assign n20811 = ~pi644 & n20640;
  assign n20812 = ~pi715 & ~n20811;
  assign n20813 = ~n20810 & n20812;
  assign n20814 = pi1160 & ~n20813;
  assign n20815 = ~n20806 & n20814;
  assign n20816 = ~pi644 & n20799;
  assign n20817 = pi644 & n20803;
  assign n20818 = ~pi715 & ~n20817;
  assign n20819 = ~n20816 & n20818;
  assign n20820 = ~pi644 & ~n20809;
  assign n20821 = pi644 & n20640;
  assign n20822 = pi715 & ~n20821;
  assign n20823 = ~n20820 & n20822;
  assign n20824 = ~pi1160 & ~n20823;
  assign n20825 = ~n20819 & n20824;
  assign n20826 = ~n20815 & ~n20825;
  assign n20827 = pi790 & ~n20826;
  assign n20828 = ~pi790 & n20799;
  assign n20829 = pi832 & ~n20828;
  assign n20830 = ~n20827 & n20829;
  assign po302 = ~n20639 & ~n20830;
  assign n20832 = ~pi907 & n6222;
  assign n20833 = pi146 & ~n16785;
  assign n20834 = ~n20832 & n20833;
  assign n20835 = pi146 & ~n16776;
  assign n20836 = n20832 & n20835;
  assign n20837 = pi735 & pi907;
  assign n20838 = n16785 & n20837;
  assign n20839 = ~pi947 & ~n20838;
  assign n20840 = ~n20836 & n20839;
  assign n20841 = pi743 & n16785;
  assign n20842 = pi947 & ~n20833;
  assign n20843 = ~n20841 & n20842;
  assign n20844 = ~n20840 & ~n20843;
  assign n20845 = ~n20834 & ~n20844;
  assign n20846 = ~n3461 & ~n20845;
  assign n20847 = pi743 & pi947;
  assign n20848 = pi907 & ~pi947;
  assign n20849 = pi735 & n20848;
  assign n20850 = ~n20847 & ~n20849;
  assign n20851 = n16661 & ~n20850;
  assign n20852 = pi146 & ~n16661;
  assign n20853 = ~n20851 & ~n20852;
  assign n20854 = n3461 & ~n20853;
  assign n20855 = ~pi215 & ~n20854;
  assign n20856 = ~n20846 & n20855;
  assign n20857 = pi146 & n16810;
  assign n20858 = n16704 & ~n20850;
  assign n20859 = pi215 & ~n20858;
  assign n20860 = ~n20857 & n20859;
  assign n20861 = ~n20856 & ~n20860;
  assign n20862 = pi299 & ~n20861;
  assign n20863 = n16785 & ~n20850;
  assign n20864 = ~n6197 & ~n20833;
  assign n20865 = ~n20863 & n20864;
  assign n20866 = n16776 & ~n20850;
  assign n20867 = n6197 & ~n20835;
  assign n20868 = ~n20866 & n20867;
  assign n20869 = ~n20865 & ~n20868;
  assign n20870 = ~n3053 & ~n20869;
  assign n20871 = n3053 & n20853;
  assign n20872 = ~pi223 & ~n20871;
  assign n20873 = ~n20870 & n20872;
  assign n20874 = pi146 & ~n16704;
  assign n20875 = ~n20858 & ~n20874;
  assign n20876 = ~n6197 & ~n20875;
  assign n20877 = ~pi146 & ~n16726;
  assign n20878 = n16726 & n20850;
  assign n20879 = n6197 & ~n20877;
  assign n20880 = ~n20878 & n20879;
  assign n20881 = ~n20876 & ~n20880;
  assign n20882 = pi223 & ~n20881;
  assign n20883 = ~pi299 & ~n20882;
  assign n20884 = ~n20873 & n20883;
  assign n20885 = ~n20862 & ~n20884;
  assign n20886 = pi39 & ~n20885;
  assign n20887 = ~pi146 & ~n16649;
  assign n20888 = n16649 & n20850;
  assign n20889 = pi299 & ~n20887;
  assign n20890 = ~n20888 & n20889;
  assign n20891 = ~pi146 & ~n16653;
  assign n20892 = n16653 & n20850;
  assign n20893 = ~pi299 & ~n20891;
  assign n20894 = ~n20892 & n20893;
  assign n20895 = ~pi39 & ~n20890;
  assign n20896 = ~n20894 & n20895;
  assign n20897 = ~pi38 & ~n20896;
  assign n20898 = ~n20886 & n20897;
  assign n20899 = ~pi146 & ~n16968;
  assign n20900 = n2755 & n20850;
  assign n20901 = n6250 & n20900;
  assign n20902 = pi38 & ~n20901;
  assign n20903 = ~n20899 & n20902;
  assign n20904 = n10178 & ~n20903;
  assign n20905 = ~n20898 & n20904;
  assign n20906 = ~pi146 & ~n10178;
  assign n20907 = ~pi832 & ~n20906;
  assign n20908 = ~n20905 & n20907;
  assign n20909 = ~pi146 & ~n2755;
  assign n20910 = pi832 & ~n20909;
  assign n20911 = ~n20900 & n20910;
  assign po303 = n20908 | n20911;
  assign n20913 = ~pi770 & pi947;
  assign n20914 = pi726 & n20848;
  assign n20915 = ~n20913 & ~n20914;
  assign n20916 = n2755 & ~n20915;
  assign n20917 = ~pi147 & ~n2755;
  assign n20918 = pi832 & ~n20917;
  assign n20919 = ~n20916 & n20918;
  assign n20920 = ~pi947 & n16655;
  assign n20921 = ~pi39 & ~n20920;
  assign n20922 = ~pi299 & n16792;
  assign n20923 = pi947 & n20922;
  assign n20924 = ~pi947 & n16799;
  assign n20925 = n16785 & n20848;
  assign n20926 = ~n16797 & ~n20925;
  assign n20927 = ~n3461 & ~n20926;
  assign n20928 = ~pi215 & ~n20927;
  assign n20929 = ~n20924 & n20928;
  assign n20930 = pi215 & ~n16809;
  assign n20931 = n16704 & n20848;
  assign n20932 = n20930 & ~n20931;
  assign n20933 = ~n20929 & ~n20932;
  assign n20934 = pi299 & ~n20933;
  assign n20935 = ~n16793 & ~n20934;
  assign n20936 = ~n20923 & n20935;
  assign n20937 = pi39 & ~n20936;
  assign n20938 = ~n20921 & ~n20937;
  assign n20939 = ~pi38 & n20938;
  assign n20940 = pi38 & ~pi947;
  assign n20941 = n17485 & n20940;
  assign n20942 = ~n20939 & ~n20941;
  assign n20943 = ~pi770 & n20942;
  assign n20944 = pi770 & ~n17487;
  assign n20945 = ~n20943 & ~n20944;
  assign n20946 = ~pi147 & ~n20945;
  assign n20947 = ~n17486 & ~n20941;
  assign n20948 = pi947 & n16655;
  assign n20949 = ~pi39 & ~n20948;
  assign n20950 = pi947 & n16792;
  assign n20951 = ~pi299 & ~n20950;
  assign n20952 = pi215 & pi947;
  assign n20953 = n16704 & n20952;
  assign n20954 = pi299 & ~n20953;
  assign n20955 = pi947 & n16785;
  assign n20956 = ~n3461 & ~n20955;
  assign n20957 = pi947 & n16661;
  assign n20958 = n3461 & ~n20957;
  assign n20959 = ~pi215 & ~n20958;
  assign n20960 = ~n20956 & n20959;
  assign n20961 = n20954 & ~n20960;
  assign n20962 = ~n20951 & ~n20961;
  assign n20963 = pi39 & ~n20962;
  assign n20964 = ~n20949 & ~n20963;
  assign n20965 = ~pi38 & ~n20964;
  assign n20966 = n20947 & ~n20965;
  assign n20967 = pi147 & ~pi770;
  assign n20968 = n20966 & n20967;
  assign n20969 = ~pi726 & ~n20968;
  assign n20970 = ~n20946 & n20969;
  assign n20971 = n16799 & ~n20848;
  assign n20972 = ~n16797 & ~n20955;
  assign n20973 = ~n3461 & ~n20972;
  assign n20974 = ~pi215 & ~n20973;
  assign n20975 = ~n20971 & n20974;
  assign n20976 = ~n20930 & ~n20975;
  assign n20977 = pi299 & ~n20976;
  assign n20978 = ~n16788 & ~n16789;
  assign n20979 = n6217 & ~n20978;
  assign n20980 = ~pi223 & ~n20979;
  assign n20981 = ~pi947 & n16728;
  assign n20982 = pi223 & ~n20981;
  assign n20983 = n16728 & ~n20848;
  assign n20984 = pi223 & ~n20983;
  assign n20985 = ~n20982 & ~n20984;
  assign n20986 = ~n20980 & n20985;
  assign n20987 = ~pi299 & ~n20986;
  assign n20988 = pi299 & pi947;
  assign n20989 = ~n20977 & ~n20988;
  assign n20990 = ~n20987 & n20989;
  assign n20991 = pi39 & n20990;
  assign n20992 = ~n6217 & n16655;
  assign n20993 = ~pi39 & ~n20992;
  assign n20994 = n16655 & n20993;
  assign n20995 = ~n20991 & ~n20994;
  assign n20996 = ~pi147 & n20995;
  assign n20997 = ~n6217 & n16792;
  assign n20998 = ~pi299 & n20997;
  assign n20999 = pi215 & ~n16805;
  assign n21000 = ~n6217 & n16661;
  assign n21001 = n3461 & n21000;
  assign n21002 = ~pi215 & ~n21001;
  assign n21003 = ~n16802 & n21002;
  assign n21004 = pi299 & ~n21003;
  assign n21005 = ~n20999 & n21004;
  assign n21006 = ~n20998 & ~n21005;
  assign n21007 = pi39 & n21006;
  assign n21008 = ~n20993 & ~n21007;
  assign n21009 = pi147 & n21008;
  assign n21010 = ~pi38 & ~n21009;
  assign n21011 = ~n20996 & n21010;
  assign n21012 = n6217 & n17485;
  assign n21013 = ~pi147 & ~n21012;
  assign n21014 = ~n6217 & n16968;
  assign n21015 = pi38 & ~n21014;
  assign n21016 = ~n21013 & n21015;
  assign n21017 = ~pi770 & ~n21016;
  assign n21018 = ~n21011 & n21017;
  assign n21019 = ~n20953 & ~n20976;
  assign n21020 = pi299 & ~n21019;
  assign n21021 = ~n20848 & n20922;
  assign n21022 = ~n21020 & ~n21021;
  assign n21023 = pi39 & ~n21022;
  assign n21024 = n16655 & ~n20848;
  assign n21025 = ~pi39 & n21024;
  assign n21026 = ~n21023 & ~n21025;
  assign n21027 = ~pi147 & n21026;
  assign n21028 = pi215 & ~n20931;
  assign n21029 = ~n3461 & ~n20925;
  assign n21030 = pi907 & n16661;
  assign n21031 = ~pi947 & n21030;
  assign n21032 = n3461 & ~n21031;
  assign n21033 = ~n21029 & ~n21032;
  assign n21034 = ~pi215 & ~n21033;
  assign n21035 = ~n21028 & ~n21034;
  assign n21036 = pi299 & ~n21035;
  assign n21037 = n16792 & n20848;
  assign n21038 = ~pi299 & ~n21037;
  assign n21039 = ~n21036 & ~n21038;
  assign n21040 = pi39 & ~n21039;
  assign n21041 = n16655 & n20848;
  assign n21042 = ~pi39 & ~n21041;
  assign n21043 = ~n21040 & ~n21042;
  assign n21044 = pi147 & n21043;
  assign n21045 = ~pi38 & ~n21044;
  assign n21046 = ~n21027 & n21045;
  assign n21047 = ~pi147 & ~n16968;
  assign n21048 = n16968 & n20848;
  assign n21049 = pi38 & ~n21048;
  assign n21050 = ~n21047 & n21049;
  assign n21051 = pi770 & ~n21050;
  assign n21052 = ~n21046 & n21051;
  assign n21053 = pi726 & ~n21018;
  assign n21054 = ~n21052 & n21053;
  assign n21055 = n10178 & ~n21054;
  assign n21056 = ~n20970 & n21055;
  assign n21057 = ~pi147 & ~n10178;
  assign n21058 = ~pi832 & ~n21057;
  assign n21059 = ~n21056 & n21058;
  assign po304 = ~n20919 & ~n21059;
  assign n21061 = ~n9725 & ~n21022;
  assign n21062 = ~n16793 & ~n21036;
  assign n21063 = pi148 & ~n21062;
  assign n21064 = ~pi749 & ~n21063;
  assign n21065 = ~n21061 & n21064;
  assign n21066 = ~pi148 & n20990;
  assign n21067 = pi148 & n21006;
  assign n21068 = pi749 & ~n21067;
  assign n21069 = ~n21066 & n21068;
  assign n21070 = pi39 & ~n21065;
  assign n21071 = ~n21069 & n21070;
  assign n21072 = ~pi148 & ~n16655;
  assign n21073 = ~pi39 & ~n21072;
  assign n21074 = ~pi749 & pi947;
  assign n21075 = n20992 & ~n21074;
  assign n21076 = n21073 & ~n21075;
  assign n21077 = ~pi38 & ~n21076;
  assign n21078 = ~n21071 & n21077;
  assign n21079 = n21014 & ~n21074;
  assign n21080 = ~pi148 & ~n16968;
  assign n21081 = ~n21079 & ~n21080;
  assign n21082 = pi38 & ~n21081;
  assign n21083 = pi706 & ~n21082;
  assign n21084 = ~n21078 & n21083;
  assign n21085 = n3268 & n6294;
  assign n21086 = ~pi148 & ~n20933;
  assign n21087 = ~n20953 & ~n20960;
  assign n21088 = pi148 & ~n21087;
  assign n21089 = pi299 & ~n21088;
  assign n21090 = ~n21086 & n21089;
  assign n21091 = ~pi148 & ~n16792;
  assign n21092 = n20951 & ~n21091;
  assign n21093 = pi749 & ~n21092;
  assign n21094 = ~n21090 & n21093;
  assign n21095 = ~pi148 & ~pi749;
  assign n21096 = ~n16814 & n21095;
  assign n21097 = pi39 & ~n21096;
  assign n21098 = ~n21094 & n21097;
  assign n21099 = pi749 & pi947;
  assign n21100 = n16655 & n21099;
  assign n21101 = n21073 & ~n21100;
  assign n21102 = ~pi38 & ~n21101;
  assign n21103 = ~n21098 & n21102;
  assign n21104 = pi148 & ~n17485;
  assign n21105 = n16968 & ~n21099;
  assign n21106 = pi38 & ~n21105;
  assign n21107 = ~n21104 & n21106;
  assign n21108 = ~pi706 & ~n21107;
  assign n21109 = ~n21103 & n21108;
  assign n21110 = n21085 & ~n21109;
  assign n21111 = ~n21084 & n21110;
  assign n21112 = ~pi148 & ~n21085;
  assign n21113 = ~pi57 & ~n21112;
  assign n21114 = ~n21111 & n21113;
  assign n21115 = pi57 & pi148;
  assign n21116 = ~pi832 & ~n21115;
  assign n21117 = ~n21114 & n21116;
  assign n21118 = pi706 & n20848;
  assign n21119 = n2755 & ~n21099;
  assign n21120 = ~n21118 & n21119;
  assign n21121 = pi148 & ~n2755;
  assign n21122 = pi832 & ~n21121;
  assign n21123 = ~n21120 & n21122;
  assign po305 = n21117 | n21123;
  assign n21125 = ~pi755 & pi947;
  assign n21126 = ~pi725 & n20848;
  assign n21127 = ~n21125 & ~n21126;
  assign n21128 = n2755 & ~n21127;
  assign n21129 = ~pi149 & ~n2755;
  assign n21130 = pi832 & ~n21129;
  assign n21131 = ~n21128 & n21130;
  assign n21132 = pi149 & ~n17485;
  assign n21133 = n16968 & ~n21125;
  assign n21134 = pi38 & ~n21133;
  assign n21135 = ~n21132 & n21134;
  assign n21136 = ~pi149 & ~n20933;
  assign n21137 = ~n16095 & ~n20961;
  assign n21138 = ~n21136 & ~n21137;
  assign n21139 = ~pi149 & ~n16792;
  assign n21140 = n20951 & ~n21139;
  assign n21141 = ~pi755 & ~n21140;
  assign n21142 = ~n21138 & n21141;
  assign n21143 = ~pi149 & pi755;
  assign n21144 = ~n16814 & n21143;
  assign n21145 = pi39 & ~n21144;
  assign n21146 = ~n21142 & n21145;
  assign n21147 = ~pi149 & ~n16655;
  assign n21148 = n16655 & n21125;
  assign n21149 = ~pi39 & ~n21147;
  assign n21150 = ~n21148 & n21149;
  assign n21151 = ~pi38 & ~n21150;
  assign n21152 = ~n21146 & n21151;
  assign n21153 = ~n21135 & ~n21152;
  assign n21154 = pi725 & ~n21153;
  assign n21155 = ~n21041 & n21150;
  assign n21156 = ~pi149 & n20990;
  assign n21157 = pi149 & n21006;
  assign n21158 = ~pi755 & ~n21157;
  assign n21159 = ~n21156 & n21158;
  assign n21160 = ~pi149 & n21020;
  assign n21161 = pi149 & ~n21062;
  assign n21162 = pi755 & ~n21021;
  assign n21163 = ~n21161 & n21162;
  assign n21164 = ~n21160 & n21163;
  assign n21165 = pi39 & ~n21164;
  assign n21166 = ~n21159 & n21165;
  assign n21167 = ~n21155 & ~n21166;
  assign n21168 = ~pi38 & ~n21167;
  assign n21169 = ~pi149 & ~n16968;
  assign n21170 = ~n6217 & n16665;
  assign n21171 = pi755 & pi947;
  assign n21172 = ~pi39 & ~n21171;
  assign n21173 = n21170 & n21172;
  assign n21174 = pi38 & ~n21169;
  assign n21175 = ~n21173 & n21174;
  assign n21176 = ~pi725 & ~n21175;
  assign n21177 = ~n21168 & n21176;
  assign n21178 = ~n21154 & ~n21177;
  assign n21179 = n10178 & ~n21178;
  assign n21180 = ~pi149 & ~n10178;
  assign n21181 = ~pi832 & ~n21180;
  assign n21182 = ~n21179 & n21181;
  assign po306 = ~n21131 & ~n21182;
  assign n21184 = ~pi150 & n20936;
  assign n21185 = pi150 & ~n20962;
  assign n21186 = ~pi751 & ~n21185;
  assign n21187 = ~n21184 & n21186;
  assign n21188 = ~pi150 & pi751;
  assign n21189 = ~n16814 & n21188;
  assign n21190 = ~n21187 & ~n21189;
  assign n21191 = pi39 & ~n21190;
  assign n21192 = pi150 & ~n16655;
  assign n21193 = pi751 & n16655;
  assign n21194 = ~n21192 & ~n21193;
  assign n21195 = n20921 & n21194;
  assign n21196 = ~pi38 & ~n21195;
  assign n21197 = ~n21191 & n21196;
  assign n21198 = pi150 & ~n17485;
  assign n21199 = ~pi751 & pi947;
  assign n21200 = n16968 & ~n21199;
  assign n21201 = ~n21198 & ~n21200;
  assign n21202 = pi38 & ~n21201;
  assign n21203 = pi701 & ~n21202;
  assign n21204 = ~n21197 & n21203;
  assign n21205 = ~pi150 & ~n21022;
  assign n21206 = pi150 & ~n21039;
  assign n21207 = pi751 & ~n21206;
  assign n21208 = ~n21205 & n21207;
  assign n21209 = ~pi150 & n20990;
  assign n21210 = pi150 & n21006;
  assign n21211 = ~pi751 & ~n21210;
  assign n21212 = ~n21209 & n21211;
  assign n21213 = ~n21208 & ~n21212;
  assign n21214 = pi39 & ~n21213;
  assign n21215 = n21024 & ~n21199;
  assign n21216 = ~pi39 & ~n21192;
  assign n21217 = ~n21215 & n21216;
  assign n21218 = ~pi38 & ~n21217;
  assign n21219 = ~n21214 & n21218;
  assign n21220 = ~pi150 & ~n16968;
  assign n21221 = pi751 & pi947;
  assign n21222 = ~pi39 & ~n21221;
  assign n21223 = n21170 & n21222;
  assign n21224 = pi38 & ~n21220;
  assign n21225 = ~n21223 & n21224;
  assign n21226 = ~pi701 & ~n21225;
  assign n21227 = ~n21219 & n21226;
  assign n21228 = ~n21204 & ~n21227;
  assign n21229 = n10178 & ~n21228;
  assign n21230 = ~pi150 & ~n10178;
  assign n21231 = ~pi832 & ~n21230;
  assign n21232 = ~n21229 & n21231;
  assign n21233 = ~pi701 & n20848;
  assign n21234 = ~n21199 & ~n21233;
  assign n21235 = n2755 & ~n21234;
  assign n21236 = ~pi150 & ~n2755;
  assign n21237 = pi832 & ~n21236;
  assign n21238 = ~n21235 & n21237;
  assign po307 = ~n21232 & ~n21238;
  assign n21240 = ~pi745 & pi947;
  assign n21241 = ~pi723 & n20848;
  assign n21242 = ~n21240 & ~n21241;
  assign n21243 = n2755 & ~n21242;
  assign n21244 = ~pi151 & ~n2755;
  assign n21245 = pi832 & ~n21244;
  assign n21246 = ~n21243 & n21245;
  assign n21247 = ~pi151 & ~n16655;
  assign n21248 = ~pi745 & n20948;
  assign n21249 = ~n21247 & ~n21248;
  assign n21250 = n21042 & n21249;
  assign n21251 = ~n16809 & ~n20931;
  assign n21252 = ~pi151 & n21251;
  assign n21253 = ~n16805 & ~n21252;
  assign n21254 = pi215 & ~n21253;
  assign n21255 = pi151 & ~n3461;
  assign n21256 = ~n16801 & n21255;
  assign n21257 = ~n16798 & ~n21256;
  assign n21258 = ~pi151 & ~n16661;
  assign n21259 = n21032 & ~n21258;
  assign n21260 = ~n21000 & n21259;
  assign n21261 = ~pi215 & ~n21260;
  assign n21262 = n21257 & n21261;
  assign n21263 = ~n21254 & ~n21262;
  assign n21264 = pi299 & ~n21263;
  assign n21265 = pi151 & ~n20997;
  assign n21266 = n20987 & ~n21265;
  assign n21267 = ~n21264 & ~n21266;
  assign n21268 = ~pi745 & ~n21267;
  assign n21269 = n21257 & ~n21259;
  assign n21270 = n20974 & n21269;
  assign n21271 = ~n21254 & ~n21270;
  assign n21272 = ~n20953 & ~n21271;
  assign n21273 = pi299 & ~n21272;
  assign n21274 = ~pi151 & ~n16792;
  assign n21275 = n21038 & ~n21274;
  assign n21276 = pi745 & ~n21275;
  assign n21277 = ~n21273 & n21276;
  assign n21278 = pi39 & ~n21277;
  assign n21279 = ~n21268 & n21278;
  assign n21280 = ~n21250 & ~n21279;
  assign n21281 = ~pi38 & ~n21280;
  assign n21282 = ~pi151 & ~n16968;
  assign n21283 = pi745 & pi947;
  assign n21284 = ~pi39 & ~n21283;
  assign n21285 = n21170 & n21284;
  assign n21286 = pi38 & ~n21282;
  assign n21287 = ~n21285 & n21286;
  assign n21288 = ~pi723 & ~n21287;
  assign n21289 = ~n21281 & n21288;
  assign n21290 = ~pi745 & ~n16793;
  assign n21291 = ~pi151 & ~n16814;
  assign n21292 = ~n21290 & n21291;
  assign n21293 = n20958 & ~n21258;
  assign n21294 = n21257 & ~n21293;
  assign n21295 = n20928 & n21294;
  assign n21296 = n21028 & ~n21253;
  assign n21297 = pi299 & ~n21296;
  assign n21298 = ~n21295 & n21297;
  assign n21299 = ~pi745 & ~n20951;
  assign n21300 = ~n21298 & n21299;
  assign n21301 = ~n21292 & ~n21300;
  assign n21302 = pi39 & ~n21301;
  assign n21303 = ~pi39 & ~n21249;
  assign n21304 = ~pi38 & ~n21303;
  assign n21305 = ~n21302 & n21304;
  assign n21306 = pi151 & ~n17485;
  assign n21307 = n16968 & ~n21240;
  assign n21308 = ~n21306 & ~n21307;
  assign n21309 = pi38 & ~n21308;
  assign n21310 = pi723 & ~n21309;
  assign n21311 = ~n21305 & n21310;
  assign n21312 = ~n21289 & ~n21311;
  assign n21313 = n10178 & ~n21312;
  assign n21314 = ~pi151 & ~n10178;
  assign n21315 = ~pi832 & ~n21314;
  assign n21316 = ~n21313 & n21315;
  assign po308 = ~n21246 & ~n21316;
  assign n21318 = pi152 & ~n16661;
  assign n21319 = ~n21000 & ~n21318;
  assign n21320 = n3461 & n21319;
  assign n21321 = ~pi215 & ~n21320;
  assign n21322 = pi152 & n20972;
  assign n21323 = n21029 & ~n21322;
  assign n21324 = ~n16801 & n21323;
  assign n21325 = n21321 & ~n21324;
  assign n21326 = ~pi152 & ~n16805;
  assign n21327 = n20930 & ~n21326;
  assign n21328 = pi299 & ~n21327;
  assign n21329 = ~n21325 & n21328;
  assign n21330 = ~pi152 & ~n16787;
  assign n21331 = ~pi947 & n16787;
  assign n21332 = ~n3053 & ~n21331;
  assign n21333 = ~n21330 & n21332;
  assign n21334 = ~n6217 & n16787;
  assign n21335 = ~n3053 & ~n21334;
  assign n21336 = ~n21333 & n21335;
  assign n21337 = n3053 & n21319;
  assign n21338 = ~pi223 & ~n21337;
  assign n21339 = ~n21336 & n21338;
  assign n21340 = ~pi152 & ~n16728;
  assign n21341 = n20984 & ~n21340;
  assign n21342 = n20982 & ~n21340;
  assign n21343 = ~pi299 & ~n21342;
  assign n21344 = ~n21341 & n21343;
  assign n21345 = ~n21339 & n21344;
  assign n21346 = pi759 & ~n21329;
  assign n21347 = ~n21345 & n21346;
  assign n21348 = ~n21031 & ~n21318;
  assign n21349 = n3053 & ~n21348;
  assign n21350 = n16787 & ~n20848;
  assign n21351 = ~n3053 & ~n21350;
  assign n21352 = ~n21330 & n21351;
  assign n21353 = ~n21349 & ~n21352;
  assign n21354 = ~pi223 & ~n21353;
  assign n21355 = ~pi299 & ~n21341;
  assign n21356 = ~n21354 & n21355;
  assign n21357 = ~n20971 & n21321;
  assign n21358 = ~n21323 & n21357;
  assign n21359 = ~n20848 & ~n20999;
  assign n21360 = n21327 & ~n21359;
  assign n21361 = pi299 & ~n21360;
  assign n21362 = ~n21358 & n21361;
  assign n21363 = ~pi759 & ~n21362;
  assign n21364 = ~n21356 & n21363;
  assign n21365 = pi39 & ~n21364;
  assign n21366 = ~n21347 & n21365;
  assign n21367 = pi152 & ~n16655;
  assign n21368 = pi759 & pi947;
  assign n21369 = ~pi39 & ~n21368;
  assign n21370 = ~n16656 & ~n21369;
  assign n21371 = ~n21367 & ~n21370;
  assign n21372 = ~n21041 & n21371;
  assign n21373 = ~pi38 & ~n21372;
  assign n21374 = ~n21366 & n21373;
  assign n21375 = ~pi152 & ~n16968;
  assign n21376 = n16665 & ~n20848;
  assign n21377 = n21369 & n21376;
  assign n21378 = pi38 & ~n21375;
  assign n21379 = ~n21377 & n21378;
  assign n21380 = pi696 & ~n21379;
  assign n21381 = ~n21374 & n21380;
  assign n21382 = ~n20927 & ~n21323;
  assign n21383 = ~n20955 & ~n21382;
  assign n21384 = ~n20957 & ~n21318;
  assign n21385 = n3461 & n21384;
  assign n21386 = ~pi215 & ~n21385;
  assign n21387 = ~n21383 & n21386;
  assign n21388 = pi152 & n20932;
  assign n21389 = n20954 & ~n21388;
  assign n21390 = ~n21387 & n21389;
  assign n21391 = n3053 & ~n21384;
  assign n21392 = ~n21333 & ~n21391;
  assign n21393 = ~pi223 & ~n21392;
  assign n21394 = n21343 & ~n21393;
  assign n21395 = pi759 & ~n21394;
  assign n21396 = ~n21390 & n21395;
  assign n21397 = ~pi759 & ~n16814;
  assign n21398 = pi152 & n21397;
  assign n21399 = pi39 & ~n21398;
  assign n21400 = ~n21396 & n21399;
  assign n21401 = ~pi38 & ~n21371;
  assign n21402 = ~n21400 & n21401;
  assign n21403 = ~pi152 & ~n17485;
  assign n21404 = n16968 & ~n21368;
  assign n21405 = pi38 & ~n21404;
  assign n21406 = ~n21403 & n21405;
  assign n21407 = ~pi696 & ~n21406;
  assign n21408 = ~n21402 & n21407;
  assign n21409 = ~n21381 & ~n21408;
  assign n21410 = n10178 & ~n21409;
  assign n21411 = ~pi152 & ~n10178;
  assign n21412 = ~pi832 & ~n21411;
  assign n21413 = ~n21410 & n21412;
  assign n21414 = pi696 & n20848;
  assign n21415 = n2755 & ~n21368;
  assign n21416 = ~n21414 & n21415;
  assign n21417 = ~pi152 & ~n2755;
  assign n21418 = pi832 & ~n21417;
  assign n21419 = ~n21416 & n21418;
  assign po309 = n21413 | n21419;
  assign n21421 = pi766 & pi947;
  assign n21422 = n2755 & ~n21421;
  assign n21423 = pi700 & n20848;
  assign n21424 = n21422 & ~n21423;
  assign n21425 = pi153 & ~n2755;
  assign n21426 = pi832 & ~n21425;
  assign n21427 = ~n21424 & n21426;
  assign n21428 = ~pi153 & ~n16655;
  assign n21429 = ~pi766 & n18015;
  assign n21430 = ~n20949 & ~n21429;
  assign n21431 = ~n21428 & ~n21430;
  assign n21432 = ~n21041 & n21431;
  assign n21433 = pi153 & ~n16805;
  assign n21434 = n20930 & ~n21433;
  assign n21435 = pi153 & ~n3461;
  assign n21436 = ~n16801 & n21435;
  assign n21437 = ~n16798 & ~n21436;
  assign n21438 = ~pi153 & ~n16661;
  assign n21439 = n20958 & ~n21438;
  assign n21440 = ~n21030 & n21439;
  assign n21441 = ~pi215 & ~n21440;
  assign n21442 = n21437 & n21441;
  assign n21443 = ~n21434 & ~n21442;
  assign n21444 = pi299 & ~n21443;
  assign n21445 = pi153 & ~n20997;
  assign n21446 = n20987 & ~n21445;
  assign n21447 = ~n21444 & ~n21446;
  assign n21448 = pi766 & ~n21447;
  assign n21449 = n21032 & ~n21438;
  assign n21450 = ~n20973 & ~n21449;
  assign n21451 = n21437 & n21450;
  assign n21452 = ~pi215 & ~n21451;
  assign n21453 = n20999 & ~n21434;
  assign n21454 = ~n20953 & ~n21453;
  assign n21455 = ~n21452 & n21454;
  assign n21456 = pi299 & ~n21455;
  assign n21457 = ~pi153 & ~n16792;
  assign n21458 = n21038 & ~n21457;
  assign n21459 = ~pi766 & ~n21458;
  assign n21460 = ~n21456 & n21459;
  assign n21461 = pi39 & ~n21460;
  assign n21462 = ~n21448 & n21461;
  assign n21463 = ~n21432 & ~n21462;
  assign n21464 = ~pi38 & ~n21463;
  assign n21465 = ~pi153 & ~n16968;
  assign n21466 = ~pi766 & pi947;
  assign n21467 = ~pi39 & ~n21466;
  assign n21468 = n21170 & n21467;
  assign n21469 = pi38 & ~n21465;
  assign n21470 = ~n21468 & n21469;
  assign n21471 = ~n21464 & ~n21470;
  assign n21472 = pi700 & ~n21471;
  assign n21473 = n20951 & ~n21457;
  assign n21474 = n21437 & ~n21439;
  assign n21475 = n20928 & n21474;
  assign n21476 = n20932 & ~n21433;
  assign n21477 = pi299 & ~n21476;
  assign n21478 = ~n21475 & n21477;
  assign n21479 = pi766 & ~n21478;
  assign n21480 = ~n21473 & n21479;
  assign n21481 = ~pi153 & ~pi766;
  assign n21482 = ~n16814 & n21481;
  assign n21483 = pi39 & ~n21482;
  assign n21484 = ~n21480 & n21483;
  assign n21485 = ~pi38 & ~n21431;
  assign n21486 = ~n21484 & n21485;
  assign n21487 = pi153 & ~n17485;
  assign n21488 = n6250 & n21422;
  assign n21489 = pi38 & ~n21488;
  assign n21490 = ~n21487 & n21489;
  assign n21491 = ~pi700 & ~n21490;
  assign n21492 = ~n21486 & n21491;
  assign n21493 = n21085 & ~n21492;
  assign n21494 = ~n21472 & n21493;
  assign n21495 = ~pi153 & ~n21085;
  assign n21496 = ~pi57 & ~n21495;
  assign n21497 = ~n21494 & n21496;
  assign n21498 = pi57 & pi153;
  assign n21499 = ~pi832 & ~n21498;
  assign n21500 = ~n21497 & n21499;
  assign po310 = n21427 | n21500;
  assign n21502 = ~pi742 & pi947;
  assign n21503 = ~pi704 & n20848;
  assign n21504 = ~n21502 & ~n21503;
  assign n21505 = n2755 & ~n21504;
  assign n21506 = ~pi154 & ~n2755;
  assign n21507 = pi832 & ~n21506;
  assign n21508 = ~n21505 & n21507;
  assign n21509 = ~pi154 & ~n16655;
  assign n21510 = n21042 & ~n21509;
  assign n21511 = ~pi154 & n21022;
  assign n21512 = pi154 & n21039;
  assign n21513 = pi39 & ~n21512;
  assign n21514 = ~n21511 & n21513;
  assign n21515 = ~n21510 & ~n21514;
  assign n21516 = ~pi38 & ~n21515;
  assign n21517 = ~pi154 & ~n16968;
  assign n21518 = n21049 & ~n21517;
  assign n21519 = pi742 & ~n21518;
  assign n21520 = ~n21516 & n21519;
  assign n21521 = ~n20992 & n21510;
  assign n21522 = ~pi154 & ~n20990;
  assign n21523 = pi154 & ~n21006;
  assign n21524 = pi39 & ~n21523;
  assign n21525 = ~n21522 & n21524;
  assign n21526 = ~n21521 & ~n21525;
  assign n21527 = ~pi38 & ~n21526;
  assign n21528 = n21015 & ~n21517;
  assign n21529 = ~pi742 & ~n21528;
  assign n21530 = ~n21527 & n21529;
  assign n21531 = ~pi704 & ~n21520;
  assign n21532 = ~n21530 & n21531;
  assign n21533 = n20949 & ~n21509;
  assign n21534 = ~pi154 & ~n20936;
  assign n21535 = pi154 & n20962;
  assign n21536 = pi39 & ~n21535;
  assign n21537 = ~n21534 & n21536;
  assign n21538 = ~n21533 & ~n21537;
  assign n21539 = ~pi38 & ~n21538;
  assign n21540 = ~pi154 & ~n17485;
  assign n21541 = ~n20947 & ~n21540;
  assign n21542 = ~pi742 & ~n21541;
  assign n21543 = ~n21539 & n21542;
  assign n21544 = ~pi154 & pi742;
  assign n21545 = ~n17487 & n21544;
  assign n21546 = pi704 & ~n21545;
  assign n21547 = ~n21543 & n21546;
  assign n21548 = n10178 & ~n21547;
  assign n21549 = ~n21532 & n21548;
  assign n21550 = ~pi154 & ~n10178;
  assign n21551 = ~pi832 & ~n21550;
  assign n21552 = ~n21549 & n21551;
  assign po311 = ~n21508 & ~n21552;
  assign n21554 = ~pi38 & ~n21008;
  assign n21555 = ~n21015 & ~n21554;
  assign n21556 = ~pi757 & n21555;
  assign n21557 = ~pi38 & ~n21043;
  assign n21558 = ~n21049 & ~n21557;
  assign n21559 = pi757 & n21558;
  assign n21560 = ~pi686 & ~n21556;
  assign n21561 = ~n21559 & n21560;
  assign n21562 = ~pi757 & n20966;
  assign n21563 = pi686 & ~n21562;
  assign n21564 = n10178 & ~n21563;
  assign n21565 = ~n21561 & n21564;
  assign n21566 = pi155 & ~n21565;
  assign n21567 = ~pi38 & ~n20995;
  assign n21568 = pi38 & n21012;
  assign n21569 = ~n21567 & ~n21568;
  assign n21570 = ~pi757 & n21569;
  assign n21571 = ~pi38 & ~n21026;
  assign n21572 = n16968 & n21049;
  assign n21573 = ~n21571 & ~n21572;
  assign n21574 = pi757 & n21573;
  assign n21575 = ~pi686 & ~n21570;
  assign n21576 = ~n21574 & n21575;
  assign n21577 = ~pi757 & n20942;
  assign n21578 = pi757 & ~n17487;
  assign n21579 = pi686 & ~n21578;
  assign n21580 = ~n21577 & n21579;
  assign n21581 = ~n21576 & ~n21580;
  assign n21582 = ~pi155 & n10178;
  assign n21583 = ~n21581 & n21582;
  assign n21584 = ~n21566 & ~n21583;
  assign n21585 = ~pi832 & ~n21584;
  assign n21586 = ~pi757 & pi947;
  assign n21587 = ~pi686 & n20848;
  assign n21588 = ~n21586 & ~n21587;
  assign n21589 = n2755 & ~n21588;
  assign n21590 = ~pi155 & ~n2755;
  assign n21591 = pi832 & ~n21590;
  assign n21592 = ~n21589 & n21591;
  assign po312 = ~n21585 & ~n21592;
  assign n21594 = ~pi741 & pi947;
  assign n21595 = ~pi724 & n20848;
  assign n21596 = ~n21594 & ~n21595;
  assign n21597 = n2755 & ~n21596;
  assign n21598 = ~pi156 & ~n2755;
  assign n21599 = pi832 & ~n21598;
  assign n21600 = ~n21597 & n21599;
  assign n21601 = ~pi741 & ~n21569;
  assign n21602 = pi741 & ~n21573;
  assign n21603 = ~pi724 & ~n21601;
  assign n21604 = ~n21602 & n21603;
  assign n21605 = ~pi741 & ~n20942;
  assign n21606 = pi741 & n17487;
  assign n21607 = pi724 & ~n21606;
  assign n21608 = ~n21605 & n21607;
  assign n21609 = n10178 & ~n21608;
  assign n21610 = ~n21604 & n21609;
  assign n21611 = ~pi156 & ~n21610;
  assign n21612 = ~pi741 & ~n21555;
  assign n21613 = pi741 & ~n21558;
  assign n21614 = ~pi724 & ~n21612;
  assign n21615 = ~n21613 & n21614;
  assign n21616 = pi724 & ~pi741;
  assign n21617 = n20966 & n21616;
  assign n21618 = ~n21615 & ~n21617;
  assign n21619 = pi156 & n10178;
  assign n21620 = ~n21618 & n21619;
  assign n21621 = ~pi832 & ~n21620;
  assign n21622 = ~n21611 & n21621;
  assign po313 = ~n21600 & ~n21622;
  assign n21624 = ~pi760 & pi947;
  assign n21625 = ~pi688 & n20848;
  assign n21626 = ~n21624 & ~n21625;
  assign n21627 = n2755 & ~n21626;
  assign n21628 = ~pi157 & ~n2755;
  assign n21629 = pi832 & ~n21628;
  assign n21630 = ~n21627 & n21629;
  assign n21631 = pi157 & ~n17485;
  assign n21632 = n16968 & ~n21624;
  assign n21633 = pi38 & ~n21632;
  assign n21634 = ~n21631 & n21633;
  assign n21635 = ~pi157 & ~n20933;
  assign n21636 = ~n13776 & ~n20961;
  assign n21637 = ~n21635 & ~n21636;
  assign n21638 = ~pi157 & ~n16792;
  assign n21639 = n20951 & ~n21638;
  assign n21640 = ~pi760 & ~n21639;
  assign n21641 = ~n21637 & n21640;
  assign n21642 = ~pi157 & pi760;
  assign n21643 = ~n16814 & n21642;
  assign n21644 = pi39 & ~n21643;
  assign n21645 = ~n21641 & n21644;
  assign n21646 = ~pi157 & ~n16655;
  assign n21647 = n16655 & n21624;
  assign n21648 = ~pi39 & ~n21646;
  assign n21649 = ~n21647 & n21648;
  assign n21650 = ~pi38 & ~n21649;
  assign n21651 = ~n21645 & n21650;
  assign n21652 = ~n21634 & ~n21651;
  assign n21653 = pi688 & ~n21652;
  assign n21654 = ~n21041 & n21649;
  assign n21655 = pi760 & ~n21022;
  assign n21656 = ~pi760 & n20990;
  assign n21657 = ~pi157 & ~n21655;
  assign n21658 = ~n21656 & n21657;
  assign n21659 = ~pi760 & n21006;
  assign n21660 = pi760 & ~n21039;
  assign n21661 = pi157 & ~n21659;
  assign n21662 = ~n21660 & n21661;
  assign n21663 = pi39 & ~n21662;
  assign n21664 = ~n21658 & n21663;
  assign n21665 = ~n21654 & ~n21664;
  assign n21666 = ~pi38 & ~n21665;
  assign n21667 = ~pi157 & ~n16968;
  assign n21668 = pi760 & pi947;
  assign n21669 = ~pi39 & ~n21668;
  assign n21670 = n21170 & n21669;
  assign n21671 = pi38 & ~n21667;
  assign n21672 = ~n21670 & n21671;
  assign n21673 = ~pi688 & ~n21672;
  assign n21674 = ~n21666 & n21673;
  assign n21675 = ~n21653 & ~n21674;
  assign n21676 = n10178 & ~n21675;
  assign n21677 = ~pi157 & ~n10178;
  assign n21678 = ~pi832 & ~n21677;
  assign n21679 = ~n21676 & n21678;
  assign po314 = ~n21630 & ~n21679;
  assign n21681 = ~pi158 & n20936;
  assign n21682 = pi158 & ~n20962;
  assign n21683 = ~pi753 & ~n21682;
  assign n21684 = ~n21681 & n21683;
  assign n21685 = ~pi158 & pi753;
  assign n21686 = ~n16814 & n21685;
  assign n21687 = ~n21684 & ~n21686;
  assign n21688 = pi39 & ~n21687;
  assign n21689 = pi158 & ~n16655;
  assign n21690 = pi753 & n16655;
  assign n21691 = ~n21689 & ~n21690;
  assign n21692 = n20921 & n21691;
  assign n21693 = ~pi38 & ~n21692;
  assign n21694 = ~n21688 & n21693;
  assign n21695 = pi158 & ~n17485;
  assign n21696 = ~pi753 & pi947;
  assign n21697 = n16968 & ~n21696;
  assign n21698 = ~n21695 & ~n21697;
  assign n21699 = pi38 & ~n21698;
  assign n21700 = pi702 & ~n21699;
  assign n21701 = ~n21694 & n21700;
  assign n21702 = ~pi158 & ~n21022;
  assign n21703 = pi158 & ~n21039;
  assign n21704 = pi753 & ~n21703;
  assign n21705 = ~n21702 & n21704;
  assign n21706 = ~pi158 & n20990;
  assign n21707 = pi158 & n21006;
  assign n21708 = ~pi753 & ~n21707;
  assign n21709 = ~n21706 & n21708;
  assign n21710 = ~n21705 & ~n21709;
  assign n21711 = pi39 & ~n21710;
  assign n21712 = n21024 & ~n21696;
  assign n21713 = ~pi39 & ~n21689;
  assign n21714 = ~n21712 & n21713;
  assign n21715 = ~pi38 & ~n21714;
  assign n21716 = ~n21711 & n21715;
  assign n21717 = ~pi158 & ~n16968;
  assign n21718 = pi753 & pi947;
  assign n21719 = ~pi39 & ~n21718;
  assign n21720 = n21170 & n21719;
  assign n21721 = pi38 & ~n21717;
  assign n21722 = ~n21720 & n21721;
  assign n21723 = ~pi702 & ~n21722;
  assign n21724 = ~n21716 & n21723;
  assign n21725 = ~n21701 & ~n21724;
  assign n21726 = n10178 & ~n21725;
  assign n21727 = ~pi158 & ~n10178;
  assign n21728 = ~pi832 & ~n21727;
  assign n21729 = ~n21726 & n21728;
  assign n21730 = ~pi702 & n20848;
  assign n21731 = ~n21696 & ~n21730;
  assign n21732 = n2755 & ~n21731;
  assign n21733 = ~pi158 & ~n2755;
  assign n21734 = pi832 & ~n21733;
  assign n21735 = ~n21732 & n21734;
  assign po315 = ~n21729 & ~n21735;
  assign n21737 = ~pi159 & n20936;
  assign n21738 = pi159 & ~n20962;
  assign n21739 = ~pi754 & ~n21738;
  assign n21740 = ~n21737 & n21739;
  assign n21741 = ~pi159 & pi754;
  assign n21742 = ~n16814 & n21741;
  assign n21743 = ~n21740 & ~n21742;
  assign n21744 = pi39 & ~n21743;
  assign n21745 = pi159 & ~n16655;
  assign n21746 = pi754 & n16655;
  assign n21747 = ~n21745 & ~n21746;
  assign n21748 = n20921 & n21747;
  assign n21749 = ~pi38 & ~n21748;
  assign n21750 = ~n21744 & n21749;
  assign n21751 = pi159 & ~n17485;
  assign n21752 = ~pi754 & pi947;
  assign n21753 = n16968 & ~n21752;
  assign n21754 = ~n21751 & ~n21753;
  assign n21755 = pi38 & ~n21754;
  assign n21756 = pi709 & ~n21755;
  assign n21757 = ~n21750 & n21756;
  assign n21758 = ~pi159 & ~n21022;
  assign n21759 = pi159 & ~n21039;
  assign n21760 = pi754 & ~n21759;
  assign n21761 = ~n21758 & n21760;
  assign n21762 = ~pi159 & n20990;
  assign n21763 = pi159 & n21006;
  assign n21764 = ~pi754 & ~n21763;
  assign n21765 = ~n21762 & n21764;
  assign n21766 = ~n21761 & ~n21765;
  assign n21767 = pi39 & ~n21766;
  assign n21768 = n21024 & ~n21752;
  assign n21769 = ~pi39 & ~n21745;
  assign n21770 = ~n21768 & n21769;
  assign n21771 = ~pi38 & ~n21770;
  assign n21772 = ~n21767 & n21771;
  assign n21773 = ~pi159 & ~n16968;
  assign n21774 = pi754 & pi947;
  assign n21775 = ~pi39 & ~n21774;
  assign n21776 = n21170 & n21775;
  assign n21777 = pi38 & ~n21773;
  assign n21778 = ~n21776 & n21777;
  assign n21779 = ~pi709 & ~n21778;
  assign n21780 = ~n21772 & n21779;
  assign n21781 = ~n21757 & ~n21780;
  assign n21782 = n10178 & ~n21781;
  assign n21783 = ~pi159 & ~n10178;
  assign n21784 = ~pi832 & ~n21783;
  assign n21785 = ~n21782 & n21784;
  assign n21786 = ~pi709 & n20848;
  assign n21787 = ~n21752 & ~n21786;
  assign n21788 = n2755 & ~n21787;
  assign n21789 = ~pi159 & ~n2755;
  assign n21790 = pi832 & ~n21789;
  assign n21791 = ~n21788 & n21790;
  assign po316 = ~n21785 & ~n21791;
  assign n21793 = ~pi756 & pi947;
  assign n21794 = ~pi734 & n20848;
  assign n21795 = ~n21793 & ~n21794;
  assign n21796 = n2755 & ~n21795;
  assign n21797 = ~pi160 & ~n2755;
  assign n21798 = pi832 & ~n21797;
  assign n21799 = ~n21796 & n21798;
  assign n21800 = pi160 & ~n17485;
  assign n21801 = n16968 & ~n21793;
  assign n21802 = pi38 & ~n21801;
  assign n21803 = ~n21800 & n21802;
  assign n21804 = ~pi160 & ~n20933;
  assign n21805 = pi160 & ~n21087;
  assign n21806 = pi299 & ~n21805;
  assign n21807 = ~n21804 & n21806;
  assign n21808 = ~pi160 & ~n16792;
  assign n21809 = n20951 & ~n21808;
  assign n21810 = ~pi756 & ~n21809;
  assign n21811 = ~n21807 & n21810;
  assign n21812 = ~pi160 & pi756;
  assign n21813 = ~n16814 & n21812;
  assign n21814 = pi39 & ~n21813;
  assign n21815 = ~n21811 & n21814;
  assign n21816 = ~pi160 & ~n16655;
  assign n21817 = n16655 & n21793;
  assign n21818 = ~pi39 & ~n21816;
  assign n21819 = ~n21817 & n21818;
  assign n21820 = ~pi38 & ~n21819;
  assign n21821 = ~n21815 & n21820;
  assign n21822 = ~n21803 & ~n21821;
  assign n21823 = pi734 & ~n21822;
  assign n21824 = ~n21041 & n21819;
  assign n21825 = ~pi160 & n20990;
  assign n21826 = pi160 & n21006;
  assign n21827 = ~pi756 & ~n21826;
  assign n21828 = ~n21825 & n21827;
  assign n21829 = ~pi160 & n21020;
  assign n21830 = pi160 & ~n21062;
  assign n21831 = pi756 & ~n21021;
  assign n21832 = ~n21830 & n21831;
  assign n21833 = ~n21829 & n21832;
  assign n21834 = pi39 & ~n21833;
  assign n21835 = ~n21828 & n21834;
  assign n21836 = ~n21824 & ~n21835;
  assign n21837 = ~pi38 & ~n21836;
  assign n21838 = ~pi160 & ~n16968;
  assign n21839 = pi756 & pi947;
  assign n21840 = ~pi39 & ~n21839;
  assign n21841 = n21170 & n21840;
  assign n21842 = pi38 & ~n21838;
  assign n21843 = ~n21841 & n21842;
  assign n21844 = ~pi734 & ~n21843;
  assign n21845 = ~n21837 & n21844;
  assign n21846 = ~n21823 & ~n21845;
  assign n21847 = n10178 & ~n21846;
  assign n21848 = ~pi160 & ~n10178;
  assign n21849 = ~pi832 & ~n21848;
  assign n21850 = ~n21847 & n21849;
  assign po317 = ~n21799 & ~n21850;
  assign n21852 = pi161 & ~n16661;
  assign n21853 = ~n21000 & ~n21852;
  assign n21854 = n3461 & n21853;
  assign n21855 = ~pi215 & ~n21854;
  assign n21856 = pi161 & n20972;
  assign n21857 = n21029 & ~n21856;
  assign n21858 = ~n16801 & n21857;
  assign n21859 = n21855 & ~n21858;
  assign n21860 = ~pi161 & ~n16805;
  assign n21861 = n20930 & ~n21860;
  assign n21862 = pi299 & ~n21861;
  assign n21863 = ~n21859 & n21862;
  assign n21864 = ~pi161 & ~n16787;
  assign n21865 = n21332 & ~n21864;
  assign n21866 = n21335 & ~n21865;
  assign n21867 = n3053 & n21853;
  assign n21868 = ~pi223 & ~n21867;
  assign n21869 = ~n21866 & n21868;
  assign n21870 = ~pi161 & ~n16728;
  assign n21871 = n20984 & ~n21870;
  assign n21872 = n20982 & ~n21870;
  assign n21873 = ~pi299 & ~n21872;
  assign n21874 = ~n21871 & n21873;
  assign n21875 = ~n21869 & n21874;
  assign n21876 = pi758 & ~n21863;
  assign n21877 = ~n21875 & n21876;
  assign n21878 = ~n21031 & ~n21852;
  assign n21879 = n3053 & ~n21878;
  assign n21880 = n21351 & ~n21864;
  assign n21881 = ~n21879 & ~n21880;
  assign n21882 = ~pi223 & ~n21881;
  assign n21883 = ~pi299 & ~n21871;
  assign n21884 = ~n21882 & n21883;
  assign n21885 = ~n20971 & n21855;
  assign n21886 = ~n21857 & n21885;
  assign n21887 = ~n21359 & n21861;
  assign n21888 = pi299 & ~n21887;
  assign n21889 = ~n21886 & n21888;
  assign n21890 = ~pi758 & ~n21889;
  assign n21891 = ~n21884 & n21890;
  assign n21892 = pi39 & ~n21891;
  assign n21893 = ~n21877 & n21892;
  assign n21894 = pi161 & ~n16655;
  assign n21895 = pi758 & pi947;
  assign n21896 = ~pi39 & ~n21895;
  assign n21897 = ~n16656 & ~n21896;
  assign n21898 = ~n21894 & ~n21897;
  assign n21899 = ~n21041 & n21898;
  assign n21900 = ~pi38 & ~n21899;
  assign n21901 = ~n21893 & n21900;
  assign n21902 = ~pi161 & ~n16968;
  assign n21903 = n21376 & n21896;
  assign n21904 = pi38 & ~n21902;
  assign n21905 = ~n21903 & n21904;
  assign n21906 = pi736 & ~n21905;
  assign n21907 = ~n21901 & n21906;
  assign n21908 = ~n20927 & ~n21857;
  assign n21909 = ~n20955 & ~n21908;
  assign n21910 = ~n20957 & ~n21852;
  assign n21911 = n3461 & n21910;
  assign n21912 = ~pi215 & ~n21911;
  assign n21913 = ~n21909 & n21912;
  assign n21914 = pi161 & n20932;
  assign n21915 = n20954 & ~n21914;
  assign n21916 = ~n21913 & n21915;
  assign n21917 = n3053 & ~n21910;
  assign n21918 = ~n21865 & ~n21917;
  assign n21919 = ~pi223 & ~n21918;
  assign n21920 = n21873 & ~n21919;
  assign n21921 = pi758 & ~n21920;
  assign n21922 = ~n21916 & n21921;
  assign n21923 = pi161 & n19829;
  assign n21924 = pi39 & ~n21923;
  assign n21925 = ~n21922 & n21924;
  assign n21926 = ~pi38 & ~n21898;
  assign n21927 = ~n21925 & n21926;
  assign n21928 = ~pi161 & ~n17485;
  assign n21929 = n16968 & ~n21895;
  assign n21930 = pi38 & ~n21929;
  assign n21931 = ~n21928 & n21930;
  assign n21932 = ~pi736 & ~n21931;
  assign n21933 = ~n21927 & n21932;
  assign n21934 = ~n21907 & ~n21933;
  assign n21935 = n10178 & ~n21934;
  assign n21936 = ~pi161 & ~n10178;
  assign n21937 = ~pi832 & ~n21936;
  assign n21938 = ~n21935 & n21937;
  assign n21939 = pi736 & n20848;
  assign n21940 = n2755 & ~n21895;
  assign n21941 = ~n21939 & n21940;
  assign n21942 = ~pi161 & ~n2755;
  assign n21943 = pi832 & ~n21942;
  assign n21944 = ~n21941 & n21943;
  assign po318 = n21938 | n21944;
  assign n21946 = pi162 & ~n17485;
  assign n21947 = ~pi761 & pi947;
  assign n21948 = n16968 & ~n21947;
  assign n21949 = pi38 & ~n21948;
  assign n21950 = ~n21946 & n21949;
  assign n21951 = ~pi761 & n20935;
  assign n21952 = pi761 & n16814;
  assign n21953 = ~pi162 & ~n21952;
  assign n21954 = ~n21951 & n21953;
  assign n21955 = n15080 & ~n21087;
  assign n21956 = ~n20923 & ~n21955;
  assign n21957 = ~pi761 & ~n21956;
  assign n21958 = pi39 & ~n21957;
  assign n21959 = ~n21954 & n21958;
  assign n21960 = ~pi162 & ~n16655;
  assign n21961 = n16655 & n21947;
  assign n21962 = ~pi39 & ~n21960;
  assign n21963 = ~n21961 & n21962;
  assign n21964 = ~pi38 & ~n21963;
  assign n21965 = ~n21959 & n21964;
  assign n21966 = ~n21950 & ~n21965;
  assign n21967 = pi738 & ~n21966;
  assign n21968 = ~n21041 & n21963;
  assign n21969 = ~n15080 & ~n21022;
  assign n21970 = pi162 & ~n21062;
  assign n21971 = pi761 & ~n21970;
  assign n21972 = ~n21969 & n21971;
  assign n21973 = ~pi162 & n20990;
  assign n21974 = pi162 & n21006;
  assign n21975 = ~pi761 & ~n21974;
  assign n21976 = ~n21973 & n21975;
  assign n21977 = pi39 & ~n21972;
  assign n21978 = ~n21976 & n21977;
  assign n21979 = ~n21968 & ~n21978;
  assign n21980 = ~pi38 & ~n21979;
  assign n21981 = ~pi162 & ~n16968;
  assign n21982 = pi761 & pi947;
  assign n21983 = ~pi39 & ~n21982;
  assign n21984 = n21170 & n21983;
  assign n21985 = pi38 & ~n21981;
  assign n21986 = ~n21984 & n21985;
  assign n21987 = ~pi738 & ~n21986;
  assign n21988 = ~n21980 & n21987;
  assign n21989 = ~n21967 & ~n21988;
  assign n21990 = n10178 & ~n21989;
  assign n21991 = ~pi162 & ~n10178;
  assign n21992 = ~pi832 & ~n21991;
  assign n21993 = ~n21990 & n21992;
  assign n21994 = ~pi738 & n20848;
  assign n21995 = ~n21947 & ~n21994;
  assign n21996 = n2755 & ~n21995;
  assign n21997 = ~pi162 & ~n2755;
  assign n21998 = pi832 & ~n21997;
  assign n21999 = ~n21996 & n21998;
  assign po319 = ~n21993 & ~n21999;
  assign n22001 = ~pi777 & pi947;
  assign n22002 = ~pi737 & n20848;
  assign n22003 = ~n22001 & ~n22002;
  assign n22004 = n2755 & ~n22003;
  assign n22005 = ~pi163 & ~n2755;
  assign n22006 = pi832 & ~n22005;
  assign n22007 = ~n22004 & n22006;
  assign n22008 = pi163 & ~n17485;
  assign n22009 = n16968 & ~n22001;
  assign n22010 = pi38 & ~n22009;
  assign n22011 = ~n22008 & n22010;
  assign n22012 = ~pi163 & ~n20933;
  assign n22013 = ~n14689 & ~n20961;
  assign n22014 = ~n22012 & ~n22013;
  assign n22015 = ~pi163 & ~n16792;
  assign n22016 = n20951 & ~n22015;
  assign n22017 = ~pi777 & ~n22016;
  assign n22018 = ~n22014 & n22017;
  assign n22019 = ~pi163 & pi777;
  assign n22020 = ~n16814 & n22019;
  assign n22021 = pi39 & ~n22020;
  assign n22022 = ~n22018 & n22021;
  assign n22023 = ~pi163 & ~n16655;
  assign n22024 = n16655 & n22001;
  assign n22025 = ~pi39 & ~n22023;
  assign n22026 = ~n22024 & n22025;
  assign n22027 = ~pi38 & ~n22026;
  assign n22028 = ~n22022 & n22027;
  assign n22029 = ~n22011 & ~n22028;
  assign n22030 = pi737 & ~n22029;
  assign n22031 = ~n21041 & n22026;
  assign n22032 = ~pi163 & n20990;
  assign n22033 = pi163 & n21006;
  assign n22034 = ~pi777 & ~n22033;
  assign n22035 = ~n22032 & n22034;
  assign n22036 = ~pi163 & n21020;
  assign n22037 = pi163 & ~n21062;
  assign n22038 = pi777 & ~n21021;
  assign n22039 = ~n22037 & n22038;
  assign n22040 = ~n22036 & n22039;
  assign n22041 = pi39 & ~n22040;
  assign n22042 = ~n22035 & n22041;
  assign n22043 = ~n22031 & ~n22042;
  assign n22044 = ~pi38 & ~n22043;
  assign n22045 = ~pi163 & ~n16968;
  assign n22046 = pi777 & pi947;
  assign n22047 = ~pi39 & ~n22046;
  assign n22048 = n21170 & n22047;
  assign n22049 = pi38 & ~n22045;
  assign n22050 = ~n22048 & n22049;
  assign n22051 = ~pi737 & ~n22050;
  assign n22052 = ~n22044 & n22051;
  assign n22053 = ~n22030 & ~n22052;
  assign n22054 = n10178 & ~n22053;
  assign n22055 = ~pi163 & ~n10178;
  assign n22056 = ~pi832 & ~n22055;
  assign n22057 = ~n22054 & n22056;
  assign po320 = ~n22007 & ~n22057;
  assign n22059 = ~pi752 & pi947;
  assign n22060 = pi703 & n20848;
  assign n22061 = ~n22059 & ~n22060;
  assign n22062 = n2755 & ~n22061;
  assign n22063 = ~pi164 & ~n2755;
  assign n22064 = pi832 & ~n22063;
  assign n22065 = ~n22062 & n22064;
  assign n22066 = ~pi164 & n20995;
  assign n22067 = pi164 & n21008;
  assign n22068 = ~pi38 & ~n22067;
  assign n22069 = ~n22066 & n22068;
  assign n22070 = ~pi164 & ~n21012;
  assign n22071 = n21015 & ~n22070;
  assign n22072 = ~pi752 & ~n22071;
  assign n22073 = ~n22069 & n22072;
  assign n22074 = ~pi164 & n21026;
  assign n22075 = pi164 & n21043;
  assign n22076 = ~pi38 & ~n22075;
  assign n22077 = ~n22074 & n22076;
  assign n22078 = ~pi164 & ~n16968;
  assign n22079 = n21049 & ~n22078;
  assign n22080 = pi752 & ~n22079;
  assign n22081 = ~n22077 & n22080;
  assign n22082 = ~n22073 & ~n22081;
  assign n22083 = pi703 & ~n22082;
  assign n22084 = pi164 & ~n20941;
  assign n22085 = ~pi752 & ~n22084;
  assign n22086 = ~n20942 & n22085;
  assign n22087 = ~pi752 & n20966;
  assign n22088 = pi164 & ~n22087;
  assign n22089 = pi752 & n17487;
  assign n22090 = ~pi703 & ~n22089;
  assign n22091 = ~n22088 & n22090;
  assign n22092 = ~n22086 & n22091;
  assign n22093 = ~n22083 & ~n22092;
  assign n22094 = n10178 & ~n22093;
  assign n22095 = ~pi164 & ~n10178;
  assign n22096 = ~pi832 & ~n22095;
  assign n22097 = ~n22094 & n22096;
  assign po321 = ~n22065 & ~n22097;
  assign n22099 = ~pi774 & pi947;
  assign n22100 = pi687 & n20848;
  assign n22101 = ~n22099 & ~n22100;
  assign n22102 = n2755 & ~n22101;
  assign n22103 = ~pi165 & ~n2755;
  assign n22104 = pi832 & ~n22103;
  assign n22105 = ~n22102 & n22104;
  assign n22106 = ~pi165 & n20995;
  assign n22107 = pi165 & n21008;
  assign n22108 = ~pi38 & ~n22107;
  assign n22109 = ~n22106 & n22108;
  assign n22110 = ~pi165 & ~n21012;
  assign n22111 = n21015 & ~n22110;
  assign n22112 = ~pi774 & ~n22111;
  assign n22113 = ~n22109 & n22112;
  assign n22114 = ~pi165 & n21026;
  assign n22115 = pi165 & n21043;
  assign n22116 = ~pi38 & ~n22115;
  assign n22117 = ~n22114 & n22116;
  assign n22118 = ~pi165 & ~n16968;
  assign n22119 = n21049 & ~n22118;
  assign n22120 = pi774 & ~n22119;
  assign n22121 = ~n22117 & n22120;
  assign n22122 = ~n22113 & ~n22121;
  assign n22123 = pi687 & ~n22122;
  assign n22124 = pi165 & ~n20941;
  assign n22125 = ~pi774 & ~n22124;
  assign n22126 = ~n20942 & n22125;
  assign n22127 = ~pi774 & n20966;
  assign n22128 = pi165 & ~n22127;
  assign n22129 = pi774 & n17487;
  assign n22130 = ~pi687 & ~n22129;
  assign n22131 = ~n22128 & n22130;
  assign n22132 = ~n22126 & n22131;
  assign n22133 = ~n22123 & ~n22132;
  assign n22134 = n10178 & ~n22133;
  assign n22135 = ~pi165 & ~n10178;
  assign n22136 = ~pi832 & ~n22135;
  assign n22137 = ~n22134 & n22136;
  assign po322 = ~n22105 & ~n22137;
  assign n22139 = pi166 & n20972;
  assign n22140 = n21029 & ~n22139;
  assign n22141 = ~n20927 & ~n22140;
  assign n22142 = ~n20955 & ~n22141;
  assign n22143 = pi166 & ~n16661;
  assign n22144 = ~n20957 & ~n22143;
  assign n22145 = n3461 & n22144;
  assign n22146 = ~pi215 & ~n22145;
  assign n22147 = ~n22142 & n22146;
  assign n22148 = pi166 & n20932;
  assign n22149 = n20954 & ~n22148;
  assign n22150 = ~n22147 & n22149;
  assign n22151 = ~pi166 & ~n16728;
  assign n22152 = n20982 & ~n22151;
  assign n22153 = ~pi299 & ~n22152;
  assign n22154 = n3053 & ~n22144;
  assign n22155 = ~pi166 & ~n16787;
  assign n22156 = n21332 & ~n22155;
  assign n22157 = ~n22154 & ~n22156;
  assign n22158 = ~pi223 & ~n22157;
  assign n22159 = n22153 & ~n22158;
  assign n22160 = pi772 & ~n22159;
  assign n22161 = ~n22150 & n22160;
  assign n22162 = ~pi772 & ~n16814;
  assign n22163 = pi166 & n22162;
  assign n22164 = pi39 & ~n22163;
  assign n22165 = ~n22161 & n22164;
  assign n22166 = pi166 & ~n16655;
  assign n22167 = pi772 & pi947;
  assign n22168 = ~pi39 & ~n22167;
  assign n22169 = ~n16656 & ~n22168;
  assign n22170 = ~n22166 & ~n22169;
  assign n22171 = ~pi38 & ~n22170;
  assign n22172 = ~n22165 & n22171;
  assign n22173 = ~pi166 & ~n17485;
  assign n22174 = n16968 & ~n22167;
  assign n22175 = pi38 & ~n22174;
  assign n22176 = ~n22173 & n22175;
  assign n22177 = ~pi727 & ~n22176;
  assign n22178 = ~n22172 & n22177;
  assign n22179 = ~n21000 & ~n22143;
  assign n22180 = n3461 & n22179;
  assign n22181 = ~pi215 & ~n22180;
  assign n22182 = ~n16801 & n22140;
  assign n22183 = n22181 & ~n22182;
  assign n22184 = ~pi166 & ~n16805;
  assign n22185 = n20930 & ~n22184;
  assign n22186 = pi299 & ~n22185;
  assign n22187 = ~n22183 & n22186;
  assign n22188 = n3053 & n22179;
  assign n22189 = ~pi223 & ~n22188;
  assign n22190 = ~n21350 & ~n22155;
  assign n22191 = n21335 & ~n22190;
  assign n22192 = n22189 & ~n22191;
  assign n22193 = ~n6217 & n16728;
  assign n22194 = ~pi166 & ~n22193;
  assign n22195 = n20984 & ~n22194;
  assign n22196 = n22153 & ~n22195;
  assign n22197 = ~n22192 & n22196;
  assign n22198 = pi772 & ~n22197;
  assign n22199 = ~n22187 & n22198;
  assign n22200 = ~n3053 & ~n22190;
  assign n22201 = n3053 & n20957;
  assign n22202 = n22189 & ~n22201;
  assign n22203 = ~n22200 & n22202;
  assign n22204 = ~pi299 & ~n22195;
  assign n22205 = ~n22203 & n22204;
  assign n22206 = ~n20971 & n22181;
  assign n22207 = ~n22140 & n22206;
  assign n22208 = ~n21359 & n22185;
  assign n22209 = pi299 & ~n22208;
  assign n22210 = ~n22207 & n22209;
  assign n22211 = ~pi772 & ~n22205;
  assign n22212 = ~n22210 & n22211;
  assign n22213 = pi39 & ~n22199;
  assign n22214 = ~n22212 & n22213;
  assign n22215 = ~n21041 & n22170;
  assign n22216 = ~pi38 & ~n22215;
  assign n22217 = ~n22214 & n22216;
  assign n22218 = n21376 & n22168;
  assign n22219 = ~pi166 & ~n16968;
  assign n22220 = pi38 & ~n22218;
  assign n22221 = ~n22219 & n22220;
  assign n22222 = pi727 & ~n22221;
  assign n22223 = ~n22217 & n22222;
  assign n22224 = ~n22178 & ~n22223;
  assign n22225 = n10178 & ~n22224;
  assign n22226 = ~pi166 & ~n10178;
  assign n22227 = ~pi832 & ~n22226;
  assign n22228 = ~n22225 & n22227;
  assign n22229 = pi727 & n20848;
  assign n22230 = n2755 & ~n22167;
  assign n22231 = ~n22229 & n22230;
  assign n22232 = ~pi166 & ~n2755;
  assign n22233 = pi832 & ~n22232;
  assign n22234 = ~n22231 & n22233;
  assign po323 = n22228 | n22234;
  assign n22236 = ~pi768 & pi947;
  assign n22237 = pi705 & n20848;
  assign n22238 = ~n22236 & ~n22237;
  assign n22239 = n2755 & ~n22238;
  assign n22240 = ~pi167 & ~n2755;
  assign n22241 = pi832 & ~n22240;
  assign n22242 = ~n22239 & n22241;
  assign n22243 = ~pi167 & n21026;
  assign n22244 = pi167 & n21043;
  assign n22245 = ~pi38 & ~n22244;
  assign n22246 = ~n22243 & n22245;
  assign n22247 = ~pi167 & ~n16968;
  assign n22248 = n21049 & ~n22247;
  assign n22249 = pi768 & ~n22248;
  assign n22250 = ~n22246 & n22249;
  assign n22251 = ~pi167 & n20995;
  assign n22252 = pi167 & n21008;
  assign n22253 = ~pi38 & ~n22252;
  assign n22254 = ~n22251 & n22253;
  assign n22255 = ~pi167 & ~n21012;
  assign n22256 = n21015 & ~n22255;
  assign n22257 = ~pi768 & ~n22256;
  assign n22258 = ~n22254 & n22257;
  assign n22259 = pi705 & ~n22250;
  assign n22260 = ~n22258 & n22259;
  assign n22261 = ~pi167 & ~n20938;
  assign n22262 = pi167 & n20964;
  assign n22263 = ~pi38 & ~n22262;
  assign n22264 = ~n22261 & n22263;
  assign n22265 = ~pi167 & ~n17485;
  assign n22266 = ~n20947 & ~n22265;
  assign n22267 = ~pi768 & ~n22266;
  assign n22268 = ~n22264 & n22267;
  assign n22269 = pi768 & ~n17487;
  assign n22270 = ~pi167 & n22269;
  assign n22271 = ~pi705 & ~n22270;
  assign n22272 = ~n22268 & n22271;
  assign n22273 = n10178 & ~n22272;
  assign n22274 = ~n22260 & n22273;
  assign n22275 = ~pi167 & ~n10178;
  assign n22276 = ~pi832 & ~n22275;
  assign n22277 = ~n22274 & n22276;
  assign po324 = ~n22242 & ~n22277;
  assign n22279 = pi763 & pi947;
  assign n22280 = n2755 & ~n22279;
  assign n22281 = pi699 & n20848;
  assign n22282 = n22280 & ~n22281;
  assign n22283 = pi168 & ~n2755;
  assign n22284 = pi832 & ~n22283;
  assign n22285 = ~n22282 & n22284;
  assign n22286 = ~pi168 & ~n16655;
  assign n22287 = ~pi763 & n18015;
  assign n22288 = ~n20949 & ~n22287;
  assign n22289 = ~n22286 & ~n22288;
  assign n22290 = ~n21041 & n22289;
  assign n22291 = pi168 & ~n16805;
  assign n22292 = n20930 & ~n22291;
  assign n22293 = pi168 & ~n3461;
  assign n22294 = ~n16801 & n22293;
  assign n22295 = ~n16798 & ~n22294;
  assign n22296 = ~pi168 & ~n16661;
  assign n22297 = n20958 & ~n22296;
  assign n22298 = ~n21030 & n22297;
  assign n22299 = ~pi215 & ~n22298;
  assign n22300 = n22295 & n22299;
  assign n22301 = ~n22292 & ~n22300;
  assign n22302 = pi299 & ~n22301;
  assign n22303 = pi168 & ~n20997;
  assign n22304 = n20987 & ~n22303;
  assign n22305 = ~n22302 & ~n22304;
  assign n22306 = pi763 & ~n22305;
  assign n22307 = n21032 & ~n22296;
  assign n22308 = ~n20973 & ~n22307;
  assign n22309 = n22295 & n22308;
  assign n22310 = ~pi215 & ~n22309;
  assign n22311 = n20999 & ~n22292;
  assign n22312 = ~n20953 & ~n22311;
  assign n22313 = ~n22310 & n22312;
  assign n22314 = pi299 & ~n22313;
  assign n22315 = ~pi168 & ~n16792;
  assign n22316 = n21038 & ~n22315;
  assign n22317 = ~pi763 & ~n22316;
  assign n22318 = ~n22314 & n22317;
  assign n22319 = pi39 & ~n22318;
  assign n22320 = ~n22306 & n22319;
  assign n22321 = ~n22290 & ~n22320;
  assign n22322 = ~pi38 & ~n22321;
  assign n22323 = ~pi168 & ~n16968;
  assign n22324 = ~pi763 & pi947;
  assign n22325 = ~pi39 & ~n22324;
  assign n22326 = n21170 & n22325;
  assign n22327 = pi38 & ~n22323;
  assign n22328 = ~n22326 & n22327;
  assign n22329 = ~n22322 & ~n22328;
  assign n22330 = pi699 & ~n22329;
  assign n22331 = n20951 & ~n22315;
  assign n22332 = n22295 & ~n22297;
  assign n22333 = n20928 & n22332;
  assign n22334 = n20932 & ~n22291;
  assign n22335 = pi299 & ~n22334;
  assign n22336 = ~n22333 & n22335;
  assign n22337 = pi763 & ~n22336;
  assign n22338 = ~n22331 & n22337;
  assign n22339 = ~pi168 & ~pi763;
  assign n22340 = ~n16814 & n22339;
  assign n22341 = pi39 & ~n22340;
  assign n22342 = ~n22338 & n22341;
  assign n22343 = ~pi38 & ~n22289;
  assign n22344 = ~n22342 & n22343;
  assign n22345 = pi168 & ~n17485;
  assign n22346 = n6250 & n22280;
  assign n22347 = pi38 & ~n22346;
  assign n22348 = ~n22345 & n22347;
  assign n22349 = ~pi699 & ~n22348;
  assign n22350 = ~n22344 & n22349;
  assign n22351 = n21085 & ~n22350;
  assign n22352 = ~n22330 & n22351;
  assign n22353 = ~pi168 & ~n21085;
  assign n22354 = ~pi57 & ~n22353;
  assign n22355 = ~n22352 & n22354;
  assign n22356 = pi57 & pi168;
  assign n22357 = ~pi832 & ~n22356;
  assign n22358 = ~n22355 & n22357;
  assign po325 = n22285 | n22358;
  assign n22360 = pi746 & pi947;
  assign n22361 = n2755 & ~n22360;
  assign n22362 = pi729 & n20848;
  assign n22363 = n22361 & ~n22362;
  assign n22364 = pi169 & ~n2755;
  assign n22365 = pi832 & ~n22364;
  assign n22366 = ~n22363 & n22365;
  assign n22367 = ~pi169 & ~n16655;
  assign n22368 = ~pi746 & n18015;
  assign n22369 = ~n20949 & ~n22368;
  assign n22370 = ~n22367 & ~n22369;
  assign n22371 = ~n21041 & n22370;
  assign n22372 = pi169 & ~n16805;
  assign n22373 = n20930 & ~n22372;
  assign n22374 = pi169 & ~n3461;
  assign n22375 = ~n16801 & n22374;
  assign n22376 = ~n16798 & ~n22375;
  assign n22377 = ~pi169 & ~n16661;
  assign n22378 = n20958 & ~n22377;
  assign n22379 = ~n21030 & n22378;
  assign n22380 = ~pi215 & ~n22379;
  assign n22381 = n22376 & n22380;
  assign n22382 = ~n22373 & ~n22381;
  assign n22383 = pi299 & ~n22382;
  assign n22384 = pi169 & ~n20997;
  assign n22385 = n20987 & ~n22384;
  assign n22386 = ~n22383 & ~n22385;
  assign n22387 = pi746 & ~n22386;
  assign n22388 = n21032 & ~n22377;
  assign n22389 = ~n20973 & ~n22388;
  assign n22390 = n22376 & n22389;
  assign n22391 = ~pi215 & ~n22390;
  assign n22392 = n20999 & ~n22373;
  assign n22393 = ~n20953 & ~n22392;
  assign n22394 = ~n22391 & n22393;
  assign n22395 = pi299 & ~n22394;
  assign n22396 = ~pi169 & ~n16792;
  assign n22397 = n21038 & ~n22396;
  assign n22398 = ~pi746 & ~n22397;
  assign n22399 = ~n22395 & n22398;
  assign n22400 = pi39 & ~n22399;
  assign n22401 = ~n22387 & n22400;
  assign n22402 = ~n22371 & ~n22401;
  assign n22403 = ~pi38 & ~n22402;
  assign n22404 = ~pi169 & ~n16968;
  assign n22405 = ~pi746 & pi947;
  assign n22406 = ~pi39 & ~n22405;
  assign n22407 = n21170 & n22406;
  assign n22408 = pi38 & ~n22404;
  assign n22409 = ~n22407 & n22408;
  assign n22410 = ~n22403 & ~n22409;
  assign n22411 = pi729 & ~n22410;
  assign n22412 = n20951 & ~n22396;
  assign n22413 = n22376 & ~n22378;
  assign n22414 = n20928 & n22413;
  assign n22415 = n20932 & ~n22372;
  assign n22416 = pi299 & ~n22415;
  assign n22417 = ~n22414 & n22416;
  assign n22418 = pi746 & ~n22417;
  assign n22419 = ~n22412 & n22418;
  assign n22420 = ~pi169 & ~pi746;
  assign n22421 = ~n16814 & n22420;
  assign n22422 = pi39 & ~n22421;
  assign n22423 = ~n22419 & n22422;
  assign n22424 = ~pi38 & ~n22370;
  assign n22425 = ~n22423 & n22424;
  assign n22426 = pi169 & ~n17485;
  assign n22427 = n6250 & n22361;
  assign n22428 = pi38 & ~n22427;
  assign n22429 = ~n22426 & n22428;
  assign n22430 = ~pi729 & ~n22429;
  assign n22431 = ~n22425 & n22430;
  assign n22432 = n21085 & ~n22431;
  assign n22433 = ~n22411 & n22432;
  assign n22434 = ~pi169 & ~n21085;
  assign n22435 = ~pi57 & ~n22434;
  assign n22436 = ~n22433 & n22435;
  assign n22437 = pi57 & pi169;
  assign n22438 = ~pi832 & ~n22437;
  assign n22439 = ~n22436 & n22438;
  assign po326 = n22366 | n22439;
  assign n22441 = pi730 & n20848;
  assign n22442 = pi748 & pi947;
  assign n22443 = n2755 & ~n22442;
  assign n22444 = ~n22441 & n22443;
  assign n22445 = pi170 & ~n2755;
  assign n22446 = pi832 & ~n22445;
  assign n22447 = ~n22444 & n22446;
  assign n22448 = pi170 & ~n3461;
  assign n22449 = ~n16801 & n22448;
  assign n22450 = ~n16798 & ~n22449;
  assign n22451 = ~pi170 & ~n16661;
  assign n22452 = n21032 & ~n22451;
  assign n22453 = ~n20973 & ~n22452;
  assign n22454 = n22450 & n22453;
  assign n22455 = ~pi215 & ~n22454;
  assign n22456 = pi170 & ~n16805;
  assign n22457 = n20930 & ~n22456;
  assign n22458 = n20999 & ~n22457;
  assign n22459 = ~n20953 & ~n22458;
  assign n22460 = ~n22455 & n22459;
  assign n22461 = pi299 & ~n22460;
  assign n22462 = ~pi170 & ~n16792;
  assign n22463 = ~pi299 & ~n22462;
  assign n22464 = ~n21037 & n22463;
  assign n22465 = ~n22461 & ~n22464;
  assign n22466 = pi39 & ~n22465;
  assign n22467 = ~pi170 & ~n16655;
  assign n22468 = n21042 & ~n22467;
  assign n22469 = ~n22466 & ~n22468;
  assign n22470 = ~pi38 & ~n22469;
  assign n22471 = ~pi170 & ~n16968;
  assign n22472 = n21049 & ~n22471;
  assign n22473 = ~pi748 & ~n22472;
  assign n22474 = ~n22470 & n22473;
  assign n22475 = n20993 & ~n22467;
  assign n22476 = pi170 & ~n20997;
  assign n22477 = n20987 & ~n22476;
  assign n22478 = n20958 & ~n22451;
  assign n22479 = ~n21030 & n22478;
  assign n22480 = ~pi215 & ~n22479;
  assign n22481 = n22450 & n22480;
  assign n22482 = ~n22457 & ~n22481;
  assign n22483 = pi299 & ~n22482;
  assign n22484 = pi39 & ~n22483;
  assign n22485 = ~n22477 & n22484;
  assign n22486 = ~n22475 & ~n22485;
  assign n22487 = ~pi38 & ~n22486;
  assign n22488 = n21015 & ~n22471;
  assign n22489 = pi748 & ~n22488;
  assign n22490 = ~n22487 & n22489;
  assign n22491 = pi730 & ~n22490;
  assign n22492 = ~n22474 & n22491;
  assign n22493 = n20949 & ~n22467;
  assign n22494 = n22450 & ~n22478;
  assign n22495 = n20928 & n22494;
  assign n22496 = n20932 & ~n22456;
  assign n22497 = pi299 & ~n22496;
  assign n22498 = ~n22495 & n22497;
  assign n22499 = ~n20950 & n22463;
  assign n22500 = ~n22498 & ~n22499;
  assign n22501 = pi39 & ~n22500;
  assign n22502 = ~n22493 & ~n22501;
  assign n22503 = ~pi38 & ~n22502;
  assign n22504 = ~pi170 & ~n17485;
  assign n22505 = ~n20947 & ~n22504;
  assign n22506 = pi748 & ~n22505;
  assign n22507 = ~n22503 & n22506;
  assign n22508 = ~pi170 & ~pi748;
  assign n22509 = ~n17487 & n22508;
  assign n22510 = ~pi730 & ~n22509;
  assign n22511 = ~n22507 & n22510;
  assign n22512 = n21085 & ~n22511;
  assign n22513 = ~n22492 & n22512;
  assign n22514 = ~pi170 & ~n21085;
  assign n22515 = ~pi57 & ~n22514;
  assign n22516 = ~n22513 & n22515;
  assign n22517 = pi57 & pi170;
  assign n22518 = ~pi832 & ~n22517;
  assign n22519 = ~n22516 & n22518;
  assign po327 = n22447 | n22519;
  assign n22521 = pi764 & pi947;
  assign n22522 = n2755 & ~n22521;
  assign n22523 = pi691 & n20848;
  assign n22524 = n22522 & ~n22523;
  assign n22525 = pi171 & ~n2755;
  assign n22526 = pi832 & ~n22525;
  assign n22527 = ~n22524 & n22526;
  assign n22528 = ~pi171 & ~n16655;
  assign n22529 = ~pi764 & n18015;
  assign n22530 = ~n20949 & ~n22529;
  assign n22531 = ~n22528 & ~n22530;
  assign n22532 = ~n21041 & n22531;
  assign n22533 = pi171 & ~n16805;
  assign n22534 = n20930 & ~n22533;
  assign n22535 = pi171 & ~n3461;
  assign n22536 = ~n16801 & n22535;
  assign n22537 = ~n16798 & ~n22536;
  assign n22538 = ~pi171 & ~n16661;
  assign n22539 = n20958 & ~n22538;
  assign n22540 = ~n21030 & n22539;
  assign n22541 = ~pi215 & ~n22540;
  assign n22542 = n22537 & n22541;
  assign n22543 = ~n22534 & ~n22542;
  assign n22544 = pi299 & ~n22543;
  assign n22545 = pi171 & ~n20997;
  assign n22546 = n20987 & ~n22545;
  assign n22547 = ~n22544 & ~n22546;
  assign n22548 = pi764 & ~n22547;
  assign n22549 = n21032 & ~n22538;
  assign n22550 = ~n20973 & ~n22549;
  assign n22551 = n22537 & n22550;
  assign n22552 = ~pi215 & ~n22551;
  assign n22553 = n20999 & ~n22534;
  assign n22554 = ~n20953 & ~n22553;
  assign n22555 = ~n22552 & n22554;
  assign n22556 = pi299 & ~n22555;
  assign n22557 = ~pi171 & ~n16792;
  assign n22558 = n21038 & ~n22557;
  assign n22559 = ~pi764 & ~n22558;
  assign n22560 = ~n22556 & n22559;
  assign n22561 = pi39 & ~n22560;
  assign n22562 = ~n22548 & n22561;
  assign n22563 = ~n22532 & ~n22562;
  assign n22564 = ~pi38 & ~n22563;
  assign n22565 = ~pi171 & ~n16968;
  assign n22566 = ~pi764 & pi947;
  assign n22567 = ~pi39 & ~n22566;
  assign n22568 = n21170 & n22567;
  assign n22569 = pi38 & ~n22565;
  assign n22570 = ~n22568 & n22569;
  assign n22571 = ~n22564 & ~n22570;
  assign n22572 = pi691 & ~n22571;
  assign n22573 = n20951 & ~n22557;
  assign n22574 = n22537 & ~n22539;
  assign n22575 = n20928 & n22574;
  assign n22576 = n20932 & ~n22533;
  assign n22577 = pi299 & ~n22576;
  assign n22578 = ~n22575 & n22577;
  assign n22579 = pi764 & ~n22578;
  assign n22580 = ~n22573 & n22579;
  assign n22581 = ~pi171 & ~pi764;
  assign n22582 = ~n16814 & n22581;
  assign n22583 = pi39 & ~n22582;
  assign n22584 = ~n22580 & n22583;
  assign n22585 = ~pi38 & ~n22531;
  assign n22586 = ~n22584 & n22585;
  assign n22587 = pi171 & ~n17485;
  assign n22588 = n6250 & n22522;
  assign n22589 = pi38 & ~n22588;
  assign n22590 = ~n22587 & n22589;
  assign n22591 = ~pi691 & ~n22590;
  assign n22592 = ~n22586 & n22591;
  assign n22593 = n21085 & ~n22592;
  assign n22594 = ~n22572 & n22593;
  assign n22595 = ~pi171 & ~n21085;
  assign n22596 = ~pi57 & ~n22595;
  assign n22597 = ~n22594 & n22596;
  assign n22598 = pi57 & pi171;
  assign n22599 = ~pi832 & ~n22598;
  assign n22600 = ~n22597 & n22599;
  assign po328 = n22527 | n22600;
  assign n22602 = pi739 & pi947;
  assign n22603 = n2755 & ~n22602;
  assign n22604 = pi690 & n20848;
  assign n22605 = n22603 & ~n22604;
  assign n22606 = pi172 & ~n2755;
  assign n22607 = pi832 & ~n22606;
  assign n22608 = ~n22605 & n22607;
  assign n22609 = ~pi172 & ~n16655;
  assign n22610 = n16655 & n22602;
  assign n22611 = ~pi39 & ~n22609;
  assign n22612 = ~n22610 & n22611;
  assign n22613 = ~n21041 & n22612;
  assign n22614 = pi172 & ~n16805;
  assign n22615 = n20930 & ~n22614;
  assign n22616 = pi172 & ~n3461;
  assign n22617 = ~n16801 & n22616;
  assign n22618 = ~n16798 & ~n22617;
  assign n22619 = ~pi172 & ~n16661;
  assign n22620 = n20958 & ~n22619;
  assign n22621 = ~n21030 & n22620;
  assign n22622 = ~pi215 & ~n22621;
  assign n22623 = n22618 & n22622;
  assign n22624 = ~n22615 & ~n22623;
  assign n22625 = pi299 & ~n22624;
  assign n22626 = pi172 & ~n20997;
  assign n22627 = n20987 & ~n22626;
  assign n22628 = ~n22625 & ~n22627;
  assign n22629 = pi739 & ~n22628;
  assign n22630 = n21032 & ~n22619;
  assign n22631 = ~n20973 & ~n22630;
  assign n22632 = n22618 & n22631;
  assign n22633 = ~pi215 & ~n22632;
  assign n22634 = n20999 & ~n22615;
  assign n22635 = ~n20953 & ~n22634;
  assign n22636 = ~n22633 & n22635;
  assign n22637 = pi299 & ~n22636;
  assign n22638 = ~pi172 & ~n16792;
  assign n22639 = n21038 & ~n22638;
  assign n22640 = ~pi739 & ~n22639;
  assign n22641 = ~n22637 & n22640;
  assign n22642 = pi39 & ~n22641;
  assign n22643 = ~n22629 & n22642;
  assign n22644 = ~n22613 & ~n22643;
  assign n22645 = ~pi38 & ~n22644;
  assign n22646 = ~pi172 & ~n16968;
  assign n22647 = ~pi739 & pi947;
  assign n22648 = ~pi39 & ~n22647;
  assign n22649 = n21170 & n22648;
  assign n22650 = pi38 & ~n22646;
  assign n22651 = ~n22649 & n22650;
  assign n22652 = ~n22645 & ~n22651;
  assign n22653 = pi690 & ~n22652;
  assign n22654 = n20951 & ~n22638;
  assign n22655 = n22618 & ~n22620;
  assign n22656 = n20928 & n22655;
  assign n22657 = n20932 & ~n22614;
  assign n22658 = pi299 & ~n22657;
  assign n22659 = ~n22656 & n22658;
  assign n22660 = pi739 & ~n22659;
  assign n22661 = ~n22654 & n22660;
  assign n22662 = ~pi172 & ~pi739;
  assign n22663 = ~n16814 & n22662;
  assign n22664 = pi39 & ~n22663;
  assign n22665 = ~n22661 & n22664;
  assign n22666 = ~pi38 & ~n22612;
  assign n22667 = ~n22665 & n22666;
  assign n22668 = pi172 & ~n17485;
  assign n22669 = n6250 & n22603;
  assign n22670 = pi38 & ~n22669;
  assign n22671 = ~n22668 & n22670;
  assign n22672 = ~pi690 & ~n22671;
  assign n22673 = ~n22667 & n22672;
  assign n22674 = n21085 & ~n22673;
  assign n22675 = ~n22653 & n22674;
  assign n22676 = ~pi172 & ~n21085;
  assign n22677 = ~pi57 & ~n22676;
  assign n22678 = ~n22675 & n22677;
  assign n22679 = pi57 & pi172;
  assign n22680 = ~pi832 & ~n22679;
  assign n22681 = ~n22678 & n22680;
  assign po329 = n22608 | n22681;
  assign n22683 = ~pi173 & ~n17494;
  assign n22684 = n17627 & ~n22683;
  assign n22685 = ~pi723 & n3268;
  assign n22686 = n22683 & ~n22685;
  assign n22687 = pi173 & ~n18064;
  assign n22688 = ~pi38 & ~n22687;
  assign n22689 = n3268 & ~n22688;
  assign n22690 = ~pi173 & n18060;
  assign n22691 = ~n22689 & ~n22690;
  assign n22692 = ~pi173 & ~n16968;
  assign n22693 = n17480 & ~n22692;
  assign n22694 = ~pi723 & ~n22693;
  assign n22695 = ~n22691 & n22694;
  assign n22696 = ~n22686 & ~n22695;
  assign n22697 = ~pi778 & n22696;
  assign n22698 = pi625 & ~n22696;
  assign n22699 = ~pi625 & n22683;
  assign n22700 = pi1153 & ~n22699;
  assign n22701 = ~n22698 & n22700;
  assign n22702 = ~pi625 & ~n22696;
  assign n22703 = pi625 & n22683;
  assign n22704 = ~pi1153 & ~n22703;
  assign n22705 = ~n22702 & n22704;
  assign n22706 = ~n22701 & ~n22705;
  assign n22707 = pi778 & ~n22706;
  assign n22708 = ~n22697 & ~n22707;
  assign n22709 = ~n17554 & ~n22708;
  assign n22710 = n17554 & ~n22683;
  assign n22711 = ~n22709 & ~n22710;
  assign n22712 = ~n17591 & n22711;
  assign n22713 = n17591 & n22683;
  assign n22714 = ~n22712 & ~n22713;
  assign n22715 = ~n17627 & n22714;
  assign n22716 = ~n22684 & ~n22715;
  assign n22717 = ~n17670 & n22716;
  assign n22718 = n17670 & n22683;
  assign n22719 = ~n22717 & ~n22718;
  assign n22720 = ~pi792 & n22719;
  assign n22721 = pi628 & ~n22719;
  assign n22722 = ~pi628 & n22683;
  assign n22723 = pi1156 & ~n22722;
  assign n22724 = ~n22721 & n22723;
  assign n22725 = ~pi628 & ~n22719;
  assign n22726 = pi628 & n22683;
  assign n22727 = ~pi1156 & ~n22726;
  assign n22728 = ~n22725 & n22727;
  assign n22729 = ~n22724 & ~n22728;
  assign n22730 = pi792 & ~n22729;
  assign n22731 = ~n22720 & ~n22730;
  assign n22732 = ~pi647 & ~n22731;
  assign n22733 = pi647 & ~n22683;
  assign n22734 = ~n22732 & ~n22733;
  assign n22735 = ~pi1157 & n22734;
  assign n22736 = pi647 & ~n22731;
  assign n22737 = ~pi647 & ~n22683;
  assign n22738 = ~n22736 & ~n22737;
  assign n22739 = pi1157 & n22738;
  assign n22740 = ~n22735 & ~n22739;
  assign n22741 = pi787 & ~n22740;
  assign n22742 = ~pi787 & n22731;
  assign n22743 = ~n22741 & ~n22742;
  assign n22744 = ~pi644 & ~n22743;
  assign n22745 = pi715 & ~n22744;
  assign n22746 = pi173 & ~n3268;
  assign n22747 = ~pi173 & ~n16816;
  assign n22748 = pi745 & ~n22747;
  assign n22749 = pi173 & ~n16963;
  assign n22750 = ~pi173 & ~pi745;
  assign n22751 = n16907 & n22750;
  assign n22752 = ~n22749 & ~n22751;
  assign n22753 = ~n22748 & n22752;
  assign n22754 = ~pi38 & ~n22753;
  assign n22755 = ~pi745 & n16970;
  assign n22756 = pi38 & ~n22692;
  assign n22757 = ~n22755 & n22756;
  assign n22758 = ~n22754 & ~n22757;
  assign n22759 = n3268 & ~n22758;
  assign n22760 = ~n22746 & ~n22759;
  assign n22761 = ~n17526 & ~n22760;
  assign n22762 = n17526 & ~n22683;
  assign n22763 = ~n22761 & ~n22762;
  assign n22764 = ~pi785 & ~n22763;
  assign n22765 = ~n17527 & ~n22683;
  assign n22766 = pi609 & n22761;
  assign n22767 = ~n22765 & ~n22766;
  assign n22768 = pi1155 & ~n22767;
  assign n22769 = ~n17539 & ~n22683;
  assign n22770 = ~pi609 & n22761;
  assign n22771 = ~n22769 & ~n22770;
  assign n22772 = ~pi1155 & ~n22771;
  assign n22773 = ~n22768 & ~n22772;
  assign n22774 = pi785 & ~n22773;
  assign n22775 = ~n22764 & ~n22774;
  assign n22776 = ~pi781 & ~n22775;
  assign n22777 = pi618 & n22775;
  assign n22778 = ~pi618 & n22683;
  assign n22779 = pi1154 & ~n22778;
  assign n22780 = ~n22777 & n22779;
  assign n22781 = ~pi618 & n22775;
  assign n22782 = pi618 & n22683;
  assign n22783 = ~pi1154 & ~n22782;
  assign n22784 = ~n22781 & n22783;
  assign n22785 = ~n22780 & ~n22784;
  assign n22786 = pi781 & ~n22785;
  assign n22787 = ~n22776 & ~n22786;
  assign n22788 = ~pi789 & ~n22787;
  assign n22789 = pi619 & n22787;
  assign n22790 = ~pi619 & n22683;
  assign n22791 = pi1159 & ~n22790;
  assign n22792 = ~n22789 & n22791;
  assign n22793 = ~pi619 & n22787;
  assign n22794 = pi619 & n22683;
  assign n22795 = ~pi1159 & ~n22794;
  assign n22796 = ~n22793 & n22795;
  assign n22797 = ~n22792 & ~n22796;
  assign n22798 = pi789 & ~n22797;
  assign n22799 = ~n22788 & ~n22798;
  assign n22800 = ~pi788 & ~n22799;
  assign n22801 = pi626 & n22799;
  assign n22802 = ~pi626 & n22683;
  assign n22803 = pi1158 & ~n22802;
  assign n22804 = ~n22801 & n22803;
  assign n22805 = ~pi626 & n22799;
  assign n22806 = pi626 & n22683;
  assign n22807 = ~pi1158 & ~n22806;
  assign n22808 = ~n22805 & n22807;
  assign n22809 = ~n22804 & ~n22808;
  assign n22810 = pi788 & ~n22809;
  assign n22811 = ~n22800 & ~n22810;
  assign n22812 = ~n17698 & n22811;
  assign n22813 = n17698 & n22683;
  assign n22814 = ~n22812 & ~n22813;
  assign n22815 = ~n17740 & ~n22814;
  assign n22816 = n17740 & n22683;
  assign n22817 = ~n22815 & ~n22816;
  assign n22818 = pi644 & ~n22817;
  assign n22819 = ~pi644 & n22683;
  assign n22820 = ~pi715 & ~n22819;
  assign n22821 = ~n22818 & n22820;
  assign n22822 = pi1160 & ~n22821;
  assign n22823 = ~n22745 & n22822;
  assign n22824 = ~n20491 & n22814;
  assign n22825 = n17738 & ~n22734;
  assign n22826 = n17737 & ~n22738;
  assign n22827 = ~n22825 & ~n22826;
  assign n22828 = ~n22824 & n22827;
  assign n22829 = pi787 & ~n22828;
  assign n22830 = ~n20502 & ~n22811;
  assign n22831 = ~pi629 & n22724;
  assign n22832 = pi629 & n22728;
  assign n22833 = ~n22831 & ~n22832;
  assign n22834 = ~n22830 & n22833;
  assign n22835 = pi792 & ~n22834;
  assign n22836 = pi723 & n22758;
  assign n22837 = ~pi173 & n17074;
  assign n22838 = pi173 & n17166;
  assign n22839 = pi745 & ~n22838;
  assign n22840 = ~n22837 & n22839;
  assign n22841 = pi173 & n17233;
  assign n22842 = ~pi173 & ~n17295;
  assign n22843 = ~pi745 & ~n22842;
  assign n22844 = ~n22841 & n22843;
  assign n22845 = pi39 & ~n22844;
  assign n22846 = ~n22840 & n22845;
  assign n22847 = pi173 & ~n17340;
  assign n22848 = ~pi173 & ~n17317;
  assign n22849 = pi745 & ~n22847;
  assign n22850 = ~n22848 & n22849;
  assign n22851 = ~pi173 & n17344;
  assign n22852 = pi173 & n17351;
  assign n22853 = ~pi745 & ~n22852;
  assign n22854 = ~n22851 & n22853;
  assign n22855 = ~n22850 & ~n22854;
  assign n22856 = ~pi39 & ~n22855;
  assign n22857 = ~pi38 & ~n22856;
  assign n22858 = ~n22846 & n22857;
  assign n22859 = ~pi745 & ~n17259;
  assign n22860 = n19303 & ~n22859;
  assign n22861 = ~pi173 & ~n22860;
  assign n22862 = ~pi745 & n16933;
  assign n22863 = ~n17154 & ~n22862;
  assign n22864 = pi173 & ~n22863;
  assign n22865 = n6250 & n22864;
  assign n22866 = pi38 & ~n22865;
  assign n22867 = ~n22861 & n22866;
  assign n22868 = ~pi723 & ~n22867;
  assign n22869 = ~n22858 & n22868;
  assign n22870 = n3268 & ~n22869;
  assign n22871 = ~n22836 & n22870;
  assign n22872 = ~n22746 & ~n22871;
  assign n22873 = ~pi625 & n22872;
  assign n22874 = pi625 & n22760;
  assign n22875 = ~pi1153 & ~n22874;
  assign n22876 = ~n22873 & n22875;
  assign n22877 = ~pi608 & ~n22701;
  assign n22878 = ~n22876 & n22877;
  assign n22879 = pi625 & n22872;
  assign n22880 = ~pi625 & n22760;
  assign n22881 = pi1153 & ~n22880;
  assign n22882 = ~n22879 & n22881;
  assign n22883 = pi608 & ~n22705;
  assign n22884 = ~n22882 & n22883;
  assign n22885 = ~n22878 & ~n22884;
  assign n22886 = pi778 & ~n22885;
  assign n22887 = ~pi778 & n22872;
  assign n22888 = ~n22886 & ~n22887;
  assign n22889 = ~pi609 & ~n22888;
  assign n22890 = pi609 & n22708;
  assign n22891 = ~pi1155 & ~n22890;
  assign n22892 = ~n22889 & n22891;
  assign n22893 = ~pi660 & ~n22768;
  assign n22894 = ~n22892 & n22893;
  assign n22895 = pi609 & ~n22888;
  assign n22896 = ~pi609 & n22708;
  assign n22897 = pi1155 & ~n22896;
  assign n22898 = ~n22895 & n22897;
  assign n22899 = pi660 & ~n22772;
  assign n22900 = ~n22898 & n22899;
  assign n22901 = ~n22894 & ~n22900;
  assign n22902 = pi785 & ~n22901;
  assign n22903 = ~pi785 & ~n22888;
  assign n22904 = ~n22902 & ~n22903;
  assign n22905 = ~pi618 & ~n22904;
  assign n22906 = pi618 & n22711;
  assign n22907 = ~pi1154 & ~n22906;
  assign n22908 = ~n22905 & n22907;
  assign n22909 = ~pi627 & ~n22780;
  assign n22910 = ~n22908 & n22909;
  assign n22911 = pi618 & ~n22904;
  assign n22912 = ~pi618 & n22711;
  assign n22913 = pi1154 & ~n22912;
  assign n22914 = ~n22911 & n22913;
  assign n22915 = pi627 & ~n22784;
  assign n22916 = ~n22914 & n22915;
  assign n22917 = ~n22910 & ~n22916;
  assign n22918 = pi781 & ~n22917;
  assign n22919 = ~pi781 & ~n22904;
  assign n22920 = ~n22918 & ~n22919;
  assign n22921 = ~pi619 & ~n22920;
  assign n22922 = pi619 & ~n22714;
  assign n22923 = ~pi1159 & ~n22922;
  assign n22924 = ~n22921 & n22923;
  assign n22925 = ~pi648 & ~n22792;
  assign n22926 = ~n22924 & n22925;
  assign n22927 = pi619 & ~n22920;
  assign n22928 = ~pi619 & ~n22714;
  assign n22929 = pi1159 & ~n22928;
  assign n22930 = ~n22927 & n22929;
  assign n22931 = pi648 & ~n22796;
  assign n22932 = ~n22930 & n22931;
  assign n22933 = pi789 & ~n22926;
  assign n22934 = ~n22932 & n22933;
  assign n22935 = ~pi789 & n22920;
  assign n22936 = n17905 & ~n22935;
  assign n22937 = ~n22934 & n22936;
  assign n22938 = n17792 & n22716;
  assign n22939 = ~n17669 & n22809;
  assign n22940 = ~n22938 & ~n22939;
  assign n22941 = pi788 & ~n22940;
  assign n22942 = ~n20298 & ~n22941;
  assign n22943 = ~n22937 & n22942;
  assign n22944 = ~n22835 & ~n22943;
  assign n22945 = n20300 & ~n22944;
  assign n22946 = ~n22829 & ~n22945;
  assign n22947 = ~pi644 & n22946;
  assign n22948 = pi644 & ~n22743;
  assign n22949 = ~pi715 & ~n22948;
  assign n22950 = ~n22947 & n22949;
  assign n22951 = ~pi644 & ~n22817;
  assign n22952 = pi644 & n22683;
  assign n22953 = pi715 & ~n22952;
  assign n22954 = ~n22951 & n22953;
  assign n22955 = ~pi1160 & ~n22954;
  assign n22956 = ~n22950 & n22955;
  assign n22957 = ~n22823 & ~n22956;
  assign n22958 = pi790 & ~n22957;
  assign n22959 = pi644 & n22822;
  assign n22960 = pi790 & ~n22959;
  assign n22961 = n22946 & ~n22960;
  assign n22962 = ~n22958 & ~n22961;
  assign n22963 = ~po1038 & ~n22962;
  assign n22964 = ~pi173 & po1038;
  assign n22965 = ~pi832 & ~n22964;
  assign n22966 = ~n22963 & n22965;
  assign n22967 = ~pi173 & ~n2755;
  assign n22968 = ~n22862 & ~n22967;
  assign n22969 = ~n17794 & ~n22968;
  assign n22970 = ~pi785 & ~n22969;
  assign n22971 = n17539 & n22862;
  assign n22972 = n22969 & ~n22971;
  assign n22973 = pi1155 & ~n22972;
  assign n22974 = ~pi1155 & ~n22967;
  assign n22975 = ~n22971 & n22974;
  assign n22976 = ~n22973 & ~n22975;
  assign n22977 = pi785 & ~n22976;
  assign n22978 = ~n22970 & ~n22977;
  assign n22979 = ~pi781 & ~n22978;
  assign n22980 = ~n17809 & n22978;
  assign n22981 = pi1154 & ~n22980;
  assign n22982 = ~n17812 & n22978;
  assign n22983 = ~pi1154 & ~n22982;
  assign n22984 = ~n22981 & ~n22983;
  assign n22985 = pi781 & ~n22984;
  assign n22986 = ~n22979 & ~n22985;
  assign n22987 = ~pi789 & ~n22986;
  assign n22988 = ~pi619 & n2755;
  assign n22989 = n22986 & ~n22988;
  assign n22990 = pi1159 & ~n22989;
  assign n22991 = pi619 & n2755;
  assign n22992 = n22986 & ~n22991;
  assign n22993 = ~pi1159 & ~n22992;
  assign n22994 = ~n22990 & ~n22993;
  assign n22995 = pi789 & ~n22994;
  assign n22996 = ~n22987 & ~n22995;
  assign n22997 = ~pi788 & ~n22996;
  assign n22998 = pi626 & n22996;
  assign n22999 = ~pi626 & n22967;
  assign n23000 = pi1158 & ~n22999;
  assign n23001 = ~n22998 & n23000;
  assign n23002 = ~pi626 & n22996;
  assign n23003 = pi626 & n22967;
  assign n23004 = ~pi1158 & ~n23003;
  assign n23005 = ~n23002 & n23004;
  assign n23006 = ~n23001 & ~n23005;
  assign n23007 = pi788 & ~n23006;
  assign n23008 = ~n22997 & ~n23007;
  assign n23009 = ~n17698 & n23008;
  assign n23010 = n17698 & n22967;
  assign n23011 = ~n23009 & ~n23010;
  assign n23012 = ~n20491 & n23011;
  assign n23013 = ~pi723 & n17153;
  assign n23014 = ~n22967 & ~n23013;
  assign n23015 = ~pi778 & ~n23014;
  assign n23016 = ~pi625 & n23013;
  assign n23017 = ~n23014 & ~n23016;
  assign n23018 = pi1153 & ~n23017;
  assign n23019 = ~pi1153 & ~n22967;
  assign n23020 = ~n23016 & n23019;
  assign n23021 = pi778 & ~n23020;
  assign n23022 = ~n23018 & n23021;
  assign n23023 = ~n23015 & ~n23022;
  assign n23024 = ~n17780 & ~n23023;
  assign n23025 = ~n17782 & n23024;
  assign n23026 = ~n17784 & n23025;
  assign n23027 = ~n17916 & n23026;
  assign n23028 = ~n17947 & n23027;
  assign n23029 = ~pi647 & n23028;
  assign n23030 = pi647 & n22967;
  assign n23031 = ~pi1157 & ~n23030;
  assign n23032 = ~n23029 & n23031;
  assign n23033 = pi647 & ~n23028;
  assign n23034 = ~pi647 & ~n22967;
  assign n23035 = ~n23033 & ~n23034;
  assign n23036 = pi1157 & ~n23035;
  assign n23037 = ~n23032 & ~n23036;
  assign n23038 = ~n17739 & ~n23037;
  assign n23039 = ~n23012 & ~n23038;
  assign n23040 = pi787 & ~n23039;
  assign n23041 = n17792 & n23026;
  assign n23042 = ~n17669 & n23006;
  assign n23043 = ~n23041 & ~n23042;
  assign n23044 = pi788 & ~n23043;
  assign n23045 = ~n16842 & ~n23014;
  assign n23046 = pi625 & n23045;
  assign n23047 = n22968 & ~n23045;
  assign n23048 = ~n23046 & ~n23047;
  assign n23049 = n23019 & ~n23048;
  assign n23050 = ~pi608 & ~n23018;
  assign n23051 = ~n23049 & n23050;
  assign n23052 = pi1153 & n22968;
  assign n23053 = ~n23046 & n23052;
  assign n23054 = pi608 & ~n23020;
  assign n23055 = ~n23053 & n23054;
  assign n23056 = ~n23051 & ~n23055;
  assign n23057 = pi778 & ~n23056;
  assign n23058 = ~pi778 & ~n23047;
  assign n23059 = ~n23057 & ~n23058;
  assign n23060 = ~pi609 & ~n23059;
  assign n23061 = pi609 & ~n23023;
  assign n23062 = ~pi1155 & ~n23061;
  assign n23063 = ~n23060 & n23062;
  assign n23064 = ~pi660 & ~n22973;
  assign n23065 = ~n23063 & n23064;
  assign n23066 = pi609 & ~n23059;
  assign n23067 = ~pi609 & ~n23023;
  assign n23068 = pi1155 & ~n23067;
  assign n23069 = ~n23066 & n23068;
  assign n23070 = pi660 & ~n22975;
  assign n23071 = ~n23069 & n23070;
  assign n23072 = ~n23065 & ~n23071;
  assign n23073 = pi785 & ~n23072;
  assign n23074 = ~pi785 & ~n23059;
  assign n23075 = ~n23073 & ~n23074;
  assign n23076 = ~pi618 & ~n23075;
  assign n23077 = pi618 & n23024;
  assign n23078 = ~pi1154 & ~n23077;
  assign n23079 = ~n23076 & n23078;
  assign n23080 = ~pi627 & ~n22981;
  assign n23081 = ~n23079 & n23080;
  assign n23082 = pi618 & ~n23075;
  assign n23083 = ~pi618 & n23024;
  assign n23084 = pi1154 & ~n23083;
  assign n23085 = ~n23082 & n23084;
  assign n23086 = pi627 & ~n22983;
  assign n23087 = ~n23085 & n23086;
  assign n23088 = ~n23081 & ~n23087;
  assign n23089 = pi781 & ~n23088;
  assign n23090 = ~pi781 & ~n23075;
  assign n23091 = ~n23089 & ~n23090;
  assign n23092 = ~pi619 & ~n23091;
  assign n23093 = pi619 & n23025;
  assign n23094 = ~pi1159 & ~n23093;
  assign n23095 = ~n23092 & n23094;
  assign n23096 = ~pi648 & ~n22990;
  assign n23097 = ~n23095 & n23096;
  assign n23098 = pi619 & ~n23091;
  assign n23099 = ~pi619 & n23025;
  assign n23100 = pi1159 & ~n23099;
  assign n23101 = ~n23098 & n23100;
  assign n23102 = pi648 & ~n22993;
  assign n23103 = ~n23101 & n23102;
  assign n23104 = pi789 & ~n23097;
  assign n23105 = ~n23103 & n23104;
  assign n23106 = ~pi789 & n23091;
  assign n23107 = n17905 & ~n23106;
  assign n23108 = ~n23105 & n23107;
  assign n23109 = ~n23044 & ~n23108;
  assign n23110 = ~n20298 & ~n23109;
  assign n23111 = n17944 & n23008;
  assign n23112 = n20786 & n23027;
  assign n23113 = ~n23111 & ~n23112;
  assign n23114 = ~pi629 & ~n23113;
  assign n23115 = n20790 & n23027;
  assign n23116 = n17943 & n23008;
  assign n23117 = ~n23115 & ~n23116;
  assign n23118 = pi629 & ~n23117;
  assign n23119 = ~n23114 & ~n23118;
  assign n23120 = pi792 & ~n23119;
  assign n23121 = n20300 & ~n23120;
  assign n23122 = ~n23110 & n23121;
  assign n23123 = ~n23040 & ~n23122;
  assign n23124 = pi644 & n23123;
  assign n23125 = ~pi787 & ~n23028;
  assign n23126 = pi787 & ~n23037;
  assign n23127 = ~n23125 & ~n23126;
  assign n23128 = ~pi644 & n23127;
  assign n23129 = pi715 & ~n23128;
  assign n23130 = ~n23124 & n23129;
  assign n23131 = ~n17740 & ~n23011;
  assign n23132 = n17740 & n22967;
  assign n23133 = ~n23131 & ~n23132;
  assign n23134 = pi644 & ~n23133;
  assign n23135 = ~pi644 & n22967;
  assign n23136 = ~pi715 & ~n23135;
  assign n23137 = ~n23134 & n23136;
  assign n23138 = pi1160 & ~n23137;
  assign n23139 = ~n23130 & n23138;
  assign n23140 = ~pi644 & n23123;
  assign n23141 = pi644 & n23127;
  assign n23142 = ~pi715 & ~n23141;
  assign n23143 = ~n23140 & n23142;
  assign n23144 = ~pi644 & ~n23133;
  assign n23145 = pi644 & n22967;
  assign n23146 = pi715 & ~n23145;
  assign n23147 = ~n23144 & n23146;
  assign n23148 = ~pi1160 & ~n23147;
  assign n23149 = ~n23143 & n23148;
  assign n23150 = ~n23139 & ~n23149;
  assign n23151 = pi790 & ~n23150;
  assign n23152 = ~pi790 & n23123;
  assign n23153 = pi832 & ~n23152;
  assign n23154 = ~n23151 & n23153;
  assign po330 = ~n22966 & ~n23154;
  assign n23156 = pi174 & ~n3268;
  assign n23157 = pi759 & n16905;
  assign n23158 = ~n21397 & ~n23157;
  assign n23159 = pi39 & ~n23158;
  assign n23160 = pi759 & n16839;
  assign n23161 = ~pi759 & n16655;
  assign n23162 = ~pi39 & ~n23161;
  assign n23163 = ~n23160 & n23162;
  assign n23164 = ~n23159 & ~n23163;
  assign n23165 = pi174 & ~n23164;
  assign n23166 = ~pi174 & pi759;
  assign n23167 = n16963 & n23166;
  assign n23168 = ~n23165 & ~n23167;
  assign n23169 = ~pi38 & ~n23168;
  assign n23170 = ~pi174 & ~n16968;
  assign n23171 = pi759 & n16842;
  assign n23172 = n16968 & ~n23171;
  assign n23173 = pi38 & ~n23170;
  assign n23174 = ~n23172 & n23173;
  assign n23175 = ~n23169 & ~n23174;
  assign n23176 = ~pi696 & n23175;
  assign n23177 = pi174 & ~n17074;
  assign n23178 = ~pi174 & ~n17166;
  assign n23179 = ~pi759 & ~n23178;
  assign n23180 = ~n23177 & n23179;
  assign n23181 = ~pi174 & ~n17233;
  assign n23182 = pi174 & n17295;
  assign n23183 = pi759 & ~n23182;
  assign n23184 = ~n23181 & n23183;
  assign n23185 = pi39 & ~n23184;
  assign n23186 = ~n23180 & n23185;
  assign n23187 = ~pi174 & ~n17340;
  assign n23188 = pi174 & ~n17317;
  assign n23189 = ~pi759 & ~n23187;
  assign n23190 = ~n23188 & n23189;
  assign n23191 = pi174 & n17344;
  assign n23192 = ~pi174 & n17351;
  assign n23193 = pi759 & ~n23192;
  assign n23194 = ~n23191 & n23193;
  assign n23195 = ~pi39 & ~n23194;
  assign n23196 = ~n23190 & n23195;
  assign n23197 = ~pi38 & ~n23196;
  assign n23198 = ~n23186 & n23197;
  assign n23199 = pi696 & ~n19316;
  assign n23200 = ~n23174 & n23199;
  assign n23201 = ~n23198 & n23200;
  assign n23202 = n3268 & ~n23201;
  assign n23203 = ~n23176 & n23202;
  assign n23204 = ~n23156 & ~n23203;
  assign n23205 = ~pi625 & n23204;
  assign n23206 = n3268 & ~n23175;
  assign n23207 = ~n23156 & ~n23206;
  assign n23208 = pi625 & n23207;
  assign n23209 = ~pi1153 & ~n23208;
  assign n23210 = ~n23205 & n23209;
  assign n23211 = pi174 & ~n17494;
  assign n23212 = pi696 & n3268;
  assign n23213 = ~n23211 & ~n23212;
  assign n23214 = pi174 & ~n18060;
  assign n23215 = ~pi174 & n18064;
  assign n23216 = ~pi38 & ~n23215;
  assign n23217 = ~n23214 & n23216;
  assign n23218 = n19892 & ~n23170;
  assign n23219 = n23212 & ~n23218;
  assign n23220 = ~n23217 & n23219;
  assign n23221 = ~n23213 & ~n23220;
  assign n23222 = pi625 & ~n23221;
  assign n23223 = ~pi625 & ~n23211;
  assign n23224 = pi1153 & ~n23223;
  assign n23225 = ~n23222 & n23224;
  assign n23226 = ~pi608 & ~n23225;
  assign n23227 = ~n23210 & n23226;
  assign n23228 = pi625 & n23204;
  assign n23229 = ~pi625 & n23207;
  assign n23230 = pi1153 & ~n23229;
  assign n23231 = ~n23228 & n23230;
  assign n23232 = ~pi625 & ~n23221;
  assign n23233 = pi625 & ~n23211;
  assign n23234 = ~pi1153 & ~n23233;
  assign n23235 = ~n23232 & n23234;
  assign n23236 = pi608 & ~n23235;
  assign n23237 = ~n23231 & n23236;
  assign n23238 = ~n23227 & ~n23237;
  assign n23239 = pi778 & ~n23238;
  assign n23240 = ~pi778 & n23204;
  assign n23241 = ~n23239 & ~n23240;
  assign n23242 = ~pi609 & ~n23241;
  assign n23243 = ~pi778 & n23221;
  assign n23244 = ~n23225 & ~n23235;
  assign n23245 = pi778 & ~n23244;
  assign n23246 = ~n23243 & ~n23245;
  assign n23247 = pi609 & n23246;
  assign n23248 = ~pi1155 & ~n23247;
  assign n23249 = ~n23242 & n23248;
  assign n23250 = n17526 & ~n23211;
  assign n23251 = ~n17526 & n23207;
  assign n23252 = ~n23250 & ~n23251;
  assign n23253 = pi609 & ~n23252;
  assign n23254 = ~pi609 & ~n23211;
  assign n23255 = pi1155 & ~n23254;
  assign n23256 = ~n23253 & n23255;
  assign n23257 = ~pi660 & ~n23256;
  assign n23258 = ~n23249 & n23257;
  assign n23259 = pi609 & ~n23241;
  assign n23260 = ~pi609 & n23246;
  assign n23261 = pi1155 & ~n23260;
  assign n23262 = ~n23259 & n23261;
  assign n23263 = ~pi609 & ~n23252;
  assign n23264 = pi609 & ~n23211;
  assign n23265 = ~pi1155 & ~n23264;
  assign n23266 = ~n23263 & n23265;
  assign n23267 = pi660 & ~n23266;
  assign n23268 = ~n23262 & n23267;
  assign n23269 = ~n23258 & ~n23268;
  assign n23270 = pi785 & ~n23269;
  assign n23271 = ~pi785 & ~n23241;
  assign n23272 = ~n23270 & ~n23271;
  assign n23273 = ~pi618 & ~n23272;
  assign n23274 = n17554 & ~n23211;
  assign n23275 = ~n17554 & n23246;
  assign n23276 = ~n23274 & ~n23275;
  assign n23277 = pi618 & ~n23276;
  assign n23278 = ~pi1154 & ~n23277;
  assign n23279 = ~n23273 & n23278;
  assign n23280 = ~pi785 & n23252;
  assign n23281 = ~n23256 & ~n23266;
  assign n23282 = pi785 & ~n23281;
  assign n23283 = ~n23280 & ~n23282;
  assign n23284 = pi618 & n23283;
  assign n23285 = ~pi618 & ~n23211;
  assign n23286 = pi1154 & ~n23285;
  assign n23287 = ~n23284 & n23286;
  assign n23288 = ~pi627 & ~n23287;
  assign n23289 = ~n23279 & n23288;
  assign n23290 = pi618 & ~n23272;
  assign n23291 = ~pi618 & ~n23276;
  assign n23292 = pi1154 & ~n23291;
  assign n23293 = ~n23290 & n23292;
  assign n23294 = ~pi618 & n23283;
  assign n23295 = pi618 & ~n23211;
  assign n23296 = ~pi1154 & ~n23295;
  assign n23297 = ~n23294 & n23296;
  assign n23298 = pi627 & ~n23297;
  assign n23299 = ~n23293 & n23298;
  assign n23300 = ~n23289 & ~n23299;
  assign n23301 = pi781 & ~n23300;
  assign n23302 = ~pi781 & ~n23272;
  assign n23303 = ~n23301 & ~n23302;
  assign n23304 = ~pi619 & ~n23303;
  assign n23305 = ~n17591 & n23276;
  assign n23306 = n17591 & n23211;
  assign n23307 = ~n23305 & ~n23306;
  assign n23308 = pi619 & n23307;
  assign n23309 = ~pi1159 & ~n23308;
  assign n23310 = ~n23304 & n23309;
  assign n23311 = ~pi781 & ~n23283;
  assign n23312 = ~n23287 & ~n23297;
  assign n23313 = pi781 & ~n23312;
  assign n23314 = ~n23311 & ~n23313;
  assign n23315 = pi619 & n23314;
  assign n23316 = ~pi619 & ~n23211;
  assign n23317 = pi1159 & ~n23316;
  assign n23318 = ~n23315 & n23317;
  assign n23319 = ~pi648 & ~n23318;
  assign n23320 = ~n23310 & n23319;
  assign n23321 = pi619 & ~n23303;
  assign n23322 = ~pi619 & n23307;
  assign n23323 = pi1159 & ~n23322;
  assign n23324 = ~n23321 & n23323;
  assign n23325 = ~pi619 & n23314;
  assign n23326 = pi619 & ~n23211;
  assign n23327 = ~pi1159 & ~n23326;
  assign n23328 = ~n23325 & n23327;
  assign n23329 = pi648 & ~n23328;
  assign n23330 = ~n23324 & n23329;
  assign n23331 = ~n23320 & ~n23330;
  assign n23332 = pi789 & ~n23331;
  assign n23333 = ~pi789 & ~n23303;
  assign n23334 = ~n23332 & ~n23333;
  assign n23335 = ~pi788 & n23334;
  assign n23336 = ~pi626 & n23334;
  assign n23337 = n17627 & ~n23211;
  assign n23338 = ~n17627 & n23307;
  assign n23339 = ~n23337 & ~n23338;
  assign n23340 = pi626 & n23339;
  assign n23341 = ~pi641 & ~n23340;
  assign n23342 = ~n23336 & n23341;
  assign n23343 = ~pi789 & ~n23314;
  assign n23344 = ~n23318 & ~n23328;
  assign n23345 = pi789 & ~n23344;
  assign n23346 = ~n23343 & ~n23345;
  assign n23347 = ~pi626 & ~n23346;
  assign n23348 = pi626 & n23211;
  assign n23349 = pi641 & ~n23348;
  assign n23350 = ~n23347 & n23349;
  assign n23351 = ~pi1158 & ~n23350;
  assign n23352 = ~n23342 & n23351;
  assign n23353 = pi626 & n23334;
  assign n23354 = ~pi626 & n23339;
  assign n23355 = pi641 & ~n23354;
  assign n23356 = ~n23353 & n23355;
  assign n23357 = pi626 & ~n23346;
  assign n23358 = ~pi626 & n23211;
  assign n23359 = ~pi641 & ~n23358;
  assign n23360 = ~n23357 & n23359;
  assign n23361 = pi1158 & ~n23360;
  assign n23362 = ~n23356 & n23361;
  assign n23363 = ~n23352 & ~n23362;
  assign n23364 = pi788 & ~n23363;
  assign n23365 = ~n23335 & ~n23364;
  assign n23366 = ~pi628 & n23365;
  assign n23367 = ~n17904 & ~n23346;
  assign n23368 = n17904 & n23211;
  assign n23369 = ~n23367 & ~n23368;
  assign n23370 = pi628 & n23369;
  assign n23371 = ~pi1156 & ~n23370;
  assign n23372 = ~n23366 & n23371;
  assign n23373 = ~n17670 & n23339;
  assign n23374 = n17670 & n23211;
  assign n23375 = ~n23373 & ~n23374;
  assign n23376 = pi628 & n23375;
  assign n23377 = ~pi628 & ~n23211;
  assign n23378 = pi1156 & ~n23377;
  assign n23379 = ~n23376 & n23378;
  assign n23380 = ~pi629 & ~n23379;
  assign n23381 = ~n23372 & n23380;
  assign n23382 = pi628 & n23365;
  assign n23383 = ~pi628 & n23369;
  assign n23384 = pi1156 & ~n23383;
  assign n23385 = ~n23382 & n23384;
  assign n23386 = ~pi628 & n23375;
  assign n23387 = pi628 & ~n23211;
  assign n23388 = ~pi1156 & ~n23387;
  assign n23389 = ~n23386 & n23388;
  assign n23390 = pi629 & ~n23389;
  assign n23391 = ~n23385 & n23390;
  assign n23392 = ~n23381 & ~n23391;
  assign n23393 = pi792 & ~n23392;
  assign n23394 = ~pi792 & n23365;
  assign n23395 = ~n23393 & ~n23394;
  assign n23396 = ~pi647 & ~n23395;
  assign n23397 = ~n17698 & ~n23369;
  assign n23398 = n17698 & n23211;
  assign n23399 = ~n23397 & ~n23398;
  assign n23400 = pi647 & n23399;
  assign n23401 = ~pi1157 & ~n23400;
  assign n23402 = ~n23396 & n23401;
  assign n23403 = ~pi792 & ~n23375;
  assign n23404 = ~n23379 & ~n23389;
  assign n23405 = pi792 & ~n23404;
  assign n23406 = ~n23403 & ~n23405;
  assign n23407 = pi647 & n23406;
  assign n23408 = ~pi647 & ~n23211;
  assign n23409 = pi1157 & ~n23408;
  assign n23410 = ~n23407 & n23409;
  assign n23411 = ~pi630 & ~n23410;
  assign n23412 = ~n23402 & n23411;
  assign n23413 = pi647 & ~n23395;
  assign n23414 = ~pi647 & n23399;
  assign n23415 = pi1157 & ~n23414;
  assign n23416 = ~n23413 & n23415;
  assign n23417 = ~pi647 & n23406;
  assign n23418 = pi647 & ~n23211;
  assign n23419 = ~pi1157 & ~n23418;
  assign n23420 = ~n23417 & n23419;
  assign n23421 = pi630 & ~n23420;
  assign n23422 = ~n23416 & n23421;
  assign n23423 = ~n23412 & ~n23422;
  assign n23424 = pi787 & ~n23423;
  assign n23425 = ~pi787 & ~n23395;
  assign n23426 = ~n23424 & ~n23425;
  assign n23427 = pi644 & ~n23426;
  assign n23428 = ~pi787 & ~n23406;
  assign n23429 = ~n23410 & ~n23420;
  assign n23430 = pi787 & ~n23429;
  assign n23431 = ~n23428 & ~n23430;
  assign n23432 = ~pi644 & n23431;
  assign n23433 = pi715 & ~n23432;
  assign n23434 = ~n23427 & n23433;
  assign n23435 = n17740 & ~n23211;
  assign n23436 = ~n17740 & n23399;
  assign n23437 = ~n23435 & ~n23436;
  assign n23438 = pi644 & ~n23437;
  assign n23439 = ~pi644 & ~n23211;
  assign n23440 = ~pi715 & ~n23439;
  assign n23441 = ~n23438 & n23440;
  assign n23442 = pi1160 & ~n23441;
  assign n23443 = ~n23434 & n23442;
  assign n23444 = ~pi644 & ~n23426;
  assign n23445 = pi644 & n23431;
  assign n23446 = ~pi715 & ~n23445;
  assign n23447 = ~n23444 & n23446;
  assign n23448 = ~pi644 & ~n23437;
  assign n23449 = pi644 & ~n23211;
  assign n23450 = pi715 & ~n23449;
  assign n23451 = ~n23448 & n23450;
  assign n23452 = ~pi1160 & ~n23451;
  assign n23453 = ~n23447 & n23452;
  assign n23454 = pi790 & ~n23443;
  assign n23455 = ~n23453 & n23454;
  assign n23456 = ~pi790 & n23426;
  assign n23457 = n6294 & ~n23456;
  assign n23458 = ~n23455 & n23457;
  assign n23459 = ~pi174 & ~n6294;
  assign n23460 = ~pi57 & ~n23459;
  assign n23461 = ~n23458 & n23460;
  assign n23462 = pi57 & pi174;
  assign n23463 = ~pi832 & ~n23462;
  assign n23464 = ~n23461 & n23463;
  assign n23465 = pi174 & ~n2755;
  assign n23466 = pi759 & n16933;
  assign n23467 = ~n23465 & ~n23466;
  assign n23468 = pi696 & n17154;
  assign n23469 = n23467 & ~n23468;
  assign n23470 = pi625 & n23468;
  assign n23471 = ~n23469 & ~n23470;
  assign n23472 = ~pi1153 & ~n23471;
  assign n23473 = pi696 & n17153;
  assign n23474 = pi625 & n23473;
  assign n23475 = pi1153 & ~n23465;
  assign n23476 = ~n23474 & n23475;
  assign n23477 = ~pi608 & ~n23476;
  assign n23478 = ~n23472 & n23477;
  assign n23479 = ~n23465 & ~n23473;
  assign n23480 = ~n23474 & ~n23479;
  assign n23481 = ~pi1153 & ~n23480;
  assign n23482 = pi1153 & n23467;
  assign n23483 = ~n23470 & n23482;
  assign n23484 = pi608 & ~n23481;
  assign n23485 = ~n23483 & n23484;
  assign n23486 = ~n23478 & ~n23485;
  assign n23487 = pi778 & ~n23486;
  assign n23488 = ~pi778 & ~n23469;
  assign n23489 = ~n23487 & ~n23488;
  assign n23490 = ~pi609 & ~n23489;
  assign n23491 = ~pi778 & n23479;
  assign n23492 = ~n23476 & ~n23481;
  assign n23493 = pi778 & ~n23492;
  assign n23494 = ~n23491 & ~n23493;
  assign n23495 = pi609 & n23494;
  assign n23496 = ~pi1155 & ~n23495;
  assign n23497 = ~n23490 & n23496;
  assign n23498 = n17527 & n23466;
  assign n23499 = pi1155 & ~n23465;
  assign n23500 = ~n23498 & n23499;
  assign n23501 = ~pi660 & ~n23500;
  assign n23502 = ~n23497 & n23501;
  assign n23503 = pi609 & ~n23489;
  assign n23504 = ~pi609 & n23494;
  assign n23505 = pi1155 & ~n23504;
  assign n23506 = ~n23503 & n23505;
  assign n23507 = n17539 & n23466;
  assign n23508 = ~pi1155 & ~n23465;
  assign n23509 = ~n23507 & n23508;
  assign n23510 = pi660 & ~n23509;
  assign n23511 = ~n23506 & n23510;
  assign n23512 = ~n23502 & ~n23511;
  assign n23513 = pi785 & ~n23512;
  assign n23514 = ~pi785 & ~n23489;
  assign n23515 = ~n23513 & ~n23514;
  assign n23516 = ~pi618 & ~n23515;
  assign n23517 = ~n17554 & n23494;
  assign n23518 = ~n23465 & ~n23517;
  assign n23519 = pi618 & ~n23518;
  assign n23520 = ~pi1154 & ~n23519;
  assign n23521 = ~n23516 & n23520;
  assign n23522 = ~n20159 & n23466;
  assign n23523 = n20247 & n23522;
  assign n23524 = pi1154 & ~n23465;
  assign n23525 = ~n23523 & n23524;
  assign n23526 = ~pi627 & ~n23525;
  assign n23527 = ~n23521 & n23526;
  assign n23528 = pi618 & ~n23515;
  assign n23529 = ~pi618 & ~n23518;
  assign n23530 = pi1154 & ~n23529;
  assign n23531 = ~n23528 & n23530;
  assign n23532 = n20257 & n23522;
  assign n23533 = ~pi1154 & ~n23465;
  assign n23534 = ~n23532 & n23533;
  assign n23535 = pi627 & ~n23534;
  assign n23536 = ~n23531 & n23535;
  assign n23537 = ~n23527 & ~n23536;
  assign n23538 = pi781 & ~n23537;
  assign n23539 = ~pi781 & ~n23515;
  assign n23540 = pi648 & n20162;
  assign n23541 = ~pi648 & n20163;
  assign n23542 = ~n23540 & ~n23541;
  assign n23543 = n17626 & n23542;
  assign n23544 = pi789 & ~n23543;
  assign n23545 = ~n23539 & ~n23544;
  assign n23546 = ~n23538 & n23545;
  assign n23547 = n19216 & n23494;
  assign n23548 = ~n23542 & ~n23547;
  assign n23549 = ~n20169 & n23522;
  assign n23550 = n20282 & n23549;
  assign n23551 = n17625 & ~n23550;
  assign n23552 = n20272 & n23549;
  assign n23553 = n17624 & ~n23552;
  assign n23554 = ~n23551 & ~n23553;
  assign n23555 = ~n23548 & n23554;
  assign n23556 = pi789 & ~n23465;
  assign n23557 = ~n23555 & n23556;
  assign n23558 = n17905 & ~n23557;
  assign n23559 = ~n23546 & n23558;
  assign n23560 = ~n17627 & n23547;
  assign n23561 = ~n23465 & ~n23560;
  assign n23562 = n17786 & ~n23561;
  assign n23563 = n20171 & n23522;
  assign n23564 = ~pi626 & n23563;
  assign n23565 = ~n23465 & ~n23564;
  assign n23566 = ~pi1158 & ~n23565;
  assign n23567 = pi641 & ~n23566;
  assign n23568 = ~n23562 & n23567;
  assign n23569 = n17787 & ~n23561;
  assign n23570 = pi626 & n23563;
  assign n23571 = ~n23465 & ~n23570;
  assign n23572 = pi1158 & ~n23571;
  assign n23573 = ~pi641 & ~n23572;
  assign n23574 = ~n23569 & n23573;
  assign n23575 = pi788 & ~n23568;
  assign n23576 = ~n23574 & n23575;
  assign n23577 = ~n20298 & ~n23576;
  assign n23578 = ~n23559 & n23577;
  assign n23579 = ~n17904 & n23563;
  assign n23580 = ~pi629 & n23579;
  assign n23581 = pi628 & ~n23580;
  assign n23582 = n19217 & n23494;
  assign n23583 = pi629 & ~n23582;
  assign n23584 = ~n23581 & ~n23583;
  assign n23585 = ~pi1156 & ~n23584;
  assign n23586 = pi628 & n23582;
  assign n23587 = ~pi628 & ~n23579;
  assign n23588 = pi629 & ~n23587;
  assign n23589 = pi1156 & ~n23588;
  assign n23590 = ~n23586 & n23589;
  assign n23591 = ~n23585 & ~n23590;
  assign n23592 = pi792 & ~n23465;
  assign n23593 = ~n23591 & n23592;
  assign n23594 = ~n23578 & ~n23593;
  assign n23595 = n20300 & ~n23594;
  assign n23596 = ~n17698 & n23579;
  assign n23597 = ~pi630 & n23596;
  assign n23598 = pi647 & ~n23597;
  assign n23599 = ~n19247 & n23582;
  assign n23600 = pi630 & ~n23599;
  assign n23601 = ~n23598 & ~n23600;
  assign n23602 = ~pi1157 & ~n23601;
  assign n23603 = ~pi630 & ~n23599;
  assign n23604 = pi647 & ~n23603;
  assign n23605 = pi630 & n23596;
  assign n23606 = pi1157 & ~n23605;
  assign n23607 = ~n23604 & n23606;
  assign n23608 = ~n23602 & ~n23607;
  assign n23609 = pi787 & ~n23465;
  assign n23610 = ~n23608 & n23609;
  assign n23611 = ~n23595 & ~n23610;
  assign n23612 = pi644 & n23611;
  assign n23613 = ~n19271 & n23599;
  assign n23614 = ~n23465 & ~n23613;
  assign n23615 = ~pi644 & ~n23614;
  assign n23616 = pi715 & ~n23615;
  assign n23617 = ~n23612 & n23616;
  assign n23618 = ~n17698 & ~n17740;
  assign n23619 = n23579 & n23618;
  assign n23620 = pi644 & n23619;
  assign n23621 = ~pi715 & ~n23465;
  assign n23622 = ~n23620 & n23621;
  assign n23623 = pi1160 & ~n23622;
  assign n23624 = ~n23617 & n23623;
  assign n23625 = ~pi644 & n23611;
  assign n23626 = pi644 & ~n23614;
  assign n23627 = ~pi715 & ~n23626;
  assign n23628 = ~n23625 & n23627;
  assign n23629 = ~pi644 & n23619;
  assign n23630 = pi715 & ~n23465;
  assign n23631 = ~n23629 & n23630;
  assign n23632 = ~pi1160 & ~n23631;
  assign n23633 = ~n23628 & n23632;
  assign n23634 = ~n23624 & ~n23633;
  assign n23635 = pi790 & ~n23634;
  assign n23636 = ~pi790 & n23611;
  assign n23637 = pi832 & ~n23636;
  assign n23638 = ~n23635 & n23637;
  assign po331 = ~n23464 & ~n23638;
  assign n23640 = ~pi175 & ~n2755;
  assign n23641 = pi766 & n16933;
  assign n23642 = ~n23640 & ~n23641;
  assign n23643 = ~n17794 & ~n23642;
  assign n23644 = ~pi785 & ~n23643;
  assign n23645 = n17539 & n23641;
  assign n23646 = n23643 & ~n23645;
  assign n23647 = pi1155 & ~n23646;
  assign n23648 = ~pi1155 & ~n23640;
  assign n23649 = ~n23645 & n23648;
  assign n23650 = ~n23647 & ~n23649;
  assign n23651 = pi785 & ~n23650;
  assign n23652 = ~n23644 & ~n23651;
  assign n23653 = ~pi781 & ~n23652;
  assign n23654 = ~n17809 & n23652;
  assign n23655 = pi1154 & ~n23654;
  assign n23656 = ~n17812 & n23652;
  assign n23657 = ~pi1154 & ~n23656;
  assign n23658 = ~n23655 & ~n23657;
  assign n23659 = pi781 & ~n23658;
  assign n23660 = ~n23653 & ~n23659;
  assign n23661 = ~pi789 & ~n23660;
  assign n23662 = ~n22988 & n23660;
  assign n23663 = pi1159 & ~n23662;
  assign n23664 = ~n22991 & n23660;
  assign n23665 = ~pi1159 & ~n23664;
  assign n23666 = ~n23663 & ~n23665;
  assign n23667 = pi789 & ~n23666;
  assign n23668 = ~n23661 & ~n23667;
  assign n23669 = ~n17904 & n23668;
  assign n23670 = n17904 & n23640;
  assign n23671 = ~n23669 & ~n23670;
  assign n23672 = ~n17698 & ~n23671;
  assign n23673 = n17698 & n23640;
  assign n23674 = ~n23672 & ~n23673;
  assign n23675 = ~n20491 & n23674;
  assign n23676 = pi700 & n17153;
  assign n23677 = ~n23640 & ~n23676;
  assign n23678 = ~pi778 & ~n23677;
  assign n23679 = ~pi625 & n23676;
  assign n23680 = ~n23677 & ~n23679;
  assign n23681 = pi1153 & ~n23680;
  assign n23682 = ~pi1153 & ~n23640;
  assign n23683 = ~n23679 & n23682;
  assign n23684 = pi778 & ~n23683;
  assign n23685 = ~n23681 & n23684;
  assign n23686 = ~n23678 & ~n23685;
  assign n23687 = ~n17780 & ~n23686;
  assign n23688 = ~n17782 & n23687;
  assign n23689 = ~n17784 & n23688;
  assign n23690 = ~n17916 & n23689;
  assign n23691 = ~n17947 & n23690;
  assign n23692 = ~pi647 & n23691;
  assign n23693 = pi647 & n23640;
  assign n23694 = ~pi1157 & ~n23693;
  assign n23695 = ~n23692 & n23694;
  assign n23696 = pi647 & ~n23691;
  assign n23697 = ~pi647 & ~n23640;
  assign n23698 = ~n23696 & ~n23697;
  assign n23699 = pi1157 & ~n23698;
  assign n23700 = ~n23695 & ~n23699;
  assign n23701 = ~n17739 & ~n23700;
  assign n23702 = ~n23675 & ~n23701;
  assign n23703 = pi787 & ~n23702;
  assign n23704 = ~pi626 & ~n23668;
  assign n23705 = pi626 & ~n23640;
  assign n23706 = n17668 & ~n23705;
  assign n23707 = ~n23704 & n23706;
  assign n23708 = pi626 & ~n23668;
  assign n23709 = ~pi626 & ~n23640;
  assign n23710 = n17667 & ~n23709;
  assign n23711 = ~n23708 & n23710;
  assign n23712 = n17792 & n23689;
  assign n23713 = ~n23707 & ~n23712;
  assign n23714 = ~n23711 & n23713;
  assign n23715 = pi788 & ~n23714;
  assign n23716 = ~n16842 & ~n23677;
  assign n23717 = pi625 & n23716;
  assign n23718 = n23642 & ~n23716;
  assign n23719 = ~n23717 & ~n23718;
  assign n23720 = n23682 & ~n23719;
  assign n23721 = ~pi608 & ~n23681;
  assign n23722 = ~n23720 & n23721;
  assign n23723 = pi1153 & n23642;
  assign n23724 = ~n23717 & n23723;
  assign n23725 = pi608 & ~n23683;
  assign n23726 = ~n23724 & n23725;
  assign n23727 = ~n23722 & ~n23726;
  assign n23728 = pi778 & ~n23727;
  assign n23729 = ~pi778 & ~n23718;
  assign n23730 = ~n23728 & ~n23729;
  assign n23731 = ~pi609 & ~n23730;
  assign n23732 = pi609 & ~n23686;
  assign n23733 = ~pi1155 & ~n23732;
  assign n23734 = ~n23731 & n23733;
  assign n23735 = ~pi660 & ~n23647;
  assign n23736 = ~n23734 & n23735;
  assign n23737 = pi609 & ~n23730;
  assign n23738 = ~pi609 & ~n23686;
  assign n23739 = pi1155 & ~n23738;
  assign n23740 = ~n23737 & n23739;
  assign n23741 = pi660 & ~n23649;
  assign n23742 = ~n23740 & n23741;
  assign n23743 = ~n23736 & ~n23742;
  assign n23744 = pi785 & ~n23743;
  assign n23745 = ~pi785 & ~n23730;
  assign n23746 = ~n23744 & ~n23745;
  assign n23747 = ~pi618 & ~n23746;
  assign n23748 = pi618 & n23687;
  assign n23749 = ~pi1154 & ~n23748;
  assign n23750 = ~n23747 & n23749;
  assign n23751 = ~pi627 & ~n23655;
  assign n23752 = ~n23750 & n23751;
  assign n23753 = pi618 & ~n23746;
  assign n23754 = ~pi618 & n23687;
  assign n23755 = pi1154 & ~n23754;
  assign n23756 = ~n23753 & n23755;
  assign n23757 = pi627 & ~n23657;
  assign n23758 = ~n23756 & n23757;
  assign n23759 = ~n23752 & ~n23758;
  assign n23760 = pi781 & ~n23759;
  assign n23761 = ~pi781 & ~n23746;
  assign n23762 = ~n23760 & ~n23761;
  assign n23763 = ~pi619 & ~n23762;
  assign n23764 = pi619 & n23688;
  assign n23765 = ~pi1159 & ~n23764;
  assign n23766 = ~n23763 & n23765;
  assign n23767 = ~pi648 & ~n23663;
  assign n23768 = ~n23766 & n23767;
  assign n23769 = pi619 & ~n23762;
  assign n23770 = ~pi619 & n23688;
  assign n23771 = pi1159 & ~n23770;
  assign n23772 = ~n23769 & n23771;
  assign n23773 = pi648 & ~n23665;
  assign n23774 = ~n23772 & n23773;
  assign n23775 = pi789 & ~n23768;
  assign n23776 = ~n23774 & n23775;
  assign n23777 = ~pi789 & n23762;
  assign n23778 = n17905 & ~n23777;
  assign n23779 = ~n23776 & n23778;
  assign n23780 = ~n23715 & ~n23779;
  assign n23781 = ~n20298 & ~n23780;
  assign n23782 = n17944 & ~n23671;
  assign n23783 = n20786 & n23690;
  assign n23784 = ~n23782 & ~n23783;
  assign n23785 = ~pi629 & ~n23784;
  assign n23786 = n20790 & n23690;
  assign n23787 = n17943 & ~n23671;
  assign n23788 = ~n23786 & ~n23787;
  assign n23789 = pi629 & ~n23788;
  assign n23790 = ~n23785 & ~n23789;
  assign n23791 = pi792 & ~n23790;
  assign n23792 = n20300 & ~n23791;
  assign n23793 = ~n23781 & n23792;
  assign n23794 = ~n23703 & ~n23793;
  assign n23795 = pi644 & n23794;
  assign n23796 = ~pi787 & ~n23691;
  assign n23797 = pi787 & ~n23700;
  assign n23798 = ~n23796 & ~n23797;
  assign n23799 = ~pi644 & n23798;
  assign n23800 = pi715 & ~n23799;
  assign n23801 = ~n23795 & n23800;
  assign n23802 = ~n17740 & ~n23674;
  assign n23803 = n17740 & n23640;
  assign n23804 = ~n23802 & ~n23803;
  assign n23805 = pi644 & ~n23804;
  assign n23806 = ~pi644 & n23640;
  assign n23807 = ~pi715 & ~n23806;
  assign n23808 = ~n23805 & n23807;
  assign n23809 = pi1160 & ~n23808;
  assign n23810 = ~n23801 & n23809;
  assign n23811 = ~pi644 & n23794;
  assign n23812 = pi644 & n23798;
  assign n23813 = ~pi715 & ~n23812;
  assign n23814 = ~n23811 & n23813;
  assign n23815 = ~pi644 & ~n23804;
  assign n23816 = pi644 & n23640;
  assign n23817 = pi715 & ~n23816;
  assign n23818 = ~n23815 & n23817;
  assign n23819 = ~pi1160 & ~n23818;
  assign n23820 = ~n23814 & n23819;
  assign n23821 = ~n23810 & ~n23820;
  assign n23822 = pi790 & ~n23821;
  assign n23823 = ~pi790 & n23794;
  assign n23824 = pi832 & ~n23823;
  assign n23825 = ~n23822 & n23824;
  assign n23826 = ~pi175 & ~n17494;
  assign n23827 = n17627 & ~n23826;
  assign n23828 = pi175 & ~n3268;
  assign n23829 = ~pi175 & n18060;
  assign n23830 = pi175 & ~n18064;
  assign n23831 = ~pi38 & ~n23830;
  assign n23832 = ~n23829 & n23831;
  assign n23833 = ~pi175 & ~n16968;
  assign n23834 = n17480 & ~n23833;
  assign n23835 = pi700 & ~n23834;
  assign n23836 = ~n23832 & n23835;
  assign n23837 = ~pi175 & ~pi700;
  assign n23838 = ~n17487 & n23837;
  assign n23839 = n3268 & ~n23838;
  assign n23840 = ~n23836 & n23839;
  assign n23841 = ~n23828 & ~n23840;
  assign n23842 = ~pi778 & ~n23841;
  assign n23843 = pi625 & n23841;
  assign n23844 = ~pi625 & n23826;
  assign n23845 = pi1153 & ~n23844;
  assign n23846 = ~n23843 & n23845;
  assign n23847 = ~pi625 & n23841;
  assign n23848 = pi625 & n23826;
  assign n23849 = ~pi1153 & ~n23848;
  assign n23850 = ~n23847 & n23849;
  assign n23851 = ~n23846 & ~n23850;
  assign n23852 = pi778 & ~n23851;
  assign n23853 = ~n23842 & ~n23852;
  assign n23854 = ~n17554 & ~n23853;
  assign n23855 = n17554 & ~n23826;
  assign n23856 = ~n23854 & ~n23855;
  assign n23857 = ~n17591 & n23856;
  assign n23858 = n17591 & n23826;
  assign n23859 = ~n23857 & ~n23858;
  assign n23860 = ~n17627 & n23859;
  assign n23861 = ~n23827 & ~n23860;
  assign n23862 = ~n17670 & n23861;
  assign n23863 = n17670 & n23826;
  assign n23864 = ~n23862 & ~n23863;
  assign n23865 = ~pi628 & ~n23864;
  assign n23866 = pi628 & n23826;
  assign n23867 = ~n23865 & ~n23866;
  assign n23868 = ~pi1156 & ~n23867;
  assign n23869 = pi628 & ~n23864;
  assign n23870 = ~pi628 & n23826;
  assign n23871 = ~n23869 & ~n23870;
  assign n23872 = pi1156 & ~n23871;
  assign n23873 = ~n23868 & ~n23872;
  assign n23874 = pi792 & ~n23873;
  assign n23875 = ~pi792 & ~n23864;
  assign n23876 = ~n23874 & ~n23875;
  assign n23877 = ~pi647 & ~n23876;
  assign n23878 = pi647 & n23826;
  assign n23879 = ~n23877 & ~n23878;
  assign n23880 = ~pi1157 & ~n23879;
  assign n23881 = pi647 & ~n23876;
  assign n23882 = ~pi647 & n23826;
  assign n23883 = ~n23881 & ~n23882;
  assign n23884 = pi1157 & ~n23883;
  assign n23885 = ~n23880 & ~n23884;
  assign n23886 = pi787 & ~n23885;
  assign n23887 = ~pi787 & ~n23876;
  assign n23888 = ~n23886 & ~n23887;
  assign n23889 = ~pi644 & ~n23888;
  assign n23890 = pi715 & ~n23889;
  assign n23891 = ~pi766 & n16814;
  assign n23892 = pi175 & n16961;
  assign n23893 = ~n23891 & ~n23892;
  assign n23894 = pi39 & ~n23893;
  assign n23895 = ~pi175 & pi766;
  assign n23896 = n16907 & n23895;
  assign n23897 = pi766 & ~n16919;
  assign n23898 = pi175 & ~n23897;
  assign n23899 = ~n21429 & ~n23898;
  assign n23900 = ~n23896 & n23899;
  assign n23901 = ~n23894 & n23900;
  assign n23902 = ~pi38 & ~n23901;
  assign n23903 = pi766 & n16970;
  assign n23904 = pi38 & ~n23833;
  assign n23905 = ~n23903 & n23904;
  assign n23906 = ~n23902 & ~n23905;
  assign n23907 = n3268 & ~n23906;
  assign n23908 = ~n23828 & ~n23907;
  assign n23909 = ~n17526 & ~n23908;
  assign n23910 = n17526 & ~n23826;
  assign n23911 = ~n23909 & ~n23910;
  assign n23912 = ~pi785 & ~n23911;
  assign n23913 = ~n17527 & ~n23826;
  assign n23914 = pi609 & n23909;
  assign n23915 = ~n23913 & ~n23914;
  assign n23916 = pi1155 & ~n23915;
  assign n23917 = ~n17539 & ~n23826;
  assign n23918 = ~pi609 & n23909;
  assign n23919 = ~n23917 & ~n23918;
  assign n23920 = ~pi1155 & ~n23919;
  assign n23921 = ~n23916 & ~n23920;
  assign n23922 = pi785 & ~n23921;
  assign n23923 = ~n23912 & ~n23922;
  assign n23924 = ~pi781 & ~n23923;
  assign n23925 = pi618 & n23923;
  assign n23926 = ~pi618 & n23826;
  assign n23927 = pi1154 & ~n23926;
  assign n23928 = ~n23925 & n23927;
  assign n23929 = ~pi618 & n23923;
  assign n23930 = pi618 & n23826;
  assign n23931 = ~pi1154 & ~n23930;
  assign n23932 = ~n23929 & n23931;
  assign n23933 = ~n23928 & ~n23932;
  assign n23934 = pi781 & ~n23933;
  assign n23935 = ~n23924 & ~n23934;
  assign n23936 = ~pi789 & ~n23935;
  assign n23937 = pi619 & n23935;
  assign n23938 = ~pi619 & n23826;
  assign n23939 = pi1159 & ~n23938;
  assign n23940 = ~n23937 & n23939;
  assign n23941 = ~pi619 & n23935;
  assign n23942 = pi619 & n23826;
  assign n23943 = ~pi1159 & ~n23942;
  assign n23944 = ~n23941 & n23943;
  assign n23945 = ~n23940 & ~n23944;
  assign n23946 = pi789 & ~n23945;
  assign n23947 = ~n23936 & ~n23946;
  assign n23948 = ~n17904 & n23947;
  assign n23949 = n17904 & n23826;
  assign n23950 = ~n23948 & ~n23949;
  assign n23951 = ~n17698 & ~n23950;
  assign n23952 = n17698 & n23826;
  assign n23953 = ~n23951 & ~n23952;
  assign n23954 = ~n17740 & ~n23953;
  assign n23955 = n17740 & n23826;
  assign n23956 = ~n23954 & ~n23955;
  assign n23957 = pi644 & ~n23956;
  assign n23958 = ~pi644 & n23826;
  assign n23959 = ~pi715 & ~n23958;
  assign n23960 = ~n23957 & n23959;
  assign n23961 = pi1160 & ~n23960;
  assign n23962 = ~n23890 & n23961;
  assign n23963 = pi644 & ~n23888;
  assign n23964 = ~pi715 & ~n23963;
  assign n23965 = ~pi644 & ~n23956;
  assign n23966 = pi644 & n23826;
  assign n23967 = pi715 & ~n23966;
  assign n23968 = ~n23965 & n23967;
  assign n23969 = ~pi1160 & ~n23968;
  assign n23970 = ~n23964 & n23969;
  assign n23971 = ~n23962 & ~n23970;
  assign n23972 = pi790 & ~n23971;
  assign n23973 = ~pi644 & n23969;
  assign n23974 = pi644 & n23961;
  assign n23975 = pi790 & ~n23973;
  assign n23976 = ~n23974 & n23975;
  assign n23977 = ~n20502 & n23950;
  assign n23978 = n17696 & n23867;
  assign n23979 = n17695 & n23871;
  assign n23980 = ~n23978 & ~n23979;
  assign n23981 = ~n23977 & n23980;
  assign n23982 = pi792 & ~n23981;
  assign n23983 = ~pi700 & n23906;
  assign n23984 = ~pi175 & n17074;
  assign n23985 = pi175 & n17166;
  assign n23986 = ~pi766 & ~n23985;
  assign n23987 = ~n23984 & n23986;
  assign n23988 = pi175 & n17233;
  assign n23989 = ~pi175 & ~n17295;
  assign n23990 = pi766 & ~n23989;
  assign n23991 = ~n23988 & n23990;
  assign n23992 = pi39 & ~n23991;
  assign n23993 = ~n23987 & n23992;
  assign n23994 = ~pi175 & n17317;
  assign n23995 = pi175 & n17340;
  assign n23996 = ~pi766 & ~n23994;
  assign n23997 = ~n23995 & n23996;
  assign n23998 = ~pi175 & ~n17344;
  assign n23999 = pi175 & ~n17351;
  assign n24000 = pi766 & ~n23999;
  assign n24001 = ~n23998 & n24000;
  assign n24002 = ~pi39 & ~n24001;
  assign n24003 = ~n23997 & n24002;
  assign n24004 = ~pi38 & ~n24003;
  assign n24005 = ~n23993 & n24004;
  assign n24006 = n16665 & ~n16978;
  assign n24007 = ~pi766 & n24006;
  assign n24008 = ~n17259 & ~n24007;
  assign n24009 = ~pi39 & ~n24008;
  assign n24010 = ~pi175 & ~n24009;
  assign n24011 = ~n17154 & ~n23641;
  assign n24012 = pi175 & ~n24011;
  assign n24013 = n6250 & n24012;
  assign n24014 = pi38 & ~n24013;
  assign n24015 = ~n24010 & n24014;
  assign n24016 = pi700 & ~n24015;
  assign n24017 = ~n24005 & n24016;
  assign n24018 = n3268 & ~n24017;
  assign n24019 = ~n23983 & n24018;
  assign n24020 = ~n23828 & ~n24019;
  assign n24021 = ~pi625 & n24020;
  assign n24022 = pi625 & n23908;
  assign n24023 = ~pi1153 & ~n24022;
  assign n24024 = ~n24021 & n24023;
  assign n24025 = ~pi608 & ~n23846;
  assign n24026 = ~n24024 & n24025;
  assign n24027 = pi625 & n24020;
  assign n24028 = ~pi625 & n23908;
  assign n24029 = pi1153 & ~n24028;
  assign n24030 = ~n24027 & n24029;
  assign n24031 = pi608 & ~n23850;
  assign n24032 = ~n24030 & n24031;
  assign n24033 = ~n24026 & ~n24032;
  assign n24034 = pi778 & ~n24033;
  assign n24035 = ~pi778 & n24020;
  assign n24036 = ~n24034 & ~n24035;
  assign n24037 = ~pi609 & ~n24036;
  assign n24038 = pi609 & n23853;
  assign n24039 = ~pi1155 & ~n24038;
  assign n24040 = ~n24037 & n24039;
  assign n24041 = ~pi660 & ~n23916;
  assign n24042 = ~n24040 & n24041;
  assign n24043 = pi609 & ~n24036;
  assign n24044 = ~pi609 & n23853;
  assign n24045 = pi1155 & ~n24044;
  assign n24046 = ~n24043 & n24045;
  assign n24047 = pi660 & ~n23920;
  assign n24048 = ~n24046 & n24047;
  assign n24049 = ~n24042 & ~n24048;
  assign n24050 = pi785 & ~n24049;
  assign n24051 = ~pi785 & ~n24036;
  assign n24052 = ~n24050 & ~n24051;
  assign n24053 = ~pi618 & ~n24052;
  assign n24054 = pi618 & n23856;
  assign n24055 = ~pi1154 & ~n24054;
  assign n24056 = ~n24053 & n24055;
  assign n24057 = ~pi627 & ~n23928;
  assign n24058 = ~n24056 & n24057;
  assign n24059 = pi618 & ~n24052;
  assign n24060 = ~pi618 & n23856;
  assign n24061 = pi1154 & ~n24060;
  assign n24062 = ~n24059 & n24061;
  assign n24063 = pi627 & ~n23932;
  assign n24064 = ~n24062 & n24063;
  assign n24065 = ~n24058 & ~n24064;
  assign n24066 = pi781 & ~n24065;
  assign n24067 = ~pi781 & ~n24052;
  assign n24068 = ~n24066 & ~n24067;
  assign n24069 = ~pi619 & ~n24068;
  assign n24070 = pi619 & ~n23859;
  assign n24071 = ~pi1159 & ~n24070;
  assign n24072 = ~n24069 & n24071;
  assign n24073 = ~pi648 & ~n23940;
  assign n24074 = ~n24072 & n24073;
  assign n24075 = pi619 & ~n24068;
  assign n24076 = ~pi619 & ~n23859;
  assign n24077 = pi1159 & ~n24076;
  assign n24078 = ~n24075 & n24077;
  assign n24079 = pi648 & ~n23944;
  assign n24080 = ~n24078 & n24079;
  assign n24081 = pi789 & ~n24074;
  assign n24082 = ~n24080 & n24081;
  assign n24083 = ~pi789 & n24068;
  assign n24084 = n17905 & ~n24083;
  assign n24085 = ~n24082 & n24084;
  assign n24086 = ~pi626 & ~n23947;
  assign n24087 = pi626 & ~n23826;
  assign n24088 = n17668 & ~n24087;
  assign n24089 = ~n24086 & n24088;
  assign n24090 = pi626 & ~n23947;
  assign n24091 = ~pi626 & ~n23826;
  assign n24092 = n17667 & ~n24091;
  assign n24093 = ~n24090 & n24092;
  assign n24094 = n17792 & n23861;
  assign n24095 = ~n24089 & ~n24094;
  assign n24096 = ~n24093 & n24095;
  assign n24097 = pi788 & ~n24096;
  assign n24098 = ~n20298 & ~n24097;
  assign n24099 = ~n24085 & n24098;
  assign n24100 = ~n23982 & ~n24099;
  assign n24101 = n20300 & ~n24100;
  assign n24102 = n17737 & n23883;
  assign n24103 = n17738 & n23879;
  assign n24104 = ~n20491 & n23953;
  assign n24105 = ~n24102 & ~n24103;
  assign n24106 = ~n24104 & n24105;
  assign n24107 = pi787 & ~n24106;
  assign n24108 = ~n24101 & ~n24107;
  assign n24109 = ~n23976 & n24108;
  assign n24110 = ~n23972 & ~n24109;
  assign n24111 = ~po1038 & ~n24110;
  assign n24112 = ~pi175 & po1038;
  assign n24113 = ~pi832 & ~n24112;
  assign n24114 = ~n24111 & n24113;
  assign po332 = ~n23825 & ~n24114;
  assign n24116 = ~pi176 & ~n2755;
  assign n24117 = ~pi742 & n16933;
  assign n24118 = ~n24116 & ~n24117;
  assign n24119 = ~n17794 & ~n24118;
  assign n24120 = ~pi785 & ~n24119;
  assign n24121 = ~n17799 & ~n24118;
  assign n24122 = pi1155 & ~n24121;
  assign n24123 = ~n17802 & n24119;
  assign n24124 = ~pi1155 & ~n24123;
  assign n24125 = ~n24122 & ~n24124;
  assign n24126 = pi785 & ~n24125;
  assign n24127 = ~n24120 & ~n24126;
  assign n24128 = ~pi781 & ~n24127;
  assign n24129 = ~n17809 & n24127;
  assign n24130 = pi1154 & ~n24129;
  assign n24131 = ~n17812 & n24127;
  assign n24132 = ~pi1154 & ~n24131;
  assign n24133 = ~n24130 & ~n24132;
  assign n24134 = pi781 & ~n24133;
  assign n24135 = ~n24128 & ~n24134;
  assign n24136 = ~pi789 & ~n24135;
  assign n24137 = pi619 & n24135;
  assign n24138 = ~pi619 & n24116;
  assign n24139 = pi1159 & ~n24138;
  assign n24140 = ~n24137 & n24139;
  assign n24141 = ~pi619 & n24135;
  assign n24142 = pi619 & n24116;
  assign n24143 = ~pi1159 & ~n24142;
  assign n24144 = ~n24141 & n24143;
  assign n24145 = ~n24140 & ~n24144;
  assign n24146 = pi789 & ~n24145;
  assign n24147 = ~n24136 & ~n24146;
  assign n24148 = ~n17904 & n24147;
  assign n24149 = n17904 & n24116;
  assign n24150 = ~n24148 & ~n24149;
  assign n24151 = ~n17698 & ~n24150;
  assign n24152 = n17698 & n24116;
  assign n24153 = ~n24151 & ~n24152;
  assign n24154 = ~n20491 & n24153;
  assign n24155 = ~pi704 & n17153;
  assign n24156 = ~n24116 & ~n24155;
  assign n24157 = ~pi778 & n24156;
  assign n24158 = ~pi625 & n24155;
  assign n24159 = ~n24156 & ~n24158;
  assign n24160 = pi1153 & ~n24159;
  assign n24161 = ~pi1153 & ~n24116;
  assign n24162 = ~n24158 & n24161;
  assign n24163 = ~n24160 & ~n24162;
  assign n24164 = pi778 & ~n24163;
  assign n24165 = ~n24157 & ~n24164;
  assign n24166 = ~n17780 & n24165;
  assign n24167 = ~n17782 & n24166;
  assign n24168 = ~n17784 & n24167;
  assign n24169 = ~n17916 & n24168;
  assign n24170 = ~n17947 & n24169;
  assign n24171 = ~pi647 & n24170;
  assign n24172 = pi647 & n24116;
  assign n24173 = ~pi1157 & ~n24172;
  assign n24174 = ~n24171 & n24173;
  assign n24175 = pi647 & ~n24170;
  assign n24176 = ~pi647 & ~n24116;
  assign n24177 = ~n24175 & ~n24176;
  assign n24178 = pi1157 & ~n24177;
  assign n24179 = ~n24174 & ~n24178;
  assign n24180 = ~n17739 & ~n24179;
  assign n24181 = ~n24154 & ~n24180;
  assign n24182 = pi787 & ~n24181;
  assign n24183 = ~pi626 & ~n24147;
  assign n24184 = pi626 & ~n24116;
  assign n24185 = n17668 & ~n24184;
  assign n24186 = ~n24183 & n24185;
  assign n24187 = pi626 & ~n24147;
  assign n24188 = ~pi626 & ~n24116;
  assign n24189 = n17667 & ~n24188;
  assign n24190 = ~n24187 & n24189;
  assign n24191 = n17792 & n24168;
  assign n24192 = ~n24186 & ~n24191;
  assign n24193 = ~n24190 & n24192;
  assign n24194 = pi788 & ~n24193;
  assign n24195 = ~n16842 & ~n24156;
  assign n24196 = pi625 & n24195;
  assign n24197 = n24118 & ~n24195;
  assign n24198 = ~n24196 & ~n24197;
  assign n24199 = n24161 & ~n24198;
  assign n24200 = ~pi608 & ~n24160;
  assign n24201 = ~n24199 & n24200;
  assign n24202 = pi1153 & n24118;
  assign n24203 = ~n24196 & n24202;
  assign n24204 = pi608 & ~n24162;
  assign n24205 = ~n24203 & n24204;
  assign n24206 = ~n24201 & ~n24205;
  assign n24207 = pi778 & ~n24206;
  assign n24208 = ~pi778 & ~n24197;
  assign n24209 = ~n24207 & ~n24208;
  assign n24210 = ~pi609 & ~n24209;
  assign n24211 = pi609 & n24165;
  assign n24212 = ~pi1155 & ~n24211;
  assign n24213 = ~n24210 & n24212;
  assign n24214 = ~pi660 & ~n24122;
  assign n24215 = ~n24213 & n24214;
  assign n24216 = pi609 & ~n24209;
  assign n24217 = ~pi609 & n24165;
  assign n24218 = pi1155 & ~n24217;
  assign n24219 = ~n24216 & n24218;
  assign n24220 = pi660 & ~n24124;
  assign n24221 = ~n24219 & n24220;
  assign n24222 = ~n24215 & ~n24221;
  assign n24223 = pi785 & ~n24222;
  assign n24224 = ~pi785 & ~n24209;
  assign n24225 = ~n24223 & ~n24224;
  assign n24226 = ~pi618 & ~n24225;
  assign n24227 = pi618 & n24166;
  assign n24228 = ~pi1154 & ~n24227;
  assign n24229 = ~n24226 & n24228;
  assign n24230 = ~pi627 & ~n24130;
  assign n24231 = ~n24229 & n24230;
  assign n24232 = pi618 & ~n24225;
  assign n24233 = ~pi618 & n24166;
  assign n24234 = pi1154 & ~n24233;
  assign n24235 = ~n24232 & n24234;
  assign n24236 = pi627 & ~n24132;
  assign n24237 = ~n24235 & n24236;
  assign n24238 = ~n24231 & ~n24237;
  assign n24239 = pi781 & ~n24238;
  assign n24240 = ~pi781 & ~n24225;
  assign n24241 = ~n24239 & ~n24240;
  assign n24242 = ~pi619 & ~n24241;
  assign n24243 = pi619 & n24167;
  assign n24244 = ~pi1159 & ~n24243;
  assign n24245 = ~n24242 & n24244;
  assign n24246 = ~pi648 & ~n24140;
  assign n24247 = ~n24245 & n24246;
  assign n24248 = pi619 & ~n24241;
  assign n24249 = ~pi619 & n24167;
  assign n24250 = pi1159 & ~n24249;
  assign n24251 = ~n24248 & n24250;
  assign n24252 = pi648 & ~n24144;
  assign n24253 = ~n24251 & n24252;
  assign n24254 = pi789 & ~n24247;
  assign n24255 = ~n24253 & n24254;
  assign n24256 = ~pi789 & n24241;
  assign n24257 = n17905 & ~n24256;
  assign n24258 = ~n24255 & n24257;
  assign n24259 = ~n24194 & ~n24258;
  assign n24260 = ~n20298 & ~n24259;
  assign n24261 = n17944 & ~n24150;
  assign n24262 = n20786 & n24169;
  assign n24263 = ~n24261 & ~n24262;
  assign n24264 = ~pi629 & ~n24263;
  assign n24265 = n20790 & n24169;
  assign n24266 = n17943 & ~n24150;
  assign n24267 = ~n24265 & ~n24266;
  assign n24268 = pi629 & ~n24267;
  assign n24269 = ~n24264 & ~n24268;
  assign n24270 = pi792 & ~n24269;
  assign n24271 = n20300 & ~n24270;
  assign n24272 = ~n24260 & n24271;
  assign n24273 = ~n24182 & ~n24272;
  assign n24274 = pi644 & n24273;
  assign n24275 = ~pi787 & ~n24170;
  assign n24276 = pi787 & ~n24179;
  assign n24277 = ~n24275 & ~n24276;
  assign n24278 = ~pi644 & n24277;
  assign n24279 = pi715 & ~n24278;
  assign n24280 = ~n24274 & n24279;
  assign n24281 = ~n17740 & ~n24153;
  assign n24282 = n17740 & n24116;
  assign n24283 = ~n24281 & ~n24282;
  assign n24284 = pi644 & ~n24283;
  assign n24285 = ~pi644 & n24116;
  assign n24286 = ~pi715 & ~n24285;
  assign n24287 = ~n24284 & n24286;
  assign n24288 = pi1160 & ~n24287;
  assign n24289 = ~n24280 & n24288;
  assign n24290 = ~pi644 & n24273;
  assign n24291 = pi644 & n24277;
  assign n24292 = ~pi715 & ~n24291;
  assign n24293 = ~n24290 & n24292;
  assign n24294 = ~pi644 & ~n24283;
  assign n24295 = pi644 & n24116;
  assign n24296 = pi715 & ~n24295;
  assign n24297 = ~n24294 & n24296;
  assign n24298 = ~pi1160 & ~n24297;
  assign n24299 = ~n24293 & n24298;
  assign n24300 = ~n24289 & ~n24299;
  assign n24301 = pi790 & ~n24300;
  assign n24302 = ~pi790 & n24273;
  assign n24303 = pi832 & ~n24302;
  assign n24304 = ~n24301 & n24303;
  assign n24305 = ~pi176 & ~n17494;
  assign n24306 = n17627 & ~n24305;
  assign n24307 = ~pi38 & n18064;
  assign n24308 = n3268 & ~n17480;
  assign n24309 = ~n24307 & n24308;
  assign n24310 = pi176 & ~n24309;
  assign n24311 = ~pi38 & n18060;
  assign n24312 = ~n19892 & ~n24311;
  assign n24313 = ~pi176 & n24312;
  assign n24314 = ~pi704 & ~n24313;
  assign n24315 = ~pi176 & ~n17487;
  assign n24316 = pi704 & n24315;
  assign n24317 = n3268 & ~n24316;
  assign n24318 = ~n24314 & n24317;
  assign n24319 = ~n24310 & ~n24318;
  assign n24320 = ~pi778 & ~n24319;
  assign n24321 = pi625 & n24319;
  assign n24322 = ~pi625 & n24305;
  assign n24323 = pi1153 & ~n24322;
  assign n24324 = ~n24321 & n24323;
  assign n24325 = ~pi625 & n24319;
  assign n24326 = pi625 & n24305;
  assign n24327 = ~pi1153 & ~n24326;
  assign n24328 = ~n24325 & n24327;
  assign n24329 = ~n24324 & ~n24328;
  assign n24330 = pi778 & ~n24329;
  assign n24331 = ~n24320 & ~n24330;
  assign n24332 = ~n17554 & ~n24331;
  assign n24333 = n17554 & ~n24305;
  assign n24334 = ~n24332 & ~n24333;
  assign n24335 = ~n17591 & n24334;
  assign n24336 = n17591 & n24305;
  assign n24337 = ~n24335 & ~n24336;
  assign n24338 = ~n17627 & n24337;
  assign n24339 = ~n24306 & ~n24338;
  assign n24340 = ~n17670 & n24339;
  assign n24341 = n17670 & n24305;
  assign n24342 = ~n24340 & ~n24341;
  assign n24343 = ~pi628 & ~n24342;
  assign n24344 = pi628 & n24305;
  assign n24345 = ~n24343 & ~n24344;
  assign n24346 = ~pi1156 & ~n24345;
  assign n24347 = pi628 & ~n24342;
  assign n24348 = ~pi628 & n24305;
  assign n24349 = ~n24347 & ~n24348;
  assign n24350 = pi1156 & ~n24349;
  assign n24351 = ~n24346 & ~n24350;
  assign n24352 = pi792 & ~n24351;
  assign n24353 = ~pi792 & ~n24342;
  assign n24354 = ~n24352 & ~n24353;
  assign n24355 = ~pi647 & ~n24354;
  assign n24356 = pi647 & n24305;
  assign n24357 = ~n24355 & ~n24356;
  assign n24358 = ~pi1157 & ~n24357;
  assign n24359 = pi647 & ~n24354;
  assign n24360 = ~pi647 & n24305;
  assign n24361 = ~n24359 & ~n24360;
  assign n24362 = pi1157 & ~n24361;
  assign n24363 = ~n24358 & ~n24362;
  assign n24364 = pi787 & ~n24363;
  assign n24365 = ~pi787 & ~n24354;
  assign n24366 = ~n24364 & ~n24365;
  assign n24367 = ~pi644 & ~n24366;
  assign n24368 = pi715 & ~n24367;
  assign n24369 = pi176 & ~n3268;
  assign n24370 = ~pi176 & n19349;
  assign n24371 = ~n19343 & ~n19344;
  assign n24372 = pi176 & n24371;
  assign n24373 = ~n24370 & ~n24372;
  assign n24374 = ~pi742 & ~n24373;
  assign n24375 = pi742 & ~n24315;
  assign n24376 = ~n24374 & ~n24375;
  assign n24377 = n3268 & ~n24376;
  assign n24378 = ~n24369 & ~n24377;
  assign n24379 = ~n17526 & ~n24378;
  assign n24380 = n17526 & ~n24305;
  assign n24381 = ~n24379 & ~n24380;
  assign n24382 = ~pi785 & ~n24381;
  assign n24383 = ~n17527 & ~n24305;
  assign n24384 = pi609 & n24379;
  assign n24385 = ~n24383 & ~n24384;
  assign n24386 = pi1155 & ~n24385;
  assign n24387 = ~n17539 & ~n24305;
  assign n24388 = ~pi609 & n24379;
  assign n24389 = ~n24387 & ~n24388;
  assign n24390 = ~pi1155 & ~n24389;
  assign n24391 = ~n24386 & ~n24390;
  assign n24392 = pi785 & ~n24391;
  assign n24393 = ~n24382 & ~n24392;
  assign n24394 = ~pi781 & ~n24393;
  assign n24395 = pi618 & n24393;
  assign n24396 = ~pi618 & n24305;
  assign n24397 = pi1154 & ~n24396;
  assign n24398 = ~n24395 & n24397;
  assign n24399 = ~pi618 & n24393;
  assign n24400 = pi618 & n24305;
  assign n24401 = ~pi1154 & ~n24400;
  assign n24402 = ~n24399 & n24401;
  assign n24403 = ~n24398 & ~n24402;
  assign n24404 = pi781 & ~n24403;
  assign n24405 = ~n24394 & ~n24404;
  assign n24406 = ~pi789 & ~n24405;
  assign n24407 = pi619 & n24405;
  assign n24408 = ~pi619 & n24305;
  assign n24409 = pi1159 & ~n24408;
  assign n24410 = ~n24407 & n24409;
  assign n24411 = ~pi619 & n24405;
  assign n24412 = pi619 & n24305;
  assign n24413 = ~pi1159 & ~n24412;
  assign n24414 = ~n24411 & n24413;
  assign n24415 = ~n24410 & ~n24414;
  assign n24416 = pi789 & ~n24415;
  assign n24417 = ~n24406 & ~n24416;
  assign n24418 = ~n17904 & n24417;
  assign n24419 = n17904 & n24305;
  assign n24420 = ~n24418 & ~n24419;
  assign n24421 = ~n17698 & ~n24420;
  assign n24422 = n17698 & n24305;
  assign n24423 = ~n24421 & ~n24422;
  assign n24424 = ~n17740 & ~n24423;
  assign n24425 = n17740 & n24305;
  assign n24426 = ~n24424 & ~n24425;
  assign n24427 = pi644 & ~n24426;
  assign n24428 = ~pi644 & n24305;
  assign n24429 = ~pi715 & ~n24428;
  assign n24430 = ~n24427 & n24429;
  assign n24431 = pi1160 & ~n24430;
  assign n24432 = ~n24368 & n24431;
  assign n24433 = pi644 & ~n24366;
  assign n24434 = ~pi715 & ~n24433;
  assign n24435 = ~pi644 & ~n24426;
  assign n24436 = pi644 & n24305;
  assign n24437 = pi715 & ~n24436;
  assign n24438 = ~n24435 & n24437;
  assign n24439 = ~pi1160 & ~n24438;
  assign n24440 = ~n24434 & n24439;
  assign n24441 = ~n24432 & ~n24440;
  assign n24442 = pi790 & ~n24441;
  assign n24443 = ~n20502 & n24420;
  assign n24444 = n17696 & n24345;
  assign n24445 = n17695 & n24349;
  assign n24446 = ~n24444 & ~n24445;
  assign n24447 = ~n24443 & n24446;
  assign n24448 = pi792 & ~n24447;
  assign n24449 = ~pi626 & ~n24417;
  assign n24450 = pi626 & ~n24305;
  assign n24451 = n17668 & ~n24450;
  assign n24452 = ~n24449 & n24451;
  assign n24453 = pi626 & ~n24417;
  assign n24454 = ~pi626 & ~n24305;
  assign n24455 = n17667 & ~n24454;
  assign n24456 = ~n24453 & n24455;
  assign n24457 = n17792 & n24339;
  assign n24458 = ~n24452 & ~n24457;
  assign n24459 = ~n24456 & n24458;
  assign n24460 = pi788 & ~n24459;
  assign n24461 = ~pi176 & n19309;
  assign n24462 = ~n19314 & ~n19316;
  assign n24463 = pi176 & ~n24462;
  assign n24464 = pi742 & ~n24463;
  assign n24465 = ~n24461 & n24464;
  assign n24466 = pi176 & n19326;
  assign n24467 = ~pi176 & ~n19334;
  assign n24468 = ~pi742 & ~n24467;
  assign n24469 = ~n24466 & n24468;
  assign n24470 = ~pi704 & ~n24469;
  assign n24471 = ~n24465 & n24470;
  assign n24472 = pi704 & n24376;
  assign n24473 = n3268 & ~n24471;
  assign n24474 = ~n24472 & n24473;
  assign n24475 = ~n24369 & ~n24474;
  assign n24476 = ~pi625 & n24475;
  assign n24477 = pi625 & n24378;
  assign n24478 = ~pi1153 & ~n24477;
  assign n24479 = ~n24476 & n24478;
  assign n24480 = ~pi608 & ~n24324;
  assign n24481 = ~n24479 & n24480;
  assign n24482 = pi625 & n24475;
  assign n24483 = ~pi625 & n24378;
  assign n24484 = pi1153 & ~n24483;
  assign n24485 = ~n24482 & n24484;
  assign n24486 = pi608 & ~n24328;
  assign n24487 = ~n24485 & n24486;
  assign n24488 = ~n24481 & ~n24487;
  assign n24489 = pi778 & ~n24488;
  assign n24490 = ~pi778 & n24475;
  assign n24491 = ~n24489 & ~n24490;
  assign n24492 = ~pi609 & ~n24491;
  assign n24493 = pi609 & n24331;
  assign n24494 = ~pi1155 & ~n24493;
  assign n24495 = ~n24492 & n24494;
  assign n24496 = ~pi660 & ~n24386;
  assign n24497 = ~n24495 & n24496;
  assign n24498 = pi609 & ~n24491;
  assign n24499 = ~pi609 & n24331;
  assign n24500 = pi1155 & ~n24499;
  assign n24501 = ~n24498 & n24500;
  assign n24502 = pi660 & ~n24390;
  assign n24503 = ~n24501 & n24502;
  assign n24504 = ~n24497 & ~n24503;
  assign n24505 = pi785 & ~n24504;
  assign n24506 = ~pi785 & ~n24491;
  assign n24507 = ~n24505 & ~n24506;
  assign n24508 = ~pi618 & ~n24507;
  assign n24509 = pi618 & n24334;
  assign n24510 = ~pi1154 & ~n24509;
  assign n24511 = ~n24508 & n24510;
  assign n24512 = ~pi627 & ~n24398;
  assign n24513 = ~n24511 & n24512;
  assign n24514 = pi618 & ~n24507;
  assign n24515 = ~pi618 & n24334;
  assign n24516 = pi1154 & ~n24515;
  assign n24517 = ~n24514 & n24516;
  assign n24518 = pi627 & ~n24402;
  assign n24519 = ~n24517 & n24518;
  assign n24520 = ~n24513 & ~n24519;
  assign n24521 = pi781 & ~n24520;
  assign n24522 = ~pi781 & ~n24507;
  assign n24523 = ~n24521 & ~n24522;
  assign n24524 = ~pi619 & ~n24523;
  assign n24525 = pi619 & ~n24337;
  assign n24526 = ~pi1159 & ~n24525;
  assign n24527 = ~n24524 & n24526;
  assign n24528 = ~pi648 & ~n24410;
  assign n24529 = ~n24527 & n24528;
  assign n24530 = pi619 & ~n24523;
  assign n24531 = ~pi619 & ~n24337;
  assign n24532 = pi1159 & ~n24531;
  assign n24533 = ~n24530 & n24532;
  assign n24534 = pi648 & ~n24414;
  assign n24535 = ~n24533 & n24534;
  assign n24536 = pi789 & ~n24529;
  assign n24537 = ~n24535 & n24536;
  assign n24538 = ~pi789 & n24523;
  assign n24539 = n17905 & ~n24538;
  assign n24540 = ~n24537 & n24539;
  assign n24541 = ~n24460 & ~n24540;
  assign n24542 = ~n24448 & ~n24541;
  assign n24543 = n20298 & n24447;
  assign n24544 = n20300 & ~n24543;
  assign n24545 = ~n24542 & n24544;
  assign n24546 = ~pi644 & n24439;
  assign n24547 = pi644 & n24431;
  assign n24548 = pi790 & ~n24546;
  assign n24549 = ~n24547 & n24548;
  assign n24550 = n17737 & n24361;
  assign n24551 = n17738 & n24357;
  assign n24552 = ~n20491 & n24423;
  assign n24553 = ~n24550 & ~n24551;
  assign n24554 = ~n24552 & n24553;
  assign n24555 = pi787 & ~n24554;
  assign n24556 = ~n24545 & ~n24555;
  assign n24557 = ~n24549 & n24556;
  assign n24558 = ~n24442 & ~n24557;
  assign n24559 = ~po1038 & ~n24558;
  assign n24560 = ~pi176 & po1038;
  assign n24561 = ~pi832 & ~n24560;
  assign n24562 = ~n24559 & n24561;
  assign po333 = ~n24304 & ~n24562;
  assign n24564 = pi177 & ~n3268;
  assign n24565 = ~pi757 & ~n19349;
  assign n24566 = ~n21578 & ~n24565;
  assign n24567 = ~pi177 & ~n24566;
  assign n24568 = ~pi177 & ~n19343;
  assign n24569 = ~pi757 & ~n24568;
  assign n24570 = ~n24371 & n24569;
  assign n24571 = ~n24567 & ~n24570;
  assign n24572 = pi686 & ~n24571;
  assign n24573 = ~pi177 & n19307;
  assign n24574 = pi177 & n19313;
  assign n24575 = ~pi38 & ~n24574;
  assign n24576 = ~n24573 & n24575;
  assign n24577 = ~pi177 & ~n16968;
  assign n24578 = n18046 & ~n24577;
  assign n24579 = pi757 & ~n24578;
  assign n24580 = ~n24576 & n24579;
  assign n24581 = pi177 & n19324;
  assign n24582 = ~n19328 & ~n19329;
  assign n24583 = ~pi177 & ~n24582;
  assign n24584 = ~pi38 & ~n24583;
  assign n24585 = ~n24581 & n24584;
  assign n24586 = ~pi177 & ~n19331;
  assign n24587 = pi177 & n19320;
  assign n24588 = pi38 & ~n24587;
  assign n24589 = ~n24586 & n24588;
  assign n24590 = ~pi757 & ~n24589;
  assign n24591 = ~n24585 & n24590;
  assign n24592 = ~n24580 & ~n24591;
  assign n24593 = ~pi686 & ~n24592;
  assign n24594 = n3268 & ~n24593;
  assign n24595 = ~n24572 & n24594;
  assign n24596 = ~n24564 & ~n24595;
  assign n24597 = ~pi625 & n24596;
  assign n24598 = n3268 & n24571;
  assign n24599 = ~n24564 & ~n24598;
  assign n24600 = pi625 & n24599;
  assign n24601 = ~pi1153 & ~n24600;
  assign n24602 = ~n24597 & n24601;
  assign n24603 = ~pi177 & n18060;
  assign n24604 = pi177 & ~n18064;
  assign n24605 = ~pi38 & ~n24604;
  assign n24606 = ~n24603 & n24605;
  assign n24607 = n17480 & ~n24577;
  assign n24608 = ~pi686 & ~n24607;
  assign n24609 = ~n24606 & n24608;
  assign n24610 = ~pi177 & pi686;
  assign n24611 = ~n17487 & n24610;
  assign n24612 = n3268 & ~n24611;
  assign n24613 = ~n24609 & n24612;
  assign n24614 = ~n24564 & ~n24613;
  assign n24615 = pi625 & n24614;
  assign n24616 = ~pi177 & ~n17494;
  assign n24617 = ~pi625 & n24616;
  assign n24618 = pi1153 & ~n24617;
  assign n24619 = ~n24615 & n24618;
  assign n24620 = ~pi608 & ~n24619;
  assign n24621 = ~n24602 & n24620;
  assign n24622 = pi625 & n24596;
  assign n24623 = ~pi625 & n24599;
  assign n24624 = pi1153 & ~n24623;
  assign n24625 = ~n24622 & n24624;
  assign n24626 = ~pi625 & n24614;
  assign n24627 = pi625 & n24616;
  assign n24628 = ~pi1153 & ~n24627;
  assign n24629 = ~n24626 & n24628;
  assign n24630 = pi608 & ~n24629;
  assign n24631 = ~n24625 & n24630;
  assign n24632 = ~n24621 & ~n24631;
  assign n24633 = pi778 & ~n24632;
  assign n24634 = ~pi778 & n24596;
  assign n24635 = ~n24633 & ~n24634;
  assign n24636 = ~pi609 & ~n24635;
  assign n24637 = ~pi778 & ~n24614;
  assign n24638 = ~n24619 & ~n24629;
  assign n24639 = pi778 & ~n24638;
  assign n24640 = ~n24637 & ~n24639;
  assign n24641 = pi609 & n24640;
  assign n24642 = ~pi1155 & ~n24641;
  assign n24643 = ~n24636 & n24642;
  assign n24644 = ~n17527 & ~n24616;
  assign n24645 = ~n17526 & ~n24599;
  assign n24646 = pi609 & n24645;
  assign n24647 = ~n24644 & ~n24646;
  assign n24648 = pi1155 & ~n24647;
  assign n24649 = ~pi660 & ~n24648;
  assign n24650 = ~n24643 & n24649;
  assign n24651 = pi609 & ~n24635;
  assign n24652 = ~pi609 & n24640;
  assign n24653 = pi1155 & ~n24652;
  assign n24654 = ~n24651 & n24653;
  assign n24655 = ~n17539 & ~n24616;
  assign n24656 = ~pi609 & n24645;
  assign n24657 = ~n24655 & ~n24656;
  assign n24658 = ~pi1155 & ~n24657;
  assign n24659 = pi660 & ~n24658;
  assign n24660 = ~n24654 & n24659;
  assign n24661 = ~n24650 & ~n24660;
  assign n24662 = pi785 & ~n24661;
  assign n24663 = ~pi785 & ~n24635;
  assign n24664 = ~n24662 & ~n24663;
  assign n24665 = ~pi618 & ~n24664;
  assign n24666 = ~n17554 & ~n24640;
  assign n24667 = n17554 & ~n24616;
  assign n24668 = ~n24666 & ~n24667;
  assign n24669 = pi618 & n24668;
  assign n24670 = ~pi1154 & ~n24669;
  assign n24671 = ~n24665 & n24670;
  assign n24672 = n17526 & ~n24616;
  assign n24673 = ~n24645 & ~n24672;
  assign n24674 = ~pi785 & ~n24673;
  assign n24675 = ~n24648 & ~n24658;
  assign n24676 = pi785 & ~n24675;
  assign n24677 = ~n24674 & ~n24676;
  assign n24678 = pi618 & n24677;
  assign n24679 = ~pi618 & n24616;
  assign n24680 = pi1154 & ~n24679;
  assign n24681 = ~n24678 & n24680;
  assign n24682 = ~pi627 & ~n24681;
  assign n24683 = ~n24671 & n24682;
  assign n24684 = pi618 & ~n24664;
  assign n24685 = ~pi618 & n24668;
  assign n24686 = pi1154 & ~n24685;
  assign n24687 = ~n24684 & n24686;
  assign n24688 = ~pi618 & n24677;
  assign n24689 = pi618 & n24616;
  assign n24690 = ~pi1154 & ~n24689;
  assign n24691 = ~n24688 & n24690;
  assign n24692 = pi627 & ~n24691;
  assign n24693 = ~n24687 & n24692;
  assign n24694 = ~n24683 & ~n24693;
  assign n24695 = pi781 & ~n24694;
  assign n24696 = ~pi781 & ~n24664;
  assign n24697 = ~n24695 & ~n24696;
  assign n24698 = ~pi619 & ~n24697;
  assign n24699 = ~n17591 & n24668;
  assign n24700 = n17591 & n24616;
  assign n24701 = ~n24699 & ~n24700;
  assign n24702 = pi619 & ~n24701;
  assign n24703 = ~pi1159 & ~n24702;
  assign n24704 = ~n24698 & n24703;
  assign n24705 = ~pi781 & ~n24677;
  assign n24706 = ~n24681 & ~n24691;
  assign n24707 = pi781 & ~n24706;
  assign n24708 = ~n24705 & ~n24707;
  assign n24709 = pi619 & n24708;
  assign n24710 = ~pi619 & n24616;
  assign n24711 = pi1159 & ~n24710;
  assign n24712 = ~n24709 & n24711;
  assign n24713 = ~pi648 & ~n24712;
  assign n24714 = ~n24704 & n24713;
  assign n24715 = pi619 & ~n24697;
  assign n24716 = ~pi619 & ~n24701;
  assign n24717 = pi1159 & ~n24716;
  assign n24718 = ~n24715 & n24717;
  assign n24719 = ~pi619 & n24708;
  assign n24720 = pi619 & n24616;
  assign n24721 = ~pi1159 & ~n24720;
  assign n24722 = ~n24719 & n24721;
  assign n24723 = pi648 & ~n24722;
  assign n24724 = ~n24718 & n24723;
  assign n24725 = ~n24714 & ~n24724;
  assign n24726 = pi789 & ~n24725;
  assign n24727 = ~pi789 & ~n24697;
  assign n24728 = ~n24726 & ~n24727;
  assign n24729 = ~pi788 & n24728;
  assign n24730 = ~pi626 & n24728;
  assign n24731 = n17627 & ~n24616;
  assign n24732 = ~n17627 & n24701;
  assign n24733 = ~n24731 & ~n24732;
  assign n24734 = pi626 & ~n24733;
  assign n24735 = ~pi641 & ~n24734;
  assign n24736 = ~n24730 & n24735;
  assign n24737 = ~pi789 & ~n24708;
  assign n24738 = ~n24712 & ~n24722;
  assign n24739 = pi789 & ~n24738;
  assign n24740 = ~n24737 & ~n24739;
  assign n24741 = ~pi626 & ~n24740;
  assign n24742 = pi626 & ~n24616;
  assign n24743 = pi641 & ~n24742;
  assign n24744 = ~n24741 & n24743;
  assign n24745 = ~pi1158 & ~n24744;
  assign n24746 = ~n24736 & n24745;
  assign n24747 = pi626 & n24728;
  assign n24748 = ~pi626 & ~n24733;
  assign n24749 = pi641 & ~n24748;
  assign n24750 = ~n24747 & n24749;
  assign n24751 = pi626 & ~n24740;
  assign n24752 = ~pi626 & ~n24616;
  assign n24753 = ~pi641 & ~n24752;
  assign n24754 = ~n24751 & n24753;
  assign n24755 = pi1158 & ~n24754;
  assign n24756 = ~n24750 & n24755;
  assign n24757 = ~n24746 & ~n24756;
  assign n24758 = pi788 & ~n24757;
  assign n24759 = ~n24729 & ~n24758;
  assign n24760 = ~pi628 & n24759;
  assign n24761 = ~n17904 & n24740;
  assign n24762 = n17904 & n24616;
  assign n24763 = ~n24761 & ~n24762;
  assign n24764 = pi628 & ~n24763;
  assign n24765 = ~pi1156 & ~n24764;
  assign n24766 = ~n24760 & n24765;
  assign n24767 = ~n17670 & n24733;
  assign n24768 = n17670 & n24616;
  assign n24769 = ~n24767 & ~n24768;
  assign n24770 = pi628 & ~n24769;
  assign n24771 = ~pi628 & n24616;
  assign n24772 = pi1156 & ~n24771;
  assign n24773 = ~n24770 & n24772;
  assign n24774 = ~pi629 & ~n24773;
  assign n24775 = ~n24766 & n24774;
  assign n24776 = pi628 & n24759;
  assign n24777 = ~pi628 & ~n24763;
  assign n24778 = pi1156 & ~n24777;
  assign n24779 = ~n24776 & n24778;
  assign n24780 = ~pi628 & ~n24769;
  assign n24781 = pi628 & n24616;
  assign n24782 = ~pi1156 & ~n24781;
  assign n24783 = ~n24780 & n24782;
  assign n24784 = pi629 & ~n24783;
  assign n24785 = ~n24779 & n24784;
  assign n24786 = ~n24775 & ~n24785;
  assign n24787 = pi792 & ~n24786;
  assign n24788 = ~pi792 & n24759;
  assign n24789 = ~n24787 & ~n24788;
  assign n24790 = ~pi647 & ~n24789;
  assign n24791 = ~n17698 & ~n24763;
  assign n24792 = n17698 & n24616;
  assign n24793 = ~n24791 & ~n24792;
  assign n24794 = pi647 & ~n24793;
  assign n24795 = ~pi1157 & ~n24794;
  assign n24796 = ~n24790 & n24795;
  assign n24797 = ~pi792 & n24769;
  assign n24798 = ~n24773 & ~n24783;
  assign n24799 = pi792 & ~n24798;
  assign n24800 = ~n24797 & ~n24799;
  assign n24801 = pi647 & n24800;
  assign n24802 = ~pi647 & n24616;
  assign n24803 = pi1157 & ~n24802;
  assign n24804 = ~n24801 & n24803;
  assign n24805 = ~pi630 & ~n24804;
  assign n24806 = ~n24796 & n24805;
  assign n24807 = pi647 & ~n24789;
  assign n24808 = ~pi647 & ~n24793;
  assign n24809 = pi1157 & ~n24808;
  assign n24810 = ~n24807 & n24809;
  assign n24811 = ~pi647 & n24800;
  assign n24812 = pi647 & n24616;
  assign n24813 = ~pi1157 & ~n24812;
  assign n24814 = ~n24811 & n24813;
  assign n24815 = pi630 & ~n24814;
  assign n24816 = ~n24810 & n24815;
  assign n24817 = ~n24806 & ~n24816;
  assign n24818 = pi787 & ~n24817;
  assign n24819 = ~pi787 & ~n24789;
  assign n24820 = ~n24818 & ~n24819;
  assign n24821 = pi644 & ~n24820;
  assign n24822 = ~pi787 & ~n24800;
  assign n24823 = ~n24804 & ~n24814;
  assign n24824 = pi787 & ~n24823;
  assign n24825 = ~n24822 & ~n24824;
  assign n24826 = ~pi644 & n24825;
  assign n24827 = pi715 & ~n24826;
  assign n24828 = ~n24821 & n24827;
  assign n24829 = n17740 & ~n24616;
  assign n24830 = ~n17740 & n24793;
  assign n24831 = ~n24829 & ~n24830;
  assign n24832 = pi644 & n24831;
  assign n24833 = ~pi644 & n24616;
  assign n24834 = ~pi715 & ~n24833;
  assign n24835 = ~n24832 & n24834;
  assign n24836 = pi1160 & ~n24835;
  assign n24837 = ~n24828 & n24836;
  assign n24838 = ~pi644 & ~n24820;
  assign n24839 = pi644 & n24825;
  assign n24840 = ~pi715 & ~n24839;
  assign n24841 = ~n24838 & n24840;
  assign n24842 = ~pi644 & n24831;
  assign n24843 = pi644 & n24616;
  assign n24844 = pi715 & ~n24843;
  assign n24845 = ~n24842 & n24844;
  assign n24846 = ~pi1160 & ~n24845;
  assign n24847 = ~n24841 & n24846;
  assign n24848 = pi790 & ~n24837;
  assign n24849 = ~n24847 & n24848;
  assign n24850 = ~pi790 & n24820;
  assign n24851 = ~po1038 & ~n24850;
  assign n24852 = ~n24849 & n24851;
  assign n24853 = ~pi177 & po1038;
  assign n24854 = ~pi832 & ~n24853;
  assign n24855 = ~n24852 & n24854;
  assign n24856 = ~pi177 & ~n2755;
  assign n24857 = ~pi757 & n16933;
  assign n24858 = ~n24856 & ~n24857;
  assign n24859 = ~n17794 & ~n24858;
  assign n24860 = ~pi785 & ~n24859;
  assign n24861 = ~n17799 & ~n24858;
  assign n24862 = pi1155 & ~n24861;
  assign n24863 = ~n17802 & n24859;
  assign n24864 = ~pi1155 & ~n24863;
  assign n24865 = ~n24862 & ~n24864;
  assign n24866 = pi785 & ~n24865;
  assign n24867 = ~n24860 & ~n24866;
  assign n24868 = ~pi781 & ~n24867;
  assign n24869 = ~n17809 & n24867;
  assign n24870 = pi1154 & ~n24869;
  assign n24871 = ~n17812 & n24867;
  assign n24872 = ~pi1154 & ~n24871;
  assign n24873 = ~n24870 & ~n24872;
  assign n24874 = pi781 & ~n24873;
  assign n24875 = ~n24868 & ~n24874;
  assign n24876 = ~pi789 & ~n24875;
  assign n24877 = pi619 & n24875;
  assign n24878 = ~pi619 & n24856;
  assign n24879 = pi1159 & ~n24878;
  assign n24880 = ~n24877 & n24879;
  assign n24881 = ~pi619 & n24875;
  assign n24882 = pi619 & n24856;
  assign n24883 = ~pi1159 & ~n24882;
  assign n24884 = ~n24881 & n24883;
  assign n24885 = ~n24880 & ~n24884;
  assign n24886 = pi789 & ~n24885;
  assign n24887 = ~n24876 & ~n24886;
  assign n24888 = ~n17904 & n24887;
  assign n24889 = n17904 & n24856;
  assign n24890 = ~n24888 & ~n24889;
  assign n24891 = ~n17698 & ~n24890;
  assign n24892 = n17698 & n24856;
  assign n24893 = ~n24891 & ~n24892;
  assign n24894 = ~n20491 & n24893;
  assign n24895 = ~pi686 & n17153;
  assign n24896 = ~n24856 & ~n24895;
  assign n24897 = ~pi778 & n24896;
  assign n24898 = ~pi625 & n24895;
  assign n24899 = ~n24896 & ~n24898;
  assign n24900 = pi1153 & ~n24899;
  assign n24901 = ~pi1153 & ~n24856;
  assign n24902 = ~n24898 & n24901;
  assign n24903 = ~n24900 & ~n24902;
  assign n24904 = pi778 & ~n24903;
  assign n24905 = ~n24897 & ~n24904;
  assign n24906 = ~n17780 & n24905;
  assign n24907 = ~n17782 & n24906;
  assign n24908 = ~n17784 & n24907;
  assign n24909 = ~n17916 & n24908;
  assign n24910 = ~n17947 & n24909;
  assign n24911 = ~pi647 & n24910;
  assign n24912 = pi647 & n24856;
  assign n24913 = ~pi1157 & ~n24912;
  assign n24914 = ~n24911 & n24913;
  assign n24915 = pi647 & ~n24910;
  assign n24916 = ~pi647 & ~n24856;
  assign n24917 = ~n24915 & ~n24916;
  assign n24918 = pi1157 & ~n24917;
  assign n24919 = ~n24914 & ~n24918;
  assign n24920 = ~n17739 & ~n24919;
  assign n24921 = ~n24894 & ~n24920;
  assign n24922 = pi787 & ~n24921;
  assign n24923 = ~pi626 & ~n24887;
  assign n24924 = pi626 & ~n24856;
  assign n24925 = n17668 & ~n24924;
  assign n24926 = ~n24923 & n24925;
  assign n24927 = pi626 & ~n24887;
  assign n24928 = ~pi626 & ~n24856;
  assign n24929 = n17667 & ~n24928;
  assign n24930 = ~n24927 & n24929;
  assign n24931 = n17792 & n24908;
  assign n24932 = ~n24926 & ~n24931;
  assign n24933 = ~n24930 & n24932;
  assign n24934 = pi788 & ~n24933;
  assign n24935 = ~n16842 & ~n24896;
  assign n24936 = pi625 & n24935;
  assign n24937 = n24858 & ~n24935;
  assign n24938 = ~n24936 & ~n24937;
  assign n24939 = n24901 & ~n24938;
  assign n24940 = ~pi608 & ~n24900;
  assign n24941 = ~n24939 & n24940;
  assign n24942 = pi1153 & n24858;
  assign n24943 = ~n24936 & n24942;
  assign n24944 = pi608 & ~n24902;
  assign n24945 = ~n24943 & n24944;
  assign n24946 = ~n24941 & ~n24945;
  assign n24947 = pi778 & ~n24946;
  assign n24948 = ~pi778 & ~n24937;
  assign n24949 = ~n24947 & ~n24948;
  assign n24950 = ~pi609 & ~n24949;
  assign n24951 = pi609 & n24905;
  assign n24952 = ~pi1155 & ~n24951;
  assign n24953 = ~n24950 & n24952;
  assign n24954 = ~pi660 & ~n24862;
  assign n24955 = ~n24953 & n24954;
  assign n24956 = pi609 & ~n24949;
  assign n24957 = ~pi609 & n24905;
  assign n24958 = pi1155 & ~n24957;
  assign n24959 = ~n24956 & n24958;
  assign n24960 = pi660 & ~n24864;
  assign n24961 = ~n24959 & n24960;
  assign n24962 = ~n24955 & ~n24961;
  assign n24963 = pi785 & ~n24962;
  assign n24964 = ~pi785 & ~n24949;
  assign n24965 = ~n24963 & ~n24964;
  assign n24966 = ~pi618 & ~n24965;
  assign n24967 = pi618 & n24906;
  assign n24968 = ~pi1154 & ~n24967;
  assign n24969 = ~n24966 & n24968;
  assign n24970 = ~pi627 & ~n24870;
  assign n24971 = ~n24969 & n24970;
  assign n24972 = pi618 & ~n24965;
  assign n24973 = ~pi618 & n24906;
  assign n24974 = pi1154 & ~n24973;
  assign n24975 = ~n24972 & n24974;
  assign n24976 = pi627 & ~n24872;
  assign n24977 = ~n24975 & n24976;
  assign n24978 = ~n24971 & ~n24977;
  assign n24979 = pi781 & ~n24978;
  assign n24980 = ~pi781 & ~n24965;
  assign n24981 = ~n24979 & ~n24980;
  assign n24982 = ~pi619 & ~n24981;
  assign n24983 = pi619 & n24907;
  assign n24984 = ~pi1159 & ~n24983;
  assign n24985 = ~n24982 & n24984;
  assign n24986 = ~pi648 & ~n24880;
  assign n24987 = ~n24985 & n24986;
  assign n24988 = pi619 & ~n24981;
  assign n24989 = ~pi619 & n24907;
  assign n24990 = pi1159 & ~n24989;
  assign n24991 = ~n24988 & n24990;
  assign n24992 = pi648 & ~n24884;
  assign n24993 = ~n24991 & n24992;
  assign n24994 = pi789 & ~n24987;
  assign n24995 = ~n24993 & n24994;
  assign n24996 = ~pi789 & n24981;
  assign n24997 = n17905 & ~n24996;
  assign n24998 = ~n24995 & n24997;
  assign n24999 = ~n24934 & ~n24998;
  assign n25000 = ~n20298 & ~n24999;
  assign n25001 = n17944 & ~n24890;
  assign n25002 = n20786 & n24909;
  assign n25003 = ~n25001 & ~n25002;
  assign n25004 = ~pi629 & ~n25003;
  assign n25005 = n20790 & n24909;
  assign n25006 = n17943 & ~n24890;
  assign n25007 = ~n25005 & ~n25006;
  assign n25008 = pi629 & ~n25007;
  assign n25009 = ~n25004 & ~n25008;
  assign n25010 = pi792 & ~n25009;
  assign n25011 = n20300 & ~n25010;
  assign n25012 = ~n25000 & n25011;
  assign n25013 = ~n24922 & ~n25012;
  assign n25014 = pi644 & n25013;
  assign n25015 = ~pi787 & ~n24910;
  assign n25016 = pi787 & ~n24919;
  assign n25017 = ~n25015 & ~n25016;
  assign n25018 = ~pi644 & n25017;
  assign n25019 = pi715 & ~n25018;
  assign n25020 = ~n25014 & n25019;
  assign n25021 = ~n17740 & ~n24893;
  assign n25022 = n17740 & n24856;
  assign n25023 = ~n25021 & ~n25022;
  assign n25024 = pi644 & ~n25023;
  assign n25025 = ~pi644 & n24856;
  assign n25026 = ~pi715 & ~n25025;
  assign n25027 = ~n25024 & n25026;
  assign n25028 = pi1160 & ~n25027;
  assign n25029 = ~n25020 & n25028;
  assign n25030 = ~pi644 & n25013;
  assign n25031 = pi644 & n25017;
  assign n25032 = ~pi715 & ~n25031;
  assign n25033 = ~n25030 & n25032;
  assign n25034 = ~pi644 & ~n25023;
  assign n25035 = pi644 & n24856;
  assign n25036 = pi715 & ~n25035;
  assign n25037 = ~n25034 & n25036;
  assign n25038 = ~pi1160 & ~n25037;
  assign n25039 = ~n25033 & n25038;
  assign n25040 = ~n25029 & ~n25039;
  assign n25041 = pi790 & ~n25040;
  assign n25042 = ~pi790 & n25013;
  assign n25043 = pi832 & ~n25042;
  assign n25044 = ~n25041 & n25043;
  assign po334 = ~n24855 & ~n25044;
  assign n25046 = ~pi178 & ~n2755;
  assign n25047 = ~pi760 & n16933;
  assign n25048 = ~n25046 & ~n25047;
  assign n25049 = ~n17794 & ~n25048;
  assign n25050 = ~pi785 & ~n25049;
  assign n25051 = n17539 & n25047;
  assign n25052 = n25049 & ~n25051;
  assign n25053 = pi1155 & ~n25052;
  assign n25054 = ~pi1155 & ~n25046;
  assign n25055 = ~n25051 & n25054;
  assign n25056 = ~n25053 & ~n25055;
  assign n25057 = pi785 & ~n25056;
  assign n25058 = ~n25050 & ~n25057;
  assign n25059 = ~pi781 & ~n25058;
  assign n25060 = ~n17809 & n25058;
  assign n25061 = pi1154 & ~n25060;
  assign n25062 = ~n17812 & n25058;
  assign n25063 = ~pi1154 & ~n25062;
  assign n25064 = ~n25061 & ~n25063;
  assign n25065 = pi781 & ~n25064;
  assign n25066 = ~n25059 & ~n25065;
  assign n25067 = ~pi789 & ~n25066;
  assign n25068 = ~n22988 & n25066;
  assign n25069 = pi1159 & ~n25068;
  assign n25070 = ~n22991 & n25066;
  assign n25071 = ~pi1159 & ~n25070;
  assign n25072 = ~n25069 & ~n25071;
  assign n25073 = pi789 & ~n25072;
  assign n25074 = ~n25067 & ~n25073;
  assign n25075 = ~n17904 & n25074;
  assign n25076 = n17904 & n25046;
  assign n25077 = ~n25075 & ~n25076;
  assign n25078 = ~n17698 & ~n25077;
  assign n25079 = n17698 & n25046;
  assign n25080 = ~n25078 & ~n25079;
  assign n25081 = ~n20491 & n25080;
  assign n25082 = ~pi688 & n17153;
  assign n25083 = ~n25046 & ~n25082;
  assign n25084 = ~pi778 & ~n25083;
  assign n25085 = ~pi625 & n25082;
  assign n25086 = ~n25083 & ~n25085;
  assign n25087 = pi1153 & ~n25086;
  assign n25088 = ~pi1153 & ~n25046;
  assign n25089 = ~n25085 & n25088;
  assign n25090 = pi778 & ~n25089;
  assign n25091 = ~n25087 & n25090;
  assign n25092 = ~n25084 & ~n25091;
  assign n25093 = ~n17780 & ~n25092;
  assign n25094 = ~n17782 & n25093;
  assign n25095 = ~n17784 & n25094;
  assign n25096 = ~n17916 & n25095;
  assign n25097 = ~n17947 & n25096;
  assign n25098 = ~pi647 & n25097;
  assign n25099 = pi647 & n25046;
  assign n25100 = ~pi1157 & ~n25099;
  assign n25101 = ~n25098 & n25100;
  assign n25102 = pi647 & ~n25097;
  assign n25103 = ~pi647 & ~n25046;
  assign n25104 = ~n25102 & ~n25103;
  assign n25105 = pi1157 & ~n25104;
  assign n25106 = ~n25101 & ~n25105;
  assign n25107 = ~n17739 & ~n25106;
  assign n25108 = ~n25081 & ~n25107;
  assign n25109 = pi787 & ~n25108;
  assign n25110 = ~pi626 & ~n25074;
  assign n25111 = pi626 & ~n25046;
  assign n25112 = n17668 & ~n25111;
  assign n25113 = ~n25110 & n25112;
  assign n25114 = pi626 & ~n25074;
  assign n25115 = ~pi626 & ~n25046;
  assign n25116 = n17667 & ~n25115;
  assign n25117 = ~n25114 & n25116;
  assign n25118 = n17792 & n25095;
  assign n25119 = ~n25113 & ~n25118;
  assign n25120 = ~n25117 & n25119;
  assign n25121 = pi788 & ~n25120;
  assign n25122 = ~n16842 & ~n25083;
  assign n25123 = pi625 & n25122;
  assign n25124 = n25048 & ~n25122;
  assign n25125 = ~n25123 & ~n25124;
  assign n25126 = n25088 & ~n25125;
  assign n25127 = ~pi608 & ~n25087;
  assign n25128 = ~n25126 & n25127;
  assign n25129 = pi1153 & n25048;
  assign n25130 = ~n25123 & n25129;
  assign n25131 = pi608 & ~n25089;
  assign n25132 = ~n25130 & n25131;
  assign n25133 = ~n25128 & ~n25132;
  assign n25134 = pi778 & ~n25133;
  assign n25135 = ~pi778 & ~n25124;
  assign n25136 = ~n25134 & ~n25135;
  assign n25137 = ~pi609 & ~n25136;
  assign n25138 = pi609 & ~n25092;
  assign n25139 = ~pi1155 & ~n25138;
  assign n25140 = ~n25137 & n25139;
  assign n25141 = ~pi660 & ~n25053;
  assign n25142 = ~n25140 & n25141;
  assign n25143 = pi609 & ~n25136;
  assign n25144 = ~pi609 & ~n25092;
  assign n25145 = pi1155 & ~n25144;
  assign n25146 = ~n25143 & n25145;
  assign n25147 = pi660 & ~n25055;
  assign n25148 = ~n25146 & n25147;
  assign n25149 = ~n25142 & ~n25148;
  assign n25150 = pi785 & ~n25149;
  assign n25151 = ~pi785 & ~n25136;
  assign n25152 = ~n25150 & ~n25151;
  assign n25153 = ~pi618 & ~n25152;
  assign n25154 = pi618 & n25093;
  assign n25155 = ~pi1154 & ~n25154;
  assign n25156 = ~n25153 & n25155;
  assign n25157 = ~pi627 & ~n25061;
  assign n25158 = ~n25156 & n25157;
  assign n25159 = pi618 & ~n25152;
  assign n25160 = ~pi618 & n25093;
  assign n25161 = pi1154 & ~n25160;
  assign n25162 = ~n25159 & n25161;
  assign n25163 = pi627 & ~n25063;
  assign n25164 = ~n25162 & n25163;
  assign n25165 = ~n25158 & ~n25164;
  assign n25166 = pi781 & ~n25165;
  assign n25167 = ~pi781 & ~n25152;
  assign n25168 = ~n25166 & ~n25167;
  assign n25169 = ~pi619 & ~n25168;
  assign n25170 = pi619 & n25094;
  assign n25171 = ~pi1159 & ~n25170;
  assign n25172 = ~n25169 & n25171;
  assign n25173 = ~pi648 & ~n25069;
  assign n25174 = ~n25172 & n25173;
  assign n25175 = pi619 & ~n25168;
  assign n25176 = ~pi619 & n25094;
  assign n25177 = pi1159 & ~n25176;
  assign n25178 = ~n25175 & n25177;
  assign n25179 = pi648 & ~n25071;
  assign n25180 = ~n25178 & n25179;
  assign n25181 = pi789 & ~n25174;
  assign n25182 = ~n25180 & n25181;
  assign n25183 = ~pi789 & n25168;
  assign n25184 = n17905 & ~n25183;
  assign n25185 = ~n25182 & n25184;
  assign n25186 = ~n25121 & ~n25185;
  assign n25187 = ~n20298 & ~n25186;
  assign n25188 = n17944 & ~n25077;
  assign n25189 = n20786 & n25096;
  assign n25190 = ~n25188 & ~n25189;
  assign n25191 = ~pi629 & ~n25190;
  assign n25192 = n20790 & n25096;
  assign n25193 = n17943 & ~n25077;
  assign n25194 = ~n25192 & ~n25193;
  assign n25195 = pi629 & ~n25194;
  assign n25196 = ~n25191 & ~n25195;
  assign n25197 = pi792 & ~n25196;
  assign n25198 = n20300 & ~n25197;
  assign n25199 = ~n25187 & n25198;
  assign n25200 = ~n25109 & ~n25199;
  assign n25201 = pi644 & n25200;
  assign n25202 = ~pi787 & ~n25097;
  assign n25203 = pi787 & ~n25106;
  assign n25204 = ~n25202 & ~n25203;
  assign n25205 = ~pi644 & n25204;
  assign n25206 = pi715 & ~n25205;
  assign n25207 = ~n25201 & n25206;
  assign n25208 = ~n17740 & ~n25080;
  assign n25209 = n17740 & n25046;
  assign n25210 = ~n25208 & ~n25209;
  assign n25211 = pi644 & ~n25210;
  assign n25212 = ~pi644 & n25046;
  assign n25213 = ~pi715 & ~n25212;
  assign n25214 = ~n25211 & n25213;
  assign n25215 = pi1160 & ~n25214;
  assign n25216 = ~n25207 & n25215;
  assign n25217 = ~pi644 & n25200;
  assign n25218 = pi644 & n25204;
  assign n25219 = ~pi715 & ~n25218;
  assign n25220 = ~n25217 & n25219;
  assign n25221 = ~pi644 & ~n25210;
  assign n25222 = pi644 & n25046;
  assign n25223 = pi715 & ~n25222;
  assign n25224 = ~n25221 & n25223;
  assign n25225 = ~pi1160 & ~n25224;
  assign n25226 = ~n25220 & n25225;
  assign n25227 = ~n25216 & ~n25226;
  assign n25228 = pi790 & ~n25227;
  assign n25229 = ~pi790 & n25200;
  assign n25230 = pi832 & ~n25229;
  assign n25231 = ~n25228 & n25230;
  assign n25232 = ~pi178 & ~n17494;
  assign n25233 = n17627 & ~n25232;
  assign n25234 = ~pi688 & n3268;
  assign n25235 = n25232 & ~n25234;
  assign n25236 = pi178 & ~n18064;
  assign n25237 = ~pi38 & ~n25236;
  assign n25238 = n3268 & ~n25237;
  assign n25239 = ~pi178 & n18060;
  assign n25240 = ~n25238 & ~n25239;
  assign n25241 = ~pi178 & ~n16968;
  assign n25242 = n17480 & ~n25241;
  assign n25243 = ~pi688 & ~n25242;
  assign n25244 = ~n25240 & n25243;
  assign n25245 = ~n25235 & ~n25244;
  assign n25246 = ~pi778 & n25245;
  assign n25247 = pi625 & ~n25245;
  assign n25248 = ~pi625 & n25232;
  assign n25249 = pi1153 & ~n25248;
  assign n25250 = ~n25247 & n25249;
  assign n25251 = ~pi625 & ~n25245;
  assign n25252 = pi625 & n25232;
  assign n25253 = ~pi1153 & ~n25252;
  assign n25254 = ~n25251 & n25253;
  assign n25255 = ~n25250 & ~n25254;
  assign n25256 = pi778 & ~n25255;
  assign n25257 = ~n25246 & ~n25256;
  assign n25258 = ~n17554 & ~n25257;
  assign n25259 = n17554 & ~n25232;
  assign n25260 = ~n25258 & ~n25259;
  assign n25261 = ~n17591 & n25260;
  assign n25262 = n17591 & n25232;
  assign n25263 = ~n25261 & ~n25262;
  assign n25264 = ~n17627 & n25263;
  assign n25265 = ~n25233 & ~n25264;
  assign n25266 = ~n17670 & n25265;
  assign n25267 = n17670 & n25232;
  assign n25268 = ~n25266 & ~n25267;
  assign n25269 = ~pi792 & n25268;
  assign n25270 = pi628 & ~n25268;
  assign n25271 = ~pi628 & n25232;
  assign n25272 = pi1156 & ~n25271;
  assign n25273 = ~n25270 & n25272;
  assign n25274 = ~pi628 & ~n25268;
  assign n25275 = pi628 & n25232;
  assign n25276 = ~pi1156 & ~n25275;
  assign n25277 = ~n25274 & n25276;
  assign n25278 = ~n25273 & ~n25277;
  assign n25279 = pi792 & ~n25278;
  assign n25280 = ~n25269 & ~n25279;
  assign n25281 = ~pi647 & ~n25280;
  assign n25282 = pi647 & ~n25232;
  assign n25283 = ~n25281 & ~n25282;
  assign n25284 = ~pi1157 & n25283;
  assign n25285 = pi647 & ~n25280;
  assign n25286 = ~pi647 & ~n25232;
  assign n25287 = ~n25285 & ~n25286;
  assign n25288 = pi1157 & n25287;
  assign n25289 = ~n25284 & ~n25288;
  assign n25290 = pi787 & ~n25289;
  assign n25291 = ~pi787 & n25280;
  assign n25292 = ~n25290 & ~n25291;
  assign n25293 = ~pi644 & ~n25292;
  assign n25294 = pi715 & ~n25293;
  assign n25295 = pi178 & ~n3268;
  assign n25296 = ~pi760 & n16970;
  assign n25297 = ~n25241 & ~n25296;
  assign n25298 = pi38 & ~n25297;
  assign n25299 = ~pi178 & n16907;
  assign n25300 = pi178 & ~n16963;
  assign n25301 = ~pi760 & ~n25300;
  assign n25302 = ~n25299 & n25301;
  assign n25303 = ~pi178 & pi760;
  assign n25304 = ~n16816 & n25303;
  assign n25305 = ~n25302 & ~n25304;
  assign n25306 = ~pi38 & ~n25305;
  assign n25307 = ~n25298 & ~n25306;
  assign n25308 = n3268 & n25307;
  assign n25309 = ~n25295 & ~n25308;
  assign n25310 = ~n17526 & ~n25309;
  assign n25311 = n17526 & ~n25232;
  assign n25312 = ~n25310 & ~n25311;
  assign n25313 = ~pi785 & ~n25312;
  assign n25314 = ~n17527 & ~n25232;
  assign n25315 = pi609 & n25310;
  assign n25316 = ~n25314 & ~n25315;
  assign n25317 = pi1155 & ~n25316;
  assign n25318 = ~n17539 & ~n25232;
  assign n25319 = ~pi609 & n25310;
  assign n25320 = ~n25318 & ~n25319;
  assign n25321 = ~pi1155 & ~n25320;
  assign n25322 = ~n25317 & ~n25321;
  assign n25323 = pi785 & ~n25322;
  assign n25324 = ~n25313 & ~n25323;
  assign n25325 = ~pi781 & ~n25324;
  assign n25326 = pi618 & n25324;
  assign n25327 = ~pi618 & n25232;
  assign n25328 = pi1154 & ~n25327;
  assign n25329 = ~n25326 & n25328;
  assign n25330 = ~pi618 & n25324;
  assign n25331 = pi618 & n25232;
  assign n25332 = ~pi1154 & ~n25331;
  assign n25333 = ~n25330 & n25332;
  assign n25334 = ~n25329 & ~n25333;
  assign n25335 = pi781 & ~n25334;
  assign n25336 = ~n25325 & ~n25335;
  assign n25337 = ~pi789 & ~n25336;
  assign n25338 = pi619 & n25336;
  assign n25339 = ~pi619 & n25232;
  assign n25340 = pi1159 & ~n25339;
  assign n25341 = ~n25338 & n25340;
  assign n25342 = ~pi619 & n25336;
  assign n25343 = pi619 & n25232;
  assign n25344 = ~pi1159 & ~n25343;
  assign n25345 = ~n25342 & n25344;
  assign n25346 = ~n25341 & ~n25345;
  assign n25347 = pi789 & ~n25346;
  assign n25348 = ~n25337 & ~n25347;
  assign n25349 = ~n17904 & n25348;
  assign n25350 = n17904 & n25232;
  assign n25351 = ~n25349 & ~n25350;
  assign n25352 = ~n17698 & ~n25351;
  assign n25353 = n17698 & n25232;
  assign n25354 = ~n25352 & ~n25353;
  assign n25355 = ~n17740 & ~n25354;
  assign n25356 = n17740 & n25232;
  assign n25357 = ~n25355 & ~n25356;
  assign n25358 = pi644 & ~n25357;
  assign n25359 = ~pi644 & n25232;
  assign n25360 = ~pi715 & ~n25359;
  assign n25361 = ~n25358 & n25360;
  assign n25362 = pi1160 & ~n25361;
  assign n25363 = ~n25294 & n25362;
  assign n25364 = pi644 & ~n25292;
  assign n25365 = ~pi715 & ~n25364;
  assign n25366 = ~pi644 & ~n25357;
  assign n25367 = pi644 & n25232;
  assign n25368 = pi715 & ~n25367;
  assign n25369 = ~n25366 & n25368;
  assign n25370 = ~pi1160 & ~n25369;
  assign n25371 = ~n25365 & n25370;
  assign n25372 = ~n25363 & ~n25371;
  assign n25373 = pi790 & ~n25372;
  assign n25374 = ~pi644 & n25370;
  assign n25375 = pi644 & n25362;
  assign n25376 = pi790 & ~n25374;
  assign n25377 = ~n25375 & n25376;
  assign n25378 = ~n20502 & n25351;
  assign n25379 = ~pi629 & n25273;
  assign n25380 = pi629 & n25277;
  assign n25381 = ~n25379 & ~n25380;
  assign n25382 = ~n25378 & n25381;
  assign n25383 = pi792 & ~n25382;
  assign n25384 = pi688 & ~n25307;
  assign n25385 = ~pi178 & n17074;
  assign n25386 = pi178 & n17166;
  assign n25387 = pi760 & ~n25386;
  assign n25388 = ~n25385 & n25387;
  assign n25389 = pi178 & n17233;
  assign n25390 = ~pi178 & ~n17295;
  assign n25391 = ~pi760 & ~n25390;
  assign n25392 = ~n25389 & n25391;
  assign n25393 = pi39 & ~n25392;
  assign n25394 = ~n25388 & n25393;
  assign n25395 = pi178 & ~n17340;
  assign n25396 = ~pi178 & ~n17317;
  assign n25397 = pi760 & ~n25395;
  assign n25398 = ~n25396 & n25397;
  assign n25399 = ~pi178 & n17344;
  assign n25400 = pi178 & n17351;
  assign n25401 = ~pi760 & ~n25400;
  assign n25402 = ~n25399 & n25401;
  assign n25403 = ~n25398 & ~n25402;
  assign n25404 = ~pi39 & ~n25403;
  assign n25405 = ~pi38 & ~n25404;
  assign n25406 = ~n25394 & n25405;
  assign n25407 = ~pi760 & ~n17259;
  assign n25408 = n19303 & ~n25407;
  assign n25409 = ~pi178 & ~n25408;
  assign n25410 = ~n17154 & ~n25047;
  assign n25411 = pi178 & ~n25410;
  assign n25412 = n6250 & n25411;
  assign n25413 = pi38 & ~n25412;
  assign n25414 = ~n25409 & n25413;
  assign n25415 = ~pi688 & ~n25414;
  assign n25416 = ~n25406 & n25415;
  assign n25417 = n3268 & ~n25416;
  assign n25418 = ~n25384 & n25417;
  assign n25419 = ~n25295 & ~n25418;
  assign n25420 = ~pi625 & n25419;
  assign n25421 = pi625 & n25309;
  assign n25422 = ~pi1153 & ~n25421;
  assign n25423 = ~n25420 & n25422;
  assign n25424 = ~pi608 & ~n25250;
  assign n25425 = ~n25423 & n25424;
  assign n25426 = pi625 & n25419;
  assign n25427 = ~pi625 & n25309;
  assign n25428 = pi1153 & ~n25427;
  assign n25429 = ~n25426 & n25428;
  assign n25430 = pi608 & ~n25254;
  assign n25431 = ~n25429 & n25430;
  assign n25432 = ~n25425 & ~n25431;
  assign n25433 = pi778 & ~n25432;
  assign n25434 = ~pi778 & n25419;
  assign n25435 = ~n25433 & ~n25434;
  assign n25436 = ~pi609 & ~n25435;
  assign n25437 = pi609 & n25257;
  assign n25438 = ~pi1155 & ~n25437;
  assign n25439 = ~n25436 & n25438;
  assign n25440 = ~pi660 & ~n25317;
  assign n25441 = ~n25439 & n25440;
  assign n25442 = pi609 & ~n25435;
  assign n25443 = ~pi609 & n25257;
  assign n25444 = pi1155 & ~n25443;
  assign n25445 = ~n25442 & n25444;
  assign n25446 = pi660 & ~n25321;
  assign n25447 = ~n25445 & n25446;
  assign n25448 = ~n25441 & ~n25447;
  assign n25449 = pi785 & ~n25448;
  assign n25450 = ~pi785 & ~n25435;
  assign n25451 = ~n25449 & ~n25450;
  assign n25452 = ~pi618 & ~n25451;
  assign n25453 = pi618 & n25260;
  assign n25454 = ~pi1154 & ~n25453;
  assign n25455 = ~n25452 & n25454;
  assign n25456 = ~pi627 & ~n25329;
  assign n25457 = ~n25455 & n25456;
  assign n25458 = pi618 & ~n25451;
  assign n25459 = ~pi618 & n25260;
  assign n25460 = pi1154 & ~n25459;
  assign n25461 = ~n25458 & n25460;
  assign n25462 = pi627 & ~n25333;
  assign n25463 = ~n25461 & n25462;
  assign n25464 = ~n25457 & ~n25463;
  assign n25465 = pi781 & ~n25464;
  assign n25466 = ~pi781 & ~n25451;
  assign n25467 = ~n25465 & ~n25466;
  assign n25468 = ~pi619 & ~n25467;
  assign n25469 = pi619 & ~n25263;
  assign n25470 = ~pi1159 & ~n25469;
  assign n25471 = ~n25468 & n25470;
  assign n25472 = ~pi648 & ~n25341;
  assign n25473 = ~n25471 & n25472;
  assign n25474 = pi619 & ~n25467;
  assign n25475 = ~pi619 & ~n25263;
  assign n25476 = pi1159 & ~n25475;
  assign n25477 = ~n25474 & n25476;
  assign n25478 = pi648 & ~n25345;
  assign n25479 = ~n25477 & n25478;
  assign n25480 = pi789 & ~n25473;
  assign n25481 = ~n25479 & n25480;
  assign n25482 = ~pi789 & n25467;
  assign n25483 = n17905 & ~n25482;
  assign n25484 = ~n25481 & n25483;
  assign n25485 = ~pi626 & ~n25348;
  assign n25486 = pi626 & ~n25232;
  assign n25487 = n17668 & ~n25486;
  assign n25488 = ~n25485 & n25487;
  assign n25489 = pi626 & ~n25348;
  assign n25490 = ~pi626 & ~n25232;
  assign n25491 = n17667 & ~n25490;
  assign n25492 = ~n25489 & n25491;
  assign n25493 = n17792 & n25265;
  assign n25494 = ~n25488 & ~n25493;
  assign n25495 = ~n25492 & n25494;
  assign n25496 = pi788 & ~n25495;
  assign n25497 = ~n20298 & ~n25496;
  assign n25498 = ~n25484 & n25497;
  assign n25499 = ~n25383 & ~n25498;
  assign n25500 = n20300 & ~n25499;
  assign n25501 = ~n20491 & n25354;
  assign n25502 = n17738 & ~n25283;
  assign n25503 = n17737 & ~n25287;
  assign n25504 = ~n25502 & ~n25503;
  assign n25505 = ~n25501 & n25504;
  assign n25506 = pi787 & ~n25505;
  assign n25507 = ~n25500 & ~n25506;
  assign n25508 = ~n25377 & n25507;
  assign n25509 = ~n25373 & ~n25508;
  assign n25510 = ~po1038 & ~n25509;
  assign n25511 = ~pi178 & po1038;
  assign n25512 = ~pi832 & ~n25511;
  assign n25513 = ~n25510 & n25512;
  assign po335 = ~n25231 & ~n25513;
  assign n25515 = pi179 & ~n3268;
  assign n25516 = ~pi179 & ~n16968;
  assign n25517 = n18046 & ~n25516;
  assign n25518 = ~pi179 & n17074;
  assign n25519 = pi179 & n17166;
  assign n25520 = pi39 & ~n25519;
  assign n25521 = ~n25518 & n25520;
  assign n25522 = ~pi179 & n17317;
  assign n25523 = pi179 & n17340;
  assign n25524 = ~pi39 & ~n25522;
  assign n25525 = ~n25523 & n25524;
  assign n25526 = ~n25521 & ~n25525;
  assign n25527 = ~pi38 & ~n25526;
  assign n25528 = ~n25517 & ~n25527;
  assign n25529 = pi741 & ~n25528;
  assign n25530 = pi179 & n19326;
  assign n25531 = ~pi179 & ~n19334;
  assign n25532 = ~pi741 & ~n25531;
  assign n25533 = ~n25530 & n25532;
  assign n25534 = ~pi724 & ~n25533;
  assign n25535 = ~n25529 & n25534;
  assign n25536 = ~pi741 & ~n24371;
  assign n25537 = pi179 & ~n25536;
  assign n25538 = ~pi179 & ~pi741;
  assign n25539 = ~n19343 & n25538;
  assign n25540 = n19349 & n25539;
  assign n25541 = ~n25537 & ~n25540;
  assign n25542 = ~n21606 & n25541;
  assign n25543 = n3268 & ~n25542;
  assign n25544 = ~pi724 & n3268;
  assign n25545 = ~n25543 & ~n25544;
  assign n25546 = ~n25535 & ~n25545;
  assign n25547 = ~n25515 & ~n25546;
  assign n25548 = ~pi625 & n25547;
  assign n25549 = ~n25515 & ~n25543;
  assign n25550 = pi625 & n25549;
  assign n25551 = ~pi1153 & ~n25550;
  assign n25552 = ~n25548 & n25551;
  assign n25553 = ~pi179 & ~n17494;
  assign n25554 = ~n25544 & n25553;
  assign n25555 = ~pi179 & n18060;
  assign n25556 = pi179 & ~n18064;
  assign n25557 = ~pi38 & ~n25556;
  assign n25558 = n3268 & ~n25557;
  assign n25559 = ~n25555 & ~n25558;
  assign n25560 = n17480 & ~n25516;
  assign n25561 = ~pi724 & ~n25560;
  assign n25562 = ~n25559 & n25561;
  assign n25563 = ~n25554 & ~n25562;
  assign n25564 = pi625 & ~n25563;
  assign n25565 = ~pi625 & n25553;
  assign n25566 = pi1153 & ~n25565;
  assign n25567 = ~n25564 & n25566;
  assign n25568 = ~pi608 & ~n25567;
  assign n25569 = ~n25552 & n25568;
  assign n25570 = pi625 & n25547;
  assign n25571 = ~pi625 & n25549;
  assign n25572 = pi1153 & ~n25571;
  assign n25573 = ~n25570 & n25572;
  assign n25574 = ~pi625 & ~n25563;
  assign n25575 = pi625 & n25553;
  assign n25576 = ~pi1153 & ~n25575;
  assign n25577 = ~n25574 & n25576;
  assign n25578 = pi608 & ~n25577;
  assign n25579 = ~n25573 & n25578;
  assign n25580 = ~n25569 & ~n25579;
  assign n25581 = pi778 & ~n25580;
  assign n25582 = ~pi778 & n25547;
  assign n25583 = ~n25581 & ~n25582;
  assign n25584 = ~pi609 & ~n25583;
  assign n25585 = ~pi778 & n25563;
  assign n25586 = ~n25567 & ~n25577;
  assign n25587 = pi778 & ~n25586;
  assign n25588 = ~n25585 & ~n25587;
  assign n25589 = pi609 & n25588;
  assign n25590 = ~pi1155 & ~n25589;
  assign n25591 = ~n25584 & n25590;
  assign n25592 = ~n17527 & ~n25553;
  assign n25593 = ~n17526 & ~n25549;
  assign n25594 = pi609 & n25593;
  assign n25595 = ~n25592 & ~n25594;
  assign n25596 = pi1155 & ~n25595;
  assign n25597 = ~pi660 & ~n25596;
  assign n25598 = ~n25591 & n25597;
  assign n25599 = pi609 & ~n25583;
  assign n25600 = ~pi609 & n25588;
  assign n25601 = pi1155 & ~n25600;
  assign n25602 = ~n25599 & n25601;
  assign n25603 = ~n17539 & ~n25553;
  assign n25604 = ~pi609 & n25593;
  assign n25605 = ~n25603 & ~n25604;
  assign n25606 = ~pi1155 & ~n25605;
  assign n25607 = pi660 & ~n25606;
  assign n25608 = ~n25602 & n25607;
  assign n25609 = ~n25598 & ~n25608;
  assign n25610 = pi785 & ~n25609;
  assign n25611 = ~pi785 & ~n25583;
  assign n25612 = ~n25610 & ~n25611;
  assign n25613 = ~pi618 & ~n25612;
  assign n25614 = ~n17554 & ~n25588;
  assign n25615 = n17554 & ~n25553;
  assign n25616 = ~n25614 & ~n25615;
  assign n25617 = pi618 & n25616;
  assign n25618 = ~pi1154 & ~n25617;
  assign n25619 = ~n25613 & n25618;
  assign n25620 = n17526 & ~n25553;
  assign n25621 = ~n25593 & ~n25620;
  assign n25622 = ~pi785 & ~n25621;
  assign n25623 = ~n25596 & ~n25606;
  assign n25624 = pi785 & ~n25623;
  assign n25625 = ~n25622 & ~n25624;
  assign n25626 = pi618 & n25625;
  assign n25627 = ~pi618 & n25553;
  assign n25628 = pi1154 & ~n25627;
  assign n25629 = ~n25626 & n25628;
  assign n25630 = ~pi627 & ~n25629;
  assign n25631 = ~n25619 & n25630;
  assign n25632 = pi618 & ~n25612;
  assign n25633 = ~pi618 & n25616;
  assign n25634 = pi1154 & ~n25633;
  assign n25635 = ~n25632 & n25634;
  assign n25636 = ~pi618 & n25625;
  assign n25637 = pi618 & n25553;
  assign n25638 = ~pi1154 & ~n25637;
  assign n25639 = ~n25636 & n25638;
  assign n25640 = pi627 & ~n25639;
  assign n25641 = ~n25635 & n25640;
  assign n25642 = ~n25631 & ~n25641;
  assign n25643 = pi781 & ~n25642;
  assign n25644 = ~pi781 & ~n25612;
  assign n25645 = ~n25643 & ~n25644;
  assign n25646 = ~pi619 & ~n25645;
  assign n25647 = ~n17591 & n25616;
  assign n25648 = n17591 & n25553;
  assign n25649 = ~n25647 & ~n25648;
  assign n25650 = pi619 & ~n25649;
  assign n25651 = ~pi1159 & ~n25650;
  assign n25652 = ~n25646 & n25651;
  assign n25653 = ~pi781 & ~n25625;
  assign n25654 = ~n25629 & ~n25639;
  assign n25655 = pi781 & ~n25654;
  assign n25656 = ~n25653 & ~n25655;
  assign n25657 = pi619 & n25656;
  assign n25658 = ~pi619 & n25553;
  assign n25659 = pi1159 & ~n25658;
  assign n25660 = ~n25657 & n25659;
  assign n25661 = ~pi648 & ~n25660;
  assign n25662 = ~n25652 & n25661;
  assign n25663 = pi619 & ~n25645;
  assign n25664 = ~pi619 & ~n25649;
  assign n25665 = pi1159 & ~n25664;
  assign n25666 = ~n25663 & n25665;
  assign n25667 = ~pi619 & n25656;
  assign n25668 = pi619 & n25553;
  assign n25669 = ~pi1159 & ~n25668;
  assign n25670 = ~n25667 & n25669;
  assign n25671 = pi648 & ~n25670;
  assign n25672 = ~n25666 & n25671;
  assign n25673 = ~n25662 & ~n25672;
  assign n25674 = pi789 & ~n25673;
  assign n25675 = ~pi789 & ~n25645;
  assign n25676 = ~n25674 & ~n25675;
  assign n25677 = ~pi788 & n25676;
  assign n25678 = ~pi626 & n25676;
  assign n25679 = n17627 & ~n25553;
  assign n25680 = ~n17627 & n25649;
  assign n25681 = ~n25679 & ~n25680;
  assign n25682 = pi626 & ~n25681;
  assign n25683 = ~pi641 & ~n25682;
  assign n25684 = ~n25678 & n25683;
  assign n25685 = ~pi789 & ~n25656;
  assign n25686 = ~n25660 & ~n25670;
  assign n25687 = pi789 & ~n25686;
  assign n25688 = ~n25685 & ~n25687;
  assign n25689 = ~pi626 & ~n25688;
  assign n25690 = pi626 & ~n25553;
  assign n25691 = pi641 & ~n25690;
  assign n25692 = ~n25689 & n25691;
  assign n25693 = ~pi1158 & ~n25692;
  assign n25694 = ~n25684 & n25693;
  assign n25695 = pi626 & n25676;
  assign n25696 = ~pi626 & ~n25681;
  assign n25697 = pi641 & ~n25696;
  assign n25698 = ~n25695 & n25697;
  assign n25699 = pi626 & ~n25688;
  assign n25700 = ~pi626 & ~n25553;
  assign n25701 = ~pi641 & ~n25700;
  assign n25702 = ~n25699 & n25701;
  assign n25703 = pi1158 & ~n25702;
  assign n25704 = ~n25698 & n25703;
  assign n25705 = ~n25694 & ~n25704;
  assign n25706 = pi788 & ~n25705;
  assign n25707 = ~n25677 & ~n25706;
  assign n25708 = ~pi628 & n25707;
  assign n25709 = ~n17904 & n25688;
  assign n25710 = n17904 & n25553;
  assign n25711 = ~n25709 & ~n25710;
  assign n25712 = pi628 & ~n25711;
  assign n25713 = ~pi1156 & ~n25712;
  assign n25714 = ~n25708 & n25713;
  assign n25715 = ~n17670 & n25681;
  assign n25716 = n17670 & n25553;
  assign n25717 = ~n25715 & ~n25716;
  assign n25718 = pi628 & ~n25717;
  assign n25719 = ~pi628 & n25553;
  assign n25720 = pi1156 & ~n25719;
  assign n25721 = ~n25718 & n25720;
  assign n25722 = ~pi629 & ~n25721;
  assign n25723 = ~n25714 & n25722;
  assign n25724 = pi628 & n25707;
  assign n25725 = ~pi628 & ~n25711;
  assign n25726 = pi1156 & ~n25725;
  assign n25727 = ~n25724 & n25726;
  assign n25728 = ~pi628 & ~n25717;
  assign n25729 = pi628 & n25553;
  assign n25730 = ~pi1156 & ~n25729;
  assign n25731 = ~n25728 & n25730;
  assign n25732 = pi629 & ~n25731;
  assign n25733 = ~n25727 & n25732;
  assign n25734 = ~n25723 & ~n25733;
  assign n25735 = pi792 & ~n25734;
  assign n25736 = ~pi792 & n25707;
  assign n25737 = ~n25735 & ~n25736;
  assign n25738 = ~pi647 & ~n25737;
  assign n25739 = ~n17698 & ~n25711;
  assign n25740 = n17698 & n25553;
  assign n25741 = ~n25739 & ~n25740;
  assign n25742 = pi647 & ~n25741;
  assign n25743 = ~pi1157 & ~n25742;
  assign n25744 = ~n25738 & n25743;
  assign n25745 = ~pi792 & n25717;
  assign n25746 = ~n25721 & ~n25731;
  assign n25747 = pi792 & ~n25746;
  assign n25748 = ~n25745 & ~n25747;
  assign n25749 = pi647 & n25748;
  assign n25750 = ~pi647 & n25553;
  assign n25751 = pi1157 & ~n25750;
  assign n25752 = ~n25749 & n25751;
  assign n25753 = ~pi630 & ~n25752;
  assign n25754 = ~n25744 & n25753;
  assign n25755 = pi647 & ~n25737;
  assign n25756 = ~pi647 & ~n25741;
  assign n25757 = pi1157 & ~n25756;
  assign n25758 = ~n25755 & n25757;
  assign n25759 = ~pi647 & n25748;
  assign n25760 = pi647 & n25553;
  assign n25761 = ~pi1157 & ~n25760;
  assign n25762 = ~n25759 & n25761;
  assign n25763 = pi630 & ~n25762;
  assign n25764 = ~n25758 & n25763;
  assign n25765 = ~n25754 & ~n25764;
  assign n25766 = pi787 & ~n25765;
  assign n25767 = ~pi787 & ~n25737;
  assign n25768 = ~n25766 & ~n25767;
  assign n25769 = pi644 & ~n25768;
  assign n25770 = ~pi787 & ~n25748;
  assign n25771 = ~n25752 & ~n25762;
  assign n25772 = pi787 & ~n25771;
  assign n25773 = ~n25770 & ~n25772;
  assign n25774 = ~pi644 & n25773;
  assign n25775 = pi715 & ~n25774;
  assign n25776 = ~n25769 & n25775;
  assign n25777 = n17740 & ~n25553;
  assign n25778 = ~n17740 & n25741;
  assign n25779 = ~n25777 & ~n25778;
  assign n25780 = pi644 & n25779;
  assign n25781 = ~pi644 & n25553;
  assign n25782 = ~pi715 & ~n25781;
  assign n25783 = ~n25780 & n25782;
  assign n25784 = pi1160 & ~n25783;
  assign n25785 = ~n25776 & n25784;
  assign n25786 = ~pi644 & ~n25768;
  assign n25787 = pi644 & n25773;
  assign n25788 = ~pi715 & ~n25787;
  assign n25789 = ~n25786 & n25788;
  assign n25790 = ~pi644 & n25779;
  assign n25791 = pi644 & n25553;
  assign n25792 = pi715 & ~n25791;
  assign n25793 = ~n25790 & n25792;
  assign n25794 = ~pi1160 & ~n25793;
  assign n25795 = ~n25789 & n25794;
  assign n25796 = pi790 & ~n25785;
  assign n25797 = ~n25795 & n25796;
  assign n25798 = ~pi790 & n25768;
  assign n25799 = ~po1038 & ~n25798;
  assign n25800 = ~n25797 & n25799;
  assign n25801 = ~pi179 & po1038;
  assign n25802 = ~pi832 & ~n25801;
  assign n25803 = ~n25800 & n25802;
  assign n25804 = ~pi179 & ~n2755;
  assign n25805 = ~pi741 & n16933;
  assign n25806 = ~n25804 & ~n25805;
  assign n25807 = ~n17794 & ~n25806;
  assign n25808 = ~pi785 & ~n25807;
  assign n25809 = ~n17799 & ~n25806;
  assign n25810 = pi1155 & ~n25809;
  assign n25811 = ~n17802 & n25807;
  assign n25812 = ~pi1155 & ~n25811;
  assign n25813 = ~n25810 & ~n25812;
  assign n25814 = pi785 & ~n25813;
  assign n25815 = ~n25808 & ~n25814;
  assign n25816 = ~pi781 & ~n25815;
  assign n25817 = ~n17809 & n25815;
  assign n25818 = pi1154 & ~n25817;
  assign n25819 = ~n17812 & n25815;
  assign n25820 = ~pi1154 & ~n25819;
  assign n25821 = ~n25818 & ~n25820;
  assign n25822 = pi781 & ~n25821;
  assign n25823 = ~n25816 & ~n25822;
  assign n25824 = ~pi789 & ~n25823;
  assign n25825 = pi619 & n25823;
  assign n25826 = ~pi619 & n25804;
  assign n25827 = pi1159 & ~n25826;
  assign n25828 = ~n25825 & n25827;
  assign n25829 = ~pi619 & n25823;
  assign n25830 = pi619 & n25804;
  assign n25831 = ~pi1159 & ~n25830;
  assign n25832 = ~n25829 & n25831;
  assign n25833 = ~n25828 & ~n25832;
  assign n25834 = pi789 & ~n25833;
  assign n25835 = ~n25824 & ~n25834;
  assign n25836 = ~n17904 & n25835;
  assign n25837 = n17904 & n25804;
  assign n25838 = ~n25836 & ~n25837;
  assign n25839 = ~n17698 & ~n25838;
  assign n25840 = n17698 & n25804;
  assign n25841 = ~n25839 & ~n25840;
  assign n25842 = ~n20491 & n25841;
  assign n25843 = ~pi724 & n17153;
  assign n25844 = ~n25804 & ~n25843;
  assign n25845 = ~pi778 & n25844;
  assign n25846 = ~pi625 & n25843;
  assign n25847 = ~n25844 & ~n25846;
  assign n25848 = pi1153 & ~n25847;
  assign n25849 = ~pi1153 & ~n25804;
  assign n25850 = ~n25846 & n25849;
  assign n25851 = ~n25848 & ~n25850;
  assign n25852 = pi778 & ~n25851;
  assign n25853 = ~n25845 & ~n25852;
  assign n25854 = ~n17780 & n25853;
  assign n25855 = ~n17782 & n25854;
  assign n25856 = ~n17784 & n25855;
  assign n25857 = ~n17916 & n25856;
  assign n25858 = ~n17947 & n25857;
  assign n25859 = ~pi647 & n25858;
  assign n25860 = pi647 & n25804;
  assign n25861 = ~pi1157 & ~n25860;
  assign n25862 = ~n25859 & n25861;
  assign n25863 = pi647 & ~n25858;
  assign n25864 = ~pi647 & ~n25804;
  assign n25865 = ~n25863 & ~n25864;
  assign n25866 = pi1157 & ~n25865;
  assign n25867 = ~n25862 & ~n25866;
  assign n25868 = ~n17739 & ~n25867;
  assign n25869 = ~n25842 & ~n25868;
  assign n25870 = pi787 & ~n25869;
  assign n25871 = ~pi626 & ~n25835;
  assign n25872 = pi626 & ~n25804;
  assign n25873 = n17668 & ~n25872;
  assign n25874 = ~n25871 & n25873;
  assign n25875 = pi626 & ~n25835;
  assign n25876 = ~pi626 & ~n25804;
  assign n25877 = n17667 & ~n25876;
  assign n25878 = ~n25875 & n25877;
  assign n25879 = n17792 & n25856;
  assign n25880 = ~n25874 & ~n25879;
  assign n25881 = ~n25878 & n25880;
  assign n25882 = pi788 & ~n25881;
  assign n25883 = ~n16842 & ~n25844;
  assign n25884 = pi625 & n25883;
  assign n25885 = n25806 & ~n25883;
  assign n25886 = ~n25884 & ~n25885;
  assign n25887 = n25849 & ~n25886;
  assign n25888 = ~pi608 & ~n25848;
  assign n25889 = ~n25887 & n25888;
  assign n25890 = pi1153 & n25806;
  assign n25891 = ~n25884 & n25890;
  assign n25892 = pi608 & ~n25850;
  assign n25893 = ~n25891 & n25892;
  assign n25894 = ~n25889 & ~n25893;
  assign n25895 = pi778 & ~n25894;
  assign n25896 = ~pi778 & ~n25885;
  assign n25897 = ~n25895 & ~n25896;
  assign n25898 = ~pi609 & ~n25897;
  assign n25899 = pi609 & n25853;
  assign n25900 = ~pi1155 & ~n25899;
  assign n25901 = ~n25898 & n25900;
  assign n25902 = ~pi660 & ~n25810;
  assign n25903 = ~n25901 & n25902;
  assign n25904 = pi609 & ~n25897;
  assign n25905 = ~pi609 & n25853;
  assign n25906 = pi1155 & ~n25905;
  assign n25907 = ~n25904 & n25906;
  assign n25908 = pi660 & ~n25812;
  assign n25909 = ~n25907 & n25908;
  assign n25910 = ~n25903 & ~n25909;
  assign n25911 = pi785 & ~n25910;
  assign n25912 = ~pi785 & ~n25897;
  assign n25913 = ~n25911 & ~n25912;
  assign n25914 = ~pi618 & ~n25913;
  assign n25915 = pi618 & n25854;
  assign n25916 = ~pi1154 & ~n25915;
  assign n25917 = ~n25914 & n25916;
  assign n25918 = ~pi627 & ~n25818;
  assign n25919 = ~n25917 & n25918;
  assign n25920 = pi618 & ~n25913;
  assign n25921 = ~pi618 & n25854;
  assign n25922 = pi1154 & ~n25921;
  assign n25923 = ~n25920 & n25922;
  assign n25924 = pi627 & ~n25820;
  assign n25925 = ~n25923 & n25924;
  assign n25926 = ~n25919 & ~n25925;
  assign n25927 = pi781 & ~n25926;
  assign n25928 = ~pi781 & ~n25913;
  assign n25929 = ~n25927 & ~n25928;
  assign n25930 = ~pi619 & ~n25929;
  assign n25931 = pi619 & n25855;
  assign n25932 = ~pi1159 & ~n25931;
  assign n25933 = ~n25930 & n25932;
  assign n25934 = ~pi648 & ~n25828;
  assign n25935 = ~n25933 & n25934;
  assign n25936 = pi619 & ~n25929;
  assign n25937 = ~pi619 & n25855;
  assign n25938 = pi1159 & ~n25937;
  assign n25939 = ~n25936 & n25938;
  assign n25940 = pi648 & ~n25832;
  assign n25941 = ~n25939 & n25940;
  assign n25942 = pi789 & ~n25935;
  assign n25943 = ~n25941 & n25942;
  assign n25944 = ~pi789 & n25929;
  assign n25945 = n17905 & ~n25944;
  assign n25946 = ~n25943 & n25945;
  assign n25947 = ~n25882 & ~n25946;
  assign n25948 = ~n20298 & ~n25947;
  assign n25949 = n17944 & ~n25838;
  assign n25950 = n20786 & n25857;
  assign n25951 = ~n25949 & ~n25950;
  assign n25952 = ~pi629 & ~n25951;
  assign n25953 = n20790 & n25857;
  assign n25954 = n17943 & ~n25838;
  assign n25955 = ~n25953 & ~n25954;
  assign n25956 = pi629 & ~n25955;
  assign n25957 = ~n25952 & ~n25956;
  assign n25958 = pi792 & ~n25957;
  assign n25959 = n20300 & ~n25958;
  assign n25960 = ~n25948 & n25959;
  assign n25961 = ~n25870 & ~n25960;
  assign n25962 = pi644 & n25961;
  assign n25963 = ~pi787 & ~n25858;
  assign n25964 = pi787 & ~n25867;
  assign n25965 = ~n25963 & ~n25964;
  assign n25966 = ~pi644 & n25965;
  assign n25967 = pi715 & ~n25966;
  assign n25968 = ~n25962 & n25967;
  assign n25969 = ~n17740 & ~n25841;
  assign n25970 = n17740 & n25804;
  assign n25971 = ~n25969 & ~n25970;
  assign n25972 = pi644 & ~n25971;
  assign n25973 = ~pi644 & n25804;
  assign n25974 = ~pi715 & ~n25973;
  assign n25975 = ~n25972 & n25974;
  assign n25976 = pi1160 & ~n25975;
  assign n25977 = ~n25968 & n25976;
  assign n25978 = ~pi644 & n25961;
  assign n25979 = pi644 & n25965;
  assign n25980 = ~pi715 & ~n25979;
  assign n25981 = ~n25978 & n25980;
  assign n25982 = ~pi644 & ~n25971;
  assign n25983 = pi644 & n25804;
  assign n25984 = pi715 & ~n25983;
  assign n25985 = ~n25982 & n25984;
  assign n25986 = ~pi1160 & ~n25985;
  assign n25987 = ~n25981 & n25986;
  assign n25988 = ~n25977 & ~n25987;
  assign n25989 = pi790 & ~n25988;
  assign n25990 = ~pi790 & n25961;
  assign n25991 = pi832 & ~n25990;
  assign n25992 = ~n25989 & n25991;
  assign po336 = ~n25803 & ~n25992;
  assign n25994 = ~pi180 & ~n2755;
  assign n25995 = ~pi753 & n16933;
  assign n25996 = ~n25994 & ~n25995;
  assign n25997 = ~n17794 & ~n25996;
  assign n25998 = ~pi785 & ~n25997;
  assign n25999 = n17539 & n25995;
  assign n26000 = n25997 & ~n25999;
  assign n26001 = pi1155 & ~n26000;
  assign n26002 = ~pi1155 & ~n25994;
  assign n26003 = ~n25999 & n26002;
  assign n26004 = ~n26001 & ~n26003;
  assign n26005 = pi785 & ~n26004;
  assign n26006 = ~n25998 & ~n26005;
  assign n26007 = ~pi781 & ~n26006;
  assign n26008 = ~n17809 & n26006;
  assign n26009 = pi1154 & ~n26008;
  assign n26010 = ~n17812 & n26006;
  assign n26011 = ~pi1154 & ~n26010;
  assign n26012 = ~n26009 & ~n26011;
  assign n26013 = pi781 & ~n26012;
  assign n26014 = ~n26007 & ~n26013;
  assign n26015 = ~pi789 & ~n26014;
  assign n26016 = ~n22988 & n26014;
  assign n26017 = pi1159 & ~n26016;
  assign n26018 = ~n22991 & n26014;
  assign n26019 = ~pi1159 & ~n26018;
  assign n26020 = ~n26017 & ~n26019;
  assign n26021 = pi789 & ~n26020;
  assign n26022 = ~n26015 & ~n26021;
  assign n26023 = ~n17904 & n26022;
  assign n26024 = n17904 & n25994;
  assign n26025 = ~n26023 & ~n26024;
  assign n26026 = ~n17698 & ~n26025;
  assign n26027 = n17698 & n25994;
  assign n26028 = ~n26026 & ~n26027;
  assign n26029 = ~n20491 & n26028;
  assign n26030 = ~pi702 & n17153;
  assign n26031 = ~n25994 & ~n26030;
  assign n26032 = ~pi778 & ~n26031;
  assign n26033 = ~pi625 & n26030;
  assign n26034 = ~n26031 & ~n26033;
  assign n26035 = pi1153 & ~n26034;
  assign n26036 = ~pi1153 & ~n25994;
  assign n26037 = ~n26033 & n26036;
  assign n26038 = pi778 & ~n26037;
  assign n26039 = ~n26035 & n26038;
  assign n26040 = ~n26032 & ~n26039;
  assign n26041 = ~n17780 & ~n26040;
  assign n26042 = ~n17782 & n26041;
  assign n26043 = ~n17784 & n26042;
  assign n26044 = ~n17916 & n26043;
  assign n26045 = ~n17947 & n26044;
  assign n26046 = ~pi647 & n26045;
  assign n26047 = pi647 & n25994;
  assign n26048 = ~pi1157 & ~n26047;
  assign n26049 = ~n26046 & n26048;
  assign n26050 = pi647 & ~n26045;
  assign n26051 = ~pi647 & ~n25994;
  assign n26052 = ~n26050 & ~n26051;
  assign n26053 = pi1157 & ~n26052;
  assign n26054 = ~n26049 & ~n26053;
  assign n26055 = ~n17739 & ~n26054;
  assign n26056 = ~n26029 & ~n26055;
  assign n26057 = pi787 & ~n26056;
  assign n26058 = ~pi626 & ~n26022;
  assign n26059 = pi626 & ~n25994;
  assign n26060 = n17668 & ~n26059;
  assign n26061 = ~n26058 & n26060;
  assign n26062 = pi626 & ~n26022;
  assign n26063 = ~pi626 & ~n25994;
  assign n26064 = n17667 & ~n26063;
  assign n26065 = ~n26062 & n26064;
  assign n26066 = n17792 & n26043;
  assign n26067 = ~n26061 & ~n26066;
  assign n26068 = ~n26065 & n26067;
  assign n26069 = pi788 & ~n26068;
  assign n26070 = ~n16842 & ~n26031;
  assign n26071 = pi625 & n26070;
  assign n26072 = n25996 & ~n26070;
  assign n26073 = ~n26071 & ~n26072;
  assign n26074 = n26036 & ~n26073;
  assign n26075 = ~pi608 & ~n26035;
  assign n26076 = ~n26074 & n26075;
  assign n26077 = pi1153 & n25996;
  assign n26078 = ~n26071 & n26077;
  assign n26079 = pi608 & ~n26037;
  assign n26080 = ~n26078 & n26079;
  assign n26081 = ~n26076 & ~n26080;
  assign n26082 = pi778 & ~n26081;
  assign n26083 = ~pi778 & ~n26072;
  assign n26084 = ~n26082 & ~n26083;
  assign n26085 = ~pi609 & ~n26084;
  assign n26086 = pi609 & ~n26040;
  assign n26087 = ~pi1155 & ~n26086;
  assign n26088 = ~n26085 & n26087;
  assign n26089 = ~pi660 & ~n26001;
  assign n26090 = ~n26088 & n26089;
  assign n26091 = pi609 & ~n26084;
  assign n26092 = ~pi609 & ~n26040;
  assign n26093 = pi1155 & ~n26092;
  assign n26094 = ~n26091 & n26093;
  assign n26095 = pi660 & ~n26003;
  assign n26096 = ~n26094 & n26095;
  assign n26097 = ~n26090 & ~n26096;
  assign n26098 = pi785 & ~n26097;
  assign n26099 = ~pi785 & ~n26084;
  assign n26100 = ~n26098 & ~n26099;
  assign n26101 = ~pi618 & ~n26100;
  assign n26102 = pi618 & n26041;
  assign n26103 = ~pi1154 & ~n26102;
  assign n26104 = ~n26101 & n26103;
  assign n26105 = ~pi627 & ~n26009;
  assign n26106 = ~n26104 & n26105;
  assign n26107 = pi618 & ~n26100;
  assign n26108 = ~pi618 & n26041;
  assign n26109 = pi1154 & ~n26108;
  assign n26110 = ~n26107 & n26109;
  assign n26111 = pi627 & ~n26011;
  assign n26112 = ~n26110 & n26111;
  assign n26113 = ~n26106 & ~n26112;
  assign n26114 = pi781 & ~n26113;
  assign n26115 = ~pi781 & ~n26100;
  assign n26116 = ~n26114 & ~n26115;
  assign n26117 = ~pi619 & ~n26116;
  assign n26118 = pi619 & n26042;
  assign n26119 = ~pi1159 & ~n26118;
  assign n26120 = ~n26117 & n26119;
  assign n26121 = ~pi648 & ~n26017;
  assign n26122 = ~n26120 & n26121;
  assign n26123 = pi619 & ~n26116;
  assign n26124 = ~pi619 & n26042;
  assign n26125 = pi1159 & ~n26124;
  assign n26126 = ~n26123 & n26125;
  assign n26127 = pi648 & ~n26019;
  assign n26128 = ~n26126 & n26127;
  assign n26129 = pi789 & ~n26122;
  assign n26130 = ~n26128 & n26129;
  assign n26131 = ~pi789 & n26116;
  assign n26132 = n17905 & ~n26131;
  assign n26133 = ~n26130 & n26132;
  assign n26134 = ~n26069 & ~n26133;
  assign n26135 = ~n20298 & ~n26134;
  assign n26136 = n17944 & ~n26025;
  assign n26137 = n20786 & n26044;
  assign n26138 = ~n26136 & ~n26137;
  assign n26139 = ~pi629 & ~n26138;
  assign n26140 = n20790 & n26044;
  assign n26141 = n17943 & ~n26025;
  assign n26142 = ~n26140 & ~n26141;
  assign n26143 = pi629 & ~n26142;
  assign n26144 = ~n26139 & ~n26143;
  assign n26145 = pi792 & ~n26144;
  assign n26146 = n20300 & ~n26145;
  assign n26147 = ~n26135 & n26146;
  assign n26148 = ~n26057 & ~n26147;
  assign n26149 = pi644 & n26148;
  assign n26150 = ~pi787 & ~n26045;
  assign n26151 = pi787 & ~n26054;
  assign n26152 = ~n26150 & ~n26151;
  assign n26153 = ~pi644 & n26152;
  assign n26154 = pi715 & ~n26153;
  assign n26155 = ~n26149 & n26154;
  assign n26156 = ~n17740 & ~n26028;
  assign n26157 = n17740 & n25994;
  assign n26158 = ~n26156 & ~n26157;
  assign n26159 = pi644 & ~n26158;
  assign n26160 = ~pi644 & n25994;
  assign n26161 = ~pi715 & ~n26160;
  assign n26162 = ~n26159 & n26161;
  assign n26163 = pi1160 & ~n26162;
  assign n26164 = ~n26155 & n26163;
  assign n26165 = ~pi644 & n26148;
  assign n26166 = pi644 & n26152;
  assign n26167 = ~pi715 & ~n26166;
  assign n26168 = ~n26165 & n26167;
  assign n26169 = ~pi644 & ~n26158;
  assign n26170 = pi644 & n25994;
  assign n26171 = pi715 & ~n26170;
  assign n26172 = ~n26169 & n26171;
  assign n26173 = ~pi1160 & ~n26172;
  assign n26174 = ~n26168 & n26173;
  assign n26175 = ~n26164 & ~n26174;
  assign n26176 = pi790 & ~n26175;
  assign n26177 = ~pi790 & n26148;
  assign n26178 = pi832 & ~n26177;
  assign n26179 = ~n26176 & n26178;
  assign n26180 = ~pi180 & ~n17494;
  assign n26181 = n17627 & ~n26180;
  assign n26182 = ~pi702 & n3268;
  assign n26183 = n26180 & ~n26182;
  assign n26184 = pi180 & ~n18064;
  assign n26185 = ~pi38 & ~n26184;
  assign n26186 = n3268 & ~n26185;
  assign n26187 = ~pi180 & n18060;
  assign n26188 = ~n26186 & ~n26187;
  assign n26189 = ~pi180 & ~n16968;
  assign n26190 = n17480 & ~n26189;
  assign n26191 = ~pi702 & ~n26190;
  assign n26192 = ~n26188 & n26191;
  assign n26193 = ~n26183 & ~n26192;
  assign n26194 = ~pi778 & n26193;
  assign n26195 = pi625 & ~n26193;
  assign n26196 = ~pi625 & n26180;
  assign n26197 = pi1153 & ~n26196;
  assign n26198 = ~n26195 & n26197;
  assign n26199 = ~pi625 & ~n26193;
  assign n26200 = pi625 & n26180;
  assign n26201 = ~pi1153 & ~n26200;
  assign n26202 = ~n26199 & n26201;
  assign n26203 = ~n26198 & ~n26202;
  assign n26204 = pi778 & ~n26203;
  assign n26205 = ~n26194 & ~n26204;
  assign n26206 = ~n17554 & ~n26205;
  assign n26207 = n17554 & ~n26180;
  assign n26208 = ~n26206 & ~n26207;
  assign n26209 = ~n17591 & n26208;
  assign n26210 = n17591 & n26180;
  assign n26211 = ~n26209 & ~n26210;
  assign n26212 = ~n17627 & n26211;
  assign n26213 = ~n26181 & ~n26212;
  assign n26214 = ~n17670 & n26213;
  assign n26215 = n17670 & n26180;
  assign n26216 = ~n26214 & ~n26215;
  assign n26217 = ~pi792 & n26216;
  assign n26218 = pi628 & ~n26216;
  assign n26219 = ~pi628 & n26180;
  assign n26220 = pi1156 & ~n26219;
  assign n26221 = ~n26218 & n26220;
  assign n26222 = ~pi628 & ~n26216;
  assign n26223 = pi628 & n26180;
  assign n26224 = ~pi1156 & ~n26223;
  assign n26225 = ~n26222 & n26224;
  assign n26226 = ~n26221 & ~n26225;
  assign n26227 = pi792 & ~n26226;
  assign n26228 = ~n26217 & ~n26227;
  assign n26229 = ~pi647 & ~n26228;
  assign n26230 = pi647 & ~n26180;
  assign n26231 = ~n26229 & ~n26230;
  assign n26232 = ~pi1157 & n26231;
  assign n26233 = pi647 & ~n26228;
  assign n26234 = ~pi647 & ~n26180;
  assign n26235 = ~n26233 & ~n26234;
  assign n26236 = pi1157 & n26235;
  assign n26237 = ~n26232 & ~n26236;
  assign n26238 = pi787 & ~n26237;
  assign n26239 = ~pi787 & n26228;
  assign n26240 = ~n26238 & ~n26239;
  assign n26241 = ~pi644 & ~n26240;
  assign n26242 = pi715 & ~n26241;
  assign n26243 = pi180 & ~n3268;
  assign n26244 = pi753 & n16814;
  assign n26245 = pi180 & n16961;
  assign n26246 = ~n26244 & ~n26245;
  assign n26247 = pi39 & ~n26246;
  assign n26248 = ~pi180 & ~pi753;
  assign n26249 = n16907 & n26248;
  assign n26250 = pi180 & pi753;
  assign n26251 = pi180 & ~n16918;
  assign n26252 = ~n21690 & ~n26251;
  assign n26253 = ~pi39 & ~n26252;
  assign n26254 = ~n26250 & ~n26253;
  assign n26255 = ~n26249 & n26254;
  assign n26256 = ~n26247 & n26255;
  assign n26257 = ~pi38 & ~n26256;
  assign n26258 = ~pi753 & n16970;
  assign n26259 = pi38 & ~n26189;
  assign n26260 = ~n26258 & n26259;
  assign n26261 = ~n26257 & ~n26260;
  assign n26262 = n3268 & ~n26261;
  assign n26263 = ~n26243 & ~n26262;
  assign n26264 = ~n17526 & ~n26263;
  assign n26265 = n17526 & ~n26180;
  assign n26266 = ~n26264 & ~n26265;
  assign n26267 = ~pi785 & ~n26266;
  assign n26268 = ~n17527 & ~n26180;
  assign n26269 = pi609 & n26264;
  assign n26270 = ~n26268 & ~n26269;
  assign n26271 = pi1155 & ~n26270;
  assign n26272 = ~n17539 & ~n26180;
  assign n26273 = ~pi609 & n26264;
  assign n26274 = ~n26272 & ~n26273;
  assign n26275 = ~pi1155 & ~n26274;
  assign n26276 = ~n26271 & ~n26275;
  assign n26277 = pi785 & ~n26276;
  assign n26278 = ~n26267 & ~n26277;
  assign n26279 = ~pi781 & ~n26278;
  assign n26280 = pi618 & n26278;
  assign n26281 = ~pi618 & n26180;
  assign n26282 = pi1154 & ~n26281;
  assign n26283 = ~n26280 & n26282;
  assign n26284 = ~pi618 & n26278;
  assign n26285 = pi618 & n26180;
  assign n26286 = ~pi1154 & ~n26285;
  assign n26287 = ~n26284 & n26286;
  assign n26288 = ~n26283 & ~n26287;
  assign n26289 = pi781 & ~n26288;
  assign n26290 = ~n26279 & ~n26289;
  assign n26291 = ~pi789 & ~n26290;
  assign n26292 = pi619 & n26290;
  assign n26293 = ~pi619 & n26180;
  assign n26294 = pi1159 & ~n26293;
  assign n26295 = ~n26292 & n26294;
  assign n26296 = ~pi619 & n26290;
  assign n26297 = pi619 & n26180;
  assign n26298 = ~pi1159 & ~n26297;
  assign n26299 = ~n26296 & n26298;
  assign n26300 = ~n26295 & ~n26299;
  assign n26301 = pi789 & ~n26300;
  assign n26302 = ~n26291 & ~n26301;
  assign n26303 = ~n17904 & n26302;
  assign n26304 = n17904 & n26180;
  assign n26305 = ~n26303 & ~n26304;
  assign n26306 = ~n17698 & ~n26305;
  assign n26307 = n17698 & n26180;
  assign n26308 = ~n26306 & ~n26307;
  assign n26309 = ~n17740 & ~n26308;
  assign n26310 = n17740 & n26180;
  assign n26311 = ~n26309 & ~n26310;
  assign n26312 = pi644 & ~n26311;
  assign n26313 = ~pi644 & n26180;
  assign n26314 = ~pi715 & ~n26313;
  assign n26315 = ~n26312 & n26314;
  assign n26316 = pi1160 & ~n26315;
  assign n26317 = ~n26242 & n26316;
  assign n26318 = pi644 & ~n26240;
  assign n26319 = ~pi715 & ~n26318;
  assign n26320 = ~pi644 & ~n26311;
  assign n26321 = pi644 & n26180;
  assign n26322 = pi715 & ~n26321;
  assign n26323 = ~n26320 & n26322;
  assign n26324 = ~pi1160 & ~n26323;
  assign n26325 = ~n26319 & n26324;
  assign n26326 = ~n26317 & ~n26325;
  assign n26327 = pi790 & ~n26326;
  assign n26328 = ~pi644 & n26324;
  assign n26329 = pi644 & n26316;
  assign n26330 = pi790 & ~n26328;
  assign n26331 = ~n26329 & n26330;
  assign n26332 = ~n20502 & n26305;
  assign n26333 = ~pi629 & n26221;
  assign n26334 = pi629 & n26225;
  assign n26335 = ~n26333 & ~n26334;
  assign n26336 = ~n26332 & n26335;
  assign n26337 = pi792 & ~n26336;
  assign n26338 = pi702 & n26261;
  assign n26339 = ~pi180 & n17074;
  assign n26340 = pi180 & n17166;
  assign n26341 = pi753 & ~n26340;
  assign n26342 = ~n26339 & n26341;
  assign n26343 = pi180 & n17233;
  assign n26344 = ~pi180 & ~n17295;
  assign n26345 = ~pi753 & ~n26344;
  assign n26346 = ~n26343 & n26345;
  assign n26347 = pi39 & ~n26346;
  assign n26348 = ~n26342 & n26347;
  assign n26349 = pi180 & ~n17340;
  assign n26350 = ~pi180 & ~n17317;
  assign n26351 = pi753 & ~n26349;
  assign n26352 = ~n26350 & n26351;
  assign n26353 = ~pi180 & n17344;
  assign n26354 = pi180 & n17351;
  assign n26355 = ~pi753 & ~n26354;
  assign n26356 = ~n26353 & n26355;
  assign n26357 = ~n26352 & ~n26356;
  assign n26358 = ~pi39 & ~n26357;
  assign n26359 = ~pi38 & ~n26358;
  assign n26360 = ~n26348 & n26359;
  assign n26361 = ~pi753 & ~n17259;
  assign n26362 = n19303 & ~n26361;
  assign n26363 = ~pi180 & ~n26362;
  assign n26364 = ~n17154 & ~n25995;
  assign n26365 = pi180 & ~n26364;
  assign n26366 = n6250 & n26365;
  assign n26367 = pi38 & ~n26366;
  assign n26368 = ~n26363 & n26367;
  assign n26369 = ~pi702 & ~n26368;
  assign n26370 = ~n26360 & n26369;
  assign n26371 = n3268 & ~n26370;
  assign n26372 = ~n26338 & n26371;
  assign n26373 = ~n26243 & ~n26372;
  assign n26374 = ~pi625 & n26373;
  assign n26375 = pi625 & n26263;
  assign n26376 = ~pi1153 & ~n26375;
  assign n26377 = ~n26374 & n26376;
  assign n26378 = ~pi608 & ~n26198;
  assign n26379 = ~n26377 & n26378;
  assign n26380 = pi625 & n26373;
  assign n26381 = ~pi625 & n26263;
  assign n26382 = pi1153 & ~n26381;
  assign n26383 = ~n26380 & n26382;
  assign n26384 = pi608 & ~n26202;
  assign n26385 = ~n26383 & n26384;
  assign n26386 = ~n26379 & ~n26385;
  assign n26387 = pi778 & ~n26386;
  assign n26388 = ~pi778 & n26373;
  assign n26389 = ~n26387 & ~n26388;
  assign n26390 = ~pi609 & ~n26389;
  assign n26391 = pi609 & n26205;
  assign n26392 = ~pi1155 & ~n26391;
  assign n26393 = ~n26390 & n26392;
  assign n26394 = ~pi660 & ~n26271;
  assign n26395 = ~n26393 & n26394;
  assign n26396 = pi609 & ~n26389;
  assign n26397 = ~pi609 & n26205;
  assign n26398 = pi1155 & ~n26397;
  assign n26399 = ~n26396 & n26398;
  assign n26400 = pi660 & ~n26275;
  assign n26401 = ~n26399 & n26400;
  assign n26402 = ~n26395 & ~n26401;
  assign n26403 = pi785 & ~n26402;
  assign n26404 = ~pi785 & ~n26389;
  assign n26405 = ~n26403 & ~n26404;
  assign n26406 = ~pi618 & ~n26405;
  assign n26407 = pi618 & n26208;
  assign n26408 = ~pi1154 & ~n26407;
  assign n26409 = ~n26406 & n26408;
  assign n26410 = ~pi627 & ~n26283;
  assign n26411 = ~n26409 & n26410;
  assign n26412 = pi618 & ~n26405;
  assign n26413 = ~pi618 & n26208;
  assign n26414 = pi1154 & ~n26413;
  assign n26415 = ~n26412 & n26414;
  assign n26416 = pi627 & ~n26287;
  assign n26417 = ~n26415 & n26416;
  assign n26418 = ~n26411 & ~n26417;
  assign n26419 = pi781 & ~n26418;
  assign n26420 = ~pi781 & ~n26405;
  assign n26421 = ~n26419 & ~n26420;
  assign n26422 = ~pi619 & ~n26421;
  assign n26423 = pi619 & ~n26211;
  assign n26424 = ~pi1159 & ~n26423;
  assign n26425 = ~n26422 & n26424;
  assign n26426 = ~pi648 & ~n26295;
  assign n26427 = ~n26425 & n26426;
  assign n26428 = pi619 & ~n26421;
  assign n26429 = ~pi619 & ~n26211;
  assign n26430 = pi1159 & ~n26429;
  assign n26431 = ~n26428 & n26430;
  assign n26432 = pi648 & ~n26299;
  assign n26433 = ~n26431 & n26432;
  assign n26434 = pi789 & ~n26427;
  assign n26435 = ~n26433 & n26434;
  assign n26436 = ~pi789 & n26421;
  assign n26437 = n17905 & ~n26436;
  assign n26438 = ~n26435 & n26437;
  assign n26439 = ~pi626 & ~n26302;
  assign n26440 = pi626 & ~n26180;
  assign n26441 = n17668 & ~n26440;
  assign n26442 = ~n26439 & n26441;
  assign n26443 = pi626 & ~n26302;
  assign n26444 = ~pi626 & ~n26180;
  assign n26445 = n17667 & ~n26444;
  assign n26446 = ~n26443 & n26445;
  assign n26447 = n17792 & n26213;
  assign n26448 = ~n26442 & ~n26447;
  assign n26449 = ~n26446 & n26448;
  assign n26450 = pi788 & ~n26449;
  assign n26451 = ~n20298 & ~n26450;
  assign n26452 = ~n26438 & n26451;
  assign n26453 = ~n26337 & ~n26452;
  assign n26454 = n20300 & ~n26453;
  assign n26455 = ~n20491 & n26308;
  assign n26456 = n17738 & ~n26231;
  assign n26457 = n17737 & ~n26235;
  assign n26458 = ~n26456 & ~n26457;
  assign n26459 = ~n26455 & n26458;
  assign n26460 = pi787 & ~n26459;
  assign n26461 = ~n26454 & ~n26460;
  assign n26462 = ~n26331 & n26461;
  assign n26463 = ~n26327 & ~n26462;
  assign n26464 = ~po1038 & ~n26463;
  assign n26465 = ~pi180 & po1038;
  assign n26466 = ~pi832 & ~n26465;
  assign n26467 = ~n26464 & n26466;
  assign po337 = ~n26179 & ~n26467;
  assign n26469 = ~pi181 & ~n2755;
  assign n26470 = ~pi754 & n16933;
  assign n26471 = ~n26469 & ~n26470;
  assign n26472 = ~n17794 & ~n26471;
  assign n26473 = ~pi785 & ~n26472;
  assign n26474 = n17539 & n26470;
  assign n26475 = n26472 & ~n26474;
  assign n26476 = pi1155 & ~n26475;
  assign n26477 = ~pi1155 & ~n26469;
  assign n26478 = ~n26474 & n26477;
  assign n26479 = ~n26476 & ~n26478;
  assign n26480 = pi785 & ~n26479;
  assign n26481 = ~n26473 & ~n26480;
  assign n26482 = ~pi781 & ~n26481;
  assign n26483 = ~n17809 & n26481;
  assign n26484 = pi1154 & ~n26483;
  assign n26485 = ~n17812 & n26481;
  assign n26486 = ~pi1154 & ~n26485;
  assign n26487 = ~n26484 & ~n26486;
  assign n26488 = pi781 & ~n26487;
  assign n26489 = ~n26482 & ~n26488;
  assign n26490 = ~pi789 & ~n26489;
  assign n26491 = ~n22988 & n26489;
  assign n26492 = pi1159 & ~n26491;
  assign n26493 = ~n22991 & n26489;
  assign n26494 = ~pi1159 & ~n26493;
  assign n26495 = ~n26492 & ~n26494;
  assign n26496 = pi789 & ~n26495;
  assign n26497 = ~n26490 & ~n26496;
  assign n26498 = ~n17904 & n26497;
  assign n26499 = n17904 & n26469;
  assign n26500 = ~n26498 & ~n26499;
  assign n26501 = ~n17698 & ~n26500;
  assign n26502 = n17698 & n26469;
  assign n26503 = ~n26501 & ~n26502;
  assign n26504 = ~n20491 & n26503;
  assign n26505 = ~pi709 & n17153;
  assign n26506 = ~n26469 & ~n26505;
  assign n26507 = ~pi778 & ~n26506;
  assign n26508 = ~pi625 & n26505;
  assign n26509 = ~n26506 & ~n26508;
  assign n26510 = pi1153 & ~n26509;
  assign n26511 = ~pi1153 & ~n26469;
  assign n26512 = ~n26508 & n26511;
  assign n26513 = pi778 & ~n26512;
  assign n26514 = ~n26510 & n26513;
  assign n26515 = ~n26507 & ~n26514;
  assign n26516 = ~n17780 & ~n26515;
  assign n26517 = ~n17782 & n26516;
  assign n26518 = ~n17784 & n26517;
  assign n26519 = ~n17916 & n26518;
  assign n26520 = ~n17947 & n26519;
  assign n26521 = ~pi647 & n26520;
  assign n26522 = pi647 & n26469;
  assign n26523 = ~pi1157 & ~n26522;
  assign n26524 = ~n26521 & n26523;
  assign n26525 = pi647 & ~n26520;
  assign n26526 = ~pi647 & ~n26469;
  assign n26527 = ~n26525 & ~n26526;
  assign n26528 = pi1157 & ~n26527;
  assign n26529 = ~n26524 & ~n26528;
  assign n26530 = ~n17739 & ~n26529;
  assign n26531 = ~n26504 & ~n26530;
  assign n26532 = pi787 & ~n26531;
  assign n26533 = ~pi626 & ~n26497;
  assign n26534 = pi626 & ~n26469;
  assign n26535 = n17668 & ~n26534;
  assign n26536 = ~n26533 & n26535;
  assign n26537 = pi626 & ~n26497;
  assign n26538 = ~pi626 & ~n26469;
  assign n26539 = n17667 & ~n26538;
  assign n26540 = ~n26537 & n26539;
  assign n26541 = n17792 & n26518;
  assign n26542 = ~n26536 & ~n26541;
  assign n26543 = ~n26540 & n26542;
  assign n26544 = pi788 & ~n26543;
  assign n26545 = ~n16842 & ~n26506;
  assign n26546 = pi625 & n26545;
  assign n26547 = n26471 & ~n26545;
  assign n26548 = ~n26546 & ~n26547;
  assign n26549 = n26511 & ~n26548;
  assign n26550 = ~pi608 & ~n26510;
  assign n26551 = ~n26549 & n26550;
  assign n26552 = pi1153 & n26471;
  assign n26553 = ~n26546 & n26552;
  assign n26554 = pi608 & ~n26512;
  assign n26555 = ~n26553 & n26554;
  assign n26556 = ~n26551 & ~n26555;
  assign n26557 = pi778 & ~n26556;
  assign n26558 = ~pi778 & ~n26547;
  assign n26559 = ~n26557 & ~n26558;
  assign n26560 = ~pi609 & ~n26559;
  assign n26561 = pi609 & ~n26515;
  assign n26562 = ~pi1155 & ~n26561;
  assign n26563 = ~n26560 & n26562;
  assign n26564 = ~pi660 & ~n26476;
  assign n26565 = ~n26563 & n26564;
  assign n26566 = pi609 & ~n26559;
  assign n26567 = ~pi609 & ~n26515;
  assign n26568 = pi1155 & ~n26567;
  assign n26569 = ~n26566 & n26568;
  assign n26570 = pi660 & ~n26478;
  assign n26571 = ~n26569 & n26570;
  assign n26572 = ~n26565 & ~n26571;
  assign n26573 = pi785 & ~n26572;
  assign n26574 = ~pi785 & ~n26559;
  assign n26575 = ~n26573 & ~n26574;
  assign n26576 = ~pi618 & ~n26575;
  assign n26577 = pi618 & n26516;
  assign n26578 = ~pi1154 & ~n26577;
  assign n26579 = ~n26576 & n26578;
  assign n26580 = ~pi627 & ~n26484;
  assign n26581 = ~n26579 & n26580;
  assign n26582 = pi618 & ~n26575;
  assign n26583 = ~pi618 & n26516;
  assign n26584 = pi1154 & ~n26583;
  assign n26585 = ~n26582 & n26584;
  assign n26586 = pi627 & ~n26486;
  assign n26587 = ~n26585 & n26586;
  assign n26588 = ~n26581 & ~n26587;
  assign n26589 = pi781 & ~n26588;
  assign n26590 = ~pi781 & ~n26575;
  assign n26591 = ~n26589 & ~n26590;
  assign n26592 = ~pi619 & ~n26591;
  assign n26593 = pi619 & n26517;
  assign n26594 = ~pi1159 & ~n26593;
  assign n26595 = ~n26592 & n26594;
  assign n26596 = ~pi648 & ~n26492;
  assign n26597 = ~n26595 & n26596;
  assign n26598 = pi619 & ~n26591;
  assign n26599 = ~pi619 & n26517;
  assign n26600 = pi1159 & ~n26599;
  assign n26601 = ~n26598 & n26600;
  assign n26602 = pi648 & ~n26494;
  assign n26603 = ~n26601 & n26602;
  assign n26604 = pi789 & ~n26597;
  assign n26605 = ~n26603 & n26604;
  assign n26606 = ~pi789 & n26591;
  assign n26607 = n17905 & ~n26606;
  assign n26608 = ~n26605 & n26607;
  assign n26609 = ~n26544 & ~n26608;
  assign n26610 = ~n20298 & ~n26609;
  assign n26611 = n17944 & ~n26500;
  assign n26612 = n20786 & n26519;
  assign n26613 = ~n26611 & ~n26612;
  assign n26614 = ~pi629 & ~n26613;
  assign n26615 = n20790 & n26519;
  assign n26616 = n17943 & ~n26500;
  assign n26617 = ~n26615 & ~n26616;
  assign n26618 = pi629 & ~n26617;
  assign n26619 = ~n26614 & ~n26618;
  assign n26620 = pi792 & ~n26619;
  assign n26621 = n20300 & ~n26620;
  assign n26622 = ~n26610 & n26621;
  assign n26623 = ~n26532 & ~n26622;
  assign n26624 = pi644 & n26623;
  assign n26625 = ~pi787 & ~n26520;
  assign n26626 = pi787 & ~n26529;
  assign n26627 = ~n26625 & ~n26626;
  assign n26628 = ~pi644 & n26627;
  assign n26629 = pi715 & ~n26628;
  assign n26630 = ~n26624 & n26629;
  assign n26631 = ~n17740 & ~n26503;
  assign n26632 = n17740 & n26469;
  assign n26633 = ~n26631 & ~n26632;
  assign n26634 = pi644 & ~n26633;
  assign n26635 = ~pi644 & n26469;
  assign n26636 = ~pi715 & ~n26635;
  assign n26637 = ~n26634 & n26636;
  assign n26638 = pi1160 & ~n26637;
  assign n26639 = ~n26630 & n26638;
  assign n26640 = ~pi644 & n26623;
  assign n26641 = pi644 & n26627;
  assign n26642 = ~pi715 & ~n26641;
  assign n26643 = ~n26640 & n26642;
  assign n26644 = ~pi644 & ~n26633;
  assign n26645 = pi644 & n26469;
  assign n26646 = pi715 & ~n26645;
  assign n26647 = ~n26644 & n26646;
  assign n26648 = ~pi1160 & ~n26647;
  assign n26649 = ~n26643 & n26648;
  assign n26650 = ~n26639 & ~n26649;
  assign n26651 = pi790 & ~n26650;
  assign n26652 = ~pi790 & n26623;
  assign n26653 = pi832 & ~n26652;
  assign n26654 = ~n26651 & n26653;
  assign n26655 = ~pi181 & ~n17494;
  assign n26656 = n17627 & ~n26655;
  assign n26657 = ~pi709 & n3268;
  assign n26658 = n26655 & ~n26657;
  assign n26659 = pi181 & ~n18064;
  assign n26660 = ~pi38 & ~n26659;
  assign n26661 = n3268 & ~n26660;
  assign n26662 = ~pi181 & n18060;
  assign n26663 = ~n26661 & ~n26662;
  assign n26664 = ~pi181 & ~n16968;
  assign n26665 = n17480 & ~n26664;
  assign n26666 = ~pi709 & ~n26665;
  assign n26667 = ~n26663 & n26666;
  assign n26668 = ~n26658 & ~n26667;
  assign n26669 = ~pi778 & n26668;
  assign n26670 = pi625 & ~n26668;
  assign n26671 = ~pi625 & n26655;
  assign n26672 = pi1153 & ~n26671;
  assign n26673 = ~n26670 & n26672;
  assign n26674 = ~pi625 & ~n26668;
  assign n26675 = pi625 & n26655;
  assign n26676 = ~pi1153 & ~n26675;
  assign n26677 = ~n26674 & n26676;
  assign n26678 = ~n26673 & ~n26677;
  assign n26679 = pi778 & ~n26678;
  assign n26680 = ~n26669 & ~n26679;
  assign n26681 = ~n17554 & ~n26680;
  assign n26682 = n17554 & ~n26655;
  assign n26683 = ~n26681 & ~n26682;
  assign n26684 = ~n17591 & n26683;
  assign n26685 = n17591 & n26655;
  assign n26686 = ~n26684 & ~n26685;
  assign n26687 = ~n17627 & n26686;
  assign n26688 = ~n26656 & ~n26687;
  assign n26689 = ~n17670 & n26688;
  assign n26690 = n17670 & n26655;
  assign n26691 = ~n26689 & ~n26690;
  assign n26692 = ~pi792 & n26691;
  assign n26693 = pi628 & ~n26691;
  assign n26694 = ~pi628 & n26655;
  assign n26695 = pi1156 & ~n26694;
  assign n26696 = ~n26693 & n26695;
  assign n26697 = ~pi628 & ~n26691;
  assign n26698 = pi628 & n26655;
  assign n26699 = ~pi1156 & ~n26698;
  assign n26700 = ~n26697 & n26699;
  assign n26701 = ~n26696 & ~n26700;
  assign n26702 = pi792 & ~n26701;
  assign n26703 = ~n26692 & ~n26702;
  assign n26704 = ~pi647 & ~n26703;
  assign n26705 = pi647 & ~n26655;
  assign n26706 = ~n26704 & ~n26705;
  assign n26707 = ~pi1157 & n26706;
  assign n26708 = pi647 & ~n26703;
  assign n26709 = ~pi647 & ~n26655;
  assign n26710 = ~n26708 & ~n26709;
  assign n26711 = pi1157 & n26710;
  assign n26712 = ~n26707 & ~n26711;
  assign n26713 = pi787 & ~n26712;
  assign n26714 = ~pi787 & n26703;
  assign n26715 = ~n26713 & ~n26714;
  assign n26716 = ~pi644 & ~n26715;
  assign n26717 = pi715 & ~n26716;
  assign n26718 = pi181 & ~n3268;
  assign n26719 = pi754 & n16814;
  assign n26720 = pi181 & n16961;
  assign n26721 = ~n26719 & ~n26720;
  assign n26722 = pi39 & ~n26721;
  assign n26723 = ~pi181 & ~pi754;
  assign n26724 = n16907 & n26723;
  assign n26725 = pi181 & pi754;
  assign n26726 = pi181 & ~n16918;
  assign n26727 = ~n21746 & ~n26726;
  assign n26728 = ~pi39 & ~n26727;
  assign n26729 = ~n26725 & ~n26728;
  assign n26730 = ~n26724 & n26729;
  assign n26731 = ~n26722 & n26730;
  assign n26732 = ~pi38 & ~n26731;
  assign n26733 = ~pi754 & n16970;
  assign n26734 = pi38 & ~n26664;
  assign n26735 = ~n26733 & n26734;
  assign n26736 = ~n26732 & ~n26735;
  assign n26737 = n3268 & ~n26736;
  assign n26738 = ~n26718 & ~n26737;
  assign n26739 = ~n17526 & ~n26738;
  assign n26740 = n17526 & ~n26655;
  assign n26741 = ~n26739 & ~n26740;
  assign n26742 = ~pi785 & ~n26741;
  assign n26743 = ~n17527 & ~n26655;
  assign n26744 = pi609 & n26739;
  assign n26745 = ~n26743 & ~n26744;
  assign n26746 = pi1155 & ~n26745;
  assign n26747 = ~n17539 & ~n26655;
  assign n26748 = ~pi609 & n26739;
  assign n26749 = ~n26747 & ~n26748;
  assign n26750 = ~pi1155 & ~n26749;
  assign n26751 = ~n26746 & ~n26750;
  assign n26752 = pi785 & ~n26751;
  assign n26753 = ~n26742 & ~n26752;
  assign n26754 = ~pi781 & ~n26753;
  assign n26755 = pi618 & n26753;
  assign n26756 = ~pi618 & n26655;
  assign n26757 = pi1154 & ~n26756;
  assign n26758 = ~n26755 & n26757;
  assign n26759 = ~pi618 & n26753;
  assign n26760 = pi618 & n26655;
  assign n26761 = ~pi1154 & ~n26760;
  assign n26762 = ~n26759 & n26761;
  assign n26763 = ~n26758 & ~n26762;
  assign n26764 = pi781 & ~n26763;
  assign n26765 = ~n26754 & ~n26764;
  assign n26766 = ~pi789 & ~n26765;
  assign n26767 = pi619 & n26765;
  assign n26768 = ~pi619 & n26655;
  assign n26769 = pi1159 & ~n26768;
  assign n26770 = ~n26767 & n26769;
  assign n26771 = ~pi619 & n26765;
  assign n26772 = pi619 & n26655;
  assign n26773 = ~pi1159 & ~n26772;
  assign n26774 = ~n26771 & n26773;
  assign n26775 = ~n26770 & ~n26774;
  assign n26776 = pi789 & ~n26775;
  assign n26777 = ~n26766 & ~n26776;
  assign n26778 = ~n17904 & n26777;
  assign n26779 = n17904 & n26655;
  assign n26780 = ~n26778 & ~n26779;
  assign n26781 = ~n17698 & ~n26780;
  assign n26782 = n17698 & n26655;
  assign n26783 = ~n26781 & ~n26782;
  assign n26784 = ~n17740 & ~n26783;
  assign n26785 = n17740 & n26655;
  assign n26786 = ~n26784 & ~n26785;
  assign n26787 = pi644 & ~n26786;
  assign n26788 = ~pi644 & n26655;
  assign n26789 = ~pi715 & ~n26788;
  assign n26790 = ~n26787 & n26789;
  assign n26791 = pi1160 & ~n26790;
  assign n26792 = ~n26717 & n26791;
  assign n26793 = pi644 & ~n26715;
  assign n26794 = ~pi715 & ~n26793;
  assign n26795 = ~pi644 & ~n26786;
  assign n26796 = pi644 & n26655;
  assign n26797 = pi715 & ~n26796;
  assign n26798 = ~n26795 & n26797;
  assign n26799 = ~pi1160 & ~n26798;
  assign n26800 = ~n26794 & n26799;
  assign n26801 = ~n26792 & ~n26800;
  assign n26802 = pi790 & ~n26801;
  assign n26803 = ~pi644 & n26799;
  assign n26804 = pi644 & n26791;
  assign n26805 = pi790 & ~n26803;
  assign n26806 = ~n26804 & n26805;
  assign n26807 = ~n20502 & n26780;
  assign n26808 = ~pi629 & n26696;
  assign n26809 = pi629 & n26700;
  assign n26810 = ~n26808 & ~n26809;
  assign n26811 = ~n26807 & n26810;
  assign n26812 = pi792 & ~n26811;
  assign n26813 = pi709 & n26736;
  assign n26814 = ~pi181 & n17074;
  assign n26815 = pi181 & n17166;
  assign n26816 = pi754 & ~n26815;
  assign n26817 = ~n26814 & n26816;
  assign n26818 = pi181 & n17233;
  assign n26819 = ~pi181 & ~n17295;
  assign n26820 = ~pi754 & ~n26819;
  assign n26821 = ~n26818 & n26820;
  assign n26822 = pi39 & ~n26821;
  assign n26823 = ~n26817 & n26822;
  assign n26824 = pi181 & ~n17340;
  assign n26825 = ~pi181 & ~n17317;
  assign n26826 = pi754 & ~n26824;
  assign n26827 = ~n26825 & n26826;
  assign n26828 = ~pi181 & n17344;
  assign n26829 = pi181 & n17351;
  assign n26830 = ~pi754 & ~n26829;
  assign n26831 = ~n26828 & n26830;
  assign n26832 = ~n26827 & ~n26831;
  assign n26833 = ~pi39 & ~n26832;
  assign n26834 = ~pi38 & ~n26833;
  assign n26835 = ~n26823 & n26834;
  assign n26836 = ~pi754 & ~n17259;
  assign n26837 = n19303 & ~n26836;
  assign n26838 = ~pi181 & ~n26837;
  assign n26839 = ~n17154 & ~n26470;
  assign n26840 = pi181 & ~n26839;
  assign n26841 = n6250 & n26840;
  assign n26842 = pi38 & ~n26841;
  assign n26843 = ~n26838 & n26842;
  assign n26844 = ~pi709 & ~n26843;
  assign n26845 = ~n26835 & n26844;
  assign n26846 = n3268 & ~n26845;
  assign n26847 = ~n26813 & n26846;
  assign n26848 = ~n26718 & ~n26847;
  assign n26849 = ~pi625 & n26848;
  assign n26850 = pi625 & n26738;
  assign n26851 = ~pi1153 & ~n26850;
  assign n26852 = ~n26849 & n26851;
  assign n26853 = ~pi608 & ~n26673;
  assign n26854 = ~n26852 & n26853;
  assign n26855 = pi625 & n26848;
  assign n26856 = ~pi625 & n26738;
  assign n26857 = pi1153 & ~n26856;
  assign n26858 = ~n26855 & n26857;
  assign n26859 = pi608 & ~n26677;
  assign n26860 = ~n26858 & n26859;
  assign n26861 = ~n26854 & ~n26860;
  assign n26862 = pi778 & ~n26861;
  assign n26863 = ~pi778 & n26848;
  assign n26864 = ~n26862 & ~n26863;
  assign n26865 = ~pi609 & ~n26864;
  assign n26866 = pi609 & n26680;
  assign n26867 = ~pi1155 & ~n26866;
  assign n26868 = ~n26865 & n26867;
  assign n26869 = ~pi660 & ~n26746;
  assign n26870 = ~n26868 & n26869;
  assign n26871 = pi609 & ~n26864;
  assign n26872 = ~pi609 & n26680;
  assign n26873 = pi1155 & ~n26872;
  assign n26874 = ~n26871 & n26873;
  assign n26875 = pi660 & ~n26750;
  assign n26876 = ~n26874 & n26875;
  assign n26877 = ~n26870 & ~n26876;
  assign n26878 = pi785 & ~n26877;
  assign n26879 = ~pi785 & ~n26864;
  assign n26880 = ~n26878 & ~n26879;
  assign n26881 = ~pi618 & ~n26880;
  assign n26882 = pi618 & n26683;
  assign n26883 = ~pi1154 & ~n26882;
  assign n26884 = ~n26881 & n26883;
  assign n26885 = ~pi627 & ~n26758;
  assign n26886 = ~n26884 & n26885;
  assign n26887 = pi618 & ~n26880;
  assign n26888 = ~pi618 & n26683;
  assign n26889 = pi1154 & ~n26888;
  assign n26890 = ~n26887 & n26889;
  assign n26891 = pi627 & ~n26762;
  assign n26892 = ~n26890 & n26891;
  assign n26893 = ~n26886 & ~n26892;
  assign n26894 = pi781 & ~n26893;
  assign n26895 = ~pi781 & ~n26880;
  assign n26896 = ~n26894 & ~n26895;
  assign n26897 = ~pi619 & ~n26896;
  assign n26898 = pi619 & ~n26686;
  assign n26899 = ~pi1159 & ~n26898;
  assign n26900 = ~n26897 & n26899;
  assign n26901 = ~pi648 & ~n26770;
  assign n26902 = ~n26900 & n26901;
  assign n26903 = pi619 & ~n26896;
  assign n26904 = ~pi619 & ~n26686;
  assign n26905 = pi1159 & ~n26904;
  assign n26906 = ~n26903 & n26905;
  assign n26907 = pi648 & ~n26774;
  assign n26908 = ~n26906 & n26907;
  assign n26909 = pi789 & ~n26902;
  assign n26910 = ~n26908 & n26909;
  assign n26911 = ~pi789 & n26896;
  assign n26912 = n17905 & ~n26911;
  assign n26913 = ~n26910 & n26912;
  assign n26914 = ~pi626 & ~n26777;
  assign n26915 = pi626 & ~n26655;
  assign n26916 = n17668 & ~n26915;
  assign n26917 = ~n26914 & n26916;
  assign n26918 = pi626 & ~n26777;
  assign n26919 = ~pi626 & ~n26655;
  assign n26920 = n17667 & ~n26919;
  assign n26921 = ~n26918 & n26920;
  assign n26922 = n17792 & n26688;
  assign n26923 = ~n26917 & ~n26922;
  assign n26924 = ~n26921 & n26923;
  assign n26925 = pi788 & ~n26924;
  assign n26926 = ~n20298 & ~n26925;
  assign n26927 = ~n26913 & n26926;
  assign n26928 = ~n26812 & ~n26927;
  assign n26929 = n20300 & ~n26928;
  assign n26930 = ~n20491 & n26783;
  assign n26931 = n17738 & ~n26706;
  assign n26932 = n17737 & ~n26710;
  assign n26933 = ~n26931 & ~n26932;
  assign n26934 = ~n26930 & n26933;
  assign n26935 = pi787 & ~n26934;
  assign n26936 = ~n26929 & ~n26935;
  assign n26937 = ~n26806 & n26936;
  assign n26938 = ~n26802 & ~n26937;
  assign n26939 = ~po1038 & ~n26938;
  assign n26940 = ~pi181 & po1038;
  assign n26941 = ~pi832 & ~n26940;
  assign n26942 = ~n26939 & n26941;
  assign po338 = ~n26654 & ~n26942;
  assign n26944 = ~pi182 & ~n2755;
  assign n26945 = ~pi756 & n16933;
  assign n26946 = ~n26944 & ~n26945;
  assign n26947 = ~n17794 & ~n26946;
  assign n26948 = ~pi785 & ~n26947;
  assign n26949 = n17539 & n26945;
  assign n26950 = n26947 & ~n26949;
  assign n26951 = pi1155 & ~n26950;
  assign n26952 = ~pi1155 & ~n26944;
  assign n26953 = ~n26949 & n26952;
  assign n26954 = ~n26951 & ~n26953;
  assign n26955 = pi785 & ~n26954;
  assign n26956 = ~n26948 & ~n26955;
  assign n26957 = ~pi781 & ~n26956;
  assign n26958 = ~n17809 & n26956;
  assign n26959 = pi1154 & ~n26958;
  assign n26960 = ~n17812 & n26956;
  assign n26961 = ~pi1154 & ~n26960;
  assign n26962 = ~n26959 & ~n26961;
  assign n26963 = pi781 & ~n26962;
  assign n26964 = ~n26957 & ~n26963;
  assign n26965 = ~pi789 & ~n26964;
  assign n26966 = ~n22988 & n26964;
  assign n26967 = pi1159 & ~n26966;
  assign n26968 = ~n22991 & n26964;
  assign n26969 = ~pi1159 & ~n26968;
  assign n26970 = ~n26967 & ~n26969;
  assign n26971 = pi789 & ~n26970;
  assign n26972 = ~n26965 & ~n26971;
  assign n26973 = ~n17904 & n26972;
  assign n26974 = n17904 & n26944;
  assign n26975 = ~n26973 & ~n26974;
  assign n26976 = ~n17698 & ~n26975;
  assign n26977 = n17698 & n26944;
  assign n26978 = ~n26976 & ~n26977;
  assign n26979 = ~n20491 & n26978;
  assign n26980 = ~pi734 & n17153;
  assign n26981 = ~n26944 & ~n26980;
  assign n26982 = ~pi778 & ~n26981;
  assign n26983 = ~pi625 & n26980;
  assign n26984 = ~n26981 & ~n26983;
  assign n26985 = pi1153 & ~n26984;
  assign n26986 = ~pi1153 & ~n26944;
  assign n26987 = ~n26983 & n26986;
  assign n26988 = pi778 & ~n26987;
  assign n26989 = ~n26985 & n26988;
  assign n26990 = ~n26982 & ~n26989;
  assign n26991 = ~n17780 & ~n26990;
  assign n26992 = ~n17782 & n26991;
  assign n26993 = ~n17784 & n26992;
  assign n26994 = ~n17916 & n26993;
  assign n26995 = ~n17947 & n26994;
  assign n26996 = ~pi647 & n26995;
  assign n26997 = pi647 & n26944;
  assign n26998 = ~pi1157 & ~n26997;
  assign n26999 = ~n26996 & n26998;
  assign n27000 = pi647 & ~n26995;
  assign n27001 = ~pi647 & ~n26944;
  assign n27002 = ~n27000 & ~n27001;
  assign n27003 = pi1157 & ~n27002;
  assign n27004 = ~n26999 & ~n27003;
  assign n27005 = ~n17739 & ~n27004;
  assign n27006 = ~n26979 & ~n27005;
  assign n27007 = pi787 & ~n27006;
  assign n27008 = ~pi626 & ~n26972;
  assign n27009 = pi626 & ~n26944;
  assign n27010 = n17668 & ~n27009;
  assign n27011 = ~n27008 & n27010;
  assign n27012 = pi626 & ~n26972;
  assign n27013 = ~pi626 & ~n26944;
  assign n27014 = n17667 & ~n27013;
  assign n27015 = ~n27012 & n27014;
  assign n27016 = n17792 & n26993;
  assign n27017 = ~n27011 & ~n27016;
  assign n27018 = ~n27015 & n27017;
  assign n27019 = pi788 & ~n27018;
  assign n27020 = ~n16842 & ~n26981;
  assign n27021 = pi625 & n27020;
  assign n27022 = n26946 & ~n27020;
  assign n27023 = ~n27021 & ~n27022;
  assign n27024 = n26986 & ~n27023;
  assign n27025 = ~pi608 & ~n26985;
  assign n27026 = ~n27024 & n27025;
  assign n27027 = pi1153 & n26946;
  assign n27028 = ~n27021 & n27027;
  assign n27029 = pi608 & ~n26987;
  assign n27030 = ~n27028 & n27029;
  assign n27031 = ~n27026 & ~n27030;
  assign n27032 = pi778 & ~n27031;
  assign n27033 = ~pi778 & ~n27022;
  assign n27034 = ~n27032 & ~n27033;
  assign n27035 = ~pi609 & ~n27034;
  assign n27036 = pi609 & ~n26990;
  assign n27037 = ~pi1155 & ~n27036;
  assign n27038 = ~n27035 & n27037;
  assign n27039 = ~pi660 & ~n26951;
  assign n27040 = ~n27038 & n27039;
  assign n27041 = pi609 & ~n27034;
  assign n27042 = ~pi609 & ~n26990;
  assign n27043 = pi1155 & ~n27042;
  assign n27044 = ~n27041 & n27043;
  assign n27045 = pi660 & ~n26953;
  assign n27046 = ~n27044 & n27045;
  assign n27047 = ~n27040 & ~n27046;
  assign n27048 = pi785 & ~n27047;
  assign n27049 = ~pi785 & ~n27034;
  assign n27050 = ~n27048 & ~n27049;
  assign n27051 = ~pi618 & ~n27050;
  assign n27052 = pi618 & n26991;
  assign n27053 = ~pi1154 & ~n27052;
  assign n27054 = ~n27051 & n27053;
  assign n27055 = ~pi627 & ~n26959;
  assign n27056 = ~n27054 & n27055;
  assign n27057 = pi618 & ~n27050;
  assign n27058 = ~pi618 & n26991;
  assign n27059 = pi1154 & ~n27058;
  assign n27060 = ~n27057 & n27059;
  assign n27061 = pi627 & ~n26961;
  assign n27062 = ~n27060 & n27061;
  assign n27063 = ~n27056 & ~n27062;
  assign n27064 = pi781 & ~n27063;
  assign n27065 = ~pi781 & ~n27050;
  assign n27066 = ~n27064 & ~n27065;
  assign n27067 = ~pi619 & ~n27066;
  assign n27068 = pi619 & n26992;
  assign n27069 = ~pi1159 & ~n27068;
  assign n27070 = ~n27067 & n27069;
  assign n27071 = ~pi648 & ~n26967;
  assign n27072 = ~n27070 & n27071;
  assign n27073 = pi619 & ~n27066;
  assign n27074 = ~pi619 & n26992;
  assign n27075 = pi1159 & ~n27074;
  assign n27076 = ~n27073 & n27075;
  assign n27077 = pi648 & ~n26969;
  assign n27078 = ~n27076 & n27077;
  assign n27079 = pi789 & ~n27072;
  assign n27080 = ~n27078 & n27079;
  assign n27081 = ~pi789 & n27066;
  assign n27082 = n17905 & ~n27081;
  assign n27083 = ~n27080 & n27082;
  assign n27084 = ~n27019 & ~n27083;
  assign n27085 = ~n20298 & ~n27084;
  assign n27086 = n17944 & ~n26975;
  assign n27087 = n20786 & n26994;
  assign n27088 = ~n27086 & ~n27087;
  assign n27089 = ~pi629 & ~n27088;
  assign n27090 = n20790 & n26994;
  assign n27091 = n17943 & ~n26975;
  assign n27092 = ~n27090 & ~n27091;
  assign n27093 = pi629 & ~n27092;
  assign n27094 = ~n27089 & ~n27093;
  assign n27095 = pi792 & ~n27094;
  assign n27096 = n20300 & ~n27095;
  assign n27097 = ~n27085 & n27096;
  assign n27098 = ~n27007 & ~n27097;
  assign n27099 = pi644 & n27098;
  assign n27100 = ~pi787 & ~n26995;
  assign n27101 = pi787 & ~n27004;
  assign n27102 = ~n27100 & ~n27101;
  assign n27103 = ~pi644 & n27102;
  assign n27104 = pi715 & ~n27103;
  assign n27105 = ~n27099 & n27104;
  assign n27106 = ~n17740 & ~n26978;
  assign n27107 = n17740 & n26944;
  assign n27108 = ~n27106 & ~n27107;
  assign n27109 = pi644 & ~n27108;
  assign n27110 = ~pi644 & n26944;
  assign n27111 = ~pi715 & ~n27110;
  assign n27112 = ~n27109 & n27111;
  assign n27113 = pi1160 & ~n27112;
  assign n27114 = ~n27105 & n27113;
  assign n27115 = ~pi644 & n27098;
  assign n27116 = pi644 & n27102;
  assign n27117 = ~pi715 & ~n27116;
  assign n27118 = ~n27115 & n27117;
  assign n27119 = ~pi644 & ~n27108;
  assign n27120 = pi644 & n26944;
  assign n27121 = pi715 & ~n27120;
  assign n27122 = ~n27119 & n27121;
  assign n27123 = ~pi1160 & ~n27122;
  assign n27124 = ~n27118 & n27123;
  assign n27125 = ~n27114 & ~n27124;
  assign n27126 = pi790 & ~n27125;
  assign n27127 = ~pi790 & n27098;
  assign n27128 = pi832 & ~n27127;
  assign n27129 = ~n27126 & n27128;
  assign n27130 = ~pi182 & ~n17494;
  assign n27131 = n17627 & ~n27130;
  assign n27132 = ~pi734 & n3268;
  assign n27133 = n27130 & ~n27132;
  assign n27134 = pi182 & ~n18064;
  assign n27135 = ~pi38 & ~n27134;
  assign n27136 = n3268 & ~n27135;
  assign n27137 = ~pi182 & n18060;
  assign n27138 = ~n27136 & ~n27137;
  assign n27139 = ~pi182 & ~n16968;
  assign n27140 = n17480 & ~n27139;
  assign n27141 = ~pi734 & ~n27140;
  assign n27142 = ~n27138 & n27141;
  assign n27143 = ~n27133 & ~n27142;
  assign n27144 = ~pi778 & n27143;
  assign n27145 = pi625 & ~n27143;
  assign n27146 = ~pi625 & n27130;
  assign n27147 = pi1153 & ~n27146;
  assign n27148 = ~n27145 & n27147;
  assign n27149 = ~pi625 & ~n27143;
  assign n27150 = pi625 & n27130;
  assign n27151 = ~pi1153 & ~n27150;
  assign n27152 = ~n27149 & n27151;
  assign n27153 = ~n27148 & ~n27152;
  assign n27154 = pi778 & ~n27153;
  assign n27155 = ~n27144 & ~n27154;
  assign n27156 = ~n17554 & ~n27155;
  assign n27157 = n17554 & ~n27130;
  assign n27158 = ~n27156 & ~n27157;
  assign n27159 = ~n17591 & n27158;
  assign n27160 = n17591 & n27130;
  assign n27161 = ~n27159 & ~n27160;
  assign n27162 = ~n17627 & n27161;
  assign n27163 = ~n27131 & ~n27162;
  assign n27164 = ~n17670 & n27163;
  assign n27165 = n17670 & n27130;
  assign n27166 = ~n27164 & ~n27165;
  assign n27167 = ~pi792 & n27166;
  assign n27168 = pi628 & ~n27166;
  assign n27169 = ~pi628 & n27130;
  assign n27170 = pi1156 & ~n27169;
  assign n27171 = ~n27168 & n27170;
  assign n27172 = ~pi628 & ~n27166;
  assign n27173 = pi628 & n27130;
  assign n27174 = ~pi1156 & ~n27173;
  assign n27175 = ~n27172 & n27174;
  assign n27176 = ~n27171 & ~n27175;
  assign n27177 = pi792 & ~n27176;
  assign n27178 = ~n27167 & ~n27177;
  assign n27179 = ~pi647 & ~n27178;
  assign n27180 = pi647 & ~n27130;
  assign n27181 = ~n27179 & ~n27180;
  assign n27182 = ~pi1157 & n27181;
  assign n27183 = pi647 & ~n27178;
  assign n27184 = ~pi647 & ~n27130;
  assign n27185 = ~n27183 & ~n27184;
  assign n27186 = pi1157 & n27185;
  assign n27187 = ~n27182 & ~n27186;
  assign n27188 = pi787 & ~n27187;
  assign n27189 = ~pi787 & n27178;
  assign n27190 = ~n27188 & ~n27189;
  assign n27191 = ~pi644 & ~n27190;
  assign n27192 = pi715 & ~n27191;
  assign n27193 = pi182 & ~n3268;
  assign n27194 = ~pi756 & n16970;
  assign n27195 = ~n27139 & ~n27194;
  assign n27196 = pi38 & ~n27195;
  assign n27197 = ~pi182 & n16907;
  assign n27198 = pi182 & ~n16963;
  assign n27199 = ~pi756 & ~n27198;
  assign n27200 = ~n27197 & n27199;
  assign n27201 = ~pi182 & pi756;
  assign n27202 = ~n16816 & n27201;
  assign n27203 = ~n27200 & ~n27202;
  assign n27204 = ~pi38 & ~n27203;
  assign n27205 = ~n27196 & ~n27204;
  assign n27206 = n3268 & n27205;
  assign n27207 = ~n27193 & ~n27206;
  assign n27208 = ~n17526 & ~n27207;
  assign n27209 = n17526 & ~n27130;
  assign n27210 = ~n27208 & ~n27209;
  assign n27211 = ~pi785 & ~n27210;
  assign n27212 = ~n17527 & ~n27130;
  assign n27213 = pi609 & n27208;
  assign n27214 = ~n27212 & ~n27213;
  assign n27215 = pi1155 & ~n27214;
  assign n27216 = ~n17539 & ~n27130;
  assign n27217 = ~pi609 & n27208;
  assign n27218 = ~n27216 & ~n27217;
  assign n27219 = ~pi1155 & ~n27218;
  assign n27220 = ~n27215 & ~n27219;
  assign n27221 = pi785 & ~n27220;
  assign n27222 = ~n27211 & ~n27221;
  assign n27223 = ~pi781 & ~n27222;
  assign n27224 = pi618 & n27222;
  assign n27225 = ~pi618 & n27130;
  assign n27226 = pi1154 & ~n27225;
  assign n27227 = ~n27224 & n27226;
  assign n27228 = ~pi618 & n27222;
  assign n27229 = pi618 & n27130;
  assign n27230 = ~pi1154 & ~n27229;
  assign n27231 = ~n27228 & n27230;
  assign n27232 = ~n27227 & ~n27231;
  assign n27233 = pi781 & ~n27232;
  assign n27234 = ~n27223 & ~n27233;
  assign n27235 = ~pi789 & ~n27234;
  assign n27236 = pi619 & n27234;
  assign n27237 = ~pi619 & n27130;
  assign n27238 = pi1159 & ~n27237;
  assign n27239 = ~n27236 & n27238;
  assign n27240 = ~pi619 & n27234;
  assign n27241 = pi619 & n27130;
  assign n27242 = ~pi1159 & ~n27241;
  assign n27243 = ~n27240 & n27242;
  assign n27244 = ~n27239 & ~n27243;
  assign n27245 = pi789 & ~n27244;
  assign n27246 = ~n27235 & ~n27245;
  assign n27247 = ~n17904 & n27246;
  assign n27248 = n17904 & n27130;
  assign n27249 = ~n27247 & ~n27248;
  assign n27250 = ~n17698 & ~n27249;
  assign n27251 = n17698 & n27130;
  assign n27252 = ~n27250 & ~n27251;
  assign n27253 = ~n17740 & ~n27252;
  assign n27254 = n17740 & n27130;
  assign n27255 = ~n27253 & ~n27254;
  assign n27256 = pi644 & ~n27255;
  assign n27257 = ~pi644 & n27130;
  assign n27258 = ~pi715 & ~n27257;
  assign n27259 = ~n27256 & n27258;
  assign n27260 = pi1160 & ~n27259;
  assign n27261 = ~n27192 & n27260;
  assign n27262 = pi644 & ~n27190;
  assign n27263 = ~pi715 & ~n27262;
  assign n27264 = ~pi644 & ~n27255;
  assign n27265 = pi644 & n27130;
  assign n27266 = pi715 & ~n27265;
  assign n27267 = ~n27264 & n27266;
  assign n27268 = ~pi1160 & ~n27267;
  assign n27269 = ~n27263 & n27268;
  assign n27270 = ~n27261 & ~n27269;
  assign n27271 = pi790 & ~n27270;
  assign n27272 = ~pi644 & n27268;
  assign n27273 = pi644 & n27260;
  assign n27274 = pi790 & ~n27272;
  assign n27275 = ~n27273 & n27274;
  assign n27276 = ~n20502 & n27249;
  assign n27277 = ~pi629 & n27171;
  assign n27278 = pi629 & n27175;
  assign n27279 = ~n27277 & ~n27278;
  assign n27280 = ~n27276 & n27279;
  assign n27281 = pi792 & ~n27280;
  assign n27282 = pi734 & ~n27205;
  assign n27283 = ~pi182 & n17074;
  assign n27284 = pi182 & n17166;
  assign n27285 = pi756 & ~n27284;
  assign n27286 = ~n27283 & n27285;
  assign n27287 = pi182 & n17233;
  assign n27288 = ~pi182 & ~n17295;
  assign n27289 = ~pi756 & ~n27288;
  assign n27290 = ~n27287 & n27289;
  assign n27291 = pi39 & ~n27290;
  assign n27292 = ~n27286 & n27291;
  assign n27293 = pi182 & ~n17340;
  assign n27294 = ~pi182 & ~n17317;
  assign n27295 = pi756 & ~n27293;
  assign n27296 = ~n27294 & n27295;
  assign n27297 = ~pi182 & n17344;
  assign n27298 = pi182 & n17351;
  assign n27299 = ~pi756 & ~n27298;
  assign n27300 = ~n27297 & n27299;
  assign n27301 = ~n27296 & ~n27300;
  assign n27302 = ~pi39 & ~n27301;
  assign n27303 = ~pi38 & ~n27302;
  assign n27304 = ~n27292 & n27303;
  assign n27305 = ~pi756 & ~n17259;
  assign n27306 = n19303 & ~n27305;
  assign n27307 = ~pi182 & ~n27306;
  assign n27308 = ~n17154 & ~n26945;
  assign n27309 = pi182 & ~n27308;
  assign n27310 = n6250 & n27309;
  assign n27311 = pi38 & ~n27310;
  assign n27312 = ~n27307 & n27311;
  assign n27313 = ~pi734 & ~n27312;
  assign n27314 = ~n27304 & n27313;
  assign n27315 = n3268 & ~n27314;
  assign n27316 = ~n27282 & n27315;
  assign n27317 = ~n27193 & ~n27316;
  assign n27318 = ~pi625 & n27317;
  assign n27319 = pi625 & n27207;
  assign n27320 = ~pi1153 & ~n27319;
  assign n27321 = ~n27318 & n27320;
  assign n27322 = ~pi608 & ~n27148;
  assign n27323 = ~n27321 & n27322;
  assign n27324 = pi625 & n27317;
  assign n27325 = ~pi625 & n27207;
  assign n27326 = pi1153 & ~n27325;
  assign n27327 = ~n27324 & n27326;
  assign n27328 = pi608 & ~n27152;
  assign n27329 = ~n27327 & n27328;
  assign n27330 = ~n27323 & ~n27329;
  assign n27331 = pi778 & ~n27330;
  assign n27332 = ~pi778 & n27317;
  assign n27333 = ~n27331 & ~n27332;
  assign n27334 = ~pi609 & ~n27333;
  assign n27335 = pi609 & n27155;
  assign n27336 = ~pi1155 & ~n27335;
  assign n27337 = ~n27334 & n27336;
  assign n27338 = ~pi660 & ~n27215;
  assign n27339 = ~n27337 & n27338;
  assign n27340 = pi609 & ~n27333;
  assign n27341 = ~pi609 & n27155;
  assign n27342 = pi1155 & ~n27341;
  assign n27343 = ~n27340 & n27342;
  assign n27344 = pi660 & ~n27219;
  assign n27345 = ~n27343 & n27344;
  assign n27346 = ~n27339 & ~n27345;
  assign n27347 = pi785 & ~n27346;
  assign n27348 = ~pi785 & ~n27333;
  assign n27349 = ~n27347 & ~n27348;
  assign n27350 = ~pi618 & ~n27349;
  assign n27351 = pi618 & n27158;
  assign n27352 = ~pi1154 & ~n27351;
  assign n27353 = ~n27350 & n27352;
  assign n27354 = ~pi627 & ~n27227;
  assign n27355 = ~n27353 & n27354;
  assign n27356 = pi618 & ~n27349;
  assign n27357 = ~pi618 & n27158;
  assign n27358 = pi1154 & ~n27357;
  assign n27359 = ~n27356 & n27358;
  assign n27360 = pi627 & ~n27231;
  assign n27361 = ~n27359 & n27360;
  assign n27362 = ~n27355 & ~n27361;
  assign n27363 = pi781 & ~n27362;
  assign n27364 = ~pi781 & ~n27349;
  assign n27365 = ~n27363 & ~n27364;
  assign n27366 = ~pi619 & ~n27365;
  assign n27367 = pi619 & ~n27161;
  assign n27368 = ~pi1159 & ~n27367;
  assign n27369 = ~n27366 & n27368;
  assign n27370 = ~pi648 & ~n27239;
  assign n27371 = ~n27369 & n27370;
  assign n27372 = pi619 & ~n27365;
  assign n27373 = ~pi619 & ~n27161;
  assign n27374 = pi1159 & ~n27373;
  assign n27375 = ~n27372 & n27374;
  assign n27376 = pi648 & ~n27243;
  assign n27377 = ~n27375 & n27376;
  assign n27378 = pi789 & ~n27371;
  assign n27379 = ~n27377 & n27378;
  assign n27380 = ~pi789 & n27365;
  assign n27381 = n17905 & ~n27380;
  assign n27382 = ~n27379 & n27381;
  assign n27383 = ~pi626 & ~n27246;
  assign n27384 = pi626 & ~n27130;
  assign n27385 = n17668 & ~n27384;
  assign n27386 = ~n27383 & n27385;
  assign n27387 = pi626 & ~n27246;
  assign n27388 = ~pi626 & ~n27130;
  assign n27389 = n17667 & ~n27388;
  assign n27390 = ~n27387 & n27389;
  assign n27391 = n17792 & n27163;
  assign n27392 = ~n27386 & ~n27391;
  assign n27393 = ~n27390 & n27392;
  assign n27394 = pi788 & ~n27393;
  assign n27395 = ~n20298 & ~n27394;
  assign n27396 = ~n27382 & n27395;
  assign n27397 = ~n27281 & ~n27396;
  assign n27398 = n20300 & ~n27397;
  assign n27399 = ~n20491 & n27252;
  assign n27400 = n17738 & ~n27181;
  assign n27401 = n17737 & ~n27185;
  assign n27402 = ~n27400 & ~n27401;
  assign n27403 = ~n27399 & n27402;
  assign n27404 = pi787 & ~n27403;
  assign n27405 = ~n27398 & ~n27404;
  assign n27406 = ~n27275 & n27405;
  assign n27407 = ~n27271 & ~n27406;
  assign n27408 = ~po1038 & ~n27407;
  assign n27409 = ~pi182 & po1038;
  assign n27410 = ~pi832 & ~n27409;
  assign n27411 = ~n27408 & n27410;
  assign po339 = ~n27129 & ~n27411;
  assign n27413 = ~pi183 & ~n2755;
  assign n27414 = ~pi755 & n16933;
  assign n27415 = ~n27413 & ~n27414;
  assign n27416 = ~n17794 & ~n27415;
  assign n27417 = ~pi785 & ~n27416;
  assign n27418 = n17539 & n27414;
  assign n27419 = n27416 & ~n27418;
  assign n27420 = pi1155 & ~n27419;
  assign n27421 = ~pi1155 & ~n27413;
  assign n27422 = ~n27418 & n27421;
  assign n27423 = ~n27420 & ~n27422;
  assign n27424 = pi785 & ~n27423;
  assign n27425 = ~n27417 & ~n27424;
  assign n27426 = ~pi781 & ~n27425;
  assign n27427 = ~n17809 & n27425;
  assign n27428 = pi1154 & ~n27427;
  assign n27429 = ~n17812 & n27425;
  assign n27430 = ~pi1154 & ~n27429;
  assign n27431 = ~n27428 & ~n27430;
  assign n27432 = pi781 & ~n27431;
  assign n27433 = ~n27426 & ~n27432;
  assign n27434 = ~pi789 & ~n27433;
  assign n27435 = ~n22988 & n27433;
  assign n27436 = pi1159 & ~n27435;
  assign n27437 = ~n22991 & n27433;
  assign n27438 = ~pi1159 & ~n27437;
  assign n27439 = ~n27436 & ~n27438;
  assign n27440 = pi789 & ~n27439;
  assign n27441 = ~n27434 & ~n27440;
  assign n27442 = ~n17904 & n27441;
  assign n27443 = n17904 & n27413;
  assign n27444 = ~n27442 & ~n27443;
  assign n27445 = ~n17698 & ~n27444;
  assign n27446 = n17698 & n27413;
  assign n27447 = ~n27445 & ~n27446;
  assign n27448 = ~n20491 & n27447;
  assign n27449 = ~pi725 & n17153;
  assign n27450 = ~n27413 & ~n27449;
  assign n27451 = ~pi778 & ~n27450;
  assign n27452 = ~pi625 & n27449;
  assign n27453 = ~n27450 & ~n27452;
  assign n27454 = pi1153 & ~n27453;
  assign n27455 = ~pi1153 & ~n27413;
  assign n27456 = ~n27452 & n27455;
  assign n27457 = pi778 & ~n27456;
  assign n27458 = ~n27454 & n27457;
  assign n27459 = ~n27451 & ~n27458;
  assign n27460 = ~n17780 & ~n27459;
  assign n27461 = ~n17782 & n27460;
  assign n27462 = ~n17784 & n27461;
  assign n27463 = ~n17916 & n27462;
  assign n27464 = ~n17947 & n27463;
  assign n27465 = ~pi647 & n27464;
  assign n27466 = pi647 & n27413;
  assign n27467 = ~pi1157 & ~n27466;
  assign n27468 = ~n27465 & n27467;
  assign n27469 = pi647 & ~n27464;
  assign n27470 = ~pi647 & ~n27413;
  assign n27471 = ~n27469 & ~n27470;
  assign n27472 = pi1157 & ~n27471;
  assign n27473 = ~n27468 & ~n27472;
  assign n27474 = ~n17739 & ~n27473;
  assign n27475 = ~n27448 & ~n27474;
  assign n27476 = pi787 & ~n27475;
  assign n27477 = ~pi626 & ~n27441;
  assign n27478 = pi626 & ~n27413;
  assign n27479 = n17668 & ~n27478;
  assign n27480 = ~n27477 & n27479;
  assign n27481 = pi626 & ~n27441;
  assign n27482 = ~pi626 & ~n27413;
  assign n27483 = n17667 & ~n27482;
  assign n27484 = ~n27481 & n27483;
  assign n27485 = n17792 & n27462;
  assign n27486 = ~n27480 & ~n27485;
  assign n27487 = ~n27484 & n27486;
  assign n27488 = pi788 & ~n27487;
  assign n27489 = ~n16842 & ~n27450;
  assign n27490 = pi625 & n27489;
  assign n27491 = n27415 & ~n27489;
  assign n27492 = ~n27490 & ~n27491;
  assign n27493 = n27455 & ~n27492;
  assign n27494 = ~pi608 & ~n27454;
  assign n27495 = ~n27493 & n27494;
  assign n27496 = pi1153 & n27415;
  assign n27497 = ~n27490 & n27496;
  assign n27498 = pi608 & ~n27456;
  assign n27499 = ~n27497 & n27498;
  assign n27500 = ~n27495 & ~n27499;
  assign n27501 = pi778 & ~n27500;
  assign n27502 = ~pi778 & ~n27491;
  assign n27503 = ~n27501 & ~n27502;
  assign n27504 = ~pi609 & ~n27503;
  assign n27505 = pi609 & ~n27459;
  assign n27506 = ~pi1155 & ~n27505;
  assign n27507 = ~n27504 & n27506;
  assign n27508 = ~pi660 & ~n27420;
  assign n27509 = ~n27507 & n27508;
  assign n27510 = pi609 & ~n27503;
  assign n27511 = ~pi609 & ~n27459;
  assign n27512 = pi1155 & ~n27511;
  assign n27513 = ~n27510 & n27512;
  assign n27514 = pi660 & ~n27422;
  assign n27515 = ~n27513 & n27514;
  assign n27516 = ~n27509 & ~n27515;
  assign n27517 = pi785 & ~n27516;
  assign n27518 = ~pi785 & ~n27503;
  assign n27519 = ~n27517 & ~n27518;
  assign n27520 = ~pi618 & ~n27519;
  assign n27521 = pi618 & n27460;
  assign n27522 = ~pi1154 & ~n27521;
  assign n27523 = ~n27520 & n27522;
  assign n27524 = ~pi627 & ~n27428;
  assign n27525 = ~n27523 & n27524;
  assign n27526 = pi618 & ~n27519;
  assign n27527 = ~pi618 & n27460;
  assign n27528 = pi1154 & ~n27527;
  assign n27529 = ~n27526 & n27528;
  assign n27530 = pi627 & ~n27430;
  assign n27531 = ~n27529 & n27530;
  assign n27532 = ~n27525 & ~n27531;
  assign n27533 = pi781 & ~n27532;
  assign n27534 = ~pi781 & ~n27519;
  assign n27535 = ~n27533 & ~n27534;
  assign n27536 = ~pi619 & ~n27535;
  assign n27537 = pi619 & n27461;
  assign n27538 = ~pi1159 & ~n27537;
  assign n27539 = ~n27536 & n27538;
  assign n27540 = ~pi648 & ~n27436;
  assign n27541 = ~n27539 & n27540;
  assign n27542 = pi619 & ~n27535;
  assign n27543 = ~pi619 & n27461;
  assign n27544 = pi1159 & ~n27543;
  assign n27545 = ~n27542 & n27544;
  assign n27546 = pi648 & ~n27438;
  assign n27547 = ~n27545 & n27546;
  assign n27548 = pi789 & ~n27541;
  assign n27549 = ~n27547 & n27548;
  assign n27550 = ~pi789 & n27535;
  assign n27551 = n17905 & ~n27550;
  assign n27552 = ~n27549 & n27551;
  assign n27553 = ~n27488 & ~n27552;
  assign n27554 = ~n20298 & ~n27553;
  assign n27555 = n17944 & ~n27444;
  assign n27556 = n20786 & n27463;
  assign n27557 = ~n27555 & ~n27556;
  assign n27558 = ~pi629 & ~n27557;
  assign n27559 = n20790 & n27463;
  assign n27560 = n17943 & ~n27444;
  assign n27561 = ~n27559 & ~n27560;
  assign n27562 = pi629 & ~n27561;
  assign n27563 = ~n27558 & ~n27562;
  assign n27564 = pi792 & ~n27563;
  assign n27565 = n20300 & ~n27564;
  assign n27566 = ~n27554 & n27565;
  assign n27567 = ~n27476 & ~n27566;
  assign n27568 = pi644 & n27567;
  assign n27569 = ~pi787 & ~n27464;
  assign n27570 = pi787 & ~n27473;
  assign n27571 = ~n27569 & ~n27570;
  assign n27572 = ~pi644 & n27571;
  assign n27573 = pi715 & ~n27572;
  assign n27574 = ~n27568 & n27573;
  assign n27575 = ~n17740 & ~n27447;
  assign n27576 = n17740 & n27413;
  assign n27577 = ~n27575 & ~n27576;
  assign n27578 = pi644 & ~n27577;
  assign n27579 = ~pi644 & n27413;
  assign n27580 = ~pi715 & ~n27579;
  assign n27581 = ~n27578 & n27580;
  assign n27582 = pi1160 & ~n27581;
  assign n27583 = ~n27574 & n27582;
  assign n27584 = ~pi644 & n27567;
  assign n27585 = pi644 & n27571;
  assign n27586 = ~pi715 & ~n27585;
  assign n27587 = ~n27584 & n27586;
  assign n27588 = ~pi644 & ~n27577;
  assign n27589 = pi644 & n27413;
  assign n27590 = pi715 & ~n27589;
  assign n27591 = ~n27588 & n27590;
  assign n27592 = ~pi1160 & ~n27591;
  assign n27593 = ~n27587 & n27592;
  assign n27594 = ~n27583 & ~n27593;
  assign n27595 = pi790 & ~n27594;
  assign n27596 = ~pi790 & n27567;
  assign n27597 = pi832 & ~n27596;
  assign n27598 = ~n27595 & n27597;
  assign n27599 = ~pi183 & ~n17494;
  assign n27600 = n17627 & ~n27599;
  assign n27601 = ~pi725 & n3268;
  assign n27602 = n27599 & ~n27601;
  assign n27603 = pi183 & ~n18064;
  assign n27604 = ~pi38 & ~n27603;
  assign n27605 = n3268 & ~n27604;
  assign n27606 = ~pi183 & n18060;
  assign n27607 = ~n27605 & ~n27606;
  assign n27608 = ~pi183 & ~n16968;
  assign n27609 = n17480 & ~n27608;
  assign n27610 = ~pi725 & ~n27609;
  assign n27611 = ~n27607 & n27610;
  assign n27612 = ~n27602 & ~n27611;
  assign n27613 = ~pi778 & n27612;
  assign n27614 = pi625 & ~n27612;
  assign n27615 = ~pi625 & n27599;
  assign n27616 = pi1153 & ~n27615;
  assign n27617 = ~n27614 & n27616;
  assign n27618 = ~pi625 & ~n27612;
  assign n27619 = pi625 & n27599;
  assign n27620 = ~pi1153 & ~n27619;
  assign n27621 = ~n27618 & n27620;
  assign n27622 = ~n27617 & ~n27621;
  assign n27623 = pi778 & ~n27622;
  assign n27624 = ~n27613 & ~n27623;
  assign n27625 = ~n17554 & ~n27624;
  assign n27626 = n17554 & ~n27599;
  assign n27627 = ~n27625 & ~n27626;
  assign n27628 = ~n17591 & n27627;
  assign n27629 = n17591 & n27599;
  assign n27630 = ~n27628 & ~n27629;
  assign n27631 = ~n17627 & n27630;
  assign n27632 = ~n27600 & ~n27631;
  assign n27633 = ~n17670 & n27632;
  assign n27634 = n17670 & n27599;
  assign n27635 = ~n27633 & ~n27634;
  assign n27636 = ~pi792 & n27635;
  assign n27637 = pi628 & ~n27635;
  assign n27638 = ~pi628 & n27599;
  assign n27639 = pi1156 & ~n27638;
  assign n27640 = ~n27637 & n27639;
  assign n27641 = ~pi628 & ~n27635;
  assign n27642 = pi628 & n27599;
  assign n27643 = ~pi1156 & ~n27642;
  assign n27644 = ~n27641 & n27643;
  assign n27645 = ~n27640 & ~n27644;
  assign n27646 = pi792 & ~n27645;
  assign n27647 = ~n27636 & ~n27646;
  assign n27648 = ~pi647 & ~n27647;
  assign n27649 = pi647 & ~n27599;
  assign n27650 = ~n27648 & ~n27649;
  assign n27651 = ~pi1157 & n27650;
  assign n27652 = pi647 & ~n27647;
  assign n27653 = ~pi647 & ~n27599;
  assign n27654 = ~n27652 & ~n27653;
  assign n27655 = pi1157 & n27654;
  assign n27656 = ~n27651 & ~n27655;
  assign n27657 = pi787 & ~n27656;
  assign n27658 = ~pi787 & n27647;
  assign n27659 = ~n27657 & ~n27658;
  assign n27660 = ~pi644 & ~n27659;
  assign n27661 = pi715 & ~n27660;
  assign n27662 = pi183 & ~n3268;
  assign n27663 = ~pi755 & n16970;
  assign n27664 = ~n27608 & ~n27663;
  assign n27665 = pi38 & ~n27664;
  assign n27666 = ~pi183 & n16907;
  assign n27667 = pi183 & ~n16963;
  assign n27668 = ~pi755 & ~n27667;
  assign n27669 = ~n27666 & n27668;
  assign n27670 = ~pi183 & pi755;
  assign n27671 = ~n16816 & n27670;
  assign n27672 = ~n27669 & ~n27671;
  assign n27673 = ~pi38 & ~n27672;
  assign n27674 = ~n27665 & ~n27673;
  assign n27675 = n3268 & n27674;
  assign n27676 = ~n27662 & ~n27675;
  assign n27677 = ~n17526 & ~n27676;
  assign n27678 = n17526 & ~n27599;
  assign n27679 = ~n27677 & ~n27678;
  assign n27680 = ~pi785 & ~n27679;
  assign n27681 = ~n17527 & ~n27599;
  assign n27682 = pi609 & n27677;
  assign n27683 = ~n27681 & ~n27682;
  assign n27684 = pi1155 & ~n27683;
  assign n27685 = ~n17539 & ~n27599;
  assign n27686 = ~pi609 & n27677;
  assign n27687 = ~n27685 & ~n27686;
  assign n27688 = ~pi1155 & ~n27687;
  assign n27689 = ~n27684 & ~n27688;
  assign n27690 = pi785 & ~n27689;
  assign n27691 = ~n27680 & ~n27690;
  assign n27692 = ~pi781 & ~n27691;
  assign n27693 = pi618 & n27691;
  assign n27694 = ~pi618 & n27599;
  assign n27695 = pi1154 & ~n27694;
  assign n27696 = ~n27693 & n27695;
  assign n27697 = ~pi618 & n27691;
  assign n27698 = pi618 & n27599;
  assign n27699 = ~pi1154 & ~n27698;
  assign n27700 = ~n27697 & n27699;
  assign n27701 = ~n27696 & ~n27700;
  assign n27702 = pi781 & ~n27701;
  assign n27703 = ~n27692 & ~n27702;
  assign n27704 = ~pi789 & ~n27703;
  assign n27705 = pi619 & n27703;
  assign n27706 = ~pi619 & n27599;
  assign n27707 = pi1159 & ~n27706;
  assign n27708 = ~n27705 & n27707;
  assign n27709 = ~pi619 & n27703;
  assign n27710 = pi619 & n27599;
  assign n27711 = ~pi1159 & ~n27710;
  assign n27712 = ~n27709 & n27711;
  assign n27713 = ~n27708 & ~n27712;
  assign n27714 = pi789 & ~n27713;
  assign n27715 = ~n27704 & ~n27714;
  assign n27716 = ~n17904 & n27715;
  assign n27717 = n17904 & n27599;
  assign n27718 = ~n27716 & ~n27717;
  assign n27719 = ~n17698 & ~n27718;
  assign n27720 = n17698 & n27599;
  assign n27721 = ~n27719 & ~n27720;
  assign n27722 = ~n17740 & ~n27721;
  assign n27723 = n17740 & n27599;
  assign n27724 = ~n27722 & ~n27723;
  assign n27725 = pi644 & ~n27724;
  assign n27726 = ~pi644 & n27599;
  assign n27727 = ~pi715 & ~n27726;
  assign n27728 = ~n27725 & n27727;
  assign n27729 = pi1160 & ~n27728;
  assign n27730 = ~n27661 & n27729;
  assign n27731 = pi644 & ~n27659;
  assign n27732 = ~pi715 & ~n27731;
  assign n27733 = ~pi644 & ~n27724;
  assign n27734 = pi644 & n27599;
  assign n27735 = pi715 & ~n27734;
  assign n27736 = ~n27733 & n27735;
  assign n27737 = ~pi1160 & ~n27736;
  assign n27738 = ~n27732 & n27737;
  assign n27739 = ~n27730 & ~n27738;
  assign n27740 = pi790 & ~n27739;
  assign n27741 = ~pi644 & n27737;
  assign n27742 = pi644 & n27729;
  assign n27743 = pi790 & ~n27741;
  assign n27744 = ~n27742 & n27743;
  assign n27745 = ~n20502 & n27718;
  assign n27746 = ~pi629 & n27640;
  assign n27747 = pi629 & n27644;
  assign n27748 = ~n27746 & ~n27747;
  assign n27749 = ~n27745 & n27748;
  assign n27750 = pi792 & ~n27749;
  assign n27751 = pi725 & ~n27674;
  assign n27752 = ~pi183 & n17074;
  assign n27753 = pi183 & n17166;
  assign n27754 = pi755 & ~n27753;
  assign n27755 = ~n27752 & n27754;
  assign n27756 = pi183 & n17233;
  assign n27757 = ~pi183 & ~n17295;
  assign n27758 = ~pi755 & ~n27757;
  assign n27759 = ~n27756 & n27758;
  assign n27760 = pi39 & ~n27759;
  assign n27761 = ~n27755 & n27760;
  assign n27762 = pi183 & ~n17340;
  assign n27763 = ~pi183 & ~n17317;
  assign n27764 = pi755 & ~n27762;
  assign n27765 = ~n27763 & n27764;
  assign n27766 = ~pi183 & n17344;
  assign n27767 = pi183 & n17351;
  assign n27768 = ~pi755 & ~n27767;
  assign n27769 = ~n27766 & n27768;
  assign n27770 = ~n27765 & ~n27769;
  assign n27771 = ~pi39 & ~n27770;
  assign n27772 = ~pi38 & ~n27771;
  assign n27773 = ~n27761 & n27772;
  assign n27774 = ~pi755 & ~n17259;
  assign n27775 = n19303 & ~n27774;
  assign n27776 = ~pi183 & ~n27775;
  assign n27777 = ~n17154 & ~n27414;
  assign n27778 = pi183 & ~n27777;
  assign n27779 = n6250 & n27778;
  assign n27780 = pi38 & ~n27779;
  assign n27781 = ~n27776 & n27780;
  assign n27782 = ~pi725 & ~n27781;
  assign n27783 = ~n27773 & n27782;
  assign n27784 = n3268 & ~n27783;
  assign n27785 = ~n27751 & n27784;
  assign n27786 = ~n27662 & ~n27785;
  assign n27787 = ~pi625 & n27786;
  assign n27788 = pi625 & n27676;
  assign n27789 = ~pi1153 & ~n27788;
  assign n27790 = ~n27787 & n27789;
  assign n27791 = ~pi608 & ~n27617;
  assign n27792 = ~n27790 & n27791;
  assign n27793 = pi625 & n27786;
  assign n27794 = ~pi625 & n27676;
  assign n27795 = pi1153 & ~n27794;
  assign n27796 = ~n27793 & n27795;
  assign n27797 = pi608 & ~n27621;
  assign n27798 = ~n27796 & n27797;
  assign n27799 = ~n27792 & ~n27798;
  assign n27800 = pi778 & ~n27799;
  assign n27801 = ~pi778 & n27786;
  assign n27802 = ~n27800 & ~n27801;
  assign n27803 = ~pi609 & ~n27802;
  assign n27804 = pi609 & n27624;
  assign n27805 = ~pi1155 & ~n27804;
  assign n27806 = ~n27803 & n27805;
  assign n27807 = ~pi660 & ~n27684;
  assign n27808 = ~n27806 & n27807;
  assign n27809 = pi609 & ~n27802;
  assign n27810 = ~pi609 & n27624;
  assign n27811 = pi1155 & ~n27810;
  assign n27812 = ~n27809 & n27811;
  assign n27813 = pi660 & ~n27688;
  assign n27814 = ~n27812 & n27813;
  assign n27815 = ~n27808 & ~n27814;
  assign n27816 = pi785 & ~n27815;
  assign n27817 = ~pi785 & ~n27802;
  assign n27818 = ~n27816 & ~n27817;
  assign n27819 = ~pi618 & ~n27818;
  assign n27820 = pi618 & n27627;
  assign n27821 = ~pi1154 & ~n27820;
  assign n27822 = ~n27819 & n27821;
  assign n27823 = ~pi627 & ~n27696;
  assign n27824 = ~n27822 & n27823;
  assign n27825 = pi618 & ~n27818;
  assign n27826 = ~pi618 & n27627;
  assign n27827 = pi1154 & ~n27826;
  assign n27828 = ~n27825 & n27827;
  assign n27829 = pi627 & ~n27700;
  assign n27830 = ~n27828 & n27829;
  assign n27831 = ~n27824 & ~n27830;
  assign n27832 = pi781 & ~n27831;
  assign n27833 = ~pi781 & ~n27818;
  assign n27834 = ~n27832 & ~n27833;
  assign n27835 = ~pi619 & ~n27834;
  assign n27836 = pi619 & ~n27630;
  assign n27837 = ~pi1159 & ~n27836;
  assign n27838 = ~n27835 & n27837;
  assign n27839 = ~pi648 & ~n27708;
  assign n27840 = ~n27838 & n27839;
  assign n27841 = pi619 & ~n27834;
  assign n27842 = ~pi619 & ~n27630;
  assign n27843 = pi1159 & ~n27842;
  assign n27844 = ~n27841 & n27843;
  assign n27845 = pi648 & ~n27712;
  assign n27846 = ~n27844 & n27845;
  assign n27847 = pi789 & ~n27840;
  assign n27848 = ~n27846 & n27847;
  assign n27849 = ~pi789 & n27834;
  assign n27850 = n17905 & ~n27849;
  assign n27851 = ~n27848 & n27850;
  assign n27852 = ~pi626 & ~n27715;
  assign n27853 = pi626 & ~n27599;
  assign n27854 = n17668 & ~n27853;
  assign n27855 = ~n27852 & n27854;
  assign n27856 = pi626 & ~n27715;
  assign n27857 = ~pi626 & ~n27599;
  assign n27858 = n17667 & ~n27857;
  assign n27859 = ~n27856 & n27858;
  assign n27860 = n17792 & n27632;
  assign n27861 = ~n27855 & ~n27860;
  assign n27862 = ~n27859 & n27861;
  assign n27863 = pi788 & ~n27862;
  assign n27864 = ~n20298 & ~n27863;
  assign n27865 = ~n27851 & n27864;
  assign n27866 = ~n27750 & ~n27865;
  assign n27867 = n20300 & ~n27866;
  assign n27868 = ~n20491 & n27721;
  assign n27869 = n17738 & ~n27650;
  assign n27870 = n17737 & ~n27654;
  assign n27871 = ~n27869 & ~n27870;
  assign n27872 = ~n27868 & n27871;
  assign n27873 = pi787 & ~n27872;
  assign n27874 = ~n27867 & ~n27873;
  assign n27875 = ~n27744 & n27874;
  assign n27876 = ~n27740 & ~n27875;
  assign n27877 = ~po1038 & ~n27876;
  assign n27878 = ~pi183 & po1038;
  assign n27879 = ~pi832 & ~n27878;
  assign n27880 = ~n27877 & n27879;
  assign po340 = ~n27598 & ~n27880;
  assign n27882 = ~pi184 & ~n2755;
  assign n27883 = ~pi777 & n16933;
  assign n27884 = ~n27882 & ~n27883;
  assign n27885 = ~n17794 & ~n27884;
  assign n27886 = ~pi785 & ~n27885;
  assign n27887 = n17539 & n27883;
  assign n27888 = n27885 & ~n27887;
  assign n27889 = pi1155 & ~n27888;
  assign n27890 = ~pi1155 & ~n27882;
  assign n27891 = ~n27887 & n27890;
  assign n27892 = ~n27889 & ~n27891;
  assign n27893 = pi785 & ~n27892;
  assign n27894 = ~n27886 & ~n27893;
  assign n27895 = ~pi781 & ~n27894;
  assign n27896 = ~n17809 & n27894;
  assign n27897 = pi1154 & ~n27896;
  assign n27898 = ~n17812 & n27894;
  assign n27899 = ~pi1154 & ~n27898;
  assign n27900 = ~n27897 & ~n27899;
  assign n27901 = pi781 & ~n27900;
  assign n27902 = ~n27895 & ~n27901;
  assign n27903 = ~pi789 & ~n27902;
  assign n27904 = ~n22988 & n27902;
  assign n27905 = pi1159 & ~n27904;
  assign n27906 = ~n22991 & n27902;
  assign n27907 = ~pi1159 & ~n27906;
  assign n27908 = ~n27905 & ~n27907;
  assign n27909 = pi789 & ~n27908;
  assign n27910 = ~n27903 & ~n27909;
  assign n27911 = ~n17904 & n27910;
  assign n27912 = n17904 & n27882;
  assign n27913 = ~n27911 & ~n27912;
  assign n27914 = ~n17698 & ~n27913;
  assign n27915 = n17698 & n27882;
  assign n27916 = ~n27914 & ~n27915;
  assign n27917 = ~n20491 & n27916;
  assign n27918 = ~pi737 & n17153;
  assign n27919 = ~n27882 & ~n27918;
  assign n27920 = ~pi778 & ~n27919;
  assign n27921 = ~pi625 & n27918;
  assign n27922 = ~n27919 & ~n27921;
  assign n27923 = pi1153 & ~n27922;
  assign n27924 = ~pi1153 & ~n27882;
  assign n27925 = ~n27921 & n27924;
  assign n27926 = pi778 & ~n27925;
  assign n27927 = ~n27923 & n27926;
  assign n27928 = ~n27920 & ~n27927;
  assign n27929 = ~n17780 & ~n27928;
  assign n27930 = ~n17782 & n27929;
  assign n27931 = ~n17784 & n27930;
  assign n27932 = ~n17916 & n27931;
  assign n27933 = ~n17947 & n27932;
  assign n27934 = ~pi647 & n27933;
  assign n27935 = pi647 & n27882;
  assign n27936 = ~pi1157 & ~n27935;
  assign n27937 = ~n27934 & n27936;
  assign n27938 = pi647 & ~n27933;
  assign n27939 = ~pi647 & ~n27882;
  assign n27940 = ~n27938 & ~n27939;
  assign n27941 = pi1157 & ~n27940;
  assign n27942 = ~n27937 & ~n27941;
  assign n27943 = ~n17739 & ~n27942;
  assign n27944 = ~n27917 & ~n27943;
  assign n27945 = pi787 & ~n27944;
  assign n27946 = ~pi626 & ~n27910;
  assign n27947 = pi626 & ~n27882;
  assign n27948 = n17668 & ~n27947;
  assign n27949 = ~n27946 & n27948;
  assign n27950 = pi626 & ~n27910;
  assign n27951 = ~pi626 & ~n27882;
  assign n27952 = n17667 & ~n27951;
  assign n27953 = ~n27950 & n27952;
  assign n27954 = n17792 & n27931;
  assign n27955 = ~n27949 & ~n27954;
  assign n27956 = ~n27953 & n27955;
  assign n27957 = pi788 & ~n27956;
  assign n27958 = ~n16842 & ~n27919;
  assign n27959 = pi625 & n27958;
  assign n27960 = n27884 & ~n27958;
  assign n27961 = ~n27959 & ~n27960;
  assign n27962 = n27924 & ~n27961;
  assign n27963 = ~pi608 & ~n27923;
  assign n27964 = ~n27962 & n27963;
  assign n27965 = pi1153 & n27884;
  assign n27966 = ~n27959 & n27965;
  assign n27967 = pi608 & ~n27925;
  assign n27968 = ~n27966 & n27967;
  assign n27969 = ~n27964 & ~n27968;
  assign n27970 = pi778 & ~n27969;
  assign n27971 = ~pi778 & ~n27960;
  assign n27972 = ~n27970 & ~n27971;
  assign n27973 = ~pi609 & ~n27972;
  assign n27974 = pi609 & ~n27928;
  assign n27975 = ~pi1155 & ~n27974;
  assign n27976 = ~n27973 & n27975;
  assign n27977 = ~pi660 & ~n27889;
  assign n27978 = ~n27976 & n27977;
  assign n27979 = pi609 & ~n27972;
  assign n27980 = ~pi609 & ~n27928;
  assign n27981 = pi1155 & ~n27980;
  assign n27982 = ~n27979 & n27981;
  assign n27983 = pi660 & ~n27891;
  assign n27984 = ~n27982 & n27983;
  assign n27985 = ~n27978 & ~n27984;
  assign n27986 = pi785 & ~n27985;
  assign n27987 = ~pi785 & ~n27972;
  assign n27988 = ~n27986 & ~n27987;
  assign n27989 = ~pi618 & ~n27988;
  assign n27990 = pi618 & n27929;
  assign n27991 = ~pi1154 & ~n27990;
  assign n27992 = ~n27989 & n27991;
  assign n27993 = ~pi627 & ~n27897;
  assign n27994 = ~n27992 & n27993;
  assign n27995 = pi618 & ~n27988;
  assign n27996 = ~pi618 & n27929;
  assign n27997 = pi1154 & ~n27996;
  assign n27998 = ~n27995 & n27997;
  assign n27999 = pi627 & ~n27899;
  assign n28000 = ~n27998 & n27999;
  assign n28001 = ~n27994 & ~n28000;
  assign n28002 = pi781 & ~n28001;
  assign n28003 = ~pi781 & ~n27988;
  assign n28004 = ~n28002 & ~n28003;
  assign n28005 = ~pi619 & ~n28004;
  assign n28006 = pi619 & n27930;
  assign n28007 = ~pi1159 & ~n28006;
  assign n28008 = ~n28005 & n28007;
  assign n28009 = ~pi648 & ~n27905;
  assign n28010 = ~n28008 & n28009;
  assign n28011 = pi619 & ~n28004;
  assign n28012 = ~pi619 & n27930;
  assign n28013 = pi1159 & ~n28012;
  assign n28014 = ~n28011 & n28013;
  assign n28015 = pi648 & ~n27907;
  assign n28016 = ~n28014 & n28015;
  assign n28017 = pi789 & ~n28010;
  assign n28018 = ~n28016 & n28017;
  assign n28019 = ~pi789 & n28004;
  assign n28020 = n17905 & ~n28019;
  assign n28021 = ~n28018 & n28020;
  assign n28022 = ~n27957 & ~n28021;
  assign n28023 = ~n20298 & ~n28022;
  assign n28024 = n17944 & ~n27913;
  assign n28025 = n20786 & n27932;
  assign n28026 = ~n28024 & ~n28025;
  assign n28027 = ~pi629 & ~n28026;
  assign n28028 = n20790 & n27932;
  assign n28029 = n17943 & ~n27913;
  assign n28030 = ~n28028 & ~n28029;
  assign n28031 = pi629 & ~n28030;
  assign n28032 = ~n28027 & ~n28031;
  assign n28033 = pi792 & ~n28032;
  assign n28034 = n20300 & ~n28033;
  assign n28035 = ~n28023 & n28034;
  assign n28036 = ~n27945 & ~n28035;
  assign n28037 = pi644 & n28036;
  assign n28038 = ~pi787 & ~n27933;
  assign n28039 = pi787 & ~n27942;
  assign n28040 = ~n28038 & ~n28039;
  assign n28041 = ~pi644 & n28040;
  assign n28042 = pi715 & ~n28041;
  assign n28043 = ~n28037 & n28042;
  assign n28044 = ~n17740 & ~n27916;
  assign n28045 = n17740 & n27882;
  assign n28046 = ~n28044 & ~n28045;
  assign n28047 = pi644 & ~n28046;
  assign n28048 = ~pi644 & n27882;
  assign n28049 = ~pi715 & ~n28048;
  assign n28050 = ~n28047 & n28049;
  assign n28051 = pi1160 & ~n28050;
  assign n28052 = ~n28043 & n28051;
  assign n28053 = ~pi644 & n28036;
  assign n28054 = pi644 & n28040;
  assign n28055 = ~pi715 & ~n28054;
  assign n28056 = ~n28053 & n28055;
  assign n28057 = ~pi644 & ~n28046;
  assign n28058 = pi644 & n27882;
  assign n28059 = pi715 & ~n28058;
  assign n28060 = ~n28057 & n28059;
  assign n28061 = ~pi1160 & ~n28060;
  assign n28062 = ~n28056 & n28061;
  assign n28063 = ~n28052 & ~n28062;
  assign n28064 = pi790 & ~n28063;
  assign n28065 = ~pi790 & n28036;
  assign n28066 = pi832 & ~n28065;
  assign n28067 = ~n28064 & n28066;
  assign n28068 = ~pi184 & ~n17494;
  assign n28069 = n17627 & ~n28068;
  assign n28070 = ~pi737 & n3268;
  assign n28071 = n28068 & ~n28070;
  assign n28072 = pi184 & ~n18064;
  assign n28073 = ~pi38 & ~n28072;
  assign n28074 = n3268 & ~n28073;
  assign n28075 = ~pi184 & n18060;
  assign n28076 = ~n28074 & ~n28075;
  assign n28077 = ~pi184 & ~n16968;
  assign n28078 = n17480 & ~n28077;
  assign n28079 = ~pi737 & ~n28078;
  assign n28080 = ~n28076 & n28079;
  assign n28081 = ~n28071 & ~n28080;
  assign n28082 = ~pi778 & n28081;
  assign n28083 = pi625 & ~n28081;
  assign n28084 = ~pi625 & n28068;
  assign n28085 = pi1153 & ~n28084;
  assign n28086 = ~n28083 & n28085;
  assign n28087 = ~pi625 & ~n28081;
  assign n28088 = pi625 & n28068;
  assign n28089 = ~pi1153 & ~n28088;
  assign n28090 = ~n28087 & n28089;
  assign n28091 = ~n28086 & ~n28090;
  assign n28092 = pi778 & ~n28091;
  assign n28093 = ~n28082 & ~n28092;
  assign n28094 = ~n17554 & ~n28093;
  assign n28095 = n17554 & ~n28068;
  assign n28096 = ~n28094 & ~n28095;
  assign n28097 = ~n17591 & n28096;
  assign n28098 = n17591 & n28068;
  assign n28099 = ~n28097 & ~n28098;
  assign n28100 = ~n17627 & n28099;
  assign n28101 = ~n28069 & ~n28100;
  assign n28102 = ~n17670 & n28101;
  assign n28103 = n17670 & n28068;
  assign n28104 = ~n28102 & ~n28103;
  assign n28105 = ~pi792 & n28104;
  assign n28106 = pi628 & ~n28104;
  assign n28107 = ~pi628 & n28068;
  assign n28108 = pi1156 & ~n28107;
  assign n28109 = ~n28106 & n28108;
  assign n28110 = ~pi628 & ~n28104;
  assign n28111 = pi628 & n28068;
  assign n28112 = ~pi1156 & ~n28111;
  assign n28113 = ~n28110 & n28112;
  assign n28114 = ~n28109 & ~n28113;
  assign n28115 = pi792 & ~n28114;
  assign n28116 = ~n28105 & ~n28115;
  assign n28117 = ~pi647 & ~n28116;
  assign n28118 = pi647 & ~n28068;
  assign n28119 = ~n28117 & ~n28118;
  assign n28120 = ~pi1157 & n28119;
  assign n28121 = pi647 & ~n28116;
  assign n28122 = ~pi647 & ~n28068;
  assign n28123 = ~n28121 & ~n28122;
  assign n28124 = pi1157 & n28123;
  assign n28125 = ~n28120 & ~n28124;
  assign n28126 = pi787 & ~n28125;
  assign n28127 = ~pi787 & n28116;
  assign n28128 = ~n28126 & ~n28127;
  assign n28129 = ~pi644 & ~n28128;
  assign n28130 = pi715 & ~n28129;
  assign n28131 = pi184 & ~n3268;
  assign n28132 = ~pi777 & n16970;
  assign n28133 = ~n28077 & ~n28132;
  assign n28134 = pi38 & ~n28133;
  assign n28135 = ~pi184 & n16907;
  assign n28136 = pi184 & ~n16963;
  assign n28137 = ~pi777 & ~n28136;
  assign n28138 = ~n28135 & n28137;
  assign n28139 = ~pi184 & pi777;
  assign n28140 = ~n16816 & n28139;
  assign n28141 = ~n28138 & ~n28140;
  assign n28142 = ~pi38 & ~n28141;
  assign n28143 = ~n28134 & ~n28142;
  assign n28144 = n3268 & n28143;
  assign n28145 = ~n28131 & ~n28144;
  assign n28146 = ~n17526 & ~n28145;
  assign n28147 = n17526 & ~n28068;
  assign n28148 = ~n28146 & ~n28147;
  assign n28149 = ~pi785 & ~n28148;
  assign n28150 = ~n17527 & ~n28068;
  assign n28151 = pi609 & n28146;
  assign n28152 = ~n28150 & ~n28151;
  assign n28153 = pi1155 & ~n28152;
  assign n28154 = ~n17539 & ~n28068;
  assign n28155 = ~pi609 & n28146;
  assign n28156 = ~n28154 & ~n28155;
  assign n28157 = ~pi1155 & ~n28156;
  assign n28158 = ~n28153 & ~n28157;
  assign n28159 = pi785 & ~n28158;
  assign n28160 = ~n28149 & ~n28159;
  assign n28161 = ~pi781 & ~n28160;
  assign n28162 = pi618 & n28160;
  assign n28163 = ~pi618 & n28068;
  assign n28164 = pi1154 & ~n28163;
  assign n28165 = ~n28162 & n28164;
  assign n28166 = ~pi618 & n28160;
  assign n28167 = pi618 & n28068;
  assign n28168 = ~pi1154 & ~n28167;
  assign n28169 = ~n28166 & n28168;
  assign n28170 = ~n28165 & ~n28169;
  assign n28171 = pi781 & ~n28170;
  assign n28172 = ~n28161 & ~n28171;
  assign n28173 = ~pi789 & ~n28172;
  assign n28174 = pi619 & n28172;
  assign n28175 = ~pi619 & n28068;
  assign n28176 = pi1159 & ~n28175;
  assign n28177 = ~n28174 & n28176;
  assign n28178 = ~pi619 & n28172;
  assign n28179 = pi619 & n28068;
  assign n28180 = ~pi1159 & ~n28179;
  assign n28181 = ~n28178 & n28180;
  assign n28182 = ~n28177 & ~n28181;
  assign n28183 = pi789 & ~n28182;
  assign n28184 = ~n28173 & ~n28183;
  assign n28185 = ~n17904 & n28184;
  assign n28186 = n17904 & n28068;
  assign n28187 = ~n28185 & ~n28186;
  assign n28188 = ~n17698 & ~n28187;
  assign n28189 = n17698 & n28068;
  assign n28190 = ~n28188 & ~n28189;
  assign n28191 = ~n17740 & ~n28190;
  assign n28192 = n17740 & n28068;
  assign n28193 = ~n28191 & ~n28192;
  assign n28194 = pi644 & ~n28193;
  assign n28195 = ~pi644 & n28068;
  assign n28196 = ~pi715 & ~n28195;
  assign n28197 = ~n28194 & n28196;
  assign n28198 = pi1160 & ~n28197;
  assign n28199 = ~n28130 & n28198;
  assign n28200 = pi644 & ~n28128;
  assign n28201 = ~pi715 & ~n28200;
  assign n28202 = ~pi644 & ~n28193;
  assign n28203 = pi644 & n28068;
  assign n28204 = pi715 & ~n28203;
  assign n28205 = ~n28202 & n28204;
  assign n28206 = ~pi1160 & ~n28205;
  assign n28207 = ~n28201 & n28206;
  assign n28208 = ~n28199 & ~n28207;
  assign n28209 = pi790 & ~n28208;
  assign n28210 = ~pi644 & n28206;
  assign n28211 = pi644 & n28198;
  assign n28212 = pi790 & ~n28210;
  assign n28213 = ~n28211 & n28212;
  assign n28214 = ~n20502 & n28187;
  assign n28215 = ~pi629 & n28109;
  assign n28216 = pi629 & n28113;
  assign n28217 = ~n28215 & ~n28216;
  assign n28218 = ~n28214 & n28217;
  assign n28219 = pi792 & ~n28218;
  assign n28220 = pi737 & ~n28143;
  assign n28221 = ~pi184 & n17074;
  assign n28222 = pi184 & n17166;
  assign n28223 = pi777 & ~n28222;
  assign n28224 = ~n28221 & n28223;
  assign n28225 = pi184 & n17233;
  assign n28226 = ~pi184 & ~n17295;
  assign n28227 = ~pi777 & ~n28226;
  assign n28228 = ~n28225 & n28227;
  assign n28229 = pi39 & ~n28228;
  assign n28230 = ~n28224 & n28229;
  assign n28231 = pi184 & ~n17340;
  assign n28232 = ~pi184 & ~n17317;
  assign n28233 = pi777 & ~n28231;
  assign n28234 = ~n28232 & n28233;
  assign n28235 = ~pi184 & n17344;
  assign n28236 = pi184 & n17351;
  assign n28237 = ~pi777 & ~n28236;
  assign n28238 = ~n28235 & n28237;
  assign n28239 = ~n28234 & ~n28238;
  assign n28240 = ~pi39 & ~n28239;
  assign n28241 = ~pi38 & ~n28240;
  assign n28242 = ~n28230 & n28241;
  assign n28243 = ~pi777 & ~n17259;
  assign n28244 = n19303 & ~n28243;
  assign n28245 = ~pi184 & ~n28244;
  assign n28246 = ~n17154 & ~n27883;
  assign n28247 = pi184 & ~n28246;
  assign n28248 = n6250 & n28247;
  assign n28249 = pi38 & ~n28248;
  assign n28250 = ~n28245 & n28249;
  assign n28251 = ~pi737 & ~n28250;
  assign n28252 = ~n28242 & n28251;
  assign n28253 = n3268 & ~n28252;
  assign n28254 = ~n28220 & n28253;
  assign n28255 = ~n28131 & ~n28254;
  assign n28256 = ~pi625 & n28255;
  assign n28257 = pi625 & n28145;
  assign n28258 = ~pi1153 & ~n28257;
  assign n28259 = ~n28256 & n28258;
  assign n28260 = ~pi608 & ~n28086;
  assign n28261 = ~n28259 & n28260;
  assign n28262 = pi625 & n28255;
  assign n28263 = ~pi625 & n28145;
  assign n28264 = pi1153 & ~n28263;
  assign n28265 = ~n28262 & n28264;
  assign n28266 = pi608 & ~n28090;
  assign n28267 = ~n28265 & n28266;
  assign n28268 = ~n28261 & ~n28267;
  assign n28269 = pi778 & ~n28268;
  assign n28270 = ~pi778 & n28255;
  assign n28271 = ~n28269 & ~n28270;
  assign n28272 = ~pi609 & ~n28271;
  assign n28273 = pi609 & n28093;
  assign n28274 = ~pi1155 & ~n28273;
  assign n28275 = ~n28272 & n28274;
  assign n28276 = ~pi660 & ~n28153;
  assign n28277 = ~n28275 & n28276;
  assign n28278 = pi609 & ~n28271;
  assign n28279 = ~pi609 & n28093;
  assign n28280 = pi1155 & ~n28279;
  assign n28281 = ~n28278 & n28280;
  assign n28282 = pi660 & ~n28157;
  assign n28283 = ~n28281 & n28282;
  assign n28284 = ~n28277 & ~n28283;
  assign n28285 = pi785 & ~n28284;
  assign n28286 = ~pi785 & ~n28271;
  assign n28287 = ~n28285 & ~n28286;
  assign n28288 = ~pi618 & ~n28287;
  assign n28289 = pi618 & n28096;
  assign n28290 = ~pi1154 & ~n28289;
  assign n28291 = ~n28288 & n28290;
  assign n28292 = ~pi627 & ~n28165;
  assign n28293 = ~n28291 & n28292;
  assign n28294 = pi618 & ~n28287;
  assign n28295 = ~pi618 & n28096;
  assign n28296 = pi1154 & ~n28295;
  assign n28297 = ~n28294 & n28296;
  assign n28298 = pi627 & ~n28169;
  assign n28299 = ~n28297 & n28298;
  assign n28300 = ~n28293 & ~n28299;
  assign n28301 = pi781 & ~n28300;
  assign n28302 = ~pi781 & ~n28287;
  assign n28303 = ~n28301 & ~n28302;
  assign n28304 = ~pi619 & ~n28303;
  assign n28305 = pi619 & ~n28099;
  assign n28306 = ~pi1159 & ~n28305;
  assign n28307 = ~n28304 & n28306;
  assign n28308 = ~pi648 & ~n28177;
  assign n28309 = ~n28307 & n28308;
  assign n28310 = pi619 & ~n28303;
  assign n28311 = ~pi619 & ~n28099;
  assign n28312 = pi1159 & ~n28311;
  assign n28313 = ~n28310 & n28312;
  assign n28314 = pi648 & ~n28181;
  assign n28315 = ~n28313 & n28314;
  assign n28316 = pi789 & ~n28309;
  assign n28317 = ~n28315 & n28316;
  assign n28318 = ~pi789 & n28303;
  assign n28319 = n17905 & ~n28318;
  assign n28320 = ~n28317 & n28319;
  assign n28321 = ~pi626 & ~n28184;
  assign n28322 = pi626 & ~n28068;
  assign n28323 = n17668 & ~n28322;
  assign n28324 = ~n28321 & n28323;
  assign n28325 = pi626 & ~n28184;
  assign n28326 = ~pi626 & ~n28068;
  assign n28327 = n17667 & ~n28326;
  assign n28328 = ~n28325 & n28327;
  assign n28329 = n17792 & n28101;
  assign n28330 = ~n28324 & ~n28329;
  assign n28331 = ~n28328 & n28330;
  assign n28332 = pi788 & ~n28331;
  assign n28333 = ~n20298 & ~n28332;
  assign n28334 = ~n28320 & n28333;
  assign n28335 = ~n28219 & ~n28334;
  assign n28336 = n20300 & ~n28335;
  assign n28337 = ~n20491 & n28190;
  assign n28338 = n17738 & ~n28119;
  assign n28339 = n17737 & ~n28123;
  assign n28340 = ~n28338 & ~n28339;
  assign n28341 = ~n28337 & n28340;
  assign n28342 = pi787 & ~n28341;
  assign n28343 = ~n28336 & ~n28342;
  assign n28344 = ~n28213 & n28343;
  assign n28345 = ~n28209 & ~n28344;
  assign n28346 = ~po1038 & ~n28345;
  assign n28347 = ~pi184 & po1038;
  assign n28348 = ~pi832 & ~n28347;
  assign n28349 = ~n28346 & n28348;
  assign po341 = ~n28067 & ~n28349;
  assign n28351 = ~pi185 & ~n2755;
  assign n28352 = ~pi751 & n16933;
  assign n28353 = ~n28351 & ~n28352;
  assign n28354 = ~n17794 & ~n28353;
  assign n28355 = ~pi785 & ~n28354;
  assign n28356 = n17539 & n28352;
  assign n28357 = n28354 & ~n28356;
  assign n28358 = pi1155 & ~n28357;
  assign n28359 = ~pi1155 & ~n28351;
  assign n28360 = ~n28356 & n28359;
  assign n28361 = ~n28358 & ~n28360;
  assign n28362 = pi785 & ~n28361;
  assign n28363 = ~n28355 & ~n28362;
  assign n28364 = ~pi781 & ~n28363;
  assign n28365 = ~n17809 & n28363;
  assign n28366 = pi1154 & ~n28365;
  assign n28367 = ~n17812 & n28363;
  assign n28368 = ~pi1154 & ~n28367;
  assign n28369 = ~n28366 & ~n28368;
  assign n28370 = pi781 & ~n28369;
  assign n28371 = ~n28364 & ~n28370;
  assign n28372 = ~pi789 & ~n28371;
  assign n28373 = ~n22988 & n28371;
  assign n28374 = pi1159 & ~n28373;
  assign n28375 = ~n22991 & n28371;
  assign n28376 = ~pi1159 & ~n28375;
  assign n28377 = ~n28374 & ~n28376;
  assign n28378 = pi789 & ~n28377;
  assign n28379 = ~n28372 & ~n28378;
  assign n28380 = ~n17904 & n28379;
  assign n28381 = n17904 & n28351;
  assign n28382 = ~n28380 & ~n28381;
  assign n28383 = ~n17698 & ~n28382;
  assign n28384 = n17698 & n28351;
  assign n28385 = ~n28383 & ~n28384;
  assign n28386 = ~n20491 & n28385;
  assign n28387 = ~pi701 & n17153;
  assign n28388 = ~n28351 & ~n28387;
  assign n28389 = ~pi778 & ~n28388;
  assign n28390 = ~pi625 & n28387;
  assign n28391 = ~n28388 & ~n28390;
  assign n28392 = pi1153 & ~n28391;
  assign n28393 = ~pi1153 & ~n28351;
  assign n28394 = ~n28390 & n28393;
  assign n28395 = pi778 & ~n28394;
  assign n28396 = ~n28392 & n28395;
  assign n28397 = ~n28389 & ~n28396;
  assign n28398 = ~n17780 & ~n28397;
  assign n28399 = ~n17782 & n28398;
  assign n28400 = ~n17784 & n28399;
  assign n28401 = ~n17916 & n28400;
  assign n28402 = ~n17947 & n28401;
  assign n28403 = ~pi647 & n28402;
  assign n28404 = pi647 & n28351;
  assign n28405 = ~pi1157 & ~n28404;
  assign n28406 = ~n28403 & n28405;
  assign n28407 = pi647 & ~n28402;
  assign n28408 = ~pi647 & ~n28351;
  assign n28409 = ~n28407 & ~n28408;
  assign n28410 = pi1157 & ~n28409;
  assign n28411 = ~n28406 & ~n28410;
  assign n28412 = ~n17739 & ~n28411;
  assign n28413 = ~n28386 & ~n28412;
  assign n28414 = pi787 & ~n28413;
  assign n28415 = ~pi626 & ~n28379;
  assign n28416 = pi626 & ~n28351;
  assign n28417 = n17668 & ~n28416;
  assign n28418 = ~n28415 & n28417;
  assign n28419 = pi626 & ~n28379;
  assign n28420 = ~pi626 & ~n28351;
  assign n28421 = n17667 & ~n28420;
  assign n28422 = ~n28419 & n28421;
  assign n28423 = n17792 & n28400;
  assign n28424 = ~n28418 & ~n28423;
  assign n28425 = ~n28422 & n28424;
  assign n28426 = pi788 & ~n28425;
  assign n28427 = ~n16842 & ~n28388;
  assign n28428 = pi625 & n28427;
  assign n28429 = n28353 & ~n28427;
  assign n28430 = ~n28428 & ~n28429;
  assign n28431 = n28393 & ~n28430;
  assign n28432 = ~pi608 & ~n28392;
  assign n28433 = ~n28431 & n28432;
  assign n28434 = pi1153 & n28353;
  assign n28435 = ~n28428 & n28434;
  assign n28436 = pi608 & ~n28394;
  assign n28437 = ~n28435 & n28436;
  assign n28438 = ~n28433 & ~n28437;
  assign n28439 = pi778 & ~n28438;
  assign n28440 = ~pi778 & ~n28429;
  assign n28441 = ~n28439 & ~n28440;
  assign n28442 = ~pi609 & ~n28441;
  assign n28443 = pi609 & ~n28397;
  assign n28444 = ~pi1155 & ~n28443;
  assign n28445 = ~n28442 & n28444;
  assign n28446 = ~pi660 & ~n28358;
  assign n28447 = ~n28445 & n28446;
  assign n28448 = pi609 & ~n28441;
  assign n28449 = ~pi609 & ~n28397;
  assign n28450 = pi1155 & ~n28449;
  assign n28451 = ~n28448 & n28450;
  assign n28452 = pi660 & ~n28360;
  assign n28453 = ~n28451 & n28452;
  assign n28454 = ~n28447 & ~n28453;
  assign n28455 = pi785 & ~n28454;
  assign n28456 = ~pi785 & ~n28441;
  assign n28457 = ~n28455 & ~n28456;
  assign n28458 = ~pi618 & ~n28457;
  assign n28459 = pi618 & n28398;
  assign n28460 = ~pi1154 & ~n28459;
  assign n28461 = ~n28458 & n28460;
  assign n28462 = ~pi627 & ~n28366;
  assign n28463 = ~n28461 & n28462;
  assign n28464 = pi618 & ~n28457;
  assign n28465 = ~pi618 & n28398;
  assign n28466 = pi1154 & ~n28465;
  assign n28467 = ~n28464 & n28466;
  assign n28468 = pi627 & ~n28368;
  assign n28469 = ~n28467 & n28468;
  assign n28470 = ~n28463 & ~n28469;
  assign n28471 = pi781 & ~n28470;
  assign n28472 = ~pi781 & ~n28457;
  assign n28473 = ~n28471 & ~n28472;
  assign n28474 = ~pi619 & ~n28473;
  assign n28475 = pi619 & n28399;
  assign n28476 = ~pi1159 & ~n28475;
  assign n28477 = ~n28474 & n28476;
  assign n28478 = ~pi648 & ~n28374;
  assign n28479 = ~n28477 & n28478;
  assign n28480 = pi619 & ~n28473;
  assign n28481 = ~pi619 & n28399;
  assign n28482 = pi1159 & ~n28481;
  assign n28483 = ~n28480 & n28482;
  assign n28484 = pi648 & ~n28376;
  assign n28485 = ~n28483 & n28484;
  assign n28486 = pi789 & ~n28479;
  assign n28487 = ~n28485 & n28486;
  assign n28488 = ~pi789 & n28473;
  assign n28489 = n17905 & ~n28488;
  assign n28490 = ~n28487 & n28489;
  assign n28491 = ~n28426 & ~n28490;
  assign n28492 = ~n20298 & ~n28491;
  assign n28493 = n17944 & ~n28382;
  assign n28494 = n20786 & n28401;
  assign n28495 = ~n28493 & ~n28494;
  assign n28496 = ~pi629 & ~n28495;
  assign n28497 = n20790 & n28401;
  assign n28498 = n17943 & ~n28382;
  assign n28499 = ~n28497 & ~n28498;
  assign n28500 = pi629 & ~n28499;
  assign n28501 = ~n28496 & ~n28500;
  assign n28502 = pi792 & ~n28501;
  assign n28503 = n20300 & ~n28502;
  assign n28504 = ~n28492 & n28503;
  assign n28505 = ~n28414 & ~n28504;
  assign n28506 = pi644 & n28505;
  assign n28507 = ~pi787 & ~n28402;
  assign n28508 = pi787 & ~n28411;
  assign n28509 = ~n28507 & ~n28508;
  assign n28510 = ~pi644 & n28509;
  assign n28511 = pi715 & ~n28510;
  assign n28512 = ~n28506 & n28511;
  assign n28513 = ~n17740 & ~n28385;
  assign n28514 = n17740 & n28351;
  assign n28515 = ~n28513 & ~n28514;
  assign n28516 = pi644 & ~n28515;
  assign n28517 = ~pi644 & n28351;
  assign n28518 = ~pi715 & ~n28517;
  assign n28519 = ~n28516 & n28518;
  assign n28520 = pi1160 & ~n28519;
  assign n28521 = ~n28512 & n28520;
  assign n28522 = ~pi644 & n28505;
  assign n28523 = pi644 & n28509;
  assign n28524 = ~pi715 & ~n28523;
  assign n28525 = ~n28522 & n28524;
  assign n28526 = ~pi644 & ~n28515;
  assign n28527 = pi644 & n28351;
  assign n28528 = pi715 & ~n28527;
  assign n28529 = ~n28526 & n28528;
  assign n28530 = ~pi1160 & ~n28529;
  assign n28531 = ~n28525 & n28530;
  assign n28532 = ~n28521 & ~n28531;
  assign n28533 = pi790 & ~n28532;
  assign n28534 = ~pi790 & n28505;
  assign n28535 = pi832 & ~n28534;
  assign n28536 = ~n28533 & n28535;
  assign n28537 = ~pi185 & ~n17494;
  assign n28538 = n17627 & ~n28537;
  assign n28539 = ~pi701 & n3268;
  assign n28540 = n28537 & ~n28539;
  assign n28541 = pi185 & ~n18064;
  assign n28542 = ~pi38 & ~n28541;
  assign n28543 = n3268 & ~n28542;
  assign n28544 = ~pi185 & n18060;
  assign n28545 = ~n28543 & ~n28544;
  assign n28546 = ~pi185 & ~n16968;
  assign n28547 = n17480 & ~n28546;
  assign n28548 = ~pi701 & ~n28547;
  assign n28549 = ~n28545 & n28548;
  assign n28550 = ~n28540 & ~n28549;
  assign n28551 = ~pi778 & n28550;
  assign n28552 = pi625 & ~n28550;
  assign n28553 = ~pi625 & n28537;
  assign n28554 = pi1153 & ~n28553;
  assign n28555 = ~n28552 & n28554;
  assign n28556 = ~pi625 & ~n28550;
  assign n28557 = pi625 & n28537;
  assign n28558 = ~pi1153 & ~n28557;
  assign n28559 = ~n28556 & n28558;
  assign n28560 = ~n28555 & ~n28559;
  assign n28561 = pi778 & ~n28560;
  assign n28562 = ~n28551 & ~n28561;
  assign n28563 = ~n17554 & ~n28562;
  assign n28564 = n17554 & ~n28537;
  assign n28565 = ~n28563 & ~n28564;
  assign n28566 = ~n17591 & n28565;
  assign n28567 = n17591 & n28537;
  assign n28568 = ~n28566 & ~n28567;
  assign n28569 = ~n17627 & n28568;
  assign n28570 = ~n28538 & ~n28569;
  assign n28571 = ~n17670 & n28570;
  assign n28572 = n17670 & n28537;
  assign n28573 = ~n28571 & ~n28572;
  assign n28574 = ~pi792 & n28573;
  assign n28575 = pi628 & ~n28573;
  assign n28576 = ~pi628 & n28537;
  assign n28577 = pi1156 & ~n28576;
  assign n28578 = ~n28575 & n28577;
  assign n28579 = ~pi628 & ~n28573;
  assign n28580 = pi628 & n28537;
  assign n28581 = ~pi1156 & ~n28580;
  assign n28582 = ~n28579 & n28581;
  assign n28583 = ~n28578 & ~n28582;
  assign n28584 = pi792 & ~n28583;
  assign n28585 = ~n28574 & ~n28584;
  assign n28586 = ~pi647 & ~n28585;
  assign n28587 = pi647 & ~n28537;
  assign n28588 = ~n28586 & ~n28587;
  assign n28589 = ~pi1157 & n28588;
  assign n28590 = pi647 & ~n28585;
  assign n28591 = ~pi647 & ~n28537;
  assign n28592 = ~n28590 & ~n28591;
  assign n28593 = pi1157 & n28592;
  assign n28594 = ~n28589 & ~n28593;
  assign n28595 = pi787 & ~n28594;
  assign n28596 = ~pi787 & n28585;
  assign n28597 = ~n28595 & ~n28596;
  assign n28598 = ~pi644 & ~n28597;
  assign n28599 = pi715 & ~n28598;
  assign n28600 = pi185 & ~n3268;
  assign n28601 = pi751 & n16814;
  assign n28602 = pi185 & n16961;
  assign n28603 = ~n28601 & ~n28602;
  assign n28604 = pi39 & ~n28603;
  assign n28605 = ~pi185 & ~pi751;
  assign n28606 = n16907 & n28605;
  assign n28607 = pi185 & pi751;
  assign n28608 = pi185 & ~n16918;
  assign n28609 = ~n21193 & ~n28608;
  assign n28610 = ~pi39 & ~n28609;
  assign n28611 = ~n28607 & ~n28610;
  assign n28612 = ~n28606 & n28611;
  assign n28613 = ~n28604 & n28612;
  assign n28614 = ~pi38 & ~n28613;
  assign n28615 = ~pi751 & n16970;
  assign n28616 = pi38 & ~n28546;
  assign n28617 = ~n28615 & n28616;
  assign n28618 = ~n28614 & ~n28617;
  assign n28619 = n3268 & ~n28618;
  assign n28620 = ~n28600 & ~n28619;
  assign n28621 = ~n17526 & ~n28620;
  assign n28622 = n17526 & ~n28537;
  assign n28623 = ~n28621 & ~n28622;
  assign n28624 = ~pi785 & ~n28623;
  assign n28625 = ~n17527 & ~n28537;
  assign n28626 = pi609 & n28621;
  assign n28627 = ~n28625 & ~n28626;
  assign n28628 = pi1155 & ~n28627;
  assign n28629 = ~n17539 & ~n28537;
  assign n28630 = ~pi609 & n28621;
  assign n28631 = ~n28629 & ~n28630;
  assign n28632 = ~pi1155 & ~n28631;
  assign n28633 = ~n28628 & ~n28632;
  assign n28634 = pi785 & ~n28633;
  assign n28635 = ~n28624 & ~n28634;
  assign n28636 = ~pi781 & ~n28635;
  assign n28637 = pi618 & n28635;
  assign n28638 = ~pi618 & n28537;
  assign n28639 = pi1154 & ~n28638;
  assign n28640 = ~n28637 & n28639;
  assign n28641 = ~pi618 & n28635;
  assign n28642 = pi618 & n28537;
  assign n28643 = ~pi1154 & ~n28642;
  assign n28644 = ~n28641 & n28643;
  assign n28645 = ~n28640 & ~n28644;
  assign n28646 = pi781 & ~n28645;
  assign n28647 = ~n28636 & ~n28646;
  assign n28648 = ~pi789 & ~n28647;
  assign n28649 = pi619 & n28647;
  assign n28650 = ~pi619 & n28537;
  assign n28651 = pi1159 & ~n28650;
  assign n28652 = ~n28649 & n28651;
  assign n28653 = ~pi619 & n28647;
  assign n28654 = pi619 & n28537;
  assign n28655 = ~pi1159 & ~n28654;
  assign n28656 = ~n28653 & n28655;
  assign n28657 = ~n28652 & ~n28656;
  assign n28658 = pi789 & ~n28657;
  assign n28659 = ~n28648 & ~n28658;
  assign n28660 = ~n17904 & n28659;
  assign n28661 = n17904 & n28537;
  assign n28662 = ~n28660 & ~n28661;
  assign n28663 = ~n17698 & ~n28662;
  assign n28664 = n17698 & n28537;
  assign n28665 = ~n28663 & ~n28664;
  assign n28666 = ~n17740 & ~n28665;
  assign n28667 = n17740 & n28537;
  assign n28668 = ~n28666 & ~n28667;
  assign n28669 = pi644 & ~n28668;
  assign n28670 = ~pi644 & n28537;
  assign n28671 = ~pi715 & ~n28670;
  assign n28672 = ~n28669 & n28671;
  assign n28673 = pi1160 & ~n28672;
  assign n28674 = ~n28599 & n28673;
  assign n28675 = pi644 & ~n28597;
  assign n28676 = ~pi715 & ~n28675;
  assign n28677 = ~pi644 & ~n28668;
  assign n28678 = pi644 & n28537;
  assign n28679 = pi715 & ~n28678;
  assign n28680 = ~n28677 & n28679;
  assign n28681 = ~pi1160 & ~n28680;
  assign n28682 = ~n28676 & n28681;
  assign n28683 = ~n28674 & ~n28682;
  assign n28684 = pi790 & ~n28683;
  assign n28685 = ~pi644 & n28681;
  assign n28686 = pi644 & n28673;
  assign n28687 = pi790 & ~n28685;
  assign n28688 = ~n28686 & n28687;
  assign n28689 = ~n20502 & n28662;
  assign n28690 = ~pi629 & n28578;
  assign n28691 = pi629 & n28582;
  assign n28692 = ~n28690 & ~n28691;
  assign n28693 = ~n28689 & n28692;
  assign n28694 = pi792 & ~n28693;
  assign n28695 = pi701 & n28618;
  assign n28696 = ~pi185 & n17074;
  assign n28697 = pi185 & n17166;
  assign n28698 = pi751 & ~n28697;
  assign n28699 = ~n28696 & n28698;
  assign n28700 = pi185 & n17233;
  assign n28701 = ~pi185 & ~n17295;
  assign n28702 = ~pi751 & ~n28701;
  assign n28703 = ~n28700 & n28702;
  assign n28704 = pi39 & ~n28703;
  assign n28705 = ~n28699 & n28704;
  assign n28706 = pi185 & ~n17340;
  assign n28707 = ~pi185 & ~n17317;
  assign n28708 = pi751 & ~n28706;
  assign n28709 = ~n28707 & n28708;
  assign n28710 = ~pi185 & n17344;
  assign n28711 = pi185 & n17351;
  assign n28712 = ~pi751 & ~n28711;
  assign n28713 = ~n28710 & n28712;
  assign n28714 = ~n28709 & ~n28713;
  assign n28715 = ~pi39 & ~n28714;
  assign n28716 = ~pi38 & ~n28715;
  assign n28717 = ~n28705 & n28716;
  assign n28718 = ~pi751 & ~n17259;
  assign n28719 = n19303 & ~n28718;
  assign n28720 = ~pi185 & ~n28719;
  assign n28721 = ~n17154 & ~n28352;
  assign n28722 = pi185 & ~n28721;
  assign n28723 = n6250 & n28722;
  assign n28724 = pi38 & ~n28723;
  assign n28725 = ~n28720 & n28724;
  assign n28726 = ~pi701 & ~n28725;
  assign n28727 = ~n28717 & n28726;
  assign n28728 = n3268 & ~n28727;
  assign n28729 = ~n28695 & n28728;
  assign n28730 = ~n28600 & ~n28729;
  assign n28731 = ~pi625 & n28730;
  assign n28732 = pi625 & n28620;
  assign n28733 = ~pi1153 & ~n28732;
  assign n28734 = ~n28731 & n28733;
  assign n28735 = ~pi608 & ~n28555;
  assign n28736 = ~n28734 & n28735;
  assign n28737 = pi625 & n28730;
  assign n28738 = ~pi625 & n28620;
  assign n28739 = pi1153 & ~n28738;
  assign n28740 = ~n28737 & n28739;
  assign n28741 = pi608 & ~n28559;
  assign n28742 = ~n28740 & n28741;
  assign n28743 = ~n28736 & ~n28742;
  assign n28744 = pi778 & ~n28743;
  assign n28745 = ~pi778 & n28730;
  assign n28746 = ~n28744 & ~n28745;
  assign n28747 = ~pi609 & ~n28746;
  assign n28748 = pi609 & n28562;
  assign n28749 = ~pi1155 & ~n28748;
  assign n28750 = ~n28747 & n28749;
  assign n28751 = ~pi660 & ~n28628;
  assign n28752 = ~n28750 & n28751;
  assign n28753 = pi609 & ~n28746;
  assign n28754 = ~pi609 & n28562;
  assign n28755 = pi1155 & ~n28754;
  assign n28756 = ~n28753 & n28755;
  assign n28757 = pi660 & ~n28632;
  assign n28758 = ~n28756 & n28757;
  assign n28759 = ~n28752 & ~n28758;
  assign n28760 = pi785 & ~n28759;
  assign n28761 = ~pi785 & ~n28746;
  assign n28762 = ~n28760 & ~n28761;
  assign n28763 = ~pi618 & ~n28762;
  assign n28764 = pi618 & n28565;
  assign n28765 = ~pi1154 & ~n28764;
  assign n28766 = ~n28763 & n28765;
  assign n28767 = ~pi627 & ~n28640;
  assign n28768 = ~n28766 & n28767;
  assign n28769 = pi618 & ~n28762;
  assign n28770 = ~pi618 & n28565;
  assign n28771 = pi1154 & ~n28770;
  assign n28772 = ~n28769 & n28771;
  assign n28773 = pi627 & ~n28644;
  assign n28774 = ~n28772 & n28773;
  assign n28775 = ~n28768 & ~n28774;
  assign n28776 = pi781 & ~n28775;
  assign n28777 = ~pi781 & ~n28762;
  assign n28778 = ~n28776 & ~n28777;
  assign n28779 = ~pi619 & ~n28778;
  assign n28780 = pi619 & ~n28568;
  assign n28781 = ~pi1159 & ~n28780;
  assign n28782 = ~n28779 & n28781;
  assign n28783 = ~pi648 & ~n28652;
  assign n28784 = ~n28782 & n28783;
  assign n28785 = pi619 & ~n28778;
  assign n28786 = ~pi619 & ~n28568;
  assign n28787 = pi1159 & ~n28786;
  assign n28788 = ~n28785 & n28787;
  assign n28789 = pi648 & ~n28656;
  assign n28790 = ~n28788 & n28789;
  assign n28791 = pi789 & ~n28784;
  assign n28792 = ~n28790 & n28791;
  assign n28793 = ~pi789 & n28778;
  assign n28794 = n17905 & ~n28793;
  assign n28795 = ~n28792 & n28794;
  assign n28796 = ~pi626 & ~n28659;
  assign n28797 = pi626 & ~n28537;
  assign n28798 = n17668 & ~n28797;
  assign n28799 = ~n28796 & n28798;
  assign n28800 = pi626 & ~n28659;
  assign n28801 = ~pi626 & ~n28537;
  assign n28802 = n17667 & ~n28801;
  assign n28803 = ~n28800 & n28802;
  assign n28804 = n17792 & n28570;
  assign n28805 = ~n28799 & ~n28804;
  assign n28806 = ~n28803 & n28805;
  assign n28807 = pi788 & ~n28806;
  assign n28808 = ~n20298 & ~n28807;
  assign n28809 = ~n28795 & n28808;
  assign n28810 = ~n28694 & ~n28809;
  assign n28811 = n20300 & ~n28810;
  assign n28812 = ~n20491 & n28665;
  assign n28813 = n17738 & ~n28588;
  assign n28814 = n17737 & ~n28592;
  assign n28815 = ~n28813 & ~n28814;
  assign n28816 = ~n28812 & n28815;
  assign n28817 = pi787 & ~n28816;
  assign n28818 = ~n28811 & ~n28817;
  assign n28819 = ~n28688 & n28818;
  assign n28820 = ~n28684 & ~n28819;
  assign n28821 = ~po1038 & ~n28820;
  assign n28822 = ~pi185 & po1038;
  assign n28823 = ~pi832 & ~n28822;
  assign n28824 = ~n28821 & n28823;
  assign po342 = ~n28536 & ~n28824;
  assign n28826 = pi186 & ~n3268;
  assign n28827 = ~pi186 & n19309;
  assign n28828 = pi186 & n19314;
  assign n28829 = pi752 & ~n19316;
  assign n28830 = ~n28828 & n28829;
  assign n28831 = ~n28827 & n28830;
  assign n28832 = pi186 & n19326;
  assign n28833 = ~pi186 & ~n19334;
  assign n28834 = ~pi752 & ~n28833;
  assign n28835 = ~n28832 & n28834;
  assign n28836 = pi703 & ~n28835;
  assign n28837 = ~n28831 & n28836;
  assign n28838 = ~pi186 & ~n17487;
  assign n28839 = pi752 & ~n28838;
  assign n28840 = pi186 & ~n19344;
  assign n28841 = ~pi186 & ~pi752;
  assign n28842 = n19349 & n28841;
  assign n28843 = ~n28840 & ~n28842;
  assign n28844 = ~n19343 & ~n28843;
  assign n28845 = ~n28839 & ~n28844;
  assign n28846 = ~pi703 & n28845;
  assign n28847 = n3268 & ~n28837;
  assign n28848 = ~n28846 & n28847;
  assign n28849 = ~n28826 & ~n28848;
  assign n28850 = ~pi625 & n28849;
  assign n28851 = n3268 & ~n28845;
  assign n28852 = ~n28826 & ~n28851;
  assign n28853 = pi625 & n28852;
  assign n28854 = ~pi1153 & ~n28853;
  assign n28855 = ~n28850 & n28854;
  assign n28856 = ~pi703 & n28838;
  assign n28857 = ~pi186 & n18060;
  assign n28858 = pi186 & ~n18064;
  assign n28859 = ~pi38 & ~n28858;
  assign n28860 = ~n28857 & n28859;
  assign n28861 = ~pi186 & ~n16968;
  assign n28862 = n17480 & ~n28861;
  assign n28863 = pi703 & ~n28862;
  assign n28864 = ~n28860 & n28863;
  assign n28865 = n3268 & ~n28856;
  assign n28866 = ~n28864 & n28865;
  assign n28867 = ~n28826 & ~n28866;
  assign n28868 = pi625 & n28867;
  assign n28869 = ~pi186 & ~n17494;
  assign n28870 = ~pi625 & n28869;
  assign n28871 = pi1153 & ~n28870;
  assign n28872 = ~n28868 & n28871;
  assign n28873 = ~pi608 & ~n28872;
  assign n28874 = ~n28855 & n28873;
  assign n28875 = pi625 & n28849;
  assign n28876 = ~pi625 & n28852;
  assign n28877 = pi1153 & ~n28876;
  assign n28878 = ~n28875 & n28877;
  assign n28879 = ~pi625 & n28867;
  assign n28880 = pi625 & n28869;
  assign n28881 = ~pi1153 & ~n28880;
  assign n28882 = ~n28879 & n28881;
  assign n28883 = pi608 & ~n28882;
  assign n28884 = ~n28878 & n28883;
  assign n28885 = ~n28874 & ~n28884;
  assign n28886 = pi778 & ~n28885;
  assign n28887 = ~pi778 & n28849;
  assign n28888 = ~n28886 & ~n28887;
  assign n28889 = ~pi609 & ~n28888;
  assign n28890 = ~pi778 & ~n28867;
  assign n28891 = ~n28872 & ~n28882;
  assign n28892 = pi778 & ~n28891;
  assign n28893 = ~n28890 & ~n28892;
  assign n28894 = pi609 & n28893;
  assign n28895 = ~pi1155 & ~n28894;
  assign n28896 = ~n28889 & n28895;
  assign n28897 = ~n17527 & ~n28869;
  assign n28898 = ~n17526 & ~n28852;
  assign n28899 = pi609 & n28898;
  assign n28900 = ~n28897 & ~n28899;
  assign n28901 = pi1155 & ~n28900;
  assign n28902 = ~pi660 & ~n28901;
  assign n28903 = ~n28896 & n28902;
  assign n28904 = pi609 & ~n28888;
  assign n28905 = ~pi609 & n28893;
  assign n28906 = pi1155 & ~n28905;
  assign n28907 = ~n28904 & n28906;
  assign n28908 = ~n17539 & ~n28869;
  assign n28909 = ~pi609 & n28898;
  assign n28910 = ~n28908 & ~n28909;
  assign n28911 = ~pi1155 & ~n28910;
  assign n28912 = pi660 & ~n28911;
  assign n28913 = ~n28907 & n28912;
  assign n28914 = ~n28903 & ~n28913;
  assign n28915 = pi785 & ~n28914;
  assign n28916 = ~pi785 & ~n28888;
  assign n28917 = ~n28915 & ~n28916;
  assign n28918 = ~pi618 & ~n28917;
  assign n28919 = ~n17554 & ~n28893;
  assign n28920 = n17554 & ~n28869;
  assign n28921 = ~n28919 & ~n28920;
  assign n28922 = pi618 & n28921;
  assign n28923 = ~pi1154 & ~n28922;
  assign n28924 = ~n28918 & n28923;
  assign n28925 = n17526 & ~n28869;
  assign n28926 = ~n28898 & ~n28925;
  assign n28927 = ~pi785 & ~n28926;
  assign n28928 = ~n28901 & ~n28911;
  assign n28929 = pi785 & ~n28928;
  assign n28930 = ~n28927 & ~n28929;
  assign n28931 = pi618 & n28930;
  assign n28932 = ~pi618 & n28869;
  assign n28933 = pi1154 & ~n28932;
  assign n28934 = ~n28931 & n28933;
  assign n28935 = ~pi627 & ~n28934;
  assign n28936 = ~n28924 & n28935;
  assign n28937 = pi618 & ~n28917;
  assign n28938 = ~pi618 & n28921;
  assign n28939 = pi1154 & ~n28938;
  assign n28940 = ~n28937 & n28939;
  assign n28941 = ~pi618 & n28930;
  assign n28942 = pi618 & n28869;
  assign n28943 = ~pi1154 & ~n28942;
  assign n28944 = ~n28941 & n28943;
  assign n28945 = pi627 & ~n28944;
  assign n28946 = ~n28940 & n28945;
  assign n28947 = ~n28936 & ~n28946;
  assign n28948 = pi781 & ~n28947;
  assign n28949 = ~pi781 & ~n28917;
  assign n28950 = ~n28948 & ~n28949;
  assign n28951 = ~pi619 & ~n28950;
  assign n28952 = ~n17591 & n28921;
  assign n28953 = n17591 & n28869;
  assign n28954 = ~n28952 & ~n28953;
  assign n28955 = pi619 & ~n28954;
  assign n28956 = ~pi1159 & ~n28955;
  assign n28957 = ~n28951 & n28956;
  assign n28958 = ~pi781 & ~n28930;
  assign n28959 = ~n28934 & ~n28944;
  assign n28960 = pi781 & ~n28959;
  assign n28961 = ~n28958 & ~n28960;
  assign n28962 = pi619 & n28961;
  assign n28963 = ~pi619 & n28869;
  assign n28964 = pi1159 & ~n28963;
  assign n28965 = ~n28962 & n28964;
  assign n28966 = ~pi648 & ~n28965;
  assign n28967 = ~n28957 & n28966;
  assign n28968 = pi619 & ~n28950;
  assign n28969 = ~pi619 & ~n28954;
  assign n28970 = pi1159 & ~n28969;
  assign n28971 = ~n28968 & n28970;
  assign n28972 = ~pi619 & n28961;
  assign n28973 = pi619 & n28869;
  assign n28974 = ~pi1159 & ~n28973;
  assign n28975 = ~n28972 & n28974;
  assign n28976 = pi648 & ~n28975;
  assign n28977 = ~n28971 & n28976;
  assign n28978 = ~n28967 & ~n28977;
  assign n28979 = pi789 & ~n28978;
  assign n28980 = ~pi789 & ~n28950;
  assign n28981 = ~n28979 & ~n28980;
  assign n28982 = ~pi788 & n28981;
  assign n28983 = ~pi626 & n28981;
  assign n28984 = n17627 & ~n28869;
  assign n28985 = ~n17627 & n28954;
  assign n28986 = ~n28984 & ~n28985;
  assign n28987 = pi626 & ~n28986;
  assign n28988 = ~pi641 & ~n28987;
  assign n28989 = ~n28983 & n28988;
  assign n28990 = ~pi789 & ~n28961;
  assign n28991 = ~n28965 & ~n28975;
  assign n28992 = pi789 & ~n28991;
  assign n28993 = ~n28990 & ~n28992;
  assign n28994 = ~pi626 & ~n28993;
  assign n28995 = pi626 & ~n28869;
  assign n28996 = pi641 & ~n28995;
  assign n28997 = ~n28994 & n28996;
  assign n28998 = ~pi1158 & ~n28997;
  assign n28999 = ~n28989 & n28998;
  assign n29000 = pi626 & n28981;
  assign n29001 = ~pi626 & ~n28986;
  assign n29002 = pi641 & ~n29001;
  assign n29003 = ~n29000 & n29002;
  assign n29004 = pi626 & ~n28993;
  assign n29005 = ~pi626 & ~n28869;
  assign n29006 = ~pi641 & ~n29005;
  assign n29007 = ~n29004 & n29006;
  assign n29008 = pi1158 & ~n29007;
  assign n29009 = ~n29003 & n29008;
  assign n29010 = ~n28999 & ~n29009;
  assign n29011 = pi788 & ~n29010;
  assign n29012 = ~n28982 & ~n29011;
  assign n29013 = ~pi628 & n29012;
  assign n29014 = ~n17904 & n28993;
  assign n29015 = n17904 & n28869;
  assign n29016 = ~n29014 & ~n29015;
  assign n29017 = pi628 & ~n29016;
  assign n29018 = ~pi1156 & ~n29017;
  assign n29019 = ~n29013 & n29018;
  assign n29020 = ~n17670 & n28986;
  assign n29021 = n17670 & n28869;
  assign n29022 = ~n29020 & ~n29021;
  assign n29023 = pi628 & ~n29022;
  assign n29024 = ~pi628 & n28869;
  assign n29025 = pi1156 & ~n29024;
  assign n29026 = ~n29023 & n29025;
  assign n29027 = ~pi629 & ~n29026;
  assign n29028 = ~n29019 & n29027;
  assign n29029 = pi628 & n29012;
  assign n29030 = ~pi628 & ~n29016;
  assign n29031 = pi1156 & ~n29030;
  assign n29032 = ~n29029 & n29031;
  assign n29033 = ~pi628 & ~n29022;
  assign n29034 = pi628 & n28869;
  assign n29035 = ~pi1156 & ~n29034;
  assign n29036 = ~n29033 & n29035;
  assign n29037 = pi629 & ~n29036;
  assign n29038 = ~n29032 & n29037;
  assign n29039 = ~n29028 & ~n29038;
  assign n29040 = pi792 & ~n29039;
  assign n29041 = ~pi792 & n29012;
  assign n29042 = ~n29040 & ~n29041;
  assign n29043 = ~pi647 & ~n29042;
  assign n29044 = ~n17698 & ~n29016;
  assign n29045 = n17698 & n28869;
  assign n29046 = ~n29044 & ~n29045;
  assign n29047 = pi647 & ~n29046;
  assign n29048 = ~pi1157 & ~n29047;
  assign n29049 = ~n29043 & n29048;
  assign n29050 = ~pi792 & n29022;
  assign n29051 = ~n29026 & ~n29036;
  assign n29052 = pi792 & ~n29051;
  assign n29053 = ~n29050 & ~n29052;
  assign n29054 = pi647 & n29053;
  assign n29055 = ~pi647 & n28869;
  assign n29056 = pi1157 & ~n29055;
  assign n29057 = ~n29054 & n29056;
  assign n29058 = ~pi630 & ~n29057;
  assign n29059 = ~n29049 & n29058;
  assign n29060 = pi647 & ~n29042;
  assign n29061 = ~pi647 & ~n29046;
  assign n29062 = pi1157 & ~n29061;
  assign n29063 = ~n29060 & n29062;
  assign n29064 = ~pi647 & n29053;
  assign n29065 = pi647 & n28869;
  assign n29066 = ~pi1157 & ~n29065;
  assign n29067 = ~n29064 & n29066;
  assign n29068 = pi630 & ~n29067;
  assign n29069 = ~n29063 & n29068;
  assign n29070 = ~n29059 & ~n29069;
  assign n29071 = pi787 & ~n29070;
  assign n29072 = ~pi787 & ~n29042;
  assign n29073 = ~n29071 & ~n29072;
  assign n29074 = pi644 & ~n29073;
  assign n29075 = ~pi787 & ~n29053;
  assign n29076 = ~n29057 & ~n29067;
  assign n29077 = pi787 & ~n29076;
  assign n29078 = ~n29075 & ~n29077;
  assign n29079 = ~pi644 & n29078;
  assign n29080 = pi715 & ~n29079;
  assign n29081 = ~n29074 & n29080;
  assign n29082 = n17740 & ~n28869;
  assign n29083 = ~n17740 & n29046;
  assign n29084 = ~n29082 & ~n29083;
  assign n29085 = pi644 & n29084;
  assign n29086 = ~pi644 & n28869;
  assign n29087 = ~pi715 & ~n29086;
  assign n29088 = ~n29085 & n29087;
  assign n29089 = pi1160 & ~n29088;
  assign n29090 = ~n29081 & n29089;
  assign n29091 = ~pi644 & ~n29073;
  assign n29092 = pi644 & n29078;
  assign n29093 = ~pi715 & ~n29092;
  assign n29094 = ~n29091 & n29093;
  assign n29095 = ~pi644 & n29084;
  assign n29096 = pi644 & n28869;
  assign n29097 = pi715 & ~n29096;
  assign n29098 = ~n29095 & n29097;
  assign n29099 = ~pi1160 & ~n29098;
  assign n29100 = ~n29094 & n29099;
  assign n29101 = pi790 & ~n29090;
  assign n29102 = ~n29100 & n29101;
  assign n29103 = ~pi790 & n29073;
  assign n29104 = ~po1038 & ~n29103;
  assign n29105 = ~n29102 & n29104;
  assign n29106 = ~pi186 & po1038;
  assign n29107 = ~pi832 & ~n29106;
  assign n29108 = ~n29105 & n29107;
  assign n29109 = ~pi186 & ~n2755;
  assign n29110 = ~pi752 & n16933;
  assign n29111 = ~n29109 & ~n29110;
  assign n29112 = ~n17794 & ~n29111;
  assign n29113 = ~pi785 & ~n29112;
  assign n29114 = ~n17799 & ~n29111;
  assign n29115 = pi1155 & ~n29114;
  assign n29116 = ~n17802 & n29112;
  assign n29117 = ~pi1155 & ~n29116;
  assign n29118 = ~n29115 & ~n29117;
  assign n29119 = pi785 & ~n29118;
  assign n29120 = ~n29113 & ~n29119;
  assign n29121 = ~pi781 & ~n29120;
  assign n29122 = ~n17809 & n29120;
  assign n29123 = pi1154 & ~n29122;
  assign n29124 = ~n17812 & n29120;
  assign n29125 = ~pi1154 & ~n29124;
  assign n29126 = ~n29123 & ~n29125;
  assign n29127 = pi781 & ~n29126;
  assign n29128 = ~n29121 & ~n29127;
  assign n29129 = ~pi789 & ~n29128;
  assign n29130 = pi619 & n29128;
  assign n29131 = ~pi619 & n29109;
  assign n29132 = pi1159 & ~n29131;
  assign n29133 = ~n29130 & n29132;
  assign n29134 = ~pi619 & n29128;
  assign n29135 = pi619 & n29109;
  assign n29136 = ~pi1159 & ~n29135;
  assign n29137 = ~n29134 & n29136;
  assign n29138 = ~n29133 & ~n29137;
  assign n29139 = pi789 & ~n29138;
  assign n29140 = ~n29129 & ~n29139;
  assign n29141 = ~n17904 & n29140;
  assign n29142 = n17904 & n29109;
  assign n29143 = ~n29141 & ~n29142;
  assign n29144 = ~n17698 & ~n29143;
  assign n29145 = n17698 & n29109;
  assign n29146 = ~n29144 & ~n29145;
  assign n29147 = ~n20491 & n29146;
  assign n29148 = pi703 & n17153;
  assign n29149 = ~n29109 & ~n29148;
  assign n29150 = ~pi778 & n29149;
  assign n29151 = ~pi625 & n29148;
  assign n29152 = ~n29149 & ~n29151;
  assign n29153 = pi1153 & ~n29152;
  assign n29154 = ~pi1153 & ~n29109;
  assign n29155 = ~n29151 & n29154;
  assign n29156 = ~n29153 & ~n29155;
  assign n29157 = pi778 & ~n29156;
  assign n29158 = ~n29150 & ~n29157;
  assign n29159 = ~n17780 & n29158;
  assign n29160 = ~n17782 & n29159;
  assign n29161 = ~n17784 & n29160;
  assign n29162 = ~n17916 & n29161;
  assign n29163 = ~n17947 & n29162;
  assign n29164 = ~pi647 & n29163;
  assign n29165 = pi647 & n29109;
  assign n29166 = ~pi1157 & ~n29165;
  assign n29167 = ~n29164 & n29166;
  assign n29168 = pi647 & ~n29163;
  assign n29169 = ~pi647 & ~n29109;
  assign n29170 = ~n29168 & ~n29169;
  assign n29171 = pi1157 & ~n29170;
  assign n29172 = ~n29167 & ~n29171;
  assign n29173 = ~n17739 & ~n29172;
  assign n29174 = ~n29147 & ~n29173;
  assign n29175 = pi787 & ~n29174;
  assign n29176 = ~pi626 & ~n29140;
  assign n29177 = pi626 & ~n29109;
  assign n29178 = n17668 & ~n29177;
  assign n29179 = ~n29176 & n29178;
  assign n29180 = pi626 & ~n29140;
  assign n29181 = ~pi626 & ~n29109;
  assign n29182 = n17667 & ~n29181;
  assign n29183 = ~n29180 & n29182;
  assign n29184 = n17792 & n29161;
  assign n29185 = ~n29179 & ~n29184;
  assign n29186 = ~n29183 & n29185;
  assign n29187 = pi788 & ~n29186;
  assign n29188 = ~n16842 & ~n29149;
  assign n29189 = pi625 & n29188;
  assign n29190 = n29111 & ~n29188;
  assign n29191 = ~n29189 & ~n29190;
  assign n29192 = n29154 & ~n29191;
  assign n29193 = ~pi608 & ~n29153;
  assign n29194 = ~n29192 & n29193;
  assign n29195 = pi1153 & n29111;
  assign n29196 = ~n29189 & n29195;
  assign n29197 = pi608 & ~n29155;
  assign n29198 = ~n29196 & n29197;
  assign n29199 = ~n29194 & ~n29198;
  assign n29200 = pi778 & ~n29199;
  assign n29201 = ~pi778 & ~n29190;
  assign n29202 = ~n29200 & ~n29201;
  assign n29203 = ~pi609 & ~n29202;
  assign n29204 = pi609 & n29158;
  assign n29205 = ~pi1155 & ~n29204;
  assign n29206 = ~n29203 & n29205;
  assign n29207 = ~pi660 & ~n29115;
  assign n29208 = ~n29206 & n29207;
  assign n29209 = pi609 & ~n29202;
  assign n29210 = ~pi609 & n29158;
  assign n29211 = pi1155 & ~n29210;
  assign n29212 = ~n29209 & n29211;
  assign n29213 = pi660 & ~n29117;
  assign n29214 = ~n29212 & n29213;
  assign n29215 = ~n29208 & ~n29214;
  assign n29216 = pi785 & ~n29215;
  assign n29217 = ~pi785 & ~n29202;
  assign n29218 = ~n29216 & ~n29217;
  assign n29219 = ~pi618 & ~n29218;
  assign n29220 = pi618 & n29159;
  assign n29221 = ~pi1154 & ~n29220;
  assign n29222 = ~n29219 & n29221;
  assign n29223 = ~pi627 & ~n29123;
  assign n29224 = ~n29222 & n29223;
  assign n29225 = pi618 & ~n29218;
  assign n29226 = ~pi618 & n29159;
  assign n29227 = pi1154 & ~n29226;
  assign n29228 = ~n29225 & n29227;
  assign n29229 = pi627 & ~n29125;
  assign n29230 = ~n29228 & n29229;
  assign n29231 = ~n29224 & ~n29230;
  assign n29232 = pi781 & ~n29231;
  assign n29233 = ~pi781 & ~n29218;
  assign n29234 = ~n29232 & ~n29233;
  assign n29235 = ~pi619 & ~n29234;
  assign n29236 = pi619 & n29160;
  assign n29237 = ~pi1159 & ~n29236;
  assign n29238 = ~n29235 & n29237;
  assign n29239 = ~pi648 & ~n29133;
  assign n29240 = ~n29238 & n29239;
  assign n29241 = pi619 & ~n29234;
  assign n29242 = ~pi619 & n29160;
  assign n29243 = pi1159 & ~n29242;
  assign n29244 = ~n29241 & n29243;
  assign n29245 = pi648 & ~n29137;
  assign n29246 = ~n29244 & n29245;
  assign n29247 = pi789 & ~n29240;
  assign n29248 = ~n29246 & n29247;
  assign n29249 = ~pi789 & n29234;
  assign n29250 = n17905 & ~n29249;
  assign n29251 = ~n29248 & n29250;
  assign n29252 = ~n29187 & ~n29251;
  assign n29253 = ~n20298 & ~n29252;
  assign n29254 = n17944 & ~n29143;
  assign n29255 = n20786 & n29162;
  assign n29256 = ~n29254 & ~n29255;
  assign n29257 = ~pi629 & ~n29256;
  assign n29258 = n20790 & n29162;
  assign n29259 = n17943 & ~n29143;
  assign n29260 = ~n29258 & ~n29259;
  assign n29261 = pi629 & ~n29260;
  assign n29262 = ~n29257 & ~n29261;
  assign n29263 = pi792 & ~n29262;
  assign n29264 = n20300 & ~n29263;
  assign n29265 = ~n29253 & n29264;
  assign n29266 = ~n29175 & ~n29265;
  assign n29267 = pi644 & n29266;
  assign n29268 = ~pi787 & ~n29163;
  assign n29269 = pi787 & ~n29172;
  assign n29270 = ~n29268 & ~n29269;
  assign n29271 = ~pi644 & n29270;
  assign n29272 = pi715 & ~n29271;
  assign n29273 = ~n29267 & n29272;
  assign n29274 = ~n17740 & ~n29146;
  assign n29275 = n17740 & n29109;
  assign n29276 = ~n29274 & ~n29275;
  assign n29277 = pi644 & ~n29276;
  assign n29278 = ~pi644 & n29109;
  assign n29279 = ~pi715 & ~n29278;
  assign n29280 = ~n29277 & n29279;
  assign n29281 = pi1160 & ~n29280;
  assign n29282 = ~n29273 & n29281;
  assign n29283 = ~pi644 & n29266;
  assign n29284 = pi644 & n29270;
  assign n29285 = ~pi715 & ~n29284;
  assign n29286 = ~n29283 & n29285;
  assign n29287 = ~pi644 & ~n29276;
  assign n29288 = pi644 & n29109;
  assign n29289 = pi715 & ~n29288;
  assign n29290 = ~n29287 & n29289;
  assign n29291 = ~pi1160 & ~n29290;
  assign n29292 = ~n29286 & n29291;
  assign n29293 = ~n29282 & ~n29292;
  assign n29294 = pi790 & ~n29293;
  assign n29295 = ~pi790 & n29266;
  assign n29296 = pi832 & ~n29295;
  assign n29297 = ~n29294 & n29296;
  assign po343 = ~n29108 & ~n29297;
  assign n29299 = pi187 & ~n3268;
  assign n29300 = ~pi770 & ~n19349;
  assign n29301 = ~n20944 & ~n29300;
  assign n29302 = ~pi187 & ~n29301;
  assign n29303 = ~pi187 & ~n19343;
  assign n29304 = ~pi770 & ~n29303;
  assign n29305 = ~n24371 & n29304;
  assign n29306 = ~n29302 & ~n29305;
  assign n29307 = ~pi726 & ~n29306;
  assign n29308 = ~pi187 & n19309;
  assign n29309 = pi187 & n19314;
  assign n29310 = pi770 & ~n19316;
  assign n29311 = ~n29309 & n29310;
  assign n29312 = ~n29308 & n29311;
  assign n29313 = pi187 & n19326;
  assign n29314 = ~pi187 & ~n19334;
  assign n29315 = ~pi770 & ~n29314;
  assign n29316 = ~n29313 & n29315;
  assign n29317 = pi726 & ~n29316;
  assign n29318 = ~n29312 & n29317;
  assign n29319 = n3268 & ~n29318;
  assign n29320 = ~n29307 & n29319;
  assign n29321 = ~n29299 & ~n29320;
  assign n29322 = ~pi625 & n29321;
  assign n29323 = n3268 & n29306;
  assign n29324 = ~n29299 & ~n29323;
  assign n29325 = pi625 & n29324;
  assign n29326 = ~pi1153 & ~n29325;
  assign n29327 = ~n29322 & n29326;
  assign n29328 = ~pi187 & n18060;
  assign n29329 = pi187 & ~n18064;
  assign n29330 = ~pi38 & ~n29329;
  assign n29331 = ~n29328 & n29330;
  assign n29332 = ~pi187 & ~n16968;
  assign n29333 = n17480 & ~n29332;
  assign n29334 = pi726 & ~n29333;
  assign n29335 = ~n29331 & n29334;
  assign n29336 = ~pi187 & ~pi726;
  assign n29337 = ~n17487 & n29336;
  assign n29338 = n3268 & ~n29337;
  assign n29339 = ~n29335 & n29338;
  assign n29340 = ~n29299 & ~n29339;
  assign n29341 = pi625 & n29340;
  assign n29342 = ~pi187 & ~n17494;
  assign n29343 = ~pi625 & n29342;
  assign n29344 = pi1153 & ~n29343;
  assign n29345 = ~n29341 & n29344;
  assign n29346 = ~pi608 & ~n29345;
  assign n29347 = ~n29327 & n29346;
  assign n29348 = pi625 & n29321;
  assign n29349 = ~pi625 & n29324;
  assign n29350 = pi1153 & ~n29349;
  assign n29351 = ~n29348 & n29350;
  assign n29352 = ~pi625 & n29340;
  assign n29353 = pi625 & n29342;
  assign n29354 = ~pi1153 & ~n29353;
  assign n29355 = ~n29352 & n29354;
  assign n29356 = pi608 & ~n29355;
  assign n29357 = ~n29351 & n29356;
  assign n29358 = ~n29347 & ~n29357;
  assign n29359 = pi778 & ~n29358;
  assign n29360 = ~pi778 & n29321;
  assign n29361 = ~n29359 & ~n29360;
  assign n29362 = ~pi609 & ~n29361;
  assign n29363 = ~pi778 & ~n29340;
  assign n29364 = ~n29345 & ~n29355;
  assign n29365 = pi778 & ~n29364;
  assign n29366 = ~n29363 & ~n29365;
  assign n29367 = pi609 & n29366;
  assign n29368 = ~pi1155 & ~n29367;
  assign n29369 = ~n29362 & n29368;
  assign n29370 = ~n17527 & ~n29342;
  assign n29371 = ~n17526 & ~n29324;
  assign n29372 = pi609 & n29371;
  assign n29373 = ~n29370 & ~n29372;
  assign n29374 = pi1155 & ~n29373;
  assign n29375 = ~pi660 & ~n29374;
  assign n29376 = ~n29369 & n29375;
  assign n29377 = pi609 & ~n29361;
  assign n29378 = ~pi609 & n29366;
  assign n29379 = pi1155 & ~n29378;
  assign n29380 = ~n29377 & n29379;
  assign n29381 = ~n17539 & ~n29342;
  assign n29382 = ~pi609 & n29371;
  assign n29383 = ~n29381 & ~n29382;
  assign n29384 = ~pi1155 & ~n29383;
  assign n29385 = pi660 & ~n29384;
  assign n29386 = ~n29380 & n29385;
  assign n29387 = ~n29376 & ~n29386;
  assign n29388 = pi785 & ~n29387;
  assign n29389 = ~pi785 & ~n29361;
  assign n29390 = ~n29388 & ~n29389;
  assign n29391 = ~pi618 & ~n29390;
  assign n29392 = ~n17554 & ~n29366;
  assign n29393 = n17554 & ~n29342;
  assign n29394 = ~n29392 & ~n29393;
  assign n29395 = pi618 & n29394;
  assign n29396 = ~pi1154 & ~n29395;
  assign n29397 = ~n29391 & n29396;
  assign n29398 = n17526 & ~n29342;
  assign n29399 = ~n29371 & ~n29398;
  assign n29400 = ~pi785 & ~n29399;
  assign n29401 = ~n29374 & ~n29384;
  assign n29402 = pi785 & ~n29401;
  assign n29403 = ~n29400 & ~n29402;
  assign n29404 = pi618 & n29403;
  assign n29405 = ~pi618 & n29342;
  assign n29406 = pi1154 & ~n29405;
  assign n29407 = ~n29404 & n29406;
  assign n29408 = ~pi627 & ~n29407;
  assign n29409 = ~n29397 & n29408;
  assign n29410 = pi618 & ~n29390;
  assign n29411 = ~pi618 & n29394;
  assign n29412 = pi1154 & ~n29411;
  assign n29413 = ~n29410 & n29412;
  assign n29414 = ~pi618 & n29403;
  assign n29415 = pi618 & n29342;
  assign n29416 = ~pi1154 & ~n29415;
  assign n29417 = ~n29414 & n29416;
  assign n29418 = pi627 & ~n29417;
  assign n29419 = ~n29413 & n29418;
  assign n29420 = ~n29409 & ~n29419;
  assign n29421 = pi781 & ~n29420;
  assign n29422 = ~pi781 & ~n29390;
  assign n29423 = ~n29421 & ~n29422;
  assign n29424 = ~pi619 & ~n29423;
  assign n29425 = ~n17591 & n29394;
  assign n29426 = n17591 & n29342;
  assign n29427 = ~n29425 & ~n29426;
  assign n29428 = pi619 & ~n29427;
  assign n29429 = ~pi1159 & ~n29428;
  assign n29430 = ~n29424 & n29429;
  assign n29431 = ~pi781 & ~n29403;
  assign n29432 = ~n29407 & ~n29417;
  assign n29433 = pi781 & ~n29432;
  assign n29434 = ~n29431 & ~n29433;
  assign n29435 = pi619 & n29434;
  assign n29436 = ~pi619 & n29342;
  assign n29437 = pi1159 & ~n29436;
  assign n29438 = ~n29435 & n29437;
  assign n29439 = ~pi648 & ~n29438;
  assign n29440 = ~n29430 & n29439;
  assign n29441 = pi619 & ~n29423;
  assign n29442 = ~pi619 & ~n29427;
  assign n29443 = pi1159 & ~n29442;
  assign n29444 = ~n29441 & n29443;
  assign n29445 = ~pi619 & n29434;
  assign n29446 = pi619 & n29342;
  assign n29447 = ~pi1159 & ~n29446;
  assign n29448 = ~n29445 & n29447;
  assign n29449 = pi648 & ~n29448;
  assign n29450 = ~n29444 & n29449;
  assign n29451 = ~n29440 & ~n29450;
  assign n29452 = pi789 & ~n29451;
  assign n29453 = ~pi789 & ~n29423;
  assign n29454 = ~n29452 & ~n29453;
  assign n29455 = ~pi788 & n29454;
  assign n29456 = ~pi626 & n29454;
  assign n29457 = n17627 & ~n29342;
  assign n29458 = ~n17627 & n29427;
  assign n29459 = ~n29457 & ~n29458;
  assign n29460 = pi626 & ~n29459;
  assign n29461 = ~pi641 & ~n29460;
  assign n29462 = ~n29456 & n29461;
  assign n29463 = ~pi789 & ~n29434;
  assign n29464 = ~n29438 & ~n29448;
  assign n29465 = pi789 & ~n29464;
  assign n29466 = ~n29463 & ~n29465;
  assign n29467 = ~pi626 & ~n29466;
  assign n29468 = pi626 & ~n29342;
  assign n29469 = pi641 & ~n29468;
  assign n29470 = ~n29467 & n29469;
  assign n29471 = ~pi1158 & ~n29470;
  assign n29472 = ~n29462 & n29471;
  assign n29473 = pi626 & n29454;
  assign n29474 = ~pi626 & ~n29459;
  assign n29475 = pi641 & ~n29474;
  assign n29476 = ~n29473 & n29475;
  assign n29477 = pi626 & ~n29466;
  assign n29478 = ~pi626 & ~n29342;
  assign n29479 = ~pi641 & ~n29478;
  assign n29480 = ~n29477 & n29479;
  assign n29481 = pi1158 & ~n29480;
  assign n29482 = ~n29476 & n29481;
  assign n29483 = ~n29472 & ~n29482;
  assign n29484 = pi788 & ~n29483;
  assign n29485 = ~n29455 & ~n29484;
  assign n29486 = ~pi628 & n29485;
  assign n29487 = ~n17904 & n29466;
  assign n29488 = n17904 & n29342;
  assign n29489 = ~n29487 & ~n29488;
  assign n29490 = pi628 & ~n29489;
  assign n29491 = ~pi1156 & ~n29490;
  assign n29492 = ~n29486 & n29491;
  assign n29493 = ~n17670 & n29459;
  assign n29494 = n17670 & n29342;
  assign n29495 = ~n29493 & ~n29494;
  assign n29496 = pi628 & ~n29495;
  assign n29497 = ~pi628 & n29342;
  assign n29498 = pi1156 & ~n29497;
  assign n29499 = ~n29496 & n29498;
  assign n29500 = ~pi629 & ~n29499;
  assign n29501 = ~n29492 & n29500;
  assign n29502 = pi628 & n29485;
  assign n29503 = ~pi628 & ~n29489;
  assign n29504 = pi1156 & ~n29503;
  assign n29505 = ~n29502 & n29504;
  assign n29506 = ~pi628 & ~n29495;
  assign n29507 = pi628 & n29342;
  assign n29508 = ~pi1156 & ~n29507;
  assign n29509 = ~n29506 & n29508;
  assign n29510 = pi629 & ~n29509;
  assign n29511 = ~n29505 & n29510;
  assign n29512 = ~n29501 & ~n29511;
  assign n29513 = pi792 & ~n29512;
  assign n29514 = ~pi792 & n29485;
  assign n29515 = ~n29513 & ~n29514;
  assign n29516 = ~pi647 & ~n29515;
  assign n29517 = ~n17698 & ~n29489;
  assign n29518 = n17698 & n29342;
  assign n29519 = ~n29517 & ~n29518;
  assign n29520 = pi647 & ~n29519;
  assign n29521 = ~pi1157 & ~n29520;
  assign n29522 = ~n29516 & n29521;
  assign n29523 = ~pi792 & n29495;
  assign n29524 = ~n29499 & ~n29509;
  assign n29525 = pi792 & ~n29524;
  assign n29526 = ~n29523 & ~n29525;
  assign n29527 = pi647 & n29526;
  assign n29528 = ~pi647 & n29342;
  assign n29529 = pi1157 & ~n29528;
  assign n29530 = ~n29527 & n29529;
  assign n29531 = ~pi630 & ~n29530;
  assign n29532 = ~n29522 & n29531;
  assign n29533 = pi647 & ~n29515;
  assign n29534 = ~pi647 & ~n29519;
  assign n29535 = pi1157 & ~n29534;
  assign n29536 = ~n29533 & n29535;
  assign n29537 = ~pi647 & n29526;
  assign n29538 = pi647 & n29342;
  assign n29539 = ~pi1157 & ~n29538;
  assign n29540 = ~n29537 & n29539;
  assign n29541 = pi630 & ~n29540;
  assign n29542 = ~n29536 & n29541;
  assign n29543 = ~n29532 & ~n29542;
  assign n29544 = pi787 & ~n29543;
  assign n29545 = ~pi787 & ~n29515;
  assign n29546 = ~n29544 & ~n29545;
  assign n29547 = pi644 & ~n29546;
  assign n29548 = ~pi787 & ~n29526;
  assign n29549 = ~n29530 & ~n29540;
  assign n29550 = pi787 & ~n29549;
  assign n29551 = ~n29548 & ~n29550;
  assign n29552 = ~pi644 & n29551;
  assign n29553 = pi715 & ~n29552;
  assign n29554 = ~n29547 & n29553;
  assign n29555 = n17740 & ~n29342;
  assign n29556 = ~n17740 & n29519;
  assign n29557 = ~n29555 & ~n29556;
  assign n29558 = pi644 & n29557;
  assign n29559 = ~pi644 & n29342;
  assign n29560 = ~pi715 & ~n29559;
  assign n29561 = ~n29558 & n29560;
  assign n29562 = pi1160 & ~n29561;
  assign n29563 = ~n29554 & n29562;
  assign n29564 = ~pi644 & ~n29546;
  assign n29565 = pi644 & n29551;
  assign n29566 = ~pi715 & ~n29565;
  assign n29567 = ~n29564 & n29566;
  assign n29568 = ~pi644 & n29557;
  assign n29569 = pi644 & n29342;
  assign n29570 = pi715 & ~n29569;
  assign n29571 = ~n29568 & n29570;
  assign n29572 = ~pi1160 & ~n29571;
  assign n29573 = ~n29567 & n29572;
  assign n29574 = pi790 & ~n29563;
  assign n29575 = ~n29573 & n29574;
  assign n29576 = ~pi790 & n29546;
  assign n29577 = ~po1038 & ~n29576;
  assign n29578 = ~n29575 & n29577;
  assign n29579 = ~pi187 & po1038;
  assign n29580 = ~pi832 & ~n29579;
  assign n29581 = ~n29578 & n29580;
  assign n29582 = ~pi187 & ~n2755;
  assign n29583 = ~pi770 & n16933;
  assign n29584 = ~n29582 & ~n29583;
  assign n29585 = ~n17794 & ~n29584;
  assign n29586 = ~pi785 & ~n29585;
  assign n29587 = ~n17799 & ~n29584;
  assign n29588 = pi1155 & ~n29587;
  assign n29589 = ~n17802 & n29585;
  assign n29590 = ~pi1155 & ~n29589;
  assign n29591 = ~n29588 & ~n29590;
  assign n29592 = pi785 & ~n29591;
  assign n29593 = ~n29586 & ~n29592;
  assign n29594 = ~pi781 & ~n29593;
  assign n29595 = ~n17809 & n29593;
  assign n29596 = pi1154 & ~n29595;
  assign n29597 = ~n17812 & n29593;
  assign n29598 = ~pi1154 & ~n29597;
  assign n29599 = ~n29596 & ~n29598;
  assign n29600 = pi781 & ~n29599;
  assign n29601 = ~n29594 & ~n29600;
  assign n29602 = ~pi789 & ~n29601;
  assign n29603 = pi619 & n29601;
  assign n29604 = ~pi619 & n29582;
  assign n29605 = pi1159 & ~n29604;
  assign n29606 = ~n29603 & n29605;
  assign n29607 = ~pi619 & n29601;
  assign n29608 = pi619 & n29582;
  assign n29609 = ~pi1159 & ~n29608;
  assign n29610 = ~n29607 & n29609;
  assign n29611 = ~n29606 & ~n29610;
  assign n29612 = pi789 & ~n29611;
  assign n29613 = ~n29602 & ~n29612;
  assign n29614 = ~n17904 & n29613;
  assign n29615 = n17904 & n29582;
  assign n29616 = ~n29614 & ~n29615;
  assign n29617 = ~n17698 & ~n29616;
  assign n29618 = n17698 & n29582;
  assign n29619 = ~n29617 & ~n29618;
  assign n29620 = ~n20491 & n29619;
  assign n29621 = pi726 & n17153;
  assign n29622 = ~n29582 & ~n29621;
  assign n29623 = ~pi778 & n29622;
  assign n29624 = ~pi625 & n29621;
  assign n29625 = ~n29622 & ~n29624;
  assign n29626 = pi1153 & ~n29625;
  assign n29627 = ~pi1153 & ~n29582;
  assign n29628 = ~n29624 & n29627;
  assign n29629 = ~n29626 & ~n29628;
  assign n29630 = pi778 & ~n29629;
  assign n29631 = ~n29623 & ~n29630;
  assign n29632 = ~n17780 & n29631;
  assign n29633 = ~n17782 & n29632;
  assign n29634 = ~n17784 & n29633;
  assign n29635 = ~n17916 & n29634;
  assign n29636 = ~n17947 & n29635;
  assign n29637 = ~pi647 & n29636;
  assign n29638 = pi647 & n29582;
  assign n29639 = ~pi1157 & ~n29638;
  assign n29640 = ~n29637 & n29639;
  assign n29641 = pi647 & ~n29636;
  assign n29642 = ~pi647 & ~n29582;
  assign n29643 = ~n29641 & ~n29642;
  assign n29644 = pi1157 & ~n29643;
  assign n29645 = ~n29640 & ~n29644;
  assign n29646 = ~n17739 & ~n29645;
  assign n29647 = ~n29620 & ~n29646;
  assign n29648 = pi787 & ~n29647;
  assign n29649 = ~pi626 & ~n29613;
  assign n29650 = pi626 & ~n29582;
  assign n29651 = n17668 & ~n29650;
  assign n29652 = ~n29649 & n29651;
  assign n29653 = pi626 & ~n29613;
  assign n29654 = ~pi626 & ~n29582;
  assign n29655 = n17667 & ~n29654;
  assign n29656 = ~n29653 & n29655;
  assign n29657 = n17792 & n29634;
  assign n29658 = ~n29652 & ~n29657;
  assign n29659 = ~n29656 & n29658;
  assign n29660 = pi788 & ~n29659;
  assign n29661 = ~n16842 & ~n29622;
  assign n29662 = pi625 & n29661;
  assign n29663 = n29584 & ~n29661;
  assign n29664 = ~n29662 & ~n29663;
  assign n29665 = n29627 & ~n29664;
  assign n29666 = ~pi608 & ~n29626;
  assign n29667 = ~n29665 & n29666;
  assign n29668 = pi1153 & n29584;
  assign n29669 = ~n29662 & n29668;
  assign n29670 = pi608 & ~n29628;
  assign n29671 = ~n29669 & n29670;
  assign n29672 = ~n29667 & ~n29671;
  assign n29673 = pi778 & ~n29672;
  assign n29674 = ~pi778 & ~n29663;
  assign n29675 = ~n29673 & ~n29674;
  assign n29676 = ~pi609 & ~n29675;
  assign n29677 = pi609 & n29631;
  assign n29678 = ~pi1155 & ~n29677;
  assign n29679 = ~n29676 & n29678;
  assign n29680 = ~pi660 & ~n29588;
  assign n29681 = ~n29679 & n29680;
  assign n29682 = pi609 & ~n29675;
  assign n29683 = ~pi609 & n29631;
  assign n29684 = pi1155 & ~n29683;
  assign n29685 = ~n29682 & n29684;
  assign n29686 = pi660 & ~n29590;
  assign n29687 = ~n29685 & n29686;
  assign n29688 = ~n29681 & ~n29687;
  assign n29689 = pi785 & ~n29688;
  assign n29690 = ~pi785 & ~n29675;
  assign n29691 = ~n29689 & ~n29690;
  assign n29692 = ~pi618 & ~n29691;
  assign n29693 = pi618 & n29632;
  assign n29694 = ~pi1154 & ~n29693;
  assign n29695 = ~n29692 & n29694;
  assign n29696 = ~pi627 & ~n29596;
  assign n29697 = ~n29695 & n29696;
  assign n29698 = pi618 & ~n29691;
  assign n29699 = ~pi618 & n29632;
  assign n29700 = pi1154 & ~n29699;
  assign n29701 = ~n29698 & n29700;
  assign n29702 = pi627 & ~n29598;
  assign n29703 = ~n29701 & n29702;
  assign n29704 = ~n29697 & ~n29703;
  assign n29705 = pi781 & ~n29704;
  assign n29706 = ~pi781 & ~n29691;
  assign n29707 = ~n29705 & ~n29706;
  assign n29708 = ~pi619 & ~n29707;
  assign n29709 = pi619 & n29633;
  assign n29710 = ~pi1159 & ~n29709;
  assign n29711 = ~n29708 & n29710;
  assign n29712 = ~pi648 & ~n29606;
  assign n29713 = ~n29711 & n29712;
  assign n29714 = pi619 & ~n29707;
  assign n29715 = ~pi619 & n29633;
  assign n29716 = pi1159 & ~n29715;
  assign n29717 = ~n29714 & n29716;
  assign n29718 = pi648 & ~n29610;
  assign n29719 = ~n29717 & n29718;
  assign n29720 = pi789 & ~n29713;
  assign n29721 = ~n29719 & n29720;
  assign n29722 = ~pi789 & n29707;
  assign n29723 = n17905 & ~n29722;
  assign n29724 = ~n29721 & n29723;
  assign n29725 = ~n29660 & ~n29724;
  assign n29726 = ~n20298 & ~n29725;
  assign n29727 = n17944 & ~n29616;
  assign n29728 = n20786 & n29635;
  assign n29729 = ~n29727 & ~n29728;
  assign n29730 = ~pi629 & ~n29729;
  assign n29731 = n20790 & n29635;
  assign n29732 = n17943 & ~n29616;
  assign n29733 = ~n29731 & ~n29732;
  assign n29734 = pi629 & ~n29733;
  assign n29735 = ~n29730 & ~n29734;
  assign n29736 = pi792 & ~n29735;
  assign n29737 = n20300 & ~n29736;
  assign n29738 = ~n29726 & n29737;
  assign n29739 = ~n29648 & ~n29738;
  assign n29740 = pi644 & n29739;
  assign n29741 = ~pi787 & ~n29636;
  assign n29742 = pi787 & ~n29645;
  assign n29743 = ~n29741 & ~n29742;
  assign n29744 = ~pi644 & n29743;
  assign n29745 = pi715 & ~n29744;
  assign n29746 = ~n29740 & n29745;
  assign n29747 = ~n17740 & ~n29619;
  assign n29748 = n17740 & n29582;
  assign n29749 = ~n29747 & ~n29748;
  assign n29750 = pi644 & ~n29749;
  assign n29751 = ~pi644 & n29582;
  assign n29752 = ~pi715 & ~n29751;
  assign n29753 = ~n29750 & n29752;
  assign n29754 = pi1160 & ~n29753;
  assign n29755 = ~n29746 & n29754;
  assign n29756 = ~pi644 & n29739;
  assign n29757 = pi644 & n29743;
  assign n29758 = ~pi715 & ~n29757;
  assign n29759 = ~n29756 & n29758;
  assign n29760 = ~pi644 & ~n29749;
  assign n29761 = pi644 & n29582;
  assign n29762 = pi715 & ~n29761;
  assign n29763 = ~n29760 & n29762;
  assign n29764 = ~pi1160 & ~n29763;
  assign n29765 = ~n29759 & n29764;
  assign n29766 = ~n29755 & ~n29765;
  assign n29767 = pi790 & ~n29766;
  assign n29768 = ~pi790 & n29739;
  assign n29769 = pi832 & ~n29768;
  assign n29770 = ~n29767 & n29769;
  assign po344 = ~n29581 & ~n29770;
  assign n29772 = pi188 & ~n3268;
  assign n29773 = ~pi768 & ~n19349;
  assign n29774 = ~n22269 & ~n29773;
  assign n29775 = ~pi188 & ~n29774;
  assign n29776 = ~pi188 & ~n19343;
  assign n29777 = ~pi768 & ~n29776;
  assign n29778 = ~n24371 & n29777;
  assign n29779 = ~n29775 & ~n29778;
  assign n29780 = ~pi705 & ~n29779;
  assign n29781 = ~pi188 & n19309;
  assign n29782 = pi188 & n19314;
  assign n29783 = pi768 & ~n19316;
  assign n29784 = ~n29782 & n29783;
  assign n29785 = ~n29781 & n29784;
  assign n29786 = pi188 & n19326;
  assign n29787 = ~pi188 & ~n19334;
  assign n29788 = ~pi768 & ~n29787;
  assign n29789 = ~n29786 & n29788;
  assign n29790 = pi705 & ~n29789;
  assign n29791 = ~n29785 & n29790;
  assign n29792 = n3268 & ~n29791;
  assign n29793 = ~n29780 & n29792;
  assign n29794 = ~n29772 & ~n29793;
  assign n29795 = ~pi625 & n29794;
  assign n29796 = n3268 & n29779;
  assign n29797 = ~n29772 & ~n29796;
  assign n29798 = pi625 & n29797;
  assign n29799 = ~pi1153 & ~n29798;
  assign n29800 = ~n29795 & n29799;
  assign n29801 = ~pi188 & n18060;
  assign n29802 = pi188 & ~n18064;
  assign n29803 = ~pi38 & ~n29802;
  assign n29804 = ~n29801 & n29803;
  assign n29805 = ~pi188 & ~n16968;
  assign n29806 = n17480 & ~n29805;
  assign n29807 = pi705 & ~n29806;
  assign n29808 = ~n29804 & n29807;
  assign n29809 = ~pi188 & ~pi705;
  assign n29810 = ~n17487 & n29809;
  assign n29811 = n3268 & ~n29810;
  assign n29812 = ~n29808 & n29811;
  assign n29813 = ~n29772 & ~n29812;
  assign n29814 = pi625 & n29813;
  assign n29815 = ~pi188 & ~n17494;
  assign n29816 = ~pi625 & n29815;
  assign n29817 = pi1153 & ~n29816;
  assign n29818 = ~n29814 & n29817;
  assign n29819 = ~pi608 & ~n29818;
  assign n29820 = ~n29800 & n29819;
  assign n29821 = pi625 & n29794;
  assign n29822 = ~pi625 & n29797;
  assign n29823 = pi1153 & ~n29822;
  assign n29824 = ~n29821 & n29823;
  assign n29825 = ~pi625 & n29813;
  assign n29826 = pi625 & n29815;
  assign n29827 = ~pi1153 & ~n29826;
  assign n29828 = ~n29825 & n29827;
  assign n29829 = pi608 & ~n29828;
  assign n29830 = ~n29824 & n29829;
  assign n29831 = ~n29820 & ~n29830;
  assign n29832 = pi778 & ~n29831;
  assign n29833 = ~pi778 & n29794;
  assign n29834 = ~n29832 & ~n29833;
  assign n29835 = ~pi609 & ~n29834;
  assign n29836 = ~pi778 & ~n29813;
  assign n29837 = ~n29818 & ~n29828;
  assign n29838 = pi778 & ~n29837;
  assign n29839 = ~n29836 & ~n29838;
  assign n29840 = pi609 & n29839;
  assign n29841 = ~pi1155 & ~n29840;
  assign n29842 = ~n29835 & n29841;
  assign n29843 = ~n17527 & ~n29815;
  assign n29844 = ~n17526 & ~n29797;
  assign n29845 = pi609 & n29844;
  assign n29846 = ~n29843 & ~n29845;
  assign n29847 = pi1155 & ~n29846;
  assign n29848 = ~pi660 & ~n29847;
  assign n29849 = ~n29842 & n29848;
  assign n29850 = pi609 & ~n29834;
  assign n29851 = ~pi609 & n29839;
  assign n29852 = pi1155 & ~n29851;
  assign n29853 = ~n29850 & n29852;
  assign n29854 = ~n17539 & ~n29815;
  assign n29855 = ~pi609 & n29844;
  assign n29856 = ~n29854 & ~n29855;
  assign n29857 = ~pi1155 & ~n29856;
  assign n29858 = pi660 & ~n29857;
  assign n29859 = ~n29853 & n29858;
  assign n29860 = ~n29849 & ~n29859;
  assign n29861 = pi785 & ~n29860;
  assign n29862 = ~pi785 & ~n29834;
  assign n29863 = ~n29861 & ~n29862;
  assign n29864 = ~pi618 & ~n29863;
  assign n29865 = ~n17554 & ~n29839;
  assign n29866 = n17554 & ~n29815;
  assign n29867 = ~n29865 & ~n29866;
  assign n29868 = pi618 & n29867;
  assign n29869 = ~pi1154 & ~n29868;
  assign n29870 = ~n29864 & n29869;
  assign n29871 = n17526 & ~n29815;
  assign n29872 = ~n29844 & ~n29871;
  assign n29873 = ~pi785 & ~n29872;
  assign n29874 = ~n29847 & ~n29857;
  assign n29875 = pi785 & ~n29874;
  assign n29876 = ~n29873 & ~n29875;
  assign n29877 = pi618 & n29876;
  assign n29878 = ~pi618 & n29815;
  assign n29879 = pi1154 & ~n29878;
  assign n29880 = ~n29877 & n29879;
  assign n29881 = ~pi627 & ~n29880;
  assign n29882 = ~n29870 & n29881;
  assign n29883 = pi618 & ~n29863;
  assign n29884 = ~pi618 & n29867;
  assign n29885 = pi1154 & ~n29884;
  assign n29886 = ~n29883 & n29885;
  assign n29887 = ~pi618 & n29876;
  assign n29888 = pi618 & n29815;
  assign n29889 = ~pi1154 & ~n29888;
  assign n29890 = ~n29887 & n29889;
  assign n29891 = pi627 & ~n29890;
  assign n29892 = ~n29886 & n29891;
  assign n29893 = ~n29882 & ~n29892;
  assign n29894 = pi781 & ~n29893;
  assign n29895 = ~pi781 & ~n29863;
  assign n29896 = ~n29894 & ~n29895;
  assign n29897 = ~pi619 & ~n29896;
  assign n29898 = ~n17591 & n29867;
  assign n29899 = n17591 & n29815;
  assign n29900 = ~n29898 & ~n29899;
  assign n29901 = pi619 & ~n29900;
  assign n29902 = ~pi1159 & ~n29901;
  assign n29903 = ~n29897 & n29902;
  assign n29904 = ~pi781 & ~n29876;
  assign n29905 = ~n29880 & ~n29890;
  assign n29906 = pi781 & ~n29905;
  assign n29907 = ~n29904 & ~n29906;
  assign n29908 = pi619 & n29907;
  assign n29909 = ~pi619 & n29815;
  assign n29910 = pi1159 & ~n29909;
  assign n29911 = ~n29908 & n29910;
  assign n29912 = ~pi648 & ~n29911;
  assign n29913 = ~n29903 & n29912;
  assign n29914 = pi619 & ~n29896;
  assign n29915 = ~pi619 & ~n29900;
  assign n29916 = pi1159 & ~n29915;
  assign n29917 = ~n29914 & n29916;
  assign n29918 = ~pi619 & n29907;
  assign n29919 = pi619 & n29815;
  assign n29920 = ~pi1159 & ~n29919;
  assign n29921 = ~n29918 & n29920;
  assign n29922 = pi648 & ~n29921;
  assign n29923 = ~n29917 & n29922;
  assign n29924 = ~n29913 & ~n29923;
  assign n29925 = pi789 & ~n29924;
  assign n29926 = ~pi789 & ~n29896;
  assign n29927 = ~n29925 & ~n29926;
  assign n29928 = ~pi788 & n29927;
  assign n29929 = ~pi626 & n29927;
  assign n29930 = n17627 & ~n29815;
  assign n29931 = ~n17627 & n29900;
  assign n29932 = ~n29930 & ~n29931;
  assign n29933 = pi626 & ~n29932;
  assign n29934 = ~pi641 & ~n29933;
  assign n29935 = ~n29929 & n29934;
  assign n29936 = ~pi789 & ~n29907;
  assign n29937 = ~n29911 & ~n29921;
  assign n29938 = pi789 & ~n29937;
  assign n29939 = ~n29936 & ~n29938;
  assign n29940 = ~pi626 & ~n29939;
  assign n29941 = pi626 & ~n29815;
  assign n29942 = pi641 & ~n29941;
  assign n29943 = ~n29940 & n29942;
  assign n29944 = ~pi1158 & ~n29943;
  assign n29945 = ~n29935 & n29944;
  assign n29946 = pi626 & n29927;
  assign n29947 = ~pi626 & ~n29932;
  assign n29948 = pi641 & ~n29947;
  assign n29949 = ~n29946 & n29948;
  assign n29950 = pi626 & ~n29939;
  assign n29951 = ~pi626 & ~n29815;
  assign n29952 = ~pi641 & ~n29951;
  assign n29953 = ~n29950 & n29952;
  assign n29954 = pi1158 & ~n29953;
  assign n29955 = ~n29949 & n29954;
  assign n29956 = ~n29945 & ~n29955;
  assign n29957 = pi788 & ~n29956;
  assign n29958 = ~n29928 & ~n29957;
  assign n29959 = ~pi628 & n29958;
  assign n29960 = ~n17904 & n29939;
  assign n29961 = n17904 & n29815;
  assign n29962 = ~n29960 & ~n29961;
  assign n29963 = pi628 & ~n29962;
  assign n29964 = ~pi1156 & ~n29963;
  assign n29965 = ~n29959 & n29964;
  assign n29966 = ~n17670 & n29932;
  assign n29967 = n17670 & n29815;
  assign n29968 = ~n29966 & ~n29967;
  assign n29969 = pi628 & ~n29968;
  assign n29970 = ~pi628 & n29815;
  assign n29971 = pi1156 & ~n29970;
  assign n29972 = ~n29969 & n29971;
  assign n29973 = ~pi629 & ~n29972;
  assign n29974 = ~n29965 & n29973;
  assign n29975 = pi628 & n29958;
  assign n29976 = ~pi628 & ~n29962;
  assign n29977 = pi1156 & ~n29976;
  assign n29978 = ~n29975 & n29977;
  assign n29979 = ~pi628 & ~n29968;
  assign n29980 = pi628 & n29815;
  assign n29981 = ~pi1156 & ~n29980;
  assign n29982 = ~n29979 & n29981;
  assign n29983 = pi629 & ~n29982;
  assign n29984 = ~n29978 & n29983;
  assign n29985 = ~n29974 & ~n29984;
  assign n29986 = pi792 & ~n29985;
  assign n29987 = ~pi792 & n29958;
  assign n29988 = ~n29986 & ~n29987;
  assign n29989 = ~pi647 & ~n29988;
  assign n29990 = ~n17698 & ~n29962;
  assign n29991 = n17698 & n29815;
  assign n29992 = ~n29990 & ~n29991;
  assign n29993 = pi647 & ~n29992;
  assign n29994 = ~pi1157 & ~n29993;
  assign n29995 = ~n29989 & n29994;
  assign n29996 = ~pi792 & n29968;
  assign n29997 = ~n29972 & ~n29982;
  assign n29998 = pi792 & ~n29997;
  assign n29999 = ~n29996 & ~n29998;
  assign n30000 = pi647 & n29999;
  assign n30001 = ~pi647 & n29815;
  assign n30002 = pi1157 & ~n30001;
  assign n30003 = ~n30000 & n30002;
  assign n30004 = ~pi630 & ~n30003;
  assign n30005 = ~n29995 & n30004;
  assign n30006 = pi647 & ~n29988;
  assign n30007 = ~pi647 & ~n29992;
  assign n30008 = pi1157 & ~n30007;
  assign n30009 = ~n30006 & n30008;
  assign n30010 = ~pi647 & n29999;
  assign n30011 = pi647 & n29815;
  assign n30012 = ~pi1157 & ~n30011;
  assign n30013 = ~n30010 & n30012;
  assign n30014 = pi630 & ~n30013;
  assign n30015 = ~n30009 & n30014;
  assign n30016 = ~n30005 & ~n30015;
  assign n30017 = pi787 & ~n30016;
  assign n30018 = ~pi787 & ~n29988;
  assign n30019 = ~n30017 & ~n30018;
  assign n30020 = pi644 & ~n30019;
  assign n30021 = ~pi787 & ~n29999;
  assign n30022 = ~n30003 & ~n30013;
  assign n30023 = pi787 & ~n30022;
  assign n30024 = ~n30021 & ~n30023;
  assign n30025 = ~pi644 & n30024;
  assign n30026 = pi715 & ~n30025;
  assign n30027 = ~n30020 & n30026;
  assign n30028 = n17740 & ~n29815;
  assign n30029 = ~n17740 & n29992;
  assign n30030 = ~n30028 & ~n30029;
  assign n30031 = pi644 & n30030;
  assign n30032 = ~pi644 & n29815;
  assign n30033 = ~pi715 & ~n30032;
  assign n30034 = ~n30031 & n30033;
  assign n30035 = pi1160 & ~n30034;
  assign n30036 = ~n30027 & n30035;
  assign n30037 = ~pi644 & ~n30019;
  assign n30038 = pi644 & n30024;
  assign n30039 = ~pi715 & ~n30038;
  assign n30040 = ~n30037 & n30039;
  assign n30041 = ~pi644 & n30030;
  assign n30042 = pi644 & n29815;
  assign n30043 = pi715 & ~n30042;
  assign n30044 = ~n30041 & n30043;
  assign n30045 = ~pi1160 & ~n30044;
  assign n30046 = ~n30040 & n30045;
  assign n30047 = pi790 & ~n30036;
  assign n30048 = ~n30046 & n30047;
  assign n30049 = ~pi790 & n30019;
  assign n30050 = ~po1038 & ~n30049;
  assign n30051 = ~n30048 & n30050;
  assign n30052 = ~pi188 & po1038;
  assign n30053 = ~pi832 & ~n30052;
  assign n30054 = ~n30051 & n30053;
  assign n30055 = ~pi188 & ~n2755;
  assign n30056 = ~pi768 & n16933;
  assign n30057 = ~n30055 & ~n30056;
  assign n30058 = ~n17794 & ~n30057;
  assign n30059 = ~pi785 & ~n30058;
  assign n30060 = ~n17799 & ~n30057;
  assign n30061 = pi1155 & ~n30060;
  assign n30062 = ~n17802 & n30058;
  assign n30063 = ~pi1155 & ~n30062;
  assign n30064 = ~n30061 & ~n30063;
  assign n30065 = pi785 & ~n30064;
  assign n30066 = ~n30059 & ~n30065;
  assign n30067 = ~pi781 & ~n30066;
  assign n30068 = ~n17809 & n30066;
  assign n30069 = pi1154 & ~n30068;
  assign n30070 = ~n17812 & n30066;
  assign n30071 = ~pi1154 & ~n30070;
  assign n30072 = ~n30069 & ~n30071;
  assign n30073 = pi781 & ~n30072;
  assign n30074 = ~n30067 & ~n30073;
  assign n30075 = ~pi789 & ~n30074;
  assign n30076 = pi619 & n30074;
  assign n30077 = ~pi619 & n30055;
  assign n30078 = pi1159 & ~n30077;
  assign n30079 = ~n30076 & n30078;
  assign n30080 = ~pi619 & n30074;
  assign n30081 = pi619 & n30055;
  assign n30082 = ~pi1159 & ~n30081;
  assign n30083 = ~n30080 & n30082;
  assign n30084 = ~n30079 & ~n30083;
  assign n30085 = pi789 & ~n30084;
  assign n30086 = ~n30075 & ~n30085;
  assign n30087 = ~n17904 & n30086;
  assign n30088 = n17904 & n30055;
  assign n30089 = ~n30087 & ~n30088;
  assign n30090 = ~n17698 & ~n30089;
  assign n30091 = n17698 & n30055;
  assign n30092 = ~n30090 & ~n30091;
  assign n30093 = ~n20491 & n30092;
  assign n30094 = pi705 & n17153;
  assign n30095 = ~n30055 & ~n30094;
  assign n30096 = ~pi778 & n30095;
  assign n30097 = ~pi625 & n30094;
  assign n30098 = ~n30095 & ~n30097;
  assign n30099 = pi1153 & ~n30098;
  assign n30100 = ~pi1153 & ~n30055;
  assign n30101 = ~n30097 & n30100;
  assign n30102 = ~n30099 & ~n30101;
  assign n30103 = pi778 & ~n30102;
  assign n30104 = ~n30096 & ~n30103;
  assign n30105 = ~n17780 & n30104;
  assign n30106 = ~n17782 & n30105;
  assign n30107 = ~n17784 & n30106;
  assign n30108 = ~n17916 & n30107;
  assign n30109 = ~n17947 & n30108;
  assign n30110 = ~pi647 & n30109;
  assign n30111 = pi647 & n30055;
  assign n30112 = ~pi1157 & ~n30111;
  assign n30113 = ~n30110 & n30112;
  assign n30114 = pi647 & ~n30109;
  assign n30115 = ~pi647 & ~n30055;
  assign n30116 = ~n30114 & ~n30115;
  assign n30117 = pi1157 & ~n30116;
  assign n30118 = ~n30113 & ~n30117;
  assign n30119 = ~n17739 & ~n30118;
  assign n30120 = ~n30093 & ~n30119;
  assign n30121 = pi787 & ~n30120;
  assign n30122 = ~pi626 & ~n30086;
  assign n30123 = pi626 & ~n30055;
  assign n30124 = n17668 & ~n30123;
  assign n30125 = ~n30122 & n30124;
  assign n30126 = pi626 & ~n30086;
  assign n30127 = ~pi626 & ~n30055;
  assign n30128 = n17667 & ~n30127;
  assign n30129 = ~n30126 & n30128;
  assign n30130 = n17792 & n30107;
  assign n30131 = ~n30125 & ~n30130;
  assign n30132 = ~n30129 & n30131;
  assign n30133 = pi788 & ~n30132;
  assign n30134 = ~n16842 & ~n30095;
  assign n30135 = pi625 & n30134;
  assign n30136 = n30057 & ~n30134;
  assign n30137 = ~n30135 & ~n30136;
  assign n30138 = n30100 & ~n30137;
  assign n30139 = ~pi608 & ~n30099;
  assign n30140 = ~n30138 & n30139;
  assign n30141 = pi1153 & n30057;
  assign n30142 = ~n30135 & n30141;
  assign n30143 = pi608 & ~n30101;
  assign n30144 = ~n30142 & n30143;
  assign n30145 = ~n30140 & ~n30144;
  assign n30146 = pi778 & ~n30145;
  assign n30147 = ~pi778 & ~n30136;
  assign n30148 = ~n30146 & ~n30147;
  assign n30149 = ~pi609 & ~n30148;
  assign n30150 = pi609 & n30104;
  assign n30151 = ~pi1155 & ~n30150;
  assign n30152 = ~n30149 & n30151;
  assign n30153 = ~pi660 & ~n30061;
  assign n30154 = ~n30152 & n30153;
  assign n30155 = pi609 & ~n30148;
  assign n30156 = ~pi609 & n30104;
  assign n30157 = pi1155 & ~n30156;
  assign n30158 = ~n30155 & n30157;
  assign n30159 = pi660 & ~n30063;
  assign n30160 = ~n30158 & n30159;
  assign n30161 = ~n30154 & ~n30160;
  assign n30162 = pi785 & ~n30161;
  assign n30163 = ~pi785 & ~n30148;
  assign n30164 = ~n30162 & ~n30163;
  assign n30165 = ~pi618 & ~n30164;
  assign n30166 = pi618 & n30105;
  assign n30167 = ~pi1154 & ~n30166;
  assign n30168 = ~n30165 & n30167;
  assign n30169 = ~pi627 & ~n30069;
  assign n30170 = ~n30168 & n30169;
  assign n30171 = pi618 & ~n30164;
  assign n30172 = ~pi618 & n30105;
  assign n30173 = pi1154 & ~n30172;
  assign n30174 = ~n30171 & n30173;
  assign n30175 = pi627 & ~n30071;
  assign n30176 = ~n30174 & n30175;
  assign n30177 = ~n30170 & ~n30176;
  assign n30178 = pi781 & ~n30177;
  assign n30179 = ~pi781 & ~n30164;
  assign n30180 = ~n30178 & ~n30179;
  assign n30181 = ~pi619 & ~n30180;
  assign n30182 = pi619 & n30106;
  assign n30183 = ~pi1159 & ~n30182;
  assign n30184 = ~n30181 & n30183;
  assign n30185 = ~pi648 & ~n30079;
  assign n30186 = ~n30184 & n30185;
  assign n30187 = pi619 & ~n30180;
  assign n30188 = ~pi619 & n30106;
  assign n30189 = pi1159 & ~n30188;
  assign n30190 = ~n30187 & n30189;
  assign n30191 = pi648 & ~n30083;
  assign n30192 = ~n30190 & n30191;
  assign n30193 = pi789 & ~n30186;
  assign n30194 = ~n30192 & n30193;
  assign n30195 = ~pi789 & n30180;
  assign n30196 = n17905 & ~n30195;
  assign n30197 = ~n30194 & n30196;
  assign n30198 = ~n30133 & ~n30197;
  assign n30199 = ~n20298 & ~n30198;
  assign n30200 = n17944 & ~n30089;
  assign n30201 = n20786 & n30108;
  assign n30202 = ~n30200 & ~n30201;
  assign n30203 = ~pi629 & ~n30202;
  assign n30204 = n20790 & n30108;
  assign n30205 = n17943 & ~n30089;
  assign n30206 = ~n30204 & ~n30205;
  assign n30207 = pi629 & ~n30206;
  assign n30208 = ~n30203 & ~n30207;
  assign n30209 = pi792 & ~n30208;
  assign n30210 = n20300 & ~n30209;
  assign n30211 = ~n30199 & n30210;
  assign n30212 = ~n30121 & ~n30211;
  assign n30213 = pi644 & n30212;
  assign n30214 = ~pi787 & ~n30109;
  assign n30215 = pi787 & ~n30118;
  assign n30216 = ~n30214 & ~n30215;
  assign n30217 = ~pi644 & n30216;
  assign n30218 = pi715 & ~n30217;
  assign n30219 = ~n30213 & n30218;
  assign n30220 = ~n17740 & ~n30092;
  assign n30221 = n17740 & n30055;
  assign n30222 = ~n30220 & ~n30221;
  assign n30223 = pi644 & ~n30222;
  assign n30224 = ~pi644 & n30055;
  assign n30225 = ~pi715 & ~n30224;
  assign n30226 = ~n30223 & n30225;
  assign n30227 = pi1160 & ~n30226;
  assign n30228 = ~n30219 & n30227;
  assign n30229 = ~pi644 & n30212;
  assign n30230 = pi644 & n30216;
  assign n30231 = ~pi715 & ~n30230;
  assign n30232 = ~n30229 & n30231;
  assign n30233 = ~pi644 & ~n30222;
  assign n30234 = pi644 & n30055;
  assign n30235 = pi715 & ~n30234;
  assign n30236 = ~n30233 & n30235;
  assign n30237 = ~pi1160 & ~n30236;
  assign n30238 = ~n30232 & n30237;
  assign n30239 = ~n30228 & ~n30238;
  assign n30240 = pi790 & ~n30239;
  assign n30241 = ~pi790 & n30212;
  assign n30242 = pi832 & ~n30241;
  assign n30243 = ~n30240 & n30242;
  assign po345 = ~n30054 & ~n30243;
  assign n30245 = pi189 & ~n3268;
  assign n30246 = pi772 & n16905;
  assign n30247 = ~n22162 & ~n30246;
  assign n30248 = pi39 & ~n30247;
  assign n30249 = pi772 & n16839;
  assign n30250 = ~pi772 & n16655;
  assign n30251 = ~pi39 & ~n30250;
  assign n30252 = ~n30249 & n30251;
  assign n30253 = ~n30248 & ~n30252;
  assign n30254 = pi189 & ~n30253;
  assign n30255 = ~pi189 & pi772;
  assign n30256 = n16963 & n30255;
  assign n30257 = ~n30254 & ~n30256;
  assign n30258 = ~pi38 & ~n30257;
  assign n30259 = ~pi189 & ~n16968;
  assign n30260 = pi772 & n16842;
  assign n30261 = n16968 & ~n30260;
  assign n30262 = pi38 & ~n30259;
  assign n30263 = ~n30261 & n30262;
  assign n30264 = ~n30258 & ~n30263;
  assign n30265 = ~pi727 & n30264;
  assign n30266 = pi189 & ~n17074;
  assign n30267 = ~pi189 & ~n17166;
  assign n30268 = ~pi772 & ~n30267;
  assign n30269 = ~n30266 & n30268;
  assign n30270 = ~pi189 & ~n17233;
  assign n30271 = pi189 & n17295;
  assign n30272 = pi772 & ~n30271;
  assign n30273 = ~n30270 & n30272;
  assign n30274 = pi39 & ~n30273;
  assign n30275 = ~n30269 & n30274;
  assign n30276 = ~pi189 & ~n17340;
  assign n30277 = pi189 & ~n17317;
  assign n30278 = ~pi772 & ~n30276;
  assign n30279 = ~n30277 & n30278;
  assign n30280 = pi189 & n17344;
  assign n30281 = ~pi189 & n17351;
  assign n30282 = pi772 & ~n30281;
  assign n30283 = ~n30280 & n30282;
  assign n30284 = ~pi39 & ~n30283;
  assign n30285 = ~n30279 & n30284;
  assign n30286 = ~pi38 & ~n30285;
  assign n30287 = ~n30275 & n30286;
  assign n30288 = pi727 & ~n19316;
  assign n30289 = ~n30263 & n30288;
  assign n30290 = ~n30287 & n30289;
  assign n30291 = n3268 & ~n30290;
  assign n30292 = ~n30265 & n30291;
  assign n30293 = ~n30245 & ~n30292;
  assign n30294 = ~pi625 & n30293;
  assign n30295 = n3268 & ~n30264;
  assign n30296 = ~n30245 & ~n30295;
  assign n30297 = pi625 & n30296;
  assign n30298 = ~pi1153 & ~n30297;
  assign n30299 = ~n30294 & n30298;
  assign n30300 = pi189 & ~n17494;
  assign n30301 = pi727 & n3268;
  assign n30302 = ~n30300 & ~n30301;
  assign n30303 = pi189 & ~n18060;
  assign n30304 = ~pi189 & n18064;
  assign n30305 = ~pi38 & ~n30304;
  assign n30306 = ~n30303 & n30305;
  assign n30307 = n19892 & ~n30259;
  assign n30308 = n30301 & ~n30307;
  assign n30309 = ~n30306 & n30308;
  assign n30310 = ~n30302 & ~n30309;
  assign n30311 = pi625 & ~n30310;
  assign n30312 = ~pi625 & ~n30300;
  assign n30313 = pi1153 & ~n30312;
  assign n30314 = ~n30311 & n30313;
  assign n30315 = ~pi608 & ~n30314;
  assign n30316 = ~n30299 & n30315;
  assign n30317 = pi625 & n30293;
  assign n30318 = ~pi625 & n30296;
  assign n30319 = pi1153 & ~n30318;
  assign n30320 = ~n30317 & n30319;
  assign n30321 = ~pi625 & ~n30310;
  assign n30322 = pi625 & ~n30300;
  assign n30323 = ~pi1153 & ~n30322;
  assign n30324 = ~n30321 & n30323;
  assign n30325 = pi608 & ~n30324;
  assign n30326 = ~n30320 & n30325;
  assign n30327 = ~n30316 & ~n30326;
  assign n30328 = pi778 & ~n30327;
  assign n30329 = ~pi778 & n30293;
  assign n30330 = ~n30328 & ~n30329;
  assign n30331 = ~pi609 & ~n30330;
  assign n30332 = ~pi778 & n30310;
  assign n30333 = ~n30314 & ~n30324;
  assign n30334 = pi778 & ~n30333;
  assign n30335 = ~n30332 & ~n30334;
  assign n30336 = pi609 & n30335;
  assign n30337 = ~pi1155 & ~n30336;
  assign n30338 = ~n30331 & n30337;
  assign n30339 = n17526 & ~n30300;
  assign n30340 = ~n17526 & n30296;
  assign n30341 = ~n30339 & ~n30340;
  assign n30342 = pi609 & ~n30341;
  assign n30343 = ~pi609 & ~n30300;
  assign n30344 = pi1155 & ~n30343;
  assign n30345 = ~n30342 & n30344;
  assign n30346 = ~pi660 & ~n30345;
  assign n30347 = ~n30338 & n30346;
  assign n30348 = pi609 & ~n30330;
  assign n30349 = ~pi609 & n30335;
  assign n30350 = pi1155 & ~n30349;
  assign n30351 = ~n30348 & n30350;
  assign n30352 = ~pi609 & ~n30341;
  assign n30353 = pi609 & ~n30300;
  assign n30354 = ~pi1155 & ~n30353;
  assign n30355 = ~n30352 & n30354;
  assign n30356 = pi660 & ~n30355;
  assign n30357 = ~n30351 & n30356;
  assign n30358 = ~n30347 & ~n30357;
  assign n30359 = pi785 & ~n30358;
  assign n30360 = ~pi785 & ~n30330;
  assign n30361 = ~n30359 & ~n30360;
  assign n30362 = ~pi618 & ~n30361;
  assign n30363 = n17554 & ~n30300;
  assign n30364 = ~n17554 & n30335;
  assign n30365 = ~n30363 & ~n30364;
  assign n30366 = pi618 & ~n30365;
  assign n30367 = ~pi1154 & ~n30366;
  assign n30368 = ~n30362 & n30367;
  assign n30369 = ~pi785 & n30341;
  assign n30370 = ~n30345 & ~n30355;
  assign n30371 = pi785 & ~n30370;
  assign n30372 = ~n30369 & ~n30371;
  assign n30373 = pi618 & n30372;
  assign n30374 = ~pi618 & ~n30300;
  assign n30375 = pi1154 & ~n30374;
  assign n30376 = ~n30373 & n30375;
  assign n30377 = ~pi627 & ~n30376;
  assign n30378 = ~n30368 & n30377;
  assign n30379 = pi618 & ~n30361;
  assign n30380 = ~pi618 & ~n30365;
  assign n30381 = pi1154 & ~n30380;
  assign n30382 = ~n30379 & n30381;
  assign n30383 = ~pi618 & n30372;
  assign n30384 = pi618 & ~n30300;
  assign n30385 = ~pi1154 & ~n30384;
  assign n30386 = ~n30383 & n30385;
  assign n30387 = pi627 & ~n30386;
  assign n30388 = ~n30382 & n30387;
  assign n30389 = ~n30378 & ~n30388;
  assign n30390 = pi781 & ~n30389;
  assign n30391 = ~pi781 & ~n30361;
  assign n30392 = ~n30390 & ~n30391;
  assign n30393 = ~pi619 & ~n30392;
  assign n30394 = ~n17591 & n30365;
  assign n30395 = n17591 & n30300;
  assign n30396 = ~n30394 & ~n30395;
  assign n30397 = pi619 & n30396;
  assign n30398 = ~pi1159 & ~n30397;
  assign n30399 = ~n30393 & n30398;
  assign n30400 = ~pi781 & ~n30372;
  assign n30401 = ~n30376 & ~n30386;
  assign n30402 = pi781 & ~n30401;
  assign n30403 = ~n30400 & ~n30402;
  assign n30404 = pi619 & n30403;
  assign n30405 = ~pi619 & ~n30300;
  assign n30406 = pi1159 & ~n30405;
  assign n30407 = ~n30404 & n30406;
  assign n30408 = ~pi648 & ~n30407;
  assign n30409 = ~n30399 & n30408;
  assign n30410 = pi619 & ~n30392;
  assign n30411 = ~pi619 & n30396;
  assign n30412 = pi1159 & ~n30411;
  assign n30413 = ~n30410 & n30412;
  assign n30414 = ~pi619 & n30403;
  assign n30415 = pi619 & ~n30300;
  assign n30416 = ~pi1159 & ~n30415;
  assign n30417 = ~n30414 & n30416;
  assign n30418 = pi648 & ~n30417;
  assign n30419 = ~n30413 & n30418;
  assign n30420 = ~n30409 & ~n30419;
  assign n30421 = pi789 & ~n30420;
  assign n30422 = ~pi789 & ~n30392;
  assign n30423 = ~n30421 & ~n30422;
  assign n30424 = ~pi788 & n30423;
  assign n30425 = ~pi626 & n30423;
  assign n30426 = n17627 & ~n30300;
  assign n30427 = ~n17627 & n30396;
  assign n30428 = ~n30426 & ~n30427;
  assign n30429 = pi626 & n30428;
  assign n30430 = ~pi641 & ~n30429;
  assign n30431 = ~n30425 & n30430;
  assign n30432 = ~pi789 & ~n30403;
  assign n30433 = ~n30407 & ~n30417;
  assign n30434 = pi789 & ~n30433;
  assign n30435 = ~n30432 & ~n30434;
  assign n30436 = ~pi626 & ~n30435;
  assign n30437 = pi626 & n30300;
  assign n30438 = pi641 & ~n30437;
  assign n30439 = ~n30436 & n30438;
  assign n30440 = ~pi1158 & ~n30439;
  assign n30441 = ~n30431 & n30440;
  assign n30442 = pi626 & n30423;
  assign n30443 = ~pi626 & n30428;
  assign n30444 = pi641 & ~n30443;
  assign n30445 = ~n30442 & n30444;
  assign n30446 = pi626 & ~n30435;
  assign n30447 = ~pi626 & n30300;
  assign n30448 = ~pi641 & ~n30447;
  assign n30449 = ~n30446 & n30448;
  assign n30450 = pi1158 & ~n30449;
  assign n30451 = ~n30445 & n30450;
  assign n30452 = ~n30441 & ~n30451;
  assign n30453 = pi788 & ~n30452;
  assign n30454 = ~n30424 & ~n30453;
  assign n30455 = ~pi628 & n30454;
  assign n30456 = ~n17904 & ~n30435;
  assign n30457 = n17904 & n30300;
  assign n30458 = ~n30456 & ~n30457;
  assign n30459 = pi628 & n30458;
  assign n30460 = ~pi1156 & ~n30459;
  assign n30461 = ~n30455 & n30460;
  assign n30462 = ~n17670 & n30428;
  assign n30463 = n17670 & n30300;
  assign n30464 = ~n30462 & ~n30463;
  assign n30465 = pi628 & n30464;
  assign n30466 = ~pi628 & ~n30300;
  assign n30467 = pi1156 & ~n30466;
  assign n30468 = ~n30465 & n30467;
  assign n30469 = ~pi629 & ~n30468;
  assign n30470 = ~n30461 & n30469;
  assign n30471 = pi628 & n30454;
  assign n30472 = ~pi628 & n30458;
  assign n30473 = pi1156 & ~n30472;
  assign n30474 = ~n30471 & n30473;
  assign n30475 = ~pi628 & n30464;
  assign n30476 = pi628 & ~n30300;
  assign n30477 = ~pi1156 & ~n30476;
  assign n30478 = ~n30475 & n30477;
  assign n30479 = pi629 & ~n30478;
  assign n30480 = ~n30474 & n30479;
  assign n30481 = ~n30470 & ~n30480;
  assign n30482 = pi792 & ~n30481;
  assign n30483 = ~pi792 & n30454;
  assign n30484 = ~n30482 & ~n30483;
  assign n30485 = ~pi647 & ~n30484;
  assign n30486 = ~n17698 & ~n30458;
  assign n30487 = n17698 & n30300;
  assign n30488 = ~n30486 & ~n30487;
  assign n30489 = pi647 & n30488;
  assign n30490 = ~pi1157 & ~n30489;
  assign n30491 = ~n30485 & n30490;
  assign n30492 = ~pi792 & ~n30464;
  assign n30493 = ~n30468 & ~n30478;
  assign n30494 = pi792 & ~n30493;
  assign n30495 = ~n30492 & ~n30494;
  assign n30496 = pi647 & n30495;
  assign n30497 = ~pi647 & ~n30300;
  assign n30498 = pi1157 & ~n30497;
  assign n30499 = ~n30496 & n30498;
  assign n30500 = ~pi630 & ~n30499;
  assign n30501 = ~n30491 & n30500;
  assign n30502 = pi647 & ~n30484;
  assign n30503 = ~pi647 & n30488;
  assign n30504 = pi1157 & ~n30503;
  assign n30505 = ~n30502 & n30504;
  assign n30506 = ~pi647 & n30495;
  assign n30507 = pi647 & ~n30300;
  assign n30508 = ~pi1157 & ~n30507;
  assign n30509 = ~n30506 & n30508;
  assign n30510 = pi630 & ~n30509;
  assign n30511 = ~n30505 & n30510;
  assign n30512 = ~n30501 & ~n30511;
  assign n30513 = pi787 & ~n30512;
  assign n30514 = ~pi787 & ~n30484;
  assign n30515 = ~n30513 & ~n30514;
  assign n30516 = pi644 & ~n30515;
  assign n30517 = ~pi787 & ~n30495;
  assign n30518 = ~n30499 & ~n30509;
  assign n30519 = pi787 & ~n30518;
  assign n30520 = ~n30517 & ~n30519;
  assign n30521 = ~pi644 & n30520;
  assign n30522 = pi715 & ~n30521;
  assign n30523 = ~n30516 & n30522;
  assign n30524 = n17740 & ~n30300;
  assign n30525 = ~n17740 & n30488;
  assign n30526 = ~n30524 & ~n30525;
  assign n30527 = pi644 & ~n30526;
  assign n30528 = ~pi644 & ~n30300;
  assign n30529 = ~pi715 & ~n30528;
  assign n30530 = ~n30527 & n30529;
  assign n30531 = pi1160 & ~n30530;
  assign n30532 = ~n30523 & n30531;
  assign n30533 = ~pi644 & ~n30515;
  assign n30534 = pi644 & n30520;
  assign n30535 = ~pi715 & ~n30534;
  assign n30536 = ~n30533 & n30535;
  assign n30537 = ~pi644 & ~n30526;
  assign n30538 = pi644 & ~n30300;
  assign n30539 = pi715 & ~n30538;
  assign n30540 = ~n30537 & n30539;
  assign n30541 = ~pi1160 & ~n30540;
  assign n30542 = ~n30536 & n30541;
  assign n30543 = pi790 & ~n30532;
  assign n30544 = ~n30542 & n30543;
  assign n30545 = ~pi790 & n30515;
  assign n30546 = n6294 & ~n30545;
  assign n30547 = ~n30544 & n30546;
  assign n30548 = ~pi189 & ~n6294;
  assign n30549 = ~pi57 & ~n30548;
  assign n30550 = ~n30547 & n30549;
  assign n30551 = pi57 & pi189;
  assign n30552 = ~pi832 & ~n30551;
  assign n30553 = ~n30550 & n30552;
  assign n30554 = pi189 & ~n2755;
  assign n30555 = pi772 & n16933;
  assign n30556 = ~n30554 & ~n30555;
  assign n30557 = pi727 & n17154;
  assign n30558 = n30556 & ~n30557;
  assign n30559 = pi625 & n30557;
  assign n30560 = ~n30558 & ~n30559;
  assign n30561 = ~pi1153 & ~n30560;
  assign n30562 = pi727 & n17153;
  assign n30563 = pi625 & n30562;
  assign n30564 = pi1153 & ~n30554;
  assign n30565 = ~n30563 & n30564;
  assign n30566 = ~pi608 & ~n30565;
  assign n30567 = ~n30561 & n30566;
  assign n30568 = ~n30554 & ~n30562;
  assign n30569 = ~n30563 & ~n30568;
  assign n30570 = ~pi1153 & ~n30569;
  assign n30571 = pi1153 & n30556;
  assign n30572 = ~n30559 & n30571;
  assign n30573 = pi608 & ~n30570;
  assign n30574 = ~n30572 & n30573;
  assign n30575 = ~n30567 & ~n30574;
  assign n30576 = pi778 & ~n30575;
  assign n30577 = ~pi778 & ~n30558;
  assign n30578 = ~n30576 & ~n30577;
  assign n30579 = ~pi609 & ~n30578;
  assign n30580 = ~pi778 & n30568;
  assign n30581 = ~n30565 & ~n30570;
  assign n30582 = pi778 & ~n30581;
  assign n30583 = ~n30580 & ~n30582;
  assign n30584 = pi609 & n30583;
  assign n30585 = ~pi1155 & ~n30584;
  assign n30586 = ~n30579 & n30585;
  assign n30587 = n17527 & n30555;
  assign n30588 = pi1155 & ~n30554;
  assign n30589 = ~n30587 & n30588;
  assign n30590 = ~pi660 & ~n30589;
  assign n30591 = ~n30586 & n30590;
  assign n30592 = pi609 & ~n30578;
  assign n30593 = ~pi609 & n30583;
  assign n30594 = pi1155 & ~n30593;
  assign n30595 = ~n30592 & n30594;
  assign n30596 = n17539 & n30555;
  assign n30597 = ~pi1155 & ~n30554;
  assign n30598 = ~n30596 & n30597;
  assign n30599 = pi660 & ~n30598;
  assign n30600 = ~n30595 & n30599;
  assign n30601 = ~n30591 & ~n30600;
  assign n30602 = pi785 & ~n30601;
  assign n30603 = ~pi785 & ~n30578;
  assign n30604 = ~n30602 & ~n30603;
  assign n30605 = pi618 & ~n30604;
  assign n30606 = ~n17554 & n30583;
  assign n30607 = ~n30554 & ~n30606;
  assign n30608 = ~pi618 & ~n30607;
  assign n30609 = pi1154 & ~n30608;
  assign n30610 = ~n30605 & n30609;
  assign n30611 = ~n20159 & n30555;
  assign n30612 = n20257 & n30611;
  assign n30613 = ~pi1154 & ~n30554;
  assign n30614 = ~n30612 & n30613;
  assign n30615 = pi627 & ~n30614;
  assign n30616 = ~n30610 & n30615;
  assign n30617 = ~pi618 & ~n30604;
  assign n30618 = pi618 & ~n30607;
  assign n30619 = ~pi1154 & ~n30618;
  assign n30620 = ~n30617 & n30619;
  assign n30621 = n20247 & n30611;
  assign n30622 = pi1154 & ~n30554;
  assign n30623 = ~n30621 & n30622;
  assign n30624 = ~pi627 & ~n30623;
  assign n30625 = ~n30620 & n30624;
  assign n30626 = ~n30616 & ~n30625;
  assign n30627 = pi781 & ~n30626;
  assign n30628 = ~pi781 & ~n30604;
  assign n30629 = ~n23544 & ~n30628;
  assign n30630 = ~n30627 & n30629;
  assign n30631 = n19216 & n30583;
  assign n30632 = ~n23542 & ~n30631;
  assign n30633 = ~n20169 & n30611;
  assign n30634 = n20282 & n30633;
  assign n30635 = n17625 & ~n30634;
  assign n30636 = n20272 & n30633;
  assign n30637 = n17624 & ~n30636;
  assign n30638 = ~n30635 & ~n30637;
  assign n30639 = ~n30632 & n30638;
  assign n30640 = pi789 & ~n30554;
  assign n30641 = ~n30639 & n30640;
  assign n30642 = n17905 & ~n30641;
  assign n30643 = ~n30630 & n30642;
  assign n30644 = ~n17627 & n30631;
  assign n30645 = ~n30554 & ~n30644;
  assign n30646 = n17786 & ~n30645;
  assign n30647 = n20171 & n30611;
  assign n30648 = ~pi626 & n30647;
  assign n30649 = ~n30554 & ~n30648;
  assign n30650 = ~pi1158 & ~n30649;
  assign n30651 = pi641 & ~n30650;
  assign n30652 = ~n30646 & n30651;
  assign n30653 = n17787 & ~n30645;
  assign n30654 = pi626 & n30647;
  assign n30655 = ~n30554 & ~n30654;
  assign n30656 = pi1158 & ~n30655;
  assign n30657 = ~pi641 & ~n30656;
  assign n30658 = ~n30653 & n30657;
  assign n30659 = pi788 & ~n30652;
  assign n30660 = ~n30658 & n30659;
  assign n30661 = ~n20298 & ~n30660;
  assign n30662 = ~n30643 & n30661;
  assign n30663 = ~n17904 & n30647;
  assign n30664 = ~pi629 & n30663;
  assign n30665 = pi628 & ~n30664;
  assign n30666 = n19217 & n30583;
  assign n30667 = pi629 & ~n30666;
  assign n30668 = ~n30665 & ~n30667;
  assign n30669 = ~pi1156 & ~n30668;
  assign n30670 = pi628 & n30666;
  assign n30671 = ~pi628 & ~n30663;
  assign n30672 = pi629 & ~n30671;
  assign n30673 = pi1156 & ~n30672;
  assign n30674 = ~n30670 & n30673;
  assign n30675 = ~n30669 & ~n30674;
  assign n30676 = pi792 & ~n30554;
  assign n30677 = ~n30675 & n30676;
  assign n30678 = ~n30662 & ~n30677;
  assign n30679 = n20300 & ~n30678;
  assign n30680 = ~n17698 & n30663;
  assign n30681 = ~pi630 & n30680;
  assign n30682 = pi647 & ~n30681;
  assign n30683 = ~n19247 & n30666;
  assign n30684 = pi630 & ~n30683;
  assign n30685 = ~n30682 & ~n30684;
  assign n30686 = ~pi1157 & ~n30685;
  assign n30687 = ~pi630 & ~n30683;
  assign n30688 = pi647 & ~n30687;
  assign n30689 = pi630 & n30680;
  assign n30690 = pi1157 & ~n30689;
  assign n30691 = ~n30688 & n30690;
  assign n30692 = ~n30686 & ~n30691;
  assign n30693 = pi787 & ~n30554;
  assign n30694 = ~n30692 & n30693;
  assign n30695 = ~n30679 & ~n30694;
  assign n30696 = pi644 & n30695;
  assign n30697 = ~n19271 & n30683;
  assign n30698 = ~n30554 & ~n30697;
  assign n30699 = ~pi644 & ~n30698;
  assign n30700 = pi715 & ~n30699;
  assign n30701 = ~n30696 & n30700;
  assign n30702 = ~n17904 & n23618;
  assign n30703 = n30647 & n30702;
  assign n30704 = pi644 & n30703;
  assign n30705 = ~pi715 & ~n30554;
  assign n30706 = ~n30704 & n30705;
  assign n30707 = pi1160 & ~n30706;
  assign n30708 = ~n30701 & n30707;
  assign n30709 = ~pi644 & n30695;
  assign n30710 = pi644 & ~n30698;
  assign n30711 = ~pi715 & ~n30710;
  assign n30712 = ~n30709 & n30711;
  assign n30713 = ~pi644 & n30703;
  assign n30714 = pi715 & ~n30554;
  assign n30715 = ~n30713 & n30714;
  assign n30716 = ~pi1160 & ~n30715;
  assign n30717 = ~n30712 & n30716;
  assign n30718 = ~n30708 & ~n30717;
  assign n30719 = pi790 & ~n30718;
  assign n30720 = ~pi790 & n30695;
  assign n30721 = pi832 & ~n30720;
  assign n30722 = ~n30719 & n30721;
  assign po346 = ~n30553 & ~n30722;
  assign n30724 = ~pi190 & ~n2755;
  assign n30725 = pi763 & n16933;
  assign n30726 = ~n30724 & ~n30725;
  assign n30727 = ~n17794 & ~n30726;
  assign n30728 = ~pi785 & ~n30727;
  assign n30729 = n17539 & n30725;
  assign n30730 = n30727 & ~n30729;
  assign n30731 = pi1155 & ~n30730;
  assign n30732 = ~pi1155 & ~n30724;
  assign n30733 = ~n30729 & n30732;
  assign n30734 = ~n30731 & ~n30733;
  assign n30735 = pi785 & ~n30734;
  assign n30736 = ~n30728 & ~n30735;
  assign n30737 = ~pi781 & ~n30736;
  assign n30738 = ~n17809 & n30736;
  assign n30739 = pi1154 & ~n30738;
  assign n30740 = ~n17812 & n30736;
  assign n30741 = ~pi1154 & ~n30740;
  assign n30742 = ~n30739 & ~n30741;
  assign n30743 = pi781 & ~n30742;
  assign n30744 = ~n30737 & ~n30743;
  assign n30745 = ~pi789 & ~n30744;
  assign n30746 = ~n22988 & n30744;
  assign n30747 = pi1159 & ~n30746;
  assign n30748 = ~n22991 & n30744;
  assign n30749 = ~pi1159 & ~n30748;
  assign n30750 = ~n30747 & ~n30749;
  assign n30751 = pi789 & ~n30750;
  assign n30752 = ~n30745 & ~n30751;
  assign n30753 = ~n17904 & n30752;
  assign n30754 = n17904 & n30724;
  assign n30755 = ~n30753 & ~n30754;
  assign n30756 = ~n17698 & ~n30755;
  assign n30757 = n17698 & n30724;
  assign n30758 = ~n30756 & ~n30757;
  assign n30759 = ~n20491 & n30758;
  assign n30760 = pi699 & n17153;
  assign n30761 = ~n30724 & ~n30760;
  assign n30762 = ~pi778 & ~n30761;
  assign n30763 = ~pi625 & n30760;
  assign n30764 = ~n30761 & ~n30763;
  assign n30765 = pi1153 & ~n30764;
  assign n30766 = ~pi1153 & ~n30724;
  assign n30767 = ~n30763 & n30766;
  assign n30768 = pi778 & ~n30767;
  assign n30769 = ~n30765 & n30768;
  assign n30770 = ~n30762 & ~n30769;
  assign n30771 = ~n17780 & ~n30770;
  assign n30772 = ~n17782 & n30771;
  assign n30773 = ~n17784 & n30772;
  assign n30774 = ~n17916 & n30773;
  assign n30775 = ~n17947 & n30774;
  assign n30776 = ~pi647 & n30775;
  assign n30777 = pi647 & n30724;
  assign n30778 = ~pi1157 & ~n30777;
  assign n30779 = ~n30776 & n30778;
  assign n30780 = pi647 & ~n30775;
  assign n30781 = ~pi647 & ~n30724;
  assign n30782 = ~n30780 & ~n30781;
  assign n30783 = pi1157 & ~n30782;
  assign n30784 = ~n30779 & ~n30783;
  assign n30785 = ~n17739 & ~n30784;
  assign n30786 = ~n30759 & ~n30785;
  assign n30787 = pi787 & ~n30786;
  assign n30788 = ~pi626 & ~n30752;
  assign n30789 = pi626 & ~n30724;
  assign n30790 = n17668 & ~n30789;
  assign n30791 = ~n30788 & n30790;
  assign n30792 = pi626 & ~n30752;
  assign n30793 = ~pi626 & ~n30724;
  assign n30794 = n17667 & ~n30793;
  assign n30795 = ~n30792 & n30794;
  assign n30796 = n17792 & n30773;
  assign n30797 = ~n30791 & ~n30796;
  assign n30798 = ~n30795 & n30797;
  assign n30799 = pi788 & ~n30798;
  assign n30800 = ~n16842 & ~n30761;
  assign n30801 = pi625 & n30800;
  assign n30802 = n30726 & ~n30800;
  assign n30803 = ~n30801 & ~n30802;
  assign n30804 = n30766 & ~n30803;
  assign n30805 = ~pi608 & ~n30765;
  assign n30806 = ~n30804 & n30805;
  assign n30807 = pi1153 & n30726;
  assign n30808 = ~n30801 & n30807;
  assign n30809 = pi608 & ~n30767;
  assign n30810 = ~n30808 & n30809;
  assign n30811 = ~n30806 & ~n30810;
  assign n30812 = pi778 & ~n30811;
  assign n30813 = ~pi778 & ~n30802;
  assign n30814 = ~n30812 & ~n30813;
  assign n30815 = ~pi609 & ~n30814;
  assign n30816 = pi609 & ~n30770;
  assign n30817 = ~pi1155 & ~n30816;
  assign n30818 = ~n30815 & n30817;
  assign n30819 = ~pi660 & ~n30731;
  assign n30820 = ~n30818 & n30819;
  assign n30821 = pi609 & ~n30814;
  assign n30822 = ~pi609 & ~n30770;
  assign n30823 = pi1155 & ~n30822;
  assign n30824 = ~n30821 & n30823;
  assign n30825 = pi660 & ~n30733;
  assign n30826 = ~n30824 & n30825;
  assign n30827 = ~n30820 & ~n30826;
  assign n30828 = pi785 & ~n30827;
  assign n30829 = ~pi785 & ~n30814;
  assign n30830 = ~n30828 & ~n30829;
  assign n30831 = ~pi618 & ~n30830;
  assign n30832 = pi618 & n30771;
  assign n30833 = ~pi1154 & ~n30832;
  assign n30834 = ~n30831 & n30833;
  assign n30835 = ~pi627 & ~n30739;
  assign n30836 = ~n30834 & n30835;
  assign n30837 = pi618 & ~n30830;
  assign n30838 = ~pi618 & n30771;
  assign n30839 = pi1154 & ~n30838;
  assign n30840 = ~n30837 & n30839;
  assign n30841 = pi627 & ~n30741;
  assign n30842 = ~n30840 & n30841;
  assign n30843 = ~n30836 & ~n30842;
  assign n30844 = pi781 & ~n30843;
  assign n30845 = ~pi781 & ~n30830;
  assign n30846 = ~n30844 & ~n30845;
  assign n30847 = ~pi619 & ~n30846;
  assign n30848 = pi619 & n30772;
  assign n30849 = ~pi1159 & ~n30848;
  assign n30850 = ~n30847 & n30849;
  assign n30851 = ~pi648 & ~n30747;
  assign n30852 = ~n30850 & n30851;
  assign n30853 = pi619 & ~n30846;
  assign n30854 = ~pi619 & n30772;
  assign n30855 = pi1159 & ~n30854;
  assign n30856 = ~n30853 & n30855;
  assign n30857 = pi648 & ~n30749;
  assign n30858 = ~n30856 & n30857;
  assign n30859 = pi789 & ~n30852;
  assign n30860 = ~n30858 & n30859;
  assign n30861 = ~pi789 & n30846;
  assign n30862 = n17905 & ~n30861;
  assign n30863 = ~n30860 & n30862;
  assign n30864 = ~n30799 & ~n30863;
  assign n30865 = ~n20298 & ~n30864;
  assign n30866 = n17944 & ~n30755;
  assign n30867 = n20786 & n30774;
  assign n30868 = ~n30866 & ~n30867;
  assign n30869 = ~pi629 & ~n30868;
  assign n30870 = n20790 & n30774;
  assign n30871 = n17943 & ~n30755;
  assign n30872 = ~n30870 & ~n30871;
  assign n30873 = pi629 & ~n30872;
  assign n30874 = ~n30869 & ~n30873;
  assign n30875 = pi792 & ~n30874;
  assign n30876 = n20300 & ~n30875;
  assign n30877 = ~n30865 & n30876;
  assign n30878 = ~n30787 & ~n30877;
  assign n30879 = pi644 & n30878;
  assign n30880 = ~pi787 & ~n30775;
  assign n30881 = pi787 & ~n30784;
  assign n30882 = ~n30880 & ~n30881;
  assign n30883 = ~pi644 & n30882;
  assign n30884 = pi715 & ~n30883;
  assign n30885 = ~n30879 & n30884;
  assign n30886 = ~n17740 & ~n30758;
  assign n30887 = n17740 & n30724;
  assign n30888 = ~n30886 & ~n30887;
  assign n30889 = pi644 & ~n30888;
  assign n30890 = ~pi644 & n30724;
  assign n30891 = ~pi715 & ~n30890;
  assign n30892 = ~n30889 & n30891;
  assign n30893 = pi1160 & ~n30892;
  assign n30894 = ~n30885 & n30893;
  assign n30895 = ~pi644 & n30878;
  assign n30896 = pi644 & n30882;
  assign n30897 = ~pi715 & ~n30896;
  assign n30898 = ~n30895 & n30897;
  assign n30899 = ~pi644 & ~n30888;
  assign n30900 = pi644 & n30724;
  assign n30901 = pi715 & ~n30900;
  assign n30902 = ~n30899 & n30901;
  assign n30903 = ~pi1160 & ~n30902;
  assign n30904 = ~n30898 & n30903;
  assign n30905 = ~n30894 & ~n30904;
  assign n30906 = pi790 & ~n30905;
  assign n30907 = ~pi790 & n30878;
  assign n30908 = pi832 & ~n30907;
  assign n30909 = ~n30906 & n30908;
  assign n30910 = ~pi190 & ~n17494;
  assign n30911 = n17627 & ~n30910;
  assign n30912 = pi190 & ~n3268;
  assign n30913 = ~pi190 & n18060;
  assign n30914 = pi190 & ~n18064;
  assign n30915 = ~pi38 & ~n30914;
  assign n30916 = ~n30913 & n30915;
  assign n30917 = ~pi190 & ~n16968;
  assign n30918 = n17480 & ~n30917;
  assign n30919 = pi699 & ~n30918;
  assign n30920 = ~n30916 & n30919;
  assign n30921 = ~pi190 & ~pi699;
  assign n30922 = ~n17487 & n30921;
  assign n30923 = n3268 & ~n30922;
  assign n30924 = ~n30920 & n30923;
  assign n30925 = ~n30912 & ~n30924;
  assign n30926 = ~pi778 & ~n30925;
  assign n30927 = pi625 & n30925;
  assign n30928 = ~pi625 & n30910;
  assign n30929 = pi1153 & ~n30928;
  assign n30930 = ~n30927 & n30929;
  assign n30931 = ~pi625 & n30925;
  assign n30932 = pi625 & n30910;
  assign n30933 = ~pi1153 & ~n30932;
  assign n30934 = ~n30931 & n30933;
  assign n30935 = ~n30930 & ~n30934;
  assign n30936 = pi778 & ~n30935;
  assign n30937 = ~n30926 & ~n30936;
  assign n30938 = ~n17554 & ~n30937;
  assign n30939 = n17554 & ~n30910;
  assign n30940 = ~n30938 & ~n30939;
  assign n30941 = ~n17591 & n30940;
  assign n30942 = n17591 & n30910;
  assign n30943 = ~n30941 & ~n30942;
  assign n30944 = ~n17627 & n30943;
  assign n30945 = ~n30911 & ~n30944;
  assign n30946 = ~n17670 & n30945;
  assign n30947 = n17670 & n30910;
  assign n30948 = ~n30946 & ~n30947;
  assign n30949 = ~pi628 & ~n30948;
  assign n30950 = pi628 & n30910;
  assign n30951 = ~n30949 & ~n30950;
  assign n30952 = ~pi1156 & ~n30951;
  assign n30953 = pi628 & ~n30948;
  assign n30954 = ~pi628 & n30910;
  assign n30955 = ~n30953 & ~n30954;
  assign n30956 = pi1156 & ~n30955;
  assign n30957 = ~n30952 & ~n30956;
  assign n30958 = pi792 & ~n30957;
  assign n30959 = ~pi792 & ~n30948;
  assign n30960 = ~n30958 & ~n30959;
  assign n30961 = ~pi647 & ~n30960;
  assign n30962 = pi647 & n30910;
  assign n30963 = ~n30961 & ~n30962;
  assign n30964 = ~pi1157 & ~n30963;
  assign n30965 = pi647 & ~n30960;
  assign n30966 = ~pi647 & n30910;
  assign n30967 = ~n30965 & ~n30966;
  assign n30968 = pi1157 & ~n30967;
  assign n30969 = ~n30964 & ~n30968;
  assign n30970 = pi787 & ~n30969;
  assign n30971 = ~pi787 & ~n30960;
  assign n30972 = ~n30970 & ~n30971;
  assign n30973 = ~pi644 & ~n30972;
  assign n30974 = pi715 & ~n30973;
  assign n30975 = ~pi763 & n16814;
  assign n30976 = pi190 & n16961;
  assign n30977 = ~n30975 & ~n30976;
  assign n30978 = pi39 & ~n30977;
  assign n30979 = ~pi190 & pi763;
  assign n30980 = n16907 & n30979;
  assign n30981 = pi763 & ~n16919;
  assign n30982 = pi190 & ~n30981;
  assign n30983 = ~n22287 & ~n30982;
  assign n30984 = ~n30980 & n30983;
  assign n30985 = ~n30978 & n30984;
  assign n30986 = ~pi38 & ~n30985;
  assign n30987 = pi763 & n16970;
  assign n30988 = pi38 & ~n30917;
  assign n30989 = ~n30987 & n30988;
  assign n30990 = ~n30986 & ~n30989;
  assign n30991 = n3268 & ~n30990;
  assign n30992 = ~n30912 & ~n30991;
  assign n30993 = ~n17526 & ~n30992;
  assign n30994 = n17526 & ~n30910;
  assign n30995 = ~n30993 & ~n30994;
  assign n30996 = ~pi785 & ~n30995;
  assign n30997 = ~n17527 & ~n30910;
  assign n30998 = pi609 & n30993;
  assign n30999 = ~n30997 & ~n30998;
  assign n31000 = pi1155 & ~n30999;
  assign n31001 = ~n17539 & ~n30910;
  assign n31002 = ~pi609 & n30993;
  assign n31003 = ~n31001 & ~n31002;
  assign n31004 = ~pi1155 & ~n31003;
  assign n31005 = ~n31000 & ~n31004;
  assign n31006 = pi785 & ~n31005;
  assign n31007 = ~n30996 & ~n31006;
  assign n31008 = ~pi781 & ~n31007;
  assign n31009 = pi618 & n31007;
  assign n31010 = ~pi618 & n30910;
  assign n31011 = pi1154 & ~n31010;
  assign n31012 = ~n31009 & n31011;
  assign n31013 = ~pi618 & n31007;
  assign n31014 = pi618 & n30910;
  assign n31015 = ~pi1154 & ~n31014;
  assign n31016 = ~n31013 & n31015;
  assign n31017 = ~n31012 & ~n31016;
  assign n31018 = pi781 & ~n31017;
  assign n31019 = ~n31008 & ~n31018;
  assign n31020 = ~pi789 & ~n31019;
  assign n31021 = pi619 & n31019;
  assign n31022 = ~pi619 & n30910;
  assign n31023 = pi1159 & ~n31022;
  assign n31024 = ~n31021 & n31023;
  assign n31025 = ~pi619 & n31019;
  assign n31026 = pi619 & n30910;
  assign n31027 = ~pi1159 & ~n31026;
  assign n31028 = ~n31025 & n31027;
  assign n31029 = ~n31024 & ~n31028;
  assign n31030 = pi789 & ~n31029;
  assign n31031 = ~n31020 & ~n31030;
  assign n31032 = ~n17904 & n31031;
  assign n31033 = n17904 & n30910;
  assign n31034 = ~n31032 & ~n31033;
  assign n31035 = ~n17698 & ~n31034;
  assign n31036 = n17698 & n30910;
  assign n31037 = ~n31035 & ~n31036;
  assign n31038 = ~n17740 & ~n31037;
  assign n31039 = n17740 & n30910;
  assign n31040 = ~n31038 & ~n31039;
  assign n31041 = pi644 & ~n31040;
  assign n31042 = ~pi644 & n30910;
  assign n31043 = ~pi715 & ~n31042;
  assign n31044 = ~n31041 & n31043;
  assign n31045 = pi1160 & ~n31044;
  assign n31046 = ~n30974 & n31045;
  assign n31047 = pi644 & ~n30972;
  assign n31048 = ~pi715 & ~n31047;
  assign n31049 = ~pi644 & ~n31040;
  assign n31050 = pi644 & n30910;
  assign n31051 = pi715 & ~n31050;
  assign n31052 = ~n31049 & n31051;
  assign n31053 = ~pi1160 & ~n31052;
  assign n31054 = ~n31048 & n31053;
  assign n31055 = ~n31046 & ~n31054;
  assign n31056 = pi790 & ~n31055;
  assign n31057 = ~pi644 & n31053;
  assign n31058 = pi644 & n31045;
  assign n31059 = pi790 & ~n31057;
  assign n31060 = ~n31058 & n31059;
  assign n31061 = ~n20502 & n31034;
  assign n31062 = n17696 & n30951;
  assign n31063 = n17695 & n30955;
  assign n31064 = ~n31062 & ~n31063;
  assign n31065 = ~n31061 & n31064;
  assign n31066 = pi792 & ~n31065;
  assign n31067 = ~pi699 & n30990;
  assign n31068 = ~pi190 & n17074;
  assign n31069 = pi190 & n17166;
  assign n31070 = ~pi763 & ~n31069;
  assign n31071 = ~n31068 & n31070;
  assign n31072 = pi190 & n17233;
  assign n31073 = ~pi190 & ~n17295;
  assign n31074 = pi763 & ~n31073;
  assign n31075 = ~n31072 & n31074;
  assign n31076 = pi39 & ~n31075;
  assign n31077 = ~n31071 & n31076;
  assign n31078 = ~pi190 & n17317;
  assign n31079 = pi190 & n17340;
  assign n31080 = ~pi763 & ~n31078;
  assign n31081 = ~n31079 & n31080;
  assign n31082 = ~pi190 & ~n17344;
  assign n31083 = pi190 & ~n17351;
  assign n31084 = pi763 & ~n31083;
  assign n31085 = ~n31082 & n31084;
  assign n31086 = ~pi39 & ~n31085;
  assign n31087 = ~n31081 & n31086;
  assign n31088 = ~pi38 & ~n31087;
  assign n31089 = ~n31077 & n31088;
  assign n31090 = ~pi763 & n24006;
  assign n31091 = ~n17259 & ~n31090;
  assign n31092 = ~pi39 & ~n31091;
  assign n31093 = ~pi190 & ~n31092;
  assign n31094 = ~n17154 & ~n30725;
  assign n31095 = pi190 & ~n31094;
  assign n31096 = n6250 & n31095;
  assign n31097 = pi38 & ~n31096;
  assign n31098 = ~n31093 & n31097;
  assign n31099 = pi699 & ~n31098;
  assign n31100 = ~n31089 & n31099;
  assign n31101 = n3268 & ~n31100;
  assign n31102 = ~n31067 & n31101;
  assign n31103 = ~n30912 & ~n31102;
  assign n31104 = ~pi625 & n31103;
  assign n31105 = pi625 & n30992;
  assign n31106 = ~pi1153 & ~n31105;
  assign n31107 = ~n31104 & n31106;
  assign n31108 = ~pi608 & ~n30930;
  assign n31109 = ~n31107 & n31108;
  assign n31110 = pi625 & n31103;
  assign n31111 = ~pi625 & n30992;
  assign n31112 = pi1153 & ~n31111;
  assign n31113 = ~n31110 & n31112;
  assign n31114 = pi608 & ~n30934;
  assign n31115 = ~n31113 & n31114;
  assign n31116 = ~n31109 & ~n31115;
  assign n31117 = pi778 & ~n31116;
  assign n31118 = ~pi778 & n31103;
  assign n31119 = ~n31117 & ~n31118;
  assign n31120 = ~pi609 & ~n31119;
  assign n31121 = pi609 & n30937;
  assign n31122 = ~pi1155 & ~n31121;
  assign n31123 = ~n31120 & n31122;
  assign n31124 = ~pi660 & ~n31000;
  assign n31125 = ~n31123 & n31124;
  assign n31126 = pi609 & ~n31119;
  assign n31127 = ~pi609 & n30937;
  assign n31128 = pi1155 & ~n31127;
  assign n31129 = ~n31126 & n31128;
  assign n31130 = pi660 & ~n31004;
  assign n31131 = ~n31129 & n31130;
  assign n31132 = ~n31125 & ~n31131;
  assign n31133 = pi785 & ~n31132;
  assign n31134 = ~pi785 & ~n31119;
  assign n31135 = ~n31133 & ~n31134;
  assign n31136 = ~pi618 & ~n31135;
  assign n31137 = pi618 & n30940;
  assign n31138 = ~pi1154 & ~n31137;
  assign n31139 = ~n31136 & n31138;
  assign n31140 = ~pi627 & ~n31012;
  assign n31141 = ~n31139 & n31140;
  assign n31142 = pi618 & ~n31135;
  assign n31143 = ~pi618 & n30940;
  assign n31144 = pi1154 & ~n31143;
  assign n31145 = ~n31142 & n31144;
  assign n31146 = pi627 & ~n31016;
  assign n31147 = ~n31145 & n31146;
  assign n31148 = ~n31141 & ~n31147;
  assign n31149 = pi781 & ~n31148;
  assign n31150 = ~pi781 & ~n31135;
  assign n31151 = ~n31149 & ~n31150;
  assign n31152 = ~pi619 & ~n31151;
  assign n31153 = pi619 & ~n30943;
  assign n31154 = ~pi1159 & ~n31153;
  assign n31155 = ~n31152 & n31154;
  assign n31156 = ~pi648 & ~n31024;
  assign n31157 = ~n31155 & n31156;
  assign n31158 = pi619 & ~n31151;
  assign n31159 = ~pi619 & ~n30943;
  assign n31160 = pi1159 & ~n31159;
  assign n31161 = ~n31158 & n31160;
  assign n31162 = pi648 & ~n31028;
  assign n31163 = ~n31161 & n31162;
  assign n31164 = pi789 & ~n31157;
  assign n31165 = ~n31163 & n31164;
  assign n31166 = ~pi789 & n31151;
  assign n31167 = n17905 & ~n31166;
  assign n31168 = ~n31165 & n31167;
  assign n31169 = ~pi626 & ~n31031;
  assign n31170 = pi626 & ~n30910;
  assign n31171 = n17668 & ~n31170;
  assign n31172 = ~n31169 & n31171;
  assign n31173 = pi626 & ~n31031;
  assign n31174 = ~pi626 & ~n30910;
  assign n31175 = n17667 & ~n31174;
  assign n31176 = ~n31173 & n31175;
  assign n31177 = n17792 & n30945;
  assign n31178 = ~n31172 & ~n31177;
  assign n31179 = ~n31176 & n31178;
  assign n31180 = pi788 & ~n31179;
  assign n31181 = ~n20298 & ~n31180;
  assign n31182 = ~n31168 & n31181;
  assign n31183 = ~n31066 & ~n31182;
  assign n31184 = n20300 & ~n31183;
  assign n31185 = n17737 & n30967;
  assign n31186 = n17738 & n30963;
  assign n31187 = ~n20491 & n31037;
  assign n31188 = ~n31185 & ~n31186;
  assign n31189 = ~n31187 & n31188;
  assign n31190 = pi787 & ~n31189;
  assign n31191 = ~n31184 & ~n31190;
  assign n31192 = ~n31060 & n31191;
  assign n31193 = ~n31056 & ~n31192;
  assign n31194 = ~po1038 & ~n31193;
  assign n31195 = ~pi190 & po1038;
  assign n31196 = ~pi832 & ~n31195;
  assign n31197 = ~n31194 & n31196;
  assign po347 = ~n30909 & ~n31197;
  assign n31199 = ~pi191 & ~n2755;
  assign n31200 = pi746 & n16933;
  assign n31201 = ~n31199 & ~n31200;
  assign n31202 = ~n17794 & ~n31201;
  assign n31203 = ~pi785 & ~n31202;
  assign n31204 = n17539 & n31200;
  assign n31205 = n31202 & ~n31204;
  assign n31206 = pi1155 & ~n31205;
  assign n31207 = ~pi1155 & ~n31199;
  assign n31208 = ~n31204 & n31207;
  assign n31209 = ~n31206 & ~n31208;
  assign n31210 = pi785 & ~n31209;
  assign n31211 = ~n31203 & ~n31210;
  assign n31212 = ~pi781 & ~n31211;
  assign n31213 = ~n17809 & n31211;
  assign n31214 = pi1154 & ~n31213;
  assign n31215 = ~n17812 & n31211;
  assign n31216 = ~pi1154 & ~n31215;
  assign n31217 = ~n31214 & ~n31216;
  assign n31218 = pi781 & ~n31217;
  assign n31219 = ~n31212 & ~n31218;
  assign n31220 = ~pi789 & ~n31219;
  assign n31221 = ~n22988 & n31219;
  assign n31222 = pi1159 & ~n31221;
  assign n31223 = ~n22991 & n31219;
  assign n31224 = ~pi1159 & ~n31223;
  assign n31225 = ~n31222 & ~n31224;
  assign n31226 = pi789 & ~n31225;
  assign n31227 = ~n31220 & ~n31226;
  assign n31228 = ~n17904 & n31227;
  assign n31229 = n17904 & n31199;
  assign n31230 = ~n31228 & ~n31229;
  assign n31231 = ~n17698 & ~n31230;
  assign n31232 = n17698 & n31199;
  assign n31233 = ~n31231 & ~n31232;
  assign n31234 = ~n20491 & n31233;
  assign n31235 = pi729 & n17153;
  assign n31236 = ~n31199 & ~n31235;
  assign n31237 = ~pi778 & ~n31236;
  assign n31238 = ~pi625 & n31235;
  assign n31239 = ~n31236 & ~n31238;
  assign n31240 = pi1153 & ~n31239;
  assign n31241 = ~pi1153 & ~n31199;
  assign n31242 = ~n31238 & n31241;
  assign n31243 = pi778 & ~n31242;
  assign n31244 = ~n31240 & n31243;
  assign n31245 = ~n31237 & ~n31244;
  assign n31246 = ~n17780 & ~n31245;
  assign n31247 = ~n17782 & n31246;
  assign n31248 = ~n17784 & n31247;
  assign n31249 = ~n17916 & n31248;
  assign n31250 = ~n17947 & n31249;
  assign n31251 = ~pi647 & n31250;
  assign n31252 = pi647 & n31199;
  assign n31253 = ~pi1157 & ~n31252;
  assign n31254 = ~n31251 & n31253;
  assign n31255 = pi647 & ~n31250;
  assign n31256 = ~pi647 & ~n31199;
  assign n31257 = ~n31255 & ~n31256;
  assign n31258 = pi1157 & ~n31257;
  assign n31259 = ~n31254 & ~n31258;
  assign n31260 = ~n17739 & ~n31259;
  assign n31261 = ~n31234 & ~n31260;
  assign n31262 = pi787 & ~n31261;
  assign n31263 = ~pi626 & ~n31227;
  assign n31264 = pi626 & ~n31199;
  assign n31265 = n17668 & ~n31264;
  assign n31266 = ~n31263 & n31265;
  assign n31267 = pi626 & ~n31227;
  assign n31268 = ~pi626 & ~n31199;
  assign n31269 = n17667 & ~n31268;
  assign n31270 = ~n31267 & n31269;
  assign n31271 = n17792 & n31248;
  assign n31272 = ~n31266 & ~n31271;
  assign n31273 = ~n31270 & n31272;
  assign n31274 = pi788 & ~n31273;
  assign n31275 = ~n16842 & ~n31236;
  assign n31276 = pi625 & n31275;
  assign n31277 = n31201 & ~n31275;
  assign n31278 = ~n31276 & ~n31277;
  assign n31279 = n31241 & ~n31278;
  assign n31280 = ~pi608 & ~n31240;
  assign n31281 = ~n31279 & n31280;
  assign n31282 = pi1153 & n31201;
  assign n31283 = ~n31276 & n31282;
  assign n31284 = pi608 & ~n31242;
  assign n31285 = ~n31283 & n31284;
  assign n31286 = ~n31281 & ~n31285;
  assign n31287 = pi778 & ~n31286;
  assign n31288 = ~pi778 & ~n31277;
  assign n31289 = ~n31287 & ~n31288;
  assign n31290 = ~pi609 & ~n31289;
  assign n31291 = pi609 & ~n31245;
  assign n31292 = ~pi1155 & ~n31291;
  assign n31293 = ~n31290 & n31292;
  assign n31294 = ~pi660 & ~n31206;
  assign n31295 = ~n31293 & n31294;
  assign n31296 = pi609 & ~n31289;
  assign n31297 = ~pi609 & ~n31245;
  assign n31298 = pi1155 & ~n31297;
  assign n31299 = ~n31296 & n31298;
  assign n31300 = pi660 & ~n31208;
  assign n31301 = ~n31299 & n31300;
  assign n31302 = ~n31295 & ~n31301;
  assign n31303 = pi785 & ~n31302;
  assign n31304 = ~pi785 & ~n31289;
  assign n31305 = ~n31303 & ~n31304;
  assign n31306 = ~pi618 & ~n31305;
  assign n31307 = pi618 & n31246;
  assign n31308 = ~pi1154 & ~n31307;
  assign n31309 = ~n31306 & n31308;
  assign n31310 = ~pi627 & ~n31214;
  assign n31311 = ~n31309 & n31310;
  assign n31312 = pi618 & ~n31305;
  assign n31313 = ~pi618 & n31246;
  assign n31314 = pi1154 & ~n31313;
  assign n31315 = ~n31312 & n31314;
  assign n31316 = pi627 & ~n31216;
  assign n31317 = ~n31315 & n31316;
  assign n31318 = ~n31311 & ~n31317;
  assign n31319 = pi781 & ~n31318;
  assign n31320 = ~pi781 & ~n31305;
  assign n31321 = ~n31319 & ~n31320;
  assign n31322 = ~pi619 & ~n31321;
  assign n31323 = pi619 & n31247;
  assign n31324 = ~pi1159 & ~n31323;
  assign n31325 = ~n31322 & n31324;
  assign n31326 = ~pi648 & ~n31222;
  assign n31327 = ~n31325 & n31326;
  assign n31328 = pi619 & ~n31321;
  assign n31329 = ~pi619 & n31247;
  assign n31330 = pi1159 & ~n31329;
  assign n31331 = ~n31328 & n31330;
  assign n31332 = pi648 & ~n31224;
  assign n31333 = ~n31331 & n31332;
  assign n31334 = pi789 & ~n31327;
  assign n31335 = ~n31333 & n31334;
  assign n31336 = ~pi789 & n31321;
  assign n31337 = n17905 & ~n31336;
  assign n31338 = ~n31335 & n31337;
  assign n31339 = ~n31274 & ~n31338;
  assign n31340 = ~n20298 & ~n31339;
  assign n31341 = n17944 & ~n31230;
  assign n31342 = n20786 & n31249;
  assign n31343 = ~n31341 & ~n31342;
  assign n31344 = ~pi629 & ~n31343;
  assign n31345 = n20790 & n31249;
  assign n31346 = n17943 & ~n31230;
  assign n31347 = ~n31345 & ~n31346;
  assign n31348 = pi629 & ~n31347;
  assign n31349 = ~n31344 & ~n31348;
  assign n31350 = pi792 & ~n31349;
  assign n31351 = n20300 & ~n31350;
  assign n31352 = ~n31340 & n31351;
  assign n31353 = ~n31262 & ~n31352;
  assign n31354 = pi644 & n31353;
  assign n31355 = ~pi787 & ~n31250;
  assign n31356 = pi787 & ~n31259;
  assign n31357 = ~n31355 & ~n31356;
  assign n31358 = ~pi644 & n31357;
  assign n31359 = pi715 & ~n31358;
  assign n31360 = ~n31354 & n31359;
  assign n31361 = ~n17740 & ~n31233;
  assign n31362 = n17740 & n31199;
  assign n31363 = ~n31361 & ~n31362;
  assign n31364 = pi644 & ~n31363;
  assign n31365 = ~pi644 & n31199;
  assign n31366 = ~pi715 & ~n31365;
  assign n31367 = ~n31364 & n31366;
  assign n31368 = pi1160 & ~n31367;
  assign n31369 = ~n31360 & n31368;
  assign n31370 = ~pi644 & n31353;
  assign n31371 = pi644 & n31357;
  assign n31372 = ~pi715 & ~n31371;
  assign n31373 = ~n31370 & n31372;
  assign n31374 = ~pi644 & ~n31363;
  assign n31375 = pi644 & n31199;
  assign n31376 = pi715 & ~n31375;
  assign n31377 = ~n31374 & n31376;
  assign n31378 = ~pi1160 & ~n31377;
  assign n31379 = ~n31373 & n31378;
  assign n31380 = ~n31369 & ~n31379;
  assign n31381 = pi790 & ~n31380;
  assign n31382 = ~pi790 & n31353;
  assign n31383 = pi832 & ~n31382;
  assign n31384 = ~n31381 & n31383;
  assign n31385 = ~pi191 & ~n17494;
  assign n31386 = n17627 & ~n31385;
  assign n31387 = pi191 & ~n3268;
  assign n31388 = ~pi191 & n18060;
  assign n31389 = pi191 & ~n18064;
  assign n31390 = ~pi38 & ~n31389;
  assign n31391 = ~n31388 & n31390;
  assign n31392 = ~pi191 & ~n16968;
  assign n31393 = n17480 & ~n31392;
  assign n31394 = pi729 & ~n31393;
  assign n31395 = ~n31391 & n31394;
  assign n31396 = ~pi191 & ~pi729;
  assign n31397 = ~n17487 & n31396;
  assign n31398 = n3268 & ~n31397;
  assign n31399 = ~n31395 & n31398;
  assign n31400 = ~n31387 & ~n31399;
  assign n31401 = ~pi778 & ~n31400;
  assign n31402 = pi625 & n31400;
  assign n31403 = ~pi625 & n31385;
  assign n31404 = pi1153 & ~n31403;
  assign n31405 = ~n31402 & n31404;
  assign n31406 = ~pi625 & n31400;
  assign n31407 = pi625 & n31385;
  assign n31408 = ~pi1153 & ~n31407;
  assign n31409 = ~n31406 & n31408;
  assign n31410 = ~n31405 & ~n31409;
  assign n31411 = pi778 & ~n31410;
  assign n31412 = ~n31401 & ~n31411;
  assign n31413 = ~n17554 & ~n31412;
  assign n31414 = n17554 & ~n31385;
  assign n31415 = ~n31413 & ~n31414;
  assign n31416 = ~n17591 & n31415;
  assign n31417 = n17591 & n31385;
  assign n31418 = ~n31416 & ~n31417;
  assign n31419 = ~n17627 & n31418;
  assign n31420 = ~n31386 & ~n31419;
  assign n31421 = ~n17670 & n31420;
  assign n31422 = n17670 & n31385;
  assign n31423 = ~n31421 & ~n31422;
  assign n31424 = ~pi628 & ~n31423;
  assign n31425 = pi628 & n31385;
  assign n31426 = ~n31424 & ~n31425;
  assign n31427 = ~pi1156 & ~n31426;
  assign n31428 = pi628 & ~n31423;
  assign n31429 = ~pi628 & n31385;
  assign n31430 = ~n31428 & ~n31429;
  assign n31431 = pi1156 & ~n31430;
  assign n31432 = ~n31427 & ~n31431;
  assign n31433 = pi792 & ~n31432;
  assign n31434 = ~pi792 & ~n31423;
  assign n31435 = ~n31433 & ~n31434;
  assign n31436 = ~pi647 & ~n31435;
  assign n31437 = pi647 & n31385;
  assign n31438 = ~n31436 & ~n31437;
  assign n31439 = ~pi1157 & ~n31438;
  assign n31440 = pi647 & ~n31435;
  assign n31441 = ~pi647 & n31385;
  assign n31442 = ~n31440 & ~n31441;
  assign n31443 = pi1157 & ~n31442;
  assign n31444 = ~n31439 & ~n31443;
  assign n31445 = pi787 & ~n31444;
  assign n31446 = ~pi787 & ~n31435;
  assign n31447 = ~n31445 & ~n31446;
  assign n31448 = ~pi644 & ~n31447;
  assign n31449 = pi715 & ~n31448;
  assign n31450 = ~pi746 & n16814;
  assign n31451 = pi191 & n16961;
  assign n31452 = ~n31450 & ~n31451;
  assign n31453 = pi39 & ~n31452;
  assign n31454 = ~pi191 & pi746;
  assign n31455 = n16907 & n31454;
  assign n31456 = pi746 & ~n16919;
  assign n31457 = pi191 & ~n31456;
  assign n31458 = ~n22368 & ~n31457;
  assign n31459 = ~n31455 & n31458;
  assign n31460 = ~n31453 & n31459;
  assign n31461 = ~pi38 & ~n31460;
  assign n31462 = pi746 & n16970;
  assign n31463 = pi38 & ~n31392;
  assign n31464 = ~n31462 & n31463;
  assign n31465 = ~n31461 & ~n31464;
  assign n31466 = n3268 & ~n31465;
  assign n31467 = ~n31387 & ~n31466;
  assign n31468 = ~n17526 & ~n31467;
  assign n31469 = n17526 & ~n31385;
  assign n31470 = ~n31468 & ~n31469;
  assign n31471 = ~pi785 & ~n31470;
  assign n31472 = ~n17527 & ~n31385;
  assign n31473 = pi609 & n31468;
  assign n31474 = ~n31472 & ~n31473;
  assign n31475 = pi1155 & ~n31474;
  assign n31476 = ~n17539 & ~n31385;
  assign n31477 = ~pi609 & n31468;
  assign n31478 = ~n31476 & ~n31477;
  assign n31479 = ~pi1155 & ~n31478;
  assign n31480 = ~n31475 & ~n31479;
  assign n31481 = pi785 & ~n31480;
  assign n31482 = ~n31471 & ~n31481;
  assign n31483 = ~pi781 & ~n31482;
  assign n31484 = pi618 & n31482;
  assign n31485 = ~pi618 & n31385;
  assign n31486 = pi1154 & ~n31485;
  assign n31487 = ~n31484 & n31486;
  assign n31488 = ~pi618 & n31482;
  assign n31489 = pi618 & n31385;
  assign n31490 = ~pi1154 & ~n31489;
  assign n31491 = ~n31488 & n31490;
  assign n31492 = ~n31487 & ~n31491;
  assign n31493 = pi781 & ~n31492;
  assign n31494 = ~n31483 & ~n31493;
  assign n31495 = ~pi789 & ~n31494;
  assign n31496 = pi619 & n31494;
  assign n31497 = ~pi619 & n31385;
  assign n31498 = pi1159 & ~n31497;
  assign n31499 = ~n31496 & n31498;
  assign n31500 = ~pi619 & n31494;
  assign n31501 = pi619 & n31385;
  assign n31502 = ~pi1159 & ~n31501;
  assign n31503 = ~n31500 & n31502;
  assign n31504 = ~n31499 & ~n31503;
  assign n31505 = pi789 & ~n31504;
  assign n31506 = ~n31495 & ~n31505;
  assign n31507 = ~n17904 & n31506;
  assign n31508 = n17904 & n31385;
  assign n31509 = ~n31507 & ~n31508;
  assign n31510 = ~n17698 & ~n31509;
  assign n31511 = n17698 & n31385;
  assign n31512 = ~n31510 & ~n31511;
  assign n31513 = ~n17740 & ~n31512;
  assign n31514 = n17740 & n31385;
  assign n31515 = ~n31513 & ~n31514;
  assign n31516 = pi644 & ~n31515;
  assign n31517 = ~pi644 & n31385;
  assign n31518 = ~pi715 & ~n31517;
  assign n31519 = ~n31516 & n31518;
  assign n31520 = pi1160 & ~n31519;
  assign n31521 = ~n31449 & n31520;
  assign n31522 = pi644 & ~n31447;
  assign n31523 = ~pi715 & ~n31522;
  assign n31524 = ~pi644 & ~n31515;
  assign n31525 = pi644 & n31385;
  assign n31526 = pi715 & ~n31525;
  assign n31527 = ~n31524 & n31526;
  assign n31528 = ~pi1160 & ~n31527;
  assign n31529 = ~n31523 & n31528;
  assign n31530 = ~n31521 & ~n31529;
  assign n31531 = pi790 & ~n31530;
  assign n31532 = ~pi644 & n31528;
  assign n31533 = pi644 & n31520;
  assign n31534 = pi790 & ~n31532;
  assign n31535 = ~n31533 & n31534;
  assign n31536 = ~n20502 & n31509;
  assign n31537 = n17696 & n31426;
  assign n31538 = n17695 & n31430;
  assign n31539 = ~n31537 & ~n31538;
  assign n31540 = ~n31536 & n31539;
  assign n31541 = pi792 & ~n31540;
  assign n31542 = ~pi729 & n31465;
  assign n31543 = ~pi191 & n17074;
  assign n31544 = pi191 & n17166;
  assign n31545 = ~pi746 & ~n31544;
  assign n31546 = ~n31543 & n31545;
  assign n31547 = pi191 & n17233;
  assign n31548 = ~pi191 & ~n17295;
  assign n31549 = pi746 & ~n31548;
  assign n31550 = ~n31547 & n31549;
  assign n31551 = pi39 & ~n31550;
  assign n31552 = ~n31546 & n31551;
  assign n31553 = ~pi191 & n17317;
  assign n31554 = pi191 & n17340;
  assign n31555 = ~pi746 & ~n31553;
  assign n31556 = ~n31554 & n31555;
  assign n31557 = ~pi191 & ~n17344;
  assign n31558 = pi191 & ~n17351;
  assign n31559 = pi746 & ~n31558;
  assign n31560 = ~n31557 & n31559;
  assign n31561 = ~pi39 & ~n31560;
  assign n31562 = ~n31556 & n31561;
  assign n31563 = ~pi38 & ~n31562;
  assign n31564 = ~n31552 & n31563;
  assign n31565 = ~pi746 & n24006;
  assign n31566 = ~n17259 & ~n31565;
  assign n31567 = ~pi39 & ~n31566;
  assign n31568 = ~pi191 & ~n31567;
  assign n31569 = ~n17154 & ~n31200;
  assign n31570 = pi191 & ~n31569;
  assign n31571 = n6250 & n31570;
  assign n31572 = pi38 & ~n31571;
  assign n31573 = ~n31568 & n31572;
  assign n31574 = pi729 & ~n31573;
  assign n31575 = ~n31564 & n31574;
  assign n31576 = n3268 & ~n31575;
  assign n31577 = ~n31542 & n31576;
  assign n31578 = ~n31387 & ~n31577;
  assign n31579 = ~pi625 & n31578;
  assign n31580 = pi625 & n31467;
  assign n31581 = ~pi1153 & ~n31580;
  assign n31582 = ~n31579 & n31581;
  assign n31583 = ~pi608 & ~n31405;
  assign n31584 = ~n31582 & n31583;
  assign n31585 = pi625 & n31578;
  assign n31586 = ~pi625 & n31467;
  assign n31587 = pi1153 & ~n31586;
  assign n31588 = ~n31585 & n31587;
  assign n31589 = pi608 & ~n31409;
  assign n31590 = ~n31588 & n31589;
  assign n31591 = ~n31584 & ~n31590;
  assign n31592 = pi778 & ~n31591;
  assign n31593 = ~pi778 & n31578;
  assign n31594 = ~n31592 & ~n31593;
  assign n31595 = ~pi609 & ~n31594;
  assign n31596 = pi609 & n31412;
  assign n31597 = ~pi1155 & ~n31596;
  assign n31598 = ~n31595 & n31597;
  assign n31599 = ~pi660 & ~n31475;
  assign n31600 = ~n31598 & n31599;
  assign n31601 = pi609 & ~n31594;
  assign n31602 = ~pi609 & n31412;
  assign n31603 = pi1155 & ~n31602;
  assign n31604 = ~n31601 & n31603;
  assign n31605 = pi660 & ~n31479;
  assign n31606 = ~n31604 & n31605;
  assign n31607 = ~n31600 & ~n31606;
  assign n31608 = pi785 & ~n31607;
  assign n31609 = ~pi785 & ~n31594;
  assign n31610 = ~n31608 & ~n31609;
  assign n31611 = ~pi618 & ~n31610;
  assign n31612 = pi618 & n31415;
  assign n31613 = ~pi1154 & ~n31612;
  assign n31614 = ~n31611 & n31613;
  assign n31615 = ~pi627 & ~n31487;
  assign n31616 = ~n31614 & n31615;
  assign n31617 = pi618 & ~n31610;
  assign n31618 = ~pi618 & n31415;
  assign n31619 = pi1154 & ~n31618;
  assign n31620 = ~n31617 & n31619;
  assign n31621 = pi627 & ~n31491;
  assign n31622 = ~n31620 & n31621;
  assign n31623 = ~n31616 & ~n31622;
  assign n31624 = pi781 & ~n31623;
  assign n31625 = ~pi781 & ~n31610;
  assign n31626 = ~n31624 & ~n31625;
  assign n31627 = ~pi619 & ~n31626;
  assign n31628 = pi619 & ~n31418;
  assign n31629 = ~pi1159 & ~n31628;
  assign n31630 = ~n31627 & n31629;
  assign n31631 = ~pi648 & ~n31499;
  assign n31632 = ~n31630 & n31631;
  assign n31633 = pi619 & ~n31626;
  assign n31634 = ~pi619 & ~n31418;
  assign n31635 = pi1159 & ~n31634;
  assign n31636 = ~n31633 & n31635;
  assign n31637 = pi648 & ~n31503;
  assign n31638 = ~n31636 & n31637;
  assign n31639 = pi789 & ~n31632;
  assign n31640 = ~n31638 & n31639;
  assign n31641 = ~pi789 & n31626;
  assign n31642 = n17905 & ~n31641;
  assign n31643 = ~n31640 & n31642;
  assign n31644 = ~pi626 & ~n31506;
  assign n31645 = pi626 & ~n31385;
  assign n31646 = n17668 & ~n31645;
  assign n31647 = ~n31644 & n31646;
  assign n31648 = pi626 & ~n31506;
  assign n31649 = ~pi626 & ~n31385;
  assign n31650 = n17667 & ~n31649;
  assign n31651 = ~n31648 & n31650;
  assign n31652 = n17792 & n31420;
  assign n31653 = ~n31647 & ~n31652;
  assign n31654 = ~n31651 & n31653;
  assign n31655 = pi788 & ~n31654;
  assign n31656 = ~n20298 & ~n31655;
  assign n31657 = ~n31643 & n31656;
  assign n31658 = ~n31541 & ~n31657;
  assign n31659 = n20300 & ~n31658;
  assign n31660 = n17737 & n31442;
  assign n31661 = n17738 & n31438;
  assign n31662 = ~n20491 & n31512;
  assign n31663 = ~n31660 & ~n31661;
  assign n31664 = ~n31662 & n31663;
  assign n31665 = pi787 & ~n31664;
  assign n31666 = ~n31659 & ~n31665;
  assign n31667 = ~n31535 & n31666;
  assign n31668 = ~n31531 & ~n31667;
  assign n31669 = ~po1038 & ~n31668;
  assign n31670 = ~pi191 & po1038;
  assign n31671 = ~pi832 & ~n31670;
  assign n31672 = ~n31669 & n31671;
  assign po348 = ~n31384 & ~n31672;
  assign n31674 = ~pi192 & ~n2755;
  assign n31675 = pi764 & n16933;
  assign n31676 = ~n31674 & ~n31675;
  assign n31677 = ~n17794 & ~n31676;
  assign n31678 = ~pi785 & ~n31677;
  assign n31679 = n17539 & n31675;
  assign n31680 = n31677 & ~n31679;
  assign n31681 = pi1155 & ~n31680;
  assign n31682 = ~pi1155 & ~n31674;
  assign n31683 = ~n31679 & n31682;
  assign n31684 = ~n31681 & ~n31683;
  assign n31685 = pi785 & ~n31684;
  assign n31686 = ~n31678 & ~n31685;
  assign n31687 = ~pi781 & ~n31686;
  assign n31688 = ~n17809 & n31686;
  assign n31689 = pi1154 & ~n31688;
  assign n31690 = ~n17812 & n31686;
  assign n31691 = ~pi1154 & ~n31690;
  assign n31692 = ~n31689 & ~n31691;
  assign n31693 = pi781 & ~n31692;
  assign n31694 = ~n31687 & ~n31693;
  assign n31695 = ~pi789 & ~n31694;
  assign n31696 = ~n22988 & n31694;
  assign n31697 = pi1159 & ~n31696;
  assign n31698 = ~n22991 & n31694;
  assign n31699 = ~pi1159 & ~n31698;
  assign n31700 = ~n31697 & ~n31699;
  assign n31701 = pi789 & ~n31700;
  assign n31702 = ~n31695 & ~n31701;
  assign n31703 = ~n17904 & n31702;
  assign n31704 = n17904 & n31674;
  assign n31705 = ~n31703 & ~n31704;
  assign n31706 = ~n17698 & ~n31705;
  assign n31707 = n17698 & n31674;
  assign n31708 = ~n31706 & ~n31707;
  assign n31709 = ~n20491 & n31708;
  assign n31710 = pi691 & n17153;
  assign n31711 = ~n31674 & ~n31710;
  assign n31712 = ~pi778 & ~n31711;
  assign n31713 = ~pi625 & n31710;
  assign n31714 = ~n31711 & ~n31713;
  assign n31715 = pi1153 & ~n31714;
  assign n31716 = ~pi1153 & ~n31674;
  assign n31717 = ~n31713 & n31716;
  assign n31718 = pi778 & ~n31717;
  assign n31719 = ~n31715 & n31718;
  assign n31720 = ~n31712 & ~n31719;
  assign n31721 = ~n17780 & ~n31720;
  assign n31722 = ~n17782 & n31721;
  assign n31723 = ~n17784 & n31722;
  assign n31724 = ~n17916 & n31723;
  assign n31725 = ~n17947 & n31724;
  assign n31726 = ~pi647 & n31725;
  assign n31727 = pi647 & n31674;
  assign n31728 = ~pi1157 & ~n31727;
  assign n31729 = ~n31726 & n31728;
  assign n31730 = pi647 & ~n31725;
  assign n31731 = ~pi647 & ~n31674;
  assign n31732 = ~n31730 & ~n31731;
  assign n31733 = pi1157 & ~n31732;
  assign n31734 = ~n31729 & ~n31733;
  assign n31735 = ~n17739 & ~n31734;
  assign n31736 = ~n31709 & ~n31735;
  assign n31737 = pi787 & ~n31736;
  assign n31738 = ~pi626 & ~n31702;
  assign n31739 = pi626 & ~n31674;
  assign n31740 = n17668 & ~n31739;
  assign n31741 = ~n31738 & n31740;
  assign n31742 = pi626 & ~n31702;
  assign n31743 = ~pi626 & ~n31674;
  assign n31744 = n17667 & ~n31743;
  assign n31745 = ~n31742 & n31744;
  assign n31746 = n17792 & n31723;
  assign n31747 = ~n31741 & ~n31746;
  assign n31748 = ~n31745 & n31747;
  assign n31749 = pi788 & ~n31748;
  assign n31750 = ~n16842 & ~n31711;
  assign n31751 = pi625 & n31750;
  assign n31752 = n31676 & ~n31750;
  assign n31753 = ~n31751 & ~n31752;
  assign n31754 = n31716 & ~n31753;
  assign n31755 = ~pi608 & ~n31715;
  assign n31756 = ~n31754 & n31755;
  assign n31757 = pi1153 & n31676;
  assign n31758 = ~n31751 & n31757;
  assign n31759 = pi608 & ~n31717;
  assign n31760 = ~n31758 & n31759;
  assign n31761 = ~n31756 & ~n31760;
  assign n31762 = pi778 & ~n31761;
  assign n31763 = ~pi778 & ~n31752;
  assign n31764 = ~n31762 & ~n31763;
  assign n31765 = ~pi609 & ~n31764;
  assign n31766 = pi609 & ~n31720;
  assign n31767 = ~pi1155 & ~n31766;
  assign n31768 = ~n31765 & n31767;
  assign n31769 = ~pi660 & ~n31681;
  assign n31770 = ~n31768 & n31769;
  assign n31771 = pi609 & ~n31764;
  assign n31772 = ~pi609 & ~n31720;
  assign n31773 = pi1155 & ~n31772;
  assign n31774 = ~n31771 & n31773;
  assign n31775 = pi660 & ~n31683;
  assign n31776 = ~n31774 & n31775;
  assign n31777 = ~n31770 & ~n31776;
  assign n31778 = pi785 & ~n31777;
  assign n31779 = ~pi785 & ~n31764;
  assign n31780 = ~n31778 & ~n31779;
  assign n31781 = ~pi618 & ~n31780;
  assign n31782 = pi618 & n31721;
  assign n31783 = ~pi1154 & ~n31782;
  assign n31784 = ~n31781 & n31783;
  assign n31785 = ~pi627 & ~n31689;
  assign n31786 = ~n31784 & n31785;
  assign n31787 = pi618 & ~n31780;
  assign n31788 = ~pi618 & n31721;
  assign n31789 = pi1154 & ~n31788;
  assign n31790 = ~n31787 & n31789;
  assign n31791 = pi627 & ~n31691;
  assign n31792 = ~n31790 & n31791;
  assign n31793 = ~n31786 & ~n31792;
  assign n31794 = pi781 & ~n31793;
  assign n31795 = ~pi781 & ~n31780;
  assign n31796 = ~n31794 & ~n31795;
  assign n31797 = ~pi619 & ~n31796;
  assign n31798 = pi619 & n31722;
  assign n31799 = ~pi1159 & ~n31798;
  assign n31800 = ~n31797 & n31799;
  assign n31801 = ~pi648 & ~n31697;
  assign n31802 = ~n31800 & n31801;
  assign n31803 = pi619 & ~n31796;
  assign n31804 = ~pi619 & n31722;
  assign n31805 = pi1159 & ~n31804;
  assign n31806 = ~n31803 & n31805;
  assign n31807 = pi648 & ~n31699;
  assign n31808 = ~n31806 & n31807;
  assign n31809 = pi789 & ~n31802;
  assign n31810 = ~n31808 & n31809;
  assign n31811 = ~pi789 & n31796;
  assign n31812 = n17905 & ~n31811;
  assign n31813 = ~n31810 & n31812;
  assign n31814 = ~n31749 & ~n31813;
  assign n31815 = ~n20298 & ~n31814;
  assign n31816 = n17944 & ~n31705;
  assign n31817 = n20786 & n31724;
  assign n31818 = ~n31816 & ~n31817;
  assign n31819 = ~pi629 & ~n31818;
  assign n31820 = n20790 & n31724;
  assign n31821 = n17943 & ~n31705;
  assign n31822 = ~n31820 & ~n31821;
  assign n31823 = pi629 & ~n31822;
  assign n31824 = ~n31819 & ~n31823;
  assign n31825 = pi792 & ~n31824;
  assign n31826 = n20300 & ~n31825;
  assign n31827 = ~n31815 & n31826;
  assign n31828 = ~n31737 & ~n31827;
  assign n31829 = pi644 & n31828;
  assign n31830 = ~pi787 & ~n31725;
  assign n31831 = pi787 & ~n31734;
  assign n31832 = ~n31830 & ~n31831;
  assign n31833 = ~pi644 & n31832;
  assign n31834 = pi715 & ~n31833;
  assign n31835 = ~n31829 & n31834;
  assign n31836 = ~n17740 & ~n31708;
  assign n31837 = n17740 & n31674;
  assign n31838 = ~n31836 & ~n31837;
  assign n31839 = pi644 & ~n31838;
  assign n31840 = ~pi644 & n31674;
  assign n31841 = ~pi715 & ~n31840;
  assign n31842 = ~n31839 & n31841;
  assign n31843 = pi1160 & ~n31842;
  assign n31844 = ~n31835 & n31843;
  assign n31845 = ~pi644 & n31828;
  assign n31846 = pi644 & n31832;
  assign n31847 = ~pi715 & ~n31846;
  assign n31848 = ~n31845 & n31847;
  assign n31849 = ~pi644 & ~n31838;
  assign n31850 = pi644 & n31674;
  assign n31851 = pi715 & ~n31850;
  assign n31852 = ~n31849 & n31851;
  assign n31853 = ~pi1160 & ~n31852;
  assign n31854 = ~n31848 & n31853;
  assign n31855 = ~n31844 & ~n31854;
  assign n31856 = pi790 & ~n31855;
  assign n31857 = ~pi790 & n31828;
  assign n31858 = pi832 & ~n31857;
  assign n31859 = ~n31856 & n31858;
  assign n31860 = ~pi192 & ~n17494;
  assign n31861 = n17627 & ~n31860;
  assign n31862 = pi192 & ~n3268;
  assign n31863 = ~pi192 & n18060;
  assign n31864 = pi192 & ~n18064;
  assign n31865 = ~pi38 & ~n31864;
  assign n31866 = ~n31863 & n31865;
  assign n31867 = ~pi192 & ~n16968;
  assign n31868 = n17480 & ~n31867;
  assign n31869 = pi691 & ~n31868;
  assign n31870 = ~n31866 & n31869;
  assign n31871 = ~pi192 & ~pi691;
  assign n31872 = ~n17487 & n31871;
  assign n31873 = n3268 & ~n31872;
  assign n31874 = ~n31870 & n31873;
  assign n31875 = ~n31862 & ~n31874;
  assign n31876 = ~pi778 & ~n31875;
  assign n31877 = pi625 & n31875;
  assign n31878 = ~pi625 & n31860;
  assign n31879 = pi1153 & ~n31878;
  assign n31880 = ~n31877 & n31879;
  assign n31881 = ~pi625 & n31875;
  assign n31882 = pi625 & n31860;
  assign n31883 = ~pi1153 & ~n31882;
  assign n31884 = ~n31881 & n31883;
  assign n31885 = ~n31880 & ~n31884;
  assign n31886 = pi778 & ~n31885;
  assign n31887 = ~n31876 & ~n31886;
  assign n31888 = ~n17554 & ~n31887;
  assign n31889 = n17554 & ~n31860;
  assign n31890 = ~n31888 & ~n31889;
  assign n31891 = ~n17591 & n31890;
  assign n31892 = n17591 & n31860;
  assign n31893 = ~n31891 & ~n31892;
  assign n31894 = ~n17627 & n31893;
  assign n31895 = ~n31861 & ~n31894;
  assign n31896 = ~n17670 & n31895;
  assign n31897 = n17670 & n31860;
  assign n31898 = ~n31896 & ~n31897;
  assign n31899 = ~pi628 & ~n31898;
  assign n31900 = pi628 & n31860;
  assign n31901 = ~n31899 & ~n31900;
  assign n31902 = ~pi1156 & ~n31901;
  assign n31903 = pi628 & ~n31898;
  assign n31904 = ~pi628 & n31860;
  assign n31905 = ~n31903 & ~n31904;
  assign n31906 = pi1156 & ~n31905;
  assign n31907 = ~n31902 & ~n31906;
  assign n31908 = pi792 & ~n31907;
  assign n31909 = ~pi792 & ~n31898;
  assign n31910 = ~n31908 & ~n31909;
  assign n31911 = ~pi647 & ~n31910;
  assign n31912 = pi647 & n31860;
  assign n31913 = ~n31911 & ~n31912;
  assign n31914 = ~pi1157 & ~n31913;
  assign n31915 = pi647 & ~n31910;
  assign n31916 = ~pi647 & n31860;
  assign n31917 = ~n31915 & ~n31916;
  assign n31918 = pi1157 & ~n31917;
  assign n31919 = ~n31914 & ~n31918;
  assign n31920 = pi787 & ~n31919;
  assign n31921 = ~pi787 & ~n31910;
  assign n31922 = ~n31920 & ~n31921;
  assign n31923 = ~pi644 & ~n31922;
  assign n31924 = pi715 & ~n31923;
  assign n31925 = ~pi764 & n16814;
  assign n31926 = pi192 & n16961;
  assign n31927 = ~n31925 & ~n31926;
  assign n31928 = pi39 & ~n31927;
  assign n31929 = ~pi192 & pi764;
  assign n31930 = n16907 & n31929;
  assign n31931 = pi764 & ~n16919;
  assign n31932 = pi192 & ~n31931;
  assign n31933 = ~n22529 & ~n31932;
  assign n31934 = ~n31930 & n31933;
  assign n31935 = ~n31928 & n31934;
  assign n31936 = ~pi38 & ~n31935;
  assign n31937 = pi764 & n16970;
  assign n31938 = pi38 & ~n31867;
  assign n31939 = ~n31937 & n31938;
  assign n31940 = ~n31936 & ~n31939;
  assign n31941 = n3268 & ~n31940;
  assign n31942 = ~n31862 & ~n31941;
  assign n31943 = ~n17526 & ~n31942;
  assign n31944 = n17526 & ~n31860;
  assign n31945 = ~n31943 & ~n31944;
  assign n31946 = ~pi785 & ~n31945;
  assign n31947 = ~n17527 & ~n31860;
  assign n31948 = pi609 & n31943;
  assign n31949 = ~n31947 & ~n31948;
  assign n31950 = pi1155 & ~n31949;
  assign n31951 = ~n17539 & ~n31860;
  assign n31952 = ~pi609 & n31943;
  assign n31953 = ~n31951 & ~n31952;
  assign n31954 = ~pi1155 & ~n31953;
  assign n31955 = ~n31950 & ~n31954;
  assign n31956 = pi785 & ~n31955;
  assign n31957 = ~n31946 & ~n31956;
  assign n31958 = ~pi781 & ~n31957;
  assign n31959 = pi618 & n31957;
  assign n31960 = ~pi618 & n31860;
  assign n31961 = pi1154 & ~n31960;
  assign n31962 = ~n31959 & n31961;
  assign n31963 = ~pi618 & n31957;
  assign n31964 = pi618 & n31860;
  assign n31965 = ~pi1154 & ~n31964;
  assign n31966 = ~n31963 & n31965;
  assign n31967 = ~n31962 & ~n31966;
  assign n31968 = pi781 & ~n31967;
  assign n31969 = ~n31958 & ~n31968;
  assign n31970 = ~pi789 & ~n31969;
  assign n31971 = pi619 & n31969;
  assign n31972 = ~pi619 & n31860;
  assign n31973 = pi1159 & ~n31972;
  assign n31974 = ~n31971 & n31973;
  assign n31975 = ~pi619 & n31969;
  assign n31976 = pi619 & n31860;
  assign n31977 = ~pi1159 & ~n31976;
  assign n31978 = ~n31975 & n31977;
  assign n31979 = ~n31974 & ~n31978;
  assign n31980 = pi789 & ~n31979;
  assign n31981 = ~n31970 & ~n31980;
  assign n31982 = ~n17904 & n31981;
  assign n31983 = n17904 & n31860;
  assign n31984 = ~n31982 & ~n31983;
  assign n31985 = ~n17698 & ~n31984;
  assign n31986 = n17698 & n31860;
  assign n31987 = ~n31985 & ~n31986;
  assign n31988 = ~n17740 & ~n31987;
  assign n31989 = n17740 & n31860;
  assign n31990 = ~n31988 & ~n31989;
  assign n31991 = pi644 & ~n31990;
  assign n31992 = ~pi644 & n31860;
  assign n31993 = ~pi715 & ~n31992;
  assign n31994 = ~n31991 & n31993;
  assign n31995 = pi1160 & ~n31994;
  assign n31996 = ~n31924 & n31995;
  assign n31997 = pi644 & ~n31922;
  assign n31998 = ~pi715 & ~n31997;
  assign n31999 = ~pi644 & ~n31990;
  assign n32000 = pi644 & n31860;
  assign n32001 = pi715 & ~n32000;
  assign n32002 = ~n31999 & n32001;
  assign n32003 = ~pi1160 & ~n32002;
  assign n32004 = ~n31998 & n32003;
  assign n32005 = ~n31996 & ~n32004;
  assign n32006 = pi790 & ~n32005;
  assign n32007 = ~pi644 & n32003;
  assign n32008 = pi644 & n31995;
  assign n32009 = pi790 & ~n32007;
  assign n32010 = ~n32008 & n32009;
  assign n32011 = ~n20502 & n31984;
  assign n32012 = n17696 & n31901;
  assign n32013 = n17695 & n31905;
  assign n32014 = ~n32012 & ~n32013;
  assign n32015 = ~n32011 & n32014;
  assign n32016 = pi792 & ~n32015;
  assign n32017 = ~pi691 & n31940;
  assign n32018 = ~pi192 & n17074;
  assign n32019 = pi192 & n17166;
  assign n32020 = ~pi764 & ~n32019;
  assign n32021 = ~n32018 & n32020;
  assign n32022 = pi192 & n17233;
  assign n32023 = ~pi192 & ~n17295;
  assign n32024 = pi764 & ~n32023;
  assign n32025 = ~n32022 & n32024;
  assign n32026 = pi39 & ~n32025;
  assign n32027 = ~n32021 & n32026;
  assign n32028 = ~pi192 & n17317;
  assign n32029 = pi192 & n17340;
  assign n32030 = ~pi764 & ~n32028;
  assign n32031 = ~n32029 & n32030;
  assign n32032 = ~pi192 & ~n17344;
  assign n32033 = pi192 & ~n17351;
  assign n32034 = pi764 & ~n32033;
  assign n32035 = ~n32032 & n32034;
  assign n32036 = ~pi39 & ~n32035;
  assign n32037 = ~n32031 & n32036;
  assign n32038 = ~pi38 & ~n32037;
  assign n32039 = ~n32027 & n32038;
  assign n32040 = ~pi764 & n24006;
  assign n32041 = ~n17259 & ~n32040;
  assign n32042 = ~pi39 & ~n32041;
  assign n32043 = ~pi192 & ~n32042;
  assign n32044 = ~n17154 & ~n31675;
  assign n32045 = pi192 & ~n32044;
  assign n32046 = n6250 & n32045;
  assign n32047 = pi38 & ~n32046;
  assign n32048 = ~n32043 & n32047;
  assign n32049 = pi691 & ~n32048;
  assign n32050 = ~n32039 & n32049;
  assign n32051 = n3268 & ~n32050;
  assign n32052 = ~n32017 & n32051;
  assign n32053 = ~n31862 & ~n32052;
  assign n32054 = ~pi625 & n32053;
  assign n32055 = pi625 & n31942;
  assign n32056 = ~pi1153 & ~n32055;
  assign n32057 = ~n32054 & n32056;
  assign n32058 = ~pi608 & ~n31880;
  assign n32059 = ~n32057 & n32058;
  assign n32060 = pi625 & n32053;
  assign n32061 = ~pi625 & n31942;
  assign n32062 = pi1153 & ~n32061;
  assign n32063 = ~n32060 & n32062;
  assign n32064 = pi608 & ~n31884;
  assign n32065 = ~n32063 & n32064;
  assign n32066 = ~n32059 & ~n32065;
  assign n32067 = pi778 & ~n32066;
  assign n32068 = ~pi778 & n32053;
  assign n32069 = ~n32067 & ~n32068;
  assign n32070 = ~pi609 & ~n32069;
  assign n32071 = pi609 & n31887;
  assign n32072 = ~pi1155 & ~n32071;
  assign n32073 = ~n32070 & n32072;
  assign n32074 = ~pi660 & ~n31950;
  assign n32075 = ~n32073 & n32074;
  assign n32076 = pi609 & ~n32069;
  assign n32077 = ~pi609 & n31887;
  assign n32078 = pi1155 & ~n32077;
  assign n32079 = ~n32076 & n32078;
  assign n32080 = pi660 & ~n31954;
  assign n32081 = ~n32079 & n32080;
  assign n32082 = ~n32075 & ~n32081;
  assign n32083 = pi785 & ~n32082;
  assign n32084 = ~pi785 & ~n32069;
  assign n32085 = ~n32083 & ~n32084;
  assign n32086 = ~pi618 & ~n32085;
  assign n32087 = pi618 & n31890;
  assign n32088 = ~pi1154 & ~n32087;
  assign n32089 = ~n32086 & n32088;
  assign n32090 = ~pi627 & ~n31962;
  assign n32091 = ~n32089 & n32090;
  assign n32092 = pi618 & ~n32085;
  assign n32093 = ~pi618 & n31890;
  assign n32094 = pi1154 & ~n32093;
  assign n32095 = ~n32092 & n32094;
  assign n32096 = pi627 & ~n31966;
  assign n32097 = ~n32095 & n32096;
  assign n32098 = ~n32091 & ~n32097;
  assign n32099 = pi781 & ~n32098;
  assign n32100 = ~pi781 & ~n32085;
  assign n32101 = ~n32099 & ~n32100;
  assign n32102 = ~pi619 & ~n32101;
  assign n32103 = pi619 & ~n31893;
  assign n32104 = ~pi1159 & ~n32103;
  assign n32105 = ~n32102 & n32104;
  assign n32106 = ~pi648 & ~n31974;
  assign n32107 = ~n32105 & n32106;
  assign n32108 = pi619 & ~n32101;
  assign n32109 = ~pi619 & ~n31893;
  assign n32110 = pi1159 & ~n32109;
  assign n32111 = ~n32108 & n32110;
  assign n32112 = pi648 & ~n31978;
  assign n32113 = ~n32111 & n32112;
  assign n32114 = pi789 & ~n32107;
  assign n32115 = ~n32113 & n32114;
  assign n32116 = ~pi789 & n32101;
  assign n32117 = n17905 & ~n32116;
  assign n32118 = ~n32115 & n32117;
  assign n32119 = ~pi626 & ~n31981;
  assign n32120 = pi626 & ~n31860;
  assign n32121 = n17668 & ~n32120;
  assign n32122 = ~n32119 & n32121;
  assign n32123 = pi626 & ~n31981;
  assign n32124 = ~pi626 & ~n31860;
  assign n32125 = n17667 & ~n32124;
  assign n32126 = ~n32123 & n32125;
  assign n32127 = n17792 & n31895;
  assign n32128 = ~n32122 & ~n32127;
  assign n32129 = ~n32126 & n32128;
  assign n32130 = pi788 & ~n32129;
  assign n32131 = ~n20298 & ~n32130;
  assign n32132 = ~n32118 & n32131;
  assign n32133 = ~n32016 & ~n32132;
  assign n32134 = n20300 & ~n32133;
  assign n32135 = n17737 & n31917;
  assign n32136 = n17738 & n31913;
  assign n32137 = ~n20491 & n31987;
  assign n32138 = ~n32135 & ~n32136;
  assign n32139 = ~n32137 & n32138;
  assign n32140 = pi787 & ~n32139;
  assign n32141 = ~n32134 & ~n32140;
  assign n32142 = ~n32010 & n32141;
  assign n32143 = ~n32006 & ~n32142;
  assign n32144 = ~po1038 & ~n32143;
  assign n32145 = ~pi192 & po1038;
  assign n32146 = ~pi832 & ~n32145;
  assign n32147 = ~n32144 & n32146;
  assign po349 = ~n31859 & ~n32147;
  assign n32149 = ~pi193 & ~n2755;
  assign n32150 = pi739 & n16933;
  assign n32151 = ~n32149 & ~n32150;
  assign n32152 = ~n17794 & ~n32151;
  assign n32153 = ~pi785 & ~n32152;
  assign n32154 = n17539 & n32150;
  assign n32155 = n32152 & ~n32154;
  assign n32156 = pi1155 & ~n32155;
  assign n32157 = ~pi1155 & ~n32149;
  assign n32158 = ~n32154 & n32157;
  assign n32159 = ~n32156 & ~n32158;
  assign n32160 = pi785 & ~n32159;
  assign n32161 = ~n32153 & ~n32160;
  assign n32162 = ~pi781 & ~n32161;
  assign n32163 = ~n17809 & n32161;
  assign n32164 = pi1154 & ~n32163;
  assign n32165 = ~n17812 & n32161;
  assign n32166 = ~pi1154 & ~n32165;
  assign n32167 = ~n32164 & ~n32166;
  assign n32168 = pi781 & ~n32167;
  assign n32169 = ~n32162 & ~n32168;
  assign n32170 = ~pi789 & ~n32169;
  assign n32171 = ~n22988 & n32169;
  assign n32172 = pi1159 & ~n32171;
  assign n32173 = ~n22991 & n32169;
  assign n32174 = ~pi1159 & ~n32173;
  assign n32175 = ~n32172 & ~n32174;
  assign n32176 = pi789 & ~n32175;
  assign n32177 = ~n32170 & ~n32176;
  assign n32178 = ~n17904 & n32177;
  assign n32179 = n17904 & n32149;
  assign n32180 = ~n32178 & ~n32179;
  assign n32181 = ~n17698 & ~n32180;
  assign n32182 = n17698 & n32149;
  assign n32183 = ~n32181 & ~n32182;
  assign n32184 = ~n20491 & n32183;
  assign n32185 = pi690 & n17153;
  assign n32186 = ~n32149 & ~n32185;
  assign n32187 = ~pi778 & ~n32186;
  assign n32188 = ~pi625 & n32185;
  assign n32189 = ~n32186 & ~n32188;
  assign n32190 = pi1153 & ~n32189;
  assign n32191 = ~pi1153 & ~n32149;
  assign n32192 = ~n32188 & n32191;
  assign n32193 = pi778 & ~n32192;
  assign n32194 = ~n32190 & n32193;
  assign n32195 = ~n32187 & ~n32194;
  assign n32196 = ~n17780 & ~n32195;
  assign n32197 = ~n17782 & n32196;
  assign n32198 = ~n17784 & n32197;
  assign n32199 = ~n17916 & n32198;
  assign n32200 = ~n17947 & n32199;
  assign n32201 = ~pi647 & n32200;
  assign n32202 = pi647 & n32149;
  assign n32203 = ~pi1157 & ~n32202;
  assign n32204 = ~n32201 & n32203;
  assign n32205 = pi647 & ~n32200;
  assign n32206 = ~pi647 & ~n32149;
  assign n32207 = ~n32205 & ~n32206;
  assign n32208 = pi1157 & ~n32207;
  assign n32209 = ~n32204 & ~n32208;
  assign n32210 = ~n17739 & ~n32209;
  assign n32211 = ~n32184 & ~n32210;
  assign n32212 = pi787 & ~n32211;
  assign n32213 = ~pi626 & ~n32177;
  assign n32214 = pi626 & ~n32149;
  assign n32215 = n17668 & ~n32214;
  assign n32216 = ~n32213 & n32215;
  assign n32217 = pi626 & ~n32177;
  assign n32218 = ~pi626 & ~n32149;
  assign n32219 = n17667 & ~n32218;
  assign n32220 = ~n32217 & n32219;
  assign n32221 = n17792 & n32198;
  assign n32222 = ~n32216 & ~n32221;
  assign n32223 = ~n32220 & n32222;
  assign n32224 = pi788 & ~n32223;
  assign n32225 = ~n16842 & ~n32186;
  assign n32226 = pi625 & n32225;
  assign n32227 = n32151 & ~n32225;
  assign n32228 = ~n32226 & ~n32227;
  assign n32229 = n32191 & ~n32228;
  assign n32230 = ~pi608 & ~n32190;
  assign n32231 = ~n32229 & n32230;
  assign n32232 = pi1153 & n32151;
  assign n32233 = ~n32226 & n32232;
  assign n32234 = pi608 & ~n32192;
  assign n32235 = ~n32233 & n32234;
  assign n32236 = ~n32231 & ~n32235;
  assign n32237 = pi778 & ~n32236;
  assign n32238 = ~pi778 & ~n32227;
  assign n32239 = ~n32237 & ~n32238;
  assign n32240 = ~pi609 & ~n32239;
  assign n32241 = pi609 & ~n32195;
  assign n32242 = ~pi1155 & ~n32241;
  assign n32243 = ~n32240 & n32242;
  assign n32244 = ~pi660 & ~n32156;
  assign n32245 = ~n32243 & n32244;
  assign n32246 = pi609 & ~n32239;
  assign n32247 = ~pi609 & ~n32195;
  assign n32248 = pi1155 & ~n32247;
  assign n32249 = ~n32246 & n32248;
  assign n32250 = pi660 & ~n32158;
  assign n32251 = ~n32249 & n32250;
  assign n32252 = ~n32245 & ~n32251;
  assign n32253 = pi785 & ~n32252;
  assign n32254 = ~pi785 & ~n32239;
  assign n32255 = ~n32253 & ~n32254;
  assign n32256 = ~pi618 & ~n32255;
  assign n32257 = pi618 & n32196;
  assign n32258 = ~pi1154 & ~n32257;
  assign n32259 = ~n32256 & n32258;
  assign n32260 = ~pi627 & ~n32164;
  assign n32261 = ~n32259 & n32260;
  assign n32262 = pi618 & ~n32255;
  assign n32263 = ~pi618 & n32196;
  assign n32264 = pi1154 & ~n32263;
  assign n32265 = ~n32262 & n32264;
  assign n32266 = pi627 & ~n32166;
  assign n32267 = ~n32265 & n32266;
  assign n32268 = ~n32261 & ~n32267;
  assign n32269 = pi781 & ~n32268;
  assign n32270 = ~pi781 & ~n32255;
  assign n32271 = ~n32269 & ~n32270;
  assign n32272 = ~pi619 & ~n32271;
  assign n32273 = pi619 & n32197;
  assign n32274 = ~pi1159 & ~n32273;
  assign n32275 = ~n32272 & n32274;
  assign n32276 = ~pi648 & ~n32172;
  assign n32277 = ~n32275 & n32276;
  assign n32278 = pi619 & ~n32271;
  assign n32279 = ~pi619 & n32197;
  assign n32280 = pi1159 & ~n32279;
  assign n32281 = ~n32278 & n32280;
  assign n32282 = pi648 & ~n32174;
  assign n32283 = ~n32281 & n32282;
  assign n32284 = pi789 & ~n32277;
  assign n32285 = ~n32283 & n32284;
  assign n32286 = ~pi789 & n32271;
  assign n32287 = n17905 & ~n32286;
  assign n32288 = ~n32285 & n32287;
  assign n32289 = ~n32224 & ~n32288;
  assign n32290 = ~n20298 & ~n32289;
  assign n32291 = n17944 & ~n32180;
  assign n32292 = n20786 & n32199;
  assign n32293 = ~n32291 & ~n32292;
  assign n32294 = ~pi629 & ~n32293;
  assign n32295 = n20790 & n32199;
  assign n32296 = n17943 & ~n32180;
  assign n32297 = ~n32295 & ~n32296;
  assign n32298 = pi629 & ~n32297;
  assign n32299 = ~n32294 & ~n32298;
  assign n32300 = pi792 & ~n32299;
  assign n32301 = n20300 & ~n32300;
  assign n32302 = ~n32290 & n32301;
  assign n32303 = ~n32212 & ~n32302;
  assign n32304 = pi644 & n32303;
  assign n32305 = ~pi787 & ~n32200;
  assign n32306 = pi787 & ~n32209;
  assign n32307 = ~n32305 & ~n32306;
  assign n32308 = ~pi644 & n32307;
  assign n32309 = pi715 & ~n32308;
  assign n32310 = ~n32304 & n32309;
  assign n32311 = ~n17740 & ~n32183;
  assign n32312 = n17740 & n32149;
  assign n32313 = ~n32311 & ~n32312;
  assign n32314 = pi644 & ~n32313;
  assign n32315 = ~pi644 & n32149;
  assign n32316 = ~pi715 & ~n32315;
  assign n32317 = ~n32314 & n32316;
  assign n32318 = pi1160 & ~n32317;
  assign n32319 = ~n32310 & n32318;
  assign n32320 = ~pi644 & n32303;
  assign n32321 = pi644 & n32307;
  assign n32322 = ~pi715 & ~n32321;
  assign n32323 = ~n32320 & n32322;
  assign n32324 = ~pi644 & ~n32313;
  assign n32325 = pi644 & n32149;
  assign n32326 = pi715 & ~n32325;
  assign n32327 = ~n32324 & n32326;
  assign n32328 = ~pi1160 & ~n32327;
  assign n32329 = ~n32323 & n32328;
  assign n32330 = ~n32319 & ~n32329;
  assign n32331 = pi790 & ~n32330;
  assign n32332 = ~pi790 & n32303;
  assign n32333 = pi832 & ~n32332;
  assign n32334 = ~n32331 & n32333;
  assign n32335 = ~pi193 & ~n17494;
  assign n32336 = n17627 & ~n32335;
  assign n32337 = pi690 & n3268;
  assign n32338 = n32335 & ~n32337;
  assign n32339 = pi193 & ~n18064;
  assign n32340 = ~pi38 & ~n32339;
  assign n32341 = n3268 & ~n32340;
  assign n32342 = ~pi193 & n18060;
  assign n32343 = ~n32341 & ~n32342;
  assign n32344 = ~pi193 & ~n16968;
  assign n32345 = n17480 & ~n32344;
  assign n32346 = pi690 & ~n32345;
  assign n32347 = ~n32343 & n32346;
  assign n32348 = ~n32338 & ~n32347;
  assign n32349 = ~pi778 & n32348;
  assign n32350 = pi625 & ~n32348;
  assign n32351 = ~pi625 & n32335;
  assign n32352 = pi1153 & ~n32351;
  assign n32353 = ~n32350 & n32352;
  assign n32354 = ~pi625 & ~n32348;
  assign n32355 = pi625 & n32335;
  assign n32356 = ~pi1153 & ~n32355;
  assign n32357 = ~n32354 & n32356;
  assign n32358 = ~n32353 & ~n32357;
  assign n32359 = pi778 & ~n32358;
  assign n32360 = ~n32349 & ~n32359;
  assign n32361 = ~n17554 & ~n32360;
  assign n32362 = n17554 & ~n32335;
  assign n32363 = ~n32361 & ~n32362;
  assign n32364 = ~n17591 & n32363;
  assign n32365 = n17591 & n32335;
  assign n32366 = ~n32364 & ~n32365;
  assign n32367 = ~n17627 & n32366;
  assign n32368 = ~n32336 & ~n32367;
  assign n32369 = ~n17670 & n32368;
  assign n32370 = n17670 & n32335;
  assign n32371 = ~n32369 & ~n32370;
  assign n32372 = ~pi792 & n32371;
  assign n32373 = pi628 & ~n32371;
  assign n32374 = ~pi628 & n32335;
  assign n32375 = pi1156 & ~n32374;
  assign n32376 = ~n32373 & n32375;
  assign n32377 = ~pi628 & ~n32371;
  assign n32378 = pi628 & n32335;
  assign n32379 = ~pi1156 & ~n32378;
  assign n32380 = ~n32377 & n32379;
  assign n32381 = ~n32376 & ~n32380;
  assign n32382 = pi792 & ~n32381;
  assign n32383 = ~n32372 & ~n32382;
  assign n32384 = ~pi647 & ~n32383;
  assign n32385 = pi647 & ~n32335;
  assign n32386 = ~n32384 & ~n32385;
  assign n32387 = ~pi1157 & n32386;
  assign n32388 = pi647 & ~n32383;
  assign n32389 = ~pi647 & ~n32335;
  assign n32390 = ~n32388 & ~n32389;
  assign n32391 = pi1157 & n32390;
  assign n32392 = ~n32387 & ~n32391;
  assign n32393 = pi787 & ~n32392;
  assign n32394 = ~pi787 & n32383;
  assign n32395 = ~n32393 & ~n32394;
  assign n32396 = ~pi644 & ~n32395;
  assign n32397 = pi715 & ~n32396;
  assign n32398 = pi193 & ~n3268;
  assign n32399 = pi739 & n16970;
  assign n32400 = ~n32344 & ~n32399;
  assign n32401 = pi38 & ~n32400;
  assign n32402 = ~pi193 & n16907;
  assign n32403 = pi193 & ~n16963;
  assign n32404 = pi739 & ~n32403;
  assign n32405 = ~n32402 & n32404;
  assign n32406 = ~pi193 & ~pi739;
  assign n32407 = ~n16816 & n32406;
  assign n32408 = ~n32405 & ~n32407;
  assign n32409 = ~pi38 & ~n32408;
  assign n32410 = ~n32401 & ~n32409;
  assign n32411 = n3268 & n32410;
  assign n32412 = ~n32398 & ~n32411;
  assign n32413 = ~n17526 & ~n32412;
  assign n32414 = n17526 & ~n32335;
  assign n32415 = ~n32413 & ~n32414;
  assign n32416 = ~pi785 & ~n32415;
  assign n32417 = ~n17527 & ~n32335;
  assign n32418 = pi609 & n32413;
  assign n32419 = ~n32417 & ~n32418;
  assign n32420 = pi1155 & ~n32419;
  assign n32421 = ~n17539 & ~n32335;
  assign n32422 = ~pi609 & n32413;
  assign n32423 = ~n32421 & ~n32422;
  assign n32424 = ~pi1155 & ~n32423;
  assign n32425 = ~n32420 & ~n32424;
  assign n32426 = pi785 & ~n32425;
  assign n32427 = ~n32416 & ~n32426;
  assign n32428 = ~pi781 & ~n32427;
  assign n32429 = pi618 & n32427;
  assign n32430 = ~pi618 & n32335;
  assign n32431 = pi1154 & ~n32430;
  assign n32432 = ~n32429 & n32431;
  assign n32433 = ~pi618 & n32427;
  assign n32434 = pi618 & n32335;
  assign n32435 = ~pi1154 & ~n32434;
  assign n32436 = ~n32433 & n32435;
  assign n32437 = ~n32432 & ~n32436;
  assign n32438 = pi781 & ~n32437;
  assign n32439 = ~n32428 & ~n32438;
  assign n32440 = ~pi789 & ~n32439;
  assign n32441 = pi619 & n32439;
  assign n32442 = ~pi619 & n32335;
  assign n32443 = pi1159 & ~n32442;
  assign n32444 = ~n32441 & n32443;
  assign n32445 = ~pi619 & n32439;
  assign n32446 = pi619 & n32335;
  assign n32447 = ~pi1159 & ~n32446;
  assign n32448 = ~n32445 & n32447;
  assign n32449 = ~n32444 & ~n32448;
  assign n32450 = pi789 & ~n32449;
  assign n32451 = ~n32440 & ~n32450;
  assign n32452 = ~n17904 & n32451;
  assign n32453 = n17904 & n32335;
  assign n32454 = ~n32452 & ~n32453;
  assign n32455 = ~n17698 & ~n32454;
  assign n32456 = n17698 & n32335;
  assign n32457 = ~n32455 & ~n32456;
  assign n32458 = ~n17740 & ~n32457;
  assign n32459 = n17740 & n32335;
  assign n32460 = ~n32458 & ~n32459;
  assign n32461 = pi644 & ~n32460;
  assign n32462 = ~pi644 & n32335;
  assign n32463 = ~pi715 & ~n32462;
  assign n32464 = ~n32461 & n32463;
  assign n32465 = pi1160 & ~n32464;
  assign n32466 = ~n32397 & n32465;
  assign n32467 = pi644 & ~n32395;
  assign n32468 = ~pi715 & ~n32467;
  assign n32469 = ~pi644 & ~n32460;
  assign n32470 = pi644 & n32335;
  assign n32471 = pi715 & ~n32470;
  assign n32472 = ~n32469 & n32471;
  assign n32473 = ~pi1160 & ~n32472;
  assign n32474 = ~n32468 & n32473;
  assign n32475 = ~n32466 & ~n32474;
  assign n32476 = pi790 & ~n32475;
  assign n32477 = ~pi644 & n32473;
  assign n32478 = pi644 & n32465;
  assign n32479 = pi790 & ~n32477;
  assign n32480 = ~n32478 & n32479;
  assign n32481 = ~n20502 & n32454;
  assign n32482 = ~pi629 & n32376;
  assign n32483 = pi629 & n32380;
  assign n32484 = ~n32482 & ~n32483;
  assign n32485 = ~n32481 & n32484;
  assign n32486 = pi792 & ~n32485;
  assign n32487 = ~pi690 & ~n32410;
  assign n32488 = ~pi193 & n17074;
  assign n32489 = pi193 & n17166;
  assign n32490 = ~pi739 & ~n32489;
  assign n32491 = ~n32488 & n32490;
  assign n32492 = pi193 & n17233;
  assign n32493 = ~pi193 & ~n17295;
  assign n32494 = pi739 & ~n32493;
  assign n32495 = ~n32492 & n32494;
  assign n32496 = pi39 & ~n32495;
  assign n32497 = ~n32491 & n32496;
  assign n32498 = ~pi193 & n17344;
  assign n32499 = pi193 & n17351;
  assign n32500 = pi739 & ~n32499;
  assign n32501 = ~n32498 & n32500;
  assign n32502 = pi193 & ~n17340;
  assign n32503 = ~pi193 & ~n17317;
  assign n32504 = ~pi739 & ~n32502;
  assign n32505 = ~n32503 & n32504;
  assign n32506 = ~n32501 & ~n32505;
  assign n32507 = ~pi39 & ~n32506;
  assign n32508 = ~pi38 & ~n32507;
  assign n32509 = ~n32497 & n32508;
  assign n32510 = ~pi739 & n24006;
  assign n32511 = ~n17259 & ~n32510;
  assign n32512 = ~pi39 & ~n32511;
  assign n32513 = ~pi193 & ~n32512;
  assign n32514 = ~n17154 & ~n32150;
  assign n32515 = pi193 & ~n32514;
  assign n32516 = n6250 & n32515;
  assign n32517 = pi38 & ~n32516;
  assign n32518 = ~n32513 & n32517;
  assign n32519 = pi690 & ~n32518;
  assign n32520 = ~n32509 & n32519;
  assign n32521 = n3268 & ~n32520;
  assign n32522 = ~n32487 & n32521;
  assign n32523 = ~n32398 & ~n32522;
  assign n32524 = ~pi625 & n32523;
  assign n32525 = pi625 & n32412;
  assign n32526 = ~pi1153 & ~n32525;
  assign n32527 = ~n32524 & n32526;
  assign n32528 = ~pi608 & ~n32353;
  assign n32529 = ~n32527 & n32528;
  assign n32530 = pi625 & n32523;
  assign n32531 = ~pi625 & n32412;
  assign n32532 = pi1153 & ~n32531;
  assign n32533 = ~n32530 & n32532;
  assign n32534 = pi608 & ~n32357;
  assign n32535 = ~n32533 & n32534;
  assign n32536 = ~n32529 & ~n32535;
  assign n32537 = pi778 & ~n32536;
  assign n32538 = ~pi778 & n32523;
  assign n32539 = ~n32537 & ~n32538;
  assign n32540 = ~pi609 & ~n32539;
  assign n32541 = pi609 & n32360;
  assign n32542 = ~pi1155 & ~n32541;
  assign n32543 = ~n32540 & n32542;
  assign n32544 = ~pi660 & ~n32420;
  assign n32545 = ~n32543 & n32544;
  assign n32546 = pi609 & ~n32539;
  assign n32547 = ~pi609 & n32360;
  assign n32548 = pi1155 & ~n32547;
  assign n32549 = ~n32546 & n32548;
  assign n32550 = pi660 & ~n32424;
  assign n32551 = ~n32549 & n32550;
  assign n32552 = ~n32545 & ~n32551;
  assign n32553 = pi785 & ~n32552;
  assign n32554 = ~pi785 & ~n32539;
  assign n32555 = ~n32553 & ~n32554;
  assign n32556 = ~pi618 & ~n32555;
  assign n32557 = pi618 & n32363;
  assign n32558 = ~pi1154 & ~n32557;
  assign n32559 = ~n32556 & n32558;
  assign n32560 = ~pi627 & ~n32432;
  assign n32561 = ~n32559 & n32560;
  assign n32562 = pi618 & ~n32555;
  assign n32563 = ~pi618 & n32363;
  assign n32564 = pi1154 & ~n32563;
  assign n32565 = ~n32562 & n32564;
  assign n32566 = pi627 & ~n32436;
  assign n32567 = ~n32565 & n32566;
  assign n32568 = ~n32561 & ~n32567;
  assign n32569 = pi781 & ~n32568;
  assign n32570 = ~pi781 & ~n32555;
  assign n32571 = ~n32569 & ~n32570;
  assign n32572 = ~pi619 & ~n32571;
  assign n32573 = pi619 & ~n32366;
  assign n32574 = ~pi1159 & ~n32573;
  assign n32575 = ~n32572 & n32574;
  assign n32576 = ~pi648 & ~n32444;
  assign n32577 = ~n32575 & n32576;
  assign n32578 = pi619 & ~n32571;
  assign n32579 = ~pi619 & ~n32366;
  assign n32580 = pi1159 & ~n32579;
  assign n32581 = ~n32578 & n32580;
  assign n32582 = pi648 & ~n32448;
  assign n32583 = ~n32581 & n32582;
  assign n32584 = pi789 & ~n32577;
  assign n32585 = ~n32583 & n32584;
  assign n32586 = ~pi789 & n32571;
  assign n32587 = n17905 & ~n32586;
  assign n32588 = ~n32585 & n32587;
  assign n32589 = ~pi626 & ~n32451;
  assign n32590 = pi626 & ~n32335;
  assign n32591 = n17668 & ~n32590;
  assign n32592 = ~n32589 & n32591;
  assign n32593 = pi626 & ~n32451;
  assign n32594 = ~pi626 & ~n32335;
  assign n32595 = n17667 & ~n32594;
  assign n32596 = ~n32593 & n32595;
  assign n32597 = n17792 & n32368;
  assign n32598 = ~n32592 & ~n32597;
  assign n32599 = ~n32596 & n32598;
  assign n32600 = pi788 & ~n32599;
  assign n32601 = ~n20298 & ~n32600;
  assign n32602 = ~n32588 & n32601;
  assign n32603 = ~n32486 & ~n32602;
  assign n32604 = n20300 & ~n32603;
  assign n32605 = ~n20491 & n32457;
  assign n32606 = n17738 & ~n32386;
  assign n32607 = n17737 & ~n32390;
  assign n32608 = ~n32606 & ~n32607;
  assign n32609 = ~n32605 & n32608;
  assign n32610 = pi787 & ~n32609;
  assign n32611 = ~n32604 & ~n32610;
  assign n32612 = ~n32480 & n32611;
  assign n32613 = ~n32476 & ~n32612;
  assign n32614 = ~po1038 & ~n32613;
  assign n32615 = ~pi193 & po1038;
  assign n32616 = ~pi832 & ~n32615;
  assign n32617 = ~n32614 & n32616;
  assign po350 = ~n32334 & ~n32617;
  assign n32619 = pi194 & ~n3268;
  assign n32620 = ~pi194 & n19349;
  assign n32621 = pi194 & n24371;
  assign n32622 = ~n32620 & ~n32621;
  assign n32623 = pi748 & ~n32622;
  assign n32624 = ~pi194 & ~n17487;
  assign n32625 = ~pi748 & ~n32624;
  assign n32626 = ~n32623 & ~n32625;
  assign n32627 = ~pi730 & n32626;
  assign n32628 = ~pi194 & n19309;
  assign n32629 = pi194 & ~n24462;
  assign n32630 = ~pi748 & ~n32629;
  assign n32631 = ~n32628 & n32630;
  assign n32632 = pi194 & n19326;
  assign n32633 = ~pi194 & ~n19334;
  assign n32634 = pi748 & ~n32633;
  assign n32635 = ~n32632 & n32634;
  assign n32636 = pi730 & ~n32635;
  assign n32637 = ~n32631 & n32636;
  assign n32638 = n3268 & ~n32627;
  assign n32639 = ~n32637 & n32638;
  assign n32640 = ~n32619 & ~n32639;
  assign n32641 = ~pi625 & n32640;
  assign n32642 = n3268 & ~n32626;
  assign n32643 = ~n32619 & ~n32642;
  assign n32644 = pi625 & n32643;
  assign n32645 = ~pi1153 & ~n32644;
  assign n32646 = ~n32641 & n32645;
  assign n32647 = pi194 & ~n24309;
  assign n32648 = ~pi194 & n24312;
  assign n32649 = pi730 & ~n32648;
  assign n32650 = ~pi730 & n32624;
  assign n32651 = n3268 & ~n32650;
  assign n32652 = ~n32649 & n32651;
  assign n32653 = ~n32647 & ~n32652;
  assign n32654 = pi625 & n32653;
  assign n32655 = ~pi194 & ~n17494;
  assign n32656 = ~pi625 & n32655;
  assign n32657 = pi1153 & ~n32656;
  assign n32658 = ~n32654 & n32657;
  assign n32659 = ~pi608 & ~n32658;
  assign n32660 = ~n32646 & n32659;
  assign n32661 = pi625 & n32640;
  assign n32662 = ~pi625 & n32643;
  assign n32663 = pi1153 & ~n32662;
  assign n32664 = ~n32661 & n32663;
  assign n32665 = ~pi625 & n32653;
  assign n32666 = pi625 & n32655;
  assign n32667 = ~pi1153 & ~n32666;
  assign n32668 = ~n32665 & n32667;
  assign n32669 = pi608 & ~n32668;
  assign n32670 = ~n32664 & n32669;
  assign n32671 = ~n32660 & ~n32670;
  assign n32672 = pi778 & ~n32671;
  assign n32673 = ~pi778 & n32640;
  assign n32674 = ~n32672 & ~n32673;
  assign n32675 = ~pi609 & ~n32674;
  assign n32676 = ~pi778 & ~n32653;
  assign n32677 = ~n32658 & ~n32668;
  assign n32678 = pi778 & ~n32677;
  assign n32679 = ~n32676 & ~n32678;
  assign n32680 = pi609 & n32679;
  assign n32681 = ~pi1155 & ~n32680;
  assign n32682 = ~n32675 & n32681;
  assign n32683 = ~n17527 & ~n32655;
  assign n32684 = ~n17526 & ~n32643;
  assign n32685 = pi609 & n32684;
  assign n32686 = ~n32683 & ~n32685;
  assign n32687 = pi1155 & ~n32686;
  assign n32688 = ~pi660 & ~n32687;
  assign n32689 = ~n32682 & n32688;
  assign n32690 = pi609 & ~n32674;
  assign n32691 = ~pi609 & n32679;
  assign n32692 = pi1155 & ~n32691;
  assign n32693 = ~n32690 & n32692;
  assign n32694 = ~n17539 & ~n32655;
  assign n32695 = ~pi609 & n32684;
  assign n32696 = ~n32694 & ~n32695;
  assign n32697 = ~pi1155 & ~n32696;
  assign n32698 = pi660 & ~n32697;
  assign n32699 = ~n32693 & n32698;
  assign n32700 = ~n32689 & ~n32699;
  assign n32701 = pi785 & ~n32700;
  assign n32702 = ~pi785 & ~n32674;
  assign n32703 = ~n32701 & ~n32702;
  assign n32704 = ~pi618 & ~n32703;
  assign n32705 = ~n17554 & ~n32679;
  assign n32706 = n17554 & ~n32655;
  assign n32707 = ~n32705 & ~n32706;
  assign n32708 = pi618 & n32707;
  assign n32709 = ~pi1154 & ~n32708;
  assign n32710 = ~n32704 & n32709;
  assign n32711 = n17526 & ~n32655;
  assign n32712 = ~n32684 & ~n32711;
  assign n32713 = ~pi785 & ~n32712;
  assign n32714 = ~n32687 & ~n32697;
  assign n32715 = pi785 & ~n32714;
  assign n32716 = ~n32713 & ~n32715;
  assign n32717 = pi618 & n32716;
  assign n32718 = ~pi618 & n32655;
  assign n32719 = pi1154 & ~n32718;
  assign n32720 = ~n32717 & n32719;
  assign n32721 = ~pi627 & ~n32720;
  assign n32722 = ~n32710 & n32721;
  assign n32723 = pi618 & ~n32703;
  assign n32724 = ~pi618 & n32707;
  assign n32725 = pi1154 & ~n32724;
  assign n32726 = ~n32723 & n32725;
  assign n32727 = ~pi618 & n32716;
  assign n32728 = pi618 & n32655;
  assign n32729 = ~pi1154 & ~n32728;
  assign n32730 = ~n32727 & n32729;
  assign n32731 = pi627 & ~n32730;
  assign n32732 = ~n32726 & n32731;
  assign n32733 = ~n32722 & ~n32732;
  assign n32734 = pi781 & ~n32733;
  assign n32735 = ~pi781 & ~n32703;
  assign n32736 = ~n32734 & ~n32735;
  assign n32737 = ~pi619 & ~n32736;
  assign n32738 = ~n17591 & n32707;
  assign n32739 = n17591 & n32655;
  assign n32740 = ~n32738 & ~n32739;
  assign n32741 = pi619 & ~n32740;
  assign n32742 = ~pi1159 & ~n32741;
  assign n32743 = ~n32737 & n32742;
  assign n32744 = ~pi781 & ~n32716;
  assign n32745 = ~n32720 & ~n32730;
  assign n32746 = pi781 & ~n32745;
  assign n32747 = ~n32744 & ~n32746;
  assign n32748 = pi619 & n32747;
  assign n32749 = ~pi619 & n32655;
  assign n32750 = pi1159 & ~n32749;
  assign n32751 = ~n32748 & n32750;
  assign n32752 = ~pi648 & ~n32751;
  assign n32753 = ~n32743 & n32752;
  assign n32754 = pi619 & ~n32736;
  assign n32755 = ~pi619 & ~n32740;
  assign n32756 = pi1159 & ~n32755;
  assign n32757 = ~n32754 & n32756;
  assign n32758 = ~pi619 & n32747;
  assign n32759 = pi619 & n32655;
  assign n32760 = ~pi1159 & ~n32759;
  assign n32761 = ~n32758 & n32760;
  assign n32762 = pi648 & ~n32761;
  assign n32763 = ~n32757 & n32762;
  assign n32764 = ~n32753 & ~n32763;
  assign n32765 = pi789 & ~n32764;
  assign n32766 = ~pi789 & ~n32736;
  assign n32767 = ~n32765 & ~n32766;
  assign n32768 = ~pi788 & n32767;
  assign n32769 = ~pi626 & n32767;
  assign n32770 = n17627 & ~n32655;
  assign n32771 = ~n17627 & n32740;
  assign n32772 = ~n32770 & ~n32771;
  assign n32773 = pi626 & ~n32772;
  assign n32774 = ~pi641 & ~n32773;
  assign n32775 = ~n32769 & n32774;
  assign n32776 = ~pi789 & ~n32747;
  assign n32777 = ~n32751 & ~n32761;
  assign n32778 = pi789 & ~n32777;
  assign n32779 = ~n32776 & ~n32778;
  assign n32780 = ~pi626 & ~n32779;
  assign n32781 = pi626 & ~n32655;
  assign n32782 = pi641 & ~n32781;
  assign n32783 = ~n32780 & n32782;
  assign n32784 = ~pi1158 & ~n32783;
  assign n32785 = ~n32775 & n32784;
  assign n32786 = pi626 & n32767;
  assign n32787 = ~pi626 & ~n32772;
  assign n32788 = pi641 & ~n32787;
  assign n32789 = ~n32786 & n32788;
  assign n32790 = pi626 & ~n32779;
  assign n32791 = ~pi626 & ~n32655;
  assign n32792 = ~pi641 & ~n32791;
  assign n32793 = ~n32790 & n32792;
  assign n32794 = pi1158 & ~n32793;
  assign n32795 = ~n32789 & n32794;
  assign n32796 = ~n32785 & ~n32795;
  assign n32797 = pi788 & ~n32796;
  assign n32798 = ~n32768 & ~n32797;
  assign n32799 = ~pi628 & n32798;
  assign n32800 = ~n17904 & n32779;
  assign n32801 = n17904 & n32655;
  assign n32802 = ~n32800 & ~n32801;
  assign n32803 = pi628 & ~n32802;
  assign n32804 = ~pi1156 & ~n32803;
  assign n32805 = ~n32799 & n32804;
  assign n32806 = ~n17670 & n32772;
  assign n32807 = n17670 & n32655;
  assign n32808 = ~n32806 & ~n32807;
  assign n32809 = pi628 & ~n32808;
  assign n32810 = ~pi628 & n32655;
  assign n32811 = pi1156 & ~n32810;
  assign n32812 = ~n32809 & n32811;
  assign n32813 = ~pi629 & ~n32812;
  assign n32814 = ~n32805 & n32813;
  assign n32815 = pi628 & n32798;
  assign n32816 = ~pi628 & ~n32802;
  assign n32817 = pi1156 & ~n32816;
  assign n32818 = ~n32815 & n32817;
  assign n32819 = ~pi628 & ~n32808;
  assign n32820 = pi628 & n32655;
  assign n32821 = ~pi1156 & ~n32820;
  assign n32822 = ~n32819 & n32821;
  assign n32823 = pi629 & ~n32822;
  assign n32824 = ~n32818 & n32823;
  assign n32825 = ~n32814 & ~n32824;
  assign n32826 = pi792 & ~n32825;
  assign n32827 = ~pi792 & n32798;
  assign n32828 = ~n32826 & ~n32827;
  assign n32829 = ~pi647 & ~n32828;
  assign n32830 = ~n17698 & ~n32802;
  assign n32831 = n17698 & n32655;
  assign n32832 = ~n32830 & ~n32831;
  assign n32833 = pi647 & ~n32832;
  assign n32834 = ~pi1157 & ~n32833;
  assign n32835 = ~n32829 & n32834;
  assign n32836 = ~pi792 & n32808;
  assign n32837 = ~n32812 & ~n32822;
  assign n32838 = pi792 & ~n32837;
  assign n32839 = ~n32836 & ~n32838;
  assign n32840 = pi647 & n32839;
  assign n32841 = ~pi647 & n32655;
  assign n32842 = pi1157 & ~n32841;
  assign n32843 = ~n32840 & n32842;
  assign n32844 = ~pi630 & ~n32843;
  assign n32845 = ~n32835 & n32844;
  assign n32846 = pi647 & ~n32828;
  assign n32847 = ~pi647 & ~n32832;
  assign n32848 = pi1157 & ~n32847;
  assign n32849 = ~n32846 & n32848;
  assign n32850 = ~pi647 & n32839;
  assign n32851 = pi647 & n32655;
  assign n32852 = ~pi1157 & ~n32851;
  assign n32853 = ~n32850 & n32852;
  assign n32854 = pi630 & ~n32853;
  assign n32855 = ~n32849 & n32854;
  assign n32856 = ~n32845 & ~n32855;
  assign n32857 = pi787 & ~n32856;
  assign n32858 = ~pi787 & ~n32828;
  assign n32859 = ~n32857 & ~n32858;
  assign n32860 = pi644 & ~n32859;
  assign n32861 = ~pi787 & ~n32839;
  assign n32862 = ~n32843 & ~n32853;
  assign n32863 = pi787 & ~n32862;
  assign n32864 = ~n32861 & ~n32863;
  assign n32865 = ~pi644 & n32864;
  assign n32866 = pi715 & ~n32865;
  assign n32867 = ~n32860 & n32866;
  assign n32868 = n17740 & ~n32655;
  assign n32869 = ~n17740 & n32832;
  assign n32870 = ~n32868 & ~n32869;
  assign n32871 = pi644 & n32870;
  assign n32872 = ~pi644 & n32655;
  assign n32873 = ~pi715 & ~n32872;
  assign n32874 = ~n32871 & n32873;
  assign n32875 = pi1160 & ~n32874;
  assign n32876 = ~n32867 & n32875;
  assign n32877 = ~pi644 & ~n32859;
  assign n32878 = pi644 & n32864;
  assign n32879 = ~pi715 & ~n32878;
  assign n32880 = ~n32877 & n32879;
  assign n32881 = ~pi644 & n32870;
  assign n32882 = pi644 & n32655;
  assign n32883 = pi715 & ~n32882;
  assign n32884 = ~n32881 & n32883;
  assign n32885 = ~pi1160 & ~n32884;
  assign n32886 = ~n32880 & n32885;
  assign n32887 = pi790 & ~n32876;
  assign n32888 = ~n32886 & n32887;
  assign n32889 = ~pi790 & n32859;
  assign n32890 = ~po1038 & ~n32889;
  assign n32891 = ~n32888 & n32890;
  assign n32892 = ~pi194 & po1038;
  assign n32893 = ~pi832 & ~n32892;
  assign n32894 = ~n32891 & n32893;
  assign n32895 = ~pi194 & ~n2755;
  assign n32896 = pi748 & n16933;
  assign n32897 = ~n32895 & ~n32896;
  assign n32898 = ~n17794 & ~n32897;
  assign n32899 = ~pi785 & ~n32898;
  assign n32900 = ~n17799 & ~n32897;
  assign n32901 = pi1155 & ~n32900;
  assign n32902 = ~n17802 & n32898;
  assign n32903 = ~pi1155 & ~n32902;
  assign n32904 = ~n32901 & ~n32903;
  assign n32905 = pi785 & ~n32904;
  assign n32906 = ~n32899 & ~n32905;
  assign n32907 = ~pi781 & ~n32906;
  assign n32908 = ~n17809 & n32906;
  assign n32909 = pi1154 & ~n32908;
  assign n32910 = ~n17812 & n32906;
  assign n32911 = ~pi1154 & ~n32910;
  assign n32912 = ~n32909 & ~n32911;
  assign n32913 = pi781 & ~n32912;
  assign n32914 = ~n32907 & ~n32913;
  assign n32915 = ~pi789 & ~n32914;
  assign n32916 = pi619 & n32914;
  assign n32917 = ~pi619 & n32895;
  assign n32918 = pi1159 & ~n32917;
  assign n32919 = ~n32916 & n32918;
  assign n32920 = ~pi619 & n32914;
  assign n32921 = pi619 & n32895;
  assign n32922 = ~pi1159 & ~n32921;
  assign n32923 = ~n32920 & n32922;
  assign n32924 = ~n32919 & ~n32923;
  assign n32925 = pi789 & ~n32924;
  assign n32926 = ~n32915 & ~n32925;
  assign n32927 = ~n17904 & n32926;
  assign n32928 = n17904 & n32895;
  assign n32929 = ~n32927 & ~n32928;
  assign n32930 = ~n17698 & ~n32929;
  assign n32931 = n17698 & n32895;
  assign n32932 = ~n32930 & ~n32931;
  assign n32933 = ~n20491 & n32932;
  assign n32934 = pi730 & n17153;
  assign n32935 = ~n32895 & ~n32934;
  assign n32936 = ~pi778 & n32935;
  assign n32937 = ~pi625 & n32934;
  assign n32938 = ~n32935 & ~n32937;
  assign n32939 = pi1153 & ~n32938;
  assign n32940 = ~pi1153 & ~n32895;
  assign n32941 = ~n32937 & n32940;
  assign n32942 = ~n32939 & ~n32941;
  assign n32943 = pi778 & ~n32942;
  assign n32944 = ~n32936 & ~n32943;
  assign n32945 = ~n17780 & n32944;
  assign n32946 = ~n17782 & n32945;
  assign n32947 = ~n17784 & n32946;
  assign n32948 = ~n17916 & n32947;
  assign n32949 = ~n17947 & n32948;
  assign n32950 = ~pi647 & n32949;
  assign n32951 = pi647 & n32895;
  assign n32952 = ~pi1157 & ~n32951;
  assign n32953 = ~n32950 & n32952;
  assign n32954 = pi647 & ~n32949;
  assign n32955 = ~pi647 & ~n32895;
  assign n32956 = ~n32954 & ~n32955;
  assign n32957 = pi1157 & ~n32956;
  assign n32958 = ~n32953 & ~n32957;
  assign n32959 = ~n17739 & ~n32958;
  assign n32960 = ~n32933 & ~n32959;
  assign n32961 = pi787 & ~n32960;
  assign n32962 = ~pi626 & ~n32926;
  assign n32963 = pi626 & ~n32895;
  assign n32964 = n17668 & ~n32963;
  assign n32965 = ~n32962 & n32964;
  assign n32966 = pi626 & ~n32926;
  assign n32967 = ~pi626 & ~n32895;
  assign n32968 = n17667 & ~n32967;
  assign n32969 = ~n32966 & n32968;
  assign n32970 = n17792 & n32947;
  assign n32971 = ~n32965 & ~n32970;
  assign n32972 = ~n32969 & n32971;
  assign n32973 = pi788 & ~n32972;
  assign n32974 = ~n16842 & ~n32935;
  assign n32975 = pi625 & n32974;
  assign n32976 = n32897 & ~n32974;
  assign n32977 = ~n32975 & ~n32976;
  assign n32978 = n32940 & ~n32977;
  assign n32979 = ~pi608 & ~n32939;
  assign n32980 = ~n32978 & n32979;
  assign n32981 = pi1153 & n32897;
  assign n32982 = ~n32975 & n32981;
  assign n32983 = pi608 & ~n32941;
  assign n32984 = ~n32982 & n32983;
  assign n32985 = ~n32980 & ~n32984;
  assign n32986 = pi778 & ~n32985;
  assign n32987 = ~pi778 & ~n32976;
  assign n32988 = ~n32986 & ~n32987;
  assign n32989 = ~pi609 & ~n32988;
  assign n32990 = pi609 & n32944;
  assign n32991 = ~pi1155 & ~n32990;
  assign n32992 = ~n32989 & n32991;
  assign n32993 = ~pi660 & ~n32901;
  assign n32994 = ~n32992 & n32993;
  assign n32995 = pi609 & ~n32988;
  assign n32996 = ~pi609 & n32944;
  assign n32997 = pi1155 & ~n32996;
  assign n32998 = ~n32995 & n32997;
  assign n32999 = pi660 & ~n32903;
  assign n33000 = ~n32998 & n32999;
  assign n33001 = ~n32994 & ~n33000;
  assign n33002 = pi785 & ~n33001;
  assign n33003 = ~pi785 & ~n32988;
  assign n33004 = ~n33002 & ~n33003;
  assign n33005 = ~pi618 & ~n33004;
  assign n33006 = pi618 & n32945;
  assign n33007 = ~pi1154 & ~n33006;
  assign n33008 = ~n33005 & n33007;
  assign n33009 = ~pi627 & ~n32909;
  assign n33010 = ~n33008 & n33009;
  assign n33011 = pi618 & ~n33004;
  assign n33012 = ~pi618 & n32945;
  assign n33013 = pi1154 & ~n33012;
  assign n33014 = ~n33011 & n33013;
  assign n33015 = pi627 & ~n32911;
  assign n33016 = ~n33014 & n33015;
  assign n33017 = ~n33010 & ~n33016;
  assign n33018 = pi781 & ~n33017;
  assign n33019 = ~pi781 & ~n33004;
  assign n33020 = ~n33018 & ~n33019;
  assign n33021 = ~pi619 & ~n33020;
  assign n33022 = pi619 & n32946;
  assign n33023 = ~pi1159 & ~n33022;
  assign n33024 = ~n33021 & n33023;
  assign n33025 = ~pi648 & ~n32919;
  assign n33026 = ~n33024 & n33025;
  assign n33027 = pi619 & ~n33020;
  assign n33028 = ~pi619 & n32946;
  assign n33029 = pi1159 & ~n33028;
  assign n33030 = ~n33027 & n33029;
  assign n33031 = pi648 & ~n32923;
  assign n33032 = ~n33030 & n33031;
  assign n33033 = pi789 & ~n33026;
  assign n33034 = ~n33032 & n33033;
  assign n33035 = ~pi789 & n33020;
  assign n33036 = n17905 & ~n33035;
  assign n33037 = ~n33034 & n33036;
  assign n33038 = ~n32973 & ~n33037;
  assign n33039 = ~n20298 & ~n33038;
  assign n33040 = n17944 & ~n32929;
  assign n33041 = n20786 & n32948;
  assign n33042 = ~n33040 & ~n33041;
  assign n33043 = ~pi629 & ~n33042;
  assign n33044 = n20790 & n32948;
  assign n33045 = n17943 & ~n32929;
  assign n33046 = ~n33044 & ~n33045;
  assign n33047 = pi629 & ~n33046;
  assign n33048 = ~n33043 & ~n33047;
  assign n33049 = pi792 & ~n33048;
  assign n33050 = n20300 & ~n33049;
  assign n33051 = ~n33039 & n33050;
  assign n33052 = ~n32961 & ~n33051;
  assign n33053 = pi644 & n33052;
  assign n33054 = ~pi787 & ~n32949;
  assign n33055 = pi787 & ~n32958;
  assign n33056 = ~n33054 & ~n33055;
  assign n33057 = ~pi644 & n33056;
  assign n33058 = pi715 & ~n33057;
  assign n33059 = ~n33053 & n33058;
  assign n33060 = ~n17740 & ~n32932;
  assign n33061 = n17740 & n32895;
  assign n33062 = ~n33060 & ~n33061;
  assign n33063 = pi644 & ~n33062;
  assign n33064 = ~pi644 & n32895;
  assign n33065 = ~pi715 & ~n33064;
  assign n33066 = ~n33063 & n33065;
  assign n33067 = pi1160 & ~n33066;
  assign n33068 = ~n33059 & n33067;
  assign n33069 = ~pi644 & n33052;
  assign n33070 = pi644 & n33056;
  assign n33071 = ~pi715 & ~n33070;
  assign n33072 = ~n33069 & n33071;
  assign n33073 = ~pi644 & ~n33062;
  assign n33074 = pi644 & n32895;
  assign n33075 = pi715 & ~n33074;
  assign n33076 = ~n33073 & n33075;
  assign n33077 = ~pi1160 & ~n33076;
  assign n33078 = ~n33072 & n33077;
  assign n33079 = ~n33068 & ~n33078;
  assign n33080 = pi790 & ~n33079;
  assign n33081 = ~pi790 & n33052;
  assign n33082 = pi832 & ~n33081;
  assign n33083 = ~n33080 & n33082;
  assign po351 = ~n32894 & ~n33083;
  assign n33085 = ~n6206 & n16144;
  assign n33086 = ~n11448 & n16121;
  assign n33087 = n16118 & ~n16501;
  assign n33088 = ~n11451 & ~n33085;
  assign n33089 = ~n33086 & ~n33087;
  assign n33090 = n33088 & n33089;
  assign n33091 = pi232 & ~n33090;
  assign n33092 = ~n16498 & ~n33091;
  assign n33093 = pi39 & ~n33092;
  assign n33094 = n13862 & ~n16146;
  assign n33095 = ~pi39 & ~n33094;
  assign n33096 = ~pi138 & n16515;
  assign n33097 = ~pi196 & n33096;
  assign n33098 = pi195 & ~n33097;
  assign n33099 = n10181 & ~n33098;
  assign n33100 = ~n33095 & n33099;
  assign n33101 = ~n33093 & n33100;
  assign n33102 = pi192 & n16450;
  assign n33103 = ~n9384 & ~n16112;
  assign n33104 = pi171 & n13683;
  assign n33105 = ~n33103 & ~n33104;
  assign n33106 = pi299 & ~n33105;
  assign n33107 = ~pi192 & n16444;
  assign n33108 = pi232 & ~n33107;
  assign n33109 = ~n33102 & n33108;
  assign n33110 = ~n33106 & n33109;
  assign n33111 = n16447 & ~n33110;
  assign n33112 = ~pi171 & n9064;
  assign n33113 = ~n16471 & ~n33112;
  assign n33114 = n9055 & ~n33113;
  assign n33115 = n9057 & ~n33114;
  assign n33116 = pi192 & n16478;
  assign n33117 = ~pi192 & n16464;
  assign n33118 = ~n33115 & ~n33117;
  assign n33119 = ~n33116 & n33118;
  assign n33120 = pi232 & ~n33119;
  assign n33121 = ~n16470 & ~n33120;
  assign n33122 = pi39 & ~n33121;
  assign n33123 = n3207 & ~n33122;
  assign n33124 = ~n33111 & n33123;
  assign n33125 = ~pi87 & ~n33124;
  assign n33126 = n16442 & ~n33125;
  assign n33127 = ~pi92 & ~n33126;
  assign n33128 = n16441 & ~n33127;
  assign n33129 = ~pi55 & ~n33128;
  assign n33130 = ~n16493 & ~n33129;
  assign n33131 = n3294 & ~n33130;
  assign n33132 = n9707 & n33098;
  assign n33133 = ~n33131 & n33132;
  assign po352 = n33101 | n33133;
  assign n33135 = ~pi170 & n9064;
  assign n33136 = ~n16471 & ~n33135;
  assign n33137 = n9055 & ~n33136;
  assign n33138 = n9057 & ~n33137;
  assign n33139 = ~n16464 & ~n33138;
  assign n33140 = pi232 & ~n33139;
  assign n33141 = ~n16470 & ~n33140;
  assign n33142 = pi232 & n16478;
  assign n33143 = n33141 & ~n33142;
  assign n33144 = pi39 & ~n33143;
  assign n33145 = ~pi38 & pi194;
  assign n33146 = ~n33144 & n33145;
  assign n33147 = pi39 & ~n33141;
  assign n33148 = ~pi38 & ~pi194;
  assign n33149 = ~n33147 & n33148;
  assign n33150 = ~n33146 & ~n33149;
  assign n33151 = ~n16447 & ~n33150;
  assign n33152 = ~n16450 & n33146;
  assign n33153 = ~n16444 & n33149;
  assign n33154 = ~n33152 & ~n33153;
  assign n33155 = ~n9384 & ~n16221;
  assign n33156 = pi170 & n13683;
  assign n33157 = ~n33155 & ~n33156;
  assign n33158 = pi299 & ~n33157;
  assign n33159 = pi232 & ~n33158;
  assign n33160 = ~n33154 & n33159;
  assign n33161 = ~n33151 & ~n33160;
  assign n33162 = ~pi100 & ~n33161;
  assign n33163 = ~pi87 & ~n33162;
  assign n33164 = n16442 & ~n33163;
  assign n33165 = ~pi92 & ~n33164;
  assign n33166 = n16441 & ~n33165;
  assign n33167 = ~pi55 & ~n33166;
  assign n33168 = ~n16493 & ~n33167;
  assign n33169 = n3294 & ~n33168;
  assign n33170 = n9707 & ~n33169;
  assign n33171 = pi196 & ~n33170;
  assign n33172 = ~pi170 & n9514;
  assign n33173 = ~n16500 & ~n33172;
  assign n33174 = n13094 & ~n33173;
  assign n33175 = n13096 & n16500;
  assign n33176 = pi232 & ~n33175;
  assign n33177 = ~n33174 & n33176;
  assign n33178 = ~n16498 & ~n33177;
  assign n33179 = pi299 & ~n33178;
  assign n33180 = ~n11449 & ~n33179;
  assign n33181 = pi39 & ~n33180;
  assign n33182 = n13862 & ~n16222;
  assign n33183 = ~pi39 & ~n33182;
  assign n33184 = ~pi38 & ~n33183;
  assign n33185 = ~n33181 & n33184;
  assign n33186 = ~pi194 & ~n33185;
  assign n33187 = pi39 & ~n33178;
  assign n33188 = n13862 & n16281;
  assign n33189 = ~pi39 & ~n33188;
  assign n33190 = ~pi38 & ~n33189;
  assign n33191 = ~n33187 & n33190;
  assign n33192 = pi194 & ~n33191;
  assign n33193 = n10178 & ~n33192;
  assign n33194 = ~n33186 & n33193;
  assign n33195 = ~pi196 & ~n33194;
  assign n33196 = ~n33096 & ~n33195;
  assign n33197 = ~n33171 & n33196;
  assign n33198 = pi195 & ~pi196;
  assign n33199 = ~n33170 & n33198;
  assign n33200 = ~n33194 & ~n33198;
  assign n33201 = n33096 & ~n33200;
  assign n33202 = ~n33199 & n33201;
  assign po353 = n33197 | n33202;
  assign n33204 = ~pi767 & pi947;
  assign n33205 = ~pi698 & n20848;
  assign n33206 = ~n33204 & ~n33205;
  assign n33207 = n2755 & ~n33206;
  assign n33208 = ~pi197 & ~n2755;
  assign n33209 = pi832 & ~n33208;
  assign n33210 = ~n33207 & n33209;
  assign n33211 = pi197 & ~n17485;
  assign n33212 = n16968 & ~n33204;
  assign n33213 = pi38 & ~n33212;
  assign n33214 = ~n33211 & n33213;
  assign n33215 = ~pi197 & ~n20933;
  assign n33216 = pi197 & ~n21087;
  assign n33217 = pi299 & ~n33216;
  assign n33218 = ~n33215 & n33217;
  assign n33219 = ~pi197 & ~n16792;
  assign n33220 = n20951 & ~n33219;
  assign n33221 = ~pi767 & ~n33220;
  assign n33222 = ~n33218 & n33221;
  assign n33223 = ~pi197 & pi767;
  assign n33224 = ~n16814 & n33223;
  assign n33225 = pi39 & ~n33224;
  assign n33226 = ~n33222 & n33225;
  assign n33227 = ~pi197 & ~n16655;
  assign n33228 = n16655 & n33204;
  assign n33229 = ~pi39 & ~n33227;
  assign n33230 = ~n33228 & n33229;
  assign n33231 = ~pi38 & ~n33230;
  assign n33232 = ~n33226 & n33231;
  assign n33233 = ~n33214 & ~n33232;
  assign n33234 = pi698 & ~n33233;
  assign n33235 = ~n21041 & n33230;
  assign n33236 = ~pi197 & n20990;
  assign n33237 = pi197 & n21006;
  assign n33238 = ~pi767 & ~n33237;
  assign n33239 = ~n33236 & n33238;
  assign n33240 = ~pi197 & n21019;
  assign n33241 = pi197 & n21035;
  assign n33242 = pi299 & ~n33241;
  assign n33243 = ~n33240 & n33242;
  assign n33244 = n21038 & ~n33219;
  assign n33245 = pi767 & ~n33244;
  assign n33246 = ~n33243 & n33245;
  assign n33247 = pi39 & ~n33246;
  assign n33248 = ~n33239 & n33247;
  assign n33249 = ~n33235 & ~n33248;
  assign n33250 = ~pi38 & ~n33249;
  assign n33251 = ~pi197 & ~n16968;
  assign n33252 = pi767 & pi947;
  assign n33253 = ~pi39 & ~n33252;
  assign n33254 = n21170 & n33253;
  assign n33255 = pi38 & ~n33251;
  assign n33256 = ~n33254 & n33255;
  assign n33257 = ~pi698 & ~n33256;
  assign n33258 = ~n33250 & n33257;
  assign n33259 = ~n33234 & ~n33258;
  assign n33260 = n10178 & ~n33259;
  assign n33261 = ~pi197 & ~n10178;
  assign n33262 = ~pi832 & ~n33261;
  assign n33263 = ~n33260 & n33262;
  assign po354 = ~n33210 & ~n33263;
  assign n33265 = n3182 & ~n16655;
  assign n33266 = n18809 & ~n33265;
  assign n33267 = pi198 & ~n33266;
  assign n33268 = pi198 & ~n16785;
  assign n33269 = ~n6223 & n33268;
  assign n33270 = pi198 & ~n16661;
  assign n33271 = ~po1101 & ~n33270;
  assign n33272 = pi198 & ~n16750;
  assign n33273 = po1101 & ~n33272;
  assign n33274 = ~n33271 & ~n33273;
  assign n33275 = n6223 & n33274;
  assign n33276 = ~n3461 & ~n33275;
  assign n33277 = ~n33269 & n33276;
  assign n33278 = n3461 & ~n33270;
  assign n33279 = ~pi215 & ~n33278;
  assign n33280 = ~n33277 & n33279;
  assign n33281 = pi198 & ~n16683;
  assign n33282 = ~n33271 & n33281;
  assign n33283 = ~n6165 & ~n16679;
  assign n33284 = n6165 & ~n16677;
  assign n33285 = pi198 & ~n33284;
  assign n33286 = ~n33283 & n33285;
  assign n33287 = ~n6223 & n33286;
  assign n33288 = ~n33282 & ~n33287;
  assign n33289 = pi215 & ~n33288;
  assign n33290 = pi299 & ~n33289;
  assign n33291 = ~n33280 & n33290;
  assign n33292 = ~n6197 & n33268;
  assign n33293 = n6197 & n33274;
  assign n33294 = ~n3053 & ~n33293;
  assign n33295 = ~n33292 & n33294;
  assign n33296 = n3053 & ~n33270;
  assign n33297 = ~pi223 & ~n33296;
  assign n33298 = ~n33295 & n33297;
  assign n33299 = ~n6197 & n33286;
  assign n33300 = ~n33282 & ~n33299;
  assign n33301 = pi223 & ~n33300;
  assign n33302 = ~pi299 & ~n33301;
  assign n33303 = ~n33298 & n33302;
  assign n33304 = n3268 & n10959;
  assign n33305 = ~n33291 & n33304;
  assign n33306 = ~n33303 & n33305;
  assign n33307 = ~n33267 & ~n33306;
  assign n33308 = n17698 & ~n33307;
  assign n33309 = pi198 & ~n3268;
  assign n33310 = pi198 & ~n16649;
  assign n33311 = pi603 & pi633;
  assign n33312 = ~n33310 & ~n33311;
  assign n33313 = pi198 & ~n16822;
  assign n33314 = ~pi198 & n16915;
  assign n33315 = ~n33313 & ~n33314;
  assign n33316 = n33311 & n33315;
  assign n33317 = ~n33312 & ~n33316;
  assign n33318 = pi299 & n33317;
  assign n33319 = ~n16827 & ~n16831;
  assign n33320 = pi633 & ~n33319;
  assign n33321 = ~n16652 & ~n33320;
  assign n33322 = ~n16836 & ~n33321;
  assign n33323 = ~pi299 & n33322;
  assign n33324 = ~pi39 & ~n33323;
  assign n33325 = ~n33318 & n33324;
  assign n33326 = pi633 & n16661;
  assign n33327 = ~n16841 & n33326;
  assign n33328 = ~n33270 & ~n33327;
  assign n33329 = pi603 & ~n33328;
  assign n33330 = ~pi603 & n33270;
  assign n33331 = ~n33329 & ~n33330;
  assign n33332 = ~n16854 & n33331;
  assign n33333 = n6170 & ~n33328;
  assign n33334 = ~n16677 & n33327;
  assign n33335 = ~n33281 & ~n33334;
  assign n33336 = ~n33333 & n33335;
  assign n33337 = pi603 & ~n33336;
  assign n33338 = n16854 & ~n33330;
  assign n33339 = ~n33337 & n33338;
  assign n33340 = ~n33332 & ~n33339;
  assign n33341 = ~n6168 & n33340;
  assign n33342 = ~n33281 & ~n33337;
  assign n33343 = n6168 & ~n33342;
  assign n33344 = ~n33341 & ~n33343;
  assign n33345 = n6197 & n33344;
  assign n33346 = pi633 & n16941;
  assign n33347 = ~n33286 & ~n33346;
  assign n33348 = ~n6168 & ~n33347;
  assign n33349 = pi198 & n16677;
  assign n33350 = ~n33334 & ~n33349;
  assign n33351 = n16885 & ~n33350;
  assign n33352 = ~n33348 & ~n33351;
  assign n33353 = ~n6197 & n33352;
  assign n33354 = pi223 & ~n33353;
  assign n33355 = ~n33345 & n33354;
  assign n33356 = pi198 & n16748;
  assign n33357 = pi633 & n17043;
  assign n33358 = ~n33356 & ~n33357;
  assign n33359 = ~n6170 & ~n33358;
  assign n33360 = ~n33333 & ~n33359;
  assign n33361 = pi603 & ~n33360;
  assign n33362 = ~pi642 & ~n33361;
  assign n33363 = pi642 & ~n33329;
  assign n33364 = n6164 & ~n33363;
  assign n33365 = ~n33362 & n33364;
  assign n33366 = ~n6164 & n33329;
  assign n33367 = ~n33330 & ~n33366;
  assign n33368 = ~n33365 & n33367;
  assign n33369 = ~n6168 & n33368;
  assign n33370 = ~pi603 & n33272;
  assign n33371 = n6168 & ~n33370;
  assign n33372 = ~n33361 & n33371;
  assign n33373 = ~n33369 & ~n33372;
  assign n33374 = n6197 & n33373;
  assign n33375 = pi603 & ~n33358;
  assign n33376 = n16854 & n33375;
  assign n33377 = n6170 & n33358;
  assign n33378 = ~n6170 & n33328;
  assign n33379 = pi603 & ~n16854;
  assign n33380 = ~n33378 & n33379;
  assign n33381 = ~n33377 & n33380;
  assign n33382 = pi198 & n17079;
  assign n33383 = ~n33376 & ~n33382;
  assign n33384 = ~n33381 & n33383;
  assign n33385 = ~n6168 & n33384;
  assign n33386 = n6168 & ~n33356;
  assign n33387 = ~n33375 & n33386;
  assign n33388 = ~n33385 & ~n33387;
  assign n33389 = ~n6197 & n33388;
  assign n33390 = ~n3053 & ~n33389;
  assign n33391 = ~n33374 & n33390;
  assign n33392 = n3053 & n33331;
  assign n33393 = ~pi223 & ~n33392;
  assign n33394 = ~n33391 & n33393;
  assign n33395 = ~n33355 & ~n33394;
  assign n33396 = ~pi299 & ~n33395;
  assign n33397 = n6223 & n33344;
  assign n33398 = ~n6223 & n33352;
  assign n33399 = pi215 & ~n33398;
  assign n33400 = ~n33397 & n33399;
  assign n33401 = n6223 & n33373;
  assign n33402 = ~n6223 & n33388;
  assign n33403 = ~n3461 & ~n33402;
  assign n33404 = ~n33401 & n33403;
  assign n33405 = n3461 & n33331;
  assign n33406 = ~pi215 & ~n33405;
  assign n33407 = ~n33404 & n33406;
  assign n33408 = ~n33400 & ~n33407;
  assign n33409 = pi299 & ~n33408;
  assign n33410 = pi39 & ~n33396;
  assign n33411 = ~n33409 & n33410;
  assign n33412 = ~n33325 & ~n33411;
  assign n33413 = ~pi38 & ~n33412;
  assign n33414 = pi39 & pi198;
  assign n33415 = pi38 & ~n33414;
  assign n33416 = pi198 & ~n16665;
  assign n33417 = pi633 & n16842;
  assign n33418 = n16665 & n33417;
  assign n33419 = ~n33416 & ~n33418;
  assign n33420 = ~pi39 & ~n33419;
  assign n33421 = n33415 & ~n33420;
  assign n33422 = n3268 & ~n33421;
  assign n33423 = ~n33413 & n33422;
  assign n33424 = ~n33309 & ~n33423;
  assign n33425 = ~n17526 & ~n33424;
  assign n33426 = n17526 & ~n33307;
  assign n33427 = ~n33425 & ~n33426;
  assign n33428 = ~pi785 & ~n33427;
  assign n33429 = ~n17527 & ~n33307;
  assign n33430 = pi609 & n33425;
  assign n33431 = ~n33429 & ~n33430;
  assign n33432 = pi1155 & ~n33431;
  assign n33433 = ~n17539 & ~n33307;
  assign n33434 = ~pi609 & n33425;
  assign n33435 = ~n33433 & ~n33434;
  assign n33436 = ~pi1155 & ~n33435;
  assign n33437 = ~n33432 & ~n33436;
  assign n33438 = pi785 & ~n33437;
  assign n33439 = ~n33428 & ~n33438;
  assign n33440 = ~pi781 & ~n33439;
  assign n33441 = pi618 & n33439;
  assign n33442 = ~pi618 & n33307;
  assign n33443 = pi1154 & ~n33442;
  assign n33444 = ~n33441 & n33443;
  assign n33445 = ~pi618 & n33439;
  assign n33446 = pi618 & n33307;
  assign n33447 = ~pi1154 & ~n33446;
  assign n33448 = ~n33445 & n33447;
  assign n33449 = ~n33444 & ~n33448;
  assign n33450 = pi781 & ~n33449;
  assign n33451 = ~n33440 & ~n33450;
  assign n33452 = ~pi789 & ~n33451;
  assign n33453 = pi619 & n33451;
  assign n33454 = ~pi619 & n33307;
  assign n33455 = pi1159 & ~n33454;
  assign n33456 = ~n33453 & n33455;
  assign n33457 = ~pi619 & n33451;
  assign n33458 = pi619 & n33307;
  assign n33459 = ~pi1159 & ~n33458;
  assign n33460 = ~n33457 & n33459;
  assign n33461 = ~n33456 & ~n33460;
  assign n33462 = pi789 & ~n33461;
  assign n33463 = ~n33452 & ~n33462;
  assign n33464 = ~n17904 & n33463;
  assign n33465 = n17904 & n33307;
  assign n33466 = ~n33464 & ~n33465;
  assign n33467 = ~n17698 & n33466;
  assign n33468 = ~n33308 & ~n33467;
  assign n33469 = ~n20491 & ~n33468;
  assign n33470 = ~n19215 & n33307;
  assign n33471 = n17591 & ~n33307;
  assign n33472 = ~n17076 & ~n33270;
  assign n33473 = pi634 & ~n33472;
  assign n33474 = ~n33270 & ~n33473;
  assign n33475 = ~n6165 & n33474;
  assign n33476 = n16976 & ~n33475;
  assign n33477 = n6170 & ~n33474;
  assign n33478 = pi634 & n17077;
  assign n33479 = ~n33356 & ~n33478;
  assign n33480 = ~n6170 & ~n33479;
  assign n33481 = ~n33477 & ~n33480;
  assign n33482 = n6165 & n33481;
  assign n33483 = n33476 & ~n33482;
  assign n33484 = n6168 & ~n33481;
  assign n33485 = n6165 & ~n33272;
  assign n33486 = ~n6165 & ~n33270;
  assign n33487 = ~pi680 & ~n33486;
  assign n33488 = ~n33485 & n33487;
  assign n33489 = ~n33484 & ~n33488;
  assign n33490 = ~n33483 & n33489;
  assign n33491 = n6197 & ~n33490;
  assign n33492 = ~n6170 & n33474;
  assign n33493 = n6170 & n33479;
  assign n33494 = ~n33492 & ~n33493;
  assign n33495 = ~n6165 & ~n33494;
  assign n33496 = n6165 & n33479;
  assign n33497 = n16976 & ~n33496;
  assign n33498 = ~n33495 & n33497;
  assign n33499 = pi198 & n17042;
  assign n33500 = n6168 & ~n33479;
  assign n33501 = ~n33499 & ~n33500;
  assign n33502 = ~n33498 & n33501;
  assign n33503 = ~n6197 & ~n33502;
  assign n33504 = ~n3053 & ~n33491;
  assign n33505 = ~n33503 & n33504;
  assign n33506 = pi680 & n33473;
  assign n33507 = ~n33270 & ~n33506;
  assign n33508 = n3053 & n33507;
  assign n33509 = ~pi223 & ~n33508;
  assign n33510 = ~n33505 & n33509;
  assign n33511 = pi634 & ~n16677;
  assign n33512 = n17076 & n33511;
  assign n33513 = ~n33349 & ~n33512;
  assign n33514 = n6170 & n33513;
  assign n33515 = ~n33492 & ~n33514;
  assign n33516 = ~n6165 & ~n33515;
  assign n33517 = n6165 & n33513;
  assign n33518 = n16976 & ~n33517;
  assign n33519 = ~n33516 & n33518;
  assign n33520 = ~pi680 & n33286;
  assign n33521 = n6168 & ~n33513;
  assign n33522 = ~n33520 & ~n33521;
  assign n33523 = ~n33519 & n33522;
  assign n33524 = ~n6197 & n33523;
  assign n33525 = ~n6170 & ~n33513;
  assign n33526 = ~n33477 & ~n33525;
  assign n33527 = n6165 & n33526;
  assign n33528 = n33476 & ~n33527;
  assign n33529 = n33281 & n33520;
  assign n33530 = n6168 & ~n33526;
  assign n33531 = ~n33529 & ~n33530;
  assign n33532 = ~n33528 & n33531;
  assign n33533 = n6197 & n33532;
  assign n33534 = pi223 & ~n33524;
  assign n33535 = ~n33533 & n33534;
  assign n33536 = ~pi299 & ~n33535;
  assign n33537 = ~n33510 & n33536;
  assign n33538 = ~n6223 & ~n33502;
  assign n33539 = n6223 & ~n33490;
  assign n33540 = ~n3461 & ~n33538;
  assign n33541 = ~n33539 & n33540;
  assign n33542 = n3461 & n33507;
  assign n33543 = ~pi215 & ~n33542;
  assign n33544 = ~n33541 & n33543;
  assign n33545 = ~n6223 & n33523;
  assign n33546 = n6223 & n33532;
  assign n33547 = pi215 & ~n33545;
  assign n33548 = ~n33546 & n33547;
  assign n33549 = pi299 & ~n33548;
  assign n33550 = ~n33544 & n33549;
  assign n33551 = ~n33537 & ~n33550;
  assign n33552 = pi39 & ~n33551;
  assign n33553 = pi634 & pi680;
  assign n33554 = ~pi198 & n17334;
  assign n33555 = pi198 & ~n17311;
  assign n33556 = ~n33554 & ~n33555;
  assign n33557 = n33553 & ~n33556;
  assign n33558 = n33310 & ~n33553;
  assign n33559 = ~n33557 & ~n33558;
  assign n33560 = pi299 & ~n33559;
  assign n33561 = pi198 & n17301;
  assign n33562 = ~n17321 & n33553;
  assign n33563 = ~n33561 & n33562;
  assign n33564 = ~n16652 & ~n33563;
  assign n33565 = ~pi299 & ~n33564;
  assign n33566 = ~pi39 & ~n33565;
  assign n33567 = ~n33560 & n33566;
  assign n33568 = ~n33552 & ~n33567;
  assign n33569 = ~pi38 & ~n33568;
  assign n33570 = pi634 & n17152;
  assign n33571 = n16665 & n33570;
  assign n33572 = ~n33416 & ~n33571;
  assign n33573 = ~pi39 & ~n33572;
  assign n33574 = n33415 & ~n33573;
  assign n33575 = n3268 & ~n33574;
  assign n33576 = ~n33569 & n33575;
  assign n33577 = ~n33309 & ~n33576;
  assign n33578 = ~pi778 & ~n33577;
  assign n33579 = pi625 & n33577;
  assign n33580 = ~pi625 & n33307;
  assign n33581 = pi1153 & ~n33580;
  assign n33582 = ~n33579 & n33581;
  assign n33583 = ~pi625 & n33577;
  assign n33584 = pi625 & n33307;
  assign n33585 = ~pi1153 & ~n33584;
  assign n33586 = ~n33583 & n33585;
  assign n33587 = ~n33582 & ~n33586;
  assign n33588 = pi778 & ~n33587;
  assign n33589 = ~n33578 & ~n33588;
  assign n33590 = ~n17554 & n33589;
  assign n33591 = n17554 & n33307;
  assign n33592 = ~n33590 & ~n33591;
  assign n33593 = ~n17591 & n33592;
  assign n33594 = ~n33471 & ~n33593;
  assign n33595 = ~n17627 & n33594;
  assign n33596 = ~n17670 & n33595;
  assign n33597 = ~n33470 & ~n33596;
  assign n33598 = ~pi792 & n33597;
  assign n33599 = pi628 & ~n33597;
  assign n33600 = ~pi628 & n33307;
  assign n33601 = ~n33599 & ~n33600;
  assign n33602 = pi1156 & n33601;
  assign n33603 = ~pi628 & ~n33597;
  assign n33604 = pi628 & n33307;
  assign n33605 = ~pi1156 & ~n33604;
  assign n33606 = ~n33603 & n33605;
  assign n33607 = ~n33602 & ~n33606;
  assign n33608 = pi792 & ~n33607;
  assign n33609 = ~n33598 & ~n33608;
  assign n33610 = ~pi647 & n33609;
  assign n33611 = pi647 & n33307;
  assign n33612 = ~pi1157 & ~n33611;
  assign n33613 = ~n33610 & n33612;
  assign n33614 = pi647 & ~n33609;
  assign n33615 = ~pi647 & ~n33307;
  assign n33616 = ~n33614 & ~n33615;
  assign n33617 = pi1157 & ~n33616;
  assign n33618 = ~n33613 & ~n33617;
  assign n33619 = ~n17739 & ~n33618;
  assign n33620 = ~n33469 & ~n33619;
  assign n33621 = pi787 & ~n33620;
  assign n33622 = ~n20502 & n33466;
  assign n33623 = pi629 & n33606;
  assign n33624 = n17695 & n33601;
  assign n33625 = ~n33623 & ~n33624;
  assign n33626 = ~n33622 & n33625;
  assign n33627 = pi792 & ~n33626;
  assign n33628 = ~pi626 & ~n33463;
  assign n33629 = pi626 & ~n33307;
  assign n33630 = n17668 & ~n33629;
  assign n33631 = ~n33628 & n33630;
  assign n33632 = pi626 & ~n33463;
  assign n33633 = ~pi626 & ~n33307;
  assign n33634 = n17667 & ~n33633;
  assign n33635 = ~n33632 & n33634;
  assign n33636 = n17627 & n33307;
  assign n33637 = ~n33595 & ~n33636;
  assign n33638 = n17792 & ~n33637;
  assign n33639 = ~n33631 & ~n33638;
  assign n33640 = ~n33635 & n33639;
  assign n33641 = pi788 & ~n33640;
  assign n33642 = ~pi603 & ~n33556;
  assign n33643 = pi198 & ~pi665;
  assign n33644 = pi633 & ~n33643;
  assign n33645 = ~n33554 & n33644;
  assign n33646 = n33315 & n33645;
  assign n33647 = ~n16915 & n33555;
  assign n33648 = ~pi198 & ~pi665;
  assign n33649 = n16822 & n33648;
  assign n33650 = ~pi633 & ~n33649;
  assign n33651 = ~n33647 & n33650;
  assign n33652 = pi603 & ~n33651;
  assign n33653 = ~n33646 & n33652;
  assign n33654 = ~n33642 & ~n33653;
  assign n33655 = n33553 & ~n33654;
  assign n33656 = n33317 & ~n33553;
  assign n33657 = pi299 & ~n33656;
  assign n33658 = ~n33655 & n33657;
  assign n33659 = ~pi634 & n16652;
  assign n33660 = pi634 & ~n16833;
  assign n33661 = n17302 & n33660;
  assign n33662 = ~n33659 & ~n33661;
  assign n33663 = ~pi633 & ~n33662;
  assign n33664 = pi198 & ~pi633;
  assign n33665 = pi634 & ~pi665;
  assign n33666 = ~n33664 & n33665;
  assign n33667 = ~n16826 & n33666;
  assign n33668 = pi603 & ~n33667;
  assign n33669 = ~n33320 & n33668;
  assign n33670 = ~n33663 & n33669;
  assign n33671 = ~pi603 & n33564;
  assign n33672 = pi680 & ~n33671;
  assign n33673 = ~n33670 & n33672;
  assign n33674 = ~pi680 & n33322;
  assign n33675 = ~pi299 & ~n33674;
  assign n33676 = ~n33673 & n33675;
  assign n33677 = ~n33658 & ~n33676;
  assign n33678 = ~pi39 & ~n33677;
  assign n33679 = ~pi680 & n33368;
  assign n33680 = n16845 & n33665;
  assign n33681 = n33328 & ~n33680;
  assign n33682 = n6170 & ~n33681;
  assign n33683 = pi634 & n17087;
  assign n33684 = n33358 & ~n33683;
  assign n33685 = ~n6170 & ~n33684;
  assign n33686 = ~n33682 & ~n33685;
  assign n33687 = pi603 & ~n33686;
  assign n33688 = ~pi642 & n33687;
  assign n33689 = ~pi603 & ~n33474;
  assign n33690 = pi603 & ~n33681;
  assign n33691 = pi642 & n33690;
  assign n33692 = ~n33689 & ~n33691;
  assign n33693 = ~n33688 & n33692;
  assign n33694 = n6164 & ~n33693;
  assign n33695 = ~n33689 & ~n33690;
  assign n33696 = ~n6164 & ~n33695;
  assign n33697 = ~n16708 & ~n33696;
  assign n33698 = ~n33694 & n33697;
  assign n33699 = ~pi603 & ~n33481;
  assign n33700 = n16708 & ~n33699;
  assign n33701 = ~n33687 & n33700;
  assign n33702 = ~n33698 & ~n33701;
  assign n33703 = pi680 & ~n33702;
  assign n33704 = ~n33679 & ~n33703;
  assign n33705 = n6197 & n33704;
  assign n33706 = ~pi680 & ~n33384;
  assign n33707 = ~pi603 & n33494;
  assign n33708 = ~n16854 & n33690;
  assign n33709 = ~n33380 & ~n33708;
  assign n33710 = ~n6165 & n33709;
  assign n33711 = ~n6170 & ~n33709;
  assign n33712 = n33684 & ~n33711;
  assign n33713 = ~n33710 & ~n33712;
  assign n33714 = ~n33707 & ~n33713;
  assign n33715 = n16976 & ~n33714;
  assign n33716 = ~n16842 & ~n33479;
  assign n33717 = ~n33375 & ~n33716;
  assign n33718 = n6168 & ~n33717;
  assign n33719 = ~n33706 & ~n33718;
  assign n33720 = ~n33715 & n33719;
  assign n33721 = ~n6197 & ~n33720;
  assign n33722 = ~n3053 & ~n33721;
  assign n33723 = ~n33705 & n33722;
  assign n33724 = n17054 & n33473;
  assign n33725 = n33331 & ~n33724;
  assign n33726 = n3053 & n33725;
  assign n33727 = ~pi223 & ~n33726;
  assign n33728 = ~n33723 & n33727;
  assign n33729 = n16868 & n33648;
  assign n33730 = n16841 & n33643;
  assign n33731 = ~n33349 & ~n33730;
  assign n33732 = ~n33729 & n33731;
  assign n33733 = pi634 & ~n33732;
  assign n33734 = ~pi634 & n33349;
  assign n33735 = ~n33334 & ~n33734;
  assign n33736 = ~n33733 & n33735;
  assign n33737 = ~n6170 & ~n33736;
  assign n33738 = ~n33682 & ~n33737;
  assign n33739 = pi603 & ~n33738;
  assign n33740 = ~pi603 & ~n33526;
  assign n33741 = ~n33739 & ~n33740;
  assign n33742 = n6168 & ~n33741;
  assign n33743 = n16854 & ~n33689;
  assign n33744 = ~n33739 & n33743;
  assign n33745 = ~n16854 & n33695;
  assign n33746 = n16976 & ~n33745;
  assign n33747 = ~n33744 & n33746;
  assign n33748 = ~pi680 & n33340;
  assign n33749 = ~n33742 & ~n33748;
  assign n33750 = ~n33747 & n33749;
  assign n33751 = n6197 & n33750;
  assign n33752 = ~pi603 & n33515;
  assign n33753 = pi603 & ~n33736;
  assign n33754 = n16854 & n33753;
  assign n33755 = ~n33709 & ~n33736;
  assign n33756 = ~n33711 & ~n33752;
  assign n33757 = ~n33754 & ~n33755;
  assign n33758 = n33756 & n33757;
  assign n33759 = n16976 & ~n33758;
  assign n33760 = ~pi680 & ~n33347;
  assign n33761 = ~pi603 & ~n33513;
  assign n33762 = ~n33753 & ~n33761;
  assign n33763 = n6168 & ~n33762;
  assign n33764 = ~n33760 & ~n33763;
  assign n33765 = ~n33759 & n33764;
  assign n33766 = ~n6197 & n33765;
  assign n33767 = pi223 & ~n33766;
  assign n33768 = ~n33751 & n33767;
  assign n33769 = ~n33728 & ~n33768;
  assign n33770 = ~pi299 & ~n33769;
  assign n33771 = n6223 & n33704;
  assign n33772 = ~n6223 & ~n33720;
  assign n33773 = ~n3461 & ~n33772;
  assign n33774 = ~n33771 & n33773;
  assign n33775 = n3461 & n33725;
  assign n33776 = ~pi215 & ~n33775;
  assign n33777 = ~n33774 & n33776;
  assign n33778 = n6223 & n33750;
  assign n33779 = ~n6223 & n33765;
  assign n33780 = pi215 & ~n33779;
  assign n33781 = ~n33778 & n33780;
  assign n33782 = ~n33777 & ~n33781;
  assign n33783 = pi299 & ~n33782;
  assign n33784 = pi39 & ~n33770;
  assign n33785 = ~n33783 & n33784;
  assign n33786 = ~n33678 & ~n33785;
  assign n33787 = ~pi38 & ~n33786;
  assign n33788 = pi634 & n17365;
  assign n33789 = n33419 & ~n33788;
  assign n33790 = ~pi39 & ~n33789;
  assign n33791 = n33415 & ~n33790;
  assign n33792 = n3268 & ~n33791;
  assign n33793 = ~n33787 & n33792;
  assign n33794 = ~n33309 & ~n33793;
  assign n33795 = ~pi625 & n33794;
  assign n33796 = pi625 & n33424;
  assign n33797 = ~pi1153 & ~n33796;
  assign n33798 = ~n33795 & n33797;
  assign n33799 = ~pi608 & ~n33582;
  assign n33800 = ~n33798 & n33799;
  assign n33801 = pi625 & n33794;
  assign n33802 = ~pi625 & n33424;
  assign n33803 = pi1153 & ~n33802;
  assign n33804 = ~n33801 & n33803;
  assign n33805 = pi608 & ~n33586;
  assign n33806 = ~n33804 & n33805;
  assign n33807 = ~n33800 & ~n33806;
  assign n33808 = pi778 & ~n33807;
  assign n33809 = ~pi778 & n33794;
  assign n33810 = ~n33808 & ~n33809;
  assign n33811 = ~pi609 & ~n33810;
  assign n33812 = pi609 & n33589;
  assign n33813 = ~pi1155 & ~n33812;
  assign n33814 = ~n33811 & n33813;
  assign n33815 = ~pi660 & ~n33432;
  assign n33816 = ~n33814 & n33815;
  assign n33817 = pi609 & ~n33810;
  assign n33818 = ~pi609 & n33589;
  assign n33819 = pi1155 & ~n33818;
  assign n33820 = ~n33817 & n33819;
  assign n33821 = pi660 & ~n33436;
  assign n33822 = ~n33820 & n33821;
  assign n33823 = ~n33816 & ~n33822;
  assign n33824 = pi785 & ~n33823;
  assign n33825 = ~pi785 & ~n33810;
  assign n33826 = ~n33824 & ~n33825;
  assign n33827 = ~pi618 & ~n33826;
  assign n33828 = pi618 & ~n33592;
  assign n33829 = ~pi1154 & ~n33828;
  assign n33830 = ~n33827 & n33829;
  assign n33831 = ~pi627 & ~n33444;
  assign n33832 = ~n33830 & n33831;
  assign n33833 = pi618 & ~n33826;
  assign n33834 = ~pi618 & ~n33592;
  assign n33835 = pi1154 & ~n33834;
  assign n33836 = ~n33833 & n33835;
  assign n33837 = pi627 & ~n33448;
  assign n33838 = ~n33836 & n33837;
  assign n33839 = ~n33832 & ~n33838;
  assign n33840 = pi781 & ~n33839;
  assign n33841 = ~pi781 & ~n33826;
  assign n33842 = ~n33840 & ~n33841;
  assign n33843 = ~pi619 & ~n33842;
  assign n33844 = pi619 & n33594;
  assign n33845 = ~pi1159 & ~n33844;
  assign n33846 = ~n33843 & n33845;
  assign n33847 = ~pi648 & ~n33456;
  assign n33848 = ~n33846 & n33847;
  assign n33849 = pi619 & ~n33842;
  assign n33850 = ~pi619 & n33594;
  assign n33851 = pi1159 & ~n33850;
  assign n33852 = ~n33849 & n33851;
  assign n33853 = pi648 & ~n33460;
  assign n33854 = ~n33852 & n33853;
  assign n33855 = pi789 & ~n33848;
  assign n33856 = ~n33854 & n33855;
  assign n33857 = ~pi789 & n33842;
  assign n33858 = n17905 & ~n33857;
  assign n33859 = ~n33856 & n33858;
  assign n33860 = ~n33641 & ~n33859;
  assign n33861 = ~n33627 & ~n33860;
  assign n33862 = n20298 & n33626;
  assign n33863 = n20300 & ~n33862;
  assign n33864 = ~n33861 & n33863;
  assign n33865 = ~n33621 & ~n33864;
  assign n33866 = ~pi790 & ~n33865;
  assign n33867 = pi644 & n33865;
  assign n33868 = ~pi787 & ~n33609;
  assign n33869 = pi787 & ~n33618;
  assign n33870 = ~n33868 & ~n33869;
  assign n33871 = ~pi644 & n33870;
  assign n33872 = pi715 & ~n33871;
  assign n33873 = ~n33867 & n33872;
  assign n33874 = ~n17740 & n33468;
  assign n33875 = n17740 & n33307;
  assign n33876 = ~n33874 & ~n33875;
  assign n33877 = pi644 & ~n33876;
  assign n33878 = ~pi644 & n33307;
  assign n33879 = ~pi715 & ~n33878;
  assign n33880 = ~n33877 & n33879;
  assign n33881 = pi1160 & ~n33880;
  assign n33882 = ~n33873 & n33881;
  assign n33883 = ~pi644 & n33865;
  assign n33884 = pi644 & n33870;
  assign n33885 = ~pi715 & ~n33884;
  assign n33886 = ~n33883 & n33885;
  assign n33887 = ~pi644 & ~n33876;
  assign n33888 = pi644 & n33307;
  assign n33889 = pi715 & ~n33888;
  assign n33890 = ~n33887 & n33889;
  assign n33891 = ~pi1160 & ~n33890;
  assign n33892 = ~n33886 & n33891;
  assign n33893 = pi790 & ~n33882;
  assign n33894 = ~n33892 & n33893;
  assign n33895 = ~n33866 & ~n33894;
  assign n33896 = ~po1038 & ~n33895;
  assign n33897 = pi198 & po1038;
  assign po355 = n33896 | n33897;
  assign n33899 = pi199 & ~n17494;
  assign n33900 = ~pi617 & ~n33899;
  assign n33901 = ~pi199 & ~n19342;
  assign n33902 = n19348 & ~n33901;
  assign n33903 = pi199 & n16907;
  assign n33904 = ~pi199 & ~n16963;
  assign n33905 = ~pi38 & ~n33904;
  assign n33906 = ~n33903 & n33905;
  assign n33907 = ~n33902 & ~n33906;
  assign n33908 = n3268 & ~n33907;
  assign n33909 = pi199 & ~n3268;
  assign n33910 = pi617 & ~n33909;
  assign n33911 = ~n33908 & n33910;
  assign n33912 = ~n33900 & ~n33911;
  assign n33913 = ~pi637 & n33912;
  assign n33914 = pi199 & n19308;
  assign n33915 = n3268 & ~n24462;
  assign n33916 = ~pi199 & ~n33915;
  assign n33917 = ~pi617 & ~n19304;
  assign n33918 = ~n33916 & n33917;
  assign n33919 = ~n33914 & n33918;
  assign n33920 = n3268 & n19326;
  assign n33921 = ~pi199 & ~n33920;
  assign n33922 = pi199 & n19334;
  assign n33923 = pi617 & ~n33922;
  assign n33924 = ~n33921 & n33923;
  assign n33925 = ~n33909 & ~n33924;
  assign n33926 = ~n33919 & n33925;
  assign n33927 = pi637 & ~n33926;
  assign n33928 = ~n33913 & ~n33927;
  assign n33929 = ~pi625 & n33928;
  assign n33930 = pi625 & ~n33912;
  assign n33931 = ~pi1153 & ~n33930;
  assign n33932 = ~n33929 & n33931;
  assign n33933 = ~pi637 & ~n33899;
  assign n33934 = ~pi199 & ~n16968;
  assign n33935 = n19892 & ~n33934;
  assign n33936 = pi199 & ~n17469;
  assign n33937 = ~pi199 & ~n17419;
  assign n33938 = pi39 & ~n33937;
  assign n33939 = ~n33936 & n33938;
  assign n33940 = pi199 & ~n17315;
  assign n33941 = ~pi199 & n17350;
  assign n33942 = ~pi39 & ~n33940;
  assign n33943 = ~n33941 & n33942;
  assign n33944 = ~pi38 & ~n33943;
  assign n33945 = ~n33939 & n33944;
  assign n33946 = ~n33935 & ~n33945;
  assign n33947 = n3268 & ~n33946;
  assign n33948 = pi637 & ~n33909;
  assign n33949 = ~n33947 & n33948;
  assign n33950 = ~n33933 & ~n33949;
  assign n33951 = pi625 & ~n33950;
  assign n33952 = ~pi625 & ~n33899;
  assign n33953 = pi1153 & ~n33952;
  assign n33954 = ~n33951 & n33953;
  assign n33955 = ~pi608 & ~n33954;
  assign n33956 = ~n33932 & n33955;
  assign n33957 = pi625 & n33928;
  assign n33958 = ~pi625 & ~n33912;
  assign n33959 = pi1153 & ~n33958;
  assign n33960 = ~n33957 & n33959;
  assign n33961 = ~pi625 & ~n33950;
  assign n33962 = pi625 & ~n33899;
  assign n33963 = ~pi1153 & ~n33962;
  assign n33964 = ~n33961 & n33963;
  assign n33965 = pi608 & ~n33964;
  assign n33966 = ~n33960 & n33965;
  assign n33967 = ~n33956 & ~n33966;
  assign n33968 = pi778 & ~n33967;
  assign n33969 = ~pi778 & n33928;
  assign n33970 = ~n33968 & ~n33969;
  assign n33971 = ~pi609 & ~n33970;
  assign n33972 = ~pi778 & n33950;
  assign n33973 = ~n33954 & ~n33964;
  assign n33974 = pi778 & ~n33973;
  assign n33975 = ~n33972 & ~n33974;
  assign n33976 = pi609 & n33975;
  assign n33977 = ~pi1155 & ~n33976;
  assign n33978 = ~n33971 & n33977;
  assign n33979 = ~n17526 & ~n33912;
  assign n33980 = n17526 & ~n33899;
  assign n33981 = ~n33979 & ~n33980;
  assign n33982 = pi609 & ~n33981;
  assign n33983 = ~pi609 & ~n33899;
  assign n33984 = pi1155 & ~n33983;
  assign n33985 = ~n33982 & n33984;
  assign n33986 = ~pi660 & ~n33985;
  assign n33987 = ~n33978 & n33986;
  assign n33988 = pi609 & ~n33970;
  assign n33989 = ~pi609 & n33975;
  assign n33990 = pi1155 & ~n33989;
  assign n33991 = ~n33988 & n33990;
  assign n33992 = ~pi609 & ~n33981;
  assign n33993 = pi609 & ~n33899;
  assign n33994 = ~pi1155 & ~n33993;
  assign n33995 = ~n33992 & n33994;
  assign n33996 = pi660 & ~n33995;
  assign n33997 = ~n33991 & n33996;
  assign n33998 = ~n33987 & ~n33997;
  assign n33999 = pi785 & ~n33998;
  assign n34000 = ~pi785 & ~n33970;
  assign n34001 = ~n33999 & ~n34000;
  assign n34002 = ~pi618 & ~n34001;
  assign n34003 = n17554 & ~n33899;
  assign n34004 = ~n17554 & n33975;
  assign n34005 = ~n34003 & ~n34004;
  assign n34006 = pi618 & ~n34005;
  assign n34007 = ~pi1154 & ~n34006;
  assign n34008 = ~n34002 & n34007;
  assign n34009 = ~pi785 & n33981;
  assign n34010 = ~n33985 & ~n33995;
  assign n34011 = pi785 & ~n34010;
  assign n34012 = ~n34009 & ~n34011;
  assign n34013 = pi618 & n34012;
  assign n34014 = ~pi618 & ~n33899;
  assign n34015 = pi1154 & ~n34014;
  assign n34016 = ~n34013 & n34015;
  assign n34017 = ~pi627 & ~n34016;
  assign n34018 = ~n34008 & n34017;
  assign n34019 = pi618 & ~n34001;
  assign n34020 = ~pi618 & ~n34005;
  assign n34021 = pi1154 & ~n34020;
  assign n34022 = ~n34019 & n34021;
  assign n34023 = ~pi618 & n34012;
  assign n34024 = pi618 & ~n33899;
  assign n34025 = ~pi1154 & ~n34024;
  assign n34026 = ~n34023 & n34025;
  assign n34027 = pi627 & ~n34026;
  assign n34028 = ~n34022 & n34027;
  assign n34029 = ~n34018 & ~n34028;
  assign n34030 = pi781 & ~n34029;
  assign n34031 = ~pi781 & ~n34001;
  assign n34032 = ~n34030 & ~n34031;
  assign n34033 = ~pi619 & ~n34032;
  assign n34034 = ~n17591 & n34005;
  assign n34035 = n17591 & n33899;
  assign n34036 = ~n34034 & ~n34035;
  assign n34037 = pi619 & n34036;
  assign n34038 = ~pi1159 & ~n34037;
  assign n34039 = ~n34033 & n34038;
  assign n34040 = ~pi781 & ~n34012;
  assign n34041 = ~n34016 & ~n34026;
  assign n34042 = pi781 & ~n34041;
  assign n34043 = ~n34040 & ~n34042;
  assign n34044 = pi619 & n34043;
  assign n34045 = ~pi619 & ~n33899;
  assign n34046 = pi1159 & ~n34045;
  assign n34047 = ~n34044 & n34046;
  assign n34048 = ~pi648 & ~n34047;
  assign n34049 = ~n34039 & n34048;
  assign n34050 = pi619 & ~n34032;
  assign n34051 = ~pi619 & n34036;
  assign n34052 = pi1159 & ~n34051;
  assign n34053 = ~n34050 & n34052;
  assign n34054 = ~pi619 & n34043;
  assign n34055 = pi619 & ~n33899;
  assign n34056 = ~pi1159 & ~n34055;
  assign n34057 = ~n34054 & n34056;
  assign n34058 = pi648 & ~n34057;
  assign n34059 = ~n34053 & n34058;
  assign n34060 = ~n34049 & ~n34059;
  assign n34061 = pi789 & ~n34060;
  assign n34062 = ~pi789 & ~n34032;
  assign n34063 = ~n34061 & ~n34062;
  assign n34064 = ~pi788 & n34063;
  assign n34065 = ~pi626 & n34063;
  assign n34066 = n17627 & ~n33899;
  assign n34067 = ~n17627 & n34036;
  assign n34068 = ~n34066 & ~n34067;
  assign n34069 = pi626 & n34068;
  assign n34070 = ~pi641 & ~n34069;
  assign n34071 = ~n34065 & n34070;
  assign n34072 = ~pi789 & ~n34043;
  assign n34073 = ~n34047 & ~n34057;
  assign n34074 = pi789 & ~n34073;
  assign n34075 = ~n34072 & ~n34074;
  assign n34076 = ~pi626 & ~n34075;
  assign n34077 = pi626 & n33899;
  assign n34078 = pi641 & ~n34077;
  assign n34079 = ~n34076 & n34078;
  assign n34080 = ~pi1158 & ~n34079;
  assign n34081 = ~n34071 & n34080;
  assign n34082 = pi626 & n34063;
  assign n34083 = ~pi626 & n34068;
  assign n34084 = pi641 & ~n34083;
  assign n34085 = ~n34082 & n34084;
  assign n34086 = pi626 & ~n34075;
  assign n34087 = ~pi626 & n33899;
  assign n34088 = ~pi641 & ~n34087;
  assign n34089 = ~n34086 & n34088;
  assign n34090 = pi1158 & ~n34089;
  assign n34091 = ~n34085 & n34090;
  assign n34092 = ~n34081 & ~n34091;
  assign n34093 = pi788 & ~n34092;
  assign n34094 = ~n34064 & ~n34093;
  assign n34095 = ~pi628 & n34094;
  assign n34096 = ~n17904 & ~n34075;
  assign n34097 = n17904 & n33899;
  assign n34098 = ~n34096 & ~n34097;
  assign n34099 = pi628 & n34098;
  assign n34100 = ~pi1156 & ~n34099;
  assign n34101 = ~n34095 & n34100;
  assign n34102 = ~n17670 & n34068;
  assign n34103 = n17670 & n33899;
  assign n34104 = ~n34102 & ~n34103;
  assign n34105 = pi628 & n34104;
  assign n34106 = ~pi628 & ~n33899;
  assign n34107 = pi1156 & ~n34106;
  assign n34108 = ~n34105 & n34107;
  assign n34109 = ~pi629 & ~n34108;
  assign n34110 = ~n34101 & n34109;
  assign n34111 = pi628 & n34094;
  assign n34112 = ~pi628 & n34098;
  assign n34113 = pi1156 & ~n34112;
  assign n34114 = ~n34111 & n34113;
  assign n34115 = ~pi628 & n34104;
  assign n34116 = pi628 & ~n33899;
  assign n34117 = ~pi1156 & ~n34116;
  assign n34118 = ~n34115 & n34117;
  assign n34119 = pi629 & ~n34118;
  assign n34120 = ~n34114 & n34119;
  assign n34121 = ~n34110 & ~n34120;
  assign n34122 = pi792 & ~n34121;
  assign n34123 = ~pi792 & n34094;
  assign n34124 = ~n34122 & ~n34123;
  assign n34125 = ~pi647 & ~n34124;
  assign n34126 = ~n17698 & ~n34098;
  assign n34127 = n17698 & n33899;
  assign n34128 = ~n34126 & ~n34127;
  assign n34129 = pi647 & n34128;
  assign n34130 = ~pi1157 & ~n34129;
  assign n34131 = ~n34125 & n34130;
  assign n34132 = ~pi792 & ~n34104;
  assign n34133 = ~n34108 & ~n34118;
  assign n34134 = pi792 & ~n34133;
  assign n34135 = ~n34132 & ~n34134;
  assign n34136 = pi647 & n34135;
  assign n34137 = ~pi647 & ~n33899;
  assign n34138 = pi1157 & ~n34137;
  assign n34139 = ~n34136 & n34138;
  assign n34140 = ~pi630 & ~n34139;
  assign n34141 = ~n34131 & n34140;
  assign n34142 = pi647 & ~n34124;
  assign n34143 = ~pi647 & n34128;
  assign n34144 = pi1157 & ~n34143;
  assign n34145 = ~n34142 & n34144;
  assign n34146 = ~pi647 & n34135;
  assign n34147 = pi647 & ~n33899;
  assign n34148 = ~pi1157 & ~n34147;
  assign n34149 = ~n34146 & n34148;
  assign n34150 = pi630 & ~n34149;
  assign n34151 = ~n34145 & n34150;
  assign n34152 = ~n34141 & ~n34151;
  assign n34153 = pi787 & ~n34152;
  assign n34154 = ~pi787 & ~n34124;
  assign n34155 = ~n34153 & ~n34154;
  assign n34156 = ~pi790 & n34155;
  assign n34157 = pi644 & ~n34155;
  assign n34158 = ~pi787 & ~n34135;
  assign n34159 = ~n34139 & ~n34149;
  assign n34160 = pi787 & ~n34159;
  assign n34161 = ~n34158 & ~n34160;
  assign n34162 = ~pi644 & n34161;
  assign n34163 = pi715 & ~n34162;
  assign n34164 = ~n34157 & n34163;
  assign n34165 = n17740 & ~n33899;
  assign n34166 = ~n17740 & n34128;
  assign n34167 = ~n34165 & ~n34166;
  assign n34168 = pi644 & ~n34167;
  assign n34169 = ~pi644 & ~n33899;
  assign n34170 = ~pi715 & ~n34169;
  assign n34171 = ~n34168 & n34170;
  assign n34172 = pi1160 & ~n34171;
  assign n34173 = ~n34164 & n34172;
  assign n34174 = ~pi644 & ~n34155;
  assign n34175 = pi644 & n34161;
  assign n34176 = ~pi715 & ~n34175;
  assign n34177 = ~n34174 & n34176;
  assign n34178 = ~pi644 & ~n34167;
  assign n34179 = pi644 & ~n33899;
  assign n34180 = pi715 & ~n34179;
  assign n34181 = ~n34178 & n34180;
  assign n34182 = ~pi1160 & ~n34181;
  assign n34183 = ~n34177 & n34182;
  assign n34184 = pi790 & ~n34173;
  assign n34185 = ~n34183 & n34184;
  assign n34186 = ~n34156 & ~n34185;
  assign n34187 = ~po1038 & ~n34186;
  assign n34188 = pi199 & po1038;
  assign po356 = n34187 | n34188;
  assign n34190 = pi200 & ~n17494;
  assign n34191 = ~pi606 & ~n34190;
  assign n34192 = ~pi200 & ~n19342;
  assign n34193 = n19348 & ~n34192;
  assign n34194 = pi200 & n16907;
  assign n34195 = ~pi200 & ~n16963;
  assign n34196 = ~pi38 & ~n34195;
  assign n34197 = ~n34194 & n34196;
  assign n34198 = ~n34193 & ~n34197;
  assign n34199 = n3268 & ~n34198;
  assign n34200 = pi200 & ~n3268;
  assign n34201 = pi606 & ~n34200;
  assign n34202 = ~n34199 & n34201;
  assign n34203 = ~n34191 & ~n34202;
  assign n34204 = ~n17526 & ~n34203;
  assign n34205 = n17526 & ~n34190;
  assign n34206 = ~n34204 & ~n34205;
  assign n34207 = ~pi785 & n34206;
  assign n34208 = pi609 & ~n34206;
  assign n34209 = ~pi609 & ~n34190;
  assign n34210 = pi1155 & ~n34209;
  assign n34211 = ~n34208 & n34210;
  assign n34212 = ~pi609 & ~n34206;
  assign n34213 = pi609 & ~n34190;
  assign n34214 = ~pi1155 & ~n34213;
  assign n34215 = ~n34212 & n34214;
  assign n34216 = ~n34211 & ~n34215;
  assign n34217 = pi785 & ~n34216;
  assign n34218 = ~n34207 & ~n34217;
  assign n34219 = ~pi781 & ~n34218;
  assign n34220 = pi618 & n34218;
  assign n34221 = ~pi618 & ~n34190;
  assign n34222 = pi1154 & ~n34221;
  assign n34223 = ~n34220 & n34222;
  assign n34224 = ~pi618 & n34218;
  assign n34225 = pi618 & ~n34190;
  assign n34226 = ~pi1154 & ~n34225;
  assign n34227 = ~n34224 & n34226;
  assign n34228 = ~n34223 & ~n34227;
  assign n34229 = pi781 & ~n34228;
  assign n34230 = ~n34219 & ~n34229;
  assign n34231 = ~pi789 & ~n34230;
  assign n34232 = pi619 & n34230;
  assign n34233 = ~pi619 & ~n34190;
  assign n34234 = pi1159 & ~n34233;
  assign n34235 = ~n34232 & n34234;
  assign n34236 = ~pi619 & n34230;
  assign n34237 = pi619 & ~n34190;
  assign n34238 = ~pi1159 & ~n34237;
  assign n34239 = ~n34236 & n34238;
  assign n34240 = ~n34235 & ~n34239;
  assign n34241 = pi789 & ~n34240;
  assign n34242 = ~n34231 & ~n34241;
  assign n34243 = ~n17904 & ~n34242;
  assign n34244 = n17904 & n34190;
  assign n34245 = ~n34243 & ~n34244;
  assign n34246 = ~n20502 & ~n34245;
  assign n34247 = n17627 & ~n34190;
  assign n34248 = n17554 & ~n34190;
  assign n34249 = ~pi643 & ~n34190;
  assign n34250 = ~pi200 & ~n16968;
  assign n34251 = n19892 & ~n34250;
  assign n34252 = pi200 & n17453;
  assign n34253 = ~pi200 & n17404;
  assign n34254 = ~pi299 & ~n34253;
  assign n34255 = ~n34252 & n34254;
  assign n34256 = pi200 & n17467;
  assign n34257 = ~pi200 & n17417;
  assign n34258 = pi299 & ~n34257;
  assign n34259 = ~n34256 & n34258;
  assign n34260 = ~n34255 & ~n34259;
  assign n34261 = pi39 & ~n34260;
  assign n34262 = ~pi200 & ~n17350;
  assign n34263 = pi200 & n17315;
  assign n34264 = ~pi39 & ~n34262;
  assign n34265 = ~n34263 & n34264;
  assign n34266 = ~n34261 & ~n34265;
  assign n34267 = ~pi38 & ~n34266;
  assign n34268 = ~n34251 & ~n34267;
  assign n34269 = n3268 & ~n34268;
  assign n34270 = pi643 & ~n34200;
  assign n34271 = ~n34269 & n34270;
  assign n34272 = ~n34249 & ~n34271;
  assign n34273 = ~pi778 & n34272;
  assign n34274 = pi625 & ~n34272;
  assign n34275 = ~pi625 & ~n34190;
  assign n34276 = pi1153 & ~n34275;
  assign n34277 = ~n34274 & n34276;
  assign n34278 = ~pi625 & ~n34272;
  assign n34279 = pi625 & ~n34190;
  assign n34280 = ~pi1153 & ~n34279;
  assign n34281 = ~n34278 & n34280;
  assign n34282 = ~n34277 & ~n34281;
  assign n34283 = pi778 & ~n34282;
  assign n34284 = ~n34273 & ~n34283;
  assign n34285 = ~n17554 & n34284;
  assign n34286 = ~n34248 & ~n34285;
  assign n34287 = ~n17591 & n34286;
  assign n34288 = n17591 & n34190;
  assign n34289 = ~n34287 & ~n34288;
  assign n34290 = ~n17627 & n34289;
  assign n34291 = ~n34247 & ~n34290;
  assign n34292 = ~n17670 & n34291;
  assign n34293 = n17670 & n34190;
  assign n34294 = ~n34292 & ~n34293;
  assign n34295 = pi628 & n34294;
  assign n34296 = ~pi628 & ~n34190;
  assign n34297 = pi1156 & ~n34296;
  assign n34298 = ~n34295 & n34297;
  assign n34299 = ~pi629 & n34298;
  assign n34300 = ~pi628 & n34294;
  assign n34301 = pi628 & ~n34190;
  assign n34302 = ~pi1156 & ~n34301;
  assign n34303 = ~n34300 & n34302;
  assign n34304 = pi629 & n34303;
  assign n34305 = ~n34299 & ~n34304;
  assign n34306 = ~n34246 & n34305;
  assign n34307 = pi792 & ~n34306;
  assign n34308 = ~pi643 & n34203;
  assign n34309 = pi200 & ~n19307;
  assign n34310 = ~pi200 & ~n19313;
  assign n34311 = ~pi38 & ~n34310;
  assign n34312 = ~n34309 & n34311;
  assign n34313 = ~n19303 & n34251;
  assign n34314 = ~n34312 & ~n34313;
  assign n34315 = ~pi606 & n3268;
  assign n34316 = ~n34314 & n34315;
  assign n34317 = ~n19321 & ~n19322;
  assign n34318 = ~pi200 & ~n34317;
  assign n34319 = pi200 & ~n24582;
  assign n34320 = ~pi200 & ~n19323;
  assign n34321 = ~pi38 & ~n34320;
  assign n34322 = ~n34319 & n34321;
  assign n34323 = pi38 & pi200;
  assign n34324 = n19331 & n34323;
  assign n34325 = pi606 & n3268;
  assign n34326 = ~n34324 & n34325;
  assign n34327 = ~n34318 & n34326;
  assign n34328 = ~n34322 & n34327;
  assign n34329 = ~n34200 & ~n34328;
  assign n34330 = ~n34316 & n34329;
  assign n34331 = pi643 & ~n34330;
  assign n34332 = ~n34308 & ~n34331;
  assign n34333 = ~pi625 & n34332;
  assign n34334 = pi625 & ~n34203;
  assign n34335 = ~pi1153 & ~n34334;
  assign n34336 = ~n34333 & n34335;
  assign n34337 = ~pi608 & ~n34277;
  assign n34338 = ~n34336 & n34337;
  assign n34339 = pi625 & n34332;
  assign n34340 = ~pi625 & ~n34203;
  assign n34341 = pi1153 & ~n34340;
  assign n34342 = ~n34339 & n34341;
  assign n34343 = pi608 & ~n34281;
  assign n34344 = ~n34342 & n34343;
  assign n34345 = ~n34338 & ~n34344;
  assign n34346 = pi778 & ~n34345;
  assign n34347 = ~pi778 & n34332;
  assign n34348 = ~n34346 & ~n34347;
  assign n34349 = ~pi609 & ~n34348;
  assign n34350 = pi609 & n34284;
  assign n34351 = ~pi1155 & ~n34350;
  assign n34352 = ~n34349 & n34351;
  assign n34353 = ~pi660 & ~n34211;
  assign n34354 = ~n34352 & n34353;
  assign n34355 = pi609 & ~n34348;
  assign n34356 = ~pi609 & n34284;
  assign n34357 = pi1155 & ~n34356;
  assign n34358 = ~n34355 & n34357;
  assign n34359 = pi660 & ~n34215;
  assign n34360 = ~n34358 & n34359;
  assign n34361 = ~n34354 & ~n34360;
  assign n34362 = pi785 & ~n34361;
  assign n34363 = ~pi785 & ~n34348;
  assign n34364 = ~n34362 & ~n34363;
  assign n34365 = ~pi618 & ~n34364;
  assign n34366 = pi618 & ~n34286;
  assign n34367 = ~pi1154 & ~n34366;
  assign n34368 = ~n34365 & n34367;
  assign n34369 = ~pi627 & ~n34223;
  assign n34370 = ~n34368 & n34369;
  assign n34371 = pi618 & ~n34364;
  assign n34372 = ~pi618 & ~n34286;
  assign n34373 = pi1154 & ~n34372;
  assign n34374 = ~n34371 & n34373;
  assign n34375 = pi627 & ~n34227;
  assign n34376 = ~n34374 & n34375;
  assign n34377 = ~n34370 & ~n34376;
  assign n34378 = pi781 & ~n34377;
  assign n34379 = ~pi781 & ~n34364;
  assign n34380 = ~n34378 & ~n34379;
  assign n34381 = ~pi619 & ~n34380;
  assign n34382 = pi619 & n34289;
  assign n34383 = ~pi1159 & ~n34382;
  assign n34384 = ~n34381 & n34383;
  assign n34385 = ~pi648 & ~n34235;
  assign n34386 = ~n34384 & n34385;
  assign n34387 = pi619 & ~n34380;
  assign n34388 = ~pi619 & n34289;
  assign n34389 = pi1159 & ~n34388;
  assign n34390 = ~n34387 & n34389;
  assign n34391 = pi648 & ~n34239;
  assign n34392 = ~n34390 & n34391;
  assign n34393 = pi789 & ~n34386;
  assign n34394 = ~n34392 & n34393;
  assign n34395 = ~pi789 & n34380;
  assign n34396 = n17905 & ~n34395;
  assign n34397 = ~n34394 & n34396;
  assign n34398 = ~pi626 & ~n34242;
  assign n34399 = pi626 & n34190;
  assign n34400 = n17668 & ~n34399;
  assign n34401 = ~n34398 & n34400;
  assign n34402 = pi626 & ~n34242;
  assign n34403 = ~pi626 & n34190;
  assign n34404 = n17667 & ~n34403;
  assign n34405 = ~n34402 & n34404;
  assign n34406 = n17792 & ~n34291;
  assign n34407 = ~n34401 & ~n34406;
  assign n34408 = ~n34405 & n34407;
  assign n34409 = pi788 & ~n34408;
  assign n34410 = ~n20298 & ~n34409;
  assign n34411 = ~n34397 & n34410;
  assign n34412 = ~n34307 & ~n34411;
  assign n34413 = n20300 & ~n34412;
  assign n34414 = ~n17698 & ~n34245;
  assign n34415 = n17698 & n34190;
  assign n34416 = ~n34414 & ~n34415;
  assign n34417 = ~n20491 & ~n34416;
  assign n34418 = ~pi792 & ~n34294;
  assign n34419 = ~n34298 & ~n34303;
  assign n34420 = pi792 & ~n34419;
  assign n34421 = ~n34418 & ~n34420;
  assign n34422 = ~pi647 & n34421;
  assign n34423 = pi647 & ~n34190;
  assign n34424 = ~pi1157 & ~n34423;
  assign n34425 = ~n34422 & n34424;
  assign n34426 = pi647 & ~n34421;
  assign n34427 = ~pi647 & n34190;
  assign n34428 = ~n34426 & ~n34427;
  assign n34429 = pi1157 & ~n34428;
  assign n34430 = ~n34425 & ~n34429;
  assign n34431 = ~n17739 & ~n34430;
  assign n34432 = ~n34417 & ~n34431;
  assign n34433 = pi787 & ~n34432;
  assign n34434 = ~n34413 & ~n34433;
  assign n34435 = ~pi644 & n34434;
  assign n34436 = ~pi787 & ~n34421;
  assign n34437 = pi787 & ~n34430;
  assign n34438 = ~n34436 & ~n34437;
  assign n34439 = pi644 & n34438;
  assign n34440 = ~pi715 & ~n34439;
  assign n34441 = ~n34435 & n34440;
  assign n34442 = ~n17740 & ~n34416;
  assign n34443 = n17740 & n34190;
  assign n34444 = ~n34442 & ~n34443;
  assign n34445 = ~pi644 & n34444;
  assign n34446 = pi644 & ~n34190;
  assign n34447 = pi715 & ~n34446;
  assign n34448 = ~n34445 & n34447;
  assign n34449 = ~pi1160 & ~n34448;
  assign n34450 = ~n34441 & n34449;
  assign n34451 = pi644 & n34434;
  assign n34452 = ~pi644 & n34438;
  assign n34453 = pi715 & ~n34452;
  assign n34454 = ~n34451 & n34453;
  assign n34455 = pi644 & n34444;
  assign n34456 = ~pi644 & ~n34190;
  assign n34457 = ~pi715 & ~n34456;
  assign n34458 = ~n34455 & n34457;
  assign n34459 = pi1160 & ~n34458;
  assign n34460 = ~n34454 & n34459;
  assign n34461 = ~n34450 & ~n34460;
  assign n34462 = pi790 & ~n34461;
  assign n34463 = ~pi790 & n34434;
  assign n34464 = ~n34462 & ~n34463;
  assign n34465 = ~po1038 & ~n34464;
  assign n34466 = ~pi200 & po1038;
  assign po357 = ~n34465 & ~n34466;
  assign n34468 = pi233 & pi237;
  assign n34469 = pi57 & pi332;
  assign n34470 = pi332 & ~n3294;
  assign n34471 = ~pi59 & ~n34470;
  assign n34472 = pi74 & pi332;
  assign n34473 = ~pi55 & ~n34472;
  assign n34474 = n2516 & n11063;
  assign n34475 = pi468 & n6165;
  assign n34476 = ~pi299 & pi587;
  assign n34477 = ~n20988 & ~n34476;
  assign n34478 = ~pi468 & ~n34477;
  assign n34479 = ~n34475 & ~n34478;
  assign n34480 = n34474 & ~n34479;
  assign n34481 = ~pi332 & ~n34480;
  assign n34482 = n7380 & ~n34481;
  assign n34483 = n3096 & n6607;
  assign n34484 = ~pi332 & ~n34483;
  assign n34485 = n15643 & ~n34484;
  assign n34486 = pi332 & ~n3239;
  assign n34487 = ~n34485 & ~n34486;
  assign n34488 = ~n34482 & n34487;
  assign n34489 = ~pi74 & ~n34488;
  assign n34490 = n34473 & ~n34489;
  assign n34491 = n3269 & n6563;
  assign n34492 = n3096 & n34491;
  assign n34493 = ~pi332 & ~n34492;
  assign n34494 = pi55 & n34493;
  assign n34495 = n3294 & ~n34494;
  assign n34496 = ~n34490 & n34495;
  assign n34497 = n34471 & ~n34496;
  assign n34498 = n6293 & ~n34493;
  assign n34499 = pi332 & ~n6293;
  assign n34500 = pi59 & ~n34499;
  assign n34501 = ~n34498 & n34500;
  assign n34502 = ~pi57 & ~n34501;
  assign n34503 = ~n34497 & n34502;
  assign n34504 = ~n34469 & ~n34503;
  assign n34505 = ~n34468 & ~n34504;
  assign n34506 = ~pi332 & ~n6165;
  assign n34507 = ~pi947 & ~n34506;
  assign n34508 = pi96 & pi210;
  assign n34509 = pi332 & n34508;
  assign n34510 = ~pi32 & pi70;
  assign n34511 = ~pi70 & ~pi841;
  assign n34512 = pi32 & n34511;
  assign n34513 = ~n34510 & ~n34512;
  assign n34514 = ~pi210 & ~n34513;
  assign n34515 = ~pi32 & ~pi96;
  assign n34516 = pi70 & n34515;
  assign n34517 = ~pi332 & ~n34516;
  assign n34518 = ~n34514 & n34517;
  assign n34519 = ~n34509 & ~n34518;
  assign n34520 = ~n6170 & n34519;
  assign n34521 = n6165 & ~n34520;
  assign n34522 = n34507 & ~n34521;
  assign n34523 = pi332 & pi468;
  assign n34524 = ~pi468 & ~n34518;
  assign n34525 = ~n34523 & ~n34524;
  assign n34526 = ~n6165 & n34525;
  assign n34527 = n6165 & ~n34519;
  assign n34528 = pi947 & ~n34527;
  assign n34529 = ~n34526 & n34528;
  assign n34530 = ~n34522 & ~n34529;
  assign n34531 = pi57 & ~n34530;
  assign n34532 = ~n3269 & n34530;
  assign n34533 = ~pi95 & n2720;
  assign n34534 = ~pi70 & ~n34533;
  assign n34535 = n34515 & ~n34534;
  assign n34536 = pi210 & n34535;
  assign n34537 = pi32 & ~n34511;
  assign n34538 = ~pi95 & n2783;
  assign n34539 = ~n34537 & n34538;
  assign n34540 = n2495 & n34539;
  assign n34541 = n2523 & n34540;
  assign n34542 = n34513 & ~n34541;
  assign n34543 = ~pi210 & ~n34542;
  assign n34544 = ~pi332 & ~n34543;
  assign n34545 = ~n34536 & n34544;
  assign n34546 = ~n34509 & ~n34545;
  assign n34547 = ~n6170 & n34546;
  assign n34548 = n6165 & ~n34547;
  assign n34549 = n34507 & ~n34548;
  assign n34550 = ~pi468 & ~n34545;
  assign n34551 = ~n34523 & ~n34550;
  assign n34552 = ~n6165 & n34551;
  assign n34553 = n6165 & ~n34546;
  assign n34554 = pi947 & ~n34553;
  assign n34555 = ~n34552 & n34554;
  assign n34556 = ~n34549 & ~n34555;
  assign n34557 = n3269 & n34556;
  assign n34558 = ~n34532 & ~n34557;
  assign n34559 = n6293 & ~n34558;
  assign n34560 = ~n6293 & n34530;
  assign n34561 = pi59 & ~n34560;
  assign n34562 = ~n34559 & n34561;
  assign n34563 = n2516 & n2536;
  assign n34564 = ~pi95 & n2450;
  assign n34565 = n34563 & n34564;
  assign n34566 = ~pi70 & ~n34565;
  assign n34567 = n34515 & ~n34566;
  assign n34568 = pi210 & n34567;
  assign n34569 = n34539 & n34563;
  assign n34570 = n34513 & ~n34569;
  assign n34571 = ~pi210 & ~n34570;
  assign n34572 = ~pi332 & ~n34571;
  assign n34573 = ~n34568 & n34572;
  assign n34574 = ~n34509 & ~n34573;
  assign n34575 = ~n6170 & n34574;
  assign n34576 = n6165 & ~n34575;
  assign n34577 = n34507 & ~n34576;
  assign n34578 = ~pi468 & ~n34573;
  assign n34579 = ~n34523 & ~n34578;
  assign n34580 = ~n6165 & n34579;
  assign n34581 = n6165 & ~n34574;
  assign n34582 = pi947 & ~n34581;
  assign n34583 = ~n34580 & n34582;
  assign n34584 = pi299 & ~n34577;
  assign n34585 = ~n34583 & n34584;
  assign n34586 = ~pi587 & ~n34506;
  assign n34587 = pi198 & n34567;
  assign n34588 = ~pi198 & ~n34570;
  assign n34589 = ~pi332 & ~n34588;
  assign n34590 = ~n34587 & n34589;
  assign n34591 = pi96 & pi198;
  assign n34592 = pi332 & n34591;
  assign n34593 = ~n34590 & ~n34592;
  assign n34594 = ~n6170 & n34593;
  assign n34595 = n6165 & ~n34594;
  assign n34596 = n34586 & ~n34595;
  assign n34597 = n6165 & ~n34593;
  assign n34598 = ~pi468 & ~n34590;
  assign n34599 = ~n6165 & ~n34523;
  assign n34600 = ~n34598 & n34599;
  assign n34601 = pi587 & ~n34597;
  assign n34602 = ~n34600 & n34601;
  assign n34603 = ~pi299 & ~n34596;
  assign n34604 = ~n34602 & n34603;
  assign n34605 = ~n34585 & ~n34604;
  assign n34606 = n7380 & ~n34605;
  assign n34607 = pi299 & ~n34556;
  assign n34608 = pi198 & n34535;
  assign n34609 = ~pi198 & ~n34542;
  assign n34610 = ~pi332 & ~n34609;
  assign n34611 = ~n34608 & n34610;
  assign n34612 = ~n34592 & ~n34611;
  assign n34613 = ~n6170 & n34612;
  assign n34614 = n6165 & ~n34613;
  assign n34615 = n34586 & ~n34614;
  assign n34616 = n6165 & ~n34612;
  assign n34617 = ~pi468 & ~n34611;
  assign n34618 = n34599 & ~n34617;
  assign n34619 = pi587 & ~n34616;
  assign n34620 = ~n34618 & n34619;
  assign n34621 = ~n34615 & ~n34620;
  assign n34622 = ~pi299 & ~n34621;
  assign n34623 = n15643 & ~n34607;
  assign n34624 = ~n34622 & n34623;
  assign n34625 = ~n34606 & ~n34624;
  assign n34626 = ~pi74 & ~n34625;
  assign n34627 = pi299 & ~n34530;
  assign n34628 = ~pi74 & n3239;
  assign n34629 = ~pi198 & ~n34513;
  assign n34630 = n34517 & ~n34629;
  assign n34631 = ~n34592 & ~n34630;
  assign n34632 = n6165 & ~n34631;
  assign n34633 = n6576 & ~n34630;
  assign n34634 = n34506 & ~n34633;
  assign n34635 = ~pi299 & ~n6575;
  assign n34636 = ~n34632 & n34635;
  assign n34637 = ~n34634 & n34636;
  assign n34638 = ~n34628 & ~n34637;
  assign n34639 = ~n34627 & n34638;
  assign n34640 = ~pi55 & ~n34639;
  assign n34641 = ~n34626 & n34640;
  assign n34642 = pi55 & n34558;
  assign n34643 = n3294 & ~n34642;
  assign n34644 = ~n34641 & n34643;
  assign n34645 = ~n3294 & n34530;
  assign n34646 = ~pi59 & ~n34645;
  assign n34647 = ~n34644 & n34646;
  assign n34648 = ~n34562 & ~n34647;
  assign n34649 = ~pi57 & ~n34648;
  assign n34650 = ~n34531 & ~n34649;
  assign n34651 = n34468 & ~n34650;
  assign n34652 = ~n34505 & ~n34651;
  assign n34653 = ~pi201 & ~n34652;
  assign n34654 = ~n16429 & ~n34508;
  assign n34655 = ~n6563 & ~n16429;
  assign n34656 = n6576 & n34591;
  assign n34657 = n16429 & ~n34656;
  assign n34658 = ~n34654 & ~n34655;
  assign n34659 = ~n34657 & n34658;
  assign n34660 = n34468 & n34659;
  assign n34661 = pi201 & ~n34660;
  assign po358 = ~n34653 & ~n34661;
  assign n34663 = ~pi233 & pi237;
  assign n34664 = ~n34504 & ~n34663;
  assign n34665 = ~n34650 & n34663;
  assign n34666 = ~n34664 & ~n34665;
  assign n34667 = ~pi202 & ~n34666;
  assign n34668 = n34659 & n34663;
  assign n34669 = pi202 & ~n34668;
  assign po359 = ~n34667 & ~n34669;
  assign n34671 = ~pi233 & ~pi237;
  assign n34672 = ~n34504 & ~n34671;
  assign n34673 = ~n34650 & n34671;
  assign n34674 = ~n34672 & ~n34673;
  assign n34675 = ~pi203 & ~n34674;
  assign n34676 = n34659 & n34671;
  assign n34677 = pi203 & ~n34676;
  assign po360 = ~n34675 & ~n34677;
  assign n34679 = ~pi468 & pi602;
  assign n34680 = pi468 & n6168;
  assign n34681 = ~n34679 & ~n34680;
  assign n34682 = ~pi299 & ~n34681;
  assign n34683 = ~n6481 & ~n34682;
  assign n34684 = n3096 & ~n34683;
  assign n34685 = ~pi332 & ~n34684;
  assign n34686 = n15643 & ~n34685;
  assign n34687 = ~pi299 & ~pi602;
  assign n34688 = pi299 & ~pi907;
  assign n34689 = ~pi468 & ~n34687;
  assign n34690 = ~n34688 & n34689;
  assign n34691 = ~n34680 & ~n34690;
  assign n34692 = n34474 & ~n34691;
  assign n34693 = ~pi332 & ~n34692;
  assign n34694 = n7380 & ~n34693;
  assign n34695 = ~n34686 & ~n34694;
  assign n34696 = ~pi74 & ~n34695;
  assign n34697 = n34473 & ~n34486;
  assign n34698 = ~n34696 & n34697;
  assign n34699 = n3269 & n6299;
  assign n34700 = n3096 & n34699;
  assign n34701 = ~pi332 & ~n34700;
  assign n34702 = pi55 & n34701;
  assign n34703 = n3294 & ~n34702;
  assign n34704 = ~n34698 & n34703;
  assign n34705 = n34471 & ~n34704;
  assign n34706 = n6293 & ~n34701;
  assign n34707 = n34500 & ~n34706;
  assign n34708 = ~pi57 & ~n34707;
  assign n34709 = ~n34705 & n34708;
  assign n34710 = ~n34469 & ~n34709;
  assign n34711 = ~n34468 & ~n34710;
  assign n34712 = ~pi332 & ~n6168;
  assign n34713 = ~pi907 & ~n34712;
  assign n34714 = n6168 & ~n34520;
  assign n34715 = n34713 & ~n34714;
  assign n34716 = ~n6168 & n34525;
  assign n34717 = n6168 & ~n34519;
  assign n34718 = pi907 & ~n34717;
  assign n34719 = ~n34716 & n34718;
  assign n34720 = ~n34715 & ~n34719;
  assign n34721 = pi57 & ~n34720;
  assign n34722 = ~n3269 & n34720;
  assign n34723 = ~n6168 & n34551;
  assign n34724 = n6168 & ~n34546;
  assign n34725 = pi907 & ~n34724;
  assign n34726 = ~n34723 & n34725;
  assign n34727 = pi332 & ~n16708;
  assign n34728 = pi680 & ~n34727;
  assign n34729 = ~n34547 & n34728;
  assign n34730 = n34713 & ~n34729;
  assign n34731 = ~n34726 & ~n34730;
  assign n34732 = n3269 & n34731;
  assign n34733 = ~n34722 & ~n34732;
  assign n34734 = n6293 & ~n34733;
  assign n34735 = ~n6293 & n34720;
  assign n34736 = pi59 & ~n34735;
  assign n34737 = ~n34734 & n34736;
  assign n34738 = pi299 & n34731;
  assign n34739 = n6168 & n34591;
  assign n34740 = pi332 & ~n34739;
  assign n34741 = ~pi299 & ~n34740;
  assign n34742 = n6412 & n34612;
  assign n34743 = n34741 & ~n34742;
  assign n34744 = ~n34738 & ~n34743;
  assign n34745 = n15643 & ~n34744;
  assign n34746 = n6412 & n34593;
  assign n34747 = n34741 & ~n34746;
  assign n34748 = n6168 & ~n34575;
  assign n34749 = n34713 & ~n34748;
  assign n34750 = ~n6168 & n34579;
  assign n34751 = n6168 & ~n34574;
  assign n34752 = pi907 & ~n34751;
  assign n34753 = ~n34750 & n34752;
  assign n34754 = pi299 & ~n34749;
  assign n34755 = ~n34753 & n34754;
  assign n34756 = ~n34747 & ~n34755;
  assign n34757 = n7380 & ~n34756;
  assign n34758 = ~n34745 & ~n34757;
  assign n34759 = ~pi74 & ~n34758;
  assign n34760 = pi299 & ~n34720;
  assign n34761 = n34631 & ~n34681;
  assign n34762 = ~n34740 & ~n34761;
  assign n34763 = ~pi299 & ~n34762;
  assign n34764 = ~n34628 & ~n34763;
  assign n34765 = ~n34760 & n34764;
  assign n34766 = ~pi55 & ~n34765;
  assign n34767 = ~n34759 & n34766;
  assign n34768 = pi55 & n34733;
  assign n34769 = n3294 & ~n34768;
  assign n34770 = ~n34767 & n34769;
  assign n34771 = ~n3294 & n34720;
  assign n34772 = ~pi59 & ~n34771;
  assign n34773 = ~n34770 & n34772;
  assign n34774 = ~n34737 & ~n34773;
  assign n34775 = ~pi57 & ~n34774;
  assign n34776 = ~n34721 & ~n34775;
  assign n34777 = n34468 & ~n34776;
  assign n34778 = ~n34711 & ~n34777;
  assign n34779 = ~pi204 & ~n34778;
  assign n34780 = n6412 & n34591;
  assign n34781 = n16429 & ~n34780;
  assign n34782 = ~n6299 & ~n16429;
  assign n34783 = ~n34654 & ~n34782;
  assign n34784 = ~n34781 & n34783;
  assign n34785 = n34468 & n34784;
  assign n34786 = pi204 & ~n34785;
  assign po361 = ~n34779 & ~n34786;
  assign n34788 = ~n34663 & ~n34710;
  assign n34789 = n34663 & ~n34776;
  assign n34790 = ~n34788 & ~n34789;
  assign n34791 = ~pi205 & ~n34790;
  assign n34792 = n34663 & n34784;
  assign n34793 = pi205 & ~n34792;
  assign po362 = ~n34791 & ~n34793;
  assign n34795 = pi233 & ~pi237;
  assign n34796 = ~n34710 & ~n34795;
  assign n34797 = ~n34776 & n34795;
  assign n34798 = ~n34796 & ~n34797;
  assign n34799 = ~pi206 & ~n34798;
  assign n34800 = n34784 & n34795;
  assign n34801 = pi206 & ~n34800;
  assign po363 = ~n34799 & ~n34801;
  assign n34803 = ~n19124 & n24309;
  assign n34804 = n19217 & n34803;
  assign n34805 = ~n19247 & n34804;
  assign n34806 = pi207 & ~n34805;
  assign n34807 = ~n17494 & n17627;
  assign n34808 = n3268 & n24312;
  assign n34809 = ~pi778 & ~n34808;
  assign n34810 = ~pi625 & ~n17494;
  assign n34811 = pi625 & ~n34808;
  assign n34812 = ~n34810 & ~n34811;
  assign n34813 = pi1153 & ~n34812;
  assign n34814 = pi625 & ~n17494;
  assign n34815 = ~pi625 & ~n34808;
  assign n34816 = ~n34814 & ~n34815;
  assign n34817 = ~pi1153 & ~n34816;
  assign n34818 = ~n34813 & ~n34817;
  assign n34819 = pi778 & ~n34818;
  assign n34820 = ~n34809 & ~n34819;
  assign n34821 = ~n17554 & ~n34820;
  assign n34822 = ~n17494 & n17554;
  assign n34823 = ~n34821 & ~n34822;
  assign n34824 = ~n17591 & n34823;
  assign n34825 = n17494 & n17591;
  assign n34826 = ~n34824 & ~n34825;
  assign n34827 = ~n17627 & n34826;
  assign n34828 = ~n34807 & ~n34827;
  assign n34829 = ~n17670 & n34828;
  assign n34830 = n17494 & n17670;
  assign n34831 = ~n34829 & ~n34830;
  assign n34832 = ~n19247 & ~n34831;
  assign n34833 = n17494 & n17946;
  assign n34834 = ~n34832 & ~n34833;
  assign n34835 = ~pi207 & ~n34834;
  assign n34836 = ~n34806 & ~n34835;
  assign n34837 = pi710 & ~n34836;
  assign n34838 = ~pi207 & ~n17494;
  assign n34839 = ~pi710 & ~n34838;
  assign n34840 = ~n34837 & ~n34839;
  assign n34841 = ~pi647 & n34840;
  assign n34842 = pi647 & n34838;
  assign n34843 = ~pi1157 & ~n34842;
  assign n34844 = ~n34841 & n34843;
  assign n34845 = pi630 & n34844;
  assign n34846 = pi647 & n34840;
  assign n34847 = ~pi647 & n34838;
  assign n34848 = pi1157 & ~n34847;
  assign n34849 = ~n34846 & n34848;
  assign n34850 = ~pi630 & n34849;
  assign n34851 = ~n17494 & n17526;
  assign n34852 = n3268 & n19349;
  assign n34853 = ~n17526 & ~n34852;
  assign n34854 = ~n34851 & ~n34853;
  assign n34855 = ~pi785 & ~n34854;
  assign n34856 = ~n17494 & ~n17539;
  assign n34857 = ~pi609 & n34853;
  assign n34858 = ~n34856 & ~n34857;
  assign n34859 = ~pi1155 & ~n34858;
  assign n34860 = ~n17494 & ~n17527;
  assign n34861 = pi609 & n34853;
  assign n34862 = ~n34860 & ~n34861;
  assign n34863 = pi1155 & ~n34862;
  assign n34864 = ~n34859 & ~n34863;
  assign n34865 = pi785 & ~n34864;
  assign n34866 = ~n34855 & ~n34865;
  assign n34867 = ~pi781 & ~n34866;
  assign n34868 = ~pi618 & n34866;
  assign n34869 = pi618 & n17494;
  assign n34870 = ~pi1154 & ~n34869;
  assign n34871 = ~n34868 & n34870;
  assign n34872 = pi618 & n34866;
  assign n34873 = ~pi618 & n17494;
  assign n34874 = pi1154 & ~n34873;
  assign n34875 = ~n34872 & n34874;
  assign n34876 = ~n34871 & ~n34875;
  assign n34877 = pi781 & ~n34876;
  assign n34878 = ~n34867 & ~n34877;
  assign n34879 = ~pi789 & ~n34878;
  assign n34880 = ~pi619 & n34878;
  assign n34881 = pi619 & n17494;
  assign n34882 = ~pi1159 & ~n34881;
  assign n34883 = ~n34880 & n34882;
  assign n34884 = pi619 & n34878;
  assign n34885 = ~pi619 & n17494;
  assign n34886 = pi1159 & ~n34885;
  assign n34887 = ~n34884 & n34886;
  assign n34888 = ~n34883 & ~n34887;
  assign n34889 = pi789 & ~n34888;
  assign n34890 = ~n34879 & ~n34889;
  assign n34891 = ~n17904 & n34890;
  assign n34892 = n17494 & n17904;
  assign n34893 = ~n34891 & ~n34892;
  assign n34894 = ~n17698 & ~n34893;
  assign n34895 = n17494 & n17698;
  assign n34896 = ~n34894 & ~n34895;
  assign n34897 = ~pi207 & ~n34896;
  assign n34898 = n3268 & ~n24371;
  assign n34899 = ~n17526 & n34898;
  assign n34900 = ~n20159 & n34899;
  assign n34901 = ~n20169 & n34900;
  assign n34902 = ~n20165 & n34901;
  assign n34903 = ~n17904 & n34902;
  assign n34904 = ~n17698 & n34903;
  assign n34905 = pi207 & ~n34904;
  assign n34906 = pi623 & ~n34905;
  assign n34907 = ~n34897 & n34906;
  assign n34908 = ~pi623 & n34838;
  assign n34909 = ~n34907 & ~n34908;
  assign n34910 = ~n20491 & n34909;
  assign n34911 = ~n34845 & ~n34850;
  assign n34912 = ~n34910 & n34911;
  assign n34913 = pi787 & ~n34912;
  assign n34914 = ~pi628 & ~n17494;
  assign n34915 = pi628 & n34831;
  assign n34916 = ~n34914 & ~n34915;
  assign n34917 = ~pi629 & ~n34916;
  assign n34918 = ~n34914 & ~n34917;
  assign n34919 = pi1156 & ~n34918;
  assign n34920 = pi628 & ~n17494;
  assign n34921 = ~pi1156 & n34920;
  assign n34922 = ~pi628 & n34831;
  assign n34923 = ~n34920 & ~n34922;
  assign n34924 = n17696 & ~n34923;
  assign n34925 = ~n34921 & ~n34924;
  assign n34926 = ~n34919 & n34925;
  assign n34927 = pi792 & ~n34926;
  assign n34928 = pi619 & n34826;
  assign n34929 = pi618 & ~n34823;
  assign n34930 = pi609 & ~n34820;
  assign n34931 = n3268 & ~n19309;
  assign n34932 = ~pi778 & ~n34931;
  assign n34933 = ~pi625 & ~n34931;
  assign n34934 = ~n34814 & ~n34933;
  assign n34935 = ~pi1153 & ~n34934;
  assign n34936 = ~pi608 & ~n34813;
  assign n34937 = ~n34935 & n34936;
  assign n34938 = pi625 & ~n34931;
  assign n34939 = ~n34810 & ~n34938;
  assign n34940 = pi1153 & ~n34939;
  assign n34941 = pi608 & ~n34817;
  assign n34942 = ~n34940 & n34941;
  assign n34943 = pi778 & ~n34937;
  assign n34944 = ~n34942 & n34943;
  assign n34945 = ~n34932 & ~n34944;
  assign n34946 = ~pi609 & ~n34945;
  assign n34947 = ~n34930 & ~n34946;
  assign n34948 = ~pi1155 & ~n34947;
  assign n34949 = pi1155 & ~n17494;
  assign n34950 = ~pi660 & ~n34949;
  assign n34951 = ~n34948 & n34950;
  assign n34952 = ~pi609 & ~n34820;
  assign n34953 = pi609 & ~n34945;
  assign n34954 = ~n34952 & ~n34953;
  assign n34955 = pi1155 & ~n34954;
  assign n34956 = ~pi1155 & ~n17494;
  assign n34957 = pi660 & ~n34956;
  assign n34958 = ~n34955 & n34957;
  assign n34959 = ~n34951 & ~n34958;
  assign n34960 = pi785 & ~n34959;
  assign n34961 = ~pi785 & n34945;
  assign n34962 = ~n34960 & ~n34961;
  assign n34963 = ~pi618 & n34962;
  assign n34964 = ~n34929 & ~n34963;
  assign n34965 = ~pi1154 & ~n34964;
  assign n34966 = pi1154 & ~n17494;
  assign n34967 = ~pi627 & ~n34966;
  assign n34968 = ~n34965 & n34967;
  assign n34969 = ~pi618 & ~n34823;
  assign n34970 = pi618 & n34962;
  assign n34971 = ~n34969 & ~n34970;
  assign n34972 = pi1154 & ~n34971;
  assign n34973 = ~pi1154 & ~n17494;
  assign n34974 = pi627 & ~n34973;
  assign n34975 = ~n34972 & n34974;
  assign n34976 = ~n34968 & ~n34975;
  assign n34977 = pi781 & ~n34976;
  assign n34978 = ~pi781 & ~n34962;
  assign n34979 = ~n34977 & ~n34978;
  assign n34980 = ~pi619 & n34979;
  assign n34981 = ~n34928 & ~n34980;
  assign n34982 = ~pi1159 & ~n34981;
  assign n34983 = pi1159 & ~n17494;
  assign n34984 = ~pi648 & ~n34983;
  assign n34985 = ~n34982 & n34984;
  assign n34986 = ~pi619 & n34826;
  assign n34987 = pi619 & n34979;
  assign n34988 = ~n34986 & ~n34987;
  assign n34989 = pi1159 & ~n34988;
  assign n34990 = ~pi1159 & ~n17494;
  assign n34991 = pi648 & ~n34990;
  assign n34992 = ~n34989 & n34991;
  assign n34993 = ~n34985 & ~n34992;
  assign n34994 = pi789 & ~n34993;
  assign n34995 = ~pi789 & ~n34979;
  assign n34996 = ~n34994 & ~n34995;
  assign n34997 = ~pi626 & ~n34996;
  assign n34998 = pi626 & n34828;
  assign n34999 = ~pi641 & ~n34998;
  assign n35000 = ~n34997 & n34999;
  assign n35001 = pi641 & ~n17494;
  assign n35002 = ~pi1158 & ~n35001;
  assign n35003 = ~n35000 & n35002;
  assign n35004 = pi626 & ~n34996;
  assign n35005 = ~pi626 & n34828;
  assign n35006 = pi641 & ~n35005;
  assign n35007 = ~n35004 & n35006;
  assign n35008 = ~pi641 & ~n17494;
  assign n35009 = pi1158 & ~n35008;
  assign n35010 = ~n35007 & n35009;
  assign n35011 = ~n35003 & ~n35010;
  assign n35012 = pi788 & ~n35011;
  assign n35013 = ~pi788 & ~n34996;
  assign n35014 = ~n20298 & ~n35013;
  assign n35015 = ~n35012 & n35014;
  assign n35016 = ~n34927 & ~n35015;
  assign n35017 = ~pi207 & ~n35016;
  assign n35018 = ~pi778 & ~n33915;
  assign n35019 = ~pi625 & n33915;
  assign n35020 = ~pi1153 & ~n35019;
  assign n35021 = pi625 & n24309;
  assign n35022 = pi1153 & ~n35021;
  assign n35023 = ~pi608 & ~n35022;
  assign n35024 = ~n35020 & n35023;
  assign n35025 = pi625 & n33915;
  assign n35026 = pi1153 & ~n35025;
  assign n35027 = ~pi625 & n24309;
  assign n35028 = ~pi1153 & ~n35027;
  assign n35029 = pi608 & ~n35028;
  assign n35030 = ~n35026 & n35029;
  assign n35031 = pi778 & ~n35024;
  assign n35032 = ~n35030 & n35031;
  assign n35033 = ~n35018 & ~n35032;
  assign n35034 = ~pi609 & ~n35033;
  assign n35035 = pi609 & ~n34803;
  assign n35036 = n17552 & ~n35035;
  assign n35037 = ~n35034 & n35036;
  assign n35038 = pi609 & ~n35033;
  assign n35039 = ~pi609 & ~n34803;
  assign n35040 = n17551 & ~n35039;
  assign n35041 = ~n35038 & n35040;
  assign n35042 = ~n35037 & ~n35041;
  assign n35043 = pi785 & ~n35042;
  assign n35044 = ~pi785 & n35033;
  assign n35045 = ~n35043 & ~n35044;
  assign n35046 = ~pi618 & n35045;
  assign n35047 = ~n17554 & n34803;
  assign n35048 = pi618 & ~n35047;
  assign n35049 = n17589 & ~n35048;
  assign n35050 = ~n35046 & n35049;
  assign n35051 = pi618 & n35045;
  assign n35052 = ~pi618 & ~n35047;
  assign n35053 = n17588 & ~n35052;
  assign n35054 = ~n35051 & n35053;
  assign n35055 = pi781 & ~n35050;
  assign n35056 = ~n35054 & n35055;
  assign n35057 = ~pi781 & n35045;
  assign n35058 = ~n23544 & ~n35057;
  assign n35059 = ~n35056 & n35058;
  assign n35060 = n19216 & n34803;
  assign n35061 = n17626 & n20165;
  assign n35062 = n35060 & n35061;
  assign n35063 = ~n35059 & ~n35062;
  assign n35064 = ~pi626 & n35063;
  assign n35065 = ~n17627 & n35060;
  assign n35066 = pi626 & ~n35065;
  assign n35067 = ~pi641 & ~n35066;
  assign n35068 = ~pi1158 & n35067;
  assign n35069 = ~n35064 & n35068;
  assign n35070 = pi626 & n35063;
  assign n35071 = ~pi626 & ~n35065;
  assign n35072 = pi641 & ~n35071;
  assign n35073 = pi1158 & n35072;
  assign n35074 = ~n35070 & n35073;
  assign n35075 = pi788 & ~n35069;
  assign n35076 = ~n35074 & n35075;
  assign n35077 = ~pi788 & n35063;
  assign n35078 = ~n20298 & ~n35077;
  assign n35079 = ~n35076 & n35078;
  assign n35080 = n17698 & n17945;
  assign n35081 = n34804 & n35080;
  assign n35082 = ~n35079 & ~n35081;
  assign n35083 = pi207 & ~n35082;
  assign n35084 = ~pi623 & ~n35083;
  assign n35085 = ~n35017 & n35084;
  assign n35086 = n3268 & n19334;
  assign n35087 = ~pi778 & ~n35086;
  assign n35088 = ~pi625 & n34852;
  assign n35089 = pi625 & n35086;
  assign n35090 = pi1153 & ~n35089;
  assign n35091 = ~n35088 & n35090;
  assign n35092 = n34941 & ~n35091;
  assign n35093 = pi625 & n34852;
  assign n35094 = ~pi625 & n35086;
  assign n35095 = ~pi1153 & ~n35094;
  assign n35096 = ~n35093 & n35095;
  assign n35097 = n34936 & ~n35096;
  assign n35098 = pi778 & ~n35092;
  assign n35099 = ~n35097 & n35098;
  assign n35100 = ~n35087 & ~n35099;
  assign n35101 = ~pi609 & ~n35100;
  assign n35102 = ~n34930 & ~n35101;
  assign n35103 = ~pi1155 & ~n35102;
  assign n35104 = ~pi660 & ~n34863;
  assign n35105 = ~n35103 & n35104;
  assign n35106 = pi609 & ~n35100;
  assign n35107 = ~n34952 & ~n35106;
  assign n35108 = pi1155 & ~n35107;
  assign n35109 = pi660 & ~n34859;
  assign n35110 = ~n35108 & n35109;
  assign n35111 = ~n35105 & ~n35110;
  assign n35112 = pi785 & ~n35111;
  assign n35113 = ~pi785 & n35100;
  assign n35114 = ~n35112 & ~n35113;
  assign n35115 = ~pi618 & n35114;
  assign n35116 = ~n34929 & ~n35115;
  assign n35117 = ~pi1154 & ~n35116;
  assign n35118 = ~pi627 & ~n34875;
  assign n35119 = ~n35117 & n35118;
  assign n35120 = pi618 & n35114;
  assign n35121 = ~n34969 & ~n35120;
  assign n35122 = pi1154 & ~n35121;
  assign n35123 = pi627 & ~n34871;
  assign n35124 = ~n35122 & n35123;
  assign n35125 = ~n35119 & ~n35124;
  assign n35126 = pi781 & ~n35125;
  assign n35127 = ~pi781 & ~n35114;
  assign n35128 = ~n35126 & ~n35127;
  assign n35129 = ~pi619 & n35128;
  assign n35130 = ~n34928 & ~n35129;
  assign n35131 = ~pi1159 & ~n35130;
  assign n35132 = ~pi648 & ~n34887;
  assign n35133 = ~n35131 & n35132;
  assign n35134 = pi619 & n35128;
  assign n35135 = ~n34986 & ~n35134;
  assign n35136 = pi1159 & ~n35135;
  assign n35137 = pi648 & ~n34883;
  assign n35138 = ~n35136 & n35137;
  assign n35139 = pi789 & ~n35133;
  assign n35140 = ~n35138 & n35139;
  assign n35141 = ~pi789 & n35128;
  assign n35142 = n17905 & ~n35141;
  assign n35143 = ~n35140 & n35142;
  assign n35144 = ~n17669 & ~n17791;
  assign n35145 = n34890 & n35144;
  assign n35146 = pi641 & ~n34828;
  assign n35147 = n17786 & ~n35008;
  assign n35148 = ~n35146 & n35147;
  assign n35149 = ~pi641 & ~n34828;
  assign n35150 = n17787 & ~n35001;
  assign n35151 = ~n35149 & n35150;
  assign n35152 = ~n35148 & ~n35151;
  assign n35153 = ~n35145 & n35152;
  assign n35154 = pi788 & ~n35153;
  assign n35155 = ~n20298 & ~n35154;
  assign n35156 = ~n35143 & n35155;
  assign n35157 = ~n20502 & n34893;
  assign n35158 = pi1156 & n34917;
  assign n35159 = ~n34924 & ~n35157;
  assign n35160 = ~n35158 & n35159;
  assign n35161 = pi792 & ~n35160;
  assign n35162 = ~n35156 & ~n35161;
  assign n35163 = ~pi207 & ~n35162;
  assign n35164 = pi1156 & ~n34903;
  assign n35165 = ~pi1156 & ~n34804;
  assign n35166 = n20498 & ~n35165;
  assign n35167 = ~n35164 & n35166;
  assign n35168 = ~pi1156 & ~n34903;
  assign n35169 = pi1156 & ~n34804;
  assign n35170 = n20500 & ~n35169;
  assign n35171 = ~n35168 & n35170;
  assign n35172 = ~n35167 & ~n35171;
  assign n35173 = pi792 & ~n35172;
  assign n35174 = ~pi1159 & ~n34901;
  assign n35175 = pi1159 & ~n35060;
  assign n35176 = ~pi619 & pi648;
  assign n35177 = ~n35174 & n35176;
  assign n35178 = ~n35175 & n35177;
  assign n35179 = pi1159 & ~n34901;
  assign n35180 = ~pi1159 & ~n35060;
  assign n35181 = pi619 & ~pi648;
  assign n35182 = ~n35179 & n35181;
  assign n35183 = ~n35180 & n35182;
  assign n35184 = pi789 & ~n35178;
  assign n35185 = ~n35183 & n35184;
  assign n35186 = pi789 & ~n35185;
  assign n35187 = ~pi1154 & ~n35048;
  assign n35188 = n20167 & n34900;
  assign n35189 = ~pi627 & ~n35188;
  assign n35190 = ~n35187 & n35189;
  assign n35191 = ~pi778 & ~n33920;
  assign n35192 = ~pi625 & n33920;
  assign n35193 = pi625 & n34898;
  assign n35194 = ~pi1153 & ~n35193;
  assign n35195 = ~n35192 & n35194;
  assign n35196 = n35023 & ~n35195;
  assign n35197 = pi625 & n33920;
  assign n35198 = ~pi625 & n34898;
  assign n35199 = pi1153 & ~n35198;
  assign n35200 = ~n35197 & n35199;
  assign n35201 = n35029 & ~n35200;
  assign n35202 = pi778 & ~n35196;
  assign n35203 = ~n35201 & n35202;
  assign n35204 = ~n35191 & ~n35203;
  assign n35205 = ~pi785 & ~n35204;
  assign n35206 = ~pi609 & ~n35204;
  assign n35207 = ~pi1155 & ~n35035;
  assign n35208 = ~n35206 & n35207;
  assign n35209 = n20157 & n34899;
  assign n35210 = ~pi660 & ~n35209;
  assign n35211 = ~n35208 & n35210;
  assign n35212 = pi609 & ~n35204;
  assign n35213 = pi1155 & ~n35039;
  assign n35214 = ~n35212 & n35213;
  assign n35215 = n20156 & n34899;
  assign n35216 = pi660 & ~n35215;
  assign n35217 = ~n35214 & n35216;
  assign n35218 = ~n35211 & ~n35217;
  assign n35219 = pi785 & ~n35218;
  assign n35220 = ~n35205 & ~n35219;
  assign n35221 = pi618 & ~n35220;
  assign n35222 = pi1154 & ~n35052;
  assign n35223 = ~n35221 & n35222;
  assign n35224 = n20166 & n34900;
  assign n35225 = pi627 & ~n35224;
  assign n35226 = ~n35223 & n35225;
  assign n35227 = ~n35190 & ~n35226;
  assign n35228 = pi781 & ~n35227;
  assign n35229 = ~pi618 & ~pi627;
  assign n35230 = pi781 & ~n35229;
  assign n35231 = ~n35220 & ~n35230;
  assign n35232 = ~n23543 & n35185;
  assign n35233 = ~n35231 & ~n35232;
  assign n35234 = ~n35228 & n35233;
  assign n35235 = ~n35186 & ~n35234;
  assign n35236 = ~pi626 & n35235;
  assign n35237 = n35067 & ~n35236;
  assign n35238 = n17789 & n34902;
  assign n35239 = ~pi1158 & ~n35238;
  assign n35240 = ~n35237 & n35239;
  assign n35241 = pi626 & n35235;
  assign n35242 = n35072 & ~n35241;
  assign n35243 = n17790 & n34902;
  assign n35244 = pi1158 & ~n35243;
  assign n35245 = ~n35242 & n35244;
  assign n35246 = ~n35240 & ~n35245;
  assign n35247 = pi788 & ~n35246;
  assign n35248 = ~pi788 & n35235;
  assign n35249 = ~n20298 & ~n35248;
  assign n35250 = ~n35247 & n35249;
  assign n35251 = ~n35173 & ~n35250;
  assign n35252 = pi207 & ~n35251;
  assign n35253 = pi623 & ~n35252;
  assign n35254 = ~n35163 & n35253;
  assign n35255 = pi710 & ~n35254;
  assign n35256 = ~n35085 & n35255;
  assign n35257 = ~pi710 & ~n34909;
  assign n35258 = n20300 & ~n35257;
  assign n35259 = ~n35256 & n35258;
  assign n35260 = ~n34913 & ~n35259;
  assign n35261 = pi644 & n35260;
  assign n35262 = ~pi787 & ~n34840;
  assign n35263 = ~n34844 & ~n34849;
  assign n35264 = pi787 & ~n35263;
  assign n35265 = ~n35262 & ~n35264;
  assign n35266 = ~pi644 & n35265;
  assign n35267 = pi715 & ~n35266;
  assign n35268 = ~n35261 & n35267;
  assign n35269 = n17740 & ~n34838;
  assign n35270 = ~n17740 & n34909;
  assign n35271 = ~n35269 & ~n35270;
  assign n35272 = pi644 & n35271;
  assign n35273 = ~pi644 & n34838;
  assign n35274 = ~pi715 & ~n35273;
  assign n35275 = ~n35272 & n35274;
  assign n35276 = pi1160 & ~n35275;
  assign n35277 = ~n35268 & n35276;
  assign n35278 = ~pi644 & n35260;
  assign n35279 = pi644 & n35265;
  assign n35280 = ~pi715 & ~n35279;
  assign n35281 = ~n35278 & n35280;
  assign n35282 = ~pi644 & n35271;
  assign n35283 = pi644 & n34838;
  assign n35284 = pi715 & ~n35283;
  assign n35285 = ~n35282 & n35284;
  assign n35286 = ~pi1160 & ~n35285;
  assign n35287 = ~n35281 & n35286;
  assign n35288 = ~n35277 & ~n35287;
  assign n35289 = pi790 & ~n35288;
  assign n35290 = ~pi790 & n35260;
  assign n35291 = ~n35289 & ~n35290;
  assign n35292 = ~po1038 & ~n35291;
  assign n35293 = ~pi207 & po1038;
  assign po364 = n35292 | n35293;
  assign n35295 = pi208 & ~n34805;
  assign n35296 = ~pi208 & ~n34834;
  assign n35297 = ~n35295 & ~n35296;
  assign n35298 = pi638 & ~n35297;
  assign n35299 = ~pi208 & ~n17494;
  assign n35300 = ~pi638 & ~n35299;
  assign n35301 = ~n35298 & ~n35300;
  assign n35302 = ~pi647 & n35301;
  assign n35303 = pi647 & n35299;
  assign n35304 = ~pi1157 & ~n35303;
  assign n35305 = ~n35302 & n35304;
  assign n35306 = pi630 & n35305;
  assign n35307 = pi647 & n35301;
  assign n35308 = ~pi647 & n35299;
  assign n35309 = pi1157 & ~n35308;
  assign n35310 = ~n35307 & n35309;
  assign n35311 = ~pi630 & n35310;
  assign n35312 = ~pi208 & ~n34896;
  assign n35313 = pi208 & ~n34904;
  assign n35314 = pi607 & ~n35313;
  assign n35315 = ~n35312 & n35314;
  assign n35316 = ~pi607 & n35299;
  assign n35317 = ~n35315 & ~n35316;
  assign n35318 = ~n20491 & n35317;
  assign n35319 = ~n35306 & ~n35311;
  assign n35320 = ~n35318 & n35319;
  assign n35321 = pi787 & ~n35320;
  assign n35322 = ~pi208 & ~n35016;
  assign n35323 = pi208 & ~n35082;
  assign n35324 = ~pi607 & ~n35323;
  assign n35325 = ~n35322 & n35324;
  assign n35326 = ~pi208 & ~n35162;
  assign n35327 = pi208 & ~n35251;
  assign n35328 = pi607 & ~n35327;
  assign n35329 = ~n35326 & n35328;
  assign n35330 = pi638 & ~n35329;
  assign n35331 = ~n35325 & n35330;
  assign n35332 = ~pi638 & ~n35317;
  assign n35333 = n20300 & ~n35332;
  assign n35334 = ~n35331 & n35333;
  assign n35335 = ~n35321 & ~n35334;
  assign n35336 = pi644 & n35335;
  assign n35337 = ~pi787 & ~n35301;
  assign n35338 = ~n35305 & ~n35310;
  assign n35339 = pi787 & ~n35338;
  assign n35340 = ~n35337 & ~n35339;
  assign n35341 = ~pi644 & n35340;
  assign n35342 = pi715 & ~n35341;
  assign n35343 = ~n35336 & n35342;
  assign n35344 = n17740 & ~n35299;
  assign n35345 = ~n17740 & n35317;
  assign n35346 = ~n35344 & ~n35345;
  assign n35347 = pi644 & n35346;
  assign n35348 = ~pi644 & n35299;
  assign n35349 = ~pi715 & ~n35348;
  assign n35350 = ~n35347 & n35349;
  assign n35351 = pi1160 & ~n35350;
  assign n35352 = ~n35343 & n35351;
  assign n35353 = ~pi644 & n35335;
  assign n35354 = pi644 & n35340;
  assign n35355 = ~pi715 & ~n35354;
  assign n35356 = ~n35353 & n35355;
  assign n35357 = ~pi644 & n35346;
  assign n35358 = pi644 & n35299;
  assign n35359 = pi715 & ~n35358;
  assign n35360 = ~n35357 & n35359;
  assign n35361 = ~pi1160 & ~n35360;
  assign n35362 = ~n35356 & n35361;
  assign n35363 = ~n35352 & ~n35362;
  assign n35364 = pi790 & ~n35363;
  assign n35365 = ~pi790 & n35335;
  assign n35366 = ~n35364 & ~n35365;
  assign n35367 = ~po1038 & ~n35366;
  assign n35368 = ~pi208 & po1038;
  assign po365 = n35367 | n35368;
  assign n35370 = n20300 & ~n35016;
  assign n35371 = ~pi647 & ~n17494;
  assign n35372 = pi647 & n34834;
  assign n35373 = ~n35371 & ~n35372;
  assign n35374 = ~pi630 & ~n35373;
  assign n35375 = ~n35371 & ~n35374;
  assign n35376 = pi1157 & ~n35375;
  assign n35377 = pi647 & ~n17494;
  assign n35378 = ~pi1157 & n35377;
  assign n35379 = ~pi647 & n34834;
  assign n35380 = ~n35377 & ~n35379;
  assign n35381 = n17738 & ~n35380;
  assign n35382 = ~n35378 & ~n35381;
  assign n35383 = ~n35376 & n35382;
  assign n35384 = pi787 & ~n35383;
  assign n35385 = ~n35370 & ~n35384;
  assign n35386 = ~pi644 & ~n35385;
  assign n35387 = ~n19271 & n34834;
  assign n35388 = ~n17494 & n19271;
  assign n35389 = ~n35387 & ~n35388;
  assign n35390 = pi644 & ~n35389;
  assign n35391 = ~pi715 & ~n35390;
  assign n35392 = ~n35386 & n35391;
  assign n35393 = pi715 & n17494;
  assign n35394 = ~pi1160 & ~n35393;
  assign n35395 = ~n35392 & n35394;
  assign n35396 = pi644 & ~n35385;
  assign n35397 = ~pi644 & ~n35389;
  assign n35398 = pi715 & ~n35397;
  assign n35399 = ~n35396 & n35398;
  assign n35400 = ~pi715 & n17494;
  assign n35401 = pi1160 & ~n35400;
  assign n35402 = ~n35399 & n35401;
  assign n35403 = ~n35395 & ~n35402;
  assign n35404 = pi790 & ~n35403;
  assign n35405 = ~pi790 & ~n35385;
  assign n35406 = ~po1038 & ~n35405;
  assign n35407 = ~n35404 & n35406;
  assign n35408 = pi639 & n35407;
  assign n35409 = n10178 & n17487;
  assign n35410 = ~pi639 & n35409;
  assign n35411 = ~pi622 & ~n35410;
  assign n35412 = ~n35408 & n35411;
  assign n35413 = n20300 & ~n35162;
  assign n35414 = ~n20491 & n34896;
  assign n35415 = ~n17739 & ~n35383;
  assign n35416 = ~n35414 & ~n35415;
  assign n35417 = pi787 & ~n35416;
  assign n35418 = ~n35413 & ~n35417;
  assign n35419 = ~pi644 & ~n35418;
  assign n35420 = n35391 & ~n35419;
  assign n35421 = ~n17494 & n17740;
  assign n35422 = ~n17740 & n34896;
  assign n35423 = ~n35421 & ~n35422;
  assign n35424 = ~pi644 & ~n35423;
  assign n35425 = pi644 & ~n17494;
  assign n35426 = ~n35424 & ~n35425;
  assign n35427 = pi715 & n35426;
  assign n35428 = ~pi1160 & ~n35427;
  assign n35429 = ~n35420 & n35428;
  assign n35430 = pi644 & ~n35418;
  assign n35431 = n35398 & ~n35430;
  assign n35432 = pi644 & ~n35423;
  assign n35433 = ~pi644 & ~n17494;
  assign n35434 = ~n35432 & ~n35433;
  assign n35435 = ~pi715 & n35434;
  assign n35436 = pi1160 & ~n35435;
  assign n35437 = ~n35431 & n35436;
  assign n35438 = ~n35429 & ~n35437;
  assign n35439 = pi790 & ~n35438;
  assign n35440 = ~pi790 & ~n35418;
  assign n35441 = ~po1038 & ~n35440;
  assign n35442 = ~n35439 & n35441;
  assign n35443 = pi639 & n35442;
  assign n35444 = pi1160 & n35434;
  assign n35445 = ~pi1160 & n35426;
  assign n35446 = pi790 & ~n35444;
  assign n35447 = ~n35445 & n35446;
  assign n35448 = ~pi790 & ~n35423;
  assign n35449 = ~po1038 & ~n35448;
  assign n35450 = ~n35447 & n35449;
  assign n35451 = ~pi639 & n35450;
  assign n35452 = pi622 & ~n35451;
  assign n35453 = ~n35443 & n35452;
  assign n35454 = ~n35412 & ~n35453;
  assign n35455 = ~pi209 & ~n35454;
  assign n35456 = ~n19271 & n34805;
  assign n35457 = pi644 & ~n35456;
  assign n35458 = ~pi715 & ~n35457;
  assign n35459 = ~pi647 & ~n35251;
  assign n35460 = pi647 & n34904;
  assign n35461 = ~pi1157 & ~n35460;
  assign n35462 = ~n35459 & n35461;
  assign n35463 = pi647 & n34805;
  assign n35464 = pi1157 & ~n35463;
  assign n35465 = ~pi630 & ~n35464;
  assign n35466 = ~n35462 & n35465;
  assign n35467 = pi647 & ~n35251;
  assign n35468 = ~pi647 & n34904;
  assign n35469 = pi1157 & ~n35468;
  assign n35470 = ~n35467 & n35469;
  assign n35471 = ~pi647 & n34805;
  assign n35472 = ~pi1157 & ~n35471;
  assign n35473 = pi630 & ~n35472;
  assign n35474 = ~n35470 & n35473;
  assign n35475 = ~n35466 & ~n35474;
  assign n35476 = pi787 & ~n35475;
  assign n35477 = ~pi787 & ~n35251;
  assign n35478 = ~n35476 & ~n35477;
  assign n35479 = ~pi644 & n35478;
  assign n35480 = n35458 & ~n35479;
  assign n35481 = n23618 & n34903;
  assign n35482 = ~pi644 & pi715;
  assign n35483 = n35481 & n35482;
  assign n35484 = ~pi1160 & ~n35483;
  assign n35485 = ~n35480 & n35484;
  assign n35486 = ~pi644 & ~n35456;
  assign n35487 = pi715 & ~n35486;
  assign n35488 = pi644 & n35478;
  assign n35489 = n35487 & ~n35488;
  assign n35490 = pi644 & ~pi715;
  assign n35491 = n35481 & n35490;
  assign n35492 = pi1160 & ~n35491;
  assign n35493 = ~n35489 & n35492;
  assign n35494 = ~n35485 & ~n35493;
  assign n35495 = pi790 & ~n35494;
  assign n35496 = ~pi790 & n35478;
  assign n35497 = ~po1038 & ~n35496;
  assign n35498 = ~n35495 & n35497;
  assign n35499 = pi622 & pi639;
  assign n35500 = ~n35498 & n35499;
  assign n35501 = n20300 & ~n35082;
  assign n35502 = n17740 & n19270;
  assign n35503 = n34805 & n35502;
  assign n35504 = ~n35501 & ~n35503;
  assign n35505 = pi644 & n35504;
  assign n35506 = pi1160 & n35487;
  assign n35507 = ~n35505 & n35506;
  assign n35508 = ~pi644 & n35504;
  assign n35509 = ~pi1160 & n35458;
  assign n35510 = ~n35508 & n35509;
  assign n35511 = pi790 & ~n35507;
  assign n35512 = ~n35510 & n35511;
  assign n35513 = ~pi790 & n35504;
  assign n35514 = ~po1038 & ~n35513;
  assign n35515 = ~n35512 & n35514;
  assign n35516 = ~pi622 & ~n35515;
  assign n35517 = ~pi644 & pi1160;
  assign n35518 = pi644 & ~pi1160;
  assign n35519 = ~n35517 & ~n35518;
  assign n35520 = pi790 & ~n35519;
  assign n35521 = ~po1038 & ~n35520;
  assign n35522 = n35481 & n35521;
  assign n35523 = pi622 & n35522;
  assign n35524 = ~pi639 & ~n35523;
  assign n35525 = pi209 & ~n35524;
  assign n35526 = ~n35516 & n35525;
  assign n35527 = ~n35500 & n35526;
  assign po366 = n35455 | n35527;
  assign n35529 = pi210 & ~n16968;
  assign n35530 = pi634 & n20848;
  assign n35531 = pi633 & pi947;
  assign n35532 = ~n35530 & ~n35531;
  assign n35533 = n16968 & ~n35532;
  assign n35534 = pi38 & ~n35529;
  assign n35535 = ~n35533 & n35534;
  assign n35536 = pi210 & ~n16661;
  assign n35537 = ~po1101 & n35536;
  assign n35538 = pi210 & po1101;
  assign n35539 = ~n16750 & n35538;
  assign n35540 = ~n35537 & ~n35539;
  assign n35541 = ~pi907 & n35540;
  assign n35542 = pi634 & n16661;
  assign n35543 = ~n35536 & ~n35542;
  assign n35544 = ~n6206 & ~n35543;
  assign n35545 = pi907 & ~n35544;
  assign n35546 = pi210 & n16748;
  assign n35547 = pi634 & ~n16748;
  assign n35548 = ~n35546 & ~n35547;
  assign n35549 = n6206 & ~n35548;
  assign n35550 = n35545 & ~n35549;
  assign n35551 = ~pi947 & ~n35550;
  assign n35552 = ~n35541 & n35551;
  assign n35553 = ~n33326 & ~n35536;
  assign n35554 = ~po1101 & n35553;
  assign n35555 = pi947 & ~n35554;
  assign n35556 = po1101 & n35553;
  assign n35557 = ~n6206 & ~n35556;
  assign n35558 = pi633 & ~n16748;
  assign n35559 = ~n35546 & ~n35558;
  assign n35560 = ~n6170 & ~n35559;
  assign n35561 = ~n35557 & ~n35560;
  assign n35562 = n35555 & ~n35561;
  assign n35563 = n6197 & ~n35562;
  assign n35564 = ~n35552 & n35563;
  assign n35565 = n6200 & n35543;
  assign n35566 = pi907 & ~n35565;
  assign n35567 = ~n6200 & n35548;
  assign n35568 = n35566 & ~n35567;
  assign n35569 = pi210 & ~n16785;
  assign n35570 = ~pi907 & n35569;
  assign n35571 = ~n35568 & ~n35570;
  assign n35572 = ~pi947 & ~n35571;
  assign n35573 = n6200 & n35553;
  assign n35574 = pi947 & ~n35573;
  assign n35575 = ~n6200 & n35559;
  assign n35576 = n35574 & ~n35575;
  assign n35577 = ~n6197 & ~n35576;
  assign n35578 = ~n35572 & n35577;
  assign n35579 = ~n35564 & ~n35578;
  assign n35580 = ~n3053 & ~n35579;
  assign n35581 = n16661 & ~n35532;
  assign n35582 = ~n35536 & ~n35581;
  assign n35583 = n3053 & n35582;
  assign n35584 = ~pi223 & ~n35583;
  assign n35585 = ~n35580 & n35584;
  assign n35586 = pi210 & n16677;
  assign n35587 = ~n33511 & ~n35586;
  assign n35588 = ~n6200 & n35587;
  assign n35589 = n35566 & ~n35588;
  assign n35590 = n6200 & n16660;
  assign n35591 = n2755 & n35590;
  assign n35592 = n35586 & ~n35591;
  assign n35593 = ~n35589 & ~n35592;
  assign n35594 = ~pi947 & ~n35593;
  assign n35595 = pi633 & ~n16677;
  assign n35596 = ~n35586 & ~n35595;
  assign n35597 = ~n6200 & n35596;
  assign n35598 = n35574 & ~n35597;
  assign n35599 = ~n6197 & ~n35598;
  assign n35600 = ~n35594 & n35599;
  assign n35601 = ~n16683 & n35538;
  assign n35602 = ~n35537 & ~n35601;
  assign n35603 = ~pi907 & n35602;
  assign n35604 = n6206 & ~n35587;
  assign n35605 = n35545 & ~n35604;
  assign n35606 = ~pi947 & ~n35605;
  assign n35607 = ~n35603 & n35606;
  assign n35608 = ~n6170 & ~n35596;
  assign n35609 = ~n35557 & ~n35608;
  assign n35610 = n35555 & ~n35609;
  assign n35611 = n6197 & ~n35610;
  assign n35612 = ~n35607 & n35611;
  assign n35613 = pi223 & ~n35600;
  assign n35614 = ~n35612 & n35613;
  assign n35615 = ~pi299 & ~n35614;
  assign n35616 = ~n35585 & n35615;
  assign n35617 = ~n6222 & ~n35569;
  assign n35618 = n6222 & n35540;
  assign n35619 = ~pi907 & ~n35618;
  assign n35620 = ~n35617 & n35619;
  assign n35621 = ~n35568 & ~n35620;
  assign n35622 = ~pi947 & ~n35621;
  assign n35623 = ~n3461 & ~n35576;
  assign n35624 = ~n35622 & n35623;
  assign n35625 = n3461 & n35582;
  assign n35626 = ~pi215 & ~n35625;
  assign n35627 = ~n35624 & n35626;
  assign n35628 = n6222 & n35602;
  assign n35629 = ~n6222 & ~n35592;
  assign n35630 = ~pi907 & ~n35629;
  assign n35631 = ~n35628 & n35630;
  assign n35632 = ~n35589 & ~n35631;
  assign n35633 = ~pi947 & ~n35632;
  assign n35634 = ~n35598 & ~n35633;
  assign n35635 = pi215 & ~n35634;
  assign n35636 = pi299 & ~n35635;
  assign n35637 = ~n35627 & n35636;
  assign n35638 = pi39 & ~n35637;
  assign n35639 = ~n35616 & n35638;
  assign n35640 = pi210 & ~n16653;
  assign n35641 = n16653 & ~n35532;
  assign n35642 = ~pi299 & ~n35640;
  assign n35643 = ~n35641 & n35642;
  assign n35644 = ~n16629 & ~n35532;
  assign n35645 = pi299 & ~n35644;
  assign n35646 = ~n16648 & n35645;
  assign n35647 = ~pi39 & ~n35646;
  assign n35648 = ~n35643 & n35647;
  assign n35649 = ~pi38 & ~n35648;
  assign n35650 = ~n35639 & n35649;
  assign n35651 = ~n35535 & ~n35650;
  assign n35652 = n10178 & ~n35651;
  assign n35653 = ~pi210 & ~n10178;
  assign po367 = ~n35652 & ~n35653;
  assign n35655 = n3268 & ~n21573;
  assign n35656 = ~pi606 & n35655;
  assign n35657 = n3268 & ~n21569;
  assign n35658 = pi606 & n35657;
  assign n35659 = pi643 & ~n35656;
  assign n35660 = ~n35658 & n35659;
  assign n35661 = n3268 & ~n20942;
  assign n35662 = pi606 & n35661;
  assign n35663 = ~pi606 & n17494;
  assign n35664 = ~pi643 & ~n35663;
  assign n35665 = ~n35662 & n35664;
  assign n35666 = ~po1038 & ~n35665;
  assign n35667 = ~n35660 & n35666;
  assign n35668 = pi211 & ~n35667;
  assign n35669 = n3268 & n21558;
  assign n35670 = ~pi606 & ~n35669;
  assign n35671 = n3268 & n21555;
  assign n35672 = pi606 & ~n35671;
  assign n35673 = pi643 & ~n35670;
  assign n35674 = ~n35672 & n35673;
  assign n35675 = n3268 & n20966;
  assign n35676 = pi606 & ~pi643;
  assign n35677 = n35675 & n35676;
  assign n35678 = ~n35674 & ~n35677;
  assign n35679 = ~pi211 & ~po1038;
  assign n35680 = ~n35678 & n35679;
  assign po368 = n35668 | n35680;
  assign n35682 = ~pi607 & n35655;
  assign n35683 = pi607 & n35657;
  assign n35684 = pi638 & ~n35682;
  assign n35685 = ~n35683 & n35684;
  assign n35686 = pi607 & n35661;
  assign n35687 = ~pi607 & n17494;
  assign n35688 = ~pi638 & ~n35687;
  assign n35689 = ~n35686 & n35688;
  assign n35690 = ~po1038 & ~n35689;
  assign n35691 = ~n35685 & n35690;
  assign n35692 = ~pi212 & ~n35691;
  assign n35693 = pi607 & ~n35671;
  assign n35694 = ~pi607 & ~n35669;
  assign n35695 = pi638 & ~n35693;
  assign n35696 = ~n35694 & n35695;
  assign n35697 = pi607 & ~pi638;
  assign n35698 = n35675 & n35697;
  assign n35699 = ~n35696 & ~n35698;
  assign n35700 = pi212 & ~po1038;
  assign n35701 = ~n35699 & n35700;
  assign po369 = n35692 | n35701;
  assign n35703 = pi213 & ~po1038;
  assign n35704 = pi622 & ~n35671;
  assign n35705 = ~pi622 & ~n35669;
  assign n35706 = pi639 & ~n35704;
  assign n35707 = ~n35705 & n35706;
  assign n35708 = pi622 & ~pi639;
  assign n35709 = n35675 & n35708;
  assign n35710 = ~n35707 & ~n35709;
  assign n35711 = n35703 & ~n35710;
  assign n35712 = ~pi639 & n35661;
  assign n35713 = pi639 & n35657;
  assign n35714 = pi622 & ~n35712;
  assign n35715 = ~n35713 & n35714;
  assign n35716 = pi639 & n35655;
  assign n35717 = ~pi639 & n17494;
  assign n35718 = ~pi622 & ~n35717;
  assign n35719 = ~n35716 & n35718;
  assign n35720 = ~po1038 & ~n35719;
  assign n35721 = ~n35715 & n35720;
  assign n35722 = ~pi213 & ~n35721;
  assign po370 = n35711 | n35722;
  assign n35724 = ~pi623 & n35655;
  assign n35725 = pi623 & n35657;
  assign n35726 = pi710 & ~n35724;
  assign n35727 = ~n35725 & n35726;
  assign n35728 = pi623 & n35661;
  assign n35729 = ~pi623 & n17494;
  assign n35730 = ~pi710 & ~n35729;
  assign n35731 = ~n35728 & n35730;
  assign n35732 = ~po1038 & ~n35731;
  assign n35733 = ~n35727 & n35732;
  assign n35734 = ~pi214 & ~n35733;
  assign n35735 = pi623 & ~n35671;
  assign n35736 = ~pi623 & ~n35669;
  assign n35737 = pi710 & ~n35735;
  assign n35738 = ~n35736 & n35737;
  assign n35739 = pi623 & ~pi710;
  assign n35740 = n35675 & n35739;
  assign n35741 = ~n35738 & ~n35740;
  assign n35742 = pi214 & ~po1038;
  assign n35743 = ~n35741 & n35742;
  assign po371 = n35734 | n35743;
  assign n35745 = pi215 & ~n10178;
  assign n35746 = ~pi947 & n21251;
  assign n35747 = pi681 & pi907;
  assign n35748 = ~pi947 & n35747;
  assign n35749 = ~n6168 & ~n16688;
  assign n35750 = n16696 & n16707;
  assign n35751 = ~pi642 & ~n35750;
  assign n35752 = ~n35749 & n35751;
  assign n35753 = pi947 & ~n35752;
  assign n35754 = ~n35748 & ~n35753;
  assign n35755 = ~n35746 & n35754;
  assign n35756 = pi299 & ~n35755;
  assign n35757 = n21331 & ~n35747;
  assign n35758 = ~pi642 & n16785;
  assign n35759 = ~n6197 & ~n35758;
  assign n35760 = ~pi642 & n16750;
  assign n35761 = n6168 & ~n35760;
  assign n35762 = n16752 & n16854;
  assign n35763 = ~n6164 & n16661;
  assign n35764 = ~pi642 & n35763;
  assign n35765 = ~n6168 & ~n35764;
  assign n35766 = ~n35762 & n35765;
  assign n35767 = ~n35761 & ~n35766;
  assign n35768 = n6197 & ~n35767;
  assign n35769 = pi947 & ~n35759;
  assign n35770 = ~n35768 & n35769;
  assign n35771 = ~n3053 & ~n35770;
  assign n35772 = ~n35757 & n35771;
  assign n35773 = n3053 & ~n16661;
  assign n35774 = pi642 & pi947;
  assign n35775 = ~n35748 & ~n35774;
  assign n35776 = n3053 & ~n35775;
  assign n35777 = ~pi223 & ~n35776;
  assign n35778 = ~n35773 & n35777;
  assign n35779 = ~n35772 & n35778;
  assign n35780 = ~n6168 & ~n16694;
  assign n35781 = n6168 & ~n16683;
  assign n35782 = ~pi642 & ~n35781;
  assign n35783 = ~n35780 & n35782;
  assign n35784 = n6197 & ~n35783;
  assign n35785 = ~n6197 & ~n35752;
  assign n35786 = pi947 & ~n35785;
  assign n35787 = ~n35784 & n35786;
  assign n35788 = ~n20981 & ~n35787;
  assign n35789 = pi223 & ~n35748;
  assign n35790 = ~n35788 & n35789;
  assign n35791 = ~pi299 & ~n35790;
  assign n35792 = ~n35779 & n35791;
  assign n35793 = ~n35756 & ~n35792;
  assign n35794 = pi215 & ~n35793;
  assign n35795 = n16758 & n35748;
  assign n35796 = pi642 & ~n16708;
  assign n35797 = n16661 & n35796;
  assign n35798 = pi642 & n16708;
  assign n35799 = ~n16717 & n35798;
  assign n35800 = ~n16767 & n35799;
  assign n35801 = ~n35797 & ~n35800;
  assign n35802 = pi947 & ~n35801;
  assign n35803 = n6197 & ~n35802;
  assign n35804 = ~n35795 & n35803;
  assign n35805 = n16782 & n35747;
  assign n35806 = ~pi947 & ~n35805;
  assign n35807 = ~n6168 & n16779;
  assign n35808 = ~n16784 & ~n35807;
  assign n35809 = n35798 & n35808;
  assign n35810 = ~n16779 & n35796;
  assign n35811 = pi947 & ~n35810;
  assign n35812 = ~n35809 & n35811;
  assign n35813 = ~n35806 & ~n35812;
  assign n35814 = ~n6197 & ~n35813;
  assign n35815 = ~n3053 & ~n35814;
  assign n35816 = ~n35804 & n35815;
  assign n35817 = n16661 & n35776;
  assign n35818 = ~pi223 & ~n35817;
  assign n35819 = ~n35816 & n35818;
  assign n35820 = n6197 & ~n16694;
  assign n35821 = n35747 & ~n35820;
  assign n35822 = ~pi947 & ~n35821;
  assign n35823 = pi947 & ~n16679;
  assign n35824 = ~n16688 & ~n35823;
  assign n35825 = ~n6197 & n35824;
  assign n35826 = ~n16712 & n35799;
  assign n35827 = pi947 & ~n35797;
  assign n35828 = ~n35826 & n35827;
  assign n35829 = ~n35825 & ~n35828;
  assign n35830 = ~n35822 & n35829;
  assign n35831 = pi223 & ~n35830;
  assign n35832 = ~n35819 & ~n35831;
  assign n35833 = ~pi299 & ~n35832;
  assign n35834 = ~n3461 & n35813;
  assign n35835 = n16799 & ~n35775;
  assign n35836 = pi299 & ~n35835;
  assign n35837 = ~n35834 & n35836;
  assign n35838 = ~pi215 & ~n35837;
  assign n35839 = ~n35833 & n35838;
  assign n35840 = ~n35794 & ~n35839;
  assign n35841 = pi39 & ~n35840;
  assign n35842 = pi215 & ~n16649;
  assign n35843 = n16649 & ~n35775;
  assign n35844 = pi299 & ~n35842;
  assign n35845 = ~n35843 & n35844;
  assign n35846 = n16653 & ~n35775;
  assign n35847 = pi215 & ~n16653;
  assign n35848 = ~pi299 & ~n35846;
  assign n35849 = ~n35847 & n35848;
  assign n35850 = ~pi39 & ~n35845;
  assign n35851 = ~n35849 & n35850;
  assign n35852 = ~pi38 & ~n35851;
  assign n35853 = ~n35841 & n35852;
  assign n35854 = n16968 & ~n35775;
  assign n35855 = pi215 & ~n16968;
  assign n35856 = pi38 & ~n35854;
  assign n35857 = ~n35855 & n35856;
  assign n35858 = n10178 & ~n35857;
  assign n35859 = ~n35853 & n35858;
  assign po372 = n35745 | n35859;
  assign n35861 = pi662 & pi907;
  assign n35862 = ~pi947 & n35861;
  assign n35863 = pi614 & pi947;
  assign n35864 = ~n35862 & ~n35863;
  assign n35865 = n16968 & ~n35864;
  assign n35866 = pi216 & ~n16968;
  assign n35867 = pi38 & ~n35865;
  assign n35868 = ~n35866 & n35867;
  assign n35869 = ~pi947 & n20926;
  assign n35870 = ~pi614 & n16785;
  assign n35871 = pi947 & ~n35870;
  assign n35872 = ~n35862 & ~n35871;
  assign n35873 = ~n35869 & n35872;
  assign n35874 = pi216 & ~n35873;
  assign n35875 = n35808 & n35863;
  assign n35876 = n16782 & n35862;
  assign n35877 = ~n35875 & ~n35876;
  assign n35878 = n5752 & ~n35877;
  assign n35879 = n16799 & ~n35864;
  assign n35880 = ~n35878 & ~n35879;
  assign n35881 = ~n35874 & n35880;
  assign n35882 = ~pi215 & ~n35881;
  assign n35883 = ~n17125 & ~n33284;
  assign n35884 = ~n33283 & n35883;
  assign n35885 = n16761 & ~n35884;
  assign n35886 = ~pi614 & ~n16677;
  assign n35887 = n6168 & n35886;
  assign n35888 = ~n35885 & ~n35887;
  assign n35889 = pi947 & n35888;
  assign n35890 = pi216 & ~n35862;
  assign n35891 = ~n35889 & n35890;
  assign n35892 = ~n35746 & n35891;
  assign n35893 = n16688 & n35861;
  assign n35894 = ~pi947 & ~n35893;
  assign n35895 = ~n16712 & n16769;
  assign n35896 = pi947 & ~n16772;
  assign n35897 = ~n35895 & n35896;
  assign n35898 = pi947 & n16679;
  assign n35899 = ~n35897 & ~n35898;
  assign n35900 = ~n35894 & n35899;
  assign n35901 = ~pi216 & ~n35900;
  assign n35902 = pi215 & ~n35901;
  assign n35903 = ~n35892 & n35902;
  assign n35904 = pi299 & ~n35903;
  assign n35905 = ~n35882 & n35904;
  assign n35906 = pi947 & ~n16766;
  assign n35907 = ~pi947 & n16776;
  assign n35908 = ~n35861 & n35907;
  assign n35909 = ~n35906 & ~n35908;
  assign n35910 = n6197 & ~n35909;
  assign n35911 = ~pi947 & ~n16785;
  assign n35912 = ~n6197 & ~n35862;
  assign n35913 = ~n35911 & n35912;
  assign n35914 = ~n35871 & n35913;
  assign n35915 = ~n3053 & ~n35914;
  assign n35916 = ~n35910 & n35915;
  assign n35917 = n3053 & ~n35864;
  assign n35918 = ~pi223 & ~n35917;
  assign n35919 = ~n35773 & n35918;
  assign n35920 = ~n35916 & n35919;
  assign n35921 = ~pi616 & n16685;
  assign n35922 = ~n6168 & ~n16721;
  assign n35923 = ~n35921 & n35922;
  assign n35924 = ~pi614 & ~n35781;
  assign n35925 = ~n35923 & n35924;
  assign n35926 = n6197 & ~n35925;
  assign n35927 = ~n6197 & n35888;
  assign n35928 = pi947 & ~n35927;
  assign n35929 = ~n35926 & n35928;
  assign n35930 = ~n20981 & ~n35929;
  assign n35931 = pi223 & ~n35862;
  assign n35932 = ~n35930 & n35931;
  assign n35933 = pi216 & ~n35932;
  assign n35934 = ~n35920 & n35933;
  assign n35935 = n16758 & n35862;
  assign n35936 = pi947 & ~n16773;
  assign n35937 = n6197 & ~n35936;
  assign n35938 = ~n35935 & n35937;
  assign n35939 = ~n6197 & n35877;
  assign n35940 = ~n3053 & ~n35939;
  assign n35941 = ~n35938 & n35940;
  assign n35942 = n16661 & n35917;
  assign n35943 = ~pi223 & ~n35942;
  assign n35944 = ~n35941 & n35943;
  assign n35945 = ~n35820 & n35861;
  assign n35946 = ~pi947 & ~n35945;
  assign n35947 = ~n35825 & ~n35897;
  assign n35948 = ~n35946 & n35947;
  assign n35949 = pi223 & ~n35948;
  assign n35950 = ~pi216 & ~n35949;
  assign n35951 = ~n35944 & n35950;
  assign n35952 = ~pi299 & ~n35951;
  assign n35953 = ~n35934 & n35952;
  assign n35954 = pi39 & ~n35953;
  assign n35955 = ~n35905 & n35954;
  assign n35956 = pi216 & ~n16649;
  assign n35957 = n16649 & ~n35864;
  assign n35958 = pi299 & ~n35956;
  assign n35959 = ~n35957 & n35958;
  assign n35960 = n16653 & ~n35864;
  assign n35961 = pi216 & ~n16653;
  assign n35962 = ~pi299 & ~n35960;
  assign n35963 = ~n35961 & n35962;
  assign n35964 = ~pi39 & ~n35959;
  assign n35965 = ~n35963 & n35964;
  assign n35966 = ~pi38 & ~n35965;
  assign n35967 = ~n35955 & n35966;
  assign n35968 = ~n35868 & ~n35967;
  assign n35969 = n10178 & ~n35968;
  assign n35970 = ~pi216 & ~n10178;
  assign po373 = ~n35969 & ~n35970;
  assign n35972 = ~pi695 & ~n35407;
  assign n35973 = pi695 & ~n35409;
  assign n35974 = ~pi217 & ~n35973;
  assign n35975 = ~n35972 & n35974;
  assign n35976 = ~pi695 & n35515;
  assign n35977 = pi217 & ~n35976;
  assign n35978 = ~pi612 & ~n35977;
  assign n35979 = ~n35975 & n35978;
  assign n35980 = ~pi695 & ~n35442;
  assign n35981 = pi695 & ~n35450;
  assign n35982 = ~pi217 & ~n35981;
  assign n35983 = ~n35980 & n35982;
  assign n35984 = ~pi695 & n35498;
  assign n35985 = pi695 & n35522;
  assign n35986 = pi217 & ~n35985;
  assign n35987 = ~n35984 & n35986;
  assign n35988 = pi612 & ~n35987;
  assign n35989 = ~n35983 & n35988;
  assign po374 = n35979 | n35989;
  assign n35991 = ~n34671 & ~n34710;
  assign n35992 = n34671 & ~n34776;
  assign n35993 = ~n35991 & ~n35992;
  assign n35994 = ~pi218 & ~n35993;
  assign n35995 = n34671 & n34784;
  assign n35996 = pi218 & ~n35995;
  assign po375 = ~n35994 & ~n35996;
  assign n35998 = ~pi219 & ~po1038;
  assign n35999 = pi617 & ~n35671;
  assign n36000 = ~pi617 & ~n35669;
  assign n36001 = pi637 & ~n35999;
  assign n36002 = ~n36000 & n36001;
  assign n36003 = pi617 & ~pi637;
  assign n36004 = n35675 & n36003;
  assign n36005 = ~n36002 & ~n36004;
  assign n36006 = n35998 & ~n36005;
  assign n36007 = ~pi617 & n35655;
  assign n36008 = pi617 & n35657;
  assign n36009 = pi637 & ~n36007;
  assign n36010 = ~n36008 & n36009;
  assign n36011 = pi617 & n35661;
  assign n36012 = ~pi617 & n17494;
  assign n36013 = ~pi637 & ~n36012;
  assign n36014 = ~n36011 & n36013;
  assign n36015 = ~po1038 & ~n36014;
  assign n36016 = ~n36010 & n36015;
  assign n36017 = pi219 & ~n36016;
  assign po376 = n36006 | n36017;
  assign n36019 = ~n34504 & ~n34795;
  assign n36020 = ~n34650 & n34795;
  assign n36021 = ~n36019 & ~n36020;
  assign n36022 = ~pi220 & ~n36021;
  assign n36023 = n34659 & n34795;
  assign n36024 = pi220 & ~n36023;
  assign po377 = ~n36022 & ~n36024;
  assign n36026 = pi661 & pi907;
  assign n36027 = ~pi947 & n36026;
  assign n36028 = pi616 & pi947;
  assign n36029 = ~n36027 & ~n36028;
  assign n36030 = n16968 & ~n36029;
  assign n36031 = pi221 & ~n16968;
  assign n36032 = pi38 & ~n36030;
  assign n36033 = ~n36031 & n36032;
  assign n36034 = n16709 & n16756;
  assign n36035 = n16766 & ~n16770;
  assign n36036 = n16713 & ~n36035;
  assign n36037 = ~n36034 & ~n36036;
  assign n36038 = pi947 & ~n36037;
  assign n36039 = n6197 & ~n35907;
  assign n36040 = ~n36038 & n36039;
  assign n36041 = ~n6170 & n16756;
  assign n36042 = ~n16778 & ~n36041;
  assign n36043 = n16709 & ~n36042;
  assign n36044 = ~n35758 & ~n35809;
  assign n36045 = n16713 & ~n36044;
  assign n36046 = pi947 & ~n36045;
  assign n36047 = ~n36043 & n36046;
  assign n36048 = ~n35911 & ~n36047;
  assign n36049 = ~n6197 & ~n36048;
  assign n36050 = ~n36027 & ~n36049;
  assign n36051 = ~n36040 & n36050;
  assign n36052 = ~n3053 & ~n36051;
  assign n36053 = n16661 & ~n36029;
  assign n36054 = n3053 & n36053;
  assign n36055 = ~pi223 & ~n36054;
  assign n36056 = ~n35773 & n36055;
  assign n36057 = ~n36052 & n36056;
  assign n36058 = ~n16679 & ~n16686;
  assign n36059 = ~n6168 & ~n36058;
  assign n36060 = ~pi616 & ~n35750;
  assign n36061 = ~n36059 & n36060;
  assign n36062 = pi947 & ~n36061;
  assign n36063 = ~pi947 & ~n16704;
  assign n36064 = ~n36062 & ~n36063;
  assign n36065 = ~n6197 & ~n36064;
  assign n36066 = ~pi947 & n16726;
  assign n36067 = pi947 & ~n16716;
  assign n36068 = n6197 & ~n36067;
  assign n36069 = ~n36066 & n36068;
  assign n36070 = pi223 & ~n36027;
  assign n36071 = ~n36069 & n36070;
  assign n36072 = ~n36065 & n36071;
  assign n36073 = pi221 & ~n36072;
  assign n36074 = ~n36057 & n36073;
  assign n36075 = n16758 & n36027;
  assign n36076 = n16719 & ~n16767;
  assign n36077 = ~n16722 & ~n36076;
  assign n36078 = pi947 & ~n36077;
  assign n36079 = n6197 & ~n36078;
  assign n36080 = ~n36075 & n36079;
  assign n36081 = n35808 & n36028;
  assign n36082 = n16782 & n36027;
  assign n36083 = ~n36081 & ~n36082;
  assign n36084 = ~n6197 & n36083;
  assign n36085 = ~n3053 & ~n36084;
  assign n36086 = ~n36080 & n36085;
  assign n36087 = n36055 & ~n36086;
  assign n36088 = pi947 & ~n16723;
  assign n36089 = n35820 & ~n36088;
  assign n36090 = ~n36027 & ~n36088;
  assign n36091 = ~n35825 & ~n36090;
  assign n36092 = ~n36089 & n36091;
  assign n36093 = pi223 & ~n36092;
  assign n36094 = ~pi221 & ~n36093;
  assign n36095 = ~n36087 & n36094;
  assign n36096 = ~pi299 & ~n36095;
  assign n36097 = ~n36074 & n36096;
  assign n36098 = ~n20926 & ~n36026;
  assign n36099 = ~pi947 & ~n36098;
  assign n36100 = pi221 & ~n36047;
  assign n36101 = ~n36099 & n36100;
  assign n36102 = pi216 & ~n36083;
  assign n36103 = ~pi216 & n36053;
  assign n36104 = ~pi221 & ~n36103;
  assign n36105 = ~n36102 & n36104;
  assign n36106 = ~pi215 & ~n36105;
  assign n36107 = ~n36101 & n36106;
  assign n36108 = pi221 & ~n36027;
  assign n36109 = ~n36062 & n36108;
  assign n36110 = ~n35746 & n36109;
  assign n36111 = ~n35824 & ~n36090;
  assign n36112 = ~pi221 & ~n36111;
  assign n36113 = pi215 & ~n36112;
  assign n36114 = ~n36110 & n36113;
  assign n36115 = pi299 & ~n36114;
  assign n36116 = ~n36107 & n36115;
  assign n36117 = pi39 & ~n36097;
  assign n36118 = ~n36116 & n36117;
  assign n36119 = pi221 & ~n16649;
  assign n36120 = n16649 & ~n36029;
  assign n36121 = pi299 & ~n36119;
  assign n36122 = ~n36120 & n36121;
  assign n36123 = n16653 & ~n36029;
  assign n36124 = pi221 & ~n16653;
  assign n36125 = ~pi299 & ~n36123;
  assign n36126 = ~n36124 & n36125;
  assign n36127 = ~pi39 & ~n36122;
  assign n36128 = ~n36126 & n36127;
  assign n36129 = ~pi38 & ~n36128;
  assign n36130 = ~n36118 & n36129;
  assign n36131 = ~n36033 & ~n36130;
  assign n36132 = n10178 & ~n36131;
  assign n36133 = ~pi221 & ~n10178;
  assign po378 = ~n36132 & ~n36133;
  assign n36135 = ~pi223 & ~n16787;
  assign n36136 = ~n16729 & ~n36135;
  assign n36137 = ~pi299 & ~n36136;
  assign n36138 = pi39 & ~n36137;
  assign n36139 = ~n16813 & n36138;
  assign n36140 = ~pi38 & ~n18015;
  assign n36141 = ~n36139 & n36140;
  assign n36142 = n18809 & ~n36141;
  assign n36143 = pi222 & ~n36142;
  assign n36144 = n17904 & ~n36143;
  assign n36145 = pi222 & ~n3268;
  assign n36146 = pi616 & ~n17084;
  assign n36147 = ~pi616 & n36042;
  assign n36148 = ~n36146 & ~n36147;
  assign n36149 = ~n16707 & ~n36148;
  assign n36150 = ~n6166 & n36148;
  assign n36151 = pi616 & n16842;
  assign n36152 = n17043 & ~n36151;
  assign n36153 = ~n16847 & ~n36152;
  assign n36154 = n6166 & ~n36153;
  assign n36155 = n16707 & ~n36154;
  assign n36156 = ~n36150 & n36155;
  assign n36157 = ~n36149 & ~n36156;
  assign n36158 = ~n6223 & n36157;
  assign n36159 = pi616 & ~n16855;
  assign n36160 = ~n16757 & ~n36159;
  assign n36161 = ~n16707 & ~n36160;
  assign n36162 = ~n6166 & n36160;
  assign n36163 = n6166 & ~n36151;
  assign n36164 = n16750 & n36163;
  assign n36165 = n16707 & ~n36164;
  assign n36166 = ~n36162 & n36165;
  assign n36167 = ~n36161 & ~n36166;
  assign n36168 = n6223 & n36167;
  assign n36169 = pi222 & ~n36168;
  assign n36170 = ~n36158 & n36169;
  assign n36171 = ~n6168 & n16922;
  assign n36172 = ~n16921 & ~n36171;
  assign n36173 = pi616 & ~n36172;
  assign n36174 = n6223 & ~n36173;
  assign n36175 = ~n16779 & n36151;
  assign n36176 = ~n16707 & ~n36175;
  assign n36177 = ~n6166 & n36175;
  assign n36178 = pi616 & n6166;
  assign n36179 = n17044 & n36178;
  assign n36180 = n16707 & ~n36179;
  assign n36181 = ~n36177 & n36180;
  assign n36182 = ~n36176 & ~n36181;
  assign n36183 = ~n6223 & ~n36182;
  assign n36184 = ~pi222 & ~n36174;
  assign n36185 = ~n36183 & n36184;
  assign n36186 = ~n3461 & ~n36185;
  assign n36187 = ~n36170 & n36186;
  assign n36188 = n16721 & n16842;
  assign n36189 = pi222 & ~n16661;
  assign n36190 = n3461 & ~n36189;
  assign n36191 = ~n36188 & n36190;
  assign n36192 = ~pi215 & ~n36191;
  assign n36193 = ~n36187 & n36192;
  assign n36194 = ~n16938 & ~n36171;
  assign n36195 = pi616 & ~n36194;
  assign n36196 = ~pi222 & n36195;
  assign n36197 = ~n16944 & n36196;
  assign n36198 = pi616 & ~n16879;
  assign n36199 = n16688 & ~n36198;
  assign n36200 = ~n16707 & ~n36199;
  assign n36201 = ~n6166 & ~n16688;
  assign n36202 = ~n16696 & ~n36198;
  assign n36203 = ~n36201 & n36202;
  assign n36204 = n16707 & ~n36203;
  assign n36205 = ~n36200 & ~n36204;
  assign n36206 = ~n6223 & n36205;
  assign n36207 = ~n16693 & ~n36159;
  assign n36208 = ~n16707 & ~n36207;
  assign n36209 = ~n6166 & n36207;
  assign n36210 = n16683 & n36163;
  assign n36211 = n16707 & ~n36210;
  assign n36212 = ~n36209 & n36211;
  assign n36213 = ~n36208 & ~n36212;
  assign n36214 = n6223 & n36213;
  assign n36215 = pi222 & ~n36206;
  assign n36216 = ~n36214 & n36215;
  assign n36217 = ~n36197 & ~n36216;
  assign n36218 = pi215 & ~n36217;
  assign n36219 = pi299 & ~n36218;
  assign n36220 = ~n36193 & n36219;
  assign n36221 = ~n6197 & n36157;
  assign n36222 = n6197 & n36167;
  assign n36223 = pi222 & ~n36222;
  assign n36224 = ~n36221 & n36223;
  assign n36225 = n6197 & n36173;
  assign n36226 = ~n6197 & n36182;
  assign n36227 = pi224 & ~n36225;
  assign n36228 = ~n36226 & n36227;
  assign n36229 = ~pi224 & ~n36188;
  assign n36230 = ~pi222 & ~n36229;
  assign n36231 = ~n36228 & n36230;
  assign n36232 = ~pi223 & ~n36231;
  assign n36233 = ~n36224 & n36232;
  assign n36234 = ~n6197 & n36205;
  assign n36235 = n6197 & n36213;
  assign n36236 = pi222 & ~n36234;
  assign n36237 = ~n36235 & n36236;
  assign n36238 = ~n16956 & n36196;
  assign n36239 = pi223 & ~n36238;
  assign n36240 = ~n36237 & n36239;
  assign n36241 = ~n36233 & ~n36240;
  assign n36242 = ~pi299 & ~n36241;
  assign n36243 = pi39 & ~n36220;
  assign n36244 = ~n36242 & n36243;
  assign n36245 = pi222 & n16839;
  assign n36246 = ~pi616 & n16918;
  assign n36247 = ~pi222 & ~n16918;
  assign n36248 = ~pi39 & ~n36246;
  assign n36249 = ~n36247 & n36248;
  assign n36250 = ~n36245 & n36249;
  assign n36251 = ~pi38 & ~n36250;
  assign n36252 = ~n36244 & n36251;
  assign n36253 = pi222 & ~n16968;
  assign n36254 = pi38 & ~n36253;
  assign n36255 = pi616 & n16970;
  assign n36256 = n36254 & ~n36255;
  assign n36257 = n3268 & ~n36256;
  assign n36258 = ~n36252 & n36257;
  assign n36259 = ~n36145 & ~n36258;
  assign n36260 = ~n17526 & ~n36259;
  assign n36261 = n17526 & n36143;
  assign n36262 = ~n36260 & ~n36261;
  assign n36263 = ~pi785 & ~n36262;
  assign n36264 = pi609 & n36262;
  assign n36265 = ~pi609 & ~n36143;
  assign n36266 = pi1155 & ~n36265;
  assign n36267 = ~n36264 & n36266;
  assign n36268 = ~pi609 & n36262;
  assign n36269 = pi609 & ~n36143;
  assign n36270 = ~pi1155 & ~n36269;
  assign n36271 = ~n36268 & n36270;
  assign n36272 = ~n36267 & ~n36271;
  assign n36273 = pi785 & ~n36272;
  assign n36274 = ~n36263 & ~n36273;
  assign n36275 = ~pi781 & ~n36274;
  assign n36276 = pi618 & n36274;
  assign n36277 = ~pi618 & ~n36143;
  assign n36278 = pi1154 & ~n36277;
  assign n36279 = ~n36276 & n36278;
  assign n36280 = ~pi618 & n36274;
  assign n36281 = pi618 & ~n36143;
  assign n36282 = ~pi1154 & ~n36281;
  assign n36283 = ~n36280 & n36282;
  assign n36284 = ~n36279 & ~n36283;
  assign n36285 = pi781 & ~n36284;
  assign n36286 = ~n36275 & ~n36285;
  assign n36287 = ~pi789 & ~n36286;
  assign n36288 = pi619 & n36286;
  assign n36289 = ~pi619 & ~n36143;
  assign n36290 = pi1159 & ~n36289;
  assign n36291 = ~n36288 & n36290;
  assign n36292 = ~pi619 & n36286;
  assign n36293 = pi619 & ~n36143;
  assign n36294 = ~pi1159 & ~n36293;
  assign n36295 = ~n36292 & n36294;
  assign n36296 = ~n36291 & ~n36295;
  assign n36297 = pi789 & ~n36296;
  assign n36298 = ~n36287 & ~n36297;
  assign n36299 = ~n17904 & n36298;
  assign n36300 = ~n36144 & ~n36299;
  assign n36301 = ~n20502 & n36300;
  assign n36302 = ~n19215 & ~n36143;
  assign n36303 = pi661 & pi680;
  assign n36304 = n17325 & ~n36303;
  assign n36305 = ~pi222 & ~n17325;
  assign n36306 = pi222 & n17305;
  assign n36307 = ~pi299 & ~n36306;
  assign n36308 = ~n36304 & n36307;
  assign n36309 = ~n36305 & n36308;
  assign n36310 = n17334 & ~n36303;
  assign n36311 = ~pi222 & ~n17334;
  assign n36312 = pi222 & n17311;
  assign n36313 = pi299 & ~n36312;
  assign n36314 = ~n36310 & n36313;
  assign n36315 = ~n36311 & n36314;
  assign n36316 = ~pi39 & ~n36309;
  assign n36317 = ~n36315 & n36316;
  assign n36318 = ~n6166 & ~n16758;
  assign n36319 = ~pi662 & n16767;
  assign n36320 = ~n36318 & ~n36319;
  assign n36321 = n16707 & ~n36320;
  assign n36322 = pi661 & ~n17425;
  assign n36323 = ~pi661 & n16759;
  assign n36324 = ~n36321 & ~n36323;
  assign n36325 = ~n36322 & n36324;
  assign n36326 = n6197 & n36325;
  assign n36327 = ~pi661 & ~n16785;
  assign n36328 = pi680 & n17239;
  assign n36329 = ~n17042 & ~n36328;
  assign n36330 = pi661 & ~n36329;
  assign n36331 = ~n36327 & ~n36330;
  assign n36332 = ~n6197 & n36331;
  assign n36333 = pi222 & ~n36332;
  assign n36334 = ~n36326 & n36333;
  assign n36335 = ~n17386 & n36303;
  assign n36336 = n6197 & n36335;
  assign n36337 = pi661 & n17392;
  assign n36338 = ~n6197 & n36337;
  assign n36339 = pi224 & ~n36336;
  assign n36340 = ~n36338 & n36339;
  assign n36341 = pi661 & n17410;
  assign n36342 = ~pi224 & ~n36341;
  assign n36343 = ~pi222 & ~n36342;
  assign n36344 = ~n36340 & n36343;
  assign n36345 = ~pi223 & ~n36344;
  assign n36346 = ~n36334 & n36345;
  assign n36347 = ~pi661 & ~n16726;
  assign n36348 = ~n17002 & ~n17443;
  assign n36349 = pi661 & ~n36348;
  assign n36350 = ~n36347 & ~n36349;
  assign n36351 = n6197 & n36350;
  assign n36352 = n16699 & n16707;
  assign n36353 = ~pi661 & n16689;
  assign n36354 = pi661 & ~n17448;
  assign n36355 = ~n36353 & ~n36354;
  assign n36356 = ~n36352 & n36355;
  assign n36357 = ~n6197 & n36356;
  assign n36358 = pi222 & ~n36357;
  assign n36359 = ~n36351 & n36358;
  assign n36360 = ~pi222 & pi661;
  assign n36361 = n17401 & n36360;
  assign n36362 = pi223 & ~n36361;
  assign n36363 = ~n36359 & n36362;
  assign n36364 = ~n36346 & ~n36363;
  assign n36365 = ~pi299 & ~n36364;
  assign n36366 = n6223 & n36325;
  assign n36367 = ~n6223 & n36331;
  assign n36368 = pi222 & ~n36367;
  assign n36369 = ~n36366 & n36368;
  assign n36370 = ~n6223 & ~n36337;
  assign n36371 = n6223 & ~n36335;
  assign n36372 = ~pi222 & ~n36370;
  assign n36373 = ~n36371 & n36372;
  assign n36374 = ~n3461 & ~n36373;
  assign n36375 = ~n36369 & n36374;
  assign n36376 = n36190 & ~n36341;
  assign n36377 = ~pi215 & ~n36376;
  assign n36378 = ~n36375 & n36377;
  assign n36379 = n17414 & n36360;
  assign n36380 = n6223 & n36350;
  assign n36381 = ~n6223 & n36356;
  assign n36382 = pi222 & ~n36381;
  assign n36383 = ~n36380 & n36382;
  assign n36384 = ~n36379 & ~n36383;
  assign n36385 = pi215 & ~n36384;
  assign n36386 = pi299 & ~n36385;
  assign n36387 = ~n36378 & n36386;
  assign n36388 = ~n36365 & ~n36387;
  assign n36389 = pi39 & ~n36388;
  assign n36390 = ~n36317 & ~n36389;
  assign n36391 = ~pi38 & ~n36390;
  assign n36392 = pi661 & n17479;
  assign n36393 = n36254 & ~n36392;
  assign n36394 = n3268 & ~n36393;
  assign n36395 = ~n36391 & n36394;
  assign n36396 = ~n36145 & ~n36395;
  assign n36397 = ~pi778 & ~n36396;
  assign n36398 = pi625 & n36396;
  assign n36399 = ~pi625 & ~n36143;
  assign n36400 = pi1153 & ~n36399;
  assign n36401 = ~n36398 & n36400;
  assign n36402 = ~pi625 & n36396;
  assign n36403 = pi625 & ~n36143;
  assign n36404 = ~pi1153 & ~n36403;
  assign n36405 = ~n36402 & n36404;
  assign n36406 = ~n36401 & ~n36405;
  assign n36407 = pi778 & ~n36406;
  assign n36408 = ~n36397 & ~n36407;
  assign n36409 = ~n17554 & ~n36408;
  assign n36410 = n17554 & n36143;
  assign n36411 = ~n36409 & ~n36410;
  assign n36412 = ~n17591 & ~n36411;
  assign n36413 = n17591 & n36143;
  assign n36414 = ~n36412 & ~n36413;
  assign n36415 = ~n17627 & n36414;
  assign n36416 = ~n17670 & n36415;
  assign n36417 = ~n36302 & ~n36416;
  assign n36418 = ~pi628 & ~n36417;
  assign n36419 = pi628 & ~n36143;
  assign n36420 = n17696 & ~n36419;
  assign n36421 = ~n36418 & n36420;
  assign n36422 = pi628 & ~n36417;
  assign n36423 = ~pi628 & ~n36143;
  assign n36424 = n17695 & ~n36423;
  assign n36425 = ~n36422 & n36424;
  assign n36426 = ~n36421 & ~n36425;
  assign n36427 = ~n36301 & n36426;
  assign n36428 = pi792 & ~n36427;
  assign n36429 = ~pi680 & n36148;
  assign n36430 = n6170 & n17029;
  assign n36431 = ~n16986 & ~n36430;
  assign n36432 = ~pi603 & n36431;
  assign n36433 = pi603 & n16748;
  assign n36434 = ~n17033 & ~n36433;
  assign n36435 = ~n36432 & n36434;
  assign n36436 = ~pi642 & n36435;
  assign n36437 = ~n17172 & n36431;
  assign n36438 = pi642 & ~n36437;
  assign n36439 = n6164 & ~n36436;
  assign n36440 = ~n36438 & n36439;
  assign n36441 = n17125 & n36437;
  assign n36442 = n17181 & ~n36431;
  assign n36443 = pi616 & ~n36442;
  assign n36444 = pi680 & ~n36443;
  assign n36445 = ~n36441 & n36444;
  assign n36446 = ~n36440 & n36445;
  assign n36447 = pi661 & ~n36446;
  assign n36448 = ~n36429 & n36447;
  assign n36449 = ~pi661 & pi681;
  assign n36450 = ~n36148 & n36449;
  assign n36451 = ~n36156 & ~n36450;
  assign n36452 = ~n36448 & n36451;
  assign n36453 = ~n6223 & ~n36452;
  assign n36454 = ~pi680 & n36160;
  assign n36455 = pi616 & ~n17247;
  assign n36456 = pi680 & ~n36455;
  assign n36457 = ~n17025 & n36456;
  assign n36458 = pi661 & ~n36454;
  assign n36459 = ~n36457 & n36458;
  assign n36460 = ~n36160 & n36449;
  assign n36461 = ~n36166 & ~n36460;
  assign n36462 = ~n36459 & n36461;
  assign n36463 = n6223 & ~n36462;
  assign n36464 = pi222 & ~n36463;
  assign n36465 = ~n36453 & n36464;
  assign n36466 = pi616 & n17173;
  assign n36467 = pi680 & ~n36466;
  assign n36468 = ~n17096 & n36467;
  assign n36469 = ~pi680 & n36175;
  assign n36470 = pi661 & ~n36469;
  assign n36471 = ~n36468 & n36470;
  assign n36472 = ~n36175 & n36449;
  assign n36473 = ~n36181 & ~n36472;
  assign n36474 = ~n36471 & n36473;
  assign n36475 = ~n6223 & n36474;
  assign n36476 = pi616 & ~n17182;
  assign n36477 = pi680 & ~n17114;
  assign n36478 = ~n36476 & n36477;
  assign n36479 = ~pi680 & n36188;
  assign n36480 = pi661 & ~n36479;
  assign n36481 = ~n36478 & n36480;
  assign n36482 = n16920 & n36178;
  assign n36483 = ~n6166 & n36188;
  assign n36484 = n16707 & ~n36483;
  assign n36485 = ~n36482 & n36484;
  assign n36486 = ~n36188 & n36449;
  assign n36487 = ~n36485 & ~n36486;
  assign n36488 = ~n36481 & n36487;
  assign n36489 = n6223 & n36488;
  assign n36490 = ~pi222 & ~n36489;
  assign n36491 = ~n36475 & n36490;
  assign n36492 = ~n36465 & ~n36491;
  assign n36493 = ~n3461 & ~n36492;
  assign n36494 = ~n36151 & ~n36303;
  assign n36495 = ~pi616 & ~n17104;
  assign n36496 = ~n36476 & ~n36495;
  assign n36497 = ~n36494 & n36496;
  assign n36498 = n36190 & ~n36497;
  assign n36499 = ~pi215 & ~n36498;
  assign n36500 = ~n36493 & n36499;
  assign n36501 = ~n16999 & n36456;
  assign n36502 = ~pi680 & n36207;
  assign n36503 = pi661 & ~n36502;
  assign n36504 = ~n36501 & n36503;
  assign n36505 = ~n36207 & n36449;
  assign n36506 = ~n36212 & ~n36505;
  assign n36507 = ~n36504 & n36506;
  assign n36508 = n6223 & ~n36507;
  assign n36509 = ~pi680 & n36199;
  assign n36510 = ~n17010 & n17181;
  assign n36511 = pi616 & ~n36510;
  assign n36512 = pi680 & ~n36511;
  assign n36513 = n17013 & n36512;
  assign n36514 = pi661 & ~n36513;
  assign n36515 = ~n36509 & n36514;
  assign n36516 = ~n36199 & n36449;
  assign n36517 = ~n36204 & ~n36516;
  assign n36518 = ~n36515 & n36517;
  assign n36519 = ~n6223 & ~n36518;
  assign n36520 = pi222 & ~n36508;
  assign n36521 = ~n36519 & n36520;
  assign n36522 = ~n16939 & ~n17211;
  assign n36523 = pi616 & n36522;
  assign n36524 = pi680 & ~n36523;
  assign n36525 = n17131 & n36524;
  assign n36526 = pi616 & n16939;
  assign n36527 = ~pi680 & n36526;
  assign n36528 = pi661 & ~n36527;
  assign n36529 = ~n36525 & n36528;
  assign n36530 = ~pi661 & ~n36526;
  assign n36531 = ~n16677 & n36188;
  assign n36532 = n6168 & ~n36531;
  assign n36533 = ~n36530 & ~n36532;
  assign n36534 = ~n36529 & n36533;
  assign n36535 = ~n6223 & n36534;
  assign n36536 = n17138 & n36303;
  assign n36537 = ~n36195 & ~n36536;
  assign n36538 = n6223 & ~n36537;
  assign n36539 = ~pi222 & ~n36538;
  assign n36540 = ~n36535 & n36539;
  assign n36541 = pi215 & ~n36540;
  assign n36542 = ~n36521 & n36541;
  assign n36543 = pi299 & ~n36542;
  assign n36544 = ~n36500 & n36543;
  assign n36545 = n36303 & ~n36496;
  assign n36546 = ~n36188 & ~n36303;
  assign n36547 = ~pi222 & ~n36546;
  assign n36548 = ~n36545 & n36547;
  assign n36549 = ~n3305 & ~n36548;
  assign n36550 = ~n6197 & n36474;
  assign n36551 = n6197 & n36488;
  assign n36552 = pi224 & ~n36551;
  assign n36553 = ~n36550 & n36552;
  assign n36554 = ~n36549 & ~n36553;
  assign n36555 = ~n6197 & n36452;
  assign n36556 = n6197 & n36462;
  assign n36557 = pi222 & ~n36556;
  assign n36558 = ~n36555 & n36557;
  assign n36559 = ~n36554 & ~n36558;
  assign n36560 = ~pi223 & ~n36559;
  assign n36561 = n6197 & ~n36507;
  assign n36562 = ~n6197 & ~n36518;
  assign n36563 = pi222 & ~n36561;
  assign n36564 = ~n36562 & n36563;
  assign n36565 = ~n6197 & n36534;
  assign n36566 = n6197 & ~n36537;
  assign n36567 = ~pi222 & ~n36566;
  assign n36568 = ~n36565 & n36567;
  assign n36569 = pi223 & ~n36568;
  assign n36570 = ~n36564 & n36569;
  assign n36571 = ~pi299 & ~n36570;
  assign n36572 = ~n36560 & n36571;
  assign n36573 = pi39 & ~n36572;
  assign n36574 = ~n36544 & n36573;
  assign n36575 = pi661 & n17330;
  assign n36576 = pi616 & n16911;
  assign n36577 = ~pi222 & ~n36576;
  assign n36578 = ~n36575 & n36577;
  assign n36579 = n17329 & ~n36303;
  assign n36580 = ~pi616 & n16911;
  assign n36581 = n17305 & ~n17327;
  assign n36582 = ~n36580 & ~n36581;
  assign n36583 = ~n36579 & n36582;
  assign n36584 = pi222 & ~n36583;
  assign n36585 = ~n36578 & ~n36584;
  assign n36586 = ~pi299 & ~n36585;
  assign n36587 = n17337 & ~n36303;
  assign n36588 = ~pi616 & n16916;
  assign n36589 = ~n16823 & n17311;
  assign n36590 = ~n36588 & ~n36589;
  assign n36591 = ~n36587 & n36590;
  assign n36592 = pi222 & ~n36591;
  assign n36593 = pi661 & n17338;
  assign n36594 = pi616 & n16916;
  assign n36595 = ~pi222 & ~n36594;
  assign n36596 = ~n36593 & n36595;
  assign n36597 = ~n36592 & ~n36596;
  assign n36598 = pi299 & ~n36597;
  assign n36599 = ~pi39 & ~n36586;
  assign n36600 = ~n36598 & n36599;
  assign n36601 = ~pi38 & ~n36600;
  assign n36602 = ~n36574 & n36601;
  assign n36603 = n16665 & n17181;
  assign n36604 = ~pi222 & ~pi616;
  assign n36605 = ~pi39 & pi616;
  assign n36606 = n36303 & n36605;
  assign n36607 = ~n36604 & ~n36606;
  assign n36608 = n36603 & ~n36607;
  assign n36609 = ~pi616 & ~n17054;
  assign n36610 = ~n36494 & ~n36609;
  assign n36611 = n16968 & n36610;
  assign n36612 = ~n36253 & ~n36611;
  assign n36613 = ~n36608 & ~n36612;
  assign n36614 = pi38 & ~n36613;
  assign n36615 = n3268 & ~n36614;
  assign n36616 = ~n36602 & n36615;
  assign n36617 = ~n36145 & ~n36616;
  assign n36618 = ~pi625 & n36617;
  assign n36619 = pi625 & n36259;
  assign n36620 = ~pi1153 & ~n36619;
  assign n36621 = ~n36618 & n36620;
  assign n36622 = ~pi608 & ~n36401;
  assign n36623 = ~n36621 & n36622;
  assign n36624 = pi625 & n36617;
  assign n36625 = ~pi625 & n36259;
  assign n36626 = pi1153 & ~n36625;
  assign n36627 = ~n36624 & n36626;
  assign n36628 = pi608 & ~n36405;
  assign n36629 = ~n36627 & n36628;
  assign n36630 = ~n36623 & ~n36629;
  assign n36631 = pi778 & ~n36630;
  assign n36632 = ~pi778 & n36617;
  assign n36633 = ~n36631 & ~n36632;
  assign n36634 = ~pi609 & ~n36633;
  assign n36635 = pi609 & n36408;
  assign n36636 = ~pi1155 & ~n36635;
  assign n36637 = ~n36634 & n36636;
  assign n36638 = ~pi660 & ~n36267;
  assign n36639 = ~n36637 & n36638;
  assign n36640 = pi609 & ~n36633;
  assign n36641 = ~pi609 & n36408;
  assign n36642 = pi1155 & ~n36641;
  assign n36643 = ~n36640 & n36642;
  assign n36644 = pi660 & ~n36271;
  assign n36645 = ~n36643 & n36644;
  assign n36646 = ~n36639 & ~n36645;
  assign n36647 = pi785 & ~n36646;
  assign n36648 = ~pi785 & ~n36633;
  assign n36649 = ~n36647 & ~n36648;
  assign n36650 = ~pi618 & ~n36649;
  assign n36651 = pi618 & n36411;
  assign n36652 = ~pi1154 & ~n36651;
  assign n36653 = ~n36650 & n36652;
  assign n36654 = ~pi627 & ~n36279;
  assign n36655 = ~n36653 & n36654;
  assign n36656 = pi618 & ~n36649;
  assign n36657 = ~pi618 & n36411;
  assign n36658 = pi1154 & ~n36657;
  assign n36659 = ~n36656 & n36658;
  assign n36660 = pi627 & ~n36283;
  assign n36661 = ~n36659 & n36660;
  assign n36662 = ~n36655 & ~n36661;
  assign n36663 = pi781 & ~n36662;
  assign n36664 = ~pi781 & ~n36649;
  assign n36665 = ~n36663 & ~n36664;
  assign n36666 = ~pi619 & ~n36665;
  assign n36667 = pi619 & n36414;
  assign n36668 = ~pi1159 & ~n36667;
  assign n36669 = ~n36666 & n36668;
  assign n36670 = ~pi648 & ~n36291;
  assign n36671 = ~n36669 & n36670;
  assign n36672 = pi619 & ~n36665;
  assign n36673 = ~pi619 & n36414;
  assign n36674 = pi1159 & ~n36673;
  assign n36675 = ~n36672 & n36674;
  assign n36676 = pi648 & ~n36295;
  assign n36677 = ~n36675 & n36676;
  assign n36678 = pi789 & ~n36671;
  assign n36679 = ~n36677 & n36678;
  assign n36680 = ~pi789 & n36665;
  assign n36681 = ~pi626 & n36298;
  assign n36682 = pi626 & ~n36143;
  assign n36683 = n17668 & ~n36682;
  assign n36684 = ~n36681 & n36683;
  assign n36685 = pi626 & n36298;
  assign n36686 = ~pi626 & ~n36143;
  assign n36687 = n17667 & ~n36686;
  assign n36688 = ~n36685 & n36687;
  assign n36689 = n17627 & ~n36143;
  assign n36690 = n17792 & ~n36689;
  assign n36691 = ~n36415 & n36690;
  assign n36692 = ~n36684 & ~n36691;
  assign n36693 = ~n36688 & n36692;
  assign n36694 = pi788 & ~n36693;
  assign n36695 = ~n36680 & ~n36694;
  assign n36696 = ~n36679 & n36695;
  assign n36697 = ~n17905 & n36693;
  assign n36698 = ~n20298 & ~n36697;
  assign n36699 = ~n36696 & n36698;
  assign n36700 = ~n36428 & ~n36699;
  assign n36701 = n20300 & ~n36700;
  assign n36702 = ~n17698 & n36300;
  assign n36703 = n17698 & n36143;
  assign n36704 = ~n36702 & ~n36703;
  assign n36705 = ~n20491 & ~n36704;
  assign n36706 = ~n19247 & ~n36417;
  assign n36707 = n17946 & ~n36143;
  assign n36708 = ~n36706 & ~n36707;
  assign n36709 = pi647 & ~n36708;
  assign n36710 = ~pi647 & ~n36143;
  assign n36711 = pi1157 & ~n36710;
  assign n36712 = ~n36709 & n36711;
  assign n36713 = ~pi630 & n36712;
  assign n36714 = ~pi647 & ~n36708;
  assign n36715 = pi647 & ~n36143;
  assign n36716 = ~pi1157 & ~n36715;
  assign n36717 = ~n36714 & n36716;
  assign n36718 = pi630 & n36717;
  assign n36719 = ~n36713 & ~n36718;
  assign n36720 = ~n36705 & n36719;
  assign n36721 = pi787 & ~n36720;
  assign n36722 = ~n36701 & ~n36721;
  assign n36723 = pi644 & n36722;
  assign n36724 = ~pi787 & n36708;
  assign n36725 = ~n36712 & ~n36717;
  assign n36726 = pi787 & ~n36725;
  assign n36727 = ~n36724 & ~n36726;
  assign n36728 = ~pi644 & n36727;
  assign n36729 = pi715 & ~n36728;
  assign n36730 = ~n36723 & n36729;
  assign n36731 = n17740 & ~n36143;
  assign n36732 = ~n17740 & n36704;
  assign n36733 = ~n36731 & ~n36732;
  assign n36734 = pi644 & ~n36733;
  assign n36735 = ~pi644 & ~n36143;
  assign n36736 = ~pi715 & ~n36735;
  assign n36737 = ~n36734 & n36736;
  assign n36738 = pi1160 & ~n36737;
  assign n36739 = ~n36730 & n36738;
  assign n36740 = ~pi644 & n36722;
  assign n36741 = pi644 & n36727;
  assign n36742 = ~pi715 & ~n36741;
  assign n36743 = ~n36740 & n36742;
  assign n36744 = ~pi644 & ~n36733;
  assign n36745 = pi644 & ~n36143;
  assign n36746 = pi715 & ~n36745;
  assign n36747 = ~n36744 & n36746;
  assign n36748 = ~pi1160 & ~n36747;
  assign n36749 = ~n36743 & n36748;
  assign n36750 = ~n36739 & ~n36749;
  assign n36751 = pi790 & ~n36750;
  assign n36752 = ~pi790 & n36722;
  assign n36753 = ~n36751 & ~n36752;
  assign n36754 = ~po1038 & ~n36753;
  assign n36755 = ~pi222 & po1038;
  assign po379 = ~n36754 & ~n36755;
  assign n36757 = ~pi299 & ~n16728;
  assign n36758 = pi39 & ~n36757;
  assign n36759 = ~n16813 & n36758;
  assign n36760 = n14819 & ~n18015;
  assign n36761 = ~n36759 & n36760;
  assign n36762 = n18809 & ~n36761;
  assign n36763 = pi223 & ~n36762;
  assign n36764 = n17904 & ~n36763;
  assign n36765 = n17526 & ~n36763;
  assign n36766 = pi223 & ~n3268;
  assign n36767 = pi642 & n16842;
  assign n36768 = n35763 & ~n36767;
  assign n36769 = pi642 & ~n16855;
  assign n36770 = n6164 & ~n36769;
  assign n36771 = ~n16753 & n36770;
  assign n36772 = ~n36768 & ~n36771;
  assign n36773 = pi681 & n36772;
  assign n36774 = ~n6167 & ~n36772;
  assign n36775 = ~n16851 & ~n35760;
  assign n36776 = n6167 & ~n36775;
  assign n36777 = ~pi681 & ~n36776;
  assign n36778 = ~n36774 & n36777;
  assign n36779 = n6223 & ~n36778;
  assign n36780 = ~n36773 & n36779;
  assign n36781 = pi642 & ~n17084;
  assign n36782 = ~pi642 & ~n16782;
  assign n36783 = ~n36781 & ~n36782;
  assign n36784 = pi681 & ~n36783;
  assign n36785 = ~n6167 & n36783;
  assign n36786 = n6167 & ~n36767;
  assign n36787 = ~n16748 & n36786;
  assign n36788 = ~pi681 & ~n36787;
  assign n36789 = ~n36785 & n36788;
  assign n36790 = ~n6223 & ~n36789;
  assign n36791 = ~n36784 & n36790;
  assign n36792 = pi223 & ~n36791;
  assign n36793 = ~n36780 & n36792;
  assign n36794 = pi642 & n16922;
  assign n36795 = ~n6167 & n36794;
  assign n36796 = ~pi681 & ~n36795;
  assign n36797 = pi642 & n6167;
  assign n36798 = n16920 & n36797;
  assign n36799 = n36796 & ~n36798;
  assign n36800 = pi681 & ~n36794;
  assign n36801 = ~n36799 & ~n36800;
  assign n36802 = n20832 & n36801;
  assign n36803 = ~n16779 & n36767;
  assign n36804 = pi681 & ~n36803;
  assign n36805 = ~n6167 & n36803;
  assign n36806 = n17044 & n36797;
  assign n36807 = ~pi681 & ~n36806;
  assign n36808 = ~n36805 & n36807;
  assign n36809 = ~n36804 & ~n36808;
  assign n36810 = ~n20832 & n36809;
  assign n36811 = ~pi947 & ~n36802;
  assign n36812 = ~n36810 & n36811;
  assign n36813 = pi947 & ~n36809;
  assign n36814 = ~pi223 & ~n36813;
  assign n36815 = ~n36812 & n36814;
  assign n36816 = ~n3461 & ~n36815;
  assign n36817 = ~n36793 & n36816;
  assign n36818 = pi223 & ~n16661;
  assign n36819 = n3461 & ~n36818;
  assign n36820 = ~n36794 & n36819;
  assign n36821 = ~pi215 & ~n36820;
  assign n36822 = ~n36817 & n36821;
  assign n36823 = n16938 & n36797;
  assign n36824 = n36796 & ~n36823;
  assign n36825 = pi642 & ~n16879;
  assign n36826 = n6167 & ~n36825;
  assign n36827 = ~n16677 & n36826;
  assign n36828 = ~pi681 & ~n36827;
  assign n36829 = n16679 & n36828;
  assign n36830 = ~n36824 & ~n36829;
  assign n36831 = pi642 & n16939;
  assign n36832 = pi681 & ~n36831;
  assign n36833 = n36830 & ~n36832;
  assign n36834 = ~n20832 & n36833;
  assign n36835 = n6223 & ~n36824;
  assign n36836 = n36794 & n36835;
  assign n36837 = ~pi947 & ~n36836;
  assign n36838 = ~n36834 & n36837;
  assign n36839 = pi947 & ~n36833;
  assign n36840 = ~pi223 & ~n36839;
  assign n36841 = ~n36838 & n36840;
  assign n36842 = n36207 & ~n36769;
  assign n36843 = ~n36768 & ~n36842;
  assign n36844 = pi681 & n36843;
  assign n36845 = ~n6167 & ~n36843;
  assign n36846 = n16665 & ~n36767;
  assign n36847 = n6167 & n36846;
  assign n36848 = n16683 & n36847;
  assign n36849 = ~pi681 & ~n36848;
  assign n36850 = ~n36845 & n36849;
  assign n36851 = ~n36844 & ~n36850;
  assign n36852 = n6223 & n36851;
  assign n36853 = ~pi642 & ~n16688;
  assign n36854 = pi642 & ~n16880;
  assign n36855 = ~n36853 & ~n36854;
  assign n36856 = ~n6167 & n36855;
  assign n36857 = n36828 & ~n36856;
  assign n36858 = pi681 & ~n36855;
  assign n36859 = ~n36857 & ~n36858;
  assign n36860 = ~n6223 & n36859;
  assign n36861 = pi223 & ~n36860;
  assign n36862 = ~n36852 & n36861;
  assign n36863 = ~n36841 & ~n36862;
  assign n36864 = pi215 & ~n36863;
  assign n36865 = pi299 & ~n36864;
  assign n36866 = ~n36822 & n36865;
  assign n36867 = n6197 & n36801;
  assign n36868 = ~n6197 & n36809;
  assign n36869 = ~n3053 & ~n36867;
  assign n36870 = ~n36868 & n36869;
  assign n36871 = n3053 & ~n36794;
  assign n36872 = ~pi223 & ~n36871;
  assign n36873 = ~n36870 & n36872;
  assign n36874 = n6197 & n36851;
  assign n36875 = ~n6197 & n36859;
  assign n36876 = pi223 & ~n36875;
  assign n36877 = ~n36874 & n36876;
  assign n36878 = ~pi299 & ~n36877;
  assign n36879 = ~n36873 & n36878;
  assign n36880 = pi39 & ~n36879;
  assign n36881 = ~n36866 & n36880;
  assign n36882 = ~pi223 & pi642;
  assign n36883 = n16911 & n36882;
  assign n36884 = ~pi299 & ~n36883;
  assign n36885 = ~pi642 & n16911;
  assign n36886 = pi223 & ~n36885;
  assign n36887 = n16837 & n36886;
  assign n36888 = n36884 & ~n36887;
  assign n36889 = n16916 & n36882;
  assign n36890 = pi299 & ~n36889;
  assign n36891 = n6163 & n16915;
  assign n36892 = pi223 & ~n36891;
  assign n36893 = ~n16824 & n36892;
  assign n36894 = n36890 & ~n36893;
  assign n36895 = ~pi39 & ~n36894;
  assign n36896 = ~n36888 & n36895;
  assign n36897 = ~pi38 & ~n36896;
  assign n36898 = ~n36881 & n36897;
  assign n36899 = pi39 & pi223;
  assign n36900 = pi38 & ~n36899;
  assign n36901 = ~pi223 & ~n16665;
  assign n36902 = ~pi39 & ~n36901;
  assign n36903 = ~n36846 & n36902;
  assign n36904 = n36900 & ~n36903;
  assign n36905 = n3268 & ~n36904;
  assign n36906 = ~n36898 & n36905;
  assign n36907 = ~n36766 & ~n36906;
  assign n36908 = ~n17526 & n36907;
  assign n36909 = ~n36765 & ~n36908;
  assign n36910 = ~pi785 & n36909;
  assign n36911 = pi609 & ~n36909;
  assign n36912 = ~pi609 & ~n36763;
  assign n36913 = pi1155 & ~n36912;
  assign n36914 = ~n36911 & n36913;
  assign n36915 = ~pi609 & ~n36909;
  assign n36916 = pi609 & ~n36763;
  assign n36917 = ~pi1155 & ~n36916;
  assign n36918 = ~n36915 & n36917;
  assign n36919 = ~n36914 & ~n36918;
  assign n36920 = pi785 & ~n36919;
  assign n36921 = ~n36910 & ~n36920;
  assign n36922 = ~pi781 & ~n36921;
  assign n36923 = pi618 & n36921;
  assign n36924 = ~pi618 & ~n36763;
  assign n36925 = pi1154 & ~n36924;
  assign n36926 = ~n36923 & n36925;
  assign n36927 = ~pi618 & n36921;
  assign n36928 = pi618 & ~n36763;
  assign n36929 = ~pi1154 & ~n36928;
  assign n36930 = ~n36927 & n36929;
  assign n36931 = ~n36926 & ~n36930;
  assign n36932 = pi781 & ~n36931;
  assign n36933 = ~n36922 & ~n36932;
  assign n36934 = ~pi789 & ~n36933;
  assign n36935 = pi619 & n36933;
  assign n36936 = ~pi619 & ~n36763;
  assign n36937 = pi1159 & ~n36936;
  assign n36938 = ~n36935 & n36937;
  assign n36939 = ~pi619 & n36933;
  assign n36940 = pi619 & ~n36763;
  assign n36941 = ~pi1159 & ~n36940;
  assign n36942 = ~n36939 & n36941;
  assign n36943 = ~n36938 & ~n36942;
  assign n36944 = pi789 & ~n36943;
  assign n36945 = ~n36934 & ~n36944;
  assign n36946 = ~n17904 & n36945;
  assign n36947 = ~n36764 & ~n36946;
  assign n36948 = ~n17698 & n36947;
  assign n36949 = n17698 & n36763;
  assign n36950 = ~n36948 & ~n36949;
  assign n36951 = ~n20491 & ~n36950;
  assign n36952 = ~n19215 & ~n36763;
  assign n36953 = n17554 & ~n36763;
  assign n36954 = pi680 & pi681;
  assign n36955 = n17325 & ~n36954;
  assign n36956 = ~pi223 & ~n17325;
  assign n36957 = pi223 & n17305;
  assign n36958 = ~pi299 & ~n36957;
  assign n36959 = ~n36955 & n36958;
  assign n36960 = ~n36956 & n36959;
  assign n36961 = n17334 & ~n36954;
  assign n36962 = ~pi223 & ~n17334;
  assign n36963 = pi223 & n17311;
  assign n36964 = pi299 & ~n36963;
  assign n36965 = ~n36961 & n36964;
  assign n36966 = ~n36962 & n36965;
  assign n36967 = ~pi39 & ~n36960;
  assign n36968 = ~n36966 & n36967;
  assign n36969 = pi681 & n17410;
  assign n36970 = n36819 & ~n36969;
  assign n36971 = pi681 & ~n17425;
  assign n36972 = n6223 & ~n16775;
  assign n36973 = ~n36971 & n36972;
  assign n36974 = pi681 & ~n36329;
  assign n36975 = ~pi681 & ~n16785;
  assign n36976 = ~n6223 & ~n36974;
  assign n36977 = ~n36975 & n36976;
  assign n36978 = pi223 & ~n36977;
  assign n36979 = ~n36973 & n36978;
  assign n36980 = pi681 & n17392;
  assign n36981 = ~n6223 & ~n36980;
  assign n36982 = ~n17386 & n36954;
  assign n36983 = n6223 & ~n36982;
  assign n36984 = ~pi223 & ~n36981;
  assign n36985 = ~n36983 & n36984;
  assign n36986 = ~n3461 & ~n36985;
  assign n36987 = ~n36979 & n36986;
  assign n36988 = ~n36970 & ~n36987;
  assign n36989 = ~pi215 & ~n36988;
  assign n36990 = pi681 & ~n17448;
  assign n36991 = ~n16703 & ~n36990;
  assign n36992 = ~n6223 & n36991;
  assign n36993 = pi681 & ~n36348;
  assign n36994 = ~n16725 & ~n36993;
  assign n36995 = n6223 & n36994;
  assign n36996 = pi223 & ~n36995;
  assign n36997 = ~n36992 & n36996;
  assign n36998 = ~pi223 & pi681;
  assign n36999 = n17414 & n36998;
  assign n37000 = pi215 & ~n36999;
  assign n37001 = ~n36997 & n37000;
  assign n37002 = pi299 & ~n37001;
  assign n37003 = ~n36989 & n37002;
  assign n37004 = n3053 & ~n36969;
  assign n37005 = n6197 & n36982;
  assign n37006 = ~n6197 & n36980;
  assign n37007 = ~n3053 & ~n37005;
  assign n37008 = ~n37006 & n37007;
  assign n37009 = ~n37004 & ~n37008;
  assign n37010 = ~pi223 & ~n37009;
  assign n37011 = ~n6197 & ~n36991;
  assign n37012 = n6197 & ~n36994;
  assign n37013 = pi223 & ~n37012;
  assign n37014 = ~n37011 & n37013;
  assign n37015 = ~pi299 & ~n37014;
  assign n37016 = ~n37010 & n37015;
  assign n37017 = pi39 & ~n37016;
  assign n37018 = ~n37003 & n37017;
  assign n37019 = ~n36968 & ~n37018;
  assign n37020 = ~pi38 & ~n37019;
  assign n37021 = pi681 & n17479;
  assign n37022 = pi223 & ~n16968;
  assign n37023 = pi38 & ~n37021;
  assign n37024 = ~n37022 & n37023;
  assign n37025 = n3268 & ~n37024;
  assign n37026 = ~n37020 & n37025;
  assign n37027 = ~n36766 & ~n37026;
  assign n37028 = ~pi778 & ~n37027;
  assign n37029 = pi625 & n37027;
  assign n37030 = ~pi625 & ~n36763;
  assign n37031 = pi1153 & ~n37030;
  assign n37032 = ~n37029 & n37031;
  assign n37033 = ~pi625 & n37027;
  assign n37034 = pi625 & ~n36763;
  assign n37035 = ~pi1153 & ~n37034;
  assign n37036 = ~n37033 & n37035;
  assign n37037 = ~n37032 & ~n37036;
  assign n37038 = pi778 & ~n37037;
  assign n37039 = ~n37028 & ~n37038;
  assign n37040 = ~n17554 & n37039;
  assign n37041 = ~n36953 & ~n37040;
  assign n37042 = ~n17591 & n37041;
  assign n37043 = n17591 & n36763;
  assign n37044 = ~n37042 & ~n37043;
  assign n37045 = ~n17627 & n37044;
  assign n37046 = ~n17670 & n37045;
  assign n37047 = ~n36952 & ~n37046;
  assign n37048 = ~n19247 & ~n37047;
  assign n37049 = n17946 & ~n36763;
  assign n37050 = ~n37048 & ~n37049;
  assign n37051 = pi647 & ~n37050;
  assign n37052 = ~pi647 & ~n36763;
  assign n37053 = pi1157 & ~n37052;
  assign n37054 = ~n37051 & n37053;
  assign n37055 = ~pi630 & n37054;
  assign n37056 = ~pi647 & ~n37050;
  assign n37057 = pi647 & ~n36763;
  assign n37058 = ~pi1157 & ~n37057;
  assign n37059 = ~n37056 & n37058;
  assign n37060 = pi630 & n37059;
  assign n37061 = ~n37055 & ~n37060;
  assign n37062 = ~n36951 & n37061;
  assign n37063 = pi787 & ~n37062;
  assign n37064 = ~n20502 & n36947;
  assign n37065 = ~pi628 & ~n37047;
  assign n37066 = pi628 & ~n36763;
  assign n37067 = n17696 & ~n37066;
  assign n37068 = ~n37065 & n37067;
  assign n37069 = pi628 & ~n37047;
  assign n37070 = ~pi628 & ~n36763;
  assign n37071 = n17695 & ~n37070;
  assign n37072 = ~n37069 & n37071;
  assign n37073 = ~n37068 & ~n37072;
  assign n37074 = ~n37064 & n37073;
  assign n37075 = pi792 & ~n37074;
  assign n37076 = pi626 & ~n36945;
  assign n37077 = ~pi626 & n36763;
  assign n37078 = n17667 & ~n37077;
  assign n37079 = ~n37076 & n37078;
  assign n37080 = ~pi626 & ~n36945;
  assign n37081 = pi626 & n36763;
  assign n37082 = n17668 & ~n37081;
  assign n37083 = ~n37080 & n37082;
  assign n37084 = n17627 & ~n36763;
  assign n37085 = ~n37045 & ~n37084;
  assign n37086 = n17792 & ~n37085;
  assign n37087 = ~n37079 & ~n37086;
  assign n37088 = ~n37083 & n37087;
  assign n37089 = pi788 & ~n37088;
  assign n37090 = ~pi680 & ~n36794;
  assign n37091 = ~pi642 & ~n16978;
  assign n37092 = ~n17181 & ~n37091;
  assign n37093 = n35763 & n37092;
  assign n37094 = pi680 & ~n37093;
  assign n37095 = pi642 & ~n17182;
  assign n37096 = n6164 & ~n37095;
  assign n37097 = ~pi642 & ~n17110;
  assign n37098 = n37096 & ~n37097;
  assign n37099 = n37094 & ~n37098;
  assign n37100 = ~n37090 & ~n37099;
  assign n37101 = pi681 & ~n37100;
  assign n37102 = ~n36799 & ~n37101;
  assign n37103 = n6223 & ~n37102;
  assign n37104 = ~n36804 & ~n36954;
  assign n37105 = ~pi642 & ~n6164;
  assign n37106 = ~n17085 & n37105;
  assign n37107 = pi642 & n17173;
  assign n37108 = pi680 & ~n37107;
  assign n37109 = ~n17092 & n37108;
  assign n37110 = ~n37106 & n37109;
  assign n37111 = ~n37104 & ~n37110;
  assign n37112 = ~n36808 & ~n37111;
  assign n37113 = ~n6223 & ~n37112;
  assign n37114 = ~pi223 & ~n37103;
  assign n37115 = ~n37113 & n37114;
  assign n37116 = ~n36773 & ~n36954;
  assign n37117 = n16665 & ~n37092;
  assign n37118 = ~n16658 & n37117;
  assign n37119 = ~n6164 & ~n37118;
  assign n37120 = pi680 & ~n37119;
  assign n37121 = pi642 & ~n17247;
  assign n37122 = ~n17021 & ~n37121;
  assign n37123 = n6164 & ~n37122;
  assign n37124 = n37120 & ~n37123;
  assign n37125 = ~n37116 & ~n37124;
  assign n37126 = n36779 & ~n37125;
  assign n37127 = ~n36784 & ~n36954;
  assign n37128 = n16854 & ~n36435;
  assign n37129 = n36437 & n37105;
  assign n37130 = pi642 & ~n36442;
  assign n37131 = pi680 & ~n37130;
  assign n37132 = ~n37128 & n37131;
  assign n37133 = ~n37129 & n37132;
  assign n37134 = ~n37127 & ~n37133;
  assign n37135 = n36790 & ~n37134;
  assign n37136 = pi223 & ~n37135;
  assign n37137 = ~n37126 & n37136;
  assign n37138 = ~n3461 & ~n37137;
  assign n37139 = ~n37115 & n37138;
  assign n37140 = n36767 & ~n36954;
  assign n37141 = n36954 & ~n37091;
  assign n37142 = ~n36603 & n37141;
  assign n37143 = ~n37140 & ~n37142;
  assign n37144 = n16661 & ~n37143;
  assign n37145 = ~pi223 & n37144;
  assign n37146 = n36846 & ~n36954;
  assign n37147 = n36954 & n37117;
  assign n37148 = pi223 & ~n37146;
  assign n37149 = ~n37147 & n37148;
  assign n37150 = n36819 & ~n37149;
  assign n37151 = ~n37145 & n37150;
  assign n37152 = ~pi215 & ~n37151;
  assign n37153 = ~n37139 & n37152;
  assign n37154 = ~n36844 & ~n36954;
  assign n37155 = ~pi614 & n16995;
  assign n37156 = ~n37121 & ~n37155;
  assign n37157 = ~pi616 & ~n37156;
  assign n37158 = n37120 & ~n37157;
  assign n37159 = ~n37154 & ~n37158;
  assign n37160 = ~n36850 & ~n37159;
  assign n37161 = n6223 & ~n37160;
  assign n37162 = ~pi680 & n36855;
  assign n37163 = ~n6164 & n17011;
  assign n37164 = pi642 & ~n36510;
  assign n37165 = pi680 & ~n17012;
  assign n37166 = ~n37164 & n37165;
  assign n37167 = ~n37163 & n37166;
  assign n37168 = pi681 & ~n37167;
  assign n37169 = ~n37162 & n37168;
  assign n37170 = ~n36857 & ~n37169;
  assign n37171 = ~n6223 & ~n37170;
  assign n37172 = pi223 & ~n37171;
  assign n37173 = ~n37161 & n37172;
  assign n37174 = ~n17128 & n37096;
  assign n37175 = n37094 & ~n37174;
  assign n37176 = ~n37090 & ~n37175;
  assign n37177 = pi681 & ~n37176;
  assign n37178 = n36835 & ~n37177;
  assign n37179 = ~n36832 & ~n36954;
  assign n37180 = n17127 & n17211;
  assign n37181 = n16854 & ~n37180;
  assign n37182 = ~n17123 & n37105;
  assign n37183 = pi642 & n36522;
  assign n37184 = pi680 & ~n37182;
  assign n37185 = ~n37183 & n37184;
  assign n37186 = ~n37181 & n37185;
  assign n37187 = ~n37179 & ~n37186;
  assign n37188 = ~n6223 & n36830;
  assign n37189 = ~n37187 & n37188;
  assign n37190 = ~pi223 & ~n37178;
  assign n37191 = ~n37189 & n37190;
  assign n37192 = pi215 & ~n37191;
  assign n37193 = ~n37173 & n37192;
  assign n37194 = pi299 & ~n37193;
  assign n37195 = ~n37153 & n37194;
  assign n37196 = ~n6197 & n37112;
  assign n37197 = n6197 & n37102;
  assign n37198 = ~n3053 & ~n37196;
  assign n37199 = ~n37197 & n37198;
  assign n37200 = n3053 & ~n37144;
  assign n37201 = ~pi223 & ~n37200;
  assign n37202 = ~n37199 & n37201;
  assign n37203 = n6197 & n37160;
  assign n37204 = ~n6197 & n37170;
  assign n37205 = pi223 & ~n37204;
  assign n37206 = ~n37203 & n37205;
  assign n37207 = ~pi299 & ~n37206;
  assign n37208 = ~n37202 & n37207;
  assign n37209 = pi39 & ~n37208;
  assign n37210 = ~n37195 & n37209;
  assign n37211 = n17329 & ~n36954;
  assign n37212 = ~n36581 & n36886;
  assign n37213 = ~n37211 & n37212;
  assign n37214 = n17330 & n36998;
  assign n37215 = n36884 & ~n37214;
  assign n37216 = ~n37213 & n37215;
  assign n37217 = n17338 & n36998;
  assign n37218 = n17337 & ~n36954;
  assign n37219 = ~n36589 & n36892;
  assign n37220 = ~n37218 & n37219;
  assign n37221 = n36890 & ~n37217;
  assign n37222 = ~n37220 & n37221;
  assign n37223 = ~pi39 & ~n37216;
  assign n37224 = ~n37222 & n37223;
  assign n37225 = ~pi38 & ~n37224;
  assign n37226 = ~n37210 & n37225;
  assign n37227 = n37143 & ~n37149;
  assign n37228 = n36902 & ~n37227;
  assign n37229 = n36900 & ~n37228;
  assign n37230 = n3268 & ~n37229;
  assign n37231 = ~n37226 & n37230;
  assign n37232 = ~n36766 & ~n37231;
  assign n37233 = ~pi625 & n37232;
  assign n37234 = pi625 & n36907;
  assign n37235 = ~pi1153 & ~n37234;
  assign n37236 = ~n37233 & n37235;
  assign n37237 = ~pi608 & ~n37236;
  assign n37238 = ~n37032 & n37237;
  assign n37239 = pi625 & n37232;
  assign n37240 = ~pi625 & n36907;
  assign n37241 = pi1153 & ~n37240;
  assign n37242 = ~n37239 & n37241;
  assign n37243 = pi608 & ~n37242;
  assign n37244 = ~n37036 & n37243;
  assign n37245 = ~n37238 & ~n37244;
  assign n37246 = pi778 & ~n37245;
  assign n37247 = ~pi778 & n37232;
  assign n37248 = ~n37246 & ~n37247;
  assign n37249 = ~pi609 & ~n37248;
  assign n37250 = pi609 & n37039;
  assign n37251 = ~pi1155 & ~n37250;
  assign n37252 = ~n37249 & n37251;
  assign n37253 = ~pi660 & ~n36914;
  assign n37254 = ~n37252 & n37253;
  assign n37255 = pi609 & ~n37248;
  assign n37256 = ~pi609 & n37039;
  assign n37257 = pi1155 & ~n37256;
  assign n37258 = ~n37255 & n37257;
  assign n37259 = pi660 & ~n36918;
  assign n37260 = ~n37258 & n37259;
  assign n37261 = ~n37254 & ~n37260;
  assign n37262 = pi785 & ~n37261;
  assign n37263 = ~pi785 & ~n37248;
  assign n37264 = ~n37262 & ~n37263;
  assign n37265 = ~pi618 & ~n37264;
  assign n37266 = pi618 & ~n37041;
  assign n37267 = ~pi1154 & ~n37266;
  assign n37268 = ~n37265 & n37267;
  assign n37269 = ~pi627 & ~n36926;
  assign n37270 = ~n37268 & n37269;
  assign n37271 = pi618 & ~n37264;
  assign n37272 = ~pi618 & ~n37041;
  assign n37273 = pi1154 & ~n37272;
  assign n37274 = ~n37271 & n37273;
  assign n37275 = pi627 & ~n36930;
  assign n37276 = ~n37274 & n37275;
  assign n37277 = ~n37270 & ~n37276;
  assign n37278 = pi781 & ~n37277;
  assign n37279 = ~pi781 & ~n37264;
  assign n37280 = ~n37278 & ~n37279;
  assign n37281 = ~pi619 & ~n37280;
  assign n37282 = pi619 & n37044;
  assign n37283 = ~pi1159 & ~n37282;
  assign n37284 = ~n37281 & n37283;
  assign n37285 = ~pi648 & ~n36938;
  assign n37286 = ~n37284 & n37285;
  assign n37287 = pi619 & ~n37280;
  assign n37288 = ~pi619 & n37044;
  assign n37289 = pi1159 & ~n37288;
  assign n37290 = ~n37287 & n37289;
  assign n37291 = pi648 & ~n36942;
  assign n37292 = ~n37290 & n37291;
  assign n37293 = pi789 & ~n37286;
  assign n37294 = ~n37292 & n37293;
  assign n37295 = ~pi789 & n37280;
  assign n37296 = n17905 & ~n37295;
  assign n37297 = ~n37294 & n37296;
  assign n37298 = ~n37089 & ~n37297;
  assign n37299 = ~n37075 & ~n37298;
  assign n37300 = n20298 & n37074;
  assign n37301 = n20300 & ~n37300;
  assign n37302 = ~n37299 & n37301;
  assign n37303 = ~n37063 & ~n37302;
  assign n37304 = pi644 & n37303;
  assign n37305 = ~pi787 & n37050;
  assign n37306 = ~n37054 & ~n37059;
  assign n37307 = pi787 & ~n37306;
  assign n37308 = ~n37305 & ~n37307;
  assign n37309 = ~pi644 & n37308;
  assign n37310 = pi715 & ~n37309;
  assign n37311 = ~n37304 & n37310;
  assign n37312 = n17740 & ~n36763;
  assign n37313 = ~n17740 & n36950;
  assign n37314 = ~n37312 & ~n37313;
  assign n37315 = pi644 & ~n37314;
  assign n37316 = ~pi644 & ~n36763;
  assign n37317 = ~pi715 & ~n37316;
  assign n37318 = ~n37315 & n37317;
  assign n37319 = pi1160 & ~n37318;
  assign n37320 = ~n37311 & n37319;
  assign n37321 = ~pi644 & n37303;
  assign n37322 = pi644 & n37308;
  assign n37323 = ~pi715 & ~n37322;
  assign n37324 = ~n37321 & n37323;
  assign n37325 = ~pi644 & ~n37314;
  assign n37326 = pi644 & ~n36763;
  assign n37327 = pi715 & ~n37326;
  assign n37328 = ~n37325 & n37327;
  assign n37329 = ~pi1160 & ~n37328;
  assign n37330 = ~n37324 & n37329;
  assign n37331 = ~n37320 & ~n37330;
  assign n37332 = pi790 & ~n37331;
  assign n37333 = ~pi790 & n37303;
  assign n37334 = ~n37332 & ~n37333;
  assign n37335 = ~po1038 & ~n37334;
  assign n37336 = ~pi223 & po1038;
  assign po380 = ~n37335 & ~n37336;
  assign n37338 = pi224 & ~n36142;
  assign n37339 = n17904 & ~n37338;
  assign n37340 = pi224 & ~n3268;
  assign n37341 = pi614 & n16842;
  assign n37342 = n16661 & ~n37341;
  assign n37343 = ~n6165 & ~n37342;
  assign n37344 = ~n16757 & ~n37343;
  assign n37345 = ~n16708 & ~n37344;
  assign n37346 = ~pi680 & ~n37344;
  assign n37347 = pi680 & n37341;
  assign n37348 = ~n16767 & ~n37347;
  assign n37349 = ~n37346 & n37348;
  assign n37350 = n16708 & ~n37349;
  assign n37351 = ~n37345 & ~n37350;
  assign n37352 = n6223 & n37351;
  assign n37353 = pi614 & ~n17084;
  assign n37354 = n6164 & ~n16782;
  assign n37355 = ~pi614 & pi616;
  assign n37356 = n16779 & n37355;
  assign n37357 = ~n37353 & ~n37356;
  assign n37358 = ~n37354 & n37357;
  assign n37359 = ~n16708 & ~n37358;
  assign n37360 = ~pi680 & ~n37358;
  assign n37361 = pi614 & n17044;
  assign n37362 = pi680 & ~n37361;
  assign n37363 = n16748 & n37362;
  assign n37364 = ~n37347 & ~n37363;
  assign n37365 = ~n37360 & n37364;
  assign n37366 = n16708 & ~n37365;
  assign n37367 = ~n37359 & ~n37366;
  assign n37368 = ~n6223 & n37367;
  assign n37369 = pi224 & ~n37368;
  assign n37370 = ~n37352 & n37369;
  assign n37371 = ~n16779 & n37341;
  assign n37372 = ~pi680 & ~n37371;
  assign n37373 = ~n37362 & ~n37372;
  assign n37374 = n16708 & ~n37373;
  assign n37375 = ~n16708 & ~n37371;
  assign n37376 = ~n37374 & ~n37375;
  assign n37377 = ~n6223 & ~n37376;
  assign n37378 = pi614 & ~n36172;
  assign n37379 = n6223 & ~n37378;
  assign n37380 = ~pi224 & ~n37379;
  assign n37381 = ~n37377 & n37380;
  assign n37382 = ~n3461 & ~n37381;
  assign n37383 = ~n37370 & n37382;
  assign n37384 = pi224 & ~n16661;
  assign n37385 = n3461 & ~n37384;
  assign n37386 = n16771 & n16842;
  assign n37387 = n37385 & ~n37386;
  assign n37388 = ~pi215 & ~n37387;
  assign n37389 = ~n37383 & n37388;
  assign n37390 = pi614 & ~n36194;
  assign n37391 = ~pi224 & n37390;
  assign n37392 = ~n16944 & n37391;
  assign n37393 = ~n16693 & ~n37343;
  assign n37394 = ~n16708 & ~n37393;
  assign n37395 = ~pi680 & ~n37393;
  assign n37396 = ~n16712 & ~n37347;
  assign n37397 = ~n37395 & n37396;
  assign n37398 = n16708 & ~n37397;
  assign n37399 = ~n37394 & ~n37398;
  assign n37400 = n6223 & n37399;
  assign n37401 = pi614 & ~n16880;
  assign n37402 = ~n35884 & ~n37401;
  assign n37403 = ~pi680 & ~n37402;
  assign n37404 = pi680 & ~n16884;
  assign n37405 = ~n35886 & n37404;
  assign n37406 = ~n37403 & ~n37405;
  assign n37407 = n16708 & ~n37406;
  assign n37408 = ~n16708 & ~n37402;
  assign n37409 = ~n37407 & ~n37408;
  assign n37410 = ~n6223 & n37409;
  assign n37411 = pi224 & ~n37410;
  assign n37412 = ~n37400 & n37411;
  assign n37413 = ~n37392 & ~n37412;
  assign n37414 = pi215 & ~n37413;
  assign n37415 = pi299 & ~n37414;
  assign n37416 = ~n37389 & n37415;
  assign n37417 = n6197 & n37399;
  assign n37418 = ~n6197 & n37409;
  assign n37419 = pi224 & ~n37418;
  assign n37420 = ~n37417 & n37419;
  assign n37421 = ~n16956 & n37391;
  assign n37422 = pi223 & ~n37421;
  assign n37423 = ~n37420 & n37422;
  assign n37424 = n6197 & n37351;
  assign n37425 = ~n6197 & n37367;
  assign n37426 = pi224 & ~n37425;
  assign n37427 = ~n37424 & n37426;
  assign n37428 = ~n6197 & ~n37376;
  assign n37429 = n6197 & ~n37378;
  assign n37430 = n5777 & ~n37429;
  assign n37431 = ~n37428 & n37430;
  assign n37432 = pi614 & n16949;
  assign n37433 = ~pi223 & ~n37432;
  assign n37434 = ~n37431 & n37433;
  assign n37435 = ~n37427 & n37434;
  assign n37436 = ~n37423 & ~n37435;
  assign n37437 = ~pi299 & ~n37436;
  assign n37438 = pi39 & ~n37416;
  assign n37439 = ~n37437 & n37438;
  assign n37440 = ~pi614 & n16911;
  assign n37441 = pi224 & ~n37440;
  assign n37442 = n16837 & n37441;
  assign n37443 = pi614 & n16911;
  assign n37444 = ~pi224 & n37443;
  assign n37445 = ~pi299 & ~n37444;
  assign n37446 = ~n37442 & n37445;
  assign n37447 = pi614 & n16916;
  assign n37448 = pi224 & n16822;
  assign n37449 = n37447 & ~n37448;
  assign n37450 = pi224 & ~n16649;
  assign n37451 = ~n37449 & ~n37450;
  assign n37452 = pi299 & n37451;
  assign n37453 = ~pi39 & ~n37446;
  assign n37454 = ~n37452 & n37453;
  assign n37455 = ~pi38 & ~n37454;
  assign n37456 = ~n37439 & n37455;
  assign n37457 = pi224 & ~n16968;
  assign n37458 = pi38 & ~n37457;
  assign n37459 = pi614 & n16970;
  assign n37460 = n37458 & ~n37459;
  assign n37461 = n3268 & ~n37460;
  assign n37462 = ~n37456 & n37461;
  assign n37463 = ~n37340 & ~n37462;
  assign n37464 = ~n17526 & ~n37463;
  assign n37465 = n17526 & n37338;
  assign n37466 = ~n37464 & ~n37465;
  assign n37467 = ~pi785 & ~n37466;
  assign n37468 = pi609 & n37466;
  assign n37469 = ~pi609 & ~n37338;
  assign n37470 = pi1155 & ~n37469;
  assign n37471 = ~n37468 & n37470;
  assign n37472 = ~pi609 & n37466;
  assign n37473 = pi609 & ~n37338;
  assign n37474 = ~pi1155 & ~n37473;
  assign n37475 = ~n37472 & n37474;
  assign n37476 = ~n37471 & ~n37475;
  assign n37477 = pi785 & ~n37476;
  assign n37478 = ~n37467 & ~n37477;
  assign n37479 = ~pi781 & ~n37478;
  assign n37480 = pi618 & n37478;
  assign n37481 = ~pi618 & ~n37338;
  assign n37482 = pi1154 & ~n37481;
  assign n37483 = ~n37480 & n37482;
  assign n37484 = ~pi618 & n37478;
  assign n37485 = pi618 & ~n37338;
  assign n37486 = ~pi1154 & ~n37485;
  assign n37487 = ~n37484 & n37486;
  assign n37488 = ~n37483 & ~n37487;
  assign n37489 = pi781 & ~n37488;
  assign n37490 = ~n37479 & ~n37489;
  assign n37491 = ~pi789 & ~n37490;
  assign n37492 = pi619 & n37490;
  assign n37493 = ~pi619 & ~n37338;
  assign n37494 = pi1159 & ~n37493;
  assign n37495 = ~n37492 & n37494;
  assign n37496 = ~pi619 & n37490;
  assign n37497 = pi619 & ~n37338;
  assign n37498 = ~pi1159 & ~n37497;
  assign n37499 = ~n37496 & n37498;
  assign n37500 = ~n37495 & ~n37499;
  assign n37501 = pi789 & ~n37500;
  assign n37502 = ~n37491 & ~n37501;
  assign n37503 = ~n17904 & n37502;
  assign n37504 = ~n37339 & ~n37503;
  assign n37505 = ~n20502 & n37504;
  assign n37506 = ~n19215 & ~n37338;
  assign n37507 = pi662 & pi680;
  assign n37508 = n17325 & ~n37507;
  assign n37509 = ~pi224 & ~n17325;
  assign n37510 = pi224 & n17305;
  assign n37511 = ~pi299 & ~n37510;
  assign n37512 = ~n37508 & n37511;
  assign n37513 = ~n37509 & n37512;
  assign n37514 = n17334 & ~n37507;
  assign n37515 = ~pi224 & ~n17334;
  assign n37516 = pi224 & n17311;
  assign n37517 = pi299 & ~n37516;
  assign n37518 = ~n37514 & n37517;
  assign n37519 = ~n37515 & n37518;
  assign n37520 = ~pi39 & ~n37513;
  assign n37521 = ~n37519 & n37520;
  assign n37522 = n17076 & n37507;
  assign n37523 = n37385 & ~n37522;
  assign n37524 = pi662 & ~n17425;
  assign n37525 = ~pi662 & ~n16776;
  assign n37526 = ~n37524 & ~n37525;
  assign n37527 = n6223 & n37526;
  assign n37528 = ~n6166 & ~n36329;
  assign n37529 = n16785 & ~n37528;
  assign n37530 = ~n6223 & n37529;
  assign n37531 = pi224 & ~n37530;
  assign n37532 = ~n37527 & n37531;
  assign n37533 = pi662 & n17392;
  assign n37534 = ~n6223 & ~n37533;
  assign n37535 = ~n17386 & n37507;
  assign n37536 = n6223 & ~n37535;
  assign n37537 = ~pi224 & ~n37534;
  assign n37538 = ~n37536 & n37537;
  assign n37539 = ~n3461 & ~n37538;
  assign n37540 = ~n37532 & n37539;
  assign n37541 = ~n37523 & ~n37540;
  assign n37542 = ~pi215 & ~n37541;
  assign n37543 = ~pi662 & ~n16704;
  assign n37544 = pi662 & ~n17448;
  assign n37545 = ~n37543 & ~n37544;
  assign n37546 = ~n6223 & n37545;
  assign n37547 = ~pi662 & ~n16726;
  assign n37548 = pi662 & ~n36348;
  assign n37549 = ~n37547 & ~n37548;
  assign n37550 = n6223 & n37549;
  assign n37551 = pi224 & ~n37550;
  assign n37552 = ~n37546 & n37551;
  assign n37553 = ~pi224 & pi662;
  assign n37554 = n17414 & n37553;
  assign n37555 = pi215 & ~n37554;
  assign n37556 = ~n37552 & n37555;
  assign n37557 = pi299 & ~n37556;
  assign n37558 = ~n37542 & n37557;
  assign n37559 = n6197 & n37526;
  assign n37560 = ~n6197 & n37529;
  assign n37561 = pi224 & ~n37560;
  assign n37562 = ~n37559 & n37561;
  assign n37563 = ~n6197 & ~n37533;
  assign n37564 = n6197 & ~n37535;
  assign n37565 = n5777 & ~n37563;
  assign n37566 = ~n37564 & n37565;
  assign n37567 = pi662 & n17384;
  assign n37568 = ~pi223 & ~n37567;
  assign n37569 = ~n37566 & n37568;
  assign n37570 = ~n37562 & n37569;
  assign n37571 = ~n6197 & n37545;
  assign n37572 = n6197 & n37549;
  assign n37573 = pi224 & ~n37572;
  assign n37574 = ~n37571 & n37573;
  assign n37575 = n17401 & n37553;
  assign n37576 = pi223 & ~n37575;
  assign n37577 = ~n37574 & n37576;
  assign n37578 = ~pi299 & ~n37577;
  assign n37579 = ~n37570 & n37578;
  assign n37580 = pi39 & ~n37579;
  assign n37581 = ~n37558 & n37580;
  assign n37582 = ~n37521 & ~n37581;
  assign n37583 = ~pi38 & ~n37582;
  assign n37584 = pi662 & n17479;
  assign n37585 = n37458 & ~n37584;
  assign n37586 = n3268 & ~n37585;
  assign n37587 = ~n37583 & n37586;
  assign n37588 = ~n37340 & ~n37587;
  assign n37589 = ~pi778 & ~n37588;
  assign n37590 = pi625 & n37588;
  assign n37591 = ~pi625 & ~n37338;
  assign n37592 = pi1153 & ~n37591;
  assign n37593 = ~n37590 & n37592;
  assign n37594 = ~pi625 & n37588;
  assign n37595 = pi625 & ~n37338;
  assign n37596 = ~pi1153 & ~n37595;
  assign n37597 = ~n37594 & n37596;
  assign n37598 = ~n37593 & ~n37597;
  assign n37599 = pi778 & ~n37598;
  assign n37600 = ~n37589 & ~n37599;
  assign n37601 = ~n17554 & ~n37600;
  assign n37602 = n17554 & n37338;
  assign n37603 = ~n37601 & ~n37602;
  assign n37604 = ~n17591 & ~n37603;
  assign n37605 = n17591 & n37338;
  assign n37606 = ~n37604 & ~n37605;
  assign n37607 = ~n17627 & n37606;
  assign n37608 = ~n17670 & n37607;
  assign n37609 = ~n37506 & ~n37608;
  assign n37610 = ~pi628 & ~n37609;
  assign n37611 = pi628 & ~n37338;
  assign n37612 = n17696 & ~n37611;
  assign n37613 = ~n37610 & n37612;
  assign n37614 = pi628 & ~n37609;
  assign n37615 = ~pi628 & ~n37338;
  assign n37616 = n17695 & ~n37615;
  assign n37617 = ~n37614 & n37616;
  assign n37618 = ~n37613 & ~n37617;
  assign n37619 = ~n37505 & n37618;
  assign n37620 = pi792 & ~n37619;
  assign n37621 = ~pi614 & ~n24006;
  assign n37622 = pi614 & ~n36603;
  assign n37623 = ~n37621 & ~n37622;
  assign n37624 = ~n16658 & n37623;
  assign n37625 = pi616 & ~n37624;
  assign n37626 = pi614 & ~n17247;
  assign n37627 = ~n17023 & ~n37626;
  assign n37628 = ~pi616 & ~n37627;
  assign n37629 = ~n37625 & ~n37628;
  assign n37630 = pi680 & ~n37629;
  assign n37631 = ~n37346 & ~n37630;
  assign n37632 = pi662 & ~n37631;
  assign n37633 = ~pi662 & ~n16707;
  assign n37634 = ~n37344 & n37633;
  assign n37635 = ~n37350 & ~n37634;
  assign n37636 = ~n37632 & n37635;
  assign n37637 = pi224 & n37636;
  assign n37638 = ~n17104 & n37355;
  assign n37639 = ~n36476 & ~n37638;
  assign n37640 = pi680 & ~n37639;
  assign n37641 = ~n36477 & ~n37386;
  assign n37642 = ~n37640 & ~n37641;
  assign n37643 = pi662 & ~n37642;
  assign n37644 = ~pi662 & ~n37378;
  assign n37645 = ~n37643 & ~n37644;
  assign n37646 = ~pi224 & ~n37645;
  assign n37647 = n6223 & ~n37646;
  assign n37648 = ~n37637 & n37647;
  assign n37649 = ~pi614 & n17097;
  assign n37650 = pi614 & ~n17173;
  assign n37651 = pi680 & ~n37650;
  assign n37652 = ~n37649 & n37651;
  assign n37653 = ~n37372 & ~n37652;
  assign n37654 = pi662 & ~n37653;
  assign n37655 = ~n37371 & n37633;
  assign n37656 = ~n37374 & ~n37655;
  assign n37657 = ~n37654 & n37656;
  assign n37658 = ~pi224 & ~n37657;
  assign n37659 = pi614 & ~n36442;
  assign n37660 = n36437 & n37355;
  assign n37661 = ~n37659 & ~n37660;
  assign n37662 = ~n36440 & n37661;
  assign n37663 = pi680 & ~n37662;
  assign n37664 = ~n37360 & ~n37663;
  assign n37665 = pi662 & ~n37664;
  assign n37666 = ~n37358 & n37633;
  assign n37667 = ~n37366 & ~n37666;
  assign n37668 = ~n37665 & n37667;
  assign n37669 = pi224 & n37668;
  assign n37670 = ~n6223 & ~n37669;
  assign n37671 = ~n37658 & n37670;
  assign n37672 = ~n3461 & ~n37671;
  assign n37673 = ~n37648 & n37672;
  assign n37674 = n17104 & n37507;
  assign n37675 = ~n37386 & ~n37674;
  assign n37676 = ~pi224 & ~n37675;
  assign n37677 = n37507 & n37623;
  assign n37678 = ~n37341 & ~n37507;
  assign n37679 = n16665 & n37678;
  assign n37680 = pi224 & ~n37679;
  assign n37681 = ~n37677 & n37680;
  assign n37682 = n37385 & ~n37681;
  assign n37683 = ~n37676 & n37682;
  assign n37684 = ~pi215 & ~n37683;
  assign n37685 = ~n37673 & n37684;
  assign n37686 = ~n16997 & ~n37626;
  assign n37687 = ~pi616 & ~n37686;
  assign n37688 = ~n37625 & ~n37687;
  assign n37689 = pi680 & ~n37688;
  assign n37690 = ~n37395 & ~n37689;
  assign n37691 = pi662 & ~n37690;
  assign n37692 = ~n37393 & n37633;
  assign n37693 = ~n37398 & ~n37692;
  assign n37694 = ~n37691 & n37693;
  assign n37695 = n6223 & ~n37694;
  assign n37696 = pi614 & ~n36510;
  assign n37697 = n17013 & ~n37696;
  assign n37698 = pi680 & ~n37697;
  assign n37699 = ~n37403 & ~n37698;
  assign n37700 = pi662 & ~n37699;
  assign n37701 = ~n37402 & n37633;
  assign n37702 = ~n37407 & ~n37701;
  assign n37703 = ~n37700 & n37702;
  assign n37704 = ~n6223 & ~n37703;
  assign n37705 = pi224 & ~n37704;
  assign n37706 = ~n37695 & n37705;
  assign n37707 = pi680 & ~n17139;
  assign n37708 = ~n37386 & ~n37707;
  assign n37709 = ~n37640 & ~n37708;
  assign n37710 = pi662 & ~n37709;
  assign n37711 = ~pi662 & ~n37390;
  assign n37712 = ~n37710 & ~n37711;
  assign n37713 = n6223 & n37712;
  assign n37714 = ~n16679 & n37390;
  assign n37715 = ~pi662 & ~n37714;
  assign n37716 = ~pi614 & n17124;
  assign n37717 = pi614 & n36522;
  assign n37718 = pi680 & ~n37717;
  assign n37719 = ~n37716 & n37718;
  assign n37720 = ~n17130 & n37719;
  assign n37721 = pi614 & ~pi680;
  assign n37722 = n16939 & n37721;
  assign n37723 = pi662 & ~n37722;
  assign n37724 = ~n37720 & n37723;
  assign n37725 = ~n37715 & ~n37724;
  assign n37726 = ~n6223 & n37725;
  assign n37727 = ~pi224 & ~n37726;
  assign n37728 = ~n37713 & n37727;
  assign n37729 = pi215 & ~n37728;
  assign n37730 = ~n37706 & n37729;
  assign n37731 = pi299 & ~n37730;
  assign n37732 = ~n37685 & n37731;
  assign n37733 = n6197 & n37636;
  assign n37734 = ~n6197 & n37668;
  assign n37735 = pi224 & ~n37734;
  assign n37736 = ~n37733 & n37735;
  assign n37737 = ~n6197 & ~n37657;
  assign n37738 = n6197 & ~n37645;
  assign n37739 = n5777 & ~n37738;
  assign n37740 = ~n37737 & n37739;
  assign n37741 = ~pi222 & n37676;
  assign n37742 = ~pi223 & ~n37741;
  assign n37743 = ~n37740 & n37742;
  assign n37744 = ~n37736 & n37743;
  assign n37745 = pi224 & n37694;
  assign n37746 = ~pi224 & ~n37712;
  assign n37747 = n6197 & ~n37746;
  assign n37748 = ~n37745 & n37747;
  assign n37749 = pi224 & n37703;
  assign n37750 = ~pi224 & ~n37725;
  assign n37751 = ~n6197 & ~n37749;
  assign n37752 = ~n37750 & n37751;
  assign n37753 = pi223 & ~n37752;
  assign n37754 = ~n37748 & n37753;
  assign n37755 = ~n37744 & ~n37754;
  assign n37756 = ~pi299 & ~n37755;
  assign n37757 = pi39 & ~n37732;
  assign n37758 = ~n37756 & n37757;
  assign n37759 = n17329 & n37507;
  assign n37760 = ~n37443 & ~n37759;
  assign n37761 = ~pi224 & ~n37760;
  assign n37762 = n17329 & ~n37507;
  assign n37763 = ~n36581 & n37441;
  assign n37764 = ~n37762 & n37763;
  assign n37765 = ~n37761 & ~n37764;
  assign n37766 = ~pi299 & ~n37765;
  assign n37767 = ~pi614 & n16916;
  assign n37768 = ~n36589 & ~n37767;
  assign n37769 = pi224 & ~n37768;
  assign n37770 = ~pi224 & ~n17337;
  assign n37771 = ~n37447 & n37770;
  assign n37772 = ~n37769 & ~n37771;
  assign n37773 = n37507 & ~n37772;
  assign n37774 = n37451 & ~n37507;
  assign n37775 = pi299 & ~n37774;
  assign n37776 = ~n37773 & n37775;
  assign n37777 = ~n37766 & ~n37776;
  assign n37778 = ~pi39 & ~n37777;
  assign n37779 = ~pi38 & ~n37778;
  assign n37780 = ~n37758 & n37779;
  assign n37781 = pi662 & n17054;
  assign n37782 = n16968 & n37781;
  assign n37783 = n37460 & ~n37782;
  assign n37784 = n3268 & ~n37783;
  assign n37785 = ~n37780 & n37784;
  assign n37786 = ~n37340 & ~n37785;
  assign n37787 = ~pi625 & n37786;
  assign n37788 = pi625 & n37463;
  assign n37789 = ~pi1153 & ~n37788;
  assign n37790 = ~n37787 & n37789;
  assign n37791 = ~pi608 & ~n37593;
  assign n37792 = ~n37790 & n37791;
  assign n37793 = pi625 & n37786;
  assign n37794 = ~pi625 & n37463;
  assign n37795 = pi1153 & ~n37794;
  assign n37796 = ~n37793 & n37795;
  assign n37797 = pi608 & ~n37597;
  assign n37798 = ~n37796 & n37797;
  assign n37799 = ~n37792 & ~n37798;
  assign n37800 = pi778 & ~n37799;
  assign n37801 = ~pi778 & n37786;
  assign n37802 = ~n37800 & ~n37801;
  assign n37803 = ~pi609 & ~n37802;
  assign n37804 = pi609 & n37600;
  assign n37805 = ~pi1155 & ~n37804;
  assign n37806 = ~n37803 & n37805;
  assign n37807 = ~pi660 & ~n37471;
  assign n37808 = ~n37806 & n37807;
  assign n37809 = pi609 & ~n37802;
  assign n37810 = ~pi609 & n37600;
  assign n37811 = pi1155 & ~n37810;
  assign n37812 = ~n37809 & n37811;
  assign n37813 = pi660 & ~n37475;
  assign n37814 = ~n37812 & n37813;
  assign n37815 = ~n37808 & ~n37814;
  assign n37816 = pi785 & ~n37815;
  assign n37817 = ~pi785 & ~n37802;
  assign n37818 = ~n37816 & ~n37817;
  assign n37819 = ~pi618 & ~n37818;
  assign n37820 = pi618 & n37603;
  assign n37821 = ~pi1154 & ~n37820;
  assign n37822 = ~n37819 & n37821;
  assign n37823 = ~pi627 & ~n37483;
  assign n37824 = ~n37822 & n37823;
  assign n37825 = pi618 & ~n37818;
  assign n37826 = ~pi618 & n37603;
  assign n37827 = pi1154 & ~n37826;
  assign n37828 = ~n37825 & n37827;
  assign n37829 = pi627 & ~n37487;
  assign n37830 = ~n37828 & n37829;
  assign n37831 = ~n37824 & ~n37830;
  assign n37832 = pi781 & ~n37831;
  assign n37833 = ~pi781 & ~n37818;
  assign n37834 = ~n37832 & ~n37833;
  assign n37835 = ~pi619 & ~n37834;
  assign n37836 = pi619 & n37606;
  assign n37837 = ~pi1159 & ~n37836;
  assign n37838 = ~n37835 & n37837;
  assign n37839 = ~pi648 & ~n37495;
  assign n37840 = ~n37838 & n37839;
  assign n37841 = pi619 & ~n37834;
  assign n37842 = ~pi619 & n37606;
  assign n37843 = pi1159 & ~n37842;
  assign n37844 = ~n37841 & n37843;
  assign n37845 = pi648 & ~n37499;
  assign n37846 = ~n37844 & n37845;
  assign n37847 = pi789 & ~n37840;
  assign n37848 = ~n37846 & n37847;
  assign n37849 = ~pi789 & n37834;
  assign n37850 = n17905 & ~n37849;
  assign n37851 = ~n37848 & n37850;
  assign n37852 = pi626 & ~n37502;
  assign n37853 = ~pi626 & n37338;
  assign n37854 = n17667 & ~n37853;
  assign n37855 = ~n37852 & n37854;
  assign n37856 = ~pi626 & ~n37502;
  assign n37857 = pi626 & n37338;
  assign n37858 = n17668 & ~n37857;
  assign n37859 = ~n37856 & n37858;
  assign n37860 = n17627 & ~n37338;
  assign n37861 = ~n37607 & ~n37860;
  assign n37862 = n17792 & ~n37861;
  assign n37863 = ~n37855 & ~n37862;
  assign n37864 = ~n37859 & n37863;
  assign n37865 = pi788 & ~n37864;
  assign n37866 = ~n20298 & ~n37865;
  assign n37867 = ~n37851 & n37866;
  assign n37868 = ~n37620 & ~n37867;
  assign n37869 = n20300 & ~n37868;
  assign n37870 = ~n17698 & n37504;
  assign n37871 = n17698 & n37338;
  assign n37872 = ~n37870 & ~n37871;
  assign n37873 = ~n20491 & ~n37872;
  assign n37874 = ~n19247 & ~n37609;
  assign n37875 = n17946 & ~n37338;
  assign n37876 = ~n37874 & ~n37875;
  assign n37877 = pi647 & ~n37876;
  assign n37878 = ~pi647 & ~n37338;
  assign n37879 = pi1157 & ~n37878;
  assign n37880 = ~n37877 & n37879;
  assign n37881 = ~pi630 & n37880;
  assign n37882 = ~pi647 & ~n37876;
  assign n37883 = pi647 & ~n37338;
  assign n37884 = ~pi1157 & ~n37883;
  assign n37885 = ~n37882 & n37884;
  assign n37886 = pi630 & n37885;
  assign n37887 = ~n37881 & ~n37886;
  assign n37888 = ~n37873 & n37887;
  assign n37889 = pi787 & ~n37888;
  assign n37890 = ~n37869 & ~n37889;
  assign n37891 = pi644 & n37890;
  assign n37892 = ~pi787 & n37876;
  assign n37893 = ~n37880 & ~n37885;
  assign n37894 = pi787 & ~n37893;
  assign n37895 = ~n37892 & ~n37894;
  assign n37896 = ~pi644 & n37895;
  assign n37897 = pi715 & ~n37896;
  assign n37898 = ~n37891 & n37897;
  assign n37899 = n17740 & ~n37338;
  assign n37900 = ~n17740 & n37872;
  assign n37901 = ~n37899 & ~n37900;
  assign n37902 = pi644 & ~n37901;
  assign n37903 = ~pi644 & ~n37338;
  assign n37904 = ~pi715 & ~n37903;
  assign n37905 = ~n37902 & n37904;
  assign n37906 = pi1160 & ~n37905;
  assign n37907 = ~n37898 & n37906;
  assign n37908 = ~pi644 & n37890;
  assign n37909 = pi644 & n37895;
  assign n37910 = ~pi715 & ~n37909;
  assign n37911 = ~n37908 & n37910;
  assign n37912 = ~pi644 & ~n37901;
  assign n37913 = pi644 & ~n37338;
  assign n37914 = pi715 & ~n37913;
  assign n37915 = ~n37912 & n37914;
  assign n37916 = ~pi1160 & ~n37915;
  assign n37917 = ~n37911 & n37916;
  assign n37918 = ~n37907 & ~n37917;
  assign n37919 = pi790 & ~n37918;
  assign n37920 = ~pi790 & n37890;
  assign n37921 = ~n37919 & ~n37920;
  assign n37922 = ~po1038 & ~n37921;
  assign n37923 = ~pi224 & po1038;
  assign po381 = ~n37922 & ~n37923;
  assign n37925 = ~n6151 & ~n6248;
  assign n37926 = ~pi137 & ~n37925;
  assign n37927 = n6252 & ~n37926;
  assign n37928 = n2920 & ~n11392;
  assign n37929 = ~n2713 & n37928;
  assign n37930 = n2556 & ~n37929;
  assign n37931 = n2554 & ~n37930;
  assign n37932 = ~n2742 & ~n37931;
  assign n37933 = ~pi95 & ~n37932;
  assign n37934 = ~n2727 & ~n37933;
  assign n37935 = pi137 & ~n37934;
  assign n37936 = n2450 & n11392;
  assign n37937 = n2785 & ~n37936;
  assign n37938 = n2795 & ~n37937;
  assign n37939 = pi1093 & ~n37938;
  assign n37940 = n2795 & n7513;
  assign n37941 = n2450 & ~n7468;
  assign n37942 = ~n2531 & n37941;
  assign n37943 = ~pi32 & ~n37942;
  assign n37944 = n37940 & ~n37943;
  assign n37945 = ~pi1093 & ~n37944;
  assign n37946 = ~n7513 & n37938;
  assign n37947 = n11391 & n37941;
  assign n37948 = n37940 & n37947;
  assign n37949 = ~n37946 & ~n37948;
  assign n37950 = n37945 & n37949;
  assign n37951 = ~n37939 & ~n37950;
  assign n37952 = n11523 & ~n37951;
  assign n37953 = n2824 & ~n7513;
  assign n37954 = n37945 & ~n37953;
  assign n37955 = ~n2768 & n37941;
  assign n37956 = ~pi32 & ~n37955;
  assign n37957 = n37940 & ~n37956;
  assign n37958 = pi1093 & ~n37953;
  assign n37959 = ~n37957 & n37958;
  assign n37960 = ~n37954 & ~n37959;
  assign n37961 = n11490 & ~n37960;
  assign n37962 = n37949 & n37961;
  assign n37963 = ~n37952 & ~n37962;
  assign n37964 = ~n37935 & n37963;
  assign n37965 = pi332 & ~n37964;
  assign n37966 = ~n2727 & ~n2744;
  assign n37967 = pi137 & ~n37966;
  assign n37968 = pi1093 & ~n2824;
  assign n37969 = ~n37954 & ~n37968;
  assign n37970 = n11523 & ~n37969;
  assign n37971 = ~n37961 & ~n37970;
  assign n37972 = ~n37967 & n37971;
  assign n37973 = ~pi332 & ~n37972;
  assign n37974 = ~n37965 & ~n37973;
  assign n37975 = ~n2857 & n37974;
  assign n37976 = ~pi137 & ~n37938;
  assign n37977 = ~n37935 & ~n37976;
  assign n37978 = pi332 & ~n37977;
  assign n37979 = ~n2825 & ~n37967;
  assign n37980 = ~pi332 & ~n37979;
  assign n37981 = ~n37978 & ~n37980;
  assign n37982 = n2857 & n37981;
  assign n37983 = ~pi210 & ~n37975;
  assign n37984 = ~n37982 & n37983;
  assign n37985 = ~n2724 & ~n2727;
  assign n37986 = pi137 & ~n37985;
  assign n37987 = ~n2787 & ~n37986;
  assign n37988 = ~pi332 & ~n37987;
  assign n37989 = ~n2501 & ~n37931;
  assign n37990 = ~pi95 & ~n37989;
  assign n37991 = n2889 & ~n37990;
  assign n37992 = ~pi137 & n2502;
  assign n37993 = ~n37937 & n37992;
  assign n37994 = pi332 & ~n37993;
  assign n37995 = ~n37991 & n37994;
  assign n37996 = ~n37988 & ~n37995;
  assign n37997 = pi210 & ~n37996;
  assign n37998 = pi299 & ~n37997;
  assign n37999 = ~n37984 & n37998;
  assign n38000 = n6491 & n37981;
  assign n38001 = ~n6491 & n37974;
  assign n38002 = ~pi198 & ~n38000;
  assign n38003 = ~n38001 & n38002;
  assign n38004 = pi198 & ~n37996;
  assign n38005 = ~pi299 & ~n38004;
  assign n38006 = ~n38003 & n38005;
  assign n38007 = ~n37999 & ~n38006;
  assign n38008 = ~pi39 & ~n38007;
  assign n38009 = pi39 & n3111;
  assign n38010 = ~pi38 & ~n38009;
  assign n38011 = ~n38008 & n38010;
  assign n38012 = pi38 & ~pi137;
  assign n38013 = n6119 & ~n38012;
  assign n38014 = ~n38011 & n38013;
  assign n38015 = ~n37927 & ~n38014;
  assign n38016 = ~pi87 & ~n38015;
  assign n38017 = n3111 & n3208;
  assign n38018 = pi87 & n38017;
  assign n38019 = ~pi75 & ~n38018;
  assign n38020 = ~n38016 & n38019;
  assign n38021 = n7291 & ~n37926;
  assign n38022 = pi75 & ~n38021;
  assign n38023 = ~pi92 & ~n38022;
  assign n38024 = ~n38020 & n38023;
  assign n38025 = pi92 & n3231;
  assign n38026 = n38017 & n38025;
  assign n38027 = ~pi54 & ~n38026;
  assign n38028 = ~n38024 & n38027;
  assign n38029 = n3278 & n38017;
  assign n38030 = pi54 & ~n38029;
  assign n38031 = ~pi74 & ~n38030;
  assign n38032 = ~n38028 & n38031;
  assign n38033 = pi74 & n6113;
  assign n38034 = n38017 & n38033;
  assign n38035 = ~pi55 & ~n38034;
  assign n38036 = ~n38032 & n38035;
  assign n38037 = n7338 & ~n38036;
  assign n38038 = pi56 & n3280;
  assign n38039 = n38017 & n38038;
  assign n38040 = ~n38037 & ~n38039;
  assign n38041 = ~pi62 & ~n38040;
  assign n38042 = n3433 & n38017;
  assign n38043 = pi62 & n38042;
  assign n38044 = n3432 & ~n38043;
  assign n38045 = ~n38041 & n38044;
  assign n38046 = ~pi62 & n38042;
  assign n38047 = ~n3432 & ~n38046;
  assign n38048 = ~n6105 & ~n38047;
  assign po382 = ~n38045 & n38048;
  assign n38050 = pi228 & pi231;
  assign n38051 = ~n2525 & ~n2915;
  assign n38052 = ~pi70 & ~n38051;
  assign n38053 = ~pi51 & ~n38052;
  assign n38054 = n2559 & ~n38053;
  assign n38055 = n2920 & ~n38054;
  assign n38056 = n2556 & ~n38055;
  assign n38057 = n2554 & ~n38056;
  assign n38058 = ~n6158 & ~n38057;
  assign n38059 = ~pi95 & ~n38058;
  assign n38060 = n2788 & ~n38059;
  assign n38061 = ~pi39 & ~n38060;
  assign n38062 = ~pi38 & ~n3353;
  assign n38063 = ~n38061 & n38062;
  assign n38064 = ~pi228 & n38063;
  assign n38065 = ~n38050 & ~n38064;
  assign n38066 = ~pi100 & ~n38065;
  assign n38067 = ~n13967 & ~n38050;
  assign n38068 = pi100 & ~n38067;
  assign n38069 = ~pi87 & ~n38068;
  assign n38070 = ~n38066 & n38069;
  assign n38071 = pi87 & ~n38050;
  assign n38072 = ~n7346 & n38071;
  assign n38073 = ~pi75 & ~n38072;
  assign n38074 = ~n38070 & n38073;
  assign n38075 = ~n13975 & ~n38050;
  assign n38076 = pi75 & ~n38075;
  assign n38077 = ~pi92 & ~n38076;
  assign n38078 = ~n38074 & n38077;
  assign n38079 = pi92 & ~n38050;
  assign n38080 = ~n7372 & n38079;
  assign n38081 = ~n38078 & ~n38080;
  assign n38082 = ~pi54 & ~n38081;
  assign n38083 = pi54 & ~n38050;
  assign n38084 = ~pi74 & ~n38083;
  assign n38085 = ~n38082 & n38084;
  assign n38086 = ~n7381 & ~n38050;
  assign n38087 = pi74 & ~n38086;
  assign n38088 = ~pi55 & ~n38087;
  assign n38089 = ~n38085 & n38088;
  assign n38090 = pi55 & ~n38050;
  assign n38091 = ~pi56 & ~n38090;
  assign n38092 = ~n38089 & n38091;
  assign n38093 = ~n7387 & ~n38050;
  assign n38094 = pi56 & ~n38093;
  assign n38095 = ~pi62 & ~n38094;
  assign n38096 = ~n38092 & n38095;
  assign n38097 = pi62 & ~n38050;
  assign n38098 = ~n7347 & n38097;
  assign n38099 = ~n38096 & ~n38098;
  assign n38100 = n3432 & ~n38099;
  assign n38101 = ~n3432 & ~n38050;
  assign po383 = ~n38100 & ~n38101;
  assign n38103 = n2497 & n6348;
  assign n38104 = ~n6265 & n10999;
  assign n38105 = n2532 & n11009;
  assign n38106 = n11007 & n38105;
  assign n38107 = ~pi91 & ~n2570;
  assign n38108 = ~n38104 & n38107;
  assign n38109 = ~n38106 & n38108;
  assign n38110 = n38103 & ~n38109;
  assign n38111 = ~pi72 & ~n38110;
  assign n38112 = n6372 & ~n38111;
  assign n38113 = pi829 & ~n6181;
  assign n38114 = ~n38112 & n38113;
  assign n38115 = n13055 & ~n13080;
  assign n38116 = n6372 & n38115;
  assign n38117 = ~n6458 & ~n38116;
  assign n38118 = pi1093 & ~n38117;
  assign n38119 = n38103 & ~n38107;
  assign n38120 = ~pi72 & ~n38119;
  assign n38121 = n10999 & n38103;
  assign n38122 = ~n7496 & n38121;
  assign n38123 = ~n8889 & n38120;
  assign n38124 = ~n38122 & n38123;
  assign n38125 = n6372 & ~n38124;
  assign n38126 = ~n38118 & ~n38125;
  assign n38127 = n38120 & ~n38121;
  assign n38128 = n6372 & ~n38127;
  assign n38129 = n10054 & ~n38128;
  assign n38130 = ~n38126 & ~n38129;
  assign n38131 = ~n38114 & n38130;
  assign n38132 = ~pi39 & ~n38131;
  assign po384 = ~n11446 | n38132;
  assign n38134 = ~pi39 & pi228;
  assign n38135 = ~n11395 & ~n11400;
  assign n38136 = pi39 & ~n38135;
  assign n38137 = n6454 & n38136;
  assign n38138 = ~n8890 & ~n10053;
  assign n38139 = ~pi32 & n10216;
  assign n38140 = ~n38138 & n38139;
  assign n38141 = n2541 & n38140;
  assign n38142 = ~n11462 & n38141;
  assign n38143 = ~n38137 & ~n38142;
  assign n38144 = n10181 & ~n38143;
  assign po385 = n38134 | n38144;
  assign n38146 = ~n6118 & n10178;
  assign n38147 = ~n6179 & n7495;
  assign n38148 = n16732 & n38147;
  assign n38149 = n16657 & ~n38147;
  assign n38150 = pi1091 & ~n38148;
  assign n38151 = ~n38149 & n38150;
  assign n38152 = n6446 & n16732;
  assign n38153 = ~n6446 & n16657;
  assign n38154 = ~pi1091 & ~n38152;
  assign n38155 = ~n38153 & n38154;
  assign n38156 = ~n38151 & ~n38155;
  assign n38157 = ~pi120 & ~n38156;
  assign n38158 = ~n16659 & ~n38157;
  assign n38159 = ~n6200 & n38158;
  assign n38160 = ~n35590 & ~n38159;
  assign n38161 = ~n6197 & n38160;
  assign n38162 = ~n6206 & n16660;
  assign n38163 = n6206 & n38158;
  assign n38164 = ~n38162 & ~n38163;
  assign n38165 = n6197 & n38164;
  assign n38166 = ~n3053 & ~n38161;
  assign n38167 = ~n38165 & n38166;
  assign n38168 = n3053 & n16660;
  assign n38169 = ~pi223 & ~n38168;
  assign n38170 = ~n38167 & n38169;
  assign n38171 = pi120 & n6184;
  assign n38172 = n16660 & ~n38171;
  assign n38173 = ~n35590 & ~n38172;
  assign n38174 = ~n6197 & ~n38173;
  assign n38175 = ~n38162 & ~n38172;
  assign n38176 = n6197 & ~n38175;
  assign n38177 = pi223 & ~n38174;
  assign n38178 = ~n38176 & n38177;
  assign n38179 = ~pi299 & ~n38178;
  assign n38180 = ~n38170 & n38179;
  assign n38181 = ~n6223 & n38160;
  assign n38182 = n6223 & n38164;
  assign n38183 = ~n3461 & ~n38181;
  assign n38184 = ~n38182 & n38183;
  assign n38185 = ~pi215 & ~n16934;
  assign n38186 = ~n38184 & n38185;
  assign n38187 = ~n6223 & ~n38173;
  assign n38188 = n6223 & ~n38175;
  assign n38189 = pi215 & ~n38187;
  assign n38190 = ~n38188 & n38189;
  assign n38191 = pi299 & ~n38190;
  assign n38192 = ~n38186 & n38191;
  assign n38193 = ~n38180 & ~n38192;
  assign n38194 = pi39 & ~n38193;
  assign n38195 = pi829 & pi1091;
  assign n38196 = n16640 & n38195;
  assign n38197 = ~pi824 & ~n38196;
  assign n38198 = pi824 & ~n16635;
  assign n38199 = ~n6450 & ~n38197;
  assign n38200 = ~n38198 & n38199;
  assign n38201 = ~n16601 & ~n38200;
  assign n38202 = n38195 & n38197;
  assign n38203 = ~n38198 & ~n38202;
  assign n38204 = n6265 & ~n6450;
  assign n38205 = ~n38203 & n38204;
  assign n38206 = ~n6151 & ~n6450;
  assign n38207 = ~n38201 & ~n38206;
  assign n38208 = ~n38205 & n38207;
  assign n38209 = ~n7496 & n16601;
  assign n38210 = ~n16618 & ~n38209;
  assign n38211 = n38206 & ~n38210;
  assign n38212 = pi1093 & ~n38211;
  assign n38213 = ~n38208 & n38212;
  assign n38214 = ~n6266 & n16601;
  assign n38215 = n6152 & n16589;
  assign n38216 = ~n16591 & n38215;
  assign n38217 = ~pi40 & ~n38216;
  assign n38218 = n10262 & ~n38217;
  assign n38219 = pi252 & ~n38218;
  assign n38220 = n6266 & ~n16588;
  assign n38221 = ~n38219 & n38220;
  assign n38222 = ~pi1093 & ~n38221;
  assign n38223 = ~n38214 & n38222;
  assign n38224 = ~pi39 & ~n38223;
  assign n38225 = ~n38213 & n38224;
  assign n38226 = ~pi38 & ~n38194;
  assign n38227 = ~n38225 & n38226;
  assign po387 = n38146 & ~n38227;
  assign n38229 = ~pi81 & ~n2675;
  assign n38230 = n6333 & ~n38229;
  assign n38231 = n2451 & ~n38230;
  assign n38232 = n2683 & ~n38231;
  assign n38233 = n2594 & ~n38232;
  assign n38234 = n2687 & ~n38233;
  assign n38235 = n2504 & ~n38234;
  assign n38236 = ~n2507 & ~n38235;
  assign n38237 = ~pi86 & ~n38236;
  assign n38238 = n2592 & ~n38237;
  assign n38239 = n2590 & ~n38238;
  assign n38240 = ~n2585 & ~n38239;
  assign n38241 = ~pi108 & ~n38240;
  assign n38242 = n2584 & ~n38241;
  assign n38243 = n2699 & ~n38242;
  assign n38244 = ~n2575 & ~n38243;
  assign n38245 = n2574 & ~n38244;
  assign n38246 = n2573 & ~n38245;
  assign n38247 = n2566 & ~n38246;
  assign n38248 = n2900 & ~n38247;
  assign n38249 = n2547 & ~n38248;
  assign n38250 = n15573 & ~n38249;
  assign n38251 = ~pi70 & ~n38250;
  assign n38252 = ~n2917 & ~n38251;
  assign n38253 = ~pi51 & ~n38252;
  assign n38254 = n2559 & ~n38253;
  assign n38255 = n2920 & ~n38254;
  assign n38256 = n2556 & ~n38255;
  assign n38257 = ~pi1082 & n2553;
  assign n38258 = ~pi32 & ~n38257;
  assign n38259 = ~n38256 & n38258;
  assign n38260 = ~n3363 & ~n38259;
  assign n38261 = ~pi95 & ~n38260;
  assign n38262 = ~n2727 & ~n38261;
  assign n38263 = ~pi39 & ~n38262;
  assign n38264 = ~n7297 & ~n7299;
  assign po950 = ~n6183 | ~n6265;
  assign n38266 = n6444 & ~po950;
  assign n38267 = ~n38264 & n38266;
  assign n38268 = n6175 & n11344;
  assign n38269 = ~n38267 & n38268;
  assign n38270 = ~n3353 & ~n38269;
  assign n38271 = ~n38263 & n38270;
  assign n38272 = ~pi38 & ~n38271;
  assign n38273 = n6119 & ~n38272;
  assign n38274 = ~pi87 & ~n6252;
  assign n38275 = ~n38273 & n38274;
  assign n38276 = ~n6277 & ~n38275;
  assign n38277 = n3238 & ~n38276;
  assign n38278 = n7296 & ~n38277;
  assign n38279 = ~pi54 & ~n38278;
  assign n38280 = ~n7331 & ~n38279;
  assign n38281 = n8865 & ~n38280;
  assign n38282 = n15663 & ~n38281;
  assign n38283 = ~pi56 & ~n38282;
  assign n38284 = ~n6112 & ~n38283;
  assign n38285 = ~pi62 & ~n38284;
  assign n38286 = ~n6288 & ~n38285;
  assign n38287 = n3432 & ~n38286;
  assign po389 = n6108 & ~n38287;
  assign n38289 = ~pi230 & ~pi233;
  assign n38290 = ~pi212 & ~pi214;
  assign n38291 = ~pi211 & ~n38290;
  assign n38292 = pi219 & ~n38291;
  assign n38293 = po1038 & ~n38292;
  assign n38294 = pi1142 & ~n10656;
  assign n38295 = pi211 & pi1143;
  assign n38296 = ~pi211 & pi1144;
  assign n38297 = ~n38295 & ~n38296;
  assign n38298 = ~pi212 & pi214;
  assign n38299 = pi212 & ~pi214;
  assign n38300 = ~n38298 & ~n38299;
  assign n38301 = ~n38297 & ~n38300;
  assign n38302 = ~pi211 & pi1143;
  assign n38303 = n10708 & n38302;
  assign n38304 = ~n38301 & ~n38303;
  assign n38305 = ~pi219 & ~n38304;
  assign n38306 = ~n38294 & ~n38305;
  assign n38307 = n38293 & ~n38306;
  assign n38308 = pi299 & ~n38297;
  assign n38309 = pi199 & pi1142;
  assign n38310 = ~pi200 & ~n38309;
  assign n38311 = ~pi199 & pi1144;
  assign n38312 = n38310 & ~n38311;
  assign n38313 = ~pi199 & pi1143;
  assign n38314 = pi200 & ~n38313;
  assign n38315 = ~n38312 & ~n38314;
  assign n38316 = ~pi299 & ~n38315;
  assign n38317 = ~pi207 & ~n38316;
  assign n38318 = n38310 & ~n38313;
  assign n38319 = pi207 & ~pi299;
  assign n38320 = ~pi199 & pi1142;
  assign n38321 = pi200 & ~n38320;
  assign n38322 = n38319 & ~n38321;
  assign n38323 = ~n38318 & n38322;
  assign n38324 = ~n38317 & ~n38323;
  assign n38325 = pi208 & ~n38324;
  assign n38326 = pi207 & ~pi208;
  assign n38327 = n38315 & n38326;
  assign n38328 = ~n38325 & ~n38327;
  assign n38329 = ~pi299 & ~n38328;
  assign n38330 = ~pi214 & ~n38329;
  assign n38331 = ~n38308 & n38330;
  assign n38332 = pi211 & pi1142;
  assign n38333 = ~n38302 & ~n38332;
  assign n38334 = pi299 & ~n38333;
  assign n38335 = pi214 & ~n38334;
  assign n38336 = ~n38329 & n38335;
  assign n38337 = pi212 & ~n38336;
  assign n38338 = ~n38331 & n38337;
  assign n38339 = ~n38308 & ~n38329;
  assign n38340 = ~pi212 & ~n38330;
  assign n38341 = ~n38339 & n38340;
  assign n38342 = ~pi219 & ~n38338;
  assign n38343 = ~n38341 & n38342;
  assign n38344 = ~n38291 & n38329;
  assign n38345 = ~pi299 & n38328;
  assign n38346 = pi299 & ~pi1142;
  assign n38347 = n38291 & ~n38346;
  assign n38348 = ~n38345 & n38347;
  assign n38349 = pi219 & ~n38344;
  assign n38350 = ~n38348 & n38349;
  assign n38351 = ~po1038 & ~n38350;
  assign n38352 = ~n38343 & n38351;
  assign n38353 = ~n38307 & ~n38352;
  assign n38354 = pi213 & n38353;
  assign n38355 = ~pi211 & pi1156;
  assign n38356 = pi211 & pi1155;
  assign n38357 = ~n38355 & ~n38356;
  assign n38358 = ~pi214 & ~n38357;
  assign n38359 = ~pi211 & pi1155;
  assign n38360 = pi211 & pi1154;
  assign n38361 = ~n38359 & ~n38360;
  assign n38362 = pi214 & ~n38361;
  assign n38363 = ~n38358 & ~n38362;
  assign n38364 = pi212 & ~n38363;
  assign n38365 = ~pi211 & pi1157;
  assign n38366 = pi211 & pi1156;
  assign n38367 = ~n38365 & ~n38366;
  assign n38368 = n38298 & ~n38367;
  assign n38369 = ~n38364 & ~n38368;
  assign n38370 = ~pi219 & n38369;
  assign n38371 = ~pi211 & pi214;
  assign n38372 = pi1155 & n38371;
  assign n38373 = ~pi212 & ~n38372;
  assign n38374 = ~pi211 & pi1154;
  assign n38375 = ~pi214 & ~n38374;
  assign n38376 = ~pi211 & pi1153;
  assign n38377 = n10708 & ~n38376;
  assign n38378 = ~n38375 & ~n38377;
  assign n38379 = ~n38373 & n38378;
  assign n38380 = pi219 & ~n38379;
  assign n38381 = po1038 & ~n38380;
  assign n38382 = ~n38370 & n38381;
  assign n38383 = ~pi213 & ~n38382;
  assign n38384 = ~pi219 & pi299;
  assign n38385 = ~n38369 & n38384;
  assign n38386 = pi299 & pi1155;
  assign n38387 = n38298 & n38386;
  assign n38388 = pi299 & pi1153;
  assign n38389 = pi214 & ~n38388;
  assign n38390 = pi299 & pi1154;
  assign n38391 = ~pi214 & ~n38390;
  assign n38392 = pi212 & ~n38389;
  assign n38393 = ~n38391 & n38392;
  assign n38394 = ~n38387 & ~n38393;
  assign n38395 = ~pi211 & pi219;
  assign n38396 = ~n38394 & n38395;
  assign n38397 = ~n38385 & ~n38396;
  assign n38398 = ~n38329 & n38397;
  assign n38399 = ~po1038 & ~n38398;
  assign n38400 = n38383 & ~n38399;
  assign n38401 = pi209 & ~n38400;
  assign n38402 = ~n38354 & n38401;
  assign n38403 = ~pi200 & pi1155;
  assign n38404 = pi199 & n38403;
  assign n38405 = ~pi299 & n38404;
  assign n38406 = ~pi1156 & ~n38405;
  assign n38407 = ~pi200 & ~pi1155;
  assign n38408 = pi199 & pi200;
  assign n38409 = ~n10793 & ~n38408;
  assign n38410 = ~pi299 & n38409;
  assign n38411 = ~n38407 & n38410;
  assign n38412 = ~n38406 & n38411;
  assign n38413 = pi207 & n38412;
  assign n38414 = ~pi208 & ~n38413;
  assign n38415 = ~pi299 & ~n38408;
  assign n38416 = pi1153 & ~n38415;
  assign n38417 = pi1154 & ~n38416;
  assign n38418 = n11348 & n38403;
  assign n38419 = ~pi1153 & ~n11348;
  assign n38420 = pi1154 & n38409;
  assign n38421 = ~n38419 & n38420;
  assign n38422 = ~n38418 & ~n38421;
  assign n38423 = n38417 & ~n38422;
  assign n38424 = ~pi200 & ~pi299;
  assign n38425 = pi199 & ~pi1153;
  assign n38426 = n38424 & ~n38425;
  assign n38427 = ~pi199 & ~pi1155;
  assign n38428 = ~pi1154 & ~n38427;
  assign n38429 = n38426 & n38428;
  assign n38430 = ~n38423 & ~n38429;
  assign n38431 = pi207 & n38430;
  assign n38432 = pi200 & ~pi299;
  assign n38433 = ~pi199 & pi1155;
  assign n38434 = n38432 & n38433;
  assign n38435 = ~pi1154 & ~n38434;
  assign n38436 = pi200 & ~n38433;
  assign n38437 = n10794 & ~n38436;
  assign n38438 = ~n38435 & n38437;
  assign n38439 = pi200 & ~pi1155;
  assign n38440 = n11348 & ~n38439;
  assign n38441 = pi1156 & n38440;
  assign n38442 = ~n38438 & ~n38441;
  assign n38443 = ~pi207 & n38442;
  assign n38444 = ~n38431 & ~n38443;
  assign n38445 = pi208 & ~n38444;
  assign n38446 = ~n38414 & ~n38445;
  assign n38447 = ~pi1157 & ~n38446;
  assign n38448 = pi199 & ~pi1155;
  assign n38449 = pi1156 & ~n38448;
  assign n38450 = n38415 & n38449;
  assign n38451 = ~pi1156 & n38424;
  assign n38452 = ~n38448 & n38451;
  assign n38453 = ~n38450 & ~n38452;
  assign n38454 = pi207 & ~n38453;
  assign n38455 = ~pi208 & ~n38454;
  assign n38456 = ~n38445 & ~n38455;
  assign n38457 = pi1157 & ~n38456;
  assign n38458 = ~n38447 & ~n38457;
  assign n38459 = pi211 & ~n38458;
  assign n38460 = ~pi214 & ~n38458;
  assign n38461 = ~pi212 & ~n38460;
  assign n38462 = n11358 & n38407;
  assign n38463 = pi1153 & n38462;
  assign n38464 = pi1153 & ~n38432;
  assign n38465 = ~pi1153 & ~n10794;
  assign n38466 = ~n38464 & ~n38465;
  assign n38467 = pi1155 & ~n38466;
  assign n38468 = ~n38463 & ~n38467;
  assign n38469 = ~pi1154 & ~n38468;
  assign n38470 = pi1155 & ~n11358;
  assign n38471 = n38410 & ~n38425;
  assign n38472 = ~n38470 & ~n38471;
  assign n38473 = pi1154 & ~n38472;
  assign n38474 = ~n38469 & ~n38473;
  assign n38475 = pi207 & n38474;
  assign n38476 = ~pi207 & ~n38386;
  assign n38477 = n38442 & n38476;
  assign n38478 = pi208 & ~n38477;
  assign n38479 = ~n38475 & n38478;
  assign n38480 = pi1155 & ~n38432;
  assign n38481 = ~n11348 & ~n38480;
  assign n38482 = pi1156 & ~n38481;
  assign n38483 = pi199 & ~pi200;
  assign n38484 = ~pi299 & ~n38483;
  assign n38485 = ~pi1155 & ~n38484;
  assign n38486 = ~pi1156 & ~n38432;
  assign n38487 = ~n38485 & n38486;
  assign n38488 = ~n38482 & ~n38487;
  assign n38489 = pi207 & n38488;
  assign n38490 = ~pi208 & ~n38476;
  assign n38491 = pi1157 & n38490;
  assign n38492 = ~n38489 & n38491;
  assign n38493 = ~pi299 & n38406;
  assign n38494 = ~pi299 & ~n38409;
  assign n38495 = ~pi1155 & ~n11348;
  assign n38496 = ~n38494 & ~n38495;
  assign n38497 = ~n38493 & n38496;
  assign n38498 = n38490 & n38497;
  assign n38499 = ~n38492 & ~n38498;
  assign n38500 = ~n38479 & n38499;
  assign n38501 = n38371 & n38500;
  assign n38502 = n38461 & ~n38501;
  assign n38503 = ~pi211 & ~pi214;
  assign n38504 = pi1155 & ~n38494;
  assign n38505 = ~n38485 & ~n38504;
  assign n38506 = pi1154 & ~n38505;
  assign n38507 = n38442 & ~n38506;
  assign n38508 = ~pi207 & ~n38507;
  assign n38509 = ~pi299 & n38472;
  assign n38510 = pi1154 & ~n38509;
  assign n38511 = ~n38429 & ~n38510;
  assign n38512 = pi207 & ~n38511;
  assign n38513 = ~n38508 & ~n38512;
  assign n38514 = pi208 & ~n38513;
  assign n38515 = ~pi1155 & ~n10794;
  assign n38516 = ~n38480 & ~n38515;
  assign n38517 = n11358 & ~n38403;
  assign n38518 = pi1156 & ~n38517;
  assign n38519 = n38516 & ~n38518;
  assign n38520 = pi207 & n38519;
  assign n38521 = ~pi207 & ~pi299;
  assign n38522 = ~pi208 & ~n38521;
  assign n38523 = ~n38520 & n38522;
  assign n38524 = pi299 & ~pi1154;
  assign n38525 = pi1157 & ~n38524;
  assign n38526 = n38523 & n38525;
  assign n38527 = ~n38390 & ~n38413;
  assign n38528 = ~pi208 & ~n38527;
  assign n38529 = ~pi1157 & n38528;
  assign n38530 = ~n38526 & ~n38529;
  assign n38531 = ~n38514 & n38530;
  assign n38532 = n38503 & n38531;
  assign n38533 = pi1153 & ~n38484;
  assign n38534 = n38422 & ~n38533;
  assign n38535 = pi207 & ~n38534;
  assign n38536 = ~n38470 & ~n38515;
  assign n38537 = pi1156 & ~n38536;
  assign n38538 = ~n38506 & ~n38537;
  assign n38539 = pi299 & ~pi1155;
  assign n38540 = ~pi299 & ~n11419;
  assign n38541 = pi1155 & ~n38540;
  assign n38542 = ~n38539 & ~n38541;
  assign n38543 = n38538 & n38542;
  assign n38544 = pi299 & ~pi1153;
  assign n38545 = ~pi207 & ~n38544;
  assign n38546 = ~n38543 & n38545;
  assign n38547 = ~n38535 & ~n38546;
  assign n38548 = pi208 & ~n38547;
  assign n38549 = pi1156 & ~n38404;
  assign n38550 = n38540 & n38549;
  assign n38551 = ~n38406 & ~n38550;
  assign n38552 = pi207 & n38551;
  assign n38553 = ~pi299 & ~n38552;
  assign n38554 = ~pi208 & ~n38553;
  assign n38555 = ~pi1157 & ~n38554;
  assign n38556 = pi1157 & ~n38523;
  assign n38557 = ~n38544 & ~n38556;
  assign n38558 = ~n38555 & n38557;
  assign n38559 = n38371 & ~n38558;
  assign n38560 = ~n38548 & n38559;
  assign n38561 = pi212 & ~n38560;
  assign n38562 = ~n38532 & n38561;
  assign n38563 = ~n38502 & ~n38562;
  assign n38564 = ~n38459 & ~n38563;
  assign n38565 = pi219 & ~n38564;
  assign n38566 = ~pi207 & n38543;
  assign n38567 = n38319 & n38534;
  assign n38568 = pi208 & ~n38567;
  assign n38569 = ~n38566 & n38568;
  assign n38570 = n38556 & ~n38569;
  assign n38571 = ~pi211 & ~n38570;
  assign n38572 = ~n38447 & n38571;
  assign n38573 = pi207 & ~n38430;
  assign n38574 = ~n38438 & ~n38537;
  assign n38575 = ~pi207 & ~n38574;
  assign n38576 = pi299 & pi1156;
  assign n38577 = pi207 & n38576;
  assign n38578 = ~n38575 & ~n38577;
  assign n38579 = ~n38573 & n38578;
  assign n38580 = pi208 & ~n38579;
  assign n38581 = ~n38406 & n38554;
  assign n38582 = ~pi208 & pi1157;
  assign n38583 = ~n38454 & ~n38576;
  assign n38584 = n38582 & ~n38583;
  assign n38585 = ~n38581 & ~n38584;
  assign n38586 = ~n38580 & n38585;
  assign n38587 = pi211 & ~n38586;
  assign n38588 = pi214 & ~n38587;
  assign n38589 = ~n38572 & n38588;
  assign n38590 = n38461 & ~n38589;
  assign n38591 = n10654 & ~n38531;
  assign n38592 = ~n10654 & ~n38503;
  assign n38593 = ~n38500 & n38592;
  assign n38594 = n38503 & ~n38586;
  assign n38595 = ~n38593 & ~n38594;
  assign n38596 = ~n38591 & n38595;
  assign n38597 = pi212 & ~n38596;
  assign n38598 = ~pi219 & ~n38597;
  assign n38599 = ~n38590 & n38598;
  assign n38600 = ~po1038 & ~n38599;
  assign n38601 = ~n38565 & n38600;
  assign n38602 = n38383 & ~n38601;
  assign n38603 = ~pi211 & n10708;
  assign n38604 = pi299 & pi1143;
  assign n38605 = n38431 & ~n38604;
  assign n38606 = pi299 & ~pi1143;
  assign n38607 = n38504 & ~n38606;
  assign n38608 = ~pi1155 & n38604;
  assign n38609 = pi1154 & ~n38462;
  assign n38610 = ~n38608 & n38609;
  assign n38611 = ~n38607 & n38610;
  assign n38612 = n38435 & ~n38604;
  assign n38613 = ~pi1156 & ~n38612;
  assign n38614 = ~n38611 & n38613;
  assign n38615 = ~n38536 & ~n38606;
  assign n38616 = ~pi1154 & ~n38615;
  assign n38617 = ~pi299 & ~n38436;
  assign n38618 = pi1154 & ~n38617;
  assign n38619 = ~n38604 & n38618;
  assign n38620 = pi1156 & ~n38619;
  assign n38621 = ~n38616 & n38620;
  assign n38622 = ~n38614 & ~n38621;
  assign n38623 = ~pi207 & n38622;
  assign n38624 = pi208 & ~n38605;
  assign n38625 = ~n38623 & n38624;
  assign n38626 = ~pi1157 & n38554;
  assign n38627 = ~n38606 & n38626;
  assign n38628 = ~n38450 & n38516;
  assign n38629 = pi207 & ~n38606;
  assign n38630 = ~n38628 & n38629;
  assign n38631 = ~n38604 & ~n38630;
  assign n38632 = n38582 & ~n38631;
  assign n38633 = ~n38627 & ~n38632;
  assign n38634 = ~n38625 & n38633;
  assign n38635 = n38603 & n38634;
  assign n38636 = pi211 & ~n38634;
  assign n38637 = pi299 & pi1144;
  assign n38638 = n38431 & ~n38637;
  assign n38639 = pi299 & ~pi1144;
  assign n38640 = n38504 & ~n38639;
  assign n38641 = ~pi1155 & n38637;
  assign n38642 = n38609 & ~n38641;
  assign n38643 = ~n38640 & n38642;
  assign n38644 = n38435 & ~n38637;
  assign n38645 = ~pi1156 & ~n38644;
  assign n38646 = ~n38643 & n38645;
  assign n38647 = ~n38536 & ~n38639;
  assign n38648 = ~pi1154 & ~n38647;
  assign n38649 = n38618 & ~n38637;
  assign n38650 = pi1156 & ~n38649;
  assign n38651 = ~n38648 & n38650;
  assign n38652 = ~n38646 & ~n38651;
  assign n38653 = ~pi207 & n38652;
  assign n38654 = pi208 & ~n38638;
  assign n38655 = ~n38653 & n38654;
  assign n38656 = n38626 & ~n38639;
  assign n38657 = pi207 & ~n38639;
  assign n38658 = ~n38628 & n38657;
  assign n38659 = ~n38637 & ~n38658;
  assign n38660 = n38582 & ~n38659;
  assign n38661 = ~n38656 & ~n38660;
  assign n38662 = ~n38655 & n38661;
  assign n38663 = ~pi211 & ~n38662;
  assign n38664 = ~n10708 & ~n38290;
  assign n38665 = ~n38636 & n38664;
  assign n38666 = ~n38663 & n38665;
  assign n38667 = ~n38635 & ~n38666;
  assign n38668 = ~pi219 & ~n38667;
  assign n38669 = ~pi219 & ~n38290;
  assign n38670 = ~n38291 & ~n38669;
  assign n38671 = ~n38458 & n38670;
  assign n38672 = ~pi299 & ~n38474;
  assign n38673 = pi299 & pi1142;
  assign n38674 = pi207 & ~n38673;
  assign n38675 = ~n38672 & n38674;
  assign n38676 = ~n38346 & ~n38538;
  assign n38677 = ~n38434 & ~n38673;
  assign n38678 = ~pi1154 & ~pi1156;
  assign n38679 = ~n38677 & n38678;
  assign n38680 = ~pi207 & ~n38679;
  assign n38681 = ~n38676 & n38680;
  assign n38682 = pi208 & ~n38681;
  assign n38683 = ~n38675 & n38682;
  assign n38684 = ~n38346 & ~n38556;
  assign n38685 = ~n38555 & n38684;
  assign n38686 = ~n10656 & ~n38670;
  assign n38687 = ~n38685 & n38686;
  assign n38688 = ~n38683 & n38687;
  assign n38689 = ~po1038 & ~n38688;
  assign n38690 = ~n38671 & n38689;
  assign n38691 = ~n38668 & n38690;
  assign n38692 = pi213 & ~n38307;
  assign n38693 = ~n38691 & n38692;
  assign n38694 = ~pi209 & ~n38693;
  assign n38695 = ~n38602 & n38694;
  assign n38696 = ~n38402 & ~n38695;
  assign n38697 = pi230 & ~n38696;
  assign po390 = n38289 | n38697;
  assign n38699 = pi211 & pi1153;
  assign n38700 = ~n38374 & ~n38699;
  assign n38701 = ~n10708 & n38700;
  assign n38702 = n38669 & ~n38701;
  assign n38703 = ~n38377 & n38702;
  assign n38704 = po1038 & n38703;
  assign n38705 = ~pi1152 & ~n38704;
  assign n38706 = ~n10463 & n38442;
  assign n38707 = ~pi207 & ~pi208;
  assign n38708 = ~n10463 & ~n38707;
  assign n38709 = ~pi1154 & ~n38418;
  assign n38710 = ~pi199 & n38407;
  assign n38711 = pi207 & n38415;
  assign n38712 = ~n38710 & n38711;
  assign n38713 = ~n38709 & n38712;
  assign n38714 = ~n38708 & ~n38713;
  assign n38715 = ~n38706 & ~n38714;
  assign n38716 = ~pi214 & ~n38715;
  assign n38717 = ~pi212 & ~n38716;
  assign n38718 = ~pi207 & n38390;
  assign n38719 = pi207 & ~n38507;
  assign n38720 = ~n38718 & ~n38719;
  assign n38721 = ~pi208 & ~n38720;
  assign n38722 = ~pi1155 & n10793;
  assign n38723 = ~n38408 & ~n38722;
  assign n38724 = ~pi299 & ~n38723;
  assign n38725 = ~n38709 & ~n38724;
  assign n38726 = pi207 & n38725;
  assign n38727 = ~n38508 & ~n38726;
  assign n38728 = pi208 & ~n38727;
  assign n38729 = ~n38721 & ~n38728;
  assign n38730 = ~pi211 & ~n38729;
  assign n38731 = pi207 & n38542;
  assign n38732 = n38538 & n38731;
  assign n38733 = n38522 & ~n38732;
  assign n38734 = n38319 & ~n38725;
  assign n38735 = pi208 & ~n38734;
  assign n38736 = ~n38566 & n38735;
  assign n38737 = ~n38733 & ~n38736;
  assign n38738 = ~n38544 & ~n38737;
  assign n38739 = pi211 & n38738;
  assign n38740 = ~n38730 & ~n38739;
  assign n38741 = pi214 & n38740;
  assign n38742 = n38717 & ~n38741;
  assign n38743 = ~pi219 & ~n38742;
  assign n38744 = ~pi214 & ~n38740;
  assign n38745 = ~pi211 & ~n38738;
  assign n38746 = pi214 & ~n38745;
  assign n38747 = pi211 & ~n38715;
  assign n38748 = n38746 & ~n38747;
  assign n38749 = ~n38744 & ~n38748;
  assign n38750 = pi212 & ~n38749;
  assign n38751 = n38743 & ~n38750;
  assign n38752 = pi219 & ~n38715;
  assign n38753 = ~po1038 & ~n38752;
  assign n38754 = ~n38751 & n38753;
  assign n38755 = n38705 & ~n38754;
  assign n38756 = pi1153 & ~n38503;
  assign n38757 = ~n38371 & ~n38375;
  assign n38758 = ~n38756 & ~n38757;
  assign n38759 = pi212 & ~n38758;
  assign n38760 = n38298 & ~n38700;
  assign n38761 = ~pi219 & ~n38760;
  assign n38762 = ~n38759 & n38761;
  assign n38763 = n38293 & ~n38762;
  assign n38764 = pi1152 & ~n38763;
  assign n38765 = ~n38737 & n38746;
  assign n38766 = ~n38744 & ~n38765;
  assign n38767 = pi212 & ~n38766;
  assign n38768 = n38743 & ~n38767;
  assign n38769 = ~n38291 & n38715;
  assign n38770 = pi219 & ~n38769;
  assign n38771 = n38291 & ~n38737;
  assign n38772 = n38770 & ~n38771;
  assign n38773 = ~po1038 & ~n38772;
  assign n38774 = ~n38768 & n38773;
  assign n38775 = n38764 & ~n38774;
  assign n38776 = ~pi213 & ~n38755;
  assign n38777 = ~n38775 & n38776;
  assign n38778 = pi207 & ~n38574;
  assign n38779 = ~n38576 & ~n38778;
  assign n38780 = ~pi208 & ~n38779;
  assign n38781 = n38578 & ~n38713;
  assign n38782 = pi208 & ~n38781;
  assign n38783 = ~n38780 & ~n38782;
  assign n38784 = ~pi211 & ~n38783;
  assign n38785 = ~n38386 & ~n38715;
  assign n38786 = pi211 & ~n38785;
  assign n38787 = ~n38784 & ~n38786;
  assign n38788 = pi214 & n38787;
  assign n38789 = n38717 & ~n38788;
  assign n38790 = ~pi214 & n38787;
  assign n38791 = pi211 & ~n38729;
  assign n38792 = ~pi211 & ~n38785;
  assign n38793 = pi214 & ~n38792;
  assign n38794 = ~n38791 & n38793;
  assign n38795 = pi212 & ~n38794;
  assign n38796 = ~n38790 & n38795;
  assign n38797 = ~pi219 & ~n38789;
  assign n38798 = ~n38796 & n38797;
  assign n38799 = ~n38290 & n38730;
  assign n38800 = n38770 & ~n38799;
  assign n38801 = n35703 & ~n38800;
  assign n38802 = ~n38798 & n38801;
  assign n38803 = pi209 & ~n38802;
  assign n38804 = ~n38777 & n38803;
  assign n38805 = ~pi199 & pi1153;
  assign n38806 = pi200 & n38805;
  assign n38807 = ~pi299 & n38806;
  assign n38808 = ~pi1154 & ~n38807;
  assign n38809 = pi1154 & n38432;
  assign n38810 = ~n38805 & n38809;
  assign n38811 = ~n38808 & ~n38810;
  assign n38812 = n38484 & ~n38811;
  assign n38813 = n38522 & ~n38812;
  assign n38814 = ~pi207 & n38812;
  assign n38815 = ~pi200 & ~pi1153;
  assign n38816 = ~pi199 & ~n38815;
  assign n38817 = ~pi299 & ~n38816;
  assign n38818 = ~n38483 & n38817;
  assign n38819 = pi207 & n38818;
  assign n38820 = pi208 & ~n38819;
  assign n38821 = ~n38814 & n38820;
  assign n38822 = ~n38813 & ~n38821;
  assign n38823 = ~pi211 & n38822;
  assign n38824 = ~pi299 & n10793;
  assign n38825 = ~pi1153 & ~n38824;
  assign n38826 = n38417 & ~n38825;
  assign n38827 = ~pi199 & ~pi1153;
  assign n38828 = n38410 & ~n38827;
  assign n38829 = ~n38826 & ~n38828;
  assign n38830 = ~n10463 & n38829;
  assign n38831 = ~pi1153 & n10793;
  assign n38832 = n38415 & ~n38831;
  assign n38833 = n10463 & ~n38832;
  assign n38834 = ~n38707 & ~n38833;
  assign n38835 = ~n38830 & n38834;
  assign n38836 = pi211 & ~n38835;
  assign n38837 = ~n38823 & ~n38836;
  assign n38838 = ~n38290 & n38837;
  assign n38839 = pi219 & ~n38290;
  assign n38840 = pi219 & ~n38835;
  assign n38841 = ~n38839 & ~n38840;
  assign n38842 = ~n38838 & ~n38841;
  assign n38843 = ~po1038 & ~n38842;
  assign n38844 = pi207 & ~n38829;
  assign n38845 = ~n38390 & ~n38844;
  assign n38846 = ~pi208 & ~n38845;
  assign n38847 = pi207 & ~n38818;
  assign n38848 = ~n38524 & n38847;
  assign n38849 = pi1154 & ~n10794;
  assign n38850 = ~n38826 & ~n38849;
  assign n38851 = ~n38828 & n38850;
  assign n38852 = ~pi207 & ~n38851;
  assign n38853 = ~n38848 & ~n38852;
  assign n38854 = pi208 & ~n38853;
  assign n38855 = ~n38846 & ~n38854;
  assign n38856 = ~pi211 & ~n38855;
  assign n38857 = ~pi207 & n38388;
  assign n38858 = ~pi1153 & ~n38424;
  assign n38859 = ~n38494 & ~n38858;
  assign n38860 = pi1154 & ~n11358;
  assign n38861 = ~n38858 & n38860;
  assign n38862 = ~n38859 & ~n38861;
  assign n38863 = pi207 & ~n38862;
  assign n38864 = ~n38857 & ~n38863;
  assign n38865 = ~pi208 & ~n38864;
  assign n38866 = ~pi207 & ~n38862;
  assign n38867 = ~pi299 & n38408;
  assign n38868 = pi207 & ~n38867;
  assign n38869 = ~n38465 & n38868;
  assign n38870 = ~n38866 & ~n38869;
  assign n38871 = pi208 & ~n38870;
  assign n38872 = ~n38865 & ~n38871;
  assign n38873 = pi211 & ~n38872;
  assign n38874 = ~n38856 & ~n38873;
  assign n38875 = ~pi214 & n38874;
  assign n38876 = ~pi211 & ~n38872;
  assign n38877 = pi211 & ~n38822;
  assign n38878 = pi214 & ~n38876;
  assign n38879 = ~n38877 & n38878;
  assign n38880 = pi212 & ~n38879;
  assign n38881 = ~n38875 & n38880;
  assign n38882 = ~pi214 & ~n38835;
  assign n38883 = ~pi212 & ~n38882;
  assign n38884 = pi214 & n38874;
  assign n38885 = n38883 & ~n38884;
  assign n38886 = ~pi219 & ~n38881;
  assign n38887 = ~n38885 & n38886;
  assign n38888 = n38843 & ~n38887;
  assign n38889 = n38764 & ~n38888;
  assign n38890 = pi1153 & ~pi1154;
  assign n38891 = ~n38540 & n38890;
  assign n38892 = ~n38861 & ~n38891;
  assign n38893 = pi207 & ~n38892;
  assign n38894 = ~n38857 & ~n38893;
  assign n38895 = ~pi208 & ~n38894;
  assign n38896 = ~pi207 & ~n38892;
  assign n38897 = pi207 & ~n10794;
  assign n38898 = pi1153 & n38897;
  assign n38899 = ~n38896 & ~n38898;
  assign n38900 = pi208 & ~n38899;
  assign n38901 = ~n38895 & ~n38900;
  assign n38902 = n38603 & n38901;
  assign n38903 = pi1153 & ~n11358;
  assign n38904 = ~n38465 & ~n38903;
  assign n38905 = pi1154 & ~n38904;
  assign n38906 = ~n38807 & ~n38905;
  assign n38907 = pi207 & ~n38906;
  assign n38908 = ~n38718 & ~n38907;
  assign n38909 = ~pi208 & ~n38908;
  assign n38910 = ~pi207 & n38906;
  assign n38911 = ~pi299 & ~pi1153;
  assign n38912 = ~n10794 & ~n38911;
  assign n38913 = ~n38524 & n38912;
  assign n38914 = pi207 & ~n38913;
  assign n38915 = pi208 & ~n38914;
  assign n38916 = ~n38910 & n38915;
  assign n38917 = ~n38909 & ~n38916;
  assign n38918 = ~pi211 & n38917;
  assign n38919 = pi211 & n38901;
  assign n38920 = ~n38918 & ~n38919;
  assign n38921 = n38664 & ~n38920;
  assign n38922 = ~n38902 & ~n38921;
  assign n38923 = ~pi219 & ~n38922;
  assign n38924 = pi200 & ~pi1153;
  assign n38925 = n11348 & ~n38924;
  assign n38926 = ~n38808 & n38925;
  assign n38927 = n38708 & n38926;
  assign n38928 = pi208 & n38319;
  assign n38929 = pi1153 & ~n10794;
  assign n38930 = n38928 & n38929;
  assign n38931 = ~n38927 & ~n38930;
  assign n38932 = pi219 & n38931;
  assign n38933 = ~po1038 & ~n38932;
  assign n38934 = ~n38371 & ~n38664;
  assign n38935 = n38931 & n38934;
  assign n38936 = n38933 & ~n38935;
  assign n38937 = ~n38923 & n38936;
  assign n38938 = n38705 & ~n38937;
  assign n38939 = ~n38889 & ~n38938;
  assign n38940 = ~pi213 & n38939;
  assign n38941 = ~pi1152 & ~po1038;
  assign n38942 = ~pi299 & ~n38806;
  assign n38943 = ~pi1154 & ~n38942;
  assign n38944 = ~n38539 & n38943;
  assign n38945 = ~n38495 & n38905;
  assign n38946 = ~n38944 & ~n38945;
  assign n38947 = pi207 & n38946;
  assign n38948 = n38490 & ~n38947;
  assign n38949 = ~pi207 & n38946;
  assign n38950 = ~n38539 & n38912;
  assign n38951 = pi207 & ~n38950;
  assign n38952 = pi208 & ~n38951;
  assign n38953 = ~n38949 & n38952;
  assign n38954 = ~n38948 & ~n38953;
  assign n38955 = ~pi211 & n38954;
  assign n38956 = pi211 & n38917;
  assign n38957 = n10708 & ~n38955;
  assign n38958 = ~n38956 & n38957;
  assign n38959 = pi211 & n38954;
  assign n38960 = ~pi211 & ~n38576;
  assign n38961 = n38931 & n38960;
  assign n38962 = ~n38300 & ~n38961;
  assign n38963 = ~n38959 & n38962;
  assign n38964 = ~n38958 & ~n38963;
  assign n38965 = ~pi219 & ~n38964;
  assign n38966 = n38290 & ~n38931;
  assign n38967 = pi211 & n38931;
  assign n38968 = n38839 & ~n38967;
  assign n38969 = ~n38918 & n38968;
  assign n38970 = ~n38966 & ~n38969;
  assign n38971 = ~n38965 & n38970;
  assign n38972 = n38941 & ~n38971;
  assign n38973 = ~n38291 & n38835;
  assign n38974 = ~n38290 & n38856;
  assign n38975 = ~n38973 & ~n38974;
  assign n38976 = pi219 & ~n38975;
  assign n38977 = pi211 & ~n38855;
  assign n38978 = n38490 & ~n38812;
  assign n38979 = ~n38821 & ~n38978;
  assign n38980 = ~pi199 & ~pi1154;
  assign n38981 = ~pi200 & n38980;
  assign n38982 = n38521 & n38981;
  assign n38983 = ~n38539 & ~n38982;
  assign n38984 = ~n38979 & n38983;
  assign n38985 = ~pi211 & n38984;
  assign n38986 = n10708 & ~n38985;
  assign n38987 = ~n38977 & n38986;
  assign n38988 = pi211 & n38984;
  assign n38989 = ~n38576 & n38829;
  assign n38990 = ~pi207 & ~n38989;
  assign n38991 = pi299 & ~pi1156;
  assign n38992 = n38847 & ~n38991;
  assign n38993 = pi208 & ~n38992;
  assign n38994 = ~n38990 & n38993;
  assign n38995 = ~pi208 & ~n38576;
  assign n38996 = ~n38844 & n38995;
  assign n38997 = ~pi211 & ~n38996;
  assign n38998 = ~n38994 & n38997;
  assign n38999 = ~n38300 & ~n38998;
  assign n39000 = ~n38988 & n38999;
  assign n39001 = ~pi212 & n38882;
  assign n39002 = ~pi219 & ~n39001;
  assign n39003 = ~n39000 & n39002;
  assign n39004 = ~n38987 & n39003;
  assign n39005 = ~n38976 & ~n39004;
  assign n39006 = pi1152 & ~po1038;
  assign n39007 = ~n39005 & n39006;
  assign n39008 = ~n38972 & ~n39007;
  assign n39009 = pi213 & ~n39008;
  assign n39010 = ~pi209 & ~n39009;
  assign n39011 = ~n38940 & n39010;
  assign n39012 = ~n38804 & ~n39011;
  assign n39013 = pi214 & ~n38357;
  assign n39014 = ~pi212 & n39013;
  assign n39015 = ~pi219 & ~n39014;
  assign n39016 = ~n38364 & n39015;
  assign n39017 = pi219 & ~n38374;
  assign n39018 = pi213 & ~n39017;
  assign n39019 = n38293 & n39018;
  assign n39020 = ~n39016 & n39019;
  assign n39021 = ~n39012 & ~n39020;
  assign n39022 = pi230 & ~n39021;
  assign n39023 = ~pi230 & pi234;
  assign po391 = n39022 | n39023;
  assign n39025 = ~n38441 & ~n38541;
  assign n39026 = pi207 & ~n39025;
  assign n39027 = ~pi207 & n38497;
  assign n39028 = ~n39026 & ~n39027;
  assign n39029 = pi208 & ~n39028;
  assign n39030 = ~n38498 & ~n39029;
  assign n39031 = ~pi1157 & ~n39030;
  assign n39032 = pi208 & pi1157;
  assign n39033 = ~pi207 & ~n38488;
  assign n39034 = ~n39026 & ~n39033;
  assign n39035 = n39032 & ~n39034;
  assign n39036 = ~n38492 & ~n39035;
  assign n39037 = ~n39031 & n39036;
  assign n39038 = pi211 & ~n39037;
  assign n39039 = ~pi1156 & n38434;
  assign n39040 = ~n38537 & ~n39039;
  assign n39041 = pi207 & ~n39040;
  assign n39042 = ~pi207 & n38551;
  assign n39043 = ~n39041 & ~n39042;
  assign n39044 = pi208 & ~n39043;
  assign n39045 = ~n38581 & ~n39044;
  assign n39046 = ~pi1157 & ~n39045;
  assign n39047 = ~n38452 & ~n38518;
  assign n39048 = ~pi207 & ~n39047;
  assign n39049 = ~n39041 & ~n39048;
  assign n39050 = n39032 & ~n39049;
  assign n39051 = ~n38584 & ~n39050;
  assign n39052 = ~n39046 & n39051;
  assign n39053 = ~pi211 & ~n39052;
  assign n39054 = n10708 & ~n39038;
  assign n39055 = ~n39053 & n39054;
  assign n39056 = n10463 & ~n38441;
  assign n39057 = ~n39039 & n39056;
  assign n39058 = ~pi207 & ~n38412;
  assign n39059 = ~n39057 & ~n39058;
  assign n39060 = ~n38414 & n39059;
  assign n39061 = ~pi1157 & ~n39060;
  assign n39062 = ~pi207 & n38453;
  assign n39063 = ~n39057 & ~n39062;
  assign n39064 = ~n38455 & n39063;
  assign n39065 = pi1157 & ~n39064;
  assign n39066 = ~n39061 & ~n39065;
  assign n39067 = n38290 & ~n39066;
  assign n39068 = pi211 & ~n39052;
  assign n39069 = ~pi207 & n38519;
  assign n39070 = pi208 & ~n39069;
  assign n39071 = ~n38537 & n38731;
  assign n39072 = n39070 & ~n39071;
  assign n39073 = ~n38523 & ~n39072;
  assign n39074 = pi1157 & n39073;
  assign n39075 = ~pi211 & ~n39061;
  assign n39076 = ~n39074 & n39075;
  assign n39077 = n38664 & ~n39076;
  assign n39078 = ~n39068 & n39077;
  assign n39079 = ~n39067 & ~n39078;
  assign n39080 = ~n39055 & n39079;
  assign n39081 = ~pi219 & ~n39080;
  assign n39082 = ~pi211 & n39037;
  assign n39083 = pi211 & ~n39066;
  assign n39084 = ~n38300 & ~n39083;
  assign n39085 = ~n39082 & n39084;
  assign n39086 = n38300 & n39066;
  assign n39087 = pi219 & ~n39086;
  assign n39088 = ~n39085 & n39087;
  assign n39089 = pi209 & ~n39088;
  assign n39090 = ~n39081 & n39089;
  assign n39091 = n38522 & ~n38567;
  assign n39092 = n38521 & n38534;
  assign n39093 = ~n38905 & ~n38943;
  assign n39094 = pi207 & n39093;
  assign n39095 = pi208 & ~n39092;
  assign n39096 = ~n39094 & n39095;
  assign n39097 = ~n39091 & ~n39096;
  assign n39098 = pi1157 & ~n39097;
  assign n39099 = n10463 & ~n38926;
  assign n39100 = ~n38430 & ~n38707;
  assign n39101 = ~n10463 & ~n39100;
  assign n39102 = ~n39099 & ~n39101;
  assign n39103 = ~pi1157 & n39102;
  assign n39104 = ~pi211 & ~n39098;
  assign n39105 = ~n39103 & n39104;
  assign n39106 = ~n38576 & ~n39102;
  assign n39107 = pi211 & n39106;
  assign n39108 = ~n39105 & ~n39107;
  assign n39109 = n38664 & ~n39108;
  assign n39110 = ~n38474 & n38490;
  assign n39111 = ~pi207 & n38474;
  assign n39112 = pi208 & ~n38947;
  assign n39113 = ~n39111 & n39112;
  assign n39114 = ~n39110 & ~n39113;
  assign n39115 = pi211 & ~n39114;
  assign n39116 = ~pi211 & ~n39106;
  assign n39117 = n10708 & ~n39115;
  assign n39118 = ~n39116 & n39117;
  assign n39119 = n38290 & ~n39102;
  assign n39120 = ~n39118 & ~n39119;
  assign n39121 = ~n39109 & n39120;
  assign n39122 = ~pi219 & ~n39121;
  assign n39123 = ~pi211 & n39114;
  assign n39124 = pi211 & ~n39102;
  assign n39125 = ~n38300 & ~n39124;
  assign n39126 = ~n39123 & n39125;
  assign n39127 = n38300 & n39102;
  assign n39128 = pi219 & ~n39127;
  assign n39129 = ~n39126 & n39128;
  assign n39130 = ~pi209 & ~n39129;
  assign n39131 = ~n39122 & n39130;
  assign n39132 = ~n39090 & ~n39131;
  assign n39133 = ~po1038 & ~n39132;
  assign n39134 = ~pi214 & ~n38367;
  assign n39135 = ~n39013 & ~n39134;
  assign n39136 = pi212 & ~n39135;
  assign n39137 = ~pi219 & ~n39136;
  assign n39138 = ~n38368 & n39137;
  assign n39139 = pi219 & ~n38359;
  assign n39140 = pi219 & ~n38664;
  assign n39141 = ~n39139 & ~n39140;
  assign n39142 = po1038 & n39141;
  assign n39143 = ~n39138 & n39142;
  assign n39144 = pi213 & ~n39143;
  assign n39145 = ~n39133 & n39144;
  assign n39146 = pi1157 & ~n39073;
  assign n39147 = pi299 & ~pi1157;
  assign n39148 = ~n39146 & ~n39147;
  assign n39149 = ~n39046 & n39148;
  assign n39150 = ~n38544 & ~n39149;
  assign n39151 = ~pi211 & ~n39150;
  assign n39152 = n39084 & ~n39151;
  assign n39153 = n39087 & ~n39152;
  assign n39154 = pi211 & n39150;
  assign n39155 = ~n38435 & ~n38542;
  assign n39156 = ~n38441 & ~n39155;
  assign n39157 = pi207 & ~n39156;
  assign n39158 = pi1154 & ~n38550;
  assign n39159 = ~n38411 & ~n39158;
  assign n39160 = ~pi207 & ~n38493;
  assign n39161 = ~n39159 & n39160;
  assign n39162 = ~n39157 & ~n39161;
  assign n39163 = pi208 & ~n39162;
  assign n39164 = ~n38528 & ~n39163;
  assign n39165 = ~pi1157 & ~n39164;
  assign n39166 = n38525 & ~n39073;
  assign n39167 = ~n39165 & ~n39166;
  assign n39168 = ~pi211 & ~n39167;
  assign n39169 = n10708 & ~n39168;
  assign n39170 = ~n39154 & n39169;
  assign n39171 = pi211 & n39167;
  assign n39172 = ~n39082 & ~n39171;
  assign n39173 = n38664 & ~n39172;
  assign n39174 = ~n39067 & ~n39170;
  assign n39175 = ~n39173 & n39174;
  assign n39176 = ~pi219 & ~n39175;
  assign n39177 = ~n39153 & ~n39176;
  assign n39178 = pi209 & ~n39177;
  assign n39179 = ~n38535 & ~n38857;
  assign n39180 = ~pi208 & ~n39179;
  assign n39181 = ~pi207 & ~n38534;
  assign n39182 = ~n38893 & ~n39181;
  assign n39183 = pi208 & ~n39182;
  assign n39184 = ~n39180 & ~n39183;
  assign n39185 = ~pi211 & n39184;
  assign n39186 = n39125 & ~n39185;
  assign n39187 = n39128 & ~n39186;
  assign n39188 = ~n38512 & ~n38718;
  assign n39189 = ~pi208 & ~n39188;
  assign n39190 = ~pi207 & ~n38511;
  assign n39191 = ~n38907 & ~n39190;
  assign n39192 = pi208 & ~n39191;
  assign n39193 = ~n39189 & ~n39192;
  assign n39194 = pi211 & n39193;
  assign n39195 = ~n39123 & ~n39194;
  assign n39196 = ~n38300 & ~n39195;
  assign n39197 = ~pi211 & ~n39193;
  assign n39198 = pi211 & ~n39184;
  assign n39199 = n10708 & ~n39198;
  assign n39200 = ~n39197 & n39199;
  assign n39201 = ~n39119 & ~n39200;
  assign n39202 = ~n39196 & n39201;
  assign n39203 = ~pi219 & ~n39202;
  assign n39204 = ~n39187 & ~n39203;
  assign n39205 = ~pi209 & ~n39204;
  assign n39206 = ~po1038 & ~n39205;
  assign n39207 = ~n39178 & n39206;
  assign n39208 = pi219 & ~n38376;
  assign n39209 = po1038 & ~n39208;
  assign n39210 = ~n38361 & n38664;
  assign n39211 = n10708 & ~n38700;
  assign n39212 = ~pi219 & ~n39210;
  assign n39213 = ~n39211 & n39212;
  assign n39214 = ~n39140 & n39209;
  assign n39215 = ~n39213 & n39214;
  assign n39216 = ~pi213 & ~n39215;
  assign n39217 = ~n39207 & n39216;
  assign n39218 = ~n39145 & ~n39217;
  assign n39219 = pi230 & ~n39218;
  assign n39220 = ~pi230 & ~pi235;
  assign po392 = ~n39219 & ~n39220;
  assign n39222 = ~pi100 & n38063;
  assign n39223 = n38274 & ~n39222;
  assign n39224 = ~n6277 & ~n39223;
  assign n39225 = ~pi75 & ~n39224;
  assign n39226 = ~n7292 & ~n39225;
  assign n39227 = ~pi92 & ~n39226;
  assign n39228 = n13616 & ~n39227;
  assign n39229 = ~pi74 & ~n39228;
  assign n39230 = n6116 & ~n39229;
  assign n39231 = ~pi56 & ~n39230;
  assign n39232 = ~n6112 & ~n39231;
  assign n39233 = ~pi62 & ~n39232;
  assign po393 = n13624 & ~n39233;
  assign n39235 = pi211 & pi1157;
  assign n39236 = ~pi211 & pi1158;
  assign n39237 = ~n39235 & ~n39236;
  assign n39238 = n38298 & ~n39237;
  assign n39239 = n39137 & ~n39238;
  assign n39240 = ~pi219 & po1038;
  assign n39241 = n38298 & n38355;
  assign n39242 = po1038 & n39241;
  assign n39243 = ~n39240 & ~n39242;
  assign n39244 = pi214 & n38374;
  assign n39245 = pi1155 & n38503;
  assign n39246 = ~n39244 & ~n39245;
  assign n39247 = pi212 & ~n39246;
  assign n39248 = po1038 & n39247;
  assign n39249 = n39243 & ~n39248;
  assign n39250 = ~n39239 & ~n39249;
  assign n39251 = ~pi213 & ~n39250;
  assign n39252 = n38384 & ~n39239;
  assign n39253 = pi199 & pi1143;
  assign n39254 = ~pi200 & ~n39253;
  assign n39255 = ~n38311 & n39254;
  assign n39256 = ~n38314 & n38928;
  assign n39257 = ~n39255 & n39256;
  assign n39258 = ~pi199 & pi1145;
  assign n39259 = n39254 & ~n39258;
  assign n39260 = pi200 & ~n38311;
  assign n39261 = n38708 & ~n39260;
  assign n39262 = ~n39259 & n39261;
  assign n39263 = ~n39257 & ~n39262;
  assign n39264 = ~pi299 & ~n39263;
  assign n39265 = n38298 & n38576;
  assign n39266 = pi214 & ~n38390;
  assign n39267 = ~pi214 & ~n38386;
  assign n39268 = pi212 & ~n39266;
  assign n39269 = ~n39267 & n39268;
  assign n39270 = ~n39265 & ~n39269;
  assign n39271 = n38395 & ~n39270;
  assign n39272 = ~n39264 & ~n39271;
  assign n39273 = ~n39252 & n39272;
  assign n39274 = ~po1038 & ~n39273;
  assign n39275 = n39251 & ~n39274;
  assign n39276 = n10708 & n38297;
  assign n39277 = ~pi211 & pi1145;
  assign n39278 = pi211 & pi1144;
  assign n39279 = ~n39277 & ~n39278;
  assign n39280 = ~n10708 & n39279;
  assign n39281 = ~n38290 & ~n39276;
  assign n39282 = ~n39280 & n39281;
  assign n39283 = ~pi219 & ~n39282;
  assign n39284 = pi219 & ~n38302;
  assign n39285 = n38293 & ~n39284;
  assign n39286 = ~n39283 & n39285;
  assign n39287 = n38384 & n39282;
  assign n39288 = pi299 & n38839;
  assign n39289 = n38302 & n39288;
  assign n39290 = ~n39264 & ~n39289;
  assign n39291 = ~n39287 & n39290;
  assign n39292 = ~po1038 & ~n39291;
  assign n39293 = ~n39286 & ~n39292;
  assign n39294 = pi213 & n39293;
  assign n39295 = pi209 & ~n39275;
  assign n39296 = ~n39294 & n39295;
  assign n39297 = pi1158 & n38824;
  assign n39298 = ~pi199 & ~pi1158;
  assign n39299 = pi1156 & ~n39298;
  assign n39300 = ~n39297 & ~n39299;
  assign n39301 = n38326 & n38424;
  assign n39302 = ~n39300 & n39301;
  assign n39303 = pi207 & n38442;
  assign n39304 = pi208 & ~n39058;
  assign n39305 = ~n39303 & n39304;
  assign n39306 = ~n39302 & ~n39305;
  assign n39307 = ~pi1157 & ~n39306;
  assign n39308 = pi1156 & n38483;
  assign n39309 = ~pi200 & ~pi1158;
  assign n39310 = ~pi199 & ~n39309;
  assign n39311 = ~n39308 & ~n39310;
  assign n39312 = n38319 & ~n39311;
  assign n39313 = ~pi208 & n39312;
  assign n39314 = pi208 & ~n39062;
  assign n39315 = ~n39303 & n39314;
  assign n39316 = ~n39313 & ~n39315;
  assign n39317 = pi1157 & ~n39316;
  assign n39318 = ~n39307 & ~n39317;
  assign n39319 = ~n38291 & n39318;
  assign n39320 = ~n38778 & ~n39048;
  assign n39321 = n39032 & ~n39320;
  assign n39322 = pi208 & ~n39042;
  assign n39323 = ~n38778 & n39322;
  assign n39324 = ~pi200 & pi207;
  assign n39325 = ~n39300 & n39324;
  assign n39326 = n38995 & ~n39325;
  assign n39327 = ~pi1157 & ~n39326;
  assign n39328 = ~n39323 & n39327;
  assign n39329 = ~n38576 & ~n39312;
  assign n39330 = n38582 & ~n39329;
  assign n39331 = ~n39321 & ~n39330;
  assign n39332 = ~n39328 & n39331;
  assign n39333 = n38298 & n39332;
  assign n39334 = ~n38386 & n38442;
  assign n39335 = pi207 & ~n39334;
  assign n39336 = ~n39027 & ~n39335;
  assign n39337 = pi208 & ~n39336;
  assign n39338 = ~pi208 & n38386;
  assign n39339 = ~n39302 & ~n39338;
  assign n39340 = ~n39337 & n39339;
  assign n39341 = ~pi1157 & ~n39340;
  assign n39342 = ~n39033 & ~n39335;
  assign n39343 = n39032 & ~n39342;
  assign n39344 = pi1156 & ~n38867;
  assign n39345 = ~pi1158 & ~n38410;
  assign n39346 = n39344 & ~n39345;
  assign n39347 = ~n39310 & ~n39346;
  assign n39348 = n38319 & ~n39347;
  assign n39349 = ~n38386 & ~n39348;
  assign n39350 = n38582 & ~n39349;
  assign n39351 = ~n39343 & ~n39350;
  assign n39352 = ~n39341 & n39351;
  assign n39353 = ~pi214 & ~n39352;
  assign n39354 = ~pi207 & ~n38519;
  assign n39355 = ~n38524 & n39354;
  assign n39356 = pi1157 & ~n39355;
  assign n39357 = ~pi1157 & ~n39302;
  assign n39358 = ~n39161 & n39357;
  assign n39359 = ~n39356 & ~n39358;
  assign n39360 = pi208 & ~n38719;
  assign n39361 = ~n39359 & n39360;
  assign n39362 = n39348 & ~n39357;
  assign n39363 = ~pi208 & ~n38390;
  assign n39364 = ~n39362 & n39363;
  assign n39365 = pi214 & ~n39364;
  assign n39366 = ~n39361 & n39365;
  assign n39367 = pi212 & ~n39366;
  assign n39368 = ~n39353 & n39367;
  assign n39369 = ~n39333 & ~n39368;
  assign n39370 = ~pi211 & ~n39369;
  assign n39371 = ~n39319 & ~n39370;
  assign n39372 = pi219 & ~n39371;
  assign n39373 = ~pi214 & n39318;
  assign n39374 = ~pi212 & ~n39373;
  assign n39375 = ~pi299 & n39311;
  assign n39376 = n38522 & ~n39375;
  assign n39377 = ~n38732 & n39070;
  assign n39378 = ~n39376 & ~n39377;
  assign n39379 = pi1157 & ~n39378;
  assign n39380 = ~n39307 & ~n39379;
  assign n39381 = pi211 & n39380;
  assign n39382 = pi1158 & n38543;
  assign n39383 = ~pi1158 & n38442;
  assign n39384 = pi207 & ~n39383;
  assign n39385 = ~n39382 & n39384;
  assign n39386 = ~pi299 & ~n38551;
  assign n39387 = pi299 & ~pi1158;
  assign n39388 = ~pi207 & ~n39387;
  assign n39389 = ~n39386 & n39388;
  assign n39390 = pi208 & ~n39389;
  assign n39391 = ~n39385 & n39390;
  assign n39392 = ~pi299 & ~n38897;
  assign n39393 = pi1158 & ~n39392;
  assign n39394 = n38319 & n39308;
  assign n39395 = ~pi208 & ~n39394;
  assign n39396 = ~n39393 & n39395;
  assign n39397 = ~pi1157 & ~n39396;
  assign n39398 = ~n39391 & n39397;
  assign n39399 = n39354 & ~n39387;
  assign n39400 = ~n39385 & ~n39399;
  assign n39401 = n39032 & ~n39400;
  assign n39402 = n38410 & ~n38486;
  assign n39403 = pi1157 & ~n39297;
  assign n39404 = ~n39402 & n39403;
  assign n39405 = pi207 & ~n39404;
  assign n39406 = ~n39393 & ~n39405;
  assign n39407 = n38582 & ~n39406;
  assign n39408 = ~pi211 & ~n39407;
  assign n39409 = ~n39398 & n39408;
  assign n39410 = ~n39401 & n39409;
  assign n39411 = ~n39381 & ~n39410;
  assign n39412 = pi214 & ~n39411;
  assign n39413 = n39374 & ~n39412;
  assign n39414 = n10654 & ~n39352;
  assign n39415 = n38503 & ~n39380;
  assign n39416 = n38592 & ~n39332;
  assign n39417 = ~n39414 & ~n39416;
  assign n39418 = ~n39415 & n39417;
  assign n39419 = pi212 & ~n39418;
  assign n39420 = ~pi219 & ~n39419;
  assign n39421 = ~n39413 & n39420;
  assign n39422 = ~po1038 & ~n39372;
  assign n39423 = ~n39421 & n39422;
  assign n39424 = n39251 & ~n39423;
  assign n39425 = pi299 & ~pi1145;
  assign n39426 = ~n38505 & ~n39425;
  assign n39427 = pi1154 & ~n39426;
  assign n39428 = pi299 & pi1145;
  assign n39429 = n38435 & ~n39428;
  assign n39430 = ~pi1156 & ~n39429;
  assign n39431 = ~n39427 & n39430;
  assign n39432 = ~n38536 & ~n39425;
  assign n39433 = ~pi1154 & ~n39432;
  assign n39434 = n38618 & ~n39428;
  assign n39435 = pi1156 & ~n39434;
  assign n39436 = ~n39433 & n39435;
  assign n39437 = ~n39431 & ~n39436;
  assign n39438 = pi207 & ~n39437;
  assign n39439 = ~pi200 & pi1157;
  assign n39440 = ~pi199 & n39439;
  assign n39441 = n39386 & ~n39440;
  assign n39442 = ~pi207 & ~n39425;
  assign n39443 = ~n39441 & n39442;
  assign n39444 = pi208 & ~n39443;
  assign n39445 = ~n39438 & n39444;
  assign n39446 = ~pi299 & n39308;
  assign n39447 = ~pi1157 & ~n39297;
  assign n39448 = ~n39446 & n39447;
  assign n39449 = n39405 & ~n39448;
  assign n39450 = ~pi208 & ~n39428;
  assign n39451 = ~n39449 & n39450;
  assign n39452 = ~n39445 & ~n39451;
  assign n39453 = ~pi211 & ~n39452;
  assign n39454 = ~pi1157 & ~n39325;
  assign n39455 = ~pi208 & ~n39454;
  assign n39456 = n39348 & n39455;
  assign n39457 = ~pi208 & ~n39456;
  assign n39458 = ~n38637 & n39457;
  assign n39459 = pi207 & ~n38652;
  assign n39460 = ~pi207 & ~n38639;
  assign n39461 = ~n39441 & n39460;
  assign n39462 = pi208 & ~n39461;
  assign n39463 = ~n39459 & n39462;
  assign n39464 = ~n39458 & ~n39463;
  assign n39465 = pi211 & ~n39464;
  assign n39466 = ~n39453 & ~n39465;
  assign n39467 = pi214 & ~n39466;
  assign n39468 = n39374 & ~n39467;
  assign n39469 = ~pi214 & ~n39466;
  assign n39470 = ~pi211 & n39464;
  assign n39471 = ~n38604 & n39457;
  assign n39472 = pi207 & ~n38622;
  assign n39473 = ~pi207 & ~n38606;
  assign n39474 = ~n39441 & n39473;
  assign n39475 = pi208 & ~n39474;
  assign n39476 = ~n39472 & n39475;
  assign n39477 = ~n39471 & ~n39476;
  assign n39478 = pi211 & n39477;
  assign n39479 = pi214 & ~n39470;
  assign n39480 = ~n39478 & n39479;
  assign n39481 = pi212 & ~n39480;
  assign n39482 = ~n39469 & n39481;
  assign n39483 = ~pi219 & ~n39468;
  assign n39484 = ~n39482 & n39483;
  assign n39485 = n38291 & ~n39477;
  assign n39486 = ~n39319 & ~n39485;
  assign n39487 = pi219 & ~n39486;
  assign n39488 = ~po1038 & ~n39487;
  assign n39489 = ~n39484 & n39488;
  assign n39490 = pi213 & ~n39286;
  assign n39491 = ~n39489 & n39490;
  assign n39492 = ~pi209 & ~n39491;
  assign n39493 = ~n39424 & n39492;
  assign n39494 = ~n39296 & ~n39493;
  assign n39495 = pi230 & ~n39494;
  assign n39496 = ~pi230 & ~pi237;
  assign po394 = n39495 | n39496;
  assign n39498 = ~pi211 & ~pi1153;
  assign n39499 = pi219 & n39498;
  assign n39500 = n38293 & ~n39499;
  assign n39501 = ~n39213 & n39500;
  assign n39502 = ~n10463 & n38424;
  assign n39503 = ~n38707 & n39502;
  assign n39504 = n38409 & n38928;
  assign n39505 = ~n39503 & ~n39504;
  assign n39506 = ~n38831 & ~n39505;
  assign n39507 = ~pi214 & ~n39506;
  assign n39508 = ~pi212 & ~n39507;
  assign n39509 = n38424 & ~n38827;
  assign n39510 = ~pi1153 & ~n38484;
  assign n39511 = ~n38464 & ~n39510;
  assign n39512 = pi1155 & ~n39511;
  assign n39513 = ~n39509 & ~n39512;
  assign n39514 = n38319 & ~n38409;
  assign n39515 = pi208 & ~n39514;
  assign n39516 = ~n38490 & ~n39515;
  assign n39517 = ~n39513 & ~n39516;
  assign n39518 = ~n39504 & ~n39517;
  assign n39519 = ~pi299 & ~n39518;
  assign n39520 = pi299 & ~n38361;
  assign n39521 = pi214 & ~n39520;
  assign n39522 = ~n39519 & n39521;
  assign n39523 = n39508 & ~n39522;
  assign n39524 = n38503 & n39518;
  assign n39525 = ~pi299 & ~n39324;
  assign n39526 = ~pi208 & ~n39525;
  assign n39527 = pi200 & n38521;
  assign n39528 = n39515 & ~n39527;
  assign n39529 = ~n39526 & ~n39528;
  assign n39530 = ~n38465 & ~n39529;
  assign n39531 = n10654 & ~n39530;
  assign n39532 = ~n38390 & n38592;
  assign n39533 = ~n39506 & n39532;
  assign n39534 = pi212 & ~n39533;
  assign n39535 = ~n39531 & n39534;
  assign n39536 = ~n39524 & n39535;
  assign n39537 = ~pi219 & ~n39536;
  assign n39538 = ~n39523 & n39537;
  assign n39539 = pi1151 & ~po1038;
  assign n39540 = ~pi211 & ~n39529;
  assign n39541 = pi211 & ~n39505;
  assign n39542 = ~n39540 & ~n39541;
  assign n39543 = ~n38465 & ~n39542;
  assign n39544 = n38290 & ~n39506;
  assign n39545 = n39543 & ~n39544;
  assign n39546 = pi219 & ~n39545;
  assign n39547 = n39539 & ~n39546;
  assign n39548 = ~n39538 & n39547;
  assign n39549 = n38708 & n38824;
  assign n39550 = pi1153 & n39549;
  assign n39551 = ~n38390 & ~n39550;
  assign n39552 = ~pi211 & ~n39551;
  assign n39553 = n10793 & n38708;
  assign n39554 = ~pi299 & ~n39553;
  assign n39555 = n38699 & ~n39554;
  assign n39556 = n10708 & ~n39555;
  assign n39557 = ~n39552 & n39556;
  assign n39558 = ~n38300 & ~n39520;
  assign n39559 = ~n39550 & n39558;
  assign n39560 = ~n39557 & ~n39559;
  assign n39561 = ~pi219 & ~n39560;
  assign n39562 = ~pi1151 & ~po1038;
  assign n39563 = ~n13025 & ~n39554;
  assign n39564 = ~pi214 & ~n39549;
  assign n39565 = ~pi212 & n39564;
  assign n39566 = n39563 & ~n39565;
  assign n39567 = pi1153 & n39566;
  assign n39568 = ~n38669 & ~n39567;
  assign n39569 = n39562 & ~n39568;
  assign n39570 = ~n39561 & n39569;
  assign n39571 = ~pi1152 & ~n39570;
  assign n39572 = ~n39548 & n39571;
  assign n39573 = pi1153 & ~n39554;
  assign n39574 = ~n38708 & ~n38897;
  assign n39575 = ~n10463 & n38540;
  assign n39576 = ~n39574 & ~n39575;
  assign n39577 = n39554 & n39576;
  assign n39578 = ~n39573 & ~n39577;
  assign n39579 = pi211 & ~n39578;
  assign n39580 = ~pi207 & ~n38817;
  assign n39581 = ~n38897 & ~n39580;
  assign n39582 = pi208 & ~n39581;
  assign n39583 = n38522 & ~n38817;
  assign n39584 = ~n39582 & ~n39583;
  assign n39585 = ~pi211 & ~n38524;
  assign n39586 = ~n39584 & n39585;
  assign n39587 = ~n39579 & ~n39586;
  assign n39588 = n10708 & ~n39587;
  assign n39589 = pi299 & n38361;
  assign n39590 = ~n38300 & ~n39584;
  assign n39591 = ~n39589 & n39590;
  assign n39592 = ~n39588 & ~n39591;
  assign n39593 = ~pi219 & ~n39592;
  assign n39594 = ~n10463 & n38815;
  assign n39595 = ~n38708 & ~n39324;
  assign n39596 = n11348 & ~n39595;
  assign n39597 = ~n39594 & n39596;
  assign n39598 = ~pi211 & n38388;
  assign n39599 = ~n38290 & n39598;
  assign n39600 = ~n39597 & ~n39599;
  assign n39601 = ~n38669 & ~n39600;
  assign n39602 = ~n39593 & ~n39601;
  assign n39603 = n39562 & ~n39602;
  assign n39604 = n38818 & ~n38868;
  assign n39605 = pi208 & ~n39604;
  assign n39606 = n38522 & ~n38819;
  assign n39607 = ~n39605 & ~n39606;
  assign n39608 = ~pi211 & ~n39607;
  assign n39609 = ~n38539 & n39608;
  assign n39610 = pi211 & ~n39607;
  assign n39611 = ~n38524 & n39610;
  assign n39612 = ~n39609 & ~n39611;
  assign n39613 = ~n38300 & ~n39612;
  assign n39614 = n38415 & ~n38707;
  assign n39615 = ~n39549 & n39614;
  assign n39616 = ~n39555 & ~n39615;
  assign n39617 = ~n39586 & n39616;
  assign n39618 = n10708 & ~n39617;
  assign n39619 = ~pi214 & ~n39615;
  assign n39620 = ~n39550 & n39619;
  assign n39621 = ~pi212 & ~n39620;
  assign n39622 = ~pi214 & n39621;
  assign n39623 = ~pi219 & ~n39622;
  assign n39624 = ~n39618 & n39623;
  assign n39625 = ~n39613 & n39624;
  assign n39626 = pi219 & ~n39615;
  assign n39627 = ~n39567 & n39626;
  assign n39628 = n39539 & ~n39627;
  assign n39629 = ~n39625 & n39628;
  assign n39630 = pi1152 & ~n39629;
  assign n39631 = ~n39603 & n39630;
  assign n39632 = ~n39572 & ~n39631;
  assign n39633 = ~pi209 & ~n39632;
  assign n39634 = n38410 & n38890;
  assign n39635 = n38850 & ~n39634;
  assign n39636 = pi207 & ~n39635;
  assign n39637 = ~n39190 & ~n39636;
  assign n39638 = pi208 & ~n39637;
  assign n39639 = ~n39189 & ~n39638;
  assign n39640 = pi211 & ~n39639;
  assign n39641 = ~n38415 & n38951;
  assign n39642 = ~pi1154 & ~n38911;
  assign n39643 = ~n38494 & n39642;
  assign n39644 = pi207 & ~n39643;
  assign n39645 = n38850 & n39644;
  assign n39646 = pi208 & ~n39645;
  assign n39647 = ~n39641 & n39646;
  assign n39648 = ~n39111 & n39647;
  assign n39649 = ~n39110 & ~n39648;
  assign n39650 = ~pi211 & ~n39649;
  assign n39651 = n38298 & ~n39650;
  assign n39652 = ~n39640 & n39651;
  assign n39653 = n38592 & ~n39639;
  assign n39654 = n38503 & ~n39649;
  assign n39655 = pi1153 & ~n38494;
  assign n39656 = ~n38826 & ~n39655;
  assign n39657 = pi207 & ~n39656;
  assign n39658 = ~n39181 & ~n39657;
  assign n39659 = pi208 & ~n39658;
  assign n39660 = ~n39180 & ~n39659;
  assign n39661 = n10654 & ~n39660;
  assign n39662 = pi212 & ~n39661;
  assign n39663 = ~n39654 & n39662;
  assign n39664 = ~n39653 & n39663;
  assign n39665 = ~n39652 & ~n39664;
  assign n39666 = ~pi219 & ~n39665;
  assign n39667 = n10463 & ~n39634;
  assign n39668 = ~n38826 & n39667;
  assign n39669 = ~n39101 & ~n39668;
  assign n39670 = pi211 & n39669;
  assign n39671 = ~pi211 & ~n39660;
  assign n39672 = ~n39670 & ~n39671;
  assign n39673 = n38839 & n39672;
  assign n39674 = ~pi214 & ~n39669;
  assign n39675 = ~pi212 & n39674;
  assign n39676 = ~po1038 & ~n39675;
  assign n39677 = ~n39673 & n39676;
  assign n39678 = ~n39666 & n39677;
  assign n39679 = pi209 & ~n39678;
  assign n39680 = ~n39633 & ~n39679;
  assign n39681 = ~n39501 & ~n39680;
  assign n39682 = pi213 & ~n39681;
  assign n39683 = ~pi211 & n38664;
  assign n39684 = pi1153 & n39683;
  assign n39685 = n10656 & ~n39684;
  assign n39686 = n38293 & ~n39685;
  assign n39687 = pi1151 & ~n39686;
  assign n39688 = ~n39092 & n39646;
  assign n39689 = ~n39091 & ~n39688;
  assign n39690 = ~pi211 & ~n39689;
  assign n39691 = ~n39670 & ~n39690;
  assign n39692 = ~n38290 & n39691;
  assign n39693 = ~n39675 & ~n39692;
  assign n39694 = pi219 & ~n39693;
  assign n39695 = ~po1038 & ~n39694;
  assign n39696 = pi214 & n39672;
  assign n39697 = ~n39674 & ~n39696;
  assign n39698 = ~pi212 & ~n39697;
  assign n39699 = ~pi214 & ~n39672;
  assign n39700 = pi211 & ~n39689;
  assign n39701 = ~pi211 & n39669;
  assign n39702 = ~n39700 & ~n39701;
  assign n39703 = pi214 & ~n39702;
  assign n39704 = pi212 & ~n39699;
  assign n39705 = ~n39703 & n39704;
  assign n39706 = ~n39698 & ~n39705;
  assign n39707 = ~pi219 & ~n39706;
  assign n39708 = n39695 & ~n39707;
  assign n39709 = n39687 & ~n39708;
  assign n39710 = n39240 & n39684;
  assign n39711 = ~pi1151 & ~n39710;
  assign n39712 = ~pi219 & n38664;
  assign n39713 = n39672 & n39712;
  assign n39714 = ~n39669 & ~n39712;
  assign n39715 = ~po1038 & ~n39714;
  assign n39716 = ~n39713 & n39715;
  assign n39717 = n39711 & ~n39716;
  assign n39718 = ~pi1152 & ~n39717;
  assign n39719 = ~n39709 & n39718;
  assign n39720 = ~n10655 & n38669;
  assign n39721 = po1038 & n39720;
  assign n39722 = ~n10708 & ~n39498;
  assign n39723 = ~n38603 & ~n39722;
  assign n39724 = n39721 & ~n39723;
  assign n39725 = ~pi1151 & ~n39724;
  assign n39726 = ~n39671 & ~n39700;
  assign n39727 = pi214 & n39726;
  assign n39728 = ~pi212 & ~n39674;
  assign n39729 = ~n39727 & n39728;
  assign n39730 = ~pi219 & ~n39729;
  assign n39731 = ~pi214 & ~n39726;
  assign n39732 = pi214 & ~n39691;
  assign n39733 = ~n39731 & ~n39732;
  assign n39734 = pi212 & ~n39733;
  assign n39735 = n39730 & ~n39734;
  assign n39736 = pi219 & ~n39669;
  assign n39737 = ~po1038 & ~n39736;
  assign n39738 = ~n39735 & n39737;
  assign n39739 = n39725 & ~n39738;
  assign n39740 = ~n10656 & n38293;
  assign n39741 = pi1151 & ~n39740;
  assign n39742 = ~n39724 & n39741;
  assign n39743 = pi214 & ~n39689;
  assign n39744 = ~n39731 & ~n39743;
  assign n39745 = pi212 & ~n39744;
  assign n39746 = n39730 & ~n39745;
  assign n39747 = n39695 & ~n39746;
  assign n39748 = n39742 & ~n39747;
  assign n39749 = pi1152 & ~n39739;
  assign n39750 = ~n39748 & n39749;
  assign n39751 = pi209 & ~n39719;
  assign n39752 = ~n39750 & n39751;
  assign n39753 = ~pi214 & n39543;
  assign n39754 = ~n13025 & ~n39550;
  assign n39755 = ~n39506 & n39754;
  assign n39756 = pi214 & ~n39755;
  assign n39757 = pi212 & ~n39756;
  assign n39758 = ~n39753 & n39757;
  assign n39759 = ~pi212 & ~n39545;
  assign n39760 = ~n39758 & ~n39759;
  assign n39761 = ~pi219 & ~n39760;
  assign n39762 = ~pi211 & pi299;
  assign n39763 = ~n39550 & ~n39762;
  assign n39764 = ~n39506 & n39763;
  assign n39765 = ~n39544 & ~n39764;
  assign n39766 = pi219 & ~n39765;
  assign n39767 = ~po1038 & ~n39766;
  assign n39768 = ~n39761 & n39767;
  assign n39769 = n39687 & ~n39768;
  assign n39770 = n39564 & n39567;
  assign n39771 = ~pi214 & n13025;
  assign n39772 = pi212 & ~n39771;
  assign n39773 = ~n39754 & n39772;
  assign n39774 = ~pi219 & ~n39773;
  assign n39775 = n38298 & n39598;
  assign n39776 = ~n39549 & ~n39775;
  assign n39777 = n39774 & n39776;
  assign n39778 = ~n39770 & n39777;
  assign n39779 = pi219 & ~n39549;
  assign n39780 = ~po1038 & ~n39779;
  assign n39781 = n39567 & n39780;
  assign n39782 = ~n39778 & n39781;
  assign n39783 = n39711 & ~n39782;
  assign n39784 = ~pi1152 & ~n39783;
  assign n39785 = ~n39769 & n39784;
  assign n39786 = ~n39550 & ~n39615;
  assign n39787 = ~n39608 & n39786;
  assign n39788 = pi214 & n39787;
  assign n39789 = ~n39620 & ~n39788;
  assign n39790 = ~pi212 & ~n39789;
  assign n39791 = ~n39787 & ~n39790;
  assign n39792 = pi219 & ~n39791;
  assign n39793 = ~po1038 & ~n39792;
  assign n39794 = ~n39573 & ~n39610;
  assign n39795 = pi214 & ~n39615;
  assign n39796 = n39794 & n39795;
  assign n39797 = n39621 & ~n39796;
  assign n39798 = n39619 & n39794;
  assign n39799 = pi214 & n39607;
  assign n39800 = pi212 & ~n39799;
  assign n39801 = ~n39798 & n39800;
  assign n39802 = ~pi219 & ~n39797;
  assign n39803 = ~n39801 & n39802;
  assign n39804 = n39793 & ~n39803;
  assign n39805 = n39742 & ~n39804;
  assign n39806 = pi219 & ~n39597;
  assign n39807 = ~po1038 & ~n39806;
  assign n39808 = ~pi211 & n39578;
  assign n39809 = n39590 & ~n39808;
  assign n39810 = ~n38664 & n39597;
  assign n39811 = pi299 & n38603;
  assign n39812 = ~pi219 & ~n39811;
  assign n39813 = ~n39810 & n39812;
  assign n39814 = ~n39809 & n39813;
  assign n39815 = n39807 & ~n39814;
  assign n39816 = n39725 & ~n39815;
  assign n39817 = pi1152 & ~n39816;
  assign n39818 = ~n39805 & n39817;
  assign n39819 = ~n39785 & ~n39818;
  assign n39820 = ~pi209 & n39819;
  assign n39821 = ~pi213 & ~n39820;
  assign n39822 = ~n39752 & n39821;
  assign n39823 = ~n39682 & ~n39822;
  assign n39824 = pi230 & ~n39823;
  assign n39825 = ~pi230 & pi238;
  assign po395 = n39824 | n39825;
  assign n39827 = n38326 & ~n38442;
  assign n39828 = ~pi214 & n39827;
  assign n39829 = ~pi212 & ~n39828;
  assign n39830 = ~pi219 & n39829;
  assign n39831 = pi299 & pi1158;
  assign n39832 = ~n38326 & n39831;
  assign n39833 = ~pi208 & n39385;
  assign n39834 = ~n39832 & ~n39833;
  assign n39835 = ~pi211 & ~n39834;
  assign n39836 = pi208 & pi299;
  assign n39837 = pi1157 & ~n39836;
  assign n39838 = ~n38733 & n39837;
  assign n39839 = ~pi1157 & ~n39827;
  assign n39840 = pi211 & ~n39839;
  assign n39841 = ~n39838 & n39840;
  assign n39842 = ~n39835 & ~n39841;
  assign n39843 = pi214 & ~n39842;
  assign n39844 = n39830 & ~n39843;
  assign n39845 = pi219 & n39829;
  assign n39846 = pi211 & ~n39827;
  assign n39847 = pi214 & ~n39846;
  assign n39848 = ~n38780 & n38960;
  assign n39849 = n39847 & ~n39848;
  assign n39850 = n39845 & ~n39849;
  assign n39851 = pi212 & ~n39827;
  assign n39852 = ~po1038 & ~n39851;
  assign n39853 = ~pi209 & n39852;
  assign n39854 = ~n39850 & n39853;
  assign n39855 = ~n39844 & n39854;
  assign n39856 = n39313 & ~n39357;
  assign n39857 = ~pi214 & n39856;
  assign n39858 = ~pi212 & ~n39857;
  assign n39859 = ~pi219 & n39858;
  assign n39860 = pi208 & ~n39831;
  assign n39861 = ~n38582 & ~n39860;
  assign n39862 = ~n39396 & n39861;
  assign n39863 = n39408 & ~n39862;
  assign n39864 = ~n39376 & n39837;
  assign n39865 = ~n39357 & ~n39864;
  assign n39866 = pi211 & ~n39865;
  assign n39867 = pi214 & ~n39866;
  assign n39868 = ~n39863 & n39867;
  assign n39869 = n39859 & ~n39868;
  assign n39870 = pi219 & n39858;
  assign n39871 = pi211 & ~n39856;
  assign n39872 = n38960 & ~n39856;
  assign n39873 = pi214 & ~n39872;
  assign n39874 = ~n39871 & n39873;
  assign n39875 = n39870 & ~n39874;
  assign n39876 = pi212 & ~n39856;
  assign n39877 = ~po1038 & ~n39876;
  assign n39878 = pi209 & n39877;
  assign n39879 = ~n39875 & n39878;
  assign n39880 = ~n39869 & n39879;
  assign n39881 = ~pi219 & ~n39238;
  assign n39882 = ~n39243 & ~n39881;
  assign n39883 = pi213 & ~n39882;
  assign n39884 = ~n39880 & n39883;
  assign n39885 = ~n39855 & n39884;
  assign n39886 = pi211 & ~n38386;
  assign n39887 = ~n39456 & n39886;
  assign n39888 = n39873 & ~n39887;
  assign n39889 = n39859 & ~n39888;
  assign n39890 = ~pi211 & ~n38390;
  assign n39891 = ~n39456 & n39890;
  assign n39892 = pi214 & ~n39871;
  assign n39893 = ~n39891 & n39892;
  assign n39894 = n39870 & ~n39893;
  assign n39895 = n39877 & ~n39889;
  assign n39896 = ~n39894 & n39895;
  assign n39897 = pi209 & ~n39896;
  assign n39898 = ~n38390 & ~n38721;
  assign n39899 = n39847 & ~n39898;
  assign n39900 = n39845 & ~n39899;
  assign n39901 = ~n39827 & n39886;
  assign n39902 = pi214 & ~n39901;
  assign n39903 = ~n39848 & n39902;
  assign n39904 = n39830 & ~n39903;
  assign n39905 = n39852 & ~n39904;
  assign n39906 = ~n39900 & n39905;
  assign n39907 = ~pi209 & ~n39906;
  assign n39908 = ~n39897 & ~n39907;
  assign n39909 = po1038 & ~n39017;
  assign n39910 = n38298 & ~n39015;
  assign n39911 = n39909 & n39910;
  assign n39912 = ~pi213 & ~n39911;
  assign n39913 = ~n39908 & n39912;
  assign n39914 = ~n39885 & ~n39913;
  assign n39915 = pi230 & ~n39914;
  assign n39916 = ~pi230 & ~pi239;
  assign po396 = ~n39915 & ~n39916;
  assign n39918 = ~po1038 & n39596;
  assign n39919 = ~n39780 & ~n39918;
  assign n39920 = ~pi214 & ~n39596;
  assign n39921 = ~pi212 & ~n39920;
  assign n39922 = pi200 & pi207;
  assign n39923 = ~pi199 & ~n39922;
  assign n39924 = ~pi299 & ~n39923;
  assign n39925 = pi208 & ~n39924;
  assign n39926 = n11348 & n38326;
  assign n39927 = ~pi299 & ~n39926;
  assign n39928 = ~n39925 & n39927;
  assign n39929 = pi214 & n39928;
  assign n39930 = n39921 & ~n39929;
  assign n39931 = ~pi219 & ~n39930;
  assign n39932 = ~pi211 & ~n39928;
  assign n39933 = pi211 & n39596;
  assign n39934 = pi214 & ~n39933;
  assign n39935 = ~n39932 & n39934;
  assign n39936 = pi212 & ~n39935;
  assign n39937 = ~n39928 & n39936;
  assign n39938 = n39931 & ~n39937;
  assign n39939 = ~n39919 & ~n39938;
  assign n39940 = ~n39721 & ~n39939;
  assign n39941 = ~pi1147 & n39940;
  assign n39942 = pi299 & ~n38290;
  assign n39943 = ~po1038 & ~n38292;
  assign n39944 = n39942 & n39943;
  assign n39945 = ~po1038 & n39614;
  assign n39946 = ~n39944 & ~n39945;
  assign n39947 = ~n38290 & n38293;
  assign n39948 = n39946 & ~n39947;
  assign n39949 = pi1147 & n39948;
  assign n39950 = pi1149 & ~n39949;
  assign n39951 = ~n39941 & n39950;
  assign n39952 = pi211 & n38298;
  assign n39953 = pi212 & n38592;
  assign n39954 = ~n39952 & ~n39953;
  assign n39955 = n39240 & ~n39954;
  assign n39956 = pi299 & n10654;
  assign n39957 = ~n39577 & ~n39956;
  assign n39958 = ~pi212 & ~n39957;
  assign n39959 = ~pi219 & ~n39958;
  assign n39960 = ~pi299 & ~n39576;
  assign n39961 = pi214 & ~n39960;
  assign n39962 = ~pi214 & n39577;
  assign n39963 = ~pi212 & ~n39962;
  assign n39964 = ~n39961 & n39963;
  assign n39965 = ~pi211 & ~n39960;
  assign n39966 = ~n39577 & ~n39965;
  assign n39967 = pi214 & ~n39966;
  assign n39968 = pi212 & ~n39967;
  assign n39969 = ~pi214 & ~n39960;
  assign n39970 = n39968 & ~n39969;
  assign n39971 = ~n39964 & ~n39970;
  assign n39972 = ~n13025 & ~n39577;
  assign n39973 = ~n39961 & n39972;
  assign n39974 = pi212 & ~n39973;
  assign n39975 = n39971 & n39974;
  assign n39976 = n39959 & ~n39975;
  assign n39977 = pi219 & ~n39577;
  assign n39978 = ~po1038 & ~n39977;
  assign n39979 = ~n39976 & n39978;
  assign n39980 = ~n39955 & ~n39979;
  assign n39981 = ~pi1147 & n39980;
  assign n39982 = pi212 & ~n38503;
  assign n39983 = ~pi219 & ~n39952;
  assign n39984 = ~n39982 & n39983;
  assign n39985 = n39944 & ~n39984;
  assign n39986 = ~po1038 & n39615;
  assign n39987 = n38293 & ~n39984;
  assign n39988 = ~n39986 & ~n39987;
  assign n39989 = ~n39985 & n39988;
  assign n39990 = pi1147 & n39989;
  assign n39991 = ~pi1149 & ~n39990;
  assign n39992 = ~n39981 & n39991;
  assign n39993 = ~n39951 & ~n39992;
  assign n39994 = pi1148 & ~n39993;
  assign n39995 = n10656 & ~n39683;
  assign n39996 = n38293 & ~n39995;
  assign n39997 = ~pi211 & ~n39505;
  assign n39998 = pi211 & ~n39529;
  assign n39999 = pi214 & ~n39998;
  assign n40000 = ~n39997 & n39999;
  assign n40001 = n10708 & ~n40000;
  assign n40002 = ~pi214 & n39505;
  assign n40003 = ~pi212 & ~n40002;
  assign n40004 = pi214 & n39542;
  assign n40005 = n40003 & ~n40004;
  assign n40006 = ~pi219 & ~n40005;
  assign n40007 = pi212 & ~n40000;
  assign n40008 = ~n39542 & n40007;
  assign n40009 = n40006 & ~n40008;
  assign n40010 = ~n40001 & n40009;
  assign n40011 = pi212 & ~n39542;
  assign n40012 = pi219 & ~n40011;
  assign n40013 = ~n40005 & n40012;
  assign n40014 = ~po1038 & ~n40013;
  assign n40015 = ~n40010 & n40014;
  assign n40016 = ~n39996 & ~n40015;
  assign n40017 = pi1147 & n40016;
  assign n40018 = n16429 & n39553;
  assign n40019 = ~pi219 & ~n16429;
  assign n40020 = n39683 & n40019;
  assign n40021 = ~n40018 & ~n40020;
  assign n40022 = ~pi1147 & n40021;
  assign n40023 = pi1149 & ~n40022;
  assign n40024 = ~n40017 & n40023;
  assign n40025 = ~pi212 & ~n39956;
  assign n40026 = ~n39615 & n40025;
  assign n40027 = ~n39615 & ~n39762;
  assign n40028 = ~n39619 & ~n40027;
  assign n40029 = n39772 & ~n40028;
  assign n40030 = ~n40026 & ~n40029;
  assign n40031 = ~pi219 & ~n40030;
  assign n40032 = n38484 & ~n39922;
  assign n40033 = pi208 & ~n40032;
  assign n40034 = ~pi199 & ~n40033;
  assign n40035 = n39615 & ~n40034;
  assign n40036 = ~pi299 & ~n40035;
  assign n40037 = ~pi219 & n40036;
  assign n40038 = ~n40031 & ~n40037;
  assign n40039 = ~pi211 & ~n40038;
  assign n40040 = ~n13025 & n39795;
  assign n40041 = ~pi214 & n40027;
  assign n40042 = pi212 & ~n40041;
  assign n40043 = ~n40040 & n40042;
  assign n40044 = ~pi212 & n40028;
  assign n40045 = ~pi219 & ~n40044;
  assign n40046 = ~n40043 & n40045;
  assign n40047 = pi219 & ~n39762;
  assign n40048 = n39943 & ~n40047;
  assign n40049 = ~n39986 & ~n40048;
  assign n40050 = ~n40046 & ~n40049;
  assign n40051 = ~n40036 & n40050;
  assign n40052 = ~n40039 & n40051;
  assign n40053 = ~n39740 & ~n40052;
  assign n40054 = pi1147 & ~pi1149;
  assign n40055 = ~n40053 & n40054;
  assign n40056 = ~n40024 & ~n40055;
  assign n40057 = ~pi1148 & ~n40056;
  assign n40058 = ~n39994 & ~n40057;
  assign n40059 = pi213 & ~n40058;
  assign n40060 = ~po1038 & n39577;
  assign n40061 = ~pi211 & pi1146;
  assign n40062 = pi211 & pi1145;
  assign n40063 = ~n40061 & ~n40062;
  assign n40064 = pi214 & ~n40063;
  assign n40065 = pi211 & pi1146;
  assign n40066 = ~pi214 & n40065;
  assign n40067 = ~n40064 & ~n40066;
  assign n40068 = pi212 & ~n40067;
  assign n40069 = n38298 & n40065;
  assign n40070 = ~n40068 & ~n40069;
  assign n40071 = ~n38839 & n40070;
  assign n40072 = po1038 & n39277;
  assign n40073 = ~n39240 & ~n40072;
  assign n40074 = ~n40071 & ~n40073;
  assign n40075 = ~pi1147 & ~n40074;
  assign n40076 = ~pi211 & n39428;
  assign n40077 = pi219 & ~n40076;
  assign n40078 = n39943 & ~n40077;
  assign n40079 = pi219 & n40078;
  assign n40080 = pi299 & ~n40070;
  assign n40081 = n35998 & n40080;
  assign n40082 = ~n40079 & ~n40081;
  assign n40083 = n40075 & n40082;
  assign n40084 = ~n40060 & n40083;
  assign n40085 = n10711 & n38669;
  assign n40086 = po1038 & n40085;
  assign n40087 = pi1147 & ~n40086;
  assign n40088 = ~n40074 & n40087;
  assign n40089 = ~n39986 & ~n40078;
  assign n40090 = pi299 & pi1146;
  assign n40091 = pi211 & n40090;
  assign n40092 = ~n39762 & ~n40091;
  assign n40093 = ~n39615 & n40092;
  assign n40094 = n38664 & ~n40093;
  assign n40095 = n38290 & n39615;
  assign n40096 = ~pi219 & ~n40095;
  assign n40097 = pi299 & ~n40063;
  assign n40098 = ~n39615 & ~n40097;
  assign n40099 = n10708 & ~n40098;
  assign n40100 = ~n40094 & n40096;
  assign n40101 = ~n40099 & n40100;
  assign n40102 = ~n40089 & ~n40101;
  assign n40103 = n40088 & ~n40102;
  assign n40104 = pi1148 & ~n40103;
  assign n40105 = ~n40084 & n40104;
  assign n40106 = ~pi1146 & n13025;
  assign n40107 = n38664 & ~n40106;
  assign n40108 = ~n40099 & ~n40107;
  assign n40109 = ~pi219 & ~n40036;
  assign n40110 = ~n40108 & n40109;
  assign n40111 = n39277 & n39288;
  assign n40112 = ~n38669 & n40035;
  assign n40113 = ~n40111 & ~n40112;
  assign n40114 = ~n40110 & n40113;
  assign n40115 = ~po1038 & ~n40114;
  assign n40116 = n40088 & ~n40115;
  assign n40117 = ~pi1148 & ~n40083;
  assign n40118 = ~n40116 & n40117;
  assign n40119 = ~n40105 & ~n40118;
  assign n40120 = ~pi1149 & ~n40119;
  assign n40121 = pi219 & n39505;
  assign n40122 = ~po1038 & ~n40121;
  assign n40123 = ~n40078 & ~n40122;
  assign n40124 = ~n39541 & ~n40091;
  assign n40125 = ~n39540 & n40124;
  assign n40126 = pi214 & n40125;
  assign n40127 = n40003 & ~n40126;
  assign n40128 = ~pi214 & n40125;
  assign n40129 = pi214 & ~n40097;
  assign n40130 = n39505 & n40129;
  assign n40131 = pi212 & ~n40130;
  assign n40132 = ~n40128 & n40131;
  assign n40133 = ~pi219 & ~n40127;
  assign n40134 = ~n40132 & n40133;
  assign n40135 = ~n40123 & ~n40134;
  assign n40136 = n40088 & ~n40135;
  assign n40137 = ~n40018 & n40083;
  assign n40138 = ~pi1148 & ~n40137;
  assign n40139 = ~n40136 & n40138;
  assign n40140 = ~n38290 & n39932;
  assign n40141 = ~n38291 & n39596;
  assign n40142 = pi219 & ~n40141;
  assign n40143 = ~n40140 & n40142;
  assign n40144 = ~po1038 & ~n40143;
  assign n40145 = n11348 & n40144;
  assign n40146 = ~n40078 & ~n40145;
  assign n40147 = ~n39596 & ~n40091;
  assign n40148 = n39921 & ~n40147;
  assign n40149 = pi212 & ~n39928;
  assign n40150 = ~n39596 & n40067;
  assign n40151 = n40149 & ~n40150;
  assign n40152 = ~pi219 & ~n40148;
  assign n40153 = ~n40151 & n40152;
  assign n40154 = ~n40146 & ~n40153;
  assign n40155 = n40075 & ~n40154;
  assign n40156 = pi219 & ~n39614;
  assign n40157 = ~po1038 & ~n40156;
  assign n40158 = pi211 & ~n39614;
  assign n40159 = pi214 & pi299;
  assign n40160 = ~n39614 & ~n40159;
  assign n40161 = ~pi212 & ~n40160;
  assign n40162 = ~n40158 & n40161;
  assign n40163 = ~pi299 & ~n39614;
  assign n40164 = pi212 & ~n40163;
  assign n40165 = pi299 & n39982;
  assign n40166 = n40164 & ~n40165;
  assign n40167 = ~pi219 & ~n40162;
  assign n40168 = ~n40166 & n40167;
  assign n40169 = n40157 & ~n40168;
  assign n40170 = n40082 & n40088;
  assign n40171 = ~n40169 & n40170;
  assign n40172 = pi1148 & ~n40171;
  assign n40173 = ~n40155 & n40172;
  assign n40174 = ~n40139 & ~n40173;
  assign n40175 = pi1149 & ~n40174;
  assign n40176 = ~n40120 & ~n40175;
  assign n40177 = ~pi213 & ~n40176;
  assign n40178 = pi209 & ~n40177;
  assign n40179 = ~n40059 & n40178;
  assign n40180 = ~pi199 & pi1146;
  assign n40181 = pi200 & ~n40180;
  assign n40182 = ~pi299 & ~n40181;
  assign n40183 = pi199 & pi1145;
  assign n40184 = n38483 & ~n40183;
  assign n40185 = n40182 & ~n40184;
  assign n40186 = ~pi207 & n40185;
  assign n40187 = ~pi200 & ~n40183;
  assign n40188 = ~n40180 & n40187;
  assign n40189 = pi200 & ~n39258;
  assign n40190 = n38319 & ~n40189;
  assign n40191 = ~n40188 & n40190;
  assign n40192 = ~n40090 & ~n40191;
  assign n40193 = ~n40186 & n40192;
  assign n40194 = pi208 & ~n40193;
  assign n40195 = n38326 & n40185;
  assign n40196 = ~n40194 & ~n40195;
  assign n40197 = ~pi299 & n40196;
  assign n40198 = pi211 & ~n40197;
  assign n40199 = n40186 & n40187;
  assign n40200 = n40194 & ~n40199;
  assign n40201 = n40182 & ~n40187;
  assign n40202 = n38326 & n40201;
  assign n40203 = ~n40200 & ~n40202;
  assign n40204 = ~pi299 & n40203;
  assign n40205 = pi214 & ~n40204;
  assign n40206 = ~n40198 & ~n40205;
  assign n40207 = pi212 & ~n40206;
  assign n40208 = n10654 & ~n40197;
  assign n40209 = ~n38708 & ~n40191;
  assign n40210 = ~n10463 & ~n40185;
  assign n40211 = ~n40209 & ~n40210;
  assign n40212 = ~pi219 & ~n40211;
  assign n40213 = ~n40208 & n40212;
  assign n40214 = ~n40207 & n40213;
  assign n40215 = ~n10463 & ~n40201;
  assign n40216 = ~n40209 & ~n40215;
  assign n40217 = n38290 & n40216;
  assign n40218 = n40214 & ~n40217;
  assign n40219 = ~pi211 & ~n40197;
  assign n40220 = ~n40211 & ~n40219;
  assign n40221 = pi214 & n40220;
  assign n40222 = ~n40204 & ~n40221;
  assign n40223 = pi212 & ~n40222;
  assign n40224 = ~pi214 & n40216;
  assign n40225 = ~pi212 & ~n40224;
  assign n40226 = ~n40205 & n40225;
  assign n40227 = ~n40223 & ~n40226;
  assign n40228 = ~pi219 & ~n40227;
  assign n40229 = pi219 & ~n40216;
  assign n40230 = ~po1038 & ~n40229;
  assign n40231 = ~n40228 & n40230;
  assign n40232 = ~n40218 & n40231;
  assign n40233 = ~pi1147 & ~n39955;
  assign n40234 = ~n40232 & n40233;
  assign n40235 = ~n38291 & n40211;
  assign n40236 = pi219 & ~n40235;
  assign n40237 = ~n38290 & n40219;
  assign n40238 = n40236 & ~n40237;
  assign n40239 = ~po1038 & ~n40238;
  assign n40240 = ~n40214 & n40239;
  assign n40241 = pi1147 & ~n39987;
  assign n40242 = ~n40240 & n40241;
  assign n40243 = ~pi1149 & ~n40242;
  assign n40244 = ~n40234 & n40243;
  assign n40245 = ~pi1147 & ~n39721;
  assign n40246 = ~n40231 & n40245;
  assign n40247 = ~n39942 & n40212;
  assign n40248 = n40239 & ~n40247;
  assign n40249 = pi1147 & ~n39947;
  assign n40250 = ~n40248 & n40249;
  assign n40251 = pi1149 & ~n40250;
  assign n40252 = ~n40246 & n40251;
  assign n40253 = pi1148 & ~n40252;
  assign n40254 = ~n40244 & n40253;
  assign n40255 = ~pi1147 & ~po1038;
  assign n40256 = n40216 & n40255;
  assign n40257 = pi214 & ~n40211;
  assign n40258 = ~n40198 & n40257;
  assign n40259 = ~pi214 & ~n40211;
  assign n40260 = ~n40219 & n40259;
  assign n40261 = pi212 & ~n40258;
  assign n40262 = ~n40260 & n40261;
  assign n40263 = ~pi212 & ~n40259;
  assign n40264 = ~n40220 & n40263;
  assign n40265 = ~pi219 & ~n40264;
  assign n40266 = ~n40262 & n40265;
  assign n40267 = n40240 & ~n40266;
  assign n40268 = ~n39740 & ~n40267;
  assign n40269 = pi1147 & ~n40268;
  assign n40270 = ~n40256 & ~n40269;
  assign n40271 = ~pi1149 & ~n40270;
  assign n40272 = n40239 & ~n40266;
  assign n40273 = ~n39996 & ~n40272;
  assign n40274 = pi1147 & ~n40273;
  assign n40275 = ~pi1147 & n40085;
  assign n40276 = ~n40256 & ~n40275;
  assign n40277 = n16429 & n40085;
  assign n40278 = n40203 & n40277;
  assign n40279 = ~n40276 & ~n40278;
  assign n40280 = ~n40274 & ~n40279;
  assign n40281 = pi1149 & ~n40280;
  assign n40282 = ~pi1148 & ~n40281;
  assign n40283 = ~n40271 & n40282;
  assign n40284 = pi213 & ~n40254;
  assign n40285 = ~n40283 & n40284;
  assign n40286 = pi219 & ~n40217;
  assign n40287 = ~n38290 & n40216;
  assign n40288 = ~n38291 & ~n40287;
  assign n40289 = ~pi299 & ~n40203;
  assign n40290 = ~pi211 & ~n39428;
  assign n40291 = ~n40289 & n40290;
  assign n40292 = ~n40288 & ~n40291;
  assign n40293 = n40286 & ~n40292;
  assign n40294 = ~n40091 & ~n40216;
  assign n40295 = ~pi214 & ~n40216;
  assign n40296 = ~pi212 & ~n40295;
  assign n40297 = ~n40294 & n40296;
  assign n40298 = ~pi219 & ~n40297;
  assign n40299 = n40129 & ~n40289;
  assign n40300 = ~pi214 & n40294;
  assign n40301 = pi212 & ~n40300;
  assign n40302 = ~n40299 & n40301;
  assign n40303 = n40298 & ~n40302;
  assign n40304 = ~po1038 & ~n40293;
  assign n40305 = ~n40303 & n40304;
  assign n40306 = n40075 & ~n40305;
  assign n40307 = ~n39425 & n40198;
  assign n40308 = n40129 & n40196;
  assign n40309 = ~n40208 & ~n40308;
  assign n40310 = ~n40307 & ~n40309;
  assign n40311 = ~pi214 & n40092;
  assign n40312 = n40196 & n40311;
  assign n40313 = pi212 & ~n40312;
  assign n40314 = ~n40310 & n40313;
  assign n40315 = ~n40264 & n40298;
  assign n40316 = ~n40314 & n40315;
  assign n40317 = ~n39425 & n40219;
  assign n40318 = ~n38290 & n40317;
  assign n40319 = n40236 & ~n40318;
  assign n40320 = ~po1038 & ~n40319;
  assign n40321 = ~n40316 & n40320;
  assign n40322 = n40088 & ~n40321;
  assign n40323 = ~n40306 & ~n40322;
  assign n40324 = ~pi213 & n40323;
  assign n40325 = ~pi209 & ~n40324;
  assign n40326 = ~n40285 & n40325;
  assign n40327 = ~n40179 & ~n40326;
  assign n40328 = pi230 & ~n40327;
  assign n40329 = ~pi230 & ~pi240;
  assign po397 = ~n40328 & ~n40329;
  assign n40331 = po1038 & ~n40085;
  assign n40332 = pi1151 & ~n40331;
  assign n40333 = ~n39607 & n40085;
  assign n40334 = n39786 & ~n40333;
  assign n40335 = pi1152 & ~n40334;
  assign n40336 = ~po1038 & ~n40335;
  assign n40337 = n40332 & ~n40336;
  assign n40338 = n39550 & n39562;
  assign n40339 = n38384 & n39683;
  assign n40340 = ~n39506 & ~n40339;
  assign n40341 = n40332 & ~n40340;
  assign n40342 = ~n40338 & ~n40341;
  assign n40343 = ~pi1152 & ~n40342;
  assign n40344 = pi1152 & n39562;
  assign n40345 = n39597 & n40344;
  assign n40346 = ~n40343 & ~n40345;
  assign n40347 = ~n40337 & n40346;
  assign n40348 = ~pi1150 & ~n40347;
  assign n40349 = pi1151 & ~n39721;
  assign n40350 = pi219 & ~n39550;
  assign n40351 = ~po1038 & ~n40350;
  assign n40352 = ~n39986 & ~n40351;
  assign n40353 = n39621 & ~n39799;
  assign n40354 = ~pi219 & ~n40353;
  assign n40355 = ~pi214 & n39607;
  assign n40356 = pi212 & ~n40355;
  assign n40357 = ~n39788 & n40356;
  assign n40358 = n40354 & ~n40357;
  assign n40359 = pi1152 & ~n40358;
  assign n40360 = ~pi299 & ~n39530;
  assign n40361 = ~pi214 & n39529;
  assign n40362 = pi212 & ~n40361;
  assign n40363 = ~n40004 & n40362;
  assign n40364 = ~n39508 & ~n40363;
  assign n40365 = ~n40360 & ~n40364;
  assign n40366 = ~pi219 & ~n40365;
  assign n40367 = ~pi1152 & ~n40121;
  assign n40368 = ~n40366 & n40367;
  assign n40369 = ~n40359 & ~n40368;
  assign n40370 = ~n40352 & ~n40369;
  assign n40371 = n40349 & ~n40370;
  assign n40372 = ~pi1151 & ~n39955;
  assign n40373 = ~pi212 & ~n39554;
  assign n40374 = ~n39564 & n40373;
  assign n40375 = ~n39762 & n40374;
  assign n40376 = ~pi219 & ~n40375;
  assign n40377 = pi214 & ~n39563;
  assign n40378 = ~pi211 & n39564;
  assign n40379 = pi212 & ~n39554;
  assign n40380 = ~n40378 & n40379;
  assign n40381 = ~n40377 & n40380;
  assign n40382 = n40376 & ~n40381;
  assign n40383 = ~n39550 & n39774;
  assign n40384 = ~pi299 & n40383;
  assign n40385 = ~n40382 & ~n40384;
  assign n40386 = n40351 & n40385;
  assign n40387 = ~pi1152 & ~n40386;
  assign n40388 = ~n39597 & ~n40385;
  assign n40389 = n39807 & ~n40388;
  assign n40390 = pi1152 & ~n40389;
  assign n40391 = ~n40387 & ~n40390;
  assign n40392 = n40372 & ~n40391;
  assign n40393 = pi1150 & ~n40392;
  assign n40394 = ~n40371 & n40393;
  assign n40395 = ~n40348 & ~n40394;
  assign n40396 = ~pi1149 & ~n40395;
  assign n40397 = ~n38592 & ~n39607;
  assign n40398 = pi212 & n39786;
  assign n40399 = ~n40397 & n40398;
  assign n40400 = ~n39790 & ~n40399;
  assign n40401 = ~pi219 & ~n40400;
  assign n40402 = pi1152 & ~n40401;
  assign n40403 = n39793 & n40402;
  assign n40404 = pi1151 & ~n39996;
  assign n40405 = ~pi214 & ~n39764;
  assign n40406 = n39757 & ~n40405;
  assign n40407 = ~pi212 & ~n39765;
  assign n40408 = ~n40406 & ~n40407;
  assign n40409 = ~pi219 & ~n40408;
  assign n40410 = ~pi1152 & n39767;
  assign n40411 = ~n40409 & n40410;
  assign n40412 = n40404 & ~n40411;
  assign n40413 = ~n40403 & n40412;
  assign n40414 = ~n40048 & ~n40351;
  assign n40415 = ~n40383 & ~n40414;
  assign n40416 = ~pi1152 & n40415;
  assign n40417 = ~n39807 & n40414;
  assign n40418 = ~n39597 & n39774;
  assign n40419 = pi1152 & ~n40417;
  assign n40420 = ~n40418 & n40419;
  assign n40421 = ~pi1151 & ~n39740;
  assign n40422 = ~n40416 & n40421;
  assign n40423 = ~n40420 & n40422;
  assign n40424 = ~pi1150 & ~n40423;
  assign n40425 = ~n40413 & n40424;
  assign n40426 = pi212 & ~n39607;
  assign n40427 = n40354 & ~n40426;
  assign n40428 = pi1152 & ~n40427;
  assign n40429 = n39793 & n40428;
  assign n40430 = pi1151 & ~n39947;
  assign n40431 = ~n39544 & ~n40360;
  assign n40432 = ~pi219 & ~n40431;
  assign n40433 = n40410 & ~n40432;
  assign n40434 = n40430 & ~n40433;
  assign n40435 = ~n40429 & n40434;
  assign n40436 = ~pi1151 & ~n39987;
  assign n40437 = n10708 & n39584;
  assign n40438 = ~n39565 & ~n39754;
  assign n40439 = ~n10708 & ~n39597;
  assign n40440 = ~n40438 & n40439;
  assign n40441 = ~n40437 & ~n40440;
  assign n40442 = ~pi219 & ~n40441;
  assign n40443 = ~n40417 & ~n40442;
  assign n40444 = pi1152 & ~n40443;
  assign n40445 = n40387 & ~n40415;
  assign n40446 = ~n40444 & ~n40445;
  assign n40447 = n40436 & ~n40446;
  assign n40448 = pi1150 & ~n40447;
  assign n40449 = ~n40435 & n40448;
  assign n40450 = ~n40425 & ~n40449;
  assign n40451 = pi1149 & ~n40450;
  assign n40452 = ~n40396 & ~n40451;
  assign n40453 = ~pi213 & ~n40452;
  assign n40454 = pi213 & ~n39819;
  assign n40455 = pi209 & ~n40454;
  assign n40456 = ~n40453 & n40455;
  assign n40457 = ~n39979 & n40372;
  assign n40458 = ~n39939 & n40349;
  assign n40459 = pi1150 & ~n40458;
  assign n40460 = ~n40457 & n40459;
  assign n40461 = ~pi1150 & pi1151;
  assign n40462 = ~n40021 & n40461;
  assign n40463 = ~pi1149 & ~n40462;
  assign n40464 = ~n40460 & n40463;
  assign n40465 = ~n40015 & n40404;
  assign n40466 = ~n40052 & n40421;
  assign n40467 = ~pi1150 & ~n40466;
  assign n40468 = ~n40465 & n40467;
  assign n40469 = ~pi1151 & n39989;
  assign n40470 = n39946 & n40430;
  assign n40471 = pi1150 & ~n40470;
  assign n40472 = ~n40469 & n40471;
  assign n40473 = pi1149 & ~n40472;
  assign n40474 = ~n40468 & n40473;
  assign n40475 = ~n40464 & ~n40474;
  assign n40476 = ~pi213 & n40475;
  assign n40477 = ~n40003 & ~n40007;
  assign n40478 = ~n38544 & n39540;
  assign n40479 = ~n39541 & ~n40478;
  assign n40480 = ~n40001 & n40479;
  assign n40481 = ~n40477 & ~n40480;
  assign n40482 = ~pi219 & ~n40481;
  assign n40483 = n40014 & ~n40482;
  assign n40484 = n39687 & ~n40483;
  assign n40485 = pi299 & n39498;
  assign n40486 = ~n40035 & ~n40339;
  assign n40487 = ~po1038 & ~n40486;
  assign n40488 = ~n40485 & n40487;
  assign n40489 = n39711 & ~n40488;
  assign n40490 = ~pi1152 & ~n40489;
  assign n40491 = ~n40484 & n40490;
  assign n40492 = ~n40000 & ~n40002;
  assign n40493 = ~pi219 & ~n40165;
  assign n40494 = ~n39545 & n40493;
  assign n40495 = ~n40492 & n40494;
  assign n40496 = n40014 & ~n40495;
  assign n40497 = n39742 & ~n40496;
  assign n40498 = ~n39942 & ~n40035;
  assign n40499 = ~n38410 & n39723;
  assign n40500 = ~n40498 & ~n40499;
  assign n40501 = ~pi219 & ~n40500;
  assign n40502 = pi219 & ~n40035;
  assign n40503 = ~po1038 & ~n40502;
  assign n40504 = ~n40501 & n40503;
  assign n40505 = n39725 & ~n40504;
  assign n40506 = pi1152 & ~n40505;
  assign n40507 = ~n40497 & n40506;
  assign n40508 = ~pi1150 & ~n40507;
  assign n40509 = ~n40491 & n40508;
  assign n40510 = ~pi219 & ~n39614;
  assign n40511 = ~n40165 & n40510;
  assign n40512 = ~pi1153 & n40511;
  assign n40513 = pi299 & n10655;
  assign n40514 = ~pi219 & ~n40513;
  assign n40515 = n40048 & ~n40514;
  assign n40516 = ~n40169 & ~n40515;
  assign n40517 = ~n40512 & ~n40516;
  assign n40518 = n39687 & ~n40517;
  assign n40519 = pi1153 & n40339;
  assign n40520 = n39711 & ~n40519;
  assign n40521 = ~pi1152 & ~n40520;
  assign n40522 = ~pi1151 & ~n39986;
  assign n40523 = ~pi1152 & ~n40522;
  assign n40524 = ~n40521 & ~n40523;
  assign n40525 = ~n40518 & ~n40524;
  assign n40526 = ~pi211 & n40511;
  assign n40527 = ~n39946 & ~n40526;
  assign n40528 = n39742 & ~n40527;
  assign n40529 = ~n40517 & n40528;
  assign n40530 = ~po1038 & ~n39626;
  assign n40531 = n10708 & ~n40027;
  assign n40532 = ~pi299 & ~n39615;
  assign n40533 = ~n38300 & ~n40485;
  assign n40534 = ~n40532 & n40533;
  assign n40535 = n40096 & ~n40531;
  assign n40536 = ~n40534 & n40535;
  assign n40537 = n40530 & ~n40536;
  assign n40538 = n39725 & ~n40537;
  assign n40539 = pi1152 & ~n40538;
  assign n40540 = ~n40529 & n40539;
  assign n40541 = pi1150 & ~n40525;
  assign n40542 = ~n40540 & n40541;
  assign n40543 = pi1149 & ~n40542;
  assign n40544 = ~n40509 & n40543;
  assign n40545 = ~n39960 & ~n40485;
  assign n40546 = pi214 & n40545;
  assign n40547 = n39963 & ~n40546;
  assign n40548 = ~pi214 & n40545;
  assign n40549 = n39968 & ~n40548;
  assign n40550 = ~n40547 & ~n40549;
  assign n40551 = ~pi219 & ~n40550;
  assign n40552 = n39978 & ~n40551;
  assign n40553 = n39725 & ~n40552;
  assign n40554 = pi211 & ~n39928;
  assign n40555 = ~n11358 & n38522;
  assign n40556 = ~n39925 & ~n40555;
  assign n40557 = ~pi211 & ~n38544;
  assign n40558 = ~n40556 & n40557;
  assign n40559 = ~n40554 & ~n40558;
  assign n40560 = pi214 & n40559;
  assign n40561 = n39921 & ~n40560;
  assign n40562 = ~pi214 & n40559;
  assign n40563 = n40149 & ~n40562;
  assign n40564 = ~pi219 & ~n40561;
  assign n40565 = ~n40563 & n40564;
  assign n40566 = n40144 & ~n40565;
  assign n40567 = n39742 & ~n40566;
  assign n40568 = pi1152 & ~n40567;
  assign n40569 = ~n40553 & n40568;
  assign n40570 = n39577 & ~n39712;
  assign n40571 = ~n38544 & ~n39960;
  assign n40572 = ~pi211 & ~n40571;
  assign n40573 = n39712 & ~n39966;
  assign n40574 = ~n40572 & n40573;
  assign n40575 = ~n40570 & ~n40574;
  assign n40576 = ~po1038 & ~n40575;
  assign n40577 = n39711 & ~n40576;
  assign n40578 = ~n39596 & ~n40554;
  assign n40579 = pi214 & n40578;
  assign n40580 = n39920 & ~n39932;
  assign n40581 = pi212 & ~n40580;
  assign n40582 = ~n40579 & n40581;
  assign n40583 = ~n40559 & n40582;
  assign n40584 = ~n39933 & ~n40558;
  assign n40585 = n39921 & ~n40584;
  assign n40586 = ~pi219 & ~n40585;
  assign n40587 = ~n40583 & n40586;
  assign n40588 = n40144 & ~n40587;
  assign n40589 = n39687 & ~n40588;
  assign n40590 = ~pi1152 & ~n40577;
  assign n40591 = ~n40589 & n40590;
  assign n40592 = pi1150 & ~n40591;
  assign n40593 = ~n40569 & n40592;
  assign n40594 = pi219 & ~n39566;
  assign n40595 = ~po1038 & ~n40594;
  assign n40596 = ~n39778 & n40595;
  assign n40597 = n40376 & ~n40380;
  assign n40598 = n40595 & ~n40597;
  assign n40599 = n39742 & ~n40596;
  assign n40600 = ~n40598 & n40599;
  assign n40601 = pi299 & n39720;
  assign n40602 = ~n39723 & n40601;
  assign n40603 = n39725 & ~n40602;
  assign n40604 = pi1152 & ~n40603;
  assign n40605 = ~n40600 & n40604;
  assign n40606 = n39687 & ~n40596;
  assign n40607 = n40521 & ~n40606;
  assign n40608 = ~pi1150 & ~n40607;
  assign n40609 = ~n40605 & n40608;
  assign n40610 = ~pi1149 & ~n40609;
  assign n40611 = ~n40593 & n40610;
  assign n40612 = ~n40544 & ~n40611;
  assign n40613 = pi213 & ~n40612;
  assign n40614 = ~pi209 & ~n40476;
  assign n40615 = ~n40613 & n40614;
  assign n40616 = ~n40456 & ~n40615;
  assign n40617 = pi230 & ~n40616;
  assign n40618 = ~pi230 & ~pi241;
  assign po398 = ~n40617 & ~n40618;
  assign n40620 = ~pi230 & ~pi242;
  assign n40621 = pi214 & ~n39279;
  assign n40622 = ~pi214 & ~n40063;
  assign n40623 = ~n40621 & ~n40622;
  assign n40624 = pi212 & ~n40623;
  assign n40625 = ~pi212 & n40064;
  assign n40626 = ~pi219 & ~n40625;
  assign n40627 = ~n40624 & n40626;
  assign n40628 = pi219 & ~n38296;
  assign n40629 = n38293 & ~n40628;
  assign n40630 = ~n40627 & n40629;
  assign n40631 = pi199 & pi1144;
  assign n40632 = ~pi200 & ~n40631;
  assign n40633 = ~n40180 & n40632;
  assign n40634 = ~pi299 & ~n40189;
  assign n40635 = ~n40633 & n40634;
  assign n40636 = ~pi207 & ~n40635;
  assign n40637 = ~pi299 & ~n39260;
  assign n40638 = ~n39258 & n40632;
  assign n40639 = n40637 & ~n40638;
  assign n40640 = pi207 & ~n40639;
  assign n40641 = pi208 & ~n40636;
  assign n40642 = ~n40640 & n40641;
  assign n40643 = n38708 & n40635;
  assign n40644 = ~n40642 & ~n40643;
  assign n40645 = ~n39428 & n40644;
  assign n40646 = ~pi211 & ~n40645;
  assign n40647 = ~n38637 & n40644;
  assign n40648 = pi211 & ~n40647;
  assign n40649 = pi214 & ~n40646;
  assign n40650 = ~n40648 & n40649;
  assign n40651 = ~n40090 & n40644;
  assign n40652 = ~pi211 & ~n40651;
  assign n40653 = pi211 & ~n40645;
  assign n40654 = ~n40652 & ~n40653;
  assign n40655 = ~pi214 & n40654;
  assign n40656 = pi212 & ~n40650;
  assign n40657 = ~n40655 & n40656;
  assign n40658 = ~pi214 & n40644;
  assign n40659 = ~pi212 & ~n40658;
  assign n40660 = ~n40654 & n40659;
  assign n40661 = ~pi219 & ~n40660;
  assign n40662 = ~n40657 & n40661;
  assign n40663 = ~n38291 & ~n40644;
  assign n40664 = pi219 & ~n40663;
  assign n40665 = n38291 & ~n40647;
  assign n40666 = n40664 & ~n40665;
  assign n40667 = ~po1038 & ~n40666;
  assign n40668 = ~n40662 & n40667;
  assign n40669 = ~n40630 & ~n40668;
  assign n40670 = pi213 & n40669;
  assign n40671 = pi211 & ~n40643;
  assign n40672 = n38326 & n40635;
  assign n40673 = n38291 & ~n38673;
  assign n40674 = ~n40672 & n40673;
  assign n40675 = ~n40671 & ~n40674;
  assign n40676 = pi219 & ~n40675;
  assign n40677 = n38290 & ~n40643;
  assign n40678 = n10708 & ~n38334;
  assign n40679 = ~n38308 & n38664;
  assign n40680 = ~n40678 & ~n40679;
  assign n40681 = ~pi219 & ~n40672;
  assign n40682 = ~n40680 & n40681;
  assign n40683 = ~n40677 & ~n40682;
  assign n40684 = ~n40676 & n40683;
  assign n40685 = ~n40642 & ~n40684;
  assign n40686 = ~po1038 & ~n40685;
  assign n40687 = ~pi213 & ~n38307;
  assign n40688 = ~n40686 & n40687;
  assign n40689 = ~n40670 & ~n40688;
  assign n40690 = pi209 & ~n40689;
  assign n40691 = ~pi213 & ~n38353;
  assign n40692 = ~n38292 & ~n40628;
  assign n40693 = ~n40627 & n40692;
  assign n40694 = pi299 & ~n40693;
  assign n40695 = ~po1038 & ~n40694;
  assign n40696 = ~n38345 & n40695;
  assign n40697 = ~n40630 & ~n40696;
  assign n40698 = pi213 & ~n40697;
  assign n40699 = ~pi209 & ~n40698;
  assign n40700 = ~n40691 & n40699;
  assign n40701 = ~n40690 & ~n40700;
  assign n40702 = pi230 & ~n40701;
  assign po399 = ~n40620 & ~n40702;
  assign n40704 = pi243 & ~pi1091;
  assign n40705 = ~pi83 & ~pi85;
  assign n40706 = pi314 & ~n40705;
  assign n40707 = pi802 & n40706;
  assign n40708 = pi276 & n40707;
  assign n40709 = ~pi1091 & ~n40708;
  assign n40710 = pi271 & ~n40709;
  assign n40711 = ~pi1091 & ~n40710;
  assign n40712 = pi273 & ~n40711;
  assign n40713 = ~pi1091 & ~n40712;
  assign n40714 = ~pi200 & ~n40713;
  assign n40715 = pi199 & ~n40713;
  assign n40716 = ~pi81 & n40705;
  assign n40717 = pi314 & ~n40716;
  assign n40718 = pi802 & n40717;
  assign n40719 = pi276 & n40718;
  assign n40720 = ~pi1091 & n40719;
  assign n40721 = pi271 & n40720;
  assign n40722 = pi273 & n40721;
  assign n40723 = ~n40712 & ~n40722;
  assign n40724 = ~pi1091 & n40723;
  assign n40725 = ~pi199 & ~n40724;
  assign n40726 = ~n40715 & ~n40725;
  assign n40727 = n40720 & ~n40726;
  assign n40728 = ~pi299 & ~n40727;
  assign n40729 = ~n40715 & n40728;
  assign n40730 = ~n40714 & n40729;
  assign n40731 = pi299 & ~n40722;
  assign n40732 = ~n40730 & ~n40731;
  assign n40733 = ~n40704 & ~n40732;
  assign n40734 = ~pi200 & ~n40720;
  assign n40735 = ~n40726 & ~n40734;
  assign n40736 = ~pi299 & ~n40735;
  assign n40737 = ~n40715 & n40736;
  assign n40738 = ~pi1091 & n40708;
  assign n40739 = pi271 & n40738;
  assign n40740 = pi273 & n40739;
  assign n40741 = pi299 & ~n40740;
  assign n40742 = ~n40714 & n40728;
  assign n40743 = ~n40725 & n40742;
  assign n40744 = ~n40741 & ~n40743;
  assign n40745 = ~n40737 & n40744;
  assign n40746 = pi299 & n40713;
  assign n40747 = ~n40742 & ~n40746;
  assign n40748 = pi243 & ~n40747;
  assign n40749 = ~n40745 & n40748;
  assign n40750 = pi1155 & ~n40749;
  assign n40751 = ~n40722 & n40746;
  assign n40752 = ~n40743 & ~n40751;
  assign n40753 = pi1155 & n40752;
  assign n40754 = ~n40750 & ~n40753;
  assign n40755 = ~n40731 & ~n40736;
  assign n40756 = ~pi243 & n40755;
  assign n40757 = ~n40730 & n40756;
  assign n40758 = ~n40754 & ~n40757;
  assign n40759 = ~n40725 & n40736;
  assign n40760 = ~n40730 & ~n40759;
  assign n40761 = ~n40751 & n40760;
  assign n40762 = ~pi243 & ~n40761;
  assign n40763 = ~n40731 & ~n40737;
  assign n40764 = pi243 & ~n40743;
  assign n40765 = n40763 & n40764;
  assign n40766 = ~n40762 & ~n40765;
  assign n40767 = ~pi1155 & ~n40766;
  assign n40768 = ~n40758 & ~n40767;
  assign n40769 = ~n40733 & n40768;
  assign n40770 = pi1156 & ~n40769;
  assign n40771 = ~n40746 & ~n40759;
  assign n40772 = ~pi243 & ~n40771;
  assign n40773 = ~pi1155 & ~n40772;
  assign n40774 = ~n40728 & ~n40731;
  assign n40775 = ~pi1155 & n40774;
  assign n40776 = ~n40773 & ~n40775;
  assign n40777 = ~n40731 & ~n40742;
  assign n40778 = pi243 & n40777;
  assign n40779 = ~n40729 & n40778;
  assign n40780 = ~n40776 & ~n40779;
  assign n40781 = ~pi1156 & ~n40780;
  assign n40782 = ~n40736 & ~n40751;
  assign n40783 = ~pi243 & ~n40782;
  assign n40784 = pi1155 & ~n40783;
  assign n40785 = ~n40778 & n40784;
  assign n40786 = n40781 & ~n40785;
  assign n40787 = pi1157 & ~n40786;
  assign n40788 = ~n40770 & n40787;
  assign n40789 = pi243 & n40774;
  assign n40790 = ~pi243 & ~pi1091;
  assign n40791 = ~n40728 & ~n40741;
  assign n40792 = n40790 & ~n40791;
  assign n40793 = ~pi1155 & ~n40792;
  assign n40794 = ~n40775 & ~n40793;
  assign n40795 = ~n40789 & ~n40794;
  assign n40796 = ~pi1156 & ~n40795;
  assign n40797 = pi1155 & ~n40704;
  assign n40798 = n40715 & n40797;
  assign n40799 = ~n40785 & ~n40798;
  assign n40800 = n40796 & n40799;
  assign n40801 = ~pi1155 & n40777;
  assign n40802 = ~n40720 & n40801;
  assign n40803 = ~n40725 & n40728;
  assign n40804 = ~n40751 & ~n40803;
  assign n40805 = pi243 & ~n40804;
  assign n40806 = ~n40729 & ~n40731;
  assign n40807 = ~pi243 & n40806;
  assign n40808 = ~n40805 & ~n40807;
  assign n40809 = pi1156 & ~n40802;
  assign n40810 = n40808 & n40809;
  assign n40811 = ~pi1157 & ~n40810;
  assign n40812 = ~n40800 & n40811;
  assign n40813 = pi211 & ~n40812;
  assign n40814 = ~n40788 & n40813;
  assign n40815 = pi1156 & ~n40768;
  assign n40816 = ~n40742 & ~n40751;
  assign n40817 = pi243 & ~n40816;
  assign n40818 = ~n40756 & ~n40817;
  assign n40819 = n40781 & n40818;
  assign n40820 = pi1157 & ~n40819;
  assign n40821 = ~n40815 & n40820;
  assign n40822 = ~pi1155 & n40816;
  assign n40823 = ~n40755 & n40822;
  assign n40824 = n40810 & ~n40823;
  assign n40825 = n40808 & n40818;
  assign n40826 = pi1155 & ~n40825;
  assign n40827 = n40796 & ~n40826;
  assign n40828 = ~pi1157 & ~n40824;
  assign n40829 = ~n40827 & n40828;
  assign n40830 = ~pi211 & ~n40829;
  assign n40831 = ~n40821 & n40830;
  assign n40832 = ~pi219 & ~n40831;
  assign n40833 = ~n40814 & n40832;
  assign n40834 = pi253 & pi254;
  assign n40835 = pi267 & n40834;
  assign n40836 = ~pi263 & n40835;
  assign n40837 = ~n40730 & ~n40746;
  assign n40838 = ~pi243 & n40837;
  assign n40839 = ~n40736 & ~n40741;
  assign n40840 = n40838 & n40839;
  assign n40841 = n40750 & ~n40840;
  assign n40842 = pi243 & ~n40745;
  assign n40843 = ~n40838 & ~n40842;
  assign n40844 = ~n40733 & ~n40772;
  assign n40845 = ~n40843 & n40844;
  assign n40846 = ~pi1155 & ~n40845;
  assign n40847 = ~n40841 & ~n40846;
  assign n40848 = pi1156 & ~n40847;
  assign n40849 = ~n40741 & ~n40759;
  assign n40850 = ~pi243 & ~n40849;
  assign n40851 = pi243 & ~n40729;
  assign n40852 = ~pi1155 & ~n40851;
  assign n40853 = ~n40850 & n40852;
  assign n40854 = ~pi243 & pi1155;
  assign n40855 = n40839 & n40854;
  assign n40856 = ~pi1156 & ~n40855;
  assign n40857 = ~n40748 & n40856;
  assign n40858 = ~n40853 & n40857;
  assign n40859 = n38365 & ~n40858;
  assign n40860 = ~n40848 & n40859;
  assign n40861 = pi243 & n40744;
  assign n40862 = n40784 & ~n40861;
  assign n40863 = ~n40773 & ~n40862;
  assign n40864 = ~n40843 & ~n40863;
  assign n40865 = pi1156 & ~n40864;
  assign n40866 = ~n40741 & ~n40742;
  assign n40867 = pi243 & n40866;
  assign n40868 = ~n40783 & ~n40867;
  assign n40869 = pi1155 & ~n40868;
  assign n40870 = ~n40729 & n40866;
  assign n40871 = pi243 & n40870;
  assign n40872 = ~n40772 & ~n40871;
  assign n40873 = ~n40869 & n40872;
  assign n40874 = ~pi1156 & ~n40873;
  assign n40875 = n39235 & ~n40874;
  assign n40876 = ~n40865 & n40875;
  assign n40877 = ~n40741 & ~n40803;
  assign n40878 = pi1155 & n40877;
  assign n40879 = ~n40736 & n40877;
  assign n40880 = ~n40878 & ~n40879;
  assign n40881 = pi243 & ~n40880;
  assign n40882 = ~n40729 & ~n40746;
  assign n40883 = ~pi243 & ~n40882;
  assign n40884 = ~n40802 & n40883;
  assign n40885 = ~n40881 & ~n40884;
  assign n40886 = pi1156 & ~n40885;
  assign n40887 = ~n40803 & n40867;
  assign n40888 = ~n40737 & ~n40746;
  assign n40889 = ~pi243 & ~n40888;
  assign n40890 = pi1155 & ~n40889;
  assign n40891 = ~n40887 & n40890;
  assign n40892 = pi243 & n40791;
  assign n40893 = n40793 & ~n40892;
  assign n40894 = ~pi1156 & ~n40893;
  assign n40895 = ~n40891 & n40894;
  assign n40896 = ~pi1157 & ~n40895;
  assign n40897 = ~n40886 & n40896;
  assign n40898 = ~n40876 & ~n40897;
  assign n40899 = ~n40860 & n40898;
  assign n40900 = pi219 & ~n40899;
  assign n40901 = n40836 & ~n40900;
  assign n40902 = ~n40833 & n40901;
  assign n40903 = ~pi299 & pi1091;
  assign n40904 = n38723 & n40903;
  assign n40905 = ~n40790 & ~n40904;
  assign n40906 = pi1156 & ~n40905;
  assign n40907 = pi1091 & ~n38824;
  assign n40908 = n39344 & n40907;
  assign n40909 = ~n40906 & ~n40908;
  assign n40910 = ~pi299 & n38483;
  assign n40911 = pi1091 & ~n40910;
  assign n40912 = ~n40704 & ~n40911;
  assign n40913 = ~n40790 & ~n40797;
  assign n40914 = n38424 & ~n40913;
  assign n40915 = ~n40912 & ~n40914;
  assign n40916 = ~pi1156 & ~n40915;
  assign n40917 = n40909 & ~n40916;
  assign n40918 = pi1157 & ~n40917;
  assign n40919 = ~n40907 & ~n40913;
  assign n40920 = ~pi1156 & ~n40919;
  assign n40921 = pi199 & pi1091;
  assign n40922 = ~pi299 & n40921;
  assign n40923 = n40797 & ~n40922;
  assign n40924 = pi1156 & ~n40923;
  assign n40925 = ~pi1155 & ~n40704;
  assign n40926 = ~n11419 & n40903;
  assign n40927 = n40925 & ~n40926;
  assign n40928 = n40924 & ~n40927;
  assign n40929 = ~pi1157 & ~n40920;
  assign n40930 = ~n40928 & n40929;
  assign n40931 = ~n40918 & ~n40930;
  assign n40932 = pi211 & ~n40931;
  assign n40933 = n40905 & n40924;
  assign n40934 = ~pi1155 & n40912;
  assign n40935 = pi200 & pi1091;
  assign n40936 = ~pi299 & n40935;
  assign n40937 = n40797 & ~n40936;
  assign n40938 = ~pi1156 & ~n40937;
  assign n40939 = ~n40934 & n40938;
  assign n40940 = ~n40933 & ~n40939;
  assign n40941 = pi1157 & ~n40940;
  assign n40942 = pi1091 & ~n11420;
  assign n40943 = n40925 & ~n40942;
  assign n40944 = ~n40923 & ~n40943;
  assign n40945 = pi200 & ~pi1156;
  assign n40946 = n40903 & n40945;
  assign n40947 = ~n40944 & ~n40946;
  assign n40948 = ~pi1157 & ~n40947;
  assign n40949 = ~pi211 & ~n40948;
  assign n40950 = ~n40941 & n40949;
  assign n40951 = ~n40932 & ~n40950;
  assign n40952 = ~pi219 & ~n40951;
  assign n40953 = n39235 & ~n40906;
  assign n40954 = ~n40916 & n40953;
  assign n40955 = pi299 & pi1091;
  assign n40956 = n40947 & ~n40955;
  assign n40957 = ~pi1157 & ~n40956;
  assign n40958 = pi1091 & n38484;
  assign n40959 = n40925 & ~n40958;
  assign n40960 = ~n40937 & ~n40959;
  assign n40961 = ~pi1156 & ~n40960;
  assign n40962 = n38365 & ~n40961;
  assign n40963 = n40909 & n40962;
  assign n40964 = pi219 & ~n40954;
  assign n40965 = ~n40957 & ~n40963;
  assign n40966 = n40964 & n40965;
  assign n40967 = ~n40952 & ~n40966;
  assign n40968 = ~n40836 & ~n40967;
  assign n40969 = ~po1038 & ~n40968;
  assign n40970 = ~n40902 & n40969;
  assign n40971 = ~pi243 & n40713;
  assign n40972 = pi243 & n40740;
  assign n40973 = n38365 & ~n40704;
  assign n40974 = ~n40738 & n40973;
  assign n40975 = ~n40972 & ~n40974;
  assign n40976 = ~n40971 & n40975;
  assign n40977 = pi219 & ~n40976;
  assign n40978 = n40704 & n40723;
  assign n40979 = ~pi243 & n40722;
  assign n40980 = ~n38359 & ~n38366;
  assign n40981 = pi1091 & n40980;
  assign n40982 = ~pi219 & ~n40981;
  assign n40983 = ~n40979 & n40982;
  assign n40984 = ~n40978 & n40983;
  assign n40985 = ~n40977 & ~n40984;
  assign n40986 = n40836 & ~n40985;
  assign n40987 = ~pi219 & ~n40980;
  assign n40988 = pi1157 & n38395;
  assign n40989 = ~n40987 & ~n40988;
  assign n40990 = pi1091 & ~n40989;
  assign n40991 = ~n40790 & ~n40990;
  assign n40992 = ~n40836 & ~n40991;
  assign n40993 = po1038 & ~n40992;
  assign n40994 = ~n40986 & n40993;
  assign n40995 = pi272 & pi283;
  assign n40996 = pi275 & n40995;
  assign n40997 = pi268 & n40996;
  assign n40998 = ~n40994 & n40997;
  assign n40999 = ~n40970 & n40998;
  assign n41000 = ~po1038 & n40967;
  assign n41001 = po1038 & n40991;
  assign n41002 = ~n40997 & ~n41001;
  assign n41003 = ~n41000 & n41002;
  assign n41004 = ~pi230 & ~n41003;
  assign n41005 = ~n40999 & n41004;
  assign n41006 = ~n16429 & ~n40989;
  assign n41007 = pi199 & ~n39439;
  assign n41008 = ~n38722 & ~n40945;
  assign n41009 = ~n41007 & n41008;
  assign n41010 = n16429 & n41009;
  assign n41011 = pi230 & ~n41006;
  assign n41012 = ~n41010 & n41011;
  assign po400 = ~n41005 & ~n41012;
  assign n41014 = ~pi230 & ~pi244;
  assign n41015 = pi213 & ~n40323;
  assign n41016 = ~n38639 & n40198;
  assign n41017 = ~n40317 & ~n41016;
  assign n41018 = ~n40204 & ~n41017;
  assign n41019 = pi214 & ~n41018;
  assign n41020 = n40296 & ~n41019;
  assign n41021 = ~pi214 & n41017;
  assign n41022 = n38297 & n40159;
  assign n41023 = pi212 & ~n41022;
  assign n41024 = ~n41021 & n41023;
  assign n41025 = ~n40204 & n41024;
  assign n41026 = ~pi219 & ~n41020;
  assign n41027 = ~n41025 & n41026;
  assign n41028 = ~pi211 & ~n38604;
  assign n41029 = ~n40289 & n41028;
  assign n41030 = ~n40288 & ~n41029;
  assign n41031 = n40286 & ~n41030;
  assign n41032 = n40255 & ~n41031;
  assign n41033 = ~n41027 & n41032;
  assign n41034 = ~n40197 & n41024;
  assign n41035 = pi214 & n41017;
  assign n41036 = n40263 & ~n41035;
  assign n41037 = ~pi219 & ~n41036;
  assign n41038 = ~n41034 & n41037;
  assign n41039 = pi299 & n39284;
  assign n41040 = pi1147 & ~n41039;
  assign n41041 = n40239 & n41040;
  assign n41042 = ~n41038 & n41041;
  assign n41043 = ~pi213 & ~n39286;
  assign n41044 = ~n41042 & n41043;
  assign n41045 = ~n41033 & n41044;
  assign n41046 = ~n41015 & ~n41045;
  assign n41047 = pi209 & ~n41046;
  assign n41048 = n40075 & ~n40081;
  assign n41049 = ~n40088 & ~n41048;
  assign n41050 = n40075 & ~n40080;
  assign n41051 = ~n10708 & n40092;
  assign n41052 = n10708 & ~n40097;
  assign n41053 = n38669 & ~n41051;
  assign n41054 = ~n41052 & n41053;
  assign n41055 = ~n41050 & n41054;
  assign n41056 = ~n39264 & ~n40111;
  assign n41057 = ~n41055 & n41056;
  assign n41058 = ~po1038 & ~n41057;
  assign n41059 = ~n41049 & ~n41058;
  assign n41060 = pi213 & ~n41059;
  assign n41061 = ~pi213 & ~n39293;
  assign n41062 = ~pi209 & ~n41061;
  assign n41063 = ~n41060 & n41062;
  assign n41064 = ~n41047 & ~n41063;
  assign n41065 = pi230 & ~n41064;
  assign po401 = ~n41014 & ~n41065;
  assign n41067 = pi1146 & n39740;
  assign n41068 = ~pi1147 & ~n41067;
  assign n41069 = n39721 & ~n39995;
  assign n41070 = n41068 & ~n41069;
  assign n41071 = ~n38290 & n40652;
  assign n41072 = n40664 & ~n41071;
  assign n41073 = ~po1038 & ~n41072;
  assign n41074 = pi214 & ~n40091;
  assign n41075 = ~pi299 & ~n40654;
  assign n41076 = n41074 & ~n41075;
  assign n41077 = pi212 & ~n41076;
  assign n41078 = ~pi299 & n40645;
  assign n41079 = ~pi211 & ~n41078;
  assign n41080 = n40644 & ~n41079;
  assign n41081 = ~pi214 & n41080;
  assign n41082 = n41077 & ~n41081;
  assign n41083 = n40659 & ~n41080;
  assign n41084 = ~pi219 & ~n41083;
  assign n41085 = ~n41082 & n41084;
  assign n41086 = n41073 & ~n41085;
  assign n41087 = n41070 & ~n41086;
  assign n41088 = pi1147 & ~n39721;
  assign n41089 = ~n41067 & n41088;
  assign n41090 = n40651 & ~n41079;
  assign n41091 = pi214 & ~n41090;
  assign n41092 = ~pi214 & ~n41078;
  assign n41093 = ~n41091 & ~n41092;
  assign n41094 = pi212 & ~n41093;
  assign n41095 = n40659 & ~n41078;
  assign n41096 = ~pi219 & ~n41095;
  assign n41097 = ~n41094 & n41096;
  assign n41098 = n41073 & ~n41097;
  assign n41099 = n41089 & ~n41098;
  assign n41100 = pi1148 & ~n41087;
  assign n41101 = ~n41099 & n41100;
  assign n41102 = ~n40241 & ~n41089;
  assign n41103 = ~n13025 & n40644;
  assign n41104 = ~pi214 & ~n41103;
  assign n41105 = ~n41091 & ~n41104;
  assign n41106 = pi212 & ~n41105;
  assign n41107 = n40659 & ~n41103;
  assign n41108 = ~pi219 & ~n41107;
  assign n41109 = ~n41106 & n41108;
  assign n41110 = n41073 & ~n41109;
  assign n41111 = ~n41102 & ~n41110;
  assign n41112 = ~n40658 & n41077;
  assign n41113 = ~pi212 & ~n40644;
  assign n41114 = ~pi219 & ~n41113;
  assign n41115 = ~n41112 & n41114;
  assign n41116 = n41073 & ~n41115;
  assign n41117 = n41068 & ~n41116;
  assign n41118 = ~pi1148 & ~n41111;
  assign n41119 = ~n41117 & n41118;
  assign n41120 = ~n41101 & ~n41119;
  assign n41121 = pi213 & ~n41120;
  assign n41122 = ~pi213 & ~n40669;
  assign n41123 = ~pi209 & ~n41122;
  assign n41124 = ~n41121 & n41123;
  assign n41125 = pi199 & pi1146;
  assign n41126 = ~pi200 & ~n41125;
  assign n41127 = n40182 & ~n41126;
  assign n41128 = pi207 & n41127;
  assign n41129 = pi1146 & ~n38484;
  assign n41130 = ~n41128 & ~n41129;
  assign n41131 = pi208 & ~n41130;
  assign n41132 = n38483 & ~n41125;
  assign n41133 = n40182 & ~n41132;
  assign n41134 = pi208 & n41133;
  assign n41135 = ~pi207 & ~n41134;
  assign n41136 = n39502 & ~n41132;
  assign n41137 = ~n41135 & n41136;
  assign n41138 = ~pi208 & n40090;
  assign n41139 = ~n41131 & ~n41138;
  assign n41140 = ~n41137 & n41139;
  assign n41141 = ~pi299 & ~n41140;
  assign n41142 = ~pi214 & ~n41141;
  assign n41143 = ~pi212 & ~n41142;
  assign n41144 = ~n10463 & ~n39503;
  assign n41145 = n41127 & ~n41144;
  assign n41146 = pi211 & ~n41145;
  assign n41147 = ~pi299 & ~n41127;
  assign n41148 = ~n41140 & ~n41147;
  assign n41149 = ~pi299 & ~n41148;
  assign n41150 = ~pi211 & n41149;
  assign n41151 = ~n41146 & ~n41150;
  assign n41152 = ~n41141 & ~n41151;
  assign n41153 = n41143 & ~n41152;
  assign n41154 = ~pi219 & ~n41153;
  assign n41155 = n41074 & ~n41141;
  assign n41156 = ~pi214 & n41152;
  assign n41157 = pi212 & ~n41156;
  assign n41158 = ~n41155 & n41157;
  assign n41159 = n41154 & ~n41158;
  assign n41160 = ~n38291 & n41141;
  assign n41161 = pi219 & ~n41160;
  assign n41162 = n38291 & ~n41140;
  assign n41163 = n41161 & ~n41162;
  assign n41164 = ~po1038 & ~n41163;
  assign n41165 = ~n41159 & n41164;
  assign n41166 = n41070 & ~n41165;
  assign n41167 = pi207 & n41133;
  assign n41168 = n38415 & ~n41126;
  assign n41169 = ~pi207 & n41168;
  assign n41170 = ~n40090 & ~n41169;
  assign n41171 = ~n41167 & n41170;
  assign n41172 = pi208 & ~pi299;
  assign n41173 = ~n41171 & n41172;
  assign n41174 = n38326 & n38415;
  assign n41175 = ~n41132 & n41174;
  assign n41176 = ~n41134 & ~n41175;
  assign n41177 = ~n41173 & n41176;
  assign n41178 = ~pi214 & n41177;
  assign n41179 = ~pi212 & ~n41178;
  assign n41180 = ~pi299 & n41177;
  assign n41181 = n41179 & ~n41180;
  assign n41182 = ~pi219 & ~n41181;
  assign n41183 = pi212 & ~n41180;
  assign n41184 = ~n40090 & n41177;
  assign n41185 = n10654 & n41184;
  assign n41186 = n41183 & ~n41185;
  assign n41187 = n41182 & ~n41186;
  assign n41188 = ~n38291 & ~n41177;
  assign n41189 = pi219 & ~n41188;
  assign n41190 = n38291 & ~n41184;
  assign n41191 = n41189 & ~n41190;
  assign n41192 = ~po1038 & ~n41191;
  assign n41193 = ~n41187 & n41192;
  assign n41194 = n41089 & ~n41193;
  assign n41195 = pi1148 & ~n41194;
  assign n41196 = ~n41166 & n41195;
  assign n41197 = n38326 & n41168;
  assign n41198 = ~n41173 & ~n41197;
  assign n41199 = ~n13025 & n41198;
  assign n41200 = pi214 & ~n41199;
  assign n41201 = ~pi214 & ~n41198;
  assign n41202 = ~pi212 & ~n41201;
  assign n41203 = ~n41200 & n41202;
  assign n41204 = ~pi214 & ~n41199;
  assign n41205 = ~n40090 & n41198;
  assign n41206 = ~pi299 & n41205;
  assign n41207 = pi214 & ~n41206;
  assign n41208 = ~pi211 & ~n41180;
  assign n41209 = n41177 & ~n41208;
  assign n41210 = n41207 & ~n41209;
  assign n41211 = pi212 & ~n41210;
  assign n41212 = ~n41204 & n41211;
  assign n41213 = ~n41203 & ~n41212;
  assign n41214 = ~pi219 & ~n41213;
  assign n41215 = ~pi1146 & ~n38592;
  assign n41216 = n40165 & ~n41215;
  assign n41217 = n41214 & ~n41216;
  assign n41218 = ~n38290 & ~n41198;
  assign n41219 = ~n38291 & ~n41218;
  assign n41220 = ~n41205 & ~n41219;
  assign n41221 = ~pi212 & n41201;
  assign n41222 = pi219 & ~n41221;
  assign n41223 = ~n41220 & n41222;
  assign n41224 = ~po1038 & ~n41223;
  assign n41225 = ~n41217 & n41224;
  assign n41226 = ~n41102 & ~n41225;
  assign n41227 = ~n40513 & ~n41141;
  assign n41228 = ~n41130 & ~n41227;
  assign n41229 = ~pi219 & ~n41228;
  assign n41230 = pi219 & ~n41145;
  assign n41231 = ~n38839 & ~n41230;
  assign n41232 = ~n38290 & ~n41146;
  assign n41233 = n41148 & n41232;
  assign n41234 = ~n41231 & ~n41233;
  assign n41235 = ~po1038 & ~n41234;
  assign n41236 = ~n41229 & n41235;
  assign n41237 = n41068 & ~n41236;
  assign n41238 = ~pi1148 & ~n41237;
  assign n41239 = ~n41226 & n41238;
  assign n41240 = ~n41196 & ~n41239;
  assign n41241 = pi213 & ~n41240;
  assign n41242 = ~pi214 & n41145;
  assign n41243 = ~n40097 & ~n41141;
  assign n41244 = pi214 & ~n41149;
  assign n41245 = ~n41243 & n41244;
  assign n41246 = ~n41242 & ~n41245;
  assign n41247 = ~pi212 & ~n41246;
  assign n41248 = pi299 & ~n40623;
  assign n41249 = ~n41141 & ~n41248;
  assign n41250 = pi212 & ~n41249;
  assign n41251 = ~n41147 & n41250;
  assign n41252 = ~pi219 & ~n41251;
  assign n41253 = ~n41247 & n41252;
  assign n41254 = ~n38639 & ~n41149;
  assign n41255 = ~pi211 & ~n41254;
  assign n41256 = n41232 & ~n41255;
  assign n41257 = ~n41231 & ~n41256;
  assign n41258 = n40255 & ~n41257;
  assign n41259 = ~n41253 & n41258;
  assign n41260 = ~n40097 & n41177;
  assign n41261 = n41207 & ~n41260;
  assign n41262 = ~n41201 & ~n41261;
  assign n41263 = ~pi212 & ~n41262;
  assign n41264 = n41177 & ~n41248;
  assign n41265 = pi212 & ~n41264;
  assign n41266 = ~n41206 & n41265;
  assign n41267 = ~pi219 & ~n41266;
  assign n41268 = ~n41263 & n41267;
  assign n41269 = ~n38637 & n41177;
  assign n41270 = ~n41206 & ~n41269;
  assign n41271 = ~pi211 & ~n41270;
  assign n41272 = ~n41219 & ~n41271;
  assign n41273 = n41222 & ~n41272;
  assign n41274 = pi1147 & ~po1038;
  assign n41275 = ~n41273 & n41274;
  assign n41276 = ~n41268 & n41275;
  assign n41277 = ~pi1148 & ~n40630;
  assign n41278 = ~n41276 & n41277;
  assign n41279 = ~n41259 & n41278;
  assign n41280 = n41143 & ~n41243;
  assign n41281 = ~pi219 & ~n41250;
  assign n41282 = ~n41280 & n41281;
  assign n41283 = ~pi299 & n41140;
  assign n41284 = n38291 & ~n41283;
  assign n41285 = ~n38639 & n41284;
  assign n41286 = n41161 & ~n41285;
  assign n41287 = n40255 & ~n41286;
  assign n41288 = ~n41282 & n41287;
  assign n41289 = n41179 & ~n41260;
  assign n41290 = ~pi219 & ~n41265;
  assign n41291 = ~n41289 & n41290;
  assign n41292 = n38291 & ~n41269;
  assign n41293 = n41189 & ~n41292;
  assign n41294 = n41274 & ~n41293;
  assign n41295 = ~n41291 & n41294;
  assign n41296 = pi1148 & ~n40630;
  assign n41297 = ~n41295 & n41296;
  assign n41298 = ~n41288 & n41297;
  assign n41299 = ~pi213 & ~n41298;
  assign n41300 = ~n41279 & n41299;
  assign n41301 = pi209 & ~n41300;
  assign n41302 = ~n41241 & n41301;
  assign n41303 = ~n41124 & ~n41302;
  assign n41304 = pi230 & ~n41303;
  assign n41305 = ~pi230 & ~pi245;
  assign po402 = ~n41304 & ~n41305;
  assign n41307 = ~pi1150 & n39989;
  assign n41308 = pi1150 & n39948;
  assign n41309 = pi1149 & ~n41307;
  assign n41310 = ~n41308 & n41309;
  assign n41311 = pi1150 & n40016;
  assign n41312 = ~pi1150 & n40053;
  assign n41313 = ~pi1149 & ~n41312;
  assign n41314 = ~n41311 & n41313;
  assign n41315 = ~n41310 & ~n41314;
  assign n41316 = pi1148 & ~n41315;
  assign n41317 = ~pi1150 & n39980;
  assign n41318 = pi1150 & n39940;
  assign n41319 = pi1149 & ~n41318;
  assign n41320 = ~n41317 & n41319;
  assign n41321 = ~pi1149 & pi1150;
  assign n41322 = ~n40021 & n41321;
  assign n41323 = ~n41320 & ~n41322;
  assign n41324 = ~pi1148 & ~n41323;
  assign n41325 = ~n41316 & ~n41324;
  assign n41326 = pi213 & ~n41325;
  assign n41327 = ~n41070 & ~n41089;
  assign n41328 = pi219 & ~n40090;
  assign n41329 = n39943 & ~n41328;
  assign n41330 = n39986 & ~n40034;
  assign n41331 = ~n41329 & ~n41330;
  assign n41332 = ~n40036 & ~n40106;
  assign n41333 = n38300 & ~n41332;
  assign n41334 = ~n40498 & ~n41333;
  assign n41335 = ~pi219 & ~n41334;
  assign n41336 = ~n41331 & ~n41335;
  assign n41337 = ~n41327 & ~n41336;
  assign n41338 = ~n40037 & ~n40046;
  assign n41339 = n41070 & ~n41338;
  assign n41340 = ~pi1150 & ~n41339;
  assign n41341 = ~n41337 & n41340;
  assign n41342 = ~n40122 & ~n41329;
  assign n41343 = ~pi214 & n39542;
  assign n41344 = pi214 & ~n39997;
  assign n41345 = n40124 & n41344;
  assign n41346 = pi212 & ~n41345;
  assign n41347 = ~n41343 & n41346;
  assign n41348 = n40006 & ~n41347;
  assign n41349 = ~n41342 & ~n41348;
  assign n41350 = n41070 & ~n41349;
  assign n41351 = ~n40126 & n40362;
  assign n41352 = ~pi212 & ~n39505;
  assign n41353 = ~pi219 & ~n41352;
  assign n41354 = ~n40374 & n41353;
  assign n41355 = ~n41351 & n41354;
  assign n41356 = ~n41342 & ~n41355;
  assign n41357 = n41089 & ~n41356;
  assign n41358 = pi1150 & ~n41357;
  assign n41359 = ~n41350 & n41358;
  assign n41360 = ~n41341 & ~n41359;
  assign n41361 = pi1148 & ~n41360;
  assign n41362 = ~pi219 & ~n40065;
  assign n41363 = ~n40514 & ~n41362;
  assign n41364 = n41329 & n41363;
  assign n41365 = n41068 & ~n41364;
  assign n41366 = ~n41102 & ~n41329;
  assign n41367 = ~n41365 & ~n41366;
  assign n41368 = pi1150 & n40018;
  assign n41369 = ~n41367 & ~n41368;
  assign n41370 = pi1150 & n39549;
  assign n41371 = pi299 & n39952;
  assign n41372 = ~pi219 & ~n41371;
  assign n41373 = ~n41216 & n41372;
  assign n41374 = ~n41370 & n41373;
  assign n41375 = ~n41102 & n41374;
  assign n41376 = ~pi1148 & ~n41375;
  assign n41377 = ~n41369 & n41376;
  assign n41378 = ~n41361 & ~n41377;
  assign n41379 = ~pi1149 & ~n41378;
  assign n41380 = n40065 & n40159;
  assign n41381 = ~n39577 & ~n41380;
  assign n41382 = n39976 & n41381;
  assign n41383 = ~pi1146 & n39977;
  assign n41384 = n39943 & ~n39960;
  assign n41385 = ~n39978 & ~n41384;
  assign n41386 = ~n41383 & ~n41385;
  assign n41387 = ~n41382 & n41386;
  assign n41388 = ~n41102 & ~n41387;
  assign n41389 = ~n39577 & n40514;
  assign n41390 = ~n41385 & ~n41389;
  assign n41391 = ~pi1146 & ~n39577;
  assign n41392 = n41390 & ~n41391;
  assign n41393 = n41068 & ~n41392;
  assign n41394 = ~pi1150 & ~n41393;
  assign n41395 = ~n41388 & n41394;
  assign n41396 = ~pi214 & n40578;
  assign n41397 = n39936 & ~n41396;
  assign n41398 = ~pi219 & ~n41397;
  assign n41399 = ~n39920 & ~n40578;
  assign n41400 = ~pi212 & n41399;
  assign n41401 = n41398 & ~n41400;
  assign n41402 = ~pi299 & n39925;
  assign n41403 = ~n39926 & ~n40090;
  assign n41404 = ~n41402 & n41403;
  assign n41405 = n41401 & n41404;
  assign n41406 = ~n40145 & ~n41329;
  assign n41407 = n41398 & ~n41399;
  assign n41408 = ~n41406 & ~n41407;
  assign n41409 = ~n41405 & n41408;
  assign n41410 = ~n39918 & ~n41409;
  assign n41411 = n39921 & ~n39935;
  assign n41412 = ~pi219 & ~n41411;
  assign n41413 = ~n40582 & n41412;
  assign n41414 = n40144 & ~n41413;
  assign n41415 = ~n41410 & n41414;
  assign n41416 = n41068 & ~n41415;
  assign n41417 = ~n41102 & ~n41409;
  assign n41418 = pi1150 & ~n41417;
  assign n41419 = ~n41416 & n41418;
  assign n41420 = ~pi1148 & ~n41419;
  assign n41421 = ~n41395 & n41420;
  assign n41422 = ~n39986 & ~n41329;
  assign n41423 = ~n40027 & n40043;
  assign n41424 = ~n40030 & ~n41423;
  assign n41425 = ~n41070 & ~n41424;
  assign n41426 = ~n39615 & n41074;
  assign n41427 = n40042 & ~n41426;
  assign n41428 = n40045 & ~n41427;
  assign n41429 = ~n41425 & n41428;
  assign n41430 = ~n41422 & ~n41429;
  assign n41431 = ~n41327 & ~n41430;
  assign n41432 = ~pi1150 & ~n41431;
  assign n41433 = ~n40169 & ~n41364;
  assign n41434 = n41070 & n41433;
  assign n41435 = pi214 & n40158;
  assign n41436 = n40164 & ~n41435;
  assign n41437 = ~pi219 & ~n40161;
  assign n41438 = ~n41436 & n41437;
  assign n41439 = n40157 & ~n41438;
  assign n41440 = pi1146 & n39944;
  assign n41441 = n41089 & ~n41440;
  assign n41442 = ~n41439 & n41441;
  assign n41443 = pi1150 & ~n41442;
  assign n41444 = ~n41434 & n41443;
  assign n41445 = pi1148 & ~n41444;
  assign n41446 = ~n41432 & n41445;
  assign n41447 = pi1149 & ~n41446;
  assign n41448 = ~n41421 & n41447;
  assign n41449 = ~n41379 & ~n41448;
  assign n41450 = ~pi213 & ~n41449;
  assign n41451 = pi209 & ~n41326;
  assign n41452 = ~n41450 & n41451;
  assign n41453 = ~pi212 & ~n41242;
  assign n41454 = ~n13025 & ~n41145;
  assign n41455 = pi214 & ~n41454;
  assign n41456 = n41453 & ~n41455;
  assign n41457 = ~pi214 & ~n41454;
  assign n41458 = pi214 & n41151;
  assign n41459 = pi212 & ~n41458;
  assign n41460 = ~n41457 & n41459;
  assign n41461 = ~n41456 & ~n41460;
  assign n41462 = ~pi219 & ~n41461;
  assign n41463 = n40255 & ~n41230;
  assign n41464 = ~n41462 & n41463;
  assign n41465 = pi219 & n41198;
  assign n41466 = n41274 & ~n41465;
  assign n41467 = ~n41214 & n41466;
  assign n41468 = ~pi1150 & ~n39955;
  assign n41469 = ~n41467 & n41468;
  assign n41470 = ~n41464 & n41469;
  assign n41471 = ~n41244 & n41453;
  assign n41472 = ~pi214 & ~n41149;
  assign n41473 = n41459 & ~n41472;
  assign n41474 = ~n41471 & ~n41473;
  assign n41475 = ~pi219 & ~n41474;
  assign n41476 = ~n41230 & ~n41475;
  assign n41477 = ~pi1147 & ~n41476;
  assign n41478 = n41202 & ~n41207;
  assign n41479 = ~pi214 & ~n41206;
  assign n41480 = n41211 & ~n41479;
  assign n41481 = ~n41478 & ~n41480;
  assign n41482 = ~pi219 & ~n41481;
  assign n41483 = ~n41465 & ~n41482;
  assign n41484 = pi1147 & ~n41483;
  assign n41485 = ~po1038 & ~n41484;
  assign n41486 = ~n41477 & n41485;
  assign n41487 = pi1150 & ~n39721;
  assign n41488 = ~n41486 & n41487;
  assign n41489 = ~n41470 & ~n41488;
  assign n41490 = pi1149 & ~n41489;
  assign n41491 = pi1150 & n40085;
  assign n41492 = ~pi1147 & n41148;
  assign n41493 = n16429 & ~n41492;
  assign n41494 = n41491 & ~n41493;
  assign n41495 = pi1147 & n41198;
  assign n41496 = n41145 & ~n41491;
  assign n41497 = ~pi1147 & ~n41496;
  assign n41498 = ~po1038 & ~n41497;
  assign n41499 = ~n41495 & n41498;
  assign n41500 = ~pi1149 & ~n41499;
  assign n41501 = ~n41494 & n41500;
  assign n41502 = ~n41490 & ~n41501;
  assign n41503 = ~pi1148 & ~n41502;
  assign n41504 = n41161 & ~n41284;
  assign n41505 = n40255 & ~n41504;
  assign n41506 = ~n41141 & n41454;
  assign n41507 = pi214 & n41506;
  assign n41508 = n41157 & ~n41507;
  assign n41509 = n41154 & ~n41508;
  assign n41510 = n41505 & ~n41509;
  assign n41511 = ~n38290 & n41208;
  assign n41512 = n41189 & ~n41511;
  assign n41513 = n41274 & ~n41512;
  assign n41514 = pi214 & ~n13025;
  assign n41515 = n41177 & n41514;
  assign n41516 = pi212 & ~n41515;
  assign n41517 = ~pi214 & n41209;
  assign n41518 = n41516 & ~n41517;
  assign n41519 = n41179 & ~n41209;
  assign n41520 = ~pi219 & ~n41519;
  assign n41521 = ~n41518 & n41520;
  assign n41522 = n41513 & ~n41521;
  assign n41523 = pi1150 & ~n39996;
  assign n41524 = ~n41522 & n41523;
  assign n41525 = ~n41510 & n41524;
  assign n41526 = ~pi219 & n41227;
  assign n41527 = n41505 & ~n41526;
  assign n41528 = ~n41178 & n41516;
  assign n41529 = ~pi212 & ~n41177;
  assign n41530 = ~pi219 & ~n41529;
  assign n41531 = ~n41528 & n41530;
  assign n41532 = n41513 & ~n41531;
  assign n41533 = ~pi1150 & ~n39740;
  assign n41534 = ~n41532 & n41533;
  assign n41535 = ~n41527 & n41534;
  assign n41536 = ~pi1149 & ~n41535;
  assign n41537 = ~n41525 & n41536;
  assign n41538 = n41182 & ~n41183;
  assign n41539 = ~n41512 & ~n41538;
  assign n41540 = n6294 & n41539;
  assign n41541 = ~n6294 & ~n38670;
  assign n41542 = ~pi57 & pi1147;
  assign n41543 = ~n41541 & n41542;
  assign n41544 = ~n41540 & n41543;
  assign n41545 = pi57 & n38670;
  assign n41546 = n6294 & ~n38669;
  assign n41547 = n41160 & n41546;
  assign n41548 = ~n38670 & ~n41283;
  assign n41549 = ~pi57 & ~pi1147;
  assign n41550 = ~n41541 & n41549;
  assign n41551 = ~n41548 & n41550;
  assign n41552 = ~n41547 & n41551;
  assign n41553 = ~n41545 & ~n41552;
  assign n41554 = ~n41544 & n41553;
  assign n41555 = pi1150 & ~n41554;
  assign n41556 = ~n41244 & n41506;
  assign n41557 = pi212 & ~n41556;
  assign n41558 = n41143 & ~n41507;
  assign n41559 = ~pi219 & ~n41558;
  assign n41560 = ~n41557 & n41559;
  assign n41561 = n41505 & ~n41560;
  assign n41562 = ~n40526 & n41274;
  assign n41563 = n41539 & n41562;
  assign n41564 = ~pi1150 & ~n39987;
  assign n41565 = ~n41563 & n41564;
  assign n41566 = ~n41561 & n41565;
  assign n41567 = pi1149 & ~n41566;
  assign n41568 = ~n41555 & n41567;
  assign n41569 = pi1148 & ~n41568;
  assign n41570 = ~n41537 & n41569;
  assign n41571 = pi213 & ~n41570;
  assign n41572 = ~n41503 & n41571;
  assign n41573 = ~pi213 & ~n41240;
  assign n41574 = ~pi209 & ~n41573;
  assign n41575 = ~n41572 & n41574;
  assign n41576 = ~n41452 & ~n41575;
  assign n41577 = pi230 & ~n41576;
  assign n41578 = ~pi230 & ~pi246;
  assign po403 = ~n41577 & ~n41578;
  assign n41580 = ~pi1147 & ~n40457;
  assign n41581 = pi1151 & ~n39955;
  assign n41582 = ~n39919 & ~n41401;
  assign n41583 = n41581 & ~n41582;
  assign n41584 = n41580 & ~n41583;
  assign n41585 = pi1151 & ~n39987;
  assign n41586 = n40144 & ~n41407;
  assign n41587 = n41585 & ~n41586;
  assign n41588 = n39959 & ~n39974;
  assign n41589 = ~n41385 & ~n41588;
  assign n41590 = ~n39987 & ~n41589;
  assign n41591 = ~pi1151 & n41590;
  assign n41592 = pi1147 & ~n41587;
  assign n41593 = ~n41591 & n41592;
  assign n41594 = ~pi1149 & ~n41593;
  assign n41595 = ~n41584 & n41594;
  assign n41596 = ~pi1151 & ~n39721;
  assign n41597 = n40045 & ~n41423;
  assign n41598 = n40530 & ~n41597;
  assign n41599 = ~n40031 & n40530;
  assign n41600 = ~n41598 & ~n41599;
  assign n41601 = n41596 & n41600;
  assign n41602 = n40349 & ~n41439;
  assign n41603 = ~pi1147 & ~n41602;
  assign n41604 = ~n41601 & n41603;
  assign n41605 = pi1147 & ~n40470;
  assign n41606 = ~n39944 & ~n39947;
  assign n41607 = n40522 & n41606;
  assign n41608 = n41605 & ~n41607;
  assign n41609 = pi1149 & ~n41608;
  assign n41610 = ~n41604 & n41609;
  assign n41611 = pi1150 & ~n41610;
  assign n41612 = ~n41595 & n41611;
  assign n41613 = pi212 & ~n39529;
  assign n41614 = n41354 & ~n41613;
  assign n41615 = n40014 & ~n41614;
  assign n41616 = n40430 & ~n41615;
  assign n41617 = pi1147 & ~n41616;
  assign n41618 = n38300 & ~n40028;
  assign n41619 = ~n40036 & ~n41618;
  assign n41620 = n40503 & n41619;
  assign n41621 = ~pi1151 & ~n39947;
  assign n41622 = ~n41620 & n41621;
  assign n41623 = ~n40051 & n41622;
  assign n41624 = n41617 & ~n41623;
  assign n41625 = ~n40363 & n41354;
  assign n41626 = n40122 & ~n41625;
  assign n41627 = ~n39721 & ~n41626;
  assign n41628 = pi1151 & n41627;
  assign n41629 = n41596 & ~n41620;
  assign n41630 = ~pi1147 & ~n41629;
  assign n41631 = ~n41628 & n41630;
  assign n41632 = pi1149 & ~n41631;
  assign n41633 = ~n41624 & n41632;
  assign n41634 = ~n39954 & n40019;
  assign n41635 = ~pi1151 & ~n41634;
  assign n41636 = ~pi1147 & ~n41635;
  assign n41637 = n39780 & ~n40382;
  assign n41638 = n41581 & ~n41637;
  assign n41639 = n41636 & ~n41638;
  assign n41640 = ~n40598 & n41585;
  assign n41641 = ~n39985 & n40436;
  assign n41642 = pi1147 & ~n41641;
  assign n41643 = ~n41640 & n41642;
  assign n41644 = ~pi1149 & ~n41639;
  assign n41645 = ~n41643 & n41644;
  assign n41646 = ~pi1150 & ~n41645;
  assign n41647 = ~n41633 & n41646;
  assign n41648 = ~n41612 & ~n41647;
  assign n41649 = pi1148 & ~n41648;
  assign n41650 = pi1147 & ~n40465;
  assign n41651 = ~pi1151 & ~n39996;
  assign n41652 = ~n40051 & n41651;
  assign n41653 = n41650 & ~n41652;
  assign n41654 = ~n40009 & n40122;
  assign n41655 = ~n40086 & ~n41654;
  assign n41656 = pi1151 & n41655;
  assign n41657 = ~pi1151 & ~n40086;
  assign n41658 = ~n40487 & n41657;
  assign n41659 = ~pi1147 & ~n41658;
  assign n41660 = ~n41656 & n41659;
  assign n41661 = ~pi1150 & ~n41660;
  assign n41662 = ~n41653 & n41661;
  assign n41663 = n40404 & n40516;
  assign n41664 = pi1147 & ~n41663;
  assign n41665 = ~n39996 & ~n40050;
  assign n41666 = ~pi1151 & n41665;
  assign n41667 = n41664 & ~n41666;
  assign n41668 = ~n41598 & n41657;
  assign n41669 = pi1151 & ~n40086;
  assign n41670 = ~n40169 & n41669;
  assign n41671 = ~pi1147 & ~n41670;
  assign n41672 = ~n41668 & n41671;
  assign n41673 = pi1150 & ~n41667;
  assign n41674 = ~n41672 & n41673;
  assign n41675 = ~n41662 & ~n41674;
  assign n41676 = pi1149 & ~n41675;
  assign n41677 = ~n41413 & n41586;
  assign n41678 = n39741 & ~n41677;
  assign n41679 = ~n39740 & ~n41390;
  assign n41680 = ~pi1151 & n41679;
  assign n41681 = pi1147 & ~n41680;
  assign n41682 = ~n41678 & n41681;
  assign n41683 = ~pi1151 & ~n40060;
  assign n41684 = ~pi1147 & ~n41683;
  assign n41685 = pi1151 & ~n39918;
  assign n41686 = n41684 & ~n41685;
  assign n41687 = pi1150 & ~n41686;
  assign n41688 = ~n41682 & n41687;
  assign n41689 = ~n39549 & n40514;
  assign n41690 = n40595 & ~n41689;
  assign n41691 = n39741 & ~n41690;
  assign n41692 = n40421 & ~n40515;
  assign n41693 = pi1147 & ~n41692;
  assign n41694 = ~n41691 & n41693;
  assign n41695 = ~pi1147 & pi1151;
  assign n41696 = n40018 & n41695;
  assign n41697 = ~pi1150 & ~n41696;
  assign n41698 = ~n41694 & n41697;
  assign n41699 = ~n41688 & ~n41698;
  assign n41700 = ~pi1149 & ~n41699;
  assign n41701 = ~pi1148 & ~n41700;
  assign n41702 = ~n41676 & n41701;
  assign n41703 = ~n41649 & ~n41702;
  assign n41704 = ~pi213 & ~n41703;
  assign n41705 = pi213 & n40475;
  assign n41706 = pi209 & ~n41705;
  assign n41707 = ~n41704 & n41706;
  assign n41708 = ~n41598 & n41669;
  assign n41709 = pi1147 & ~n40522;
  assign n41710 = ~n41708 & n41709;
  assign n41711 = ~po1038 & ~n40570;
  assign n41712 = ~n40573 & n41711;
  assign n41713 = ~n40331 & ~n41712;
  assign n41714 = n41684 & n41713;
  assign n41715 = ~pi1150 & ~n41714;
  assign n41716 = ~n41710 & n41715;
  assign n41717 = n39971 & n39978;
  assign n41718 = n40349 & ~n41717;
  assign n41719 = n41580 & ~n41718;
  assign n41720 = n40349 & n41600;
  assign n41721 = n40372 & ~n41599;
  assign n41722 = pi1147 & ~n41721;
  assign n41723 = ~n41720 & n41722;
  assign n41724 = pi1150 & ~n41723;
  assign n41725 = ~n41719 & n41724;
  assign n41726 = ~n41716 & ~n41725;
  assign n41727 = ~pi1149 & ~n41726;
  assign n41728 = n40421 & ~n41677;
  assign n41729 = ~n39996 & ~n41414;
  assign n41730 = pi1151 & n41729;
  assign n41731 = ~pi1147 & ~n41730;
  assign n41732 = ~n41728 & n41731;
  assign n41733 = ~n39945 & n41692;
  assign n41734 = n41664 & ~n41733;
  assign n41735 = ~pi1150 & ~n41734;
  assign n41736 = ~n41732 & n41735;
  assign n41737 = n40436 & ~n41586;
  assign n41738 = n39931 & ~n40149;
  assign n41739 = n40144 & ~n41738;
  assign n41740 = n40430 & ~n41739;
  assign n41741 = ~pi1147 & ~n41740;
  assign n41742 = ~n41737 & n41741;
  assign n41743 = ~n39987 & ~n40527;
  assign n41744 = ~pi1151 & n41743;
  assign n41745 = n41605 & ~n41744;
  assign n41746 = pi1150 & ~n41745;
  assign n41747 = ~n41742 & n41746;
  assign n41748 = ~n41736 & ~n41747;
  assign n41749 = pi1149 & ~n41748;
  assign n41750 = pi1148 & ~n41749;
  assign n41751 = ~n41727 & n41750;
  assign n41752 = ~pi219 & ~n40380;
  assign n41753 = ~n40492 & n41752;
  assign n41754 = n40014 & ~n41753;
  assign n41755 = ~n40010 & n41754;
  assign n41756 = n40421 & ~n41755;
  assign n41757 = n41650 & ~n41756;
  assign n41758 = n39566 & n39780;
  assign n41759 = ~n10708 & n41758;
  assign n41760 = ~n41690 & ~n41759;
  assign n41761 = n40404 & n41760;
  assign n41762 = n40421 & ~n41690;
  assign n41763 = ~pi1147 & ~n41762;
  assign n41764 = ~n41761 & n41763;
  assign n41765 = ~pi1150 & ~n41764;
  assign n41766 = ~n41757 & n41765;
  assign n41767 = ~n39987 & ~n41754;
  assign n41768 = ~pi1151 & n41767;
  assign n41769 = n41617 & ~n41768;
  assign n41770 = n40430 & ~n41758;
  assign n41771 = ~n40598 & n41770;
  assign n41772 = n40436 & ~n40598;
  assign n41773 = ~pi1147 & ~n41771;
  assign n41774 = ~n41772 & n41773;
  assign n41775 = pi1150 & ~n41774;
  assign n41776 = ~n41769 & n41775;
  assign n41777 = ~n41766 & ~n41776;
  assign n41778 = pi1149 & ~n41777;
  assign n41779 = n40038 & n40503;
  assign n41780 = ~n39955 & ~n41779;
  assign n41781 = ~pi1151 & n41780;
  assign n41782 = n40349 & ~n41620;
  assign n41783 = pi1147 & ~n41782;
  assign n41784 = ~n41781 & n41783;
  assign n41785 = ~n16429 & n39720;
  assign n41786 = pi1151 & ~n41785;
  assign n41787 = n41636 & ~n41786;
  assign n41788 = pi1150 & ~n41787;
  assign n41789 = ~n41784 & n41788;
  assign n41790 = ~n40086 & ~n40487;
  assign n41791 = ~pi1151 & ~n41330;
  assign n41792 = pi1147 & ~n41791;
  assign n41793 = ~n41790 & n41792;
  assign n41794 = n40020 & n41695;
  assign n41795 = ~pi1150 & ~n41794;
  assign n41796 = ~n41793 & n41795;
  assign n41797 = ~n41789 & ~n41796;
  assign n41798 = ~pi1149 & ~n41797;
  assign n41799 = ~pi1148 & ~n41798;
  assign n41800 = ~n41778 & n41799;
  assign n41801 = ~n41751 & ~n41800;
  assign n41802 = pi213 & ~n41801;
  assign n41803 = ~pi213 & ~n40058;
  assign n41804 = ~pi209 & ~n41803;
  assign n41805 = ~n41802 & n41804;
  assign n41806 = ~n41707 & ~n41805;
  assign n41807 = pi230 & ~n41806;
  assign n41808 = ~pi230 & ~pi247;
  assign po404 = ~n41807 & ~n41808;
  assign n41810 = pi1152 & ~n41772;
  assign n41811 = ~n41587 & n41810;
  assign n41812 = pi1151 & n41590;
  assign n41813 = ~pi1152 & ~n41641;
  assign n41814 = ~n41812 & n41813;
  assign n41815 = ~pi1150 & ~n41811;
  assign n41816 = ~n41814 & n41815;
  assign n41817 = pi1152 & ~n40470;
  assign n41818 = ~n41615 & n41621;
  assign n41819 = n41817 & ~n41818;
  assign n41820 = pi1151 & ~n39986;
  assign n41821 = n41606 & n41820;
  assign n41822 = ~pi1152 & ~n41821;
  assign n41823 = ~n41623 & n41822;
  assign n41824 = pi1150 & ~n41823;
  assign n41825 = ~n41819 & n41824;
  assign n41826 = pi1148 & ~n41816;
  assign n41827 = ~n41825 & n41826;
  assign n41828 = ~n39979 & n41581;
  assign n41829 = ~pi1152 & ~n41828;
  assign n41830 = ~n41635 & n41829;
  assign n41831 = n40372 & ~n41637;
  assign n41832 = pi1152 & ~n41831;
  assign n41833 = ~n41583 & n41832;
  assign n41834 = ~pi1150 & ~n41833;
  assign n41835 = ~n41830 & n41834;
  assign n41836 = ~pi1151 & n41627;
  assign n41837 = pi1152 & ~n41602;
  assign n41838 = ~n41836 & n41837;
  assign n41839 = ~pi1152 & ~n41629;
  assign n41840 = ~n41720 & n41839;
  assign n41841 = pi1150 & ~n41840;
  assign n41842 = ~n41838 & n41841;
  assign n41843 = ~pi1148 & ~n41842;
  assign n41844 = ~n41835 & n41843;
  assign n41845 = ~n41827 & ~n41844;
  assign n41846 = pi1149 & ~n41845;
  assign n41847 = ~n40015 & n41651;
  assign n41848 = pi1152 & ~n41847;
  assign n41849 = ~n41663 & n41848;
  assign n41850 = pi1151 & n41665;
  assign n41851 = ~pi1152 & ~n41652;
  assign n41852 = ~n41850 & n41851;
  assign n41853 = ~n41849 & ~n41852;
  assign n41854 = pi1150 & ~n41853;
  assign n41855 = ~n41678 & ~n41762;
  assign n41856 = pi1152 & ~n41855;
  assign n41857 = pi1151 & n41679;
  assign n41858 = ~n41692 & ~n41857;
  assign n41859 = ~pi1152 & ~n41858;
  assign n41860 = ~pi1150 & ~n41859;
  assign n41861 = ~n41856 & n41860;
  assign n41862 = pi1148 & ~n41861;
  assign n41863 = ~n41854 & n41862;
  assign n41864 = ~pi1151 & n41655;
  assign n41865 = pi1152 & ~n41670;
  assign n41866 = ~n41864 & n41865;
  assign n41867 = ~pi1152 & ~n41658;
  assign n41868 = ~n41708 & n41867;
  assign n41869 = pi1150 & ~n41868;
  assign n41870 = ~n41866 & n41869;
  assign n41871 = pi1151 & ~pi1152;
  assign n41872 = n40060 & n41871;
  assign n41873 = ~pi1151 & ~n40018;
  assign n41874 = pi1152 & ~n41685;
  assign n41875 = ~n41873 & n41874;
  assign n41876 = ~pi1150 & ~n41872;
  assign n41877 = ~n41875 & n41876;
  assign n41878 = ~n41870 & ~n41877;
  assign n41879 = ~pi1148 & ~n41878;
  assign n41880 = ~pi1149 & ~n41879;
  assign n41881 = ~n41863 & n41880;
  assign n41882 = ~n41846 & ~n41881;
  assign n41883 = ~pi213 & ~n41882;
  assign n41884 = ~n39980 & n41871;
  assign n41885 = ~pi1151 & ~n40020;
  assign n41886 = ~n40018 & n41885;
  assign n41887 = pi1152 & ~n41886;
  assign n41888 = ~n40458 & n41887;
  assign n41889 = ~pi1150 & ~n41888;
  assign n41890 = ~n41884 & n41889;
  assign n41891 = n41817 & ~n41847;
  assign n41892 = pi1151 & n39989;
  assign n41893 = ~pi1152 & ~n41892;
  assign n41894 = ~n40466 & n41893;
  assign n41895 = pi1150 & ~n41894;
  assign n41896 = ~n41891 & n41895;
  assign n41897 = ~n41890 & ~n41896;
  assign n41898 = pi213 & n41897;
  assign n41899 = pi209 & ~n41898;
  assign n41900 = ~n41883 & n41899;
  assign n41901 = ~n41683 & n41829;
  assign n41902 = ~pi1151 & ~n41713;
  assign n41903 = pi1152 & ~n41902;
  assign n41904 = ~n41718 & n41903;
  assign n41905 = ~pi1150 & ~n41904;
  assign n41906 = ~n41901 & n41905;
  assign n41907 = ~pi1152 & ~n41587;
  assign n41908 = ~n41728 & n41907;
  assign n41909 = ~pi1151 & n41729;
  assign n41910 = pi1152 & ~n41740;
  assign n41911 = ~n41909 & n41910;
  assign n41912 = pi1150 & ~n41911;
  assign n41913 = ~n41908 & n41912;
  assign n41914 = pi1149 & ~n41913;
  assign n41915 = ~n41906 & n41914;
  assign n41916 = n41651 & n41760;
  assign n41917 = pi1152 & ~n41771;
  assign n41918 = ~n41916 & n41917;
  assign n41919 = ~pi1152 & ~n41762;
  assign n41920 = ~n41640 & n41919;
  assign n41921 = pi1150 & ~n41920;
  assign n41922 = ~n41918 & n41921;
  assign n41923 = pi1152 & ~n41786;
  assign n41924 = ~n41885 & n41923;
  assign n41925 = n41634 & n41871;
  assign n41926 = ~pi1150 & ~n41925;
  assign n41927 = ~n41924 & n41926;
  assign n41928 = ~pi1149 & ~n41927;
  assign n41929 = ~n41922 & n41928;
  assign n41930 = ~pi1148 & ~n41929;
  assign n41931 = ~n41915 & n41930;
  assign n41932 = ~n41616 & n41848;
  assign n41933 = pi1151 & n41767;
  assign n41934 = ~pi1152 & ~n41756;
  assign n41935 = ~n41933 & n41934;
  assign n41936 = pi1150 & ~n41932;
  assign n41937 = ~n41935 & n41936;
  assign n41938 = pi1151 & n41780;
  assign n41939 = ~pi1152 & ~n41791;
  assign n41940 = ~n41938 & n41939;
  assign n41941 = pi1152 & ~n41658;
  assign n41942 = ~n41782 & n41941;
  assign n41943 = ~pi1150 & ~n41942;
  assign n41944 = ~n41940 & n41943;
  assign n41945 = ~pi1149 & ~n41944;
  assign n41946 = ~n41937 & n41945;
  assign n41947 = pi1152 & ~n41668;
  assign n41948 = ~n41720 & n41947;
  assign n41949 = n41581 & ~n41599;
  assign n41950 = n40523 & ~n41949;
  assign n41951 = ~pi1150 & ~n41950;
  assign n41952 = ~n41948 & n41951;
  assign n41953 = n40516 & n41651;
  assign n41954 = n41817 & ~n41953;
  assign n41955 = pi1151 & n41743;
  assign n41956 = ~pi1152 & ~n41733;
  assign n41957 = ~n41955 & n41956;
  assign n41958 = pi1150 & ~n41957;
  assign n41959 = ~n41954 & n41958;
  assign n41960 = pi1149 & ~n41959;
  assign n41961 = ~n41952 & n41960;
  assign n41962 = pi1148 & ~n41961;
  assign n41963 = ~n41946 & n41962;
  assign n41964 = pi213 & ~n41931;
  assign n41965 = ~n41963 & n41964;
  assign n41966 = ~pi213 & ~n41325;
  assign n41967 = ~pi209 & ~n41966;
  assign n41968 = ~n41965 & n41967;
  assign n41969 = ~n41900 & ~n41968;
  assign n41970 = pi230 & ~n41969;
  assign n41971 = ~pi230 & ~pi248;
  assign po405 = ~n41970 & ~n41971;
  assign n41973 = ~pi213 & n41897;
  assign n41974 = pi299 & n38700;
  assign n41975 = ~n40036 & ~n41974;
  assign n41976 = ~n39619 & n41975;
  assign n41977 = ~pi212 & ~n41976;
  assign n41978 = ~pi214 & n41975;
  assign n41979 = ~n39762 & ~n40035;
  assign n41980 = pi214 & ~n40485;
  assign n41981 = ~n41979 & n41980;
  assign n41982 = pi212 & ~n41981;
  assign n41983 = ~n41978 & n41982;
  assign n41984 = ~n41977 & ~n41983;
  assign n41985 = ~pi219 & ~n41984;
  assign n41986 = n6294 & ~n40502;
  assign n41987 = ~n41985 & n41986;
  assign n41988 = ~n6294 & n38703;
  assign n41989 = ~pi57 & ~pi1151;
  assign n41990 = ~n41988 & n41989;
  assign n41991 = ~n41987 & n41990;
  assign n41992 = pi57 & ~n38703;
  assign n41993 = ~n40532 & ~n41974;
  assign n41994 = ~pi214 & ~n41993;
  assign n41995 = ~n39598 & n39795;
  assign n41996 = pi212 & ~n41995;
  assign n41997 = ~n41994 & n41996;
  assign n41998 = pi214 & ~n41993;
  assign n41999 = ~pi212 & ~n39619;
  assign n42000 = ~n41998 & n41999;
  assign n42001 = ~pi219 & ~n41997;
  assign n42002 = ~n42000 & n42001;
  assign n42003 = n6294 & ~n39626;
  assign n42004 = ~n42002 & n42003;
  assign n42005 = ~pi57 & pi1151;
  assign n42006 = ~n41988 & n42005;
  assign n42007 = ~n42004 & n42006;
  assign n42008 = ~n41992 & ~n42007;
  assign n42009 = ~n41991 & n42008;
  assign n42010 = ~pi1152 & ~n42009;
  assign n42011 = n39999 & ~n40478;
  assign n42012 = ~n39529 & ~n41974;
  assign n42013 = ~pi214 & ~n42012;
  assign n42014 = pi212 & ~n42013;
  assign n42015 = ~n42011 & n42014;
  assign n42016 = n40374 & ~n41974;
  assign n42017 = n41353 & ~n42016;
  assign n42018 = ~n42015 & n42017;
  assign n42019 = ~pi1151 & ~n42018;
  assign n42020 = n40014 & n42019;
  assign n42021 = pi299 & ~n38700;
  assign n42022 = ~n10708 & n42021;
  assign n42023 = ~n38759 & ~n42022;
  assign n42024 = n39942 & ~n42023;
  assign n42025 = n40510 & ~n42024;
  assign n42026 = ~n40048 & ~n40157;
  assign n42027 = pi1151 & ~n42026;
  assign n42028 = ~n42025 & n42027;
  assign n42029 = n38764 & ~n42028;
  assign n42030 = ~n42020 & n42029;
  assign n42031 = pi1150 & ~n42030;
  assign n42032 = ~n42010 & n42031;
  assign n42033 = ~n38524 & n39965;
  assign n42034 = pi211 & n40571;
  assign n42035 = n38664 & ~n42033;
  assign n42036 = ~n42034 & n42035;
  assign n42037 = n10708 & n40572;
  assign n42038 = n38934 & ~n39577;
  assign n42039 = ~n42037 & ~n42038;
  assign n42040 = ~n42036 & n42039;
  assign n42041 = ~pi219 & ~n42040;
  assign n42042 = pi1151 & n39978;
  assign n42043 = ~n42041 & n42042;
  assign n42044 = ~n39598 & ~n42022;
  assign n42045 = n38702 & n39562;
  assign n42046 = ~n42044 & n42045;
  assign n42047 = n38705 & ~n42046;
  assign n42048 = ~n42043 & n42047;
  assign n42049 = n39920 & ~n42021;
  assign n42050 = pi212 & ~n42049;
  assign n42051 = ~n40560 & n42050;
  assign n42052 = ~pi212 & n39596;
  assign n42053 = ~pi219 & ~n42052;
  assign n42054 = ~n42016 & n42053;
  assign n42055 = ~n42051 & n42054;
  assign n42056 = n39539 & ~n40143;
  assign n42057 = ~n42055 & n42056;
  assign n42058 = ~pi1151 & n41690;
  assign n42059 = n38764 & ~n42046;
  assign n42060 = ~n42058 & n42059;
  assign n42061 = ~n42057 & n42060;
  assign n42062 = ~pi1150 & ~n42061;
  assign n42063 = ~n42048 & n42062;
  assign n42064 = ~n42032 & ~n42063;
  assign n42065 = pi213 & ~n42064;
  assign n42066 = ~pi209 & ~n42065;
  assign n42067 = ~n41973 & n42066;
  assign n42068 = ~n10654 & ~n38931;
  assign n42069 = n38522 & ~n39094;
  assign n42070 = ~pi207 & n39093;
  assign n42071 = pi207 & ~n38544;
  assign n42072 = ~n38929 & n42071;
  assign n42073 = pi208 & ~n42072;
  assign n42074 = ~n42070 & n42073;
  assign n42075 = ~n42069 & ~n42074;
  assign n42076 = pi211 & ~n42075;
  assign n42077 = pi214 & n42076;
  assign n42078 = ~n42068 & ~n42077;
  assign n42079 = ~pi212 & ~n42078;
  assign n42080 = ~pi219 & ~n42079;
  assign n42081 = ~pi211 & n42075;
  assign n42082 = ~n38967 & ~n42081;
  assign n42083 = pi214 & ~n42082;
  assign n42084 = ~pi211 & ~n38931;
  assign n42085 = ~pi214 & ~n42084;
  assign n42086 = ~n42076 & n42085;
  assign n42087 = pi212 & ~n42086;
  assign n42088 = ~n42083 & n42087;
  assign n42089 = n42080 & ~n42088;
  assign n42090 = n38933 & ~n42089;
  assign n42091 = n41581 & ~n42090;
  assign n42092 = ~n38931 & n38941;
  assign n42093 = ~n41871 & ~n42092;
  assign n42094 = ~n42091 & ~n42093;
  assign n42095 = pi214 & n38822;
  assign n42096 = n38883 & ~n42095;
  assign n42097 = ~pi219 & ~n42096;
  assign n42098 = pi214 & ~n38837;
  assign n42099 = ~pi214 & n38822;
  assign n42100 = pi212 & ~n42099;
  assign n42101 = ~n42098 & n42100;
  assign n42102 = n42097 & ~n42101;
  assign n42103 = ~po1038 & ~n38840;
  assign n42104 = ~n42102 & n42103;
  assign n42105 = n40349 & ~n42104;
  assign n42106 = ~n38837 & n39712;
  assign n42107 = ~n38835 & ~n39712;
  assign n42108 = ~po1038 & ~n42107;
  assign n42109 = ~n42106 & n42108;
  assign n42110 = n41657 & ~n42109;
  assign n42111 = pi1152 & ~n42110;
  assign n42112 = ~n42105 & n42111;
  assign n42113 = ~n42094 & ~n42112;
  assign n42114 = ~pi1150 & ~n42113;
  assign n42115 = ~n38290 & n42082;
  assign n42116 = pi219 & ~n38966;
  assign n42117 = ~n42115 & n42116;
  assign n42118 = ~po1038 & ~n42117;
  assign n42119 = pi214 & n42075;
  assign n42120 = n42087 & ~n42119;
  assign n42121 = n42080 & ~n42120;
  assign n42122 = n42118 & ~n42121;
  assign n42123 = n41585 & ~n42122;
  assign n42124 = pi212 & ~n42078;
  assign n42125 = ~pi212 & ~n38931;
  assign n42126 = ~pi219 & ~n42125;
  assign n42127 = ~n42124 & n42126;
  assign n42128 = n42118 & ~n42127;
  assign n42129 = n40421 & ~n42128;
  assign n42130 = ~pi1152 & ~n42129;
  assign n42131 = ~n42123 & n42130;
  assign n42132 = ~n38882 & ~n42098;
  assign n42133 = ~pi212 & ~n42132;
  assign n42134 = ~pi211 & n38835;
  assign n42135 = ~n38877 & ~n42134;
  assign n42136 = pi214 & ~n42135;
  assign n42137 = ~pi214 & n38837;
  assign n42138 = pi212 & ~n42136;
  assign n42139 = ~n42137 & n42138;
  assign n42140 = ~n42133 & ~n42139;
  assign n42141 = ~pi219 & ~n42140;
  assign n42142 = n38843 & ~n42141;
  assign n42143 = n41651 & ~n42142;
  assign n42144 = pi212 & ~n38822;
  assign n42145 = n42097 & ~n42144;
  assign n42146 = n38843 & ~n42145;
  assign n42147 = n40430 & ~n42146;
  assign n42148 = pi1152 & ~n42147;
  assign n42149 = ~n42143 & n42148;
  assign n42150 = ~n42131 & ~n42149;
  assign n42151 = pi1150 & ~n42150;
  assign n42152 = ~n42114 & ~n42151;
  assign n42153 = ~pi213 & ~n42152;
  assign n42154 = pi213 & n38939;
  assign n42155 = pi209 & ~n42154;
  assign n42156 = ~n42153 & n42155;
  assign n42157 = ~n42067 & ~n42156;
  assign n42158 = pi230 & ~n42157;
  assign n42159 = ~pi230 & ~pi249;
  assign po406 = ~n42158 & ~n42159;
  assign n42161 = n3277 & n11486;
  assign n42162 = ~n6252 & ~n42161;
  assign n42163 = ~pi75 & ~n42162;
  assign n42164 = n7323 & n8952;
  assign n42165 = ~n42163 & ~n42164;
  assign n42166 = ~pi87 & ~pi250;
  assign n42167 = n8867 & n42166;
  assign po407 = ~n42165 & n42167;
  assign n42169 = pi897 & n10793;
  assign n42170 = ~pi476 & n11419;
  assign n42171 = ~n42169 & ~n42170;
  assign n42172 = ~pi200 & pi1053;
  assign n42173 = pi200 & pi1039;
  assign n42174 = ~pi199 & ~n42172;
  assign n42175 = ~n42173 & n42174;
  assign n42176 = ~n42171 & ~n42175;
  assign n42177 = pi251 & n42171;
  assign po408 = n42176 | n42177;
  assign n42179 = ~n6206 & n11526;
  assign n42180 = ~pi979 & ~pi984;
  assign n42181 = pi1001 & n42180;
  assign n42182 = n6176 & n42181;
  assign n42183 = ~n6179 & n42182;
  assign n42184 = n6443 & n42183;
  assign n42185 = ~pi252 & ~n42184;
  assign n42186 = pi1092 & ~pi1093;
  assign n42187 = ~n42185 & n42186;
  assign n42188 = n6455 & ~n42187;
  assign n42189 = n6454 & n42187;
  assign n42190 = ~n42188 & ~n42189;
  assign n42191 = n6206 & n42190;
  assign n42192 = ~n42179 & ~n42191;
  assign n42193 = n6223 & ~n42192;
  assign n42194 = ~n6200 & n42190;
  assign n42195 = n6200 & n11526;
  assign n42196 = ~n42194 & ~n42195;
  assign n42197 = ~n6223 & ~n42196;
  assign n42198 = pi299 & ~n42193;
  assign n42199 = ~n42197 & n42198;
  assign n42200 = n6197 & ~n42192;
  assign n42201 = ~n6197 & ~n42196;
  assign n42202 = ~pi299 & ~n42200;
  assign n42203 = ~n42201 & n42202;
  assign n42204 = n10960 & ~n42199;
  assign n42205 = ~n42203 & n42204;
  assign n42206 = ~n10960 & n11526;
  assign n42207 = ~n8856 & ~n42206;
  assign n42208 = ~n42205 & n42207;
  assign n42209 = n10959 & n42182;
  assign n42210 = n21085 & n42209;
  assign n42211 = n6183 & n42210;
  assign n42212 = ~n38264 & n42211;
  assign n42213 = n6443 & n42212;
  assign n42214 = ~pi252 & ~n42213;
  assign n42215 = ~pi57 & pi1092;
  assign n42216 = ~n42214 & n42215;
  assign n42217 = pi57 & n11525;
  assign n42218 = n8856 & ~n42217;
  assign n42219 = ~n42216 & n42218;
  assign po409 = ~n42208 & ~n42219;
  assign n42221 = ~n13025 & ~n38384;
  assign n42222 = ~n38484 & n42221;
  assign n42223 = ~po1038 & n42222;
  assign n42224 = ~pi211 & po1038;
  assign n42225 = pi219 & n42224;
  assign n42226 = ~n42223 & ~n42225;
  assign n42227 = pi1153 & ~n42226;
  assign n42228 = ~pi1151 & ~n42227;
  assign n42229 = n10709 & n38466;
  assign n42230 = pi211 & ~n38426;
  assign n42231 = ~n42229 & ~n42230;
  assign n42232 = ~n38419 & ~n38432;
  assign n42233 = n38395 & ~n42232;
  assign n42234 = ~po1038 & ~n42233;
  assign n42235 = n42231 & n42234;
  assign n42236 = ~n11421 & n39209;
  assign n42237 = pi1151 & ~n42236;
  assign n42238 = ~n42235 & n42237;
  assign n42239 = ~n42228 & ~n42238;
  assign n42240 = ~pi1152 & ~n42239;
  assign n42241 = n38395 & n39655;
  assign n42242 = ~pi1151 & ~n11422;
  assign n42243 = ~n38471 & n42242;
  assign n42244 = ~n42241 & n42243;
  assign n42245 = ~n38424 & ~n39762;
  assign n42246 = pi1153 & ~n42245;
  assign n42247 = ~n11348 & ~n38384;
  assign n42248 = pi1151 & n42247;
  assign n42249 = ~n42246 & n42248;
  assign n42250 = ~po1038 & ~n42249;
  assign n42251 = ~n42244 & n42250;
  assign n42252 = ~pi1151 & n10709;
  assign n42253 = n39209 & ~n42252;
  assign n42254 = pi1152 & ~n42253;
  assign n42255 = ~n42251 & n42254;
  assign n42256 = ~n42240 & ~n42255;
  assign n42257 = pi230 & ~n42256;
  assign n42258 = n40732 & n40782;
  assign n42259 = pi1153 & ~n42258;
  assign n42260 = ~pi1153 & ~n40806;
  assign n42261 = ~pi219 & ~n42260;
  assign n42262 = ~n42259 & n42261;
  assign n42263 = ~n40737 & ~n40751;
  assign n42264 = ~pi211 & n40731;
  assign n42265 = n42263 & ~n42264;
  assign n42266 = ~n40730 & n40771;
  assign n42267 = n42265 & n42266;
  assign n42268 = pi1153 & ~n42267;
  assign n42269 = ~pi1153 & ~n40882;
  assign n42270 = pi219 & ~n42269;
  assign n42271 = ~n42268 & n42270;
  assign n42272 = pi253 & ~n42262;
  assign n42273 = ~n42271 & n42272;
  assign n42274 = ~n40742 & n40882;
  assign n42275 = ~pi211 & n42274;
  assign n42276 = ~n40744 & ~n42275;
  assign n42277 = pi1153 & ~n42276;
  assign n42278 = ~n40877 & ~n42277;
  assign n42279 = pi219 & n42278;
  assign n42280 = pi1153 & n40752;
  assign n42281 = ~pi1153 & n40804;
  assign n42282 = ~pi219 & ~n42281;
  assign n42283 = ~n42280 & n42282;
  assign n42284 = ~pi253 & ~n42283;
  assign n42285 = ~n42279 & n42284;
  assign n42286 = ~n42273 & ~n42285;
  assign n42287 = ~po1038 & ~n42286;
  assign n42288 = ~pi219 & ~n40724;
  assign n42289 = ~pi211 & ~n40722;
  assign n42290 = n42288 & ~n42289;
  assign n42291 = ~pi219 & ~n42290;
  assign n42292 = po1038 & n42291;
  assign n42293 = ~n40713 & n42292;
  assign n42294 = pi219 & pi1091;
  assign n42295 = ~n38376 & n42294;
  assign n42296 = ~n40740 & ~n42295;
  assign n42297 = ~n42288 & n42296;
  assign n42298 = pi253 & ~n42297;
  assign n42299 = ~pi211 & ~n40713;
  assign n42300 = pi211 & n40740;
  assign n42301 = pi219 & ~n42300;
  assign n42302 = ~n42299 & n42301;
  assign n42303 = ~pi219 & ~n40722;
  assign n42304 = ~n42295 & ~n42303;
  assign n42305 = ~n42302 & n42304;
  assign n42306 = ~pi253 & ~n42305;
  assign n42307 = po1038 & ~n42298;
  assign n42308 = ~n42306 & n42307;
  assign n42309 = pi1151 & ~n42293;
  assign n42310 = ~n42308 & n42309;
  assign n42311 = ~n42287 & n42310;
  assign n42312 = ~n40751 & ~n40759;
  assign n42313 = ~pi1153 & ~n42312;
  assign n42314 = ~n40743 & n42265;
  assign n42315 = ~n42313 & n42314;
  assign n42316 = ~pi219 & ~n42315;
  assign n42317 = pi219 & n40737;
  assign n42318 = ~n42316 & ~n42317;
  assign n42319 = ~n42279 & n42318;
  assign n42320 = ~pi253 & ~n42319;
  assign n42321 = ~n40732 & ~n42275;
  assign n42322 = n42288 & ~n42321;
  assign n42323 = ~n40760 & ~n42313;
  assign n42324 = n42322 & ~n42323;
  assign n42325 = pi219 & n40837;
  assign n42326 = ~n40849 & n42268;
  assign n42327 = n42325 & ~n42326;
  assign n42328 = ~n42324 & ~n42327;
  assign n42329 = pi253 & ~n42328;
  assign n42330 = ~po1038 & ~n42329;
  assign n42331 = ~n42320 & n42330;
  assign n42332 = ~pi1151 & ~n42331;
  assign n42333 = ~n42311 & ~n42332;
  assign n42334 = ~n42299 & n42303;
  assign n42335 = n42288 & ~n42334;
  assign n42336 = pi219 & ~n40713;
  assign n42337 = po1038 & ~n42336;
  assign n42338 = ~n42335 & n42337;
  assign n42339 = ~n40713 & n42338;
  assign n42340 = ~n42308 & ~n42339;
  assign n42341 = ~n42333 & n42340;
  assign n42342 = pi1152 & ~n42341;
  assign n42343 = pi219 & ~n42278;
  assign n42344 = ~n42283 & n42322;
  assign n42345 = ~n42343 & ~n42344;
  assign n42346 = ~n40742 & ~n42345;
  assign n42347 = ~pi253 & ~n42346;
  assign n42348 = pi1153 & ~n40782;
  assign n42349 = n42265 & n42288;
  assign n42350 = ~n42348 & n42349;
  assign n42351 = ~n40839 & ~n42267;
  assign n42352 = pi1153 & n42351;
  assign n42353 = ~pi1153 & ~n40888;
  assign n42354 = pi219 & ~n42353;
  assign n42355 = ~n42352 & n42354;
  assign n42356 = ~n42350 & ~n42355;
  assign n42357 = pi253 & ~n42356;
  assign n42358 = ~po1038 & ~n42357;
  assign n42359 = ~n42347 & n42358;
  assign n42360 = n42310 & ~n42359;
  assign n42361 = ~n40729 & n42343;
  assign n42362 = ~pi1153 & ~n40774;
  assign n42363 = ~n40742 & ~n42362;
  assign n42364 = ~pi219 & n40806;
  assign n42365 = n42363 & n42364;
  assign n42366 = ~pi253 & ~n42365;
  assign n42367 = ~n42361 & n42366;
  assign n42368 = ~n40849 & ~n42267;
  assign n42369 = ~pi1091 & ~n40877;
  assign n42370 = ~pi1153 & ~n42369;
  assign n42371 = ~pi219 & n42312;
  assign n42372 = ~n42370 & ~n42371;
  assign n42373 = n42368 & n42372;
  assign n42374 = pi253 & ~n42373;
  assign n42375 = ~po1038 & ~n42374;
  assign n42376 = ~n42367 & n42375;
  assign n42377 = ~pi1151 & ~n42308;
  assign n42378 = ~n42376 & n42377;
  assign n42379 = ~pi1152 & ~n42378;
  assign n42380 = ~n42360 & n42379;
  assign n42381 = ~n42342 & ~n42380;
  assign n42382 = n40997 & ~n42381;
  assign n42383 = pi1091 & ~n42231;
  assign n42384 = ~pi1153 & ~n40907;
  assign n42385 = pi1153 & ~n40936;
  assign n42386 = n38395 & ~n42385;
  assign n42387 = ~n42384 & n42386;
  assign n42388 = ~n42383 & ~n42387;
  assign n42389 = pi253 & ~n42388;
  assign n42390 = ~n13028 & ~n42246;
  assign n42391 = pi1091 & ~n42390;
  assign n42392 = ~pi253 & ~n42391;
  assign n42393 = ~po1038 & ~n42392;
  assign n42394 = ~n42389 & n42393;
  assign n42395 = ~pi253 & ~pi1091;
  assign n42396 = po1038 & ~n42395;
  assign n42397 = pi211 & pi1091;
  assign n42398 = pi1091 & ~pi1153;
  assign n42399 = pi219 & n42398;
  assign n42400 = ~n42397 & ~n42399;
  assign n42401 = n42396 & n42400;
  assign n42402 = pi1151 & ~n42401;
  assign n42403 = ~n42394 & n42402;
  assign n42404 = ~n42295 & n42396;
  assign n42405 = pi219 & n42404;
  assign n42406 = pi1091 & pi1153;
  assign n42407 = n42223 & n42406;
  assign n42408 = pi253 & ~pi1091;
  assign n42409 = ~pi1151 & ~n42408;
  assign n42410 = ~n42407 & n42409;
  assign n42411 = ~n42405 & n42410;
  assign n42412 = ~n42403 & ~n42411;
  assign n42413 = ~pi1152 & ~n42412;
  assign n42414 = ~pi1153 & ~n40942;
  assign n42415 = ~n38409 & n40903;
  assign n42416 = pi1153 & ~n42415;
  assign n42417 = n38395 & ~n42416;
  assign n42418 = ~n42414 & n42417;
  assign n42419 = n11421 & n40903;
  assign n42420 = ~n38471 & n42419;
  assign n42421 = pi253 & ~n42420;
  assign n42422 = ~n42418 & n42421;
  assign n42423 = pi1091 & n39655;
  assign n42424 = pi1091 & n38432;
  assign n42425 = n38827 & n42424;
  assign n42426 = n38395 & ~n42425;
  assign n42427 = ~n42423 & n42426;
  assign n42428 = pi1091 & n38471;
  assign n42429 = pi211 & ~n40955;
  assign n42430 = ~n42428 & n42429;
  assign n42431 = ~pi253 & ~n42427;
  assign n42432 = ~n42430 & n42431;
  assign n42433 = ~n42422 & ~n42432;
  assign n42434 = ~n11421 & ~n38395;
  assign n42435 = ~n42408 & n42434;
  assign n42436 = ~n42428 & n42435;
  assign n42437 = n39562 & ~n42436;
  assign n42438 = ~n42433 & n42437;
  assign n42439 = n42245 & ~n42408;
  assign n42440 = ~n42398 & ~n42439;
  assign n42441 = n42247 & ~n42440;
  assign n42442 = ~po1038 & ~n42395;
  assign n42443 = ~n42441 & n42442;
  assign n42444 = ~n42404 & ~n42443;
  assign n42445 = pi1151 & ~n42444;
  assign n42446 = ~pi211 & pi1091;
  assign n42447 = ~pi219 & n42446;
  assign n42448 = n42404 & ~n42447;
  assign n42449 = pi1152 & ~n42448;
  assign n42450 = ~n42445 & n42449;
  assign n42451 = ~n42438 & n42450;
  assign n42452 = ~n40997 & ~n42451;
  assign n42453 = ~n42413 & n42452;
  assign n42454 = ~pi230 & ~n42453;
  assign n42455 = ~n42382 & n42454;
  assign po410 = ~n42257 & ~n42455;
  assign n42457 = pi1154 & n38859;
  assign n42458 = ~n38891 & ~n42457;
  assign n42459 = n11421 & ~n42458;
  assign n42460 = pi299 & n38395;
  assign n42461 = ~n11421 & n38828;
  assign n42462 = ~n42460 & ~n42461;
  assign n42463 = ~n38808 & ~n42462;
  assign n42464 = ~n42459 & ~n42463;
  assign n42465 = ~po1038 & ~n42464;
  assign n42466 = ~pi219 & ~n38699;
  assign n42467 = ~n39017 & ~n42466;
  assign n42468 = po1038 & n42467;
  assign n42469 = ~pi1152 & ~n42468;
  assign n42470 = ~n42465 & n42469;
  assign n42471 = ~n38416 & ~n38858;
  assign n42472 = n38360 & ~n42471;
  assign n42473 = ~n38811 & ~n38925;
  assign n42474 = ~n42472 & ~n42473;
  assign n42475 = pi219 & ~n42474;
  assign n42476 = ~pi200 & pi1154;
  assign n42477 = n11358 & ~n42476;
  assign n42478 = n38858 & ~n39762;
  assign n42479 = ~n42477 & ~n42478;
  assign n42480 = ~pi219 & ~n42479;
  assign n42481 = ~po1038 & ~n42480;
  assign n42482 = ~n42475 & n42481;
  assign n42483 = n11421 & ~n38699;
  assign n42484 = n39909 & ~n42483;
  assign n42485 = pi1152 & ~n42484;
  assign n42486 = ~n42482 & n42485;
  assign n42487 = ~n42470 & ~n42486;
  assign n42488 = pi230 & ~n42487;
  assign n42489 = ~pi1153 & n42315;
  assign n42490 = ~n40806 & ~n42489;
  assign n42491 = ~pi1154 & ~n42490;
  assign n42492 = pi1154 & ~n40736;
  assign n42493 = n42265 & n42492;
  assign n42494 = ~n42259 & n42493;
  assign n42495 = pi254 & ~n42494;
  assign n42496 = ~n42491 & n42495;
  assign n42497 = ~n40743 & n40888;
  assign n42498 = pi1154 & n42497;
  assign n42499 = ~n40804 & ~n42498;
  assign n42500 = ~pi1153 & ~n42264;
  assign n42501 = ~n40777 & n42500;
  assign n42502 = ~pi254 & ~n42501;
  assign n42503 = ~n42499 & n42502;
  assign n42504 = ~n42496 & ~n42503;
  assign n42505 = ~pi219 & ~n42504;
  assign n42506 = pi1154 & ~n42268;
  assign n42507 = ~n42351 & n42506;
  assign n42508 = pi1153 & ~n40882;
  assign n42509 = ~pi1154 & ~n42353;
  assign n42510 = ~n42508 & n42509;
  assign n42511 = pi254 & ~n42510;
  assign n42512 = ~n42507 & n42511;
  assign n42513 = ~n42269 & n42497;
  assign n42514 = n38374 & ~n42513;
  assign n42515 = ~n40714 & n42514;
  assign n42516 = ~pi1153 & ~n40791;
  assign n42517 = n40879 & ~n42516;
  assign n42518 = ~pi1154 & ~n42517;
  assign n42519 = ~n40742 & n40877;
  assign n42520 = n42518 & ~n42519;
  assign n42521 = pi1153 & n40744;
  assign n42522 = n38360 & ~n40866;
  assign n42523 = ~n42521 & n42522;
  assign n42524 = ~pi254 & ~n42523;
  assign n42525 = ~n42515 & n42524;
  assign n42526 = ~n42520 & n42525;
  assign n42527 = ~n42512 & ~n42526;
  assign n42528 = pi219 & ~n42527;
  assign n42529 = pi253 & ~n42528;
  assign n42530 = ~n42505 & n42529;
  assign n42531 = pi1153 & ~n40922;
  assign n42532 = ~pi1154 & ~n42531;
  assign n42533 = ~pi211 & n38465;
  assign n42534 = ~n42384 & n42532;
  assign n42535 = ~n42533 & n42534;
  assign n42536 = pi1091 & n38360;
  assign n42537 = ~n38424 & n42536;
  assign n42538 = ~n38903 & n42537;
  assign n42539 = ~n42535 & ~n42538;
  assign n42540 = ~pi219 & ~n42539;
  assign n42541 = pi1154 & n42446;
  assign n42542 = ~n42294 & ~n42541;
  assign n42543 = ~n42474 & ~n42542;
  assign n42544 = ~n42540 & ~n42543;
  assign n42545 = pi254 & ~n42544;
  assign n42546 = ~pi254 & ~pi1091;
  assign n42547 = pi1154 & ~n42245;
  assign n42548 = pi219 & ~n38925;
  assign n42549 = ~n42547 & n42548;
  assign n42550 = ~n42480 & ~n42549;
  assign n42551 = ~pi254 & ~n42550;
  assign n42552 = ~n42546 & ~n42551;
  assign n42553 = ~n42545 & n42552;
  assign n42554 = ~pi253 & ~n42553;
  assign n42555 = ~po1038 & ~n42554;
  assign n42556 = ~n42530 & n42555;
  assign n42557 = ~pi211 & ~n40738;
  assign n42558 = n42336 & ~n42557;
  assign n42559 = ~pi219 & n40722;
  assign n42560 = ~n42558 & ~n42559;
  assign n42561 = pi1091 & n39017;
  assign n42562 = n11421 & n42398;
  assign n42563 = pi254 & ~n42562;
  assign n42564 = ~n42561 & n42563;
  assign n42565 = n42560 & n42564;
  assign n42566 = n42334 & ~n42406;
  assign n42567 = ~pi254 & ~n42561;
  assign n42568 = ~n42302 & n42567;
  assign n42569 = ~n42566 & n42568;
  assign n42570 = pi253 & ~n42565;
  assign n42571 = ~n42569 & n42570;
  assign n42572 = pi1091 & ~n42467;
  assign n42573 = po1038 & ~n42546;
  assign n42574 = ~n42572 & n42573;
  assign n42575 = po1038 & n42447;
  assign n42576 = ~n42574 & ~n42575;
  assign n42577 = pi253 & po1038;
  assign n42578 = n42576 & ~n42577;
  assign n42579 = ~n42571 & ~n42578;
  assign n42580 = pi1152 & ~n42579;
  assign n42581 = ~n42556 & n42580;
  assign n42582 = ~pi1154 & ~n40870;
  assign n42583 = ~pi1154 & ~n42582;
  assign n42584 = ~pi1153 & n40771;
  assign n42585 = ~n42266 & ~n42584;
  assign n42586 = ~n42583 & n42585;
  assign n42587 = n38374 & ~n40849;
  assign n42588 = pi219 & ~n42587;
  assign n42589 = ~n42586 & n42588;
  assign n42590 = n42321 & ~n42584;
  assign n42591 = pi1154 & n40759;
  assign n42592 = ~pi219 & ~n42591;
  assign n42593 = ~n42590 & n42592;
  assign n42594 = ~n42589 & ~n42593;
  assign n42595 = pi254 & ~n42594;
  assign n42596 = n40745 & ~n42269;
  assign n42597 = n38360 & ~n42596;
  assign n42598 = pi219 & ~n42514;
  assign n42599 = ~n42518 & n42598;
  assign n42600 = ~n42597 & n42599;
  assign n42601 = ~n40736 & n40804;
  assign n42602 = ~n42362 & n42601;
  assign n42603 = ~pi1154 & ~n42602;
  assign n42604 = ~n40742 & n40806;
  assign n42605 = pi1154 & ~n42604;
  assign n42606 = ~n42602 & n42605;
  assign n42607 = pi1154 & n40737;
  assign n42608 = ~n40731 & ~n42607;
  assign n42609 = ~pi211 & ~n42608;
  assign n42610 = ~pi219 & ~n42609;
  assign n42611 = ~n42603 & n42610;
  assign n42612 = ~n42606 & n42611;
  assign n42613 = ~pi254 & ~n42612;
  assign n42614 = ~n42600 & n42613;
  assign n42615 = ~n42595 & ~n42614;
  assign n42616 = pi253 & ~n42615;
  assign n42617 = n40910 & n42398;
  assign n42618 = ~n42423 & ~n42617;
  assign n42619 = pi211 & ~n42532;
  assign n42620 = ~n42618 & n42619;
  assign n42621 = pi1091 & n38828;
  assign n42622 = pi1154 & ~n42621;
  assign n42623 = n11420 & n42406;
  assign n42624 = ~pi1154 & ~n42623;
  assign n42625 = ~pi211 & ~n42624;
  assign n42626 = ~n42622 & n42625;
  assign n42627 = ~n42620 & ~n42626;
  assign n42628 = ~pi219 & ~n42627;
  assign n42629 = pi211 & n42622;
  assign n42630 = pi1091 & n39510;
  assign n42631 = n38374 & ~n42630;
  assign n42632 = ~n42423 & n42631;
  assign n42633 = pi219 & ~n42624;
  assign n42634 = ~n42632 & n42633;
  assign n42635 = ~n42629 & n42634;
  assign n42636 = ~n42628 & ~n42635;
  assign n42637 = ~pi254 & ~n42636;
  assign n42638 = pi1091 & ~n11421;
  assign n42639 = ~n38807 & n42638;
  assign n42640 = ~pi1154 & ~n42639;
  assign n42641 = ~pi1153 & ~n40911;
  assign n42642 = ~n42416 & ~n42641;
  assign n42643 = pi1091 & ~n38410;
  assign n42644 = ~n42642 & ~n42643;
  assign n42645 = n42434 & ~n42644;
  assign n42646 = n40958 & n42417;
  assign n42647 = pi1154 & ~n42646;
  assign n42648 = ~n42645 & n42647;
  assign n42649 = ~n42640 & ~n42648;
  assign n42650 = pi1091 & ~pi1154;
  assign n42651 = n38540 & n42650;
  assign n42652 = ~n42642 & ~n42651;
  assign n42653 = n11421 & ~n42652;
  assign n42654 = pi254 & ~n42653;
  assign n42655 = ~n42649 & n42654;
  assign n42656 = ~n42637 & ~n42655;
  assign n42657 = ~pi253 & n42656;
  assign n42658 = ~po1038 & ~n42657;
  assign n42659 = ~n42616 & n42658;
  assign n42660 = ~n42574 & ~n42577;
  assign n42661 = ~n42335 & n42565;
  assign n42662 = ~n42291 & n42569;
  assign n42663 = pi253 & ~n42661;
  assign n42664 = ~n42662 & n42663;
  assign n42665 = ~n42660 & ~n42664;
  assign n42666 = ~pi1152 & ~n42665;
  assign n42667 = ~n42659 & n42666;
  assign n42668 = n40997 & ~n42667;
  assign n42669 = ~n42581 & n42668;
  assign n42670 = ~po1038 & ~n42656;
  assign n42671 = ~pi1152 & ~n42574;
  assign n42672 = ~n42670 & n42671;
  assign n42673 = ~po1038 & n42553;
  assign n42674 = pi1152 & n42576;
  assign n42675 = ~n42673 & n42674;
  assign n42676 = ~n40997 & ~n42675;
  assign n42677 = ~n42672 & n42676;
  assign n42678 = ~pi230 & ~n42677;
  assign n42679 = ~n42669 & n42678;
  assign po411 = ~n42488 & ~n42679;
  assign n42681 = ~pi200 & pi1049;
  assign n42682 = pi200 & pi1036;
  assign n42683 = ~n42681 & ~n42682;
  assign n42684 = ~n42171 & n42683;
  assign n42685 = ~pi255 & n42171;
  assign po412 = ~n42684 & ~n42685;
  assign n42687 = ~pi200 & pi1048;
  assign n42688 = pi200 & pi1070;
  assign n42689 = ~n42687 & ~n42688;
  assign n42690 = ~n42171 & n42689;
  assign n42691 = ~pi256 & n42171;
  assign po413 = ~n42690 & ~n42691;
  assign n42693 = ~pi200 & pi1084;
  assign n42694 = pi200 & pi1065;
  assign n42695 = ~n42693 & ~n42694;
  assign n42696 = ~n42171 & n42695;
  assign n42697 = ~pi257 & n42171;
  assign po414 = ~n42696 & ~n42697;
  assign n42699 = ~pi200 & pi1072;
  assign n42700 = pi200 & pi1062;
  assign n42701 = ~n42699 & ~n42700;
  assign n42702 = ~n42171 & n42701;
  assign n42703 = ~pi258 & n42171;
  assign po415 = ~n42702 & ~n42703;
  assign n42705 = ~pi200 & pi1059;
  assign n42706 = pi200 & pi1069;
  assign n42707 = ~n42705 & ~n42706;
  assign n42708 = ~n42171 & n42707;
  assign n42709 = ~pi259 & n42171;
  assign po416 = ~n42708 & ~n42709;
  assign n42711 = ~pi200 & pi1044;
  assign n42712 = pi200 & pi1067;
  assign n42713 = ~pi199 & ~n42711;
  assign n42714 = ~n42712 & n42713;
  assign n42715 = ~n42171 & ~n42714;
  assign n42716 = pi260 & n42171;
  assign po417 = n42715 | n42716;
  assign n42718 = ~pi200 & pi1037;
  assign n42719 = pi200 & pi1040;
  assign n42720 = ~pi199 & ~n42718;
  assign n42721 = ~n42719 & n42720;
  assign n42722 = ~n42171 & ~n42721;
  assign n42723 = pi261 & n42171;
  assign po418 = n42722 | n42723;
  assign n42725 = pi1093 & pi1142;
  assign n42726 = ~pi262 & ~pi1093;
  assign n42727 = ~n42725 & ~n42726;
  assign n42728 = ~pi228 & ~n42727;
  assign n42729 = ~pi123 & ~pi1142;
  assign n42730 = pi123 & pi262;
  assign n42731 = pi228 & ~n42729;
  assign n42732 = ~n42730 & n42731;
  assign n42733 = ~n42728 & ~n42732;
  assign n42734 = ~pi228 & ~pi1093;
  assign n42735 = pi123 & pi228;
  assign n42736 = ~n42734 & ~n42735;
  assign n42737 = ~pi262 & ~n42736;
  assign n42738 = ~n40601 & ~n42737;
  assign n42739 = pi199 & n42736;
  assign n42740 = n38319 & ~n42739;
  assign n42741 = n42738 & ~n42740;
  assign n42742 = ~n42733 & ~n42741;
  assign n42743 = ~pi207 & n42737;
  assign n42744 = ~pi208 & ~n42743;
  assign n42745 = ~n40601 & ~n42744;
  assign n42746 = ~n42742 & ~n42745;
  assign n42747 = pi299 & ~n42738;
  assign n42748 = ~n39923 & n42736;
  assign n42749 = ~pi299 & ~n42748;
  assign n42750 = ~n42733 & n42749;
  assign n42751 = pi208 & ~n42750;
  assign n42752 = ~n42747 & n42751;
  assign n42753 = ~po1038 & ~n42752;
  assign n42754 = ~n42746 & n42753;
  assign n42755 = ~n39720 & n42736;
  assign n42756 = po1038 & ~n42733;
  assign n42757 = ~n42755 & n42756;
  assign po419 = n42754 | n42757;
  assign n42759 = pi1154 & ~n40753;
  assign n42760 = ~n40801 & n42759;
  assign n42761 = ~pi1154 & ~n40775;
  assign n42762 = pi1155 & n42601;
  assign n42763 = n42761 & ~n42762;
  assign n42764 = ~n40822 & n42759;
  assign n42765 = ~pi1156 & ~n42591;
  assign n42766 = ~n42764 & n42765;
  assign n42767 = ~pi1156 & ~n42766;
  assign n42768 = ~n42763 & ~n42767;
  assign n42769 = pi1156 & n42604;
  assign n42770 = ~n42768 & ~n42769;
  assign n42771 = ~n42760 & ~n42770;
  assign n42772 = pi211 & ~n42771;
  assign n42773 = n40755 & ~n40803;
  assign n42774 = pi1155 & n42773;
  assign n42775 = n42761 & ~n42774;
  assign n42776 = n42766 & ~n42775;
  assign n42777 = ~n42604 & n42775;
  assign n42778 = pi1156 & ~n42777;
  assign n42779 = ~n42764 & n42778;
  assign n42780 = ~pi211 & ~n42779;
  assign n42781 = ~n42776 & n42780;
  assign n42782 = ~pi219 & ~n42781;
  assign n42783 = ~n42772 & n42782;
  assign n42784 = ~n40747 & ~n40878;
  assign n42785 = ~n40745 & ~n42607;
  assign n42786 = ~n42784 & ~n42785;
  assign n42787 = ~n40803 & n42786;
  assign n42788 = ~pi1156 & ~n42787;
  assign n42789 = pi1155 & ~n42497;
  assign n42790 = ~pi1155 & ~n42274;
  assign n42791 = ~pi1154 & ~n42789;
  assign n42792 = ~n42790 & n42791;
  assign n42793 = pi1154 & ~n42784;
  assign n42794 = n38355 & ~n42793;
  assign n42795 = ~n42792 & n42794;
  assign n42796 = n38366 & ~n42786;
  assign n42797 = pi219 & ~n42795;
  assign n42798 = ~n42796 & n42797;
  assign n42799 = ~n42788 & n42798;
  assign n42800 = pi263 & ~n42799;
  assign n42801 = ~n42783 & n42800;
  assign n42802 = ~pi1155 & n42369;
  assign n42803 = ~n40804 & n42802;
  assign n42804 = pi1155 & ~n40732;
  assign n42805 = ~pi1154 & ~n42804;
  assign n42806 = ~n42803 & n42805;
  assign n42807 = ~pi1156 & ~n42806;
  assign n42808 = pi1155 & ~n40806;
  assign n42809 = pi1154 & ~n42808;
  assign n42810 = n40763 & n42809;
  assign n42811 = pi1155 & ~n40837;
  assign n42812 = ~pi1154 & ~n42811;
  assign n42813 = ~n42802 & n42812;
  assign n42814 = ~n42810 & ~n42813;
  assign n42815 = n42807 & n42814;
  assign n42816 = ~pi1155 & n40771;
  assign n42817 = ~n40731 & n40760;
  assign n42818 = ~n42816 & ~n42817;
  assign n42819 = ~pi1154 & ~n42818;
  assign n42820 = pi1156 & ~n42819;
  assign n42821 = n40771 & n42812;
  assign n42822 = ~n40734 & n42810;
  assign n42823 = ~n42821 & ~n42822;
  assign n42824 = n42820 & n42823;
  assign n42825 = ~pi211 & ~n42815;
  assign n42826 = ~n42824 & n42825;
  assign n42827 = n40782 & n42809;
  assign n42828 = n42820 & ~n42827;
  assign n42829 = n42263 & n42809;
  assign n42830 = n42807 & ~n42829;
  assign n42831 = pi211 & ~n42828;
  assign n42832 = ~n42830 & n42831;
  assign n42833 = ~pi219 & ~n42826;
  assign n42834 = ~n42832 & n42833;
  assign n42835 = pi1155 & n40730;
  assign n42836 = pi1154 & n40888;
  assign n42837 = ~n42835 & n42836;
  assign n42838 = ~n40736 & n42837;
  assign n42839 = ~n42821 & ~n42838;
  assign n42840 = n38366 & ~n42839;
  assign n42841 = ~n42813 & ~n42837;
  assign n42842 = ~pi1156 & ~n42841;
  assign n42843 = ~pi1154 & n40877;
  assign n42844 = ~n40839 & ~n42843;
  assign n42845 = n38355 & ~n42835;
  assign n42846 = ~n42844 & n42845;
  assign n42847 = pi219 & ~n42846;
  assign n42848 = ~n42840 & n42847;
  assign n42849 = ~n42842 & n42848;
  assign n42850 = ~pi263 & ~n42849;
  assign n42851 = ~n42834 & n42850;
  assign n42852 = n40835 & ~n42851;
  assign n42853 = ~n42801 & n42852;
  assign n42854 = pi1155 & ~n38867;
  assign n42855 = n40936 & ~n42854;
  assign n42856 = ~pi1154 & n42643;
  assign n42857 = ~n42855 & ~n42856;
  assign n42858 = ~n40955 & n42857;
  assign n42859 = n38366 & ~n42858;
  assign n42860 = ~pi1154 & ~n38505;
  assign n42861 = n38432 & ~n38433;
  assign n42862 = pi1154 & ~n42861;
  assign n42863 = pi1091 & n38355;
  assign n42864 = ~n42862 & n42863;
  assign n42865 = ~n42860 & n42864;
  assign n42866 = ~n40907 & ~n42650;
  assign n42867 = ~pi1156 & ~n38434;
  assign n42868 = ~n42866 & n42867;
  assign n42869 = pi219 & ~n42868;
  assign n42870 = ~n42865 & n42869;
  assign n42871 = ~n42859 & n42870;
  assign n42872 = ~pi211 & ~n42857;
  assign n42873 = n38424 & ~n38980;
  assign n42874 = n42397 & ~n42873;
  assign n42875 = ~n38541 & n42874;
  assign n42876 = ~n42872 & ~n42875;
  assign n42877 = pi1156 & ~n42876;
  assign n42878 = ~n38541 & ~n42866;
  assign n42879 = pi211 & n42878;
  assign n42880 = ~n38434 & ~n38849;
  assign n42881 = n42446 & n42880;
  assign n42882 = ~n42879 & ~n42881;
  assign n42883 = ~pi1156 & ~n42882;
  assign n42884 = ~pi219 & ~n42883;
  assign n42885 = ~n42877 & n42884;
  assign n42886 = ~n42871 & ~n42885;
  assign n42887 = ~pi263 & ~n42886;
  assign n42888 = ~n38515 & n42860;
  assign n42889 = ~n38424 & ~n38470;
  assign n42890 = pi1154 & ~n42889;
  assign n42891 = pi1156 & ~n42890;
  assign n42892 = ~n42888 & n42891;
  assign n42893 = ~pi1156 & n42878;
  assign n42894 = pi211 & ~n42893;
  assign n42895 = ~n42892 & n42894;
  assign n42896 = ~n38439 & n39402;
  assign n42897 = ~n38849 & ~n42896;
  assign n42898 = ~pi211 & ~n42897;
  assign n42899 = ~pi219 & ~n42898;
  assign n42900 = ~n42895 & n42899;
  assign n42901 = pi1154 & ~n38436;
  assign n42902 = pi1156 & ~n42901;
  assign n42903 = ~pi299 & ~n42902;
  assign n42904 = ~pi1154 & n38437;
  assign n42905 = ~n39762 & ~n42904;
  assign n42906 = ~n42903 & n42905;
  assign n42907 = pi1156 & ~n42906;
  assign n42908 = ~n42880 & n42903;
  assign n42909 = pi219 & ~n42908;
  assign n42910 = ~n42907 & n42909;
  assign n42911 = pi263 & pi1091;
  assign n42912 = ~n42910 & n42911;
  assign n42913 = ~n42900 & n42912;
  assign n42914 = ~n42887 & ~n42913;
  assign n42915 = ~n40835 & ~n42914;
  assign n42916 = ~po1038 & ~n42915;
  assign n42917 = ~n42853 & n42916;
  assign n42918 = pi211 & n40713;
  assign n42919 = ~pi211 & ~n42650;
  assign n42920 = ~n38356 & ~n42919;
  assign n42921 = ~n42918 & n42920;
  assign n42922 = ~n40722 & ~n42921;
  assign n42923 = ~pi219 & ~n42922;
  assign n42924 = ~pi263 & ~n42558;
  assign n42925 = ~n42923 & n42924;
  assign n42926 = ~n38356 & ~n42541;
  assign n42927 = ~n42918 & ~n42926;
  assign n42928 = n42303 & ~n42927;
  assign n42929 = pi263 & ~n42302;
  assign n42930 = ~n42928 & n42929;
  assign n42931 = ~n42925 & ~n42930;
  assign n42932 = pi219 & ~n38355;
  assign n42933 = pi1091 & n42932;
  assign n42934 = n40835 & ~n42933;
  assign n42935 = ~n42931 & n42934;
  assign n42936 = ~pi219 & ~n38356;
  assign n42937 = ~n38374 & n42936;
  assign n42938 = ~n42932 & ~n42937;
  assign n42939 = pi1091 & ~n42938;
  assign n42940 = pi263 & ~pi1091;
  assign n42941 = ~n42939 & ~n42940;
  assign n42942 = ~n40835 & n42941;
  assign n42943 = po1038 & ~n42942;
  assign n42944 = ~n42935 & n42943;
  assign n42945 = n40997 & ~n42944;
  assign n42946 = ~n42917 & n42945;
  assign n42947 = ~po1038 & n42914;
  assign n42948 = po1038 & ~n42941;
  assign n42949 = ~n40997 & ~n42948;
  assign n42950 = ~n42947 & n42949;
  assign n42951 = ~pi230 & ~n42950;
  assign n42952 = ~n42946 & n42951;
  assign n42953 = ~n38435 & n38440;
  assign n42954 = ~pi1156 & ~n42953;
  assign n42955 = n38617 & ~n38981;
  assign n42956 = ~n42954 & n42955;
  assign n42957 = ~n38386 & ~n42956;
  assign n42958 = pi211 & ~n42957;
  assign n42959 = n42899 & ~n42958;
  assign n42960 = pi1156 & n39762;
  assign n42961 = pi219 & ~n42960;
  assign n42962 = ~n42956 & n42961;
  assign n42963 = ~po1038 & ~n42962;
  assign n42964 = ~n42959 & n42963;
  assign n42965 = po1038 & n42938;
  assign n42966 = pi230 & ~n42965;
  assign n42967 = ~n42964 & n42966;
  assign po420 = ~n42952 & ~n42967;
  assign n42969 = ~pi796 & n40717;
  assign n42970 = pi264 & ~n40717;
  assign n42971 = ~pi1091 & ~n42969;
  assign n42972 = ~n42970 & n42971;
  assign n42973 = pi1091 & pi1141;
  assign n42974 = ~n42972 & ~n42973;
  assign n42975 = ~pi200 & ~n42974;
  assign n42976 = pi1091 & pi1142;
  assign n42977 = ~n42972 & ~n42976;
  assign n42978 = pi200 & ~n42977;
  assign n42979 = ~pi199 & ~n42975;
  assign n42980 = ~n42978 & n42979;
  assign n42981 = ~pi796 & n40706;
  assign n42982 = pi264 & ~n40706;
  assign n42983 = ~pi1091 & ~n42981;
  assign n42984 = ~n42982 & n42983;
  assign n42985 = pi1091 & pi1143;
  assign n42986 = ~pi200 & n42985;
  assign n42987 = pi199 & ~n42986;
  assign n42988 = ~n42984 & n42987;
  assign n42989 = n16429 & ~n42988;
  assign n42990 = ~n42980 & n42989;
  assign n42991 = ~pi211 & ~n42974;
  assign n42992 = pi211 & ~n42977;
  assign n42993 = ~pi219 & ~n42991;
  assign n42994 = ~n42992 & n42993;
  assign n42995 = pi219 & ~n42446;
  assign n42996 = ~n39284 & ~n42995;
  assign n42997 = ~n42984 & ~n42996;
  assign n42998 = ~n16429 & ~n42997;
  assign n42999 = ~n42994 & n42998;
  assign n43000 = ~n42990 & ~n42999;
  assign n43001 = ~pi230 & ~n43000;
  assign n43002 = ~pi211 & pi1141;
  assign n43003 = ~pi219 & ~n38332;
  assign n43004 = ~n43002 & n43003;
  assign n43005 = ~n39284 & ~n43004;
  assign n43006 = ~n16429 & ~n43005;
  assign n43007 = ~pi199 & pi1141;
  assign n43008 = n39254 & ~n43007;
  assign n43009 = ~n38321 & ~n43008;
  assign n43010 = n16429 & ~n43009;
  assign n43011 = pi230 & ~n43006;
  assign n43012 = ~n43010 & n43011;
  assign po421 = n43001 | n43012;
  assign n43014 = ~pi819 & n40717;
  assign n43015 = pi265 & ~n40717;
  assign n43016 = ~pi1091 & ~n43014;
  assign n43017 = ~n43015 & n43016;
  assign n43018 = ~n42976 & ~n43017;
  assign n43019 = ~pi200 & ~n43018;
  assign n43020 = ~n42985 & ~n43017;
  assign n43021 = pi200 & ~n43020;
  assign n43022 = ~pi199 & ~n43019;
  assign n43023 = ~n43021 & n43022;
  assign n43024 = ~pi819 & n40706;
  assign n43025 = pi265 & ~n40706;
  assign n43026 = ~pi1091 & ~n43024;
  assign n43027 = ~n43025 & n43026;
  assign n43028 = pi1091 & pi1144;
  assign n43029 = ~pi200 & n43028;
  assign n43030 = pi199 & ~n43029;
  assign n43031 = ~n43027 & n43030;
  assign n43032 = n16429 & ~n43031;
  assign n43033 = ~n43023 & n43032;
  assign n43034 = ~pi211 & ~n43018;
  assign n43035 = pi211 & ~n43020;
  assign n43036 = ~pi219 & ~n43034;
  assign n43037 = ~n43035 & n43036;
  assign n43038 = ~n40628 & ~n42995;
  assign n43039 = ~n43027 & ~n43038;
  assign n43040 = ~n16429 & ~n43039;
  assign n43041 = ~n43037 & n43040;
  assign n43042 = ~n43033 & ~n43041;
  assign n43043 = ~pi230 & ~n43042;
  assign n43044 = ~pi211 & pi1142;
  assign n43045 = ~pi219 & ~n38295;
  assign n43046 = ~n43044 & n43045;
  assign n43047 = ~n40628 & ~n43046;
  assign n43048 = ~n16429 & ~n43047;
  assign n43049 = ~n38320 & n40632;
  assign n43050 = ~n38314 & ~n43049;
  assign n43051 = n16429 & ~n43050;
  assign n43052 = pi230 & ~n43048;
  assign n43053 = ~n43051 & n43052;
  assign po422 = n43043 | n43053;
  assign n43055 = ~pi211 & pi1136;
  assign n43056 = pi219 & ~n43055;
  assign n43057 = pi211 & ~pi1135;
  assign n43058 = ~n43056 & ~n43057;
  assign n43059 = ~n10709 & n43058;
  assign n43060 = pi299 & n43059;
  assign n43061 = ~pi199 & pi1135;
  assign n43062 = pi200 & ~n43061;
  assign n43063 = pi199 & pi1136;
  assign n43064 = ~pi200 & ~n43063;
  assign n43065 = ~pi299 & ~n43062;
  assign n43066 = ~n43064 & n43065;
  assign n43067 = ~n43060 & ~n43066;
  assign n43068 = ~po1038 & ~n43067;
  assign n43069 = po1038 & n43059;
  assign n43070 = pi230 & ~n43069;
  assign n43071 = ~n43068 & n43070;
  assign n43072 = ~pi266 & ~n40717;
  assign n43073 = ~pi948 & n40717;
  assign n43074 = ~pi1091 & ~n43072;
  assign n43075 = ~n43073 & n43074;
  assign n43076 = ~pi199 & ~n43075;
  assign n43077 = pi1091 & pi1136;
  assign n43078 = ~pi266 & ~n40706;
  assign n43079 = ~pi948 & n40706;
  assign n43080 = ~pi1091 & ~n43078;
  assign n43081 = ~n43079 & n43080;
  assign n43082 = pi199 & ~n43081;
  assign n43083 = ~n43077 & n43082;
  assign n43084 = ~n43076 & ~n43083;
  assign n43085 = ~pi200 & n43084;
  assign n43086 = pi1091 & pi1135;
  assign n43087 = n43076 & ~n43086;
  assign n43088 = pi200 & ~n43082;
  assign n43089 = ~n43087 & n43088;
  assign n43090 = ~n43085 & ~n43089;
  assign n43091 = n16429 & ~n43090;
  assign n43092 = ~n42995 & ~n43056;
  assign n43093 = ~n43081 & ~n43092;
  assign n43094 = ~n16429 & ~n43093;
  assign n43095 = ~pi219 & ~n43075;
  assign n43096 = pi1135 & n42397;
  assign n43097 = n43095 & ~n43096;
  assign n43098 = n43094 & ~n43097;
  assign n43099 = ~pi230 & ~n43098;
  assign n43100 = ~n43091 & n43099;
  assign n43101 = ~n43071 & ~n43100;
  assign n43102 = ~pi1134 & ~n43101;
  assign n43103 = n38483 & ~n43063;
  assign n43104 = ~n43062 & ~n43103;
  assign n43105 = n16429 & n43104;
  assign n43106 = ~n16429 & n43058;
  assign n43107 = pi230 & ~n43105;
  assign n43108 = ~n43106 & n43107;
  assign n43109 = ~pi199 & pi1091;
  assign n43110 = ~n43084 & ~n43109;
  assign n43111 = ~pi200 & ~n43110;
  assign n43112 = ~n43089 & ~n43111;
  assign n43113 = n16429 & ~n43112;
  assign n43114 = pi1091 & ~n43057;
  assign n43115 = n43095 & ~n43114;
  assign n43116 = n43094 & ~n43115;
  assign n43117 = ~pi230 & ~n43116;
  assign n43118 = ~n43113 & n43117;
  assign n43119 = ~n43108 & ~n43118;
  assign n43120 = pi1134 & ~n43119;
  assign po423 = ~n43102 & ~n43120;
  assign n43122 = ~n42516 & n42519;
  assign n43123 = n42582 & ~n43122;
  assign n43124 = pi1154 & pi1155;
  assign n43125 = ~n40745 & n43124;
  assign n43126 = ~n42521 & n43125;
  assign n43127 = ~n43123 & ~n43126;
  assign n43128 = pi211 & ~n43127;
  assign n43129 = pi1153 & n40747;
  assign n43130 = n38359 & ~n42274;
  assign n43131 = ~n43129 & n43130;
  assign n43132 = ~n42498 & n43131;
  assign n43133 = n40877 & n42492;
  assign n43134 = ~pi1155 & ~n43133;
  assign n43135 = ~n43122 & n43134;
  assign n43136 = ~pi267 & ~n43135;
  assign n43137 = ~n43132 & n43136;
  assign n43138 = ~n43128 & n43137;
  assign n43139 = ~n42263 & ~n42281;
  assign n43140 = n40837 & ~n43139;
  assign n43141 = pi1154 & ~n43140;
  assign n43142 = ~pi1154 & ~n40888;
  assign n43143 = ~n42370 & n43142;
  assign n43144 = ~pi1155 & ~n43143;
  assign n43145 = ~n43141 & n43144;
  assign n43146 = pi1155 & ~n42348;
  assign n43147 = n40730 & ~n42843;
  assign n43148 = n43146 & ~n43147;
  assign n43149 = ~n42368 & n43148;
  assign n43150 = pi267 & ~n43149;
  assign n43151 = ~n43145 & n43150;
  assign n43152 = ~n43138 & ~n43151;
  assign n43153 = pi219 & ~n43152;
  assign n43154 = n40732 & ~n43140;
  assign n43155 = n42789 & ~n43154;
  assign n43156 = pi1154 & ~n43155;
  assign n43157 = ~pi1154 & ~n42260;
  assign n43158 = pi1155 & ~n43157;
  assign n43159 = n40777 & ~n43158;
  assign n43160 = ~n43156 & ~n43159;
  assign n43161 = ~pi1155 & ~n42601;
  assign n43162 = ~n43122 & n43161;
  assign n43163 = pi211 & ~n43162;
  assign n43164 = ~n43160 & n43163;
  assign n43165 = pi1153 & ~n40804;
  assign n43166 = ~pi1155 & ~n43165;
  assign n43167 = n42363 & n43166;
  assign n43168 = ~n42604 & ~n43129;
  assign n43169 = pi1155 & ~n43168;
  assign n43170 = ~pi1154 & ~n43167;
  assign n43171 = ~n43169 & n43170;
  assign n43172 = ~pi1153 & ~n42773;
  assign n43173 = n43166 & ~n43172;
  assign n43174 = pi1154 & ~n42774;
  assign n43175 = ~n43169 & n43174;
  assign n43176 = ~n43173 & n43175;
  assign n43177 = ~pi211 & ~n43171;
  assign n43178 = ~n43176 & n43177;
  assign n43179 = ~pi267 & ~n43178;
  assign n43180 = ~n43164 & n43179;
  assign n43181 = ~pi1153 & n40816;
  assign n43182 = ~n40806 & ~n43181;
  assign n43183 = ~pi1155 & n40732;
  assign n43184 = ~n43182 & n43183;
  assign n43185 = n42817 & n43146;
  assign n43186 = pi1154 & ~n43184;
  assign n43187 = ~n43185 & n43186;
  assign n43188 = ~pi1154 & ~n42281;
  assign n43189 = ~n40763 & n43188;
  assign n43190 = ~pi1155 & ~n43189;
  assign n43191 = ~n40782 & n43188;
  assign n43192 = ~n43190 & n43191;
  assign n43193 = ~n43187 & ~n43192;
  assign n43194 = pi211 & ~n43193;
  assign n43195 = pi1154 & n43182;
  assign n43196 = n43190 & ~n43195;
  assign n43197 = ~n40755 & ~n42584;
  assign n43198 = pi1154 & n40730;
  assign n43199 = pi1155 & ~n43198;
  assign n43200 = ~n43197 & n43199;
  assign n43201 = ~pi211 & ~n43200;
  assign n43202 = ~n43196 & n43201;
  assign n43203 = pi267 & ~n43202;
  assign n43204 = ~n43194 & n43203;
  assign n43205 = ~pi219 & ~n43204;
  assign n43206 = ~n43180 & n43205;
  assign n43207 = ~n43153 & ~n43206;
  assign n43208 = n40834 & ~n43207;
  assign n43209 = pi1155 & ~n42385;
  assign n43210 = ~n42641 & n43209;
  assign n43211 = ~pi1155 & ~n38929;
  assign n43212 = pi1091 & n43211;
  assign n43213 = ~n43210 & ~n43212;
  assign n43214 = ~pi1154 & ~n43213;
  assign n43215 = n42643 & n43209;
  assign n43216 = ~pi1155 & ~n42531;
  assign n43217 = ~n42414 & n43216;
  assign n43218 = ~n43215 & ~n43217;
  assign n43219 = pi1154 & ~n43218;
  assign n43220 = ~pi219 & ~n43214;
  assign n43221 = ~n43219 & n43220;
  assign n43222 = pi1091 & n42854;
  assign n43223 = ~n42384 & n43222;
  assign n43224 = pi1154 & ~n43223;
  assign n43225 = ~pi299 & n38816;
  assign n43226 = pi1091 & ~n43225;
  assign n43227 = n43224 & n43226;
  assign n43228 = pi1153 & n38824;
  assign n43229 = n42650 & ~n43228;
  assign n43230 = ~n39512 & n43229;
  assign n43231 = pi219 & ~n43230;
  assign n43232 = ~n43227 & n43231;
  assign n43233 = ~n43221 & ~n43232;
  assign n43234 = ~pi211 & ~n43233;
  assign n43235 = ~pi1155 & ~n38817;
  assign n43236 = ~n38504 & ~n43235;
  assign n43237 = ~n13026 & ~n43236;
  assign n43238 = pi1155 & n38832;
  assign n43239 = pi1154 & ~n43238;
  assign n43240 = pi1091 & n43239;
  assign n43241 = ~n43237 & n43240;
  assign n43242 = ~n38485 & ~n40911;
  assign n43243 = n43229 & ~n43242;
  assign n43244 = pi211 & ~n43243;
  assign n43245 = ~n43241 & n43244;
  assign n43246 = ~n43234 & ~n43245;
  assign n43247 = pi267 & ~n43246;
  assign n43248 = pi1091 & ~pi1155;
  assign n43249 = ~n38817 & n43248;
  assign n43250 = n38360 & ~n43249;
  assign n43251 = ~n43223 & n43250;
  assign n43252 = ~pi1154 & n38432;
  assign n43253 = ~n38517 & ~n43252;
  assign n43254 = ~n38465 & n43253;
  assign n43255 = pi1091 & n43254;
  assign n43256 = ~pi211 & ~n43255;
  assign n43257 = ~pi219 & ~n43251;
  assign n43258 = ~n43256 & n43257;
  assign n43259 = n43225 & n43248;
  assign n43260 = n43224 & ~n43259;
  assign n43261 = n42854 & n43239;
  assign n43262 = ~n43260 & ~n43261;
  assign n43263 = pi211 & ~n43262;
  assign n43264 = pi1154 & ~n43260;
  assign n43265 = ~n38485 & n42650;
  assign n43266 = ~n39511 & n43265;
  assign n43267 = ~pi211 & ~n43266;
  assign n43268 = ~n43264 & n43267;
  assign n43269 = pi219 & ~n43263;
  assign n43270 = ~n43268 & n43269;
  assign n43271 = ~n43258 & ~n43270;
  assign n43272 = n38424 & n42406;
  assign n43273 = ~n42617 & ~n43272;
  assign n43274 = ~n43211 & ~n43273;
  assign n43275 = pi211 & ~pi1154;
  assign n43276 = ~n43274 & n43275;
  assign n43277 = ~pi267 & ~n43276;
  assign n43278 = ~n43271 & n43277;
  assign n43279 = ~n43247 & ~n43278;
  assign n43280 = ~n40834 & ~n43279;
  assign n43281 = ~po1038 & ~n43280;
  assign n43282 = ~n43208 & n43281;
  assign n43283 = pi267 & n42560;
  assign n43284 = ~pi267 & ~n40724;
  assign n43285 = ~n42302 & n43284;
  assign n43286 = n40834 & ~n43285;
  assign n43287 = ~n43283 & n43286;
  assign n43288 = ~pi219 & ~n38360;
  assign n43289 = ~n38376 & n43288;
  assign n43290 = ~n39139 & ~n43289;
  assign n43291 = pi1091 & ~n43290;
  assign n43292 = ~pi267 & ~pi1091;
  assign n43293 = ~n40834 & n43292;
  assign n43294 = ~n43291 & ~n43293;
  assign n43295 = ~n43287 & n43294;
  assign n43296 = po1038 & ~n43295;
  assign n43297 = n40997 & ~n43296;
  assign n43298 = ~n43282 & n43297;
  assign n43299 = ~po1038 & n43279;
  assign n43300 = ~n43291 & ~n43292;
  assign n43301 = po1038 & ~n43300;
  assign n43302 = ~n40997 & ~n43301;
  assign n43303 = ~n43299 & n43302;
  assign n43304 = ~pi230 & ~n43303;
  assign n43305 = ~n43298 & n43304;
  assign n43306 = pi219 & ~n38832;
  assign n43307 = ~pi1155 & n43228;
  assign n43308 = ~pi1154 & ~n43307;
  assign n43309 = ~n38817 & ~n43308;
  assign n43310 = pi1155 & n39509;
  assign n43311 = ~n43309 & ~n43310;
  assign n43312 = ~n43306 & ~n43311;
  assign n43313 = pi211 & ~n43312;
  assign n43314 = ~pi199 & pi1154;
  assign n43315 = pi200 & ~n43314;
  assign n43316 = ~n38495 & ~n38831;
  assign n43317 = ~n43315 & n43316;
  assign n43318 = ~n38386 & ~n43317;
  assign n43319 = pi219 & ~n43318;
  assign n43320 = ~pi219 & n43254;
  assign n43321 = ~pi211 & ~n43320;
  assign n43322 = ~n43319 & n43321;
  assign n43323 = ~po1038 & ~n43322;
  assign n43324 = ~n43313 & n43323;
  assign n43325 = po1038 & n43290;
  assign n43326 = pi230 & ~n43325;
  assign n43327 = ~n43324 & n43326;
  assign po424 = ~n43305 & ~n43327;
  assign n43329 = ~n42290 & n42337;
  assign n43330 = ~n40743 & n42349;
  assign n43331 = pi219 & ~n42276;
  assign n43332 = ~n40737 & n43331;
  assign n43333 = ~n43330 & ~n43332;
  assign n43334 = ~po1038 & ~n42267;
  assign n43335 = n43333 & n43334;
  assign n43336 = ~n43329 & ~n43335;
  assign n43337 = ~pi1151 & ~n43336;
  assign n43338 = ~po1038 & ~n42364;
  assign n43339 = pi219 & n40882;
  assign n43340 = n43338 & ~n43339;
  assign n43341 = n42337 & ~n42559;
  assign n43342 = ~n43340 & ~n43341;
  assign n43343 = pi1151 & ~n43342;
  assign n43344 = ~n43337 & ~n43343;
  assign n43345 = pi268 & ~n43344;
  assign n43346 = po1038 & ~n42302;
  assign n43347 = ~n42334 & n43346;
  assign n43348 = po1038 & ~n42558;
  assign n43349 = ~n42288 & n43348;
  assign n43350 = n43347 & ~n43349;
  assign n43351 = pi219 & ~n40741;
  assign n43352 = ~n42322 & ~n43351;
  assign n43353 = ~n40742 & ~n43352;
  assign n43354 = ~po1038 & ~n40803;
  assign n43355 = n43353 & n43354;
  assign n43356 = ~n43350 & ~n43355;
  assign n43357 = ~pi1151 & n43356;
  assign n43358 = ~n40713 & ~n43342;
  assign n43359 = ~n40791 & n43338;
  assign n43360 = pi219 & po1038;
  assign n43361 = ~n40740 & n43360;
  assign n43362 = ~n42303 & ~n43361;
  assign n43363 = ~n43359 & n43362;
  assign n43364 = ~n43358 & ~n43363;
  assign n43365 = pi1151 & n43364;
  assign n43366 = ~pi268 & ~n43365;
  assign n43367 = ~n43357 & n43366;
  assign n43368 = ~n43345 & ~n43367;
  assign n43369 = ~pi1152 & ~n43368;
  assign n43370 = ~n42290 & n43348;
  assign n43371 = ~n40839 & ~n42371;
  assign n43372 = ~n43333 & ~n43371;
  assign n43373 = ~po1038 & ~n43372;
  assign n43374 = ~n40740 & ~n42351;
  assign n43375 = n43373 & ~n43374;
  assign n43376 = ~n43370 & ~n43375;
  assign n43377 = ~pi1151 & ~n43376;
  assign n43378 = ~n40709 & n43334;
  assign n43379 = ~n42559 & n43348;
  assign n43380 = ~n43340 & ~n43379;
  assign n43381 = ~n43378 & n43380;
  assign n43382 = pi1151 & ~n43381;
  assign n43383 = pi268 & ~n43382;
  assign n43384 = ~n43377 & n43383;
  assign n43385 = ~n42275 & ~n43353;
  assign n43386 = ~po1038 & ~n43385;
  assign n43387 = ~n43347 & ~n43386;
  assign n43388 = ~pi1151 & ~n43387;
  assign n43389 = ~pi219 & n40752;
  assign n43390 = ~n43331 & ~n43389;
  assign n43391 = ~po1038 & ~n43390;
  assign n43392 = ~n42291 & n43346;
  assign n43393 = ~n43350 & ~n43392;
  assign n43394 = ~n43391 & n43393;
  assign n43395 = pi1151 & ~n43394;
  assign n43396 = ~pi268 & ~n43395;
  assign n43397 = ~n43388 & n43396;
  assign n43398 = pi1152 & ~n43397;
  assign n43399 = ~n43384 & n43398;
  assign n43400 = ~n43369 & ~n43399;
  assign n43401 = pi1150 & ~n43400;
  assign n43402 = ~n42303 & n43346;
  assign n43403 = ~pi219 & ~n40777;
  assign n43404 = ~n40729 & ~n43403;
  assign n43405 = n43391 & n43404;
  assign n43406 = ~n43402 & ~n43405;
  assign n43407 = ~pi1151 & ~n43406;
  assign n43408 = ~po1038 & ~n43333;
  assign n43409 = ~n43392 & ~n43408;
  assign n43410 = pi1151 & ~n43409;
  assign n43411 = pi1152 & ~n43407;
  assign n43412 = ~n43410 & n43411;
  assign n43413 = ~n42292 & ~n43361;
  assign n43414 = ~n43373 & n43413;
  assign n43415 = pi1151 & n43414;
  assign n43416 = ~pi1151 & n43363;
  assign n43417 = ~pi1152 & ~n43416;
  assign n43418 = ~n43415 & n43417;
  assign n43419 = ~n43412 & ~n43418;
  assign n43420 = ~pi268 & ~n43419;
  assign n43421 = ~n42335 & n43348;
  assign n43422 = pi219 & ~n42368;
  assign n43423 = ~n42322 & ~n43422;
  assign n43424 = n40760 & ~n43423;
  assign n43425 = ~po1038 & ~n43424;
  assign n43426 = ~n43421 & ~n43425;
  assign n43427 = pi1151 & n43426;
  assign n43428 = ~po1038 & ~n42371;
  assign n43429 = ~n43422 & n43428;
  assign n43430 = ~n43349 & ~n43429;
  assign n43431 = ~pi1151 & n43430;
  assign n43432 = pi1152 & ~n43431;
  assign n43433 = ~n43427 & n43432;
  assign n43434 = ~po1038 & ~n42325;
  assign n43435 = ~n42322 & n43434;
  assign n43436 = ~n42338 & ~n43435;
  assign n43437 = pi1151 & n43436;
  assign n43438 = n40713 & ~n43342;
  assign n43439 = ~pi1151 & ~n43438;
  assign n43440 = ~pi1152 & ~n43439;
  assign n43441 = ~n43437 & n43440;
  assign n43442 = pi268 & ~n43441;
  assign n43443 = ~n43433 & n43442;
  assign n43444 = ~pi1150 & ~n43443;
  assign n43445 = ~n43420 & n43444;
  assign n43446 = ~n43401 & ~n43445;
  assign n43447 = n40996 & ~n43446;
  assign n43448 = pi268 & pi1152;
  assign n43449 = ~pi199 & n16429;
  assign n43450 = ~n40019 & ~n43449;
  assign n43451 = ~pi211 & ~n16429;
  assign n43452 = ~po1038 & n38424;
  assign n43453 = ~n43451 & ~n43452;
  assign n43454 = pi1152 & ~n43453;
  assign n43455 = n43450 & ~n43454;
  assign n43456 = ~pi1151 & n43453;
  assign n43457 = pi1150 & ~n43456;
  assign n43458 = ~n43455 & n43457;
  assign n43459 = ~n43448 & n43458;
  assign n43460 = ~n16429 & n42434;
  assign n43461 = ~po1038 & n38494;
  assign n43462 = ~n43460 & ~n43461;
  assign n43463 = pi1151 & ~n43462;
  assign n43464 = pi1152 & n43463;
  assign n43465 = ~pi1151 & n42226;
  assign n43466 = ~po1038 & ~n11423;
  assign n43467 = po1038 & n11421;
  assign n43468 = ~n43466 & ~n43467;
  assign n43469 = pi1151 & ~n43468;
  assign n43470 = ~pi1152 & ~n43469;
  assign n43471 = ~pi1150 & ~n43465;
  assign n43472 = ~n43470 & n43471;
  assign n43473 = ~n43464 & n43472;
  assign n43474 = ~n43459 & ~n43473;
  assign n43475 = pi1091 & ~n43474;
  assign n43476 = pi1152 & n43458;
  assign n43477 = pi1091 & ~n43476;
  assign n43478 = pi268 & ~n43477;
  assign n43479 = ~n43475 & ~n43478;
  assign n43480 = ~n40996 & ~n43479;
  assign n43481 = ~pi230 & ~n43480;
  assign n43482 = ~n43447 & n43481;
  assign n43483 = pi230 & ~n43458;
  assign n43484 = ~n43473 & n43483;
  assign po425 = ~n43482 & ~n43484;
  assign n43486 = ~pi199 & pi1137;
  assign n43487 = pi200 & ~n43486;
  assign n43488 = pi199 & pi1138;
  assign n43489 = ~pi199 & pi1136;
  assign n43490 = ~pi200 & ~n43488;
  assign n43491 = ~n43489 & n43490;
  assign n43492 = ~n43487 & ~n43491;
  assign n43493 = n16429 & ~n43492;
  assign n43494 = ~pi211 & pi1138;
  assign n43495 = pi219 & n43494;
  assign n43496 = pi211 & pi1137;
  assign n43497 = ~n43055 & ~n43496;
  assign n43498 = ~pi219 & ~n43497;
  assign n43499 = ~n43495 & ~n43498;
  assign n43500 = ~n16429 & n43499;
  assign n43501 = ~n43493 & ~n43500;
  assign n43502 = pi230 & ~n43501;
  assign n43503 = ~pi200 & n43077;
  assign n43504 = pi1137 & n40935;
  assign n43505 = ~n43503 & ~n43504;
  assign n43506 = n43449 & n43505;
  assign n43507 = pi1091 & ~n43497;
  assign n43508 = n40019 & ~n43507;
  assign n43509 = ~n43506 & ~n43508;
  assign n43510 = ~pi817 & n40717;
  assign n43511 = pi269 & ~n40717;
  assign n43512 = ~pi1091 & ~n43510;
  assign n43513 = ~n43511 & n43512;
  assign n43514 = ~n43509 & ~n43513;
  assign n43515 = ~pi817 & n40706;
  assign n43516 = pi269 & ~n40706;
  assign n43517 = ~pi1091 & ~n43515;
  assign n43518 = ~n43516 & n43517;
  assign n43519 = pi1138 & n42446;
  assign n43520 = pi219 & ~n16429;
  assign n43521 = ~n43519 & n43520;
  assign n43522 = ~pi200 & pi1091;
  assign n43523 = pi1138 & n43522;
  assign n43524 = pi199 & ~n43523;
  assign n43525 = n16429 & n43524;
  assign n43526 = ~n43521 & ~n43525;
  assign n43527 = ~n43518 & ~n43526;
  assign n43528 = ~n43514 & ~n43527;
  assign n43529 = ~pi230 & ~n43528;
  assign po426 = ~n43502 & ~n43529;
  assign n43531 = ~pi805 & n40706;
  assign n43532 = pi270 & ~n40706;
  assign n43533 = ~pi1091 & ~n43531;
  assign n43534 = ~n43532 & n43533;
  assign n43535 = n42446 & n43002;
  assign n43536 = n43520 & ~n43535;
  assign n43537 = ~pi200 & n42973;
  assign n43538 = pi199 & ~n43537;
  assign n43539 = n16429 & n43538;
  assign n43540 = ~n43536 & ~n43539;
  assign n43541 = ~n43534 & ~n43540;
  assign n43542 = ~pi805 & n40717;
  assign n43543 = pi270 & ~n40717;
  assign n43544 = ~pi1091 & ~n43542;
  assign n43545 = ~n43543 & n43544;
  assign n43546 = ~pi211 & pi1139;
  assign n43547 = pi211 & pi1140;
  assign n43548 = ~n43546 & ~n43547;
  assign n43549 = pi1091 & ~n43548;
  assign n43550 = n40019 & ~n43549;
  assign n43551 = pi1091 & pi1140;
  assign n43552 = pi200 & n43551;
  assign n43553 = pi1139 & n43522;
  assign n43554 = ~n43552 & ~n43553;
  assign n43555 = n43449 & n43554;
  assign n43556 = ~n43550 & ~n43555;
  assign n43557 = ~n43545 & ~n43556;
  assign n43558 = ~pi230 & ~n43541;
  assign n43559 = ~n43557 & n43558;
  assign n43560 = pi219 & ~n43002;
  assign n43561 = ~pi219 & n43548;
  assign n43562 = ~n43560 & ~n43561;
  assign n43563 = ~n16429 & ~n43562;
  assign n43564 = ~pi199 & pi1140;
  assign n43565 = pi200 & ~n43564;
  assign n43566 = pi199 & pi1141;
  assign n43567 = ~pi199 & pi1139;
  assign n43568 = ~pi200 & ~n43566;
  assign n43569 = ~n43567 & n43568;
  assign n43570 = ~n43565 & ~n43569;
  assign n43571 = n16429 & ~n43570;
  assign n43572 = pi230 & ~n43563;
  assign n43573 = ~n43571 & n43572;
  assign po427 = n43559 | n43573;
  assign n43575 = ~pi271 & ~n40738;
  assign n43576 = ~n40710 & ~n43575;
  assign n43577 = pi219 & ~n43576;
  assign n43578 = ~pi1091 & ~n40719;
  assign n43579 = pi271 & ~n43578;
  assign n43580 = ~pi271 & ~n40720;
  assign n43581 = ~n43579 & ~n43580;
  assign n43582 = pi1091 & pi1146;
  assign n43583 = ~n43581 & ~n43582;
  assign n43584 = ~pi211 & n43582;
  assign n43585 = ~n43583 & ~n43584;
  assign n43586 = pi1091 & n39277;
  assign n43587 = ~pi219 & ~n43586;
  assign n43588 = ~n43585 & n43587;
  assign n43589 = ~n43577 & ~n43588;
  assign n43590 = ~pi211 & pi1147;
  assign n43591 = n42294 & n43590;
  assign n43592 = ~n16429 & ~n43591;
  assign n43593 = ~n43589 & n43592;
  assign n43594 = pi199 & ~n43576;
  assign n43595 = ~pi199 & n43583;
  assign n43596 = ~n43594 & ~n43595;
  assign n43597 = pi200 & ~n43596;
  assign n43598 = pi1091 & pi1145;
  assign n43599 = ~pi199 & ~n43598;
  assign n43600 = ~n43581 & n43599;
  assign n43601 = ~n43594 & ~n43600;
  assign n43602 = pi1147 & n40921;
  assign n43603 = ~pi200 & ~n43602;
  assign n43604 = ~n43601 & n43603;
  assign n43605 = ~n43597 & ~n43604;
  assign n43606 = n16429 & ~n43605;
  assign n43607 = ~n43593 & ~n43606;
  assign n43608 = ~pi230 & ~n43607;
  assign n43609 = ~pi200 & ~n39258;
  assign n43610 = n40182 & ~n43609;
  assign n43611 = pi1147 & n42222;
  assign n43612 = ~n40076 & ~n40091;
  assign n43613 = ~pi219 & ~n43612;
  assign n43614 = ~n43610 & ~n43611;
  assign n43615 = ~n43613 & n43614;
  assign n43616 = ~po1038 & ~n43615;
  assign n43617 = pi219 & ~n43590;
  assign n43618 = ~n39277 & n41362;
  assign n43619 = ~n43617 & ~n43618;
  assign n43620 = po1038 & n43619;
  assign n43621 = pi230 & ~n43620;
  assign n43622 = ~n43616 & n43621;
  assign po428 = ~n43608 & ~n43622;
  assign n43624 = pi1150 & n43381;
  assign n43625 = ~pi1150 & n43342;
  assign n43626 = pi1149 & ~n43625;
  assign n43627 = ~n43624 & n43626;
  assign n43628 = pi1150 & n43376;
  assign n43629 = ~pi1150 & n43336;
  assign n43630 = ~pi1149 & ~n43629;
  assign n43631 = ~n43628 & n43630;
  assign n43632 = ~n43627 & ~n43631;
  assign n43633 = pi1148 & ~n43632;
  assign n43634 = pi1150 & n43430;
  assign n43635 = ~pi1150 & ~n43438;
  assign n43636 = ~pi1149 & ~n43635;
  assign n43637 = ~n43634 & n43636;
  assign n43638 = pi1150 & n43426;
  assign n43639 = ~pi1150 & n43436;
  assign n43640 = pi1149 & ~n43639;
  assign n43641 = ~n43638 & n43640;
  assign n43642 = ~n43637 & ~n43641;
  assign n43643 = ~pi1148 & ~n43642;
  assign n43644 = pi283 & ~n43643;
  assign n43645 = ~n43633 & n43644;
  assign n43646 = po1038 & n10709;
  assign n43647 = ~n13029 & ~n43646;
  assign n43648 = ~pi1150 & n43647;
  assign n43649 = ~n43453 & ~n43648;
  assign n43650 = ~pi1149 & ~n43649;
  assign n43651 = pi1149 & ~pi1150;
  assign n43652 = ~n43453 & ~n43651;
  assign n43653 = n43450 & ~n43652;
  assign n43654 = ~n43650 & ~n43653;
  assign n43655 = pi1091 & ~n43654;
  assign n43656 = pi1148 & ~n43655;
  assign n43657 = pi1150 & ~n42226;
  assign n43658 = ~pi1149 & ~n43657;
  assign n43659 = pi1091 & n43658;
  assign n43660 = pi1150 & n43462;
  assign n43661 = ~pi1150 & ~n43468;
  assign n43662 = pi1091 & pi1149;
  assign n43663 = ~n43661 & n43662;
  assign n43664 = ~n43660 & n43663;
  assign n43665 = ~pi1148 & ~n43664;
  assign n43666 = ~n43659 & n43665;
  assign n43667 = ~pi283 & ~n43666;
  assign n43668 = ~n43656 & n43667;
  assign n43669 = pi272 & ~n43668;
  assign n43670 = ~n43645 & n43669;
  assign n43671 = pi1150 & ~n43394;
  assign n43672 = ~pi1150 & ~n43364;
  assign n43673 = pi1149 & ~n43672;
  assign n43674 = ~n43671 & n43673;
  assign n43675 = pi1150 & ~n43387;
  assign n43676 = ~pi1150 & ~n43356;
  assign n43677 = ~pi1149 & ~n43676;
  assign n43678 = ~n43675 & n43677;
  assign n43679 = ~n43674 & ~n43678;
  assign n43680 = pi1148 & ~n43679;
  assign n43681 = ~pi1150 & ~n43414;
  assign n43682 = pi1150 & n43409;
  assign n43683 = pi1149 & ~n43682;
  assign n43684 = ~n43681 & n43683;
  assign n43685 = pi1150 & n43406;
  assign n43686 = ~pi1150 & ~n43363;
  assign n43687 = ~pi1149 & ~n43686;
  assign n43688 = ~n43685 & n43687;
  assign n43689 = ~pi1148 & ~n43688;
  assign n43690 = ~n43684 & n43689;
  assign n43691 = ~n43680 & ~n43690;
  assign n43692 = pi283 & ~n43691;
  assign n43693 = ~po1038 & n38415;
  assign n43694 = ~n40019 & ~n43693;
  assign n43695 = ~n43451 & n43694;
  assign n43696 = pi1150 & ~n43695;
  assign n43697 = pi1149 & ~n43696;
  assign n43698 = n43450 & n43697;
  assign n43699 = pi1148 & ~n43650;
  assign n43700 = ~n43698 & n43699;
  assign n43701 = pi1091 & n43700;
  assign n43702 = pi1091 & n43666;
  assign n43703 = ~pi283 & ~n43702;
  assign n43704 = ~n43701 & n43703;
  assign n43705 = ~pi272 & ~n43704;
  assign n43706 = ~n43692 & n43705;
  assign n43707 = ~pi230 & ~n43670;
  assign n43708 = ~n43706 & n43707;
  assign n43709 = pi1149 & ~n43462;
  assign n43710 = ~n43697 & ~n43709;
  assign n43711 = ~n43661 & ~n43710;
  assign n43712 = ~pi1148 & ~n43658;
  assign n43713 = ~n43711 & n43712;
  assign n43714 = pi230 & ~n43700;
  assign n43715 = ~n43713 & n43714;
  assign po429 = ~n43708 & ~n43715;
  assign n43717 = ~pi273 & ~n40739;
  assign n43718 = ~n40712 & ~n43717;
  assign n43719 = pi219 & ~n43718;
  assign n43720 = ~pi273 & ~n40721;
  assign n43721 = n40723 & ~n43720;
  assign n43722 = ~pi219 & ~n43584;
  assign n43723 = ~n43721 & n43722;
  assign n43724 = ~n43719 & ~n43723;
  assign n43725 = pi299 & n43724;
  assign n43726 = ~pi200 & n43582;
  assign n43727 = ~pi199 & ~n43726;
  assign n43728 = ~n43721 & n43727;
  assign n43729 = pi199 & ~n43718;
  assign n43730 = ~pi299 & ~n43729;
  assign n43731 = ~n43728 & n43730;
  assign n43732 = ~n43725 & ~n43731;
  assign n43733 = ~n11422 & ~n40879;
  assign n43734 = pi1091 & ~n43733;
  assign n43735 = n43732 & ~n43734;
  assign n43736 = ~po1038 & ~n43735;
  assign n43737 = pi1091 & n42338;
  assign n43738 = ~n43736 & ~n43737;
  assign n43739 = pi1147 & ~n43738;
  assign n43740 = po1038 & n43724;
  assign n43741 = n40255 & ~n43732;
  assign n43742 = ~pi1148 & ~n43741;
  assign n43743 = pi1091 & n38395;
  assign n43744 = ~n43724 & ~n43743;
  assign n43745 = pi299 & ~n43744;
  assign n43746 = n40922 & ~n43597;
  assign n43747 = ~n43731 & ~n43746;
  assign n43748 = ~n43745 & n43747;
  assign n43749 = ~po1038 & ~n43748;
  assign n43750 = n42224 & n42294;
  assign n43751 = pi1148 & ~n43750;
  assign n43752 = ~n43749 & n43751;
  assign n43753 = ~n43742 & ~n43752;
  assign n43754 = ~n43740 & ~n43753;
  assign n43755 = ~n43739 & n43754;
  assign n43756 = ~pi230 & ~n43755;
  assign n43757 = ~pi211 & ~n40090;
  assign n43758 = n40019 & ~n43757;
  assign n43759 = ~pi1146 & n10793;
  assign n43760 = n43449 & ~n43759;
  assign n43761 = ~n43758 & ~n43760;
  assign n43762 = pi1147 & ~n43761;
  assign n43763 = pi1146 & ~n41274;
  assign n43764 = ~n43647 & n43763;
  assign n43765 = ~pi1148 & ~n43764;
  assign n43766 = ~n43762 & n43765;
  assign n43767 = ~pi1146 & n10709;
  assign n43768 = pi1147 & n40019;
  assign n43769 = ~n43451 & ~n43768;
  assign n43770 = ~n43767 & ~n43769;
  assign n43771 = ~pi199 & pi1147;
  assign n43772 = pi200 & ~n43771;
  assign n43773 = ~n43759 & ~n43772;
  assign n43774 = n16429 & n43773;
  assign n43775 = pi1148 & ~n43774;
  assign n43776 = ~n43770 & n43775;
  assign n43777 = pi230 & ~n43766;
  assign n43778 = ~n43776 & n43777;
  assign po430 = n43756 | n43778;
  assign n43780 = ~pi659 & n40717;
  assign n43781 = pi274 & ~n40717;
  assign n43782 = ~pi1091 & ~n43780;
  assign n43783 = ~n43781 & n43782;
  assign n43784 = ~n43028 & ~n43783;
  assign n43785 = pi200 & ~n43784;
  assign n43786 = ~n42985 & ~n43783;
  assign n43787 = ~pi200 & ~n43786;
  assign n43788 = ~pi199 & ~n43785;
  assign n43789 = ~n43787 & n43788;
  assign n43790 = ~pi659 & n40706;
  assign n43791 = pi274 & ~n40706;
  assign n43792 = ~pi1091 & ~n43790;
  assign n43793 = ~n43791 & n43792;
  assign n43794 = ~pi200 & n43598;
  assign n43795 = pi199 & ~n43794;
  assign n43796 = ~n43793 & n43795;
  assign n43797 = n16429 & ~n43796;
  assign n43798 = ~n43789 & n43797;
  assign n43799 = pi211 & ~n43784;
  assign n43800 = ~pi211 & ~n43786;
  assign n43801 = ~pi219 & ~n43799;
  assign n43802 = ~n43800 & n43801;
  assign n43803 = pi219 & ~n43586;
  assign n43804 = ~n43793 & n43803;
  assign n43805 = ~n16429 & ~n43804;
  assign n43806 = ~n43802 & n43805;
  assign n43807 = ~pi230 & ~n43798;
  assign n43808 = ~n43806 & n43807;
  assign n43809 = ~pi219 & ~n38302;
  assign n43810 = ~n39278 & n43809;
  assign n43811 = ~n40073 & ~n43810;
  assign n43812 = ~n38384 & ~n40076;
  assign n43813 = ~n43810 & ~n43812;
  assign n43814 = ~n38313 & n40187;
  assign n43815 = n40637 & ~n43814;
  assign n43816 = ~n43813 & ~n43815;
  assign n43817 = ~po1038 & ~n43816;
  assign n43818 = pi230 & ~n43817;
  assign n43819 = ~n43811 & n43818;
  assign po431 = ~n43808 & ~n43819;
  assign n43821 = pi1151 & ~n43453;
  assign n43822 = pi1149 & n43450;
  assign n43823 = ~n43821 & n43822;
  assign n43824 = ~pi1149 & n43463;
  assign n43825 = ~n43823 & ~n43824;
  assign n43826 = pi1150 & ~n43825;
  assign n43827 = ~pi1151 & n43647;
  assign n43828 = pi1149 & ~n43453;
  assign n43829 = ~n43827 & n43828;
  assign n43830 = ~pi1149 & pi1151;
  assign n43831 = ~n42226 & n43830;
  assign n43832 = ~pi1150 & ~n43831;
  assign n43833 = ~n43829 & n43832;
  assign n43834 = ~n43826 & ~n43833;
  assign n43835 = pi1091 & ~n43834;
  assign n43836 = pi1091 & ~pi1151;
  assign n43837 = n41321 & n43836;
  assign n43838 = n43468 & n43837;
  assign n43839 = ~n43835 & ~n43838;
  assign n43840 = pi275 & ~n43839;
  assign n43841 = ~pi1151 & n43468;
  assign n43842 = pi1150 & ~n43841;
  assign n43843 = ~n43463 & n43842;
  assign n43844 = n40461 & ~n42226;
  assign n43845 = ~pi1149 & ~n43844;
  assign n43846 = ~n43843 & n43845;
  assign n43847 = n43453 & n43651;
  assign n43848 = ~n43823 & ~n43847;
  assign n43849 = ~n43846 & n43848;
  assign n43850 = pi1091 & n43849;
  assign n43851 = ~pi275 & ~n43850;
  assign n43852 = ~n40995 & ~n43851;
  assign n43853 = ~n43840 & n43852;
  assign n43854 = ~pi1150 & n43406;
  assign n43855 = pi1151 & ~n43682;
  assign n43856 = ~n43854 & n43855;
  assign n43857 = pi1150 & ~n43414;
  assign n43858 = ~pi1151 & ~n43686;
  assign n43859 = ~n43857 & n43858;
  assign n43860 = ~n43856 & ~n43859;
  assign n43861 = ~pi275 & ~n43860;
  assign n43862 = ~pi1150 & n43430;
  assign n43863 = ~n43638 & ~n43862;
  assign n43864 = pi1151 & ~n43863;
  assign n43865 = pi1150 & n43436;
  assign n43866 = ~n43635 & ~n43865;
  assign n43867 = ~pi1151 & ~n43866;
  assign n43868 = pi275 & ~n43867;
  assign n43869 = ~n43864 & n43868;
  assign n43870 = ~pi1149 & ~n43869;
  assign n43871 = ~n43861 & n43870;
  assign n43872 = pi1151 & ~n43376;
  assign n43873 = ~pi1150 & ~n43337;
  assign n43874 = ~n43872 & n43873;
  assign n43875 = ~pi1151 & ~n43342;
  assign n43876 = pi1150 & ~n43875;
  assign n43877 = ~n43382 & n43876;
  assign n43878 = pi275 & ~n43877;
  assign n43879 = ~n43874 & n43878;
  assign n43880 = ~pi1150 & ~n43387;
  assign n43881 = pi1151 & ~n43671;
  assign n43882 = ~n43880 & n43881;
  assign n43883 = pi1150 & ~n43364;
  assign n43884 = ~pi1151 & ~n43883;
  assign n43885 = ~n43676 & n43884;
  assign n43886 = ~pi275 & ~n43885;
  assign n43887 = ~n43882 & n43886;
  assign n43888 = pi1149 & ~n43887;
  assign n43889 = ~n43879 & n43888;
  assign n43890 = n40995 & ~n43871;
  assign n43891 = ~n43889 & n43890;
  assign n43892 = ~n43853 & ~n43891;
  assign n43893 = ~pi230 & ~n43892;
  assign n43894 = pi230 & n43849;
  assign po432 = n43893 | n43894;
  assign n43896 = ~pi276 & ~n40718;
  assign n43897 = n43578 & ~n43896;
  assign n43898 = ~n38296 & ~n40062;
  assign n43899 = pi1091 & ~n43898;
  assign n43900 = n40019 & ~n43899;
  assign n43901 = pi1145 & n40935;
  assign n43902 = ~n43029 & ~n43901;
  assign n43903 = n43449 & n43902;
  assign n43904 = ~n43900 & ~n43903;
  assign n43905 = ~n43897 & ~n43904;
  assign n43906 = ~pi276 & ~n40707;
  assign n43907 = n40709 & ~n43906;
  assign n43908 = n43520 & ~n43584;
  assign n43909 = pi199 & ~n43726;
  assign n43910 = n16429 & n43909;
  assign n43911 = ~n43908 & ~n43910;
  assign n43912 = ~n43907 & ~n43911;
  assign n43913 = ~pi230 & ~n43905;
  assign n43914 = ~n43912 & n43913;
  assign n43915 = ~n38311 & n41126;
  assign n43916 = ~n40189 & ~n43915;
  assign n43917 = n16429 & ~n43916;
  assign n43918 = ~pi219 & ~n43898;
  assign n43919 = pi1146 & n38395;
  assign n43920 = ~n43918 & ~n43919;
  assign n43921 = ~n16429 & n43920;
  assign n43922 = pi230 & ~n43917;
  assign n43923 = ~n43921 & n43922;
  assign po433 = n43914 | n43923;
  assign n43925 = ~pi820 & n40717;
  assign n43926 = pi277 & ~n40717;
  assign n43927 = ~pi1091 & ~n43925;
  assign n43928 = ~n43926 & n43927;
  assign n43929 = ~n43551 & ~n43928;
  assign n43930 = ~pi200 & ~n43929;
  assign n43931 = ~n42973 & ~n43928;
  assign n43932 = pi200 & ~n43931;
  assign n43933 = ~pi199 & ~n43930;
  assign n43934 = ~n43932 & n43933;
  assign n43935 = ~pi820 & n40706;
  assign n43936 = pi277 & ~n40706;
  assign n43937 = ~pi1091 & ~n43935;
  assign n43938 = ~n43936 & n43937;
  assign n43939 = ~pi200 & n42976;
  assign n43940 = pi199 & ~n43939;
  assign n43941 = ~n43938 & n43940;
  assign n43942 = n16429 & ~n43941;
  assign n43943 = ~n43934 & n43942;
  assign n43944 = ~pi211 & ~n43929;
  assign n43945 = pi211 & ~n43931;
  assign n43946 = ~pi219 & ~n43944;
  assign n43947 = ~n43945 & n43946;
  assign n43948 = pi219 & ~n43044;
  assign n43949 = ~n42995 & ~n43948;
  assign n43950 = ~n43938 & ~n43949;
  assign n43951 = ~n16429 & ~n43950;
  assign n43952 = ~n43947 & n43951;
  assign n43953 = ~n43943 & ~n43952;
  assign n43954 = ~pi230 & ~n43953;
  assign n43955 = pi211 & pi1141;
  assign n43956 = ~pi211 & pi1140;
  assign n43957 = ~pi219 & ~n43955;
  assign n43958 = ~n43956 & n43957;
  assign n43959 = ~n43948 & ~n43958;
  assign n43960 = ~n16429 & ~n43959;
  assign n43961 = n38310 & ~n43564;
  assign n43962 = pi200 & ~n43007;
  assign n43963 = ~n43961 & ~n43962;
  assign n43964 = n16429 & ~n43963;
  assign n43965 = pi230 & ~n43960;
  assign n43966 = ~n43964 & n43965;
  assign po434 = n43954 | n43966;
  assign n43968 = ~pi278 & ~n40706;
  assign n43969 = ~pi976 & n40706;
  assign n43970 = ~pi1091 & ~n43968;
  assign n43971 = ~n43969 & n43970;
  assign n43972 = pi199 & ~n43971;
  assign n43973 = pi1091 & ~pi1132;
  assign n43974 = pi976 & n40717;
  assign n43975 = pi278 & ~n40717;
  assign n43976 = ~pi1091 & ~n43974;
  assign n43977 = ~n43975 & n43976;
  assign n43978 = ~n43973 & ~n43977;
  assign n43979 = ~pi199 & ~n43978;
  assign n43980 = ~n43972 & ~n43979;
  assign n43981 = ~pi200 & ~n43980;
  assign n43982 = pi1091 & ~pi1133;
  assign n43983 = ~n43977 & ~n43982;
  assign n43984 = ~pi199 & ~n43983;
  assign n43985 = ~n43972 & ~n43984;
  assign n43986 = pi200 & ~n43985;
  assign n43987 = ~pi299 & ~n43986;
  assign n43988 = ~n43981 & n43987;
  assign n43989 = pi219 & ~n43971;
  assign n43990 = pi211 & ~pi1133;
  assign n43991 = ~pi211 & ~pi1132;
  assign n43992 = ~n43990 & ~n43991;
  assign n43993 = pi1091 & ~n43992;
  assign n43994 = ~n43977 & ~n43993;
  assign n43995 = ~pi219 & ~n43994;
  assign n43996 = ~n43989 & ~n43995;
  assign n43997 = pi299 & n43996;
  assign n43998 = ~n43988 & ~n43997;
  assign n43999 = ~po1038 & ~n43998;
  assign n44000 = po1038 & n43996;
  assign n44001 = ~pi230 & ~n44000;
  assign n44002 = ~n43999 & n44001;
  assign n44003 = ~pi199 & pi1132;
  assign n44004 = ~pi200 & ~n44003;
  assign n44005 = ~pi199 & pi1133;
  assign n44006 = pi200 & ~n44005;
  assign n44007 = ~pi299 & ~n44006;
  assign n44008 = ~n44004 & n44007;
  assign n44009 = n38384 & n43992;
  assign n44010 = ~n44008 & ~n44009;
  assign n44011 = ~po1038 & ~n44010;
  assign n44012 = n39240 & n43992;
  assign n44013 = pi230 & ~n44012;
  assign n44014 = ~n44011 & n44013;
  assign n44015 = ~n44002 & ~n44014;
  assign n44016 = ~pi1134 & ~n44015;
  assign n44017 = n10793 & ~n44003;
  assign n44018 = n44007 & ~n44017;
  assign n44019 = ~n42460 & ~n44009;
  assign n44020 = ~n44018 & n44019;
  assign n44021 = ~po1038 & ~n44020;
  assign n44022 = ~n42225 & ~n44021;
  assign n44023 = n44013 & n44022;
  assign n44024 = ~n40921 & n43981;
  assign n44025 = n43987 & ~n44024;
  assign n44026 = n13026 & n42446;
  assign n44027 = ~n43997 & ~n44026;
  assign n44028 = ~n44025 & n44027;
  assign n44029 = ~po1038 & ~n44028;
  assign n44030 = ~n43750 & n44001;
  assign n44031 = ~n44029 & n44030;
  assign n44032 = ~n44023 & ~n44031;
  assign n44033 = pi1134 & ~n44032;
  assign po435 = ~n44016 & ~n44033;
  assign n44035 = ~pi279 & ~n40706;
  assign n44036 = ~pi958 & n40706;
  assign n44037 = ~pi1091 & ~n44035;
  assign n44038 = ~n44036 & n44037;
  assign n44039 = pi1135 & n43522;
  assign n44040 = ~n44038 & ~n44039;
  assign n44041 = pi199 & ~n44040;
  assign n44042 = pi958 & n40717;
  assign n44043 = pi279 & ~n40717;
  assign n44044 = ~pi1091 & ~n44042;
  assign n44045 = ~n44043 & n44044;
  assign n44046 = ~pi1133 & n43522;
  assign n44047 = ~pi199 & ~n44046;
  assign n44048 = ~n44045 & n44047;
  assign n44049 = ~n44041 & ~n44048;
  assign n44050 = n16429 & ~n44049;
  assign n44051 = ~n40935 & n44050;
  assign n44052 = ~n42397 & ~n43982;
  assign n44053 = ~n44045 & n44052;
  assign n44054 = ~pi219 & ~n44053;
  assign n44055 = pi1135 & n42446;
  assign n44056 = pi219 & ~n44055;
  assign n44057 = ~n44038 & n44056;
  assign n44058 = ~n16429 & ~n44057;
  assign n44059 = ~n44054 & n44058;
  assign n44060 = ~pi230 & ~n44059;
  assign n44061 = ~n44051 & n44060;
  assign n44062 = pi199 & pi1135;
  assign n44063 = ~n44005 & ~n44062;
  assign n44064 = n38424 & ~n44063;
  assign n44065 = pi1135 & n38395;
  assign n44066 = ~pi211 & ~pi1133;
  assign n44067 = ~pi219 & ~n44066;
  assign n44068 = ~pi211 & n44067;
  assign n44069 = ~n44065 & ~n44068;
  assign n44070 = pi299 & ~n44069;
  assign n44071 = ~n44064 & ~n44070;
  assign n44072 = ~po1038 & ~n44071;
  assign n44073 = po1038 & ~n44069;
  assign n44074 = pi230 & ~n44073;
  assign n44075 = ~n44072 & n44074;
  assign n44076 = ~n44061 & ~n44075;
  assign n44077 = ~pi1134 & ~n44076;
  assign n44078 = ~pi1133 & n10793;
  assign n44079 = ~pi200 & pi1135;
  assign n44080 = pi199 & ~n44079;
  assign n44081 = ~n44078 & ~n44080;
  assign n44082 = n16429 & ~n44081;
  assign n44083 = ~n44065 & ~n44067;
  assign n44084 = ~n16429 & n44083;
  assign n44085 = ~n44082 & ~n44084;
  assign n44086 = pi230 & ~n44085;
  assign n44087 = pi1091 & ~n44066;
  assign n44088 = n40019 & n44087;
  assign n44089 = ~n44050 & ~n44088;
  assign n44090 = n44060 & n44089;
  assign n44091 = ~n44086 & ~n44090;
  assign n44092 = pi1134 & ~n44091;
  assign po436 = ~n44077 & ~n44092;
  assign n44094 = ~pi211 & pi1135;
  assign n44095 = pi211 & pi1136;
  assign n44096 = ~n44094 & ~n44095;
  assign n44097 = pi1091 & n44096;
  assign n44098 = ~pi280 & ~n40717;
  assign n44099 = pi914 & n40717;
  assign n44100 = ~pi1091 & ~n44098;
  assign n44101 = ~n44099 & n44100;
  assign n44102 = ~n44097 & ~n44101;
  assign n44103 = ~pi219 & ~n44102;
  assign n44104 = ~pi211 & pi1137;
  assign n44105 = pi219 & ~n44104;
  assign n44106 = ~n42995 & ~n44105;
  assign n44107 = ~pi914 & n40706;
  assign n44108 = pi280 & ~n40706;
  assign n44109 = ~pi1091 & ~n44107;
  assign n44110 = ~n44108 & n44109;
  assign n44111 = ~n44106 & ~n44110;
  assign n44112 = ~n44103 & ~n44111;
  assign n44113 = ~n16429 & ~n44112;
  assign n44114 = pi1137 & n43522;
  assign n44115 = ~n44110 & ~n44114;
  assign n44116 = pi199 & ~n44115;
  assign n44117 = pi200 & pi1136;
  assign n44118 = pi1091 & ~n44079;
  assign n44119 = ~n44117 & n44118;
  assign n44120 = ~pi199 & ~n44119;
  assign n44121 = ~n44101 & n44120;
  assign n44122 = n16429 & ~n44116;
  assign n44123 = ~n44121 & n44122;
  assign n44124 = ~n44113 & ~n44123;
  assign n44125 = ~pi230 & ~n44124;
  assign n44126 = pi200 & ~n43489;
  assign n44127 = pi199 & pi1137;
  assign n44128 = ~pi200 & ~n43061;
  assign n44129 = ~n44127 & n44128;
  assign n44130 = ~n44126 & ~n44129;
  assign n44131 = n16429 & n44130;
  assign n44132 = ~pi219 & n44096;
  assign n44133 = ~n44105 & ~n44132;
  assign n44134 = ~n16429 & n44133;
  assign n44135 = pi230 & ~n44131;
  assign n44136 = ~n44134 & n44135;
  assign po437 = ~n44125 & ~n44136;
  assign n44138 = ~pi199 & pi1138;
  assign n44139 = pi200 & ~n44138;
  assign n44140 = pi199 & pi1139;
  assign n44141 = ~pi200 & ~n43486;
  assign n44142 = ~n44140 & n44141;
  assign n44143 = ~n44139 & ~n44142;
  assign n44144 = n16429 & ~n44143;
  assign n44145 = pi219 & n43546;
  assign n44146 = pi211 & pi1138;
  assign n44147 = ~n44104 & ~n44146;
  assign n44148 = ~pi219 & ~n44147;
  assign n44149 = ~n44145 & ~n44148;
  assign n44150 = ~n16429 & n44149;
  assign n44151 = ~n44144 & ~n44150;
  assign n44152 = pi230 & ~n44151;
  assign n44153 = ~pi830 & n40717;
  assign n44154 = pi281 & ~n40717;
  assign n44155 = ~pi1091 & ~n44153;
  assign n44156 = ~n44154 & n44155;
  assign n44157 = pi1091 & ~n44147;
  assign n44158 = n40019 & ~n44157;
  assign n44159 = pi1138 & n40935;
  assign n44160 = ~n44114 & ~n44159;
  assign n44161 = n43449 & n44160;
  assign n44162 = ~n44158 & ~n44161;
  assign n44163 = ~n44156 & ~n44162;
  assign n44164 = ~pi830 & n40706;
  assign n44165 = pi281 & ~n40706;
  assign n44166 = ~pi1091 & ~n44164;
  assign n44167 = ~n44165 & n44166;
  assign n44168 = pi1139 & n42446;
  assign n44169 = n43520 & ~n44168;
  assign n44170 = pi199 & ~n43553;
  assign n44171 = n16429 & n44170;
  assign n44172 = ~n44169 & ~n44171;
  assign n44173 = ~n44167 & ~n44172;
  assign n44174 = ~n44163 & ~n44173;
  assign n44175 = ~pi230 & ~n44174;
  assign po438 = ~n44152 & ~n44175;
  assign n44177 = pi200 & ~n43567;
  assign n44178 = pi199 & pi1140;
  assign n44179 = ~pi200 & ~n44138;
  assign n44180 = ~n44178 & n44179;
  assign n44181 = ~n44177 & ~n44180;
  assign n44182 = n16429 & ~n44181;
  assign n44183 = pi219 & n43956;
  assign n44184 = pi211 & pi1139;
  assign n44185 = ~n43494 & ~n44184;
  assign n44186 = ~pi219 & ~n44185;
  assign n44187 = ~n44183 & ~n44186;
  assign n44188 = ~n16429 & n44187;
  assign n44189 = ~n44182 & ~n44188;
  assign n44190 = pi230 & ~n44189;
  assign n44191 = ~pi836 & n40717;
  assign n44192 = pi282 & ~n40717;
  assign n44193 = ~pi1091 & ~n44191;
  assign n44194 = ~n44192 & n44193;
  assign n44195 = pi1091 & ~n44185;
  assign n44196 = n40019 & ~n44195;
  assign n44197 = pi1139 & n40935;
  assign n44198 = ~n43523 & ~n44197;
  assign n44199 = n43449 & n44198;
  assign n44200 = ~n44196 & ~n44199;
  assign n44201 = ~n44194 & ~n44200;
  assign n44202 = ~pi836 & n40706;
  assign n44203 = pi282 & ~n40706;
  assign n44204 = ~pi1091 & ~n44202;
  assign n44205 = ~n44203 & n44204;
  assign n44206 = pi1140 & n42446;
  assign n44207 = n43520 & ~n44206;
  assign n44208 = ~pi200 & n43551;
  assign n44209 = pi199 & ~n44208;
  assign n44210 = n16429 & n44209;
  assign n44211 = ~n44207 & ~n44210;
  assign n44212 = ~n44205 & ~n44211;
  assign n44213 = ~n44201 & ~n44212;
  assign n44214 = ~pi230 & ~n44213;
  assign po439 = ~n44190 & ~n44214;
  assign n44216 = pi1147 & ~n43647;
  assign n44217 = n43709 & ~n44216;
  assign n44218 = pi1147 & ~n43450;
  assign n44219 = ~pi1149 & n43468;
  assign n44220 = ~n44218 & n44219;
  assign n44221 = pi1148 & ~n44217;
  assign n44222 = ~n44220 & n44221;
  assign n44223 = pi1149 & ~n42226;
  assign n44224 = ~n44216 & ~n44223;
  assign n44225 = ~pi1148 & ~n44224;
  assign n44226 = pi230 & ~n44225;
  assign n44227 = ~n44222 & n44226;
  assign n44228 = pi1147 & n43376;
  assign n44229 = ~pi1147 & n43430;
  assign n44230 = ~pi1148 & ~n44229;
  assign n44231 = ~n44228 & n44230;
  assign n44232 = ~pi1147 & n43426;
  assign n44233 = pi1147 & n43381;
  assign n44234 = pi1148 & ~n44233;
  assign n44235 = ~n44232 & n44234;
  assign n44236 = pi1149 & ~n44235;
  assign n44237 = ~n44231 & n44236;
  assign n44238 = pi1147 & n43336;
  assign n44239 = ~pi1147 & ~n43438;
  assign n44240 = ~pi1148 & ~n44239;
  assign n44241 = ~n44238 & n44240;
  assign n44242 = ~pi1147 & n43436;
  assign n44243 = pi1147 & n43342;
  assign n44244 = pi1148 & ~n44243;
  assign n44245 = ~n44242 & n44244;
  assign n44246 = ~pi1149 & ~n44245;
  assign n44247 = ~n44241 & n44246;
  assign n44248 = pi283 & ~n44247;
  assign n44249 = ~n44237 & n44248;
  assign n44250 = pi1147 & n43387;
  assign n44251 = ~pi1147 & n43406;
  assign n44252 = pi1149 & ~n44251;
  assign n44253 = ~n44250 & n44252;
  assign n44254 = pi1147 & n43356;
  assign n44255 = ~pi1147 & ~n43363;
  assign n44256 = ~pi1149 & ~n44255;
  assign n44257 = ~n44254 & n44256;
  assign n44258 = ~pi1148 & ~n44257;
  assign n44259 = ~n44253 & n44258;
  assign n44260 = ~pi1147 & ~n43414;
  assign n44261 = pi1147 & n43364;
  assign n44262 = ~pi1149 & ~n44261;
  assign n44263 = ~n44260 & n44262;
  assign n44264 = ~pi1147 & n43409;
  assign n44265 = pi1147 & n43394;
  assign n44266 = pi1149 & ~n44265;
  assign n44267 = ~n44264 & n44266;
  assign n44268 = pi1148 & ~n44267;
  assign n44269 = ~n44263 & n44268;
  assign n44270 = ~pi283 & ~n44259;
  assign n44271 = ~n44269 & n44270;
  assign n44272 = ~pi230 & ~n44249;
  assign n44273 = ~n44271 & n44272;
  assign po440 = ~n44227 & ~n44273;
  assign n44275 = ~pi284 & ~n42736;
  assign n44276 = pi1143 & n42736;
  assign n44277 = ~n40021 & n44276;
  assign po441 = n44275 | n44277;
  assign n44279 = n3269 & ~n10398;
  assign n44280 = ~n8044 & n44279;
  assign n44281 = pi286 & n44280;
  assign n44282 = pi288 & pi289;
  assign n44283 = n44281 & n44282;
  assign n44284 = pi285 & n44283;
  assign n44285 = pi285 & n44279;
  assign n44286 = ~n44283 & ~n44285;
  assign n44287 = ~po1038 & ~n44284;
  assign n44288 = ~n44286 & n44287;
  assign n44289 = ~po1038 & n44283;
  assign n44290 = ~pi286 & n8044;
  assign n44291 = ~pi288 & n44290;
  assign n44292 = pi285 & ~pi289;
  assign n44293 = n44291 & n44292;
  assign n44294 = pi285 & ~n44293;
  assign n44295 = ~n44289 & n44294;
  assign n44296 = ~n44288 & ~n44295;
  assign po442 = ~pi793 & ~n44296;
  assign n44298 = ~pi288 & ~n7719;
  assign n44299 = n8044 & ~n44279;
  assign n44300 = pi286 & ~n44299;
  assign n44301 = ~n44279 & n44290;
  assign n44302 = ~n44300 & ~n44301;
  assign n44303 = n44298 & ~n44302;
  assign n44304 = ~pi286 & ~n44280;
  assign n44305 = pi288 & ~n44281;
  assign n44306 = ~n44304 & n44305;
  assign n44307 = ~po1038 & ~n44303;
  assign n44308 = ~n44306 & n44307;
  assign n44309 = n8044 & n44298;
  assign n44310 = pi286 & ~n44309;
  assign n44311 = ~pi286 & n44309;
  assign n44312 = po1038 & ~n44310;
  assign n44313 = ~n44311 & n44312;
  assign n44314 = ~pi793 & ~n44313;
  assign po443 = ~n44308 & n44314;
  assign n44316 = ~pi287 & pi457;
  assign po444 = ~pi332 & ~n44316;
  assign n44318 = pi288 & ~n8044;
  assign n44319 = ~n44309 & ~n44318;
  assign po637 = ~po1038 & n44279;
  assign n44321 = ~n44319 & po637;
  assign n44322 = n44319 & ~po637;
  assign n44323 = ~pi793 & ~n44321;
  assign po445 = ~n44322 & n44323;
  assign n44325 = ~pi289 & n44305;
  assign n44326 = n44292 & n44301;
  assign n44327 = pi289 & ~n44301;
  assign n44328 = ~pi288 & ~n44326;
  assign n44329 = ~n44327 & n44328;
  assign n44330 = ~n44283 & ~n44325;
  assign n44331 = ~n44329 & n44330;
  assign n44332 = ~po1038 & ~n44331;
  assign n44333 = pi289 & ~n44291;
  assign n44334 = po1038 & ~n44293;
  assign n44335 = ~n44333 & n44334;
  assign n44336 = ~pi793 & ~n44335;
  assign po446 = ~n44332 & n44336;
  assign n44338 = ~pi290 & pi476;
  assign n44339 = ~pi476 & ~pi1048;
  assign po447 = ~n44338 & ~n44339;
  assign n44341 = ~pi291 & pi476;
  assign n44342 = ~pi476 & ~pi1049;
  assign po448 = ~n44341 & ~n44342;
  assign n44344 = ~pi292 & pi476;
  assign n44345 = ~pi476 & ~pi1084;
  assign po449 = ~n44344 & ~n44345;
  assign n44347 = ~pi293 & pi476;
  assign n44348 = ~pi476 & ~pi1059;
  assign po450 = ~n44347 & ~n44348;
  assign n44350 = ~pi294 & pi476;
  assign n44351 = ~pi476 & ~pi1072;
  assign po451 = ~n44350 & ~n44351;
  assign n44353 = ~pi295 & pi476;
  assign n44354 = ~pi476 & ~pi1053;
  assign po452 = ~n44353 & ~n44354;
  assign n44356 = ~pi296 & pi476;
  assign n44357 = ~pi476 & ~pi1037;
  assign po453 = ~n44356 & ~n44357;
  assign n44359 = ~pi297 & pi476;
  assign n44360 = ~pi476 & ~pi1044;
  assign po454 = ~n44359 & ~n44360;
  assign n44362 = ~pi478 & pi1044;
  assign n44363 = pi298 & pi478;
  assign po455 = n44362 | n44363;
  assign n44365 = pi54 & n3096;
  assign n44366 = ~pi54 & n13116;
  assign n44367 = n13375 & n44366;
  assign n44368 = ~n44365 & ~n44367;
  assign n44369 = n3243 & n8866;
  assign n44370 = ~n44368 & n44369;
  assign n44371 = ~pi39 & ~n44370;
  assign po456 = ~n11246 & ~n44371;
  assign n44373 = pi57 & ~pi59;
  assign n44374 = n10123 & n44373;
  assign n44375 = ~pi312 & n44374;
  assign n44376 = pi300 & ~n44375;
  assign n44377 = ~pi300 & n44375;
  assign n44378 = ~pi55 & ~n44377;
  assign po457 = n44376 | ~n44378;
  assign n44380 = ~pi301 & n44378;
  assign n44381 = ~pi55 & pi301;
  assign n44382 = n44377 & n44381;
  assign po458 = n44380 | n44382;
  assign n44384 = n5784 & ~po1038;
  assign n44385 = ~pi222 & ~pi223;
  assign n44386 = pi937 & ~n44385;
  assign n44387 = pi273 & n3305;
  assign n44388 = ~n44386 & ~n44387;
  assign n44389 = n44384 & n44388;
  assign n44390 = n3462 & ~n16429;
  assign n44391 = ~n44389 & ~n44390;
  assign n44392 = pi237 & ~n44391;
  assign n44393 = n5795 & ~n16429;
  assign n44394 = ~n44384 & ~n44393;
  assign n44395 = ~pi1148 & n44394;
  assign n44396 = ~n3053 & n44389;
  assign n44397 = ~pi215 & n3325;
  assign n44398 = ~pi273 & n44397;
  assign n44399 = pi833 & n8074;
  assign n44400 = ~pi937 & n44399;
  assign n44401 = ~n44398 & ~n44400;
  assign n44402 = ~n16429 & ~n44401;
  assign n44403 = ~n44396 & ~n44402;
  assign n44404 = ~n44392 & n44403;
  assign po459 = ~n44395 & n44404;
  assign n44406 = ~pi478 & pi1049;
  assign n44407 = pi303 & pi478;
  assign po460 = n44406 | n44407;
  assign n44409 = ~pi478 & pi1048;
  assign n44410 = pi304 & pi478;
  assign po461 = n44409 | n44410;
  assign n44412 = ~pi478 & pi1084;
  assign n44413 = pi305 & pi478;
  assign po462 = n44412 | n44413;
  assign n44415 = ~pi478 & pi1059;
  assign n44416 = pi306 & pi478;
  assign po463 = n44415 | n44416;
  assign n44418 = ~pi478 & pi1053;
  assign n44419 = pi307 & pi478;
  assign po464 = n44418 | n44419;
  assign n44421 = ~pi478 & pi1037;
  assign n44422 = pi308 & pi478;
  assign po465 = n44421 | n44422;
  assign n44424 = ~pi478 & pi1072;
  assign n44425 = pi309 & pi478;
  assign po466 = n44424 | n44425;
  assign n44427 = pi1147 & n44394;
  assign n44428 = ~n3461 & n44393;
  assign n44429 = pi934 & ~n3137;
  assign n44430 = pi271 & n3325;
  assign n44431 = ~n44429 & ~n44430;
  assign n44432 = n44428 & ~n44431;
  assign n44433 = pi222 & ~pi934;
  assign n44434 = ~pi271 & n3305;
  assign n44435 = ~n44433 & ~n44434;
  assign n44436 = n44384 & n44435;
  assign n44437 = ~n44390 & ~n44436;
  assign n44438 = ~n44432 & n44437;
  assign n44439 = ~n44427 & n44438;
  assign n44440 = ~pi233 & ~n44439;
  assign n44441 = n44393 & n44431;
  assign n44442 = n3101 & n16429;
  assign n44443 = n44384 & ~n44435;
  assign n44444 = pi1147 & ~n44442;
  assign n44445 = ~n44443 & n44444;
  assign n44446 = ~n44441 & n44445;
  assign n44447 = ~n3053 & n44384;
  assign n44448 = ~n44428 & ~n44447;
  assign n44449 = ~pi1147 & ~n44448;
  assign n44450 = ~n44438 & n44449;
  assign n44451 = ~n44446 & ~n44450;
  assign n44452 = pi233 & ~n44451;
  assign po467 = n44440 | n44452;
  assign n44454 = ~pi55 & ~pi311;
  assign n44455 = ~n44382 & ~n44454;
  assign n44456 = ~pi311 & n44382;
  assign po468 = ~n44455 & ~n44456;
  assign n44458 = pi312 & ~n44374;
  assign n44459 = ~n44375 & ~n44458;
  assign po469 = ~pi55 & ~n44459;
  assign n44461 = ~n10387 & ~n13410;
  assign n44462 = po740 & ~n13417;
  assign n44463 = n10147 & ~n44462;
  assign po634 = n44461 | ~n44463;
  assign n44465 = ~pi954 & po634;
  assign n44466 = pi313 & pi954;
  assign po470 = ~n44465 & ~n44466;
  assign n44468 = n6544 & n8866;
  assign n44469 = n14395 & ~n44468;
  assign n44470 = ~pi39 & ~n14453;
  assign n44471 = pi39 & ~n15248;
  assign n44472 = n3207 & ~n44471;
  assign n44473 = ~n44470 & n44472;
  assign n44474 = ~n15543 & ~n44473;
  assign n44475 = n3278 & n10144;
  assign n44476 = ~n44474 & n44475;
  assign n44477 = ~n44469 & ~n44476;
  assign n44478 = n14387 & n14388;
  assign po471 = ~n44477 & n44478;
  assign n44480 = ~pi340 & n44279;
  assign n44481 = ~po1038 & n44480;
  assign n44482 = pi315 & ~n44481;
  assign n44483 = pi1080 & n44481;
  assign po472 = n44482 | n44483;
  assign n44485 = pi316 & ~n44481;
  assign n44486 = pi1047 & n44481;
  assign po473 = n44485 | n44486;
  assign n44488 = ~pi330 & po637;
  assign n44489 = pi317 & ~n44488;
  assign n44490 = pi1078 & n44488;
  assign po474 = n44489 | n44490;
  assign n44492 = ~pi341 & n44279;
  assign n44493 = ~po1038 & n44492;
  assign n44494 = pi318 & ~n44493;
  assign n44495 = pi1074 & n44493;
  assign po475 = n44494 | n44495;
  assign n44497 = pi319 & ~n44493;
  assign n44498 = pi1072 & n44493;
  assign po476 = n44497 | n44498;
  assign n44500 = pi320 & ~n44481;
  assign n44501 = pi1048 & n44481;
  assign po477 = n44500 | n44501;
  assign n44503 = pi321 & ~n44481;
  assign n44504 = pi1058 & n44481;
  assign po478 = n44503 | n44504;
  assign n44506 = pi322 & ~n44481;
  assign n44507 = pi1051 & n44481;
  assign po479 = n44506 | n44507;
  assign n44509 = pi323 & ~n44481;
  assign n44510 = pi1065 & n44481;
  assign po480 = n44509 | n44510;
  assign n44512 = pi324 & ~n44493;
  assign n44513 = pi1086 & n44493;
  assign po481 = n44512 | n44513;
  assign n44515 = pi325 & ~n44493;
  assign n44516 = pi1063 & n44493;
  assign po482 = n44515 | n44516;
  assign n44518 = pi326 & ~n44493;
  assign n44519 = pi1057 & n44493;
  assign po483 = n44518 | n44519;
  assign n44521 = pi327 & ~n44481;
  assign n44522 = pi1040 & n44481;
  assign po484 = n44521 | n44522;
  assign n44524 = pi328 & ~n44493;
  assign n44525 = pi1058 & n44493;
  assign po485 = n44524 | n44525;
  assign n44527 = pi329 & ~n44493;
  assign n44528 = pi1043 & n44493;
  assign po486 = n44527 | n44528;
  assign n44530 = pi1092 & ~n10053;
  assign n44531 = po1038 & n44530;
  assign n44532 = ~pi330 & n44531;
  assign n44533 = ~po1038 & n44530;
  assign n44534 = ~pi330 & ~n44279;
  assign n44535 = ~n44480 & ~n44534;
  assign n44536 = n44533 & ~n44535;
  assign po487 = n44532 | n44536;
  assign n44538 = ~pi331 & n44531;
  assign n44539 = ~pi331 & ~n44279;
  assign n44540 = ~n44492 & ~n44539;
  assign n44541 = n44533 & ~n44540;
  assign po488 = n44538 | n44541;
  assign n44543 = n10979 & n13137;
  assign n44544 = ~n10979 & ~n13067;
  assign n44545 = n7459 & ~n44544;
  assign n44546 = ~pi70 & ~n44545;
  assign n44547 = pi332 & n9552;
  assign n44548 = ~n44546 & n44547;
  assign n44549 = ~n44543 & ~n44548;
  assign n44550 = ~pi39 & ~n44549;
  assign n44551 = pi39 & n10413;
  assign n44552 = ~pi38 & ~n44551;
  assign n44553 = ~n44550 & n44552;
  assign po489 = n38146 & ~n44553;
  assign n44555 = pi333 & ~n44493;
  assign n44556 = pi1040 & n44493;
  assign po490 = n44555 | n44556;
  assign n44558 = pi334 & ~n44493;
  assign n44559 = pi1065 & n44493;
  assign po491 = n44558 | n44559;
  assign n44561 = pi335 & ~n44493;
  assign n44562 = pi1069 & n44493;
  assign po492 = n44561 | n44562;
  assign n44564 = pi336 & ~n44488;
  assign n44565 = pi1070 & n44488;
  assign po493 = n44564 | n44565;
  assign n44567 = pi337 & ~n44488;
  assign n44568 = pi1044 & n44488;
  assign po494 = n44567 | n44568;
  assign n44570 = pi338 & ~n44488;
  assign n44571 = pi1072 & n44488;
  assign po495 = n44570 | n44571;
  assign n44573 = pi339 & ~n44488;
  assign n44574 = pi1086 & n44488;
  assign po496 = n44573 | n44574;
  assign n44576 = pi340 & n44531;
  assign n44577 = ~pi340 & ~n44279;
  assign n44578 = ~pi331 & n44279;
  assign n44579 = n44533 & ~n44577;
  assign n44580 = ~n44578 & n44579;
  assign po497 = ~n44576 & ~n44580;
  assign n44582 = ~pi341 & ~po637;
  assign n44583 = ~n44488 & ~n44582;
  assign po498 = n44530 & ~n44583;
  assign n44585 = pi342 & ~n44481;
  assign n44586 = pi1049 & n44481;
  assign po499 = n44585 | n44586;
  assign n44588 = pi343 & ~n44481;
  assign n44589 = pi1062 & n44481;
  assign po500 = n44588 | n44589;
  assign n44591 = pi344 & ~n44481;
  assign n44592 = pi1069 & n44481;
  assign po501 = n44591 | n44592;
  assign n44594 = pi345 & ~n44481;
  assign n44595 = pi1039 & n44481;
  assign po502 = n44594 | n44595;
  assign n44597 = pi346 & ~n44481;
  assign n44598 = pi1067 & n44481;
  assign po503 = n44597 | n44598;
  assign n44600 = pi347 & ~n44481;
  assign n44601 = pi1055 & n44481;
  assign po504 = n44600 | n44601;
  assign n44603 = pi348 & ~n44481;
  assign n44604 = pi1087 & n44481;
  assign po505 = n44603 | n44604;
  assign n44606 = pi349 & ~n44481;
  assign n44607 = pi1043 & n44481;
  assign po506 = n44606 | n44607;
  assign n44609 = pi350 & ~n44481;
  assign n44610 = pi1035 & n44481;
  assign po507 = n44609 | n44610;
  assign n44612 = pi351 & ~n44481;
  assign n44613 = pi1079 & n44481;
  assign po508 = n44612 | n44613;
  assign n44615 = pi352 & ~n44481;
  assign n44616 = pi1078 & n44481;
  assign po509 = n44615 | n44616;
  assign n44618 = pi353 & ~n44481;
  assign n44619 = pi1063 & n44481;
  assign po510 = n44618 | n44619;
  assign n44621 = pi354 & ~n44481;
  assign n44622 = pi1045 & n44481;
  assign po511 = n44621 | n44622;
  assign n44624 = pi355 & ~n44481;
  assign n44625 = pi1084 & n44481;
  assign po512 = n44624 | n44625;
  assign n44627 = pi356 & ~n44481;
  assign n44628 = pi1081 & n44481;
  assign po513 = n44627 | n44628;
  assign n44630 = pi357 & ~n44481;
  assign n44631 = pi1076 & n44481;
  assign po514 = n44630 | n44631;
  assign n44633 = pi358 & ~n44481;
  assign n44634 = pi1071 & n44481;
  assign po515 = n44633 | n44634;
  assign n44636 = pi359 & ~n44481;
  assign n44637 = pi1068 & n44481;
  assign po516 = n44636 | n44637;
  assign n44639 = pi360 & ~n44481;
  assign n44640 = pi1042 & n44481;
  assign po517 = n44639 | n44640;
  assign n44642 = pi361 & ~n44481;
  assign n44643 = pi1059 & n44481;
  assign po518 = n44642 | n44643;
  assign n44645 = pi362 & ~n44481;
  assign n44646 = pi1070 & n44481;
  assign po519 = n44645 | n44646;
  assign n44648 = pi363 & ~n44488;
  assign n44649 = pi1049 & n44488;
  assign po520 = n44648 | n44649;
  assign n44651 = pi364 & ~n44488;
  assign n44652 = pi1062 & n44488;
  assign po521 = n44651 | n44652;
  assign n44654 = pi365 & ~n44488;
  assign n44655 = pi1065 & n44488;
  assign po522 = n44654 | n44655;
  assign n44657 = pi366 & ~n44488;
  assign n44658 = pi1069 & n44488;
  assign po523 = n44657 | n44658;
  assign n44660 = pi367 & ~n44488;
  assign n44661 = pi1039 & n44488;
  assign po524 = n44660 | n44661;
  assign n44663 = pi368 & ~n44488;
  assign n44664 = pi1067 & n44488;
  assign po525 = n44663 | n44664;
  assign n44666 = pi369 & ~n44488;
  assign n44667 = pi1080 & n44488;
  assign po526 = n44666 | n44667;
  assign n44669 = pi370 & ~n44488;
  assign n44670 = pi1055 & n44488;
  assign po527 = n44669 | n44670;
  assign n44672 = pi371 & ~n44488;
  assign n44673 = pi1051 & n44488;
  assign po528 = n44672 | n44673;
  assign n44675 = pi372 & ~n44488;
  assign n44676 = pi1048 & n44488;
  assign po529 = n44675 | n44676;
  assign n44678 = pi373 & ~n44488;
  assign n44679 = pi1087 & n44488;
  assign po530 = n44678 | n44679;
  assign n44681 = pi374 & ~n44488;
  assign n44682 = pi1035 & n44488;
  assign po531 = n44681 | n44682;
  assign n44684 = pi375 & ~n44488;
  assign n44685 = pi1047 & n44488;
  assign po532 = n44684 | n44685;
  assign n44687 = pi376 & ~n44488;
  assign n44688 = pi1079 & n44488;
  assign po533 = n44687 | n44688;
  assign n44690 = pi377 & ~n44488;
  assign n44691 = pi1074 & n44488;
  assign po534 = n44690 | n44691;
  assign n44693 = pi378 & ~n44488;
  assign n44694 = pi1063 & n44488;
  assign po535 = n44693 | n44694;
  assign n44696 = pi379 & ~n44488;
  assign n44697 = pi1045 & n44488;
  assign po536 = n44696 | n44697;
  assign n44699 = pi380 & ~n44488;
  assign n44700 = pi1084 & n44488;
  assign po537 = n44699 | n44700;
  assign n44702 = pi381 & ~n44488;
  assign n44703 = pi1081 & n44488;
  assign po538 = n44702 | n44703;
  assign n44705 = pi382 & ~n44488;
  assign n44706 = pi1076 & n44488;
  assign po539 = n44705 | n44706;
  assign n44708 = pi383 & ~n44488;
  assign n44709 = pi1071 & n44488;
  assign po540 = n44708 | n44709;
  assign n44711 = pi384 & ~n44488;
  assign n44712 = pi1068 & n44488;
  assign po541 = n44711 | n44712;
  assign n44714 = pi385 & ~n44488;
  assign n44715 = pi1042 & n44488;
  assign po542 = n44714 | n44715;
  assign n44717 = pi386 & ~n44488;
  assign n44718 = pi1059 & n44488;
  assign po543 = n44717 | n44718;
  assign n44720 = pi387 & ~n44488;
  assign n44721 = pi1053 & n44488;
  assign po544 = n44720 | n44721;
  assign n44723 = pi388 & ~n44488;
  assign n44724 = pi1037 & n44488;
  assign po545 = n44723 | n44724;
  assign n44726 = pi389 & ~n44488;
  assign n44727 = pi1036 & n44488;
  assign po546 = n44726 | n44727;
  assign n44729 = pi390 & ~n44493;
  assign n44730 = pi1049 & n44493;
  assign po547 = n44729 | n44730;
  assign n44732 = pi391 & ~n44493;
  assign n44733 = pi1062 & n44493;
  assign po548 = n44732 | n44733;
  assign n44735 = pi392 & ~n44493;
  assign n44736 = pi1039 & n44493;
  assign po549 = n44735 | n44736;
  assign n44738 = pi393 & ~n44493;
  assign n44739 = pi1067 & n44493;
  assign po550 = n44738 | n44739;
  assign n44741 = pi394 & ~n44493;
  assign n44742 = pi1080 & n44493;
  assign po551 = n44741 | n44742;
  assign n44744 = pi395 & ~n44493;
  assign n44745 = pi1055 & n44493;
  assign po552 = n44744 | n44745;
  assign n44747 = pi396 & ~n44493;
  assign n44748 = pi1051 & n44493;
  assign po553 = n44747 | n44748;
  assign n44750 = pi397 & ~n44493;
  assign n44751 = pi1048 & n44493;
  assign po554 = n44750 | n44751;
  assign n44753 = pi398 & ~n44493;
  assign n44754 = pi1087 & n44493;
  assign po555 = n44753 | n44754;
  assign n44756 = pi399 & ~n44493;
  assign n44757 = pi1047 & n44493;
  assign po556 = n44756 | n44757;
  assign n44759 = pi400 & ~n44493;
  assign n44760 = pi1035 & n44493;
  assign po557 = n44759 | n44760;
  assign n44762 = pi401 & ~n44493;
  assign n44763 = pi1079 & n44493;
  assign po558 = n44762 | n44763;
  assign n44765 = pi402 & ~n44493;
  assign n44766 = pi1078 & n44493;
  assign po559 = n44765 | n44766;
  assign n44768 = pi403 & ~n44493;
  assign n44769 = pi1045 & n44493;
  assign po560 = n44768 | n44769;
  assign n44771 = pi404 & ~n44493;
  assign n44772 = pi1084 & n44493;
  assign po561 = n44771 | n44772;
  assign n44774 = pi405 & ~n44493;
  assign n44775 = pi1081 & n44493;
  assign po562 = n44774 | n44775;
  assign n44777 = pi406 & ~n44493;
  assign n44778 = pi1076 & n44493;
  assign po563 = n44777 | n44778;
  assign n44780 = pi407 & ~n44493;
  assign n44781 = pi1071 & n44493;
  assign po564 = n44780 | n44781;
  assign n44783 = pi408 & ~n44493;
  assign n44784 = pi1068 & n44493;
  assign po565 = n44783 | n44784;
  assign n44786 = pi409 & ~n44493;
  assign n44787 = pi1042 & n44493;
  assign po566 = n44786 | n44787;
  assign n44789 = pi410 & ~n44493;
  assign n44790 = pi1059 & n44493;
  assign po567 = n44789 | n44790;
  assign n44792 = pi411 & ~n44493;
  assign n44793 = pi1053 & n44493;
  assign po568 = n44792 | n44793;
  assign n44795 = pi412 & ~n44493;
  assign n44796 = pi1037 & n44493;
  assign po569 = n44795 | n44796;
  assign n44798 = pi413 & ~n44493;
  assign n44799 = pi1036 & n44493;
  assign po570 = n44798 | n44799;
  assign n44801 = ~po1038 & n44578;
  assign n44802 = pi414 & ~n44801;
  assign n44803 = pi1049 & n44801;
  assign po571 = n44802 | n44803;
  assign n44805 = pi415 & ~n44801;
  assign n44806 = pi1062 & n44801;
  assign po572 = n44805 | n44806;
  assign n44808 = pi416 & ~n44801;
  assign n44809 = pi1069 & n44801;
  assign po573 = n44808 | n44809;
  assign n44811 = pi417 & ~n44801;
  assign n44812 = pi1039 & n44801;
  assign po574 = n44811 | n44812;
  assign n44814 = pi418 & ~n44801;
  assign n44815 = pi1067 & n44801;
  assign po575 = n44814 | n44815;
  assign n44817 = pi419 & ~n44801;
  assign n44818 = pi1080 & n44801;
  assign po576 = n44817 | n44818;
  assign n44820 = pi420 & ~n44801;
  assign n44821 = pi1055 & n44801;
  assign po577 = n44820 | n44821;
  assign n44823 = pi421 & ~n44801;
  assign n44824 = pi1051 & n44801;
  assign po578 = n44823 | n44824;
  assign n44826 = pi422 & ~n44801;
  assign n44827 = pi1048 & n44801;
  assign po579 = n44826 | n44827;
  assign n44829 = pi423 & ~n44801;
  assign n44830 = pi1087 & n44801;
  assign po580 = n44829 | n44830;
  assign n44832 = pi424 & ~n44801;
  assign n44833 = pi1047 & n44801;
  assign po581 = n44832 | n44833;
  assign n44835 = pi425 & ~n44801;
  assign n44836 = pi1035 & n44801;
  assign po582 = n44835 | n44836;
  assign n44838 = pi426 & ~n44801;
  assign n44839 = pi1079 & n44801;
  assign po583 = n44838 | n44839;
  assign n44841 = pi427 & ~n44801;
  assign n44842 = pi1078 & n44801;
  assign po584 = n44841 | n44842;
  assign n44844 = pi428 & ~n44801;
  assign n44845 = pi1045 & n44801;
  assign po585 = n44844 | n44845;
  assign n44847 = pi429 & ~n44801;
  assign n44848 = pi1084 & n44801;
  assign po586 = n44847 | n44848;
  assign n44850 = pi430 & ~n44801;
  assign n44851 = pi1076 & n44801;
  assign po587 = n44850 | n44851;
  assign n44853 = pi431 & ~n44801;
  assign n44854 = pi1071 & n44801;
  assign po588 = n44853 | n44854;
  assign n44856 = pi432 & ~n44801;
  assign n44857 = pi1068 & n44801;
  assign po589 = n44856 | n44857;
  assign n44859 = pi433 & ~n44801;
  assign n44860 = pi1042 & n44801;
  assign po590 = n44859 | n44860;
  assign n44862 = pi434 & ~n44801;
  assign n44863 = pi1059 & n44801;
  assign po591 = n44862 | n44863;
  assign n44865 = pi435 & ~n44801;
  assign n44866 = pi1053 & n44801;
  assign po592 = n44865 | n44866;
  assign n44868 = pi436 & ~n44801;
  assign n44869 = pi1037 & n44801;
  assign po593 = n44868 | n44869;
  assign n44871 = pi437 & ~n44801;
  assign n44872 = pi1070 & n44801;
  assign po594 = n44871 | n44872;
  assign n44874 = pi438 & ~n44801;
  assign n44875 = pi1036 & n44801;
  assign po595 = n44874 | n44875;
  assign n44877 = pi439 & ~n44488;
  assign n44878 = pi1057 & n44488;
  assign po596 = n44877 | n44878;
  assign n44880 = pi440 & ~n44488;
  assign n44881 = pi1043 & n44488;
  assign po597 = n44880 | n44881;
  assign n44883 = pi441 & ~n44481;
  assign n44884 = pi1044 & n44481;
  assign po598 = n44883 | n44884;
  assign n44886 = pi442 & ~n44488;
  assign n44887 = pi1058 & n44488;
  assign po599 = n44886 | n44887;
  assign n44889 = pi443 & ~n44801;
  assign n44890 = pi1044 & n44801;
  assign po600 = n44889 | n44890;
  assign n44892 = pi444 & ~n44801;
  assign n44893 = pi1072 & n44801;
  assign po601 = n44892 | n44893;
  assign n44895 = pi445 & ~n44801;
  assign n44896 = pi1081 & n44801;
  assign po602 = n44895 | n44896;
  assign n44898 = pi446 & ~n44801;
  assign n44899 = pi1086 & n44801;
  assign po603 = n44898 | n44899;
  assign n44901 = pi447 & ~n44488;
  assign n44902 = pi1040 & n44488;
  assign po604 = n44901 | n44902;
  assign n44904 = pi448 & ~n44801;
  assign n44905 = pi1074 & n44801;
  assign po605 = n44904 | n44905;
  assign n44907 = pi449 & ~n44801;
  assign n44908 = pi1057 & n44801;
  assign po606 = n44907 | n44908;
  assign n44910 = pi450 & ~n44481;
  assign n44911 = pi1036 & n44481;
  assign po607 = n44910 | n44911;
  assign n44913 = pi451 & ~n44801;
  assign n44914 = pi1063 & n44801;
  assign po608 = n44913 | n44914;
  assign n44916 = pi452 & ~n44481;
  assign n44917 = pi1053 & n44481;
  assign po609 = n44916 | n44917;
  assign n44919 = pi453 & ~n44801;
  assign n44920 = pi1040 & n44801;
  assign po610 = n44919 | n44920;
  assign n44922 = pi454 & ~n44801;
  assign n44923 = pi1043 & n44801;
  assign po611 = n44922 | n44923;
  assign n44925 = pi455 & ~n44481;
  assign n44926 = pi1037 & n44481;
  assign po612 = n44925 | n44926;
  assign n44928 = pi456 & ~n44493;
  assign n44929 = pi1044 & n44493;
  assign po613 = n44928 | n44929;
  assign n44931 = pi594 & pi600;
  assign n44932 = pi597 & n44931;
  assign n44933 = pi601 & n44932;
  assign n44934 = ~pi804 & ~pi810;
  assign n44935 = ~pi595 & n44934;
  assign n44936 = ~pi599 & pi810;
  assign n44937 = pi596 & ~n44936;
  assign n44938 = pi804 & ~n44937;
  assign n44939 = pi595 & pi815;
  assign n44940 = ~n44938 & n44939;
  assign n44941 = ~n44935 & ~n44940;
  assign n44942 = n44933 & ~n44941;
  assign n44943 = pi600 & ~pi810;
  assign n44944 = pi804 & ~n44943;
  assign n44945 = ~pi601 & ~n44934;
  assign n44946 = ~pi815 & ~n44944;
  assign n44947 = ~n44945 & n44946;
  assign n44948 = ~n44942 & ~n44947;
  assign n44949 = pi605 & ~n44948;
  assign n44950 = pi990 & n44931;
  assign n44951 = ~pi815 & n44944;
  assign n44952 = n44950 & n44951;
  assign n44953 = ~n44949 & ~n44952;
  assign po614 = pi821 & ~n44953;
  assign n44955 = pi458 & ~n44481;
  assign n44956 = pi1072 & n44481;
  assign po615 = n44955 | n44956;
  assign n44958 = pi459 & ~n44801;
  assign n44959 = pi1058 & n44801;
  assign po616 = n44958 | n44959;
  assign n44961 = pi460 & ~n44481;
  assign n44962 = pi1086 & n44481;
  assign po617 = n44961 | n44962;
  assign n44964 = pi461 & ~n44481;
  assign n44965 = pi1057 & n44481;
  assign po618 = n44964 | n44965;
  assign n44967 = pi462 & ~n44481;
  assign n44968 = pi1074 & n44481;
  assign po619 = n44967 | n44968;
  assign n44970 = pi463 & ~n44493;
  assign n44971 = pi1070 & n44493;
  assign po620 = n44970 | n44971;
  assign n44973 = pi464 & ~n44801;
  assign n44974 = pi1065 & n44801;
  assign po621 = n44973 | n44974;
  assign n44976 = ~n5775 & ~n5784;
  assign n44977 = pi926 & ~n44976;
  assign n44978 = pi1157 & n44976;
  assign n44979 = ~n11371 & ~n11374;
  assign n44980 = ~pi243 & ~n44979;
  assign n44981 = ~n44977 & ~n44980;
  assign n44982 = ~n44978 & n44981;
  assign n44983 = ~pi299 & n44385;
  assign n44984 = ~n11398 & ~n44983;
  assign n44985 = ~pi243 & pi1157;
  assign n44986 = ~n44984 & ~n44985;
  assign n44987 = ~n44980 & n44986;
  assign n44988 = ~n3484 & ~n11399;
  assign n44989 = pi926 & n44985;
  assign n44990 = ~n44988 & n44989;
  assign n44991 = ~n44987 & ~n44990;
  assign n44992 = ~n44982 & n44991;
  assign n44993 = ~po1038 & ~n44992;
  assign n44994 = ~pi243 & n44397;
  assign n44995 = pi926 & n44399;
  assign n44996 = pi1157 & ~n5795;
  assign n44997 = po1038 & ~n44994;
  assign n44998 = ~n44995 & ~n44996;
  assign n44999 = n44997 & n44998;
  assign po622 = ~n44993 & ~n44999;
  assign n45001 = po1038 & ~n44397;
  assign n45002 = ~po1038 & n44979;
  assign n45003 = ~n45001 & ~n45002;
  assign n45004 = ~pi943 & ~n45003;
  assign n45005 = pi943 & n44448;
  assign n45006 = ~n45004 & ~n45005;
  assign n45007 = ~pi1151 & ~n45006;
  assign n45008 = ~n44394 & n45004;
  assign n45009 = ~n44390 & ~n44442;
  assign n45010 = pi943 & pi1151;
  assign n45011 = ~n45009 & n45010;
  assign n45012 = ~po1038 & ~n44984;
  assign n45013 = n3137 & po1038;
  assign n45014 = ~n45012 & ~n45013;
  assign n45015 = ~pi275 & ~n45014;
  assign n45016 = ~n45008 & ~n45015;
  assign n45017 = ~n45011 & n45016;
  assign po623 = ~n45007 & n45017;
  assign n45019 = pi40 & ~pi287;
  assign n45020 = n42181 & n45019;
  assign n45021 = po950 & n45020;
  assign n45022 = ~n10146 & ~n45021;
  assign n45023 = ~pi102 & ~n13345;
  assign n45024 = n8885 & n10143;
  assign n45025 = n16582 & n45024;
  assign n45026 = ~n45023 & n45025;
  assign n45027 = n16580 & n45026;
  assign n45028 = n45020 & ~n45027;
  assign n45029 = ~n45020 & n45027;
  assign n45030 = ~n45028 & ~n45029;
  assign n45031 = ~n6266 & ~n45030;
  assign n45032 = n6266 & n45027;
  assign n45033 = ~n45031 & ~n45032;
  assign n45034 = ~n7560 & ~n45033;
  assign n45035 = n7560 & ~n45030;
  assign n45036 = pi1091 & ~n45035;
  assign n45037 = ~n45034 & n45036;
  assign n45038 = ~pi1093 & ~n45033;
  assign n45039 = ~n7496 & ~n45030;
  assign n45040 = n7496 & n45027;
  assign n45041 = ~n45039 & ~n45040;
  assign n45042 = pi1093 & ~n45041;
  assign n45043 = ~pi1091 & ~n45038;
  assign n45044 = ~n45042 & n45043;
  assign n45045 = ~n45037 & ~n45044;
  assign n45046 = n3223 & n44468;
  assign n45047 = ~n45045 & n45046;
  assign po624 = ~n45022 & ~n45047;
  assign n45049 = n10181 & n11314;
  assign n45050 = pi38 & ~pi39;
  assign n45051 = n10178 & n45050;
  assign n45052 = n8948 & n45051;
  assign n45053 = pi468 & ~n45052;
  assign po625 = n45049 | n45053;
  assign n45055 = pi942 & ~n44976;
  assign n45056 = pi1156 & n44976;
  assign n45057 = ~pi263 & ~n44979;
  assign n45058 = ~n45055 & ~n45057;
  assign n45059 = ~n45056 & n45058;
  assign n45060 = ~pi263 & pi1156;
  assign n45061 = ~n44984 & ~n45060;
  assign n45062 = ~n45057 & n45061;
  assign n45063 = pi942 & n45060;
  assign n45064 = ~n44988 & n45063;
  assign n45065 = ~n45062 & ~n45064;
  assign n45066 = ~n45059 & n45065;
  assign n45067 = ~po1038 & ~n45066;
  assign n45068 = ~pi263 & n44397;
  assign n45069 = pi1156 & ~n5795;
  assign n45070 = pi942 & n44399;
  assign n45071 = po1038 & ~n45068;
  assign n45072 = ~n45069 & ~n45070;
  assign n45073 = n45071 & n45072;
  assign po626 = ~n45067 & ~n45073;
  assign n45075 = pi925 & ~n44976;
  assign n45076 = pi1155 & n44976;
  assign n45077 = pi267 & ~n44979;
  assign n45078 = ~n45075 & ~n45077;
  assign n45079 = ~n45076 & n45078;
  assign n45080 = pi267 & pi1155;
  assign n45081 = ~n44984 & ~n45080;
  assign n45082 = ~n45077 & n45081;
  assign n45083 = pi925 & n45080;
  assign n45084 = ~n44988 & n45083;
  assign n45085 = ~n45082 & ~n45084;
  assign n45086 = ~n45079 & n45085;
  assign n45087 = ~po1038 & ~n45086;
  assign n45088 = pi267 & n44397;
  assign n45089 = pi1155 & ~n5795;
  assign n45090 = pi925 & n44399;
  assign n45091 = po1038 & ~n45088;
  assign n45092 = ~n45089 & ~n45090;
  assign n45093 = n45091 & n45092;
  assign po627 = ~n45087 & ~n45093;
  assign n45095 = pi941 & ~n44976;
  assign n45096 = pi1153 & n44976;
  assign n45097 = pi253 & ~n44979;
  assign n45098 = ~n45095 & ~n45097;
  assign n45099 = ~n45096 & n45098;
  assign n45100 = pi253 & pi1153;
  assign n45101 = ~n44984 & ~n45100;
  assign n45102 = ~n45097 & n45101;
  assign n45103 = pi941 & n45100;
  assign n45104 = ~n44988 & n45103;
  assign n45105 = ~n45102 & ~n45104;
  assign n45106 = ~n45099 & n45105;
  assign n45107 = ~po1038 & ~n45106;
  assign n45108 = pi253 & n44397;
  assign n45109 = pi1153 & ~n5795;
  assign n45110 = pi941 & n44399;
  assign n45111 = po1038 & ~n45108;
  assign n45112 = ~n45109 & ~n45110;
  assign n45113 = n45111 & n45112;
  assign po628 = ~n45107 & ~n45113;
  assign n45115 = pi923 & ~n44976;
  assign n45116 = pi1154 & n44976;
  assign n45117 = pi254 & ~n44979;
  assign n45118 = ~n45115 & ~n45117;
  assign n45119 = ~n45116 & n45118;
  assign n45120 = pi254 & pi1154;
  assign n45121 = ~n44984 & ~n45120;
  assign n45122 = ~n45117 & n45121;
  assign n45123 = pi923 & n45120;
  assign n45124 = ~n44988 & n45123;
  assign n45125 = ~n45122 & ~n45124;
  assign n45126 = ~n45119 & n45125;
  assign n45127 = ~po1038 & ~n45126;
  assign n45128 = pi254 & n44397;
  assign n45129 = pi1154 & ~n5795;
  assign n45130 = pi923 & n44399;
  assign n45131 = po1038 & ~n45128;
  assign n45132 = ~n45129 & ~n45130;
  assign n45133 = n45131 & n45132;
  assign po629 = ~n45127 & ~n45133;
  assign n45135 = ~pi922 & ~n45003;
  assign n45136 = pi922 & n44448;
  assign n45137 = ~n45135 & ~n45136;
  assign n45138 = ~pi1152 & ~n45137;
  assign n45139 = ~n44394 & n45135;
  assign n45140 = pi922 & pi1152;
  assign n45141 = ~n45009 & n45140;
  assign n45142 = ~pi268 & ~n45014;
  assign n45143 = ~n45139 & ~n45142;
  assign n45144 = ~n45141 & n45143;
  assign po630 = ~n45138 & n45144;
  assign n45146 = ~pi931 & ~n45003;
  assign n45147 = pi931 & n44448;
  assign n45148 = ~n45146 & ~n45147;
  assign n45149 = ~pi1150 & ~n45148;
  assign n45150 = ~n44394 & n45146;
  assign n45151 = pi931 & pi1150;
  assign n45152 = ~n45009 & n45151;
  assign n45153 = ~pi272 & ~n45014;
  assign n45154 = ~n45150 & ~n45153;
  assign n45155 = ~n45152 & n45154;
  assign po631 = ~n45149 & n45155;
  assign n45157 = ~pi936 & ~n45003;
  assign n45158 = pi936 & n44448;
  assign n45159 = ~n45157 & ~n45158;
  assign n45160 = ~pi1149 & ~n45159;
  assign n45161 = ~n44394 & n45157;
  assign n45162 = pi936 & pi1149;
  assign n45163 = ~n45009 & n45162;
  assign n45164 = ~pi283 & ~n45014;
  assign n45165 = ~n45161 & ~n45164;
  assign n45166 = ~n45163 & n45165;
  assign po632 = ~n45160 & n45166;
  assign n45168 = pi71 & n43467;
  assign n45169 = pi71 & ~n11423;
  assign n45170 = n11423 & n13012;
  assign n45171 = n10132 & ~n11423;
  assign n45172 = n10128 & n45171;
  assign n45173 = ~n45170 & ~n45172;
  assign n45174 = n3269 & n10143;
  assign n45175 = ~n45173 & n45174;
  assign n45176 = n13020 & n45175;
  assign n45177 = ~n45169 & ~n45176;
  assign n45178 = ~po1038 & ~n45177;
  assign po633 = n45168 | n45178;
  assign po635 = pi71 & ~n43647;
  assign n45181 = pi481 & ~n34660;
  assign n45182 = pi248 & n34660;
  assign po638 = n45181 | n45182;
  assign n45184 = pi482 & ~n34676;
  assign n45185 = pi249 & n34676;
  assign po639 = n45184 | n45185;
  assign n45187 = pi483 & ~n34800;
  assign n45188 = pi242 & n34800;
  assign po640 = n45187 | n45188;
  assign n45190 = pi484 & ~n34800;
  assign n45191 = pi249 & n34800;
  assign po641 = n45190 | n45191;
  assign n45193 = pi485 & ~n35995;
  assign n45194 = pi234 & n35995;
  assign po642 = n45193 | n45194;
  assign n45196 = pi486 & ~n35995;
  assign n45197 = pi244 & n35995;
  assign po643 = n45196 | n45197;
  assign n45199 = pi487 & ~n34660;
  assign n45200 = pi246 & n34660;
  assign po644 = n45199 | n45200;
  assign n45202 = pi488 & ~n34660;
  assign n45203 = ~pi239 & n34660;
  assign po645 = ~n45202 & ~n45203;
  assign n45205 = pi489 & ~n35995;
  assign n45206 = pi242 & n35995;
  assign po646 = n45205 | n45206;
  assign n45208 = pi490 & ~n34800;
  assign n45209 = pi241 & n34800;
  assign po647 = n45208 | n45209;
  assign n45211 = pi491 & ~n34800;
  assign n45212 = pi238 & n34800;
  assign po648 = n45211 | n45212;
  assign n45214 = pi492 & ~n34800;
  assign n45215 = pi240 & n34800;
  assign po649 = n45214 | n45215;
  assign n45217 = pi493 & ~n34800;
  assign n45218 = pi244 & n34800;
  assign po650 = n45217 | n45218;
  assign n45220 = pi494 & ~n34800;
  assign n45221 = ~pi239 & n34800;
  assign po651 = ~n45220 & ~n45221;
  assign n45223 = pi495 & ~n34800;
  assign n45224 = pi235 & n34800;
  assign po652 = n45223 | n45224;
  assign n45226 = pi496 & ~n34792;
  assign n45227 = pi249 & n34792;
  assign po653 = n45226 | n45227;
  assign n45229 = pi497 & ~n34792;
  assign n45230 = ~pi239 & n34792;
  assign po654 = ~n45229 & ~n45230;
  assign n45232 = pi498 & ~n34676;
  assign n45233 = pi238 & n34676;
  assign po655 = n45232 | n45233;
  assign n45235 = pi499 & ~n34792;
  assign n45236 = pi246 & n34792;
  assign po656 = n45235 | n45236;
  assign n45238 = pi500 & ~n34792;
  assign n45239 = pi241 & n34792;
  assign po657 = n45238 | n45239;
  assign n45241 = pi501 & ~n34792;
  assign n45242 = pi248 & n34792;
  assign po658 = n45241 | n45242;
  assign n45244 = pi502 & ~n34792;
  assign n45245 = pi247 & n34792;
  assign po659 = n45244 | n45245;
  assign n45247 = pi503 & ~n34792;
  assign n45248 = pi245 & n34792;
  assign po660 = n45247 | n45248;
  assign n45250 = pi504 & ~n34785;
  assign n45251 = pi242 & n34785;
  assign po661 = n45250 | n45251;
  assign n45253 = ~n6412 & n16429;
  assign n45254 = ~n34782 & ~n45253;
  assign n45255 = ~pi234 & n45254;
  assign n45256 = n34792 & n45255;
  assign n45257 = pi505 & ~n45256;
  assign n45258 = pi234 & n34784;
  assign n45259 = ~pi505 & n34663;
  assign n45260 = n45258 & n45259;
  assign po662 = n45257 | n45260;
  assign n45262 = pi506 & ~n34785;
  assign n45263 = pi241 & n34785;
  assign po663 = n45262 | n45263;
  assign n45265 = pi507 & ~n34785;
  assign n45266 = pi238 & n34785;
  assign po664 = n45265 | n45266;
  assign n45268 = pi508 & ~n34785;
  assign n45269 = pi247 & n34785;
  assign po665 = n45268 | n45269;
  assign n45271 = pi509 & ~n34785;
  assign n45272 = pi245 & n34785;
  assign po666 = n45271 | n45272;
  assign n45274 = pi510 & ~n34660;
  assign n45275 = pi242 & n34660;
  assign po667 = n45274 | n45275;
  assign n45277 = n6606 & ~po1038;
  assign n45278 = ~n34655 & ~n45277;
  assign n45279 = ~pi234 & n45278;
  assign n45280 = n34660 & ~n45279;
  assign n45281 = pi511 & ~n34660;
  assign po668 = n45280 | n45281;
  assign n45283 = pi512 & ~n34660;
  assign n45284 = pi235 & n34660;
  assign po669 = n45283 | n45284;
  assign n45286 = pi513 & ~n34660;
  assign n45287 = pi244 & n34660;
  assign po670 = n45286 | n45287;
  assign n45289 = pi514 & ~n34660;
  assign n45290 = pi245 & n34660;
  assign po671 = n45289 | n45290;
  assign n45292 = pi515 & ~n34660;
  assign n45293 = pi240 & n34660;
  assign po672 = n45292 | n45293;
  assign n45295 = pi516 & ~n34660;
  assign n45296 = pi247 & n34660;
  assign po673 = n45295 | n45296;
  assign n45298 = pi517 & ~n34660;
  assign n45299 = pi238 & n34660;
  assign po674 = n45298 | n45299;
  assign n45301 = n34668 & n45279;
  assign n45302 = pi518 & ~n45301;
  assign n45303 = pi234 & n34659;
  assign n45304 = ~pi518 & n34663;
  assign n45305 = n45303 & n45304;
  assign po675 = n45302 | n45305;
  assign n45307 = pi519 & ~n34668;
  assign n45308 = ~pi239 & n34668;
  assign po676 = ~n45307 & ~n45308;
  assign n45310 = pi520 & ~n34668;
  assign n45311 = pi246 & n34668;
  assign po677 = n45310 | n45311;
  assign n45313 = pi521 & ~n34668;
  assign n45314 = pi248 & n34668;
  assign po678 = n45313 | n45314;
  assign n45316 = pi522 & ~n34668;
  assign n45317 = pi238 & n34668;
  assign po679 = n45316 | n45317;
  assign n45319 = n36023 & n45279;
  assign n45320 = pi523 & ~n45319;
  assign n45321 = ~pi523 & n34795;
  assign n45322 = n45303 & n45321;
  assign po680 = n45320 | n45322;
  assign n45324 = pi524 & ~n36023;
  assign n45325 = ~pi239 & n36023;
  assign po681 = ~n45324 & ~n45325;
  assign n45327 = pi525 & ~n36023;
  assign n45328 = pi245 & n36023;
  assign po682 = n45327 | n45328;
  assign n45330 = pi526 & ~n36023;
  assign n45331 = pi246 & n36023;
  assign po683 = n45330 | n45331;
  assign n45333 = pi527 & ~n36023;
  assign n45334 = pi247 & n36023;
  assign po684 = n45333 | n45334;
  assign n45336 = pi528 & ~n36023;
  assign n45337 = pi249 & n36023;
  assign po685 = n45336 | n45337;
  assign n45339 = pi529 & ~n36023;
  assign n45340 = pi238 & n36023;
  assign po686 = n45339 | n45340;
  assign n45342 = pi530 & ~n36023;
  assign n45343 = pi240 & n36023;
  assign po687 = n45342 | n45343;
  assign n45345 = pi531 & ~n34676;
  assign n45346 = pi235 & n34676;
  assign po688 = n45345 | n45346;
  assign n45348 = pi532 & ~n34676;
  assign n45349 = pi247 & n34676;
  assign po689 = n45348 | n45349;
  assign n45351 = pi533 & ~n34785;
  assign n45352 = pi235 & n34785;
  assign po690 = n45351 | n45352;
  assign n45354 = pi534 & ~n34785;
  assign n45355 = ~pi239 & n34785;
  assign po691 = ~n45354 & ~n45355;
  assign n45357 = pi535 & ~n34785;
  assign n45358 = pi240 & n34785;
  assign po692 = n45357 | n45358;
  assign n45360 = pi536 & ~n34785;
  assign n45361 = pi246 & n34785;
  assign po693 = n45360 | n45361;
  assign n45363 = pi537 & ~n34785;
  assign n45364 = pi248 & n34785;
  assign po694 = n45363 | n45364;
  assign n45366 = pi538 & ~n34785;
  assign n45367 = pi249 & n34785;
  assign po695 = n45366 | n45367;
  assign n45369 = pi539 & ~n34792;
  assign n45370 = pi242 & n34792;
  assign po696 = n45369 | n45370;
  assign n45372 = pi540 & ~n34792;
  assign n45373 = pi235 & n34792;
  assign po697 = n45372 | n45373;
  assign n45375 = pi541 & ~n34792;
  assign n45376 = pi244 & n34792;
  assign po698 = n45375 | n45376;
  assign n45378 = pi542 & ~n34792;
  assign n45379 = pi240 & n34792;
  assign po699 = n45378 | n45379;
  assign n45381 = pi543 & ~n34792;
  assign n45382 = pi238 & n34792;
  assign po700 = n45381 | n45382;
  assign n45384 = n34800 & n45255;
  assign n45385 = pi544 & ~n45384;
  assign n45386 = ~pi544 & n34795;
  assign n45387 = n45258 & n45386;
  assign po701 = n45385 | n45387;
  assign n45389 = pi545 & ~n34800;
  assign n45390 = pi245 & n34800;
  assign po702 = n45389 | n45390;
  assign n45392 = pi546 & ~n34800;
  assign n45393 = pi246 & n34800;
  assign po703 = n45392 | n45393;
  assign n45395 = pi547 & ~n34800;
  assign n45396 = pi247 & n34800;
  assign po704 = n45395 | n45396;
  assign n45398 = pi548 & ~n34800;
  assign n45399 = pi248 & n34800;
  assign po705 = n45398 | n45399;
  assign n45401 = pi549 & ~n35995;
  assign n45402 = pi235 & n35995;
  assign po706 = n45401 | n45402;
  assign n45404 = pi550 & ~n35995;
  assign n45405 = ~pi239 & n35995;
  assign po707 = ~n45404 & ~n45405;
  assign n45407 = pi551 & ~n35995;
  assign n45408 = pi240 & n35995;
  assign po708 = n45407 | n45408;
  assign n45410 = pi552 & ~n35995;
  assign n45411 = pi247 & n35995;
  assign po709 = n45410 | n45411;
  assign n45413 = pi553 & ~n35995;
  assign n45414 = pi241 & n35995;
  assign po710 = n45413 | n45414;
  assign n45416 = pi554 & ~n35995;
  assign n45417 = pi248 & n35995;
  assign po711 = n45416 | n45417;
  assign n45419 = pi555 & ~n35995;
  assign n45420 = pi249 & n35995;
  assign po712 = n45419 | n45420;
  assign n45422 = pi556 & ~n34676;
  assign n45423 = pi242 & n34676;
  assign po713 = n45422 | n45423;
  assign n45425 = n34785 & n45255;
  assign n45426 = pi557 & ~n45425;
  assign n45427 = ~pi557 & n34468;
  assign n45428 = n45258 & n45427;
  assign po714 = n45426 | n45428;
  assign n45430 = pi558 & ~n34785;
  assign n45431 = pi244 & n34785;
  assign po715 = n45430 | n45431;
  assign n45433 = pi559 & ~n34660;
  assign n45434 = pi241 & n34660;
  assign po716 = n45433 | n45434;
  assign n45436 = pi560 & ~n34676;
  assign n45437 = pi240 & n34676;
  assign po717 = n45436 | n45437;
  assign n45439 = pi561 & ~n34668;
  assign n45440 = pi247 & n34668;
  assign po718 = n45439 | n45440;
  assign n45442 = pi562 & ~n34676;
  assign n45443 = pi241 & n34676;
  assign po719 = n45442 | n45443;
  assign n45445 = pi563 & ~n35995;
  assign n45446 = pi246 & n35995;
  assign po720 = n45445 | n45446;
  assign n45448 = pi564 & ~n34676;
  assign n45449 = pi246 & n34676;
  assign po721 = n45448 | n45449;
  assign n45451 = pi565 & ~n34676;
  assign n45452 = pi248 & n34676;
  assign po722 = n45451 | n45452;
  assign n45454 = pi566 & ~n34676;
  assign n45455 = pi244 & n34676;
  assign po723 = n45454 | n45455;
  assign n45457 = pi603 & n16879;
  assign n45458 = ~n20159 & n45457;
  assign n45459 = n20170 & n45458;
  assign n45460 = ~pi567 & pi1092;
  assign n45461 = ~pi1093 & n45460;
  assign n45462 = ~pi789 & ~n45461;
  assign n45463 = ~n45459 & n45462;
  assign n45464 = ~pi619 & n45459;
  assign n45465 = ~n45461 & ~n45464;
  assign n45466 = ~pi1159 & ~n45465;
  assign n45467 = pi619 & n45459;
  assign n45468 = ~n45461 & ~n45467;
  assign n45469 = pi1159 & ~n45468;
  assign n45470 = pi789 & ~n45466;
  assign n45471 = ~n45469 & n45470;
  assign n45472 = ~n45463 & ~n45471;
  assign n45473 = pi680 & n17459;
  assign n45474 = ~n19124 & n45473;
  assign n45475 = ~n45461 & ~n45474;
  assign n45476 = n19216 & ~n45475;
  assign n45477 = ~n17626 & n45471;
  assign n45478 = n45476 & ~n45477;
  assign n45479 = ~n45472 & ~n45478;
  assign n45480 = n17905 & ~n45479;
  assign n45481 = n35144 & n45472;
  assign n45482 = ~n17627 & n45476;
  assign n45483 = pi641 & n45482;
  assign n45484 = ~n45461 & ~n45483;
  assign n45485 = n17786 & ~n45484;
  assign n45486 = ~pi641 & n45482;
  assign n45487 = ~n45461 & ~n45486;
  assign n45488 = n17787 & ~n45487;
  assign n45489 = ~n45485 & ~n45488;
  assign n45490 = ~n45481 & n45489;
  assign n45491 = pi788 & ~n45490;
  assign n45492 = ~n45480 & ~n45491;
  assign n45493 = ~n20298 & ~n45492;
  assign n45494 = ~n17904 & n45472;
  assign n45495 = n17904 & n45461;
  assign n45496 = ~n45494 & ~n45495;
  assign n45497 = n17944 & ~n45496;
  assign n45498 = n19217 & ~n45475;
  assign n45499 = pi628 & n45498;
  assign n45500 = ~n45461 & ~n45499;
  assign n45501 = pi1156 & ~n45500;
  assign n45502 = ~pi629 & ~n45501;
  assign n45503 = ~n45497 & n45502;
  assign n45504 = n17943 & ~n45496;
  assign n45505 = ~pi628 & n45498;
  assign n45506 = ~n45461 & ~n45505;
  assign n45507 = ~pi1156 & ~n45506;
  assign n45508 = pi629 & ~n45507;
  assign n45509 = ~n45504 & n45508;
  assign n45510 = pi792 & ~n45503;
  assign n45511 = ~n45509 & n45510;
  assign n45512 = ~n45493 & ~n45511;
  assign n45513 = ~pi647 & ~n45512;
  assign n45514 = ~n17698 & ~n45496;
  assign n45515 = n17698 & n45461;
  assign n45516 = ~n45514 & ~n45515;
  assign n45517 = pi647 & ~n45516;
  assign n45518 = ~pi1157 & ~n45517;
  assign n45519 = ~n45513 & n45518;
  assign n45520 = ~n19247 & n45498;
  assign n45521 = pi647 & n45520;
  assign n45522 = pi1157 & ~n45461;
  assign n45523 = ~n45521 & n45522;
  assign n45524 = ~pi630 & ~n45523;
  assign n45525 = ~n45519 & n45524;
  assign n45526 = pi647 & ~n45512;
  assign n45527 = ~pi647 & ~n45516;
  assign n45528 = pi1157 & ~n45527;
  assign n45529 = ~n45526 & n45528;
  assign n45530 = ~pi647 & n45520;
  assign n45531 = ~pi1157 & ~n45461;
  assign n45532 = ~n45530 & n45531;
  assign n45533 = pi630 & ~n45532;
  assign n45534 = ~n45529 & n45533;
  assign n45535 = ~n45525 & ~n45534;
  assign n45536 = pi787 & ~n45535;
  assign n45537 = ~pi787 & ~n45512;
  assign n45538 = ~n45536 & ~n45537;
  assign n45539 = ~pi790 & ~n45538;
  assign n45540 = ~pi644 & ~n45538;
  assign n45541 = ~n19271 & n45520;
  assign n45542 = ~n45461 & ~n45541;
  assign n45543 = pi644 & ~n45542;
  assign n45544 = ~pi715 & ~n45543;
  assign n45545 = ~n45540 & n45544;
  assign n45546 = ~n17740 & n45514;
  assign n45547 = ~pi644 & n45546;
  assign n45548 = pi715 & ~n45461;
  assign n45549 = ~n45547 & n45548;
  assign n45550 = ~n45545 & ~n45549;
  assign n45551 = ~pi1160 & ~n45550;
  assign n45552 = pi644 & n45538;
  assign n45553 = ~pi644 & n45542;
  assign n45554 = pi715 & ~n45553;
  assign n45555 = ~n45552 & n45554;
  assign n45556 = pi644 & n45546;
  assign n45557 = ~n45461 & ~n45556;
  assign n45558 = ~pi715 & ~n45557;
  assign n45559 = pi1160 & ~n45558;
  assign n45560 = ~n45555 & n45559;
  assign n45561 = pi790 & ~n45560;
  assign n45562 = ~n45551 & n45561;
  assign n45563 = ~n45539 & ~n45562;
  assign n45564 = pi230 & ~n45563;
  assign n45565 = ~pi230 & n45460;
  assign po724 = n45564 | n45565;
  assign n45567 = pi568 & ~n34676;
  assign n45568 = pi245 & n34676;
  assign po725 = n45567 | n45568;
  assign n45570 = pi569 & ~n34676;
  assign n45571 = ~pi239 & n34676;
  assign po726 = ~n45570 & ~n45571;
  assign n45573 = n34676 & n45279;
  assign n45574 = pi570 & ~n45573;
  assign n45575 = ~pi570 & n34671;
  assign n45576 = n45303 & n45575;
  assign po727 = n45574 | n45576;
  assign n45578 = pi571 & ~n36023;
  assign n45579 = pi241 & n36023;
  assign po728 = n45578 | n45579;
  assign n45581 = pi572 & ~n36023;
  assign n45582 = pi244 & n36023;
  assign po729 = n45581 | n45582;
  assign n45584 = pi573 & ~n36023;
  assign n45585 = pi242 & n36023;
  assign po730 = n45584 | n45585;
  assign n45587 = pi574 & ~n34668;
  assign n45588 = pi241 & n34668;
  assign po731 = n45587 | n45588;
  assign n45590 = pi575 & ~n36023;
  assign n45591 = pi235 & n36023;
  assign po732 = n45590 | n45591;
  assign n45593 = pi576 & ~n36023;
  assign n45594 = pi248 & n36023;
  assign po733 = n45593 | n45594;
  assign n45596 = pi577 & ~n35995;
  assign n45597 = pi238 & n35995;
  assign po734 = n45596 | n45597;
  assign n45599 = pi578 & ~n34668;
  assign n45600 = pi249 & n34668;
  assign po735 = n45599 | n45600;
  assign n45602 = pi579 & ~n34660;
  assign n45603 = pi249 & n34660;
  assign po736 = n45602 | n45603;
  assign n45605 = pi580 & ~n35995;
  assign n45606 = pi245 & n35995;
  assign po737 = n45605 | n45606;
  assign n45608 = pi581 & ~n34668;
  assign n45609 = pi235 & n34668;
  assign po738 = n45608 | n45609;
  assign n45611 = pi582 & ~n34668;
  assign n45612 = pi240 & n34668;
  assign po739 = n45611 | n45612;
  assign n45614 = pi584 & ~n34668;
  assign n45615 = pi245 & n34668;
  assign po741 = n45614 | n45615;
  assign n45617 = pi585 & ~n34668;
  assign n45618 = pi244 & n34668;
  assign po742 = n45617 | n45618;
  assign n45620 = pi586 & ~n34668;
  assign n45621 = pi242 & n34668;
  assign po743 = n45620 | n45621;
  assign n45623 = ~pi230 & pi587;
  assign n45624 = pi230 & n16842;
  assign n45625 = ~n20159 & n45624;
  assign n45626 = ~n35520 & n45625;
  assign n45627 = n20171 & n45626;
  assign n45628 = n30702 & n45627;
  assign po744 = n45623 | n45628;
  assign n45630 = ~pi123 & n12178;
  assign n45631 = ~pi588 & ~n45630;
  assign n45632 = ~pi591 & n45630;
  assign n45633 = n44530 & ~n45631;
  assign po745 = ~n45632 & n45633;
  assign n45635 = ~pi204 & n45254;
  assign n45636 = ~pi201 & n45278;
  assign n45637 = pi233 & ~n45635;
  assign n45638 = ~n45636 & n45637;
  assign n45639 = ~pi205 & n45254;
  assign n45640 = ~pi202 & n45278;
  assign n45641 = ~pi233 & ~n45639;
  assign n45642 = ~n45640 & n45641;
  assign n45643 = ~n45638 & ~n45642;
  assign n45644 = pi237 & ~n45643;
  assign n45645 = ~pi206 & n45254;
  assign n45646 = ~pi220 & n45278;
  assign n45647 = pi233 & ~n45645;
  assign n45648 = ~n45646 & n45647;
  assign n45649 = ~pi218 & n45254;
  assign n45650 = ~pi203 & n45278;
  assign n45651 = ~pi233 & ~n45649;
  assign n45652 = ~n45650 & n45651;
  assign n45653 = ~n45648 & ~n45652;
  assign n45654 = ~pi237 & ~n45653;
  assign po746 = ~n45644 & ~n45654;
  assign n45656 = pi588 & n45630;
  assign n45657 = pi590 & ~n45630;
  assign n45658 = n44530 & ~n45656;
  assign po747 = n45657 | ~n45658;
  assign n45660 = ~pi591 & ~n45630;
  assign n45661 = ~pi592 & n45630;
  assign n45662 = n44530 & ~n45660;
  assign po748 = ~n45661 & n45662;
  assign n45664 = ~pi592 & ~n45630;
  assign n45665 = ~pi590 & n45630;
  assign n45666 = n44530 & ~n45664;
  assign po749 = ~n45665 & n45666;
  assign n45668 = ~pi557 & ~n45255;
  assign n45669 = pi234 & n45254;
  assign n45670 = pi557 & ~n45669;
  assign n45671 = pi246 & pi536;
  assign n45672 = ~pi246 & ~pi536;
  assign n45673 = ~n45671 & ~n45672;
  assign n45674 = ~n45668 & ~n45673;
  assign n45675 = ~n45670 & n45674;
  assign n45676 = ~pi538 & n45675;
  assign n45677 = ~pi249 & ~n45676;
  assign n45678 = pi538 & n45675;
  assign n45679 = pi249 & ~n45678;
  assign n45680 = ~n45677 & ~n45679;
  assign n45681 = ~pi537 & n45680;
  assign n45682 = ~pi248 & ~n45681;
  assign n45683 = pi537 & n45680;
  assign n45684 = pi248 & ~n45683;
  assign n45685 = ~n45682 & ~n45684;
  assign n45686 = pi241 & pi506;
  assign n45687 = ~pi241 & ~pi506;
  assign n45688 = ~n45686 & ~n45687;
  assign n45689 = n45685 & ~n45688;
  assign n45690 = pi240 & pi535;
  assign n45691 = ~pi240 & ~pi535;
  assign n45692 = ~n45690 & ~n45691;
  assign n45693 = n45689 & ~n45692;
  assign n45694 = pi534 & n45693;
  assign n45695 = ~pi239 & ~n45694;
  assign n45696 = ~pi534 & n45693;
  assign n45697 = pi239 & ~n45696;
  assign n45698 = ~n45695 & ~n45697;
  assign n45699 = pi504 & n45698;
  assign n45700 = pi242 & ~n45699;
  assign n45701 = ~pi504 & n45698;
  assign n45702 = ~pi242 & ~n45701;
  assign n45703 = ~n45700 & ~n45702;
  assign n45704 = pi533 & n45703;
  assign n45705 = pi235 & ~n45704;
  assign n45706 = ~pi533 & n45703;
  assign n45707 = ~pi235 & ~n45706;
  assign n45708 = ~n45705 & ~n45707;
  assign n45709 = pi558 & n45708;
  assign n45710 = pi244 & ~n45709;
  assign n45711 = ~pi558 & n45708;
  assign n45712 = ~pi244 & ~n45711;
  assign n45713 = ~n45710 & ~n45712;
  assign n45714 = pi509 & n45713;
  assign n45715 = pi245 & ~n45714;
  assign n45716 = ~pi509 & n45713;
  assign n45717 = ~pi245 & ~n45716;
  assign n45718 = ~n45715 & ~n45717;
  assign n45719 = pi508 & n45718;
  assign n45720 = pi247 & ~n45719;
  assign n45721 = pi248 & pi481;
  assign n45722 = ~pi248 & ~pi481;
  assign n45723 = ~n45721 & ~n45722;
  assign n45724 = ~pi511 & ~n45279;
  assign n45725 = pi234 & n45278;
  assign n45726 = pi511 & ~n45725;
  assign n45727 = pi246 & pi487;
  assign n45728 = ~pi246 & ~pi487;
  assign n45729 = ~n45727 & ~n45728;
  assign n45730 = ~n45724 & ~n45729;
  assign n45731 = ~n45726 & n45730;
  assign n45732 = ~pi249 & ~pi579;
  assign n45733 = pi249 & pi579;
  assign n45734 = ~n45732 & ~n45733;
  assign n45735 = n45731 & ~n45734;
  assign n45736 = ~n45723 & n45735;
  assign n45737 = pi559 & n45736;
  assign n45738 = pi241 & ~n45737;
  assign n45739 = ~pi559 & n45736;
  assign n45740 = ~pi241 & ~n45739;
  assign n45741 = ~n45738 & ~n45740;
  assign n45742 = pi515 & n45741;
  assign n45743 = pi240 & ~n45742;
  assign n45744 = ~pi579 & ~n45735;
  assign n45745 = ~n45677 & n45731;
  assign n45746 = pi579 & ~n45745;
  assign n45747 = ~n45744 & ~n45746;
  assign n45748 = ~n45680 & ~n45747;
  assign n45749 = ~pi537 & ~n45748;
  assign n45750 = pi537 & n45735;
  assign n45751 = ~pi248 & ~n45750;
  assign n45752 = ~n45749 & n45751;
  assign n45753 = ~n45684 & ~n45752;
  assign n45754 = ~pi481 & ~n45753;
  assign n45755 = pi537 & ~n45748;
  assign n45756 = ~pi537 & n45735;
  assign n45757 = pi248 & ~n45756;
  assign n45758 = ~n45755 & n45757;
  assign n45759 = ~n45682 & ~n45758;
  assign n45760 = pi481 & ~n45759;
  assign n45761 = ~n45754 & ~n45760;
  assign n45762 = ~pi559 & n45761;
  assign n45763 = pi559 & n45685;
  assign n45764 = ~pi241 & ~n45763;
  assign n45765 = ~n45762 & n45764;
  assign n45766 = ~n45738 & ~n45765;
  assign n45767 = ~pi506 & ~n45766;
  assign n45768 = pi559 & n45761;
  assign n45769 = ~pi559 & n45685;
  assign n45770 = pi241 & ~n45769;
  assign n45771 = ~n45768 & n45770;
  assign n45772 = ~n45740 & ~n45771;
  assign n45773 = pi506 & ~n45772;
  assign n45774 = ~n45767 & ~n45773;
  assign n45775 = ~pi515 & n45774;
  assign n45776 = pi515 & n45689;
  assign n45777 = ~pi240 & ~n45776;
  assign n45778 = ~n45775 & n45777;
  assign n45779 = ~n45743 & ~n45778;
  assign n45780 = ~pi535 & ~n45779;
  assign n45781 = ~pi515 & n45741;
  assign n45782 = ~pi240 & ~n45781;
  assign n45783 = pi515 & n45774;
  assign n45784 = ~pi515 & n45689;
  assign n45785 = pi240 & ~n45784;
  assign n45786 = ~n45783 & n45785;
  assign n45787 = ~n45782 & ~n45786;
  assign n45788 = pi535 & ~n45787;
  assign n45789 = ~n45780 & ~n45788;
  assign n45790 = ~pi534 & n45789;
  assign n45791 = ~n45743 & ~n45782;
  assign n45792 = pi534 & n45791;
  assign n45793 = pi239 & ~n45792;
  assign n45794 = ~n45790 & n45793;
  assign n45795 = ~n45695 & ~n45794;
  assign n45796 = ~pi488 & ~n45795;
  assign n45797 = pi534 & n45789;
  assign n45798 = ~pi534 & n45791;
  assign n45799 = ~pi239 & ~n45798;
  assign n45800 = ~n45797 & n45799;
  assign n45801 = ~n45697 & ~n45800;
  assign n45802 = pi488 & ~n45801;
  assign n45803 = ~n45796 & ~n45802;
  assign n45804 = ~pi504 & n45803;
  assign n45805 = ~pi239 & pi488;
  assign n45806 = pi239 & ~pi488;
  assign n45807 = ~n45805 & ~n45806;
  assign n45808 = n45791 & ~n45807;
  assign n45809 = pi504 & n45808;
  assign n45810 = ~pi242 & ~n45809;
  assign n45811 = ~n45804 & n45810;
  assign n45812 = ~n45700 & ~n45811;
  assign n45813 = ~pi510 & ~n45812;
  assign n45814 = pi504 & n45803;
  assign n45815 = ~pi504 & n45808;
  assign n45816 = pi242 & ~n45815;
  assign n45817 = ~n45814 & n45816;
  assign n45818 = ~n45702 & ~n45817;
  assign n45819 = pi510 & ~n45818;
  assign n45820 = ~n45813 & ~n45819;
  assign n45821 = ~pi533 & n45820;
  assign n45822 = pi242 & pi510;
  assign n45823 = ~pi242 & ~pi510;
  assign n45824 = ~n45822 & ~n45823;
  assign n45825 = n45808 & ~n45824;
  assign n45826 = pi533 & n45825;
  assign n45827 = ~pi235 & ~n45826;
  assign n45828 = ~n45821 & n45827;
  assign n45829 = ~n45705 & ~n45828;
  assign n45830 = ~pi512 & ~n45829;
  assign n45831 = pi533 & n45820;
  assign n45832 = ~pi533 & n45825;
  assign n45833 = pi235 & ~n45832;
  assign n45834 = ~n45831 & n45833;
  assign n45835 = ~n45707 & ~n45834;
  assign n45836 = pi512 & ~n45835;
  assign n45837 = ~n45830 & ~n45836;
  assign n45838 = ~pi558 & n45837;
  assign n45839 = pi235 & pi512;
  assign n45840 = ~pi235 & ~pi512;
  assign n45841 = ~n45839 & ~n45840;
  assign n45842 = n45825 & ~n45841;
  assign n45843 = pi558 & n45842;
  assign n45844 = ~pi244 & ~n45843;
  assign n45845 = ~n45838 & n45844;
  assign n45846 = ~n45710 & ~n45845;
  assign n45847 = ~pi513 & ~n45846;
  assign n45848 = pi558 & n45837;
  assign n45849 = ~pi558 & n45842;
  assign n45850 = pi244 & ~n45849;
  assign n45851 = ~n45848 & n45850;
  assign n45852 = ~n45712 & ~n45851;
  assign n45853 = pi513 & ~n45852;
  assign n45854 = ~n45847 & ~n45853;
  assign n45855 = ~pi509 & n45854;
  assign n45856 = pi244 & pi513;
  assign n45857 = ~pi244 & ~pi513;
  assign n45858 = ~n45856 & ~n45857;
  assign n45859 = n45842 & ~n45858;
  assign n45860 = pi509 & n45859;
  assign n45861 = ~pi245 & ~n45860;
  assign n45862 = ~n45855 & n45861;
  assign n45863 = ~n45715 & ~n45862;
  assign n45864 = ~pi514 & ~n45863;
  assign n45865 = pi509 & n45854;
  assign n45866 = ~pi509 & n45859;
  assign n45867 = pi245 & ~n45866;
  assign n45868 = ~n45865 & n45867;
  assign n45869 = ~n45717 & ~n45868;
  assign n45870 = pi514 & ~n45869;
  assign n45871 = ~n45864 & ~n45870;
  assign n45872 = ~pi508 & n45871;
  assign n45873 = pi245 & pi514;
  assign n45874 = ~pi245 & ~pi514;
  assign n45875 = ~n45873 & ~n45874;
  assign n45876 = n45859 & ~n45875;
  assign n45877 = pi508 & n45876;
  assign n45878 = ~pi247 & ~n45877;
  assign n45879 = ~n45872 & n45878;
  assign n45880 = ~n45720 & ~n45879;
  assign n45881 = ~pi516 & ~n45880;
  assign n45882 = ~pi508 & n45718;
  assign n45883 = ~pi247 & ~n45882;
  assign n45884 = pi508 & n45871;
  assign n45885 = ~pi508 & n45876;
  assign n45886 = pi247 & ~n45885;
  assign n45887 = ~n45884 & n45886;
  assign n45888 = ~n45883 & ~n45887;
  assign n45889 = pi516 & ~n45888;
  assign n45890 = ~n45881 & ~n45889;
  assign n45891 = ~pi238 & n45890;
  assign n45892 = ~pi517 & ~n45891;
  assign n45893 = ~n45720 & ~n45883;
  assign n45894 = ~pi238 & n45893;
  assign n45895 = pi247 & pi516;
  assign n45896 = ~pi247 & ~pi516;
  assign n45897 = ~n45895 & ~n45896;
  assign n45898 = n45876 & ~n45897;
  assign n45899 = pi238 & n45898;
  assign n45900 = pi517 & ~n45899;
  assign n45901 = ~n45894 & n45900;
  assign n45902 = ~pi507 & ~n45901;
  assign n45903 = ~n45892 & n45902;
  assign n45904 = pi238 & n45890;
  assign n45905 = pi517 & ~n45904;
  assign n45906 = pi238 & n45893;
  assign n45907 = ~pi238 & n45898;
  assign n45908 = ~pi517 & ~n45907;
  assign n45909 = ~n45906 & n45908;
  assign n45910 = pi507 & ~n45909;
  assign n45911 = ~n45905 & n45910;
  assign n45912 = ~n45903 & ~n45911;
  assign n45913 = pi233 & ~n45912;
  assign n45914 = ~pi247 & ~pi561;
  assign n45915 = pi505 & ~n45669;
  assign n45916 = ~pi505 & ~n45255;
  assign n45917 = pi240 & pi542;
  assign n45918 = ~pi240 & ~pi542;
  assign n45919 = ~n45917 & ~n45918;
  assign n45920 = pi249 & ~pi496;
  assign n45921 = ~pi249 & pi496;
  assign n45922 = ~pi246 & ~pi499;
  assign n45923 = pi246 & pi499;
  assign n45924 = ~n45922 & ~n45923;
  assign n45925 = ~pi241 & ~pi500;
  assign n45926 = pi241 & pi500;
  assign n45927 = ~n45925 & ~n45926;
  assign n45928 = ~pi248 & ~pi501;
  assign n45929 = pi248 & pi501;
  assign n45930 = ~n45928 & ~n45929;
  assign n45931 = ~n45920 & ~n45921;
  assign n45932 = ~n45919 & n45931;
  assign n45933 = ~n45924 & ~n45927;
  assign n45934 = ~n45930 & n45933;
  assign n45935 = n45932 & n45934;
  assign n45936 = ~n45915 & n45935;
  assign n45937 = ~n45916 & n45936;
  assign n45938 = pi497 & n45937;
  assign n45939 = ~pi239 & ~n45938;
  assign n45940 = ~pi497 & n45937;
  assign n45941 = pi239 & ~n45940;
  assign n45942 = ~n45939 & ~n45941;
  assign n45943 = pi539 & n45942;
  assign n45944 = pi242 & ~n45943;
  assign n45945 = ~pi539 & n45942;
  assign n45946 = ~pi242 & ~n45945;
  assign n45947 = ~n45944 & ~n45946;
  assign n45948 = pi540 & n45947;
  assign n45949 = pi235 & ~n45948;
  assign n45950 = ~pi540 & n45947;
  assign n45951 = ~pi235 & ~n45950;
  assign n45952 = ~n45949 & ~n45951;
  assign n45953 = pi244 & pi541;
  assign n45954 = ~pi244 & ~pi541;
  assign n45955 = ~n45953 & ~n45954;
  assign n45956 = n45952 & ~n45955;
  assign n45957 = pi245 & pi503;
  assign n45958 = ~pi245 & ~pi503;
  assign n45959 = ~n45957 & ~n45958;
  assign n45960 = n45956 & ~n45959;
  assign n45961 = ~pi502 & n45960;
  assign n45962 = ~pi247 & ~n45961;
  assign n45963 = ~n45914 & ~n45962;
  assign n45964 = pi518 & ~n45725;
  assign n45965 = ~pi518 & ~n45279;
  assign n45966 = pi249 & ~pi578;
  assign n45967 = ~pi249 & pi578;
  assign n45968 = pi248 & ~pi521;
  assign n45969 = ~pi248 & pi521;
  assign n45970 = pi241 & pi574;
  assign n45971 = ~pi241 & ~pi574;
  assign n45972 = ~n45970 & ~n45971;
  assign n45973 = pi246 & ~pi520;
  assign n45974 = ~pi246 & pi520;
  assign n45975 = ~n45966 & ~n45967;
  assign n45976 = ~n45968 & ~n45969;
  assign n45977 = ~n45973 & ~n45974;
  assign n45978 = n45976 & n45977;
  assign n45979 = ~n45972 & n45975;
  assign n45980 = n45978 & n45979;
  assign n45981 = ~n45964 & n45980;
  assign n45982 = ~n45965 & n45981;
  assign n45983 = pi582 & n45982;
  assign n45984 = pi240 & ~n45983;
  assign n45985 = ~pi582 & n45982;
  assign n45986 = ~pi240 & ~n45985;
  assign n45987 = pi235 & pi581;
  assign n45988 = ~pi235 & ~pi581;
  assign n45989 = ~n45987 & ~n45988;
  assign n45990 = ~pi239 & pi519;
  assign n45991 = pi239 & ~pi519;
  assign n45992 = ~n45990 & ~n45991;
  assign n45993 = pi242 & pi586;
  assign n45994 = ~pi242 & ~pi586;
  assign n45995 = ~n45993 & ~n45994;
  assign n45996 = ~n45989 & ~n45992;
  assign n45997 = ~n45995 & n45996;
  assign n45998 = ~n45984 & n45997;
  assign n45999 = ~n45986 & n45998;
  assign n46000 = pi585 & n45999;
  assign n46001 = pi244 & ~n46000;
  assign n46002 = ~pi585 & n45999;
  assign n46003 = ~pi244 & ~n46002;
  assign n46004 = ~n46001 & ~n46003;
  assign n46005 = pi584 & n46004;
  assign n46006 = pi245 & ~n46005;
  assign n46007 = ~n45952 & n46003;
  assign n46008 = ~n46001 & ~n46007;
  assign n46009 = ~pi541 & ~n46008;
  assign n46010 = ~n45952 & n46001;
  assign n46011 = ~n46003 & ~n46010;
  assign n46012 = pi541 & ~n46011;
  assign n46013 = ~n46009 & ~n46012;
  assign n46014 = ~pi584 & n46013;
  assign n46015 = pi584 & n45956;
  assign n46016 = ~pi245 & ~n46015;
  assign n46017 = ~n46014 & n46016;
  assign n46018 = ~n46006 & ~n46017;
  assign n46019 = ~pi503 & ~n46018;
  assign n46020 = ~pi584 & n46004;
  assign n46021 = ~pi245 & ~n46020;
  assign n46022 = pi584 & n46013;
  assign n46023 = ~pi584 & n45956;
  assign n46024 = pi245 & ~n46023;
  assign n46025 = ~n46022 & n46024;
  assign n46026 = ~n46021 & ~n46025;
  assign n46027 = pi503 & ~n46026;
  assign n46028 = ~n46019 & ~n46027;
  assign n46029 = ~pi502 & ~n46028;
  assign n46030 = ~n46006 & ~n46021;
  assign n46031 = pi502 & ~n46030;
  assign n46032 = ~pi561 & ~n46031;
  assign n46033 = ~n46029 & n46032;
  assign n46034 = ~n45963 & ~n46033;
  assign n46035 = pi247 & pi561;
  assign n46036 = pi502 & n45960;
  assign n46037 = pi247 & ~n46036;
  assign n46038 = ~n46035 & ~n46037;
  assign n46039 = pi502 & ~n46028;
  assign n46040 = ~pi502 & ~n46030;
  assign n46041 = pi561 & ~n46040;
  assign n46042 = ~n46039 & n46041;
  assign n46043 = ~n46038 & ~n46042;
  assign n46044 = ~n46034 & ~n46043;
  assign n46045 = ~pi238 & n46044;
  assign n46046 = ~pi522 & ~n46045;
  assign n46047 = ~n45962 & ~n46037;
  assign n46048 = ~pi238 & n46047;
  assign n46049 = ~n45914 & ~n46035;
  assign n46050 = n46030 & ~n46049;
  assign n46051 = pi238 & n46050;
  assign n46052 = pi522 & ~n46051;
  assign n46053 = ~n46048 & n46052;
  assign n46054 = ~pi543 & ~n46053;
  assign n46055 = ~n46046 & n46054;
  assign n46056 = pi238 & n46044;
  assign n46057 = pi522 & ~n46056;
  assign n46058 = pi238 & n46047;
  assign n46059 = ~pi238 & n46050;
  assign n46060 = ~pi522 & ~n46059;
  assign n46061 = ~n46058 & n46060;
  assign n46062 = pi543 & ~n46061;
  assign n46063 = ~n46057 & n46062;
  assign n46064 = ~n46055 & ~n46063;
  assign n46065 = ~pi233 & ~n46064;
  assign n46066 = pi237 & ~n46065;
  assign n46067 = ~n45913 & n46066;
  assign n46068 = pi485 & ~n45669;
  assign n46069 = ~pi485 & ~n45255;
  assign n46070 = pi249 & ~pi555;
  assign n46071 = ~pi249 & pi555;
  assign n46072 = pi241 & ~pi553;
  assign n46073 = ~pi241 & pi553;
  assign n46074 = pi240 & pi551;
  assign n46075 = ~pi240 & ~pi551;
  assign n46076 = ~n46074 & ~n46075;
  assign n46077 = pi248 & ~pi554;
  assign n46078 = ~pi248 & pi554;
  assign n46079 = ~pi246 & pi563;
  assign n46080 = pi246 & ~pi563;
  assign n46081 = ~n46070 & ~n46071;
  assign n46082 = ~n46072 & ~n46073;
  assign n46083 = ~n46077 & ~n46078;
  assign n46084 = ~n46079 & ~n46080;
  assign n46085 = n46083 & n46084;
  assign n46086 = n46081 & n46082;
  assign n46087 = ~n46076 & n46086;
  assign n46088 = n46085 & n46087;
  assign n46089 = ~n46068 & n46088;
  assign n46090 = ~n46069 & n46089;
  assign n46091 = pi550 & n46090;
  assign n46092 = ~pi239 & ~n46091;
  assign n46093 = ~pi550 & n46090;
  assign n46094 = pi239 & ~n46093;
  assign n46095 = ~n46092 & ~n46094;
  assign n46096 = ~pi489 & n46095;
  assign n46097 = ~pi242 & ~n46096;
  assign n46098 = pi489 & n46095;
  assign n46099 = pi242 & ~n46098;
  assign n46100 = ~n46097 & ~n46099;
  assign n46101 = pi549 & n46100;
  assign n46102 = pi235 & ~n46101;
  assign n46103 = ~pi549 & n46100;
  assign n46104 = ~pi235 & ~n46103;
  assign n46105 = ~n46102 & ~n46104;
  assign n46106 = pi486 & n46105;
  assign n46107 = pi244 & ~n46106;
  assign n46108 = ~pi486 & n46105;
  assign n46109 = ~pi244 & ~n46108;
  assign n46110 = ~n46107 & ~n46109;
  assign n46111 = pi245 & pi580;
  assign n46112 = ~pi245 & ~pi580;
  assign n46113 = ~n46111 & ~n46112;
  assign n46114 = n46110 & ~n46113;
  assign n46115 = pi552 & n46114;
  assign n46116 = pi247 & ~n46115;
  assign n46117 = ~pi242 & ~pi556;
  assign n46118 = pi242 & pi556;
  assign n46119 = ~n46117 & ~n46118;
  assign n46120 = pi570 & ~n45725;
  assign n46121 = ~pi570 & ~n45279;
  assign n46122 = pi241 & pi562;
  assign n46123 = ~pi241 & ~pi562;
  assign n46124 = ~n46122 & ~n46123;
  assign n46125 = ~pi249 & pi482;
  assign n46126 = ~pi246 & pi564;
  assign n46127 = pi249 & ~pi482;
  assign n46128 = ~n46125 & ~n46126;
  assign n46129 = ~n46127 & n46128;
  assign n46130 = ~n46124 & n46129;
  assign n46131 = ~n46120 & n46130;
  assign n46132 = ~n46121 & n46131;
  assign n46133 = pi240 & pi560;
  assign n46134 = ~pi240 & ~pi560;
  assign n46135 = ~n46133 & ~n46134;
  assign n46136 = pi246 & ~pi564;
  assign n46137 = pi248 & ~pi565;
  assign n46138 = ~pi248 & pi565;
  assign n46139 = ~n46136 & ~n46137;
  assign n46140 = ~n46138 & n46139;
  assign n46141 = ~n46135 & n46140;
  assign n46142 = n46132 & n46141;
  assign n46143 = ~pi240 & ~n46142;
  assign n46144 = pi560 & n46140;
  assign n46145 = n46132 & n46144;
  assign n46146 = pi240 & ~n46145;
  assign n46147 = ~n46143 & ~n46146;
  assign n46148 = ~pi239 & pi569;
  assign n46149 = pi239 & ~pi569;
  assign n46150 = ~n46148 & ~n46149;
  assign n46151 = n46147 & ~n46150;
  assign n46152 = ~n46119 & n46151;
  assign n46153 = pi235 & pi531;
  assign n46154 = ~pi235 & ~pi531;
  assign n46155 = ~n46153 & ~n46154;
  assign n46156 = n46152 & ~n46155;
  assign n46157 = pi244 & pi566;
  assign n46158 = ~pi244 & ~pi566;
  assign n46159 = ~n46157 & ~n46158;
  assign n46160 = n46156 & ~n46159;
  assign n46161 = pi568 & n46160;
  assign n46162 = pi245 & ~n46161;
  assign n46163 = ~n46097 & ~n46117;
  assign n46164 = pi569 & ~n46094;
  assign n46165 = n46147 & n46164;
  assign n46166 = n46142 & n46149;
  assign n46167 = ~n46095 & ~n46166;
  assign n46168 = ~n46165 & n46167;
  assign n46169 = ~pi489 & n46168;
  assign n46170 = pi489 & ~n46151;
  assign n46171 = ~pi556 & ~n46170;
  assign n46172 = ~n46169 & n46171;
  assign n46173 = ~n46163 & ~n46172;
  assign n46174 = ~n46099 & ~n46118;
  assign n46175 = pi489 & n46168;
  assign n46176 = ~pi489 & ~n46151;
  assign n46177 = pi556 & ~n46176;
  assign n46178 = ~n46175 & n46177;
  assign n46179 = ~n46174 & ~n46178;
  assign n46180 = ~n46173 & ~n46179;
  assign n46181 = ~pi549 & n46180;
  assign n46182 = pi549 & n46152;
  assign n46183 = ~pi235 & ~n46182;
  assign n46184 = ~n46181 & n46183;
  assign n46185 = ~n46102 & ~n46184;
  assign n46186 = ~pi531 & ~n46185;
  assign n46187 = pi549 & n46180;
  assign n46188 = ~pi549 & n46152;
  assign n46189 = pi235 & ~n46188;
  assign n46190 = ~n46187 & n46189;
  assign n46191 = ~n46104 & ~n46190;
  assign n46192 = pi531 & ~n46191;
  assign n46193 = ~n46186 & ~n46192;
  assign n46194 = ~pi486 & n46193;
  assign n46195 = pi486 & n46156;
  assign n46196 = ~pi244 & ~n46195;
  assign n46197 = ~n46194 & n46196;
  assign n46198 = ~n46107 & ~n46197;
  assign n46199 = ~pi566 & ~n46198;
  assign n46200 = pi486 & n46193;
  assign n46201 = ~pi486 & n46156;
  assign n46202 = pi244 & ~n46201;
  assign n46203 = ~n46200 & n46202;
  assign n46204 = ~n46109 & ~n46203;
  assign n46205 = pi566 & ~n46204;
  assign n46206 = ~n46199 & ~n46205;
  assign n46207 = ~pi568 & n46206;
  assign n46208 = pi568 & n46110;
  assign n46209 = ~pi245 & ~n46208;
  assign n46210 = ~n46207 & n46209;
  assign n46211 = ~n46162 & ~n46210;
  assign n46212 = ~pi580 & ~n46211;
  assign n46213 = ~pi568 & n46160;
  assign n46214 = ~pi245 & ~n46213;
  assign n46215 = pi568 & n46206;
  assign n46216 = ~pi568 & n46110;
  assign n46217 = pi245 & ~n46216;
  assign n46218 = ~n46215 & n46217;
  assign n46219 = ~n46214 & ~n46218;
  assign n46220 = pi580 & ~n46219;
  assign n46221 = ~n46212 & ~n46220;
  assign n46222 = ~pi552 & n46221;
  assign n46223 = ~n46162 & ~n46214;
  assign n46224 = pi552 & n46223;
  assign n46225 = ~pi247 & ~n46224;
  assign n46226 = ~n46222 & n46225;
  assign n46227 = ~n46116 & ~n46226;
  assign n46228 = ~pi532 & ~n46227;
  assign n46229 = ~pi552 & n46114;
  assign n46230 = ~pi247 & ~n46229;
  assign n46231 = pi552 & n46221;
  assign n46232 = ~pi552 & n46223;
  assign n46233 = pi247 & ~n46232;
  assign n46234 = ~n46231 & n46233;
  assign n46235 = ~n46230 & ~n46234;
  assign n46236 = pi532 & ~n46235;
  assign n46237 = ~n46228 & ~n46236;
  assign n46238 = ~pi238 & n46237;
  assign n46239 = ~pi577 & ~n46238;
  assign n46240 = ~n46116 & ~n46230;
  assign n46241 = pi238 & n46240;
  assign n46242 = pi247 & pi532;
  assign n46243 = ~pi247 & ~pi532;
  assign n46244 = ~n46242 & ~n46243;
  assign n46245 = n46223 & ~n46244;
  assign n46246 = ~pi238 & n46245;
  assign n46247 = pi577 & ~n46246;
  assign n46248 = ~n46241 & n46247;
  assign n46249 = ~pi498 & ~n46248;
  assign n46250 = ~n46239 & n46249;
  assign n46251 = pi238 & n46237;
  assign n46252 = pi577 & ~n46251;
  assign n46253 = ~pi238 & n46240;
  assign n46254 = pi238 & n46245;
  assign n46255 = ~pi577 & ~n46254;
  assign n46256 = ~n46253 & n46255;
  assign n46257 = pi498 & ~n46256;
  assign n46258 = ~n46252 & n46257;
  assign n46259 = ~n46250 & ~n46258;
  assign n46260 = ~pi233 & ~n46259;
  assign n46261 = ~pi544 & ~n45255;
  assign n46262 = pi544 & ~n45669;
  assign n46263 = ~pi240 & ~pi492;
  assign n46264 = pi240 & pi492;
  assign n46265 = ~n46263 & ~n46264;
  assign n46266 = pi241 & pi490;
  assign n46267 = ~pi241 & ~pi490;
  assign n46268 = ~n46266 & ~n46267;
  assign n46269 = pi246 & pi546;
  assign n46270 = ~pi246 & ~pi546;
  assign n46271 = ~n46269 & ~n46270;
  assign n46272 = pi248 & pi548;
  assign n46273 = ~pi248 & ~pi548;
  assign n46274 = ~n46272 & ~n46273;
  assign n46275 = pi249 & pi484;
  assign n46276 = ~pi249 & ~pi484;
  assign n46277 = ~n46275 & ~n46276;
  assign n46278 = ~n46265 & ~n46268;
  assign n46279 = ~n46271 & ~n46274;
  assign n46280 = ~n46277 & n46279;
  assign n46281 = n46278 & n46280;
  assign n46282 = ~n46261 & n46281;
  assign n46283 = ~n46262 & n46282;
  assign n46284 = pi494 & n46283;
  assign n46285 = ~pi239 & ~n46284;
  assign n46286 = ~pi494 & n46283;
  assign n46287 = pi239 & ~n46286;
  assign n46288 = ~n46285 & ~n46287;
  assign n46289 = pi483 & n46288;
  assign n46290 = pi242 & ~n46289;
  assign n46291 = ~pi483 & n46288;
  assign n46292 = ~pi242 & ~n46291;
  assign n46293 = ~n46290 & ~n46292;
  assign n46294 = pi495 & n46293;
  assign n46295 = pi235 & ~n46294;
  assign n46296 = ~pi495 & n46293;
  assign n46297 = ~pi235 & ~n46296;
  assign n46298 = pi244 & pi493;
  assign n46299 = ~pi244 & ~pi493;
  assign n46300 = ~n46298 & ~n46299;
  assign n46301 = ~n46295 & ~n46300;
  assign n46302 = ~n46297 & n46301;
  assign n46303 = pi545 & n46302;
  assign n46304 = pi245 & ~n46303;
  assign n46305 = ~pi545 & n46302;
  assign n46306 = ~pi245 & ~n46305;
  assign n46307 = ~n46304 & ~n46306;
  assign n46308 = pi547 & n46307;
  assign n46309 = pi247 & ~n46308;
  assign n46310 = ~pi547 & n46307;
  assign n46311 = ~pi247 & ~n46310;
  assign n46312 = ~n46309 & ~n46311;
  assign n46313 = ~pi238 & n46312;
  assign n46314 = pi523 & ~n45725;
  assign n46315 = ~pi523 & ~n45279;
  assign n46316 = pi246 & pi526;
  assign n46317 = ~pi246 & ~pi526;
  assign n46318 = ~n46316 & ~n46317;
  assign n46319 = pi248 & pi576;
  assign n46320 = ~pi248 & ~pi576;
  assign n46321 = ~n46319 & ~n46320;
  assign n46322 = pi249 & pi528;
  assign n46323 = ~pi249 & ~pi528;
  assign n46324 = ~n46322 & ~n46323;
  assign n46325 = ~n46318 & ~n46321;
  assign n46326 = ~n46324 & n46325;
  assign n46327 = ~n46314 & n46326;
  assign n46328 = ~n46315 & n46327;
  assign n46329 = pi571 & n46328;
  assign n46330 = pi241 & ~n46329;
  assign n46331 = ~pi571 & n46328;
  assign n46332 = ~pi241 & ~n46331;
  assign n46333 = ~n46330 & ~n46332;
  assign n46334 = ~pi530 & n46333;
  assign n46335 = ~pi240 & ~n46334;
  assign n46336 = pi530 & n46333;
  assign n46337 = pi240 & ~n46336;
  assign n46338 = pi242 & pi573;
  assign n46339 = ~pi242 & ~pi573;
  assign n46340 = ~n46338 & ~n46339;
  assign n46341 = pi235 & pi575;
  assign n46342 = ~pi235 & ~pi575;
  assign n46343 = ~n46341 & ~n46342;
  assign n46344 = ~pi239 & pi524;
  assign n46345 = pi239 & ~pi524;
  assign n46346 = ~n46344 & ~n46345;
  assign n46347 = ~n46340 & ~n46343;
  assign n46348 = ~n46346 & n46347;
  assign n46349 = ~n46335 & n46348;
  assign n46350 = ~n46337 & n46349;
  assign n46351 = ~pi572 & n46350;
  assign n46352 = ~pi244 & ~n46351;
  assign n46353 = pi572 & n46350;
  assign n46354 = pi244 & ~n46353;
  assign n46355 = pi245 & pi525;
  assign n46356 = ~pi245 & ~pi525;
  assign n46357 = ~n46355 & ~n46356;
  assign n46358 = pi247 & pi527;
  assign n46359 = ~pi247 & ~pi527;
  assign n46360 = ~n46358 & ~n46359;
  assign n46361 = ~n46357 & ~n46360;
  assign n46362 = ~n46352 & n46361;
  assign n46363 = ~n46354 & n46362;
  assign n46364 = ~pi238 & n46363;
  assign n46365 = ~pi529 & ~n46364;
  assign n46366 = ~n46313 & n46365;
  assign n46367 = pi238 & n46363;
  assign n46368 = pi529 & ~n46367;
  assign n46369 = ~n46313 & n46368;
  assign n46370 = ~pi491 & ~n46366;
  assign n46371 = ~n46369 & n46370;
  assign n46372 = pi238 & n46312;
  assign n46373 = n46365 & ~n46372;
  assign n46374 = n46368 & ~n46372;
  assign n46375 = pi491 & ~n46373;
  assign n46376 = ~n46374 & n46375;
  assign n46377 = ~n46371 & ~n46376;
  assign n46378 = pi233 & ~n46377;
  assign n46379 = ~pi237 & ~n46378;
  assign n46380 = ~n46260 & n46379;
  assign po750 = ~n46067 & ~n46380;
  assign n46382 = ~pi806 & n44950;
  assign n46383 = ~pi332 & ~pi806;
  assign n46384 = pi990 & n46383;
  assign n46385 = pi600 & n46384;
  assign n46386 = ~pi332 & pi594;
  assign n46387 = ~n46385 & ~n46386;
  assign po751 = ~n46382 & ~n46387;
  assign n46389 = pi605 & ~pi806;
  assign n46390 = n44933 & n46389;
  assign n46391 = ~pi595 & ~n46390;
  assign n46392 = pi595 & n46390;
  assign n46393 = ~pi332 & ~n46391;
  assign po752 = ~n46392 & n46393;
  assign n46395 = ~pi332 & pi596;
  assign n46396 = pi595 & n44932;
  assign n46397 = n46384 & n46396;
  assign n46398 = ~n46395 & ~n46397;
  assign n46399 = pi596 & n46397;
  assign po753 = ~n46398 & ~n46399;
  assign n46401 = ~pi597 & ~n46382;
  assign n46402 = pi597 & n46382;
  assign n46403 = ~pi332 & ~n46401;
  assign po754 = ~n46402 & n46403;
  assign n46405 = ~pi882 & ~po1038;
  assign n46406 = pi947 & n46405;
  assign n46407 = pi598 & ~n46406;
  assign n46408 = pi740 & pi780;
  assign n46409 = n6165 & n46408;
  assign po755 = n46407 | n46409;
  assign n46411 = ~pi332 & pi599;
  assign n46412 = ~n46399 & ~n46411;
  assign n46413 = pi599 & n46399;
  assign po756 = ~n46412 & ~n46413;
  assign n46415 = ~pi332 & pi600;
  assign n46416 = ~n46384 & ~n46415;
  assign po757 = ~n46385 & ~n46416;
  assign n46418 = ~pi806 & ~pi989;
  assign n46419 = ~pi601 & pi806;
  assign n46420 = ~pi332 & ~n46418;
  assign po758 = ~n46419 & n46420;
  assign n46422 = ~pi230 & pi602;
  assign n46423 = ~pi715 & ~pi1160;
  assign n46424 = pi715 & pi1160;
  assign n46425 = pi790 & ~n46423;
  assign n46426 = ~n46424 & n46425;
  assign n46427 = pi230 & n17152;
  assign n46428 = ~n17946 & n46427;
  assign n46429 = ~n19124 & ~n19271;
  assign n46430 = ~n46426 & n46429;
  assign n46431 = n46428 & n46430;
  assign n46432 = n19217 & n46431;
  assign po759 = n46422 | n46432;
  assign n46434 = ~pi980 & pi1038;
  assign n46435 = pi1060 & n46434;
  assign n46436 = pi952 & ~pi1061;
  assign n46437 = n46435 & n46436;
  assign po897 = pi832 & n46437;
  assign n46439 = ~pi603 & ~po897;
  assign n46440 = pi832 & ~pi1100;
  assign n46441 = n46437 & n46440;
  assign n46442 = ~pi966 & ~n46441;
  assign n46443 = ~n46439 & n46442;
  assign n46444 = pi871 & pi966;
  assign n46445 = pi872 & pi966;
  assign n46446 = ~n46444 & ~n46445;
  assign po760 = n46443 | ~n46446;
  assign n46448 = pi823 & n16708;
  assign n46449 = ~pi779 & n46448;
  assign n46450 = ~pi299 & pi983;
  assign n46451 = pi907 & n46450;
  assign n46452 = pi604 & ~n46451;
  assign n46453 = ~n46448 & n46452;
  assign po761 = n46449 | n46453;
  assign n46455 = ~pi605 & ~n46383;
  assign n46456 = ~pi332 & ~n46389;
  assign po762 = ~n46455 & n46456;
  assign n46458 = ~pi606 & ~po897;
  assign n46459 = ~pi1104 & po897;
  assign n46460 = ~n46458 & ~n46459;
  assign n46461 = ~pi966 & ~n46460;
  assign n46462 = ~pi837 & pi966;
  assign po763 = ~n46461 & ~n46462;
  assign n46464 = ~pi607 & ~po897;
  assign n46465 = ~pi1107 & po897;
  assign n46466 = ~pi966 & ~n46464;
  assign po764 = ~n46465 & n46466;
  assign n46468 = ~pi608 & ~po897;
  assign n46469 = ~pi1116 & po897;
  assign n46470 = ~pi966 & ~n46468;
  assign po765 = ~n46469 & n46470;
  assign n46472 = ~pi609 & ~po897;
  assign n46473 = ~pi1118 & po897;
  assign n46474 = ~pi966 & ~n46472;
  assign po766 = ~n46473 & n46474;
  assign n46476 = ~pi610 & ~po897;
  assign n46477 = ~pi1113 & po897;
  assign n46478 = ~pi966 & ~n46476;
  assign po767 = ~n46477 & n46478;
  assign n46480 = ~pi611 & ~po897;
  assign n46481 = ~pi1114 & po897;
  assign n46482 = ~pi966 & ~n46480;
  assign po768 = ~n46481 & n46482;
  assign n46484 = ~pi612 & ~po897;
  assign n46485 = ~pi1111 & po897;
  assign n46486 = ~pi966 & ~n46484;
  assign po769 = ~n46485 & n46486;
  assign n46488 = ~pi613 & ~po897;
  assign n46489 = ~pi1115 & po897;
  assign n46490 = ~pi966 & ~n46488;
  assign po770 = ~n46489 & n46490;
  assign n46492 = ~pi614 & ~po897;
  assign n46493 = ~pi1102 & po897;
  assign n46494 = ~pi966 & ~n46492;
  assign n46495 = ~n46493 & n46494;
  assign po771 = n46444 | n46495;
  assign n46497 = pi907 & n46405;
  assign n46498 = ~pi615 & ~n46497;
  assign n46499 = pi779 & pi797;
  assign n46500 = n6168 & n46499;
  assign po772 = n46498 | n46500;
  assign n46502 = ~pi616 & ~po897;
  assign n46503 = ~pi1101 & po897;
  assign n46504 = ~pi966 & ~n46502;
  assign n46505 = ~n46503 & n46504;
  assign po773 = n46445 | n46505;
  assign n46507 = ~pi617 & ~po897;
  assign n46508 = ~pi1105 & po897;
  assign n46509 = ~n46507 & ~n46508;
  assign n46510 = ~pi966 & ~n46509;
  assign n46511 = ~pi850 & pi966;
  assign po774 = ~n46510 & ~n46511;
  assign n46513 = ~pi618 & ~po897;
  assign n46514 = ~pi1117 & po897;
  assign n46515 = ~pi966 & ~n46513;
  assign po775 = ~n46514 & n46515;
  assign n46517 = ~pi619 & ~po897;
  assign n46518 = ~pi1122 & po897;
  assign n46519 = ~pi966 & ~n46517;
  assign po776 = ~n46518 & n46519;
  assign n46521 = ~pi620 & ~po897;
  assign n46522 = ~pi1112 & po897;
  assign n46523 = ~pi966 & ~n46521;
  assign po777 = ~n46522 & n46523;
  assign n46525 = ~pi621 & ~po897;
  assign n46526 = ~pi1108 & po897;
  assign n46527 = ~pi966 & ~n46525;
  assign po778 = ~n46526 & n46527;
  assign n46529 = ~pi622 & ~po897;
  assign n46530 = ~pi1109 & po897;
  assign n46531 = ~pi966 & ~n46529;
  assign po779 = ~n46530 & n46531;
  assign n46533 = ~pi623 & ~po897;
  assign n46534 = ~pi1106 & po897;
  assign n46535 = ~pi966 & ~n46533;
  assign po780 = ~n46534 & n46535;
  assign n46537 = pi831 & n16854;
  assign n46538 = ~pi780 & n46537;
  assign n46539 = pi947 & n46450;
  assign n46540 = pi624 & ~n46539;
  assign n46541 = ~n46537 & n46540;
  assign po781 = n46538 | n46541;
  assign n46543 = pi832 & ~pi973;
  assign n46544 = ~pi1054 & pi1066;
  assign n46545 = pi1088 & n46544;
  assign n46546 = n46543 & n46545;
  assign po954 = ~pi953 & n46546;
  assign n46548 = ~pi625 & ~po954;
  assign n46549 = ~pi1116 & po954;
  assign n46550 = ~pi962 & ~n46548;
  assign po782 = ~n46549 & n46550;
  assign n46552 = ~pi626 & ~po897;
  assign n46553 = ~pi1121 & po897;
  assign n46554 = ~pi966 & ~n46552;
  assign po783 = ~n46553 & n46554;
  assign n46556 = ~pi627 & ~po954;
  assign n46557 = ~pi1117 & po954;
  assign n46558 = ~pi962 & ~n46556;
  assign po784 = ~n46557 & n46558;
  assign n46560 = ~pi628 & ~po954;
  assign n46561 = ~pi1119 & po954;
  assign n46562 = ~pi962 & ~n46560;
  assign po785 = ~n46561 & n46562;
  assign n46564 = ~pi629 & ~po897;
  assign n46565 = ~pi1119 & po897;
  assign n46566 = ~pi966 & ~n46564;
  assign po786 = ~n46565 & n46566;
  assign n46568 = ~pi630 & ~po897;
  assign n46569 = ~pi1120 & po897;
  assign n46570 = ~pi966 & ~n46568;
  assign po787 = ~n46569 & n46570;
  assign n46572 = ~pi1113 & po954;
  assign n46573 = pi631 & ~po954;
  assign n46574 = ~pi962 & ~n46572;
  assign po788 = ~n46573 & n46574;
  assign n46576 = ~pi1115 & po954;
  assign n46577 = pi632 & ~po954;
  assign n46578 = ~pi962 & ~n46576;
  assign po789 = ~n46577 & n46578;
  assign n46580 = ~pi633 & ~po897;
  assign n46581 = ~pi1110 & po897;
  assign n46582 = ~pi966 & ~n46580;
  assign po790 = ~n46581 & n46582;
  assign n46584 = ~pi634 & ~po954;
  assign n46585 = ~pi1110 & po954;
  assign n46586 = ~pi962 & ~n46584;
  assign po791 = ~n46585 & n46586;
  assign n46588 = ~pi1112 & po954;
  assign n46589 = pi635 & ~po954;
  assign n46590 = ~pi962 & ~n46588;
  assign po792 = ~n46589 & n46590;
  assign n46592 = ~pi636 & ~po897;
  assign n46593 = ~pi1127 & po897;
  assign n46594 = ~pi966 & ~n46592;
  assign po793 = ~n46593 & n46594;
  assign n46596 = ~pi637 & ~po954;
  assign n46597 = ~pi1105 & po954;
  assign n46598 = ~pi962 & ~n46596;
  assign po794 = ~n46597 & n46598;
  assign n46600 = ~pi638 & ~po954;
  assign n46601 = ~pi1107 & po954;
  assign n46602 = ~pi962 & ~n46600;
  assign po795 = ~n46601 & n46602;
  assign n46604 = ~pi639 & ~po954;
  assign n46605 = ~pi1109 & po954;
  assign n46606 = ~pi962 & ~n46604;
  assign po796 = ~n46605 & n46606;
  assign n46608 = ~pi640 & ~po897;
  assign n46609 = ~pi1128 & po897;
  assign n46610 = ~pi966 & ~n46608;
  assign po797 = ~n46609 & n46610;
  assign n46612 = ~pi641 & ~po954;
  assign n46613 = ~pi1121 & po954;
  assign n46614 = ~pi962 & ~n46612;
  assign po798 = ~n46613 & n46614;
  assign n46616 = ~pi642 & ~po897;
  assign n46617 = ~pi1103 & po897;
  assign n46618 = ~pi966 & ~n46616;
  assign po799 = ~n46617 & n46618;
  assign n46620 = ~pi643 & ~po954;
  assign n46621 = ~pi1104 & po954;
  assign n46622 = ~pi962 & ~n46620;
  assign po800 = ~n46621 & n46622;
  assign n46624 = ~pi644 & ~po897;
  assign n46625 = ~pi1123 & po897;
  assign n46626 = ~pi966 & ~n46624;
  assign po801 = ~n46625 & n46626;
  assign n46628 = ~pi645 & ~po897;
  assign n46629 = ~pi1125 & po897;
  assign n46630 = ~pi966 & ~n46628;
  assign po802 = ~n46629 & n46630;
  assign n46632 = ~pi1114 & po954;
  assign n46633 = pi646 & ~po954;
  assign n46634 = ~pi962 & ~n46632;
  assign po803 = ~n46633 & n46634;
  assign n46636 = ~pi647 & ~po954;
  assign n46637 = ~pi1120 & po954;
  assign n46638 = ~pi962 & ~n46636;
  assign po804 = ~n46637 & n46638;
  assign n46640 = ~pi648 & ~po954;
  assign n46641 = ~pi1122 & po954;
  assign n46642 = ~pi962 & ~n46640;
  assign po805 = ~n46641 & n46642;
  assign n46644 = ~pi1126 & po954;
  assign n46645 = pi649 & ~po954;
  assign n46646 = ~pi962 & ~n46644;
  assign po806 = ~n46645 & n46646;
  assign n46648 = ~pi1127 & po954;
  assign n46649 = pi650 & ~po954;
  assign n46650 = ~pi962 & ~n46648;
  assign po807 = ~n46649 & n46650;
  assign n46652 = ~pi651 & ~po897;
  assign n46653 = ~pi1130 & po897;
  assign n46654 = ~pi966 & ~n46652;
  assign po808 = ~n46653 & n46654;
  assign n46656 = ~pi652 & ~po897;
  assign n46657 = ~pi1131 & po897;
  assign n46658 = ~pi966 & ~n46656;
  assign po809 = ~n46657 & n46658;
  assign n46660 = ~pi653 & ~po897;
  assign n46661 = ~pi1129 & po897;
  assign n46662 = ~pi966 & ~n46660;
  assign po810 = ~n46661 & n46662;
  assign n46664 = ~pi1130 & po954;
  assign n46665 = pi654 & ~po954;
  assign n46666 = ~pi962 & ~n46664;
  assign po811 = ~n46665 & n46666;
  assign n46668 = ~pi1124 & po954;
  assign n46669 = pi655 & ~po954;
  assign n46670 = ~pi962 & ~n46668;
  assign po812 = ~n46669 & n46670;
  assign n46672 = ~pi656 & ~po897;
  assign n46673 = ~pi1126 & po897;
  assign n46674 = ~pi966 & ~n46672;
  assign po813 = ~n46673 & n46674;
  assign n46676 = ~pi1131 & po954;
  assign n46677 = pi657 & ~po954;
  assign n46678 = ~pi962 & ~n46676;
  assign po814 = ~n46677 & n46678;
  assign n46680 = ~pi658 & ~po897;
  assign n46681 = ~pi1124 & po897;
  assign n46682 = ~pi966 & ~n46680;
  assign po815 = ~n46681 & n46682;
  assign n46684 = pi266 & pi992;
  assign n46685 = ~pi280 & n46684;
  assign n46686 = ~pi269 & n46685;
  assign n46687 = ~pi281 & n46686;
  assign n46688 = ~pi270 & ~pi277;
  assign n46689 = ~pi282 & n46688;
  assign n46690 = n46687 & n46689;
  assign n46691 = ~pi264 & n46690;
  assign n46692 = ~pi265 & n46691;
  assign po959 = ~pi274 & n46692;
  assign n46694 = pi274 & ~n46692;
  assign po816 = ~po959 & ~n46694;
  assign n46696 = ~pi660 & ~po954;
  assign n46697 = ~pi1118 & po954;
  assign n46698 = ~pi962 & ~n46696;
  assign po817 = ~n46697 & n46698;
  assign n46700 = ~pi661 & ~po954;
  assign n46701 = ~pi1101 & po954;
  assign n46702 = ~pi962 & ~n46700;
  assign po818 = ~n46701 & n46702;
  assign n46704 = ~pi662 & ~po954;
  assign n46705 = ~pi1102 & po954;
  assign n46706 = ~pi962 & ~n46704;
  assign po819 = ~n46705 & n46706;
  assign n46708 = pi199 & ~pi1065;
  assign n46709 = ~pi223 & ~pi224;
  assign n46710 = ~pi199 & ~pi257;
  assign n46711 = ~n46708 & ~n46709;
  assign n46712 = ~n46710 & n46711;
  assign n46713 = ~pi591 & pi592;
  assign n46714 = pi365 & n46713;
  assign n46715 = pi334 & pi591;
  assign n46716 = ~pi592 & n46715;
  assign n46717 = ~n46714 & ~n46716;
  assign n46718 = ~pi590 & ~n46717;
  assign n46719 = ~pi591 & ~pi592;
  assign n46720 = pi590 & n46719;
  assign n46721 = pi323 & n46720;
  assign n46722 = ~pi588 & ~n46721;
  assign n46723 = ~n46718 & n46722;
  assign n46724 = ~pi592 & n8585;
  assign n46725 = pi464 & n46724;
  assign n46726 = pi588 & ~n46725;
  assign n46727 = n46709 & ~n46726;
  assign n46728 = ~n46723 & n46727;
  assign n46729 = ~n46712 & ~n46728;
  assign n46730 = n8856 & ~n46729;
  assign n46731 = ~pi1137 & ~pi1138;
  assign n46732 = ~pi1134 & n46731;
  assign n46733 = ~pi784 & ~pi1136;
  assign n46734 = ~pi634 & pi1136;
  assign n46735 = pi1135 & ~n46733;
  assign n46736 = ~n46734 & n46735;
  assign n46737 = ~pi815 & ~pi1136;
  assign n46738 = ~pi633 & pi1136;
  assign n46739 = ~pi1135 & ~n46737;
  assign n46740 = ~n46738 & n46739;
  assign n46741 = ~n46736 & ~n46740;
  assign n46742 = n46732 & ~n46741;
  assign n46743 = pi1135 & n46731;
  assign n46744 = pi1136 & ~n46743;
  assign n46745 = ~pi766 & n46744;
  assign n46746 = pi1135 & ~pi1136;
  assign n46747 = pi1134 & n46731;
  assign n46748 = ~n46746 & n46747;
  assign n46749 = ~pi855 & ~pi1136;
  assign n46750 = ~pi700 & pi1135;
  assign n46751 = ~n46749 & ~n46750;
  assign n46752 = n46748 & n46751;
  assign n46753 = ~n46745 & n46752;
  assign n46754 = ~n46742 & ~n46753;
  assign n46755 = ~n8856 & ~n46754;
  assign po820 = n46730 | n46755;
  assign n46757 = ~pi590 & pi591;
  assign n46758 = pi404 & n46757;
  assign n46759 = ~pi590 & pi592;
  assign n46760 = ~pi588 & ~n46759;
  assign n46761 = ~n46758 & n46760;
  assign n46762 = pi380 & ~pi591;
  assign n46763 = pi592 & ~n46762;
  assign n46764 = ~n46761 & ~n46763;
  assign n46765 = pi355 & n46720;
  assign n46766 = ~n46764 & ~n46765;
  assign n46767 = pi429 & n46724;
  assign n46768 = pi588 & ~n46767;
  assign n46769 = n46709 & ~n46768;
  assign n46770 = ~n46766 & n46769;
  assign n46771 = ~pi199 & ~pi292;
  assign n46772 = pi199 & ~pi1084;
  assign n46773 = ~n46709 & ~n46771;
  assign n46774 = ~n46772 & n46773;
  assign n46775 = ~n46770 & ~n46774;
  assign n46776 = n8856 & ~n46775;
  assign n46777 = pi614 & ~pi1135;
  assign n46778 = pi662 & pi1135;
  assign n46779 = pi1136 & ~n46777;
  assign n46780 = ~n46778 & n46779;
  assign n46781 = pi811 & ~pi1135;
  assign n46782 = pi785 & pi1135;
  assign n46783 = ~pi1136 & ~n46781;
  assign n46784 = ~n46782 & n46783;
  assign n46785 = ~n46780 & ~n46784;
  assign n46786 = ~pi1134 & ~n46785;
  assign n46787 = ~pi772 & ~pi1135;
  assign n46788 = ~pi727 & pi1135;
  assign n46789 = pi1136 & ~n46787;
  assign n46790 = ~n46788 & n46789;
  assign n46791 = ~pi1135 & ~pi1136;
  assign n46792 = pi872 & n46791;
  assign n46793 = pi1134 & ~n46792;
  assign n46794 = ~n46790 & n46793;
  assign n46795 = ~n8856 & n46731;
  assign n46796 = ~n46794 & n46795;
  assign n46797 = ~n46786 & n46796;
  assign po821 = n46776 | n46797;
  assign n46799 = ~pi665 & ~po954;
  assign n46800 = ~pi1108 & po954;
  assign n46801 = ~pi962 & ~n46799;
  assign po822 = ~n46800 & n46801;
  assign n46803 = ~pi607 & ~pi1135;
  assign n46804 = ~pi638 & pi1135;
  assign n46805 = pi1136 & ~n46803;
  assign n46806 = ~n46804 & n46805;
  assign n46807 = ~pi790 & pi1135;
  assign n46808 = pi799 & ~pi1135;
  assign n46809 = ~pi1136 & ~n46807;
  assign n46810 = ~n46808 & n46809;
  assign n46811 = ~n46806 & ~n46810;
  assign n46812 = n46732 & ~n46811;
  assign n46813 = ~pi764 & n46744;
  assign n46814 = ~pi691 & pi1135;
  assign n46815 = ~pi873 & ~pi1136;
  assign n46816 = ~n46814 & ~n46815;
  assign n46817 = n46748 & n46816;
  assign n46818 = ~n46813 & n46817;
  assign n46819 = ~n46812 & ~n46818;
  assign n46820 = ~n8856 & ~n46819;
  assign n46821 = ~pi199 & ~pi297;
  assign n46822 = pi199 & ~pi1044;
  assign n46823 = ~n46709 & ~n46821;
  assign n46824 = ~n46822 & n46823;
  assign n46825 = pi456 & n46757;
  assign n46826 = n46760 & ~n46825;
  assign n46827 = pi337 & ~pi591;
  assign n46828 = pi592 & ~n46827;
  assign n46829 = ~n46826 & ~n46828;
  assign n46830 = pi441 & n46720;
  assign n46831 = ~n46829 & ~n46830;
  assign n46832 = pi443 & n46724;
  assign n46833 = pi588 & ~n46832;
  assign n46834 = n46709 & ~n46833;
  assign n46835 = ~n46831 & n46834;
  assign n46836 = ~n46824 & ~n46835;
  assign n46837 = n8856 & ~n46836;
  assign po823 = n46820 | n46837;
  assign n46839 = pi319 & n46757;
  assign n46840 = n46760 & ~n46839;
  assign n46841 = pi338 & ~pi591;
  assign n46842 = pi592 & ~n46841;
  assign n46843 = ~n46840 & ~n46842;
  assign n46844 = pi458 & n46720;
  assign n46845 = ~n46843 & ~n46844;
  assign n46846 = pi444 & n46724;
  assign n46847 = pi588 & ~n46846;
  assign n46848 = n46709 & ~n46847;
  assign n46849 = ~n46845 & n46848;
  assign n46850 = ~pi199 & ~pi294;
  assign n46851 = pi199 & ~pi1072;
  assign n46852 = ~n46709 & ~n46850;
  assign n46853 = ~n46851 & n46852;
  assign n46854 = ~n46849 & ~n46853;
  assign n46855 = n8856 & ~n46854;
  assign n46856 = pi792 & ~pi1136;
  assign n46857 = pi681 & pi1136;
  assign n46858 = pi1135 & ~n46856;
  assign n46859 = ~n46857 & n46858;
  assign n46860 = ~pi809 & ~pi1136;
  assign n46861 = pi642 & pi1136;
  assign n46862 = ~pi1135 & ~n46860;
  assign n46863 = ~n46861 & n46862;
  assign n46864 = ~n46859 & ~n46863;
  assign n46865 = ~pi1134 & ~n46864;
  assign n46866 = ~pi763 & ~pi1135;
  assign n46867 = ~pi699 & pi1135;
  assign n46868 = pi1136 & ~n46866;
  assign n46869 = ~n46867 & n46868;
  assign n46870 = pi871 & n46791;
  assign n46871 = pi1134 & ~n46870;
  assign n46872 = ~n46869 & n46871;
  assign n46873 = n46795 & ~n46872;
  assign n46874 = ~n46865 & n46873;
  assign po824 = n46855 | n46874;
  assign n46876 = ~pi603 & ~pi1135;
  assign n46877 = ~pi680 & pi1135;
  assign n46878 = pi1136 & ~n46876;
  assign n46879 = ~n46877 & n46878;
  assign n46880 = ~pi981 & ~pi1135;
  assign n46881 = ~pi778 & pi1135;
  assign n46882 = ~pi1136 & ~n46880;
  assign n46883 = ~n46881 & n46882;
  assign n46884 = ~n46879 & ~n46883;
  assign n46885 = n46732 & ~n46884;
  assign n46886 = ~pi759 & n46744;
  assign n46887 = ~pi696 & pi1135;
  assign n46888 = ~pi837 & ~pi1136;
  assign n46889 = ~n46887 & ~n46888;
  assign n46890 = n46748 & n46889;
  assign n46891 = ~n46886 & n46890;
  assign n46892 = ~n46885 & ~n46891;
  assign n46893 = ~n8856 & ~n46892;
  assign n46894 = ~pi199 & ~pi291;
  assign n46895 = pi199 & ~pi1049;
  assign n46896 = ~n46709 & ~n46894;
  assign n46897 = ~n46895 & n46896;
  assign n46898 = pi390 & n46757;
  assign n46899 = n46760 & ~n46898;
  assign n46900 = pi363 & ~pi591;
  assign n46901 = pi592 & ~n46900;
  assign n46902 = ~n46899 & ~n46901;
  assign n46903 = pi342 & n46720;
  assign n46904 = ~n46902 & ~n46903;
  assign n46905 = pi414 & n46724;
  assign n46906 = pi588 & ~n46905;
  assign n46907 = n46709 & ~n46906;
  assign n46908 = ~n46904 & n46907;
  assign n46909 = ~n46897 & ~n46908;
  assign n46910 = n8856 & ~n46909;
  assign po825 = n46893 | n46910;
  assign n46912 = ~pi1125 & po954;
  assign n46913 = pi669 & ~po954;
  assign n46914 = ~pi962 & ~n46912;
  assign po826 = ~n46913 & n46914;
  assign n46916 = ~pi199 & ~pi258;
  assign n46917 = pi199 & ~pi1062;
  assign n46918 = ~n46709 & ~n46916;
  assign n46919 = ~n46917 & n46918;
  assign n46920 = pi364 & n46713;
  assign n46921 = pi391 & pi591;
  assign n46922 = ~pi592 & n46921;
  assign n46923 = ~n46920 & ~n46922;
  assign n46924 = ~pi590 & ~n46923;
  assign n46925 = pi343 & n46720;
  assign n46926 = ~pi588 & ~n46925;
  assign n46927 = ~n46924 & n46926;
  assign n46928 = pi415 & n46724;
  assign n46929 = pi588 & ~n46928;
  assign n46930 = n46709 & ~n46929;
  assign n46931 = ~n46927 & n46930;
  assign n46932 = ~n46919 & ~n46931;
  assign n46933 = n8856 & ~n46932;
  assign n46934 = pi745 & n46744;
  assign n46935 = pi723 & pi1135;
  assign n46936 = ~pi852 & ~pi1136;
  assign n46937 = ~n46935 & ~n46936;
  assign n46938 = n46748 & n46937;
  assign n46939 = ~n46934 & n46938;
  assign n46940 = pi1136 & n46731;
  assign n46941 = pi695 & pi1135;
  assign n46942 = ~pi612 & ~pi1135;
  assign n46943 = ~pi1134 & ~n46941;
  assign n46944 = ~n46942 & n46943;
  assign n46945 = n46940 & n46944;
  assign n46946 = ~n46939 & ~n46945;
  assign n46947 = ~n8856 & ~n46946;
  assign po827 = n46933 | n46947;
  assign n46949 = ~pi199 & ~pi261;
  assign n46950 = pi199 & ~pi1040;
  assign n46951 = ~n46709 & ~n46949;
  assign n46952 = ~n46950 & n46951;
  assign n46953 = pi447 & n46713;
  assign n46954 = pi333 & pi591;
  assign n46955 = ~pi592 & n46954;
  assign n46956 = ~n46953 & ~n46955;
  assign n46957 = ~pi590 & ~n46956;
  assign n46958 = pi327 & n46720;
  assign n46959 = ~pi588 & ~n46958;
  assign n46960 = ~n46957 & n46959;
  assign n46961 = pi453 & n46724;
  assign n46962 = pi588 & ~n46961;
  assign n46963 = n46709 & ~n46962;
  assign n46964 = ~n46960 & n46963;
  assign n46965 = ~n46952 & ~n46964;
  assign n46966 = n8856 & ~n46965;
  assign n46967 = pi741 & n46744;
  assign n46968 = pi724 & pi1135;
  assign n46969 = ~pi865 & ~pi1136;
  assign n46970 = ~n46968 & ~n46969;
  assign n46971 = n46748 & n46970;
  assign n46972 = ~n46967 & n46971;
  assign n46973 = pi646 & pi1135;
  assign n46974 = ~pi611 & ~pi1135;
  assign n46975 = ~pi1134 & ~n46973;
  assign n46976 = ~n46974 & n46975;
  assign n46977 = n46940 & n46976;
  assign n46978 = ~n46972 & ~n46977;
  assign n46979 = ~n8856 & ~n46978;
  assign po828 = n46966 | n46979;
  assign n46981 = ~pi616 & ~pi1135;
  assign n46982 = ~pi661 & pi1135;
  assign n46983 = pi1136 & ~n46981;
  assign n46984 = ~n46982 & n46983;
  assign n46985 = ~pi808 & ~pi1135;
  assign n46986 = ~pi781 & pi1135;
  assign n46987 = ~pi1136 & ~n46985;
  assign n46988 = ~n46986 & n46987;
  assign n46989 = ~n46984 & ~n46988;
  assign n46990 = n46732 & ~n46989;
  assign n46991 = ~pi758 & n46744;
  assign n46992 = ~pi736 & pi1135;
  assign n46993 = ~pi850 & ~pi1136;
  assign n46994 = ~n46992 & ~n46993;
  assign n46995 = n46748 & n46994;
  assign n46996 = ~n46991 & n46995;
  assign n46997 = ~n46990 & ~n46996;
  assign n46998 = ~n8856 & ~n46997;
  assign n46999 = ~pi199 & ~pi290;
  assign n47000 = pi199 & ~pi1048;
  assign n47001 = ~n46709 & ~n46999;
  assign n47002 = ~n47000 & n47001;
  assign n47003 = pi397 & n46757;
  assign n47004 = n46760 & ~n47003;
  assign n47005 = pi372 & ~pi591;
  assign n47006 = pi592 & ~n47005;
  assign n47007 = ~n47004 & ~n47006;
  assign n47008 = pi320 & n46720;
  assign n47009 = ~n47007 & ~n47008;
  assign n47010 = pi422 & n46724;
  assign n47011 = pi588 & ~n47010;
  assign n47012 = n46709 & ~n47011;
  assign n47013 = ~n47009 & n47012;
  assign n47014 = ~n47002 & ~n47013;
  assign n47015 = n8856 & ~n47014;
  assign po829 = n46998 | n47015;
  assign n47017 = ~pi617 & ~pi1135;
  assign n47018 = ~pi637 & pi1135;
  assign n47019 = pi1136 & ~n47017;
  assign n47020 = ~n47018 & n47019;
  assign n47021 = ~pi788 & pi1135;
  assign n47022 = pi814 & ~pi1135;
  assign n47023 = ~pi1136 & ~n47021;
  assign n47024 = ~n47022 & n47023;
  assign n47025 = ~n47020 & ~n47024;
  assign n47026 = n46732 & ~n47025;
  assign n47027 = ~pi749 & n46744;
  assign n47028 = ~pi706 & pi1135;
  assign n47029 = ~pi866 & ~pi1136;
  assign n47030 = ~n47028 & ~n47029;
  assign n47031 = n46748 & n47030;
  assign n47032 = ~n47027 & n47031;
  assign n47033 = ~n47026 & ~n47032;
  assign n47034 = ~n8856 & ~n47033;
  assign n47035 = ~pi199 & ~pi295;
  assign n47036 = pi199 & ~pi1053;
  assign n47037 = ~n46709 & ~n47035;
  assign n47038 = ~n47036 & n47037;
  assign n47039 = pi411 & n46757;
  assign n47040 = n46760 & ~n47039;
  assign n47041 = pi387 & ~pi591;
  assign n47042 = pi592 & ~n47041;
  assign n47043 = ~n47040 & ~n47042;
  assign n47044 = pi452 & n46720;
  assign n47045 = ~n47043 & ~n47044;
  assign n47046 = pi435 & n46724;
  assign n47047 = pi588 & ~n47046;
  assign n47048 = n46709 & ~n47047;
  assign n47049 = ~n47045 & n47048;
  assign n47050 = ~n47038 & ~n47049;
  assign n47051 = n8856 & ~n47050;
  assign po830 = n47034 | n47051;
  assign n47053 = ~pi199 & ~pi256;
  assign n47054 = pi199 & ~pi1070;
  assign n47055 = ~n46709 & ~n47053;
  assign n47056 = ~n47054 & n47055;
  assign n47057 = pi336 & n46713;
  assign n47058 = pi463 & pi591;
  assign n47059 = ~pi592 & n47058;
  assign n47060 = ~n47057 & ~n47059;
  assign n47061 = ~pi590 & ~n47060;
  assign n47062 = pi362 & n46720;
  assign n47063 = ~pi588 & ~n47062;
  assign n47064 = ~n47061 & n47063;
  assign n47065 = pi437 & n46724;
  assign n47066 = pi588 & ~n47065;
  assign n47067 = n46709 & ~n47066;
  assign n47068 = ~n47064 & n47067;
  assign n47069 = ~n47056 & ~n47068;
  assign n47070 = n8856 & ~n47069;
  assign n47071 = pi622 & ~pi1135;
  assign n47072 = pi639 & pi1135;
  assign n47073 = pi1136 & ~n47071;
  assign n47074 = ~n47072 & n47073;
  assign n47075 = pi804 & ~pi1135;
  assign n47076 = pi783 & pi1135;
  assign n47077 = ~pi1136 & ~n47075;
  assign n47078 = ~n47076 & n47077;
  assign n47079 = ~n47074 & ~n47078;
  assign n47080 = ~pi1134 & ~n47079;
  assign n47081 = ~pi743 & ~pi1135;
  assign n47082 = ~pi735 & pi1135;
  assign n47083 = pi1136 & ~n47081;
  assign n47084 = ~n47082 & n47083;
  assign n47085 = pi859 & n46791;
  assign n47086 = pi1134 & ~n47085;
  assign n47087 = ~n47084 & n47086;
  assign n47088 = n46795 & ~n47087;
  assign n47089 = ~n47080 & n47088;
  assign po831 = n47070 | n47089;
  assign n47091 = pi876 & n46791;
  assign n47092 = ~pi748 & ~pi1135;
  assign n47093 = ~pi730 & pi1135;
  assign n47094 = pi1136 & ~n47092;
  assign n47095 = ~n47093 & n47094;
  assign n47096 = ~n47091 & ~n47095;
  assign n47097 = n46747 & ~n47096;
  assign n47098 = ~pi623 & n46744;
  assign n47099 = pi789 & n46746;
  assign n47100 = ~pi710 & pi1135;
  assign n47101 = pi1136 & ~n47100;
  assign n47102 = ~pi803 & ~pi1135;
  assign n47103 = ~n47099 & ~n47102;
  assign n47104 = ~n47101 & n47103;
  assign n47105 = n46732 & ~n47098;
  assign n47106 = ~n47104 & n47105;
  assign n47107 = ~n47097 & ~n47106;
  assign n47108 = ~n8856 & ~n47107;
  assign n47109 = ~pi199 & ~pi296;
  assign n47110 = pi199 & ~pi1037;
  assign n47111 = ~n46709 & ~n47109;
  assign n47112 = ~n47110 & n47111;
  assign n47113 = pi412 & n46757;
  assign n47114 = n46760 & ~n47113;
  assign n47115 = pi388 & ~pi591;
  assign n47116 = pi592 & ~n47115;
  assign n47117 = ~n47114 & ~n47116;
  assign n47118 = pi455 & n46720;
  assign n47119 = ~n47117 & ~n47118;
  assign n47120 = pi436 & n46724;
  assign n47121 = pi588 & ~n47120;
  assign n47122 = n46709 & ~n47121;
  assign n47123 = ~n47119 & n47122;
  assign n47124 = ~n47112 & ~n47123;
  assign n47125 = n8856 & ~n47124;
  assign po832 = n47108 | n47125;
  assign n47127 = ~pi606 & ~pi1135;
  assign n47128 = ~pi643 & pi1135;
  assign n47129 = pi1136 & ~n47127;
  assign n47130 = ~n47128 & n47129;
  assign n47131 = ~pi787 & pi1135;
  assign n47132 = pi812 & ~pi1135;
  assign n47133 = ~pi1136 & ~n47131;
  assign n47134 = ~n47132 & n47133;
  assign n47135 = ~n47130 & ~n47134;
  assign n47136 = n46732 & ~n47135;
  assign n47137 = ~pi746 & n46744;
  assign n47138 = ~pi729 & pi1135;
  assign n47139 = ~pi881 & ~pi1136;
  assign n47140 = ~n47138 & ~n47139;
  assign n47141 = n46748 & n47140;
  assign n47142 = ~n47137 & n47141;
  assign n47143 = ~n47136 & ~n47142;
  assign n47144 = ~n8856 & ~n47143;
  assign n47145 = ~pi199 & ~pi293;
  assign n47146 = pi199 & ~pi1059;
  assign n47147 = ~n46709 & ~n47145;
  assign n47148 = ~n47146 & n47147;
  assign n47149 = pi410 & n46757;
  assign n47150 = n46760 & ~n47149;
  assign n47151 = pi386 & ~pi591;
  assign n47152 = pi592 & ~n47151;
  assign n47153 = ~n47150 & ~n47152;
  assign n47154 = pi361 & n46720;
  assign n47155 = ~n47153 & ~n47154;
  assign n47156 = pi434 & n46724;
  assign n47157 = pi588 & ~n47156;
  assign n47158 = n46709 & ~n47157;
  assign n47159 = ~n47155 & n47158;
  assign n47160 = ~n47148 & ~n47159;
  assign n47161 = n8856 & ~n47160;
  assign po833 = n47144 | n47161;
  assign n47163 = ~pi199 & ~pi259;
  assign n47164 = pi199 & ~pi1069;
  assign n47165 = ~n46709 & ~n47163;
  assign n47166 = ~n47164 & n47165;
  assign n47167 = pi366 & n46713;
  assign n47168 = pi335 & pi591;
  assign n47169 = ~pi592 & n47168;
  assign n47170 = ~n47167 & ~n47169;
  assign n47171 = ~pi590 & ~n47170;
  assign n47172 = pi344 & n46720;
  assign n47173 = ~pi588 & ~n47172;
  assign n47174 = ~n47171 & n47173;
  assign n47175 = pi416 & n46724;
  assign n47176 = pi588 & ~n47175;
  assign n47177 = n46709 & ~n47176;
  assign n47178 = ~n47174 & n47177;
  assign n47179 = ~n47166 & ~n47178;
  assign n47180 = n8856 & ~n47179;
  assign n47181 = pi742 & n46744;
  assign n47182 = pi704 & pi1135;
  assign n47183 = ~pi870 & ~pi1136;
  assign n47184 = ~n47182 & ~n47183;
  assign n47185 = n46748 & n47184;
  assign n47186 = ~n47181 & n47185;
  assign n47187 = pi635 & pi1135;
  assign n47188 = ~pi620 & ~pi1135;
  assign n47189 = ~pi1134 & ~n47187;
  assign n47190 = ~n47188 & n47189;
  assign n47191 = n46940 & n47190;
  assign n47192 = ~n47186 & ~n47191;
  assign n47193 = ~n8856 & ~n47192;
  assign po834 = n47180 | n47193;
  assign n47195 = ~pi199 & ~pi260;
  assign n47196 = pi199 & ~pi1067;
  assign n47197 = ~n46709 & ~n47195;
  assign n47198 = ~n47196 & n47197;
  assign n47199 = pi368 & n46713;
  assign n47200 = pi393 & pi591;
  assign n47201 = ~pi592 & n47200;
  assign n47202 = ~n47199 & ~n47201;
  assign n47203 = ~pi590 & ~n47202;
  assign n47204 = pi346 & n46720;
  assign n47205 = ~pi588 & ~n47204;
  assign n47206 = ~n47203 & n47205;
  assign n47207 = pi418 & n46724;
  assign n47208 = pi588 & ~n47207;
  assign n47209 = n46709 & ~n47208;
  assign n47210 = ~n47206 & n47209;
  assign n47211 = ~n47198 & ~n47210;
  assign n47212 = n8856 & ~n47211;
  assign n47213 = pi760 & n46744;
  assign n47214 = pi688 & pi1135;
  assign n47215 = ~pi856 & ~pi1136;
  assign n47216 = ~n47214 & ~n47215;
  assign n47217 = n46748 & n47216;
  assign n47218 = ~n47213 & n47217;
  assign n47219 = pi632 & pi1135;
  assign n47220 = ~pi613 & ~pi1135;
  assign n47221 = ~pi1134 & ~n47219;
  assign n47222 = ~n47220 & n47221;
  assign n47223 = n46940 & n47222;
  assign n47224 = ~n47218 & ~n47223;
  assign n47225 = ~n8856 & ~n47224;
  assign po835 = n47212 | n47225;
  assign n47227 = ~pi199 & ~pi255;
  assign n47228 = pi199 & ~pi1036;
  assign n47229 = ~n46709 & ~n47227;
  assign n47230 = ~n47228 & n47229;
  assign n47231 = pi389 & n46713;
  assign n47232 = pi413 & pi591;
  assign n47233 = ~pi592 & n47232;
  assign n47234 = ~n47231 & ~n47233;
  assign n47235 = ~pi590 & ~n47234;
  assign n47236 = pi450 & n46720;
  assign n47237 = ~pi588 & ~n47236;
  assign n47238 = ~n47235 & n47237;
  assign n47239 = pi438 & n46724;
  assign n47240 = pi588 & ~n47239;
  assign n47241 = n46709 & ~n47240;
  assign n47242 = ~n47238 & n47241;
  assign n47243 = ~n47230 & ~n47242;
  assign n47244 = n8856 & ~n47243;
  assign n47245 = ~pi791 & ~pi1136;
  assign n47246 = ~pi665 & pi1136;
  assign n47247 = pi1135 & ~n47245;
  assign n47248 = ~n47246 & n47247;
  assign n47249 = ~pi810 & ~pi1136;
  assign n47250 = ~pi621 & pi1136;
  assign n47251 = ~pi1135 & ~n47249;
  assign n47252 = ~n47250 & n47251;
  assign n47253 = ~n47248 & ~n47252;
  assign n47254 = n46732 & ~n47253;
  assign n47255 = ~pi739 & n46744;
  assign n47256 = ~pi874 & ~pi1136;
  assign n47257 = ~pi690 & pi1135;
  assign n47258 = ~n47256 & ~n47257;
  assign n47259 = n46748 & n47258;
  assign n47260 = ~n47255 & n47259;
  assign n47261 = ~n47254 & ~n47260;
  assign n47262 = ~n8856 & ~n47261;
  assign po836 = n47244 | n47262;
  assign n47264 = ~pi680 & ~po954;
  assign n47265 = ~pi1100 & po954;
  assign n47266 = ~pi962 & ~n47264;
  assign po837 = ~n47265 & n47266;
  assign n47268 = ~pi681 & ~po954;
  assign n47269 = ~pi1103 & po954;
  assign n47270 = ~pi962 & ~n47268;
  assign po838 = ~n47269 & n47270;
  assign n47272 = ~pi199 & ~pi251;
  assign n47273 = pi199 & ~pi1039;
  assign n47274 = ~n46709 & ~n47272;
  assign n47275 = ~n47273 & n47274;
  assign n47276 = pi367 & n46713;
  assign n47277 = pi392 & pi591;
  assign n47278 = ~pi592 & n47277;
  assign n47279 = ~n47276 & ~n47278;
  assign n47280 = ~pi590 & ~n47279;
  assign n47281 = pi345 & n46720;
  assign n47282 = ~pi588 & ~n47281;
  assign n47283 = ~n47280 & n47282;
  assign n47284 = pi417 & n46724;
  assign n47285 = pi588 & ~n47284;
  assign n47286 = n46709 & ~n47285;
  assign n47287 = ~n47283 & n47286;
  assign n47288 = ~n47275 & ~n47287;
  assign n47289 = n8856 & ~n47288;
  assign n47290 = pi757 & n46744;
  assign n47291 = pi686 & pi1135;
  assign n47292 = ~pi848 & ~pi1136;
  assign n47293 = ~n47291 & ~n47292;
  assign n47294 = n46748 & n47293;
  assign n47295 = ~n47290 & n47294;
  assign n47296 = pi631 & pi1135;
  assign n47297 = ~pi610 & ~pi1135;
  assign n47298 = ~pi1134 & ~n47296;
  assign n47299 = ~n47297 & n47298;
  assign n47300 = n46940 & n47299;
  assign n47301 = ~n47295 & ~n47300;
  assign n47302 = ~n8856 & ~n47301;
  assign po839 = n47289 | n47302;
  assign po980 = pi953 & n46546;
  assign n47305 = ~pi1130 & po980;
  assign n47306 = pi684 & ~po980;
  assign n47307 = ~pi962 & ~n47305;
  assign po841 = ~n47306 & n47307;
  assign n47309 = pi590 & ~pi592;
  assign n47310 = pi357 & n47309;
  assign n47311 = pi382 & n46759;
  assign n47312 = ~n47310 & ~n47311;
  assign n47313 = ~pi591 & ~n47312;
  assign n47314 = pi406 & ~pi592;
  assign n47315 = n46757 & n47314;
  assign n47316 = ~n47313 & ~n47315;
  assign n47317 = ~pi588 & ~n47316;
  assign n47318 = pi588 & ~pi590;
  assign n47319 = pi430 & n46719;
  assign n47320 = n47318 & n47319;
  assign n47321 = ~n47317 & ~n47320;
  assign n47322 = n46709 & ~n47321;
  assign n47323 = pi199 & ~pi1076;
  assign n47324 = ~n46709 & ~n47323;
  assign n47325 = ~n42714 & n47324;
  assign n47326 = ~n47322 & ~n47325;
  assign n47327 = n8856 & ~n47326;
  assign n47328 = pi860 & n46791;
  assign n47329 = pi744 & ~pi1135;
  assign n47330 = pi728 & pi1135;
  assign n47331 = pi1136 & ~n47329;
  assign n47332 = ~n47330 & n47331;
  assign n47333 = ~n47328 & ~n47332;
  assign n47334 = n46747 & ~n47333;
  assign n47335 = pi1136 & ~n46731;
  assign n47336 = ~pi1134 & ~n47335;
  assign n47337 = ~pi652 & ~pi1135;
  assign n47338 = pi657 & pi1135;
  assign n47339 = pi1136 & ~n47337;
  assign n47340 = ~n47338 & n47339;
  assign n47341 = pi813 & n46731;
  assign n47342 = n46791 & n47341;
  assign n47343 = ~n47340 & ~n47342;
  assign n47344 = n47336 & ~n47343;
  assign n47345 = ~n47334 & ~n47344;
  assign n47346 = ~n8856 & ~n47345;
  assign po842 = n47327 | n47346;
  assign n47348 = ~pi1113 & po980;
  assign n47349 = pi686 & ~po980;
  assign n47350 = ~pi962 & ~n47348;
  assign po843 = ~n47349 & n47350;
  assign n47352 = ~pi687 & ~po980;
  assign n47353 = ~pi1127 & po980;
  assign n47354 = ~pi962 & ~n47352;
  assign po844 = ~n47353 & n47354;
  assign n47356 = ~pi1115 & po980;
  assign n47357 = pi688 & ~po980;
  assign n47358 = ~pi962 & ~n47356;
  assign po845 = ~n47357 & n47358;
  assign n47360 = pi351 & n47309;
  assign n47361 = pi376 & n46759;
  assign n47362 = ~n47360 & ~n47361;
  assign n47363 = ~pi591 & ~n47362;
  assign n47364 = pi401 & ~pi592;
  assign n47365 = n46757 & n47364;
  assign n47366 = ~n47363 & ~n47365;
  assign n47367 = ~pi588 & ~n47366;
  assign n47368 = pi426 & n46719;
  assign n47369 = n47318 & n47368;
  assign n47370 = ~n47367 & ~n47369;
  assign n47371 = n46709 & ~n47370;
  assign n47372 = ~pi199 & n42683;
  assign n47373 = pi199 & ~pi1079;
  assign n47374 = ~n46709 & ~n47373;
  assign n47375 = ~n47372 & n47374;
  assign n47376 = ~n47371 & ~n47375;
  assign n47377 = n8856 & ~n47376;
  assign n47378 = pi798 & n46791;
  assign n47379 = ~pi658 & ~pi1135;
  assign n47380 = pi655 & pi1135;
  assign n47381 = pi1136 & ~n47379;
  assign n47382 = ~n47380 & n47381;
  assign n47383 = ~n47378 & ~n47382;
  assign n47384 = n46732 & ~n47383;
  assign n47385 = pi752 & n46744;
  assign n47386 = ~pi703 & pi1135;
  assign n47387 = ~pi843 & ~pi1136;
  assign n47388 = ~n47386 & ~n47387;
  assign n47389 = n46748 & n47388;
  assign n47390 = ~n47385 & n47389;
  assign n47391 = ~n47384 & ~n47390;
  assign n47392 = ~n8856 & ~n47391;
  assign po846 = n47377 | n47392;
  assign n47394 = ~pi690 & ~po980;
  assign n47395 = ~pi1108 & po980;
  assign n47396 = ~pi962 & ~n47394;
  assign po847 = ~n47395 & n47396;
  assign n47398 = ~pi691 & ~po980;
  assign n47399 = ~pi1107 & po980;
  assign n47400 = ~pi962 & ~n47398;
  assign po848 = ~n47399 & n47400;
  assign n47402 = pi352 & n47309;
  assign n47403 = pi317 & n46759;
  assign n47404 = ~n47402 & ~n47403;
  assign n47405 = ~pi591 & ~n47404;
  assign n47406 = pi402 & ~pi592;
  assign n47407 = n46757 & n47406;
  assign n47408 = ~n47405 & ~n47407;
  assign n47409 = ~pi588 & ~n47408;
  assign n47410 = pi427 & n46719;
  assign n47411 = n47318 & n47410;
  assign n47412 = ~n47409 & ~n47411;
  assign n47413 = n46709 & ~n47412;
  assign n47414 = ~pi199 & n42695;
  assign n47415 = pi199 & ~pi1078;
  assign n47416 = ~n46709 & ~n47415;
  assign n47417 = ~n47414 & n47416;
  assign n47418 = ~n47413 & ~n47417;
  assign n47419 = n8856 & ~n47418;
  assign n47420 = ~pi726 & pi1135;
  assign n47421 = pi770 & ~pi1135;
  assign n47422 = pi1136 & ~n47420;
  assign n47423 = ~n47421 & n47422;
  assign n47424 = pi844 & n46791;
  assign n47425 = pi1134 & ~n47424;
  assign n47426 = ~n47423 & n47425;
  assign n47427 = ~pi656 & ~pi1135;
  assign n47428 = pi649 & pi1135;
  assign n47429 = pi1136 & ~n47427;
  assign n47430 = ~n47428 & n47429;
  assign n47431 = pi801 & n46791;
  assign n47432 = ~pi1134 & ~n47431;
  assign n47433 = ~n47430 & n47432;
  assign n47434 = n46795 & ~n47426;
  assign n47435 = ~n47433 & n47434;
  assign po849 = n47419 | n47435;
  assign n47437 = ~pi1129 & po954;
  assign n47438 = pi693 & ~po954;
  assign n47439 = ~pi962 & ~n47437;
  assign po850 = ~n47438 & n47439;
  assign n47441 = ~pi1128 & po980;
  assign n47442 = pi694 & ~po980;
  assign n47443 = ~pi962 & ~n47441;
  assign po851 = ~n47442 & n47443;
  assign n47445 = ~pi1111 & po954;
  assign n47446 = pi695 & ~po954;
  assign n47447 = ~pi962 & ~n47445;
  assign po852 = ~n47446 & n47447;
  assign n47449 = ~pi696 & ~po980;
  assign n47450 = ~pi1100 & po980;
  assign n47451 = ~pi962 & ~n47449;
  assign po853 = ~n47450 & n47451;
  assign n47453 = ~pi1129 & po980;
  assign n47454 = pi697 & ~po980;
  assign n47455 = ~pi962 & ~n47453;
  assign po854 = ~n47454 & n47455;
  assign n47457 = ~pi1116 & po980;
  assign n47458 = pi698 & ~po980;
  assign n47459 = ~pi962 & ~n47457;
  assign po855 = ~n47458 & n47459;
  assign n47461 = ~pi699 & ~po980;
  assign n47462 = ~pi1103 & po980;
  assign n47463 = ~pi962 & ~n47461;
  assign po856 = ~n47462 & n47463;
  assign n47465 = ~pi700 & ~po980;
  assign n47466 = ~pi1110 & po980;
  assign n47467 = ~pi962 & ~n47465;
  assign po857 = ~n47466 & n47467;
  assign n47469 = ~pi1123 & po980;
  assign n47470 = pi701 & ~po980;
  assign n47471 = ~pi962 & ~n47469;
  assign po858 = ~n47470 & n47471;
  assign n47473 = ~pi1117 & po980;
  assign n47474 = pi702 & ~po980;
  assign n47475 = ~pi962 & ~n47473;
  assign po859 = ~n47474 & n47475;
  assign n47477 = ~pi703 & ~po980;
  assign n47478 = ~pi1124 & po980;
  assign n47479 = ~pi962 & ~n47477;
  assign po860 = ~n47478 & n47479;
  assign n47481 = ~pi1112 & po980;
  assign n47482 = pi704 & ~po980;
  assign n47483 = ~pi962 & ~n47481;
  assign po861 = ~n47482 & n47483;
  assign n47485 = ~pi705 & ~po980;
  assign n47486 = ~pi1125 & po980;
  assign n47487 = ~pi962 & ~n47485;
  assign po862 = ~n47486 & n47487;
  assign n47489 = ~pi706 & ~po980;
  assign n47490 = ~pi1105 & po980;
  assign n47491 = ~pi962 & ~n47489;
  assign po863 = ~n47490 & n47491;
  assign n47493 = pi370 & n46713;
  assign n47494 = pi395 & pi591;
  assign n47495 = ~pi592 & n47494;
  assign n47496 = ~n47493 & ~n47495;
  assign n47497 = ~pi590 & ~n47496;
  assign n47498 = pi347 & n46720;
  assign n47499 = ~n47497 & ~n47498;
  assign n47500 = ~pi588 & n46709;
  assign n47501 = ~n47499 & n47500;
  assign n47502 = ~pi200 & ~pi304;
  assign n47503 = pi200 & ~pi1048;
  assign n47504 = ~n47502 & ~n47503;
  assign n47505 = ~pi199 & ~n47504;
  assign n47506 = pi199 & ~pi1055;
  assign n47507 = ~n46709 & ~n47506;
  assign n47508 = ~n47505 & n47507;
  assign n47509 = n46709 & n46724;
  assign n47510 = pi420 & pi588;
  assign n47511 = n47509 & n47510;
  assign n47512 = ~n47508 & ~n47511;
  assign n47513 = ~n47501 & n47512;
  assign n47514 = n8856 & ~n47513;
  assign n47515 = ~pi627 & pi1135;
  assign n47516 = ~pi618 & ~pi1135;
  assign n47517 = ~pi1134 & ~n47515;
  assign n47518 = ~n47516 & n47517;
  assign n47519 = n46940 & n47518;
  assign n47520 = pi753 & n46744;
  assign n47521 = pi702 & pi1135;
  assign n47522 = ~pi847 & ~pi1136;
  assign n47523 = ~n47521 & ~n47522;
  assign n47524 = n46748 & n47523;
  assign n47525 = ~n47520 & n47524;
  assign n47526 = ~n47519 & ~n47525;
  assign n47527 = ~n8856 & ~n47526;
  assign po864 = n47514 | n47527;
  assign n47529 = n46709 & n46713;
  assign n47530 = pi442 & n47529;
  assign n47531 = ~pi592 & n46709;
  assign n47532 = pi328 & pi591;
  assign n47533 = n47531 & n47532;
  assign n47534 = ~n47530 & ~n47533;
  assign n47535 = ~pi590 & ~n47534;
  assign n47536 = pi321 & n46709;
  assign n47537 = n46720 & n47536;
  assign n47538 = ~n47535 & ~n47537;
  assign n47539 = ~pi588 & ~n47538;
  assign n47540 = ~pi200 & ~pi305;
  assign n47541 = pi200 & ~pi1084;
  assign n47542 = ~n47540 & ~n47541;
  assign n47543 = ~pi199 & ~n47542;
  assign n47544 = pi199 & ~pi1058;
  assign n47545 = ~n46709 & ~n47544;
  assign n47546 = ~n47543 & n47545;
  assign n47547 = n46709 & n46719;
  assign n47548 = pi459 & n47318;
  assign n47549 = n47547 & n47548;
  assign n47550 = n8856 & ~n47549;
  assign n47551 = ~n47546 & n47550;
  assign n47552 = ~n47539 & n47551;
  assign n47553 = pi754 & n46744;
  assign n47554 = n46731 & ~n46746;
  assign n47555 = pi709 & pi1135;
  assign n47556 = ~pi857 & ~pi1136;
  assign n47557 = pi1134 & ~n47555;
  assign n47558 = ~n47556 & n47557;
  assign n47559 = n47554 & n47558;
  assign n47560 = ~n47553 & n47559;
  assign n47561 = ~pi609 & ~pi1135;
  assign n47562 = ~pi660 & pi1135;
  assign n47563 = ~pi1134 & ~n47561;
  assign n47564 = ~n47562 & n47563;
  assign n47565 = n46940 & n47564;
  assign n47566 = ~n8856 & ~n47565;
  assign n47567 = ~n47560 & n47566;
  assign po865 = ~n47552 & ~n47567;
  assign n47569 = ~pi1118 & po980;
  assign n47570 = pi709 & ~po980;
  assign n47571 = ~pi962 & ~n47569;
  assign po866 = ~n47570 & n47571;
  assign n47573 = ~pi710 & ~po954;
  assign n47574 = ~pi1106 & po954;
  assign n47575 = ~pi962 & ~n47573;
  assign po867 = ~n47574 & n47575;
  assign n47577 = pi373 & n46713;
  assign n47578 = pi398 & pi591;
  assign n47579 = ~pi592 & n47578;
  assign n47580 = ~n47577 & ~n47579;
  assign n47581 = ~pi590 & ~n47580;
  assign n47582 = pi348 & n46720;
  assign n47583 = ~n47581 & ~n47582;
  assign n47584 = n47500 & ~n47583;
  assign n47585 = ~pi200 & ~pi306;
  assign n47586 = pi200 & ~pi1059;
  assign n47587 = ~n47585 & ~n47586;
  assign n47588 = ~pi199 & ~n47587;
  assign n47589 = pi199 & ~pi1087;
  assign n47590 = ~n46709 & ~n47589;
  assign n47591 = ~n47588 & n47590;
  assign n47592 = pi423 & pi588;
  assign n47593 = n47509 & n47592;
  assign n47594 = ~n47591 & ~n47593;
  assign n47595 = ~n47584 & n47594;
  assign n47596 = n8856 & ~n47595;
  assign n47597 = ~pi647 & pi1135;
  assign n47598 = ~pi630 & ~pi1135;
  assign n47599 = ~pi1134 & ~n47597;
  assign n47600 = ~n47598 & n47599;
  assign n47601 = n46940 & n47600;
  assign n47602 = pi755 & n46744;
  assign n47603 = pi725 & pi1135;
  assign n47604 = ~pi858 & ~pi1136;
  assign n47605 = ~n47603 & ~n47604;
  assign n47606 = n46748 & n47605;
  assign n47607 = ~n47602 & n47606;
  assign n47608 = ~n47601 & ~n47607;
  assign n47609 = ~n8856 & ~n47608;
  assign po868 = n47596 | n47609;
  assign n47611 = pi751 & n46744;
  assign n47612 = pi701 & pi1135;
  assign n47613 = ~pi842 & ~pi1136;
  assign n47614 = pi1134 & ~n47612;
  assign n47615 = ~n47613 & n47614;
  assign n47616 = n47554 & n47615;
  assign n47617 = ~n47611 & n47616;
  assign n47618 = ~pi715 & pi1135;
  assign n47619 = ~pi644 & ~pi1135;
  assign n47620 = ~pi1134 & ~n47618;
  assign n47621 = ~n47619 & n47620;
  assign n47622 = n46940 & n47621;
  assign n47623 = ~n47617 & ~n47622;
  assign n47624 = ~n8856 & ~n47623;
  assign n47625 = pi374 & n46713;
  assign n47626 = pi400 & pi591;
  assign n47627 = ~pi592 & n47626;
  assign n47628 = ~n47625 & ~n47627;
  assign n47629 = ~pi590 & ~n47628;
  assign n47630 = pi350 & n46720;
  assign n47631 = ~n47629 & ~n47630;
  assign n47632 = ~pi588 & ~n47631;
  assign n47633 = pi425 & n46719;
  assign n47634 = n47318 & n47633;
  assign n47635 = n46709 & ~n47634;
  assign n47636 = ~n47632 & n47635;
  assign n47637 = pi298 & n10793;
  assign n47638 = pi1044 & n11419;
  assign n47639 = pi199 & pi1035;
  assign n47640 = ~n46709 & ~n47639;
  assign n47641 = ~n47637 & n47640;
  assign n47642 = ~n47638 & n47641;
  assign n47643 = n8856 & ~n47642;
  assign n47644 = ~n47636 & n47643;
  assign po869 = n47624 | n47644;
  assign n47646 = pi371 & n46713;
  assign n47647 = pi396 & pi591;
  assign n47648 = ~pi592 & n47647;
  assign n47649 = ~n47646 & ~n47648;
  assign n47650 = ~pi590 & ~n47649;
  assign n47651 = pi322 & n46720;
  assign n47652 = ~n47650 & ~n47651;
  assign n47653 = n47500 & ~n47652;
  assign n47654 = ~pi200 & ~pi309;
  assign n47655 = pi200 & ~pi1072;
  assign n47656 = ~n47654 & ~n47655;
  assign n47657 = ~pi199 & ~n47656;
  assign n47658 = pi199 & ~pi1051;
  assign n47659 = ~n46709 & ~n47658;
  assign n47660 = ~n47657 & n47659;
  assign n47661 = pi421 & pi588;
  assign n47662 = n47509 & n47661;
  assign n47663 = ~n47660 & ~n47662;
  assign n47664 = ~n47653 & n47663;
  assign n47665 = n8856 & ~n47664;
  assign n47666 = ~pi628 & pi1135;
  assign n47667 = ~pi629 & ~pi1135;
  assign n47668 = ~pi1134 & ~n47666;
  assign n47669 = ~n47667 & n47668;
  assign n47670 = n46940 & n47669;
  assign n47671 = pi756 & n46744;
  assign n47672 = pi734 & pi1135;
  assign n47673 = ~pi854 & ~pi1136;
  assign n47674 = ~n47672 & ~n47673;
  assign n47675 = n46748 & n47674;
  assign n47676 = ~n47671 & n47675;
  assign n47677 = ~n47670 & ~n47676;
  assign n47678 = ~n8856 & ~n47677;
  assign po870 = n47665 | n47678;
  assign n47680 = pi461 & n47309;
  assign n47681 = pi439 & n46759;
  assign n47682 = ~n47680 & ~n47681;
  assign n47683 = ~pi591 & ~n47682;
  assign n47684 = pi326 & ~pi592;
  assign n47685 = n46757 & n47684;
  assign n47686 = ~n47683 & ~n47685;
  assign n47687 = ~pi588 & ~n47686;
  assign n47688 = pi449 & n46719;
  assign n47689 = n47318 & n47688;
  assign n47690 = ~n47687 & ~n47689;
  assign n47691 = n46709 & ~n47690;
  assign n47692 = pi199 & ~pi1057;
  assign n47693 = ~n46709 & ~n47692;
  assign n47694 = ~n42175 & n47693;
  assign n47695 = ~n47691 & ~n47694;
  assign n47696 = n8856 & ~n47695;
  assign n47697 = pi867 & n46791;
  assign n47698 = pi762 & ~pi1135;
  assign n47699 = pi697 & pi1135;
  assign n47700 = pi1136 & ~n47698;
  assign n47701 = ~n47699 & n47700;
  assign n47702 = ~n47697 & ~n47701;
  assign n47703 = n46747 & ~n47702;
  assign n47704 = ~pi653 & ~pi1135;
  assign n47705 = pi693 & pi1135;
  assign n47706 = pi1136 & ~n47704;
  assign n47707 = ~n47705 & n47706;
  assign n47708 = pi816 & n46731;
  assign n47709 = n46791 & n47708;
  assign n47710 = ~n47707 & ~n47709;
  assign n47711 = n47336 & ~n47710;
  assign n47712 = ~n47703 & ~n47711;
  assign n47713 = ~n8856 & ~n47712;
  assign po871 = n47696 | n47713;
  assign n47715 = ~pi715 & ~po954;
  assign n47716 = ~pi1123 & po954;
  assign n47717 = ~pi962 & ~n47715;
  assign po872 = ~n47716 & n47717;
  assign n47719 = pi440 & n47529;
  assign n47720 = pi329 & pi591;
  assign n47721 = n47531 & n47720;
  assign n47722 = ~n47719 & ~n47721;
  assign n47723 = ~pi590 & ~n47722;
  assign n47724 = pi349 & n46709;
  assign n47725 = n46720 & n47724;
  assign n47726 = ~n47723 & ~n47725;
  assign n47727 = ~pi588 & ~n47726;
  assign n47728 = ~pi200 & ~pi307;
  assign n47729 = pi200 & ~pi1053;
  assign n47730 = ~n47728 & ~n47729;
  assign n47731 = ~pi199 & ~n47730;
  assign n47732 = pi199 & ~pi1043;
  assign n47733 = ~n46709 & ~n47732;
  assign n47734 = ~n47731 & n47733;
  assign n47735 = pi454 & n47318;
  assign n47736 = n47547 & n47735;
  assign n47737 = n8856 & ~n47736;
  assign n47738 = ~n47734 & n47737;
  assign n47739 = ~n47727 & n47738;
  assign n47740 = pi761 & n46744;
  assign n47741 = pi738 & pi1135;
  assign n47742 = ~pi845 & ~pi1136;
  assign n47743 = pi1134 & ~n47741;
  assign n47744 = ~n47742 & n47743;
  assign n47745 = n47554 & n47744;
  assign n47746 = ~n47740 & n47745;
  assign n47747 = ~pi626 & ~pi1135;
  assign n47748 = ~pi641 & pi1135;
  assign n47749 = ~pi1134 & ~n47747;
  assign n47750 = ~n47748 & n47749;
  assign n47751 = n46940 & n47750;
  assign n47752 = ~n8856 & ~n47751;
  assign n47753 = ~n47746 & n47752;
  assign po873 = ~n47739 & ~n47753;
  assign n47755 = pi318 & pi591;
  assign n47756 = ~pi592 & n47755;
  assign n47757 = ~pi591 & n7772;
  assign n47758 = ~n47756 & ~n47757;
  assign n47759 = ~pi590 & ~n47758;
  assign n47760 = pi462 & n46720;
  assign n47761 = ~n47759 & ~n47760;
  assign n47762 = n47500 & ~n47761;
  assign n47763 = ~pi199 & n42689;
  assign n47764 = pi199 & ~pi1074;
  assign n47765 = ~n46709 & ~n47764;
  assign n47766 = ~n47763 & n47765;
  assign n47767 = pi448 & pi588;
  assign n47768 = n47509 & n47767;
  assign n47769 = ~n47766 & ~n47768;
  assign n47770 = ~n47762 & n47769;
  assign n47771 = n8856 & ~n47770;
  assign n47772 = pi768 & n46744;
  assign n47773 = ~pi705 & pi1135;
  assign n47774 = ~pi839 & ~pi1136;
  assign n47775 = pi1134 & ~n47773;
  assign n47776 = ~n47774 & n47775;
  assign n47777 = n47554 & n47776;
  assign n47778 = ~n47772 & n47777;
  assign n47779 = pi800 & n46791;
  assign n47780 = ~pi645 & ~pi1135;
  assign n47781 = pi669 & pi1135;
  assign n47782 = pi1136 & ~n47780;
  assign n47783 = ~n47781 & n47782;
  assign n47784 = ~n47779 & ~n47783;
  assign n47785 = n46732 & ~n47784;
  assign n47786 = ~n47778 & ~n47785;
  assign n47787 = ~n8856 & ~n47786;
  assign po874 = n47771 | n47787;
  assign n47789 = pi369 & n47529;
  assign n47790 = pi394 & pi591;
  assign n47791 = n47531 & n47790;
  assign n47792 = ~n47789 & ~n47791;
  assign n47793 = ~pi590 & ~n47792;
  assign n47794 = pi315 & n46709;
  assign n47795 = n46720 & n47794;
  assign n47796 = ~n47793 & ~n47795;
  assign n47797 = ~pi588 & ~n47796;
  assign n47798 = ~pi200 & ~pi303;
  assign n47799 = pi200 & ~pi1049;
  assign n47800 = ~n47798 & ~n47799;
  assign n47801 = ~pi199 & ~n47800;
  assign n47802 = pi199 & ~pi1080;
  assign n47803 = ~n46709 & ~n47802;
  assign n47804 = ~n47801 & n47803;
  assign n47805 = pi419 & n47318;
  assign n47806 = n47547 & n47805;
  assign n47807 = n8856 & ~n47806;
  assign n47808 = ~n47804 & n47807;
  assign n47809 = ~n47797 & n47808;
  assign n47810 = pi767 & n46744;
  assign n47811 = pi698 & pi1135;
  assign n47812 = ~pi853 & ~pi1136;
  assign n47813 = pi1134 & ~n47811;
  assign n47814 = ~n47812 & n47813;
  assign n47815 = n47554 & n47814;
  assign n47816 = ~n47810 & n47815;
  assign n47817 = ~pi608 & ~pi1135;
  assign n47818 = ~pi625 & pi1135;
  assign n47819 = ~pi1134 & ~n47817;
  assign n47820 = ~n47818 & n47819;
  assign n47821 = n46940 & n47820;
  assign n47822 = ~n8856 & ~n47821;
  assign n47823 = ~n47816 & n47822;
  assign po875 = ~n47809 & ~n47823;
  assign n47825 = pi378 & n46713;
  assign n47826 = pi325 & pi591;
  assign n47827 = ~pi592 & n47826;
  assign n47828 = ~n47825 & ~n47827;
  assign n47829 = ~pi590 & ~n47828;
  assign n47830 = pi353 & n46720;
  assign n47831 = ~n47829 & ~n47830;
  assign n47832 = n47500 & ~n47831;
  assign n47833 = ~pi199 & n42701;
  assign n47834 = pi199 & ~pi1063;
  assign n47835 = ~n46709 & ~n47834;
  assign n47836 = ~n47833 & n47835;
  assign n47837 = pi451 & pi588;
  assign n47838 = n47509 & n47837;
  assign n47839 = ~n47836 & ~n47838;
  assign n47840 = ~n47832 & n47839;
  assign n47841 = n8856 & ~n47840;
  assign n47842 = pi774 & n46744;
  assign n47843 = ~pi687 & pi1135;
  assign n47844 = ~pi868 & ~pi1136;
  assign n47845 = pi1134 & ~n47843;
  assign n47846 = ~n47844 & n47845;
  assign n47847 = n47554 & n47846;
  assign n47848 = ~n47842 & n47847;
  assign n47849 = pi807 & n46791;
  assign n47850 = ~pi636 & ~pi1135;
  assign n47851 = pi650 & pi1135;
  assign n47852 = pi1136 & ~n47850;
  assign n47853 = ~n47851 & n47852;
  assign n47854 = ~n47849 & ~n47853;
  assign n47855 = n46732 & ~n47854;
  assign n47856 = ~n47848 & ~n47855;
  assign n47857 = ~n8856 & ~n47856;
  assign po876 = n47841 | n47857;
  assign n47859 = pi356 & n47309;
  assign n47860 = pi381 & n46759;
  assign n47861 = ~n47859 & ~n47860;
  assign n47862 = ~pi591 & ~n47861;
  assign n47863 = pi405 & ~pi592;
  assign n47864 = n46757 & n47863;
  assign n47865 = ~n47862 & ~n47864;
  assign n47866 = ~pi588 & ~n47865;
  assign n47867 = pi445 & n46719;
  assign n47868 = n47318 & n47867;
  assign n47869 = ~n47866 & ~n47868;
  assign n47870 = n46709 & ~n47869;
  assign n47871 = pi199 & ~pi1081;
  assign n47872 = ~n46709 & ~n47871;
  assign n47873 = ~n42721 & n47872;
  assign n47874 = ~n47870 & ~n47873;
  assign n47875 = n8856 & ~n47874;
  assign n47876 = pi880 & n46791;
  assign n47877 = pi750 & ~pi1135;
  assign n47878 = pi684 & pi1135;
  assign n47879 = pi1136 & ~n47877;
  assign n47880 = ~n47878 & n47879;
  assign n47881 = ~n47876 & ~n47880;
  assign n47882 = n46747 & ~n47881;
  assign n47883 = ~pi651 & ~pi1135;
  assign n47884 = pi654 & pi1135;
  assign n47885 = pi1136 & ~n47883;
  assign n47886 = ~n47884 & n47885;
  assign n47887 = pi794 & n46731;
  assign n47888 = n46791 & n47887;
  assign n47889 = ~n47886 & ~n47888;
  assign n47890 = n47336 & ~n47889;
  assign n47891 = ~n47882 & ~n47890;
  assign n47892 = ~n8856 & ~n47891;
  assign po877 = n47875 | n47892;
  assign n47894 = pi747 & pi773;
  assign n47895 = pi769 & n47894;
  assign n47896 = pi721 & n47895;
  assign n47897 = ~pi721 & ~n47895;
  assign n47898 = pi775 & ~n47896;
  assign n47899 = ~n47897 & n47898;
  assign n47900 = pi721 & pi813;
  assign n47901 = ~pi773 & ~pi801;
  assign n47902 = pi773 & pi801;
  assign n47903 = ~n47901 & ~n47902;
  assign n47904 = ~pi771 & ~pi800;
  assign n47905 = pi771 & pi800;
  assign n47906 = ~n47904 & ~n47905;
  assign n47907 = ~pi769 & ~pi794;
  assign n47908 = pi769 & pi794;
  assign n47909 = ~n47907 & ~n47908;
  assign n47910 = ~pi765 & ~pi798;
  assign n47911 = pi765 & pi798;
  assign n47912 = ~n47910 & ~n47911;
  assign n47913 = pi807 & ~n47912;
  assign n47914 = pi747 & n47913;
  assign n47915 = ~pi747 & ~pi807;
  assign n47916 = ~n47912 & n47915;
  assign n47917 = ~n47914 & ~n47916;
  assign n47918 = ~n47909 & ~n47917;
  assign n47919 = ~n47906 & n47918;
  assign n47920 = ~n47903 & n47919;
  assign n47921 = n47900 & n47920;
  assign n47922 = ~n47906 & n47913;
  assign n47923 = ~pi721 & ~pi813;
  assign n47924 = pi794 & pi801;
  assign n47925 = n47923 & n47924;
  assign n47926 = n47922 & n47925;
  assign n47927 = ~n47921 & ~n47926;
  assign n47928 = pi816 & ~n47927;
  assign n47929 = n47899 & ~n47928;
  assign n47930 = pi795 & ~n47929;
  assign n47931 = ~pi945 & pi988;
  assign n47932 = pi731 & n47931;
  assign n47933 = pi721 & ~pi775;
  assign n47934 = ~n47899 & ~n47933;
  assign n47935 = n47932 & ~n47934;
  assign n47936 = ~n47930 & n47935;
  assign n47937 = ~pi775 & ~pi816;
  assign n47938 = pi775 & pi816;
  assign n47939 = ~n47937 & ~n47938;
  assign n47940 = n47921 & ~n47939;
  assign n47941 = n47933 & ~n47940;
  assign n47942 = ~pi731 & ~pi795;
  assign n47943 = pi731 & pi795;
  assign n47944 = ~n47942 & ~n47943;
  assign n47945 = n47940 & ~n47944;
  assign n47946 = pi721 & ~n47932;
  assign n47947 = ~n47945 & n47946;
  assign n47948 = ~n47941 & ~n47947;
  assign po878 = n47936 | ~n47948;
  assign n47950 = pi379 & n46713;
  assign n47951 = pi403 & pi591;
  assign n47952 = ~pi592 & n47951;
  assign n47953 = ~n47950 & ~n47952;
  assign n47954 = ~pi590 & ~n47953;
  assign n47955 = pi354 & n46720;
  assign n47956 = ~n47954 & ~n47955;
  assign n47957 = n47500 & ~n47956;
  assign n47958 = ~pi199 & n42707;
  assign n47959 = pi199 & ~pi1045;
  assign n47960 = ~n46709 & ~n47959;
  assign n47961 = ~n47958 & n47960;
  assign n47962 = pi428 & pi588;
  assign n47963 = n47509 & n47962;
  assign n47964 = ~n47961 & ~n47963;
  assign n47965 = ~n47957 & n47964;
  assign n47966 = n8856 & ~n47965;
  assign n47967 = ~pi795 & ~pi1134;
  assign n47968 = ~pi851 & pi1134;
  assign n47969 = ~pi1136 & ~n47967;
  assign n47970 = ~n47968 & n47969;
  assign n47971 = ~pi640 & ~pi1134;
  assign n47972 = pi776 & pi1134;
  assign n47973 = pi1136 & ~n47971;
  assign n47974 = ~n47972 & n47973;
  assign n47975 = ~n47970 & ~n47974;
  assign n47976 = ~pi1135 & ~n47975;
  assign n47977 = pi694 & pi1134;
  assign n47978 = pi732 & ~pi1134;
  assign n47979 = pi1135 & pi1136;
  assign n47980 = ~n47977 & n47979;
  assign n47981 = ~n47978 & n47980;
  assign n47982 = ~n47976 & ~n47981;
  assign n47983 = n46795 & ~n47982;
  assign po879 = n47966 | n47983;
  assign n47985 = ~pi1111 & po980;
  assign n47986 = pi723 & ~po980;
  assign n47987 = ~pi962 & ~n47985;
  assign po880 = ~n47986 & n47987;
  assign n47989 = ~pi1114 & po980;
  assign n47990 = pi724 & ~po980;
  assign n47991 = ~pi962 & ~n47989;
  assign po881 = ~n47990 & n47991;
  assign n47993 = ~pi1120 & po980;
  assign n47994 = pi725 & ~po980;
  assign n47995 = ~pi962 & ~n47993;
  assign po882 = ~n47994 & n47995;
  assign n47997 = ~pi726 & ~po980;
  assign n47998 = ~pi1126 & po980;
  assign n47999 = ~pi962 & ~n47997;
  assign po883 = ~n47998 & n47999;
  assign n48001 = ~pi727 & ~po980;
  assign n48002 = ~pi1102 & po980;
  assign n48003 = ~pi962 & ~n48001;
  assign po884 = ~n48002 & n48003;
  assign n48005 = ~pi1131 & po980;
  assign n48006 = pi728 & ~po980;
  assign n48007 = ~pi962 & ~n48005;
  assign po885 = ~n48006 & n48007;
  assign n48009 = ~pi729 & ~po980;
  assign n48010 = ~pi1104 & po980;
  assign n48011 = ~pi962 & ~n48009;
  assign po886 = ~n48010 & n48011;
  assign n48013 = ~pi730 & ~po980;
  assign n48014 = ~pi1106 & po980;
  assign n48015 = ~pi962 & ~n48013;
  assign po887 = ~n48014 & n48015;
  assign n48017 = ~n47900 & ~n47923;
  assign n48018 = n47920 & ~n48017;
  assign n48019 = pi795 & ~n47939;
  assign n48020 = n48018 & n48019;
  assign n48021 = ~n47894 & ~n48020;
  assign n48022 = n47932 & ~n48021;
  assign n48023 = pi731 & ~n48020;
  assign n48024 = ~n47939 & ~n48017;
  assign n48025 = ~pi795 & pi801;
  assign n48026 = ~n47909 & n48025;
  assign n48027 = n48024 & n48026;
  assign n48028 = n47922 & n48027;
  assign n48029 = n47894 & ~n48028;
  assign n48030 = ~pi731 & ~n48029;
  assign n48031 = n47931 & ~n48030;
  assign n48032 = ~n48023 & ~n48031;
  assign po888 = ~n48022 & ~n48032;
  assign n48034 = ~pi1128 & po954;
  assign n48035 = pi732 & ~po954;
  assign n48036 = ~pi962 & ~n48034;
  assign po889 = ~n48035 & n48036;
  assign n48038 = pi375 & n47529;
  assign n48039 = pi399 & pi591;
  assign n48040 = n47531 & n48039;
  assign n48041 = ~n48038 & ~n48040;
  assign n48042 = ~pi590 & ~n48041;
  assign n48043 = pi316 & n46709;
  assign n48044 = n46720 & n48043;
  assign n48045 = ~n48042 & ~n48044;
  assign n48046 = ~pi588 & ~n48045;
  assign n48047 = ~pi200 & ~pi308;
  assign n48048 = pi200 & ~pi1037;
  assign n48049 = ~n48047 & ~n48048;
  assign n48050 = ~pi199 & ~n48049;
  assign n48051 = pi199 & ~pi1047;
  assign n48052 = ~n46709 & ~n48051;
  assign n48053 = ~n48050 & n48052;
  assign n48054 = pi424 & n47318;
  assign n48055 = n47547 & n48054;
  assign n48056 = n8856 & ~n48055;
  assign n48057 = ~n48053 & n48056;
  assign n48058 = ~n48046 & n48057;
  assign n48059 = pi777 & n46744;
  assign n48060 = pi737 & pi1135;
  assign n48061 = ~pi838 & ~pi1136;
  assign n48062 = pi1134 & ~n48060;
  assign n48063 = ~n48061 & n48062;
  assign n48064 = n47554 & n48063;
  assign n48065 = ~n48059 & n48064;
  assign n48066 = ~pi619 & ~pi1135;
  assign n48067 = ~pi648 & pi1135;
  assign n48068 = ~pi1134 & ~n48066;
  assign n48069 = ~n48067 & n48068;
  assign n48070 = n46940 & n48069;
  assign n48071 = ~n8856 & ~n48070;
  assign n48072 = ~n48065 & n48071;
  assign po890 = ~n48058 & ~n48072;
  assign n48074 = ~pi1119 & po980;
  assign n48075 = pi734 & ~po980;
  assign n48076 = ~pi962 & ~n48074;
  assign po891 = ~n48075 & n48076;
  assign n48078 = ~pi735 & ~po980;
  assign n48079 = ~pi1109 & po980;
  assign n48080 = ~pi962 & ~n48078;
  assign po892 = ~n48079 & n48080;
  assign n48082 = ~pi736 & ~po980;
  assign n48083 = ~pi1101 & po980;
  assign n48084 = ~pi962 & ~n48082;
  assign po893 = ~n48083 & n48084;
  assign n48086 = ~pi1122 & po980;
  assign n48087 = pi737 & ~po980;
  assign n48088 = ~pi962 & ~n48086;
  assign po894 = ~n48087 & n48088;
  assign n48090 = ~pi1121 & po980;
  assign n48091 = pi738 & ~po980;
  assign n48092 = ~pi962 & ~n48090;
  assign po895 = ~n48091 & n48092;
  assign n48094 = ~pi952 & ~pi1061;
  assign n48095 = n46435 & n48094;
  assign po988 = pi832 & n48095;
  assign n48097 = pi1108 & po988;
  assign n48098 = pi739 & ~po988;
  assign n48099 = ~pi966 & ~n48097;
  assign po896 = n48098 | ~n48099;
  assign n48101 = ~pi741 & ~po988;
  assign n48102 = pi1114 & po988;
  assign n48103 = ~pi966 & ~n48101;
  assign po898 = n48102 | ~n48103;
  assign n48105 = ~pi742 & ~po988;
  assign n48106 = pi1112 & po988;
  assign n48107 = ~pi966 & ~n48105;
  assign po899 = n48106 | ~n48107;
  assign n48109 = pi1109 & po988;
  assign n48110 = pi743 & ~po988;
  assign n48111 = ~pi966 & ~n48109;
  assign po900 = n48110 | ~n48111;
  assign n48113 = ~pi744 & ~po988;
  assign n48114 = pi1131 & po988;
  assign n48115 = ~pi966 & ~n48113;
  assign po901 = n48114 | ~n48115;
  assign n48117 = ~pi745 & ~po988;
  assign n48118 = pi1111 & po988;
  assign n48119 = ~pi966 & ~n48117;
  assign po902 = n48118 | ~n48119;
  assign n48121 = pi1104 & po988;
  assign n48122 = pi746 & ~po988;
  assign n48123 = ~pi966 & ~n48121;
  assign po903 = n48122 | ~n48123;
  assign n48125 = pi801 & n47916;
  assign n48126 = pi773 & n47931;
  assign n48127 = ~n47903 & ~n48126;
  assign n48128 = n47913 & n48127;
  assign n48129 = ~n48125 & ~n48128;
  assign n48130 = ~n47944 & n48024;
  assign n48131 = ~n47906 & ~n47909;
  assign n48132 = n48130 & n48131;
  assign n48133 = ~n48129 & n48132;
  assign n48134 = ~pi747 & ~n48126;
  assign n48135 = n47894 & n47931;
  assign n48136 = ~n48134 & ~n48135;
  assign po904 = ~n48133 & n48136;
  assign n48138 = pi1106 & po988;
  assign n48139 = pi748 & ~po988;
  assign n48140 = ~pi966 & ~n48138;
  assign po905 = n48139 | ~n48140;
  assign n48142 = pi1105 & po988;
  assign n48143 = pi749 & ~po988;
  assign n48144 = ~pi966 & ~n48142;
  assign po906 = n48143 | ~n48144;
  assign n48146 = ~pi750 & ~po988;
  assign n48147 = pi1130 & po988;
  assign n48148 = ~pi966 & ~n48146;
  assign po907 = n48147 | ~n48148;
  assign n48150 = ~pi751 & ~po988;
  assign n48151 = pi1123 & po988;
  assign n48152 = ~pi966 & ~n48150;
  assign po908 = n48151 | ~n48152;
  assign n48154 = ~pi752 & ~po988;
  assign n48155 = pi1124 & po988;
  assign n48156 = ~pi966 & ~n48154;
  assign po909 = n48155 | ~n48156;
  assign n48158 = ~pi753 & ~po988;
  assign n48159 = pi1117 & po988;
  assign n48160 = ~pi966 & ~n48158;
  assign po910 = n48159 | ~n48160;
  assign n48162 = ~pi754 & ~po988;
  assign n48163 = pi1118 & po988;
  assign n48164 = ~pi966 & ~n48162;
  assign po911 = n48163 | ~n48164;
  assign n48166 = ~pi755 & ~po988;
  assign n48167 = pi1120 & po988;
  assign n48168 = ~pi966 & ~n48166;
  assign po912 = n48167 | ~n48168;
  assign n48170 = ~pi756 & ~po988;
  assign n48171 = pi1119 & po988;
  assign n48172 = ~pi966 & ~n48170;
  assign po913 = n48171 | ~n48172;
  assign n48174 = ~pi757 & ~po988;
  assign n48175 = pi1113 & po988;
  assign n48176 = ~pi966 & ~n48174;
  assign po914 = n48175 | ~n48176;
  assign n48178 = pi1101 & po988;
  assign n48179 = pi758 & ~po988;
  assign n48180 = ~pi966 & ~n48178;
  assign po915 = n48179 | ~n48180;
  assign n48182 = ~pi759 & ~po988;
  assign n48183 = n46440 & n48095;
  assign n48184 = ~n48182 & ~n48183;
  assign po916 = pi966 | n48184;
  assign n48186 = ~pi760 & ~po988;
  assign n48187 = pi1115 & po988;
  assign n48188 = ~pi966 & ~n48186;
  assign po917 = n48187 | ~n48188;
  assign n48190 = ~pi761 & ~po988;
  assign n48191 = pi1121 & po988;
  assign n48192 = ~pi966 & ~n48190;
  assign po918 = n48191 | ~n48192;
  assign n48194 = ~pi762 & ~po988;
  assign n48195 = pi1129 & po988;
  assign n48196 = ~pi966 & ~n48194;
  assign po919 = n48195 | ~n48196;
  assign n48198 = pi1103 & po988;
  assign n48199 = pi763 & ~po988;
  assign n48200 = ~pi966 & ~n48198;
  assign po920 = n48199 | ~n48200;
  assign n48202 = pi1107 & po988;
  assign n48203 = pi764 & ~po988;
  assign n48204 = ~pi966 & ~n48202;
  assign po921 = n48203 | ~n48204;
  assign po978 = n47920 & n48130;
  assign n48207 = pi765 & ~po978;
  assign n48208 = pi945 & ~n48207;
  assign n48209 = ~pi765 & ~n47905;
  assign n48210 = ~n47908 & n48209;
  assign n48211 = ~n47914 & n48210;
  assign n48212 = n47901 & ~n48211;
  assign n48213 = ~n47902 & ~n48212;
  assign n48214 = n47919 & ~n48213;
  assign n48215 = ~pi721 & ~n48214;
  assign n48216 = n47937 & ~n48215;
  assign n48217 = ~n47938 & ~n48216;
  assign n48218 = n47942 & ~n48217;
  assign n48219 = ~n47939 & n47943;
  assign n48220 = ~n48218 & ~n48219;
  assign po963 = n48018 & ~n48220;
  assign n48222 = ~pi765 & ~po963;
  assign n48223 = ~pi945 & ~n48222;
  assign po922 = ~n48208 & ~n48223;
  assign n48225 = pi1110 & po988;
  assign n48226 = pi766 & ~po988;
  assign n48227 = ~pi966 & ~n48225;
  assign po923 = n48226 | ~n48227;
  assign n48229 = ~pi767 & ~po988;
  assign n48230 = pi1116 & po988;
  assign n48231 = ~pi966 & ~n48229;
  assign po924 = n48230 | ~n48231;
  assign n48233 = ~pi768 & ~po988;
  assign n48234 = pi1125 & po988;
  assign n48235 = ~pi966 & ~n48233;
  assign po925 = n48234 | ~n48235;
  assign n48237 = n47938 & n48018;
  assign n48238 = pi794 & ~n47903;
  assign n48239 = ~n47906 & n48238;
  assign n48240 = n48024 & n48239;
  assign n48241 = ~n47917 & n48240;
  assign n48242 = ~pi775 & n48241;
  assign n48243 = ~n48237 & ~n48242;
  assign n48244 = pi795 & ~n48243;
  assign n48245 = pi775 & n47894;
  assign n48246 = pi769 & ~n48245;
  assign n48247 = ~pi769 & n48245;
  assign n48248 = ~n48246 & ~n48247;
  assign n48249 = n47932 & ~n48248;
  assign n48250 = ~n48244 & n48249;
  assign n48251 = ~n47944 & n48241;
  assign n48252 = pi769 & ~n47932;
  assign n48253 = ~n48251 & n48252;
  assign po926 = n48250 | n48253;
  assign n48255 = ~pi770 & ~po988;
  assign n48256 = pi1126 & po988;
  assign n48257 = ~pi966 & ~n48255;
  assign po927 = n48256 | ~n48257;
  assign n48259 = ~pi945 & pi987;
  assign n48260 = ~po963 & n48259;
  assign n48261 = pi771 & pi945;
  assign n48262 = ~po978 & n48261;
  assign po928 = n48260 | n48262;
  assign n48264 = pi1102 & po988;
  assign n48265 = pi772 & ~po988;
  assign n48266 = ~pi966 & ~n48264;
  assign po929 = n48265 | ~n48266;
  assign n48268 = ~pi801 & n47919;
  assign n48269 = po963 & n48268;
  assign n48270 = n47931 & ~n48269;
  assign n48271 = pi801 & ~n48130;
  assign n48272 = n47920 & ~n48271;
  assign n48273 = pi773 & ~n48272;
  assign n48274 = ~n48270 & ~n48273;
  assign po930 = ~n48126 & ~n48274;
  assign n48276 = ~pi774 & ~po988;
  assign n48277 = pi1127 & po988;
  assign n48278 = ~pi966 & ~n48276;
  assign po931 = n48277 | ~n48278;
  assign n48280 = pi775 & ~po978;
  assign n48281 = pi731 & ~pi945;
  assign n48282 = pi765 & pi771;
  assign n48283 = n47894 & n48282;
  assign n48284 = pi795 & pi800;
  assign n48285 = pi801 & ~pi816;
  assign n48286 = n48284 & n48285;
  assign n48287 = ~n48017 & n48286;
  assign n48288 = n47918 & n48287;
  assign n48289 = n48283 & ~n48288;
  assign n48290 = ~pi775 & ~n48289;
  assign n48291 = n48281 & ~n48290;
  assign n48292 = ~n48280 & ~n48291;
  assign n48293 = ~n48020 & ~n48283;
  assign n48294 = pi775 & n48281;
  assign n48295 = ~n48293 & n48294;
  assign po932 = ~n48292 & ~n48295;
  assign n48297 = ~pi776 & ~po988;
  assign n48298 = pi1128 & po988;
  assign n48299 = ~pi966 & ~n48297;
  assign po933 = n48298 | ~n48299;
  assign n48301 = ~pi777 & ~po988;
  assign n48302 = pi1122 & po988;
  assign n48303 = ~pi966 & ~n48301;
  assign po934 = n48302 | ~n48303;
  assign n48305 = pi832 & pi956;
  assign n48306 = ~pi1046 & ~pi1083;
  assign n48307 = pi1085 & n48306;
  assign n48308 = n48305 & n48307;
  assign n48309 = ~pi968 & n48308;
  assign n48310 = pi778 & ~n48309;
  assign n48311 = pi1100 & n48309;
  assign po935 = n48310 | n48311;
  assign po936 = ~pi779 | n46497;
  assign po937 = ~pi780 | n46406;
  assign n48315 = pi781 & ~n48309;
  assign n48316 = pi1101 & n48309;
  assign po938 = n48315 | n48316;
  assign n48318 = ~n42180 & ~n46450;
  assign po939 = n46405 | ~n48318;
  assign n48320 = pi783 & ~n48309;
  assign n48321 = pi1109 & n48309;
  assign po940 = n48320 | n48321;
  assign n48323 = pi784 & ~n48309;
  assign n48324 = pi1110 & n48309;
  assign po941 = n48323 | n48324;
  assign n48326 = pi785 & ~n48309;
  assign n48327 = pi1102 & n48309;
  assign po942 = n48326 | n48327;
  assign n48329 = pi24 & ~pi954;
  assign n48330 = pi786 & pi954;
  assign po943 = ~n48329 & ~n48330;
  assign n48332 = pi787 & ~n48309;
  assign n48333 = pi1104 & n48309;
  assign po944 = n48332 | n48333;
  assign n48335 = pi788 & ~n48309;
  assign n48336 = pi1105 & n48309;
  assign po945 = n48335 | n48336;
  assign n48338 = pi789 & ~n48309;
  assign n48339 = pi1106 & n48309;
  assign po946 = n48338 | n48339;
  assign n48341 = pi790 & ~n48309;
  assign n48342 = pi1107 & n48309;
  assign po947 = n48341 | n48342;
  assign n48344 = pi791 & ~n48309;
  assign n48345 = pi1108 & n48309;
  assign po948 = n48344 | n48345;
  assign n48347 = pi792 & ~n48309;
  assign n48348 = pi1103 & n48309;
  assign po949 = n48347 | n48348;
  assign n48350 = pi968 & n48308;
  assign n48351 = pi794 & ~n48350;
  assign n48352 = pi1130 & n48350;
  assign po951 = n48351 | n48352;
  assign n48354 = pi795 & ~n48350;
  assign n48355 = pi1128 & n48350;
  assign po952 = n48354 | n48355;
  assign n48357 = pi266 & ~pi269;
  assign n48358 = pi278 & pi279;
  assign n48359 = ~pi280 & n48358;
  assign n48360 = n48357 & n48359;
  assign n48361 = ~pi281 & n48360;
  assign n48362 = n46689 & n48361;
  assign n48363 = pi264 & ~n48362;
  assign n48364 = ~pi264 & n48362;
  assign po953 = ~n48363 & ~n48364;
  assign n48366 = pi798 & ~n48350;
  assign n48367 = pi1124 & n48350;
  assign po955 = n48366 | n48367;
  assign n48369 = pi799 & ~n48350;
  assign n48370 = ~pi1107 & n48350;
  assign po956 = ~n48369 & ~n48370;
  assign n48372 = pi800 & ~n48350;
  assign n48373 = pi1125 & n48350;
  assign po957 = n48372 | n48373;
  assign n48375 = pi801 & ~n48350;
  assign n48376 = pi1126 & n48350;
  assign po958 = n48375 | n48376;
  assign n48378 = pi803 & ~n48350;
  assign n48379 = ~pi1106 & n48350;
  assign po960 = ~n48378 & ~n48379;
  assign n48381 = pi804 & ~n48350;
  assign n48382 = pi1109 & n48350;
  assign po961 = n48381 | n48382;
  assign n48384 = ~pi282 & n46687;
  assign n48385 = ~pi270 & n48384;
  assign n48386 = pi270 & ~n48384;
  assign po962 = ~n48385 & ~n48386;
  assign n48388 = pi807 & ~n48350;
  assign n48389 = pi1127 & n48350;
  assign po964 = n48388 | n48389;
  assign n48391 = pi808 & ~n48350;
  assign n48392 = pi1101 & n48350;
  assign po965 = n48391 | n48392;
  assign n48394 = pi809 & ~n48350;
  assign n48395 = ~pi1103 & n48350;
  assign po966 = ~n48394 & ~n48395;
  assign n48397 = pi810 & ~n48350;
  assign n48398 = pi1108 & n48350;
  assign po967 = n48397 | n48398;
  assign n48400 = pi811 & ~n48350;
  assign n48401 = pi1102 & n48350;
  assign po968 = n48400 | n48401;
  assign n48403 = pi812 & ~n48350;
  assign n48404 = ~pi1104 & n48350;
  assign po969 = ~n48403 & ~n48404;
  assign n48406 = pi813 & ~n48350;
  assign n48407 = pi1131 & n48350;
  assign po970 = n48406 | n48407;
  assign n48409 = pi814 & ~n48350;
  assign n48410 = ~pi1105 & n48350;
  assign po971 = ~n48409 & ~n48410;
  assign n48412 = pi815 & ~n48350;
  assign n48413 = pi1110 & n48350;
  assign po972 = n48412 | n48413;
  assign n48415 = pi816 & ~n48350;
  assign n48416 = pi1129 & n48350;
  assign po973 = n48415 | n48416;
  assign n48418 = pi269 & ~n46685;
  assign po974 = ~n46686 & ~n48418;
  assign n48420 = n8856 & n14132;
  assign po975 = n13986 | n48420;
  assign n48422 = pi265 & ~n46691;
  assign po976 = ~n46692 & ~n48422;
  assign n48424 = pi277 & ~n48385;
  assign po977 = ~n46690 & ~n48424;
  assign po979 = ~pi811 & ~pi893;
  assign n48427 = ~pi982 & ~n10054;
  assign n48428 = n7558 & n8856;
  assign n48429 = ~n48427 & ~n48428;
  assign po981 = n6265 & ~n48429;
  assign n48431 = pi123 & n3101;
  assign n48432 = pi1131 & ~n48431;
  assign n48433 = pi1127 & ~n48431;
  assign n48434 = ~n48432 & ~n48433;
  assign n48435 = ~pi825 & n48431;
  assign n48436 = n48434 & ~n48435;
  assign n48437 = pi1131 & n48433;
  assign n48438 = ~n48436 & ~n48437;
  assign n48439 = pi1124 & ~pi1130;
  assign n48440 = ~pi1124 & pi1130;
  assign n48441 = ~n48439 & ~n48440;
  assign n48442 = ~pi1128 & ~pi1129;
  assign n48443 = pi1128 & pi1129;
  assign n48444 = ~n48442 & ~n48443;
  assign n48445 = ~pi1125 & ~pi1126;
  assign n48446 = pi1125 & pi1126;
  assign n48447 = ~n48445 & ~n48446;
  assign n48448 = n48444 & ~n48447;
  assign n48449 = ~n48444 & n48447;
  assign n48450 = ~n48448 & ~n48449;
  assign n48451 = n48441 & n48450;
  assign n48452 = ~n48441 & ~n48450;
  assign n48453 = ~n48451 & ~n48452;
  assign n48454 = ~n48438 & ~n48453;
  assign n48455 = pi825 & n48431;
  assign n48456 = n48434 & ~n48455;
  assign n48457 = ~n48437 & n48453;
  assign n48458 = ~n48456 & n48457;
  assign po982 = ~n48454 & ~n48458;
  assign n48460 = pi1123 & ~n48431;
  assign n48461 = pi1122 & ~n48431;
  assign n48462 = ~n48460 & ~n48461;
  assign n48463 = ~pi826 & n48431;
  assign n48464 = n48462 & ~n48463;
  assign n48465 = pi1123 & n48461;
  assign n48466 = ~n48464 & ~n48465;
  assign n48467 = pi1118 & ~pi1119;
  assign n48468 = ~pi1118 & pi1119;
  assign n48469 = ~n48467 & ~n48468;
  assign n48470 = ~pi1120 & ~pi1121;
  assign n48471 = pi1120 & pi1121;
  assign n48472 = ~n48470 & ~n48471;
  assign n48473 = ~pi1116 & ~pi1117;
  assign n48474 = pi1116 & pi1117;
  assign n48475 = ~n48473 & ~n48474;
  assign n48476 = n48472 & ~n48475;
  assign n48477 = ~n48472 & n48475;
  assign n48478 = ~n48476 & ~n48477;
  assign n48479 = n48469 & n48478;
  assign n48480 = ~n48469 & ~n48478;
  assign n48481 = ~n48479 & ~n48480;
  assign n48482 = ~n48466 & ~n48481;
  assign n48483 = pi826 & n48431;
  assign n48484 = n48462 & ~n48483;
  assign n48485 = ~n48465 & n48481;
  assign n48486 = ~n48484 & n48485;
  assign po983 = ~n48482 & ~n48486;
  assign n48488 = pi1100 & ~n48431;
  assign n48489 = pi1107 & ~n48431;
  assign n48490 = ~n48488 & ~n48489;
  assign n48491 = ~pi827 & n48431;
  assign n48492 = n48490 & ~n48491;
  assign n48493 = pi1100 & n48489;
  assign n48494 = ~n48492 & ~n48493;
  assign n48495 = pi1103 & ~pi1105;
  assign n48496 = ~pi1103 & pi1105;
  assign n48497 = ~n48495 & ~n48496;
  assign n48498 = ~pi1101 & ~pi1102;
  assign n48499 = pi1101 & pi1102;
  assign n48500 = ~n48498 & ~n48499;
  assign n48501 = ~pi1104 & ~pi1106;
  assign n48502 = pi1104 & pi1106;
  assign n48503 = ~n48501 & ~n48502;
  assign n48504 = n48500 & ~n48503;
  assign n48505 = ~n48500 & n48503;
  assign n48506 = ~n48504 & ~n48505;
  assign n48507 = n48497 & n48506;
  assign n48508 = ~n48497 & ~n48506;
  assign n48509 = ~n48507 & ~n48508;
  assign n48510 = ~n48494 & ~n48509;
  assign n48511 = pi827 & n48431;
  assign n48512 = n48490 & ~n48511;
  assign n48513 = ~n48493 & n48509;
  assign n48514 = ~n48512 & n48513;
  assign po984 = ~n48510 & ~n48514;
  assign n48516 = pi1115 & ~n48431;
  assign n48517 = pi1114 & ~n48431;
  assign n48518 = ~n48516 & ~n48517;
  assign n48519 = ~pi828 & n48431;
  assign n48520 = n48518 & ~n48519;
  assign n48521 = pi1115 & n48517;
  assign n48522 = ~n48520 & ~n48521;
  assign n48523 = pi1110 & ~pi1111;
  assign n48524 = ~pi1110 & pi1111;
  assign n48525 = ~n48523 & ~n48524;
  assign n48526 = ~pi1112 & ~pi1113;
  assign n48527 = pi1112 & pi1113;
  assign n48528 = ~n48526 & ~n48527;
  assign n48529 = ~pi1108 & ~pi1109;
  assign n48530 = pi1108 & pi1109;
  assign n48531 = ~n48529 & ~n48530;
  assign n48532 = n48528 & ~n48531;
  assign n48533 = ~n48528 & n48531;
  assign n48534 = ~n48532 & ~n48533;
  assign n48535 = n48525 & n48534;
  assign n48536 = ~n48525 & ~n48534;
  assign n48537 = ~n48535 & ~n48536;
  assign n48538 = ~n48522 & ~n48537;
  assign n48539 = pi828 & n48431;
  assign n48540 = n48518 & ~n48539;
  assign n48541 = ~n48521 & n48537;
  assign n48542 = ~n48540 & n48541;
  assign po985 = ~n48538 & ~n48542;
  assign n48544 = n8856 & n10053;
  assign n48545 = pi951 & ~n48544;
  assign po986 = pi1092 & ~n48545;
  assign n48547 = pi281 & ~n48360;
  assign po987 = ~n48361 & ~n48547;
  assign n48549 = ~pi832 & pi1091;
  assign n48550 = pi1162 & n48549;
  assign po989 = n8860 & n48550;
  assign n48552 = pi833 & ~n2755;
  assign po990 = n16622 | n48552;
  assign po991 = pi946 & n2755;
  assign n48555 = pi282 & ~n46687;
  assign po992 = ~n48384 & ~n48555;
  assign n48557 = ~pi955 & pi1049;
  assign n48558 = pi837 & pi955;
  assign po993 = n48557 | n48558;
  assign n48560 = ~pi955 & pi1047;
  assign n48561 = pi838 & pi955;
  assign po994 = n48560 | n48561;
  assign n48563 = ~pi955 & pi1074;
  assign n48564 = pi839 & pi955;
  assign po995 = n48563 | n48564;
  assign n48566 = pi840 & ~n2755;
  assign n48567 = pi1196 & n2755;
  assign po996 = n48566 | n48567;
  assign po997 = ~pi33 & n8965;
  assign n48570 = ~pi955 & pi1035;
  assign n48571 = pi842 & pi955;
  assign po998 = n48570 | n48571;
  assign n48573 = ~pi955 & pi1079;
  assign n48574 = pi843 & pi955;
  assign po999 = n48573 | n48574;
  assign n48576 = ~pi955 & pi1078;
  assign n48577 = pi844 & pi955;
  assign po1000 = n48576 | n48577;
  assign n48579 = ~pi955 & pi1043;
  assign n48580 = pi845 & pi955;
  assign po1001 = n48579 | n48580;
  assign n48582 = pi846 & ~n42736;
  assign n48583 = pi1134 & n42736;
  assign po1002 = n48582 | n48583;
  assign n48585 = ~pi955 & pi1055;
  assign n48586 = pi847 & pi955;
  assign po1003 = n48585 | n48586;
  assign n48588 = ~pi955 & pi1039;
  assign n48589 = pi848 & pi955;
  assign po1004 = n48588 | n48589;
  assign n48591 = pi849 & ~n2755;
  assign n48592 = pi1198 & n2755;
  assign po1005 = n48591 | n48592;
  assign n48594 = ~pi955 & pi1048;
  assign n48595 = pi850 & pi955;
  assign po1006 = n48594 | n48595;
  assign n48597 = ~pi955 & pi1045;
  assign n48598 = pi851 & pi955;
  assign po1007 = n48597 | n48598;
  assign n48600 = ~pi955 & pi1062;
  assign n48601 = pi852 & pi955;
  assign po1008 = n48600 | n48601;
  assign n48603 = ~pi955 & pi1080;
  assign n48604 = pi853 & pi955;
  assign po1009 = n48603 | n48604;
  assign n48606 = ~pi955 & pi1051;
  assign n48607 = pi854 & pi955;
  assign po1010 = n48606 | n48607;
  assign n48609 = ~pi955 & pi1065;
  assign n48610 = pi855 & pi955;
  assign po1011 = n48609 | n48610;
  assign n48612 = ~pi955 & pi1067;
  assign n48613 = pi856 & pi955;
  assign po1012 = n48612 | n48613;
  assign n48615 = ~pi955 & pi1058;
  assign n48616 = pi857 & pi955;
  assign po1013 = n48615 | n48616;
  assign n48618 = ~pi955 & pi1087;
  assign n48619 = pi858 & pi955;
  assign po1014 = n48618 | n48619;
  assign n48621 = ~pi955 & pi1070;
  assign n48622 = pi859 & pi955;
  assign po1015 = n48621 | n48622;
  assign n48624 = ~pi955 & pi1076;
  assign n48625 = pi860 & pi955;
  assign po1016 = n48624 | n48625;
  assign n48627 = pi1093 & pi1141;
  assign n48628 = pi861 & ~pi1093;
  assign n48629 = ~n48627 & ~n48628;
  assign n48630 = ~pi228 & ~n48629;
  assign n48631 = ~pi123 & ~pi1141;
  assign n48632 = pi123 & ~pi861;
  assign n48633 = pi228 & ~n48631;
  assign n48634 = ~n48632 & n48633;
  assign po1017 = n48630 | n48634;
  assign n48636 = pi862 & ~n42736;
  assign n48637 = pi1139 & n42736;
  assign po1018 = n48636 | n48637;
  assign n48639 = pi863 & ~n2755;
  assign n48640 = pi1199 & n2755;
  assign po1019 = n48639 | n48640;
  assign n48642 = pi864 & ~n2755;
  assign n48643 = pi1197 & n2755;
  assign po1020 = n48642 | n48643;
  assign n48645 = ~pi955 & pi1040;
  assign n48646 = pi865 & pi955;
  assign po1021 = n48645 | n48646;
  assign n48648 = ~pi955 & pi1053;
  assign n48649 = pi866 & pi955;
  assign po1022 = n48648 | n48649;
  assign n48651 = ~pi955 & pi1057;
  assign n48652 = pi867 & pi955;
  assign po1023 = n48651 | n48652;
  assign n48654 = ~pi955 & pi1063;
  assign n48655 = pi868 & pi955;
  assign po1024 = n48654 | n48655;
  assign n48657 = pi1093 & pi1140;
  assign n48658 = pi869 & ~pi1093;
  assign n48659 = ~n48657 & ~n48658;
  assign n48660 = ~pi228 & ~n48659;
  assign n48661 = ~pi123 & ~pi1140;
  assign n48662 = pi123 & ~pi869;
  assign n48663 = pi228 & ~n48661;
  assign n48664 = ~n48662 & n48663;
  assign po1025 = n48660 | n48664;
  assign n48666 = ~pi955 & pi1069;
  assign n48667 = pi870 & pi955;
  assign po1026 = n48666 | n48667;
  assign n48669 = ~pi955 & pi1072;
  assign n48670 = pi871 & pi955;
  assign po1027 = n48669 | n48670;
  assign n48672 = ~pi955 & pi1084;
  assign n48673 = pi872 & pi955;
  assign po1028 = n48672 | n48673;
  assign n48675 = ~pi955 & pi1044;
  assign n48676 = pi873 & pi955;
  assign po1029 = n48675 | n48676;
  assign n48678 = ~pi955 & pi1036;
  assign n48679 = pi874 & pi955;
  assign po1030 = n48678 | n48679;
  assign n48681 = pi1093 & ~pi1136;
  assign n48682 = ~pi875 & ~pi1093;
  assign n48683 = ~n48681 & ~n48682;
  assign n48684 = ~pi228 & ~n48683;
  assign n48685 = ~pi123 & pi1136;
  assign n48686 = pi123 & pi875;
  assign n48687 = pi228 & ~n48685;
  assign n48688 = ~n48686 & n48687;
  assign po1031 = ~n48684 & ~n48688;
  assign n48690 = ~pi955 & pi1037;
  assign n48691 = pi876 & pi955;
  assign po1032 = n48690 | n48691;
  assign n48693 = pi1093 & pi1138;
  assign n48694 = pi877 & ~pi1093;
  assign n48695 = ~n48693 & ~n48694;
  assign n48696 = ~pi228 & ~n48695;
  assign n48697 = ~pi123 & ~pi1138;
  assign n48698 = pi123 & ~pi877;
  assign n48699 = pi228 & ~n48697;
  assign n48700 = ~n48698 & n48699;
  assign po1033 = n48696 | n48700;
  assign n48702 = pi1093 & pi1137;
  assign n48703 = pi878 & ~pi1093;
  assign n48704 = ~n48702 & ~n48703;
  assign n48705 = ~pi228 & ~n48704;
  assign n48706 = ~pi123 & ~pi1137;
  assign n48707 = pi123 & ~pi878;
  assign n48708 = pi228 & ~n48706;
  assign n48709 = ~n48707 & n48708;
  assign po1034 = n48705 | n48709;
  assign n48711 = pi1093 & pi1135;
  assign n48712 = pi879 & ~pi1093;
  assign n48713 = ~n48711 & ~n48712;
  assign n48714 = ~pi228 & ~n48713;
  assign n48715 = ~pi123 & ~pi1135;
  assign n48716 = pi123 & ~pi879;
  assign n48717 = pi228 & ~n48715;
  assign n48718 = ~n48716 & n48717;
  assign po1035 = n48714 | n48718;
  assign n48720 = ~pi955 & pi1081;
  assign n48721 = pi880 & pi955;
  assign po1036 = n48720 | n48721;
  assign n48723 = ~pi955 & pi1059;
  assign n48724 = pi881 & pi955;
  assign po1037 = n48723 | n48724;
  assign n48726 = ~pi883 & n48431;
  assign po1039 = n48489 | n48726;
  assign n48728 = pi1124 & ~n48431;
  assign n48729 = ~pi884 & n48431;
  assign po1040 = n48728 | n48729;
  assign n48731 = pi1125 & ~n48431;
  assign n48732 = ~pi885 & n48431;
  assign po1041 = n48731 | n48732;
  assign n48734 = pi1109 & ~n48431;
  assign n48735 = ~pi886 & n48431;
  assign po1042 = n48734 | n48735;
  assign n48737 = ~pi887 & n48431;
  assign po1043 = n48488 | n48737;
  assign n48739 = pi1120 & ~n48431;
  assign n48740 = ~pi888 & n48431;
  assign po1044 = n48739 | n48740;
  assign n48742 = pi1103 & ~n48431;
  assign n48743 = ~pi889 & n48431;
  assign po1045 = n48742 | n48743;
  assign n48745 = pi1126 & ~n48431;
  assign n48746 = ~pi890 & n48431;
  assign po1046 = n48745 | n48746;
  assign n48748 = pi1116 & ~n48431;
  assign n48749 = ~pi891 & n48431;
  assign po1047 = n48748 | n48749;
  assign n48751 = pi1101 & ~n48431;
  assign n48752 = ~pi892 & n48431;
  assign po1048 = n48751 | n48752;
  assign n48754 = pi1119 & ~n48431;
  assign n48755 = ~pi894 & n48431;
  assign po1050 = n48754 | n48755;
  assign n48757 = pi1113 & ~n48431;
  assign n48758 = ~pi895 & n48431;
  assign po1051 = n48757 | n48758;
  assign n48760 = pi1118 & ~n48431;
  assign n48761 = ~pi896 & n48431;
  assign po1052 = n48760 | n48761;
  assign n48763 = pi1129 & ~n48431;
  assign n48764 = ~pi898 & n48431;
  assign po1054 = n48763 | n48764;
  assign n48766 = ~pi899 & n48431;
  assign po1055 = n48516 | n48766;
  assign n48768 = pi1110 & ~n48431;
  assign n48769 = ~pi900 & n48431;
  assign po1056 = n48768 | n48769;
  assign n48771 = pi1111 & ~n48431;
  assign n48772 = ~pi902 & n48431;
  assign po1058 = n48771 | n48772;
  assign n48774 = pi1121 & ~n48431;
  assign n48775 = ~pi903 & n48431;
  assign po1059 = n48774 | n48775;
  assign n48777 = ~pi904 & n48431;
  assign po1060 = n48433 | n48777;
  assign n48779 = ~pi905 & n48431;
  assign po1061 = n48432 | n48779;
  assign n48781 = pi1128 & ~n48431;
  assign n48782 = ~pi906 & n48431;
  assign po1062 = n48781 | n48782;
  assign n48784 = ~pi624 & ~pi979;
  assign n48785 = ~pi598 & pi979;
  assign n48786 = pi782 & ~n48784;
  assign n48787 = ~n48785 & n48786;
  assign n48788 = ~pi604 & ~pi979;
  assign n48789 = pi615 & pi979;
  assign n48790 = ~n48788 & ~n48789;
  assign n48791 = pi782 & ~n48790;
  assign n48792 = ~pi782 & ~pi907;
  assign n48793 = ~n48787 & ~n48792;
  assign po1063 = ~n48791 & n48793;
  assign n48795 = ~pi908 & n48431;
  assign po1064 = n48461 | n48795;
  assign n48797 = pi1105 & ~n48431;
  assign n48798 = ~pi909 & n48431;
  assign po1065 = n48797 | n48798;
  assign n48800 = pi1117 & ~n48431;
  assign n48801 = ~pi910 & n48431;
  assign po1066 = n48800 | n48801;
  assign n48803 = pi1130 & ~n48431;
  assign n48804 = ~pi911 & n48431;
  assign po1067 = n48803 | n48804;
  assign n48806 = ~pi912 & n48431;
  assign po1068 = n48517 | n48806;
  assign n48808 = pi1106 & ~n48431;
  assign n48809 = ~pi913 & n48431;
  assign po1069 = n48808 | n48809;
  assign n48811 = pi280 & ~n46684;
  assign po1070 = ~n46685 & ~n48811;
  assign n48813 = pi1108 & ~n48431;
  assign n48814 = ~pi915 & n48431;
  assign po1071 = n48813 | n48814;
  assign n48816 = ~pi916 & n48431;
  assign po1072 = n48460 | n48816;
  assign n48818 = pi1112 & ~n48431;
  assign n48819 = ~pi917 & n48431;
  assign po1073 = n48818 | n48819;
  assign n48821 = pi1104 & ~n48431;
  assign n48822 = ~pi918 & n48431;
  assign po1074 = n48821 | n48822;
  assign n48824 = pi1102 & ~n48431;
  assign n48825 = ~pi919 & n48431;
  assign po1075 = n48824 | n48825;
  assign n48827 = pi1093 & pi1139;
  assign n48828 = pi920 & ~pi1093;
  assign po1076 = n48827 | n48828;
  assign n48830 = pi921 & ~pi1093;
  assign po1077 = n48657 | n48830;
  assign n48832 = ~pi922 & ~pi1093;
  assign n48833 = pi1093 & ~pi1152;
  assign po1078 = ~n48832 & ~n48833;
  assign n48835 = ~pi923 & ~pi1093;
  assign n48836 = pi1093 & ~pi1154;
  assign po1079 = ~n48835 & ~n48836;
  assign n48838 = ~pi300 & pi301;
  assign n48839 = pi311 & ~pi312;
  assign po1080 = n48838 & n48839;
  assign n48841 = ~pi925 & ~pi1093;
  assign n48842 = pi1093 & ~pi1155;
  assign po1081 = ~n48841 & ~n48842;
  assign n48844 = ~pi926 & ~pi1093;
  assign n48845 = pi1093 & ~pi1157;
  assign po1082 = ~n48844 & ~n48845;
  assign n48847 = ~pi927 & ~pi1093;
  assign n48848 = pi1093 & ~pi1145;
  assign po1083 = ~n48847 & ~n48848;
  assign n48850 = ~pi928 & ~pi1093;
  assign po1084 = ~n48681 & ~n48850;
  assign n48852 = ~pi929 & ~pi1093;
  assign n48853 = pi1093 & ~pi1144;
  assign po1085 = ~n48852 & ~n48853;
  assign n48855 = ~pi930 & ~pi1093;
  assign n48856 = pi1093 & ~pi1134;
  assign po1086 = ~n48855 & ~n48856;
  assign n48858 = ~pi931 & ~pi1093;
  assign n48859 = pi1093 & ~pi1150;
  assign po1087 = ~n48858 & ~n48859;
  assign n48861 = pi932 & ~pi1093;
  assign po1088 = n42725 | n48861;
  assign n48863 = pi933 & ~pi1093;
  assign po1089 = n48702 | n48863;
  assign n48865 = ~pi934 & ~pi1093;
  assign n48866 = pi1093 & ~pi1147;
  assign po1090 = ~n48865 & ~n48866;
  assign n48868 = pi935 & ~pi1093;
  assign po1091 = n48627 | n48868;
  assign n48870 = ~pi936 & ~pi1093;
  assign n48871 = pi1093 & ~pi1149;
  assign po1092 = ~n48870 & ~n48871;
  assign n48873 = ~pi937 & ~pi1093;
  assign n48874 = pi1093 & ~pi1148;
  assign po1093 = ~n48873 & ~n48874;
  assign n48876 = pi938 & ~pi1093;
  assign po1094 = n48711 | n48876;
  assign n48878 = ~pi939 & ~pi1093;
  assign n48879 = pi1093 & ~pi1146;
  assign po1095 = ~n48878 & ~n48879;
  assign n48881 = pi940 & ~pi1093;
  assign po1096 = n48693 | n48881;
  assign n48883 = ~pi941 & ~pi1093;
  assign n48884 = pi1093 & ~pi1153;
  assign po1097 = ~n48883 & ~n48884;
  assign n48886 = ~pi942 & ~pi1093;
  assign n48887 = pi1093 & ~pi1156;
  assign po1098 = ~n48886 & ~n48887;
  assign n48889 = ~pi943 & ~pi1093;
  assign n48890 = pi1093 & ~pi1151;
  assign po1099 = ~n48889 & ~n48890;
  assign n48892 = pi1093 & pi1143;
  assign n48893 = pi944 & ~pi1093;
  assign po1100 = n48892 | n48893;
  assign po1102 = pi230 & n2755;
  assign n48896 = ~pi782 & pi947;
  assign po1103 = n48787 | n48896;
  assign n48898 = ~pi266 & ~pi992;
  assign po1104 = ~n46684 & ~n48898;
  assign n48900 = ~pi313 & ~pi954;
  assign n48901 = pi949 & pi954;
  assign po1105 = n48900 | n48901;
  assign po1107 = ~n7558 & n14216;
  assign n48904 = pi957 & pi1092;
  assign po1112 = pi31 | n48904;
  assign po1115 = ~pi782 & pi960;
  assign po1116 = ~pi230 & pi961;
  assign po1118 = ~pi782 & pi963;
  assign po1122 = ~pi230 & pi967;
  assign po1124 = ~pi230 & pi969;
  assign po1125 = ~pi782 & pi970;
  assign po1126 = ~pi230 & pi971;
  assign po1127 = ~pi782 & pi972;
  assign po1128 = ~pi230 & pi974;
  assign po1129 = ~pi782 & pi975;
  assign po1131 = ~pi230 & pi977;
  assign po1132 = ~pi782 & pi978;
  assign po1133 = pi598 | ~pi615;
  assign po1135 = pi824 & pi1092;
  assign po1137 = pi604 | pi624;
  assign po166 = 1'b1;
  assign po170 = ~pi1090;
  assign po1110 = ~pi954;
  assign po1130 = ~pi278;
  assign po1146 = ~pi915;
  assign po1147 = ~pi825;
  assign po1148 = ~pi826;
  assign po1149 = ~pi913;
  assign po1150 = ~pi894;
  assign po1151 = ~pi905;
  assign po1153 = ~pi890;
  assign po1155 = ~pi906;
  assign po1156 = ~pi896;
  assign po1157 = ~pi909;
  assign po1158 = ~pi911;
  assign po1159 = ~pi908;
  assign po1160 = ~pi891;
  assign po1161 = ~pi902;
  assign po1162 = ~pi903;
  assign po1163 = ~pi883;
  assign po1164 = ~pi888;
  assign po1165 = ~pi919;
  assign po1166 = ~pi886;
  assign po1167 = ~pi912;
  assign po1168 = ~pi895;
  assign po1169 = ~pi916;
  assign po1170 = ~pi889;
  assign po1171 = ~pi900;
  assign po1172 = ~pi885;
  assign po1173 = ~pi904;
  assign po1174 = ~pi899;
  assign po1175 = ~pi918;
  assign po1176 = ~pi898;
  assign po1177 = ~pi917;
  assign po1178 = ~pi827;
  assign po1179 = ~pi887;
  assign po1180 = ~pi884;
  assign po1181 = ~pi910;
  assign po1182 = ~pi828;
  assign po1183 = ~pi892;
  assign po0 = pi668;
  assign po1 = pi672;
  assign po2 = pi664;
  assign po3 = pi667;
  assign po4 = pi676;
  assign po5 = pi673;
  assign po6 = pi675;
  assign po7 = pi666;
  assign po8 = pi679;
  assign po9 = pi674;
  assign po10 = pi663;
  assign po11 = pi670;
  assign po12 = pi677;
  assign po13 = pi682;
  assign po14 = pi671;
  assign po15 = pi678;
  assign po16 = pi718;
  assign po17 = pi707;
  assign po18 = pi708;
  assign po19 = pi713;
  assign po20 = pi711;
  assign po21 = pi716;
  assign po22 = pi733;
  assign po23 = pi712;
  assign po24 = pi689;
  assign po25 = pi717;
  assign po26 = pi692;
  assign po27 = pi719;
  assign po28 = pi722;
  assign po29 = pi714;
  assign po30 = pi720;
  assign po31 = pi685;
  assign po32 = pi837;
  assign po33 = pi850;
  assign po34 = pi872;
  assign po35 = pi871;
  assign po36 = pi881;
  assign po37 = pi866;
  assign po38 = pi876;
  assign po39 = pi873;
  assign po40 = pi874;
  assign po41 = pi859;
  assign po42 = pi855;
  assign po43 = pi852;
  assign po44 = pi870;
  assign po45 = pi848;
  assign po46 = pi865;
  assign po47 = pi856;
  assign po48 = pi853;
  assign po49 = pi847;
  assign po50 = pi857;
  assign po51 = pi854;
  assign po52 = pi858;
  assign po53 = pi845;
  assign po54 = pi838;
  assign po55 = pi842;
  assign po56 = pi843;
  assign po57 = pi839;
  assign po58 = pi844;
  assign po59 = pi868;
  assign po60 = pi851;
  assign po61 = pi867;
  assign po62 = pi880;
  assign po63 = pi860;
  assign po64 = pi1030;
  assign po65 = pi1034;
  assign po66 = pi1015;
  assign po67 = pi1020;
  assign po68 = pi1025;
  assign po69 = pi1005;
  assign po70 = pi996;
  assign po71 = pi1012;
  assign po72 = pi993;
  assign po73 = pi1016;
  assign po74 = pi1021;
  assign po75 = pi1010;
  assign po76 = pi1027;
  assign po77 = pi1018;
  assign po78 = pi1017;
  assign po79 = pi1024;
  assign po80 = pi1009;
  assign po81 = pi1032;
  assign po82 = pi1003;
  assign po83 = pi997;
  assign po84 = pi1013;
  assign po85 = pi1011;
  assign po86 = pi1008;
  assign po87 = pi1019;
  assign po88 = pi1031;
  assign po89 = pi1022;
  assign po90 = pi1000;
  assign po91 = pi1023;
  assign po92 = pi1002;
  assign po93 = pi1026;
  assign po94 = pi1006;
  assign po95 = pi998;
  assign po96 = pi31;
  assign po97 = pi80;
  assign po98 = pi893;
  assign po99 = pi467;
  assign po100 = pi78;
  assign po101 = pi112;
  assign po102 = pi13;
  assign po103 = pi25;
  assign po104 = pi226;
  assign po105 = pi127;
  assign po106 = pi822;
  assign po107 = pi808;
  assign po108 = pi227;
  assign po109 = pi477;
  assign po110 = pi834;
  assign po111 = pi229;
  assign po112 = pi12;
  assign po113 = pi11;
  assign po114 = pi10;
  assign po115 = pi9;
  assign po116 = pi8;
  assign po117 = pi7;
  assign po118 = pi6;
  assign po119 = pi5;
  assign po120 = pi4;
  assign po121 = pi3;
  assign po122 = pi0;
  assign po123 = pi2;
  assign po124 = pi1;
  assign po125 = pi310;
  assign po126 = pi302;
  assign po127 = pi475;
  assign po128 = pi474;
  assign po129 = pi466;
  assign po130 = pi473;
  assign po131 = pi471;
  assign po132 = pi472;
  assign po133 = pi470;
  assign po134 = pi469;
  assign po135 = pi465;
  assign po136 = pi1028;
  assign po137 = pi1033;
  assign po138 = pi995;
  assign po139 = pi994;
  assign po140 = pi28;
  assign po141 = pi27;
  assign po142 = pi26;
  assign po143 = pi29;
  assign po144 = pi15;
  assign po145 = pi14;
  assign po146 = pi21;
  assign po147 = pi20;
  assign po148 = pi19;
  assign po149 = pi18;
  assign po150 = pi17;
  assign po151 = pi16;
  assign po152 = pi1096;
  assign po168 = pi228;
  assign po169 = pi22;
  assign po179 = pi1089;
  assign po180 = pi23;
  assign po181 = po167;
  assign po188 = pi37;
  assign po263 = pi117;
  assign po285 = pi131;
  assign po386 = pi232;
  assign po388 = pi236;
  assign po636 = pi583;
  assign po1053 = pi67;
  assign po1108 = pi1134;
  assign po1109 = pi964;
  assign po1111 = pi965;
  assign po1113 = pi991;
  assign po1114 = pi985;
  assign po1117 = pi1014;
  assign po1119 = pi1029;
  assign po1120 = pi1004;
  assign po1121 = pi1007;
  assign po1123 = pi1135;
  assign po1134 = pi1064;
  assign po1136 = pi299;
  assign po1138 = pi1075;
  assign po1139 = pi1052;
  assign po1140 = pi771;
  assign po1141 = pi765;
  assign po1142 = pi605;
  assign po1143 = pi601;
  assign po1144 = pi278;
  assign po1145 = pi279;
  assign po1152 = pi1095;
  assign po1154 = pi1094;
  assign po1184 = pi1187;
  assign po1185 = pi1172;
  assign po1186 = pi1170;
  assign po1187 = pi1138;
  assign po1188 = pi1177;
  assign po1189 = pi1178;
  assign po1190 = pi863;
  assign po1191 = pi1203;
  assign po1192 = pi1185;
  assign po1193 = pi1171;
  assign po1194 = pi1192;
  assign po1195 = pi1137;
  assign po1196 = pi1186;
  assign po1197 = pi1165;
  assign po1198 = pi1164;
  assign po1199 = pi1098;
  assign po1200 = pi1183;
  assign po1201 = pi230;
  assign po1202 = pi1169;
  assign po1203 = pi1136;
  assign po1204 = pi1181;
  assign po1205 = pi849;
  assign po1206 = pi1193;
  assign po1207 = pi1182;
  assign po1208 = pi1168;
  assign po1209 = pi1175;
  assign po1210 = pi1191;
  assign po1211 = pi1099;
  assign po1212 = pi1174;
  assign po1213 = pi1179;
  assign po1214 = pi1202;
  assign po1215 = pi1176;
  assign po1216 = pi1173;
  assign po1217 = pi1201;
  assign po1218 = pi1167;
  assign po1219 = pi840;
  assign po1220 = pi1189;
  assign po1221 = pi1195;
  assign po1222 = pi864;
  assign po1223 = pi1190;
  assign po1224 = pi1188;
  assign po1225 = pi1180;
  assign po1226 = pi1194;
  assign po1227 = pi1097;
  assign po1228 = pi1166;
  assign po1229 = pi1200;
  assign po1230 = pi1184;
endmodule
