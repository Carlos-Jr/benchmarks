module alu4_cl ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13,
    po0, po1, po2, po3, po4, po5, po6, po7  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13;
  output po0, po1, po2, po3, po4, po5, po6, po7;
  wire n23, n24, n25, n26, n27, n28, n29,
    n30, n31, n32, n33, n34, n35, n36, n37,
    n38, n39, n40, n41, n42, n43, n44, n45,
    n46, n47, n48, n49, n50, n51, n52, n53,
    n54, n55, n56, n57, n58, n59, n60, n61,
    n62, n63, n64, n65, n66, n67, n68, n69,
    n70, n71, n72, n73, n74, n75, n76, n77,
    n78, n79, n80, n81, n82, n83, n84, n85,
    n86, n87, n88, n89, n90, n91, n92, n93,
    n94, n95, n96, n97, n98, n99, n100,
    n101, n102, n103, n104, n105, n106, n107,
    n108, n109, n110, n111, n112, n113, n114,
    n115, n116, n117, n118, n119, n120, n121,
    n122, n123, n124, n125, n126, n127, n128,
    n129, n130, n131, n132, n133, n134, n135,
    n136, n137, n138, n139, n140, n141, n142,
    n143, n144, n145, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156,
    n157, n158, n159, n160, n161, n162, n163,
    n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177,
    n178, n179, n180, n181, n182, n183, n184,
    n185, n186, n187, n188, n190, n191, n192,
    n193, n194, n195, n196, n197, n198, n199,
    n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213,
    n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227,
    n228, n229, n230, n231, n232, n233, n234,
    n235, n236, n237, n238, n239, n240, n241,
    n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403,
    n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416, n417,
    n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438,
    n439, n440, n441, n442, n443, n444, n445,
    n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n488,
    n489, n490, n491, n492, n493, n494, n495,
    n496, n497, n498, n499, n500, n502, n503,
    n504, n505, n506, n507, n508, n509, n510,
    n511, n512, n513, n514, n515, n516, n517,
    n518, n519, n520, n521, n522, n523, n524,
    n525, n526, n527, n528, n529, n530, n531,
    n532, n533, n534, n535, n536, n538, n539,
    n540, n541, n542, n543, n544, n545, n546,
    n547, n548, n549, n550, n551, n552, n553,
    n554, n555, n556, n557, n558, n559, n560,
    n561, n562, n563, n564, n565, n566, n567,
    n568, n569, n570, n571, n572, n573, n574,
    n575, n576, n577, n578, n579, n580, n581,
    n582, n583, n584, n585, n586, n587, n588,
    n589, n590, n591, n592, n593, n594, n595,
    n596, n597, n598, n599, n600, n601, n602,
    n603, n604, n605, n606, n607, n608, n609,
    n610, n611, n612, n613, n614, n615, n616,
    n617, n618, n619, n620, n621, n622, n623,
    n624, n625, n626, n627, n628, n629, n630,
    n631, n632, n633, n634, n635, n636, n637,
    n638, n639, n640, n641, n642, n643, n644,
    n645, n647, n648, n649, n650, n651, n652,
    n653, n654, n655, n656, n657, n658, n659,
    n660, n661, n662, n663, n664, n665, n666,
    n667, n668, n669, n670, n671, n672, n674,
    n675, n676, n677, n678, n679;
  assign n23 = ~pi08 & pi09;
  assign n24 = pi00 & ~pi04;
  assign n25 = ~pi00 & pi04;
  assign n26 = pi10 & ~pi11;
  assign n27 = n25 & n26;
  assign n28 = ~n24 & ~n27;
  assign n29 = pi13 & ~n28;
  assign n30 = n23 & n29;
  assign n31 = ~pi00 & ~pi04;
  assign n32 = pi08 & ~pi09;
  assign n33 = pi10 & pi13;
  assign n34 = ~pi10 & ~pi11;
  assign n35 = ~pi13 & n34;
  assign n36 = ~n33 & ~n35;
  assign n37 = n32 & ~n36;
  assign n38 = ~n31 & n37;
  assign n39 = pi08 & pi09;
  assign n40 = ~pi10 & n39;
  assign n41 = pi11 & n40;
  assign n42 = ~pi08 & ~pi10;
  assign n43 = ~pi09 & pi11;
  assign n44 = n42 & n43;
  assign n45 = ~n41 & ~n44;
  assign n46 = pi13 & ~n45;
  assign n47 = ~pi08 & n26;
  assign n48 = ~pi09 & n47;
  assign n49 = ~n46 & ~n48;
  assign n50 = pi00 & pi04;
  assign n51 = ~n49 & n50;
  assign n52 = ~n38 & ~n51;
  assign n53 = pi09 & pi11;
  assign n54 = ~pi10 & ~n53;
  assign n55 = ~pi13 & n54;
  assign n56 = ~pi08 & n55;
  assign n57 = ~pi00 & n56;
  assign n58 = n26 & n39;
  assign n59 = n23 & ~n26;
  assign n60 = pi13 & n59;
  assign n61 = pi08 & pi10;
  assign n62 = ~pi13 & n61;
  assign n63 = n43 & n62;
  assign n64 = ~n60 & ~n63;
  assign n65 = ~n58 & n64;
  assign n66 = ~pi04 & ~n65;
  assign n67 = ~n57 & ~n66;
  assign n68 = n52 & n67;
  assign n69 = ~n30 & n68;
  assign n70 = ~pi00 & n69;
  assign n71 = ~pi08 & pi11;
  assign n72 = pi09 & n71;
  assign n73 = pi13 & n72;
  assign n74 = ~n70 & n73;
  assign n75 = pi13 & n26;
  assign n76 = ~pi08 & ~pi09;
  assign n77 = n69 & n76;
  assign n78 = n32 & n50;
  assign n79 = pi00 & ~n69;
  assign n80 = n39 & n79;
  assign n81 = ~n78 & ~n80;
  assign n82 = ~n77 & n81;
  assign n83 = n75 & ~n82;
  assign n84 = ~n74 & ~n83;
  assign n85 = ~pi10 & ~n76;
  assign n86 = ~pi00 & ~n85;
  assign n87 = n48 & n86;
  assign n88 = pi09 & n42;
  assign n89 = ~pi10 & n73;
  assign n90 = n50 & n89;
  assign n91 = ~pi09 & n26;
  assign n92 = pi13 & n91;
  assign n93 = pi08 & n92;
  assign n94 = n84 & n93;
  assign n95 = ~n90 & ~n94;
  assign n96 = n88 & ~n95;
  assign n97 = pi11 & n88;
  assign n98 = ~n96 & n97;
  assign n99 = ~n87 & ~n98;
  assign n100 = ~n84 & ~n99;
  assign n101 = pi09 & ~n69;
  assign n102 = ~pi00 & ~n101;
  assign n103 = ~pi11 & ~n102;
  assign n104 = pi00 & ~pi09;
  assign n105 = n69 & n104;
  assign n106 = ~n103 & ~n105;
  assign n107 = n42 & ~n106;
  assign n108 = pi08 & n95;
  assign n109 = n91 & n108;
  assign n110 = pi11 & n86;
  assign n111 = ~n109 & ~n110;
  assign n112 = ~n69 & ~n111;
  assign n113 = pi09 & n47;
  assign n114 = ~n41 & ~n113;
  assign n115 = pi00 & pi11;
  assign n116 = ~n39 & n115;
  assign n117 = ~pi09 & ~pi11;
  assign n118 = pi08 & ~n95;
  assign n119 = n117 & n118;
  assign n120 = ~n116 & ~n119;
  assign n121 = pi10 & ~n120;
  assign n122 = n114 & ~n121;
  assign n123 = n69 & ~n122;
  assign n124 = pi08 & ~pi10;
  assign n125 = pi04 & n124;
  assign n126 = pi00 & ~pi08;
  assign n127 = n84 & n126;
  assign n128 = ~n125 & ~n127;
  assign n129 = n117 & ~n128;
  assign n130 = pi11 & n96;
  assign n131 = ~n58 & ~n130;
  assign n132 = n84 & ~n131;
  assign n133 = pi09 & n61;
  assign n134 = n110 & n133;
  assign n135 = ~n132 & ~n134;
  assign n136 = ~n129 & n135;
  assign n137 = ~n123 & n136;
  assign n138 = ~n112 & n137;
  assign n139 = ~n107 & n138;
  assign n140 = ~n100 & n139;
  assign n141 = ~pi09 & n124;
  assign n142 = ~n31 & ~n50;
  assign n143 = n141 & n142;
  assign n144 = n140 & ~n143;
  assign n145 = pi13 & ~n144;
  assign n146 = ~pi12 & n145;
  assign n147 = pi12 & ~n145;
  assign n148 = ~n146 & ~n147;
  assign n149 = pi13 & n148;
  assign n150 = n34 & n39;
  assign n151 = pi13 & n150;
  assign n152 = ~pi09 & pi10;
  assign n153 = n71 & n152;
  assign n154 = ~pi13 & n153;
  assign n155 = ~n151 & ~n154;
  assign n156 = pi04 & n42;
  assign n157 = ~n39 & ~n85;
  assign n158 = ~n26 & n157;
  assign n159 = ~pi09 & n158;
  assign n160 = ~n156 & ~n159;
  assign n161 = ~n69 & ~n160;
  assign n162 = pi04 & n71;
  assign n163 = n31 & n47;
  assign n164 = ~n162 & ~n163;
  assign n165 = ~pi08 & pi10;
  assign n166 = ~pi11 & ~n165;
  assign n167 = n50 & ~n166;
  assign n168 = n61 & n79;
  assign n169 = ~n167 & ~n168;
  assign n170 = n164 & n169;
  assign n171 = pi09 & ~n170;
  assign n172 = pi08 & n34;
  assign n173 = ~n165 & ~n172;
  assign n174 = n69 & ~n173;
  assign n175 = pi08 & n26;
  assign n176 = ~pi04 & n175;
  assign n177 = ~n174 & ~n176;
  assign n178 = pi11 & n124;
  assign n179 = ~n115 & ~n178;
  assign n180 = n142 & ~n179;
  assign n181 = n177 & ~n180;
  assign n182 = ~pi09 & ~n181;
  assign n183 = ~n85 & n115;
  assign n184 = ~n182 & ~n183;
  assign n185 = ~n171 & n184;
  assign n186 = ~n161 & n185;
  assign n187 = ~pi13 & ~n186;
  assign n188 = n155 & ~n187;
  assign po0 = n149 | ~n188;
  assign n190 = pi11 & ~n85;
  assign n191 = pi01 & pi05;
  assign n192 = n49 & ~n92;
  assign n193 = ~pi08 & pi13;
  assign n194 = n27 & n193;
  assign n195 = n192 & ~n194;
  assign n196 = n191 & ~n195;
  assign n197 = n115 & n152;
  assign n198 = ~pi01 & ~pi05;
  assign n199 = n25 & n198;
  assign n200 = pi01 & ~pi05;
  assign n201 = ~pi01 & pi05;
  assign n202 = n25 & ~n200;
  assign n203 = ~n201 & ~n202;
  assign n204 = n26 & ~n203;
  assign n205 = ~n200 & ~n204;
  assign n206 = ~n25 & ~n205;
  assign n207 = ~n199 & ~n206;
  assign n208 = pi09 & ~n207;
  assign n209 = ~n197 & ~n208;
  assign n210 = ~pi08 & ~n209;
  assign n211 = pi13 & n210;
  assign n212 = n37 & ~n198;
  assign n213 = ~pi01 & n56;
  assign n214 = ~pi05 & ~n65;
  assign n215 = ~n213 & ~n214;
  assign n216 = ~n212 & n215;
  assign n217 = ~n211 & n216;
  assign n218 = ~n196 & n217;
  assign n219 = n133 & ~n218;
  assign n220 = ~n190 & ~n219;
  assign n221 = pi01 & ~n220;
  assign n222 = pi05 & n42;
  assign n223 = ~n159 & ~n222;
  assign n224 = ~n218 & ~n223;
  assign n225 = pi05 & n71;
  assign n226 = ~n166 & n191;
  assign n227 = n47 & n198;
  assign n228 = ~n226 & ~n227;
  assign n229 = ~n225 & n228;
  assign n230 = pi09 & ~n229;
  assign n231 = pi11 & n200;
  assign n232 = n178 & n201;
  assign n233 = ~n231 & ~n232;
  assign n234 = ~n173 & n218;
  assign n235 = ~pi05 & n175;
  assign n236 = ~n234 & ~n235;
  assign n237 = n233 & n236;
  assign n238 = ~pi09 & ~n237;
  assign n239 = ~n230 & ~n238;
  assign n240 = ~n224 & n239;
  assign n241 = ~n221 & n240;
  assign n242 = ~pi13 & ~n241;
  assign n243 = n155 & ~n242;
  assign n244 = pi11 & n157;
  assign n245 = n79 & ~n218;
  assign n246 = ~n79 & n218;
  assign n247 = ~n245 & ~n246;
  assign n248 = n244 & n247;
  assign n249 = ~pi01 & n218;
  assign n250 = n73 & ~n249;
  assign n251 = n76 & n218;
  assign n252 = pi09 & ~n218;
  assign n253 = pi05 & ~pi09;
  assign n254 = ~n252 & ~n253;
  assign n255 = pi08 & ~n254;
  assign n256 = pi01 & n255;
  assign n257 = ~n251 & ~n256;
  assign n258 = n75 & ~n257;
  assign n259 = ~n250 & ~n258;
  assign n260 = pi00 & ~n84;
  assign n261 = n259 & n260;
  assign n262 = ~n259 & ~n260;
  assign n263 = ~n261 & ~n262;
  assign n264 = n48 & ~n263;
  assign n265 = ~n248 & ~n264;
  assign n266 = ~pi01 & ~n265;
  assign n267 = ~n69 & ~n95;
  assign n268 = n89 & n191;
  assign n269 = n93 & n259;
  assign n270 = ~n268 & ~n269;
  assign n271 = n267 & ~n270;
  assign n272 = ~n267 & n270;
  assign n273 = ~n271 & ~n272;
  assign n274 = ~n218 & ~n273;
  assign n275 = n218 & n273;
  assign n276 = ~n274 & ~n275;
  assign n277 = n61 & ~n276;
  assign n278 = pi05 & n124;
  assign n279 = ~pi08 & n263;
  assign n280 = pi01 & n279;
  assign n281 = ~n278 & ~n280;
  assign n282 = ~n277 & n281;
  assign n283 = n117 & ~n282;
  assign n284 = ~pi00 & ~pi01;
  assign n285 = n133 & n284;
  assign n286 = n50 & n198;
  assign n287 = n141 & n286;
  assign n288 = ~n285 & ~n287;
  assign n289 = pi11 & ~n288;
  assign n290 = ~n84 & ~n95;
  assign n291 = ~n270 & n290;
  assign n292 = n270 & ~n290;
  assign n293 = ~n291 & ~n292;
  assign n294 = ~n259 & ~n293;
  assign n295 = n259 & n293;
  assign n296 = ~n294 & ~n295;
  assign n297 = n97 & ~n296;
  assign n298 = n158 & ~n247;
  assign n299 = n34 & ~n39;
  assign n300 = n115 & n133;
  assign n301 = ~pi05 & ~n50;
  assign n302 = n141 & n301;
  assign n303 = ~n300 & ~n302;
  assign n304 = ~n299 & n303;
  assign n305 = ~n298 & n304;
  assign n306 = pi01 & ~n305;
  assign n307 = n84 & n259;
  assign n308 = ~n84 & ~n259;
  assign n309 = ~n307 & ~n308;
  assign n310 = n133 & ~n309;
  assign n311 = n88 & ~n218;
  assign n312 = ~n310 & ~n311;
  assign n313 = ~pi11 & ~n312;
  assign n314 = ~n50 & n201;
  assign n315 = n50 & n191;
  assign n316 = ~n314 & ~n315;
  assign n317 = n141 & ~n316;
  assign n318 = n69 & n218;
  assign n319 = ~n114 & n318;
  assign n320 = ~pi11 & n88;
  assign n321 = n114 & ~n320;
  assign n322 = ~n69 & ~n321;
  assign n323 = ~n218 & n322;
  assign n324 = ~n319 & ~n323;
  assign n325 = ~n317 & n324;
  assign n326 = ~n313 & n325;
  assign n327 = ~n306 & n326;
  assign n328 = ~n297 & n327;
  assign n329 = ~n289 & n328;
  assign n330 = ~n283 & n329;
  assign n331 = ~n266 & n330;
  assign n332 = pi13 & ~n331;
  assign n333 = n146 & n332;
  assign n334 = ~n146 & ~n332;
  assign n335 = ~n333 & ~n334;
  assign po1 = ~n243 | n335;
  assign n337 = pi02 & pi11;
  assign n338 = ~pi06 & ~pi09;
  assign n339 = n85 & ~n338;
  assign n340 = n337 & ~n339;
  assign n341 = pi06 & n204;
  assign n342 = pi09 & n203;
  assign n343 = ~pi06 & n342;
  assign n344 = ~n341 & ~n343;
  assign n345 = pi02 & ~n344;
  assign n346 = ~pi06 & ~n203;
  assign n347 = n26 & n203;
  assign n348 = pi06 & n347;
  assign n349 = ~n346 & ~n348;
  assign n350 = pi09 & ~n349;
  assign n351 = ~pi02 & n350;
  assign n352 = pi01 & pi11;
  assign n353 = n152 & n352;
  assign n354 = ~n351 & ~n353;
  assign n355 = ~n345 & n354;
  assign n356 = ~pi08 & ~n355;
  assign n357 = pi13 & n356;
  assign n358 = pi02 & pi06;
  assign n359 = ~n192 & n358;
  assign n360 = ~pi06 & ~n65;
  assign n361 = ~n359 & ~n360;
  assign n362 = ~pi02 & n56;
  assign n363 = ~pi02 & ~pi06;
  assign n364 = n37 & ~n363;
  assign n365 = ~n362 & ~n364;
  assign n366 = n361 & n365;
  assign n367 = ~n357 & n366;
  assign n368 = pi06 & n42;
  assign n369 = pi02 & n133;
  assign n370 = ~n159 & ~n369;
  assign n371 = ~n368 & n370;
  assign n372 = ~n367 & ~n371;
  assign n373 = ~pi02 & n178;
  assign n374 = ~pi09 & n373;
  assign n375 = ~n72 & ~n374;
  assign n376 = pi06 & ~n375;
  assign n377 = ~n358 & ~n363;
  assign n378 = ~n47 & ~n337;
  assign n379 = ~n377 & ~n378;
  assign n380 = pi09 & n379;
  assign n381 = ~n173 & n367;
  assign n382 = ~pi06 & n175;
  assign n383 = ~n381 & ~n382;
  assign n384 = ~pi09 & ~n383;
  assign n385 = ~n380 & ~n384;
  assign n386 = ~n376 & n385;
  assign n387 = ~n372 & n386;
  assign n388 = ~n340 & n387;
  assign n389 = ~pi13 & ~n388;
  assign n390 = n155 & ~n389;
  assign n391 = pi01 & n247;
  assign n392 = ~n245 & ~n391;
  assign n393 = n158 & n392;
  assign n394 = pi02 & n393;
  assign n395 = n244 & ~n392;
  assign n396 = ~pi02 & n395;
  assign n397 = ~n394 & ~n396;
  assign n398 = n367 & ~n397;
  assign n399 = n50 & ~n198;
  assign n400 = ~n191 & ~n399;
  assign n401 = pi11 & n363;
  assign n402 = ~n358 & ~n401;
  assign n403 = ~n400 & ~n402;
  assign n404 = n377 & n400;
  assign n405 = ~n403 & ~n404;
  assign n406 = n141 & ~n405;
  assign n407 = n244 & n392;
  assign n408 = ~n367 & n407;
  assign n409 = ~pi02 & n367;
  assign n410 = n73 & ~n409;
  assign n411 = n76 & n367;
  assign n412 = pi09 & ~n367;
  assign n413 = pi06 & ~pi09;
  assign n414 = ~n412 & ~n413;
  assign n415 = pi08 & ~n414;
  assign n416 = pi02 & n415;
  assign n417 = ~n411 & ~n416;
  assign n418 = n75 & ~n417;
  assign n419 = ~n410 & ~n418;
  assign n420 = ~pi01 & ~n260;
  assign n421 = ~n259 & ~n420;
  assign n422 = pi01 & n260;
  assign n423 = ~n421 & ~n422;
  assign n424 = ~n419 & n423;
  assign n425 = n419 & ~n423;
  assign n426 = ~n424 & ~n425;
  assign n427 = n165 & ~n426;
  assign n428 = n117 & n427;
  assign n429 = ~n408 & ~n428;
  assign n430 = ~pi02 & ~n429;
  assign n431 = n89 & n358;
  assign n432 = n93 & n419;
  assign n433 = ~n431 & ~n432;
  assign n434 = ~n292 & ~n295;
  assign n435 = ~n419 & ~n434;
  assign n436 = n419 & n434;
  assign n437 = ~n435 & ~n436;
  assign n438 = ~n433 & n437;
  assign n439 = n433 & ~n437;
  assign n440 = ~n438 & ~n439;
  assign n441 = n97 & ~n440;
  assign n442 = n367 & n433;
  assign n443 = ~n367 & ~n433;
  assign n444 = ~n442 & ~n443;
  assign n445 = ~n272 & ~n275;
  assign n446 = ~n444 & n445;
  assign n447 = n444 & ~n445;
  assign n448 = ~n446 & ~n447;
  assign n449 = n61 & ~n448;
  assign n450 = pi06 & n124;
  assign n451 = ~pi08 & n426;
  assign n452 = pi02 & n451;
  assign n453 = ~n450 & ~n452;
  assign n454 = ~n449 & n453;
  assign n455 = n117 & ~n454;
  assign n456 = n158 & ~n392;
  assign n457 = ~n367 & n456;
  assign n458 = ~n299 & ~n457;
  assign n459 = pi02 & ~n458;
  assign n460 = ~n318 & ~n321;
  assign n461 = ~n320 & ~n460;
  assign n462 = ~n367 & ~n461;
  assign n463 = n307 & n419;
  assign n464 = ~n307 & ~n419;
  assign n465 = ~n463 & ~n464;
  assign n466 = ~pi11 & ~n465;
  assign n467 = ~pi02 & n284;
  assign n468 = pi11 & n467;
  assign n469 = ~n284 & n337;
  assign n470 = ~n468 & ~n469;
  assign n471 = ~n466 & n470;
  assign n472 = n133 & ~n471;
  assign n473 = n318 & n367;
  assign n474 = ~n114 & n473;
  assign n475 = ~n472 & ~n474;
  assign n476 = ~n462 & n475;
  assign n477 = ~n459 & n476;
  assign n478 = ~n455 & n477;
  assign n479 = ~n441 & n478;
  assign n480 = ~n430 & n479;
  assign n481 = ~n406 & n480;
  assign n482 = ~n398 & n481;
  assign n483 = pi13 & ~n482;
  assign n484 = n333 & n483;
  assign n485 = ~n333 & ~n483;
  assign n486 = ~n484 & ~n485;
  assign po2 = ~n390 | n486;
  assign n488 = pi03 & pi11;
  assign n489 = ~pi07 & ~pi09;
  assign n490 = n85 & ~n489;
  assign n491 = n488 & ~n490;
  assign n492 = pi02 & ~pi06;
  assign n493 = ~pi02 & pi06;
  assign n494 = n203 & ~n493;
  assign n495 = ~n492 & ~n494;
  assign n496 = pi09 & ~n495;
  assign n497 = pi03 & n496;
  assign n498 = n193 & n497;
  assign n499 = n65 & ~n498;
  assign n500 = ~pi07 & ~n499;
  assign po5 = pi03 & pi07;
  assign n502 = n75 & n495;
  assign n503 = ~n91 & ~n502;
  assign n504 = po5 & ~n503;
  assign n505 = pi07 & n75;
  assign n506 = n496 & n505;
  assign n507 = ~n55 & ~n506;
  assign n508 = ~pi03 & ~n507;
  assign n509 = n152 & n337;
  assign n510 = ~pi03 & ~pi07;
  assign n511 = pi09 & n495;
  assign n512 = n510 & n511;
  assign n513 = ~n509 & ~n512;
  assign n514 = pi13 & ~n513;
  assign n515 = ~n508 & ~n514;
  assign n516 = ~n504 & n515;
  assign n517 = ~pi08 & ~n516;
  assign n518 = ~n46 & ~n92;
  assign n519 = po5 & ~n518;
  assign n520 = n37 & ~n510;
  assign n521 = ~n519 & ~n520;
  assign n522 = ~n517 & n521;
  assign n523 = ~n500 & n522;
  assign n524 = pi07 & n42;
  assign n525 = ~n159 & ~n524;
  assign n526 = ~n523 & ~n525;
  assign n527 = ~pi03 & n178;
  assign n528 = ~pi09 & n527;
  assign n529 = ~n72 & ~n528;
  assign n530 = pi07 & ~n529;
  assign n531 = ~n173 & n523;
  assign n532 = ~pi07 & n175;
  assign n533 = ~n531 & ~n532;
  assign n534 = ~pi09 & ~n533;
  assign n535 = pi03 & ~n523;
  assign n536 = n61 & n535;
  assign po4 = po5 | n510;
  assign n538 = ~n47 & ~n488;
  assign n539 = po4 & ~n538;
  assign n540 = ~n536 & ~n539;
  assign n541 = pi09 & ~n540;
  assign n542 = ~n534 & ~n541;
  assign n543 = ~n530 & n542;
  assign n544 = ~n526 & n543;
  assign n545 = ~n491 & n544;
  assign n546 = ~pi13 & ~n545;
  assign n547 = n155 & ~n546;
  assign n548 = ~n321 & ~n473;
  assign n549 = ~n320 & ~n548;
  assign n550 = ~n523 & ~n549;
  assign n551 = ~pi03 & n523;
  assign n552 = n73 & ~n551;
  assign n553 = n76 & n523;
  assign n554 = n39 & n535;
  assign n555 = n32 & po5;
  assign n556 = ~n554 & ~n555;
  assign n557 = ~n553 & n556;
  assign n558 = n75 & ~n557;
  assign n559 = ~n552 & ~n558;
  assign n560 = ~pi02 & n423;
  assign n561 = ~n419 & ~n560;
  assign n562 = pi02 & ~n423;
  assign n563 = ~n561 & ~n562;
  assign n564 = ~n559 & ~n563;
  assign n565 = n559 & n563;
  assign n566 = ~n564 & ~n565;
  assign n567 = ~pi08 & n566;
  assign n568 = ~pi03 & n567;
  assign n569 = ~n442 & ~n447;
  assign n570 = n89 & po5;
  assign n571 = n93 & n559;
  assign n572 = ~n570 & ~n571;
  assign n573 = n523 & n572;
  assign n574 = ~n523 & ~n572;
  assign n575 = ~n573 & ~n574;
  assign n576 = n569 & ~n575;
  assign n577 = ~n569 & n575;
  assign n578 = ~n576 & ~n577;
  assign n579 = pi08 & ~n578;
  assign n580 = ~n568 & ~n579;
  assign n581 = n91 & ~n580;
  assign n582 = n419 & ~n434;
  assign n583 = ~n439 & ~n582;
  assign n584 = ~n559 & ~n583;
  assign n585 = n559 & n583;
  assign n586 = ~n584 & ~n585;
  assign n587 = ~n572 & n586;
  assign n588 = n572 & ~n586;
  assign n589 = ~n587 & ~n588;
  assign n590 = n88 & ~n589;
  assign n591 = ~pi03 & n467;
  assign n592 = n133 & n591;
  assign n593 = ~n363 & ~n404;
  assign n594 = n510 & n593;
  assign n595 = n141 & n594;
  assign n596 = ~n592 & ~n595;
  assign n597 = ~n590 & n596;
  assign n598 = pi11 & ~n597;
  assign n599 = ~pi02 & n392;
  assign n600 = ~n367 & ~n599;
  assign n601 = pi02 & ~n392;
  assign n602 = ~n600 & ~n601;
  assign n603 = ~n523 & n602;
  assign n604 = n523 & ~n602;
  assign n605 = ~n603 & ~n604;
  assign n606 = n244 & ~n605;
  assign n607 = pi07 & ~n593;
  assign n608 = n141 & n607;
  assign n609 = ~n606 & ~n608;
  assign n610 = ~pi03 & ~n609;
  assign n611 = n463 & n559;
  assign n612 = ~n463 & ~n559;
  assign n613 = ~n611 & ~n612;
  assign n614 = n133 & ~n613;
  assign n615 = n76 & ~n566;
  assign n616 = pi03 & n615;
  assign n617 = pi07 & n141;
  assign n618 = ~n616 & ~n617;
  assign n619 = ~n614 & n618;
  assign n620 = ~pi11 & ~n619;
  assign n621 = po5 & n593;
  assign n622 = ~n510 & n593;
  assign n623 = ~po5 & ~n622;
  assign n624 = pi03 & n623;
  assign n625 = ~n621 & ~n624;
  assign n626 = n141 & ~n625;
  assign n627 = n158 & n605;
  assign n628 = ~n299 & ~n627;
  assign n629 = pi03 & ~n628;
  assign n630 = n473 & n523;
  assign n631 = ~n114 & n630;
  assign n632 = ~n467 & n488;
  assign n633 = n133 & n632;
  assign n634 = ~n631 & ~n633;
  assign n635 = ~n629 & n634;
  assign n636 = ~n626 & n635;
  assign n637 = ~n620 & n636;
  assign n638 = ~n610 & n637;
  assign n639 = ~n598 & n638;
  assign n640 = ~n581 & n639;
  assign n641 = ~n550 & n640;
  assign n642 = pi13 & ~n641;
  assign n643 = n484 & n642;
  assign n644 = ~n484 & ~n642;
  assign n645 = ~n643 & ~n644;
  assign po3 = ~n547 | n645;
  assign n647 = ~n40 & ~n113;
  assign n648 = n630 & ~n647;
  assign n649 = n559 & ~n583;
  assign n650 = ~n588 & ~n649;
  assign n651 = n88 & n650;
  assign n652 = n141 & ~n623;
  assign n653 = ~n551 & ~n602;
  assign n654 = ~n535 & ~n653;
  assign n655 = n157 & ~n654;
  assign n656 = ~n592 & ~n655;
  assign n657 = ~n652 & n656;
  assign n658 = ~n651 & n657;
  assign n659 = pi11 & ~n658;
  assign n660 = ~n573 & ~n577;
  assign n661 = pi08 & n660;
  assign n662 = ~pi08 & ~n565;
  assign n663 = ~n568 & n662;
  assign n664 = ~n661 & ~n663;
  assign n665 = n152 & ~n664;
  assign n666 = n39 & n611;
  assign n667 = ~n40 & ~n666;
  assign n668 = ~n665 & n667;
  assign n669 = ~pi11 & ~n668;
  assign n670 = ~n643 & ~n669;
  assign n671 = ~n659 & n670;
  assign n672 = ~n648 & n671;
  assign po6 = pi13 & ~n672;
  assign n674 = ~n142 & n191;
  assign n675 = ~n286 & ~n674;
  assign n676 = ~n377 & ~n675;
  assign n677 = n284 & ~n377;
  assign n678 = n203 & n677;
  assign n679 = ~n676 & ~n678;
  assign po7 = po4 & ~n679;
endmodule
