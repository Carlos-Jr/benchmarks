module top ( 
    pi0 , pi1 , pi2 , pi3 ,
    pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 ,
    po0 , po1 , po2 , po3 ,
    po4 , po5 , po6 , po7 ,
    po8 , po9 , po10   );
  input  pi0 , pi1 , pi2 ,
    pi3 , pi4 , pi5 , pi6 ,
    pi7 , pi8 , pi9 ;
  output po0 , po1 , po2 ,
    po3 , po4 , po5 , po6 ,
    po7 , po8 , po9 , po10 ;
  wire n22, n23, n24, n25, n26, n27, n28,
    n29, n30, n31, n32, n33, n34, n35, n36,
    n37, n38, n39, n40, n41, n42, n43, n44,
    n45, n46, n47, n48, n49, n50, n51, n52,
    n53, n54, n55, n56, n57, n58, n59, n60,
    n61, n62, n63, n64, n65, n66, n67, n68,
    n69, n70, n71, n72, n73, n74, n75, n76,
    n77, n78, n79, n80, n81, n82, n83, n84,
    n85, n86, n87, n88, n89, n90, n91, n92,
    n93, n94, n95, n96, n97, n98, n99,
    n100, n101, n102, n103, n104, n105, n106,
    n107, n108, n109, n110, n111, n112, n113,
    n114, n115, n116, n117, n118, n119, n120,
    n121, n122, n123, n124, n125, n126, n127,
    n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141,
    n142, n144, n145, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156,
    n157, n158, n159, n160, n161, n162, n163,
    n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177,
    n178, n179, n180, n181, n182, n183, n184,
    n185, n186, n187, n188, n189, n190, n191,
    n192, n193, n194, n195, n196, n197, n198,
    n199, n200, n201, n202, n203, n204, n205,
    n206, n207, n208, n209, n210, n211, n212,
    n213, n214, n215, n216, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226,
    n227, n228, n229, n230, n231, n232, n233,
    n234, n235, n236, n237, n238, n239, n240,
    n241, n242, n243, n244, n245, n246, n247,
    n248, n249, n250, n251, n252, n253, n255,
    n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339,
    n340, n341, n342, n343, n344, n345, n346,
    n347, n348, n349, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403,
    n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416, n417,
    n419, n420, n421, n422, n423, n424, n425,
    n427, n428, n429, n431, n432, n433, n434,
    n435, n436, n437, n438, n439, n440, n441,
    n442, n443, n444, n445, n446, n447, n448,
    n449, n450, n451, n452, n453, n454, n455,
    n456, n457, n458, n459, n460, n461, n462,
    n463, n464, n465, n466, n467, n468, n469,
    n470, n471, n472, n473, n474, n475, n476,
    n477, n478, n479, n480, n481, n482, n483,
    n484, n485, n486, n487, n488, n489, n490,
    n491, n492, n493, n494, n495, n496, n497,
    n498, n499, n500, n501, n502, n503, n504,
    n505, n506, n507, n508, n509, n510, n511,
    n512, n514, n515, n516, n517, n518, n519,
    n520, n521, n522, n523, n524, n525, n526,
    n527, n528, n529, n530, n531, n532, n533,
    n534, n535, n536, n537, n538, n539, n540,
    n541, n542, n543, n544, n545, n546, n547,
    n548, n549, n550, n551, n552, n553, n554,
    n555, n556, n557, n558, n559, n560, n561,
    n562, n563, n564, n565, n566, n567, n568,
    n569, n570, n571, n572, n573, n574, n575,
    n576, n577, n578, n579, n580, n581, n582,
    n583, n584, n585, n586, n587, n588, n589,
    n590, n591, n592, n593, n594, n596, n597,
    n598, n599, n600, n601, n602, n603, n604,
    n605, n606, n607, n608, n609, n610, n611,
    n612, n613, n614, n615, n616, n617, n618,
    n619, n620, n621, n622, n623, n624, n625,
    n626, n627, n628, n629, n630, n631, n632,
    n633, n634, n635, n636, n637, n638, n639,
    n640, n641, n642, n643, n644, n645, n646,
    n647, n648, n649, n650, n652, n653, n654,
    n655, n656, n657, n658, n659, n660, n661,
    n662, n663, n664, n665, n666, n667, n668,
    n669, n670, n671, n672, n673, n674, n675,
    n676, n677, n678, n679, n680, n681, n682,
    n683, n684, n685, n686, n687, n689, n690,
    n691, n692, n693, n694;
  assign n22 = ~pi1  & pi9 ;
  assign n23 = ~pi0  & pi9 ;
  assign n24 = pi1  & ~n23;
  assign n25 = ~pi3  & ~pi5 ;
  assign n26 = ~n24 & n25;
  assign n27 = ~n22 & n26;
  assign n28 = pi0  & ~pi9 ;
  assign n29 = ~pi1  & ~n28;
  assign n30 = pi1  & ~pi9 ;
  assign n31 = ~pi7  & ~n30;
  assign n32 = ~n29 & n31;
  assign n33 = ~n27 & ~n32;
  assign n34 = ~pi2  & ~n33;
  assign n35 = pi1  & ~pi3 ;
  assign n36 = ~pi2  & ~pi3 ;
  assign n37 = pi9  & ~n36;
  assign n38 = pi0  & pi3 ;
  assign n39 = ~n37 & ~n38;
  assign n40 = ~pi1  & ~n39;
  assign n41 = ~pi0  & pi5 ;
  assign n42 = pi0  & ~pi1 ;
  assign n43 = pi2  & ~n42;
  assign n44 = ~n41 & ~n43;
  assign n45 = ~pi9  & ~n44;
  assign n46 = ~n40 & ~n45;
  assign n47 = ~n35 & n46;
  assign n48 = ~pi7  & ~n47;
  assign n49 = ~n34 & ~n48;
  assign n50 = ~pi8  & ~n49;
  assign n51 = pi7  & pi8 ;
  assign n52 = ~pi5  & n51;
  assign n53 = ~pi7  & pi9 ;
  assign n54 = ~n52 & ~n53;
  assign n55 = pi1  & ~n54;
  assign n56 = pi1  & ~pi7 ;
  assign n57 = ~pi5  & ~pi9 ;
  assign n58 = ~n56 & n57;
  assign n59 = ~n55 & ~n58;
  assign n60 = pi0  & ~pi2 ;
  assign n61 = ~n59 & n60;
  assign n62 = ~pi0  & ~pi1 ;
  assign n63 = pi2  & ~pi9 ;
  assign n64 = n62 & n63;
  assign n65 = n52 & n64;
  assign n66 = ~n61 & ~n65;
  assign n67 = ~pi3  & ~n66;
  assign n68 = ~n50 & ~n67;
  assign n69 = ~pi6  & ~n68;
  assign n70 = ~pi0  & ~pi2 ;
  assign n71 = n22 & n70;
  assign n72 = ~pi5  & ~n71;
  assign n73 = pi6  & ~n72;
  assign n74 = pi1  & pi2 ;
  assign n75 = ~pi0  & ~pi9 ;
  assign n76 = pi0  & pi9 ;
  assign n77 = ~n75 & ~n76;
  assign n78 = pi5  & ~n77;
  assign n79 = n74 & n78;
  assign n80 = ~n73 & ~n79;
  assign n81 = pi8  & ~n80;
  assign n82 = ~pi1  & ~n23;
  assign n83 = ~pi8  & ~n82;
  assign n84 = n42 & n63;
  assign n85 = ~n83 & ~n84;
  assign n86 = ~pi5  & ~n85;
  assign n87 = ~n81 & ~n86;
  assign n88 = pi3  & ~n87;
  assign n89 = ~pi2  & ~n28;
  assign n90 = pi6  & ~n89;
  assign n91 = pi1  & ~n77;
  assign n92 = n36 & n91;
  assign n93 = ~n90 & ~n92;
  assign n94 = pi5  & ~n93;
  assign n95 = ~pi2  & pi9 ;
  assign n96 = ~n63 & ~n95;
  assign n97 = ~pi0  & ~pi3 ;
  assign n98 = ~pi1  & ~pi9 ;
  assign n99 = pi6  & ~n98;
  assign n100 = n97 & n99;
  assign n101 = n96 & n100;
  assign n102 = ~n94 & ~n101;
  assign n103 = pi8  & ~n102;
  assign n104 = pi1  & ~pi8 ;
  assign n105 = pi2  & ~pi3 ;
  assign n106 = n22 & n105;
  assign n107 = ~n104 & ~n106;
  assign n108 = ~pi0  & ~n107;
  assign n109 = pi2  & pi9 ;
  assign n110 = ~pi2  & pi6 ;
  assign n111 = pi3  & ~n110;
  assign n112 = n98 & ~n111;
  assign n113 = ~n109 & ~n112;
  assign n114 = ~pi8  & ~n113;
  assign n115 = ~n108 & ~n114;
  assign n116 = ~pi5  & ~n115;
  assign n117 = ~n103 & ~n116;
  assign n118 = ~n88 & n117;
  assign n119 = ~pi0  & ~pi8 ;
  assign n120 = n36 & n119;
  assign n121 = n98 & n120;
  assign n122 = n118 & ~n121;
  assign n123 = ~pi7  & ~n122;
  assign n124 = ~n69 & ~n123;
  assign n125 = ~pi4  & ~n124;
  assign n126 = ~pi8  & ~pi9 ;
  assign n127 = ~pi6  & n126;
  assign n128 = pi4  & pi8 ;
  assign n129 = pi6  & n128;
  assign n130 = ~n127 & ~n129;
  assign n131 = pi5  & ~n130;
  assign n132 = ~pi6  & pi9 ;
  assign n133 = ~pi5  & pi6 ;
  assign n134 = ~n132 & ~n133;
  assign n135 = ~pi4  & pi9 ;
  assign n136 = ~pi8  & ~n135;
  assign n137 = ~n134 & n136;
  assign n138 = ~n131 & ~n137;
  assign n139 = ~pi1  & ~pi3 ;
  assign n140 = ~n138 & n139;
  assign n141 = ~pi7  & n140;
  assign n142 = n70 & n141;
  assign po0  = n125 | n142;
  assign n144 = pi0  & pi8 ;
  assign n145 = n109 & n144;
  assign n146 = ~pi2  & ~pi8 ;
  assign n147 = ~pi0  & n146;
  assign n148 = ~pi9  & n147;
  assign n149 = ~n145 & ~n148;
  assign n150 = pi5  & ~n149;
  assign n151 = ~pi5  & pi8 ;
  assign n152 = pi6  & pi9 ;
  assign n153 = ~n151 & ~n152;
  assign n154 = ~pi0  & ~n153;
  assign n155 = ~pi8  & n57;
  assign n156 = pi8  & n152;
  assign n157 = ~n155 & ~n156;
  assign n158 = ~n154 & n157;
  assign n159 = pi2  & ~n158;
  assign n160 = ~n150 & ~n159;
  assign n161 = ~pi4  & ~n160;
  assign n162 = pi4  & pi9 ;
  assign n163 = pi5  & ~pi8 ;
  assign n164 = ~n128 & ~n163;
  assign n165 = ~pi6  & ~n164;
  assign n166 = ~n162 & ~n165;
  assign n167 = ~n132 & ~n166;
  assign n168 = n70 & n167;
  assign n169 = ~n161 & ~n168;
  assign n170 = ~pi1  & ~n169;
  assign n171 = ~pi8  & pi9 ;
  assign n172 = n41 & n171;
  assign n173 = pi6  & pi8 ;
  assign n174 = ~n153 & ~n173;
  assign n175 = pi0  & n174;
  assign n176 = ~n172 & ~n175;
  assign n177 = ~pi2  & ~n176;
  assign n178 = ~pi6  & ~pi8 ;
  assign n179 = ~pi0  & pi6 ;
  assign n180 = ~pi2  & ~n179;
  assign n181 = n151 & ~n180;
  assign n182 = ~n178 & ~n181;
  assign n183 = ~pi9  & ~n182;
  assign n184 = ~n177 & ~n183;
  assign n185 = pi1  & ~n184;
  assign n186 = ~pi6  & pi8 ;
  assign n187 = n63 & n186;
  assign n188 = ~n185 & ~n187;
  assign n189 = ~pi4  & ~n188;
  assign n190 = ~n170 & ~n189;
  assign n191 = ~pi3  & ~n190;
  assign n192 = ~pi2  & pi8 ;
  assign n193 = pi0  & n192;
  assign n194 = pi0  & ~pi5 ;
  assign n195 = ~n193 & ~n194;
  assign n196 = ~n41 & n195;
  assign n197 = pi1  & ~n196;
  assign n198 = pi3  & pi8 ;
  assign n199 = ~pi2  & ~n198;
  assign n200 = ~pi0  & ~n199;
  assign n201 = pi5  & n146;
  assign n202 = ~pi3  & ~pi8 ;
  assign n203 = ~n151 & ~n202;
  assign n204 = pi0  & n203;
  assign n205 = ~n201 & ~n204;
  assign n206 = ~pi1  & ~n205;
  assign n207 = ~n200 & ~n206;
  assign n208 = ~n197 & n207;
  assign n209 = ~pi6  & ~n208;
  assign n210 = ~pi1  & pi6 ;
  assign n211 = pi2  & ~n210;
  assign n212 = ~pi1  & ~pi8 ;
  assign n213 = pi3  & ~n212;
  assign n214 = ~n211 & n213;
  assign n215 = ~pi0  & pi8 ;
  assign n216 = pi0  & pi1 ;
  assign n217 = ~pi1  & ~pi6 ;
  assign n218 = ~pi2  & ~n217;
  assign n219 = ~n216 & n218;
  assign n220 = ~n215 & n219;
  assign n221 = ~n214 & ~n220;
  assign n222 = ~pi5  & ~n221;
  assign n223 = ~pi9  & ~n222;
  assign n224 = ~n209 & n223;
  assign n225 = ~pi4  & ~n224;
  assign n226 = pi1  & pi5 ;
  assign n227 = ~pi1  & ~pi2 ;
  assign n228 = pi3  & ~pi8 ;
  assign n229 = n227 & n228;
  assign n230 = ~n226 & ~n229;
  assign n231 = pi0  & ~n230;
  assign n232 = pi5  & ~n36;
  assign n233 = ~n231 & ~n232;
  assign n234 = pi6  & ~n233;
  assign n235 = pi3  & n74;
  assign n236 = ~pi6  & ~n163;
  assign n237 = n235 & ~n236;
  assign n238 = pi9  & ~n237;
  assign n239 = ~n234 & n238;
  assign n240 = n225 & ~n239;
  assign n241 = ~n191 & ~n240;
  assign n242 = ~pi7  & ~n241;
  assign n243 = n30 & n192;
  assign n244 = n89 & ~n216;
  assign n245 = pi2  & ~n62;
  assign n246 = ~pi8  & ~n245;
  assign n247 = ~n244 & n246;
  assign n248 = ~n243 & ~n247;
  assign n249 = pi7  & ~n248;
  assign n250 = ~n64 & ~n249;
  assign n251 = n25 & ~n250;
  assign n252 = ~pi4  & n251;
  assign n253 = ~pi6  & n252;
  assign po1  = n242 | n253;
  assign n255 = pi3  & ~n192;
  assign n256 = pi5  & ~n255;
  assign n257 = pi2  & ~pi5 ;
  assign n258 = pi3  & ~n257;
  assign n259 = pi8  & ~n258;
  assign n260 = ~n256 & ~n259;
  assign n261 = pi1  & ~n260;
  assign n262 = ~pi3  & n133;
  assign n263 = n212 & n262;
  assign n264 = ~n261 & ~n263;
  assign n265 = ~pi9  & ~n264;
  assign n266 = pi1  & pi8 ;
  assign n267 = pi6  & ~n266;
  assign n268 = ~pi9  & ~n267;
  assign n269 = ~pi2  & ~n268;
  assign n270 = ~pi8  & n22;
  assign n271 = ~n269 & ~n270;
  assign n272 = pi3  & ~n271;
  assign n273 = pi6  & ~pi8 ;
  assign n274 = ~pi3  & pi9 ;
  assign n275 = pi1  & n274;
  assign n276 = n273 & n275;
  assign n277 = ~n272 & ~n276;
  assign n278 = pi2  & ~n186;
  assign n279 = pi1  & ~n278;
  assign n280 = ~n199 & ~n279;
  assign n281 = pi5  & n280;
  assign n282 = n277 & ~n281;
  assign n283 = ~n265 & n282;
  assign n284 = ~n98 & ~n274;
  assign n285 = pi3  & ~n171;
  assign n286 = ~pi6  & ~n285;
  assign n287 = n284 & n286;
  assign n288 = n283 & ~n287;
  assign n289 = ~pi4  & ~n288;
  assign n290 = ~pi3  & pi4 ;
  assign n291 = pi8  & ~pi9 ;
  assign n292 = ~pi5  & ~n291;
  assign n293 = ~n178 & n292;
  assign n294 = n290 & ~n293;
  assign n295 = n227 & n294;
  assign n296 = ~n289 & ~n295;
  assign n297 = ~pi0  & ~n296;
  assign n298 = ~pi5  & n109;
  assign n299 = ~n171 & ~n291;
  assign n300 = pi5  & ~n215;
  assign n301 = n299 & n300;
  assign n302 = ~n298 & ~n301;
  assign n303 = pi1  & ~n302;
  assign n304 = ~n98 & n299;
  assign n305 = pi2  & ~n304;
  assign n306 = ~n303 & ~n305;
  assign n307 = ~pi3  & ~n306;
  assign n308 = ~pi1  & pi8 ;
  assign n309 = n37 & n308;
  assign n310 = ~pi1  & pi3 ;
  assign n311 = pi5  & ~n310;
  assign n312 = ~pi2  & ~n311;
  assign n313 = n126 & n312;
  assign n314 = ~n309 & ~n313;
  assign n315 = pi0  & ~n314;
  assign n316 = ~n307 & ~n315;
  assign n317 = ~pi6  & ~n316;
  assign n318 = pi6  & ~n22;
  assign n319 = ~n30 & ~n318;
  assign n320 = pi8  & ~n319;
  assign n321 = pi1  & pi9 ;
  assign n322 = ~n98 & ~n321;
  assign n323 = n202 & ~n322;
  assign n324 = ~n320 & ~n323;
  assign n325 = ~pi2  & ~n324;
  assign n326 = pi2  & n321;
  assign n327 = ~n308 & ~n326;
  assign n328 = pi6  & ~n327;
  assign n329 = pi8  & ~n63;
  assign n330 = pi2  & n126;
  assign n331 = ~n329 & ~n330;
  assign n332 = ~n328 & n331;
  assign n333 = pi3  & ~n332;
  assign n334 = ~n325 & ~n333;
  assign n335 = n194 & ~n334;
  assign n336 = ~n317 & ~n335;
  assign n337 = ~pi4  & ~n336;
  assign n338 = ~n297 & ~n337;
  assign n339 = ~pi7  & ~n338;
  assign n340 = ~pi5  & ~pi6 ;
  assign n341 = pi8  & pi9 ;
  assign n342 = pi7  & n341;
  assign n343 = pi0  & ~n342;
  assign n344 = n24 & ~n343;
  assign n345 = n28 & n212;
  assign n346 = ~n344 & ~n345;
  assign n347 = n340 & ~n346;
  assign n348 = ~pi4  & n347;
  assign n349 = n36 & n348;
  assign po2  = n339 | n349;
  assign n351 = pi6  & ~n36;
  assign n352 = pi3  & ~pi9 ;
  assign n353 = ~n351 & ~n352;
  assign n354 = ~pi4  & ~n353;
  assign n355 = pi5  & pi6 ;
  assign n356 = ~n340 & ~n355;
  assign n357 = ~pi2  & n290;
  assign n358 = ~pi6  & ~n341;
  assign n359 = n357 & ~n358;
  assign n360 = ~n356 & n359;
  assign n361 = ~n354 & ~n360;
  assign n362 = ~pi1  & ~n361;
  assign n363 = pi5  & ~n186;
  assign n364 = ~pi3  & ~n273;
  assign n365 = pi5  & pi9 ;
  assign n366 = ~n126 & ~n365;
  assign n367 = pi2  & ~n366;
  assign n368 = n364 & ~n367;
  assign n369 = pi1  & ~n368;
  assign n370 = ~n363 & n369;
  assign n371 = pi2  & n133;
  assign n372 = ~n370 & ~n371;
  assign n373 = ~pi4  & ~n372;
  assign n374 = ~n362 & ~n373;
  assign n375 = ~pi0  & ~n374;
  assign n376 = pi2  & ~n203;
  assign n377 = pi5  & n192;
  assign n378 = ~n376 & ~n377;
  assign n379 = ~pi9  & ~n378;
  assign n380 = pi5  & n171;
  assign n381 = ~pi3  & ~n380;
  assign n382 = ~pi2  & ~n381;
  assign n383 = ~pi6  & ~n228;
  assign n384 = pi3  & ~pi5 ;
  assign n385 = ~n383 & ~n384;
  assign n386 = ~n382 & ~n385;
  assign n387 = ~n379 & n386;
  assign n388 = pi1  & ~n387;
  assign n389 = n201 & n217;
  assign n390 = ~n262 & ~n389;
  assign n391 = ~pi9  & ~n390;
  assign n392 = ~n388 & ~n391;
  assign n393 = pi0  & ~n392;
  assign n394 = ~pi9  & n133;
  assign n395 = n266 & n394;
  assign n396 = pi3  & ~pi6 ;
  assign n397 = pi2  & n396;
  assign n398 = ~n36 & n133;
  assign n399 = ~n397 & ~n398;
  assign n400 = pi9  & ~n399;
  assign n401 = ~n394 & ~n396;
  assign n402 = ~pi8  & ~n401;
  assign n403 = ~n400 & ~n402;
  assign n404 = ~pi1  & ~n403;
  assign n405 = ~n57 & ~n178;
  assign n406 = ~pi2  & ~n405;
  assign n407 = ~pi6  & ~n365;
  assign n408 = pi5  & pi8 ;
  assign n409 = ~n321 & ~n408;
  assign n410 = n407 & ~n409;
  assign n411 = ~n406 & ~n410;
  assign n412 = pi3  & ~n411;
  assign n413 = ~n404 & ~n412;
  assign n414 = ~n395 & n413;
  assign n415 = ~n393 & n414;
  assign n416 = ~pi4  & ~n415;
  assign n417 = ~n375 & ~n416;
  assign po3  = ~pi7  & ~n417;
  assign n419 = ~pi4  & n245;
  assign n420 = pi3  & ~pi4 ;
  assign n421 = ~n290 & ~n420;
  assign n422 = ~pi0  & n227;
  assign n423 = ~n421 & n422;
  assign n424 = ~n419 & ~n423;
  assign n425 = ~pi7  & n355;
  assign po4  = ~n424 & n425;
  assign n427 = n420 & ~n422;
  assign n428 = n62 & n357;
  assign n429 = ~n427 & ~n428;
  assign po5  = n425 & ~n429;
  assign n431 = ~pi0  & n109;
  assign n432 = ~pi9  & n212;
  assign n433 = ~n431 & ~n432;
  assign n434 = pi5  & ~n433;
  assign n435 = pi5  & n321;
  assign n436 = ~pi1  & ~pi5 ;
  assign n437 = pi2  & ~n436;
  assign n438 = ~pi6  & ~n437;
  assign n439 = ~pi9  & n438;
  assign n440 = ~n435 & ~n439;
  assign n441 = pi0  & ~n440;
  assign n442 = ~pi0  & pi2 ;
  assign n443 = ~n57 & n442;
  assign n444 = ~n441 & ~n443;
  assign n445 = pi8  & ~n444;
  assign n446 = pi2  & pi8 ;
  assign n447 = ~n146 & ~n446;
  assign n448 = pi6  & ~n447;
  assign n449 = n96 & n448;
  assign n450 = ~n445 & ~n449;
  assign n451 = ~n434 & n450;
  assign n452 = ~pi7  & ~n451;
  assign n453 = pi7  & ~pi9 ;
  assign n454 = pi8  & ~n453;
  assign n455 = pi2  & ~n454;
  assign n456 = ~n30 & ~n455;
  assign n457 = ~pi0  & ~n456;
  assign n458 = ~n74 & n457;
  assign n459 = pi8  & n76;
  assign n460 = pi1  & n459;
  assign n461 = ~n126 & ~n460;
  assign n462 = ~pi2  & ~n461;
  assign n463 = pi7  & n462;
  assign n464 = ~n458 & ~n463;
  assign n465 = n340 & ~n464;
  assign n466 = ~n452 & ~n465;
  assign n467 = ~pi3  & ~n466;
  assign n468 = pi2  & n30;
  assign n469 = ~pi1  & ~n126;
  assign n470 = ~n30 & ~n469;
  assign n471 = pi0  & n470;
  assign n472 = ~n468 & ~n471;
  assign n473 = ~pi0  & ~pi6 ;
  assign n474 = ~n212 & n322;
  assign n475 = n473 & n474;
  assign n476 = n472 & ~n475;
  assign n477 = ~pi5  & ~n476;
  assign n478 = n104 & ~n442;
  assign n479 = pi0  & n173;
  assign n480 = ~pi2  & n479;
  assign n481 = ~n478 & ~n480;
  assign n482 = pi9  & ~n481;
  assign n483 = ~n119 & ~n194;
  assign n484 = n30 & n483;
  assign n485 = ~n482 & ~n484;
  assign n486 = ~n477 & n485;
  assign n487 = pi3  & ~n486;
  assign n488 = ~pi6  & ~n257;
  assign n489 = n23 & ~n488;
  assign n490 = ~pi2  & pi5 ;
  assign n491 = ~n77 & n490;
  assign n492 = ~n489 & ~n491;
  assign n493 = ~pi8  & ~n492;
  assign n494 = pi2  & ~n126;
  assign n495 = ~n459 & ~n494;
  assign n496 = pi6  & ~n495;
  assign n497 = ~n493 & ~n496;
  assign n498 = pi1  & ~n497;
  assign n499 = pi8  & ~n194;
  assign n500 = ~pi9  & ~n473;
  assign n501 = ~pi2  & n500;
  assign n502 = ~n499 & n501;
  assign n503 = n23 & n446;
  assign n504 = ~n502 & ~n503;
  assign n505 = ~pi1  & ~n504;
  assign n506 = ~n498 & ~n505;
  assign n507 = ~n487 & n506;
  assign n508 = ~pi7  & ~n507;
  assign n509 = ~n467 & ~n508;
  assign n510 = ~pi4  & ~n509;
  assign n511 = ~n355 & ~n428;
  assign n512 = ~pi7  & ~n511;
  assign po6  = ~n510 & ~n512;
  assign n514 = pi3  & ~n341;
  assign n515 = ~n144 & ~n514;
  assign n516 = ~pi6  & ~n515;
  assign n517 = ~pi3  & n341;
  assign n518 = ~n516 & ~n517;
  assign n519 = pi2  & ~n518;
  assign n520 = ~pi3  & n127;
  assign n521 = ~n126 & ~n178;
  assign n522 = pi3  & ~n152;
  assign n523 = pi0  & ~n522;
  assign n524 = n521 & n523;
  assign n525 = pi6  & n291;
  assign n526 = n215 & n396;
  assign n527 = ~n273 & ~n526;
  assign n528 = pi9  & ~n527;
  assign n529 = ~n525 & ~n528;
  assign n530 = ~n524 & n529;
  assign n531 = ~pi2  & ~n530;
  assign n532 = ~n520 & ~n531;
  assign n533 = ~n519 & n532;
  assign n534 = pi1  & ~n533;
  assign n535 = n89 & n358;
  assign n536 = n179 & n299;
  assign n537 = ~n535 & ~n536;
  assign n538 = pi3  & ~n537;
  assign n539 = ~n147 & ~n479;
  assign n540 = ~pi9  & ~n539;
  assign n541 = ~pi6  & ~n202;
  assign n542 = n494 & ~n541;
  assign n543 = ~n540 & ~n542;
  assign n544 = ~n538 & n543;
  assign n545 = ~pi1  & ~n544;
  assign n546 = ~pi2  & pi3 ;
  assign n547 = ~pi9  & n273;
  assign n548 = n546 & n547;
  assign n549 = ~n545 & ~n548;
  assign n550 = ~n534 & n549;
  assign n551 = ~pi5  & ~n550;
  assign n552 = n38 & n330;
  assign n553 = pi2  & pi3 ;
  assign n554 = ~n299 & ~n553;
  assign n555 = ~pi2  & ~n38;
  assign n556 = pi5  & ~n555;
  assign n557 = ~n554 & n556;
  assign n558 = ~n552 & ~n557;
  assign n559 = ~pi1  & ~n558;
  assign n560 = pi8  & n365;
  assign n561 = n553 & n560;
  assign n562 = pi3  & pi5 ;
  assign n563 = ~n63 & ~n562;
  assign n564 = ~pi0  & ~n563;
  assign n565 = pi5  & n546;
  assign n566 = ~n564 & ~n565;
  assign n567 = ~pi8  & ~n566;
  assign n568 = pi0  & ~n96;
  assign n569 = ~pi9  & n41;
  assign n570 = ~n568 & ~n569;
  assign n571 = pi8  & ~n570;
  assign n572 = n109 & n163;
  assign n573 = ~n571 & ~n572;
  assign n574 = ~pi3  & ~n573;
  assign n575 = ~pi9  & n565;
  assign n576 = ~n574 & ~n575;
  assign n577 = ~n567 & n576;
  assign n578 = pi1  & ~n577;
  assign n579 = ~n561 & ~n578;
  assign n580 = ~n559 & n579;
  assign n581 = ~pi6  & ~n580;
  assign n582 = ~n551 & ~n581;
  assign n583 = ~pi7  & ~n582;
  assign n584 = ~n299 & n442;
  assign n585 = n193 & n453;
  assign n586 = ~n584 & ~n585;
  assign n587 = n25 & ~n586;
  assign n588 = n217 & n587;
  assign n589 = ~n583 & ~n588;
  assign n590 = ~pi4  & ~n589;
  assign n591 = pi4  & ~pi7 ;
  assign n592 = n25 & n591;
  assign n593 = n70 & n592;
  assign n594 = n217 & n593;
  assign po7  = ~n590 & ~n594;
  assign n596 = ~pi2  & ~n384;
  assign n597 = ~n226 & n596;
  assign n598 = n284 & n597;
  assign n599 = n98 & n490;
  assign n600 = ~n275 & ~n599;
  assign n601 = ~pi0  & ~n600;
  assign n602 = n322 & ~n436;
  assign n603 = n105 & ~n602;
  assign n604 = ~n601 & ~n603;
  assign n605 = ~n598 & n604;
  assign n606 = ~pi8  & ~n605;
  assign n607 = ~n97 & n597;
  assign n608 = n25 & n42;
  assign n609 = ~n607 & ~n608;
  assign n610 = pi8  & ~n609;
  assign n611 = ~pi5  & ~n215;
  assign n612 = ~n562 & ~n611;
  assign n613 = n74 & n612;
  assign n614 = ~n610 & ~n613;
  assign n615 = ~pi9  & ~n614;
  assign n616 = ~n25 & ~n490;
  assign n617 = pi1  & ~n616;
  assign n618 = ~n199 & n617;
  assign n619 = ~n41 & n310;
  assign n620 = n192 & n619;
  assign n621 = ~n618 & ~n620;
  assign n622 = pi9  & ~n621;
  assign n623 = ~n615 & ~n622;
  assign n624 = ~n606 & n623;
  assign n625 = ~pi6  & ~n624;
  assign n626 = pi2  & ~n469;
  assign n627 = ~n318 & ~n626;
  assign n628 = pi0  & ~n627;
  assign n629 = ~pi6  & ~n104;
  assign n630 = pi2  & ~n629;
  assign n631 = ~n341 & ~n469;
  assign n632 = pi6  & n631;
  assign n633 = ~n630 & ~n632;
  assign n634 = ~n628 & n633;
  assign n635 = n384 & ~n634;
  assign n636 = ~n625 & ~n635;
  assign n637 = ~pi7  & ~n636;
  assign n638 = ~pi0  & ~n447;
  assign n639 = ~n193 & ~n638;
  assign n640 = ~pi9  & ~n639;
  assign n641 = ~pi8  & n431;
  assign n642 = ~n640 & ~n641;
  assign n643 = ~pi1  & ~n642;
  assign n644 = n147 & n321;
  assign n645 = ~n643 & ~n644;
  assign n646 = ~pi6  & ~n645;
  assign n647 = n25 & n646;
  assign n648 = ~n637 & ~n647;
  assign n649 = ~pi4  & ~n648;
  assign n650 = ~pi1  & n593;
  assign po8  = ~n649 & ~n650;
  assign n652 = n194 & n397;
  assign n653 = ~pi7  & ~n652;
  assign n654 = ~n469 & ~n653;
  assign n655 = ~pi2  & n139;
  assign n656 = ~pi7  & ~n655;
  assign n657 = pi0  & ~n656;
  assign n658 = pi4  & ~n655;
  assign n659 = ~pi3  & ~n57;
  assign n660 = n215 & ~n522;
  assign n661 = ~n659 & ~n660;
  assign n662 = ~pi2  & ~n661;
  assign n663 = ~pi6  & ~n560;
  assign n664 = ~pi3  & ~n663;
  assign n665 = n340 & ~n341;
  assign n666 = n553 & n665;
  assign n667 = ~n664 & ~n666;
  assign n668 = ~n662 & n667;
  assign n669 = pi1  & ~n668;
  assign n670 = ~pi5  & ~n105;
  assign n671 = pi6  & ~n670;
  assign n672 = pi7  & ~n105;
  assign n673 = n215 & ~n407;
  assign n674 = n522 & ~n673;
  assign n675 = n290 & ~n340;
  assign n676 = ~pi2  & ~n675;
  assign n677 = ~n674 & n676;
  assign n678 = ~pi8  & ~n365;
  assign n679 = pi2  & ~n678;
  assign n680 = n659 & n679;
  assign n681 = ~n677 & ~n680;
  assign n682 = ~pi1  & ~n681;
  assign n683 = ~n672 & ~n682;
  assign n684 = ~n671 & n683;
  assign n685 = ~n669 & n684;
  assign n686 = ~n658 & n685;
  assign n687 = ~n657 & n686;
  assign po9  = ~n654 & n687;
  assign n689 = pi8  & ~n24;
  assign n690 = pi2  & ~n689;
  assign n691 = ~n29 & n690;
  assign n692 = n420 & n691;
  assign n693 = ~n428 & ~n692;
  assign n694 = n340 & ~n693;
  assign po10  = ~pi7  & n694;
endmodule
