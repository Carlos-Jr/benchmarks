module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 , pi32 ,
    pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 , pi40 ,
    pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 , pi56 ,
    pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 , pi64 ,
    pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 ,
    pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 ,
    pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 ,
    pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 ,
    pi97 , pi98 , pi99 , pi100 , pi101 , pi102 , pi103 ,
    pi104 , pi105 , pi106 , pi107 , pi108 , pi109 , pi110 ,
    pi111 , pi112 , pi113 , pi114 , pi115 , pi116 , pi117 ,
    pi118 , pi119 , pi120 , pi121 , pi122 , pi123 , pi124 ,
    pi125 , pi126 , pi127 ,
    po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7  );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    pi32 , pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 ,
    pi56 , pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 ,
    pi64 , pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 ,
    pi72 , pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 ,
    pi80 , pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 ,
    pi88 , pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 ,
    pi96 , pi97 , pi98 , pi99 , pi100 , pi101 , pi102 ,
    pi103 , pi104 , pi105 , pi106 , pi107 , pi108 , pi109 ,
    pi110 , pi111 , pi112 , pi113 , pi114 , pi115 , pi116 ,
    pi117 , pi118 , pi119 , pi120 , pi121 , pi122 , pi123 ,
    pi124 , pi125 , pi126 , pi127 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7;
  wire n137, n138, n139, n140, n141, n142, n143,
    n144, n145, n146, n147, n148, n149, n150,
    n151, n152, n153, n154, n155, n156, n157,
    n158, n159, n160, n161, n162, n163, n164,
    n165, n166, n167, n168, n169, n170, n171,
    n172, n173, n174, n175, n176, n177, n178,
    n179, n180, n181, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192,
    n193, n194, n195, n196, n197, n198, n199,
    n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213,
    n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227,
    n228, n229, n230, n231, n232, n233, n234,
    n235, n236, n237, n238, n239, n240, n241,
    n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339,
    n340, n341, n342, n343, n344, n345, n346,
    n347, n348, n349, n350, n351, n352, n353,
    n354, n355, n356, n357, n358, n359, n360,
    n361, n362, n363, n364, n365, n366, n367,
    n368, n369, n370, n371, n372, n373, n374,
    n375, n376, n377, n378, n379, n380, n381,
    n382, n383, n384, n385, n386, n387, n388,
    n389, n390, n391, n392, n393, n394, n395,
    n396, n397, n398, n399, n400, n401, n402,
    n403, n404, n405, n406, n407, n408, n409,
    n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423,
    n424, n425, n426, n427, n428, n429, n430,
    n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444,
    n445, n446, n447, n448, n449, n450, n451,
    n452, n453, n454, n455, n456, n457, n458,
    n459, n460, n461, n462, n463, n464, n465,
    n466, n467, n468, n469, n470, n471, n472,
    n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487,
    n488, n489, n490, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501,
    n502, n503, n504, n505, n506, n507, n508,
    n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n541, n542, n543,
    n544, n545, n546, n547, n548, n549, n550,
    n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564,
    n565, n566, n567, n568, n569, n570, n571,
    n572, n573, n574, n575, n576, n577, n578,
    n579, n580, n581, n582, n583, n584, n585,
    n586, n587, n588, n589, n590, n591, n592,
    n593, n594, n595, n596, n597, n598, n599,
    n600, n601, n602, n603, n604, n605, n606,
    n607, n608, n609, n610, n611, n612, n613,
    n614, n615, n616, n617, n618, n619, n620,
    n621, n622, n623, n624, n625, n626, n627,
    n628, n629, n630, n631, n632, n633, n634,
    n635, n636, n637, n638, n639, n640, n641,
    n642, n643, n644, n645, n646, n647, n648,
    n649, n650, n651, n652, n653, n654, n655,
    n656, n657, n658, n659, n660, n661, n662,
    n663, n664, n665, n666, n667, n668, n669,
    n670, n671, n672, n673, n674, n675, n676,
    n677, n678, n679, n680, n681, n682, n684,
    n685, n686, n687, n688, n689, n690, n691,
    n692, n693, n694, n695, n696, n697, n698,
    n699, n700, n701, n702, n703, n704, n705,
    n706, n707, n708, n709, n710, n711, n712,
    n713, n714, n715, n716, n717, n718, n719,
    n720, n721, n722, n723, n724, n725, n726,
    n727, n728, n729, n730, n731, n732, n733,
    n734, n735, n736, n737, n738, n739, n740,
    n741, n742, n743, n744, n745, n746, n747,
    n748, n749, n750, n751, n752, n753, n754,
    n755, n756, n757, n758, n759, n761, n762,
    n763, n764, n765, n766, n767, n768, n769,
    n770, n771, n772, n773, n774, n775, n776,
    n777, n778, n779, n780, n781, n782, n783,
    n784, n785, n786, n787, n788, n789, n790,
    n791, n792, n794, n795, n796, n797, n798,
    n799, n800, n801, n802, n803, n804, n805,
    n807, n808, n809, n810, n813, n814, n815,
    n816, n817, n818;
  assign n137 = pi1  & ~pi2 ;
  assign n138 = ~pi3  & ~n137;
  assign n139 = ~pi4  & ~n138;
  assign n140 = ~pi5  & ~n139;
  assign n141 = ~pi6  & ~n140;
  assign n142 = ~pi7  & ~n141;
  assign n143 = ~pi8  & ~n142;
  assign n144 = ~pi9  & ~n143;
  assign n145 = ~pi10  & ~n144;
  assign n146 = ~pi11  & ~n145;
  assign n147 = ~pi12  & ~n146;
  assign n148 = ~pi13  & ~n147;
  assign n149 = ~pi116  & pi118 ;
  assign n150 = ~pi119  & n149;
  assign n151 = pi117  & ~pi118 ;
  assign n152 = ~pi119  & ~n151;
  assign n153 = pi116  & n152;
  assign n154 = ~pi120  & ~n150;
  assign n155 = ~n153 & n154;
  assign n156 = ~pi114  & ~n155;
  assign n157 = ~pi120  & ~n152;
  assign n158 = ~pi115  & ~n157;
  assign n159 = pi115  & ~n155;
  assign n160 = ~n158 & ~n159;
  assign n161 = pi114  & ~n160;
  assign n162 = ~n156 & ~n161;
  assign n163 = ~pi112  & ~n162;
  assign n164 = ~pi113  & ~n160;
  assign n165 = pi113  & ~n162;
  assign n166 = ~n164 & ~n165;
  assign n167 = pi112  & ~n166;
  assign n168 = ~n163 & ~n167;
  assign n169 = ~pi110  & ~n168;
  assign n170 = ~pi111  & ~n166;
  assign n171 = pi111  & ~n168;
  assign n172 = ~n170 & ~n171;
  assign n173 = pi110  & ~n172;
  assign n174 = ~n169 & ~n173;
  assign n175 = ~pi108  & ~n174;
  assign n176 = ~pi109  & ~n172;
  assign n177 = pi109  & ~n174;
  assign n178 = ~n176 & ~n177;
  assign n179 = pi108  & ~n178;
  assign n180 = ~n175 & ~n179;
  assign n181 = ~pi106  & ~n180;
  assign n182 = ~pi107  & ~n178;
  assign n183 = pi107  & ~n180;
  assign n184 = ~n182 & ~n183;
  assign n185 = pi106  & ~n184;
  assign n186 = ~n181 & ~n185;
  assign n187 = ~pi104  & ~n186;
  assign n188 = ~pi105  & ~n184;
  assign n189 = pi105  & ~n186;
  assign n190 = ~n188 & ~n189;
  assign n191 = pi104  & ~n190;
  assign n192 = ~n187 & ~n191;
  assign n193 = ~pi102  & ~n192;
  assign n194 = ~pi103  & ~n190;
  assign n195 = pi103  & ~n192;
  assign n196 = ~n194 & ~n195;
  assign n197 = pi102  & ~n196;
  assign n198 = ~n193 & ~n197;
  assign n199 = ~pi100  & ~n198;
  assign n200 = ~pi101  & ~n196;
  assign n201 = pi101  & ~n198;
  assign n202 = ~n200 & ~n201;
  assign n203 = pi100  & ~n202;
  assign n204 = ~n199 & ~n203;
  assign n205 = ~pi98  & ~n204;
  assign n206 = ~pi99  & ~n202;
  assign n207 = pi99  & ~n204;
  assign n208 = ~n206 & ~n207;
  assign n209 = pi98  & ~n208;
  assign n210 = ~n205 & ~n209;
  assign n211 = ~pi96  & ~n210;
  assign n212 = ~pi97  & ~n208;
  assign n213 = pi97  & ~n210;
  assign n214 = ~n212 & ~n213;
  assign n215 = pi96  & ~n214;
  assign n216 = ~n211 & ~n215;
  assign n217 = ~pi94  & ~n216;
  assign n218 = ~pi95  & ~n214;
  assign n219 = pi95  & ~n216;
  assign n220 = ~n218 & ~n219;
  assign n221 = pi94  & ~n220;
  assign n222 = ~n217 & ~n221;
  assign n223 = ~pi92  & ~n222;
  assign n224 = ~pi93  & ~n220;
  assign n225 = pi93  & ~n222;
  assign n226 = ~n224 & ~n225;
  assign n227 = pi92  & ~n226;
  assign n228 = ~n223 & ~n227;
  assign n229 = ~pi90  & ~n228;
  assign n230 = ~pi91  & ~n226;
  assign n231 = pi91  & ~n228;
  assign n232 = ~n230 & ~n231;
  assign n233 = pi90  & ~n232;
  assign n234 = ~n229 & ~n233;
  assign n235 = ~pi88  & ~n234;
  assign n236 = ~pi89  & ~n232;
  assign n237 = pi89  & ~n234;
  assign n238 = ~n236 & ~n237;
  assign n239 = pi88  & ~n238;
  assign n240 = ~n235 & ~n239;
  assign n241 = ~pi86  & ~n240;
  assign n242 = ~pi87  & ~n238;
  assign n243 = pi87  & ~n240;
  assign n244 = ~n242 & ~n243;
  assign n245 = pi86  & ~n244;
  assign n246 = ~n241 & ~n245;
  assign n247 = ~pi84  & ~n246;
  assign n248 = ~pi85  & ~n244;
  assign n249 = pi85  & ~n246;
  assign n250 = ~n248 & ~n249;
  assign n251 = pi84  & ~n250;
  assign n252 = ~n247 & ~n251;
  assign n253 = ~pi82  & ~n252;
  assign n254 = ~pi83  & ~n250;
  assign n255 = pi83  & ~n252;
  assign n256 = ~n254 & ~n255;
  assign n257 = pi82  & ~n256;
  assign n258 = ~n253 & ~n257;
  assign n259 = ~pi80  & ~n258;
  assign n260 = ~pi81  & ~n256;
  assign n261 = pi81  & ~n258;
  assign n262 = ~n260 & ~n261;
  assign n263 = pi80  & ~n262;
  assign n264 = ~n259 & ~n263;
  assign n265 = ~pi78  & ~n264;
  assign n266 = ~pi79  & ~n262;
  assign n267 = pi79  & ~n264;
  assign n268 = ~n266 & ~n267;
  assign n269 = pi78  & ~n268;
  assign n270 = ~n265 & ~n269;
  assign n271 = ~pi76  & ~n270;
  assign n272 = ~pi77  & ~n268;
  assign n273 = pi77  & ~n270;
  assign n274 = ~n272 & ~n273;
  assign n275 = pi76  & ~n274;
  assign n276 = ~n271 & ~n275;
  assign n277 = ~pi74  & ~n276;
  assign n278 = ~pi75  & ~n274;
  assign n279 = pi75  & ~n276;
  assign n280 = ~n278 & ~n279;
  assign n281 = pi74  & ~n280;
  assign n282 = ~n277 & ~n281;
  assign n283 = ~pi72  & ~n282;
  assign n284 = ~pi73  & ~n280;
  assign n285 = pi73  & ~n282;
  assign n286 = ~n284 & ~n285;
  assign n287 = pi72  & ~n286;
  assign n288 = ~n283 & ~n287;
  assign n289 = ~pi70  & ~n288;
  assign n290 = ~pi71  & ~n286;
  assign n291 = pi71  & ~n288;
  assign n292 = ~n290 & ~n291;
  assign n293 = pi70  & ~n292;
  assign n294 = ~n289 & ~n293;
  assign n295 = ~pi68  & ~n294;
  assign n296 = ~pi69  & ~n292;
  assign n297 = pi69  & ~n294;
  assign n298 = ~n296 & ~n297;
  assign n299 = pi68  & ~n298;
  assign n300 = ~n295 & ~n299;
  assign n301 = ~pi66  & ~n300;
  assign n302 = ~pi67  & ~n298;
  assign n303 = pi67  & ~n300;
  assign n304 = ~n302 & ~n303;
  assign n305 = pi66  & ~n304;
  assign n306 = ~n301 & ~n305;
  assign n307 = ~pi64  & ~n306;
  assign n308 = ~pi65  & ~n304;
  assign n309 = pi65  & ~n306;
  assign n310 = ~n308 & ~n309;
  assign n311 = pi64  & ~n310;
  assign n312 = ~n307 & ~n311;
  assign n313 = ~pi62  & ~n312;
  assign n314 = ~pi63  & ~n310;
  assign n315 = pi63  & ~n312;
  assign n316 = ~n314 & ~n315;
  assign n317 = pi62  & ~n316;
  assign n318 = ~n313 & ~n317;
  assign n319 = ~pi60  & ~n318;
  assign n320 = ~pi61  & ~n316;
  assign n321 = pi61  & ~n318;
  assign n322 = ~n320 & ~n321;
  assign n323 = pi60  & ~n322;
  assign n324 = ~n319 & ~n323;
  assign n325 = ~pi58  & ~n324;
  assign n326 = ~pi59  & ~n322;
  assign n327 = pi59  & ~n324;
  assign n328 = ~n326 & ~n327;
  assign n329 = pi58  & ~n328;
  assign n330 = ~n325 & ~n329;
  assign n331 = ~pi56  & ~n330;
  assign n332 = ~pi57  & ~n328;
  assign n333 = pi57  & ~n330;
  assign n334 = ~n332 & ~n333;
  assign n335 = pi56  & ~n334;
  assign n336 = ~n331 & ~n335;
  assign n337 = ~pi54  & ~n336;
  assign n338 = ~pi55  & ~n334;
  assign n339 = pi55  & ~n336;
  assign n340 = ~n338 & ~n339;
  assign n341 = pi54  & ~n340;
  assign n342 = ~n337 & ~n341;
  assign n343 = ~pi52  & ~n342;
  assign n344 = ~pi53  & ~n340;
  assign n345 = pi53  & ~n342;
  assign n346 = ~n344 & ~n345;
  assign n347 = pi52  & ~n346;
  assign n348 = ~n343 & ~n347;
  assign n349 = ~pi50  & ~n348;
  assign n350 = ~pi51  & ~n346;
  assign n351 = pi51  & ~n348;
  assign n352 = ~n350 & ~n351;
  assign n353 = pi50  & ~n352;
  assign n354 = ~n349 & ~n353;
  assign n355 = ~pi48  & ~n354;
  assign n356 = ~pi49  & ~n352;
  assign n357 = pi49  & ~n354;
  assign n358 = ~n356 & ~n357;
  assign n359 = pi48  & ~n358;
  assign n360 = ~n355 & ~n359;
  assign n361 = ~pi46  & ~n360;
  assign n362 = ~pi47  & ~n358;
  assign n363 = pi47  & ~n360;
  assign n364 = ~n362 & ~n363;
  assign n365 = pi46  & ~n364;
  assign n366 = ~n361 & ~n365;
  assign n367 = ~pi44  & ~n366;
  assign n368 = ~pi45  & ~n364;
  assign n369 = pi45  & ~n366;
  assign n370 = ~n368 & ~n369;
  assign n371 = pi44  & ~n370;
  assign n372 = ~n367 & ~n371;
  assign n373 = ~pi42  & ~n372;
  assign n374 = ~pi43  & ~n370;
  assign n375 = pi43  & ~n372;
  assign n376 = ~n374 & ~n375;
  assign n377 = pi42  & ~n376;
  assign n378 = ~n373 & ~n377;
  assign n379 = ~pi40  & ~n378;
  assign n380 = ~pi41  & ~n376;
  assign n381 = pi41  & ~n378;
  assign n382 = ~n380 & ~n381;
  assign n383 = pi40  & ~n382;
  assign n384 = ~n379 & ~n383;
  assign n385 = ~pi38  & ~n384;
  assign n386 = ~pi39  & ~n382;
  assign n387 = pi39  & ~n384;
  assign n388 = ~n386 & ~n387;
  assign n389 = pi38  & ~n388;
  assign n390 = ~n385 & ~n389;
  assign n391 = ~pi36  & ~n390;
  assign n392 = ~pi37  & ~n388;
  assign n393 = pi37  & ~n390;
  assign n394 = ~n392 & ~n393;
  assign n395 = pi36  & ~n394;
  assign n396 = ~n391 & ~n395;
  assign n397 = ~pi34  & ~n396;
  assign n398 = ~pi35  & ~n394;
  assign n399 = pi35  & ~n396;
  assign n400 = ~n398 & ~n399;
  assign n401 = pi34  & ~n400;
  assign n402 = ~n397 & ~n401;
  assign n403 = ~pi32  & ~n402;
  assign n404 = ~pi33  & ~n400;
  assign n405 = pi33  & ~n402;
  assign n406 = ~n404 & ~n405;
  assign n407 = pi32  & ~n406;
  assign n408 = ~n403 & ~n407;
  assign n409 = ~pi30  & ~n408;
  assign n410 = ~pi31  & ~n406;
  assign n411 = pi31  & ~n408;
  assign n412 = ~n410 & ~n411;
  assign n413 = pi30  & ~n412;
  assign n414 = ~n409 & ~n413;
  assign n415 = ~pi28  & ~n414;
  assign n416 = ~pi29  & ~n412;
  assign n417 = pi29  & ~n414;
  assign n418 = ~n416 & ~n417;
  assign n419 = pi28  & ~n418;
  assign n420 = ~n415 & ~n419;
  assign n421 = ~pi26  & ~n420;
  assign n422 = ~pi27  & ~n418;
  assign n423 = pi27  & ~n420;
  assign n424 = ~n422 & ~n423;
  assign n425 = pi26  & ~n424;
  assign n426 = ~n421 & ~n425;
  assign n427 = ~pi24  & ~n426;
  assign n428 = ~pi25  & ~n424;
  assign n429 = pi25  & ~n426;
  assign n430 = ~n428 & ~n429;
  assign n431 = pi24  & ~n430;
  assign n432 = ~n427 & ~n431;
  assign n433 = ~pi22  & ~n432;
  assign n434 = ~pi23  & ~n430;
  assign n435 = pi23  & ~n432;
  assign n436 = ~n434 & ~n435;
  assign n437 = pi22  & ~n436;
  assign n438 = ~n433 & ~n437;
  assign n439 = ~pi20  & ~n438;
  assign n440 = ~pi21  & ~n436;
  assign n441 = pi21  & ~n438;
  assign n442 = ~n440 & ~n441;
  assign n443 = pi20  & ~n442;
  assign n444 = ~n439 & ~n443;
  assign n445 = ~pi18  & ~n444;
  assign n446 = ~pi19  & ~n442;
  assign n447 = pi19  & ~n444;
  assign n448 = ~n446 & ~n447;
  assign n449 = pi18  & ~n448;
  assign n450 = ~n445 & ~n449;
  assign n451 = ~pi16  & ~n450;
  assign n452 = ~pi17  & ~n448;
  assign n453 = pi17  & ~n450;
  assign n454 = ~n452 & ~n453;
  assign n455 = pi16  & ~n454;
  assign n456 = ~n451 & ~n455;
  assign n457 = ~pi14  & n456;
  assign n458 = ~pi15  & ~n454;
  assign n459 = pi15  & ~n456;
  assign n460 = ~n458 & ~n459;
  assign n461 = pi14  & n460;
  assign n462 = ~pi121  & ~n148;
  assign n463 = ~n457 & n462;
  assign n464 = ~n461 & n463;
  assign n465 = ~pi121  & n148;
  assign n466 = ~n460 & n465;
  assign n467 = ~pi122  & ~n466;
  assign n468 = ~n464 & n467;
  assign n469 = ~pi123  & ~n468;
  assign n470 = ~pi124  & ~n469;
  assign n471 = ~pi125  & ~n470;
  assign n472 = ~pi126  & ~n471;
  assign po0  = pi127  | n472;
  assign n474 = ~pi126  & ~pi127 ;
  assign n475 = ~pi124  & ~pi125 ;
  assign n476 = ~pi122  & ~pi123 ;
  assign n477 = ~pi120  & ~pi121 ;
  assign n478 = ~pi118  & ~pi119 ;
  assign n479 = ~pi116  & ~pi117 ;
  assign n480 = ~pi24  & ~pi25 ;
  assign n481 = ~pi22  & ~pi23 ;
  assign n482 = ~pi20  & ~pi21 ;
  assign n483 = ~pi18  & ~pi19 ;
  assign n484 = ~pi16  & ~pi17 ;
  assign n485 = ~pi14  & ~pi15 ;
  assign n486 = ~pi12  & ~pi13 ;
  assign n487 = ~pi10  & ~pi11 ;
  assign n488 = ~pi8  & ~pi9 ;
  assign n489 = ~pi6  & ~pi7 ;
  assign n490 = ~pi4  & ~pi5 ;
  assign n491 = ~pi2  & ~pi3 ;
  assign n492 = n490 & ~n491;
  assign n493 = n489 & ~n492;
  assign n494 = n488 & ~n493;
  assign n495 = n487 & ~n494;
  assign n496 = n486 & ~n495;
  assign n497 = n485 & ~n496;
  assign n498 = n484 & ~n497;
  assign n499 = n483 & ~n498;
  assign n500 = n482 & ~n499;
  assign n501 = n481 & ~n500;
  assign n502 = n480 & ~n501;
  assign n503 = ~pi26  & ~pi27 ;
  assign n504 = ~pi30  & ~pi31 ;
  assign n505 = ~pi32  & ~pi33 ;
  assign n506 = ~pi34  & ~pi35 ;
  assign n507 = ~pi36  & ~pi37 ;
  assign n508 = ~pi38  & ~pi39 ;
  assign n509 = ~pi40  & ~pi41 ;
  assign n510 = ~pi42  & ~pi43 ;
  assign n511 = ~pi44  & ~pi45 ;
  assign n512 = ~pi46  & ~pi47 ;
  assign n513 = ~pi48  & ~pi49 ;
  assign n514 = ~pi50  & ~pi51 ;
  assign n515 = ~pi52  & ~pi53 ;
  assign n516 = ~pi54  & ~pi55 ;
  assign n517 = ~pi56  & ~pi57 ;
  assign n518 = ~pi58  & ~pi59 ;
  assign n519 = ~pi60  & ~pi61 ;
  assign n520 = ~pi62  & ~pi63 ;
  assign n521 = ~pi64  & ~pi65 ;
  assign n522 = ~pi66  & ~pi67 ;
  assign n523 = ~pi68  & ~pi69 ;
  assign n524 = ~pi70  & ~pi71 ;
  assign n525 = ~pi72  & ~pi73 ;
  assign n526 = ~pi74  & ~pi75 ;
  assign n527 = ~pi76  & ~pi77 ;
  assign n528 = ~pi78  & ~pi79 ;
  assign n529 = ~pi80  & ~pi81 ;
  assign n530 = ~pi82  & ~pi83 ;
  assign n531 = ~pi84  & ~pi85 ;
  assign n532 = ~pi86  & ~pi87 ;
  assign n533 = ~pi88  & ~pi89 ;
  assign n534 = ~pi90  & ~pi91 ;
  assign n535 = ~pi92  & ~pi93 ;
  assign n536 = ~pi94  & ~pi95 ;
  assign n537 = ~pi96  & ~pi97 ;
  assign n538 = ~pi98  & ~pi99 ;
  assign n539 = ~pi102  & ~pi103 ;
  assign n540 = ~pi112  & ~pi113 ;
  assign n541 = ~pi110  & ~pi111 ;
  assign n542 = ~pi106  & ~pi107 ;
  assign n543 = ~pi108  & ~pi109 ;
  assign n544 = ~n542 & n543;
  assign n545 = n541 & ~n544;
  assign n546 = n540 & ~n545;
  assign n547 = n539 & ~n546;
  assign n548 = ~pi104  & ~pi105 ;
  assign n549 = n545 & ~n548;
  assign n550 = n541 & ~n543;
  assign n551 = n548 & n550;
  assign n552 = n540 & ~n551;
  assign n553 = ~n549 & n552;
  assign n554 = ~n539 & ~n553;
  assign n555 = ~n547 & ~n554;
  assign n556 = ~pi100  & ~pi101 ;
  assign n557 = n555 & ~n556;
  assign n558 = n553 & n556;
  assign n559 = ~n557 & ~n558;
  assign n560 = ~n538 & ~n559;
  assign n561 = n538 & n555;
  assign n562 = ~n560 & ~n561;
  assign n563 = ~n537 & ~n562;
  assign n564 = n537 & ~n559;
  assign n565 = ~n563 & ~n564;
  assign n566 = ~n536 & ~n565;
  assign n567 = n536 & ~n562;
  assign n568 = ~n566 & ~n567;
  assign n569 = ~n535 & ~n568;
  assign n570 = n535 & ~n565;
  assign n571 = ~n569 & ~n570;
  assign n572 = ~n534 & ~n571;
  assign n573 = n534 & ~n568;
  assign n574 = ~n572 & ~n573;
  assign n575 = ~n533 & ~n574;
  assign n576 = n533 & ~n571;
  assign n577 = ~n575 & ~n576;
  assign n578 = ~n532 & ~n577;
  assign n579 = n532 & ~n574;
  assign n580 = ~n578 & ~n579;
  assign n581 = ~n531 & ~n580;
  assign n582 = n531 & ~n577;
  assign n583 = ~n581 & ~n582;
  assign n584 = ~n530 & ~n583;
  assign n585 = n530 & ~n580;
  assign n586 = ~n584 & ~n585;
  assign n587 = ~n529 & ~n586;
  assign n588 = n529 & ~n583;
  assign n589 = ~n587 & ~n588;
  assign n590 = ~n528 & ~n589;
  assign n591 = n528 & ~n586;
  assign n592 = ~n590 & ~n591;
  assign n593 = ~n527 & ~n592;
  assign n594 = n527 & ~n589;
  assign n595 = ~n593 & ~n594;
  assign n596 = ~n526 & ~n595;
  assign n597 = n526 & ~n592;
  assign n598 = ~n596 & ~n597;
  assign n599 = ~n525 & ~n598;
  assign n600 = n525 & ~n595;
  assign n601 = ~n599 & ~n600;
  assign n602 = ~n524 & ~n601;
  assign n603 = n524 & ~n598;
  assign n604 = ~n602 & ~n603;
  assign n605 = ~n523 & ~n604;
  assign n606 = n523 & ~n601;
  assign n607 = ~n605 & ~n606;
  assign n608 = ~n522 & ~n607;
  assign n609 = n522 & ~n604;
  assign n610 = ~n608 & ~n609;
  assign n611 = ~n521 & ~n610;
  assign n612 = n521 & ~n607;
  assign n613 = ~n611 & ~n612;
  assign n614 = ~n520 & ~n613;
  assign n615 = n520 & ~n610;
  assign n616 = ~n614 & ~n615;
  assign n617 = ~n519 & ~n616;
  assign n618 = n519 & ~n613;
  assign n619 = ~n617 & ~n618;
  assign n620 = ~n518 & ~n619;
  assign n621 = n518 & ~n616;
  assign n622 = ~n620 & ~n621;
  assign n623 = ~n517 & ~n622;
  assign n624 = n517 & ~n619;
  assign n625 = ~n623 & ~n624;
  assign n626 = ~n516 & ~n625;
  assign n627 = n516 & ~n622;
  assign n628 = ~n626 & ~n627;
  assign n629 = ~n515 & ~n628;
  assign n630 = n515 & ~n625;
  assign n631 = ~n629 & ~n630;
  assign n632 = ~n514 & ~n631;
  assign n633 = n514 & ~n628;
  assign n634 = ~n632 & ~n633;
  assign n635 = ~n513 & ~n634;
  assign n636 = n513 & ~n631;
  assign n637 = ~n635 & ~n636;
  assign n638 = ~n512 & ~n637;
  assign n639 = n512 & ~n634;
  assign n640 = ~n638 & ~n639;
  assign n641 = ~n511 & ~n640;
  assign n642 = n511 & ~n637;
  assign n643 = ~n641 & ~n642;
  assign n644 = ~n510 & ~n643;
  assign n645 = n510 & ~n640;
  assign n646 = ~n644 & ~n645;
  assign n647 = ~n509 & ~n646;
  assign n648 = n509 & ~n643;
  assign n649 = ~n647 & ~n648;
  assign n650 = ~n508 & ~n649;
  assign n651 = n508 & ~n646;
  assign n652 = ~n650 & ~n651;
  assign n653 = ~n507 & ~n652;
  assign n654 = n507 & ~n649;
  assign n655 = ~n653 & ~n654;
  assign n656 = ~n506 & ~n655;
  assign n657 = n506 & ~n652;
  assign n658 = ~n656 & ~n657;
  assign n659 = ~n505 & ~n658;
  assign n660 = n505 & ~n655;
  assign n661 = ~n659 & ~n660;
  assign n662 = ~n504 & ~n661;
  assign n663 = n504 & ~n658;
  assign n664 = ~n662 & ~n663;
  assign n665 = n503 & ~n664;
  assign n666 = ~pi114  & ~pi115 ;
  assign n667 = ~pi28  & ~pi29 ;
  assign n668 = ~n664 & ~n667;
  assign n669 = ~n661 & n667;
  assign n670 = ~n668 & ~n669;
  assign n671 = ~n503 & ~n670;
  assign n672 = ~n502 & n666;
  assign n673 = ~n665 & n672;
  assign n674 = ~n671 & n673;
  assign n675 = n502 & n666;
  assign n676 = n670 & n675;
  assign n677 = n479 & ~n676;
  assign n678 = ~n674 & n677;
  assign n679 = n478 & ~n678;
  assign n680 = n477 & ~n679;
  assign n681 = n476 & ~n680;
  assign n682 = n475 & ~n681;
  assign po1  = ~n474 | n682;
  assign n684 = n474 & n475;
  assign n685 = n476 & n477;
  assign n686 = n478 & n479;
  assign n687 = n540 & n666;
  assign n688 = n531 & n532;
  assign n689 = n542 & n548;
  assign n690 = n533 & n534;
  assign n691 = n539 & n556;
  assign n692 = n537 & n538;
  assign n693 = n535 & n536;
  assign n694 = n692 & ~n693;
  assign n695 = n691 & ~n694;
  assign n696 = ~n690 & n695;
  assign n697 = n690 & n691;
  assign n698 = ~n692 & n697;
  assign n699 = n689 & ~n698;
  assign n700 = ~n696 & n699;
  assign n701 = ~n688 & n700;
  assign n702 = n541 & n543;
  assign n703 = n688 & n689;
  assign n704 = ~n695 & n703;
  assign n705 = n702 & ~n704;
  assign n706 = ~n701 & n705;
  assign n707 = n687 & ~n706;
  assign n708 = n686 & ~n707;
  assign n709 = n685 & ~n708;
  assign n710 = n529 & n530;
  assign n711 = n709 & ~n710;
  assign n712 = ~n700 & n702;
  assign n713 = n687 & ~n712;
  assign n714 = n686 & ~n713;
  assign n715 = n685 & n710;
  assign n716 = ~n714 & n715;
  assign n717 = n527 & n528;
  assign n718 = n525 & n526;
  assign n719 = n523 & n524;
  assign n720 = n521 & n522;
  assign n721 = n519 & n520;
  assign n722 = n517 & n518;
  assign n723 = n515 & n516;
  assign n724 = n513 & n514;
  assign n725 = n511 & n512;
  assign n726 = n509 & n510;
  assign n727 = n507 & n508;
  assign n728 = n505 & n506;
  assign n729 = n504 & n667;
  assign n730 = n480 & n503;
  assign n731 = n481 & n482;
  assign n732 = n483 & n484;
  assign n733 = n485 & n486;
  assign n734 = n487 & n488;
  assign n735 = n489 & n490;
  assign n736 = n734 & ~n735;
  assign n737 = n733 & ~n736;
  assign n738 = n732 & ~n737;
  assign n739 = n731 & ~n738;
  assign n740 = n730 & ~n739;
  assign n741 = n729 & ~n740;
  assign n742 = n728 & ~n741;
  assign n743 = n727 & ~n742;
  assign n744 = n726 & ~n743;
  assign n745 = n725 & ~n744;
  assign n746 = n724 & ~n745;
  assign n747 = n723 & ~n746;
  assign n748 = n722 & ~n747;
  assign n749 = n721 & ~n748;
  assign n750 = n720 & ~n749;
  assign n751 = n719 & ~n750;
  assign n752 = n718 & ~n751;
  assign n753 = n717 & ~n752;
  assign n754 = n684 & ~n716;
  assign n755 = ~n711 & n754;
  assign n756 = ~n753 & n755;
  assign n757 = n684 & n717;
  assign n758 = ~n709 & n757;
  assign n759 = ~n752 & n758;
  assign po2  = ~n756 & ~n759;
  assign n761 = n684 & n685;
  assign n762 = n688 & n710;
  assign n763 = n717 & n718;
  assign n764 = n719 & n720;
  assign n765 = n721 & n722;
  assign n766 = n723 & n724;
  assign n767 = n725 & n726;
  assign n768 = n727 & n728;
  assign n769 = n729 & n730;
  assign n770 = n731 & n732;
  assign n771 = n733 & n734;
  assign n772 = n770 & ~n771;
  assign n773 = n769 & ~n772;
  assign n774 = n768 & ~n773;
  assign n775 = n767 & ~n774;
  assign n776 = n766 & ~n775;
  assign n777 = n765 & ~n776;
  assign n778 = n764 & ~n777;
  assign n779 = n763 & ~n778;
  assign n780 = n762 & ~n779;
  assign n781 = n686 & n687;
  assign n782 = n689 & n702;
  assign n783 = n690 & n693;
  assign n784 = n691 & n692;
  assign n785 = ~n783 & n784;
  assign n786 = n782 & ~n785;
  assign n787 = n781 & ~n786;
  assign n788 = ~n780 & n787;
  assign n789 = n782 & ~n784;
  assign n790 = n781 & ~n789;
  assign n791 = n780 & n790;
  assign n792 = n761 & ~n788;
  assign po3  = n791 | ~n792;
  assign n794 = n761 & n781;
  assign n795 = n782 & n784;
  assign n796 = n762 & n783;
  assign n797 = n765 & n766;
  assign n798 = n769 & n770;
  assign n799 = n767 & n768;
  assign n800 = ~n798 & n799;
  assign n801 = n797 & ~n800;
  assign n802 = n763 & n764;
  assign n803 = ~n801 & n802;
  assign n804 = n796 & ~n803;
  assign n805 = n795 & ~n804;
  assign po4  = ~n794 | n805;
  assign n807 = n794 & n795;
  assign n808 = n796 & n802;
  assign n809 = n797 & n799;
  assign n810 = n808 & ~n809;
  assign po5  = ~n807 | n810;
  assign po6  = ~n807 | ~n808;
  assign n813 = ~pi0  & ~pi1 ;
  assign n814 = n491 & n813;
  assign n815 = n735 & n814;
  assign n816 = n771 & n815;
  assign n817 = n798 & n816;
  assign n818 = n809 & n817;
  assign po7 = po6  | ~n818;
endmodule
