module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 , pi32 ,
    pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 , pi40 ,
    pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 , pi56 ,
    pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 , pi64 ,
    pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 ,
    pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 ,
    pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 ,
    pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 ,
    pi97 , pi98 , pi99 , pi100 , pi101 , pi102 , pi103 ,
    pi104 , pi105 , pi106 , pi107 , pi108 , pi109 , pi110 ,
    pi111 , pi112 , pi113 , pi114 , pi115 , pi116 , pi117 ,
    pi118 , pi119 , pi120 , pi121 , pi122 , pi123 , pi124 ,
    pi125 , pi126 , pi127 , pi128 , pi129 , pi130 , pi131 , pi132 ,
    pi133 , pi134 , pi135 , pi136 , pi137 , pi138 , pi139 , pi140 ,
    pi141 , pi142 , pi143 , pi144 , pi145 , pi146 , pi147 , pi148 ,
    pi149 , pi150 , pi151 , pi152 , pi153 , pi154 , pi155 , pi156 ,
    pi157 , pi158 , pi159 , pi160 , pi161 , pi162 , pi163 , pi164 ,
    pi165 , pi166 , pi167 , pi168 , pi169 , pi170 , pi171 , pi172 ,
    pi173 , pi174 , pi175 , pi176 , pi177 , pi178 , pi179 , pi180 ,
    pi181 , pi182 , pi183 , pi184 , pi185 , pi186 , pi187 , pi188 ,
    pi189 , pi190 , pi191 , pi192 , pi193 , pi194 , pi195 , pi196 ,
    pi197 , pi198 , pi199 , pi200 , pi201 , pi202 , pi203 , pi204 ,
    pi205 , pi206 , pi207 , pi208 , pi209 , pi210 , pi211 , pi212 ,
    pi213 , pi214 , pi215 , pi216 , pi217 , pi218 , pi219 , pi220 ,
    pi221 , pi222 , pi223 , pi224 , pi225 , pi226 , pi227 ,
    pi228 , pi229 , pi230 , pi231 , pi232 , pi233 , pi234 ,
    pi235 , pi236 , pi237 , pi238 , pi239 , pi240 , pi241 ,
    pi242 , pi243 , pi244 , pi245 , pi246 , pi247 , pi248 ,
    pi249 , pi250 , pi251 , pi252 , pi253 , pi254 , pi255 ,
    po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7 , po8 ,
    po9 , po10 , po11 , po12 , po13 , po14 , po15 , po16 ,
    po17 , po18 , po19 , po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 , po30 , po31 , po32 ,
    po33 , po34 , po35 , po36 , po37 , po38 , po39 , po40 ,
    po41 , po42 , po43 , po44 , po45 , po46 , po47 , po48 ,
    po49 , po50 , po51 , po52 , po53 , po54 , po55 , po56 ,
    po57 , po58 , po59 , po60 , po61 , po62 , po63 , po64 ,
    po65 , po66 , po67 , po68 , po69 , po70 , po71 , po72 ,
    po73 , po74 , po75 , po76 , po77 , po78 , po79 , po80 ,
    po81 , po82 , po83 , po84 , po85 , po86 , po87 , po88 ,
    po89 , po90 , po91 , po92 , po93 , po94 , po95 , po96 ,
    po97 , po98 , po99 , po100 , po101 , po102 , po103 ,
    po104 , po105 , po106 , po107 , po108 , po109 , po110 ,
    po111 , po112 , po113 , po114 , po115 , po116 , po117 ,
    po118 , po119 , po120 , po121 , po122 , po123 , po124 ,
    po125 , po126 , po127 , po128  );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    pi32 , pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 ,
    pi56 , pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 ,
    pi64 , pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 ,
    pi72 , pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 ,
    pi80 , pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 ,
    pi88 , pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 ,
    pi96 , pi97 , pi98 , pi99 , pi100 , pi101 , pi102 ,
    pi103 , pi104 , pi105 , pi106 , pi107 , pi108 , pi109 ,
    pi110 , pi111 , pi112 , pi113 , pi114 , pi115 , pi116 ,
    pi117 , pi118 , pi119 , pi120 , pi121 , pi122 , pi123 ,
    pi124 , pi125 , pi126 , pi127 , pi128 , pi129 , pi130 , pi131 ,
    pi132 , pi133 , pi134 , pi135 , pi136 , pi137 , pi138 , pi139 ,
    pi140 , pi141 , pi142 , pi143 , pi144 , pi145 , pi146 , pi147 ,
    pi148 , pi149 , pi150 , pi151 , pi152 , pi153 , pi154 , pi155 ,
    pi156 , pi157 , pi158 , pi159 , pi160 , pi161 , pi162 , pi163 ,
    pi164 , pi165 , pi166 , pi167 , pi168 , pi169 , pi170 , pi171 ,
    pi172 , pi173 , pi174 , pi175 , pi176 , pi177 , pi178 , pi179 ,
    pi180 , pi181 , pi182 , pi183 , pi184 , pi185 , pi186 , pi187 ,
    pi188 , pi189 , pi190 , pi191 , pi192 , pi193 , pi194 , pi195 ,
    pi196 , pi197 , pi198 , pi199 , pi200 , pi201 , pi202 , pi203 ,
    pi204 , pi205 , pi206 , pi207 , pi208 , pi209 , pi210 , pi211 ,
    pi212 , pi213 , pi214 , pi215 , pi216 , pi217 , pi218 , pi219 ,
    pi220 , pi221 , pi222 , pi223 , pi224 , pi225 , pi226 , pi227 ,
    pi228 , pi229 , pi230 , pi231 , pi232 , pi233 , pi234 ,
    pi235 , pi236 , pi237 , pi238 , pi239 , pi240 , pi241 ,
    pi242 , pi243 , pi244 , pi245 , pi246 , pi247 , pi248 ,
    pi249 , pi250 , pi251 , pi252 , pi253 , pi254 , pi255 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7 ,
    po8 , po9 , po10 , po11 , po12 , po13 , po14 , po15 ,
    po16 , po17 , po18 , po19 , po20 , po21 , po22 , po23 ,
    po24 , po25 , po26 , po27 , po28 , po29 , po30 , po31 ,
    po32 , po33 , po34 , po35 , po36 , po37 , po38 , po39 ,
    po40 , po41 , po42 , po43 , po44 , po45 , po46 , po47 ,
    po48 , po49 , po50 , po51 , po52 , po53 , po54 , po55 ,
    po56 , po57 , po58 , po59 , po60 , po61 , po62 , po63 ,
    po64 , po65 , po66 , po67 , po68 , po69 , po70 , po71 ,
    po72 , po73 , po74 , po75 , po76 , po77 , po78 , po79 ,
    po80 , po81 , po82 , po83 , po84 , po85 , po86 , po87 ,
    po88 , po89 , po90 , po91 , po92 , po93 , po94 , po95 ,
    po96 , po97 , po98 , po99 , po100 , po101 , po102 ,
    po103 , po104 , po105 , po106 , po107 , po108 , po109 ,
    po110 , po111 , po112 , po113 , po114 , po115 , po116 ,
    po117 , po118 , po119 , po120 , po121 , po122 , po123 ,
    po124 , po125 , po126 , po127 , po128;
  wire n386, n387, n389, n390, n391, n392, n393,
    n395, n396, n397, n398, n399, n400, n401,
    n403, n404, n405, n406, n407, n408, n409,
    n411, n412, n413, n414, n415, n416, n417,
    n419, n420, n421, n422, n423, n424, n425,
    n427, n428, n429, n430, n431, n432, n433,
    n435, n436, n437, n438, n439, n440, n441,
    n443, n444, n445, n446, n447, n448, n449,
    n451, n452, n453, n454, n455, n456, n457,
    n459, n460, n461, n462, n463, n464, n465,
    n467, n468, n469, n470, n471, n472, n473,
    n475, n476, n477, n478, n479, n480, n481,
    n483, n484, n485, n486, n487, n488, n489,
    n491, n492, n493, n494, n495, n496, n497,
    n499, n500, n501, n502, n503, n504, n505,
    n507, n508, n509, n510, n511, n512, n513,
    n515, n516, n517, n518, n519, n520, n521,
    n523, n524, n525, n526, n527, n528, n529,
    n531, n532, n533, n534, n535, n536, n537,
    n539, n540, n541, n542, n543, n544, n545,
    n547, n548, n549, n550, n551, n552, n553,
    n555, n556, n557, n558, n559, n560, n561,
    n563, n564, n565, n566, n567, n568, n569,
    n571, n572, n573, n574, n575, n576, n577,
    n579, n580, n581, n582, n583, n584, n585,
    n587, n588, n589, n590, n591, n592, n593,
    n595, n596, n597, n598, n599, n600, n601,
    n603, n604, n605, n606, n607, n608, n609,
    n611, n612, n613, n614, n615, n616, n617,
    n619, n620, n621, n622, n623, n624, n625,
    n627, n628, n629, n630, n631, n632, n633,
    n635, n636, n637, n638, n639, n640, n641,
    n643, n644, n645, n646, n647, n648, n649,
    n651, n652, n653, n654, n655, n656, n657,
    n659, n660, n661, n662, n663, n664, n665,
    n667, n668, n669, n670, n671, n672, n673,
    n675, n676, n677, n678, n679, n680, n681,
    n683, n684, n685, n686, n687, n688, n689,
    n691, n692, n693, n694, n695, n696, n697,
    n699, n700, n701, n702, n703, n704, n705,
    n707, n708, n709, n710, n711, n712, n713,
    n715, n716, n717, n718, n719, n720, n721,
    n723, n724, n725, n726, n727, n728, n729,
    n731, n732, n733, n734, n735, n736, n737,
    n739, n740, n741, n742, n743, n744, n745,
    n747, n748, n749, n750, n751, n752, n753,
    n755, n756, n757, n758, n759, n760, n761,
    n763, n764, n765, n766, n767, n768, n769,
    n771, n772, n773, n774, n775, n776, n777,
    n779, n780, n781, n782, n783, n784, n785,
    n787, n788, n789, n790, n791, n792, n793,
    n795, n796, n797, n798, n799, n800, n801,
    n803, n804, n805, n806, n807, n808, n809,
    n811, n812, n813, n814, n815, n816, n817,
    n819, n820, n821, n822, n823, n824, n825,
    n827, n828, n829, n830, n831, n832, n833,
    n835, n836, n837, n838, n839, n840, n841,
    n843, n844, n845, n846, n847, n848, n849,
    n851, n852, n853, n854, n855, n856, n857,
    n859, n860, n861, n862, n863, n864, n865,
    n867, n868, n869, n870, n871, n872, n873,
    n875, n876, n877, n878, n879, n880, n881,
    n883, n884, n885, n886, n887, n888, n889,
    n891, n892, n893, n894, n895, n896, n897,
    n899, n900, n901, n902, n903, n904, n905,
    n907, n908, n909, n910, n911, n912, n913,
    n915, n916, n917, n918, n919, n920, n921,
    n923, n924, n925, n926, n927, n928, n929,
    n931, n932, n933, n934, n935, n936, n937,
    n939, n940, n941, n942, n943, n944, n945,
    n947, n948, n949, n950, n951, n952, n953,
    n955, n956, n957, n958, n959, n960, n961,
    n963, n964, n965, n966, n967, n968, n969,
    n971, n972, n973, n974, n975, n976, n977,
    n979, n980, n981, n982, n983, n984, n985,
    n987, n988, n989, n990, n991, n992, n993,
    n995, n996, n997, n998, n999, n1000, n1001,
    n1003, n1004, n1005, n1006, n1007, n1008,
    n1009, n1011, n1012, n1013, n1014, n1015,
    n1016, n1017, n1019, n1020, n1021, n1022,
    n1023, n1024, n1025, n1027, n1028, n1029,
    n1030, n1031, n1032, n1033, n1035, n1036,
    n1037, n1038, n1039, n1040, n1041, n1043,
    n1044, n1045, n1046, n1047, n1048, n1049,
    n1051, n1052, n1053, n1054, n1055, n1056,
    n1057, n1059, n1060, n1061, n1062, n1063,
    n1064, n1065, n1067, n1068, n1069, n1070,
    n1071, n1072, n1073, n1075, n1076, n1077,
    n1078, n1079, n1080, n1081, n1083, n1084,
    n1085, n1086, n1087, n1088, n1089, n1091,
    n1092, n1093, n1094, n1095, n1096, n1097,
    n1099, n1100, n1101, n1102, n1103, n1104,
    n1105, n1107, n1108, n1109, n1110, n1111,
    n1112, n1113, n1115, n1116, n1117, n1118,
    n1119, n1120, n1121, n1123, n1124, n1125,
    n1126, n1127, n1128, n1129, n1131, n1132,
    n1133, n1134, n1135, n1136, n1137, n1139,
    n1140, n1141, n1142, n1143, n1144, n1145,
    n1147, n1148, n1149, n1150, n1151, n1152,
    n1153, n1155, n1156, n1157, n1158, n1159,
    n1160, n1161, n1163, n1164, n1165, n1166,
    n1167, n1168, n1169, n1171, n1172, n1173,
    n1174, n1175, n1176, n1177, n1179, n1180,
    n1181, n1182, n1183, n1184, n1185, n1187,
    n1188, n1189, n1190, n1191, n1192, n1193,
    n1195, n1196, n1197, n1198, n1199, n1200,
    n1201, n1203, n1204, n1205, n1206, n1207,
    n1208, n1209, n1211, n1212, n1213, n1214,
    n1215, n1216, n1217, n1219, n1220, n1221,
    n1222, n1223, n1224, n1225, n1227, n1228,
    n1229, n1230, n1231, n1232, n1233, n1235,
    n1236, n1237, n1238, n1239, n1240, n1241,
    n1243, n1244, n1245, n1246, n1247, n1248,
    n1249, n1251, n1252, n1253, n1254, n1255,
    n1256, n1257, n1259, n1260, n1261, n1262,
    n1263, n1264, n1265, n1267, n1268, n1269,
    n1270, n1271, n1272, n1273, n1275, n1276,
    n1277, n1278, n1279, n1280, n1281, n1283,
    n1284, n1285, n1286, n1287, n1288, n1289,
    n1291, n1292, n1293, n1294, n1295, n1296,
    n1297, n1299, n1300, n1301, n1302, n1303,
    n1304, n1305, n1307, n1308, n1309, n1310,
    n1311, n1312, n1313, n1315, n1316, n1317,
    n1318, n1319, n1320, n1321, n1323, n1324,
    n1325, n1326, n1327, n1328, n1329, n1331,
    n1332, n1333, n1334, n1335, n1336, n1337,
    n1339, n1340, n1341, n1342, n1343, n1344,
    n1345, n1347, n1348, n1349, n1350, n1351,
    n1352, n1353, n1355, n1356, n1357, n1358,
    n1359, n1360, n1361, n1363, n1364, n1365,
    n1366, n1367, n1368, n1369, n1371, n1372,
    n1373, n1374, n1375, n1376, n1377, n1379,
    n1380, n1381, n1382, n1383, n1384, n1385,
    n1387, n1388, n1389, n1390, n1391, n1392,
    n1393, n1395, n1396, n1397, n1398, n1399,
    n1400, n1401, n1403;
  assign n386 = pi0  & pi128 ;
  assign n387 = ~pi0  & ~pi128 ;
  assign po0  = ~n386 & ~n387;
  assign n389 = ~pi1  & ~pi129 ;
  assign n390 = pi1  & pi129 ;
  assign n391 = ~n389 & ~n390;
  assign n392 = n386 & ~n391;
  assign n393 = ~n386 & n391;
  assign po1  = n392 | n393;
  assign n395 = ~pi2  & ~pi130 ;
  assign n396 = pi2  & pi130 ;
  assign n397 = ~n395 & ~n396;
  assign n398 = ~n386 & ~n390;
  assign n399 = ~n389 & ~n398;
  assign n400 = n397 & ~n399;
  assign n401 = ~n397 & n399;
  assign po2  = n400 | n401;
  assign n403 = ~pi3  & ~pi131 ;
  assign n404 = pi3  & pi131 ;
  assign n405 = ~n403 & ~n404;
  assign n406 = ~n396 & ~n399;
  assign n407 = ~n395 & ~n406;
  assign n408 = n405 & ~n407;
  assign n409 = ~n405 & n407;
  assign po3  = n408 | n409;
  assign n411 = ~pi4  & ~pi132 ;
  assign n412 = pi4  & pi132 ;
  assign n413 = ~n411 & ~n412;
  assign n414 = ~n404 & ~n407;
  assign n415 = ~n403 & ~n414;
  assign n416 = n413 & ~n415;
  assign n417 = ~n413 & n415;
  assign po4  = n416 | n417;
  assign n419 = ~pi5  & ~pi133 ;
  assign n420 = pi5  & pi133 ;
  assign n421 = ~n419 & ~n420;
  assign n422 = ~n412 & ~n415;
  assign n423 = ~n411 & ~n422;
  assign n424 = n421 & ~n423;
  assign n425 = ~n421 & n423;
  assign po5  = n424 | n425;
  assign n427 = ~pi6  & ~pi134 ;
  assign n428 = pi6  & pi134 ;
  assign n429 = ~n427 & ~n428;
  assign n430 = ~n420 & ~n423;
  assign n431 = ~n419 & ~n430;
  assign n432 = n429 & ~n431;
  assign n433 = ~n429 & n431;
  assign po6  = n432 | n433;
  assign n435 = ~pi7  & ~pi135 ;
  assign n436 = pi7  & pi135 ;
  assign n437 = ~n435 & ~n436;
  assign n438 = ~n428 & ~n431;
  assign n439 = ~n427 & ~n438;
  assign n440 = n437 & ~n439;
  assign n441 = ~n437 & n439;
  assign po7  = n440 | n441;
  assign n443 = ~pi8  & ~pi136 ;
  assign n444 = pi8  & pi136 ;
  assign n445 = ~n443 & ~n444;
  assign n446 = ~n436 & ~n439;
  assign n447 = ~n435 & ~n446;
  assign n448 = n445 & ~n447;
  assign n449 = ~n445 & n447;
  assign po8  = n448 | n449;
  assign n451 = ~pi9  & ~pi137 ;
  assign n452 = pi9  & pi137 ;
  assign n453 = ~n451 & ~n452;
  assign n454 = ~n444 & ~n447;
  assign n455 = ~n443 & ~n454;
  assign n456 = n453 & ~n455;
  assign n457 = ~n453 & n455;
  assign po9  = n456 | n457;
  assign n459 = ~pi10  & ~pi138 ;
  assign n460 = pi10  & pi138 ;
  assign n461 = ~n459 & ~n460;
  assign n462 = ~n452 & ~n455;
  assign n463 = ~n451 & ~n462;
  assign n464 = n461 & ~n463;
  assign n465 = ~n461 & n463;
  assign po10  = n464 | n465;
  assign n467 = ~pi11  & ~pi139 ;
  assign n468 = pi11  & pi139 ;
  assign n469 = ~n467 & ~n468;
  assign n470 = ~n460 & ~n463;
  assign n471 = ~n459 & ~n470;
  assign n472 = n469 & ~n471;
  assign n473 = ~n469 & n471;
  assign po11  = n472 | n473;
  assign n475 = ~pi12  & ~pi140 ;
  assign n476 = pi12  & pi140 ;
  assign n477 = ~n475 & ~n476;
  assign n478 = ~n468 & ~n471;
  assign n479 = ~n467 & ~n478;
  assign n480 = n477 & ~n479;
  assign n481 = ~n477 & n479;
  assign po12  = n480 | n481;
  assign n483 = ~pi13  & ~pi141 ;
  assign n484 = pi13  & pi141 ;
  assign n485 = ~n483 & ~n484;
  assign n486 = ~n476 & ~n479;
  assign n487 = ~n475 & ~n486;
  assign n488 = n485 & ~n487;
  assign n489 = ~n485 & n487;
  assign po13  = n488 | n489;
  assign n491 = ~pi14  & ~pi142 ;
  assign n492 = pi14  & pi142 ;
  assign n493 = ~n491 & ~n492;
  assign n494 = ~n484 & ~n487;
  assign n495 = ~n483 & ~n494;
  assign n496 = n493 & ~n495;
  assign n497 = ~n493 & n495;
  assign po14  = n496 | n497;
  assign n499 = ~pi15  & ~pi143 ;
  assign n500 = pi15  & pi143 ;
  assign n501 = ~n499 & ~n500;
  assign n502 = ~n492 & ~n495;
  assign n503 = ~n491 & ~n502;
  assign n504 = n501 & ~n503;
  assign n505 = ~n501 & n503;
  assign po15  = n504 | n505;
  assign n507 = ~pi16  & ~pi144 ;
  assign n508 = pi16  & pi144 ;
  assign n509 = ~n507 & ~n508;
  assign n510 = ~n500 & ~n503;
  assign n511 = ~n499 & ~n510;
  assign n512 = n509 & ~n511;
  assign n513 = ~n509 & n511;
  assign po16  = n512 | n513;
  assign n515 = ~pi17  & ~pi145 ;
  assign n516 = pi17  & pi145 ;
  assign n517 = ~n515 & ~n516;
  assign n518 = ~n508 & ~n511;
  assign n519 = ~n507 & ~n518;
  assign n520 = n517 & ~n519;
  assign n521 = ~n517 & n519;
  assign po17  = n520 | n521;
  assign n523 = ~pi18  & ~pi146 ;
  assign n524 = pi18  & pi146 ;
  assign n525 = ~n523 & ~n524;
  assign n526 = ~n516 & ~n519;
  assign n527 = ~n515 & ~n526;
  assign n528 = n525 & ~n527;
  assign n529 = ~n525 & n527;
  assign po18  = n528 | n529;
  assign n531 = ~pi19  & ~pi147 ;
  assign n532 = pi19  & pi147 ;
  assign n533 = ~n531 & ~n532;
  assign n534 = ~n524 & ~n527;
  assign n535 = ~n523 & ~n534;
  assign n536 = n533 & ~n535;
  assign n537 = ~n533 & n535;
  assign po19  = n536 | n537;
  assign n539 = ~pi20  & ~pi148 ;
  assign n540 = pi20  & pi148 ;
  assign n541 = ~n539 & ~n540;
  assign n542 = ~n532 & ~n535;
  assign n543 = ~n531 & ~n542;
  assign n544 = n541 & ~n543;
  assign n545 = ~n541 & n543;
  assign po20  = n544 | n545;
  assign n547 = ~pi21  & ~pi149 ;
  assign n548 = pi21  & pi149 ;
  assign n549 = ~n547 & ~n548;
  assign n550 = ~n540 & ~n543;
  assign n551 = ~n539 & ~n550;
  assign n552 = n549 & ~n551;
  assign n553 = ~n549 & n551;
  assign po21  = n552 | n553;
  assign n555 = ~pi22  & ~pi150 ;
  assign n556 = pi22  & pi150 ;
  assign n557 = ~n555 & ~n556;
  assign n558 = ~n548 & ~n551;
  assign n559 = ~n547 & ~n558;
  assign n560 = n557 & ~n559;
  assign n561 = ~n557 & n559;
  assign po22  = n560 | n561;
  assign n563 = ~pi23  & ~pi151 ;
  assign n564 = pi23  & pi151 ;
  assign n565 = ~n563 & ~n564;
  assign n566 = ~n556 & ~n559;
  assign n567 = ~n555 & ~n566;
  assign n568 = n565 & ~n567;
  assign n569 = ~n565 & n567;
  assign po23  = n568 | n569;
  assign n571 = ~pi24  & ~pi152 ;
  assign n572 = pi24  & pi152 ;
  assign n573 = ~n571 & ~n572;
  assign n574 = ~n564 & ~n567;
  assign n575 = ~n563 & ~n574;
  assign n576 = n573 & ~n575;
  assign n577 = ~n573 & n575;
  assign po24  = n576 | n577;
  assign n579 = ~pi25  & ~pi153 ;
  assign n580 = pi25  & pi153 ;
  assign n581 = ~n579 & ~n580;
  assign n582 = ~n572 & ~n575;
  assign n583 = ~n571 & ~n582;
  assign n584 = n581 & ~n583;
  assign n585 = ~n581 & n583;
  assign po25  = n584 | n585;
  assign n587 = ~pi26  & ~pi154 ;
  assign n588 = pi26  & pi154 ;
  assign n589 = ~n587 & ~n588;
  assign n590 = ~n580 & ~n583;
  assign n591 = ~n579 & ~n590;
  assign n592 = n589 & ~n591;
  assign n593 = ~n589 & n591;
  assign po26  = n592 | n593;
  assign n595 = ~pi27  & ~pi155 ;
  assign n596 = pi27  & pi155 ;
  assign n597 = ~n595 & ~n596;
  assign n598 = ~n588 & ~n591;
  assign n599 = ~n587 & ~n598;
  assign n600 = n597 & ~n599;
  assign n601 = ~n597 & n599;
  assign po27  = n600 | n601;
  assign n603 = ~pi28  & ~pi156 ;
  assign n604 = pi28  & pi156 ;
  assign n605 = ~n603 & ~n604;
  assign n606 = ~n596 & ~n599;
  assign n607 = ~n595 & ~n606;
  assign n608 = n605 & ~n607;
  assign n609 = ~n605 & n607;
  assign po28  = n608 | n609;
  assign n611 = ~pi29  & ~pi157 ;
  assign n612 = pi29  & pi157 ;
  assign n613 = ~n611 & ~n612;
  assign n614 = ~n604 & ~n607;
  assign n615 = ~n603 & ~n614;
  assign n616 = n613 & ~n615;
  assign n617 = ~n613 & n615;
  assign po29  = n616 | n617;
  assign n619 = ~pi30  & ~pi158 ;
  assign n620 = pi30  & pi158 ;
  assign n621 = ~n619 & ~n620;
  assign n622 = ~n612 & ~n615;
  assign n623 = ~n611 & ~n622;
  assign n624 = n621 & ~n623;
  assign n625 = ~n621 & n623;
  assign po30  = n624 | n625;
  assign n627 = ~pi31  & ~pi159 ;
  assign n628 = pi31  & pi159 ;
  assign n629 = ~n627 & ~n628;
  assign n630 = ~n620 & ~n623;
  assign n631 = ~n619 & ~n630;
  assign n632 = n629 & ~n631;
  assign n633 = ~n629 & n631;
  assign po31  = n632 | n633;
  assign n635 = ~pi32  & ~pi160 ;
  assign n636 = pi32  & pi160 ;
  assign n637 = ~n635 & ~n636;
  assign n638 = ~n628 & ~n631;
  assign n639 = ~n627 & ~n638;
  assign n640 = n637 & ~n639;
  assign n641 = ~n637 & n639;
  assign po32  = n640 | n641;
  assign n643 = ~pi33  & ~pi161 ;
  assign n644 = pi33  & pi161 ;
  assign n645 = ~n643 & ~n644;
  assign n646 = ~n636 & ~n639;
  assign n647 = ~n635 & ~n646;
  assign n648 = n645 & ~n647;
  assign n649 = ~n645 & n647;
  assign po33  = n648 | n649;
  assign n651 = ~pi34  & ~pi162 ;
  assign n652 = pi34  & pi162 ;
  assign n653 = ~n651 & ~n652;
  assign n654 = ~n644 & ~n647;
  assign n655 = ~n643 & ~n654;
  assign n656 = n653 & ~n655;
  assign n657 = ~n653 & n655;
  assign po34  = n656 | n657;
  assign n659 = ~pi35  & ~pi163 ;
  assign n660 = pi35  & pi163 ;
  assign n661 = ~n659 & ~n660;
  assign n662 = ~n652 & ~n655;
  assign n663 = ~n651 & ~n662;
  assign n664 = n661 & ~n663;
  assign n665 = ~n661 & n663;
  assign po35  = n664 | n665;
  assign n667 = ~pi36  & ~pi164 ;
  assign n668 = pi36  & pi164 ;
  assign n669 = ~n667 & ~n668;
  assign n670 = ~n660 & ~n663;
  assign n671 = ~n659 & ~n670;
  assign n672 = n669 & ~n671;
  assign n673 = ~n669 & n671;
  assign po36  = n672 | n673;
  assign n675 = ~pi37  & ~pi165 ;
  assign n676 = pi37  & pi165 ;
  assign n677 = ~n675 & ~n676;
  assign n678 = ~n668 & ~n671;
  assign n679 = ~n667 & ~n678;
  assign n680 = n677 & ~n679;
  assign n681 = ~n677 & n679;
  assign po37  = n680 | n681;
  assign n683 = ~pi38  & ~pi166 ;
  assign n684 = pi38  & pi166 ;
  assign n685 = ~n683 & ~n684;
  assign n686 = ~n676 & ~n679;
  assign n687 = ~n675 & ~n686;
  assign n688 = n685 & ~n687;
  assign n689 = ~n685 & n687;
  assign po38  = n688 | n689;
  assign n691 = ~pi39  & ~pi167 ;
  assign n692 = pi39  & pi167 ;
  assign n693 = ~n691 & ~n692;
  assign n694 = ~n684 & ~n687;
  assign n695 = ~n683 & ~n694;
  assign n696 = n693 & ~n695;
  assign n697 = ~n693 & n695;
  assign po39  = n696 | n697;
  assign n699 = ~pi40  & ~pi168 ;
  assign n700 = pi40  & pi168 ;
  assign n701 = ~n699 & ~n700;
  assign n702 = ~n692 & ~n695;
  assign n703 = ~n691 & ~n702;
  assign n704 = n701 & ~n703;
  assign n705 = ~n701 & n703;
  assign po40  = n704 | n705;
  assign n707 = ~pi41  & ~pi169 ;
  assign n708 = pi41  & pi169 ;
  assign n709 = ~n707 & ~n708;
  assign n710 = ~n700 & ~n703;
  assign n711 = ~n699 & ~n710;
  assign n712 = n709 & ~n711;
  assign n713 = ~n709 & n711;
  assign po41  = n712 | n713;
  assign n715 = ~pi42  & ~pi170 ;
  assign n716 = pi42  & pi170 ;
  assign n717 = ~n715 & ~n716;
  assign n718 = ~n708 & ~n711;
  assign n719 = ~n707 & ~n718;
  assign n720 = n717 & ~n719;
  assign n721 = ~n717 & n719;
  assign po42  = n720 | n721;
  assign n723 = ~pi43  & ~pi171 ;
  assign n724 = pi43  & pi171 ;
  assign n725 = ~n723 & ~n724;
  assign n726 = ~n716 & ~n719;
  assign n727 = ~n715 & ~n726;
  assign n728 = n725 & ~n727;
  assign n729 = ~n725 & n727;
  assign po43  = n728 | n729;
  assign n731 = ~pi44  & ~pi172 ;
  assign n732 = pi44  & pi172 ;
  assign n733 = ~n731 & ~n732;
  assign n734 = ~n724 & ~n727;
  assign n735 = ~n723 & ~n734;
  assign n736 = n733 & ~n735;
  assign n737 = ~n733 & n735;
  assign po44  = n736 | n737;
  assign n739 = ~pi45  & ~pi173 ;
  assign n740 = pi45  & pi173 ;
  assign n741 = ~n739 & ~n740;
  assign n742 = ~n732 & ~n735;
  assign n743 = ~n731 & ~n742;
  assign n744 = n741 & ~n743;
  assign n745 = ~n741 & n743;
  assign po45  = n744 | n745;
  assign n747 = ~pi46  & ~pi174 ;
  assign n748 = pi46  & pi174 ;
  assign n749 = ~n747 & ~n748;
  assign n750 = ~n740 & ~n743;
  assign n751 = ~n739 & ~n750;
  assign n752 = n749 & ~n751;
  assign n753 = ~n749 & n751;
  assign po46  = n752 | n753;
  assign n755 = ~pi47  & ~pi175 ;
  assign n756 = pi47  & pi175 ;
  assign n757 = ~n755 & ~n756;
  assign n758 = ~n748 & ~n751;
  assign n759 = ~n747 & ~n758;
  assign n760 = n757 & ~n759;
  assign n761 = ~n757 & n759;
  assign po47  = n760 | n761;
  assign n763 = ~pi48  & ~pi176 ;
  assign n764 = pi48  & pi176 ;
  assign n765 = ~n763 & ~n764;
  assign n766 = ~n756 & ~n759;
  assign n767 = ~n755 & ~n766;
  assign n768 = n765 & ~n767;
  assign n769 = ~n765 & n767;
  assign po48  = n768 | n769;
  assign n771 = ~pi49  & ~pi177 ;
  assign n772 = pi49  & pi177 ;
  assign n773 = ~n771 & ~n772;
  assign n774 = ~n764 & ~n767;
  assign n775 = ~n763 & ~n774;
  assign n776 = n773 & ~n775;
  assign n777 = ~n773 & n775;
  assign po49  = n776 | n777;
  assign n779 = ~pi50  & ~pi178 ;
  assign n780 = pi50  & pi178 ;
  assign n781 = ~n779 & ~n780;
  assign n782 = ~n772 & ~n775;
  assign n783 = ~n771 & ~n782;
  assign n784 = n781 & ~n783;
  assign n785 = ~n781 & n783;
  assign po50  = n784 | n785;
  assign n787 = ~pi51  & ~pi179 ;
  assign n788 = pi51  & pi179 ;
  assign n789 = ~n787 & ~n788;
  assign n790 = ~n780 & ~n783;
  assign n791 = ~n779 & ~n790;
  assign n792 = n789 & ~n791;
  assign n793 = ~n789 & n791;
  assign po51  = n792 | n793;
  assign n795 = ~pi52  & ~pi180 ;
  assign n796 = pi52  & pi180 ;
  assign n797 = ~n795 & ~n796;
  assign n798 = ~n788 & ~n791;
  assign n799 = ~n787 & ~n798;
  assign n800 = n797 & ~n799;
  assign n801 = ~n797 & n799;
  assign po52  = n800 | n801;
  assign n803 = ~pi53  & ~pi181 ;
  assign n804 = pi53  & pi181 ;
  assign n805 = ~n803 & ~n804;
  assign n806 = ~n796 & ~n799;
  assign n807 = ~n795 & ~n806;
  assign n808 = n805 & ~n807;
  assign n809 = ~n805 & n807;
  assign po53  = n808 | n809;
  assign n811 = ~pi54  & ~pi182 ;
  assign n812 = pi54  & pi182 ;
  assign n813 = ~n811 & ~n812;
  assign n814 = ~n804 & ~n807;
  assign n815 = ~n803 & ~n814;
  assign n816 = n813 & ~n815;
  assign n817 = ~n813 & n815;
  assign po54  = n816 | n817;
  assign n819 = ~pi55  & ~pi183 ;
  assign n820 = pi55  & pi183 ;
  assign n821 = ~n819 & ~n820;
  assign n822 = ~n812 & ~n815;
  assign n823 = ~n811 & ~n822;
  assign n824 = n821 & ~n823;
  assign n825 = ~n821 & n823;
  assign po55  = n824 | n825;
  assign n827 = ~pi56  & ~pi184 ;
  assign n828 = pi56  & pi184 ;
  assign n829 = ~n827 & ~n828;
  assign n830 = ~n820 & ~n823;
  assign n831 = ~n819 & ~n830;
  assign n832 = n829 & ~n831;
  assign n833 = ~n829 & n831;
  assign po56  = n832 | n833;
  assign n835 = ~pi57  & ~pi185 ;
  assign n836 = pi57  & pi185 ;
  assign n837 = ~n835 & ~n836;
  assign n838 = ~n828 & ~n831;
  assign n839 = ~n827 & ~n838;
  assign n840 = n837 & ~n839;
  assign n841 = ~n837 & n839;
  assign po57  = n840 | n841;
  assign n843 = ~pi58  & ~pi186 ;
  assign n844 = pi58  & pi186 ;
  assign n845 = ~n843 & ~n844;
  assign n846 = ~n836 & ~n839;
  assign n847 = ~n835 & ~n846;
  assign n848 = n845 & ~n847;
  assign n849 = ~n845 & n847;
  assign po58  = n848 | n849;
  assign n851 = ~pi59  & ~pi187 ;
  assign n852 = pi59  & pi187 ;
  assign n853 = ~n851 & ~n852;
  assign n854 = ~n844 & ~n847;
  assign n855 = ~n843 & ~n854;
  assign n856 = n853 & ~n855;
  assign n857 = ~n853 & n855;
  assign po59  = n856 | n857;
  assign n859 = ~pi60  & ~pi188 ;
  assign n860 = pi60  & pi188 ;
  assign n861 = ~n859 & ~n860;
  assign n862 = ~n852 & ~n855;
  assign n863 = ~n851 & ~n862;
  assign n864 = n861 & ~n863;
  assign n865 = ~n861 & n863;
  assign po60  = n864 | n865;
  assign n867 = ~pi61  & ~pi189 ;
  assign n868 = pi61  & pi189 ;
  assign n869 = ~n867 & ~n868;
  assign n870 = ~n860 & ~n863;
  assign n871 = ~n859 & ~n870;
  assign n872 = n869 & ~n871;
  assign n873 = ~n869 & n871;
  assign po61  = n872 | n873;
  assign n875 = ~pi62  & ~pi190 ;
  assign n876 = pi62  & pi190 ;
  assign n877 = ~n875 & ~n876;
  assign n878 = ~n868 & ~n871;
  assign n879 = ~n867 & ~n878;
  assign n880 = n877 & ~n879;
  assign n881 = ~n877 & n879;
  assign po62  = n880 | n881;
  assign n883 = ~pi63  & ~pi191 ;
  assign n884 = pi63  & pi191 ;
  assign n885 = ~n883 & ~n884;
  assign n886 = ~n876 & ~n879;
  assign n887 = ~n875 & ~n886;
  assign n888 = n885 & ~n887;
  assign n889 = ~n885 & n887;
  assign po63  = n888 | n889;
  assign n891 = ~pi64  & ~pi192 ;
  assign n892 = pi64  & pi192 ;
  assign n893 = ~n891 & ~n892;
  assign n894 = ~n884 & ~n887;
  assign n895 = ~n883 & ~n894;
  assign n896 = n893 & ~n895;
  assign n897 = ~n893 & n895;
  assign po64  = n896 | n897;
  assign n899 = ~pi65  & ~pi193 ;
  assign n900 = pi65  & pi193 ;
  assign n901 = ~n899 & ~n900;
  assign n902 = ~n892 & ~n895;
  assign n903 = ~n891 & ~n902;
  assign n904 = n901 & ~n903;
  assign n905 = ~n901 & n903;
  assign po65  = n904 | n905;
  assign n907 = ~pi66  & ~pi194 ;
  assign n908 = pi66  & pi194 ;
  assign n909 = ~n907 & ~n908;
  assign n910 = ~n900 & ~n903;
  assign n911 = ~n899 & ~n910;
  assign n912 = n909 & ~n911;
  assign n913 = ~n909 & n911;
  assign po66  = n912 | n913;
  assign n915 = ~pi67  & ~pi195 ;
  assign n916 = pi67  & pi195 ;
  assign n917 = ~n915 & ~n916;
  assign n918 = ~n908 & ~n911;
  assign n919 = ~n907 & ~n918;
  assign n920 = n917 & ~n919;
  assign n921 = ~n917 & n919;
  assign po67  = n920 | n921;
  assign n923 = ~pi68  & ~pi196 ;
  assign n924 = pi68  & pi196 ;
  assign n925 = ~n923 & ~n924;
  assign n926 = ~n916 & ~n919;
  assign n927 = ~n915 & ~n926;
  assign n928 = n925 & ~n927;
  assign n929 = ~n925 & n927;
  assign po68  = n928 | n929;
  assign n931 = ~pi69  & ~pi197 ;
  assign n932 = pi69  & pi197 ;
  assign n933 = ~n931 & ~n932;
  assign n934 = ~n924 & ~n927;
  assign n935 = ~n923 & ~n934;
  assign n936 = n933 & ~n935;
  assign n937 = ~n933 & n935;
  assign po69  = n936 | n937;
  assign n939 = ~pi70  & ~pi198 ;
  assign n940 = pi70  & pi198 ;
  assign n941 = ~n939 & ~n940;
  assign n942 = ~n932 & ~n935;
  assign n943 = ~n931 & ~n942;
  assign n944 = n941 & ~n943;
  assign n945 = ~n941 & n943;
  assign po70  = n944 | n945;
  assign n947 = ~pi71  & ~pi199 ;
  assign n948 = pi71  & pi199 ;
  assign n949 = ~n947 & ~n948;
  assign n950 = ~n940 & ~n943;
  assign n951 = ~n939 & ~n950;
  assign n952 = n949 & ~n951;
  assign n953 = ~n949 & n951;
  assign po71  = n952 | n953;
  assign n955 = ~pi72  & ~pi200 ;
  assign n956 = pi72  & pi200 ;
  assign n957 = ~n955 & ~n956;
  assign n958 = ~n948 & ~n951;
  assign n959 = ~n947 & ~n958;
  assign n960 = n957 & ~n959;
  assign n961 = ~n957 & n959;
  assign po72  = n960 | n961;
  assign n963 = ~pi73  & ~pi201 ;
  assign n964 = pi73  & pi201 ;
  assign n965 = ~n963 & ~n964;
  assign n966 = ~n956 & ~n959;
  assign n967 = ~n955 & ~n966;
  assign n968 = n965 & ~n967;
  assign n969 = ~n965 & n967;
  assign po73  = n968 | n969;
  assign n971 = ~pi74  & ~pi202 ;
  assign n972 = pi74  & pi202 ;
  assign n973 = ~n971 & ~n972;
  assign n974 = ~n964 & ~n967;
  assign n975 = ~n963 & ~n974;
  assign n976 = n973 & ~n975;
  assign n977 = ~n973 & n975;
  assign po74  = n976 | n977;
  assign n979 = ~pi75  & ~pi203 ;
  assign n980 = pi75  & pi203 ;
  assign n981 = ~n979 & ~n980;
  assign n982 = ~n972 & ~n975;
  assign n983 = ~n971 & ~n982;
  assign n984 = n981 & ~n983;
  assign n985 = ~n981 & n983;
  assign po75  = n984 | n985;
  assign n987 = ~pi76  & ~pi204 ;
  assign n988 = pi76  & pi204 ;
  assign n989 = ~n987 & ~n988;
  assign n990 = ~n980 & ~n983;
  assign n991 = ~n979 & ~n990;
  assign n992 = n989 & ~n991;
  assign n993 = ~n989 & n991;
  assign po76  = n992 | n993;
  assign n995 = ~pi77  & ~pi205 ;
  assign n996 = pi77  & pi205 ;
  assign n997 = ~n995 & ~n996;
  assign n998 = ~n988 & ~n991;
  assign n999 = ~n987 & ~n998;
  assign n1000 = n997 & ~n999;
  assign n1001 = ~n997 & n999;
  assign po77  = n1000 | n1001;
  assign n1003 = ~pi78  & ~pi206 ;
  assign n1004 = pi78  & pi206 ;
  assign n1005 = ~n1003 & ~n1004;
  assign n1006 = ~n996 & ~n999;
  assign n1007 = ~n995 & ~n1006;
  assign n1008 = n1005 & ~n1007;
  assign n1009 = ~n1005 & n1007;
  assign po78  = n1008 | n1009;
  assign n1011 = ~pi79  & ~pi207 ;
  assign n1012 = pi79  & pi207 ;
  assign n1013 = ~n1011 & ~n1012;
  assign n1014 = ~n1004 & ~n1007;
  assign n1015 = ~n1003 & ~n1014;
  assign n1016 = n1013 & ~n1015;
  assign n1017 = ~n1013 & n1015;
  assign po79  = n1016 | n1017;
  assign n1019 = ~pi80  & ~pi208 ;
  assign n1020 = pi80  & pi208 ;
  assign n1021 = ~n1019 & ~n1020;
  assign n1022 = ~n1012 & ~n1015;
  assign n1023 = ~n1011 & ~n1022;
  assign n1024 = n1021 & ~n1023;
  assign n1025 = ~n1021 & n1023;
  assign po80  = n1024 | n1025;
  assign n1027 = ~pi81  & ~pi209 ;
  assign n1028 = pi81  & pi209 ;
  assign n1029 = ~n1027 & ~n1028;
  assign n1030 = ~n1020 & ~n1023;
  assign n1031 = ~n1019 & ~n1030;
  assign n1032 = n1029 & ~n1031;
  assign n1033 = ~n1029 & n1031;
  assign po81  = n1032 | n1033;
  assign n1035 = ~pi82  & ~pi210 ;
  assign n1036 = pi82  & pi210 ;
  assign n1037 = ~n1035 & ~n1036;
  assign n1038 = ~n1028 & ~n1031;
  assign n1039 = ~n1027 & ~n1038;
  assign n1040 = n1037 & ~n1039;
  assign n1041 = ~n1037 & n1039;
  assign po82  = n1040 | n1041;
  assign n1043 = ~pi83  & ~pi211 ;
  assign n1044 = pi83  & pi211 ;
  assign n1045 = ~n1043 & ~n1044;
  assign n1046 = ~n1036 & ~n1039;
  assign n1047 = ~n1035 & ~n1046;
  assign n1048 = n1045 & ~n1047;
  assign n1049 = ~n1045 & n1047;
  assign po83  = n1048 | n1049;
  assign n1051 = ~pi84  & ~pi212 ;
  assign n1052 = pi84  & pi212 ;
  assign n1053 = ~n1051 & ~n1052;
  assign n1054 = ~n1044 & ~n1047;
  assign n1055 = ~n1043 & ~n1054;
  assign n1056 = n1053 & ~n1055;
  assign n1057 = ~n1053 & n1055;
  assign po84  = n1056 | n1057;
  assign n1059 = ~pi85  & ~pi213 ;
  assign n1060 = pi85  & pi213 ;
  assign n1061 = ~n1059 & ~n1060;
  assign n1062 = ~n1052 & ~n1055;
  assign n1063 = ~n1051 & ~n1062;
  assign n1064 = n1061 & ~n1063;
  assign n1065 = ~n1061 & n1063;
  assign po85  = n1064 | n1065;
  assign n1067 = ~pi86  & ~pi214 ;
  assign n1068 = pi86  & pi214 ;
  assign n1069 = ~n1067 & ~n1068;
  assign n1070 = ~n1060 & ~n1063;
  assign n1071 = ~n1059 & ~n1070;
  assign n1072 = n1069 & ~n1071;
  assign n1073 = ~n1069 & n1071;
  assign po86  = n1072 | n1073;
  assign n1075 = ~pi87  & ~pi215 ;
  assign n1076 = pi87  & pi215 ;
  assign n1077 = ~n1075 & ~n1076;
  assign n1078 = ~n1068 & ~n1071;
  assign n1079 = ~n1067 & ~n1078;
  assign n1080 = n1077 & ~n1079;
  assign n1081 = ~n1077 & n1079;
  assign po87  = n1080 | n1081;
  assign n1083 = ~pi88  & ~pi216 ;
  assign n1084 = pi88  & pi216 ;
  assign n1085 = ~n1083 & ~n1084;
  assign n1086 = ~n1076 & ~n1079;
  assign n1087 = ~n1075 & ~n1086;
  assign n1088 = n1085 & ~n1087;
  assign n1089 = ~n1085 & n1087;
  assign po88  = n1088 | n1089;
  assign n1091 = ~pi89  & ~pi217 ;
  assign n1092 = pi89  & pi217 ;
  assign n1093 = ~n1091 & ~n1092;
  assign n1094 = ~n1084 & ~n1087;
  assign n1095 = ~n1083 & ~n1094;
  assign n1096 = n1093 & ~n1095;
  assign n1097 = ~n1093 & n1095;
  assign po89  = n1096 | n1097;
  assign n1099 = ~pi90  & ~pi218 ;
  assign n1100 = pi90  & pi218 ;
  assign n1101 = ~n1099 & ~n1100;
  assign n1102 = ~n1092 & ~n1095;
  assign n1103 = ~n1091 & ~n1102;
  assign n1104 = n1101 & ~n1103;
  assign n1105 = ~n1101 & n1103;
  assign po90  = n1104 | n1105;
  assign n1107 = ~pi91  & ~pi219 ;
  assign n1108 = pi91  & pi219 ;
  assign n1109 = ~n1107 & ~n1108;
  assign n1110 = ~n1100 & ~n1103;
  assign n1111 = ~n1099 & ~n1110;
  assign n1112 = n1109 & ~n1111;
  assign n1113 = ~n1109 & n1111;
  assign po91  = n1112 | n1113;
  assign n1115 = ~pi92  & ~pi220 ;
  assign n1116 = pi92  & pi220 ;
  assign n1117 = ~n1115 & ~n1116;
  assign n1118 = ~n1108 & ~n1111;
  assign n1119 = ~n1107 & ~n1118;
  assign n1120 = n1117 & ~n1119;
  assign n1121 = ~n1117 & n1119;
  assign po92  = n1120 | n1121;
  assign n1123 = ~pi93  & ~pi221 ;
  assign n1124 = pi93  & pi221 ;
  assign n1125 = ~n1123 & ~n1124;
  assign n1126 = ~n1116 & ~n1119;
  assign n1127 = ~n1115 & ~n1126;
  assign n1128 = n1125 & ~n1127;
  assign n1129 = ~n1125 & n1127;
  assign po93  = n1128 | n1129;
  assign n1131 = ~pi94  & ~pi222 ;
  assign n1132 = pi94  & pi222 ;
  assign n1133 = ~n1131 & ~n1132;
  assign n1134 = ~n1124 & ~n1127;
  assign n1135 = ~n1123 & ~n1134;
  assign n1136 = n1133 & ~n1135;
  assign n1137 = ~n1133 & n1135;
  assign po94  = n1136 | n1137;
  assign n1139 = ~pi95  & ~pi223 ;
  assign n1140 = pi95  & pi223 ;
  assign n1141 = ~n1139 & ~n1140;
  assign n1142 = ~n1132 & ~n1135;
  assign n1143 = ~n1131 & ~n1142;
  assign n1144 = n1141 & ~n1143;
  assign n1145 = ~n1141 & n1143;
  assign po95  = n1144 | n1145;
  assign n1147 = ~pi96  & ~pi224 ;
  assign n1148 = pi96  & pi224 ;
  assign n1149 = ~n1147 & ~n1148;
  assign n1150 = ~n1140 & ~n1143;
  assign n1151 = ~n1139 & ~n1150;
  assign n1152 = n1149 & ~n1151;
  assign n1153 = ~n1149 & n1151;
  assign po96  = n1152 | n1153;
  assign n1155 = ~pi97  & ~pi225 ;
  assign n1156 = pi97  & pi225 ;
  assign n1157 = ~n1155 & ~n1156;
  assign n1158 = ~n1148 & ~n1151;
  assign n1159 = ~n1147 & ~n1158;
  assign n1160 = n1157 & ~n1159;
  assign n1161 = ~n1157 & n1159;
  assign po97  = n1160 | n1161;
  assign n1163 = ~pi98  & ~pi226 ;
  assign n1164 = pi98  & pi226 ;
  assign n1165 = ~n1163 & ~n1164;
  assign n1166 = ~n1156 & ~n1159;
  assign n1167 = ~n1155 & ~n1166;
  assign n1168 = n1165 & ~n1167;
  assign n1169 = ~n1165 & n1167;
  assign po98  = n1168 | n1169;
  assign n1171 = ~pi99  & ~pi227 ;
  assign n1172 = pi99  & pi227 ;
  assign n1173 = ~n1171 & ~n1172;
  assign n1174 = ~n1164 & ~n1167;
  assign n1175 = ~n1163 & ~n1174;
  assign n1176 = n1173 & ~n1175;
  assign n1177 = ~n1173 & n1175;
  assign po99  = n1176 | n1177;
  assign n1179 = ~pi100  & ~pi228 ;
  assign n1180 = pi100  & pi228 ;
  assign n1181 = ~n1179 & ~n1180;
  assign n1182 = ~n1172 & ~n1175;
  assign n1183 = ~n1171 & ~n1182;
  assign n1184 = n1181 & ~n1183;
  assign n1185 = ~n1181 & n1183;
  assign po100  = n1184 | n1185;
  assign n1187 = ~pi101  & ~pi229 ;
  assign n1188 = pi101  & pi229 ;
  assign n1189 = ~n1187 & ~n1188;
  assign n1190 = ~n1180 & ~n1183;
  assign n1191 = ~n1179 & ~n1190;
  assign n1192 = n1189 & ~n1191;
  assign n1193 = ~n1189 & n1191;
  assign po101  = n1192 | n1193;
  assign n1195 = ~pi102  & ~pi230 ;
  assign n1196 = pi102  & pi230 ;
  assign n1197 = ~n1195 & ~n1196;
  assign n1198 = ~n1188 & ~n1191;
  assign n1199 = ~n1187 & ~n1198;
  assign n1200 = n1197 & ~n1199;
  assign n1201 = ~n1197 & n1199;
  assign po102  = n1200 | n1201;
  assign n1203 = ~pi103  & ~pi231 ;
  assign n1204 = pi103  & pi231 ;
  assign n1205 = ~n1203 & ~n1204;
  assign n1206 = ~n1196 & ~n1199;
  assign n1207 = ~n1195 & ~n1206;
  assign n1208 = n1205 & ~n1207;
  assign n1209 = ~n1205 & n1207;
  assign po103  = n1208 | n1209;
  assign n1211 = ~pi104  & ~pi232 ;
  assign n1212 = pi104  & pi232 ;
  assign n1213 = ~n1211 & ~n1212;
  assign n1214 = ~n1204 & ~n1207;
  assign n1215 = ~n1203 & ~n1214;
  assign n1216 = n1213 & ~n1215;
  assign n1217 = ~n1213 & n1215;
  assign po104  = n1216 | n1217;
  assign n1219 = ~pi105  & ~pi233 ;
  assign n1220 = pi105  & pi233 ;
  assign n1221 = ~n1219 & ~n1220;
  assign n1222 = ~n1212 & ~n1215;
  assign n1223 = ~n1211 & ~n1222;
  assign n1224 = n1221 & ~n1223;
  assign n1225 = ~n1221 & n1223;
  assign po105  = n1224 | n1225;
  assign n1227 = ~pi106  & ~pi234 ;
  assign n1228 = pi106  & pi234 ;
  assign n1229 = ~n1227 & ~n1228;
  assign n1230 = ~n1220 & ~n1223;
  assign n1231 = ~n1219 & ~n1230;
  assign n1232 = n1229 & ~n1231;
  assign n1233 = ~n1229 & n1231;
  assign po106  = n1232 | n1233;
  assign n1235 = ~pi107  & ~pi235 ;
  assign n1236 = pi107  & pi235 ;
  assign n1237 = ~n1235 & ~n1236;
  assign n1238 = ~n1228 & ~n1231;
  assign n1239 = ~n1227 & ~n1238;
  assign n1240 = n1237 & ~n1239;
  assign n1241 = ~n1237 & n1239;
  assign po107  = n1240 | n1241;
  assign n1243 = ~pi108  & ~pi236 ;
  assign n1244 = pi108  & pi236 ;
  assign n1245 = ~n1243 & ~n1244;
  assign n1246 = ~n1236 & ~n1239;
  assign n1247 = ~n1235 & ~n1246;
  assign n1248 = n1245 & ~n1247;
  assign n1249 = ~n1245 & n1247;
  assign po108  = n1248 | n1249;
  assign n1251 = ~pi109  & ~pi237 ;
  assign n1252 = pi109  & pi237 ;
  assign n1253 = ~n1251 & ~n1252;
  assign n1254 = ~n1244 & ~n1247;
  assign n1255 = ~n1243 & ~n1254;
  assign n1256 = n1253 & ~n1255;
  assign n1257 = ~n1253 & n1255;
  assign po109  = n1256 | n1257;
  assign n1259 = ~pi110  & ~pi238 ;
  assign n1260 = pi110  & pi238 ;
  assign n1261 = ~n1259 & ~n1260;
  assign n1262 = ~n1252 & ~n1255;
  assign n1263 = ~n1251 & ~n1262;
  assign n1264 = n1261 & ~n1263;
  assign n1265 = ~n1261 & n1263;
  assign po110  = n1264 | n1265;
  assign n1267 = ~pi111  & ~pi239 ;
  assign n1268 = pi111  & pi239 ;
  assign n1269 = ~n1267 & ~n1268;
  assign n1270 = ~n1260 & ~n1263;
  assign n1271 = ~n1259 & ~n1270;
  assign n1272 = n1269 & ~n1271;
  assign n1273 = ~n1269 & n1271;
  assign po111  = n1272 | n1273;
  assign n1275 = ~pi112  & ~pi240 ;
  assign n1276 = pi112  & pi240 ;
  assign n1277 = ~n1275 & ~n1276;
  assign n1278 = ~n1268 & ~n1271;
  assign n1279 = ~n1267 & ~n1278;
  assign n1280 = n1277 & ~n1279;
  assign n1281 = ~n1277 & n1279;
  assign po112  = n1280 | n1281;
  assign n1283 = ~pi113  & ~pi241 ;
  assign n1284 = pi113  & pi241 ;
  assign n1285 = ~n1283 & ~n1284;
  assign n1286 = ~n1276 & ~n1279;
  assign n1287 = ~n1275 & ~n1286;
  assign n1288 = n1285 & ~n1287;
  assign n1289 = ~n1285 & n1287;
  assign po113  = n1288 | n1289;
  assign n1291 = ~pi114  & ~pi242 ;
  assign n1292 = pi114  & pi242 ;
  assign n1293 = ~n1291 & ~n1292;
  assign n1294 = ~n1284 & ~n1287;
  assign n1295 = ~n1283 & ~n1294;
  assign n1296 = n1293 & ~n1295;
  assign n1297 = ~n1293 & n1295;
  assign po114  = n1296 | n1297;
  assign n1299 = ~pi115  & ~pi243 ;
  assign n1300 = pi115  & pi243 ;
  assign n1301 = ~n1299 & ~n1300;
  assign n1302 = ~n1292 & ~n1295;
  assign n1303 = ~n1291 & ~n1302;
  assign n1304 = n1301 & ~n1303;
  assign n1305 = ~n1301 & n1303;
  assign po115  = n1304 | n1305;
  assign n1307 = ~pi116  & ~pi244 ;
  assign n1308 = pi116  & pi244 ;
  assign n1309 = ~n1307 & ~n1308;
  assign n1310 = ~n1300 & ~n1303;
  assign n1311 = ~n1299 & ~n1310;
  assign n1312 = n1309 & ~n1311;
  assign n1313 = ~n1309 & n1311;
  assign po116  = n1312 | n1313;
  assign n1315 = ~pi117  & ~pi245 ;
  assign n1316 = pi117  & pi245 ;
  assign n1317 = ~n1315 & ~n1316;
  assign n1318 = ~n1308 & ~n1311;
  assign n1319 = ~n1307 & ~n1318;
  assign n1320 = n1317 & ~n1319;
  assign n1321 = ~n1317 & n1319;
  assign po117  = n1320 | n1321;
  assign n1323 = ~pi118  & ~pi246 ;
  assign n1324 = pi118  & pi246 ;
  assign n1325 = ~n1323 & ~n1324;
  assign n1326 = ~n1316 & ~n1319;
  assign n1327 = ~n1315 & ~n1326;
  assign n1328 = n1325 & ~n1327;
  assign n1329 = ~n1325 & n1327;
  assign po118  = n1328 | n1329;
  assign n1331 = ~pi119  & ~pi247 ;
  assign n1332 = pi119  & pi247 ;
  assign n1333 = ~n1331 & ~n1332;
  assign n1334 = ~n1324 & ~n1327;
  assign n1335 = ~n1323 & ~n1334;
  assign n1336 = n1333 & ~n1335;
  assign n1337 = ~n1333 & n1335;
  assign po119  = n1336 | n1337;
  assign n1339 = ~pi120  & ~pi248 ;
  assign n1340 = pi120  & pi248 ;
  assign n1341 = ~n1339 & ~n1340;
  assign n1342 = ~n1332 & ~n1335;
  assign n1343 = ~n1331 & ~n1342;
  assign n1344 = n1341 & ~n1343;
  assign n1345 = ~n1341 & n1343;
  assign po120  = n1344 | n1345;
  assign n1347 = ~pi121  & ~pi249 ;
  assign n1348 = pi121  & pi249 ;
  assign n1349 = ~n1347 & ~n1348;
  assign n1350 = ~n1340 & ~n1343;
  assign n1351 = ~n1339 & ~n1350;
  assign n1352 = n1349 & ~n1351;
  assign n1353 = ~n1349 & n1351;
  assign po121  = n1352 | n1353;
  assign n1355 = ~pi122  & ~pi250 ;
  assign n1356 = pi122  & pi250 ;
  assign n1357 = ~n1355 & ~n1356;
  assign n1358 = ~n1348 & ~n1351;
  assign n1359 = ~n1347 & ~n1358;
  assign n1360 = n1357 & ~n1359;
  assign n1361 = ~n1357 & n1359;
  assign po122  = n1360 | n1361;
  assign n1363 = ~pi123  & ~pi251 ;
  assign n1364 = pi123  & pi251 ;
  assign n1365 = ~n1363 & ~n1364;
  assign n1366 = ~n1356 & ~n1359;
  assign n1367 = ~n1355 & ~n1366;
  assign n1368 = n1365 & ~n1367;
  assign n1369 = ~n1365 & n1367;
  assign po123  = n1368 | n1369;
  assign n1371 = ~pi124  & ~pi252 ;
  assign n1372 = pi124  & pi252 ;
  assign n1373 = ~n1371 & ~n1372;
  assign n1374 = ~n1364 & ~n1367;
  assign n1375 = ~n1363 & ~n1374;
  assign n1376 = n1373 & ~n1375;
  assign n1377 = ~n1373 & n1375;
  assign po124  = n1376 | n1377;
  assign n1379 = ~pi125  & ~pi253 ;
  assign n1380 = pi125  & pi253 ;
  assign n1381 = ~n1379 & ~n1380;
  assign n1382 = ~n1372 & ~n1375;
  assign n1383 = ~n1371 & ~n1382;
  assign n1384 = n1381 & ~n1383;
  assign n1385 = ~n1381 & n1383;
  assign po125  = n1384 | n1385;
  assign n1387 = ~pi126  & ~pi254 ;
  assign n1388 = pi126  & pi254 ;
  assign n1389 = ~n1387 & ~n1388;
  assign n1390 = ~n1380 & ~n1383;
  assign n1391 = ~n1379 & ~n1390;
  assign n1392 = n1389 & ~n1391;
  assign n1393 = ~n1389 & n1391;
  assign po126  = n1392 | n1393;
  assign n1395 = ~pi127  & ~pi255 ;
  assign n1396 = pi127  & pi255 ;
  assign n1397 = ~n1395 & ~n1396;
  assign n1398 = ~n1388 & ~n1391;
  assign n1399 = ~n1387 & ~n1398;
  assign n1400 = n1397 & ~n1399;
  assign n1401 = ~n1397 & n1399;
  assign po127  = n1400 | n1401;
  assign n1403 = ~n1396 & ~n1399;
  assign po128 = ~n1395 & ~n1403;
endmodule
