module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 , pi32 ,
    pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 , pi40 ,
    pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 , pi56 ,
    pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 , pi64 ,
    pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 , pi73 ,
    pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 , pi81 ,
    pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 , pi89 ,
    pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 , pi97 ,
    pi98 , pi99 , pi100 , pi101 , pi102 , pi103 , pi104 , pi105 ,
    pi106 , pi107 , pi108 , pi109 , pi110 , pi111 , pi112 , pi113 ,
    pi114 , pi115 , pi116 , pi117 , pi118 , pi119 , pi120 , pi121 ,
    pi122 , pi123 , pi124 , pi125 , pi126 , pi127 ,
    po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7 , po8 ,
    po9 , po10 , po11 , po12 , po13 , po14 , po15 , po16 ,
    po17 , po18 , po19 , po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 , po30 , po31 , po32 ,
    po33 , po34 , po35 , po36 , po37 , po38 , po39 , po40 ,
    po41 , po42 , po43 , po44 , po45 , po46 , po47 , po48 ,
    po49 , po50 , po51 , po52 , po53 , po54 , po55 , po56 ,
    po57 , po58 , po59 , po60 , po61 , po62 , po63 , po64 ,
    po65 , po66 , po67 , po68 , po69 , po70 , po71 , po72 ,
    po73 , po74 , po75 , po76 , po77 , po78 , po79 , po80 ,
    po81 , po82 , po83 , po84 , po85 , po86 , po87 , po88 ,
    po89 , po90 , po91 , po92 , po93 , po94 , po95 , po96 ,
    po97 , po98 , po99 , po100 , po101 , po102 , po103 ,
    po104 , po105 , po106 , po107 , po108 , po109 , po110 ,
    po111 , po112 , po113 , po114 , po115 , po116 , po117 ,
    po118 , po119 , po120 , po121 , po122 , po123 , po124 ,
    po125 , po126 , po127   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    pi32 , pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 ,
    pi56 , pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 ,
    pi64 , pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 ,
    pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 ,
    pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 ,
    pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 ,
    pi97 , pi98 , pi99 , pi100 , pi101 , pi102 , pi103 , pi104 ,
    pi105 , pi106 , pi107 , pi108 , pi109 , pi110 , pi111 , pi112 ,
    pi113 , pi114 , pi115 , pi116 , pi117 , pi118 , pi119 , pi120 ,
    pi121 , pi122 , pi123 , pi124 , pi125 , pi126 , pi127 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7 ,
    po8 , po9 , po10 , po11 , po12 , po13 , po14 , po15 ,
    po16 , po17 , po18 , po19 , po20 , po21 , po22 , po23 ,
    po24 , po25 , po26 , po27 , po28 , po29 , po30 , po31 ,
    po32 , po33 , po34 , po35 , po36 , po37 , po38 , po39 ,
    po40 , po41 , po42 , po43 , po44 , po45 , po46 , po47 ,
    po48 , po49 , po50 , po51 , po52 , po53 , po54 , po55 ,
    po56 , po57 , po58 , po59 , po60 , po61 , po62 , po63 ,
    po64 , po65 , po66 , po67 , po68 , po69 , po70 , po71 ,
    po72 , po73 , po74 , po75 , po76 , po77 , po78 , po79 ,
    po80 , po81 , po82 , po83 , po84 , po85 , po86 , po87 ,
    po88 , po89 , po90 , po91 , po92 , po93 , po94 , po95 ,
    po96 , po97 , po98 , po99 , po100 , po101 , po102 ,
    po103 , po104 , po105 , po106 , po107 , po108 , po109 ,
    po110 , po111 , po112 , po113 , po114 , po115 , po116 ,
    po117 , po118 , po119 , po120 , po121 , po122 , po123 ,
    po124 , po125 , po126 , po127 ;
  wire n258, n259, n260, n261, n262, n263, n264,
    n265, n266, n267, n268, n269, n270, n271,
    n272, n273, n274, n275, n276, n277, n278,
    n280, n281, n282, n283, n284, n285, n286,
    n287, n288, n289, n290, n291, n292, n293,
    n294, n295, n296, n297, n298, n299, n300,
    n302, n303, n304, n305, n306, n307, n308,
    n309, n310, n311, n312, n313, n314, n315,
    n316, n317, n318, n319, n320, n321, n322,
    n323, n324, n325, n326, n327, n328, n329,
    n331, n332, n333, n334, n335, n336, n337,
    n338, n339, n340, n341, n342, n343, n344,
    n345, n346, n347, n348, n349, n350, n351,
    n352, n353, n354, n355, n356, n357, n358,
    n359, n360, n361, n362, n363, n364, n365,
    n366, n367, n368, n369, n370, n371, n372,
    n373, n374, n375, n376, n377, n379, n380,
    n381, n382, n383, n384, n385, n386, n387,
    n388, n389, n390, n391, n392, n393, n394,
    n395, n396, n397, n398, n399, n400, n401,
    n402, n403, n404, n405, n406, n407, n408,
    n409, n410, n411, n412, n413, n414, n415,
    n416, n417, n418, n419, n421, n422, n423,
    n424, n425, n426, n427, n428, n429, n430,
    n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444,
    n445, n446, n447, n448, n449, n450, n451,
    n452, n453, n454, n455, n456, n457, n458,
    n459, n460, n461, n462, n463, n464, n465,
    n466, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487,
    n488, n489, n490, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501,
    n502, n503, n504, n505, n506, n507, n508,
    n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n532, n533, n535, n536, n537,
    n538, n539, n540, n541, n542, n543, n544,
    n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n557, n558,
    n559, n560, n561, n562, n563, n564, n565,
    n566, n567, n568, n569, n570, n571, n572,
    n573, n574, n575, n576, n577, n578, n579,
    n580, n581, n582, n583, n584, n585, n586,
    n587, n588, n589, n590, n591, n592, n593,
    n594, n596, n597, n598, n599, n600, n601,
    n602, n603, n604, n605, n606, n607, n608,
    n609, n610, n611, n612, n613, n614, n615,
    n616, n617, n618, n619, n620, n621, n622,
    n623, n624, n625, n626, n627, n628, n629,
    n630, n631, n632, n633, n634, n635, n636,
    n637, n638, n639, n640, n641, n642, n643,
    n644, n645, n646, n647, n648, n649, n650,
    n651, n652, n653, n654, n655, n656, n657,
    n658, n659, n660, n662, n663, n664, n665,
    n666, n667, n668, n669, n670, n671, n672,
    n673, n674, n675, n676, n677, n678, n679,
    n680, n681, n682, n683, n684, n685, n686,
    n687, n688, n689, n690, n691, n692, n693,
    n694, n695, n696, n697, n698, n699, n700,
    n701, n702, n703, n704, n705, n706, n707,
    n708, n709, n710, n711, n712, n713, n714,
    n715, n716, n717, n718, n719, n720, n721,
    n722, n723, n724, n725, n726, n727, n728,
    n729, n730, n731, n732, n733, n734, n735,
    n736, n737, n738, n739, n740, n741, n742,
    n743, n744, n745, n747, n748, n749, n750,
    n751, n752, n753, n754, n755, n756, n757,
    n758, n759, n760, n761, n762, n763, n764,
    n765, n766, n767, n768, n769, n770, n771,
    n772, n773, n774, n775, n776, n777, n778,
    n779, n780, n781, n782, n783, n784, n785,
    n786, n787, n788, n789, n790, n791, n792,
    n793, n794, n795, n796, n797, n798, n799,
    n800, n801, n802, n803, n804, n805, n806,
    n807, n808, n809, n810, n811, n812, n813,
    n814, n815, n816, n817, n818, n819, n820,
    n821, n822, n823, n824, n825, n827, n828,
    n829, n830, n831, n832, n833, n834, n835,
    n836, n837, n838, n839, n840, n841, n842,
    n843, n844, n845, n846, n847, n848, n849,
    n850, n851, n852, n853, n854, n855, n856,
    n857, n858, n859, n860, n861, n862, n863,
    n864, n865, n866, n867, n868, n869, n870,
    n871, n872, n873, n874, n875, n876, n877,
    n878, n879, n880, n881, n882, n883, n884,
    n885, n886, n887, n888, n889, n890, n891,
    n892, n893, n894, n895, n896, n897, n898,
    n899, n900, n901, n902, n903, n904, n905,
    n906, n907, n908, n909, n910, n912, n913,
    n914, n915, n916, n917, n918, n919, n920,
    n921, n922, n923, n924, n925, n926, n927,
    n928, n929, n930, n931, n932, n933, n934,
    n935, n936, n937, n938, n939, n940, n941,
    n942, n943, n944, n945, n946, n947, n948,
    n949, n950, n951, n952, n953, n954, n955,
    n956, n957, n958, n959, n960, n961, n962,
    n963, n964, n965, n966, n967, n968, n969,
    n970, n971, n972, n973, n974, n975, n976,
    n977, n978, n979, n980, n981, n982, n983,
    n984, n985, n986, n987, n988, n989, n990,
    n991, n992, n993, n994, n995, n996, n997,
    n998, n999, n1000, n1001, n1002, n1003,
    n1004, n1005, n1006, n1007, n1008, n1009,
    n1010, n1011, n1012, n1013, n1014, n1015,
    n1017, n1018, n1019, n1020, n1021, n1022,
    n1023, n1024, n1025, n1026, n1027, n1028,
    n1029, n1030, n1031, n1032, n1033, n1034,
    n1035, n1036, n1037, n1038, n1039, n1040,
    n1041, n1042, n1043, n1044, n1045, n1046,
    n1047, n1048, n1049, n1050, n1051, n1052,
    n1053, n1054, n1055, n1056, n1057, n1058,
    n1059, n1060, n1061, n1062, n1063, n1064,
    n1065, n1066, n1067, n1068, n1069, n1070,
    n1071, n1072, n1073, n1074, n1075, n1076,
    n1077, n1078, n1079, n1080, n1081, n1082,
    n1083, n1084, n1085, n1086, n1087, n1088,
    n1089, n1090, n1091, n1092, n1093, n1094,
    n1095, n1096, n1097, n1098, n1099, n1100,
    n1101, n1102, n1103, n1104, n1105, n1106,
    n1107, n1108, n1109, n1110, n1111, n1112,
    n1114, n1115, n1116, n1117, n1118, n1119,
    n1120, n1121, n1122, n1123, n1124, n1125,
    n1126, n1127, n1128, n1129, n1130, n1131,
    n1132, n1133, n1134, n1135, n1136, n1137,
    n1138, n1139, n1140, n1141, n1142, n1143,
    n1144, n1145, n1146, n1147, n1148, n1149,
    n1150, n1151, n1152, n1153, n1154, n1155,
    n1156, n1157, n1158, n1159, n1160, n1161,
    n1162, n1163, n1164, n1165, n1166, n1167,
    n1168, n1169, n1170, n1171, n1172, n1173,
    n1174, n1175, n1176, n1177, n1178, n1179,
    n1180, n1181, n1182, n1183, n1184, n1185,
    n1186, n1187, n1188, n1189, n1190, n1191,
    n1192, n1193, n1194, n1195, n1196, n1197,
    n1198, n1199, n1200, n1201, n1202, n1203,
    n1204, n1205, n1206, n1207, n1208, n1209,
    n1210, n1211, n1212, n1213, n1214, n1215,
    n1216, n1218, n1219, n1220, n1221, n1222,
    n1223, n1224, n1225, n1226, n1227, n1228,
    n1229, n1230, n1231, n1232, n1233, n1234,
    n1235, n1236, n1237, n1238, n1239, n1240,
    n1241, n1242, n1243, n1244, n1245, n1246,
    n1247, n1248, n1249, n1250, n1251, n1252,
    n1253, n1254, n1255, n1256, n1257, n1258,
    n1259, n1260, n1261, n1262, n1263, n1264,
    n1265, n1266, n1267, n1268, n1269, n1270,
    n1271, n1272, n1273, n1274, n1275, n1276,
    n1277, n1278, n1279, n1280, n1281, n1282,
    n1283, n1284, n1285, n1286, n1287, n1288,
    n1289, n1290, n1291, n1292, n1293, n1294,
    n1295, n1296, n1297, n1298, n1299, n1300,
    n1301, n1302, n1303, n1304, n1305, n1306,
    n1307, n1308, n1309, n1310, n1311, n1312,
    n1313, n1314, n1315, n1316, n1317, n1318,
    n1319, n1320, n1321, n1322, n1323, n1324,
    n1325, n1326, n1327, n1328, n1329, n1330,
    n1331, n1332, n1333, n1334, n1335, n1336,
    n1338, n1339, n1340, n1341, n1342, n1343,
    n1344, n1345, n1346, n1347, n1348, n1349,
    n1350, n1351, n1352, n1353, n1354, n1355,
    n1356, n1357, n1358, n1359, n1360, n1361,
    n1362, n1363, n1364, n1365, n1366, n1367,
    n1368, n1369, n1370, n1371, n1372, n1373,
    n1374, n1375, n1376, n1377, n1378, n1379,
    n1380, n1381, n1382, n1383, n1384, n1385,
    n1386, n1387, n1388, n1389, n1390, n1391,
    n1392, n1393, n1394, n1395, n1396, n1397,
    n1398, n1399, n1400, n1401, n1402, n1403,
    n1404, n1405, n1406, n1407, n1408, n1409,
    n1410, n1411, n1412, n1413, n1414, n1415,
    n1416, n1417, n1418, n1419, n1420, n1421,
    n1422, n1423, n1424, n1425, n1426, n1427,
    n1428, n1429, n1430, n1431, n1432, n1433,
    n1434, n1435, n1436, n1437, n1438, n1439,
    n1440, n1441, n1442, n1443, n1444, n1445,
    n1446, n1447, n1448, n1449, n1450, n1451,
    n1452, n1453, n1455, n1456, n1457, n1458,
    n1459, n1460, n1461, n1462, n1463, n1464,
    n1465, n1466, n1467, n1468, n1469, n1470,
    n1471, n1472, n1473, n1474, n1475, n1476,
    n1477, n1478, n1479, n1480, n1481, n1482,
    n1483, n1484, n1485, n1486, n1487, n1488,
    n1489, n1490, n1491, n1492, n1493, n1494,
    n1495, n1496, n1497, n1498, n1499, n1500,
    n1501, n1502, n1503, n1504, n1505, n1506,
    n1507, n1508, n1509, n1510, n1511, n1512,
    n1513, n1514, n1515, n1516, n1517, n1518,
    n1519, n1520, n1521, n1522, n1523, n1524,
    n1525, n1526, n1527, n1528, n1529, n1530,
    n1531, n1532, n1533, n1534, n1535, n1536,
    n1537, n1538, n1539, n1540, n1541, n1542,
    n1543, n1544, n1545, n1546, n1547, n1548,
    n1549, n1550, n1551, n1552, n1553, n1554,
    n1555, n1556, n1557, n1558, n1559, n1560,
    n1561, n1562, n1563, n1564, n1565, n1566,
    n1567, n1568, n1569, n1570, n1571, n1572,
    n1574, n1575, n1576, n1577, n1578, n1579,
    n1580, n1581, n1582, n1583, n1584, n1585,
    n1586, n1587, n1588, n1589, n1590, n1591,
    n1592, n1593, n1594, n1595, n1596, n1597,
    n1598, n1599, n1600, n1601, n1602, n1603,
    n1604, n1605, n1606, n1607, n1608, n1609,
    n1610, n1611, n1612, n1613, n1614, n1615,
    n1616, n1617, n1618, n1619, n1620, n1621,
    n1622, n1623, n1624, n1625, n1626, n1627,
    n1628, n1629, n1630, n1631, n1632, n1633,
    n1634, n1635, n1636, n1637, n1638, n1639,
    n1640, n1641, n1642, n1643, n1644, n1645,
    n1646, n1647, n1648, n1649, n1650, n1651,
    n1652, n1653, n1654, n1655, n1656, n1657,
    n1658, n1659, n1660, n1661, n1662, n1663,
    n1664, n1665, n1666, n1667, n1668, n1669,
    n1670, n1671, n1672, n1673, n1674, n1675,
    n1676, n1677, n1678, n1679, n1680, n1681,
    n1682, n1683, n1684, n1685, n1686, n1687,
    n1688, n1689, n1690, n1691, n1692, n1693,
    n1694, n1695, n1696, n1697, n1698, n1699,
    n1700, n1701, n1702, n1703, n1704, n1705,
    n1706, n1707, n1708, n1709, n1710, n1711,
    n1712, n1713, n1714, n1716, n1717, n1718,
    n1719, n1720, n1721, n1722, n1723, n1724,
    n1725, n1726, n1727, n1728, n1729, n1730,
    n1731, n1732, n1733, n1734, n1735, n1736,
    n1737, n1738, n1739, n1740, n1741, n1742,
    n1743, n1744, n1745, n1746, n1747, n1748,
    n1749, n1750, n1751, n1752, n1753, n1754,
    n1755, n1756, n1757, n1758, n1759, n1760,
    n1761, n1762, n1763, n1764, n1765, n1766,
    n1767, n1768, n1769, n1770, n1771, n1772,
    n1773, n1774, n1775, n1776, n1777, n1778,
    n1779, n1780, n1781, n1782, n1783, n1784,
    n1785, n1786, n1787, n1788, n1789, n1790,
    n1791, n1792, n1793, n1794, n1795, n1796,
    n1797, n1798, n1799, n1800, n1801, n1802,
    n1803, n1804, n1805, n1806, n1807, n1808,
    n1809, n1810, n1811, n1812, n1813, n1814,
    n1815, n1816, n1817, n1818, n1819, n1820,
    n1821, n1822, n1823, n1824, n1825, n1826,
    n1827, n1828, n1829, n1830, n1831, n1832,
    n1833, n1834, n1835, n1836, n1837, n1838,
    n1839, n1840, n1841, n1842, n1843, n1844,
    n1845, n1846, n1847, n1848, n1849, n1850,
    n1851, n1852, n1854, n1855, n1856, n1857,
    n1858, n1859, n1860, n1861, n1862, n1863,
    n1864, n1865, n1866, n1867, n1868, n1869,
    n1870, n1871, n1872, n1873, n1874, n1875,
    n1876, n1877, n1878, n1879, n1880, n1881,
    n1882, n1883, n1884, n1885, n1886, n1887,
    n1888, n1889, n1890, n1891, n1892, n1893,
    n1894, n1895, n1896, n1897, n1898, n1899,
    n1900, n1901, n1902, n1903, n1904, n1905,
    n1906, n1907, n1908, n1909, n1910, n1911,
    n1912, n1913, n1914, n1915, n1916, n1917,
    n1918, n1919, n1920, n1921, n1922, n1923,
    n1924, n1925, n1926, n1927, n1928, n1929,
    n1930, n1931, n1932, n1933, n1934, n1935,
    n1936, n1937, n1938, n1939, n1940, n1941,
    n1942, n1943, n1944, n1945, n1946, n1947,
    n1948, n1949, n1950, n1951, n1952, n1953,
    n1954, n1955, n1956, n1957, n1958, n1959,
    n1960, n1961, n1962, n1963, n1964, n1965,
    n1966, n1967, n1968, n1969, n1970, n1971,
    n1972, n1973, n1974, n1975, n1976, n1977,
    n1978, n1979, n1980, n1981, n1982, n1983,
    n1984, n1985, n1986, n1987, n1988, n1989,
    n1990, n1992, n1993, n1994, n1995, n1996,
    n1997, n1998, n1999, n2000, n2001, n2002,
    n2003, n2004, n2005, n2006, n2007, n2008,
    n2009, n2010, n2011, n2012, n2013, n2014,
    n2015, n2016, n2017, n2018, n2019, n2020,
    n2021, n2022, n2023, n2024, n2025, n2026,
    n2027, n2028, n2029, n2030, n2031, n2032,
    n2033, n2034, n2035, n2036, n2037, n2038,
    n2039, n2040, n2041, n2042, n2043, n2044,
    n2045, n2046, n2047, n2048, n2049, n2050,
    n2051, n2052, n2053, n2054, n2055, n2056,
    n2057, n2058, n2059, n2060, n2061, n2062,
    n2063, n2064, n2065, n2066, n2067, n2068,
    n2069, n2070, n2071, n2072, n2073, n2074,
    n2075, n2076, n2077, n2078, n2079, n2080,
    n2081, n2082, n2083, n2084, n2085, n2086,
    n2087, n2088, n2089, n2090, n2091, n2092,
    n2093, n2094, n2095, n2096, n2097, n2098,
    n2099, n2100, n2101, n2102, n2103, n2104,
    n2105, n2106, n2107, n2108, n2109, n2110,
    n2111, n2112, n2113, n2114, n2115, n2116,
    n2117, n2118, n2119, n2120, n2121, n2122,
    n2123, n2124, n2125, n2126, n2127, n2128,
    n2129, n2130, n2131, n2132, n2133, n2134,
    n2135, n2136, n2137, n2138, n2139, n2140,
    n2141, n2142, n2143, n2144, n2145, n2146,
    n2147, n2148, n2149, n2151, n2152, n2153,
    n2154, n2155, n2156, n2157, n2158, n2159,
    n2160, n2161, n2162, n2163, n2164, n2165,
    n2166, n2167, n2168, n2169, n2170, n2171,
    n2172, n2173, n2174, n2175, n2176, n2177,
    n2178, n2179, n2180, n2181, n2182, n2183,
    n2184, n2185, n2186, n2187, n2188, n2189,
    n2190, n2191, n2192, n2193, n2194, n2195,
    n2196, n2197, n2198, n2199, n2200, n2201,
    n2202, n2203, n2204, n2205, n2206, n2207,
    n2208, n2209, n2210, n2211, n2212, n2213,
    n2214, n2215, n2216, n2217, n2218, n2219,
    n2220, n2221, n2222, n2223, n2224, n2225,
    n2226, n2227, n2228, n2229, n2230, n2231,
    n2232, n2233, n2234, n2235, n2236, n2237,
    n2238, n2239, n2240, n2241, n2242, n2243,
    n2244, n2245, n2246, n2247, n2248, n2249,
    n2250, n2251, n2252, n2253, n2254, n2255,
    n2256, n2257, n2258, n2259, n2260, n2261,
    n2262, n2263, n2264, n2265, n2266, n2267,
    n2268, n2269, n2270, n2271, n2272, n2273,
    n2274, n2275, n2276, n2277, n2278, n2279,
    n2280, n2281, n2282, n2283, n2284, n2285,
    n2286, n2287, n2288, n2289, n2290, n2291,
    n2292, n2293, n2294, n2295, n2296, n2297,
    n2298, n2299, n2300, n2301, n2302, n2303,
    n2304, n2305, n2306, n2308, n2309, n2310,
    n2311, n2312, n2313, n2314, n2315, n2316,
    n2317, n2318, n2319, n2320, n2321, n2322,
    n2323, n2324, n2325, n2326, n2327, n2328,
    n2329, n2330, n2331, n2332, n2333, n2334,
    n2335, n2336, n2337, n2338, n2339, n2340,
    n2341, n2342, n2343, n2344, n2345, n2346,
    n2347, n2348, n2349, n2350, n2351, n2352,
    n2353, n2354, n2355, n2356, n2357, n2358,
    n2359, n2360, n2361, n2362, n2363, n2364,
    n2365, n2366, n2367, n2368, n2369, n2370,
    n2371, n2372, n2373, n2374, n2375, n2376,
    n2377, n2378, n2379, n2380, n2381, n2382,
    n2383, n2384, n2385, n2386, n2387, n2388,
    n2389, n2390, n2391, n2392, n2393, n2394,
    n2395, n2396, n2397, n2398, n2399, n2400,
    n2401, n2402, n2403, n2404, n2405, n2406,
    n2407, n2408, n2409, n2410, n2411, n2412,
    n2413, n2414, n2415, n2416, n2417, n2418,
    n2419, n2420, n2421, n2422, n2423, n2424,
    n2425, n2426, n2427, n2428, n2429, n2430,
    n2431, n2432, n2433, n2434, n2435, n2436,
    n2437, n2438, n2439, n2440, n2441, n2442,
    n2443, n2444, n2445, n2446, n2447, n2448,
    n2449, n2450, n2451, n2452, n2453, n2454,
    n2455, n2456, n2457, n2458, n2459, n2460,
    n2461, n2462, n2463, n2464, n2466, n2467,
    n2468, n2469, n2470, n2471, n2472, n2473,
    n2474, n2475, n2476, n2477, n2478, n2479,
    n2480, n2481, n2482, n2483, n2484, n2485,
    n2486, n2487, n2488, n2489, n2490, n2491,
    n2492, n2493, n2494, n2495, n2496, n2497,
    n2498, n2499, n2500, n2501, n2502, n2503,
    n2504, n2505, n2506, n2507, n2508, n2509,
    n2510, n2511, n2512, n2513, n2514, n2515,
    n2516, n2517, n2518, n2519, n2520, n2521,
    n2522, n2523, n2524, n2525, n2526, n2527,
    n2528, n2529, n2530, n2531, n2532, n2533,
    n2534, n2535, n2536, n2537, n2538, n2539,
    n2540, n2541, n2542, n2543, n2544, n2545,
    n2546, n2547, n2548, n2549, n2550, n2551,
    n2552, n2553, n2554, n2555, n2556, n2557,
    n2558, n2559, n2560, n2561, n2562, n2563,
    n2564, n2565, n2566, n2567, n2568, n2569,
    n2570, n2571, n2572, n2573, n2574, n2575,
    n2576, n2577, n2578, n2579, n2580, n2581,
    n2582, n2583, n2584, n2585, n2586, n2587,
    n2588, n2589, n2590, n2591, n2592, n2593,
    n2594, n2595, n2596, n2597, n2598, n2599,
    n2600, n2601, n2602, n2603, n2604, n2605,
    n2606, n2607, n2608, n2609, n2610, n2611,
    n2612, n2613, n2614, n2615, n2616, n2617,
    n2618, n2619, n2620, n2621, n2622, n2623,
    n2624, n2625, n2626, n2627, n2628, n2629,
    n2630, n2631, n2632, n2633, n2634, n2635,
    n2636, n2637, n2638, n2639, n2640, n2641,
    n2642, n2643, n2645, n2646, n2647, n2648,
    n2649, n2650, n2651, n2652, n2653, n2654,
    n2655, n2656, n2657, n2658, n2659, n2660,
    n2661, n2662, n2663, n2664, n2665, n2666,
    n2667, n2668, n2669, n2670, n2671, n2672,
    n2673, n2674, n2675, n2676, n2677, n2678,
    n2679, n2680, n2681, n2682, n2683, n2684,
    n2685, n2686, n2687, n2688, n2689, n2690,
    n2691, n2692, n2693, n2694, n2695, n2696,
    n2697, n2698, n2699, n2700, n2701, n2702,
    n2703, n2704, n2705, n2706, n2707, n2708,
    n2709, n2710, n2711, n2712, n2713, n2714,
    n2715, n2716, n2717, n2718, n2719, n2720,
    n2721, n2722, n2723, n2724, n2725, n2726,
    n2727, n2728, n2729, n2730, n2731, n2732,
    n2733, n2734, n2735, n2736, n2737, n2738,
    n2739, n2740, n2741, n2742, n2743, n2744,
    n2745, n2746, n2747, n2748, n2749, n2750,
    n2751, n2752, n2753, n2754, n2755, n2756,
    n2757, n2758, n2759, n2760, n2761, n2762,
    n2763, n2764, n2765, n2766, n2767, n2768,
    n2769, n2770, n2771, n2772, n2773, n2774,
    n2775, n2776, n2777, n2778, n2779, n2780,
    n2781, n2782, n2783, n2784, n2785, n2786,
    n2787, n2788, n2789, n2790, n2791, n2792,
    n2793, n2794, n2795, n2796, n2797, n2798,
    n2799, n2800, n2801, n2802, n2803, n2804,
    n2805, n2806, n2807, n2808, n2809, n2810,
    n2811, n2812, n2813, n2814, n2815, n2816,
    n2817, n2819, n2820, n2821, n2822, n2823,
    n2824, n2825, n2826, n2827, n2828, n2829,
    n2830, n2831, n2832, n2833, n2834, n2835,
    n2836, n2837, n2838, n2839, n2840, n2841,
    n2842, n2843, n2844, n2845, n2846, n2847,
    n2848, n2849, n2850, n2851, n2852, n2853,
    n2854, n2855, n2856, n2857, n2858, n2859,
    n2860, n2861, n2862, n2863, n2864, n2865,
    n2866, n2867, n2868, n2869, n2870, n2871,
    n2872, n2873, n2874, n2875, n2876, n2877,
    n2878, n2879, n2880, n2881, n2882, n2883,
    n2884, n2885, n2886, n2887, n2888, n2889,
    n2890, n2891, n2892, n2893, n2894, n2895,
    n2896, n2897, n2898, n2899, n2900, n2901,
    n2902, n2903, n2904, n2905, n2906, n2907,
    n2908, n2909, n2910, n2911, n2912, n2913,
    n2914, n2915, n2916, n2917, n2918, n2919,
    n2920, n2921, n2922, n2923, n2924, n2925,
    n2926, n2927, n2928, n2929, n2930, n2931,
    n2932, n2933, n2934, n2935, n2936, n2937,
    n2938, n2939, n2940, n2941, n2942, n2943,
    n2944, n2945, n2946, n2947, n2948, n2949,
    n2950, n2951, n2952, n2953, n2954, n2955,
    n2956, n2957, n2958, n2959, n2960, n2961,
    n2962, n2963, n2964, n2965, n2966, n2967,
    n2968, n2969, n2970, n2971, n2972, n2973,
    n2974, n2975, n2976, n2977, n2978, n2979,
    n2980, n2981, n2982, n2983, n2984, n2985,
    n2986, n2987, n2988, n2989, n2990, n2991,
    n2992, n2993, n2994, n2996, n2997, n2998,
    n2999, n3000, n3001, n3002, n3003, n3004,
    n3005, n3006, n3007, n3008, n3009, n3010,
    n3011, n3012, n3013, n3014, n3015, n3016,
    n3017, n3018, n3019, n3020, n3021, n3022,
    n3023, n3024, n3025, n3026, n3027, n3028,
    n3029, n3030, n3031, n3032, n3033, n3034,
    n3035, n3036, n3037, n3038, n3039, n3040,
    n3041, n3042, n3043, n3044, n3045, n3046,
    n3047, n3048, n3049, n3050, n3051, n3052,
    n3053, n3054, n3055, n3056, n3057, n3058,
    n3059, n3060, n3061, n3062, n3063, n3064,
    n3065, n3066, n3067, n3068, n3069, n3070,
    n3071, n3072, n3073, n3074, n3075, n3076,
    n3077, n3078, n3079, n3080, n3081, n3082,
    n3083, n3084, n3085, n3086, n3087, n3088,
    n3089, n3090, n3091, n3092, n3093, n3094,
    n3095, n3096, n3097, n3098, n3099, n3100,
    n3101, n3102, n3103, n3104, n3105, n3106,
    n3107, n3108, n3109, n3110, n3111, n3112,
    n3113, n3114, n3115, n3116, n3117, n3118,
    n3119, n3120, n3121, n3122, n3123, n3124,
    n3125, n3126, n3127, n3128, n3129, n3130,
    n3131, n3132, n3133, n3134, n3135, n3136,
    n3137, n3138, n3139, n3140, n3141, n3142,
    n3143, n3144, n3145, n3146, n3147, n3148,
    n3149, n3150, n3151, n3152, n3153, n3154,
    n3155, n3156, n3157, n3158, n3159, n3160,
    n3161, n3162, n3163, n3164, n3165, n3166,
    n3167, n3168, n3169, n3170, n3171, n3172,
    n3173, n3174, n3175, n3176, n3177, n3178,
    n3179, n3180, n3181, n3182, n3183, n3184,
    n3185, n3186, n3187, n3188, n3189, n3190,
    n3191, n3192, n3193, n3195, n3196, n3197,
    n3198, n3199, n3200, n3201, n3202, n3203,
    n3204, n3205, n3206, n3207, n3208, n3209,
    n3210, n3211, n3212, n3213, n3214, n3215,
    n3216, n3217, n3218, n3219, n3220, n3221,
    n3222, n3223, n3224, n3225, n3226, n3227,
    n3228, n3229, n3230, n3231, n3232, n3233,
    n3234, n3235, n3236, n3237, n3238, n3239,
    n3240, n3241, n3242, n3243, n3244, n3245,
    n3246, n3247, n3248, n3249, n3250, n3251,
    n3252, n3253, n3254, n3255, n3256, n3257,
    n3258, n3259, n3260, n3261, n3262, n3263,
    n3264, n3265, n3266, n3267, n3268, n3269,
    n3270, n3271, n3272, n3273, n3274, n3275,
    n3276, n3277, n3278, n3279, n3280, n3281,
    n3282, n3283, n3284, n3285, n3286, n3287,
    n3288, n3289, n3290, n3291, n3292, n3293,
    n3294, n3295, n3296, n3297, n3298, n3299,
    n3300, n3301, n3302, n3303, n3304, n3305,
    n3306, n3307, n3308, n3309, n3310, n3311,
    n3312, n3313, n3314, n3315, n3316, n3317,
    n3318, n3319, n3320, n3321, n3322, n3323,
    n3324, n3325, n3326, n3327, n3328, n3329,
    n3330, n3331, n3332, n3333, n3334, n3335,
    n3336, n3337, n3338, n3339, n3340, n3341,
    n3342, n3343, n3344, n3345, n3346, n3347,
    n3348, n3349, n3350, n3351, n3352, n3353,
    n3354, n3355, n3356, n3357, n3358, n3359,
    n3360, n3361, n3362, n3363, n3364, n3365,
    n3366, n3367, n3368, n3369, n3370, n3371,
    n3372, n3373, n3374, n3375, n3376, n3377,
    n3378, n3379, n3380, n3381, n3382, n3383,
    n3384, n3385, n3386, n3387, n3388, n3389,
    n3391, n3392, n3393, n3394, n3395, n3396,
    n3397, n3398, n3399, n3400, n3401, n3402,
    n3403, n3404, n3405, n3406, n3407, n3408,
    n3409, n3410, n3411, n3412, n3413, n3414,
    n3415, n3416, n3417, n3418, n3419, n3420,
    n3421, n3422, n3423, n3424, n3425, n3426,
    n3427, n3428, n3429, n3430, n3431, n3432,
    n3433, n3434, n3435, n3436, n3437, n3438,
    n3439, n3440, n3441, n3442, n3443, n3444,
    n3445, n3446, n3447, n3448, n3449, n3450,
    n3451, n3452, n3453, n3454, n3455, n3456,
    n3457, n3458, n3459, n3460, n3461, n3462,
    n3463, n3464, n3465, n3466, n3467, n3468,
    n3469, n3470, n3471, n3472, n3473, n3474,
    n3475, n3476, n3477, n3478, n3479, n3480,
    n3481, n3482, n3483, n3484, n3485, n3486,
    n3487, n3488, n3489, n3490, n3491, n3492,
    n3493, n3494, n3495, n3496, n3497, n3498,
    n3499, n3500, n3501, n3502, n3503, n3504,
    n3505, n3506, n3507, n3508, n3509, n3510,
    n3511, n3512, n3513, n3514, n3515, n3516,
    n3517, n3518, n3519, n3520, n3521, n3522,
    n3523, n3524, n3525, n3526, n3527, n3528,
    n3529, n3530, n3531, n3532, n3533, n3534,
    n3535, n3536, n3537, n3538, n3539, n3540,
    n3541, n3542, n3543, n3544, n3545, n3546,
    n3547, n3548, n3549, n3550, n3551, n3552,
    n3553, n3554, n3555, n3556, n3557, n3558,
    n3559, n3560, n3561, n3562, n3563, n3564,
    n3565, n3566, n3567, n3568, n3569, n3570,
    n3571, n3572, n3573, n3574, n3575, n3576,
    n3577, n3578, n3579, n3580, n3581, n3582,
    n3583, n3585, n3586, n3587, n3588, n3589,
    n3590, n3591, n3592, n3593, n3594, n3595,
    n3596, n3597, n3598, n3599, n3600, n3601,
    n3602, n3603, n3604, n3605, n3606, n3607,
    n3608, n3609, n3610, n3611, n3612, n3613,
    n3614, n3615, n3616, n3617, n3618, n3619,
    n3620, n3621, n3622, n3623, n3624, n3625,
    n3626, n3627, n3628, n3629, n3630, n3631,
    n3632, n3633, n3634, n3635, n3636, n3637,
    n3638, n3639, n3640, n3641, n3642, n3643,
    n3644, n3645, n3646, n3647, n3648, n3649,
    n3650, n3651, n3652, n3653, n3654, n3655,
    n3656, n3657, n3658, n3659, n3660, n3661,
    n3662, n3663, n3664, n3665, n3666, n3667,
    n3668, n3669, n3670, n3671, n3672, n3673,
    n3674, n3675, n3676, n3677, n3678, n3679,
    n3680, n3681, n3682, n3683, n3684, n3685,
    n3686, n3687, n3688, n3689, n3690, n3691,
    n3692, n3693, n3694, n3695, n3696, n3697,
    n3698, n3699, n3700, n3701, n3702, n3703,
    n3704, n3705, n3706, n3707, n3708, n3709,
    n3710, n3711, n3712, n3713, n3714, n3715,
    n3716, n3717, n3718, n3719, n3720, n3721,
    n3722, n3723, n3724, n3725, n3726, n3727,
    n3728, n3729, n3730, n3731, n3732, n3733,
    n3734, n3735, n3736, n3737, n3738, n3739,
    n3740, n3741, n3742, n3743, n3744, n3745,
    n3746, n3747, n3748, n3749, n3750, n3751,
    n3752, n3753, n3754, n3755, n3756, n3757,
    n3758, n3759, n3760, n3761, n3762, n3763,
    n3764, n3765, n3766, n3767, n3768, n3769,
    n3770, n3771, n3772, n3773, n3774, n3775,
    n3776, n3777, n3778, n3779, n3780, n3781,
    n3782, n3783, n3784, n3785, n3786, n3787,
    n3788, n3789, n3790, n3791, n3792, n3793,
    n3794, n3795, n3796, n3797, n3798, n3799,
    n3800, n3801, n3802, n3804, n3805, n3806,
    n3807, n3808, n3809, n3810, n3811, n3812,
    n3813, n3814, n3815, n3816, n3817, n3818,
    n3819, n3820, n3821, n3822, n3823, n3824,
    n3825, n3826, n3827, n3828, n3829, n3830,
    n3831, n3832, n3833, n3834, n3835, n3836,
    n3837, n3838, n3839, n3840, n3841, n3842,
    n3843, n3844, n3845, n3846, n3847, n3848,
    n3849, n3850, n3851, n3852, n3853, n3854,
    n3855, n3856, n3857, n3858, n3859, n3860,
    n3861, n3862, n3863, n3864, n3865, n3866,
    n3867, n3868, n3869, n3870, n3871, n3872,
    n3873, n3874, n3875, n3876, n3877, n3878,
    n3879, n3880, n3881, n3882, n3883, n3884,
    n3885, n3886, n3887, n3888, n3889, n3890,
    n3891, n3892, n3893, n3894, n3895, n3896,
    n3897, n3898, n3899, n3900, n3901, n3902,
    n3903, n3904, n3905, n3906, n3907, n3908,
    n3909, n3910, n3911, n3912, n3913, n3914,
    n3915, n3916, n3917, n3918, n3919, n3920,
    n3921, n3922, n3923, n3924, n3925, n3926,
    n3927, n3928, n3929, n3930, n3931, n3932,
    n3933, n3934, n3935, n3936, n3937, n3938,
    n3939, n3940, n3941, n3942, n3943, n3944,
    n3945, n3946, n3947, n3948, n3949, n3950,
    n3951, n3952, n3953, n3954, n3955, n3956,
    n3957, n3958, n3959, n3960, n3961, n3962,
    n3963, n3964, n3965, n3966, n3967, n3968,
    n3969, n3970, n3971, n3972, n3973, n3974,
    n3975, n3976, n3977, n3978, n3979, n3980,
    n3981, n3982, n3983, n3984, n3985, n3986,
    n3987, n3988, n3989, n3990, n3991, n3992,
    n3993, n3994, n3995, n3996, n3997, n3998,
    n3999, n4000, n4001, n4002, n4003, n4004,
    n4005, n4006, n4007, n4008, n4009, n4010,
    n4011, n4012, n4013, n4014, n4015, n4016,
    n4017, n4019, n4020, n4021, n4022, n4023,
    n4024, n4025, n4026, n4027, n4028, n4029,
    n4030, n4031, n4032, n4033, n4034, n4035,
    n4036, n4037, n4038, n4039, n4040, n4041,
    n4042, n4043, n4044, n4045, n4046, n4047,
    n4048, n4049, n4050, n4051, n4052, n4053,
    n4054, n4055, n4056, n4057, n4058, n4059,
    n4060, n4061, n4062, n4063, n4064, n4065,
    n4066, n4067, n4068, n4069, n4070, n4071,
    n4072, n4073, n4074, n4075, n4076, n4077,
    n4078, n4079, n4080, n4081, n4082, n4083,
    n4084, n4085, n4086, n4087, n4088, n4089,
    n4090, n4091, n4092, n4093, n4094, n4095,
    n4096, n4097, n4098, n4099, n4100, n4101,
    n4102, n4103, n4104, n4105, n4106, n4107,
    n4108, n4109, n4110, n4111, n4112, n4113,
    n4114, n4115, n4116, n4117, n4118, n4119,
    n4120, n4121, n4122, n4123, n4124, n4125,
    n4126, n4127, n4128, n4129, n4130, n4131,
    n4132, n4133, n4134, n4135, n4136, n4137,
    n4138, n4139, n4140, n4141, n4142, n4143,
    n4144, n4145, n4146, n4147, n4148, n4149,
    n4150, n4151, n4152, n4153, n4154, n4155,
    n4156, n4157, n4158, n4159, n4160, n4161,
    n4162, n4163, n4164, n4165, n4166, n4167,
    n4168, n4169, n4170, n4171, n4172, n4173,
    n4174, n4175, n4176, n4177, n4178, n4179,
    n4180, n4181, n4182, n4183, n4184, n4185,
    n4186, n4187, n4188, n4189, n4190, n4191,
    n4192, n4193, n4194, n4195, n4196, n4197,
    n4198, n4199, n4200, n4201, n4202, n4203,
    n4204, n4205, n4206, n4207, n4208, n4209,
    n4210, n4211, n4212, n4213, n4214, n4215,
    n4216, n4217, n4218, n4219, n4220, n4221,
    n4222, n4223, n4224, n4225, n4226, n4227,
    n4229, n4230, n4231, n4232, n4233, n4234,
    n4235, n4236, n4237, n4238, n4239, n4240,
    n4241, n4242, n4243, n4244, n4245, n4246,
    n4247, n4248, n4249, n4250, n4251, n4252,
    n4253, n4254, n4255, n4256, n4257, n4258,
    n4259, n4260, n4261, n4262, n4263, n4264,
    n4265, n4266, n4267, n4268, n4269, n4270,
    n4271, n4272, n4273, n4274, n4275, n4276,
    n4277, n4278, n4279, n4280, n4281, n4282,
    n4283, n4284, n4285, n4286, n4287, n4288,
    n4289, n4290, n4291, n4292, n4293, n4294,
    n4295, n4296, n4297, n4298, n4299, n4300,
    n4301, n4302, n4303, n4304, n4305, n4306,
    n4307, n4308, n4309, n4310, n4311, n4312,
    n4313, n4314, n4315, n4316, n4317, n4318,
    n4319, n4320, n4321, n4322, n4323, n4324,
    n4325, n4326, n4327, n4328, n4329, n4330,
    n4331, n4332, n4333, n4334, n4335, n4336,
    n4337, n4338, n4339, n4340, n4341, n4342,
    n4343, n4344, n4345, n4346, n4347, n4348,
    n4349, n4350, n4351, n4352, n4353, n4354,
    n4355, n4356, n4357, n4358, n4359, n4360,
    n4361, n4362, n4363, n4364, n4365, n4366,
    n4367, n4368, n4369, n4370, n4371, n4372,
    n4373, n4374, n4375, n4376, n4377, n4378,
    n4379, n4380, n4381, n4382, n4383, n4384,
    n4385, n4386, n4387, n4388, n4389, n4390,
    n4391, n4392, n4393, n4394, n4395, n4396,
    n4397, n4398, n4399, n4400, n4401, n4402,
    n4403, n4404, n4405, n4406, n4407, n4408,
    n4409, n4410, n4411, n4412, n4413, n4414,
    n4415, n4416, n4417, n4418, n4419, n4420,
    n4421, n4422, n4423, n4424, n4425, n4426,
    n4427, n4428, n4429, n4430, n4431, n4432,
    n4433, n4434, n4435, n4436, n4437, n4438,
    n4439, n4440, n4441, n4442, n4443, n4444,
    n4445, n4446, n4447, n4448, n4449, n4450,
    n4451, n4452, n4453, n4454, n4455, n4456,
    n4457, n4458, n4459, n4460, n4461, n4462,
    n4463, n4464, n4465, n4466, n4467, n4468,
    n4469, n4470, n4472, n4473, n4474, n4475,
    n4476, n4477, n4478, n4479, n4480, n4481,
    n4482, n4483, n4484, n4485, n4486, n4487,
    n4488, n4489, n4490, n4491, n4492, n4493,
    n4494, n4495, n4496, n4497, n4498, n4499,
    n4500, n4501, n4502, n4503, n4504, n4505,
    n4506, n4507, n4508, n4509, n4510, n4511,
    n4512, n4513, n4514, n4515, n4516, n4517,
    n4518, n4519, n4520, n4521, n4522, n4523,
    n4524, n4525, n4526, n4527, n4528, n4529,
    n4530, n4531, n4532, n4533, n4534, n4535,
    n4536, n4537, n4538, n4539, n4540, n4541,
    n4542, n4543, n4544, n4545, n4546, n4547,
    n4548, n4549, n4550, n4551, n4552, n4553,
    n4554, n4555, n4556, n4557, n4558, n4559,
    n4560, n4561, n4562, n4563, n4564, n4565,
    n4566, n4567, n4568, n4569, n4570, n4571,
    n4572, n4573, n4574, n4575, n4576, n4577,
    n4578, n4579, n4580, n4581, n4582, n4583,
    n4584, n4585, n4586, n4587, n4588, n4589,
    n4590, n4591, n4592, n4593, n4594, n4595,
    n4596, n4597, n4598, n4599, n4600, n4601,
    n4602, n4603, n4604, n4605, n4606, n4607,
    n4608, n4609, n4610, n4611, n4612, n4613,
    n4614, n4615, n4616, n4617, n4618, n4619,
    n4620, n4621, n4622, n4623, n4624, n4625,
    n4626, n4627, n4628, n4629, n4630, n4631,
    n4632, n4633, n4634, n4635, n4636, n4637,
    n4638, n4639, n4640, n4641, n4642, n4643,
    n4644, n4645, n4646, n4647, n4648, n4649,
    n4650, n4651, n4652, n4653, n4654, n4655,
    n4656, n4657, n4658, n4659, n4660, n4661,
    n4662, n4663, n4664, n4665, n4666, n4667,
    n4668, n4669, n4670, n4671, n4672, n4673,
    n4674, n4675, n4676, n4677, n4678, n4679,
    n4680, n4681, n4682, n4683, n4684, n4685,
    n4686, n4687, n4688, n4689, n4690, n4691,
    n4692, n4693, n4694, n4695, n4696, n4697,
    n4698, n4699, n4700, n4702, n4703, n4704,
    n4705, n4706, n4707, n4708, n4709, n4710,
    n4711, n4712, n4713, n4714, n4715, n4716,
    n4717, n4718, n4719, n4720, n4721, n4722,
    n4723, n4724, n4725, n4726, n4727, n4728,
    n4729, n4730, n4731, n4732, n4733, n4734,
    n4735, n4736, n4737, n4738, n4739, n4740,
    n4741, n4742, n4743, n4744, n4745, n4746,
    n4747, n4748, n4749, n4750, n4751, n4752,
    n4753, n4754, n4755, n4756, n4757, n4758,
    n4759, n4760, n4761, n4762, n4763, n4764,
    n4765, n4766, n4767, n4768, n4769, n4770,
    n4771, n4772, n4773, n4774, n4775, n4776,
    n4777, n4778, n4779, n4780, n4781, n4782,
    n4783, n4784, n4785, n4786, n4787, n4788,
    n4789, n4790, n4791, n4792, n4793, n4794,
    n4795, n4796, n4797, n4798, n4799, n4800,
    n4801, n4802, n4803, n4804, n4805, n4806,
    n4807, n4808, n4809, n4810, n4811, n4812,
    n4813, n4814, n4815, n4816, n4817, n4818,
    n4819, n4820, n4821, n4822, n4823, n4824,
    n4825, n4826, n4827, n4828, n4829, n4830,
    n4831, n4832, n4833, n4834, n4835, n4836,
    n4837, n4838, n4839, n4840, n4841, n4842,
    n4843, n4844, n4845, n4846, n4847, n4848,
    n4849, n4850, n4851, n4852, n4853, n4854,
    n4855, n4856, n4857, n4858, n4859, n4860,
    n4861, n4862, n4863, n4864, n4865, n4866,
    n4867, n4868, n4869, n4870, n4871, n4872,
    n4873, n4874, n4875, n4876, n4877, n4878,
    n4879, n4880, n4881, n4882, n4883, n4884,
    n4885, n4886, n4887, n4888, n4889, n4890,
    n4891, n4892, n4893, n4894, n4895, n4896,
    n4897, n4898, n4899, n4900, n4901, n4902,
    n4903, n4904, n4905, n4906, n4907, n4908,
    n4909, n4910, n4911, n4912, n4913, n4914,
    n4915, n4916, n4917, n4918, n4919, n4920,
    n4921, n4922, n4923, n4924, n4925, n4926,
    n4927, n4928, n4929, n4931, n4932, n4933,
    n4934, n4935, n4936, n4937, n4938, n4939,
    n4940, n4941, n4942, n4943, n4944, n4945,
    n4946, n4947, n4948, n4949, n4950, n4951,
    n4952, n4953, n4954, n4955, n4956, n4957,
    n4958, n4959, n4960, n4961, n4962, n4963,
    n4964, n4965, n4966, n4967, n4968, n4969,
    n4970, n4971, n4972, n4973, n4974, n4975,
    n4976, n4977, n4978, n4979, n4980, n4981,
    n4982, n4983, n4984, n4985, n4986, n4987,
    n4988, n4989, n4990, n4991, n4992, n4993,
    n4994, n4995, n4996, n4997, n4998, n4999,
    n5000, n5001, n5002, n5003, n5004, n5005,
    n5006, n5007, n5008, n5009, n5010, n5011,
    n5012, n5013, n5014, n5015, n5016, n5017,
    n5018, n5019, n5020, n5021, n5022, n5023,
    n5024, n5025, n5026, n5027, n5028, n5029,
    n5030, n5031, n5032, n5033, n5034, n5035,
    n5036, n5037, n5038, n5039, n5040, n5041,
    n5042, n5043, n5044, n5045, n5046, n5047,
    n5048, n5049, n5050, n5051, n5052, n5053,
    n5054, n5055, n5056, n5057, n5058, n5059,
    n5060, n5061, n5062, n5063, n5064, n5065,
    n5066, n5067, n5068, n5069, n5070, n5071,
    n5072, n5073, n5074, n5075, n5076, n5077,
    n5078, n5079, n5080, n5081, n5082, n5083,
    n5084, n5085, n5086, n5087, n5088, n5089,
    n5090, n5091, n5092, n5093, n5094, n5095,
    n5096, n5097, n5098, n5099, n5100, n5101,
    n5102, n5103, n5104, n5105, n5106, n5107,
    n5108, n5109, n5110, n5111, n5112, n5113,
    n5114, n5115, n5116, n5117, n5118, n5119,
    n5120, n5121, n5122, n5123, n5124, n5125,
    n5126, n5127, n5128, n5129, n5130, n5131,
    n5132, n5133, n5134, n5135, n5136, n5137,
    n5138, n5139, n5140, n5141, n5142, n5143,
    n5144, n5145, n5146, n5147, n5148, n5149,
    n5150, n5151, n5152, n5153, n5154, n5155,
    n5156, n5157, n5158, n5159, n5160, n5161,
    n5162, n5163, n5164, n5165, n5166, n5167,
    n5168, n5169, n5170, n5171, n5172, n5173,
    n5174, n5175, n5176, n5177, n5178, n5179,
    n5180, n5181, n5182, n5183, n5184, n5185,
    n5187, n5188, n5189, n5190, n5191, n5192,
    n5193, n5194, n5195, n5196, n5197, n5198,
    n5199, n5200, n5201, n5202, n5203, n5204,
    n5205, n5206, n5207, n5208, n5209, n5210,
    n5211, n5212, n5213, n5214, n5215, n5216,
    n5217, n5218, n5219, n5220, n5221, n5222,
    n5223, n5224, n5225, n5226, n5227, n5228,
    n5229, n5230, n5231, n5232, n5233, n5234,
    n5235, n5236, n5237, n5238, n5239, n5240,
    n5241, n5242, n5243, n5244, n5245, n5246,
    n5247, n5248, n5249, n5250, n5251, n5252,
    n5253, n5254, n5255, n5256, n5257, n5258,
    n5259, n5260, n5261, n5262, n5263, n5264,
    n5265, n5266, n5267, n5268, n5269, n5270,
    n5271, n5272, n5273, n5274, n5275, n5276,
    n5277, n5278, n5279, n5280, n5281, n5282,
    n5283, n5284, n5285, n5286, n5287, n5288,
    n5289, n5290, n5291, n5292, n5293, n5294,
    n5295, n5296, n5297, n5298, n5299, n5300,
    n5301, n5302, n5303, n5304, n5305, n5306,
    n5307, n5308, n5309, n5310, n5311, n5312,
    n5313, n5314, n5315, n5316, n5317, n5318,
    n5319, n5320, n5321, n5322, n5323, n5324,
    n5325, n5326, n5327, n5328, n5329, n5330,
    n5331, n5332, n5333, n5334, n5335, n5336,
    n5337, n5338, n5339, n5340, n5341, n5342,
    n5343, n5344, n5345, n5346, n5347, n5348,
    n5349, n5350, n5351, n5352, n5353, n5354,
    n5355, n5356, n5357, n5358, n5359, n5360,
    n5361, n5362, n5363, n5364, n5365, n5366,
    n5367, n5368, n5369, n5370, n5371, n5372,
    n5373, n5374, n5375, n5376, n5377, n5378,
    n5379, n5380, n5381, n5382, n5383, n5384,
    n5385, n5386, n5387, n5388, n5389, n5390,
    n5391, n5392, n5393, n5394, n5395, n5396,
    n5397, n5398, n5399, n5400, n5401, n5402,
    n5403, n5404, n5405, n5406, n5407, n5408,
    n5409, n5410, n5411, n5412, n5413, n5414,
    n5415, n5416, n5417, n5418, n5419, n5420,
    n5421, n5422, n5423, n5424, n5425, n5426,
    n5427, n5428, n5429, n5430, n5431, n5433,
    n5434, n5435, n5436, n5437, n5438, n5439,
    n5440, n5441, n5442, n5443, n5444, n5445,
    n5446, n5447, n5448, n5449, n5450, n5451,
    n5452, n5453, n5454, n5455, n5456, n5457,
    n5458, n5459, n5460, n5461, n5462, n5463,
    n5464, n5465, n5466, n5467, n5468, n5469,
    n5470, n5471, n5472, n5473, n5474, n5475,
    n5476, n5477, n5478, n5479, n5480, n5481,
    n5482, n5483, n5484, n5485, n5486, n5487,
    n5488, n5489, n5490, n5491, n5492, n5493,
    n5494, n5495, n5496, n5497, n5498, n5499,
    n5500, n5501, n5502, n5503, n5504, n5505,
    n5506, n5507, n5508, n5509, n5510, n5511,
    n5512, n5513, n5514, n5515, n5516, n5517,
    n5518, n5519, n5520, n5521, n5522, n5523,
    n5524, n5525, n5526, n5527, n5528, n5529,
    n5530, n5531, n5532, n5533, n5534, n5535,
    n5536, n5537, n5538, n5539, n5540, n5541,
    n5542, n5543, n5544, n5545, n5546, n5547,
    n5548, n5549, n5550, n5551, n5552, n5553,
    n5554, n5555, n5556, n5557, n5558, n5559,
    n5560, n5561, n5562, n5563, n5564, n5565,
    n5566, n5567, n5568, n5569, n5570, n5571,
    n5572, n5573, n5574, n5575, n5576, n5577,
    n5578, n5579, n5580, n5581, n5582, n5583,
    n5584, n5585, n5586, n5587, n5588, n5589,
    n5590, n5591, n5592, n5593, n5594, n5595,
    n5596, n5597, n5598, n5599, n5600, n5601,
    n5602, n5603, n5604, n5605, n5606, n5607,
    n5608, n5609, n5610, n5611, n5612, n5613,
    n5614, n5615, n5616, n5617, n5618, n5619,
    n5620, n5621, n5622, n5623, n5624, n5625,
    n5626, n5627, n5628, n5629, n5630, n5631,
    n5632, n5633, n5634, n5635, n5636, n5637,
    n5638, n5639, n5640, n5641, n5642, n5643,
    n5644, n5645, n5646, n5647, n5648, n5649,
    n5650, n5651, n5652, n5653, n5654, n5655,
    n5656, n5657, n5658, n5659, n5660, n5661,
    n5662, n5663, n5664, n5665, n5666, n5667,
    n5668, n5669, n5670, n5671, n5672, n5673,
    n5674, n5675, n5676, n5677, n5678, n5679,
    n5680, n5681, n5682, n5684, n5685, n5686,
    n5687, n5688, n5689, n5690, n5691, n5692,
    n5693, n5694, n5695, n5696, n5697, n5698,
    n5699, n5700, n5701, n5702, n5703, n5704,
    n5705, n5706, n5707, n5708, n5709, n5710,
    n5711, n5712, n5713, n5714, n5715, n5716,
    n5717, n5718, n5719, n5720, n5721, n5722,
    n5723, n5724, n5725, n5726, n5727, n5728,
    n5729, n5730, n5731, n5732, n5733, n5734,
    n5735, n5736, n5737, n5738, n5739, n5740,
    n5741, n5742, n5743, n5744, n5745, n5746,
    n5747, n5748, n5749, n5750, n5751, n5752,
    n5753, n5754, n5755, n5756, n5757, n5758,
    n5759, n5760, n5761, n5762, n5763, n5764,
    n5765, n5766, n5767, n5768, n5769, n5770,
    n5771, n5772, n5773, n5774, n5775, n5776,
    n5777, n5778, n5779, n5780, n5781, n5782,
    n5783, n5784, n5785, n5786, n5787, n5788,
    n5789, n5790, n5791, n5792, n5793, n5794,
    n5795, n5796, n5797, n5798, n5799, n5800,
    n5801, n5802, n5803, n5804, n5805, n5806,
    n5807, n5808, n5809, n5810, n5811, n5812,
    n5813, n5814, n5815, n5816, n5817, n5818,
    n5819, n5820, n5821, n5822, n5823, n5824,
    n5825, n5826, n5827, n5828, n5829, n5830,
    n5831, n5832, n5833, n5834, n5835, n5836,
    n5837, n5838, n5839, n5840, n5841, n5842,
    n5843, n5844, n5845, n5846, n5847, n5848,
    n5849, n5850, n5851, n5852, n5853, n5854,
    n5855, n5856, n5857, n5858, n5859, n5860,
    n5861, n5862, n5863, n5864, n5865, n5866,
    n5867, n5868, n5869, n5870, n5871, n5872,
    n5873, n5874, n5875, n5876, n5877, n5878,
    n5879, n5880, n5881, n5882, n5883, n5884,
    n5885, n5886, n5887, n5888, n5889, n5890,
    n5891, n5892, n5893, n5894, n5895, n5896,
    n5897, n5898, n5899, n5900, n5901, n5902,
    n5903, n5904, n5905, n5906, n5907, n5908,
    n5909, n5910, n5911, n5912, n5913, n5914,
    n5915, n5916, n5917, n5918, n5919, n5920,
    n5921, n5922, n5923, n5924, n5925, n5926,
    n5927, n5928, n5929, n5930, n5931, n5932,
    n5933, n5934, n5935, n5936, n5937, n5938,
    n5939, n5940, n5941, n5942, n5943, n5944,
    n5945, n5946, n5947, n5948, n5949, n5950,
    n5951, n5952, n5953, n5954, n5955, n5956,
    n5957, n5958, n5959, n5961, n5962, n5963,
    n5964, n5965, n5966, n5967, n5968, n5969,
    n5970, n5971, n5972, n5973, n5974, n5975,
    n5976, n5977, n5978, n5979, n5980, n5981,
    n5982, n5983, n5984, n5985, n5986, n5987,
    n5988, n5989, n5990, n5991, n5992, n5993,
    n5994, n5995, n5996, n5997, n5998, n5999,
    n6000, n6001, n6002, n6003, n6004, n6005,
    n6006, n6007, n6008, n6009, n6010, n6011,
    n6012, n6013, n6014, n6015, n6016, n6017,
    n6018, n6019, n6020, n6021, n6022, n6023,
    n6024, n6025, n6026, n6027, n6028, n6029,
    n6030, n6031, n6032, n6033, n6034, n6035,
    n6036, n6037, n6038, n6039, n6040, n6041,
    n6042, n6043, n6044, n6045, n6046, n6047,
    n6048, n6049, n6050, n6051, n6052, n6053,
    n6054, n6055, n6056, n6057, n6058, n6059,
    n6060, n6061, n6062, n6063, n6064, n6065,
    n6066, n6067, n6068, n6069, n6070, n6071,
    n6072, n6073, n6074, n6075, n6076, n6077,
    n6078, n6079, n6080, n6081, n6082, n6083,
    n6084, n6085, n6086, n6087, n6088, n6089,
    n6090, n6091, n6092, n6093, n6094, n6095,
    n6096, n6097, n6098, n6099, n6100, n6101,
    n6102, n6103, n6104, n6105, n6106, n6107,
    n6108, n6109, n6110, n6111, n6112, n6113,
    n6114, n6115, n6116, n6117, n6118, n6119,
    n6120, n6121, n6122, n6123, n6124, n6125,
    n6126, n6127, n6128, n6129, n6130, n6131,
    n6132, n6133, n6134, n6135, n6136, n6137,
    n6138, n6139, n6140, n6141, n6142, n6143,
    n6144, n6145, n6146, n6147, n6148, n6149,
    n6150, n6151, n6152, n6153, n6154, n6155,
    n6156, n6157, n6158, n6159, n6160, n6161,
    n6162, n6163, n6164, n6165, n6166, n6167,
    n6168, n6169, n6170, n6171, n6172, n6173,
    n6174, n6175, n6176, n6177, n6178, n6179,
    n6180, n6181, n6182, n6183, n6184, n6185,
    n6186, n6187, n6188, n6189, n6190, n6191,
    n6192, n6193, n6194, n6195, n6196, n6197,
    n6198, n6199, n6200, n6201, n6202, n6203,
    n6204, n6205, n6206, n6207, n6208, n6209,
    n6210, n6211, n6212, n6213, n6214, n6215,
    n6216, n6217, n6218, n6219, n6220, n6221,
    n6222, n6223, n6225, n6226, n6227, n6228,
    n6229, n6230, n6231, n6232, n6233, n6234,
    n6235, n6236, n6237, n6238, n6239, n6240,
    n6241, n6242, n6243, n6244, n6245, n6246,
    n6247, n6248, n6249, n6250, n6251, n6252,
    n6253, n6254, n6255, n6256, n6257, n6258,
    n6259, n6260, n6261, n6262, n6263, n6264,
    n6265, n6266, n6267, n6268, n6269, n6270,
    n6271, n6272, n6273, n6274, n6275, n6276,
    n6277, n6278, n6279, n6280, n6281, n6282,
    n6283, n6284, n6285, n6286, n6287, n6288,
    n6289, n6290, n6291, n6292, n6293, n6294,
    n6295, n6296, n6297, n6298, n6299, n6300,
    n6301, n6302, n6303, n6304, n6305, n6306,
    n6307, n6308, n6309, n6310, n6311, n6312,
    n6313, n6314, n6315, n6316, n6317, n6318,
    n6319, n6320, n6321, n6322, n6323, n6324,
    n6325, n6326, n6327, n6328, n6329, n6330,
    n6331, n6332, n6333, n6334, n6335, n6336,
    n6337, n6338, n6339, n6340, n6341, n6342,
    n6343, n6344, n6345, n6346, n6347, n6348,
    n6349, n6350, n6351, n6352, n6353, n6354,
    n6355, n6356, n6357, n6358, n6359, n6360,
    n6361, n6362, n6363, n6364, n6365, n6366,
    n6367, n6368, n6369, n6370, n6371, n6372,
    n6373, n6374, n6375, n6376, n6377, n6378,
    n6379, n6380, n6381, n6382, n6383, n6384,
    n6385, n6386, n6387, n6388, n6389, n6390,
    n6391, n6392, n6393, n6394, n6395, n6396,
    n6397, n6398, n6399, n6400, n6401, n6402,
    n6403, n6404, n6405, n6406, n6407, n6408,
    n6409, n6410, n6411, n6412, n6413, n6414,
    n6415, n6416, n6417, n6418, n6419, n6420,
    n6421, n6422, n6423, n6424, n6425, n6426,
    n6427, n6428, n6429, n6430, n6431, n6432,
    n6433, n6434, n6435, n6436, n6437, n6438,
    n6439, n6440, n6441, n6442, n6443, n6444,
    n6445, n6446, n6447, n6448, n6449, n6450,
    n6451, n6452, n6453, n6454, n6455, n6456,
    n6457, n6458, n6459, n6460, n6461, n6462,
    n6463, n6464, n6465, n6466, n6467, n6468,
    n6469, n6470, n6471, n6472, n6473, n6474,
    n6475, n6476, n6477, n6478, n6479, n6480,
    n6481, n6482, n6483, n6484, n6485, n6486,
    n6487, n6488, n6489, n6490, n6491, n6492,
    n6493, n6494, n6495, n6497, n6498, n6499,
    n6500, n6501, n6502, n6503, n6504, n6505,
    n6506, n6507, n6508, n6509, n6510, n6511,
    n6512, n6513, n6514, n6515, n6516, n6517,
    n6518, n6519, n6520, n6521, n6522, n6523,
    n6524, n6525, n6526, n6527, n6528, n6529,
    n6530, n6531, n6532, n6533, n6534, n6535,
    n6536, n6537, n6538, n6539, n6540, n6541,
    n6542, n6543, n6544, n6545, n6546, n6547,
    n6548, n6549, n6550, n6551, n6552, n6553,
    n6554, n6555, n6556, n6557, n6558, n6559,
    n6560, n6561, n6562, n6563, n6564, n6565,
    n6566, n6567, n6568, n6569, n6570, n6571,
    n6572, n6573, n6574, n6575, n6576, n6577,
    n6578, n6579, n6580, n6581, n6582, n6583,
    n6584, n6585, n6586, n6587, n6588, n6589,
    n6590, n6591, n6592, n6593, n6594, n6595,
    n6596, n6597, n6598, n6599, n6600, n6601,
    n6602, n6603, n6604, n6605, n6606, n6607,
    n6608, n6609, n6610, n6611, n6612, n6613,
    n6614, n6615, n6616, n6617, n6618, n6619,
    n6620, n6621, n6622, n6623, n6624, n6625,
    n6626, n6627, n6628, n6629, n6630, n6631,
    n6632, n6633, n6634, n6635, n6636, n6637,
    n6638, n6639, n6640, n6641, n6642, n6643,
    n6644, n6645, n6646, n6647, n6648, n6649,
    n6650, n6651, n6652, n6653, n6654, n6655,
    n6656, n6657, n6658, n6659, n6660, n6661,
    n6662, n6663, n6664, n6665, n6666, n6667,
    n6668, n6669, n6670, n6671, n6672, n6673,
    n6674, n6675, n6676, n6677, n6678, n6679,
    n6680, n6681, n6682, n6683, n6684, n6685,
    n6686, n6687, n6688, n6689, n6690, n6691,
    n6692, n6693, n6694, n6695, n6696, n6697,
    n6698, n6699, n6700, n6701, n6702, n6703,
    n6704, n6705, n6706, n6707, n6708, n6709,
    n6710, n6711, n6712, n6713, n6714, n6715,
    n6716, n6717, n6718, n6719, n6720, n6721,
    n6722, n6723, n6724, n6725, n6726, n6727,
    n6728, n6729, n6730, n6731, n6732, n6733,
    n6734, n6735, n6736, n6737, n6738, n6739,
    n6740, n6741, n6742, n6743, n6744, n6745,
    n6746, n6747, n6748, n6749, n6750, n6751,
    n6752, n6753, n6754, n6755, n6756, n6757,
    n6758, n6759, n6760, n6761, n6762, n6763,
    n6764, n6765, n6766, n6767, n6768, n6769,
    n6770, n6771, n6772, n6773, n6774, n6775,
    n6776, n6777, n6778, n6779, n6780, n6781,
    n6782, n6783, n6784, n6785, n6786, n6787,
    n6788, n6789, n6790, n6791, n6792, n6793,
    n6795, n6796, n6797, n6798, n6799, n6800,
    n6801, n6802, n6803, n6804, n6805, n6806,
    n6807, n6808, n6809, n6810, n6811, n6812,
    n6813, n6814, n6815, n6816, n6817, n6818,
    n6819, n6820, n6821, n6822, n6823, n6824,
    n6825, n6826, n6827, n6828, n6829, n6830,
    n6831, n6832, n6833, n6834, n6835, n6836,
    n6837, n6838, n6839, n6840, n6841, n6842,
    n6843, n6844, n6845, n6846, n6847, n6848,
    n6849, n6850, n6851, n6852, n6853, n6854,
    n6855, n6856, n6857, n6858, n6859, n6860,
    n6861, n6862, n6863, n6864, n6865, n6866,
    n6867, n6868, n6869, n6870, n6871, n6872,
    n6873, n6874, n6875, n6876, n6877, n6878,
    n6879, n6880, n6881, n6882, n6883, n6884,
    n6885, n6886, n6887, n6888, n6889, n6890,
    n6891, n6892, n6893, n6894, n6895, n6896,
    n6897, n6898, n6899, n6900, n6901, n6902,
    n6903, n6904, n6905, n6906, n6907, n6908,
    n6909, n6910, n6911, n6912, n6913, n6914,
    n6915, n6916, n6917, n6918, n6919, n6920,
    n6921, n6922, n6923, n6924, n6925, n6926,
    n6927, n6928, n6929, n6930, n6931, n6932,
    n6933, n6934, n6935, n6936, n6937, n6938,
    n6939, n6940, n6941, n6942, n6943, n6944,
    n6945, n6946, n6947, n6948, n6949, n6950,
    n6951, n6952, n6953, n6954, n6955, n6956,
    n6957, n6958, n6959, n6960, n6961, n6962,
    n6963, n6964, n6965, n6966, n6967, n6968,
    n6969, n6970, n6971, n6972, n6973, n6974,
    n6975, n6976, n6977, n6978, n6979, n6980,
    n6981, n6982, n6983, n6984, n6985, n6986,
    n6987, n6988, n6989, n6990, n6991, n6992,
    n6993, n6994, n6995, n6996, n6997, n6998,
    n6999, n7000, n7001, n7002, n7003, n7004,
    n7005, n7006, n7007, n7008, n7009, n7010,
    n7011, n7012, n7013, n7014, n7015, n7016,
    n7017, n7018, n7019, n7020, n7021, n7022,
    n7023, n7024, n7025, n7026, n7027, n7028,
    n7029, n7030, n7031, n7032, n7033, n7034,
    n7035, n7036, n7037, n7038, n7039, n7040,
    n7041, n7042, n7043, n7044, n7045, n7046,
    n7047, n7048, n7049, n7050, n7051, n7052,
    n7053, n7054, n7055, n7056, n7057, n7058,
    n7059, n7060, n7061, n7062, n7063, n7064,
    n7065, n7066, n7067, n7068, n7069, n7070,
    n7071, n7072, n7073, n7074, n7075, n7076,
    n7078, n7079, n7080, n7081, n7082, n7083,
    n7084, n7085, n7086, n7087, n7088, n7089,
    n7090, n7091, n7092, n7093, n7094, n7095,
    n7096, n7097, n7098, n7099, n7100, n7101,
    n7102, n7103, n7104, n7105, n7106, n7107,
    n7108, n7109, n7110, n7111, n7112, n7113,
    n7114, n7115, n7116, n7117, n7118, n7119,
    n7120, n7121, n7122, n7123, n7124, n7125,
    n7126, n7127, n7128, n7129, n7130, n7131,
    n7132, n7133, n7134, n7135, n7136, n7137,
    n7138, n7139, n7140, n7141, n7142, n7143,
    n7144, n7145, n7146, n7147, n7148, n7149,
    n7150, n7151, n7152, n7153, n7154, n7155,
    n7156, n7157, n7158, n7159, n7160, n7161,
    n7162, n7163, n7164, n7165, n7166, n7167,
    n7168, n7169, n7170, n7171, n7172, n7173,
    n7174, n7175, n7176, n7177, n7178, n7179,
    n7180, n7181, n7182, n7183, n7184, n7185,
    n7186, n7187, n7188, n7189, n7190, n7191,
    n7192, n7193, n7194, n7195, n7196, n7197,
    n7198, n7199, n7200, n7201, n7202, n7203,
    n7204, n7205, n7206, n7207, n7208, n7209,
    n7210, n7211, n7212, n7213, n7214, n7215,
    n7216, n7217, n7218, n7219, n7220, n7221,
    n7222, n7223, n7224, n7225, n7226, n7227,
    n7228, n7229, n7230, n7231, n7232, n7233,
    n7234, n7235, n7236, n7237, n7238, n7239,
    n7240, n7241, n7242, n7243, n7244, n7245,
    n7246, n7247, n7248, n7249, n7250, n7251,
    n7252, n7253, n7254, n7255, n7256, n7257,
    n7258, n7259, n7260, n7261, n7262, n7263,
    n7264, n7265, n7266, n7267, n7268, n7269,
    n7270, n7271, n7272, n7273, n7274, n7275,
    n7276, n7277, n7278, n7279, n7280, n7281,
    n7282, n7283, n7284, n7285, n7286, n7287,
    n7288, n7289, n7290, n7291, n7292, n7293,
    n7294, n7295, n7296, n7297, n7298, n7299,
    n7300, n7301, n7302, n7303, n7304, n7305,
    n7306, n7307, n7308, n7309, n7310, n7311,
    n7312, n7313, n7314, n7315, n7316, n7317,
    n7318, n7319, n7320, n7321, n7322, n7323,
    n7324, n7325, n7326, n7327, n7328, n7329,
    n7330, n7331, n7332, n7333, n7334, n7335,
    n7336, n7337, n7338, n7339, n7340, n7341,
    n7342, n7343, n7344, n7345, n7346, n7347,
    n7348, n7349, n7350, n7351, n7352, n7353,
    n7354, n7355, n7356, n7357, n7358, n7359,
    n7360, n7361, n7362, n7363, n7364, n7365,
    n7367, n7368, n7369, n7370, n7371, n7372,
    n7373, n7374, n7375, n7376, n7377, n7378,
    n7379, n7380, n7381, n7382, n7383, n7384,
    n7385, n7386, n7387, n7388, n7389, n7390,
    n7391, n7392, n7393, n7394, n7395, n7396,
    n7397, n7398, n7399, n7400, n7401, n7402,
    n7403, n7404, n7405, n7406, n7407, n7408,
    n7409, n7410, n7411, n7412, n7413, n7414,
    n7415, n7416, n7417, n7418, n7419, n7420,
    n7421, n7422, n7423, n7424, n7425, n7426,
    n7427, n7428, n7429, n7430, n7431, n7432,
    n7433, n7434, n7435, n7436, n7437, n7438,
    n7439, n7440, n7441, n7442, n7443, n7444,
    n7445, n7446, n7447, n7448, n7449, n7450,
    n7451, n7452, n7453, n7454, n7455, n7456,
    n7457, n7458, n7459, n7460, n7461, n7462,
    n7463, n7464, n7465, n7466, n7467, n7468,
    n7469, n7470, n7471, n7472, n7473, n7474,
    n7475, n7476, n7477, n7478, n7479, n7480,
    n7481, n7482, n7483, n7484, n7485, n7486,
    n7487, n7488, n7489, n7490, n7491, n7492,
    n7493, n7494, n7495, n7496, n7497, n7498,
    n7499, n7500, n7501, n7502, n7503, n7504,
    n7505, n7506, n7507, n7508, n7509, n7510,
    n7511, n7512, n7513, n7514, n7515, n7516,
    n7517, n7518, n7519, n7520, n7521, n7522,
    n7523, n7524, n7525, n7526, n7527, n7528,
    n7529, n7530, n7531, n7532, n7533, n7534,
    n7535, n7536, n7537, n7538, n7539, n7540,
    n7541, n7542, n7543, n7544, n7545, n7546,
    n7547, n7548, n7549, n7550, n7551, n7552,
    n7553, n7554, n7555, n7556, n7557, n7558,
    n7559, n7560, n7561, n7562, n7563, n7564,
    n7565, n7566, n7567, n7568, n7569, n7570,
    n7571, n7572, n7573, n7574, n7575, n7576,
    n7577, n7578, n7579, n7580, n7581, n7582,
    n7583, n7584, n7585, n7586, n7587, n7588,
    n7589, n7590, n7591, n7592, n7593, n7594,
    n7595, n7596, n7597, n7598, n7599, n7600,
    n7601, n7602, n7603, n7604, n7605, n7606,
    n7607, n7608, n7609, n7610, n7611, n7612,
    n7613, n7614, n7615, n7616, n7617, n7618,
    n7619, n7620, n7621, n7622, n7623, n7624,
    n7625, n7626, n7627, n7628, n7629, n7630,
    n7631, n7632, n7633, n7634, n7635, n7636,
    n7637, n7638, n7639, n7640, n7641, n7642,
    n7643, n7644, n7645, n7646, n7647, n7648,
    n7649, n7650, n7651, n7652, n7653, n7654,
    n7655, n7656, n7657, n7658, n7659, n7660,
    n7661, n7662, n7663, n7664, n7665, n7666,
    n7667, n7668, n7669, n7670, n7671, n7672,
    n7673, n7674, n7675, n7676, n7677, n7678,
    n7679, n7680, n7681, n7682, n7683, n7685,
    n7686, n7687, n7688, n7689, n7690, n7691,
    n7692, n7693, n7694, n7695, n7696, n7697,
    n7698, n7699, n7700, n7701, n7702, n7703,
    n7704, n7705, n7706, n7707, n7708, n7709,
    n7710, n7711, n7712, n7713, n7714, n7715,
    n7716, n7717, n7718, n7719, n7720, n7721,
    n7722, n7723, n7724, n7725, n7726, n7727,
    n7728, n7729, n7730, n7731, n7732, n7733,
    n7734, n7735, n7736, n7737, n7738, n7739,
    n7740, n7741, n7742, n7743, n7744, n7745,
    n7746, n7747, n7748, n7749, n7750, n7751,
    n7752, n7753, n7754, n7755, n7756, n7757,
    n7758, n7759, n7760, n7761, n7762, n7763,
    n7764, n7765, n7766, n7767, n7768, n7769,
    n7770, n7771, n7772, n7773, n7774, n7775,
    n7776, n7777, n7778, n7779, n7780, n7781,
    n7782, n7783, n7784, n7785, n7786, n7787,
    n7788, n7789, n7790, n7791, n7792, n7793,
    n7794, n7795, n7796, n7797, n7798, n7799,
    n7800, n7801, n7802, n7803, n7804, n7805,
    n7806, n7807, n7808, n7809, n7810, n7811,
    n7812, n7813, n7814, n7815, n7816, n7817,
    n7818, n7819, n7820, n7821, n7822, n7823,
    n7824, n7825, n7826, n7827, n7828, n7829,
    n7830, n7831, n7832, n7833, n7834, n7835,
    n7836, n7837, n7838, n7839, n7840, n7841,
    n7842, n7843, n7844, n7845, n7846, n7847,
    n7848, n7849, n7850, n7851, n7852, n7853,
    n7854, n7855, n7856, n7857, n7858, n7859,
    n7860, n7861, n7862, n7863, n7864, n7865,
    n7866, n7867, n7868, n7869, n7870, n7871,
    n7872, n7873, n7874, n7875, n7876, n7877,
    n7878, n7879, n7880, n7881, n7882, n7883,
    n7884, n7885, n7886, n7887, n7888, n7889,
    n7890, n7891, n7892, n7893, n7894, n7895,
    n7896, n7897, n7898, n7899, n7900, n7901,
    n7902, n7903, n7904, n7905, n7906, n7907,
    n7908, n7909, n7910, n7911, n7912, n7913,
    n7914, n7915, n7916, n7917, n7918, n7919,
    n7920, n7921, n7922, n7923, n7924, n7925,
    n7926, n7927, n7928, n7929, n7930, n7931,
    n7932, n7933, n7934, n7935, n7936, n7937,
    n7938, n7939, n7940, n7941, n7942, n7943,
    n7944, n7945, n7946, n7947, n7948, n7949,
    n7950, n7951, n7952, n7953, n7954, n7955,
    n7956, n7957, n7958, n7959, n7960, n7961,
    n7962, n7963, n7964, n7965, n7966, n7967,
    n7968, n7969, n7970, n7971, n7972, n7973,
    n7974, n7975, n7976, n7977, n7978, n7979,
    n7980, n7981, n7982, n7983, n7984, n7985,
    n7986, n7987, n7988, n7990, n7991, n7992,
    n7993, n7994, n7995, n7996, n7997, n7998,
    n7999, n8000, n8001, n8002, n8003, n8004,
    n8005, n8006, n8007, n8008, n8009, n8010,
    n8011, n8012, n8013, n8014, n8015, n8016,
    n8017, n8018, n8019, n8020, n8021, n8022,
    n8023, n8024, n8025, n8026, n8027, n8028,
    n8029, n8030, n8031, n8032, n8033, n8034,
    n8035, n8036, n8037, n8038, n8039, n8040,
    n8041, n8042, n8043, n8044, n8045, n8046,
    n8047, n8048, n8049, n8050, n8051, n8052,
    n8053, n8054, n8055, n8056, n8057, n8058,
    n8059, n8060, n8061, n8062, n8063, n8064,
    n8065, n8066, n8067, n8068, n8069, n8070,
    n8071, n8072, n8073, n8074, n8075, n8076,
    n8077, n8078, n8079, n8080, n8081, n8082,
    n8083, n8084, n8085, n8086, n8087, n8088,
    n8089, n8090, n8091, n8092, n8093, n8094,
    n8095, n8096, n8097, n8098, n8099, n8100,
    n8101, n8102, n8103, n8104, n8105, n8106,
    n8107, n8108, n8109, n8110, n8111, n8112,
    n8113, n8114, n8115, n8116, n8117, n8118,
    n8119, n8120, n8121, n8122, n8123, n8124,
    n8125, n8126, n8127, n8128, n8129, n8130,
    n8131, n8132, n8133, n8134, n8135, n8136,
    n8137, n8138, n8139, n8140, n8141, n8142,
    n8143, n8144, n8145, n8146, n8147, n8148,
    n8149, n8150, n8151, n8152, n8153, n8154,
    n8155, n8156, n8157, n8158, n8159, n8160,
    n8161, n8162, n8163, n8164, n8165, n8166,
    n8167, n8168, n8169, n8170, n8171, n8172,
    n8173, n8174, n8175, n8176, n8177, n8178,
    n8179, n8180, n8181, n8182, n8183, n8184,
    n8185, n8186, n8187, n8188, n8189, n8190,
    n8191, n8192, n8193, n8194, n8195, n8196,
    n8197, n8198, n8199, n8200, n8201, n8202,
    n8203, n8204, n8205, n8206, n8207, n8208,
    n8209, n8210, n8211, n8212, n8213, n8214,
    n8215, n8216, n8217, n8218, n8219, n8220,
    n8221, n8222, n8223, n8224, n8225, n8226,
    n8227, n8228, n8229, n8230, n8231, n8232,
    n8233, n8234, n8235, n8236, n8237, n8238,
    n8239, n8240, n8241, n8242, n8243, n8244,
    n8245, n8246, n8247, n8248, n8249, n8250,
    n8251, n8252, n8253, n8254, n8255, n8256,
    n8257, n8258, n8259, n8260, n8261, n8262,
    n8263, n8264, n8265, n8266, n8267, n8268,
    n8269, n8270, n8271, n8272, n8273, n8274,
    n8275, n8276, n8277, n8278, n8279, n8280,
    n8281, n8282, n8283, n8284, n8285, n8286,
    n8287, n8288, n8289, n8290, n8291, n8292,
    n8294, n8295, n8296, n8297, n8298, n8299,
    n8300, n8301, n8302, n8303, n8304, n8305,
    n8306, n8307, n8308, n8309, n8310, n8311,
    n8312, n8313, n8314, n8315, n8316, n8317,
    n8318, n8319, n8320, n8321, n8322, n8323,
    n8324, n8325, n8326, n8327, n8328, n8329,
    n8330, n8331, n8332, n8333, n8334, n8335,
    n8336, n8337, n8338, n8339, n8340, n8341,
    n8342, n8343, n8344, n8345, n8346, n8347,
    n8348, n8349, n8350, n8351, n8352, n8353,
    n8354, n8355, n8356, n8357, n8358, n8359,
    n8360, n8361, n8362, n8363, n8364, n8365,
    n8366, n8367, n8368, n8369, n8370, n8371,
    n8372, n8373, n8374, n8375, n8376, n8377,
    n8378, n8379, n8380, n8381, n8382, n8383,
    n8384, n8385, n8386, n8387, n8388, n8389,
    n8390, n8391, n8392, n8393, n8394, n8395,
    n8396, n8397, n8398, n8399, n8400, n8401,
    n8402, n8403, n8404, n8405, n8406, n8407,
    n8408, n8409, n8410, n8411, n8412, n8413,
    n8414, n8415, n8416, n8417, n8418, n8419,
    n8420, n8421, n8422, n8423, n8424, n8425,
    n8426, n8427, n8428, n8429, n8430, n8431,
    n8432, n8433, n8434, n8435, n8436, n8437,
    n8438, n8439, n8440, n8441, n8442, n8443,
    n8444, n8445, n8446, n8447, n8448, n8449,
    n8450, n8451, n8452, n8453, n8454, n8455,
    n8456, n8457, n8458, n8459, n8460, n8461,
    n8462, n8463, n8464, n8465, n8466, n8467,
    n8468, n8469, n8470, n8471, n8472, n8473,
    n8474, n8475, n8476, n8477, n8478, n8479,
    n8480, n8481, n8482, n8483, n8484, n8485,
    n8486, n8487, n8488, n8489, n8490, n8491,
    n8492, n8493, n8494, n8495, n8496, n8497,
    n8498, n8499, n8500, n8501, n8502, n8503,
    n8504, n8505, n8506, n8507, n8508, n8509,
    n8510, n8511, n8512, n8513, n8514, n8515,
    n8516, n8517, n8518, n8519, n8520, n8521,
    n8522, n8523, n8524, n8525, n8526, n8527,
    n8528, n8529, n8530, n8531, n8532, n8533,
    n8534, n8535, n8536, n8537, n8538, n8539,
    n8540, n8541, n8542, n8543, n8544, n8545,
    n8546, n8547, n8548, n8549, n8550, n8551,
    n8552, n8553, n8554, n8555, n8556, n8557,
    n8558, n8559, n8560, n8561, n8562, n8563,
    n8564, n8565, n8566, n8567, n8568, n8569,
    n8570, n8571, n8572, n8573, n8574, n8575,
    n8576, n8577, n8578, n8579, n8580, n8581,
    n8582, n8583, n8584, n8585, n8586, n8587,
    n8588, n8589, n8590, n8591, n8592, n8593,
    n8594, n8595, n8596, n8597, n8598, n8599,
    n8600, n8601, n8602, n8603, n8604, n8605,
    n8606, n8607, n8608, n8609, n8610, n8611,
    n8612, n8613, n8614, n8615, n8616, n8617,
    n8618, n8619, n8620, n8621, n8622, n8623,
    n8624, n8625, n8626, n8627, n8628, n8630,
    n8631, n8632, n8633, n8634, n8635, n8636,
    n8637, n8638, n8639, n8640, n8641, n8642,
    n8643, n8644, n8645, n8646, n8647, n8648,
    n8649, n8650, n8651, n8652, n8653, n8654,
    n8655, n8656, n8657, n8658, n8659, n8660,
    n8661, n8662, n8663, n8664, n8665, n8666,
    n8667, n8668, n8669, n8670, n8671, n8672,
    n8673, n8674, n8675, n8676, n8677, n8678,
    n8679, n8680, n8681, n8682, n8683, n8684,
    n8685, n8686, n8687, n8688, n8689, n8690,
    n8691, n8692, n8693, n8694, n8695, n8696,
    n8697, n8698, n8699, n8700, n8701, n8702,
    n8703, n8704, n8705, n8706, n8707, n8708,
    n8709, n8710, n8711, n8712, n8713, n8714,
    n8715, n8716, n8717, n8718, n8719, n8720,
    n8721, n8722, n8723, n8724, n8725, n8726,
    n8727, n8728, n8729, n8730, n8731, n8732,
    n8733, n8734, n8735, n8736, n8737, n8738,
    n8739, n8740, n8741, n8742, n8743, n8744,
    n8745, n8746, n8747, n8748, n8749, n8750,
    n8751, n8752, n8753, n8754, n8755, n8756,
    n8757, n8758, n8759, n8760, n8761, n8762,
    n8763, n8764, n8765, n8766, n8767, n8768,
    n8769, n8770, n8771, n8772, n8773, n8774,
    n8775, n8776, n8777, n8778, n8779, n8780,
    n8781, n8782, n8783, n8784, n8785, n8786,
    n8787, n8788, n8789, n8790, n8791, n8792,
    n8793, n8794, n8795, n8796, n8797, n8798,
    n8799, n8800, n8801, n8802, n8803, n8804,
    n8805, n8806, n8807, n8808, n8809, n8810,
    n8811, n8812, n8813, n8814, n8815, n8816,
    n8817, n8818, n8819, n8820, n8821, n8822,
    n8823, n8824, n8825, n8826, n8827, n8828,
    n8829, n8830, n8831, n8832, n8833, n8834,
    n8835, n8836, n8837, n8838, n8839, n8840,
    n8841, n8842, n8843, n8844, n8845, n8846,
    n8847, n8848, n8849, n8850, n8851, n8852,
    n8853, n8854, n8855, n8856, n8857, n8858,
    n8859, n8860, n8861, n8862, n8863, n8864,
    n8865, n8866, n8867, n8868, n8869, n8870,
    n8871, n8872, n8873, n8874, n8875, n8876,
    n8877, n8878, n8879, n8880, n8881, n8882,
    n8883, n8884, n8885, n8886, n8887, n8888,
    n8889, n8890, n8891, n8892, n8893, n8894,
    n8895, n8896, n8897, n8898, n8899, n8900,
    n8901, n8902, n8903, n8904, n8905, n8906,
    n8907, n8908, n8909, n8910, n8911, n8912,
    n8913, n8914, n8915, n8916, n8917, n8918,
    n8919, n8920, n8921, n8922, n8923, n8924,
    n8925, n8926, n8927, n8928, n8929, n8930,
    n8931, n8932, n8933, n8934, n8935, n8936,
    n8937, n8938, n8939, n8940, n8941, n8942,
    n8943, n8944, n8945, n8946, n8947, n8948,
    n8949, n8950, n8951, n8952, n8953, n8954,
    n8956, n8957, n8958, n8959, n8960, n8961,
    n8962, n8963, n8964, n8965, n8966, n8967,
    n8968, n8969, n8970, n8971, n8972, n8973,
    n8974, n8975, n8976, n8977, n8978, n8979,
    n8980, n8981, n8982, n8983, n8984, n8985,
    n8986, n8987, n8988, n8989, n8990, n8991,
    n8992, n8993, n8994, n8995, n8996, n8997,
    n8998, n8999, n9000, n9001, n9002, n9003,
    n9004, n9005, n9006, n9007, n9008, n9009,
    n9010, n9011, n9012, n9013, n9014, n9015,
    n9016, n9017, n9018, n9019, n9020, n9021,
    n9022, n9023, n9024, n9025, n9026, n9027,
    n9028, n9029, n9030, n9031, n9032, n9033,
    n9034, n9035, n9036, n9037, n9038, n9039,
    n9040, n9041, n9042, n9043, n9044, n9045,
    n9046, n9047, n9048, n9049, n9050, n9051,
    n9052, n9053, n9054, n9055, n9056, n9057,
    n9058, n9059, n9060, n9061, n9062, n9063,
    n9064, n9065, n9066, n9067, n9068, n9069,
    n9070, n9071, n9072, n9073, n9074, n9075,
    n9076, n9077, n9078, n9079, n9080, n9081,
    n9082, n9083, n9084, n9085, n9086, n9087,
    n9088, n9089, n9090, n9091, n9092, n9093,
    n9094, n9095, n9096, n9097, n9098, n9099,
    n9100, n9101, n9102, n9103, n9104, n9105,
    n9106, n9107, n9108, n9109, n9110, n9111,
    n9112, n9113, n9114, n9115, n9116, n9117,
    n9118, n9119, n9120, n9121, n9122, n9123,
    n9124, n9125, n9126, n9127, n9128, n9129,
    n9130, n9131, n9132, n9133, n9134, n9135,
    n9136, n9137, n9138, n9139, n9140, n9141,
    n9142, n9143, n9144, n9145, n9146, n9147,
    n9148, n9149, n9150, n9151, n9152, n9153,
    n9154, n9155, n9156, n9157, n9158, n9159,
    n9160, n9161, n9162, n9163, n9164, n9165,
    n9166, n9167, n9168, n9169, n9170, n9171,
    n9172, n9173, n9174, n9175, n9176, n9177,
    n9178, n9179, n9180, n9181, n9182, n9183,
    n9184, n9185, n9186, n9187, n9188, n9189,
    n9190, n9191, n9192, n9193, n9194, n9195,
    n9196, n9197, n9198, n9199, n9200, n9201,
    n9202, n9203, n9204, n9205, n9206, n9207,
    n9208, n9209, n9210, n9211, n9212, n9213,
    n9214, n9215, n9216, n9217, n9218, n9219,
    n9220, n9221, n9222, n9223, n9224, n9225,
    n9226, n9227, n9228, n9229, n9230, n9231,
    n9232, n9233, n9234, n9235, n9236, n9237,
    n9238, n9239, n9240, n9241, n9242, n9243,
    n9244, n9245, n9246, n9247, n9248, n9249,
    n9250, n9251, n9252, n9253, n9254, n9255,
    n9256, n9257, n9258, n9259, n9260, n9261,
    n9262, n9263, n9264, n9265, n9266, n9267,
    n9268, n9269, n9270, n9271, n9272, n9273,
    n9274, n9275, n9277, n9278, n9279, n9280,
    n9281, n9282, n9283, n9284, n9285, n9286,
    n9287, n9288, n9289, n9290, n9291, n9292,
    n9293, n9294, n9295, n9296, n9297, n9298,
    n9299, n9300, n9301, n9302, n9303, n9304,
    n9305, n9306, n9307, n9308, n9309, n9310,
    n9311, n9312, n9313, n9314, n9315, n9316,
    n9317, n9318, n9319, n9320, n9321, n9322,
    n9323, n9324, n9325, n9326, n9327, n9328,
    n9329, n9330, n9331, n9332, n9333, n9334,
    n9335, n9336, n9337, n9338, n9339, n9340,
    n9341, n9342, n9343, n9344, n9345, n9346,
    n9347, n9348, n9349, n9350, n9351, n9352,
    n9353, n9354, n9355, n9356, n9357, n9358,
    n9359, n9360, n9361, n9362, n9363, n9364,
    n9365, n9366, n9367, n9368, n9369, n9370,
    n9371, n9372, n9373, n9374, n9375, n9376,
    n9377, n9378, n9379, n9380, n9381, n9382,
    n9383, n9384, n9385, n9386, n9387, n9388,
    n9389, n9390, n9391, n9392, n9393, n9394,
    n9395, n9396, n9397, n9398, n9399, n9400,
    n9401, n9402, n9403, n9404, n9405, n9406,
    n9407, n9408, n9409, n9410, n9411, n9412,
    n9413, n9414, n9415, n9416, n9417, n9418,
    n9419, n9420, n9421, n9422, n9423, n9424,
    n9425, n9426, n9427, n9428, n9429, n9430,
    n9431, n9432, n9433, n9434, n9435, n9436,
    n9437, n9438, n9439, n9440, n9441, n9442,
    n9443, n9444, n9445, n9446, n9447, n9448,
    n9449, n9450, n9451, n9452, n9453, n9454,
    n9455, n9456, n9457, n9458, n9459, n9460,
    n9461, n9462, n9463, n9464, n9465, n9466,
    n9467, n9468, n9469, n9470, n9471, n9472,
    n9473, n9474, n9475, n9476, n9477, n9478,
    n9479, n9480, n9481, n9482, n9483, n9484,
    n9485, n9486, n9487, n9488, n9489, n9490,
    n9491, n9492, n9493, n9494, n9495, n9496,
    n9497, n9498, n9499, n9500, n9501, n9502,
    n9503, n9504, n9505, n9506, n9507, n9508,
    n9509, n9510, n9511, n9512, n9513, n9514,
    n9515, n9516, n9517, n9518, n9519, n9520,
    n9521, n9522, n9523, n9524, n9525, n9526,
    n9527, n9528, n9529, n9530, n9531, n9532,
    n9533, n9534, n9535, n9536, n9537, n9538,
    n9539, n9540, n9541, n9542, n9543, n9544,
    n9545, n9546, n9547, n9548, n9549, n9550,
    n9551, n9552, n9553, n9554, n9555, n9556,
    n9557, n9558, n9559, n9560, n9561, n9562,
    n9563, n9564, n9565, n9566, n9567, n9568,
    n9569, n9570, n9571, n9572, n9573, n9574,
    n9575, n9576, n9577, n9578, n9579, n9580,
    n9581, n9582, n9583, n9584, n9585, n9586,
    n9587, n9588, n9589, n9590, n9591, n9592,
    n9593, n9594, n9595, n9596, n9597, n9598,
    n9599, n9600, n9601, n9602, n9603, n9604,
    n9605, n9606, n9607, n9608, n9609, n9610,
    n9611, n9612, n9613, n9614, n9615, n9616,
    n9617, n9618, n9619, n9620, n9621, n9622,
    n9623, n9624, n9625, n9626, n9627, n9628,
    n9629, n9630, n9632, n9633, n9634, n9635,
    n9636, n9637, n9638, n9639, n9640, n9641,
    n9642, n9643, n9644, n9645, n9646, n9647,
    n9648, n9649, n9650, n9651, n9652, n9653,
    n9654, n9655, n9656, n9657, n9658, n9659,
    n9660, n9661, n9662, n9663, n9664, n9665,
    n9666, n9667, n9668, n9669, n9670, n9671,
    n9672, n9673, n9674, n9675, n9676, n9677,
    n9678, n9679, n9680, n9681, n9682, n9683,
    n9684, n9685, n9686, n9687, n9688, n9689,
    n9690, n9691, n9692, n9693, n9694, n9695,
    n9696, n9697, n9698, n9699, n9700, n9701,
    n9702, n9703, n9704, n9705, n9706, n9707,
    n9708, n9709, n9710, n9711, n9712, n9713,
    n9714, n9715, n9716, n9717, n9718, n9719,
    n9720, n9721, n9722, n9723, n9724, n9725,
    n9726, n9727, n9728, n9729, n9730, n9731,
    n9732, n9733, n9734, n9735, n9736, n9737,
    n9738, n9739, n9740, n9741, n9742, n9743,
    n9744, n9745, n9746, n9747, n9748, n9749,
    n9750, n9751, n9752, n9753, n9754, n9755,
    n9756, n9757, n9758, n9759, n9760, n9761,
    n9762, n9763, n9764, n9765, n9766, n9767,
    n9768, n9769, n9770, n9771, n9772, n9773,
    n9774, n9775, n9776, n9777, n9778, n9779,
    n9780, n9781, n9782, n9783, n9784, n9785,
    n9786, n9787, n9788, n9789, n9790, n9791,
    n9792, n9793, n9794, n9795, n9796, n9797,
    n9798, n9799, n9800, n9801, n9802, n9803,
    n9804, n9805, n9806, n9807, n9808, n9809,
    n9810, n9811, n9812, n9813, n9814, n9815,
    n9816, n9817, n9818, n9819, n9820, n9821,
    n9822, n9823, n9824, n9825, n9826, n9827,
    n9828, n9829, n9830, n9831, n9832, n9833,
    n9834, n9835, n9836, n9837, n9838, n9839,
    n9840, n9841, n9842, n9843, n9844, n9845,
    n9846, n9847, n9848, n9849, n9850, n9851,
    n9852, n9853, n9854, n9855, n9856, n9857,
    n9858, n9859, n9860, n9861, n9862, n9863,
    n9864, n9865, n9866, n9867, n9868, n9869,
    n9870, n9871, n9872, n9873, n9874, n9875,
    n9876, n9877, n9878, n9879, n9880, n9881,
    n9882, n9883, n9884, n9885, n9886, n9887,
    n9888, n9889, n9890, n9891, n9892, n9893,
    n9894, n9895, n9896, n9897, n9898, n9899,
    n9900, n9901, n9902, n9903, n9904, n9905,
    n9906, n9907, n9908, n9909, n9910, n9911,
    n9912, n9913, n9914, n9915, n9916, n9917,
    n9918, n9919, n9920, n9921, n9922, n9923,
    n9924, n9925, n9926, n9927, n9928, n9929,
    n9930, n9931, n9932, n9933, n9934, n9935,
    n9936, n9937, n9938, n9939, n9940, n9941,
    n9942, n9943, n9944, n9945, n9946, n9947,
    n9948, n9949, n9950, n9951, n9952, n9953,
    n9954, n9955, n9956, n9957, n9958, n9959,
    n9960, n9961, n9962, n9963, n9964, n9965,
    n9966, n9967, n9968, n9969, n9970, n9971,
    n9972, n9973, n9974, n9976, n9977, n9978,
    n9979, n9980, n9981, n9982, n9983, n9984,
    n9985, n9986, n9987, n9988, n9989, n9990,
    n9991, n9992, n9993, n9994, n9995, n9996,
    n9997, n9998, n9999, n10000, n10001, n10002,
    n10003, n10004, n10005, n10006, n10007, n10008,
    n10009, n10010, n10011, n10012, n10013, n10014,
    n10015, n10016, n10017, n10018, n10019, n10020,
    n10021, n10022, n10023, n10024, n10025, n10026,
    n10027, n10028, n10029, n10030, n10031, n10032,
    n10033, n10034, n10035, n10036, n10037, n10038,
    n10039, n10040, n10041, n10042, n10043, n10044,
    n10045, n10046, n10047, n10048, n10049, n10050,
    n10051, n10052, n10053, n10054, n10055, n10056,
    n10057, n10058, n10059, n10060, n10061, n10062,
    n10063, n10064, n10065, n10066, n10067, n10068,
    n10069, n10070, n10071, n10072, n10073, n10074,
    n10075, n10076, n10077, n10078, n10079, n10080,
    n10081, n10082, n10083, n10084, n10085, n10086,
    n10087, n10088, n10089, n10090, n10091, n10092,
    n10093, n10094, n10095, n10096, n10097, n10098,
    n10099, n10100, n10101, n10102, n10103, n10104,
    n10105, n10106, n10107, n10108, n10109, n10110,
    n10111, n10112, n10113, n10114, n10115, n10116,
    n10117, n10118, n10119, n10120, n10121, n10122,
    n10123, n10124, n10125, n10126, n10127, n10128,
    n10129, n10130, n10131, n10132, n10133, n10134,
    n10135, n10136, n10137, n10138, n10139, n10140,
    n10141, n10142, n10143, n10144, n10145, n10146,
    n10147, n10148, n10149, n10150, n10151, n10152,
    n10153, n10154, n10155, n10156, n10157, n10158,
    n10159, n10160, n10161, n10162, n10163, n10164,
    n10165, n10166, n10167, n10168, n10169, n10170,
    n10171, n10172, n10173, n10174, n10175, n10176,
    n10177, n10178, n10179, n10180, n10181, n10182,
    n10183, n10184, n10185, n10186, n10187, n10188,
    n10189, n10190, n10191, n10192, n10193, n10194,
    n10195, n10196, n10197, n10198, n10199, n10200,
    n10201, n10202, n10203, n10204, n10205, n10206,
    n10207, n10208, n10209, n10210, n10211, n10212,
    n10213, n10214, n10215, n10216, n10217, n10218,
    n10219, n10220, n10221, n10222, n10223, n10224,
    n10225, n10226, n10227, n10228, n10229, n10230,
    n10231, n10232, n10233, n10234, n10235, n10236,
    n10237, n10238, n10239, n10240, n10241, n10242,
    n10243, n10244, n10245, n10246, n10247, n10248,
    n10249, n10250, n10251, n10252, n10253, n10254,
    n10255, n10256, n10257, n10258, n10259, n10260,
    n10261, n10262, n10263, n10264, n10265, n10266,
    n10267, n10268, n10269, n10270, n10271, n10272,
    n10273, n10274, n10275, n10276, n10277, n10278,
    n10279, n10280, n10281, n10282, n10283, n10284,
    n10285, n10286, n10287, n10288, n10289, n10290,
    n10291, n10292, n10293, n10294, n10295, n10296,
    n10297, n10298, n10299, n10300, n10301, n10302,
    n10303, n10304, n10305, n10306, n10307, n10308,
    n10309, n10310, n10311, n10312, n10313, n10314,
    n10315, n10317, n10318, n10319, n10320, n10321,
    n10322, n10323, n10324, n10325, n10326, n10327,
    n10328, n10329, n10330, n10331, n10332, n10333,
    n10334, n10335, n10336, n10337, n10338, n10339,
    n10340, n10341, n10342, n10343, n10344, n10345,
    n10346, n10347, n10348, n10349, n10350, n10351,
    n10352, n10353, n10354, n10355, n10356, n10357,
    n10358, n10359, n10360, n10361, n10362, n10363,
    n10364, n10365, n10366, n10367, n10368, n10369,
    n10370, n10371, n10372, n10373, n10374, n10375,
    n10376, n10377, n10378, n10379, n10380, n10381,
    n10382, n10383, n10384, n10385, n10386, n10387,
    n10388, n10389, n10390, n10391, n10392, n10393,
    n10394, n10395, n10396, n10397, n10398, n10399,
    n10400, n10401, n10402, n10403, n10404, n10405,
    n10406, n10407, n10408, n10409, n10410, n10411,
    n10412, n10413, n10414, n10415, n10416, n10417,
    n10418, n10419, n10420, n10421, n10422, n10423,
    n10424, n10425, n10426, n10427, n10428, n10429,
    n10430, n10431, n10432, n10433, n10434, n10435,
    n10436, n10437, n10438, n10439, n10440, n10441,
    n10442, n10443, n10444, n10445, n10446, n10447,
    n10448, n10449, n10450, n10451, n10452, n10453,
    n10454, n10455, n10456, n10457, n10458, n10459,
    n10460, n10461, n10462, n10463, n10464, n10465,
    n10466, n10467, n10468, n10469, n10470, n10471,
    n10472, n10473, n10474, n10475, n10476, n10477,
    n10478, n10479, n10480, n10481, n10482, n10483,
    n10484, n10485, n10486, n10487, n10488, n10489,
    n10490, n10491, n10492, n10493, n10494, n10495,
    n10496, n10497, n10498, n10499, n10500, n10501,
    n10502, n10503, n10504, n10505, n10506, n10507,
    n10508, n10509, n10510, n10511, n10512, n10513,
    n10514, n10515, n10516, n10517, n10518, n10519,
    n10520, n10521, n10522, n10523, n10524, n10525,
    n10526, n10527, n10528, n10529, n10530, n10531,
    n10532, n10533, n10534, n10535, n10536, n10537,
    n10538, n10539, n10540, n10541, n10542, n10543,
    n10544, n10545, n10546, n10547, n10548, n10549,
    n10550, n10551, n10552, n10553, n10554, n10555,
    n10556, n10557, n10558, n10559, n10560, n10561,
    n10562, n10563, n10564, n10565, n10566, n10567,
    n10568, n10569, n10570, n10571, n10572, n10573,
    n10574, n10575, n10576, n10577, n10578, n10579,
    n10580, n10581, n10582, n10583, n10584, n10585,
    n10586, n10587, n10588, n10589, n10590, n10591,
    n10592, n10593, n10594, n10595, n10596, n10597,
    n10598, n10599, n10600, n10601, n10602, n10603,
    n10604, n10605, n10606, n10607, n10608, n10609,
    n10610, n10611, n10612, n10613, n10614, n10615,
    n10616, n10617, n10618, n10619, n10620, n10621,
    n10622, n10623, n10624, n10625, n10626, n10627,
    n10628, n10629, n10630, n10631, n10632, n10633,
    n10634, n10635, n10636, n10637, n10638, n10639,
    n10640, n10641, n10642, n10643, n10644, n10645,
    n10646, n10647, n10648, n10649, n10650, n10651,
    n10652, n10653, n10654, n10655, n10656, n10657,
    n10658, n10659, n10660, n10661, n10662, n10663,
    n10664, n10665, n10666, n10667, n10668, n10669,
    n10670, n10671, n10672, n10673, n10674, n10675,
    n10676, n10677, n10678, n10679, n10680, n10681,
    n10682, n10683, n10685, n10686, n10687, n10688,
    n10689, n10690, n10691, n10692, n10693, n10694,
    n10695, n10696, n10697, n10698, n10699, n10700,
    n10701, n10702, n10703, n10704, n10705, n10706,
    n10707, n10708, n10709, n10710, n10711, n10712,
    n10713, n10714, n10715, n10716, n10717, n10718,
    n10719, n10720, n10721, n10722, n10723, n10724,
    n10725, n10726, n10727, n10728, n10729, n10730,
    n10731, n10732, n10733, n10734, n10735, n10736,
    n10737, n10738, n10739, n10740, n10741, n10742,
    n10743, n10744, n10745, n10746, n10747, n10748,
    n10749, n10750, n10751, n10752, n10753, n10754,
    n10755, n10756, n10757, n10758, n10759, n10760,
    n10761, n10762, n10763, n10764, n10765, n10766,
    n10767, n10768, n10769, n10770, n10771, n10772,
    n10773, n10774, n10775, n10776, n10777, n10778,
    n10779, n10780, n10781, n10782, n10783, n10784,
    n10785, n10786, n10787, n10788, n10789, n10790,
    n10791, n10792, n10793, n10794, n10795, n10796,
    n10797, n10798, n10799, n10800, n10801, n10802,
    n10803, n10804, n10805, n10806, n10807, n10808,
    n10809, n10810, n10811, n10812, n10813, n10814,
    n10815, n10816, n10817, n10818, n10819, n10820,
    n10821, n10822, n10823, n10824, n10825, n10826,
    n10827, n10828, n10829, n10830, n10831, n10832,
    n10833, n10834, n10835, n10836, n10837, n10838,
    n10839, n10840, n10841, n10842, n10843, n10844,
    n10845, n10846, n10847, n10848, n10849, n10850,
    n10851, n10852, n10853, n10854, n10855, n10856,
    n10857, n10858, n10859, n10860, n10861, n10862,
    n10863, n10864, n10865, n10866, n10867, n10868,
    n10869, n10870, n10871, n10872, n10873, n10874,
    n10875, n10876, n10877, n10878, n10879, n10880,
    n10881, n10882, n10883, n10884, n10885, n10886,
    n10887, n10888, n10889, n10890, n10891, n10892,
    n10893, n10894, n10895, n10896, n10897, n10898,
    n10899, n10900, n10901, n10902, n10903, n10904,
    n10905, n10906, n10907, n10908, n10909, n10910,
    n10911, n10912, n10913, n10914, n10915, n10916,
    n10917, n10918, n10919, n10920, n10921, n10922,
    n10923, n10924, n10925, n10926, n10927, n10928,
    n10929, n10930, n10931, n10932, n10933, n10934,
    n10935, n10936, n10937, n10938, n10939, n10940,
    n10941, n10942, n10943, n10944, n10945, n10946,
    n10947, n10948, n10949, n10950, n10951, n10952,
    n10953, n10954, n10955, n10956, n10957, n10958,
    n10959, n10960, n10961, n10962, n10963, n10964,
    n10965, n10966, n10967, n10968, n10969, n10970,
    n10971, n10972, n10973, n10974, n10975, n10976,
    n10977, n10978, n10979, n10980, n10981, n10982,
    n10983, n10984, n10985, n10986, n10987, n10988,
    n10989, n10990, n10991, n10992, n10993, n10994,
    n10995, n10996, n10997, n10998, n10999, n11000,
    n11001, n11002, n11003, n11004, n11005, n11006,
    n11007, n11008, n11009, n11010, n11011, n11012,
    n11013, n11014, n11015, n11016, n11017, n11018,
    n11019, n11020, n11021, n11022, n11023, n11024,
    n11025, n11026, n11027, n11028, n11029, n11030,
    n11031, n11032, n11033, n11034, n11035, n11036,
    n11037, n11038, n11039, n11040, n11041, n11042,
    n11043, n11044, n11045, n11046, n11048, n11049,
    n11050, n11051, n11052, n11053, n11054, n11055,
    n11056, n11057, n11058, n11059, n11060, n11061,
    n11062, n11063, n11064, n11065, n11066, n11067,
    n11068, n11069, n11070, n11071, n11072, n11073,
    n11074, n11075, n11076, n11077, n11078, n11079,
    n11080, n11081, n11082, n11083, n11084, n11085,
    n11086, n11087, n11088, n11089, n11090, n11091,
    n11092, n11093, n11094, n11095, n11096, n11097,
    n11098, n11099, n11100, n11101, n11102, n11103,
    n11104, n11105, n11106, n11107, n11108, n11109,
    n11110, n11111, n11112, n11113, n11114, n11115,
    n11116, n11117, n11118, n11119, n11120, n11121,
    n11122, n11123, n11124, n11125, n11126, n11127,
    n11128, n11129, n11130, n11131, n11132, n11133,
    n11134, n11135, n11136, n11137, n11138, n11139,
    n11140, n11141, n11142, n11143, n11144, n11145,
    n11146, n11147, n11148, n11149, n11150, n11151,
    n11152, n11153, n11154, n11155, n11156, n11157,
    n11158, n11159, n11160, n11161, n11162, n11163,
    n11164, n11165, n11166, n11167, n11168, n11169,
    n11170, n11171, n11172, n11173, n11174, n11175,
    n11176, n11177, n11178, n11179, n11180, n11181,
    n11182, n11183, n11184, n11185, n11186, n11187,
    n11188, n11189, n11190, n11191, n11192, n11193,
    n11194, n11195, n11196, n11197, n11198, n11199,
    n11200, n11201, n11202, n11203, n11204, n11205,
    n11206, n11207, n11208, n11209, n11210, n11211,
    n11212, n11213, n11214, n11215, n11216, n11217,
    n11218, n11219, n11220, n11221, n11222, n11223,
    n11224, n11225, n11226, n11227, n11228, n11229,
    n11230, n11231, n11232, n11233, n11234, n11235,
    n11236, n11237, n11238, n11239, n11240, n11241,
    n11242, n11243, n11244, n11245, n11246, n11247,
    n11248, n11249, n11250, n11251, n11252, n11253,
    n11254, n11255, n11256, n11257, n11258, n11259,
    n11260, n11261, n11262, n11263, n11264, n11265,
    n11266, n11267, n11268, n11269, n11270, n11271,
    n11272, n11273, n11274, n11275, n11276, n11277,
    n11278, n11279, n11280, n11281, n11282, n11283,
    n11284, n11285, n11286, n11287, n11288, n11289,
    n11290, n11291, n11292, n11293, n11294, n11295,
    n11296, n11297, n11298, n11299, n11300, n11301,
    n11302, n11303, n11304, n11305, n11306, n11307,
    n11308, n11309, n11310, n11311, n11312, n11313,
    n11314, n11315, n11316, n11317, n11318, n11319,
    n11320, n11321, n11322, n11323, n11324, n11325,
    n11326, n11327, n11328, n11329, n11330, n11331,
    n11332, n11333, n11334, n11335, n11336, n11337,
    n11338, n11339, n11340, n11341, n11342, n11343,
    n11344, n11345, n11346, n11347, n11348, n11349,
    n11350, n11351, n11352, n11353, n11354, n11355,
    n11356, n11357, n11358, n11359, n11360, n11361,
    n11362, n11363, n11364, n11365, n11366, n11367,
    n11368, n11369, n11370, n11371, n11372, n11373,
    n11374, n11375, n11376, n11377, n11378, n11379,
    n11380, n11381, n11382, n11383, n11384, n11385,
    n11386, n11387, n11388, n11389, n11390, n11391,
    n11392, n11393, n11394, n11395, n11396, n11397,
    n11398, n11399, n11400, n11401, n11402, n11403,
    n11404, n11405, n11406, n11407, n11409, n11410,
    n11411, n11412, n11413, n11414, n11415, n11416,
    n11417, n11418, n11419, n11420, n11421, n11422,
    n11423, n11424, n11425, n11426, n11427, n11428,
    n11429, n11430, n11431, n11432, n11433, n11434,
    n11435, n11436, n11437, n11438, n11439, n11440,
    n11441, n11442, n11443, n11444, n11445, n11446,
    n11447, n11448, n11449, n11450, n11451, n11452,
    n11453, n11454, n11455, n11456, n11457, n11458,
    n11459, n11460, n11461, n11462, n11463, n11464,
    n11465, n11466, n11467, n11468, n11469, n11470,
    n11471, n11472, n11473, n11474, n11475, n11476,
    n11477, n11478, n11479, n11480, n11481, n11482,
    n11483, n11484, n11485, n11486, n11487, n11488,
    n11489, n11490, n11491, n11492, n11493, n11494,
    n11495, n11496, n11497, n11498, n11499, n11500,
    n11501, n11502, n11503, n11504, n11505, n11506,
    n11507, n11508, n11509, n11510, n11511, n11512,
    n11513, n11514, n11515, n11516, n11517, n11518,
    n11519, n11520, n11521, n11522, n11523, n11524,
    n11525, n11526, n11527, n11528, n11529, n11530,
    n11531, n11532, n11533, n11534, n11535, n11536,
    n11537, n11538, n11539, n11540, n11541, n11542,
    n11543, n11544, n11545, n11546, n11547, n11548,
    n11549, n11550, n11551, n11552, n11553, n11554,
    n11555, n11556, n11557, n11558, n11559, n11560,
    n11561, n11562, n11563, n11564, n11565, n11566,
    n11567, n11568, n11569, n11570, n11571, n11572,
    n11573, n11574, n11575, n11576, n11577, n11578,
    n11579, n11580, n11581, n11582, n11583, n11584,
    n11585, n11586, n11587, n11588, n11589, n11590,
    n11591, n11592, n11593, n11594, n11595, n11596,
    n11597, n11598, n11599, n11600, n11601, n11602,
    n11603, n11604, n11605, n11606, n11607, n11608,
    n11609, n11610, n11611, n11612, n11613, n11614,
    n11615, n11616, n11617, n11618, n11619, n11620,
    n11621, n11622, n11623, n11624, n11625, n11626,
    n11627, n11628, n11629, n11630, n11631, n11632,
    n11633, n11634, n11635, n11636, n11637, n11638,
    n11639, n11640, n11641, n11642, n11643, n11644,
    n11645, n11646, n11647, n11648, n11649, n11650,
    n11651, n11652, n11653, n11654, n11655, n11656,
    n11657, n11658, n11659, n11660, n11661, n11662,
    n11663, n11664, n11665, n11666, n11667, n11668,
    n11669, n11670, n11671, n11672, n11673, n11674,
    n11675, n11676, n11677, n11678, n11679, n11680,
    n11681, n11682, n11683, n11684, n11685, n11686,
    n11687, n11688, n11689, n11690, n11691, n11692,
    n11693, n11694, n11695, n11696, n11697, n11698,
    n11699, n11700, n11701, n11702, n11703, n11704,
    n11705, n11706, n11707, n11708, n11709, n11710,
    n11711, n11712, n11713, n11714, n11715, n11716,
    n11717, n11718, n11719, n11720, n11721, n11722,
    n11723, n11724, n11725, n11726, n11727, n11728,
    n11729, n11730, n11731, n11732, n11733, n11734,
    n11735, n11736, n11737, n11738, n11739, n11740,
    n11741, n11742, n11743, n11744, n11745, n11746,
    n11747, n11748, n11749, n11750, n11751, n11752,
    n11753, n11754, n11755, n11756, n11757, n11758,
    n11759, n11760, n11761, n11762, n11763, n11764,
    n11765, n11766, n11767, n11768, n11769, n11770,
    n11771, n11772, n11773, n11774, n11775, n11776,
    n11777, n11778, n11779, n11780, n11781, n11782,
    n11783, n11784, n11785, n11786, n11787, n11788,
    n11789, n11790, n11791, n11792, n11793, n11794,
    n11795, n11796, n11798, n11799, n11800, n11801,
    n11802, n11803, n11804, n11805, n11806, n11807,
    n11808, n11809, n11810, n11811, n11812, n11813,
    n11814, n11815, n11816, n11817, n11818, n11819,
    n11820, n11821, n11822, n11823, n11824, n11825,
    n11826, n11827, n11828, n11829, n11830, n11831,
    n11832, n11833, n11834, n11835, n11836, n11837,
    n11838, n11839, n11840, n11841, n11842, n11843,
    n11844, n11845, n11846, n11847, n11848, n11849,
    n11850, n11851, n11852, n11853, n11854, n11855,
    n11856, n11857, n11858, n11859, n11860, n11861,
    n11862, n11863, n11864, n11865, n11866, n11867,
    n11868, n11869, n11870, n11871, n11872, n11873,
    n11874, n11875, n11876, n11877, n11878, n11879,
    n11880, n11881, n11882, n11883, n11884, n11885,
    n11886, n11887, n11888, n11889, n11890, n11891,
    n11892, n11893, n11894, n11895, n11896, n11897,
    n11898, n11899, n11900, n11901, n11902, n11903,
    n11904, n11905, n11906, n11907, n11908, n11909,
    n11910, n11911, n11912, n11913, n11914, n11915,
    n11916, n11917, n11918, n11919, n11920, n11921,
    n11922, n11923, n11924, n11925, n11926, n11927,
    n11928, n11929, n11930, n11931, n11932, n11933,
    n11934, n11935, n11936, n11937, n11938, n11939,
    n11940, n11941, n11942, n11943, n11944, n11945,
    n11946, n11947, n11948, n11949, n11950, n11951,
    n11952, n11953, n11954, n11955, n11956, n11957,
    n11958, n11959, n11960, n11961, n11962, n11963,
    n11964, n11965, n11966, n11967, n11968, n11969,
    n11970, n11971, n11972, n11973, n11974, n11975,
    n11976, n11977, n11978, n11979, n11980, n11981,
    n11982, n11983, n11984, n11985, n11986, n11987,
    n11988, n11989, n11990, n11991, n11992, n11993,
    n11994, n11995, n11996, n11997, n11998, n11999,
    n12000, n12001, n12002, n12003, n12004, n12005,
    n12006, n12007, n12008, n12009, n12010, n12011,
    n12012, n12013, n12014, n12015, n12016, n12017,
    n12018, n12019, n12020, n12021, n12022, n12023,
    n12024, n12025, n12026, n12027, n12028, n12029,
    n12030, n12031, n12032, n12033, n12034, n12035,
    n12036, n12037, n12038, n12039, n12040, n12041,
    n12042, n12043, n12044, n12045, n12046, n12047,
    n12048, n12049, n12050, n12051, n12052, n12053,
    n12054, n12055, n12056, n12057, n12058, n12059,
    n12060, n12061, n12062, n12063, n12064, n12065,
    n12066, n12067, n12068, n12069, n12070, n12071,
    n12072, n12073, n12074, n12075, n12076, n12077,
    n12078, n12079, n12080, n12081, n12082, n12083,
    n12084, n12085, n12086, n12087, n12088, n12089,
    n12090, n12091, n12092, n12093, n12094, n12095,
    n12096, n12097, n12098, n12099, n12100, n12101,
    n12102, n12103, n12104, n12105, n12106, n12107,
    n12108, n12109, n12110, n12111, n12112, n12113,
    n12114, n12115, n12116, n12117, n12118, n12119,
    n12120, n12121, n12122, n12123, n12124, n12125,
    n12126, n12127, n12128, n12129, n12130, n12131,
    n12132, n12133, n12134, n12135, n12136, n12137,
    n12138, n12139, n12140, n12141, n12142, n12143,
    n12144, n12145, n12146, n12147, n12148, n12149,
    n12150, n12151, n12152, n12153, n12154, n12155,
    n12156, n12157, n12158, n12159, n12160, n12161,
    n12162, n12163, n12164, n12165, n12166, n12167,
    n12168, n12169, n12170, n12171, n12172, n12173,
    n12174, n12175, n12176, n12177, n12178, n12180,
    n12181, n12182, n12183, n12184, n12185, n12186,
    n12187, n12188, n12189, n12190, n12191, n12192,
    n12193, n12194, n12195, n12196, n12197, n12198,
    n12199, n12200, n12201, n12202, n12203, n12204,
    n12205, n12206, n12207, n12208, n12209, n12210,
    n12211, n12212, n12213, n12214, n12215, n12216,
    n12217, n12218, n12219, n12220, n12221, n12222,
    n12223, n12224, n12225, n12226, n12227, n12228,
    n12229, n12230, n12231, n12232, n12233, n12234,
    n12235, n12236, n12237, n12238, n12239, n12240,
    n12241, n12242, n12243, n12244, n12245, n12246,
    n12247, n12248, n12249, n12250, n12251, n12252,
    n12253, n12254, n12255, n12256, n12257, n12258,
    n12259, n12260, n12261, n12262, n12263, n12264,
    n12265, n12266, n12267, n12268, n12269, n12270,
    n12271, n12272, n12273, n12274, n12275, n12276,
    n12277, n12278, n12279, n12280, n12281, n12282,
    n12283, n12284, n12285, n12286, n12287, n12288,
    n12289, n12290, n12291, n12292, n12293, n12294,
    n12295, n12296, n12297, n12298, n12299, n12300,
    n12301, n12302, n12303, n12304, n12305, n12306,
    n12307, n12308, n12309, n12310, n12311, n12312,
    n12313, n12314, n12315, n12316, n12317, n12318,
    n12319, n12320, n12321, n12322, n12323, n12324,
    n12325, n12326, n12327, n12328, n12329, n12330,
    n12331, n12332, n12333, n12334, n12335, n12336,
    n12337, n12338, n12339, n12340, n12341, n12342,
    n12343, n12344, n12345, n12346, n12347, n12348,
    n12349, n12350, n12351, n12352, n12353, n12354,
    n12355, n12356, n12357, n12358, n12359, n12360,
    n12361, n12362, n12363, n12364, n12365, n12366,
    n12367, n12368, n12369, n12370, n12371, n12372,
    n12373, n12374, n12375, n12376, n12377, n12378,
    n12379, n12380, n12381, n12382, n12383, n12384,
    n12385, n12386, n12387, n12388, n12389, n12390,
    n12391, n12392, n12393, n12394, n12395, n12396,
    n12397, n12398, n12399, n12400, n12401, n12402,
    n12403, n12404, n12405, n12406, n12407, n12408,
    n12409, n12410, n12411, n12412, n12413, n12414,
    n12415, n12416, n12417, n12418, n12419, n12420,
    n12421, n12422, n12423, n12424, n12425, n12426,
    n12427, n12428, n12429, n12430, n12431, n12432,
    n12433, n12434, n12435, n12436, n12437, n12438,
    n12439, n12440, n12441, n12442, n12443, n12444,
    n12445, n12446, n12447, n12448, n12449, n12450,
    n12451, n12452, n12453, n12454, n12455, n12456,
    n12457, n12458, n12459, n12460, n12461, n12462,
    n12463, n12464, n12465, n12466, n12467, n12468,
    n12469, n12470, n12471, n12472, n12473, n12474,
    n12475, n12476, n12477, n12478, n12479, n12480,
    n12481, n12482, n12483, n12484, n12485, n12486,
    n12487, n12488, n12489, n12490, n12491, n12492,
    n12493, n12494, n12495, n12496, n12497, n12498,
    n12499, n12500, n12501, n12502, n12503, n12504,
    n12505, n12506, n12507, n12508, n12509, n12510,
    n12511, n12512, n12513, n12514, n12515, n12516,
    n12517, n12518, n12519, n12520, n12521, n12522,
    n12523, n12524, n12525, n12526, n12527, n12528,
    n12529, n12530, n12531, n12532, n12533, n12534,
    n12535, n12536, n12537, n12538, n12539, n12540,
    n12541, n12542, n12543, n12544, n12545, n12546,
    n12547, n12548, n12549, n12550, n12551, n12552,
    n12553, n12554, n12555, n12556, n12557, n12559,
    n12560, n12561, n12562, n12563, n12564, n12565,
    n12566, n12567, n12568, n12569, n12570, n12571,
    n12572, n12573, n12574, n12575, n12576, n12577,
    n12578, n12579, n12580, n12581, n12582, n12583,
    n12584, n12585, n12586, n12587, n12588, n12589,
    n12590, n12591, n12592, n12593, n12594, n12595,
    n12596, n12597, n12598, n12599, n12600, n12601,
    n12602, n12603, n12604, n12605, n12606, n12607,
    n12608, n12609, n12610, n12611, n12612, n12613,
    n12614, n12615, n12616, n12617, n12618, n12619,
    n12620, n12621, n12622, n12623, n12624, n12625,
    n12626, n12627, n12628, n12629, n12630, n12631,
    n12632, n12633, n12634, n12635, n12636, n12637,
    n12638, n12639, n12640, n12641, n12642, n12643,
    n12644, n12645, n12646, n12647, n12648, n12649,
    n12650, n12651, n12652, n12653, n12654, n12655,
    n12656, n12657, n12658, n12659, n12660, n12661,
    n12662, n12663, n12664, n12665, n12666, n12667,
    n12668, n12669, n12670, n12671, n12672, n12673,
    n12674, n12675, n12676, n12677, n12678, n12679,
    n12680, n12681, n12682, n12683, n12684, n12685,
    n12686, n12687, n12688, n12689, n12690, n12691,
    n12692, n12693, n12694, n12695, n12696, n12697,
    n12698, n12699, n12700, n12701, n12702, n12703,
    n12704, n12705, n12706, n12707, n12708, n12709,
    n12710, n12711, n12712, n12713, n12714, n12715,
    n12716, n12717, n12718, n12719, n12720, n12721,
    n12722, n12723, n12724, n12725, n12726, n12727,
    n12728, n12729, n12730, n12731, n12732, n12733,
    n12734, n12735, n12736, n12737, n12738, n12739,
    n12740, n12741, n12742, n12743, n12744, n12745,
    n12746, n12747, n12748, n12749, n12750, n12751,
    n12752, n12753, n12754, n12755, n12756, n12757,
    n12758, n12759, n12760, n12761, n12762, n12763,
    n12764, n12765, n12766, n12767, n12768, n12769,
    n12770, n12771, n12772, n12773, n12774, n12775,
    n12776, n12777, n12778, n12779, n12780, n12781,
    n12782, n12783, n12784, n12785, n12786, n12787,
    n12788, n12789, n12790, n12791, n12792, n12793,
    n12794, n12795, n12796, n12797, n12798, n12799,
    n12800, n12801, n12802, n12803, n12804, n12805,
    n12806, n12807, n12808, n12809, n12810, n12811,
    n12812, n12813, n12814, n12815, n12816, n12817,
    n12818, n12819, n12820, n12821, n12822, n12823,
    n12824, n12825, n12826, n12827, n12828, n12829,
    n12830, n12831, n12832, n12833, n12834, n12835,
    n12836, n12837, n12838, n12839, n12840, n12841,
    n12842, n12843, n12844, n12845, n12846, n12847,
    n12848, n12849, n12850, n12851, n12852, n12853,
    n12854, n12855, n12856, n12857, n12858, n12859,
    n12860, n12861, n12862, n12863, n12864, n12865,
    n12866, n12867, n12868, n12869, n12870, n12871,
    n12872, n12873, n12874, n12875, n12876, n12877,
    n12878, n12879, n12880, n12881, n12882, n12883,
    n12884, n12885, n12886, n12887, n12888, n12889,
    n12890, n12891, n12892, n12893, n12894, n12895,
    n12896, n12897, n12898, n12899, n12900, n12901,
    n12902, n12903, n12904, n12905, n12906, n12907,
    n12908, n12909, n12910, n12911, n12912, n12913,
    n12914, n12915, n12916, n12917, n12918, n12919,
    n12920, n12921, n12922, n12923, n12924, n12925,
    n12926, n12927, n12928, n12929, n12930, n12931,
    n12932, n12933, n12934, n12935, n12936, n12937,
    n12938, n12939, n12940, n12941, n12942, n12943,
    n12944, n12945, n12946, n12947, n12948, n12949,
    n12950, n12951, n12952, n12953, n12954, n12955,
    n12956, n12957, n12958, n12959, n12960, n12961,
    n12962, n12963, n12964, n12965, n12967, n12968,
    n12969, n12970, n12971, n12972, n12973, n12974,
    n12975, n12976, n12977, n12978, n12979, n12980,
    n12981, n12982, n12983, n12984, n12985, n12986,
    n12987, n12988, n12989, n12990, n12991, n12992,
    n12993, n12994, n12995, n12996, n12997, n12998,
    n12999, n13000, n13001, n13002, n13003, n13004,
    n13005, n13006, n13007, n13008, n13009, n13010,
    n13011, n13012, n13013, n13014, n13015, n13016,
    n13017, n13018, n13019, n13020, n13021, n13022,
    n13023, n13024, n13025, n13026, n13027, n13028,
    n13029, n13030, n13031, n13032, n13033, n13034,
    n13035, n13036, n13037, n13038, n13039, n13040,
    n13041, n13042, n13043, n13044, n13045, n13046,
    n13047, n13048, n13049, n13050, n13051, n13052,
    n13053, n13054, n13055, n13056, n13057, n13058,
    n13059, n13060, n13061, n13062, n13063, n13064,
    n13065, n13066, n13067, n13068, n13069, n13070,
    n13071, n13072, n13073, n13074, n13075, n13076,
    n13077, n13078, n13079, n13080, n13081, n13082,
    n13083, n13084, n13085, n13086, n13087, n13088,
    n13089, n13090, n13091, n13092, n13093, n13094,
    n13095, n13096, n13097, n13098, n13099, n13100,
    n13101, n13102, n13103, n13104, n13105, n13106,
    n13107, n13108, n13109, n13110, n13111, n13112,
    n13113, n13114, n13115, n13116, n13117, n13118,
    n13119, n13120, n13121, n13122, n13123, n13124,
    n13125, n13126, n13127, n13128, n13129, n13130,
    n13131, n13132, n13133, n13134, n13135, n13136,
    n13137, n13138, n13139, n13140, n13141, n13142,
    n13143, n13144, n13145, n13146, n13147, n13148,
    n13149, n13150, n13151, n13152, n13153, n13154,
    n13155, n13156, n13157, n13158, n13159, n13160,
    n13161, n13162, n13163, n13164, n13165, n13166,
    n13167, n13168, n13169, n13170, n13171, n13172,
    n13173, n13174, n13175, n13176, n13177, n13178,
    n13179, n13180, n13181, n13182, n13183, n13184,
    n13185, n13186, n13187, n13188, n13189, n13190,
    n13191, n13192, n13193, n13194, n13195, n13196,
    n13197, n13198, n13199, n13200, n13201, n13202,
    n13203, n13204, n13205, n13206, n13207, n13208,
    n13209, n13210, n13211, n13212, n13213, n13214,
    n13215, n13216, n13217, n13218, n13219, n13220,
    n13221, n13222, n13223, n13224, n13225, n13226,
    n13227, n13228, n13229, n13230, n13231, n13232,
    n13233, n13234, n13235, n13236, n13237, n13238,
    n13239, n13240, n13241, n13242, n13243, n13244,
    n13245, n13246, n13247, n13248, n13249, n13250,
    n13251, n13252, n13253, n13254, n13255, n13256,
    n13257, n13258, n13259, n13260, n13261, n13262,
    n13263, n13264, n13265, n13266, n13267, n13268,
    n13269, n13270, n13271, n13272, n13273, n13274,
    n13275, n13276, n13277, n13278, n13279, n13280,
    n13281, n13282, n13283, n13284, n13285, n13286,
    n13287, n13288, n13289, n13290, n13291, n13292,
    n13293, n13294, n13295, n13296, n13297, n13298,
    n13299, n13300, n13301, n13302, n13303, n13304,
    n13305, n13306, n13307, n13308, n13309, n13310,
    n13311, n13312, n13313, n13314, n13315, n13316,
    n13317, n13318, n13319, n13320, n13321, n13322,
    n13323, n13324, n13325, n13326, n13327, n13328,
    n13329, n13330, n13331, n13332, n13333, n13334,
    n13335, n13336, n13337, n13338, n13339, n13340,
    n13341, n13342, n13343, n13344, n13345, n13346,
    n13347, n13348, n13349, n13350, n13351, n13352,
    n13353, n13354, n13355, n13356, n13357, n13358,
    n13359, n13360, n13361, n13362, n13363, n13365,
    n13366, n13367, n13368, n13369, n13370, n13371,
    n13372, n13373, n13374, n13375, n13376, n13377,
    n13378, n13379, n13380, n13381, n13382, n13383,
    n13384, n13385, n13386, n13387, n13388, n13389,
    n13390, n13391, n13392, n13393, n13394, n13395,
    n13396, n13397, n13398, n13399, n13400, n13401,
    n13402, n13403, n13404, n13405, n13406, n13407,
    n13408, n13409, n13410, n13411, n13412, n13413,
    n13414, n13415, n13416, n13417, n13418, n13419,
    n13420, n13421, n13422, n13423, n13424, n13425,
    n13426, n13427, n13428, n13429, n13430, n13431,
    n13432, n13433, n13434, n13435, n13436, n13437,
    n13438, n13439, n13440, n13441, n13442, n13443,
    n13444, n13445, n13446, n13447, n13448, n13449,
    n13450, n13451, n13452, n13453, n13454, n13455,
    n13456, n13457, n13458, n13459, n13460, n13461,
    n13462, n13463, n13464, n13465, n13466, n13467,
    n13468, n13469, n13470, n13471, n13472, n13473,
    n13474, n13475, n13476, n13477, n13478, n13479,
    n13480, n13481, n13482, n13483, n13484, n13485,
    n13486, n13487, n13488, n13489, n13490, n13491,
    n13492, n13493, n13494, n13495, n13496, n13497,
    n13498, n13499, n13500, n13501, n13502, n13503,
    n13504, n13505, n13506, n13507, n13508, n13509,
    n13510, n13511, n13512, n13513, n13514, n13515,
    n13516, n13517, n13518, n13519, n13520, n13521,
    n13522, n13523, n13524, n13525, n13526, n13527,
    n13528, n13529, n13530, n13531, n13532, n13533,
    n13534, n13535, n13536, n13537, n13538, n13539,
    n13540, n13541, n13542, n13543, n13544, n13545,
    n13546, n13547, n13548, n13549, n13550, n13551,
    n13552, n13553, n13554, n13555, n13556, n13557,
    n13558, n13559, n13560, n13561, n13562, n13563,
    n13564, n13565, n13566, n13567, n13568, n13569,
    n13570, n13571, n13572, n13573, n13574, n13575,
    n13576, n13577, n13578, n13579, n13580, n13581,
    n13582, n13583, n13584, n13585, n13586, n13587,
    n13588, n13589, n13590, n13591, n13592, n13593,
    n13594, n13595, n13596, n13597, n13598, n13599,
    n13600, n13601, n13602, n13603, n13604, n13605,
    n13606, n13607, n13608, n13609, n13610, n13611,
    n13612, n13613, n13614, n13615, n13616, n13617,
    n13618, n13619, n13620, n13621, n13622, n13623,
    n13624, n13625, n13626, n13627, n13628, n13629,
    n13630, n13631, n13632, n13633, n13634, n13635,
    n13636, n13637, n13638, n13639, n13640, n13641,
    n13642, n13643, n13644, n13645, n13646, n13647,
    n13648, n13649, n13650, n13651, n13652, n13653,
    n13654, n13655, n13656, n13657, n13658, n13659,
    n13660, n13661, n13662, n13663, n13664, n13665,
    n13666, n13667, n13668, n13669, n13670, n13671,
    n13672, n13673, n13674, n13675, n13676, n13677,
    n13678, n13679, n13680, n13681, n13682, n13683,
    n13684, n13685, n13686, n13687, n13688, n13689,
    n13690, n13691, n13692, n13693, n13694, n13695,
    n13696, n13697, n13698, n13699, n13700, n13701,
    n13702, n13703, n13704, n13705, n13706, n13707,
    n13708, n13709, n13710, n13711, n13712, n13713,
    n13714, n13715, n13716, n13717, n13718, n13719,
    n13720, n13721, n13722, n13723, n13724, n13725,
    n13726, n13727, n13728, n13729, n13730, n13731,
    n13732, n13733, n13734, n13735, n13736, n13737,
    n13738, n13739, n13740, n13741, n13742, n13743,
    n13744, n13745, n13746, n13747, n13748, n13749,
    n13750, n13751, n13752, n13753, n13754, n13755,
    n13756, n13757, n13758, n13759, n13760, n13761,
    n13762, n13763, n13764, n13765, n13767, n13768,
    n13769, n13770, n13771, n13772, n13773, n13774,
    n13775, n13776, n13777, n13778, n13779, n13780,
    n13781, n13782, n13783, n13784, n13785, n13786,
    n13787, n13788, n13789, n13790, n13791, n13792,
    n13793, n13794, n13795, n13796, n13797, n13798,
    n13799, n13800, n13801, n13802, n13803, n13804,
    n13805, n13806, n13807, n13808, n13809, n13810,
    n13811, n13812, n13813, n13814, n13815, n13816,
    n13817, n13818, n13819, n13820, n13821, n13822,
    n13823, n13824, n13825, n13826, n13827, n13828,
    n13829, n13830, n13831, n13832, n13833, n13834,
    n13835, n13836, n13837, n13838, n13839, n13840,
    n13841, n13842, n13843, n13844, n13845, n13846,
    n13847, n13848, n13849, n13850, n13851, n13852,
    n13853, n13854, n13855, n13856, n13857, n13858,
    n13859, n13860, n13861, n13862, n13863, n13864,
    n13865, n13866, n13867, n13868, n13869, n13870,
    n13871, n13872, n13873, n13874, n13875, n13876,
    n13877, n13878, n13879, n13880, n13881, n13882,
    n13883, n13884, n13885, n13886, n13887, n13888,
    n13889, n13890, n13891, n13892, n13893, n13894,
    n13895, n13896, n13897, n13898, n13899, n13900,
    n13901, n13902, n13903, n13904, n13905, n13906,
    n13907, n13908, n13909, n13910, n13911, n13912,
    n13913, n13914, n13915, n13916, n13917, n13918,
    n13919, n13920, n13921, n13922, n13923, n13924,
    n13925, n13926, n13927, n13928, n13929, n13930,
    n13931, n13932, n13933, n13934, n13935, n13936,
    n13937, n13938, n13939, n13940, n13941, n13942,
    n13943, n13944, n13945, n13946, n13947, n13948,
    n13949, n13950, n13951, n13952, n13953, n13954,
    n13955, n13956, n13957, n13958, n13959, n13960,
    n13961, n13962, n13963, n13964, n13965, n13966,
    n13967, n13968, n13969, n13970, n13971, n13972,
    n13973, n13974, n13975, n13976, n13977, n13978,
    n13979, n13980, n13981, n13982, n13983, n13984,
    n13985, n13986, n13987, n13988, n13989, n13990,
    n13991, n13992, n13993, n13994, n13995, n13996,
    n13997, n13998, n13999, n14000, n14001, n14002,
    n14003, n14004, n14005, n14006, n14007, n14008,
    n14009, n14010, n14011, n14012, n14013, n14014,
    n14015, n14016, n14017, n14018, n14019, n14020,
    n14021, n14022, n14023, n14024, n14025, n14026,
    n14027, n14028, n14029, n14030, n14031, n14032,
    n14033, n14034, n14035, n14036, n14037, n14038,
    n14039, n14040, n14041, n14042, n14043, n14044,
    n14045, n14046, n14047, n14048, n14049, n14050,
    n14051, n14052, n14053, n14054, n14055, n14056,
    n14057, n14058, n14059, n14060, n14061, n14062,
    n14063, n14064, n14065, n14066, n14067, n14068,
    n14069, n14070, n14071, n14072, n14073, n14074,
    n14075, n14076, n14077, n14078, n14079, n14080,
    n14081, n14082, n14083, n14084, n14085, n14086,
    n14087, n14088, n14089, n14090, n14091, n14092,
    n14093, n14094, n14095, n14096, n14097, n14098,
    n14099, n14100, n14101, n14102, n14103, n14104,
    n14105, n14106, n14107, n14108, n14109, n14110,
    n14111, n14112, n14113, n14114, n14115, n14116,
    n14117, n14118, n14119, n14120, n14121, n14122,
    n14123, n14124, n14125, n14126, n14127, n14128,
    n14129, n14130, n14131, n14132, n14133, n14134,
    n14135, n14136, n14137, n14138, n14139, n14140,
    n14141, n14142, n14143, n14144, n14145, n14146,
    n14147, n14148, n14149, n14150, n14151, n14152,
    n14153, n14154, n14155, n14156, n14157, n14158,
    n14159, n14160, n14161, n14162, n14163, n14164,
    n14165, n14166, n14168, n14169, n14170, n14171,
    n14172, n14173, n14174, n14175, n14176, n14177,
    n14178, n14179, n14180, n14181, n14182, n14183,
    n14184, n14185, n14186, n14187, n14188, n14189,
    n14190, n14191, n14192, n14193, n14194, n14195,
    n14196, n14197, n14198, n14199, n14200, n14201,
    n14202, n14203, n14204, n14205, n14206, n14207,
    n14208, n14209, n14210, n14211, n14212, n14213,
    n14214, n14215, n14216, n14217, n14218, n14219,
    n14220, n14221, n14222, n14223, n14224, n14225,
    n14226, n14227, n14228, n14229, n14230, n14231,
    n14232, n14233, n14234, n14235, n14236, n14237,
    n14238, n14239, n14240, n14241, n14242, n14243,
    n14244, n14245, n14246, n14247, n14248, n14249,
    n14250, n14251, n14252, n14253, n14254, n14255,
    n14256, n14257, n14258, n14259, n14260, n14261,
    n14262, n14263, n14264, n14265, n14266, n14267,
    n14268, n14269, n14270, n14271, n14272, n14273,
    n14274, n14275, n14276, n14277, n14278, n14279,
    n14280, n14281, n14282, n14283, n14284, n14285,
    n14286, n14287, n14288, n14289, n14290, n14291,
    n14292, n14293, n14294, n14295, n14296, n14297,
    n14298, n14299, n14300, n14301, n14302, n14303,
    n14304, n14305, n14306, n14307, n14308, n14309,
    n14310, n14311, n14312, n14313, n14314, n14315,
    n14316, n14317, n14318, n14319, n14320, n14321,
    n14322, n14323, n14324, n14325, n14326, n14327,
    n14328, n14329, n14330, n14331, n14332, n14333,
    n14334, n14335, n14336, n14337, n14338, n14339,
    n14340, n14341, n14342, n14343, n14344, n14345,
    n14346, n14347, n14348, n14349, n14350, n14351,
    n14352, n14353, n14354, n14355, n14356, n14357,
    n14358, n14359, n14360, n14361, n14362, n14363,
    n14364, n14365, n14366, n14367, n14368, n14369,
    n14370, n14371, n14372, n14373, n14374, n14375,
    n14376, n14377, n14378, n14379, n14380, n14381,
    n14382, n14383, n14384, n14385, n14386, n14387,
    n14388, n14389, n14390, n14391, n14392, n14393,
    n14394, n14395, n14396, n14397, n14398, n14399,
    n14400, n14401, n14402, n14403, n14404, n14405,
    n14406, n14407, n14408, n14409, n14410, n14411,
    n14412, n14413, n14414, n14415, n14416, n14417,
    n14418, n14419, n14420, n14421, n14422, n14423,
    n14424, n14425, n14426, n14427, n14428, n14429,
    n14430, n14431, n14432, n14433, n14434, n14435,
    n14436, n14437, n14438, n14439, n14440, n14441,
    n14442, n14443, n14444, n14445, n14446, n14447,
    n14448, n14449, n14450, n14451, n14452, n14453,
    n14454, n14455, n14456, n14457, n14458, n14459,
    n14460, n14461, n14462, n14463, n14464, n14465,
    n14466, n14467, n14468, n14469, n14470, n14471,
    n14472, n14473, n14474, n14475, n14476, n14477,
    n14478, n14479, n14480, n14481, n14482, n14483,
    n14484, n14485, n14486, n14487, n14488, n14489,
    n14490, n14491, n14492, n14493, n14494, n14495,
    n14496, n14497, n14498, n14499, n14500, n14501,
    n14502, n14503, n14504, n14505, n14506, n14507,
    n14508, n14509, n14510, n14511, n14512, n14513,
    n14514, n14515, n14516, n14517, n14518, n14519,
    n14520, n14521, n14522, n14523, n14524, n14525,
    n14526, n14527, n14528, n14529, n14530, n14531,
    n14532, n14533, n14534, n14535, n14536, n14537,
    n14538, n14539, n14540, n14541, n14542, n14543,
    n14544, n14545, n14546, n14547, n14548, n14549,
    n14550, n14551, n14552, n14553, n14554, n14555,
    n14556, n14557, n14558, n14559, n14560, n14561,
    n14562, n14563, n14564, n14566, n14567, n14568,
    n14569, n14570, n14571, n14572, n14573, n14574,
    n14575, n14576, n14577, n14578, n14579, n14580,
    n14581, n14582, n14583, n14584, n14585, n14586,
    n14587, n14588, n14589, n14590, n14591, n14592,
    n14593, n14594, n14595, n14596, n14597, n14598,
    n14599, n14600, n14601, n14602, n14603, n14604,
    n14605, n14606, n14607, n14608, n14609, n14610,
    n14611, n14612, n14613, n14614, n14615, n14616,
    n14617, n14618, n14619, n14620, n14621, n14622,
    n14623, n14624, n14625, n14626, n14627, n14628,
    n14629, n14630, n14631, n14632, n14633, n14634,
    n14635, n14636, n14637, n14638, n14639, n14640,
    n14641, n14642, n14643, n14644, n14645, n14646,
    n14647, n14648, n14649, n14650, n14651, n14652,
    n14653, n14654, n14655, n14656, n14657, n14658,
    n14659, n14660, n14661, n14662, n14663, n14664,
    n14665, n14666, n14667, n14668, n14669, n14670,
    n14671, n14672, n14673, n14674, n14675, n14676,
    n14677, n14678, n14679, n14680, n14681, n14682,
    n14683, n14684, n14685, n14686, n14687, n14688,
    n14689, n14690, n14691, n14692, n14693, n14694,
    n14695, n14696, n14697, n14698, n14699, n14700,
    n14701, n14702, n14703, n14704, n14705, n14706,
    n14707, n14708, n14709, n14710, n14711, n14712,
    n14713, n14714, n14715, n14716, n14717, n14718,
    n14719, n14720, n14721, n14722, n14723, n14724,
    n14725, n14726, n14727, n14728, n14729, n14730,
    n14731, n14732, n14733, n14734, n14735, n14736,
    n14737, n14738, n14739, n14740, n14741, n14742,
    n14743, n14744, n14745, n14746, n14747, n14748,
    n14749, n14750, n14751, n14752, n14753, n14754,
    n14755, n14756, n14757, n14758, n14759, n14760,
    n14761, n14762, n14763, n14764, n14765, n14766,
    n14767, n14768, n14769, n14770, n14771, n14772,
    n14773, n14774, n14775, n14776, n14777, n14778,
    n14779, n14780, n14781, n14782, n14783, n14784,
    n14785, n14786, n14787, n14788, n14789, n14790,
    n14791, n14792, n14793, n14794, n14795, n14796,
    n14797, n14798, n14799, n14800, n14801, n14802,
    n14803, n14804, n14805, n14806, n14807, n14808,
    n14809, n14810, n14811, n14812, n14813, n14814,
    n14815, n14816, n14817, n14818, n14819, n14820,
    n14821, n14822, n14823, n14824, n14825, n14826,
    n14827, n14828, n14829, n14830, n14831, n14832,
    n14833, n14834, n14835, n14836, n14837, n14838,
    n14839, n14840, n14841, n14842, n14843, n14844,
    n14845, n14846, n14847, n14848, n14849, n14850,
    n14851, n14852, n14853, n14854, n14855, n14856,
    n14857, n14858, n14859, n14860, n14861, n14862,
    n14863, n14864, n14865, n14866, n14867, n14868,
    n14869, n14870, n14871, n14872, n14873, n14874,
    n14875, n14876, n14877, n14878, n14879, n14880,
    n14881, n14882, n14883, n14884, n14885, n14886,
    n14887, n14888, n14889, n14890, n14891, n14892,
    n14893, n14894, n14895, n14896, n14897, n14898,
    n14899, n14900, n14901, n14902, n14903, n14904,
    n14905, n14906, n14907, n14908, n14909, n14910,
    n14911, n14912, n14913, n14914, n14915, n14916,
    n14917, n14918, n14919, n14920, n14921, n14922,
    n14923, n14924, n14925, n14926, n14927, n14928,
    n14929, n14930, n14931, n14932, n14933, n14934,
    n14935, n14936, n14937, n14938, n14939, n14940,
    n14941, n14942, n14943, n14944, n14945, n14946,
    n14947, n14948, n14949, n14950, n14951, n14953,
    n14954, n14955, n14956, n14957, n14958, n14959,
    n14960, n14961, n14962, n14963, n14964, n14965,
    n14966, n14967, n14968, n14969, n14970, n14971,
    n14972, n14973, n14974, n14975, n14976, n14977,
    n14978, n14979, n14980, n14981, n14982, n14983,
    n14984, n14985, n14986, n14987, n14988, n14989,
    n14990, n14991, n14992, n14993, n14994, n14995,
    n14996, n14997, n14998, n14999, n15000, n15001,
    n15002, n15003, n15004, n15005, n15006, n15007,
    n15008, n15009, n15010, n15011, n15012, n15013,
    n15014, n15015, n15016, n15017, n15018, n15019,
    n15020, n15021, n15022, n15023, n15024, n15025,
    n15026, n15027, n15028, n15029, n15030, n15031,
    n15032, n15033, n15034, n15035, n15036, n15037,
    n15038, n15039, n15040, n15041, n15042, n15043,
    n15044, n15045, n15046, n15047, n15048, n15049,
    n15050, n15051, n15052, n15053, n15054, n15055,
    n15056, n15057, n15058, n15059, n15060, n15061,
    n15062, n15063, n15064, n15065, n15066, n15067,
    n15068, n15069, n15070, n15071, n15072, n15073,
    n15074, n15075, n15076, n15077, n15078, n15079,
    n15080, n15081, n15082, n15083, n15084, n15085,
    n15086, n15087, n15088, n15089, n15090, n15091,
    n15092, n15093, n15094, n15095, n15096, n15097,
    n15098, n15099, n15100, n15101, n15102, n15103,
    n15104, n15105, n15106, n15107, n15108, n15109,
    n15110, n15111, n15112, n15113, n15114, n15115,
    n15116, n15117, n15118, n15119, n15120, n15121,
    n15122, n15123, n15124, n15125, n15126, n15127,
    n15128, n15129, n15130, n15131, n15132, n15133,
    n15134, n15135, n15136, n15137, n15138, n15139,
    n15140, n15141, n15142, n15143, n15144, n15145,
    n15146, n15147, n15148, n15149, n15150, n15151,
    n15152, n15153, n15154, n15155, n15156, n15157,
    n15158, n15159, n15160, n15161, n15162, n15163,
    n15164, n15165, n15166, n15167, n15168, n15169,
    n15170, n15171, n15172, n15173, n15174, n15175,
    n15176, n15177, n15178, n15179, n15180, n15181,
    n15182, n15183, n15184, n15185, n15186, n15187,
    n15188, n15189, n15190, n15191, n15192, n15193,
    n15194, n15195, n15196, n15197, n15198, n15199,
    n15200, n15201, n15202, n15203, n15204, n15205,
    n15206, n15207, n15208, n15209, n15210, n15211,
    n15212, n15213, n15214, n15215, n15216, n15217,
    n15218, n15219, n15220, n15221, n15222, n15223,
    n15224, n15225, n15226, n15227, n15228, n15229,
    n15230, n15231, n15232, n15233, n15234, n15235,
    n15236, n15237, n15238, n15239, n15240, n15241,
    n15242, n15243, n15244, n15245, n15246, n15247,
    n15248, n15249, n15250, n15251, n15252, n15253,
    n15254, n15255, n15256, n15257, n15258, n15259,
    n15260, n15261, n15262, n15263, n15264, n15265,
    n15266, n15267, n15268, n15269, n15270, n15271,
    n15272, n15273, n15274, n15275, n15276, n15277,
    n15278, n15279, n15280, n15281, n15282, n15283,
    n15284, n15285, n15286, n15287, n15288, n15289,
    n15290, n15291, n15292, n15293, n15294, n15295,
    n15296, n15297, n15298, n15299, n15300, n15301,
    n15302, n15303, n15304, n15305, n15306, n15307,
    n15308, n15309, n15310, n15311, n15312, n15313,
    n15314, n15315, n15316, n15317, n15318, n15319,
    n15320, n15321, n15322, n15323, n15324, n15325,
    n15326, n15327, n15328, n15329, n15330, n15331,
    n15332, n15333, n15334, n15335, n15336, n15337,
    n15338, n15339, n15340, n15341, n15342, n15343,
    n15344, n15345, n15347, n15348, n15349, n15350,
    n15351, n15352, n15353, n15354, n15355, n15356,
    n15357, n15358, n15359, n15360, n15361, n15362,
    n15363, n15364, n15365, n15366, n15367, n15368,
    n15369, n15370, n15371, n15372, n15373, n15374,
    n15375, n15376, n15377, n15378, n15379, n15380,
    n15381, n15382, n15383, n15384, n15385, n15386,
    n15387, n15388, n15389, n15390, n15391, n15392,
    n15393, n15394, n15395, n15396, n15397, n15398,
    n15399, n15400, n15401, n15402, n15403, n15404,
    n15405, n15406, n15407, n15408, n15409, n15410,
    n15411, n15412, n15413, n15414, n15415, n15416,
    n15417, n15418, n15419, n15420, n15421, n15422,
    n15423, n15424, n15425, n15426, n15427, n15428,
    n15429, n15430, n15431, n15432, n15433, n15434,
    n15435, n15436, n15437, n15438, n15439, n15440,
    n15441, n15442, n15443, n15444, n15445, n15446,
    n15447, n15448, n15449, n15450, n15451, n15452,
    n15453, n15454, n15455, n15456, n15457, n15458,
    n15459, n15460, n15461, n15462, n15463, n15464,
    n15465, n15466, n15467, n15468, n15469, n15470,
    n15471, n15472, n15473, n15474, n15475, n15476,
    n15477, n15478, n15479, n15480, n15481, n15482,
    n15483, n15484, n15485, n15486, n15487, n15488,
    n15489, n15490, n15491, n15492, n15493, n15494,
    n15495, n15496, n15497, n15498, n15499, n15500,
    n15501, n15502, n15503, n15504, n15505, n15506,
    n15507, n15508, n15509, n15510, n15511, n15512,
    n15513, n15514, n15515, n15516, n15517, n15518,
    n15519, n15520, n15521, n15522, n15523, n15524,
    n15525, n15526, n15527, n15528, n15529, n15530,
    n15531, n15532, n15533, n15534, n15535, n15536,
    n15537, n15538, n15539, n15540, n15541, n15542,
    n15543, n15544, n15545, n15546, n15547, n15548,
    n15549, n15550, n15551, n15552, n15553, n15554,
    n15555, n15556, n15557, n15558, n15559, n15560,
    n15561, n15562, n15563, n15564, n15565, n15566,
    n15567, n15568, n15569, n15570, n15571, n15572,
    n15573, n15574, n15575, n15576, n15577, n15578,
    n15579, n15580, n15581, n15582, n15583, n15584,
    n15585, n15586, n15587, n15588, n15589, n15590,
    n15591, n15592, n15593, n15594, n15595, n15596,
    n15597, n15598, n15599, n15600, n15601, n15602,
    n15603, n15604, n15605, n15606, n15607, n15608,
    n15609, n15610, n15611, n15612, n15613, n15614,
    n15615, n15616, n15617, n15618, n15619, n15620,
    n15621, n15622, n15623, n15624, n15625, n15626,
    n15627, n15628, n15629, n15630, n15631, n15632,
    n15633, n15634, n15635, n15636, n15637, n15638,
    n15639, n15640, n15641, n15642, n15643, n15644,
    n15645, n15646, n15647, n15648, n15649, n15650,
    n15651, n15652, n15653, n15654, n15655, n15656,
    n15657, n15658, n15659, n15660, n15661, n15662,
    n15663, n15664, n15665, n15666, n15667, n15668,
    n15669, n15670, n15671, n15672, n15673, n15674,
    n15675, n15676, n15677, n15678, n15679, n15680,
    n15681, n15682, n15683, n15684, n15685, n15686,
    n15687, n15688, n15689, n15690, n15691, n15692,
    n15693, n15694, n15695, n15696, n15697, n15698,
    n15699, n15700, n15701, n15702, n15703, n15704,
    n15705, n15706, n15707, n15708, n15709, n15710,
    n15711, n15712, n15713, n15714, n15715, n15716,
    n15717, n15718, n15719, n15720, n15721, n15722,
    n15723, n15724, n15725, n15726, n15727, n15728,
    n15729, n15730, n15731, n15732, n15733, n15734,
    n15736, n15737, n15738, n15739, n15740, n15741,
    n15742, n15743, n15744, n15745, n15746, n15747,
    n15748, n15749, n15750, n15751, n15752, n15753,
    n15754, n15755, n15756, n15757, n15758, n15759,
    n15760, n15761, n15762, n15763, n15764, n15765,
    n15766, n15767, n15768, n15769, n15770, n15771,
    n15772, n15773, n15774, n15775, n15776, n15777,
    n15778, n15779, n15780, n15781, n15782, n15783,
    n15784, n15785, n15786, n15787, n15788, n15789,
    n15790, n15791, n15792, n15793, n15794, n15795,
    n15796, n15797, n15798, n15799, n15800, n15801,
    n15802, n15803, n15804, n15805, n15806, n15807,
    n15808, n15809, n15810, n15811, n15812, n15813,
    n15814, n15815, n15816, n15817, n15818, n15819,
    n15820, n15821, n15822, n15823, n15824, n15825,
    n15826, n15827, n15828, n15829, n15830, n15831,
    n15832, n15833, n15834, n15835, n15836, n15837,
    n15838, n15839, n15840, n15841, n15842, n15843,
    n15844, n15845, n15846, n15847, n15848, n15849,
    n15850, n15851, n15852, n15853, n15854, n15855,
    n15856, n15857, n15858, n15859, n15860, n15861,
    n15862, n15863, n15864, n15865, n15866, n15867,
    n15868, n15869, n15870, n15871, n15872, n15873,
    n15874, n15875, n15876, n15877, n15878, n15879,
    n15880, n15881, n15882, n15883, n15884, n15885,
    n15886, n15887, n15888, n15889, n15890, n15891,
    n15892, n15893, n15894, n15895, n15896, n15897,
    n15898, n15899, n15900, n15901, n15902, n15903,
    n15904, n15905, n15906, n15907, n15908, n15909,
    n15910, n15911, n15912, n15913, n15914, n15915,
    n15916, n15917, n15918, n15919, n15920, n15921,
    n15922, n15923, n15924, n15925, n15926, n15927,
    n15928, n15929, n15930, n15931, n15932, n15933,
    n15934, n15935, n15936, n15937, n15938, n15939,
    n15940, n15941, n15942, n15943, n15944, n15945,
    n15946, n15947, n15948, n15949, n15950, n15951,
    n15952, n15953, n15954, n15955, n15956, n15957,
    n15958, n15959, n15960, n15961, n15962, n15963,
    n15964, n15965, n15966, n15967, n15968, n15969,
    n15970, n15971, n15972, n15973, n15974, n15975,
    n15976, n15977, n15978, n15979, n15980, n15981,
    n15982, n15983, n15984, n15985, n15986, n15987,
    n15988, n15989, n15990, n15991, n15992, n15993,
    n15994, n15995, n15996, n15997, n15998, n15999,
    n16000, n16001, n16002, n16003, n16004, n16005,
    n16006, n16007, n16008, n16009, n16010, n16011,
    n16012, n16013, n16014, n16015, n16016, n16017,
    n16018, n16019, n16020, n16021, n16022, n16023,
    n16024, n16025, n16026, n16027, n16028, n16029,
    n16030, n16031, n16032, n16033, n16034, n16035,
    n16036, n16037, n16038, n16039, n16040, n16041,
    n16042, n16043, n16044, n16045, n16046, n16047,
    n16048, n16049, n16050, n16051, n16052, n16053,
    n16054, n16055, n16056, n16057, n16058, n16059,
    n16060, n16061, n16062, n16063, n16064, n16065,
    n16066, n16067, n16068, n16069, n16070, n16071,
    n16072, n16073, n16074, n16075, n16076, n16077,
    n16078, n16079, n16080, n16081, n16082, n16083,
    n16084, n16085, n16086, n16087, n16088, n16089,
    n16090, n16091, n16092, n16093, n16094, n16095,
    n16096, n16097, n16098, n16099, n16100, n16101,
    n16102, n16103, n16104, n16105, n16106, n16107,
    n16108, n16109, n16110, n16111, n16112, n16114,
    n16115, n16116, n16117, n16118, n16119, n16120,
    n16121, n16122, n16123, n16124, n16125, n16126,
    n16127, n16128, n16129, n16130, n16131, n16132,
    n16133, n16134, n16135, n16136, n16137, n16138,
    n16139, n16140, n16141, n16142, n16143, n16144,
    n16145, n16146, n16147, n16148, n16149, n16150,
    n16151, n16152, n16153, n16154, n16155, n16156,
    n16157, n16158, n16159, n16160, n16161, n16162,
    n16163, n16164, n16165, n16166, n16167, n16168,
    n16169, n16170, n16171, n16172, n16173, n16174,
    n16175, n16176, n16177, n16178, n16179, n16180,
    n16181, n16182, n16183, n16184, n16185, n16186,
    n16187, n16188, n16189, n16190, n16191, n16192,
    n16193, n16194, n16195, n16196, n16197, n16198,
    n16199, n16200, n16201, n16202, n16203, n16204,
    n16205, n16206, n16207, n16208, n16209, n16210,
    n16211, n16212, n16213, n16214, n16215, n16216,
    n16217, n16218, n16219, n16220, n16221, n16222,
    n16223, n16224, n16225, n16226, n16227, n16228,
    n16229, n16230, n16231, n16232, n16233, n16234,
    n16235, n16236, n16237, n16238, n16239, n16240,
    n16241, n16242, n16243, n16244, n16245, n16246,
    n16247, n16248, n16249, n16250, n16251, n16252,
    n16253, n16254, n16255, n16256, n16257, n16258,
    n16259, n16260, n16261, n16262, n16263, n16264,
    n16265, n16266, n16267, n16268, n16269, n16270,
    n16271, n16272, n16273, n16274, n16275, n16276,
    n16277, n16278, n16279, n16280, n16281, n16282,
    n16283, n16284, n16285, n16286, n16287, n16288,
    n16289, n16290, n16291, n16292, n16293, n16294,
    n16295, n16296, n16297, n16298, n16299, n16300,
    n16301, n16302, n16303, n16304, n16305, n16306,
    n16307, n16308, n16309, n16310, n16311, n16312,
    n16313, n16314, n16315, n16316, n16317, n16318,
    n16319, n16320, n16321, n16322, n16323, n16324,
    n16325, n16326, n16327, n16328, n16329, n16330,
    n16331, n16332, n16333, n16334, n16335, n16336,
    n16337, n16338, n16339, n16340, n16341, n16342,
    n16343, n16344, n16345, n16346, n16347, n16348,
    n16349, n16350, n16351, n16352, n16353, n16354,
    n16355, n16356, n16357, n16358, n16359, n16360,
    n16361, n16362, n16363, n16364, n16365, n16366,
    n16367, n16368, n16369, n16370, n16371, n16372,
    n16373, n16374, n16375, n16376, n16377, n16378,
    n16379, n16380, n16381, n16382, n16383, n16384,
    n16385, n16386, n16387, n16388, n16389, n16390,
    n16391, n16392, n16393, n16394, n16395, n16396,
    n16397, n16398, n16399, n16400, n16401, n16402,
    n16403, n16404, n16405, n16406, n16407, n16408,
    n16409, n16410, n16411, n16412, n16413, n16414,
    n16415, n16416, n16417, n16418, n16419, n16420,
    n16421, n16422, n16423, n16424, n16425, n16426,
    n16427, n16428, n16429, n16430, n16431, n16432,
    n16433, n16434, n16435, n16436, n16437, n16438,
    n16439, n16440, n16441, n16442, n16443, n16444,
    n16445, n16446, n16447, n16448, n16449, n16450,
    n16451, n16452, n16453, n16454, n16455, n16456,
    n16457, n16458, n16459, n16460, n16461, n16462,
    n16463, n16464, n16465, n16466, n16467, n16468,
    n16469, n16470, n16471, n16472, n16473, n16474,
    n16475, n16476, n16477, n16478, n16479, n16480,
    n16481, n16482, n16484, n16485, n16486, n16487,
    n16488, n16489, n16490, n16491, n16492, n16493,
    n16494, n16495, n16496, n16497, n16498, n16499,
    n16500, n16501, n16502, n16503, n16504, n16505,
    n16506, n16507, n16508, n16509, n16510, n16511,
    n16512, n16513, n16514, n16515, n16516, n16517,
    n16518, n16519, n16520, n16521, n16522, n16523,
    n16524, n16525, n16526, n16527, n16528, n16529,
    n16530, n16531, n16532, n16533, n16534, n16535,
    n16536, n16537, n16538, n16539, n16540, n16541,
    n16542, n16543, n16544, n16545, n16546, n16547,
    n16548, n16549, n16550, n16551, n16552, n16553,
    n16554, n16555, n16556, n16557, n16558, n16559,
    n16560, n16561, n16562, n16563, n16564, n16565,
    n16566, n16567, n16568, n16569, n16570, n16571,
    n16572, n16573, n16574, n16575, n16576, n16577,
    n16578, n16579, n16580, n16581, n16582, n16583,
    n16584, n16585, n16586, n16587, n16588, n16589,
    n16590, n16591, n16592, n16593, n16594, n16595,
    n16596, n16597, n16598, n16599, n16600, n16601,
    n16602, n16603, n16604, n16605, n16606, n16607,
    n16608, n16609, n16610, n16611, n16612, n16613,
    n16614, n16615, n16616, n16617, n16618, n16619,
    n16620, n16621, n16622, n16623, n16624, n16625,
    n16626, n16627, n16628, n16629, n16630, n16631,
    n16632, n16633, n16634, n16635, n16636, n16637,
    n16638, n16639, n16640, n16641, n16642, n16643,
    n16644, n16645, n16646, n16647, n16648, n16649,
    n16650, n16651, n16652, n16653, n16654, n16655,
    n16656, n16657, n16658, n16659, n16660, n16661,
    n16662, n16663, n16664, n16665, n16666, n16667,
    n16668, n16669, n16670, n16671, n16672, n16673,
    n16674, n16675, n16676, n16677, n16678, n16679,
    n16680, n16681, n16682, n16683, n16684, n16685,
    n16686, n16687, n16688, n16689, n16690, n16691,
    n16692, n16693, n16694, n16695, n16696, n16697,
    n16698, n16699, n16700, n16701, n16702, n16703,
    n16704, n16705, n16706, n16707, n16708, n16709,
    n16710, n16711, n16712, n16713, n16714, n16715,
    n16716, n16717, n16718, n16719, n16720, n16721,
    n16722, n16723, n16724, n16725, n16726, n16727,
    n16728, n16729, n16730, n16731, n16732, n16733,
    n16734, n16735, n16736, n16737, n16738, n16739,
    n16740, n16741, n16742, n16743, n16744, n16745,
    n16746, n16747, n16748, n16749, n16750, n16751,
    n16752, n16753, n16754, n16755, n16756, n16757,
    n16758, n16759, n16760, n16761, n16762, n16763,
    n16764, n16765, n16766, n16767, n16768, n16769,
    n16770, n16771, n16772, n16773, n16774, n16775,
    n16776, n16777, n16778, n16779, n16780, n16781,
    n16782, n16783, n16784, n16785, n16786, n16787,
    n16788, n16789, n16790, n16791, n16792, n16793,
    n16794, n16795, n16796, n16797, n16798, n16799,
    n16800, n16801, n16802, n16803, n16804, n16805,
    n16806, n16807, n16808, n16809, n16810, n16811,
    n16812, n16813, n16814, n16815, n16816, n16817,
    n16818, n16819, n16820, n16821, n16822, n16823,
    n16824, n16825, n16826, n16827, n16828, n16829,
    n16830, n16831, n16832, n16833, n16834, n16835,
    n16836, n16837, n16838, n16839, n16840, n16841,
    n16842, n16843, n16844, n16845, n16846, n16847,
    n16848, n16849, n16850, n16851, n16853, n16854,
    n16855, n16856, n16857, n16858, n16859, n16860,
    n16861, n16862, n16863, n16864, n16865, n16866,
    n16867, n16868, n16869, n16870, n16871, n16872,
    n16873, n16874, n16875, n16876, n16877, n16878,
    n16879, n16880, n16881, n16882, n16883, n16884,
    n16885, n16886, n16887, n16888, n16889, n16890,
    n16891, n16892, n16893, n16894, n16895, n16896,
    n16897, n16898, n16899, n16900, n16901, n16902,
    n16903, n16904, n16905, n16906, n16907, n16908,
    n16909, n16910, n16911, n16912, n16913, n16914,
    n16915, n16916, n16917, n16918, n16919, n16920,
    n16921, n16922, n16923, n16924, n16925, n16926,
    n16927, n16928, n16929, n16930, n16931, n16932,
    n16933, n16934, n16935, n16936, n16937, n16938,
    n16939, n16940, n16941, n16942, n16943, n16944,
    n16945, n16946, n16947, n16948, n16949, n16950,
    n16951, n16952, n16953, n16954, n16955, n16956,
    n16957, n16958, n16959, n16960, n16961, n16962,
    n16963, n16964, n16965, n16966, n16967, n16968,
    n16969, n16970, n16971, n16972, n16973, n16974,
    n16975, n16976, n16977, n16978, n16979, n16980,
    n16981, n16982, n16983, n16984, n16985, n16986,
    n16987, n16988, n16989, n16990, n16991, n16992,
    n16993, n16994, n16995, n16996, n16997, n16998,
    n16999, n17000, n17001, n17002, n17003, n17004,
    n17005, n17006, n17007, n17008, n17009, n17010,
    n17011, n17012, n17013, n17014, n17015, n17016,
    n17017, n17018, n17019, n17020, n17021, n17022,
    n17023, n17024, n17025, n17026, n17027, n17028,
    n17029, n17030, n17031, n17032, n17033, n17034,
    n17035, n17036, n17037, n17038, n17039, n17040,
    n17041, n17042, n17043, n17044, n17045, n17046,
    n17047, n17048, n17049, n17050, n17051, n17052,
    n17053, n17054, n17055, n17056, n17057, n17058,
    n17059, n17060, n17061, n17062, n17063, n17064,
    n17065, n17066, n17067, n17068, n17069, n17070,
    n17071, n17072, n17073, n17074, n17075, n17076,
    n17077, n17078, n17079, n17080, n17081, n17082,
    n17083, n17084, n17085, n17086, n17087, n17088,
    n17089, n17090, n17091, n17092, n17093, n17094,
    n17095, n17096, n17097, n17098, n17099, n17100,
    n17101, n17102, n17103, n17104, n17105, n17106,
    n17107, n17108, n17109, n17110, n17111, n17112,
    n17113, n17114, n17115, n17116, n17117, n17118,
    n17119, n17120, n17121, n17122, n17123, n17124,
    n17125, n17126, n17127, n17128, n17129, n17130,
    n17131, n17132, n17133, n17134, n17135, n17136,
    n17137, n17138, n17139, n17140, n17141, n17142,
    n17143, n17144, n17145, n17146, n17147, n17148,
    n17149, n17150, n17151, n17152, n17153, n17154,
    n17155, n17156, n17157, n17158, n17159, n17160,
    n17161, n17162, n17163, n17164, n17165, n17166,
    n17167, n17168, n17169, n17170, n17171, n17172,
    n17173, n17174, n17175, n17176, n17177, n17178,
    n17179, n17180, n17181, n17182, n17183, n17184,
    n17185, n17186, n17187, n17188, n17189, n17190,
    n17191, n17192, n17193, n17194, n17195, n17196,
    n17197, n17198, n17199, n17200, n17201, n17202,
    n17203, n17204, n17205, n17206, n17207, n17208,
    n17209, n17210, n17211, n17212, n17213, n17215,
    n17216, n17217, n17218, n17219, n17220, n17221,
    n17222, n17223, n17224, n17225, n17226, n17227,
    n17228, n17229, n17230, n17231, n17232, n17233,
    n17234, n17235, n17236, n17237, n17238, n17239,
    n17240, n17241, n17242, n17243, n17244, n17245,
    n17246, n17247, n17248, n17249, n17250, n17251,
    n17252, n17253, n17254, n17255, n17256, n17257,
    n17258, n17259, n17260, n17261, n17262, n17263,
    n17264, n17265, n17266, n17267, n17268, n17269,
    n17270, n17271, n17272, n17273, n17274, n17275,
    n17276, n17277, n17278, n17279, n17280, n17281,
    n17282, n17283, n17284, n17285, n17286, n17287,
    n17288, n17289, n17290, n17291, n17292, n17293,
    n17294, n17295, n17296, n17297, n17298, n17299,
    n17300, n17301, n17302, n17303, n17304, n17305,
    n17306, n17307, n17308, n17309, n17310, n17311,
    n17312, n17313, n17314, n17315, n17316, n17317,
    n17318, n17319, n17320, n17321, n17322, n17323,
    n17324, n17325, n17326, n17327, n17328, n17329,
    n17330, n17331, n17332, n17333, n17334, n17335,
    n17336, n17337, n17338, n17339, n17340, n17341,
    n17342, n17343, n17344, n17345, n17346, n17347,
    n17348, n17349, n17350, n17351, n17352, n17353,
    n17354, n17355, n17356, n17357, n17358, n17359,
    n17360, n17361, n17362, n17363, n17364, n17365,
    n17366, n17367, n17368, n17369, n17370, n17371,
    n17372, n17373, n17374, n17375, n17376, n17377,
    n17378, n17379, n17380, n17381, n17382, n17383,
    n17384, n17385, n17386, n17387, n17388, n17389,
    n17390, n17391, n17392, n17393, n17394, n17395,
    n17396, n17397, n17398, n17399, n17400, n17401,
    n17402, n17403, n17404, n17405, n17406, n17407,
    n17408, n17409, n17410, n17411, n17412, n17413,
    n17414, n17415, n17416, n17417, n17418, n17419,
    n17420, n17421, n17422, n17423, n17424, n17425,
    n17426, n17427, n17428, n17429, n17430, n17431,
    n17432, n17433, n17434, n17435, n17436, n17437,
    n17438, n17439, n17440, n17441, n17442, n17443,
    n17444, n17445, n17446, n17447, n17448, n17449,
    n17450, n17451, n17452, n17453, n17454, n17455,
    n17456, n17457, n17458, n17459, n17460, n17461,
    n17462, n17463, n17464, n17465, n17466, n17467,
    n17468, n17469, n17470, n17471, n17472, n17473,
    n17474, n17475, n17476, n17477, n17478, n17479,
    n17480, n17481, n17482, n17483, n17484, n17485,
    n17486, n17487, n17488, n17489, n17490, n17491,
    n17492, n17493, n17494, n17495, n17496, n17497,
    n17498, n17499, n17500, n17501, n17502, n17503,
    n17504, n17505, n17506, n17507, n17508, n17509,
    n17510, n17511, n17512, n17513, n17514, n17515,
    n17516, n17517, n17518, n17519, n17520, n17521,
    n17522, n17523, n17524, n17525, n17526, n17527,
    n17528, n17529, n17530, n17531, n17532, n17533,
    n17534, n17535, n17536, n17537, n17538, n17539,
    n17540, n17541, n17542, n17543, n17544, n17545,
    n17546, n17547, n17548, n17549, n17550, n17551,
    n17552, n17553, n17554, n17555, n17556, n17557,
    n17558, n17559, n17560, n17561, n17562, n17563,
    n17564, n17565, n17566, n17567, n17568, n17569,
    n17570, n17571, n17572, n17573, n17575, n17576,
    n17577, n17578, n17579, n17580, n17581, n17582,
    n17583, n17584, n17585, n17586, n17587, n17588,
    n17589, n17590, n17591, n17592, n17593, n17594,
    n17595, n17596, n17597, n17598, n17599, n17600,
    n17601, n17602, n17603, n17604, n17605, n17606,
    n17607, n17608, n17609, n17610, n17611, n17612,
    n17613, n17614, n17615, n17616, n17617, n17618,
    n17619, n17620, n17621, n17622, n17623, n17624,
    n17625, n17626, n17627, n17628, n17629, n17630,
    n17631, n17632, n17633, n17634, n17635, n17636,
    n17637, n17638, n17639, n17640, n17641, n17642,
    n17643, n17644, n17645, n17646, n17647, n17648,
    n17649, n17650, n17651, n17652, n17653, n17654,
    n17655, n17656, n17657, n17658, n17659, n17660,
    n17661, n17662, n17663, n17664, n17665, n17666,
    n17667, n17668, n17669, n17670, n17671, n17672,
    n17673, n17674, n17675, n17676, n17677, n17678,
    n17679, n17680, n17681, n17682, n17683, n17684,
    n17685, n17686, n17687, n17688, n17689, n17690,
    n17691, n17692, n17693, n17694, n17695, n17696,
    n17697, n17698, n17699, n17700, n17701, n17702,
    n17703, n17704, n17705, n17706, n17707, n17708,
    n17709, n17710, n17711, n17712, n17713, n17714,
    n17715, n17716, n17717, n17718, n17719, n17720,
    n17721, n17722, n17723, n17724, n17725, n17726,
    n17727, n17728, n17729, n17730, n17731, n17732,
    n17733, n17734, n17735, n17736, n17737, n17738,
    n17739, n17740, n17741, n17742, n17743, n17744,
    n17745, n17746, n17747, n17748, n17749, n17750,
    n17751, n17752, n17753, n17754, n17755, n17756,
    n17757, n17758, n17759, n17760, n17761, n17762,
    n17763, n17764, n17765, n17766, n17767, n17768,
    n17769, n17770, n17771, n17772, n17773, n17774,
    n17775, n17776, n17777, n17778, n17779, n17780,
    n17781, n17782, n17783, n17784, n17785, n17786,
    n17787, n17788, n17789, n17790, n17791, n17792,
    n17793, n17794, n17795, n17796, n17797, n17798,
    n17799, n17800, n17801, n17802, n17803, n17804,
    n17805, n17806, n17807, n17808, n17809, n17810,
    n17811, n17812, n17813, n17814, n17815, n17816,
    n17817, n17818, n17819, n17820, n17821, n17822,
    n17823, n17824, n17825, n17826, n17827, n17828,
    n17829, n17830, n17831, n17832, n17833, n17834,
    n17835, n17836, n17837, n17838, n17839, n17840,
    n17841, n17842, n17843, n17844, n17845, n17846,
    n17847, n17848, n17849, n17850, n17851, n17852,
    n17853, n17854, n17855, n17856, n17857, n17858,
    n17859, n17860, n17861, n17862, n17863, n17864,
    n17865, n17866, n17867, n17868, n17869, n17870,
    n17871, n17872, n17873, n17874, n17875, n17876,
    n17877, n17878, n17879, n17880, n17881, n17882,
    n17883, n17884, n17885, n17886, n17887, n17888,
    n17889, n17890, n17891, n17892, n17893, n17894,
    n17895, n17896, n17897, n17898, n17899, n17900,
    n17901, n17902, n17903, n17904, n17905, n17906,
    n17907, n17908, n17909, n17910, n17911, n17912,
    n17913, n17914, n17915, n17916, n17917, n17918,
    n17919, n17920, n17922, n17923, n17924, n17925,
    n17926, n17927, n17928, n17929, n17930, n17931,
    n17932, n17933, n17934, n17935, n17936, n17937,
    n17938, n17939, n17940, n17941, n17942, n17943,
    n17944, n17945, n17946, n17947, n17948, n17949,
    n17950, n17951, n17952, n17953, n17954, n17955,
    n17956, n17957, n17958, n17959, n17960, n17961,
    n17962, n17963, n17964, n17965, n17966, n17967,
    n17968, n17969, n17970, n17971, n17972, n17973,
    n17974, n17975, n17976, n17977, n17978, n17979,
    n17980, n17981, n17982, n17983, n17984, n17985,
    n17986, n17987, n17988, n17989, n17990, n17991,
    n17992, n17993, n17994, n17995, n17996, n17997,
    n17998, n17999, n18000, n18001, n18002, n18003,
    n18004, n18005, n18006, n18007, n18008, n18009,
    n18010, n18011, n18012, n18013, n18014, n18015,
    n18016, n18017, n18018, n18019, n18020, n18021,
    n18022, n18023, n18024, n18025, n18026, n18027,
    n18028, n18029, n18030, n18031, n18032, n18033,
    n18034, n18035, n18036, n18037, n18038, n18039,
    n18040, n18041, n18042, n18043, n18044, n18045,
    n18046, n18047, n18048, n18049, n18050, n18051,
    n18052, n18053, n18054, n18055, n18056, n18057,
    n18058, n18059, n18060, n18061, n18062, n18063,
    n18064, n18065, n18066, n18067, n18068, n18069,
    n18070, n18071, n18072, n18073, n18074, n18075,
    n18076, n18077, n18078, n18079, n18080, n18081,
    n18082, n18083, n18084, n18085, n18086, n18087,
    n18088, n18089, n18090, n18091, n18092, n18093,
    n18094, n18095, n18096, n18097, n18098, n18099,
    n18100, n18101, n18102, n18103, n18104, n18105,
    n18106, n18107, n18108, n18109, n18110, n18111,
    n18112, n18113, n18114, n18115, n18116, n18117,
    n18118, n18119, n18120, n18121, n18122, n18123,
    n18124, n18125, n18126, n18127, n18128, n18129,
    n18130, n18131, n18132, n18133, n18134, n18135,
    n18136, n18137, n18138, n18139, n18140, n18141,
    n18142, n18143, n18144, n18145, n18146, n18147,
    n18148, n18149, n18150, n18151, n18152, n18153,
    n18154, n18155, n18156, n18157, n18158, n18159,
    n18160, n18161, n18162, n18163, n18164, n18165,
    n18166, n18167, n18168, n18169, n18170, n18171,
    n18172, n18173, n18174, n18175, n18176, n18177,
    n18178, n18179, n18180, n18181, n18182, n18183,
    n18184, n18185, n18186, n18187, n18188, n18189,
    n18190, n18191, n18192, n18193, n18194, n18195,
    n18196, n18197, n18198, n18199, n18200, n18201,
    n18202, n18203, n18204, n18205, n18206, n18207,
    n18208, n18209, n18210, n18211, n18212, n18213,
    n18214, n18215, n18216, n18217, n18218, n18219,
    n18220, n18221, n18222, n18223, n18224, n18225,
    n18226, n18227, n18228, n18229, n18230, n18231,
    n18232, n18233, n18234, n18235, n18236, n18237,
    n18238, n18239, n18240, n18241, n18242, n18243,
    n18244, n18245, n18246, n18247, n18248, n18249,
    n18250, n18251, n18252, n18253, n18254, n18255,
    n18256, n18257, n18258, n18259, n18260, n18261,
    n18262, n18264, n18265, n18266, n18267, n18268,
    n18269, n18270, n18271, n18272, n18273, n18274,
    n18275, n18276, n18277, n18278, n18279, n18280,
    n18281, n18282, n18283, n18284, n18285, n18286,
    n18287, n18288, n18289, n18290, n18291, n18292,
    n18293, n18294, n18295, n18296, n18297, n18298,
    n18299, n18300, n18301, n18302, n18303, n18304,
    n18305, n18306, n18307, n18308, n18309, n18310,
    n18311, n18312, n18313, n18314, n18315, n18316,
    n18317, n18318, n18319, n18320, n18321, n18322,
    n18323, n18324, n18325, n18326, n18327, n18328,
    n18329, n18330, n18331, n18332, n18333, n18334,
    n18335, n18336, n18337, n18338, n18339, n18340,
    n18341, n18342, n18343, n18344, n18345, n18346,
    n18347, n18348, n18349, n18350, n18351, n18352,
    n18353, n18354, n18355, n18356, n18357, n18358,
    n18359, n18360, n18361, n18362, n18363, n18364,
    n18365, n18366, n18367, n18368, n18369, n18370,
    n18371, n18372, n18373, n18374, n18375, n18376,
    n18377, n18378, n18379, n18380, n18381, n18382,
    n18383, n18384, n18385, n18386, n18387, n18388,
    n18389, n18390, n18391, n18392, n18393, n18394,
    n18395, n18396, n18397, n18398, n18399, n18400,
    n18401, n18402, n18403, n18404, n18405, n18406,
    n18407, n18408, n18409, n18410, n18411, n18412,
    n18413, n18414, n18415, n18416, n18417, n18418,
    n18419, n18420, n18421, n18422, n18423, n18424,
    n18425, n18426, n18427, n18428, n18429, n18430,
    n18431, n18432, n18433, n18434, n18435, n18436,
    n18437, n18438, n18439, n18440, n18441, n18442,
    n18443, n18444, n18445, n18446, n18447, n18448,
    n18449, n18450, n18451, n18452, n18453, n18454,
    n18455, n18456, n18457, n18458, n18459, n18460,
    n18461, n18462, n18463, n18464, n18465, n18466,
    n18467, n18468, n18469, n18470, n18471, n18472,
    n18473, n18474, n18475, n18476, n18477, n18478,
    n18479, n18480, n18481, n18482, n18483, n18484,
    n18485, n18486, n18487, n18488, n18489, n18490,
    n18491, n18492, n18493, n18494, n18495, n18496,
    n18497, n18498, n18499, n18500, n18501, n18502,
    n18503, n18504, n18505, n18506, n18507, n18508,
    n18509, n18510, n18511, n18512, n18513, n18514,
    n18515, n18516, n18517, n18518, n18519, n18520,
    n18521, n18522, n18523, n18524, n18525, n18526,
    n18527, n18528, n18529, n18530, n18531, n18532,
    n18533, n18534, n18535, n18536, n18537, n18538,
    n18539, n18540, n18541, n18542, n18543, n18544,
    n18545, n18546, n18547, n18548, n18549, n18550,
    n18551, n18552, n18553, n18554, n18555, n18556,
    n18557, n18558, n18559, n18560, n18561, n18562,
    n18563, n18564, n18565, n18566, n18567, n18568,
    n18569, n18570, n18571, n18572, n18573, n18574,
    n18575, n18576, n18577, n18578, n18579, n18580,
    n18581, n18582, n18583, n18584, n18585, n18586,
    n18587, n18588, n18589, n18590, n18591, n18592,
    n18593, n18594, n18595, n18596, n18597, n18598,
    n18599, n18600, n18601, n18602, n18603, n18605,
    n18606, n18607, n18608, n18609, n18610, n18611,
    n18612, n18613, n18614, n18615, n18616, n18617,
    n18618, n18619, n18620, n18621, n18622, n18623,
    n18624, n18625, n18626, n18627, n18628, n18629,
    n18630, n18631, n18632, n18633, n18634, n18635,
    n18636, n18637, n18638, n18639, n18640, n18641,
    n18642, n18643, n18644, n18645, n18646, n18647,
    n18648, n18649, n18650, n18651, n18652, n18653,
    n18654, n18655, n18656, n18657, n18658, n18659,
    n18660, n18661, n18662, n18663, n18664, n18665,
    n18666, n18667, n18668, n18669, n18670, n18671,
    n18672, n18673, n18674, n18675, n18676, n18677,
    n18678, n18679, n18680, n18681, n18682, n18683,
    n18684, n18685, n18686, n18687, n18688, n18689,
    n18690, n18691, n18692, n18693, n18694, n18695,
    n18696, n18697, n18698, n18699, n18700, n18701,
    n18702, n18703, n18704, n18705, n18706, n18707,
    n18708, n18709, n18710, n18711, n18712, n18713,
    n18714, n18715, n18716, n18717, n18718, n18719,
    n18720, n18721, n18722, n18723, n18724, n18725,
    n18726, n18727, n18728, n18729, n18730, n18731,
    n18732, n18733, n18734, n18735, n18736, n18737,
    n18738, n18739, n18740, n18741, n18742, n18743,
    n18744, n18745, n18746, n18747, n18748, n18749,
    n18750, n18751, n18752, n18753, n18754, n18755,
    n18756, n18757, n18758, n18759, n18760, n18761,
    n18762, n18763, n18764, n18765, n18766, n18767,
    n18768, n18769, n18770, n18771, n18772, n18773,
    n18774, n18775, n18776, n18777, n18778, n18779,
    n18780, n18781, n18782, n18783, n18784, n18785,
    n18786, n18787, n18788, n18789, n18790, n18791,
    n18792, n18793, n18794, n18795, n18796, n18797,
    n18798, n18799, n18800, n18801, n18802, n18803,
    n18804, n18805, n18806, n18807, n18808, n18809,
    n18810, n18811, n18812, n18813, n18814, n18815,
    n18816, n18817, n18818, n18819, n18820, n18821,
    n18822, n18823, n18824, n18825, n18826, n18827,
    n18828, n18829, n18830, n18831, n18832, n18833,
    n18834, n18835, n18836, n18837, n18838, n18839,
    n18840, n18841, n18842, n18843, n18844, n18845,
    n18846, n18847, n18848, n18849, n18850, n18851,
    n18852, n18853, n18854, n18855, n18856, n18857,
    n18858, n18859, n18860, n18861, n18862, n18863,
    n18864, n18865, n18866, n18867, n18868, n18869,
    n18870, n18871, n18872, n18873, n18874, n18875,
    n18876, n18877, n18878, n18879, n18880, n18881,
    n18882, n18883, n18884, n18885, n18886, n18887,
    n18888, n18889, n18890, n18891, n18892, n18893,
    n18894, n18895, n18896, n18897, n18898, n18899,
    n18900, n18901, n18902, n18903, n18904, n18905,
    n18906, n18907, n18908, n18909, n18910, n18911,
    n18912, n18913, n18914, n18915, n18916, n18917,
    n18918, n18919, n18920, n18921, n18922, n18923,
    n18924, n18925, n18926, n18927, n18929, n18930,
    n18931, n18932, n18933, n18934, n18935, n18936,
    n18937, n18938, n18939, n18940, n18941, n18942,
    n18943, n18944, n18945, n18946, n18947, n18948,
    n18949, n18950, n18951, n18952, n18953, n18954,
    n18955, n18956, n18957, n18958, n18959, n18960,
    n18961, n18962, n18963, n18964, n18965, n18966,
    n18967, n18968, n18969, n18970, n18971, n18972,
    n18973, n18974, n18975, n18976, n18977, n18978,
    n18979, n18980, n18981, n18982, n18983, n18984,
    n18985, n18986, n18987, n18988, n18989, n18990,
    n18991, n18992, n18993, n18994, n18995, n18996,
    n18997, n18998, n18999, n19000, n19001, n19002,
    n19003, n19004, n19005, n19006, n19007, n19008,
    n19009, n19010, n19011, n19012, n19013, n19014,
    n19015, n19016, n19017, n19018, n19019, n19020,
    n19021, n19022, n19023, n19024, n19025, n19026,
    n19027, n19028, n19029, n19030, n19031, n19032,
    n19033, n19034, n19035, n19036, n19037, n19038,
    n19039, n19040, n19041, n19042, n19043, n19044,
    n19045, n19046, n19047, n19048, n19049, n19050,
    n19051, n19052, n19053, n19054, n19055, n19056,
    n19057, n19058, n19059, n19060, n19061, n19062,
    n19063, n19064, n19065, n19066, n19067, n19068,
    n19069, n19070, n19071, n19072, n19073, n19074,
    n19075, n19076, n19077, n19078, n19079, n19080,
    n19081, n19082, n19083, n19084, n19085, n19086,
    n19087, n19088, n19089, n19090, n19091, n19092,
    n19093, n19094, n19095, n19096, n19097, n19098,
    n19099, n19100, n19101, n19102, n19103, n19104,
    n19105, n19106, n19107, n19108, n19109, n19110,
    n19111, n19112, n19113, n19114, n19115, n19116,
    n19117, n19118, n19119, n19120, n19121, n19122,
    n19123, n19124, n19125, n19126, n19127, n19128,
    n19129, n19130, n19131, n19132, n19133, n19134,
    n19135, n19136, n19137, n19138, n19139, n19140,
    n19141, n19142, n19143, n19144, n19145, n19146,
    n19147, n19148, n19149, n19150, n19151, n19152,
    n19153, n19154, n19155, n19156, n19157, n19158,
    n19159, n19160, n19161, n19162, n19163, n19164,
    n19165, n19166, n19167, n19168, n19169, n19170,
    n19171, n19172, n19173, n19174, n19175, n19176,
    n19177, n19178, n19179, n19180, n19181, n19182,
    n19183, n19184, n19185, n19186, n19187, n19188,
    n19189, n19190, n19191, n19192, n19193, n19194,
    n19195, n19196, n19197, n19198, n19199, n19200,
    n19201, n19202, n19203, n19204, n19205, n19206,
    n19207, n19208, n19209, n19210, n19211, n19212,
    n19213, n19214, n19215, n19216, n19217, n19218,
    n19219, n19220, n19221, n19222, n19223, n19224,
    n19225, n19226, n19227, n19228, n19229, n19230,
    n19231, n19232, n19233, n19234, n19235, n19236,
    n19237, n19238, n19239, n19240, n19241, n19242,
    n19243, n19244, n19245, n19246, n19247, n19248,
    n19249, n19251, n19252, n19253, n19254, n19255,
    n19256, n19257, n19258, n19259, n19260, n19261,
    n19262, n19263, n19264, n19265, n19266, n19267,
    n19268, n19269, n19270, n19271, n19272, n19273,
    n19274, n19275, n19276, n19277, n19278, n19279,
    n19280, n19281, n19282, n19283, n19284, n19285,
    n19286, n19287, n19288, n19289, n19290, n19291,
    n19292, n19293, n19294, n19295, n19296, n19297,
    n19298, n19299, n19300, n19301, n19302, n19303,
    n19304, n19305, n19306, n19307, n19308, n19309,
    n19310, n19311, n19312, n19313, n19314, n19315,
    n19316, n19317, n19318, n19319, n19320, n19321,
    n19322, n19323, n19324, n19325, n19326, n19327,
    n19328, n19329, n19330, n19331, n19332, n19333,
    n19334, n19335, n19336, n19337, n19338, n19339,
    n19340, n19341, n19342, n19343, n19344, n19345,
    n19346, n19347, n19348, n19349, n19350, n19351,
    n19352, n19353, n19354, n19355, n19356, n19357,
    n19358, n19359, n19360, n19361, n19362, n19363,
    n19364, n19365, n19366, n19367, n19368, n19369,
    n19370, n19371, n19372, n19373, n19374, n19375,
    n19376, n19377, n19378, n19379, n19380, n19381,
    n19382, n19383, n19384, n19385, n19386, n19387,
    n19388, n19389, n19390, n19391, n19392, n19393,
    n19394, n19395, n19396, n19397, n19398, n19399,
    n19400, n19401, n19402, n19403, n19404, n19405,
    n19406, n19407, n19408, n19409, n19410, n19411,
    n19412, n19413, n19414, n19415, n19416, n19417,
    n19418, n19419, n19420, n19421, n19422, n19423,
    n19424, n19425, n19426, n19427, n19428, n19429,
    n19430, n19431, n19432, n19433, n19434, n19435,
    n19436, n19437, n19438, n19439, n19440, n19441,
    n19442, n19443, n19444, n19445, n19446, n19447,
    n19448, n19449, n19450, n19451, n19452, n19453,
    n19454, n19455, n19456, n19457, n19458, n19459,
    n19460, n19461, n19462, n19463, n19464, n19465,
    n19466, n19467, n19468, n19469, n19470, n19471,
    n19472, n19473, n19474, n19475, n19476, n19477,
    n19478, n19479, n19480, n19481, n19482, n19483,
    n19484, n19485, n19486, n19487, n19488, n19489,
    n19490, n19491, n19492, n19493, n19494, n19495,
    n19496, n19497, n19498, n19499, n19500, n19501,
    n19502, n19503, n19504, n19505, n19506, n19507,
    n19508, n19509, n19510, n19511, n19512, n19513,
    n19514, n19515, n19516, n19517, n19518, n19519,
    n19520, n19521, n19522, n19523, n19524, n19525,
    n19526, n19527, n19528, n19529, n19530, n19531,
    n19532, n19533, n19534, n19535, n19536, n19537,
    n19538, n19539, n19540, n19541, n19542, n19543,
    n19544, n19545, n19546, n19547, n19548, n19549,
    n19550, n19551, n19552, n19553, n19554, n19555,
    n19556, n19557, n19558, n19559, n19561, n19562,
    n19563, n19564, n19565, n19566, n19567, n19568,
    n19569, n19570, n19571, n19572, n19573, n19574,
    n19575, n19576, n19577, n19578, n19579, n19580,
    n19581, n19582, n19583, n19584, n19585, n19586,
    n19587, n19588, n19589, n19590, n19591, n19592,
    n19593, n19594, n19595, n19596, n19597, n19598,
    n19599, n19600, n19601, n19602, n19603, n19604,
    n19605, n19606, n19607, n19608, n19609, n19610,
    n19611, n19612, n19613, n19614, n19615, n19616,
    n19617, n19618, n19619, n19620, n19621, n19622,
    n19623, n19624, n19625, n19626, n19627, n19628,
    n19629, n19630, n19631, n19632, n19633, n19634,
    n19635, n19636, n19637, n19638, n19639, n19640,
    n19641, n19642, n19643, n19644, n19645, n19646,
    n19647, n19648, n19649, n19650, n19651, n19652,
    n19653, n19654, n19655, n19656, n19657, n19658,
    n19659, n19660, n19661, n19662, n19663, n19664,
    n19665, n19666, n19667, n19668, n19669, n19670,
    n19671, n19672, n19673, n19674, n19675, n19676,
    n19677, n19678, n19679, n19680, n19681, n19682,
    n19683, n19684, n19685, n19686, n19687, n19688,
    n19689, n19690, n19691, n19692, n19693, n19694,
    n19695, n19696, n19697, n19698, n19699, n19700,
    n19701, n19702, n19703, n19704, n19705, n19706,
    n19707, n19708, n19709, n19710, n19711, n19712,
    n19713, n19714, n19715, n19716, n19717, n19718,
    n19719, n19720, n19721, n19722, n19723, n19724,
    n19725, n19726, n19727, n19728, n19729, n19730,
    n19731, n19732, n19733, n19734, n19735, n19736,
    n19737, n19738, n19739, n19740, n19741, n19742,
    n19743, n19744, n19745, n19746, n19747, n19748,
    n19749, n19750, n19751, n19752, n19753, n19754,
    n19755, n19756, n19757, n19758, n19759, n19760,
    n19761, n19762, n19763, n19764, n19765, n19766,
    n19767, n19768, n19769, n19770, n19771, n19772,
    n19773, n19774, n19775, n19776, n19777, n19778,
    n19779, n19780, n19781, n19782, n19783, n19784,
    n19785, n19786, n19787, n19788, n19789, n19790,
    n19791, n19792, n19793, n19794, n19795, n19796,
    n19797, n19798, n19799, n19800, n19801, n19802,
    n19803, n19804, n19805, n19806, n19807, n19808,
    n19809, n19810, n19811, n19812, n19813, n19814,
    n19815, n19816, n19817, n19818, n19819, n19820,
    n19821, n19822, n19823, n19824, n19825, n19826,
    n19827, n19828, n19829, n19830, n19831, n19832,
    n19833, n19834, n19835, n19836, n19837, n19838,
    n19839, n19840, n19841, n19842, n19843, n19844,
    n19845, n19846, n19847, n19848, n19849, n19850,
    n19851, n19852, n19853, n19854, n19855, n19856,
    n19857, n19858, n19859, n19860, n19861, n19862,
    n19863, n19864, n19865, n19866, n19867, n19869,
    n19870, n19871, n19872, n19873, n19874, n19875,
    n19876, n19877, n19878, n19879, n19880, n19881,
    n19882, n19883, n19884, n19885, n19886, n19887,
    n19888, n19889, n19890, n19891, n19892, n19893,
    n19894, n19895, n19896, n19897, n19898, n19899,
    n19900, n19901, n19902, n19903, n19904, n19905,
    n19906, n19907, n19908, n19909, n19910, n19911,
    n19912, n19913, n19914, n19915, n19916, n19917,
    n19918, n19919, n19920, n19921, n19922, n19923,
    n19924, n19925, n19926, n19927, n19928, n19929,
    n19930, n19931, n19932, n19933, n19934, n19935,
    n19936, n19937, n19938, n19939, n19940, n19941,
    n19942, n19943, n19944, n19945, n19946, n19947,
    n19948, n19949, n19950, n19951, n19952, n19953,
    n19954, n19955, n19956, n19957, n19958, n19959,
    n19960, n19961, n19962, n19963, n19964, n19965,
    n19966, n19967, n19968, n19969, n19970, n19971,
    n19972, n19973, n19974, n19975, n19976, n19977,
    n19978, n19979, n19980, n19981, n19982, n19983,
    n19984, n19985, n19986, n19987, n19988, n19989,
    n19990, n19991, n19992, n19993, n19994, n19995,
    n19996, n19997, n19998, n19999, n20000, n20001,
    n20002, n20003, n20004, n20005, n20006, n20007,
    n20008, n20009, n20010, n20011, n20012, n20013,
    n20014, n20015, n20016, n20017, n20018, n20019,
    n20020, n20021, n20022, n20023, n20024, n20025,
    n20026, n20027, n20028, n20029, n20030, n20031,
    n20032, n20033, n20034, n20035, n20036, n20037,
    n20038, n20039, n20040, n20041, n20042, n20043,
    n20044, n20045, n20046, n20047, n20048, n20049,
    n20050, n20051, n20052, n20053, n20054, n20055,
    n20056, n20057, n20058, n20059, n20060, n20061,
    n20062, n20063, n20064, n20065, n20066, n20067,
    n20068, n20069, n20070, n20071, n20072, n20073,
    n20074, n20075, n20076, n20077, n20078, n20079,
    n20080, n20081, n20082, n20083, n20084, n20085,
    n20086, n20087, n20088, n20089, n20090, n20091,
    n20092, n20093, n20094, n20095, n20096, n20097,
    n20098, n20099, n20100, n20101, n20102, n20103,
    n20104, n20105, n20106, n20107, n20108, n20109,
    n20110, n20111, n20112, n20113, n20114, n20115,
    n20116, n20117, n20118, n20119, n20120, n20121,
    n20122, n20123, n20124, n20125, n20126, n20127,
    n20128, n20129, n20130, n20131, n20132, n20133,
    n20134, n20135, n20136, n20137, n20138, n20139,
    n20140, n20141, n20142, n20143, n20144, n20145,
    n20146, n20147, n20148, n20149, n20150, n20151,
    n20152, n20153, n20154, n20155, n20156, n20157,
    n20158, n20159, n20160, n20161, n20162, n20163,
    n20164, n20165, n20166, n20167, n20168, n20170,
    n20171, n20172, n20173, n20174, n20175, n20176,
    n20177, n20178, n20179, n20180, n20181, n20182,
    n20183, n20184, n20185, n20186, n20187, n20188,
    n20189, n20190, n20191, n20192, n20193, n20194,
    n20195, n20196, n20197, n20198, n20199, n20200,
    n20201, n20202, n20203, n20204, n20205, n20206,
    n20207, n20208, n20209, n20210, n20211, n20212,
    n20213, n20214, n20215, n20216, n20217, n20218,
    n20219, n20220, n20221, n20222, n20223, n20224,
    n20225, n20226, n20227, n20228, n20229, n20230,
    n20231, n20232, n20233, n20234, n20235, n20236,
    n20237, n20238, n20239, n20240, n20241, n20242,
    n20243, n20244, n20245, n20246, n20247, n20248,
    n20249, n20250, n20251, n20252, n20253, n20254,
    n20255, n20256, n20257, n20258, n20259, n20260,
    n20261, n20262, n20263, n20264, n20265, n20266,
    n20267, n20268, n20269, n20270, n20271, n20272,
    n20273, n20274, n20275, n20276, n20277, n20278,
    n20279, n20280, n20281, n20282, n20283, n20284,
    n20285, n20286, n20287, n20288, n20289, n20290,
    n20291, n20292, n20293, n20294, n20295, n20296,
    n20297, n20298, n20299, n20300, n20301, n20302,
    n20303, n20304, n20305, n20306, n20307, n20308,
    n20309, n20310, n20311, n20312, n20313, n20314,
    n20315, n20316, n20317, n20318, n20319, n20320,
    n20321, n20322, n20323, n20324, n20325, n20326,
    n20327, n20328, n20329, n20330, n20331, n20332,
    n20333, n20334, n20335, n20336, n20337, n20338,
    n20339, n20340, n20341, n20342, n20343, n20344,
    n20345, n20346, n20347, n20348, n20349, n20350,
    n20351, n20352, n20353, n20354, n20355, n20356,
    n20357, n20358, n20359, n20360, n20361, n20362,
    n20363, n20364, n20365, n20366, n20367, n20368,
    n20369, n20370, n20371, n20372, n20373, n20374,
    n20375, n20376, n20377, n20378, n20379, n20380,
    n20381, n20382, n20383, n20384, n20385, n20386,
    n20387, n20388, n20389, n20390, n20391, n20392,
    n20393, n20394, n20395, n20396, n20397, n20398,
    n20399, n20400, n20401, n20402, n20403, n20404,
    n20405, n20406, n20407, n20408, n20409, n20410,
    n20411, n20412, n20413, n20414, n20415, n20416,
    n20417, n20418, n20419, n20420, n20421, n20422,
    n20423, n20424, n20425, n20426, n20427, n20428,
    n20429, n20430, n20431, n20432, n20433, n20434,
    n20435, n20436, n20437, n20438, n20439, n20440,
    n20441, n20442, n20443, n20444, n20445, n20446,
    n20447, n20448, n20449, n20450, n20451, n20452,
    n20453, n20454, n20455, n20456, n20457, n20458,
    n20459, n20460, n20462, n20463, n20464, n20465,
    n20466, n20467, n20468, n20469, n20470, n20471,
    n20472, n20473, n20474, n20475, n20476, n20477,
    n20478, n20479, n20480, n20481, n20482, n20483,
    n20484, n20485, n20486, n20487, n20488, n20489,
    n20490, n20491, n20492, n20493, n20494, n20495,
    n20496, n20497, n20498, n20499, n20500, n20501,
    n20502, n20503, n20504, n20505, n20506, n20507,
    n20508, n20509, n20510, n20511, n20512, n20513,
    n20514, n20515, n20516, n20517, n20518, n20519,
    n20520, n20521, n20522, n20523, n20524, n20525,
    n20526, n20527, n20528, n20529, n20530, n20531,
    n20532, n20533, n20534, n20535, n20536, n20537,
    n20538, n20539, n20540, n20541, n20542, n20543,
    n20544, n20545, n20546, n20547, n20548, n20549,
    n20550, n20551, n20552, n20553, n20554, n20555,
    n20556, n20557, n20558, n20559, n20560, n20561,
    n20562, n20563, n20564, n20565, n20566, n20567,
    n20568, n20569, n20570, n20571, n20572, n20573,
    n20574, n20575, n20576, n20577, n20578, n20579,
    n20580, n20581, n20582, n20583, n20584, n20585,
    n20586, n20587, n20588, n20589, n20590, n20591,
    n20592, n20593, n20594, n20595, n20596, n20597,
    n20598, n20599, n20600, n20601, n20602, n20603,
    n20604, n20605, n20606, n20607, n20608, n20609,
    n20610, n20611, n20612, n20613, n20614, n20615,
    n20616, n20617, n20618, n20619, n20620, n20621,
    n20622, n20623, n20624, n20625, n20626, n20627,
    n20628, n20629, n20630, n20631, n20632, n20633,
    n20634, n20635, n20636, n20637, n20638, n20639,
    n20640, n20641, n20642, n20643, n20644, n20645,
    n20646, n20647, n20648, n20649, n20650, n20651,
    n20652, n20653, n20654, n20655, n20656, n20657,
    n20658, n20659, n20660, n20661, n20662, n20663,
    n20664, n20665, n20666, n20667, n20668, n20669,
    n20670, n20671, n20672, n20673, n20674, n20675,
    n20676, n20677, n20678, n20679, n20680, n20681,
    n20682, n20683, n20684, n20685, n20686, n20687,
    n20688, n20689, n20690, n20691, n20692, n20693,
    n20694, n20695, n20696, n20697, n20698, n20699,
    n20700, n20701, n20702, n20703, n20704, n20705,
    n20706, n20707, n20708, n20709, n20710, n20711,
    n20712, n20713, n20714, n20715, n20716, n20717,
    n20718, n20719, n20720, n20721, n20722, n20723,
    n20724, n20725, n20726, n20727, n20728, n20729,
    n20730, n20731, n20732, n20733, n20734, n20735,
    n20736, n20737, n20738, n20739, n20740, n20741,
    n20742, n20743, n20744, n20745, n20747, n20748,
    n20749, n20750, n20751, n20752, n20753, n20754,
    n20755, n20756, n20757, n20758, n20759, n20760,
    n20761, n20762, n20763, n20764, n20765, n20766,
    n20767, n20768, n20769, n20770, n20771, n20772,
    n20773, n20774, n20775, n20776, n20777, n20778,
    n20779, n20780, n20781, n20782, n20783, n20784,
    n20785, n20786, n20787, n20788, n20789, n20790,
    n20791, n20792, n20793, n20794, n20795, n20796,
    n20797, n20798, n20799, n20800, n20801, n20802,
    n20803, n20804, n20805, n20806, n20807, n20808,
    n20809, n20810, n20811, n20812, n20813, n20814,
    n20815, n20816, n20817, n20818, n20819, n20820,
    n20821, n20822, n20823, n20824, n20825, n20826,
    n20827, n20828, n20829, n20830, n20831, n20832,
    n20833, n20834, n20835, n20836, n20837, n20838,
    n20839, n20840, n20841, n20842, n20843, n20844,
    n20845, n20846, n20847, n20848, n20849, n20850,
    n20851, n20852, n20853, n20854, n20855, n20856,
    n20857, n20858, n20859, n20860, n20861, n20862,
    n20863, n20864, n20865, n20866, n20867, n20868,
    n20869, n20870, n20871, n20872, n20873, n20874,
    n20875, n20876, n20877, n20878, n20879, n20880,
    n20881, n20882, n20883, n20884, n20885, n20886,
    n20887, n20888, n20889, n20890, n20891, n20892,
    n20893, n20894, n20895, n20896, n20897, n20898,
    n20899, n20900, n20901, n20902, n20903, n20904,
    n20905, n20906, n20907, n20908, n20909, n20910,
    n20911, n20912, n20913, n20914, n20915, n20916,
    n20917, n20918, n20919, n20920, n20921, n20922,
    n20923, n20924, n20925, n20926, n20927, n20928,
    n20929, n20930, n20931, n20932, n20933, n20934,
    n20935, n20936, n20937, n20938, n20939, n20940,
    n20941, n20942, n20943, n20944, n20945, n20946,
    n20947, n20948, n20949, n20950, n20951, n20952,
    n20953, n20954, n20955, n20956, n20957, n20958,
    n20959, n20960, n20961, n20962, n20963, n20964,
    n20965, n20966, n20967, n20968, n20969, n20970,
    n20971, n20972, n20973, n20974, n20975, n20976,
    n20977, n20978, n20979, n20980, n20981, n20982,
    n20983, n20984, n20985, n20986, n20987, n20988,
    n20989, n20990, n20991, n20992, n20993, n20994,
    n20995, n20996, n20997, n20998, n20999, n21000,
    n21001, n21002, n21003, n21004, n21005, n21006,
    n21007, n21008, n21009, n21010, n21011, n21012,
    n21013, n21014, n21015, n21016, n21017, n21018,
    n21019, n21020, n21021, n21022, n21023, n21024,
    n21025, n21026, n21027, n21028, n21029, n21030,
    n21032, n21033, n21034, n21035, n21036, n21037,
    n21038, n21039, n21040, n21041, n21042, n21043,
    n21044, n21045, n21046, n21047, n21048, n21049,
    n21050, n21051, n21052, n21053, n21054, n21055,
    n21056, n21057, n21058, n21059, n21060, n21061,
    n21062, n21063, n21064, n21065, n21066, n21067,
    n21068, n21069, n21070, n21071, n21072, n21073,
    n21074, n21075, n21076, n21077, n21078, n21079,
    n21080, n21081, n21082, n21083, n21084, n21085,
    n21086, n21087, n21088, n21089, n21090, n21091,
    n21092, n21093, n21094, n21095, n21096, n21097,
    n21098, n21099, n21100, n21101, n21102, n21103,
    n21104, n21105, n21106, n21107, n21108, n21109,
    n21110, n21111, n21112, n21113, n21114, n21115,
    n21116, n21117, n21118, n21119, n21120, n21121,
    n21122, n21123, n21124, n21125, n21126, n21127,
    n21128, n21129, n21130, n21131, n21132, n21133,
    n21134, n21135, n21136, n21137, n21138, n21139,
    n21140, n21141, n21142, n21143, n21144, n21145,
    n21146, n21147, n21148, n21149, n21150, n21151,
    n21152, n21153, n21154, n21155, n21156, n21157,
    n21158, n21159, n21160, n21161, n21162, n21163,
    n21164, n21165, n21166, n21167, n21168, n21169,
    n21170, n21171, n21172, n21173, n21174, n21175,
    n21176, n21177, n21178, n21179, n21180, n21181,
    n21182, n21183, n21184, n21185, n21186, n21187,
    n21188, n21189, n21190, n21191, n21192, n21193,
    n21194, n21195, n21196, n21197, n21198, n21199,
    n21200, n21201, n21202, n21203, n21204, n21205,
    n21206, n21207, n21208, n21209, n21210, n21211,
    n21212, n21213, n21214, n21215, n21216, n21217,
    n21218, n21219, n21220, n21221, n21222, n21223,
    n21224, n21225, n21226, n21227, n21228, n21229,
    n21230, n21231, n21232, n21233, n21234, n21235,
    n21236, n21237, n21238, n21239, n21240, n21241,
    n21242, n21243, n21244, n21245, n21246, n21247,
    n21248, n21249, n21250, n21251, n21252, n21253,
    n21254, n21255, n21256, n21257, n21258, n21259,
    n21260, n21261, n21262, n21263, n21264, n21265,
    n21266, n21267, n21268, n21269, n21270, n21271,
    n21272, n21273, n21274, n21275, n21276, n21277,
    n21278, n21279, n21280, n21281, n21282, n21283,
    n21284, n21285, n21286, n21287, n21288, n21289,
    n21290, n21291, n21292, n21293, n21294, n21295,
    n21296, n21297, n21298, n21299, n21300, n21302,
    n21303, n21304, n21305, n21306, n21307, n21308,
    n21309, n21310, n21311, n21312, n21313, n21314,
    n21315, n21316, n21317, n21318, n21319, n21320,
    n21321, n21322, n21323, n21324, n21325, n21326,
    n21327, n21328, n21329, n21330, n21331, n21332,
    n21333, n21334, n21335, n21336, n21337, n21338,
    n21339, n21340, n21341, n21342, n21343, n21344,
    n21345, n21346, n21347, n21348, n21349, n21350,
    n21351, n21352, n21353, n21354, n21355, n21356,
    n21357, n21358, n21359, n21360, n21361, n21362,
    n21363, n21364, n21365, n21366, n21367, n21368,
    n21369, n21370, n21371, n21372, n21373, n21374,
    n21375, n21376, n21377, n21378, n21379, n21380,
    n21381, n21382, n21383, n21384, n21385, n21386,
    n21387, n21388, n21389, n21390, n21391, n21392,
    n21393, n21394, n21395, n21396, n21397, n21398,
    n21399, n21400, n21401, n21402, n21403, n21404,
    n21405, n21406, n21407, n21408, n21409, n21410,
    n21411, n21412, n21413, n21414, n21415, n21416,
    n21417, n21418, n21419, n21420, n21421, n21422,
    n21423, n21424, n21425, n21426, n21427, n21428,
    n21429, n21430, n21431, n21432, n21433, n21434,
    n21435, n21436, n21437, n21438, n21439, n21440,
    n21441, n21442, n21443, n21444, n21445, n21446,
    n21447, n21448, n21449, n21450, n21451, n21452,
    n21453, n21454, n21455, n21456, n21457, n21458,
    n21459, n21460, n21461, n21462, n21463, n21464,
    n21465, n21466, n21467, n21468, n21469, n21470,
    n21471, n21472, n21473, n21474, n21475, n21476,
    n21477, n21478, n21479, n21480, n21481, n21482,
    n21483, n21484, n21485, n21486, n21487, n21488,
    n21489, n21490, n21491, n21492, n21493, n21494,
    n21495, n21496, n21497, n21498, n21499, n21500,
    n21501, n21502, n21503, n21504, n21505, n21506,
    n21507, n21508, n21509, n21510, n21511, n21512,
    n21513, n21514, n21515, n21516, n21517, n21518,
    n21519, n21520, n21521, n21522, n21523, n21524,
    n21525, n21526, n21527, n21528, n21529, n21530,
    n21531, n21532, n21533, n21534, n21535, n21536,
    n21537, n21538, n21539, n21540, n21541, n21542,
    n21543, n21544, n21545, n21546, n21547, n21548,
    n21549, n21550, n21551, n21552, n21553, n21554,
    n21555, n21556, n21557, n21558, n21559, n21560,
    n21561, n21562, n21563, n21564, n21565, n21566,
    n21567, n21568, n21569, n21570, n21572, n21573,
    n21574, n21575, n21576, n21577, n21578, n21579,
    n21580, n21581, n21582, n21583, n21584, n21585,
    n21586, n21587, n21588, n21589, n21590, n21591,
    n21592, n21593, n21594, n21595, n21596, n21597,
    n21598, n21599, n21600, n21601, n21602, n21603,
    n21604, n21605, n21606, n21607, n21608, n21609,
    n21610, n21611, n21612, n21613, n21614, n21615,
    n21616, n21617, n21618, n21619, n21620, n21621,
    n21622, n21623, n21624, n21625, n21626, n21627,
    n21628, n21629, n21630, n21631, n21632, n21633,
    n21634, n21635, n21636, n21637, n21638, n21639,
    n21640, n21641, n21642, n21643, n21644, n21645,
    n21646, n21647, n21648, n21649, n21650, n21651,
    n21652, n21653, n21654, n21655, n21656, n21657,
    n21658, n21659, n21660, n21661, n21662, n21663,
    n21664, n21665, n21666, n21667, n21668, n21669,
    n21670, n21671, n21672, n21673, n21674, n21675,
    n21676, n21677, n21678, n21679, n21680, n21681,
    n21682, n21683, n21684, n21685, n21686, n21687,
    n21688, n21689, n21690, n21691, n21692, n21693,
    n21694, n21695, n21696, n21697, n21698, n21699,
    n21700, n21701, n21702, n21703, n21704, n21705,
    n21706, n21707, n21708, n21709, n21710, n21711,
    n21712, n21713, n21714, n21715, n21716, n21717,
    n21718, n21719, n21720, n21721, n21722, n21723,
    n21724, n21725, n21726, n21727, n21728, n21729,
    n21730, n21731, n21732, n21733, n21734, n21735,
    n21736, n21737, n21738, n21739, n21740, n21741,
    n21742, n21743, n21744, n21745, n21746, n21747,
    n21748, n21749, n21750, n21751, n21752, n21753,
    n21754, n21755, n21756, n21757, n21758, n21759,
    n21760, n21761, n21762, n21763, n21764, n21765,
    n21766, n21767, n21768, n21769, n21770, n21771,
    n21772, n21773, n21774, n21775, n21776, n21777,
    n21778, n21779, n21780, n21781, n21782, n21783,
    n21784, n21785, n21786, n21787, n21788, n21789,
    n21790, n21791, n21792, n21793, n21794, n21795,
    n21796, n21797, n21798, n21799, n21800, n21801,
    n21802, n21803, n21804, n21805, n21806, n21807,
    n21808, n21809, n21810, n21811, n21812, n21813,
    n21814, n21815, n21816, n21817, n21818, n21819,
    n21820, n21821, n21822, n21823, n21824, n21825,
    n21826, n21827, n21828, n21829, n21830, n21831,
    n21832, n21833, n21834, n21836, n21837, n21838,
    n21839, n21840, n21841, n21842, n21843, n21844,
    n21845, n21846, n21847, n21848, n21849, n21850,
    n21851, n21852, n21853, n21854, n21855, n21856,
    n21857, n21858, n21859, n21860, n21861, n21862,
    n21863, n21864, n21865, n21866, n21867, n21868,
    n21869, n21870, n21871, n21872, n21873, n21874,
    n21875, n21876, n21877, n21878, n21879, n21880,
    n21881, n21882, n21883, n21884, n21885, n21886,
    n21887, n21888, n21889, n21890, n21891, n21892,
    n21893, n21894, n21895, n21896, n21897, n21898,
    n21899, n21900, n21901, n21902, n21903, n21904,
    n21905, n21906, n21907, n21908, n21909, n21910,
    n21911, n21912, n21913, n21914, n21915, n21916,
    n21917, n21918, n21919, n21920, n21921, n21922,
    n21923, n21924, n21925, n21926, n21927, n21928,
    n21929, n21930, n21931, n21932, n21933, n21934,
    n21935, n21936, n21937, n21938, n21939, n21940,
    n21941, n21942, n21943, n21944, n21945, n21946,
    n21947, n21948, n21949, n21950, n21951, n21952,
    n21953, n21954, n21955, n21956, n21957, n21958,
    n21959, n21960, n21961, n21962, n21963, n21964,
    n21965, n21966, n21967, n21968, n21969, n21970,
    n21971, n21972, n21973, n21974, n21975, n21976,
    n21977, n21978, n21979, n21980, n21981, n21982,
    n21983, n21984, n21985, n21986, n21987, n21988,
    n21989, n21990, n21991, n21992, n21993, n21994,
    n21995, n21996, n21997, n21998, n21999, n22000,
    n22001, n22002, n22003, n22004, n22005, n22006,
    n22007, n22008, n22009, n22010, n22011, n22012,
    n22013, n22014, n22015, n22016, n22017, n22018,
    n22019, n22020, n22021, n22022, n22023, n22024,
    n22025, n22026, n22027, n22028, n22029, n22030,
    n22031, n22032, n22033, n22034, n22035, n22036,
    n22037, n22038, n22039, n22040, n22041, n22042,
    n22043, n22044, n22045, n22046, n22047, n22048,
    n22049, n22050, n22051, n22052, n22053, n22054,
    n22055, n22056, n22057, n22058, n22059, n22060,
    n22061, n22062, n22063, n22064, n22065, n22066,
    n22067, n22068, n22069, n22070, n22071, n22072,
    n22073, n22074, n22075, n22076, n22077, n22078,
    n22079, n22080, n22081, n22082, n22083, n22084,
    n22085, n22086, n22087, n22088, n22089, n22090,
    n22091, n22093, n22094, n22095, n22096, n22097,
    n22098, n22099, n22100, n22101, n22102, n22103,
    n22104, n22105, n22106, n22107, n22108, n22109,
    n22110, n22111, n22112, n22113, n22114, n22115,
    n22116, n22117, n22118, n22119, n22120, n22121,
    n22122, n22123, n22124, n22125, n22126, n22127,
    n22128, n22129, n22130, n22131, n22132, n22133,
    n22134, n22135, n22136, n22137, n22138, n22139,
    n22140, n22141, n22142, n22143, n22144, n22145,
    n22146, n22147, n22148, n22149, n22150, n22151,
    n22152, n22153, n22154, n22155, n22156, n22157,
    n22158, n22159, n22160, n22161, n22162, n22163,
    n22164, n22165, n22166, n22167, n22168, n22169,
    n22170, n22171, n22172, n22173, n22174, n22175,
    n22176, n22177, n22178, n22179, n22180, n22181,
    n22182, n22183, n22184, n22185, n22186, n22187,
    n22188, n22189, n22190, n22191, n22192, n22193,
    n22194, n22195, n22196, n22197, n22198, n22199,
    n22200, n22201, n22202, n22203, n22204, n22205,
    n22206, n22207, n22208, n22209, n22210, n22211,
    n22212, n22213, n22214, n22215, n22216, n22217,
    n22218, n22219, n22220, n22221, n22222, n22223,
    n22224, n22225, n22226, n22227, n22228, n22229,
    n22230, n22231, n22232, n22233, n22234, n22235,
    n22236, n22237, n22238, n22239, n22240, n22241,
    n22242, n22243, n22244, n22245, n22246, n22247,
    n22248, n22249, n22250, n22251, n22252, n22253,
    n22254, n22255, n22256, n22257, n22258, n22259,
    n22260, n22261, n22262, n22263, n22264, n22265,
    n22266, n22267, n22268, n22269, n22270, n22271,
    n22272, n22273, n22274, n22275, n22276, n22277,
    n22278, n22279, n22280, n22281, n22282, n22283,
    n22284, n22285, n22286, n22287, n22288, n22289,
    n22290, n22291, n22292, n22293, n22294, n22295,
    n22296, n22297, n22298, n22299, n22300, n22301,
    n22302, n22303, n22304, n22305, n22306, n22307,
    n22308, n22309, n22310, n22311, n22312, n22313,
    n22314, n22315, n22316, n22317, n22318, n22319,
    n22320, n22321, n22322, n22323, n22324, n22325,
    n22326, n22327, n22328, n22329, n22330, n22331,
    n22332, n22333, n22334, n22335, n22336, n22337,
    n22338, n22339, n22341, n22342, n22343, n22344,
    n22345, n22346, n22347, n22348, n22349, n22350,
    n22351, n22352, n22353, n22354, n22355, n22356,
    n22357, n22358, n22359, n22360, n22361, n22362,
    n22363, n22364, n22365, n22366, n22367, n22368,
    n22369, n22370, n22371, n22372, n22373, n22374,
    n22375, n22376, n22377, n22378, n22379, n22380,
    n22381, n22382, n22383, n22384, n22385, n22386,
    n22387, n22388, n22389, n22390, n22391, n22392,
    n22393, n22394, n22395, n22396, n22397, n22398,
    n22399, n22400, n22401, n22402, n22403, n22404,
    n22405, n22406, n22407, n22408, n22409, n22410,
    n22411, n22412, n22413, n22414, n22415, n22416,
    n22417, n22418, n22419, n22420, n22421, n22422,
    n22423, n22424, n22425, n22426, n22427, n22428,
    n22429, n22430, n22431, n22432, n22433, n22434,
    n22435, n22436, n22437, n22438, n22439, n22440,
    n22441, n22442, n22443, n22444, n22445, n22446,
    n22447, n22448, n22449, n22450, n22451, n22452,
    n22453, n22454, n22455, n22456, n22457, n22458,
    n22459, n22460, n22461, n22462, n22463, n22464,
    n22465, n22466, n22467, n22468, n22469, n22470,
    n22471, n22472, n22473, n22474, n22475, n22476,
    n22477, n22478, n22479, n22480, n22481, n22482,
    n22483, n22484, n22485, n22486, n22487, n22488,
    n22489, n22490, n22491, n22492, n22493, n22494,
    n22495, n22496, n22497, n22498, n22499, n22500,
    n22501, n22502, n22503, n22504, n22505, n22506,
    n22507, n22508, n22509, n22510, n22511, n22512,
    n22513, n22514, n22515, n22516, n22517, n22518,
    n22519, n22520, n22521, n22522, n22523, n22524,
    n22525, n22526, n22527, n22528, n22529, n22530,
    n22531, n22532, n22533, n22534, n22535, n22536,
    n22537, n22538, n22539, n22540, n22541, n22542,
    n22543, n22544, n22545, n22546, n22547, n22548,
    n22549, n22550, n22551, n22552, n22553, n22554,
    n22555, n22556, n22557, n22558, n22559, n22560,
    n22561, n22562, n22563, n22564, n22565, n22566,
    n22567, n22568, n22569, n22570, n22571, n22572,
    n22573, n22574, n22575, n22576, n22577, n22578,
    n22579, n22580, n22581, n22582, n22584, n22585,
    n22586, n22587, n22588, n22589, n22590, n22591,
    n22592, n22593, n22594, n22595, n22596, n22597,
    n22598, n22599, n22600, n22601, n22602, n22603,
    n22604, n22605, n22606, n22607, n22608, n22609,
    n22610, n22611, n22612, n22613, n22614, n22615,
    n22616, n22617, n22618, n22619, n22620, n22621,
    n22622, n22623, n22624, n22625, n22626, n22627,
    n22628, n22629, n22630, n22631, n22632, n22633,
    n22634, n22635, n22636, n22637, n22638, n22639,
    n22640, n22641, n22642, n22643, n22644, n22645,
    n22646, n22647, n22648, n22649, n22650, n22651,
    n22652, n22653, n22654, n22655, n22656, n22657,
    n22658, n22659, n22660, n22661, n22662, n22663,
    n22664, n22665, n22666, n22667, n22668, n22669,
    n22670, n22671, n22672, n22673, n22674, n22675,
    n22676, n22677, n22678, n22679, n22680, n22681,
    n22682, n22683, n22684, n22685, n22686, n22687,
    n22688, n22689, n22690, n22691, n22692, n22693,
    n22694, n22695, n22696, n22697, n22698, n22699,
    n22700, n22701, n22702, n22703, n22704, n22705,
    n22706, n22707, n22708, n22709, n22710, n22711,
    n22712, n22713, n22714, n22715, n22716, n22717,
    n22718, n22719, n22720, n22721, n22722, n22723,
    n22724, n22725, n22726, n22727, n22728, n22729,
    n22730, n22731, n22732, n22733, n22734, n22735,
    n22736, n22737, n22738, n22739, n22740, n22741,
    n22742, n22743, n22744, n22745, n22746, n22747,
    n22748, n22749, n22750, n22751, n22752, n22753,
    n22754, n22755, n22756, n22757, n22758, n22759,
    n22760, n22761, n22762, n22763, n22764, n22765,
    n22766, n22767, n22768, n22769, n22770, n22771,
    n22772, n22773, n22774, n22775, n22776, n22777,
    n22778, n22779, n22780, n22781, n22782, n22783,
    n22784, n22785, n22786, n22787, n22788, n22789,
    n22790, n22791, n22792, n22793, n22794, n22795,
    n22796, n22797, n22798, n22799, n22800, n22801,
    n22802, n22803, n22804, n22805, n22806, n22807,
    n22808, n22809, n22810, n22811, n22812, n22813,
    n22814, n22815, n22816, n22818, n22819, n22820,
    n22821, n22822, n22823, n22824, n22825, n22826,
    n22827, n22828, n22829, n22830, n22831, n22832,
    n22833, n22834, n22835, n22836, n22837, n22838,
    n22839, n22840, n22841, n22842, n22843, n22844,
    n22845, n22846, n22847, n22848, n22849, n22850,
    n22851, n22852, n22853, n22854, n22855, n22856,
    n22857, n22858, n22859, n22860, n22861, n22862,
    n22863, n22864, n22865, n22866, n22867, n22868,
    n22869, n22870, n22871, n22872, n22873, n22874,
    n22875, n22876, n22877, n22878, n22879, n22880,
    n22881, n22882, n22883, n22884, n22885, n22886,
    n22887, n22888, n22889, n22890, n22891, n22892,
    n22893, n22894, n22895, n22896, n22897, n22898,
    n22899, n22900, n22901, n22902, n22903, n22904,
    n22905, n22906, n22907, n22908, n22909, n22910,
    n22911, n22912, n22913, n22914, n22915, n22916,
    n22917, n22918, n22919, n22920, n22921, n22922,
    n22923, n22924, n22925, n22926, n22927, n22928,
    n22929, n22930, n22931, n22932, n22933, n22934,
    n22935, n22936, n22937, n22938, n22939, n22940,
    n22941, n22942, n22943, n22944, n22945, n22946,
    n22947, n22948, n22949, n22950, n22951, n22952,
    n22953, n22954, n22955, n22956, n22957, n22958,
    n22959, n22960, n22961, n22962, n22963, n22964,
    n22965, n22966, n22967, n22968, n22969, n22970,
    n22971, n22972, n22973, n22974, n22975, n22976,
    n22977, n22978, n22979, n22980, n22981, n22982,
    n22983, n22984, n22985, n22986, n22987, n22988,
    n22989, n22990, n22991, n22992, n22993, n22994,
    n22995, n22996, n22997, n22998, n22999, n23000,
    n23001, n23002, n23003, n23004, n23005, n23006,
    n23007, n23008, n23009, n23010, n23011, n23012,
    n23013, n23014, n23015, n23016, n23017, n23018,
    n23019, n23020, n23021, n23022, n23023, n23024,
    n23025, n23026, n23027, n23028, n23029, n23030,
    n23031, n23032, n23033, n23034, n23035, n23036,
    n23037, n23038, n23039, n23040, n23041, n23042,
    n23043, n23044, n23045, n23046, n23047, n23048,
    n23049, n23051, n23052, n23053, n23054, n23055,
    n23056, n23057, n23058, n23059, n23060, n23061,
    n23062, n23063, n23064, n23065, n23066, n23067,
    n23068, n23069, n23070, n23071, n23072, n23073,
    n23074, n23075, n23076, n23077, n23078, n23079,
    n23080, n23081, n23082, n23083, n23084, n23085,
    n23086, n23087, n23088, n23089, n23090, n23091,
    n23092, n23093, n23094, n23095, n23096, n23097,
    n23098, n23099, n23100, n23101, n23102, n23103,
    n23104, n23105, n23106, n23107, n23108, n23109,
    n23110, n23111, n23112, n23113, n23114, n23115,
    n23116, n23117, n23118, n23119, n23120, n23121,
    n23122, n23123, n23124, n23125, n23126, n23127,
    n23128, n23129, n23130, n23131, n23132, n23133,
    n23134, n23135, n23136, n23137, n23138, n23139,
    n23140, n23141, n23142, n23143, n23144, n23145,
    n23146, n23147, n23148, n23149, n23150, n23151,
    n23152, n23153, n23154, n23155, n23156, n23157,
    n23158, n23159, n23160, n23161, n23162, n23163,
    n23164, n23165, n23166, n23167, n23168, n23169,
    n23170, n23171, n23172, n23173, n23174, n23175,
    n23176, n23177, n23178, n23179, n23180, n23181,
    n23182, n23183, n23184, n23185, n23186, n23187,
    n23188, n23189, n23190, n23191, n23192, n23193,
    n23194, n23195, n23196, n23197, n23198, n23199,
    n23200, n23201, n23202, n23203, n23204, n23205,
    n23206, n23207, n23208, n23209, n23210, n23211,
    n23212, n23213, n23214, n23215, n23216, n23217,
    n23218, n23219, n23220, n23221, n23222, n23223,
    n23224, n23225, n23226, n23227, n23228, n23229,
    n23230, n23231, n23232, n23233, n23234, n23235,
    n23236, n23237, n23238, n23239, n23240, n23241,
    n23242, n23243, n23244, n23245, n23246, n23247,
    n23248, n23249, n23250, n23251, n23252, n23253,
    n23254, n23255, n23256, n23257, n23258, n23259,
    n23260, n23261, n23262, n23263, n23264, n23265,
    n23266, n23267, n23268, n23269, n23270, n23271,
    n23272, n23273, n23274, n23275, n23277, n23278,
    n23279, n23280, n23281, n23282, n23283, n23284,
    n23285, n23286, n23287, n23288, n23289, n23290,
    n23291, n23292, n23293, n23294, n23295, n23296,
    n23297, n23298, n23299, n23300, n23301, n23302,
    n23303, n23304, n23305, n23306, n23307, n23308,
    n23309, n23310, n23311, n23312, n23313, n23314,
    n23315, n23316, n23317, n23318, n23319, n23320,
    n23321, n23322, n23323, n23324, n23325, n23326,
    n23327, n23328, n23329, n23330, n23331, n23332,
    n23333, n23334, n23335, n23336, n23337, n23338,
    n23339, n23340, n23341, n23342, n23343, n23344,
    n23345, n23346, n23347, n23348, n23349, n23350,
    n23351, n23352, n23353, n23354, n23355, n23356,
    n23357, n23358, n23359, n23360, n23361, n23362,
    n23363, n23364, n23365, n23366, n23367, n23368,
    n23369, n23370, n23371, n23372, n23373, n23374,
    n23375, n23376, n23377, n23378, n23379, n23380,
    n23381, n23382, n23383, n23384, n23385, n23386,
    n23387, n23388, n23389, n23390, n23391, n23392,
    n23393, n23394, n23395, n23396, n23397, n23398,
    n23399, n23400, n23401, n23402, n23403, n23404,
    n23405, n23406, n23407, n23408, n23409, n23410,
    n23411, n23412, n23413, n23414, n23415, n23416,
    n23417, n23418, n23419, n23420, n23421, n23422,
    n23423, n23424, n23425, n23426, n23427, n23428,
    n23429, n23430, n23431, n23432, n23433, n23434,
    n23435, n23436, n23437, n23438, n23439, n23440,
    n23441, n23442, n23443, n23444, n23445, n23446,
    n23447, n23448, n23449, n23450, n23451, n23452,
    n23453, n23454, n23455, n23456, n23457, n23458,
    n23459, n23460, n23461, n23462, n23463, n23464,
    n23465, n23466, n23467, n23468, n23469, n23470,
    n23471, n23472, n23473, n23474, n23475, n23476,
    n23477, n23478, n23479, n23480, n23481, n23482,
    n23483, n23484, n23485, n23486, n23487, n23488,
    n23489, n23490, n23491, n23492, n23494, n23495,
    n23496, n23497, n23498, n23499, n23500, n23501,
    n23502, n23503, n23504, n23505, n23506, n23507,
    n23508, n23509, n23510, n23511, n23512, n23513,
    n23514, n23515, n23516, n23517, n23518, n23519,
    n23520, n23521, n23522, n23523, n23524, n23525,
    n23526, n23527, n23528, n23529, n23530, n23531,
    n23532, n23533, n23534, n23535, n23536, n23537,
    n23538, n23539, n23540, n23541, n23542, n23543,
    n23544, n23545, n23546, n23547, n23548, n23549,
    n23550, n23551, n23552, n23553, n23554, n23555,
    n23556, n23557, n23558, n23559, n23560, n23561,
    n23562, n23563, n23564, n23565, n23566, n23567,
    n23568, n23569, n23570, n23571, n23572, n23573,
    n23574, n23575, n23576, n23577, n23578, n23579,
    n23580, n23581, n23582, n23583, n23584, n23585,
    n23586, n23587, n23588, n23589, n23590, n23591,
    n23592, n23593, n23594, n23595, n23596, n23597,
    n23598, n23599, n23600, n23601, n23602, n23603,
    n23604, n23605, n23606, n23607, n23608, n23609,
    n23610, n23611, n23612, n23613, n23614, n23615,
    n23616, n23617, n23618, n23619, n23620, n23621,
    n23622, n23623, n23624, n23625, n23626, n23627,
    n23628, n23629, n23630, n23631, n23632, n23633,
    n23634, n23635, n23636, n23637, n23638, n23639,
    n23640, n23641, n23642, n23643, n23644, n23645,
    n23646, n23647, n23648, n23649, n23650, n23651,
    n23652, n23653, n23654, n23655, n23656, n23657,
    n23658, n23659, n23660, n23661, n23662, n23663,
    n23664, n23665, n23666, n23667, n23668, n23669,
    n23670, n23671, n23672, n23673, n23674, n23675,
    n23676, n23677, n23678, n23679, n23680, n23681,
    n23682, n23683, n23684, n23685, n23686, n23687,
    n23688, n23689, n23690, n23691, n23692, n23693,
    n23694, n23695, n23696, n23697, n23698, n23699,
    n23700, n23701, n23702, n23703, n23704, n23705,
    n23706, n23708, n23709, n23710, n23711, n23712,
    n23713, n23714, n23715, n23716, n23717, n23718,
    n23719, n23720, n23721, n23722, n23723, n23724,
    n23725, n23726, n23727, n23728, n23729, n23730,
    n23731, n23732, n23733, n23734, n23735, n23736,
    n23737, n23738, n23739, n23740, n23741, n23742,
    n23743, n23744, n23745, n23746, n23747, n23748,
    n23749, n23750, n23751, n23752, n23753, n23754,
    n23755, n23756, n23757, n23758, n23759, n23760,
    n23761, n23762, n23763, n23764, n23765, n23766,
    n23767, n23768, n23769, n23770, n23771, n23772,
    n23773, n23774, n23775, n23776, n23777, n23778,
    n23779, n23780, n23781, n23782, n23783, n23784,
    n23785, n23786, n23787, n23788, n23789, n23790,
    n23791, n23792, n23793, n23794, n23795, n23796,
    n23797, n23798, n23799, n23800, n23801, n23802,
    n23803, n23804, n23805, n23806, n23807, n23808,
    n23809, n23810, n23811, n23812, n23813, n23814,
    n23815, n23816, n23817, n23818, n23819, n23820,
    n23821, n23822, n23823, n23824, n23825, n23826,
    n23827, n23828, n23829, n23830, n23831, n23832,
    n23833, n23834, n23835, n23836, n23837, n23838,
    n23839, n23840, n23841, n23842, n23843, n23844,
    n23845, n23846, n23847, n23848, n23849, n23850,
    n23851, n23852, n23853, n23854, n23855, n23856,
    n23857, n23858, n23859, n23860, n23861, n23862,
    n23863, n23864, n23865, n23866, n23867, n23868,
    n23869, n23870, n23871, n23872, n23873, n23874,
    n23875, n23876, n23877, n23878, n23879, n23880,
    n23881, n23882, n23883, n23884, n23885, n23886,
    n23887, n23888, n23889, n23890, n23891, n23892,
    n23893, n23894, n23895, n23896, n23897, n23898,
    n23899, n23900, n23901, n23902, n23903, n23904,
    n23905, n23906, n23907, n23908, n23909, n23910,
    n23911, n23912, n23913, n23914, n23916, n23917,
    n23918, n23919, n23920, n23921, n23922, n23923,
    n23924, n23925, n23926, n23927, n23928, n23929,
    n23930, n23931, n23932, n23933, n23934, n23935,
    n23936, n23937, n23938, n23939, n23940, n23941,
    n23942, n23943, n23944, n23945, n23946, n23947,
    n23948, n23949, n23950, n23951, n23952, n23953,
    n23954, n23955, n23956, n23957, n23958, n23959,
    n23960, n23961, n23962, n23963, n23964, n23965,
    n23966, n23967, n23968, n23969, n23970, n23971,
    n23972, n23973, n23974, n23975, n23976, n23977,
    n23978, n23979, n23980, n23981, n23982, n23983,
    n23984, n23985, n23986, n23987, n23988, n23989,
    n23990, n23991, n23992, n23993, n23994, n23995,
    n23996, n23997, n23998, n23999, n24000, n24001,
    n24002, n24003, n24004, n24005, n24006, n24007,
    n24008, n24009, n24010, n24011, n24012, n24013,
    n24014, n24015, n24016, n24017, n24018, n24019,
    n24020, n24021, n24022, n24023, n24024, n24025,
    n24026, n24027, n24028, n24029, n24030, n24031,
    n24032, n24033, n24034, n24035, n24036, n24037,
    n24038, n24039, n24040, n24041, n24042, n24043,
    n24044, n24045, n24046, n24047, n24048, n24049,
    n24050, n24051, n24052, n24053, n24054, n24055,
    n24056, n24057, n24058, n24059, n24060, n24061,
    n24062, n24063, n24064, n24065, n24066, n24067,
    n24068, n24069, n24070, n24071, n24072, n24073,
    n24074, n24075, n24076, n24077, n24078, n24079,
    n24080, n24081, n24082, n24083, n24084, n24085,
    n24086, n24087, n24088, n24089, n24090, n24091,
    n24092, n24093, n24094, n24095, n24096, n24097,
    n24098, n24099, n24100, n24101, n24102, n24103,
    n24104, n24105, n24106, n24107, n24108, n24109,
    n24110, n24111, n24113, n24114, n24115, n24116,
    n24117, n24118, n24119, n24120, n24121, n24122,
    n24123, n24124, n24125, n24126, n24127, n24128,
    n24129, n24130, n24131, n24132, n24133, n24134,
    n24135, n24136, n24137, n24138, n24139, n24140,
    n24141, n24142, n24143, n24144, n24145, n24146,
    n24147, n24148, n24149, n24150, n24151, n24152,
    n24153, n24154, n24155, n24156, n24157, n24158,
    n24159, n24160, n24161, n24162, n24163, n24164,
    n24165, n24166, n24167, n24168, n24169, n24170,
    n24171, n24172, n24173, n24174, n24175, n24176,
    n24177, n24178, n24179, n24180, n24181, n24182,
    n24183, n24184, n24185, n24186, n24187, n24188,
    n24189, n24190, n24191, n24192, n24193, n24194,
    n24195, n24196, n24197, n24198, n24199, n24200,
    n24201, n24202, n24203, n24204, n24205, n24206,
    n24207, n24208, n24209, n24210, n24211, n24212,
    n24213, n24214, n24215, n24216, n24217, n24218,
    n24219, n24220, n24221, n24222, n24223, n24224,
    n24225, n24226, n24227, n24228, n24229, n24230,
    n24231, n24232, n24233, n24234, n24235, n24236,
    n24237, n24238, n24239, n24240, n24241, n24242,
    n24243, n24244, n24245, n24246, n24247, n24248,
    n24249, n24250, n24251, n24252, n24253, n24254,
    n24255, n24256, n24257, n24258, n24259, n24260,
    n24261, n24262, n24263, n24264, n24265, n24266,
    n24267, n24268, n24269, n24270, n24271, n24272,
    n24273, n24274, n24275, n24276, n24277, n24278,
    n24279, n24280, n24281, n24282, n24283, n24284,
    n24285, n24286, n24287, n24288, n24289, n24290,
    n24291, n24292, n24293, n24294, n24295, n24296,
    n24297, n24298, n24299, n24300, n24301, n24302,
    n24303, n24304, n24305, n24306, n24308, n24309,
    n24310, n24311, n24312, n24313, n24314, n24315,
    n24316, n24317, n24318, n24319, n24320, n24321,
    n24322, n24323, n24324, n24325, n24326, n24327,
    n24328, n24329, n24330, n24331, n24332, n24333,
    n24334, n24335, n24336, n24337, n24338, n24339,
    n24340, n24341, n24342, n24343, n24344, n24345,
    n24346, n24347, n24348, n24349, n24350, n24351,
    n24352, n24353, n24354, n24355, n24356, n24357,
    n24358, n24359, n24360, n24361, n24362, n24363,
    n24364, n24365, n24366, n24367, n24368, n24369,
    n24370, n24371, n24372, n24373, n24374, n24375,
    n24376, n24377, n24378, n24379, n24380, n24381,
    n24382, n24383, n24384, n24385, n24386, n24387,
    n24388, n24389, n24390, n24391, n24392, n24393,
    n24394, n24395, n24396, n24397, n24398, n24399,
    n24400, n24401, n24402, n24403, n24404, n24405,
    n24406, n24407, n24408, n24409, n24410, n24411,
    n24412, n24413, n24414, n24415, n24416, n24417,
    n24418, n24419, n24420, n24421, n24422, n24423,
    n24424, n24425, n24426, n24427, n24428, n24429,
    n24430, n24431, n24432, n24433, n24434, n24435,
    n24436, n24437, n24438, n24439, n24440, n24441,
    n24442, n24443, n24444, n24445, n24446, n24447,
    n24448, n24449, n24450, n24451, n24452, n24453,
    n24454, n24455, n24456, n24457, n24458, n24459,
    n24460, n24461, n24462, n24463, n24464, n24465,
    n24466, n24467, n24468, n24469, n24470, n24471,
    n24472, n24473, n24474, n24475, n24476, n24477,
    n24478, n24479, n24480, n24481, n24482, n24483,
    n24484, n24485, n24486, n24487, n24488, n24489,
    n24490, n24491, n24492, n24493, n24495, n24496,
    n24497, n24498, n24499, n24500, n24501, n24502,
    n24503, n24504, n24505, n24506, n24507, n24508,
    n24509, n24510, n24511, n24512, n24513, n24514,
    n24515, n24516, n24517, n24518, n24519, n24520,
    n24521, n24522, n24523, n24524, n24525, n24526,
    n24527, n24528, n24529, n24530, n24531, n24532,
    n24533, n24534, n24535, n24536, n24537, n24538,
    n24539, n24540, n24541, n24542, n24543, n24544,
    n24545, n24546, n24547, n24548, n24549, n24550,
    n24551, n24552, n24553, n24554, n24555, n24556,
    n24557, n24558, n24559, n24560, n24561, n24562,
    n24563, n24564, n24565, n24566, n24567, n24568,
    n24569, n24570, n24571, n24572, n24573, n24574,
    n24575, n24576, n24577, n24578, n24579, n24580,
    n24581, n24582, n24583, n24584, n24585, n24586,
    n24587, n24588, n24589, n24590, n24591, n24592,
    n24593, n24594, n24595, n24596, n24597, n24598,
    n24599, n24600, n24601, n24602, n24603, n24604,
    n24605, n24606, n24607, n24608, n24609, n24610,
    n24611, n24612, n24613, n24614, n24615, n24616,
    n24617, n24618, n24619, n24620, n24621, n24622,
    n24623, n24624, n24625, n24626, n24627, n24628,
    n24629, n24630, n24631, n24632, n24633, n24634,
    n24635, n24636, n24637, n24638, n24639, n24640,
    n24641, n24642, n24643, n24644, n24645, n24646,
    n24647, n24648, n24649, n24650, n24651, n24652,
    n24653, n24654, n24655, n24656, n24657, n24658,
    n24659, n24660, n24661, n24662, n24663, n24664,
    n24665, n24666, n24667, n24668, n24669, n24670,
    n24671, n24672, n24673, n24674, n24675, n24677,
    n24678, n24679, n24680, n24681, n24682, n24683,
    n24684, n24685, n24686, n24687, n24688, n24689,
    n24690, n24691, n24692, n24693, n24694, n24695,
    n24696, n24697, n24698, n24699, n24700, n24701,
    n24702, n24703, n24704, n24705, n24706, n24707,
    n24708, n24709, n24710, n24711, n24712, n24713,
    n24714, n24715, n24716, n24717, n24718, n24719,
    n24720, n24721, n24722, n24723, n24724, n24725,
    n24726, n24727, n24728, n24729, n24730, n24731,
    n24732, n24733, n24734, n24735, n24736, n24737,
    n24738, n24739, n24740, n24741, n24742, n24743,
    n24744, n24745, n24746, n24747, n24748, n24749,
    n24750, n24751, n24752, n24753, n24754, n24755,
    n24756, n24757, n24758, n24759, n24760, n24761,
    n24762, n24763, n24764, n24765, n24766, n24767,
    n24768, n24769, n24770, n24771, n24772, n24773,
    n24774, n24775, n24776, n24777, n24778, n24779,
    n24780, n24781, n24782, n24783, n24784, n24785,
    n24786, n24787, n24788, n24789, n24790, n24791,
    n24792, n24793, n24794, n24795, n24796, n24797,
    n24798, n24799, n24800, n24801, n24802, n24803,
    n24804, n24805, n24806, n24807, n24808, n24809,
    n24810, n24811, n24812, n24813, n24814, n24815,
    n24816, n24817, n24818, n24819, n24820, n24821,
    n24822, n24823, n24824, n24825, n24826, n24827,
    n24828, n24829, n24830, n24831, n24832, n24833,
    n24834, n24835, n24836, n24837, n24838, n24839,
    n24840, n24841, n24842, n24843, n24844, n24845,
    n24846, n24847, n24848, n24849, n24850, n24851,
    n24853, n24854, n24855, n24856, n24857, n24858,
    n24859, n24860, n24861, n24862, n24863, n24864,
    n24865, n24866, n24867, n24868, n24869, n24870,
    n24871, n24872, n24873, n24874, n24875, n24876,
    n24877, n24878, n24879, n24880, n24881, n24882,
    n24883, n24884, n24885, n24886, n24887, n24888,
    n24889, n24890, n24891, n24892, n24893, n24894,
    n24895, n24896, n24897, n24898, n24899, n24900,
    n24901, n24902, n24903, n24904, n24905, n24906,
    n24907, n24908, n24909, n24910, n24911, n24912,
    n24913, n24914, n24915, n24916, n24917, n24918,
    n24919, n24920, n24921, n24922, n24923, n24924,
    n24925, n24926, n24927, n24928, n24929, n24930,
    n24931, n24932, n24933, n24934, n24935, n24936,
    n24937, n24938, n24939, n24940, n24941, n24942,
    n24943, n24944, n24945, n24946, n24947, n24948,
    n24949, n24950, n24951, n24952, n24953, n24954,
    n24955, n24956, n24957, n24958, n24959, n24960,
    n24961, n24962, n24963, n24964, n24965, n24966,
    n24967, n24968, n24969, n24970, n24971, n24972,
    n24973, n24974, n24975, n24976, n24977, n24978,
    n24979, n24980, n24981, n24982, n24983, n24984,
    n24985, n24986, n24987, n24988, n24989, n24990,
    n24991, n24992, n24993, n24994, n24995, n24996,
    n24997, n24998, n24999, n25000, n25001, n25002,
    n25003, n25004, n25005, n25006, n25007, n25008,
    n25009, n25010, n25011, n25012, n25013, n25014,
    n25015, n25016, n25017, n25018, n25019, n25020,
    n25021, n25023, n25024, n25025, n25026, n25027,
    n25028, n25029, n25030, n25031, n25032, n25033,
    n25034, n25035, n25036, n25037, n25038, n25039,
    n25040, n25041, n25042, n25043, n25044, n25045,
    n25046, n25047, n25048, n25049, n25050, n25051,
    n25052, n25053, n25054, n25055, n25056, n25057,
    n25058, n25059, n25060, n25061, n25062, n25063,
    n25064, n25065, n25066, n25067, n25068, n25069,
    n25070, n25071, n25072, n25073, n25074, n25075,
    n25076, n25077, n25078, n25079, n25080, n25081,
    n25082, n25083, n25084, n25085, n25086, n25087,
    n25088, n25089, n25090, n25091, n25092, n25093,
    n25094, n25095, n25096, n25097, n25098, n25099,
    n25100, n25101, n25102, n25103, n25104, n25105,
    n25106, n25107, n25108, n25109, n25110, n25111,
    n25112, n25113, n25114, n25115, n25116, n25117,
    n25118, n25119, n25120, n25121, n25122, n25123,
    n25124, n25125, n25126, n25127, n25128, n25129,
    n25130, n25131, n25132, n25133, n25134, n25135,
    n25136, n25137, n25138, n25139, n25140, n25141,
    n25142, n25143, n25144, n25145, n25146, n25147,
    n25148, n25149, n25150, n25151, n25152, n25153,
    n25154, n25155, n25156, n25157, n25158, n25159,
    n25160, n25161, n25162, n25163, n25164, n25165,
    n25166, n25167, n25168, n25169, n25170, n25171,
    n25172, n25173, n25174, n25175, n25176, n25177,
    n25178, n25179, n25180, n25181, n25182, n25184,
    n25185, n25186, n25187, n25188, n25189, n25190,
    n25191, n25192, n25193, n25194, n25195, n25196,
    n25197, n25198, n25199, n25200, n25201, n25202,
    n25203, n25204, n25205, n25206, n25207, n25208,
    n25209, n25210, n25211, n25212, n25213, n25214,
    n25215, n25216, n25217, n25218, n25219, n25220,
    n25221, n25222, n25223, n25224, n25225, n25226,
    n25227, n25228, n25229, n25230, n25231, n25232,
    n25233, n25234, n25235, n25236, n25237, n25238,
    n25239, n25240, n25241, n25242, n25243, n25244,
    n25245, n25246, n25247, n25248, n25249, n25250,
    n25251, n25252, n25253, n25254, n25255, n25256,
    n25257, n25258, n25259, n25260, n25261, n25262,
    n25263, n25264, n25265, n25266, n25267, n25268,
    n25269, n25270, n25271, n25272, n25273, n25274,
    n25275, n25276, n25277, n25278, n25279, n25280,
    n25281, n25282, n25283, n25284, n25285, n25286,
    n25287, n25288, n25289, n25290, n25291, n25292,
    n25293, n25294, n25295, n25296, n25297, n25298,
    n25299, n25300, n25301, n25302, n25303, n25304,
    n25305, n25306, n25307, n25308, n25309, n25310,
    n25311, n25312, n25313, n25314, n25315, n25316,
    n25317, n25318, n25319, n25320, n25321, n25322,
    n25323, n25324, n25325, n25326, n25327, n25328,
    n25329, n25330, n25331, n25332, n25333, n25334,
    n25335, n25336, n25337, n25338, n25339, n25341,
    n25342, n25343, n25344, n25345, n25346, n25347,
    n25348, n25349, n25350, n25351, n25352, n25353,
    n25354, n25355, n25356, n25357, n25358, n25359,
    n25360, n25361, n25362, n25363, n25364, n25365,
    n25366, n25367, n25368, n25369, n25370, n25371,
    n25372, n25373, n25374, n25375, n25376, n25377,
    n25378, n25379, n25380, n25381, n25382, n25383,
    n25384, n25385, n25386, n25387, n25388, n25389,
    n25390, n25391, n25392, n25393, n25394, n25395,
    n25396, n25397, n25398, n25399, n25400, n25401,
    n25402, n25403, n25404, n25405, n25406, n25407,
    n25408, n25409, n25410, n25411, n25412, n25413,
    n25414, n25415, n25416, n25417, n25418, n25419,
    n25420, n25421, n25422, n25423, n25424, n25425,
    n25426, n25427, n25428, n25429, n25430, n25431,
    n25432, n25433, n25434, n25435, n25436, n25437,
    n25438, n25439, n25440, n25441, n25442, n25443,
    n25444, n25445, n25446, n25447, n25448, n25449,
    n25450, n25451, n25452, n25453, n25454, n25455,
    n25456, n25457, n25458, n25459, n25460, n25461,
    n25462, n25463, n25464, n25465, n25466, n25467,
    n25468, n25469, n25470, n25471, n25472, n25473,
    n25474, n25475, n25476, n25477, n25478, n25479,
    n25480, n25481, n25482, n25483, n25484, n25485,
    n25486, n25487, n25488, n25489, n25490, n25492,
    n25493, n25494, n25495, n25496, n25497, n25498,
    n25499, n25500, n25501, n25502, n25503, n25504,
    n25505, n25506, n25507, n25508, n25509, n25510,
    n25511, n25512, n25513, n25514, n25515, n25516,
    n25517, n25518, n25519, n25520, n25521, n25522,
    n25523, n25524, n25525, n25526, n25527, n25528,
    n25529, n25530, n25531, n25532, n25533, n25534,
    n25535, n25536, n25537, n25538, n25539, n25540,
    n25541, n25542, n25543, n25544, n25545, n25546,
    n25547, n25548, n25549, n25550, n25551, n25552,
    n25553, n25554, n25555, n25556, n25557, n25558,
    n25559, n25560, n25561, n25562, n25563, n25564,
    n25565, n25566, n25567, n25568, n25569, n25570,
    n25571, n25572, n25573, n25574, n25575, n25576,
    n25577, n25578, n25579, n25580, n25581, n25582,
    n25583, n25584, n25585, n25586, n25587, n25588,
    n25589, n25590, n25591, n25592, n25593, n25594,
    n25595, n25596, n25597, n25598, n25599, n25600,
    n25601, n25602, n25603, n25604, n25605, n25606,
    n25607, n25608, n25609, n25610, n25611, n25612,
    n25613, n25614, n25615, n25616, n25617, n25618,
    n25619, n25620, n25621, n25622, n25623, n25624,
    n25625, n25626, n25627, n25628, n25629, n25630,
    n25631, n25632, n25633, n25635, n25636, n25637,
    n25638, n25639, n25640, n25641, n25642, n25643,
    n25644, n25645, n25646, n25647, n25648, n25649,
    n25650, n25651, n25652, n25653, n25654, n25655,
    n25656, n25657, n25658, n25659, n25660, n25661,
    n25662, n25663, n25664, n25665, n25666, n25667,
    n25668, n25669, n25670, n25671, n25672, n25673,
    n25674, n25675, n25676, n25677, n25678, n25679,
    n25680, n25681, n25682, n25683, n25684, n25685,
    n25686, n25687, n25688, n25689, n25690, n25691,
    n25692, n25693, n25694, n25695, n25696, n25697,
    n25698, n25699, n25700, n25701, n25702, n25703,
    n25704, n25705, n25706, n25707, n25708, n25709,
    n25710, n25711, n25712, n25713, n25714, n25715,
    n25716, n25717, n25718, n25719, n25720, n25721,
    n25722, n25723, n25724, n25725, n25726, n25727,
    n25728, n25729, n25730, n25731, n25732, n25733,
    n25734, n25735, n25736, n25737, n25738, n25739,
    n25740, n25741, n25742, n25743, n25744, n25745,
    n25746, n25747, n25748, n25749, n25750, n25751,
    n25752, n25753, n25754, n25755, n25756, n25757,
    n25758, n25759, n25760, n25761, n25762, n25763,
    n25764, n25765, n25766, n25767, n25768, n25769,
    n25770, n25771, n25772, n25773, n25775, n25776,
    n25777, n25778, n25779, n25780, n25781, n25782,
    n25783, n25784, n25785, n25786, n25787, n25788,
    n25789, n25790, n25791, n25792, n25793, n25794,
    n25795, n25796, n25797, n25798, n25799, n25800,
    n25801, n25802, n25803, n25804, n25805, n25806,
    n25807, n25808, n25809, n25810, n25811, n25812,
    n25813, n25814, n25815, n25816, n25817, n25818,
    n25819, n25820, n25821, n25822, n25823, n25824,
    n25825, n25826, n25827, n25828, n25829, n25830,
    n25831, n25832, n25833, n25834, n25835, n25836,
    n25837, n25838, n25839, n25840, n25841, n25842,
    n25843, n25844, n25845, n25846, n25847, n25848,
    n25849, n25850, n25851, n25852, n25853, n25854,
    n25855, n25856, n25857, n25858, n25859, n25860,
    n25861, n25862, n25863, n25864, n25865, n25866,
    n25867, n25868, n25869, n25870, n25871, n25872,
    n25873, n25874, n25875, n25876, n25877, n25878,
    n25879, n25880, n25881, n25882, n25883, n25884,
    n25885, n25886, n25887, n25888, n25889, n25890,
    n25891, n25892, n25893, n25894, n25895, n25896,
    n25897, n25898, n25899, n25900, n25901, n25902,
    n25903, n25905, n25906, n25907, n25908, n25909,
    n25910, n25911, n25912, n25913, n25914, n25915,
    n25916, n25917, n25918, n25919, n25920, n25921,
    n25922, n25923, n25924, n25925, n25926, n25927,
    n25928, n25929, n25930, n25931, n25932, n25933,
    n25934, n25935, n25936, n25937, n25938, n25939,
    n25940, n25941, n25942, n25943, n25944, n25945,
    n25946, n25947, n25948, n25949, n25950, n25951,
    n25952, n25953, n25954, n25955, n25956, n25957,
    n25958, n25959, n25960, n25961, n25962, n25963,
    n25964, n25965, n25966, n25967, n25968, n25969,
    n25970, n25971, n25972, n25973, n25974, n25975,
    n25976, n25977, n25978, n25979, n25980, n25981,
    n25982, n25983, n25984, n25985, n25986, n25987,
    n25988, n25989, n25990, n25991, n25992, n25993,
    n25994, n25995, n25996, n25997, n25998, n25999,
    n26000, n26001, n26002, n26003, n26004, n26005,
    n26006, n26007, n26008, n26009, n26010, n26011,
    n26012, n26013, n26014, n26015, n26016, n26017,
    n26018, n26019, n26020, n26021, n26022, n26023,
    n26024, n26025, n26027, n26028, n26029, n26030,
    n26031, n26032, n26033, n26034, n26035, n26036,
    n26037, n26038, n26039, n26040, n26041, n26042,
    n26043, n26044, n26045, n26046, n26047, n26048,
    n26049, n26050, n26051, n26052, n26053, n26054,
    n26055, n26056, n26057, n26058, n26059, n26060,
    n26061, n26062, n26063, n26064, n26065, n26066,
    n26067, n26068, n26069, n26070, n26071, n26072,
    n26073, n26074, n26075, n26076, n26077, n26078,
    n26079, n26080, n26081, n26082, n26083, n26084,
    n26085, n26086, n26087, n26088, n26089, n26090,
    n26091, n26092, n26093, n26094, n26095, n26096,
    n26097, n26098, n26099, n26100, n26101, n26102,
    n26103, n26104, n26105, n26106, n26107, n26108,
    n26109, n26110, n26111, n26112, n26113, n26114,
    n26115, n26116, n26117, n26118, n26119, n26120,
    n26121, n26122, n26123, n26124, n26125, n26126,
    n26127, n26128, n26129, n26130, n26131, n26132,
    n26133, n26134, n26135, n26136, n26137, n26138,
    n26139, n26140, n26141, n26142, n26143, n26144,
    n26145, n26146, n26147, n26149, n26150, n26151,
    n26152, n26153, n26154, n26155, n26156, n26157,
    n26158, n26159, n26160, n26161, n26162, n26163,
    n26164, n26165, n26166, n26167, n26168, n26169,
    n26170, n26171, n26172, n26173, n26174, n26175,
    n26176, n26177, n26178, n26179, n26180, n26181,
    n26182, n26183, n26184, n26185, n26186, n26187,
    n26188, n26189, n26190, n26191, n26192, n26193,
    n26194, n26195, n26196, n26197, n26198, n26199,
    n26200, n26201, n26202, n26203, n26204, n26205,
    n26206, n26207, n26208, n26209, n26210, n26211,
    n26212, n26213, n26214, n26215, n26216, n26217,
    n26218, n26219, n26220, n26221, n26222, n26223,
    n26224, n26225, n26226, n26227, n26228, n26229,
    n26230, n26231, n26232, n26233, n26234, n26235,
    n26236, n26237, n26238, n26239, n26240, n26241,
    n26242, n26243, n26244, n26245, n26246, n26247,
    n26248, n26249, n26250, n26251, n26252, n26253,
    n26254, n26255, n26256, n26257, n26259, n26260,
    n26261, n26262, n26263, n26264, n26265, n26266,
    n26267, n26268, n26269, n26270, n26271, n26272,
    n26273, n26274, n26275, n26276, n26277, n26278,
    n26279, n26280, n26281, n26282, n26283, n26284,
    n26285, n26286, n26287, n26288, n26289, n26290,
    n26291, n26292, n26293, n26294, n26295, n26296,
    n26297, n26298, n26299, n26300, n26301, n26302,
    n26303, n26304, n26305, n26306, n26307, n26308,
    n26309, n26310, n26311, n26312, n26313, n26314,
    n26315, n26316, n26317, n26318, n26319, n26320,
    n26321, n26322, n26323, n26324, n26325, n26326,
    n26327, n26328, n26329, n26330, n26331, n26332,
    n26333, n26334, n26335, n26336, n26337, n26338,
    n26339, n26340, n26341, n26342, n26343, n26344,
    n26345, n26346, n26347, n26348, n26349, n26350,
    n26351, n26352, n26353, n26354, n26355, n26356,
    n26357, n26358, n26359, n26360, n26362, n26363,
    n26364, n26365, n26366, n26367, n26368, n26369,
    n26370, n26371, n26372, n26373, n26374, n26375,
    n26376, n26377, n26378, n26379, n26380, n26381,
    n26382, n26383, n26384, n26385, n26386, n26387,
    n26388, n26389, n26390, n26391, n26392, n26393,
    n26394, n26395, n26396, n26397, n26398, n26399,
    n26400, n26401, n26402, n26403, n26404, n26405,
    n26406, n26407, n26408, n26409, n26410, n26411,
    n26412, n26413, n26414, n26415, n26416, n26417,
    n26418, n26419, n26420, n26421, n26422, n26423,
    n26424, n26425, n26426, n26427, n26428, n26429,
    n26430, n26431, n26432, n26433, n26434, n26435,
    n26436, n26437, n26438, n26439, n26440, n26441,
    n26442, n26443, n26444, n26445, n26446, n26447,
    n26448, n26449, n26450, n26451, n26452, n26453,
    n26454, n26455, n26456, n26457, n26458, n26459,
    n26460, n26461, n26463, n26464, n26465, n26466,
    n26467, n26468, n26469, n26470, n26471, n26472,
    n26473, n26474, n26475, n26476, n26477, n26478,
    n26479, n26480, n26481, n26482, n26483, n26484,
    n26485, n26486, n26487, n26488, n26489, n26490,
    n26491, n26492, n26493, n26494, n26495, n26496,
    n26497, n26498, n26499, n26500, n26501, n26502,
    n26503, n26504, n26505, n26506, n26507, n26508,
    n26509, n26510, n26511, n26512, n26513, n26514,
    n26515, n26516, n26517, n26518, n26519, n26520,
    n26521, n26522, n26523, n26524, n26525, n26526,
    n26527, n26528, n26529, n26530, n26531, n26532,
    n26533, n26534, n26535, n26536, n26537, n26538,
    n26539, n26540, n26541, n26542, n26543, n26544,
    n26545, n26546, n26547, n26548, n26549, n26550,
    n26551, n26552, n26553, n26555, n26556, n26557,
    n26558, n26559, n26560, n26561, n26562, n26563,
    n26564, n26565, n26566, n26567, n26568, n26569,
    n26570, n26571, n26572, n26573, n26574, n26575,
    n26576, n26577, n26578, n26579, n26580, n26581,
    n26582, n26583, n26584, n26585, n26586, n26587,
    n26588, n26589, n26590, n26591, n26592, n26593,
    n26594, n26595, n26596, n26597, n26598, n26599,
    n26600, n26601, n26602, n26603, n26604, n26605,
    n26606, n26607, n26608, n26609, n26610, n26611,
    n26612, n26613, n26614, n26615, n26616, n26617,
    n26618, n26619, n26620, n26621, n26622, n26623,
    n26624, n26625, n26626, n26627, n26628, n26629,
    n26630, n26631, n26632, n26633, n26634, n26635,
    n26636, n26638, n26639, n26640, n26641, n26642,
    n26643, n26644, n26645, n26646, n26647, n26648,
    n26649, n26650, n26651, n26652, n26653, n26654,
    n26655, n26656, n26657, n26658, n26659, n26660,
    n26661, n26662, n26663, n26664, n26665, n26666,
    n26667, n26668, n26669, n26670, n26671, n26672,
    n26673, n26674, n26675, n26676, n26677, n26678,
    n26679, n26680, n26681, n26682, n26683, n26684,
    n26685, n26686, n26687, n26688, n26689, n26690,
    n26691, n26692, n26693, n26694, n26695, n26696,
    n26697, n26698, n26699, n26700, n26701, n26702,
    n26703, n26704, n26705, n26706, n26707, n26708,
    n26709, n26710, n26711, n26712, n26713, n26714,
    n26715, n26716, n26717, n26718, n26720, n26721,
    n26722, n26723, n26724, n26725, n26726, n26727,
    n26728, n26729, n26730, n26731, n26732, n26733,
    n26734, n26735, n26736, n26737, n26738, n26739,
    n26740, n26741, n26742, n26743, n26744, n26745,
    n26746, n26747, n26748, n26749, n26750, n26751,
    n26752, n26753, n26754, n26755, n26756, n26757,
    n26758, n26759, n26760, n26761, n26762, n26763,
    n26764, n26765, n26766, n26767, n26768, n26769,
    n26770, n26771, n26772, n26773, n26774, n26775,
    n26776, n26777, n26778, n26779, n26780, n26781,
    n26782, n26783, n26784, n26785, n26786, n26787,
    n26788, n26789, n26790, n26791, n26792, n26793,
    n26795, n26796, n26797, n26798, n26799, n26800,
    n26801, n26802, n26803, n26804, n26805, n26806,
    n26807, n26808, n26809, n26810, n26811, n26812,
    n26813, n26814, n26815, n26816, n26817, n26818,
    n26819, n26820, n26821, n26822, n26823, n26824,
    n26825, n26826, n26827, n26828, n26829, n26830,
    n26831, n26832, n26833, n26834, n26835, n26836,
    n26837, n26838, n26839, n26840, n26841, n26842,
    n26843, n26844, n26845, n26846, n26847, n26848,
    n26849, n26850, n26851, n26852, n26853, n26854,
    n26855, n26856, n26857, n26858, n26859, n26860,
    n26861, n26863, n26864, n26865, n26866, n26867,
    n26868, n26869, n26870, n26871, n26872, n26873,
    n26874, n26875, n26876, n26877, n26878, n26879,
    n26880, n26881, n26882, n26883, n26884, n26885,
    n26886, n26887, n26888, n26889, n26890, n26891,
    n26892, n26893, n26894, n26895, n26896, n26897,
    n26898, n26899, n26900, n26901, n26902, n26903,
    n26904, n26905, n26906, n26907, n26908, n26909,
    n26910, n26911, n26912, n26913, n26914, n26915,
    n26916, n26917, n26918, n26919, n26920, n26921,
    n26922, n26923, n26924, n26925, n26927, n26928,
    n26929, n26930, n26931, n26932, n26933, n26934,
    n26935, n26936, n26937, n26938, n26939, n26940,
    n26941, n26942, n26943, n26944, n26945, n26946,
    n26947, n26948, n26949, n26950, n26951, n26952,
    n26953, n26954, n26955, n26956, n26957, n26958,
    n26959, n26960, n26961, n26962, n26963, n26964,
    n26965, n26966, n26967, n26968, n26969, n26970,
    n26971, n26972, n26973, n26974, n26975, n26976,
    n26977, n26978, n26979, n26980, n26981, n26982,
    n26984, n26985, n26986, n26987, n26988, n26989,
    n26990, n26991, n26992, n26993, n26994, n26995,
    n26996, n26997, n26998, n26999, n27000, n27001,
    n27002, n27003, n27004, n27005, n27006, n27007,
    n27008, n27009, n27010, n27011, n27012, n27013,
    n27014, n27015, n27016, n27017, n27018, n27019,
    n27020, n27021, n27022, n27023, n27024, n27025,
    n27026, n27027, n27028, n27030, n27031, n27032,
    n27033, n27034, n27035, n27036, n27037, n27038,
    n27039, n27040, n27041, n27042, n27043, n27044,
    n27045, n27046, n27047, n27048, n27049, n27050,
    n27051, n27052, n27053, n27054, n27055, n27056,
    n27057, n27058, n27059, n27060, n27061, n27062,
    n27063, n27064, n27065, n27066, n27067, n27068,
    n27069, n27070, n27071, n27072, n27073, n27074,
    n27076, n27077, n27078, n27079, n27080, n27081,
    n27082, n27083, n27084, n27085, n27086, n27087,
    n27088, n27089, n27090, n27091, n27092, n27093,
    n27094, n27095, n27096, n27097, n27098, n27099,
    n27100, n27101, n27102, n27103, n27104, n27105,
    n27106, n27107, n27108, n27109, n27110, n27111,
    n27113, n27114, n27115, n27116, n27117, n27118,
    n27119, n27120, n27121, n27122, n27123, n27124,
    n27125, n27126, n27127, n27128, n27129, n27130,
    n27131, n27132, n27133, n27134, n27135, n27136,
    n27137, n27138, n27139, n27140, n27142, n27143,
    n27144, n27145, n27146, n27147, n27148, n27149,
    n27150, n27151, n27152, n27153, n27154, n27155,
    n27156, n27157, n27158, n27159, n27160, n27161,
    n27162, n27163, n27164, n27165, n27167, n27168,
    n27169, n27170, n27171, n27172, n27173, n27174,
    n27175, n27176, n27177, n27178, n27179, n27180,
    n27181, n27182, n27184, n27185, n27186, n27187,
    n27188, n27189, n27190, n27191;
  assign po0  = pi0  & pi64 ;
  assign n258 = pi2  & ~po0 ;
  assign n259 = ~pi1  & pi2 ;
  assign n260 = pi1  & ~pi2 ;
  assign n261 = ~n259 & ~n260;
  assign n262 = pi0  & ~n261;
  assign n263 = pi64  & ~pi65 ;
  assign n264 = ~pi64  & pi65 ;
  assign n265 = ~n263 & ~n264;
  assign n266 = n262 & ~n265;
  assign n267 = pi0  & n261;
  assign n268 = pi65  & n267;
  assign n269 = ~pi0  & pi1 ;
  assign n270 = pi64  & n269;
  assign n271 = ~n266 & ~n270;
  assign n272 = ~n268 & n271;
  assign n273 = pi2  & ~n272;
  assign n274 = pi2  & ~n273;
  assign n275 = ~n272 & ~n273;
  assign n276 = ~n274 & ~n275;
  assign n277 = n258 & ~n276;
  assign n278 = ~n258 & n276;
  assign po1  = ~n277 & ~n278;
  assign n280 = pi64  & pi65 ;
  assign n281 = ~pi66  & n280;
  assign n282 = ~pi65  & pi66 ;
  assign n283 = pi65  & ~pi66 ;
  assign n284 = ~n280 & ~n282;
  assign n285 = ~n283 & n284;
  assign n286 = ~n281 & ~n285;
  assign n287 = n262 & n286;
  assign n288 = n259 & ~n262;
  assign n289 = pi64  & n288;
  assign n290 = pi66  & n267;
  assign n291 = pi65  & n269;
  assign n292 = ~n290 & ~n291;
  assign n293 = ~n287 & n292;
  assign n294 = ~n289 & n293;
  assign n295 = pi2  & ~n294;
  assign n296 = pi2  & ~n295;
  assign n297 = ~n294 & ~n295;
  assign n298 = ~n296 & ~n297;
  assign n299 = n277 & ~n298;
  assign n300 = ~n277 & n298;
  assign po2  = ~n299 & ~n300;
  assign n302 = pi65  & pi66 ;
  assign n303 = ~n281 & ~n302;
  assign n304 = ~pi66  & ~pi67 ;
  assign n305 = pi66  & pi67 ;
  assign n306 = ~n304 & ~n305;
  assign n307 = ~n303 & n306;
  assign n308 = n303 & ~n306;
  assign n309 = ~n307 & ~n308;
  assign n310 = n262 & n309;
  assign n311 = pi65  & n288;
  assign n312 = pi67  & n267;
  assign n313 = pi66  & n269;
  assign n314 = ~n312 & ~n313;
  assign n315 = ~n311 & n314;
  assign n316 = ~n310 & n315;
  assign n317 = pi2  & ~n316;
  assign n318 = pi2  & ~n317;
  assign n319 = ~n316 & ~n317;
  assign n320 = ~n318 & ~n319;
  assign n321 = pi2  & ~pi3 ;
  assign n322 = ~pi2  & pi3 ;
  assign n323 = ~n321 & ~n322;
  assign n324 = pi64  & ~n323;
  assign n325 = ~n320 & n324;
  assign n326 = n320 & ~n324;
  assign n327 = ~n325 & ~n326;
  assign n328 = n299 & n327;
  assign n329 = ~n299 & ~n327;
  assign po3  = ~n328 & ~n329;
  assign n331 = pi5  & ~n324;
  assign n332 = ~pi3  & pi4 ;
  assign n333 = pi3  & ~pi4 ;
  assign n334 = ~n332 & ~n333;
  assign n335 = n323 & ~n334;
  assign n336 = pi64  & n335;
  assign n337 = ~pi4  & pi5 ;
  assign n338 = pi4  & ~pi5 ;
  assign n339 = ~n337 & ~n338;
  assign n340 = ~n323 & n339;
  assign n341 = pi65  & n340;
  assign n342 = ~n323 & ~n339;
  assign n343 = ~n265 & n342;
  assign n344 = ~n336 & ~n341;
  assign n345 = ~n343 & n344;
  assign n346 = pi5  & ~n345;
  assign n347 = pi5  & ~n346;
  assign n348 = ~n345 & ~n346;
  assign n349 = ~n347 & ~n348;
  assign n350 = n331 & ~n349;
  assign n351 = ~n331 & n349;
  assign n352 = ~n350 & ~n351;
  assign n353 = ~n305 & ~n307;
  assign n354 = ~pi67  & ~pi68 ;
  assign n355 = pi67  & pi68 ;
  assign n356 = ~n354 & ~n355;
  assign n357 = ~n353 & n356;
  assign n358 = n353 & ~n356;
  assign n359 = ~n357 & ~n358;
  assign n360 = n262 & n359;
  assign n361 = pi66  & n288;
  assign n362 = pi68  & n267;
  assign n363 = pi67  & n269;
  assign n364 = ~n362 & ~n363;
  assign n365 = ~n361 & n364;
  assign n366 = ~n360 & n365;
  assign n367 = pi2  & ~n366;
  assign n368 = pi2  & ~n367;
  assign n369 = ~n366 & ~n367;
  assign n370 = ~n368 & ~n369;
  assign n371 = n352 & ~n370;
  assign n372 = n352 & ~n371;
  assign n373 = ~n370 & ~n371;
  assign n374 = ~n372 & ~n373;
  assign n375 = ~n325 & ~n328;
  assign n376 = ~n374 & ~n375;
  assign n377 = n374 & n375;
  assign po4  = ~n376 & ~n377;
  assign n379 = n323 & n334;
  assign n380 = ~n339 & n379;
  assign n381 = pi64  & n380;
  assign n382 = pi66  & n340;
  assign n383 = pi65  & n335;
  assign n384 = ~n382 & ~n383;
  assign n385 = ~n381 & n384;
  assign n386 = ~n342 & n385;
  assign n387 = ~n286 & n385;
  assign n388 = ~n386 & ~n387;
  assign n389 = pi5  & ~n388;
  assign n390 = ~pi5  & n388;
  assign n391 = ~n389 & ~n390;
  assign n392 = n350 & ~n391;
  assign n393 = ~n350 & n391;
  assign n394 = ~n392 & ~n393;
  assign n395 = ~n355 & ~n357;
  assign n396 = ~pi68  & ~pi69 ;
  assign n397 = pi68  & pi69 ;
  assign n398 = ~n396 & ~n397;
  assign n399 = ~n395 & n398;
  assign n400 = n395 & ~n398;
  assign n401 = ~n399 & ~n400;
  assign n402 = n262 & n401;
  assign n403 = pi67  & n288;
  assign n404 = pi69  & n267;
  assign n405 = pi68  & n269;
  assign n406 = ~n404 & ~n405;
  assign n407 = ~n403 & n406;
  assign n408 = ~n402 & n407;
  assign n409 = pi2  & ~n408;
  assign n410 = pi2  & ~n409;
  assign n411 = ~n408 & ~n409;
  assign n412 = ~n410 & ~n411;
  assign n413 = n394 & ~n412;
  assign n414 = n394 & ~n413;
  assign n415 = ~n412 & ~n413;
  assign n416 = ~n414 & ~n415;
  assign n417 = ~n371 & ~n376;
  assign n418 = ~n416 & ~n417;
  assign n419 = n416 & n417;
  assign po5  = ~n418 & ~n419;
  assign n421 = ~n413 & ~n418;
  assign n422 = pi5  & ~pi6 ;
  assign n423 = ~pi5  & pi6 ;
  assign n424 = ~n422 & ~n423;
  assign n425 = pi64  & ~n424;
  assign n426 = n392 & n425;
  assign n427 = n392 & ~n426;
  assign n428 = n425 & ~n426;
  assign n429 = ~n427 & ~n428;
  assign n430 = n309 & n342;
  assign n431 = pi65  & n380;
  assign n432 = pi67  & n340;
  assign n433 = pi66  & n335;
  assign n434 = ~n432 & ~n433;
  assign n435 = ~n431 & n434;
  assign n436 = ~n430 & n435;
  assign n437 = pi5  & ~n436;
  assign n438 = pi5  & ~n437;
  assign n439 = ~n436 & ~n437;
  assign n440 = ~n438 & ~n439;
  assign n441 = ~n429 & n440;
  assign n442 = n429 & ~n440;
  assign n443 = ~n441 & ~n442;
  assign n444 = ~n397 & ~n399;
  assign n445 = ~pi69  & ~pi70 ;
  assign n446 = pi69  & pi70 ;
  assign n447 = ~n445 & ~n446;
  assign n448 = ~n444 & n447;
  assign n449 = n444 & ~n447;
  assign n450 = ~n448 & ~n449;
  assign n451 = n262 & n450;
  assign n452 = pi68  & n288;
  assign n453 = pi70  & n267;
  assign n454 = pi69  & n269;
  assign n455 = ~n453 & ~n454;
  assign n456 = ~n452 & n455;
  assign n457 = ~n451 & n456;
  assign n458 = pi2  & ~n457;
  assign n459 = pi2  & ~n458;
  assign n460 = ~n457 & ~n458;
  assign n461 = ~n459 & ~n460;
  assign n462 = ~n443 & ~n461;
  assign n463 = n443 & n461;
  assign n464 = ~n462 & ~n463;
  assign n465 = ~n421 & n464;
  assign n466 = n421 & ~n464;
  assign po6  = ~n465 & ~n466;
  assign n468 = ~n462 & ~n465;
  assign n469 = ~n446 & ~n448;
  assign n470 = ~pi70  & ~pi71 ;
  assign n471 = pi70  & pi71 ;
  assign n472 = ~n470 & ~n471;
  assign n473 = ~n469 & n472;
  assign n474 = n469 & ~n472;
  assign n475 = ~n473 & ~n474;
  assign n476 = n262 & n475;
  assign n477 = pi69  & n288;
  assign n478 = pi71  & n267;
  assign n479 = pi70  & n269;
  assign n480 = ~n478 & ~n479;
  assign n481 = ~n477 & n480;
  assign n482 = ~n476 & n481;
  assign n483 = pi2  & ~n482;
  assign n484 = pi2  & ~n483;
  assign n485 = ~n482 & ~n483;
  assign n486 = ~n484 & ~n485;
  assign n487 = pi8  & ~n425;
  assign n488 = ~pi6  & pi7 ;
  assign n489 = pi6  & ~pi7 ;
  assign n490 = ~n488 & ~n489;
  assign n491 = n424 & ~n490;
  assign n492 = pi64  & n491;
  assign n493 = ~pi7  & pi8 ;
  assign n494 = pi7  & ~pi8 ;
  assign n495 = ~n493 & ~n494;
  assign n496 = ~n424 & n495;
  assign n497 = pi65  & n496;
  assign n498 = ~n424 & ~n495;
  assign n499 = ~n265 & n498;
  assign n500 = ~n492 & ~n497;
  assign n501 = ~n499 & n500;
  assign n502 = pi8  & ~n501;
  assign n503 = pi8  & ~n502;
  assign n504 = ~n501 & ~n502;
  assign n505 = ~n503 & ~n504;
  assign n506 = n487 & ~n505;
  assign n507 = ~n487 & n505;
  assign n508 = ~n506 & ~n507;
  assign n509 = n342 & n359;
  assign n510 = pi66  & n380;
  assign n511 = pi68  & n340;
  assign n512 = pi67  & n335;
  assign n513 = ~n511 & ~n512;
  assign n514 = ~n510 & n513;
  assign n515 = ~n509 & n514;
  assign n516 = pi5  & ~n515;
  assign n517 = pi5  & ~n516;
  assign n518 = ~n515 & ~n516;
  assign n519 = ~n517 & ~n518;
  assign n520 = n508 & ~n519;
  assign n521 = n508 & ~n520;
  assign n522 = ~n519 & ~n520;
  assign n523 = ~n521 & ~n522;
  assign n524 = ~n429 & ~n440;
  assign n525 = ~n426 & ~n524;
  assign n526 = ~n523 & ~n525;
  assign n527 = n523 & n525;
  assign n528 = ~n526 & ~n527;
  assign n529 = ~n486 & n528;
  assign n530 = n486 & ~n528;
  assign n531 = ~n529 & ~n530;
  assign n532 = ~n468 & n531;
  assign n533 = n468 & ~n531;
  assign po7  = ~n532 & ~n533;
  assign n535 = n286 & n498;
  assign n536 = n424 & n490;
  assign n537 = ~n495 & n536;
  assign n538 = pi64  & n537;
  assign n539 = pi66  & n496;
  assign n540 = pi65  & n491;
  assign n541 = ~n539 & ~n540;
  assign n542 = ~n535 & n541;
  assign n543 = ~n538 & n542;
  assign n544 = pi8  & ~n543;
  assign n545 = pi8  & ~n544;
  assign n546 = ~n543 & ~n544;
  assign n547 = ~n545 & ~n546;
  assign n548 = ~n506 & n547;
  assign n549 = n506 & ~n547;
  assign n550 = ~n548 & ~n549;
  assign n551 = n342 & n401;
  assign n552 = pi67  & n380;
  assign n553 = pi69  & n340;
  assign n554 = pi68  & n335;
  assign n555 = ~n553 & ~n554;
  assign n556 = ~n552 & n555;
  assign n557 = ~n551 & n556;
  assign n558 = pi5  & ~n557;
  assign n559 = pi5  & ~n558;
  assign n560 = ~n557 & ~n558;
  assign n561 = ~n559 & ~n560;
  assign n562 = n550 & ~n561;
  assign n563 = n550 & ~n562;
  assign n564 = ~n561 & ~n562;
  assign n565 = ~n563 & ~n564;
  assign n566 = ~n520 & ~n526;
  assign n567 = n565 & n566;
  assign n568 = ~n565 & ~n566;
  assign n569 = ~n567 & ~n568;
  assign n570 = ~n471 & ~n473;
  assign n571 = ~pi71  & ~pi72 ;
  assign n572 = pi71  & pi72 ;
  assign n573 = ~n571 & ~n572;
  assign n574 = ~n570 & n573;
  assign n575 = n570 & ~n573;
  assign n576 = ~n574 & ~n575;
  assign n577 = n262 & n576;
  assign n578 = pi70  & n288;
  assign n579 = pi72  & n267;
  assign n580 = pi71  & n269;
  assign n581 = ~n579 & ~n580;
  assign n582 = ~n578 & n581;
  assign n583 = ~n577 & n582;
  assign n584 = pi2  & ~n583;
  assign n585 = pi2  & ~n584;
  assign n586 = ~n583 & ~n584;
  assign n587 = ~n585 & ~n586;
  assign n588 = n569 & ~n587;
  assign n589 = n569 & ~n588;
  assign n590 = ~n587 & ~n588;
  assign n591 = ~n589 & ~n590;
  assign n592 = ~n529 & ~n532;
  assign n593 = ~n591 & ~n592;
  assign n594 = n591 & n592;
  assign po8  = ~n593 & ~n594;
  assign n596 = pi8  & ~pi9 ;
  assign n597 = ~pi8  & pi9 ;
  assign n598 = ~n596 & ~n597;
  assign n599 = pi64  & ~n598;
  assign n600 = ~n549 & n599;
  assign n601 = n549 & ~n599;
  assign n602 = ~n600 & ~n601;
  assign n603 = n309 & n498;
  assign n604 = pi65  & n537;
  assign n605 = pi67  & n496;
  assign n606 = pi66  & n491;
  assign n607 = ~n605 & ~n606;
  assign n608 = ~n604 & n607;
  assign n609 = ~n603 & n608;
  assign n610 = pi8  & ~n609;
  assign n611 = pi8  & ~n610;
  assign n612 = ~n609 & ~n610;
  assign n613 = ~n611 & ~n612;
  assign n614 = ~n602 & ~n613;
  assign n615 = n602 & n613;
  assign n616 = ~n614 & ~n615;
  assign n617 = n342 & n450;
  assign n618 = pi68  & n380;
  assign n619 = pi70  & n340;
  assign n620 = pi69  & n335;
  assign n621 = ~n619 & ~n620;
  assign n622 = ~n618 & n621;
  assign n623 = ~n617 & n622;
  assign n624 = pi5  & ~n623;
  assign n625 = pi5  & ~n624;
  assign n626 = ~n623 & ~n624;
  assign n627 = ~n625 & ~n626;
  assign n628 = n616 & ~n627;
  assign n629 = n616 & ~n628;
  assign n630 = ~n627 & ~n628;
  assign n631 = ~n629 & ~n630;
  assign n632 = ~n562 & ~n568;
  assign n633 = n631 & n632;
  assign n634 = ~n631 & ~n632;
  assign n635 = ~n633 & ~n634;
  assign n636 = ~n572 & ~n574;
  assign n637 = ~pi72  & ~pi73 ;
  assign n638 = pi72  & pi73 ;
  assign n639 = ~n637 & ~n638;
  assign n640 = ~n636 & n639;
  assign n641 = n636 & ~n639;
  assign n642 = ~n640 & ~n641;
  assign n643 = n262 & n642;
  assign n644 = pi71  & n288;
  assign n645 = pi73  & n267;
  assign n646 = pi72  & n269;
  assign n647 = ~n645 & ~n646;
  assign n648 = ~n644 & n647;
  assign n649 = ~n643 & n648;
  assign n650 = pi2  & ~n649;
  assign n651 = pi2  & ~n650;
  assign n652 = ~n649 & ~n650;
  assign n653 = ~n651 & ~n652;
  assign n654 = n635 & ~n653;
  assign n655 = n635 & ~n654;
  assign n656 = ~n653 & ~n654;
  assign n657 = ~n655 & ~n656;
  assign n658 = ~n588 & ~n593;
  assign n659 = ~n657 & ~n658;
  assign n660 = n657 & n658;
  assign po9  = ~n659 & ~n660;
  assign n662 = ~n654 & ~n659;
  assign n663 = n549 & n599;
  assign n664 = ~n614 & ~n663;
  assign n665 = n359 & n498;
  assign n666 = pi66  & n537;
  assign n667 = pi68  & n496;
  assign n668 = pi67  & n491;
  assign n669 = ~n667 & ~n668;
  assign n670 = ~n666 & n669;
  assign n671 = ~n665 & n670;
  assign n672 = pi8  & ~n671;
  assign n673 = pi8  & ~n672;
  assign n674 = ~n671 & ~n672;
  assign n675 = ~n673 & ~n674;
  assign n676 = pi11  & ~n599;
  assign n677 = ~pi9  & pi10 ;
  assign n678 = pi9  & ~pi10 ;
  assign n679 = ~n677 & ~n678;
  assign n680 = n598 & ~n679;
  assign n681 = pi64  & n680;
  assign n682 = ~pi10  & pi11 ;
  assign n683 = pi10  & ~pi11 ;
  assign n684 = ~n682 & ~n683;
  assign n685 = ~n598 & n684;
  assign n686 = pi65  & n685;
  assign n687 = ~n598 & ~n684;
  assign n688 = ~n265 & n687;
  assign n689 = ~n681 & ~n686;
  assign n690 = ~n688 & n689;
  assign n691 = pi11  & ~n690;
  assign n692 = pi11  & ~n691;
  assign n693 = ~n690 & ~n691;
  assign n694 = ~n692 & ~n693;
  assign n695 = n676 & ~n694;
  assign n696 = ~n676 & n694;
  assign n697 = ~n695 & ~n696;
  assign n698 = n675 & ~n697;
  assign n699 = ~n675 & n697;
  assign n700 = ~n698 & ~n699;
  assign n701 = ~n664 & n700;
  assign n702 = n664 & ~n700;
  assign n703 = ~n701 & ~n702;
  assign n704 = n342 & n475;
  assign n705 = pi69  & n380;
  assign n706 = pi71  & n340;
  assign n707 = pi70  & n335;
  assign n708 = ~n706 & ~n707;
  assign n709 = ~n705 & n708;
  assign n710 = ~n704 & n709;
  assign n711 = pi5  & ~n710;
  assign n712 = pi5  & ~n711;
  assign n713 = ~n710 & ~n711;
  assign n714 = ~n712 & ~n713;
  assign n715 = n703 & ~n714;
  assign n716 = n703 & ~n715;
  assign n717 = ~n714 & ~n715;
  assign n718 = ~n716 & ~n717;
  assign n719 = ~n628 & ~n634;
  assign n720 = n718 & n719;
  assign n721 = ~n718 & ~n719;
  assign n722 = ~n720 & ~n721;
  assign n723 = ~n638 & ~n640;
  assign n724 = ~pi73  & ~pi74 ;
  assign n725 = pi73  & pi74 ;
  assign n726 = ~n724 & ~n725;
  assign n727 = ~n723 & n726;
  assign n728 = n723 & ~n726;
  assign n729 = ~n727 & ~n728;
  assign n730 = n262 & n729;
  assign n731 = pi72  & n288;
  assign n732 = pi74  & n267;
  assign n733 = pi73  & n269;
  assign n734 = ~n732 & ~n733;
  assign n735 = ~n731 & n734;
  assign n736 = ~n730 & n735;
  assign n737 = pi2  & ~n736;
  assign n738 = pi2  & ~n737;
  assign n739 = ~n736 & ~n737;
  assign n740 = ~n738 & ~n739;
  assign n741 = ~n722 & n740;
  assign n742 = n722 & ~n740;
  assign n743 = ~n741 & ~n742;
  assign n744 = ~n662 & n743;
  assign n745 = n662 & ~n743;
  assign po10  = ~n744 & ~n745;
  assign n747 = ~n742 & ~n744;
  assign n748 = ~n715 & ~n721;
  assign n749 = n342 & n576;
  assign n750 = pi70  & n380;
  assign n751 = pi72  & n340;
  assign n752 = pi71  & n335;
  assign n753 = ~n751 & ~n752;
  assign n754 = ~n750 & n753;
  assign n755 = ~n749 & n754;
  assign n756 = pi5  & ~n755;
  assign n757 = pi5  & ~n756;
  assign n758 = ~n755 & ~n756;
  assign n759 = ~n757 & ~n758;
  assign n760 = ~n699 & ~n701;
  assign n761 = n286 & n687;
  assign n762 = n598 & n679;
  assign n763 = ~n684 & n762;
  assign n764 = pi64  & n763;
  assign n765 = pi66  & n685;
  assign n766 = pi65  & n680;
  assign n767 = ~n765 & ~n766;
  assign n768 = ~n761 & n767;
  assign n769 = ~n764 & n768;
  assign n770 = pi11  & ~n769;
  assign n771 = pi11  & ~n770;
  assign n772 = ~n769 & ~n770;
  assign n773 = ~n771 & ~n772;
  assign n774 = ~n695 & n773;
  assign n775 = n695 & ~n773;
  assign n776 = ~n774 & ~n775;
  assign n777 = n401 & n498;
  assign n778 = pi67  & n537;
  assign n779 = pi69  & n496;
  assign n780 = pi68  & n491;
  assign n781 = ~n779 & ~n780;
  assign n782 = ~n778 & n781;
  assign n783 = ~n777 & n782;
  assign n784 = pi8  & ~n783;
  assign n785 = pi8  & ~n784;
  assign n786 = ~n783 & ~n784;
  assign n787 = ~n785 & ~n786;
  assign n788 = n776 & ~n787;
  assign n789 = n776 & ~n788;
  assign n790 = ~n787 & ~n788;
  assign n791 = ~n789 & ~n790;
  assign n792 = ~n760 & ~n791;
  assign n793 = n760 & n791;
  assign n794 = ~n792 & ~n793;
  assign n795 = ~n759 & n794;
  assign n796 = ~n759 & ~n795;
  assign n797 = n794 & ~n795;
  assign n798 = ~n796 & ~n797;
  assign n799 = ~n748 & ~n798;
  assign n800 = ~n748 & ~n799;
  assign n801 = ~n798 & ~n799;
  assign n802 = ~n800 & ~n801;
  assign n803 = ~n725 & ~n727;
  assign n804 = ~pi74  & ~pi75 ;
  assign n805 = pi74  & pi75 ;
  assign n806 = ~n804 & ~n805;
  assign n807 = ~n803 & n806;
  assign n808 = n803 & ~n806;
  assign n809 = ~n807 & ~n808;
  assign n810 = n262 & n809;
  assign n811 = pi73  & n288;
  assign n812 = pi75  & n267;
  assign n813 = pi74  & n269;
  assign n814 = ~n812 & ~n813;
  assign n815 = ~n811 & n814;
  assign n816 = ~n810 & n815;
  assign n817 = pi2  & ~n816;
  assign n818 = pi2  & ~n817;
  assign n819 = ~n816 & ~n817;
  assign n820 = ~n818 & ~n819;
  assign n821 = ~n802 & n820;
  assign n822 = n802 & ~n820;
  assign n823 = ~n821 & ~n822;
  assign n824 = ~n747 & ~n823;
  assign n825 = n747 & n823;
  assign po11  = ~n824 & ~n825;
  assign n827 = pi11  & ~pi12 ;
  assign n828 = ~pi11  & pi12 ;
  assign n829 = ~n827 & ~n828;
  assign n830 = pi64  & ~n829;
  assign n831 = ~n775 & n830;
  assign n832 = n775 & ~n830;
  assign n833 = ~n831 & ~n832;
  assign n834 = n309 & n687;
  assign n835 = pi65  & n763;
  assign n836 = pi67  & n685;
  assign n837 = pi66  & n680;
  assign n838 = ~n836 & ~n837;
  assign n839 = ~n835 & n838;
  assign n840 = ~n834 & n839;
  assign n841 = pi11  & ~n840;
  assign n842 = pi11  & ~n841;
  assign n843 = ~n840 & ~n841;
  assign n844 = ~n842 & ~n843;
  assign n845 = ~n833 & ~n844;
  assign n846 = n833 & n844;
  assign n847 = ~n845 & ~n846;
  assign n848 = n450 & n498;
  assign n849 = pi68  & n537;
  assign n850 = pi70  & n496;
  assign n851 = pi69  & n491;
  assign n852 = ~n850 & ~n851;
  assign n853 = ~n849 & n852;
  assign n854 = ~n848 & n853;
  assign n855 = pi8  & ~n854;
  assign n856 = pi8  & ~n855;
  assign n857 = ~n854 & ~n855;
  assign n858 = ~n856 & ~n857;
  assign n859 = n847 & ~n858;
  assign n860 = n847 & ~n859;
  assign n861 = ~n858 & ~n859;
  assign n862 = ~n860 & ~n861;
  assign n863 = ~n788 & ~n792;
  assign n864 = n862 & n863;
  assign n865 = ~n862 & ~n863;
  assign n866 = ~n864 & ~n865;
  assign n867 = n342 & n642;
  assign n868 = pi71  & n380;
  assign n869 = pi73  & n340;
  assign n870 = pi72  & n335;
  assign n871 = ~n869 & ~n870;
  assign n872 = ~n868 & n871;
  assign n873 = ~n867 & n872;
  assign n874 = pi5  & ~n873;
  assign n875 = pi5  & ~n874;
  assign n876 = ~n873 & ~n874;
  assign n877 = ~n875 & ~n876;
  assign n878 = ~n866 & n877;
  assign n879 = n866 & ~n877;
  assign n880 = ~n878 & ~n879;
  assign n881 = ~n795 & ~n799;
  assign n882 = n880 & ~n881;
  assign n883 = ~n880 & n881;
  assign n884 = ~n882 & ~n883;
  assign n885 = ~n805 & ~n807;
  assign n886 = ~pi75  & ~pi76 ;
  assign n887 = pi75  & pi76 ;
  assign n888 = ~n886 & ~n887;
  assign n889 = ~n885 & n888;
  assign n890 = n885 & ~n888;
  assign n891 = ~n889 & ~n890;
  assign n892 = n262 & n891;
  assign n893 = pi74  & n288;
  assign n894 = pi76  & n267;
  assign n895 = pi75  & n269;
  assign n896 = ~n894 & ~n895;
  assign n897 = ~n893 & n896;
  assign n898 = ~n892 & n897;
  assign n899 = pi2  & ~n898;
  assign n900 = pi2  & ~n899;
  assign n901 = ~n898 & ~n899;
  assign n902 = ~n900 & ~n901;
  assign n903 = n884 & ~n902;
  assign n904 = n884 & ~n903;
  assign n905 = ~n902 & ~n903;
  assign n906 = ~n904 & ~n905;
  assign n907 = ~n802 & ~n820;
  assign n908 = ~n824 & ~n907;
  assign n909 = ~n906 & ~n908;
  assign n910 = n906 & n908;
  assign po12  = ~n909 & ~n910;
  assign n912 = ~n903 & ~n909;
  assign n913 = ~n879 & ~n882;
  assign n914 = n775 & n830;
  assign n915 = ~n845 & ~n914;
  assign n916 = n359 & n687;
  assign n917 = pi66  & n763;
  assign n918 = pi68  & n685;
  assign n919 = pi67  & n680;
  assign n920 = ~n918 & ~n919;
  assign n921 = ~n917 & n920;
  assign n922 = ~n916 & n921;
  assign n923 = pi11  & ~n922;
  assign n924 = pi11  & ~n923;
  assign n925 = ~n922 & ~n923;
  assign n926 = ~n924 & ~n925;
  assign n927 = pi14  & ~n830;
  assign n928 = ~pi12  & pi13 ;
  assign n929 = pi12  & ~pi13 ;
  assign n930 = ~n928 & ~n929;
  assign n931 = n829 & ~n930;
  assign n932 = pi64  & n931;
  assign n933 = ~pi13  & pi14 ;
  assign n934 = pi13  & ~pi14 ;
  assign n935 = ~n933 & ~n934;
  assign n936 = ~n829 & n935;
  assign n937 = pi65  & n936;
  assign n938 = ~n829 & ~n935;
  assign n939 = ~n265 & n938;
  assign n940 = ~n932 & ~n937;
  assign n941 = ~n939 & n940;
  assign n942 = pi14  & ~n941;
  assign n943 = pi14  & ~n942;
  assign n944 = ~n941 & ~n942;
  assign n945 = ~n943 & ~n944;
  assign n946 = n927 & ~n945;
  assign n947 = ~n927 & n945;
  assign n948 = ~n946 & ~n947;
  assign n949 = n926 & ~n948;
  assign n950 = ~n926 & n948;
  assign n951 = ~n949 & ~n950;
  assign n952 = ~n915 & n951;
  assign n953 = n915 & ~n951;
  assign n954 = ~n952 & ~n953;
  assign n955 = n475 & n498;
  assign n956 = pi69  & n537;
  assign n957 = pi71  & n496;
  assign n958 = pi70  & n491;
  assign n959 = ~n957 & ~n958;
  assign n960 = ~n956 & n959;
  assign n961 = ~n955 & n960;
  assign n962 = pi8  & ~n961;
  assign n963 = pi8  & ~n962;
  assign n964 = ~n961 & ~n962;
  assign n965 = ~n963 & ~n964;
  assign n966 = n954 & ~n965;
  assign n967 = n954 & ~n966;
  assign n968 = ~n965 & ~n966;
  assign n969 = ~n967 & ~n968;
  assign n970 = ~n859 & ~n865;
  assign n971 = n969 & n970;
  assign n972 = ~n969 & ~n970;
  assign n973 = ~n971 & ~n972;
  assign n974 = n342 & n729;
  assign n975 = pi72  & n380;
  assign n976 = pi74  & n340;
  assign n977 = pi73  & n335;
  assign n978 = ~n976 & ~n977;
  assign n979 = ~n975 & n978;
  assign n980 = ~n974 & n979;
  assign n981 = pi5  & ~n980;
  assign n982 = pi5  & ~n981;
  assign n983 = ~n980 & ~n981;
  assign n984 = ~n982 & ~n983;
  assign n985 = n973 & ~n984;
  assign n986 = ~n973 & n984;
  assign n987 = ~n985 & ~n986;
  assign n988 = ~n913 & n987;
  assign n989 = ~n913 & ~n988;
  assign n990 = ~n985 & ~n988;
  assign n991 = ~n986 & n990;
  assign n992 = ~n989 & ~n991;
  assign n993 = ~n887 & ~n889;
  assign n994 = ~pi76  & ~pi77 ;
  assign n995 = pi76  & pi77 ;
  assign n996 = ~n994 & ~n995;
  assign n997 = ~n993 & n996;
  assign n998 = n993 & ~n996;
  assign n999 = ~n997 & ~n998;
  assign n1000 = n262 & n999;
  assign n1001 = pi75  & n288;
  assign n1002 = pi77  & n267;
  assign n1003 = pi76  & n269;
  assign n1004 = ~n1002 & ~n1003;
  assign n1005 = ~n1001 & n1004;
  assign n1006 = ~n1000 & n1005;
  assign n1007 = pi2  & ~n1006;
  assign n1008 = pi2  & ~n1007;
  assign n1009 = ~n1006 & ~n1007;
  assign n1010 = ~n1008 & ~n1009;
  assign n1011 = ~n992 & n1010;
  assign n1012 = n992 & ~n1010;
  assign n1013 = ~n1011 & ~n1012;
  assign n1014 = ~n912 & ~n1013;
  assign n1015 = n912 & n1013;
  assign po13  = ~n1014 & ~n1015;
  assign n1017 = ~n992 & ~n1010;
  assign n1018 = ~n1014 & ~n1017;
  assign n1019 = ~n995 & ~n997;
  assign n1020 = ~pi77  & ~pi78 ;
  assign n1021 = pi77  & pi78 ;
  assign n1022 = ~n1020 & ~n1021;
  assign n1023 = ~n1019 & n1022;
  assign n1024 = n1019 & ~n1022;
  assign n1025 = ~n1023 & ~n1024;
  assign n1026 = n262 & n1025;
  assign n1027 = pi76  & n288;
  assign n1028 = pi78  & n267;
  assign n1029 = pi77  & n269;
  assign n1030 = ~n1028 & ~n1029;
  assign n1031 = ~n1027 & n1030;
  assign n1032 = ~n1026 & n1031;
  assign n1033 = pi2  & ~n1032;
  assign n1034 = pi2  & ~n1033;
  assign n1035 = ~n1032 & ~n1033;
  assign n1036 = ~n1034 & ~n1035;
  assign n1037 = n342 & n809;
  assign n1038 = pi73  & n380;
  assign n1039 = pi75  & n340;
  assign n1040 = pi74  & n335;
  assign n1041 = ~n1039 & ~n1040;
  assign n1042 = ~n1038 & n1041;
  assign n1043 = ~n1037 & n1042;
  assign n1044 = pi5  & ~n1043;
  assign n1045 = pi5  & ~n1044;
  assign n1046 = ~n1043 & ~n1044;
  assign n1047 = ~n1045 & ~n1046;
  assign n1048 = ~n966 & ~n972;
  assign n1049 = ~n950 & ~n952;
  assign n1050 = n286 & n938;
  assign n1051 = n829 & n930;
  assign n1052 = ~n935 & n1051;
  assign n1053 = pi64  & n1052;
  assign n1054 = pi66  & n936;
  assign n1055 = pi65  & n931;
  assign n1056 = ~n1054 & ~n1055;
  assign n1057 = ~n1050 & n1056;
  assign n1058 = ~n1053 & n1057;
  assign n1059 = pi14  & ~n1058;
  assign n1060 = pi14  & ~n1059;
  assign n1061 = ~n1058 & ~n1059;
  assign n1062 = ~n1060 & ~n1061;
  assign n1063 = ~n946 & n1062;
  assign n1064 = n946 & ~n1062;
  assign n1065 = ~n1063 & ~n1064;
  assign n1066 = n401 & n687;
  assign n1067 = pi67  & n763;
  assign n1068 = pi69  & n685;
  assign n1069 = pi68  & n680;
  assign n1070 = ~n1068 & ~n1069;
  assign n1071 = ~n1067 & n1070;
  assign n1072 = ~n1066 & n1071;
  assign n1073 = pi11  & ~n1072;
  assign n1074 = pi11  & ~n1073;
  assign n1075 = ~n1072 & ~n1073;
  assign n1076 = ~n1074 & ~n1075;
  assign n1077 = n1065 & ~n1076;
  assign n1078 = ~n1065 & n1076;
  assign n1079 = ~n1077 & ~n1078;
  assign n1080 = ~n1049 & n1079;
  assign n1081 = ~n1049 & ~n1080;
  assign n1082 = ~n1077 & ~n1080;
  assign n1083 = ~n1078 & n1082;
  assign n1084 = ~n1081 & ~n1083;
  assign n1085 = n498 & n576;
  assign n1086 = pi70  & n537;
  assign n1087 = pi72  & n496;
  assign n1088 = pi71  & n491;
  assign n1089 = ~n1087 & ~n1088;
  assign n1090 = ~n1086 & n1089;
  assign n1091 = ~n1085 & n1090;
  assign n1092 = pi8  & ~n1091;
  assign n1093 = pi8  & ~n1092;
  assign n1094 = ~n1091 & ~n1092;
  assign n1095 = ~n1093 & ~n1094;
  assign n1096 = n1084 & n1095;
  assign n1097 = ~n1084 & ~n1095;
  assign n1098 = ~n1096 & ~n1097;
  assign n1099 = ~n1048 & n1098;
  assign n1100 = n1048 & ~n1098;
  assign n1101 = ~n1099 & ~n1100;
  assign n1102 = n1047 & ~n1101;
  assign n1103 = ~n1047 & n1101;
  assign n1104 = ~n1102 & ~n1103;
  assign n1105 = ~n990 & n1104;
  assign n1106 = n990 & ~n1104;
  assign n1107 = ~n1105 & ~n1106;
  assign n1108 = n1036 & n1107;
  assign n1109 = ~n1036 & ~n1107;
  assign n1110 = ~n1108 & ~n1109;
  assign n1111 = ~n1018 & ~n1110;
  assign n1112 = n1018 & n1110;
  assign po14  = ~n1111 & ~n1112;
  assign n1114 = ~n1036 & n1107;
  assign n1115 = ~n1111 & ~n1114;
  assign n1116 = ~n1021 & ~n1023;
  assign n1117 = ~pi78  & ~pi79 ;
  assign n1118 = pi78  & pi79 ;
  assign n1119 = ~n1117 & ~n1118;
  assign n1120 = ~n1116 & n1119;
  assign n1121 = n1116 & ~n1119;
  assign n1122 = ~n1120 & ~n1121;
  assign n1123 = n262 & n1122;
  assign n1124 = pi77  & n288;
  assign n1125 = pi79  & n267;
  assign n1126 = pi78  & n269;
  assign n1127 = ~n1125 & ~n1126;
  assign n1128 = ~n1124 & n1127;
  assign n1129 = ~n1123 & n1128;
  assign n1130 = pi2  & ~n1129;
  assign n1131 = pi2  & ~n1130;
  assign n1132 = ~n1129 & ~n1130;
  assign n1133 = ~n1131 & ~n1132;
  assign n1134 = ~n1103 & ~n1105;
  assign n1135 = n342 & n891;
  assign n1136 = pi74  & n380;
  assign n1137 = pi76  & n340;
  assign n1138 = pi75  & n335;
  assign n1139 = ~n1137 & ~n1138;
  assign n1140 = ~n1136 & n1139;
  assign n1141 = ~n1135 & n1140;
  assign n1142 = pi5  & ~n1141;
  assign n1143 = pi5  & ~n1142;
  assign n1144 = ~n1141 & ~n1142;
  assign n1145 = ~n1143 & ~n1144;
  assign n1146 = ~n1097 & ~n1099;
  assign n1147 = n498 & n642;
  assign n1148 = pi71  & n537;
  assign n1149 = pi73  & n496;
  assign n1150 = pi72  & n491;
  assign n1151 = ~n1149 & ~n1150;
  assign n1152 = ~n1148 & n1151;
  assign n1153 = ~n1147 & n1152;
  assign n1154 = pi8  & ~n1153;
  assign n1155 = pi8  & ~n1154;
  assign n1156 = ~n1153 & ~n1154;
  assign n1157 = ~n1155 & ~n1156;
  assign n1158 = pi14  & ~pi15 ;
  assign n1159 = ~pi14  & pi15 ;
  assign n1160 = ~n1158 & ~n1159;
  assign n1161 = pi64  & ~n1160;
  assign n1162 = ~n1064 & n1161;
  assign n1163 = n1064 & ~n1161;
  assign n1164 = ~n1162 & ~n1163;
  assign n1165 = n309 & n938;
  assign n1166 = pi65  & n1052;
  assign n1167 = pi67  & n936;
  assign n1168 = pi66  & n931;
  assign n1169 = ~n1167 & ~n1168;
  assign n1170 = ~n1166 & n1169;
  assign n1171 = ~n1165 & n1170;
  assign n1172 = pi14  & ~n1171;
  assign n1173 = pi14  & ~n1172;
  assign n1174 = ~n1171 & ~n1172;
  assign n1175 = ~n1173 & ~n1174;
  assign n1176 = ~n1164 & ~n1175;
  assign n1177 = n1164 & n1175;
  assign n1178 = ~n1176 & ~n1177;
  assign n1179 = n450 & n687;
  assign n1180 = pi68  & n763;
  assign n1181 = pi70  & n685;
  assign n1182 = pi69  & n680;
  assign n1183 = ~n1181 & ~n1182;
  assign n1184 = ~n1180 & n1183;
  assign n1185 = ~n1179 & n1184;
  assign n1186 = pi11  & ~n1185;
  assign n1187 = pi11  & ~n1186;
  assign n1188 = ~n1185 & ~n1186;
  assign n1189 = ~n1187 & ~n1188;
  assign n1190 = n1178 & ~n1189;
  assign n1191 = n1178 & ~n1190;
  assign n1192 = ~n1189 & ~n1190;
  assign n1193 = ~n1191 & ~n1192;
  assign n1194 = ~n1082 & ~n1193;
  assign n1195 = n1082 & n1193;
  assign n1196 = ~n1194 & ~n1195;
  assign n1197 = ~n1157 & n1196;
  assign n1198 = ~n1157 & ~n1197;
  assign n1199 = n1196 & ~n1197;
  assign n1200 = ~n1198 & ~n1199;
  assign n1201 = ~n1146 & ~n1200;
  assign n1202 = n1146 & n1200;
  assign n1203 = ~n1201 & ~n1202;
  assign n1204 = ~n1145 & n1203;
  assign n1205 = ~n1145 & ~n1204;
  assign n1206 = n1203 & ~n1204;
  assign n1207 = ~n1205 & ~n1206;
  assign n1208 = ~n1134 & ~n1207;
  assign n1209 = n1134 & n1207;
  assign n1210 = ~n1208 & ~n1209;
  assign n1211 = ~n1133 & n1210;
  assign n1212 = ~n1133 & ~n1211;
  assign n1213 = n1210 & ~n1211;
  assign n1214 = ~n1212 & ~n1213;
  assign n1215 = ~n1115 & ~n1214;
  assign n1216 = n1115 & n1214;
  assign po15  = ~n1215 & ~n1216;
  assign n1218 = ~n1211 & ~n1215;
  assign n1219 = ~n1118 & ~n1120;
  assign n1220 = ~pi79  & ~pi80 ;
  assign n1221 = pi79  & pi80 ;
  assign n1222 = ~n1220 & ~n1221;
  assign n1223 = ~n1219 & n1222;
  assign n1224 = n1219 & ~n1222;
  assign n1225 = ~n1223 & ~n1224;
  assign n1226 = n262 & n1225;
  assign n1227 = pi78  & n288;
  assign n1228 = pi80  & n267;
  assign n1229 = pi79  & n269;
  assign n1230 = ~n1228 & ~n1229;
  assign n1231 = ~n1227 & n1230;
  assign n1232 = ~n1226 & n1231;
  assign n1233 = pi2  & ~n1232;
  assign n1234 = pi2  & ~n1233;
  assign n1235 = ~n1232 & ~n1233;
  assign n1236 = ~n1234 & ~n1235;
  assign n1237 = ~n1204 & ~n1208;
  assign n1238 = n342 & n999;
  assign n1239 = pi75  & n380;
  assign n1240 = pi77  & n340;
  assign n1241 = pi76  & n335;
  assign n1242 = ~n1240 & ~n1241;
  assign n1243 = ~n1239 & n1242;
  assign n1244 = ~n1238 & n1243;
  assign n1245 = pi5  & ~n1244;
  assign n1246 = pi5  & ~n1245;
  assign n1247 = ~n1244 & ~n1245;
  assign n1248 = ~n1246 & ~n1247;
  assign n1249 = ~n1197 & ~n1201;
  assign n1250 = n498 & n729;
  assign n1251 = pi72  & n537;
  assign n1252 = pi74  & n496;
  assign n1253 = pi73  & n491;
  assign n1254 = ~n1252 & ~n1253;
  assign n1255 = ~n1251 & n1254;
  assign n1256 = ~n1250 & n1255;
  assign n1257 = pi8  & ~n1256;
  assign n1258 = pi8  & ~n1257;
  assign n1259 = ~n1256 & ~n1257;
  assign n1260 = ~n1258 & ~n1259;
  assign n1261 = ~n1190 & ~n1194;
  assign n1262 = n475 & n687;
  assign n1263 = pi69  & n763;
  assign n1264 = pi71  & n685;
  assign n1265 = pi70  & n680;
  assign n1266 = ~n1264 & ~n1265;
  assign n1267 = ~n1263 & n1266;
  assign n1268 = ~n1262 & n1267;
  assign n1269 = pi11  & ~n1268;
  assign n1270 = pi11  & ~n1269;
  assign n1271 = ~n1268 & ~n1269;
  assign n1272 = ~n1270 & ~n1271;
  assign n1273 = n1064 & n1161;
  assign n1274 = ~n1176 & ~n1273;
  assign n1275 = n359 & n938;
  assign n1276 = pi66  & n1052;
  assign n1277 = pi68  & n936;
  assign n1278 = pi67  & n931;
  assign n1279 = ~n1277 & ~n1278;
  assign n1280 = ~n1276 & n1279;
  assign n1281 = ~n1275 & n1280;
  assign n1282 = pi14  & ~n1281;
  assign n1283 = pi14  & ~n1282;
  assign n1284 = ~n1281 & ~n1282;
  assign n1285 = ~n1283 & ~n1284;
  assign n1286 = pi17  & ~n1161;
  assign n1287 = ~pi15  & pi16 ;
  assign n1288 = pi15  & ~pi16 ;
  assign n1289 = ~n1287 & ~n1288;
  assign n1290 = n1160 & ~n1289;
  assign n1291 = pi64  & n1290;
  assign n1292 = ~pi16  & pi17 ;
  assign n1293 = pi16  & ~pi17 ;
  assign n1294 = ~n1292 & ~n1293;
  assign n1295 = ~n1160 & n1294;
  assign n1296 = pi65  & n1295;
  assign n1297 = ~n1160 & ~n1294;
  assign n1298 = ~n265 & n1297;
  assign n1299 = ~n1291 & ~n1296;
  assign n1300 = ~n1298 & n1299;
  assign n1301 = pi17  & ~n1300;
  assign n1302 = pi17  & ~n1301;
  assign n1303 = ~n1300 & ~n1301;
  assign n1304 = ~n1302 & ~n1303;
  assign n1305 = n1286 & ~n1304;
  assign n1306 = ~n1286 & n1304;
  assign n1307 = ~n1305 & ~n1306;
  assign n1308 = n1285 & ~n1307;
  assign n1309 = ~n1285 & n1307;
  assign n1310 = ~n1308 & ~n1309;
  assign n1311 = ~n1274 & n1310;
  assign n1312 = n1274 & ~n1310;
  assign n1313 = ~n1311 & ~n1312;
  assign n1314 = n1272 & ~n1313;
  assign n1315 = ~n1272 & n1313;
  assign n1316 = ~n1314 & ~n1315;
  assign n1317 = ~n1261 & n1316;
  assign n1318 = n1261 & ~n1316;
  assign n1319 = ~n1317 & ~n1318;
  assign n1320 = n1260 & ~n1319;
  assign n1321 = ~n1260 & n1319;
  assign n1322 = ~n1320 & ~n1321;
  assign n1323 = ~n1249 & n1322;
  assign n1324 = n1249 & ~n1322;
  assign n1325 = ~n1323 & ~n1324;
  assign n1326 = n1248 & ~n1325;
  assign n1327 = ~n1248 & n1325;
  assign n1328 = ~n1326 & ~n1327;
  assign n1329 = ~n1237 & n1328;
  assign n1330 = n1237 & ~n1328;
  assign n1331 = ~n1329 & ~n1330;
  assign n1332 = n1236 & n1331;
  assign n1333 = ~n1236 & ~n1331;
  assign n1334 = ~n1332 & ~n1333;
  assign n1335 = ~n1218 & ~n1334;
  assign n1336 = n1218 & n1334;
  assign po16  = ~n1335 & ~n1336;
  assign n1338 = ~n1327 & ~n1329;
  assign n1339 = n342 & n1025;
  assign n1340 = pi76  & n380;
  assign n1341 = pi78  & n340;
  assign n1342 = pi77  & n335;
  assign n1343 = ~n1341 & ~n1342;
  assign n1344 = ~n1340 & n1343;
  assign n1345 = ~n1339 & n1344;
  assign n1346 = pi5  & ~n1345;
  assign n1347 = pi5  & ~n1346;
  assign n1348 = ~n1345 & ~n1346;
  assign n1349 = ~n1347 & ~n1348;
  assign n1350 = ~n1321 & ~n1323;
  assign n1351 = n498 & n809;
  assign n1352 = pi73  & n537;
  assign n1353 = pi75  & n496;
  assign n1354 = pi74  & n491;
  assign n1355 = ~n1353 & ~n1354;
  assign n1356 = ~n1352 & n1355;
  assign n1357 = ~n1351 & n1356;
  assign n1358 = pi8  & ~n1357;
  assign n1359 = pi8  & ~n1358;
  assign n1360 = ~n1357 & ~n1358;
  assign n1361 = ~n1359 & ~n1360;
  assign n1362 = ~n1315 & ~n1317;
  assign n1363 = ~n1309 & ~n1311;
  assign n1364 = n286 & n1297;
  assign n1365 = n1160 & n1289;
  assign n1366 = ~n1294 & n1365;
  assign n1367 = pi64  & n1366;
  assign n1368 = pi66  & n1295;
  assign n1369 = pi65  & n1290;
  assign n1370 = ~n1368 & ~n1369;
  assign n1371 = ~n1364 & n1370;
  assign n1372 = ~n1367 & n1371;
  assign n1373 = pi17  & ~n1372;
  assign n1374 = pi17  & ~n1373;
  assign n1375 = ~n1372 & ~n1373;
  assign n1376 = ~n1374 & ~n1375;
  assign n1377 = ~n1305 & n1376;
  assign n1378 = n1305 & ~n1376;
  assign n1379 = ~n1377 & ~n1378;
  assign n1380 = n401 & n938;
  assign n1381 = pi67  & n1052;
  assign n1382 = pi69  & n936;
  assign n1383 = pi68  & n931;
  assign n1384 = ~n1382 & ~n1383;
  assign n1385 = ~n1381 & n1384;
  assign n1386 = ~n1380 & n1385;
  assign n1387 = pi14  & ~n1386;
  assign n1388 = pi14  & ~n1387;
  assign n1389 = ~n1386 & ~n1387;
  assign n1390 = ~n1388 & ~n1389;
  assign n1391 = n1379 & ~n1390;
  assign n1392 = ~n1379 & n1390;
  assign n1393 = ~n1391 & ~n1392;
  assign n1394 = ~n1363 & n1393;
  assign n1395 = ~n1363 & ~n1394;
  assign n1396 = ~n1391 & ~n1394;
  assign n1397 = ~n1392 & n1396;
  assign n1398 = ~n1395 & ~n1397;
  assign n1399 = n576 & n687;
  assign n1400 = pi70  & n763;
  assign n1401 = pi72  & n685;
  assign n1402 = pi71  & n680;
  assign n1403 = ~n1401 & ~n1402;
  assign n1404 = ~n1400 & n1403;
  assign n1405 = ~n1399 & n1404;
  assign n1406 = pi11  & ~n1405;
  assign n1407 = pi11  & ~n1406;
  assign n1408 = ~n1405 & ~n1406;
  assign n1409 = ~n1407 & ~n1408;
  assign n1410 = n1398 & n1409;
  assign n1411 = ~n1398 & ~n1409;
  assign n1412 = ~n1410 & ~n1411;
  assign n1413 = ~n1362 & n1412;
  assign n1414 = n1362 & ~n1412;
  assign n1415 = ~n1413 & ~n1414;
  assign n1416 = n1361 & ~n1415;
  assign n1417 = ~n1361 & n1415;
  assign n1418 = ~n1416 & ~n1417;
  assign n1419 = ~n1350 & n1418;
  assign n1420 = n1350 & ~n1418;
  assign n1421 = ~n1419 & ~n1420;
  assign n1422 = n1349 & ~n1421;
  assign n1423 = ~n1349 & n1421;
  assign n1424 = ~n1422 & ~n1423;
  assign n1425 = ~n1338 & n1424;
  assign n1426 = n1338 & ~n1424;
  assign n1427 = ~n1425 & ~n1426;
  assign n1428 = ~n1221 & ~n1223;
  assign n1429 = ~pi80  & ~pi81 ;
  assign n1430 = pi80  & pi81 ;
  assign n1431 = ~n1429 & ~n1430;
  assign n1432 = ~n1428 & n1431;
  assign n1433 = n1428 & ~n1431;
  assign n1434 = ~n1432 & ~n1433;
  assign n1435 = n262 & n1434;
  assign n1436 = pi79  & n288;
  assign n1437 = pi81  & n267;
  assign n1438 = pi80  & n269;
  assign n1439 = ~n1437 & ~n1438;
  assign n1440 = ~n1436 & n1439;
  assign n1441 = ~n1435 & n1440;
  assign n1442 = pi2  & ~n1441;
  assign n1443 = pi2  & ~n1442;
  assign n1444 = ~n1441 & ~n1442;
  assign n1445 = ~n1443 & ~n1444;
  assign n1446 = n1427 & ~n1445;
  assign n1447 = n1427 & ~n1446;
  assign n1448 = ~n1445 & ~n1446;
  assign n1449 = ~n1447 & ~n1448;
  assign n1450 = ~n1236 & n1331;
  assign n1451 = ~n1335 & ~n1450;
  assign n1452 = ~n1449 & ~n1451;
  assign n1453 = n1449 & n1451;
  assign po17  = ~n1452 & ~n1453;
  assign n1455 = ~n1423 & ~n1425;
  assign n1456 = n342 & n1122;
  assign n1457 = pi77  & n380;
  assign n1458 = pi79  & n340;
  assign n1459 = pi78  & n335;
  assign n1460 = ~n1458 & ~n1459;
  assign n1461 = ~n1457 & n1460;
  assign n1462 = ~n1456 & n1461;
  assign n1463 = pi5  & ~n1462;
  assign n1464 = pi5  & ~n1463;
  assign n1465 = ~n1462 & ~n1463;
  assign n1466 = ~n1464 & ~n1465;
  assign n1467 = ~n1417 & ~n1419;
  assign n1468 = n498 & n891;
  assign n1469 = pi74  & n537;
  assign n1470 = pi76  & n496;
  assign n1471 = pi75  & n491;
  assign n1472 = ~n1470 & ~n1471;
  assign n1473 = ~n1469 & n1472;
  assign n1474 = ~n1468 & n1473;
  assign n1475 = pi8  & ~n1474;
  assign n1476 = pi8  & ~n1475;
  assign n1477 = ~n1474 & ~n1475;
  assign n1478 = ~n1476 & ~n1477;
  assign n1479 = ~n1411 & ~n1413;
  assign n1480 = pi17  & ~pi18 ;
  assign n1481 = ~pi17  & pi18 ;
  assign n1482 = ~n1480 & ~n1481;
  assign n1483 = pi64  & ~n1482;
  assign n1484 = ~n1378 & n1483;
  assign n1485 = n1378 & ~n1483;
  assign n1486 = ~n1484 & ~n1485;
  assign n1487 = n309 & n1297;
  assign n1488 = pi65  & n1366;
  assign n1489 = pi67  & n1295;
  assign n1490 = pi66  & n1290;
  assign n1491 = ~n1489 & ~n1490;
  assign n1492 = ~n1488 & n1491;
  assign n1493 = ~n1487 & n1492;
  assign n1494 = pi17  & ~n1493;
  assign n1495 = pi17  & ~n1494;
  assign n1496 = ~n1493 & ~n1494;
  assign n1497 = ~n1495 & ~n1496;
  assign n1498 = ~n1486 & ~n1497;
  assign n1499 = n1486 & n1497;
  assign n1500 = ~n1498 & ~n1499;
  assign n1501 = n450 & n938;
  assign n1502 = pi68  & n1052;
  assign n1503 = pi70  & n936;
  assign n1504 = pi69  & n931;
  assign n1505 = ~n1503 & ~n1504;
  assign n1506 = ~n1502 & n1505;
  assign n1507 = ~n1501 & n1506;
  assign n1508 = pi14  & ~n1507;
  assign n1509 = pi14  & ~n1508;
  assign n1510 = ~n1507 & ~n1508;
  assign n1511 = ~n1509 & ~n1510;
  assign n1512 = n1500 & ~n1511;
  assign n1513 = n1500 & ~n1512;
  assign n1514 = ~n1511 & ~n1512;
  assign n1515 = ~n1513 & ~n1514;
  assign n1516 = ~n1396 & n1515;
  assign n1517 = n1396 & ~n1515;
  assign n1518 = ~n1516 & ~n1517;
  assign n1519 = n642 & n687;
  assign n1520 = pi71  & n763;
  assign n1521 = pi73  & n685;
  assign n1522 = pi72  & n680;
  assign n1523 = ~n1521 & ~n1522;
  assign n1524 = ~n1520 & n1523;
  assign n1525 = ~n1519 & n1524;
  assign n1526 = pi11  & ~n1525;
  assign n1527 = pi11  & ~n1526;
  assign n1528 = ~n1525 & ~n1526;
  assign n1529 = ~n1527 & ~n1528;
  assign n1530 = ~n1518 & ~n1529;
  assign n1531 = n1518 & n1529;
  assign n1532 = ~n1530 & ~n1531;
  assign n1533 = ~n1479 & n1532;
  assign n1534 = n1479 & ~n1532;
  assign n1535 = ~n1533 & ~n1534;
  assign n1536 = n1478 & ~n1535;
  assign n1537 = ~n1478 & n1535;
  assign n1538 = ~n1536 & ~n1537;
  assign n1539 = ~n1467 & n1538;
  assign n1540 = n1467 & ~n1538;
  assign n1541 = ~n1539 & ~n1540;
  assign n1542 = ~n1466 & n1541;
  assign n1543 = n1466 & ~n1541;
  assign n1544 = ~n1542 & ~n1543;
  assign n1545 = ~n1455 & n1544;
  assign n1546 = n1455 & ~n1544;
  assign n1547 = ~n1545 & ~n1546;
  assign n1548 = ~n1430 & ~n1432;
  assign n1549 = ~pi81  & ~pi82 ;
  assign n1550 = pi81  & pi82 ;
  assign n1551 = ~n1549 & ~n1550;
  assign n1552 = ~n1548 & n1551;
  assign n1553 = n1548 & ~n1551;
  assign n1554 = ~n1552 & ~n1553;
  assign n1555 = n262 & n1554;
  assign n1556 = pi80  & n288;
  assign n1557 = pi82  & n267;
  assign n1558 = pi81  & n269;
  assign n1559 = ~n1557 & ~n1558;
  assign n1560 = ~n1556 & n1559;
  assign n1561 = ~n1555 & n1560;
  assign n1562 = pi2  & ~n1561;
  assign n1563 = pi2  & ~n1562;
  assign n1564 = ~n1561 & ~n1562;
  assign n1565 = ~n1563 & ~n1564;
  assign n1566 = n1547 & ~n1565;
  assign n1567 = n1547 & ~n1566;
  assign n1568 = ~n1565 & ~n1566;
  assign n1569 = ~n1567 & ~n1568;
  assign n1570 = ~n1446 & ~n1452;
  assign n1571 = ~n1569 & ~n1570;
  assign n1572 = n1569 & n1570;
  assign po18  = ~n1571 & ~n1572;
  assign n1574 = ~n1396 & ~n1515;
  assign n1575 = ~n1512 & ~n1574;
  assign n1576 = n475 & n938;
  assign n1577 = pi69  & n1052;
  assign n1578 = pi71  & n936;
  assign n1579 = pi70  & n931;
  assign n1580 = ~n1578 & ~n1579;
  assign n1581 = ~n1577 & n1580;
  assign n1582 = ~n1576 & n1581;
  assign n1583 = pi14  & ~n1582;
  assign n1584 = pi14  & ~n1583;
  assign n1585 = ~n1582 & ~n1583;
  assign n1586 = ~n1584 & ~n1585;
  assign n1587 = n1378 & n1483;
  assign n1588 = ~n1498 & ~n1587;
  assign n1589 = n359 & n1297;
  assign n1590 = pi66  & n1366;
  assign n1591 = pi68  & n1295;
  assign n1592 = pi67  & n1290;
  assign n1593 = ~n1591 & ~n1592;
  assign n1594 = ~n1590 & n1593;
  assign n1595 = ~n1589 & n1594;
  assign n1596 = pi17  & ~n1595;
  assign n1597 = pi17  & ~n1596;
  assign n1598 = ~n1595 & ~n1596;
  assign n1599 = ~n1597 & ~n1598;
  assign n1600 = pi20  & ~n1483;
  assign n1601 = ~pi18  & pi19 ;
  assign n1602 = pi18  & ~pi19 ;
  assign n1603 = ~n1601 & ~n1602;
  assign n1604 = n1482 & ~n1603;
  assign n1605 = pi64  & n1604;
  assign n1606 = ~pi19  & pi20 ;
  assign n1607 = pi19  & ~pi20 ;
  assign n1608 = ~n1606 & ~n1607;
  assign n1609 = ~n1482 & n1608;
  assign n1610 = pi65  & n1609;
  assign n1611 = ~n1482 & ~n1608;
  assign n1612 = ~n265 & n1611;
  assign n1613 = ~n1605 & ~n1610;
  assign n1614 = ~n1612 & n1613;
  assign n1615 = pi20  & ~n1614;
  assign n1616 = pi20  & ~n1615;
  assign n1617 = ~n1614 & ~n1615;
  assign n1618 = ~n1616 & ~n1617;
  assign n1619 = n1600 & ~n1618;
  assign n1620 = ~n1600 & n1618;
  assign n1621 = ~n1619 & ~n1620;
  assign n1622 = n1599 & n1621;
  assign n1623 = ~n1599 & ~n1621;
  assign n1624 = ~n1622 & ~n1623;
  assign n1625 = ~n1588 & ~n1624;
  assign n1626 = n1588 & n1624;
  assign n1627 = ~n1625 & ~n1626;
  assign n1628 = ~n1586 & n1627;
  assign n1629 = n1586 & ~n1627;
  assign n1630 = ~n1628 & ~n1629;
  assign n1631 = ~n1575 & n1630;
  assign n1632 = n1575 & ~n1630;
  assign n1633 = ~n1631 & ~n1632;
  assign n1634 = n687 & n729;
  assign n1635 = pi72  & n763;
  assign n1636 = pi74  & n685;
  assign n1637 = pi73  & n680;
  assign n1638 = ~n1636 & ~n1637;
  assign n1639 = ~n1635 & n1638;
  assign n1640 = ~n1634 & n1639;
  assign n1641 = pi11  & ~n1640;
  assign n1642 = pi11  & ~n1641;
  assign n1643 = ~n1640 & ~n1641;
  assign n1644 = ~n1642 & ~n1643;
  assign n1645 = n1633 & ~n1644;
  assign n1646 = n1633 & ~n1645;
  assign n1647 = ~n1644 & ~n1645;
  assign n1648 = ~n1646 & ~n1647;
  assign n1649 = ~n1530 & ~n1533;
  assign n1650 = n1648 & n1649;
  assign n1651 = ~n1648 & ~n1649;
  assign n1652 = ~n1650 & ~n1651;
  assign n1653 = n498 & n999;
  assign n1654 = pi75  & n537;
  assign n1655 = pi77  & n496;
  assign n1656 = pi76  & n491;
  assign n1657 = ~n1655 & ~n1656;
  assign n1658 = ~n1654 & n1657;
  assign n1659 = ~n1653 & n1658;
  assign n1660 = pi8  & ~n1659;
  assign n1661 = pi8  & ~n1660;
  assign n1662 = ~n1659 & ~n1660;
  assign n1663 = ~n1661 & ~n1662;
  assign n1664 = ~n1652 & n1663;
  assign n1665 = n1652 & ~n1663;
  assign n1666 = ~n1664 & ~n1665;
  assign n1667 = ~n1537 & ~n1539;
  assign n1668 = n1666 & ~n1667;
  assign n1669 = ~n1666 & n1667;
  assign n1670 = ~n1668 & ~n1669;
  assign n1671 = n342 & n1225;
  assign n1672 = pi78  & n380;
  assign n1673 = pi80  & n340;
  assign n1674 = pi79  & n335;
  assign n1675 = ~n1673 & ~n1674;
  assign n1676 = ~n1672 & n1675;
  assign n1677 = ~n1671 & n1676;
  assign n1678 = pi5  & ~n1677;
  assign n1679 = pi5  & ~n1678;
  assign n1680 = ~n1677 & ~n1678;
  assign n1681 = ~n1679 & ~n1680;
  assign n1682 = n1670 & ~n1681;
  assign n1683 = n1670 & ~n1682;
  assign n1684 = ~n1681 & ~n1682;
  assign n1685 = ~n1683 & ~n1684;
  assign n1686 = ~n1542 & ~n1545;
  assign n1687 = n1685 & n1686;
  assign n1688 = ~n1685 & ~n1686;
  assign n1689 = ~n1687 & ~n1688;
  assign n1690 = ~n1550 & ~n1552;
  assign n1691 = ~pi82  & ~pi83 ;
  assign n1692 = pi82  & pi83 ;
  assign n1693 = ~n1691 & ~n1692;
  assign n1694 = ~n1690 & n1693;
  assign n1695 = n1690 & ~n1693;
  assign n1696 = ~n1694 & ~n1695;
  assign n1697 = n262 & n1696;
  assign n1698 = pi81  & n288;
  assign n1699 = pi83  & n267;
  assign n1700 = pi82  & n269;
  assign n1701 = ~n1699 & ~n1700;
  assign n1702 = ~n1698 & n1701;
  assign n1703 = ~n1697 & n1702;
  assign n1704 = pi2  & ~n1703;
  assign n1705 = pi2  & ~n1704;
  assign n1706 = ~n1703 & ~n1704;
  assign n1707 = ~n1705 & ~n1706;
  assign n1708 = n1689 & ~n1707;
  assign n1709 = n1689 & ~n1708;
  assign n1710 = ~n1707 & ~n1708;
  assign n1711 = ~n1709 & ~n1710;
  assign n1712 = ~n1566 & ~n1571;
  assign n1713 = ~n1711 & ~n1712;
  assign n1714 = n1711 & n1712;
  assign po19  = ~n1713 & ~n1714;
  assign n1716 = ~n1682 & ~n1688;
  assign n1717 = n342 & n1434;
  assign n1718 = pi79  & n380;
  assign n1719 = pi81  & n340;
  assign n1720 = pi80  & n335;
  assign n1721 = ~n1719 & ~n1720;
  assign n1722 = ~n1718 & n1721;
  assign n1723 = ~n1717 & n1722;
  assign n1724 = pi5  & ~n1723;
  assign n1725 = pi5  & ~n1724;
  assign n1726 = ~n1723 & ~n1724;
  assign n1727 = ~n1725 & ~n1726;
  assign n1728 = ~n1645 & ~n1651;
  assign n1729 = n687 & n809;
  assign n1730 = pi73  & n763;
  assign n1731 = pi75  & n685;
  assign n1732 = pi74  & n680;
  assign n1733 = ~n1731 & ~n1732;
  assign n1734 = ~n1730 & n1733;
  assign n1735 = ~n1729 & n1734;
  assign n1736 = pi11  & ~n1735;
  assign n1737 = pi11  & ~n1736;
  assign n1738 = ~n1735 & ~n1736;
  assign n1739 = ~n1737 & ~n1738;
  assign n1740 = ~n1628 & ~n1631;
  assign n1741 = ~n1599 & n1621;
  assign n1742 = ~n1625 & ~n1741;
  assign n1743 = n286 & n1611;
  assign n1744 = n1482 & n1603;
  assign n1745 = ~n1608 & n1744;
  assign n1746 = pi64  & n1745;
  assign n1747 = pi66  & n1609;
  assign n1748 = pi65  & n1604;
  assign n1749 = ~n1747 & ~n1748;
  assign n1750 = ~n1743 & n1749;
  assign n1751 = ~n1746 & n1750;
  assign n1752 = pi20  & ~n1751;
  assign n1753 = pi20  & ~n1752;
  assign n1754 = ~n1751 & ~n1752;
  assign n1755 = ~n1753 & ~n1754;
  assign n1756 = ~n1619 & n1755;
  assign n1757 = n1619 & ~n1755;
  assign n1758 = ~n1756 & ~n1757;
  assign n1759 = n401 & n1297;
  assign n1760 = pi67  & n1366;
  assign n1761 = pi69  & n1295;
  assign n1762 = pi68  & n1290;
  assign n1763 = ~n1761 & ~n1762;
  assign n1764 = ~n1760 & n1763;
  assign n1765 = ~n1759 & n1764;
  assign n1766 = pi17  & ~n1765;
  assign n1767 = pi17  & ~n1766;
  assign n1768 = ~n1765 & ~n1766;
  assign n1769 = ~n1767 & ~n1768;
  assign n1770 = n1758 & ~n1769;
  assign n1771 = ~n1758 & n1769;
  assign n1772 = ~n1770 & ~n1771;
  assign n1773 = ~n1742 & n1772;
  assign n1774 = ~n1742 & ~n1773;
  assign n1775 = ~n1770 & ~n1773;
  assign n1776 = ~n1771 & n1775;
  assign n1777 = ~n1774 & ~n1776;
  assign n1778 = n576 & n938;
  assign n1779 = pi70  & n1052;
  assign n1780 = pi72  & n936;
  assign n1781 = pi71  & n931;
  assign n1782 = ~n1780 & ~n1781;
  assign n1783 = ~n1779 & n1782;
  assign n1784 = ~n1778 & n1783;
  assign n1785 = pi14  & ~n1784;
  assign n1786 = pi14  & ~n1785;
  assign n1787 = ~n1784 & ~n1785;
  assign n1788 = ~n1786 & ~n1787;
  assign n1789 = n1777 & n1788;
  assign n1790 = ~n1777 & ~n1788;
  assign n1791 = ~n1789 & ~n1790;
  assign n1792 = ~n1740 & n1791;
  assign n1793 = n1740 & ~n1791;
  assign n1794 = ~n1792 & ~n1793;
  assign n1795 = n1739 & ~n1794;
  assign n1796 = ~n1739 & n1794;
  assign n1797 = ~n1795 & ~n1796;
  assign n1798 = ~n1728 & n1797;
  assign n1799 = n1728 & ~n1797;
  assign n1800 = ~n1798 & ~n1799;
  assign n1801 = n498 & n1025;
  assign n1802 = pi76  & n537;
  assign n1803 = pi78  & n496;
  assign n1804 = pi77  & n491;
  assign n1805 = ~n1803 & ~n1804;
  assign n1806 = ~n1802 & n1805;
  assign n1807 = ~n1801 & n1806;
  assign n1808 = pi8  & ~n1807;
  assign n1809 = pi8  & ~n1808;
  assign n1810 = ~n1807 & ~n1808;
  assign n1811 = ~n1809 & ~n1810;
  assign n1812 = n1800 & ~n1811;
  assign n1813 = n1800 & ~n1812;
  assign n1814 = ~n1811 & ~n1812;
  assign n1815 = ~n1813 & ~n1814;
  assign n1816 = ~n1665 & ~n1668;
  assign n1817 = ~n1815 & ~n1816;
  assign n1818 = n1815 & n1816;
  assign n1819 = ~n1817 & ~n1818;
  assign n1820 = ~n1727 & n1819;
  assign n1821 = ~n1727 & ~n1820;
  assign n1822 = n1819 & ~n1820;
  assign n1823 = ~n1821 & ~n1822;
  assign n1824 = ~n1716 & ~n1823;
  assign n1825 = ~n1716 & ~n1824;
  assign n1826 = ~n1823 & ~n1824;
  assign n1827 = ~n1825 & ~n1826;
  assign n1828 = ~n1692 & ~n1694;
  assign n1829 = ~pi83  & ~pi84 ;
  assign n1830 = pi83  & pi84 ;
  assign n1831 = ~n1829 & ~n1830;
  assign n1832 = ~n1828 & n1831;
  assign n1833 = n1828 & ~n1831;
  assign n1834 = ~n1832 & ~n1833;
  assign n1835 = n262 & n1834;
  assign n1836 = pi82  & n288;
  assign n1837 = pi84  & n267;
  assign n1838 = pi83  & n269;
  assign n1839 = ~n1837 & ~n1838;
  assign n1840 = ~n1836 & n1839;
  assign n1841 = ~n1835 & n1840;
  assign n1842 = pi2  & ~n1841;
  assign n1843 = pi2  & ~n1842;
  assign n1844 = ~n1841 & ~n1842;
  assign n1845 = ~n1843 & ~n1844;
  assign n1846 = ~n1827 & ~n1845;
  assign n1847 = ~n1827 & ~n1846;
  assign n1848 = ~n1845 & ~n1846;
  assign n1849 = ~n1847 & ~n1848;
  assign n1850 = ~n1708 & ~n1713;
  assign n1851 = ~n1849 & ~n1850;
  assign n1852 = n1849 & n1850;
  assign po20  = ~n1851 & ~n1852;
  assign n1854 = ~n1812 & ~n1817;
  assign n1855 = n498 & n1122;
  assign n1856 = pi77  & n537;
  assign n1857 = pi79  & n496;
  assign n1858 = pi78  & n491;
  assign n1859 = ~n1857 & ~n1858;
  assign n1860 = ~n1856 & n1859;
  assign n1861 = ~n1855 & n1860;
  assign n1862 = pi8  & ~n1861;
  assign n1863 = pi8  & ~n1862;
  assign n1864 = ~n1861 & ~n1862;
  assign n1865 = ~n1863 & ~n1864;
  assign n1866 = ~n1796 & ~n1798;
  assign n1867 = n687 & n891;
  assign n1868 = pi74  & n763;
  assign n1869 = pi76  & n685;
  assign n1870 = pi75  & n680;
  assign n1871 = ~n1869 & ~n1870;
  assign n1872 = ~n1868 & n1871;
  assign n1873 = ~n1867 & n1872;
  assign n1874 = pi11  & ~n1873;
  assign n1875 = pi11  & ~n1874;
  assign n1876 = ~n1873 & ~n1874;
  assign n1877 = ~n1875 & ~n1876;
  assign n1878 = ~n1790 & ~n1792;
  assign n1879 = pi20  & ~pi21 ;
  assign n1880 = ~pi20  & pi21 ;
  assign n1881 = ~n1879 & ~n1880;
  assign n1882 = pi64  & ~n1881;
  assign n1883 = ~n1757 & n1882;
  assign n1884 = n1757 & ~n1882;
  assign n1885 = ~n1883 & ~n1884;
  assign n1886 = n309 & n1611;
  assign n1887 = pi65  & n1745;
  assign n1888 = pi67  & n1609;
  assign n1889 = pi66  & n1604;
  assign n1890 = ~n1888 & ~n1889;
  assign n1891 = ~n1887 & n1890;
  assign n1892 = ~n1886 & n1891;
  assign n1893 = pi20  & ~n1892;
  assign n1894 = pi20  & ~n1893;
  assign n1895 = ~n1892 & ~n1893;
  assign n1896 = ~n1894 & ~n1895;
  assign n1897 = ~n1885 & ~n1896;
  assign n1898 = n1885 & n1896;
  assign n1899 = ~n1897 & ~n1898;
  assign n1900 = n450 & n1297;
  assign n1901 = pi68  & n1366;
  assign n1902 = pi70  & n1295;
  assign n1903 = pi69  & n1290;
  assign n1904 = ~n1902 & ~n1903;
  assign n1905 = ~n1901 & n1904;
  assign n1906 = ~n1900 & n1905;
  assign n1907 = pi17  & ~n1906;
  assign n1908 = pi17  & ~n1907;
  assign n1909 = ~n1906 & ~n1907;
  assign n1910 = ~n1908 & ~n1909;
  assign n1911 = n1899 & ~n1910;
  assign n1912 = n1899 & ~n1911;
  assign n1913 = ~n1910 & ~n1911;
  assign n1914 = ~n1912 & ~n1913;
  assign n1915 = ~n1775 & n1914;
  assign n1916 = n1775 & ~n1914;
  assign n1917 = ~n1915 & ~n1916;
  assign n1918 = n642 & n938;
  assign n1919 = pi71  & n1052;
  assign n1920 = pi73  & n936;
  assign n1921 = pi72  & n931;
  assign n1922 = ~n1920 & ~n1921;
  assign n1923 = ~n1919 & n1922;
  assign n1924 = ~n1918 & n1923;
  assign n1925 = pi14  & ~n1924;
  assign n1926 = pi14  & ~n1925;
  assign n1927 = ~n1924 & ~n1925;
  assign n1928 = ~n1926 & ~n1927;
  assign n1929 = ~n1917 & ~n1928;
  assign n1930 = n1917 & n1928;
  assign n1931 = ~n1929 & ~n1930;
  assign n1932 = ~n1878 & n1931;
  assign n1933 = n1878 & ~n1931;
  assign n1934 = ~n1932 & ~n1933;
  assign n1935 = n1877 & ~n1934;
  assign n1936 = ~n1877 & n1934;
  assign n1937 = ~n1935 & ~n1936;
  assign n1938 = ~n1866 & n1937;
  assign n1939 = n1866 & ~n1937;
  assign n1940 = ~n1938 & ~n1939;
  assign n1941 = ~n1865 & n1940;
  assign n1942 = n1865 & ~n1940;
  assign n1943 = ~n1941 & ~n1942;
  assign n1944 = ~n1854 & n1943;
  assign n1945 = n1854 & ~n1943;
  assign n1946 = ~n1944 & ~n1945;
  assign n1947 = n342 & n1554;
  assign n1948 = pi80  & n380;
  assign n1949 = pi82  & n340;
  assign n1950 = pi81  & n335;
  assign n1951 = ~n1949 & ~n1950;
  assign n1952 = ~n1948 & n1951;
  assign n1953 = ~n1947 & n1952;
  assign n1954 = pi5  & ~n1953;
  assign n1955 = pi5  & ~n1954;
  assign n1956 = ~n1953 & ~n1954;
  assign n1957 = ~n1955 & ~n1956;
  assign n1958 = n1946 & ~n1957;
  assign n1959 = n1946 & ~n1958;
  assign n1960 = ~n1957 & ~n1958;
  assign n1961 = ~n1959 & ~n1960;
  assign n1962 = ~n1820 & ~n1824;
  assign n1963 = n1961 & n1962;
  assign n1964 = ~n1961 & ~n1962;
  assign n1965 = ~n1963 & ~n1964;
  assign n1966 = ~n1830 & ~n1832;
  assign n1967 = ~pi84  & ~pi85 ;
  assign n1968 = pi84  & pi85 ;
  assign n1969 = ~n1967 & ~n1968;
  assign n1970 = ~n1966 & n1969;
  assign n1971 = n1966 & ~n1969;
  assign n1972 = ~n1970 & ~n1971;
  assign n1973 = n262 & n1972;
  assign n1974 = pi83  & n288;
  assign n1975 = pi85  & n267;
  assign n1976 = pi84  & n269;
  assign n1977 = ~n1975 & ~n1976;
  assign n1978 = ~n1974 & n1977;
  assign n1979 = ~n1973 & n1978;
  assign n1980 = pi2  & ~n1979;
  assign n1981 = pi2  & ~n1980;
  assign n1982 = ~n1979 & ~n1980;
  assign n1983 = ~n1981 & ~n1982;
  assign n1984 = n1965 & ~n1983;
  assign n1985 = n1965 & ~n1984;
  assign n1986 = ~n1983 & ~n1984;
  assign n1987 = ~n1985 & ~n1986;
  assign n1988 = ~n1846 & ~n1851;
  assign n1989 = ~n1987 & ~n1988;
  assign n1990 = n1987 & n1988;
  assign po21  = ~n1989 & ~n1990;
  assign n1992 = ~n1984 & ~n1989;
  assign n1993 = ~n1941 & ~n1944;
  assign n1994 = n498 & n1225;
  assign n1995 = pi78  & n537;
  assign n1996 = pi80  & n496;
  assign n1997 = pi79  & n491;
  assign n1998 = ~n1996 & ~n1997;
  assign n1999 = ~n1995 & n1998;
  assign n2000 = ~n1994 & n1999;
  assign n2001 = pi8  & ~n2000;
  assign n2002 = pi8  & ~n2001;
  assign n2003 = ~n2000 & ~n2001;
  assign n2004 = ~n2002 & ~n2003;
  assign n2005 = ~n1936 & ~n1938;
  assign n2006 = ~n1775 & ~n1914;
  assign n2007 = ~n1911 & ~n2006;
  assign n2008 = n475 & n1297;
  assign n2009 = pi69  & n1366;
  assign n2010 = pi71  & n1295;
  assign n2011 = pi70  & n1290;
  assign n2012 = ~n2010 & ~n2011;
  assign n2013 = ~n2009 & n2012;
  assign n2014 = ~n2008 & n2013;
  assign n2015 = pi17  & ~n2014;
  assign n2016 = pi17  & ~n2015;
  assign n2017 = ~n2014 & ~n2015;
  assign n2018 = ~n2016 & ~n2017;
  assign n2019 = n1757 & n1882;
  assign n2020 = ~n1897 & ~n2019;
  assign n2021 = n359 & n1611;
  assign n2022 = pi66  & n1745;
  assign n2023 = pi68  & n1609;
  assign n2024 = pi67  & n1604;
  assign n2025 = ~n2023 & ~n2024;
  assign n2026 = ~n2022 & n2025;
  assign n2027 = ~n2021 & n2026;
  assign n2028 = pi20  & ~n2027;
  assign n2029 = pi20  & ~n2028;
  assign n2030 = ~n2027 & ~n2028;
  assign n2031 = ~n2029 & ~n2030;
  assign n2032 = pi23  & ~n1882;
  assign n2033 = ~pi21  & pi22 ;
  assign n2034 = pi21  & ~pi22 ;
  assign n2035 = ~n2033 & ~n2034;
  assign n2036 = n1881 & ~n2035;
  assign n2037 = pi64  & n2036;
  assign n2038 = ~pi22  & pi23 ;
  assign n2039 = pi22  & ~pi23 ;
  assign n2040 = ~n2038 & ~n2039;
  assign n2041 = ~n1881 & n2040;
  assign n2042 = pi65  & n2041;
  assign n2043 = ~n1881 & ~n2040;
  assign n2044 = ~n265 & n2043;
  assign n2045 = ~n2037 & ~n2042;
  assign n2046 = ~n2044 & n2045;
  assign n2047 = pi23  & ~n2046;
  assign n2048 = pi23  & ~n2047;
  assign n2049 = ~n2046 & ~n2047;
  assign n2050 = ~n2048 & ~n2049;
  assign n2051 = n2032 & ~n2050;
  assign n2052 = ~n2032 & n2050;
  assign n2053 = ~n2051 & ~n2052;
  assign n2054 = n2031 & n2053;
  assign n2055 = ~n2031 & ~n2053;
  assign n2056 = ~n2054 & ~n2055;
  assign n2057 = ~n2020 & ~n2056;
  assign n2058 = n2020 & n2056;
  assign n2059 = ~n2057 & ~n2058;
  assign n2060 = ~n2018 & n2059;
  assign n2061 = n2018 & ~n2059;
  assign n2062 = ~n2060 & ~n2061;
  assign n2063 = ~n2007 & n2062;
  assign n2064 = n2007 & ~n2062;
  assign n2065 = ~n2063 & ~n2064;
  assign n2066 = n729 & n938;
  assign n2067 = pi72  & n1052;
  assign n2068 = pi74  & n936;
  assign n2069 = pi73  & n931;
  assign n2070 = ~n2068 & ~n2069;
  assign n2071 = ~n2067 & n2070;
  assign n2072 = ~n2066 & n2071;
  assign n2073 = pi14  & ~n2072;
  assign n2074 = pi14  & ~n2073;
  assign n2075 = ~n2072 & ~n2073;
  assign n2076 = ~n2074 & ~n2075;
  assign n2077 = n2065 & ~n2076;
  assign n2078 = n2065 & ~n2077;
  assign n2079 = ~n2076 & ~n2077;
  assign n2080 = ~n2078 & ~n2079;
  assign n2081 = ~n1929 & ~n1932;
  assign n2082 = n2080 & n2081;
  assign n2083 = ~n2080 & ~n2081;
  assign n2084 = ~n2082 & ~n2083;
  assign n2085 = n687 & n999;
  assign n2086 = pi75  & n763;
  assign n2087 = pi77  & n685;
  assign n2088 = pi76  & n680;
  assign n2089 = ~n2087 & ~n2088;
  assign n2090 = ~n2086 & n2089;
  assign n2091 = ~n2085 & n2090;
  assign n2092 = pi11  & ~n2091;
  assign n2093 = pi11  & ~n2092;
  assign n2094 = ~n2091 & ~n2092;
  assign n2095 = ~n2093 & ~n2094;
  assign n2096 = ~n2084 & n2095;
  assign n2097 = n2084 & ~n2095;
  assign n2098 = ~n2096 & ~n2097;
  assign n2099 = ~n2005 & n2098;
  assign n2100 = n2005 & ~n2098;
  assign n2101 = ~n2099 & ~n2100;
  assign n2102 = ~n2004 & n2101;
  assign n2103 = n2004 & ~n2101;
  assign n2104 = ~n2102 & ~n2103;
  assign n2105 = ~n1993 & n2104;
  assign n2106 = n1993 & ~n2104;
  assign n2107 = ~n2105 & ~n2106;
  assign n2108 = n342 & n1696;
  assign n2109 = pi81  & n380;
  assign n2110 = pi83  & n340;
  assign n2111 = pi82  & n335;
  assign n2112 = ~n2110 & ~n2111;
  assign n2113 = ~n2109 & n2112;
  assign n2114 = ~n2108 & n2113;
  assign n2115 = pi5  & ~n2114;
  assign n2116 = pi5  & ~n2115;
  assign n2117 = ~n2114 & ~n2115;
  assign n2118 = ~n2116 & ~n2117;
  assign n2119 = n2107 & ~n2118;
  assign n2120 = n2107 & ~n2119;
  assign n2121 = ~n2118 & ~n2119;
  assign n2122 = ~n2120 & ~n2121;
  assign n2123 = ~n1958 & ~n1964;
  assign n2124 = n2122 & n2123;
  assign n2125 = ~n2122 & ~n2123;
  assign n2126 = ~n2124 & ~n2125;
  assign n2127 = ~n1968 & ~n1970;
  assign n2128 = ~pi85  & ~pi86 ;
  assign n2129 = pi85  & pi86 ;
  assign n2130 = ~n2128 & ~n2129;
  assign n2131 = ~n2127 & n2130;
  assign n2132 = n2127 & ~n2130;
  assign n2133 = ~n2131 & ~n2132;
  assign n2134 = n262 & n2133;
  assign n2135 = pi84  & n288;
  assign n2136 = pi86  & n267;
  assign n2137 = pi85  & n269;
  assign n2138 = ~n2136 & ~n2137;
  assign n2139 = ~n2135 & n2138;
  assign n2140 = ~n2134 & n2139;
  assign n2141 = pi2  & ~n2140;
  assign n2142 = pi2  & ~n2141;
  assign n2143 = ~n2140 & ~n2141;
  assign n2144 = ~n2142 & ~n2143;
  assign n2145 = ~n2126 & n2144;
  assign n2146 = n2126 & ~n2144;
  assign n2147 = ~n2145 & ~n2146;
  assign n2148 = ~n1992 & n2147;
  assign n2149 = n1992 & ~n2147;
  assign po22  = ~n2148 & ~n2149;
  assign n2151 = ~n2102 & ~n2105;
  assign n2152 = n498 & n1434;
  assign n2153 = pi79  & n537;
  assign n2154 = pi81  & n496;
  assign n2155 = pi80  & n491;
  assign n2156 = ~n2154 & ~n2155;
  assign n2157 = ~n2153 & n2156;
  assign n2158 = ~n2152 & n2157;
  assign n2159 = pi8  & ~n2158;
  assign n2160 = pi8  & ~n2159;
  assign n2161 = ~n2158 & ~n2159;
  assign n2162 = ~n2160 & ~n2161;
  assign n2163 = ~n2077 & ~n2083;
  assign n2164 = n809 & n938;
  assign n2165 = pi73  & n1052;
  assign n2166 = pi75  & n936;
  assign n2167 = pi74  & n931;
  assign n2168 = ~n2166 & ~n2167;
  assign n2169 = ~n2165 & n2168;
  assign n2170 = ~n2164 & n2169;
  assign n2171 = pi14  & ~n2170;
  assign n2172 = pi14  & ~n2171;
  assign n2173 = ~n2170 & ~n2171;
  assign n2174 = ~n2172 & ~n2173;
  assign n2175 = ~n2060 & ~n2063;
  assign n2176 = ~n2031 & n2053;
  assign n2177 = ~n2057 & ~n2176;
  assign n2178 = n286 & n2043;
  assign n2179 = n1881 & n2035;
  assign n2180 = ~n2040 & n2179;
  assign n2181 = pi64  & n2180;
  assign n2182 = pi66  & n2041;
  assign n2183 = pi65  & n2036;
  assign n2184 = ~n2182 & ~n2183;
  assign n2185 = ~n2178 & n2184;
  assign n2186 = ~n2181 & n2185;
  assign n2187 = pi23  & ~n2186;
  assign n2188 = pi23  & ~n2187;
  assign n2189 = ~n2186 & ~n2187;
  assign n2190 = ~n2188 & ~n2189;
  assign n2191 = ~n2051 & n2190;
  assign n2192 = n2051 & ~n2190;
  assign n2193 = ~n2191 & ~n2192;
  assign n2194 = n401 & n1611;
  assign n2195 = pi67  & n1745;
  assign n2196 = pi69  & n1609;
  assign n2197 = pi68  & n1604;
  assign n2198 = ~n2196 & ~n2197;
  assign n2199 = ~n2195 & n2198;
  assign n2200 = ~n2194 & n2199;
  assign n2201 = pi20  & ~n2200;
  assign n2202 = pi20  & ~n2201;
  assign n2203 = ~n2200 & ~n2201;
  assign n2204 = ~n2202 & ~n2203;
  assign n2205 = n2193 & ~n2204;
  assign n2206 = ~n2193 & n2204;
  assign n2207 = ~n2205 & ~n2206;
  assign n2208 = ~n2177 & n2207;
  assign n2209 = ~n2177 & ~n2208;
  assign n2210 = ~n2205 & ~n2208;
  assign n2211 = ~n2206 & n2210;
  assign n2212 = ~n2209 & ~n2211;
  assign n2213 = n576 & n1297;
  assign n2214 = pi70  & n1366;
  assign n2215 = pi72  & n1295;
  assign n2216 = pi71  & n1290;
  assign n2217 = ~n2215 & ~n2216;
  assign n2218 = ~n2214 & n2217;
  assign n2219 = ~n2213 & n2218;
  assign n2220 = pi17  & ~n2219;
  assign n2221 = pi17  & ~n2220;
  assign n2222 = ~n2219 & ~n2220;
  assign n2223 = ~n2221 & ~n2222;
  assign n2224 = n2212 & n2223;
  assign n2225 = ~n2212 & ~n2223;
  assign n2226 = ~n2224 & ~n2225;
  assign n2227 = ~n2175 & n2226;
  assign n2228 = n2175 & ~n2226;
  assign n2229 = ~n2227 & ~n2228;
  assign n2230 = n2174 & ~n2229;
  assign n2231 = ~n2174 & n2229;
  assign n2232 = ~n2230 & ~n2231;
  assign n2233 = ~n2163 & n2232;
  assign n2234 = n2163 & ~n2232;
  assign n2235 = ~n2233 & ~n2234;
  assign n2236 = n687 & n1025;
  assign n2237 = pi76  & n763;
  assign n2238 = pi78  & n685;
  assign n2239 = pi77  & n680;
  assign n2240 = ~n2238 & ~n2239;
  assign n2241 = ~n2237 & n2240;
  assign n2242 = ~n2236 & n2241;
  assign n2243 = pi11  & ~n2242;
  assign n2244 = pi11  & ~n2243;
  assign n2245 = ~n2242 & ~n2243;
  assign n2246 = ~n2244 & ~n2245;
  assign n2247 = n2235 & ~n2246;
  assign n2248 = n2235 & ~n2247;
  assign n2249 = ~n2246 & ~n2247;
  assign n2250 = ~n2248 & ~n2249;
  assign n2251 = ~n2097 & ~n2099;
  assign n2252 = ~n2250 & ~n2251;
  assign n2253 = n2250 & n2251;
  assign n2254 = ~n2252 & ~n2253;
  assign n2255 = ~n2162 & n2254;
  assign n2256 = ~n2162 & ~n2255;
  assign n2257 = n2254 & ~n2255;
  assign n2258 = ~n2256 & ~n2257;
  assign n2259 = ~n2151 & ~n2258;
  assign n2260 = ~n2151 & ~n2259;
  assign n2261 = ~n2258 & ~n2259;
  assign n2262 = ~n2260 & ~n2261;
  assign n2263 = n342 & n1834;
  assign n2264 = pi82  & n380;
  assign n2265 = pi84  & n340;
  assign n2266 = pi83  & n335;
  assign n2267 = ~n2265 & ~n2266;
  assign n2268 = ~n2264 & n2267;
  assign n2269 = ~n2263 & n2268;
  assign n2270 = pi5  & ~n2269;
  assign n2271 = pi5  & ~n2270;
  assign n2272 = ~n2269 & ~n2270;
  assign n2273 = ~n2271 & ~n2272;
  assign n2274 = ~n2262 & ~n2273;
  assign n2275 = ~n2262 & ~n2274;
  assign n2276 = ~n2273 & ~n2274;
  assign n2277 = ~n2275 & ~n2276;
  assign n2278 = ~n2119 & ~n2125;
  assign n2279 = n2277 & n2278;
  assign n2280 = ~n2277 & ~n2278;
  assign n2281 = ~n2279 & ~n2280;
  assign n2282 = ~n2129 & ~n2131;
  assign n2283 = ~pi86  & ~pi87 ;
  assign n2284 = pi86  & pi87 ;
  assign n2285 = ~n2283 & ~n2284;
  assign n2286 = ~n2282 & n2285;
  assign n2287 = n2282 & ~n2285;
  assign n2288 = ~n2286 & ~n2287;
  assign n2289 = n262 & n2288;
  assign n2290 = pi85  & n288;
  assign n2291 = pi87  & n267;
  assign n2292 = pi86  & n269;
  assign n2293 = ~n2291 & ~n2292;
  assign n2294 = ~n2290 & n2293;
  assign n2295 = ~n2289 & n2294;
  assign n2296 = pi2  & ~n2295;
  assign n2297 = pi2  & ~n2296;
  assign n2298 = ~n2295 & ~n2296;
  assign n2299 = ~n2297 & ~n2298;
  assign n2300 = n2281 & ~n2299;
  assign n2301 = n2281 & ~n2300;
  assign n2302 = ~n2299 & ~n2300;
  assign n2303 = ~n2301 & ~n2302;
  assign n2304 = ~n2146 & ~n2148;
  assign n2305 = ~n2303 & ~n2304;
  assign n2306 = n2303 & n2304;
  assign po23  = ~n2305 & ~n2306;
  assign n2308 = ~n2274 & ~n2280;
  assign n2309 = n342 & n1972;
  assign n2310 = pi83  & n380;
  assign n2311 = pi85  & n340;
  assign n2312 = pi84  & n335;
  assign n2313 = ~n2311 & ~n2312;
  assign n2314 = ~n2310 & n2313;
  assign n2315 = ~n2309 & n2314;
  assign n2316 = pi5  & ~n2315;
  assign n2317 = pi5  & ~n2316;
  assign n2318 = ~n2315 & ~n2316;
  assign n2319 = ~n2317 & ~n2318;
  assign n2320 = ~n2255 & ~n2259;
  assign n2321 = ~n2231 & ~n2233;
  assign n2322 = n891 & n938;
  assign n2323 = pi74  & n1052;
  assign n2324 = pi76  & n936;
  assign n2325 = pi75  & n931;
  assign n2326 = ~n2324 & ~n2325;
  assign n2327 = ~n2323 & n2326;
  assign n2328 = ~n2322 & n2327;
  assign n2329 = pi14  & ~n2328;
  assign n2330 = pi14  & ~n2329;
  assign n2331 = ~n2328 & ~n2329;
  assign n2332 = ~n2330 & ~n2331;
  assign n2333 = ~n2225 & ~n2227;
  assign n2334 = pi23  & ~pi24 ;
  assign n2335 = ~pi23  & pi24 ;
  assign n2336 = ~n2334 & ~n2335;
  assign n2337 = pi64  & ~n2336;
  assign n2338 = ~n2192 & n2337;
  assign n2339 = n2192 & ~n2337;
  assign n2340 = ~n2338 & ~n2339;
  assign n2341 = n309 & n2043;
  assign n2342 = pi65  & n2180;
  assign n2343 = pi67  & n2041;
  assign n2344 = pi66  & n2036;
  assign n2345 = ~n2343 & ~n2344;
  assign n2346 = ~n2342 & n2345;
  assign n2347 = ~n2341 & n2346;
  assign n2348 = pi23  & ~n2347;
  assign n2349 = pi23  & ~n2348;
  assign n2350 = ~n2347 & ~n2348;
  assign n2351 = ~n2349 & ~n2350;
  assign n2352 = ~n2340 & ~n2351;
  assign n2353 = n2340 & n2351;
  assign n2354 = ~n2352 & ~n2353;
  assign n2355 = n450 & n1611;
  assign n2356 = pi68  & n1745;
  assign n2357 = pi70  & n1609;
  assign n2358 = pi69  & n1604;
  assign n2359 = ~n2357 & ~n2358;
  assign n2360 = ~n2356 & n2359;
  assign n2361 = ~n2355 & n2360;
  assign n2362 = pi20  & ~n2361;
  assign n2363 = pi20  & ~n2362;
  assign n2364 = ~n2361 & ~n2362;
  assign n2365 = ~n2363 & ~n2364;
  assign n2366 = n2354 & ~n2365;
  assign n2367 = n2354 & ~n2366;
  assign n2368 = ~n2365 & ~n2366;
  assign n2369 = ~n2367 & ~n2368;
  assign n2370 = ~n2210 & n2369;
  assign n2371 = n2210 & ~n2369;
  assign n2372 = ~n2370 & ~n2371;
  assign n2373 = n642 & n1297;
  assign n2374 = pi71  & n1366;
  assign n2375 = pi73  & n1295;
  assign n2376 = pi72  & n1290;
  assign n2377 = ~n2375 & ~n2376;
  assign n2378 = ~n2374 & n2377;
  assign n2379 = ~n2373 & n2378;
  assign n2380 = pi17  & ~n2379;
  assign n2381 = pi17  & ~n2380;
  assign n2382 = ~n2379 & ~n2380;
  assign n2383 = ~n2381 & ~n2382;
  assign n2384 = ~n2372 & ~n2383;
  assign n2385 = n2372 & n2383;
  assign n2386 = ~n2384 & ~n2385;
  assign n2387 = ~n2333 & n2386;
  assign n2388 = n2333 & ~n2386;
  assign n2389 = ~n2387 & ~n2388;
  assign n2390 = n2332 & ~n2389;
  assign n2391 = ~n2332 & n2389;
  assign n2392 = ~n2390 & ~n2391;
  assign n2393 = ~n2321 & n2392;
  assign n2394 = n2321 & ~n2392;
  assign n2395 = ~n2393 & ~n2394;
  assign n2396 = n687 & n1122;
  assign n2397 = pi77  & n763;
  assign n2398 = pi79  & n685;
  assign n2399 = pi78  & n680;
  assign n2400 = ~n2398 & ~n2399;
  assign n2401 = ~n2397 & n2400;
  assign n2402 = ~n2396 & n2401;
  assign n2403 = pi11  & ~n2402;
  assign n2404 = pi11  & ~n2403;
  assign n2405 = ~n2402 & ~n2403;
  assign n2406 = ~n2404 & ~n2405;
  assign n2407 = n2395 & ~n2406;
  assign n2408 = n2395 & ~n2407;
  assign n2409 = ~n2406 & ~n2407;
  assign n2410 = ~n2408 & ~n2409;
  assign n2411 = ~n2247 & ~n2252;
  assign n2412 = n2410 & n2411;
  assign n2413 = ~n2410 & ~n2411;
  assign n2414 = ~n2412 & ~n2413;
  assign n2415 = n498 & n1554;
  assign n2416 = pi80  & n537;
  assign n2417 = pi82  & n496;
  assign n2418 = pi81  & n491;
  assign n2419 = ~n2417 & ~n2418;
  assign n2420 = ~n2416 & n2419;
  assign n2421 = ~n2415 & n2420;
  assign n2422 = pi8  & ~n2421;
  assign n2423 = pi8  & ~n2422;
  assign n2424 = ~n2421 & ~n2422;
  assign n2425 = ~n2423 & ~n2424;
  assign n2426 = ~n2414 & n2425;
  assign n2427 = n2414 & ~n2425;
  assign n2428 = ~n2426 & ~n2427;
  assign n2429 = ~n2320 & n2428;
  assign n2430 = n2320 & ~n2428;
  assign n2431 = ~n2429 & ~n2430;
  assign n2432 = ~n2319 & n2431;
  assign n2433 = ~n2319 & ~n2432;
  assign n2434 = n2431 & ~n2432;
  assign n2435 = ~n2433 & ~n2434;
  assign n2436 = ~n2308 & ~n2435;
  assign n2437 = ~n2308 & ~n2436;
  assign n2438 = ~n2435 & ~n2436;
  assign n2439 = ~n2437 & ~n2438;
  assign n2440 = ~n2284 & ~n2286;
  assign n2441 = ~pi87  & ~pi88 ;
  assign n2442 = pi87  & pi88 ;
  assign n2443 = ~n2441 & ~n2442;
  assign n2444 = ~n2440 & n2443;
  assign n2445 = n2440 & ~n2443;
  assign n2446 = ~n2444 & ~n2445;
  assign n2447 = n262 & n2446;
  assign n2448 = pi86  & n288;
  assign n2449 = pi88  & n267;
  assign n2450 = pi87  & n269;
  assign n2451 = ~n2449 & ~n2450;
  assign n2452 = ~n2448 & n2451;
  assign n2453 = ~n2447 & n2452;
  assign n2454 = pi2  & ~n2453;
  assign n2455 = pi2  & ~n2454;
  assign n2456 = ~n2453 & ~n2454;
  assign n2457 = ~n2455 & ~n2456;
  assign n2458 = ~n2439 & ~n2457;
  assign n2459 = ~n2439 & ~n2458;
  assign n2460 = ~n2457 & ~n2458;
  assign n2461 = ~n2459 & ~n2460;
  assign n2462 = ~n2300 & ~n2305;
  assign n2463 = ~n2461 & ~n2462;
  assign n2464 = n2461 & n2462;
  assign po24  = ~n2463 & ~n2464;
  assign n2466 = ~n2458 & ~n2463;
  assign n2467 = ~n2442 & ~n2444;
  assign n2468 = ~pi88  & ~pi89 ;
  assign n2469 = pi88  & pi89 ;
  assign n2470 = ~n2468 & ~n2469;
  assign n2471 = ~n2467 & n2470;
  assign n2472 = n2467 & ~n2470;
  assign n2473 = ~n2471 & ~n2472;
  assign n2474 = n262 & n2473;
  assign n2475 = pi87  & n288;
  assign n2476 = pi89  & n267;
  assign n2477 = pi88  & n269;
  assign n2478 = ~n2476 & ~n2477;
  assign n2479 = ~n2475 & n2478;
  assign n2480 = ~n2474 & n2479;
  assign n2481 = pi2  & ~n2480;
  assign n2482 = pi2  & ~n2481;
  assign n2483 = ~n2480 & ~n2481;
  assign n2484 = ~n2482 & ~n2483;
  assign n2485 = ~n2432 & ~n2436;
  assign n2486 = ~n2210 & ~n2369;
  assign n2487 = ~n2366 & ~n2486;
  assign n2488 = n475 & n1611;
  assign n2489 = pi69  & n1745;
  assign n2490 = pi71  & n1609;
  assign n2491 = pi70  & n1604;
  assign n2492 = ~n2490 & ~n2491;
  assign n2493 = ~n2489 & n2492;
  assign n2494 = ~n2488 & n2493;
  assign n2495 = pi20  & ~n2494;
  assign n2496 = pi20  & ~n2495;
  assign n2497 = ~n2494 & ~n2495;
  assign n2498 = ~n2496 & ~n2497;
  assign n2499 = n2192 & n2337;
  assign n2500 = ~n2352 & ~n2499;
  assign n2501 = n359 & n2043;
  assign n2502 = pi66  & n2180;
  assign n2503 = pi68  & n2041;
  assign n2504 = pi67  & n2036;
  assign n2505 = ~n2503 & ~n2504;
  assign n2506 = ~n2502 & n2505;
  assign n2507 = ~n2501 & n2506;
  assign n2508 = pi23  & ~n2507;
  assign n2509 = pi23  & ~n2508;
  assign n2510 = ~n2507 & ~n2508;
  assign n2511 = ~n2509 & ~n2510;
  assign n2512 = pi26  & ~n2337;
  assign n2513 = ~pi24  & pi25 ;
  assign n2514 = pi24  & ~pi25 ;
  assign n2515 = ~n2513 & ~n2514;
  assign n2516 = n2336 & ~n2515;
  assign n2517 = pi64  & n2516;
  assign n2518 = ~pi25  & pi26 ;
  assign n2519 = pi25  & ~pi26 ;
  assign n2520 = ~n2518 & ~n2519;
  assign n2521 = ~n2336 & n2520;
  assign n2522 = pi65  & n2521;
  assign n2523 = ~n2336 & ~n2520;
  assign n2524 = ~n265 & n2523;
  assign n2525 = ~n2517 & ~n2522;
  assign n2526 = ~n2524 & n2525;
  assign n2527 = pi26  & ~n2526;
  assign n2528 = pi26  & ~n2527;
  assign n2529 = ~n2526 & ~n2527;
  assign n2530 = ~n2528 & ~n2529;
  assign n2531 = n2512 & ~n2530;
  assign n2532 = ~n2512 & n2530;
  assign n2533 = ~n2531 & ~n2532;
  assign n2534 = n2511 & n2533;
  assign n2535 = ~n2511 & ~n2533;
  assign n2536 = ~n2534 & ~n2535;
  assign n2537 = ~n2500 & ~n2536;
  assign n2538 = n2500 & n2536;
  assign n2539 = ~n2537 & ~n2538;
  assign n2540 = ~n2498 & n2539;
  assign n2541 = n2498 & ~n2539;
  assign n2542 = ~n2540 & ~n2541;
  assign n2543 = ~n2487 & n2542;
  assign n2544 = n2487 & ~n2542;
  assign n2545 = ~n2543 & ~n2544;
  assign n2546 = n729 & n1297;
  assign n2547 = pi72  & n1366;
  assign n2548 = pi74  & n1295;
  assign n2549 = pi73  & n1290;
  assign n2550 = ~n2548 & ~n2549;
  assign n2551 = ~n2547 & n2550;
  assign n2552 = ~n2546 & n2551;
  assign n2553 = pi17  & ~n2552;
  assign n2554 = pi17  & ~n2553;
  assign n2555 = ~n2552 & ~n2553;
  assign n2556 = ~n2554 & ~n2555;
  assign n2557 = n2545 & ~n2556;
  assign n2558 = n2545 & ~n2557;
  assign n2559 = ~n2556 & ~n2557;
  assign n2560 = ~n2558 & ~n2559;
  assign n2561 = ~n2384 & ~n2387;
  assign n2562 = n2560 & n2561;
  assign n2563 = ~n2560 & ~n2561;
  assign n2564 = ~n2562 & ~n2563;
  assign n2565 = n938 & n999;
  assign n2566 = pi75  & n1052;
  assign n2567 = pi77  & n936;
  assign n2568 = pi76  & n931;
  assign n2569 = ~n2567 & ~n2568;
  assign n2570 = ~n2566 & n2569;
  assign n2571 = ~n2565 & n2570;
  assign n2572 = pi14  & ~n2571;
  assign n2573 = pi14  & ~n2572;
  assign n2574 = ~n2571 & ~n2572;
  assign n2575 = ~n2573 & ~n2574;
  assign n2576 = ~n2564 & n2575;
  assign n2577 = n2564 & ~n2575;
  assign n2578 = ~n2576 & ~n2577;
  assign n2579 = ~n2391 & ~n2393;
  assign n2580 = n2578 & ~n2579;
  assign n2581 = ~n2578 & n2579;
  assign n2582 = ~n2580 & ~n2581;
  assign n2583 = n687 & n1225;
  assign n2584 = pi78  & n763;
  assign n2585 = pi80  & n685;
  assign n2586 = pi79  & n680;
  assign n2587 = ~n2585 & ~n2586;
  assign n2588 = ~n2584 & n2587;
  assign n2589 = ~n2583 & n2588;
  assign n2590 = pi11  & ~n2589;
  assign n2591 = pi11  & ~n2590;
  assign n2592 = ~n2589 & ~n2590;
  assign n2593 = ~n2591 & ~n2592;
  assign n2594 = n2582 & ~n2593;
  assign n2595 = n2582 & ~n2594;
  assign n2596 = ~n2593 & ~n2594;
  assign n2597 = ~n2595 & ~n2596;
  assign n2598 = ~n2407 & ~n2413;
  assign n2599 = n2597 & n2598;
  assign n2600 = ~n2597 & ~n2598;
  assign n2601 = ~n2599 & ~n2600;
  assign n2602 = n498 & n1696;
  assign n2603 = pi81  & n537;
  assign n2604 = pi83  & n496;
  assign n2605 = pi82  & n491;
  assign n2606 = ~n2604 & ~n2605;
  assign n2607 = ~n2603 & n2606;
  assign n2608 = ~n2602 & n2607;
  assign n2609 = pi8  & ~n2608;
  assign n2610 = pi8  & ~n2609;
  assign n2611 = ~n2608 & ~n2609;
  assign n2612 = ~n2610 & ~n2611;
  assign n2613 = n2601 & ~n2612;
  assign n2614 = n2601 & ~n2613;
  assign n2615 = ~n2612 & ~n2613;
  assign n2616 = ~n2614 & ~n2615;
  assign n2617 = ~n2427 & ~n2429;
  assign n2618 = ~n2616 & ~n2617;
  assign n2619 = ~n2616 & ~n2618;
  assign n2620 = ~n2617 & ~n2618;
  assign n2621 = ~n2619 & ~n2620;
  assign n2622 = n342 & n2133;
  assign n2623 = pi84  & n380;
  assign n2624 = pi86  & n340;
  assign n2625 = pi85  & n335;
  assign n2626 = ~n2624 & ~n2625;
  assign n2627 = ~n2623 & n2626;
  assign n2628 = ~n2622 & n2627;
  assign n2629 = pi5  & ~n2628;
  assign n2630 = pi5  & ~n2629;
  assign n2631 = ~n2628 & ~n2629;
  assign n2632 = ~n2630 & ~n2631;
  assign n2633 = ~n2621 & n2632;
  assign n2634 = n2621 & ~n2632;
  assign n2635 = ~n2633 & ~n2634;
  assign n2636 = ~n2485 & ~n2635;
  assign n2637 = n2485 & n2635;
  assign n2638 = ~n2636 & ~n2637;
  assign n2639 = ~n2484 & n2638;
  assign n2640 = n2484 & ~n2638;
  assign n2641 = ~n2639 & ~n2640;
  assign n2642 = ~n2466 & n2641;
  assign n2643 = n2466 & ~n2641;
  assign po25  = ~n2642 & ~n2643;
  assign n2645 = ~n2639 & ~n2642;
  assign n2646 = ~n2621 & ~n2632;
  assign n2647 = ~n2636 & ~n2646;
  assign n2648 = ~n2594 & ~n2600;
  assign n2649 = ~n2577 & ~n2580;
  assign n2650 = ~n2557 & ~n2563;
  assign n2651 = n809 & n1297;
  assign n2652 = pi73  & n1366;
  assign n2653 = pi75  & n1295;
  assign n2654 = pi74  & n1290;
  assign n2655 = ~n2653 & ~n2654;
  assign n2656 = ~n2652 & n2655;
  assign n2657 = ~n2651 & n2656;
  assign n2658 = pi17  & ~n2657;
  assign n2659 = pi17  & ~n2658;
  assign n2660 = ~n2657 & ~n2658;
  assign n2661 = ~n2659 & ~n2660;
  assign n2662 = ~n2540 & ~n2543;
  assign n2663 = ~n2511 & n2533;
  assign n2664 = ~n2537 & ~n2663;
  assign n2665 = n286 & n2523;
  assign n2666 = n2336 & n2515;
  assign n2667 = ~n2520 & n2666;
  assign n2668 = pi64  & n2667;
  assign n2669 = pi66  & n2521;
  assign n2670 = pi65  & n2516;
  assign n2671 = ~n2669 & ~n2670;
  assign n2672 = ~n2665 & n2671;
  assign n2673 = ~n2668 & n2672;
  assign n2674 = pi26  & ~n2673;
  assign n2675 = pi26  & ~n2674;
  assign n2676 = ~n2673 & ~n2674;
  assign n2677 = ~n2675 & ~n2676;
  assign n2678 = ~n2531 & n2677;
  assign n2679 = n2531 & ~n2677;
  assign n2680 = ~n2678 & ~n2679;
  assign n2681 = n401 & n2043;
  assign n2682 = pi67  & n2180;
  assign n2683 = pi69  & n2041;
  assign n2684 = pi68  & n2036;
  assign n2685 = ~n2683 & ~n2684;
  assign n2686 = ~n2682 & n2685;
  assign n2687 = ~n2681 & n2686;
  assign n2688 = pi23  & ~n2687;
  assign n2689 = pi23  & ~n2688;
  assign n2690 = ~n2687 & ~n2688;
  assign n2691 = ~n2689 & ~n2690;
  assign n2692 = n2680 & ~n2691;
  assign n2693 = ~n2680 & n2691;
  assign n2694 = ~n2692 & ~n2693;
  assign n2695 = ~n2664 & n2694;
  assign n2696 = ~n2664 & ~n2695;
  assign n2697 = ~n2692 & ~n2695;
  assign n2698 = ~n2693 & n2697;
  assign n2699 = ~n2696 & ~n2698;
  assign n2700 = n576 & n1611;
  assign n2701 = pi70  & n1745;
  assign n2702 = pi72  & n1609;
  assign n2703 = pi71  & n1604;
  assign n2704 = ~n2702 & ~n2703;
  assign n2705 = ~n2701 & n2704;
  assign n2706 = ~n2700 & n2705;
  assign n2707 = pi20  & ~n2706;
  assign n2708 = pi20  & ~n2707;
  assign n2709 = ~n2706 & ~n2707;
  assign n2710 = ~n2708 & ~n2709;
  assign n2711 = n2699 & n2710;
  assign n2712 = ~n2699 & ~n2710;
  assign n2713 = ~n2711 & ~n2712;
  assign n2714 = ~n2662 & n2713;
  assign n2715 = n2662 & ~n2713;
  assign n2716 = ~n2714 & ~n2715;
  assign n2717 = n2661 & ~n2716;
  assign n2718 = ~n2661 & n2716;
  assign n2719 = ~n2717 & ~n2718;
  assign n2720 = ~n2650 & n2719;
  assign n2721 = n2650 & ~n2719;
  assign n2722 = ~n2720 & ~n2721;
  assign n2723 = n938 & n1025;
  assign n2724 = pi76  & n1052;
  assign n2725 = pi78  & n936;
  assign n2726 = pi77  & n931;
  assign n2727 = ~n2725 & ~n2726;
  assign n2728 = ~n2724 & n2727;
  assign n2729 = ~n2723 & n2728;
  assign n2730 = pi14  & ~n2729;
  assign n2731 = pi14  & ~n2730;
  assign n2732 = ~n2729 & ~n2730;
  assign n2733 = ~n2731 & ~n2732;
  assign n2734 = n2722 & ~n2733;
  assign n2735 = n2722 & ~n2734;
  assign n2736 = ~n2733 & ~n2734;
  assign n2737 = ~n2735 & ~n2736;
  assign n2738 = ~n2649 & n2737;
  assign n2739 = n2649 & ~n2737;
  assign n2740 = ~n2738 & ~n2739;
  assign n2741 = n687 & n1434;
  assign n2742 = pi79  & n763;
  assign n2743 = pi81  & n685;
  assign n2744 = pi80  & n680;
  assign n2745 = ~n2743 & ~n2744;
  assign n2746 = ~n2742 & n2745;
  assign n2747 = ~n2741 & n2746;
  assign n2748 = pi11  & ~n2747;
  assign n2749 = pi11  & ~n2748;
  assign n2750 = ~n2747 & ~n2748;
  assign n2751 = ~n2749 & ~n2750;
  assign n2752 = ~n2740 & ~n2751;
  assign n2753 = n2740 & n2751;
  assign n2754 = ~n2752 & ~n2753;
  assign n2755 = n2648 & ~n2754;
  assign n2756 = ~n2648 & n2754;
  assign n2757 = ~n2755 & ~n2756;
  assign n2758 = n498 & n1834;
  assign n2759 = pi82  & n537;
  assign n2760 = pi84  & n496;
  assign n2761 = pi83  & n491;
  assign n2762 = ~n2760 & ~n2761;
  assign n2763 = ~n2759 & n2762;
  assign n2764 = ~n2758 & n2763;
  assign n2765 = pi8  & ~n2764;
  assign n2766 = pi8  & ~n2765;
  assign n2767 = ~n2764 & ~n2765;
  assign n2768 = ~n2766 & ~n2767;
  assign n2769 = n2757 & ~n2768;
  assign n2770 = n2757 & ~n2769;
  assign n2771 = ~n2768 & ~n2769;
  assign n2772 = ~n2770 & ~n2771;
  assign n2773 = ~n2613 & ~n2618;
  assign n2774 = n2772 & n2773;
  assign n2775 = ~n2772 & ~n2773;
  assign n2776 = ~n2774 & ~n2775;
  assign n2777 = n342 & n2288;
  assign n2778 = pi85  & n380;
  assign n2779 = pi87  & n340;
  assign n2780 = pi86  & n335;
  assign n2781 = ~n2779 & ~n2780;
  assign n2782 = ~n2778 & n2781;
  assign n2783 = ~n2777 & n2782;
  assign n2784 = pi5  & ~n2783;
  assign n2785 = pi5  & ~n2784;
  assign n2786 = ~n2783 & ~n2784;
  assign n2787 = ~n2785 & ~n2786;
  assign n2788 = n2776 & ~n2787;
  assign n2789 = n2776 & ~n2788;
  assign n2790 = ~n2787 & ~n2788;
  assign n2791 = ~n2789 & ~n2790;
  assign n2792 = ~n2647 & n2791;
  assign n2793 = n2647 & ~n2791;
  assign n2794 = ~n2792 & ~n2793;
  assign n2795 = ~n2469 & ~n2471;
  assign n2796 = ~pi89  & ~pi90 ;
  assign n2797 = pi89  & pi90 ;
  assign n2798 = ~n2796 & ~n2797;
  assign n2799 = ~n2795 & n2798;
  assign n2800 = n2795 & ~n2798;
  assign n2801 = ~n2799 & ~n2800;
  assign n2802 = n262 & n2801;
  assign n2803 = pi88  & n288;
  assign n2804 = pi90  & n267;
  assign n2805 = pi89  & n269;
  assign n2806 = ~n2804 & ~n2805;
  assign n2807 = ~n2803 & n2806;
  assign n2808 = ~n2802 & n2807;
  assign n2809 = pi2  & ~n2808;
  assign n2810 = pi2  & ~n2809;
  assign n2811 = ~n2808 & ~n2809;
  assign n2812 = ~n2810 & ~n2811;
  assign n2813 = ~n2794 & ~n2812;
  assign n2814 = n2794 & n2812;
  assign n2815 = ~n2813 & ~n2814;
  assign n2816 = ~n2645 & n2815;
  assign n2817 = n2645 & ~n2815;
  assign po26  = ~n2816 & ~n2817;
  assign n2819 = ~n2813 & ~n2816;
  assign n2820 = ~n2718 & ~n2720;
  assign n2821 = n891 & n1297;
  assign n2822 = pi74  & n1366;
  assign n2823 = pi76  & n1295;
  assign n2824 = pi75  & n1290;
  assign n2825 = ~n2823 & ~n2824;
  assign n2826 = ~n2822 & n2825;
  assign n2827 = ~n2821 & n2826;
  assign n2828 = pi17  & ~n2827;
  assign n2829 = pi17  & ~n2828;
  assign n2830 = ~n2827 & ~n2828;
  assign n2831 = ~n2829 & ~n2830;
  assign n2832 = ~n2712 & ~n2714;
  assign n2833 = pi26  & ~pi27 ;
  assign n2834 = ~pi26  & pi27 ;
  assign n2835 = ~n2833 & ~n2834;
  assign n2836 = pi64  & ~n2835;
  assign n2837 = ~n2679 & n2836;
  assign n2838 = n2679 & ~n2836;
  assign n2839 = ~n2837 & ~n2838;
  assign n2840 = n309 & n2523;
  assign n2841 = pi65  & n2667;
  assign n2842 = pi67  & n2521;
  assign n2843 = pi66  & n2516;
  assign n2844 = ~n2842 & ~n2843;
  assign n2845 = ~n2841 & n2844;
  assign n2846 = ~n2840 & n2845;
  assign n2847 = pi26  & ~n2846;
  assign n2848 = pi26  & ~n2847;
  assign n2849 = ~n2846 & ~n2847;
  assign n2850 = ~n2848 & ~n2849;
  assign n2851 = ~n2839 & ~n2850;
  assign n2852 = n2839 & n2850;
  assign n2853 = ~n2851 & ~n2852;
  assign n2854 = n450 & n2043;
  assign n2855 = pi68  & n2180;
  assign n2856 = pi70  & n2041;
  assign n2857 = pi69  & n2036;
  assign n2858 = ~n2856 & ~n2857;
  assign n2859 = ~n2855 & n2858;
  assign n2860 = ~n2854 & n2859;
  assign n2861 = pi23  & ~n2860;
  assign n2862 = pi23  & ~n2861;
  assign n2863 = ~n2860 & ~n2861;
  assign n2864 = ~n2862 & ~n2863;
  assign n2865 = n2853 & ~n2864;
  assign n2866 = n2853 & ~n2865;
  assign n2867 = ~n2864 & ~n2865;
  assign n2868 = ~n2866 & ~n2867;
  assign n2869 = ~n2697 & n2868;
  assign n2870 = n2697 & ~n2868;
  assign n2871 = ~n2869 & ~n2870;
  assign n2872 = n642 & n1611;
  assign n2873 = pi71  & n1745;
  assign n2874 = pi73  & n1609;
  assign n2875 = pi72  & n1604;
  assign n2876 = ~n2874 & ~n2875;
  assign n2877 = ~n2873 & n2876;
  assign n2878 = ~n2872 & n2877;
  assign n2879 = pi20  & ~n2878;
  assign n2880 = pi20  & ~n2879;
  assign n2881 = ~n2878 & ~n2879;
  assign n2882 = ~n2880 & ~n2881;
  assign n2883 = ~n2871 & ~n2882;
  assign n2884 = n2871 & n2882;
  assign n2885 = ~n2883 & ~n2884;
  assign n2886 = ~n2832 & n2885;
  assign n2887 = n2832 & ~n2885;
  assign n2888 = ~n2886 & ~n2887;
  assign n2889 = n2831 & ~n2888;
  assign n2890 = ~n2831 & n2888;
  assign n2891 = ~n2889 & ~n2890;
  assign n2892 = ~n2820 & n2891;
  assign n2893 = n2820 & ~n2891;
  assign n2894 = ~n2892 & ~n2893;
  assign n2895 = n938 & n1122;
  assign n2896 = pi77  & n1052;
  assign n2897 = pi79  & n936;
  assign n2898 = pi78  & n931;
  assign n2899 = ~n2897 & ~n2898;
  assign n2900 = ~n2896 & n2899;
  assign n2901 = ~n2895 & n2900;
  assign n2902 = pi14  & ~n2901;
  assign n2903 = pi14  & ~n2902;
  assign n2904 = ~n2901 & ~n2902;
  assign n2905 = ~n2903 & ~n2904;
  assign n2906 = n2894 & ~n2905;
  assign n2907 = n2894 & ~n2906;
  assign n2908 = ~n2905 & ~n2906;
  assign n2909 = ~n2907 & ~n2908;
  assign n2910 = ~n2649 & ~n2737;
  assign n2911 = ~n2734 & ~n2910;
  assign n2912 = n2909 & n2911;
  assign n2913 = ~n2909 & ~n2911;
  assign n2914 = ~n2912 & ~n2913;
  assign n2915 = n687 & n1554;
  assign n2916 = pi80  & n763;
  assign n2917 = pi82  & n685;
  assign n2918 = pi81  & n680;
  assign n2919 = ~n2917 & ~n2918;
  assign n2920 = ~n2916 & n2919;
  assign n2921 = ~n2915 & n2920;
  assign n2922 = pi11  & ~n2921;
  assign n2923 = pi11  & ~n2922;
  assign n2924 = ~n2921 & ~n2922;
  assign n2925 = ~n2923 & ~n2924;
  assign n2926 = n2914 & ~n2925;
  assign n2927 = n2914 & ~n2926;
  assign n2928 = ~n2925 & ~n2926;
  assign n2929 = ~n2927 & ~n2928;
  assign n2930 = ~n2752 & ~n2756;
  assign n2931 = n2929 & n2930;
  assign n2932 = ~n2929 & ~n2930;
  assign n2933 = ~n2931 & ~n2932;
  assign n2934 = n498 & n1972;
  assign n2935 = pi83  & n537;
  assign n2936 = pi85  & n496;
  assign n2937 = pi84  & n491;
  assign n2938 = ~n2936 & ~n2937;
  assign n2939 = ~n2935 & n2938;
  assign n2940 = ~n2934 & n2939;
  assign n2941 = pi8  & ~n2940;
  assign n2942 = pi8  & ~n2941;
  assign n2943 = ~n2940 & ~n2941;
  assign n2944 = ~n2942 & ~n2943;
  assign n2945 = ~n2933 & n2944;
  assign n2946 = n2933 & ~n2944;
  assign n2947 = ~n2945 & ~n2946;
  assign n2948 = ~n2769 & ~n2775;
  assign n2949 = n2947 & ~n2948;
  assign n2950 = ~n2947 & n2948;
  assign n2951 = ~n2949 & ~n2950;
  assign n2952 = n342 & n2446;
  assign n2953 = pi86  & n380;
  assign n2954 = pi88  & n340;
  assign n2955 = pi87  & n335;
  assign n2956 = ~n2954 & ~n2955;
  assign n2957 = ~n2953 & n2956;
  assign n2958 = ~n2952 & n2957;
  assign n2959 = pi5  & ~n2958;
  assign n2960 = pi5  & ~n2959;
  assign n2961 = ~n2958 & ~n2959;
  assign n2962 = ~n2960 & ~n2961;
  assign n2963 = n2951 & ~n2962;
  assign n2964 = n2951 & ~n2963;
  assign n2965 = ~n2962 & ~n2963;
  assign n2966 = ~n2964 & ~n2965;
  assign n2967 = ~n2647 & ~n2791;
  assign n2968 = ~n2788 & ~n2967;
  assign n2969 = n2966 & n2968;
  assign n2970 = ~n2966 & ~n2968;
  assign n2971 = ~n2969 & ~n2970;
  assign n2972 = ~n2797 & ~n2799;
  assign n2973 = ~pi90  & ~pi91 ;
  assign n2974 = pi90  & pi91 ;
  assign n2975 = ~n2973 & ~n2974;
  assign n2976 = ~n2972 & n2975;
  assign n2977 = n2972 & ~n2975;
  assign n2978 = ~n2976 & ~n2977;
  assign n2979 = n262 & n2978;
  assign n2980 = pi89  & n288;
  assign n2981 = pi91  & n267;
  assign n2982 = pi90  & n269;
  assign n2983 = ~n2981 & ~n2982;
  assign n2984 = ~n2980 & n2983;
  assign n2985 = ~n2979 & n2984;
  assign n2986 = pi2  & ~n2985;
  assign n2987 = pi2  & ~n2986;
  assign n2988 = ~n2985 & ~n2986;
  assign n2989 = ~n2987 & ~n2988;
  assign n2990 = ~n2971 & n2989;
  assign n2991 = n2971 & ~n2989;
  assign n2992 = ~n2990 & ~n2991;
  assign n2993 = ~n2819 & n2992;
  assign n2994 = n2819 & ~n2992;
  assign po27  = ~n2993 & ~n2994;
  assign n2996 = ~n2991 & ~n2993;
  assign n2997 = ~n2697 & ~n2868;
  assign n2998 = ~n2865 & ~n2997;
  assign n2999 = n475 & n2043;
  assign n3000 = pi69  & n2180;
  assign n3001 = pi71  & n2041;
  assign n3002 = pi70  & n2036;
  assign n3003 = ~n3001 & ~n3002;
  assign n3004 = ~n3000 & n3003;
  assign n3005 = ~n2999 & n3004;
  assign n3006 = pi23  & ~n3005;
  assign n3007 = pi23  & ~n3006;
  assign n3008 = ~n3005 & ~n3006;
  assign n3009 = ~n3007 & ~n3008;
  assign n3010 = n2679 & n2836;
  assign n3011 = ~n2851 & ~n3010;
  assign n3012 = n359 & n2523;
  assign n3013 = pi66  & n2667;
  assign n3014 = pi68  & n2521;
  assign n3015 = pi67  & n2516;
  assign n3016 = ~n3014 & ~n3015;
  assign n3017 = ~n3013 & n3016;
  assign n3018 = ~n3012 & n3017;
  assign n3019 = pi26  & ~n3018;
  assign n3020 = pi26  & ~n3019;
  assign n3021 = ~n3018 & ~n3019;
  assign n3022 = ~n3020 & ~n3021;
  assign n3023 = pi29  & ~n2836;
  assign n3024 = ~pi27  & pi28 ;
  assign n3025 = pi27  & ~pi28 ;
  assign n3026 = ~n3024 & ~n3025;
  assign n3027 = n2835 & ~n3026;
  assign n3028 = pi64  & n3027;
  assign n3029 = ~pi28  & pi29 ;
  assign n3030 = pi28  & ~pi29 ;
  assign n3031 = ~n3029 & ~n3030;
  assign n3032 = ~n2835 & n3031;
  assign n3033 = pi65  & n3032;
  assign n3034 = ~n2835 & ~n3031;
  assign n3035 = ~n265 & n3034;
  assign n3036 = ~n3028 & ~n3033;
  assign n3037 = ~n3035 & n3036;
  assign n3038 = pi29  & ~n3037;
  assign n3039 = pi29  & ~n3038;
  assign n3040 = ~n3037 & ~n3038;
  assign n3041 = ~n3039 & ~n3040;
  assign n3042 = n3023 & ~n3041;
  assign n3043 = ~n3023 & n3041;
  assign n3044 = ~n3042 & ~n3043;
  assign n3045 = n3022 & n3044;
  assign n3046 = ~n3022 & ~n3044;
  assign n3047 = ~n3045 & ~n3046;
  assign n3048 = ~n3011 & ~n3047;
  assign n3049 = n3011 & n3047;
  assign n3050 = ~n3048 & ~n3049;
  assign n3051 = ~n3009 & n3050;
  assign n3052 = n3009 & ~n3050;
  assign n3053 = ~n3051 & ~n3052;
  assign n3054 = ~n2998 & n3053;
  assign n3055 = n2998 & ~n3053;
  assign n3056 = ~n3054 & ~n3055;
  assign n3057 = n729 & n1611;
  assign n3058 = pi72  & n1745;
  assign n3059 = pi74  & n1609;
  assign n3060 = pi73  & n1604;
  assign n3061 = ~n3059 & ~n3060;
  assign n3062 = ~n3058 & n3061;
  assign n3063 = ~n3057 & n3062;
  assign n3064 = pi20  & ~n3063;
  assign n3065 = pi20  & ~n3064;
  assign n3066 = ~n3063 & ~n3064;
  assign n3067 = ~n3065 & ~n3066;
  assign n3068 = n3056 & ~n3067;
  assign n3069 = n3056 & ~n3068;
  assign n3070 = ~n3067 & ~n3068;
  assign n3071 = ~n3069 & ~n3070;
  assign n3072 = ~n2883 & ~n2886;
  assign n3073 = n3071 & n3072;
  assign n3074 = ~n3071 & ~n3072;
  assign n3075 = ~n3073 & ~n3074;
  assign n3076 = n999 & n1297;
  assign n3077 = pi75  & n1366;
  assign n3078 = pi77  & n1295;
  assign n3079 = pi76  & n1290;
  assign n3080 = ~n3078 & ~n3079;
  assign n3081 = ~n3077 & n3080;
  assign n3082 = ~n3076 & n3081;
  assign n3083 = pi17  & ~n3082;
  assign n3084 = pi17  & ~n3083;
  assign n3085 = ~n3082 & ~n3083;
  assign n3086 = ~n3084 & ~n3085;
  assign n3087 = n3075 & ~n3086;
  assign n3088 = n3075 & ~n3087;
  assign n3089 = ~n3086 & ~n3087;
  assign n3090 = ~n3088 & ~n3089;
  assign n3091 = ~n2890 & ~n2892;
  assign n3092 = ~n3090 & ~n3091;
  assign n3093 = ~n3090 & ~n3092;
  assign n3094 = ~n3091 & ~n3092;
  assign n3095 = ~n3093 & ~n3094;
  assign n3096 = n938 & n1225;
  assign n3097 = pi78  & n1052;
  assign n3098 = pi80  & n936;
  assign n3099 = pi79  & n931;
  assign n3100 = ~n3098 & ~n3099;
  assign n3101 = ~n3097 & n3100;
  assign n3102 = ~n3096 & n3101;
  assign n3103 = pi14  & ~n3102;
  assign n3104 = pi14  & ~n3103;
  assign n3105 = ~n3102 & ~n3103;
  assign n3106 = ~n3104 & ~n3105;
  assign n3107 = ~n3095 & ~n3106;
  assign n3108 = ~n3095 & ~n3107;
  assign n3109 = ~n3106 & ~n3107;
  assign n3110 = ~n3108 & ~n3109;
  assign n3111 = ~n2906 & ~n2913;
  assign n3112 = n3110 & n3111;
  assign n3113 = ~n3110 & ~n3111;
  assign n3114 = ~n3112 & ~n3113;
  assign n3115 = n687 & n1696;
  assign n3116 = pi81  & n763;
  assign n3117 = pi83  & n685;
  assign n3118 = pi82  & n680;
  assign n3119 = ~n3117 & ~n3118;
  assign n3120 = ~n3116 & n3119;
  assign n3121 = ~n3115 & n3120;
  assign n3122 = pi11  & ~n3121;
  assign n3123 = pi11  & ~n3122;
  assign n3124 = ~n3121 & ~n3122;
  assign n3125 = ~n3123 & ~n3124;
  assign n3126 = n3114 & ~n3125;
  assign n3127 = n3114 & ~n3126;
  assign n3128 = ~n3125 & ~n3126;
  assign n3129 = ~n3127 & ~n3128;
  assign n3130 = ~n2926 & ~n2932;
  assign n3131 = n3129 & n3130;
  assign n3132 = ~n3129 & ~n3130;
  assign n3133 = ~n3131 & ~n3132;
  assign n3134 = n498 & n2133;
  assign n3135 = pi84  & n537;
  assign n3136 = pi86  & n496;
  assign n3137 = pi85  & n491;
  assign n3138 = ~n3136 & ~n3137;
  assign n3139 = ~n3135 & n3138;
  assign n3140 = ~n3134 & n3139;
  assign n3141 = pi8  & ~n3140;
  assign n3142 = pi8  & ~n3141;
  assign n3143 = ~n3140 & ~n3141;
  assign n3144 = ~n3142 & ~n3143;
  assign n3145 = ~n3133 & n3144;
  assign n3146 = n3133 & ~n3144;
  assign n3147 = ~n3145 & ~n3146;
  assign n3148 = ~n2946 & ~n2949;
  assign n3149 = n3147 & ~n3148;
  assign n3150 = ~n3147 & n3148;
  assign n3151 = ~n3149 & ~n3150;
  assign n3152 = n342 & n2473;
  assign n3153 = pi87  & n380;
  assign n3154 = pi89  & n340;
  assign n3155 = pi88  & n335;
  assign n3156 = ~n3154 & ~n3155;
  assign n3157 = ~n3153 & n3156;
  assign n3158 = ~n3152 & n3157;
  assign n3159 = pi5  & ~n3158;
  assign n3160 = pi5  & ~n3159;
  assign n3161 = ~n3158 & ~n3159;
  assign n3162 = ~n3160 & ~n3161;
  assign n3163 = n3151 & ~n3162;
  assign n3164 = n3151 & ~n3163;
  assign n3165 = ~n3162 & ~n3163;
  assign n3166 = ~n3164 & ~n3165;
  assign n3167 = ~n2963 & ~n2970;
  assign n3168 = n3166 & n3167;
  assign n3169 = ~n3166 & ~n3167;
  assign n3170 = ~n3168 & ~n3169;
  assign n3171 = ~n2974 & ~n2976;
  assign n3172 = ~pi91  & ~pi92 ;
  assign n3173 = pi91  & pi92 ;
  assign n3174 = ~n3172 & ~n3173;
  assign n3175 = ~n3171 & n3174;
  assign n3176 = n3171 & ~n3174;
  assign n3177 = ~n3175 & ~n3176;
  assign n3178 = n262 & n3177;
  assign n3179 = pi90  & n288;
  assign n3180 = pi92  & n267;
  assign n3181 = pi91  & n269;
  assign n3182 = ~n3180 & ~n3181;
  assign n3183 = ~n3179 & n3182;
  assign n3184 = ~n3178 & n3183;
  assign n3185 = pi2  & ~n3184;
  assign n3186 = pi2  & ~n3185;
  assign n3187 = ~n3184 & ~n3185;
  assign n3188 = ~n3186 & ~n3187;
  assign n3189 = ~n3170 & n3188;
  assign n3190 = n3170 & ~n3188;
  assign n3191 = ~n3189 & ~n3190;
  assign n3192 = ~n2996 & n3191;
  assign n3193 = n2996 & ~n3191;
  assign po28  = ~n3192 & ~n3193;
  assign n3195 = ~n3163 & ~n3169;
  assign n3196 = n342 & n2801;
  assign n3197 = pi88  & n380;
  assign n3198 = pi90  & n340;
  assign n3199 = pi89  & n335;
  assign n3200 = ~n3198 & ~n3199;
  assign n3201 = ~n3197 & n3200;
  assign n3202 = ~n3196 & n3201;
  assign n3203 = pi5  & ~n3202;
  assign n3204 = pi5  & ~n3203;
  assign n3205 = ~n3202 & ~n3203;
  assign n3206 = ~n3204 & ~n3205;
  assign n3207 = ~n3126 & ~n3132;
  assign n3208 = ~n3068 & ~n3074;
  assign n3209 = n809 & n1611;
  assign n3210 = pi73  & n1745;
  assign n3211 = pi75  & n1609;
  assign n3212 = pi74  & n1604;
  assign n3213 = ~n3211 & ~n3212;
  assign n3214 = ~n3210 & n3213;
  assign n3215 = ~n3209 & n3214;
  assign n3216 = pi20  & ~n3215;
  assign n3217 = pi20  & ~n3216;
  assign n3218 = ~n3215 & ~n3216;
  assign n3219 = ~n3217 & ~n3218;
  assign n3220 = ~n3051 & ~n3054;
  assign n3221 = ~n3022 & n3044;
  assign n3222 = ~n3048 & ~n3221;
  assign n3223 = n286 & n3034;
  assign n3224 = n2835 & n3026;
  assign n3225 = ~n3031 & n3224;
  assign n3226 = pi64  & n3225;
  assign n3227 = pi66  & n3032;
  assign n3228 = pi65  & n3027;
  assign n3229 = ~n3227 & ~n3228;
  assign n3230 = ~n3223 & n3229;
  assign n3231 = ~n3226 & n3230;
  assign n3232 = pi29  & ~n3231;
  assign n3233 = pi29  & ~n3232;
  assign n3234 = ~n3231 & ~n3232;
  assign n3235 = ~n3233 & ~n3234;
  assign n3236 = ~n3042 & n3235;
  assign n3237 = n3042 & ~n3235;
  assign n3238 = ~n3236 & ~n3237;
  assign n3239 = n401 & n2523;
  assign n3240 = pi67  & n2667;
  assign n3241 = pi69  & n2521;
  assign n3242 = pi68  & n2516;
  assign n3243 = ~n3241 & ~n3242;
  assign n3244 = ~n3240 & n3243;
  assign n3245 = ~n3239 & n3244;
  assign n3246 = pi26  & ~n3245;
  assign n3247 = pi26  & ~n3246;
  assign n3248 = ~n3245 & ~n3246;
  assign n3249 = ~n3247 & ~n3248;
  assign n3250 = n3238 & ~n3249;
  assign n3251 = ~n3238 & n3249;
  assign n3252 = ~n3250 & ~n3251;
  assign n3253 = ~n3222 & n3252;
  assign n3254 = ~n3222 & ~n3253;
  assign n3255 = ~n3250 & ~n3253;
  assign n3256 = ~n3251 & n3255;
  assign n3257 = ~n3254 & ~n3256;
  assign n3258 = n576 & n2043;
  assign n3259 = pi70  & n2180;
  assign n3260 = pi72  & n2041;
  assign n3261 = pi71  & n2036;
  assign n3262 = ~n3260 & ~n3261;
  assign n3263 = ~n3259 & n3262;
  assign n3264 = ~n3258 & n3263;
  assign n3265 = pi23  & ~n3264;
  assign n3266 = pi23  & ~n3265;
  assign n3267 = ~n3264 & ~n3265;
  assign n3268 = ~n3266 & ~n3267;
  assign n3269 = n3257 & n3268;
  assign n3270 = ~n3257 & ~n3268;
  assign n3271 = ~n3269 & ~n3270;
  assign n3272 = ~n3220 & n3271;
  assign n3273 = n3220 & ~n3271;
  assign n3274 = ~n3272 & ~n3273;
  assign n3275 = n3219 & ~n3274;
  assign n3276 = ~n3219 & n3274;
  assign n3277 = ~n3275 & ~n3276;
  assign n3278 = ~n3208 & n3277;
  assign n3279 = n3208 & ~n3277;
  assign n3280 = ~n3278 & ~n3279;
  assign n3281 = n1025 & n1297;
  assign n3282 = pi76  & n1366;
  assign n3283 = pi78  & n1295;
  assign n3284 = pi77  & n1290;
  assign n3285 = ~n3283 & ~n3284;
  assign n3286 = ~n3282 & n3285;
  assign n3287 = ~n3281 & n3286;
  assign n3288 = pi17  & ~n3287;
  assign n3289 = pi17  & ~n3288;
  assign n3290 = ~n3287 & ~n3288;
  assign n3291 = ~n3289 & ~n3290;
  assign n3292 = n3280 & ~n3291;
  assign n3293 = n3280 & ~n3292;
  assign n3294 = ~n3291 & ~n3292;
  assign n3295 = ~n3293 & ~n3294;
  assign n3296 = ~n3087 & ~n3092;
  assign n3297 = n3295 & n3296;
  assign n3298 = ~n3295 & ~n3296;
  assign n3299 = ~n3297 & ~n3298;
  assign n3300 = n938 & n1434;
  assign n3301 = pi79  & n1052;
  assign n3302 = pi81  & n936;
  assign n3303 = pi80  & n931;
  assign n3304 = ~n3302 & ~n3303;
  assign n3305 = ~n3301 & n3304;
  assign n3306 = ~n3300 & n3305;
  assign n3307 = pi14  & ~n3306;
  assign n3308 = pi14  & ~n3307;
  assign n3309 = ~n3306 & ~n3307;
  assign n3310 = ~n3308 & ~n3309;
  assign n3311 = n3299 & ~n3310;
  assign n3312 = n3299 & ~n3311;
  assign n3313 = ~n3310 & ~n3311;
  assign n3314 = ~n3312 & ~n3313;
  assign n3315 = ~n3107 & ~n3113;
  assign n3316 = n3314 & n3315;
  assign n3317 = ~n3314 & ~n3315;
  assign n3318 = ~n3316 & ~n3317;
  assign n3319 = n687 & n1834;
  assign n3320 = pi82  & n763;
  assign n3321 = pi84  & n685;
  assign n3322 = pi83  & n680;
  assign n3323 = ~n3321 & ~n3322;
  assign n3324 = ~n3320 & n3323;
  assign n3325 = ~n3319 & n3324;
  assign n3326 = pi11  & ~n3325;
  assign n3327 = pi11  & ~n3326;
  assign n3328 = ~n3325 & ~n3326;
  assign n3329 = ~n3327 & ~n3328;
  assign n3330 = n3318 & ~n3329;
  assign n3331 = ~n3318 & n3329;
  assign n3332 = ~n3330 & ~n3331;
  assign n3333 = ~n3207 & n3332;
  assign n3334 = ~n3207 & ~n3333;
  assign n3335 = ~n3330 & ~n3333;
  assign n3336 = ~n3331 & n3335;
  assign n3337 = ~n3334 & ~n3336;
  assign n3338 = n498 & n2288;
  assign n3339 = pi85  & n537;
  assign n3340 = pi87  & n496;
  assign n3341 = pi86  & n491;
  assign n3342 = ~n3340 & ~n3341;
  assign n3343 = ~n3339 & n3342;
  assign n3344 = ~n3338 & n3343;
  assign n3345 = pi8  & ~n3344;
  assign n3346 = pi8  & ~n3345;
  assign n3347 = ~n3344 & ~n3345;
  assign n3348 = ~n3346 & ~n3347;
  assign n3349 = ~n3337 & ~n3348;
  assign n3350 = ~n3337 & ~n3349;
  assign n3351 = ~n3348 & ~n3349;
  assign n3352 = ~n3350 & ~n3351;
  assign n3353 = ~n3146 & ~n3149;
  assign n3354 = ~n3352 & ~n3353;
  assign n3355 = n3352 & n3353;
  assign n3356 = ~n3354 & ~n3355;
  assign n3357 = ~n3206 & n3356;
  assign n3358 = ~n3206 & ~n3357;
  assign n3359 = n3356 & ~n3357;
  assign n3360 = ~n3358 & ~n3359;
  assign n3361 = ~n3195 & ~n3360;
  assign n3362 = ~n3195 & ~n3361;
  assign n3363 = ~n3360 & ~n3361;
  assign n3364 = ~n3362 & ~n3363;
  assign n3365 = ~n3173 & ~n3175;
  assign n3366 = ~pi92  & ~pi93 ;
  assign n3367 = pi92  & pi93 ;
  assign n3368 = ~n3366 & ~n3367;
  assign n3369 = ~n3365 & n3368;
  assign n3370 = n3365 & ~n3368;
  assign n3371 = ~n3369 & ~n3370;
  assign n3372 = n262 & n3371;
  assign n3373 = pi91  & n288;
  assign n3374 = pi93  & n267;
  assign n3375 = pi92  & n269;
  assign n3376 = ~n3374 & ~n3375;
  assign n3377 = ~n3373 & n3376;
  assign n3378 = ~n3372 & n3377;
  assign n3379 = pi2  & ~n3378;
  assign n3380 = pi2  & ~n3379;
  assign n3381 = ~n3378 & ~n3379;
  assign n3382 = ~n3380 & ~n3381;
  assign n3383 = ~n3364 & ~n3382;
  assign n3384 = ~n3364 & ~n3383;
  assign n3385 = ~n3382 & ~n3383;
  assign n3386 = ~n3384 & ~n3385;
  assign n3387 = ~n3190 & ~n3192;
  assign n3388 = ~n3386 & ~n3387;
  assign n3389 = n3386 & n3387;
  assign po29  = ~n3388 & ~n3389;
  assign n3391 = ~n3349 & ~n3354;
  assign n3392 = ~n3276 & ~n3278;
  assign n3393 = n891 & n1611;
  assign n3394 = pi74  & n1745;
  assign n3395 = pi76  & n1609;
  assign n3396 = pi75  & n1604;
  assign n3397 = ~n3395 & ~n3396;
  assign n3398 = ~n3394 & n3397;
  assign n3399 = ~n3393 & n3398;
  assign n3400 = pi20  & ~n3399;
  assign n3401 = pi20  & ~n3400;
  assign n3402 = ~n3399 & ~n3400;
  assign n3403 = ~n3401 & ~n3402;
  assign n3404 = ~n3270 & ~n3272;
  assign n3405 = pi29  & ~pi30 ;
  assign n3406 = ~pi29  & pi30 ;
  assign n3407 = ~n3405 & ~n3406;
  assign n3408 = pi64  & ~n3407;
  assign n3409 = ~n3237 & n3408;
  assign n3410 = n3237 & ~n3408;
  assign n3411 = ~n3409 & ~n3410;
  assign n3412 = n309 & n3034;
  assign n3413 = pi65  & n3225;
  assign n3414 = pi67  & n3032;
  assign n3415 = pi66  & n3027;
  assign n3416 = ~n3414 & ~n3415;
  assign n3417 = ~n3413 & n3416;
  assign n3418 = ~n3412 & n3417;
  assign n3419 = pi29  & ~n3418;
  assign n3420 = pi29  & ~n3419;
  assign n3421 = ~n3418 & ~n3419;
  assign n3422 = ~n3420 & ~n3421;
  assign n3423 = ~n3411 & ~n3422;
  assign n3424 = n3411 & n3422;
  assign n3425 = ~n3423 & ~n3424;
  assign n3426 = n450 & n2523;
  assign n3427 = pi68  & n2667;
  assign n3428 = pi70  & n2521;
  assign n3429 = pi69  & n2516;
  assign n3430 = ~n3428 & ~n3429;
  assign n3431 = ~n3427 & n3430;
  assign n3432 = ~n3426 & n3431;
  assign n3433 = pi26  & ~n3432;
  assign n3434 = pi26  & ~n3433;
  assign n3435 = ~n3432 & ~n3433;
  assign n3436 = ~n3434 & ~n3435;
  assign n3437 = n3425 & ~n3436;
  assign n3438 = n3425 & ~n3437;
  assign n3439 = ~n3436 & ~n3437;
  assign n3440 = ~n3438 & ~n3439;
  assign n3441 = ~n3255 & n3440;
  assign n3442 = n3255 & ~n3440;
  assign n3443 = ~n3441 & ~n3442;
  assign n3444 = n642 & n2043;
  assign n3445 = pi71  & n2180;
  assign n3446 = pi73  & n2041;
  assign n3447 = pi72  & n2036;
  assign n3448 = ~n3446 & ~n3447;
  assign n3449 = ~n3445 & n3448;
  assign n3450 = ~n3444 & n3449;
  assign n3451 = pi23  & ~n3450;
  assign n3452 = pi23  & ~n3451;
  assign n3453 = ~n3450 & ~n3451;
  assign n3454 = ~n3452 & ~n3453;
  assign n3455 = ~n3443 & ~n3454;
  assign n3456 = n3443 & n3454;
  assign n3457 = ~n3455 & ~n3456;
  assign n3458 = ~n3404 & n3457;
  assign n3459 = n3404 & ~n3457;
  assign n3460 = ~n3458 & ~n3459;
  assign n3461 = n3403 & ~n3460;
  assign n3462 = ~n3403 & n3460;
  assign n3463 = ~n3461 & ~n3462;
  assign n3464 = ~n3392 & n3463;
  assign n3465 = n3392 & ~n3463;
  assign n3466 = ~n3464 & ~n3465;
  assign n3467 = n1122 & n1297;
  assign n3468 = pi77  & n1366;
  assign n3469 = pi79  & n1295;
  assign n3470 = pi78  & n1290;
  assign n3471 = ~n3469 & ~n3470;
  assign n3472 = ~n3468 & n3471;
  assign n3473 = ~n3467 & n3472;
  assign n3474 = pi17  & ~n3473;
  assign n3475 = pi17  & ~n3474;
  assign n3476 = ~n3473 & ~n3474;
  assign n3477 = ~n3475 & ~n3476;
  assign n3478 = n3466 & ~n3477;
  assign n3479 = n3466 & ~n3478;
  assign n3480 = ~n3477 & ~n3478;
  assign n3481 = ~n3479 & ~n3480;
  assign n3482 = ~n3292 & ~n3298;
  assign n3483 = n3481 & n3482;
  assign n3484 = ~n3481 & ~n3482;
  assign n3485 = ~n3483 & ~n3484;
  assign n3486 = n938 & n1554;
  assign n3487 = pi80  & n1052;
  assign n3488 = pi82  & n936;
  assign n3489 = pi81  & n931;
  assign n3490 = ~n3488 & ~n3489;
  assign n3491 = ~n3487 & n3490;
  assign n3492 = ~n3486 & n3491;
  assign n3493 = pi14  & ~n3492;
  assign n3494 = pi14  & ~n3493;
  assign n3495 = ~n3492 & ~n3493;
  assign n3496 = ~n3494 & ~n3495;
  assign n3497 = n3485 & ~n3496;
  assign n3498 = n3485 & ~n3497;
  assign n3499 = ~n3496 & ~n3497;
  assign n3500 = ~n3498 & ~n3499;
  assign n3501 = ~n3311 & ~n3317;
  assign n3502 = n3500 & n3501;
  assign n3503 = ~n3500 & ~n3501;
  assign n3504 = ~n3502 & ~n3503;
  assign n3505 = n687 & n1972;
  assign n3506 = pi83  & n763;
  assign n3507 = pi85  & n685;
  assign n3508 = pi84  & n680;
  assign n3509 = ~n3507 & ~n3508;
  assign n3510 = ~n3506 & n3509;
  assign n3511 = ~n3505 & n3510;
  assign n3512 = pi11  & ~n3511;
  assign n3513 = pi11  & ~n3512;
  assign n3514 = ~n3511 & ~n3512;
  assign n3515 = ~n3513 & ~n3514;
  assign n3516 = n3504 & ~n3515;
  assign n3517 = n3504 & ~n3516;
  assign n3518 = ~n3515 & ~n3516;
  assign n3519 = ~n3517 & ~n3518;
  assign n3520 = ~n3335 & n3519;
  assign n3521 = n3335 & ~n3519;
  assign n3522 = ~n3520 & ~n3521;
  assign n3523 = n498 & n2446;
  assign n3524 = pi86  & n537;
  assign n3525 = pi88  & n496;
  assign n3526 = pi87  & n491;
  assign n3527 = ~n3525 & ~n3526;
  assign n3528 = ~n3524 & n3527;
  assign n3529 = ~n3523 & n3528;
  assign n3530 = pi8  & ~n3529;
  assign n3531 = pi8  & ~n3530;
  assign n3532 = ~n3529 & ~n3530;
  assign n3533 = ~n3531 & ~n3532;
  assign n3534 = ~n3522 & ~n3533;
  assign n3535 = n3522 & n3533;
  assign n3536 = ~n3534 & ~n3535;
  assign n3537 = n3391 & ~n3536;
  assign n3538 = ~n3391 & n3536;
  assign n3539 = ~n3537 & ~n3538;
  assign n3540 = n342 & n2978;
  assign n3541 = pi89  & n380;
  assign n3542 = pi91  & n340;
  assign n3543 = pi90  & n335;
  assign n3544 = ~n3542 & ~n3543;
  assign n3545 = ~n3541 & n3544;
  assign n3546 = ~n3540 & n3545;
  assign n3547 = pi5  & ~n3546;
  assign n3548 = pi5  & ~n3547;
  assign n3549 = ~n3546 & ~n3547;
  assign n3550 = ~n3548 & ~n3549;
  assign n3551 = n3539 & ~n3550;
  assign n3552 = n3539 & ~n3551;
  assign n3553 = ~n3550 & ~n3551;
  assign n3554 = ~n3552 & ~n3553;
  assign n3555 = ~n3357 & ~n3361;
  assign n3556 = n3554 & n3555;
  assign n3557 = ~n3554 & ~n3555;
  assign n3558 = ~n3556 & ~n3557;
  assign n3559 = ~n3367 & ~n3369;
  assign n3560 = ~pi93  & ~pi94 ;
  assign n3561 = pi93  & pi94 ;
  assign n3562 = ~n3560 & ~n3561;
  assign n3563 = ~n3559 & n3562;
  assign n3564 = n3559 & ~n3562;
  assign n3565 = ~n3563 & ~n3564;
  assign n3566 = n262 & n3565;
  assign n3567 = pi92  & n288;
  assign n3568 = pi94  & n267;
  assign n3569 = pi93  & n269;
  assign n3570 = ~n3568 & ~n3569;
  assign n3571 = ~n3567 & n3570;
  assign n3572 = ~n3566 & n3571;
  assign n3573 = pi2  & ~n3572;
  assign n3574 = pi2  & ~n3573;
  assign n3575 = ~n3572 & ~n3573;
  assign n3576 = ~n3574 & ~n3575;
  assign n3577 = n3558 & ~n3576;
  assign n3578 = n3558 & ~n3577;
  assign n3579 = ~n3576 & ~n3577;
  assign n3580 = ~n3578 & ~n3579;
  assign n3581 = ~n3383 & ~n3388;
  assign n3582 = ~n3580 & ~n3581;
  assign n3583 = n3580 & n3581;
  assign po30  = ~n3582 & ~n3583;
  assign n3585 = ~n3255 & ~n3440;
  assign n3586 = ~n3437 & ~n3585;
  assign n3587 = n475 & n2523;
  assign n3588 = pi69  & n2667;
  assign n3589 = pi71  & n2521;
  assign n3590 = pi70  & n2516;
  assign n3591 = ~n3589 & ~n3590;
  assign n3592 = ~n3588 & n3591;
  assign n3593 = ~n3587 & n3592;
  assign n3594 = pi26  & ~n3593;
  assign n3595 = pi26  & ~n3594;
  assign n3596 = ~n3593 & ~n3594;
  assign n3597 = ~n3595 & ~n3596;
  assign n3598 = n3237 & n3408;
  assign n3599 = ~n3423 & ~n3598;
  assign n3600 = n359 & n3034;
  assign n3601 = pi66  & n3225;
  assign n3602 = pi68  & n3032;
  assign n3603 = pi67  & n3027;
  assign n3604 = ~n3602 & ~n3603;
  assign n3605 = ~n3601 & n3604;
  assign n3606 = ~n3600 & n3605;
  assign n3607 = pi29  & ~n3606;
  assign n3608 = pi29  & ~n3607;
  assign n3609 = ~n3606 & ~n3607;
  assign n3610 = ~n3608 & ~n3609;
  assign n3611 = pi32  & ~n3408;
  assign n3612 = ~pi30  & pi31 ;
  assign n3613 = pi30  & ~pi31 ;
  assign n3614 = ~n3612 & ~n3613;
  assign n3615 = n3407 & ~n3614;
  assign n3616 = pi64  & n3615;
  assign n3617 = ~pi31  & pi32 ;
  assign n3618 = pi31  & ~pi32 ;
  assign n3619 = ~n3617 & ~n3618;
  assign n3620 = ~n3407 & n3619;
  assign n3621 = pi65  & n3620;
  assign n3622 = ~n3407 & ~n3619;
  assign n3623 = ~n265 & n3622;
  assign n3624 = ~n3616 & ~n3621;
  assign n3625 = ~n3623 & n3624;
  assign n3626 = pi32  & ~n3625;
  assign n3627 = pi32  & ~n3626;
  assign n3628 = ~n3625 & ~n3626;
  assign n3629 = ~n3627 & ~n3628;
  assign n3630 = n3611 & ~n3629;
  assign n3631 = ~n3611 & n3629;
  assign n3632 = ~n3630 & ~n3631;
  assign n3633 = n3610 & n3632;
  assign n3634 = ~n3610 & ~n3632;
  assign n3635 = ~n3633 & ~n3634;
  assign n3636 = ~n3599 & ~n3635;
  assign n3637 = n3599 & n3635;
  assign n3638 = ~n3636 & ~n3637;
  assign n3639 = ~n3597 & n3638;
  assign n3640 = n3597 & ~n3638;
  assign n3641 = ~n3639 & ~n3640;
  assign n3642 = ~n3586 & n3641;
  assign n3643 = n3586 & ~n3641;
  assign n3644 = ~n3642 & ~n3643;
  assign n3645 = n729 & n2043;
  assign n3646 = pi72  & n2180;
  assign n3647 = pi74  & n2041;
  assign n3648 = pi73  & n2036;
  assign n3649 = ~n3647 & ~n3648;
  assign n3650 = ~n3646 & n3649;
  assign n3651 = ~n3645 & n3650;
  assign n3652 = pi23  & ~n3651;
  assign n3653 = pi23  & ~n3652;
  assign n3654 = ~n3651 & ~n3652;
  assign n3655 = ~n3653 & ~n3654;
  assign n3656 = n3644 & ~n3655;
  assign n3657 = n3644 & ~n3656;
  assign n3658 = ~n3655 & ~n3656;
  assign n3659 = ~n3657 & ~n3658;
  assign n3660 = ~n3455 & ~n3458;
  assign n3661 = n3659 & n3660;
  assign n3662 = ~n3659 & ~n3660;
  assign n3663 = ~n3661 & ~n3662;
  assign n3664 = n999 & n1611;
  assign n3665 = pi75  & n1745;
  assign n3666 = pi77  & n1609;
  assign n3667 = pi76  & n1604;
  assign n3668 = ~n3666 & ~n3667;
  assign n3669 = ~n3665 & n3668;
  assign n3670 = ~n3664 & n3669;
  assign n3671 = pi20  & ~n3670;
  assign n3672 = pi20  & ~n3671;
  assign n3673 = ~n3670 & ~n3671;
  assign n3674 = ~n3672 & ~n3673;
  assign n3675 = ~n3663 & n3674;
  assign n3676 = n3663 & ~n3674;
  assign n3677 = ~n3675 & ~n3676;
  assign n3678 = ~n3462 & ~n3464;
  assign n3679 = n3677 & ~n3678;
  assign n3680 = ~n3677 & n3678;
  assign n3681 = ~n3679 & ~n3680;
  assign n3682 = n1225 & n1297;
  assign n3683 = pi78  & n1366;
  assign n3684 = pi80  & n1295;
  assign n3685 = pi79  & n1290;
  assign n3686 = ~n3684 & ~n3685;
  assign n3687 = ~n3683 & n3686;
  assign n3688 = ~n3682 & n3687;
  assign n3689 = pi17  & ~n3688;
  assign n3690 = pi17  & ~n3689;
  assign n3691 = ~n3688 & ~n3689;
  assign n3692 = ~n3690 & ~n3691;
  assign n3693 = n3681 & ~n3692;
  assign n3694 = n3681 & ~n3693;
  assign n3695 = ~n3692 & ~n3693;
  assign n3696 = ~n3694 & ~n3695;
  assign n3697 = ~n3478 & ~n3484;
  assign n3698 = n3696 & n3697;
  assign n3699 = ~n3696 & ~n3697;
  assign n3700 = ~n3698 & ~n3699;
  assign n3701 = n938 & n1696;
  assign n3702 = pi81  & n1052;
  assign n3703 = pi83  & n936;
  assign n3704 = pi82  & n931;
  assign n3705 = ~n3703 & ~n3704;
  assign n3706 = ~n3702 & n3705;
  assign n3707 = ~n3701 & n3706;
  assign n3708 = pi14  & ~n3707;
  assign n3709 = pi14  & ~n3708;
  assign n3710 = ~n3707 & ~n3708;
  assign n3711 = ~n3709 & ~n3710;
  assign n3712 = n3700 & ~n3711;
  assign n3713 = n3700 & ~n3712;
  assign n3714 = ~n3711 & ~n3712;
  assign n3715 = ~n3713 & ~n3714;
  assign n3716 = ~n3497 & ~n3503;
  assign n3717 = n3715 & n3716;
  assign n3718 = ~n3715 & ~n3716;
  assign n3719 = ~n3717 & ~n3718;
  assign n3720 = n687 & n2133;
  assign n3721 = pi84  & n763;
  assign n3722 = pi86  & n685;
  assign n3723 = pi85  & n680;
  assign n3724 = ~n3722 & ~n3723;
  assign n3725 = ~n3721 & n3724;
  assign n3726 = ~n3720 & n3725;
  assign n3727 = pi11  & ~n3726;
  assign n3728 = pi11  & ~n3727;
  assign n3729 = ~n3726 & ~n3727;
  assign n3730 = ~n3728 & ~n3729;
  assign n3731 = n3719 & ~n3730;
  assign n3732 = n3719 & ~n3731;
  assign n3733 = ~n3730 & ~n3731;
  assign n3734 = ~n3732 & ~n3733;
  assign n3735 = ~n3335 & ~n3519;
  assign n3736 = ~n3516 & ~n3735;
  assign n3737 = n3734 & n3736;
  assign n3738 = ~n3734 & ~n3736;
  assign n3739 = ~n3737 & ~n3738;
  assign n3740 = n498 & n2473;
  assign n3741 = pi87  & n537;
  assign n3742 = pi89  & n496;
  assign n3743 = pi88  & n491;
  assign n3744 = ~n3742 & ~n3743;
  assign n3745 = ~n3741 & n3744;
  assign n3746 = ~n3740 & n3745;
  assign n3747 = pi8  & ~n3746;
  assign n3748 = pi8  & ~n3747;
  assign n3749 = ~n3746 & ~n3747;
  assign n3750 = ~n3748 & ~n3749;
  assign n3751 = n3739 & ~n3750;
  assign n3752 = n3739 & ~n3751;
  assign n3753 = ~n3750 & ~n3751;
  assign n3754 = ~n3752 & ~n3753;
  assign n3755 = ~n3534 & ~n3538;
  assign n3756 = n3754 & n3755;
  assign n3757 = ~n3754 & ~n3755;
  assign n3758 = ~n3756 & ~n3757;
  assign n3759 = n342 & n3177;
  assign n3760 = pi90  & n380;
  assign n3761 = pi92  & n340;
  assign n3762 = pi91  & n335;
  assign n3763 = ~n3761 & ~n3762;
  assign n3764 = ~n3760 & n3763;
  assign n3765 = ~n3759 & n3764;
  assign n3766 = pi5  & ~n3765;
  assign n3767 = pi5  & ~n3766;
  assign n3768 = ~n3765 & ~n3766;
  assign n3769 = ~n3767 & ~n3768;
  assign n3770 = n3758 & ~n3769;
  assign n3771 = n3758 & ~n3770;
  assign n3772 = ~n3769 & ~n3770;
  assign n3773 = ~n3771 & ~n3772;
  assign n3774 = ~n3551 & ~n3557;
  assign n3775 = n3773 & n3774;
  assign n3776 = ~n3773 & ~n3774;
  assign n3777 = ~n3775 & ~n3776;
  assign n3778 = ~n3561 & ~n3563;
  assign n3779 = ~pi94  & ~pi95 ;
  assign n3780 = pi94  & pi95 ;
  assign n3781 = ~n3779 & ~n3780;
  assign n3782 = ~n3778 & n3781;
  assign n3783 = n3778 & ~n3781;
  assign n3784 = ~n3782 & ~n3783;
  assign n3785 = n262 & n3784;
  assign n3786 = pi93  & n288;
  assign n3787 = pi95  & n267;
  assign n3788 = pi94  & n269;
  assign n3789 = ~n3787 & ~n3788;
  assign n3790 = ~n3786 & n3789;
  assign n3791 = ~n3785 & n3790;
  assign n3792 = pi2  & ~n3791;
  assign n3793 = pi2  & ~n3792;
  assign n3794 = ~n3791 & ~n3792;
  assign n3795 = ~n3793 & ~n3794;
  assign n3796 = n3777 & ~n3795;
  assign n3797 = n3777 & ~n3796;
  assign n3798 = ~n3795 & ~n3796;
  assign n3799 = ~n3797 & ~n3798;
  assign n3800 = ~n3577 & ~n3582;
  assign n3801 = ~n3799 & ~n3800;
  assign n3802 = n3799 & n3800;
  assign po31  = ~n3801 & ~n3802;
  assign n3804 = ~n3796 & ~n3801;
  assign n3805 = ~n3770 & ~n3776;
  assign n3806 = ~n3731 & ~n3738;
  assign n3807 = ~n3712 & ~n3718;
  assign n3808 = ~n3676 & ~n3679;
  assign n3809 = ~n3656 & ~n3662;
  assign n3810 = ~n3610 & n3632;
  assign n3811 = ~n3636 & ~n3810;
  assign n3812 = n286 & n3622;
  assign n3813 = n3407 & n3614;
  assign n3814 = ~n3619 & n3813;
  assign n3815 = pi64  & n3814;
  assign n3816 = pi66  & n3620;
  assign n3817 = pi65  & n3615;
  assign n3818 = ~n3816 & ~n3817;
  assign n3819 = ~n3812 & n3818;
  assign n3820 = ~n3815 & n3819;
  assign n3821 = pi32  & ~n3820;
  assign n3822 = pi32  & ~n3821;
  assign n3823 = ~n3820 & ~n3821;
  assign n3824 = ~n3822 & ~n3823;
  assign n3825 = ~n3630 & n3824;
  assign n3826 = n3630 & ~n3824;
  assign n3827 = ~n3825 & ~n3826;
  assign n3828 = n401 & n3034;
  assign n3829 = pi67  & n3225;
  assign n3830 = pi69  & n3032;
  assign n3831 = pi68  & n3027;
  assign n3832 = ~n3830 & ~n3831;
  assign n3833 = ~n3829 & n3832;
  assign n3834 = ~n3828 & n3833;
  assign n3835 = pi29  & ~n3834;
  assign n3836 = pi29  & ~n3835;
  assign n3837 = ~n3834 & ~n3835;
  assign n3838 = ~n3836 & ~n3837;
  assign n3839 = n3827 & ~n3838;
  assign n3840 = ~n3827 & n3838;
  assign n3841 = ~n3839 & ~n3840;
  assign n3842 = ~n3811 & n3841;
  assign n3843 = ~n3811 & ~n3842;
  assign n3844 = ~n3839 & ~n3842;
  assign n3845 = ~n3840 & n3844;
  assign n3846 = ~n3843 & ~n3845;
  assign n3847 = n576 & n2523;
  assign n3848 = pi70  & n2667;
  assign n3849 = pi72  & n2521;
  assign n3850 = pi71  & n2516;
  assign n3851 = ~n3849 & ~n3850;
  assign n3852 = ~n3848 & n3851;
  assign n3853 = ~n3847 & n3852;
  assign n3854 = pi26  & ~n3853;
  assign n3855 = pi26  & ~n3854;
  assign n3856 = ~n3853 & ~n3854;
  assign n3857 = ~n3855 & ~n3856;
  assign n3858 = ~n3846 & ~n3857;
  assign n3859 = ~n3846 & ~n3858;
  assign n3860 = ~n3857 & ~n3858;
  assign n3861 = ~n3859 & ~n3860;
  assign n3862 = ~n3639 & ~n3642;
  assign n3863 = n3861 & n3862;
  assign n3864 = ~n3861 & ~n3862;
  assign n3865 = ~n3863 & ~n3864;
  assign n3866 = n809 & n2043;
  assign n3867 = pi73  & n2180;
  assign n3868 = pi75  & n2041;
  assign n3869 = pi74  & n2036;
  assign n3870 = ~n3868 & ~n3869;
  assign n3871 = ~n3867 & n3870;
  assign n3872 = ~n3866 & n3871;
  assign n3873 = pi23  & ~n3872;
  assign n3874 = pi23  & ~n3873;
  assign n3875 = ~n3872 & ~n3873;
  assign n3876 = ~n3874 & ~n3875;
  assign n3877 = n3865 & ~n3876;
  assign n3878 = ~n3865 & n3876;
  assign n3879 = ~n3877 & ~n3878;
  assign n3880 = ~n3809 & n3879;
  assign n3881 = ~n3809 & ~n3880;
  assign n3882 = ~n3877 & ~n3880;
  assign n3883 = ~n3878 & n3882;
  assign n3884 = ~n3881 & ~n3883;
  assign n3885 = n1025 & n1611;
  assign n3886 = pi76  & n1745;
  assign n3887 = pi78  & n1609;
  assign n3888 = pi77  & n1604;
  assign n3889 = ~n3887 & ~n3888;
  assign n3890 = ~n3886 & n3889;
  assign n3891 = ~n3885 & n3890;
  assign n3892 = pi20  & ~n3891;
  assign n3893 = pi20  & ~n3892;
  assign n3894 = ~n3891 & ~n3892;
  assign n3895 = ~n3893 & ~n3894;
  assign n3896 = n3884 & n3895;
  assign n3897 = ~n3884 & ~n3895;
  assign n3898 = ~n3896 & ~n3897;
  assign n3899 = ~n3808 & n3898;
  assign n3900 = n3808 & ~n3898;
  assign n3901 = ~n3899 & ~n3900;
  assign n3902 = n1297 & n1434;
  assign n3903 = pi79  & n1366;
  assign n3904 = pi81  & n1295;
  assign n3905 = pi80  & n1290;
  assign n3906 = ~n3904 & ~n3905;
  assign n3907 = ~n3903 & n3906;
  assign n3908 = ~n3902 & n3907;
  assign n3909 = pi17  & ~n3908;
  assign n3910 = pi17  & ~n3909;
  assign n3911 = ~n3908 & ~n3909;
  assign n3912 = ~n3910 & ~n3911;
  assign n3913 = n3901 & ~n3912;
  assign n3914 = n3901 & ~n3913;
  assign n3915 = ~n3912 & ~n3913;
  assign n3916 = ~n3914 & ~n3915;
  assign n3917 = ~n3693 & ~n3699;
  assign n3918 = n3916 & n3917;
  assign n3919 = ~n3916 & ~n3917;
  assign n3920 = ~n3918 & ~n3919;
  assign n3921 = n938 & n1834;
  assign n3922 = pi82  & n1052;
  assign n3923 = pi84  & n936;
  assign n3924 = pi83  & n931;
  assign n3925 = ~n3923 & ~n3924;
  assign n3926 = ~n3922 & n3925;
  assign n3927 = ~n3921 & n3926;
  assign n3928 = pi14  & ~n3927;
  assign n3929 = pi14  & ~n3928;
  assign n3930 = ~n3927 & ~n3928;
  assign n3931 = ~n3929 & ~n3930;
  assign n3932 = n3920 & ~n3931;
  assign n3933 = ~n3920 & n3931;
  assign n3934 = ~n3932 & ~n3933;
  assign n3935 = ~n3807 & n3934;
  assign n3936 = ~n3807 & ~n3935;
  assign n3937 = ~n3932 & ~n3935;
  assign n3938 = ~n3933 & n3937;
  assign n3939 = ~n3936 & ~n3938;
  assign n3940 = n687 & n2288;
  assign n3941 = pi85  & n763;
  assign n3942 = pi87  & n685;
  assign n3943 = pi86  & n680;
  assign n3944 = ~n3942 & ~n3943;
  assign n3945 = ~n3941 & n3944;
  assign n3946 = ~n3940 & n3945;
  assign n3947 = pi11  & ~n3946;
  assign n3948 = pi11  & ~n3947;
  assign n3949 = ~n3946 & ~n3947;
  assign n3950 = ~n3948 & ~n3949;
  assign n3951 = n3939 & n3950;
  assign n3952 = ~n3939 & ~n3950;
  assign n3953 = ~n3951 & ~n3952;
  assign n3954 = ~n3806 & n3953;
  assign n3955 = n3806 & ~n3953;
  assign n3956 = ~n3954 & ~n3955;
  assign n3957 = n498 & n2801;
  assign n3958 = pi88  & n537;
  assign n3959 = pi90  & n496;
  assign n3960 = pi89  & n491;
  assign n3961 = ~n3959 & ~n3960;
  assign n3962 = ~n3958 & n3961;
  assign n3963 = ~n3957 & n3962;
  assign n3964 = pi8  & ~n3963;
  assign n3965 = pi8  & ~n3964;
  assign n3966 = ~n3963 & ~n3964;
  assign n3967 = ~n3965 & ~n3966;
  assign n3968 = n3956 & ~n3967;
  assign n3969 = n3956 & ~n3968;
  assign n3970 = ~n3967 & ~n3968;
  assign n3971 = ~n3969 & ~n3970;
  assign n3972 = ~n3751 & ~n3757;
  assign n3973 = n3971 & n3972;
  assign n3974 = ~n3971 & ~n3972;
  assign n3975 = ~n3973 & ~n3974;
  assign n3976 = n342 & n3371;
  assign n3977 = pi91  & n380;
  assign n3978 = pi93  & n340;
  assign n3979 = pi92  & n335;
  assign n3980 = ~n3978 & ~n3979;
  assign n3981 = ~n3977 & n3980;
  assign n3982 = ~n3976 & n3981;
  assign n3983 = pi5  & ~n3982;
  assign n3984 = pi5  & ~n3983;
  assign n3985 = ~n3982 & ~n3983;
  assign n3986 = ~n3984 & ~n3985;
  assign n3987 = n3975 & ~n3986;
  assign n3988 = ~n3975 & n3986;
  assign n3989 = ~n3987 & ~n3988;
  assign n3990 = ~n3805 & n3989;
  assign n3991 = ~n3805 & ~n3990;
  assign n3992 = ~n3987 & ~n3990;
  assign n3993 = ~n3988 & n3992;
  assign n3994 = ~n3991 & ~n3993;
  assign n3995 = ~n3780 & ~n3782;
  assign n3996 = ~pi95  & ~pi96 ;
  assign n3997 = pi95  & pi96 ;
  assign n3998 = ~n3996 & ~n3997;
  assign n3999 = ~n3995 & n3998;
  assign n4000 = n3995 & ~n3998;
  assign n4001 = ~n3999 & ~n4000;
  assign n4002 = n262 & n4001;
  assign n4003 = pi94  & n288;
  assign n4004 = pi96  & n267;
  assign n4005 = pi95  & n269;
  assign n4006 = ~n4004 & ~n4005;
  assign n4007 = ~n4003 & n4006;
  assign n4008 = ~n4002 & n4007;
  assign n4009 = pi2  & ~n4008;
  assign n4010 = pi2  & ~n4009;
  assign n4011 = ~n4008 & ~n4009;
  assign n4012 = ~n4010 & ~n4011;
  assign n4013 = ~n3994 & n4012;
  assign n4014 = n3994 & ~n4012;
  assign n4015 = ~n4013 & ~n4014;
  assign n4016 = ~n3804 & ~n4015;
  assign n4017 = n3804 & n4015;
  assign po32  = ~n4016 & ~n4017;
  assign n4019 = ~n3994 & ~n4012;
  assign n4020 = ~n4016 & ~n4019;
  assign n4021 = ~n3952 & ~n3954;
  assign n4022 = ~n3913 & ~n3919;
  assign n4023 = ~n3897 & ~n3899;
  assign n4024 = ~n3858 & ~n3864;
  assign n4025 = pi32  & ~pi33 ;
  assign n4026 = ~pi32  & pi33 ;
  assign n4027 = ~n4025 & ~n4026;
  assign n4028 = pi64  & ~n4027;
  assign n4029 = ~n3826 & n4028;
  assign n4030 = n3826 & ~n4028;
  assign n4031 = ~n4029 & ~n4030;
  assign n4032 = n309 & n3622;
  assign n4033 = pi65  & n3814;
  assign n4034 = pi67  & n3620;
  assign n4035 = pi66  & n3615;
  assign n4036 = ~n4034 & ~n4035;
  assign n4037 = ~n4033 & n4036;
  assign n4038 = ~n4032 & n4037;
  assign n4039 = pi32  & ~n4038;
  assign n4040 = pi32  & ~n4039;
  assign n4041 = ~n4038 & ~n4039;
  assign n4042 = ~n4040 & ~n4041;
  assign n4043 = ~n4031 & ~n4042;
  assign n4044 = n4031 & n4042;
  assign n4045 = ~n4043 & ~n4044;
  assign n4046 = n450 & n3034;
  assign n4047 = pi68  & n3225;
  assign n4048 = pi70  & n3032;
  assign n4049 = pi69  & n3027;
  assign n4050 = ~n4048 & ~n4049;
  assign n4051 = ~n4047 & n4050;
  assign n4052 = ~n4046 & n4051;
  assign n4053 = pi29  & ~n4052;
  assign n4054 = pi29  & ~n4053;
  assign n4055 = ~n4052 & ~n4053;
  assign n4056 = ~n4054 & ~n4055;
  assign n4057 = n4045 & ~n4056;
  assign n4058 = n4045 & ~n4057;
  assign n4059 = ~n4056 & ~n4057;
  assign n4060 = ~n4058 & ~n4059;
  assign n4061 = ~n3844 & n4060;
  assign n4062 = n3844 & ~n4060;
  assign n4063 = ~n4061 & ~n4062;
  assign n4064 = n642 & n2523;
  assign n4065 = pi71  & n2667;
  assign n4066 = pi73  & n2521;
  assign n4067 = pi72  & n2516;
  assign n4068 = ~n4066 & ~n4067;
  assign n4069 = ~n4065 & n4068;
  assign n4070 = ~n4064 & n4069;
  assign n4071 = pi26  & ~n4070;
  assign n4072 = pi26  & ~n4071;
  assign n4073 = ~n4070 & ~n4071;
  assign n4074 = ~n4072 & ~n4073;
  assign n4075 = ~n4063 & ~n4074;
  assign n4076 = n4063 & n4074;
  assign n4077 = ~n4075 & ~n4076;
  assign n4078 = n4024 & ~n4077;
  assign n4079 = ~n4024 & n4077;
  assign n4080 = ~n4078 & ~n4079;
  assign n4081 = n891 & n2043;
  assign n4082 = pi74  & n2180;
  assign n4083 = pi76  & n2041;
  assign n4084 = pi75  & n2036;
  assign n4085 = ~n4083 & ~n4084;
  assign n4086 = ~n4082 & n4085;
  assign n4087 = ~n4081 & n4086;
  assign n4088 = pi23  & ~n4087;
  assign n4089 = pi23  & ~n4088;
  assign n4090 = ~n4087 & ~n4088;
  assign n4091 = ~n4089 & ~n4090;
  assign n4092 = ~n4080 & n4091;
  assign n4093 = n4080 & ~n4091;
  assign n4094 = ~n4092 & ~n4093;
  assign n4095 = ~n3882 & n4094;
  assign n4096 = n3882 & ~n4094;
  assign n4097 = ~n4095 & ~n4096;
  assign n4098 = n1122 & n1611;
  assign n4099 = pi77  & n1745;
  assign n4100 = pi79  & n1609;
  assign n4101 = pi78  & n1604;
  assign n4102 = ~n4100 & ~n4101;
  assign n4103 = ~n4099 & n4102;
  assign n4104 = ~n4098 & n4103;
  assign n4105 = pi20  & ~n4104;
  assign n4106 = pi20  & ~n4105;
  assign n4107 = ~n4104 & ~n4105;
  assign n4108 = ~n4106 & ~n4107;
  assign n4109 = n4097 & ~n4108;
  assign n4110 = n4097 & ~n4109;
  assign n4111 = ~n4108 & ~n4109;
  assign n4112 = ~n4110 & ~n4111;
  assign n4113 = ~n4023 & n4112;
  assign n4114 = n4023 & ~n4112;
  assign n4115 = ~n4113 & ~n4114;
  assign n4116 = n1297 & n1554;
  assign n4117 = pi80  & n1366;
  assign n4118 = pi82  & n1295;
  assign n4119 = pi81  & n1290;
  assign n4120 = ~n4118 & ~n4119;
  assign n4121 = ~n4117 & n4120;
  assign n4122 = ~n4116 & n4121;
  assign n4123 = pi17  & ~n4122;
  assign n4124 = pi17  & ~n4123;
  assign n4125 = ~n4122 & ~n4123;
  assign n4126 = ~n4124 & ~n4125;
  assign n4127 = ~n4115 & ~n4126;
  assign n4128 = n4115 & n4126;
  assign n4129 = ~n4127 & ~n4128;
  assign n4130 = n4022 & ~n4129;
  assign n4131 = ~n4022 & n4129;
  assign n4132 = ~n4130 & ~n4131;
  assign n4133 = n938 & n1972;
  assign n4134 = pi83  & n1052;
  assign n4135 = pi85  & n936;
  assign n4136 = pi84  & n931;
  assign n4137 = ~n4135 & ~n4136;
  assign n4138 = ~n4134 & n4137;
  assign n4139 = ~n4133 & n4138;
  assign n4140 = pi14  & ~n4139;
  assign n4141 = pi14  & ~n4140;
  assign n4142 = ~n4139 & ~n4140;
  assign n4143 = ~n4141 & ~n4142;
  assign n4144 = n4132 & ~n4143;
  assign n4145 = n4132 & ~n4144;
  assign n4146 = ~n4143 & ~n4144;
  assign n4147 = ~n4145 & ~n4146;
  assign n4148 = ~n3937 & n4147;
  assign n4149 = n3937 & ~n4147;
  assign n4150 = ~n4148 & ~n4149;
  assign n4151 = n687 & n2446;
  assign n4152 = pi86  & n763;
  assign n4153 = pi88  & n685;
  assign n4154 = pi87  & n680;
  assign n4155 = ~n4153 & ~n4154;
  assign n4156 = ~n4152 & n4155;
  assign n4157 = ~n4151 & n4156;
  assign n4158 = pi11  & ~n4157;
  assign n4159 = pi11  & ~n4158;
  assign n4160 = ~n4157 & ~n4158;
  assign n4161 = ~n4159 & ~n4160;
  assign n4162 = n4150 & n4161;
  assign n4163 = ~n4150 & ~n4161;
  assign n4164 = ~n4162 & ~n4163;
  assign n4165 = ~n4021 & n4164;
  assign n4166 = n4021 & ~n4164;
  assign n4167 = ~n4165 & ~n4166;
  assign n4168 = n498 & n2978;
  assign n4169 = pi89  & n537;
  assign n4170 = pi91  & n496;
  assign n4171 = pi90  & n491;
  assign n4172 = ~n4170 & ~n4171;
  assign n4173 = ~n4169 & n4172;
  assign n4174 = ~n4168 & n4173;
  assign n4175 = pi8  & ~n4174;
  assign n4176 = pi8  & ~n4175;
  assign n4177 = ~n4174 & ~n4175;
  assign n4178 = ~n4176 & ~n4177;
  assign n4179 = n4167 & ~n4178;
  assign n4180 = n4167 & ~n4179;
  assign n4181 = ~n4178 & ~n4179;
  assign n4182 = ~n4180 & ~n4181;
  assign n4183 = ~n3968 & ~n3974;
  assign n4184 = n4182 & n4183;
  assign n4185 = ~n4182 & ~n4183;
  assign n4186 = ~n4184 & ~n4185;
  assign n4187 = n342 & n3565;
  assign n4188 = pi92  & n380;
  assign n4189 = pi94  & n340;
  assign n4190 = pi93  & n335;
  assign n4191 = ~n4189 & ~n4190;
  assign n4192 = ~n4188 & n4191;
  assign n4193 = ~n4187 & n4192;
  assign n4194 = pi5  & ~n4193;
  assign n4195 = pi5  & ~n4194;
  assign n4196 = ~n4193 & ~n4194;
  assign n4197 = ~n4195 & ~n4196;
  assign n4198 = n4186 & ~n4197;
  assign n4199 = n4186 & ~n4198;
  assign n4200 = ~n4197 & ~n4198;
  assign n4201 = ~n4199 & ~n4200;
  assign n4202 = ~n3992 & n4201;
  assign n4203 = n3992 & ~n4201;
  assign n4204 = ~n4202 & ~n4203;
  assign n4205 = ~n3997 & ~n3999;
  assign n4206 = ~pi96  & ~pi97 ;
  assign n4207 = pi96  & pi97 ;
  assign n4208 = ~n4206 & ~n4207;
  assign n4209 = ~n4205 & n4208;
  assign n4210 = n4205 & ~n4208;
  assign n4211 = ~n4209 & ~n4210;
  assign n4212 = n262 & n4211;
  assign n4213 = pi95  & n288;
  assign n4214 = pi97  & n267;
  assign n4215 = pi96  & n269;
  assign n4216 = ~n4214 & ~n4215;
  assign n4217 = ~n4213 & n4216;
  assign n4218 = ~n4212 & n4217;
  assign n4219 = pi2  & ~n4218;
  assign n4220 = pi2  & ~n4219;
  assign n4221 = ~n4218 & ~n4219;
  assign n4222 = ~n4220 & ~n4221;
  assign n4223 = ~n4204 & ~n4222;
  assign n4224 = n4204 & n4222;
  assign n4225 = ~n4223 & ~n4224;
  assign n4226 = ~n4020 & n4225;
  assign n4227 = n4020 & ~n4225;
  assign po33  = ~n4226 & ~n4227;
  assign n4229 = ~n4223 & ~n4226;
  assign n4230 = ~n3992 & ~n4201;
  assign n4231 = ~n4198 & ~n4230;
  assign n4232 = ~n4163 & ~n4165;
  assign n4233 = ~n4093 & ~n4095;
  assign n4234 = ~n3844 & ~n4060;
  assign n4235 = ~n4057 & ~n4234;
  assign n4236 = n475 & n3034;
  assign n4237 = pi69  & n3225;
  assign n4238 = pi71  & n3032;
  assign n4239 = pi70  & n3027;
  assign n4240 = ~n4238 & ~n4239;
  assign n4241 = ~n4237 & n4240;
  assign n4242 = ~n4236 & n4241;
  assign n4243 = pi29  & ~n4242;
  assign n4244 = pi29  & ~n4243;
  assign n4245 = ~n4242 & ~n4243;
  assign n4246 = ~n4244 & ~n4245;
  assign n4247 = n3826 & n4028;
  assign n4248 = ~n4043 & ~n4247;
  assign n4249 = n359 & n3622;
  assign n4250 = pi66  & n3814;
  assign n4251 = pi68  & n3620;
  assign n4252 = pi67  & n3615;
  assign n4253 = ~n4251 & ~n4252;
  assign n4254 = ~n4250 & n4253;
  assign n4255 = ~n4249 & n4254;
  assign n4256 = pi32  & ~n4255;
  assign n4257 = pi32  & ~n4256;
  assign n4258 = ~n4255 & ~n4256;
  assign n4259 = ~n4257 & ~n4258;
  assign n4260 = pi35  & ~n4028;
  assign n4261 = ~pi33  & pi34 ;
  assign n4262 = pi33  & ~pi34 ;
  assign n4263 = ~n4261 & ~n4262;
  assign n4264 = n4027 & ~n4263;
  assign n4265 = pi64  & n4264;
  assign n4266 = ~pi34  & pi35 ;
  assign n4267 = pi34  & ~pi35 ;
  assign n4268 = ~n4266 & ~n4267;
  assign n4269 = ~n4027 & n4268;
  assign n4270 = pi65  & n4269;
  assign n4271 = ~n4027 & ~n4268;
  assign n4272 = ~n265 & n4271;
  assign n4273 = ~n4265 & ~n4270;
  assign n4274 = ~n4272 & n4273;
  assign n4275 = pi35  & ~n4274;
  assign n4276 = pi35  & ~n4275;
  assign n4277 = ~n4274 & ~n4275;
  assign n4278 = ~n4276 & ~n4277;
  assign n4279 = n4260 & ~n4278;
  assign n4280 = ~n4260 & n4278;
  assign n4281 = ~n4279 & ~n4280;
  assign n4282 = n4259 & ~n4281;
  assign n4283 = ~n4259 & n4281;
  assign n4284 = ~n4282 & ~n4283;
  assign n4285 = ~n4248 & n4284;
  assign n4286 = n4248 & ~n4284;
  assign n4287 = ~n4285 & ~n4286;
  assign n4288 = n4246 & ~n4287;
  assign n4289 = ~n4246 & n4287;
  assign n4290 = ~n4288 & ~n4289;
  assign n4291 = ~n4235 & n4290;
  assign n4292 = n4235 & ~n4290;
  assign n4293 = ~n4291 & ~n4292;
  assign n4294 = n729 & n2523;
  assign n4295 = pi72  & n2667;
  assign n4296 = pi74  & n2521;
  assign n4297 = pi73  & n2516;
  assign n4298 = ~n4296 & ~n4297;
  assign n4299 = ~n4295 & n4298;
  assign n4300 = ~n4294 & n4299;
  assign n4301 = pi26  & ~n4300;
  assign n4302 = pi26  & ~n4301;
  assign n4303 = ~n4300 & ~n4301;
  assign n4304 = ~n4302 & ~n4303;
  assign n4305 = n4293 & ~n4304;
  assign n4306 = n4293 & ~n4305;
  assign n4307 = ~n4304 & ~n4305;
  assign n4308 = ~n4306 & ~n4307;
  assign n4309 = ~n4075 & ~n4079;
  assign n4310 = n4308 & n4309;
  assign n4311 = ~n4308 & ~n4309;
  assign n4312 = ~n4310 & ~n4311;
  assign n4313 = n999 & n2043;
  assign n4314 = pi75  & n2180;
  assign n4315 = pi77  & n2041;
  assign n4316 = pi76  & n2036;
  assign n4317 = ~n4315 & ~n4316;
  assign n4318 = ~n4314 & n4317;
  assign n4319 = ~n4313 & n4318;
  assign n4320 = pi23  & ~n4319;
  assign n4321 = pi23  & ~n4320;
  assign n4322 = ~n4319 & ~n4320;
  assign n4323 = ~n4321 & ~n4322;
  assign n4324 = n4312 & ~n4323;
  assign n4325 = ~n4312 & n4323;
  assign n4326 = ~n4324 & ~n4325;
  assign n4327 = ~n4233 & n4326;
  assign n4328 = ~n4233 & ~n4327;
  assign n4329 = ~n4324 & ~n4327;
  assign n4330 = ~n4325 & n4329;
  assign n4331 = ~n4328 & ~n4330;
  assign n4332 = n1225 & n1611;
  assign n4333 = pi78  & n1745;
  assign n4334 = pi80  & n1609;
  assign n4335 = pi79  & n1604;
  assign n4336 = ~n4334 & ~n4335;
  assign n4337 = ~n4333 & n4336;
  assign n4338 = ~n4332 & n4337;
  assign n4339 = pi20  & ~n4338;
  assign n4340 = pi20  & ~n4339;
  assign n4341 = ~n4338 & ~n4339;
  assign n4342 = ~n4340 & ~n4341;
  assign n4343 = ~n4331 & ~n4342;
  assign n4344 = ~n4331 & ~n4343;
  assign n4345 = ~n4342 & ~n4343;
  assign n4346 = ~n4344 & ~n4345;
  assign n4347 = ~n4023 & ~n4112;
  assign n4348 = ~n4109 & ~n4347;
  assign n4349 = n4346 & n4348;
  assign n4350 = ~n4346 & ~n4348;
  assign n4351 = ~n4349 & ~n4350;
  assign n4352 = n1297 & n1696;
  assign n4353 = pi81  & n1366;
  assign n4354 = pi83  & n1295;
  assign n4355 = pi82  & n1290;
  assign n4356 = ~n4354 & ~n4355;
  assign n4357 = ~n4353 & n4356;
  assign n4358 = ~n4352 & n4357;
  assign n4359 = pi17  & ~n4358;
  assign n4360 = pi17  & ~n4359;
  assign n4361 = ~n4358 & ~n4359;
  assign n4362 = ~n4360 & ~n4361;
  assign n4363 = n4351 & ~n4362;
  assign n4364 = n4351 & ~n4363;
  assign n4365 = ~n4362 & ~n4363;
  assign n4366 = ~n4364 & ~n4365;
  assign n4367 = ~n4127 & ~n4131;
  assign n4368 = n4366 & n4367;
  assign n4369 = ~n4366 & ~n4367;
  assign n4370 = ~n4368 & ~n4369;
  assign n4371 = n938 & n2133;
  assign n4372 = pi84  & n1052;
  assign n4373 = pi86  & n936;
  assign n4374 = pi85  & n931;
  assign n4375 = ~n4373 & ~n4374;
  assign n4376 = ~n4372 & n4375;
  assign n4377 = ~n4371 & n4376;
  assign n4378 = pi14  & ~n4377;
  assign n4379 = pi14  & ~n4378;
  assign n4380 = ~n4377 & ~n4378;
  assign n4381 = ~n4379 & ~n4380;
  assign n4382 = n4370 & ~n4381;
  assign n4383 = n4370 & ~n4382;
  assign n4384 = ~n4381 & ~n4382;
  assign n4385 = ~n4383 & ~n4384;
  assign n4386 = ~n3937 & ~n4147;
  assign n4387 = ~n4144 & ~n4386;
  assign n4388 = n4385 & n4387;
  assign n4389 = ~n4385 & ~n4387;
  assign n4390 = ~n4388 & ~n4389;
  assign n4391 = n687 & n2473;
  assign n4392 = pi87  & n763;
  assign n4393 = pi89  & n685;
  assign n4394 = pi88  & n680;
  assign n4395 = ~n4393 & ~n4394;
  assign n4396 = ~n4392 & n4395;
  assign n4397 = ~n4391 & n4396;
  assign n4398 = pi11  & ~n4397;
  assign n4399 = pi11  & ~n4398;
  assign n4400 = ~n4397 & ~n4398;
  assign n4401 = ~n4399 & ~n4400;
  assign n4402 = n4390 & ~n4401;
  assign n4403 = ~n4390 & n4401;
  assign n4404 = ~n4402 & ~n4403;
  assign n4405 = ~n4232 & n4404;
  assign n4406 = ~n4232 & ~n4405;
  assign n4407 = ~n4402 & ~n4405;
  assign n4408 = ~n4403 & n4407;
  assign n4409 = ~n4406 & ~n4408;
  assign n4410 = n498 & n3177;
  assign n4411 = pi90  & n537;
  assign n4412 = pi92  & n496;
  assign n4413 = pi91  & n491;
  assign n4414 = ~n4412 & ~n4413;
  assign n4415 = ~n4411 & n4414;
  assign n4416 = ~n4410 & n4415;
  assign n4417 = pi8  & ~n4416;
  assign n4418 = pi8  & ~n4417;
  assign n4419 = ~n4416 & ~n4417;
  assign n4420 = ~n4418 & ~n4419;
  assign n4421 = ~n4409 & ~n4420;
  assign n4422 = ~n4409 & ~n4421;
  assign n4423 = ~n4420 & ~n4421;
  assign n4424 = ~n4422 & ~n4423;
  assign n4425 = ~n4179 & ~n4185;
  assign n4426 = n4424 & n4425;
  assign n4427 = ~n4424 & ~n4425;
  assign n4428 = ~n4426 & ~n4427;
  assign n4429 = n342 & n3784;
  assign n4430 = pi93  & n380;
  assign n4431 = pi95  & n340;
  assign n4432 = pi94  & n335;
  assign n4433 = ~n4431 & ~n4432;
  assign n4434 = ~n4430 & n4433;
  assign n4435 = ~n4429 & n4434;
  assign n4436 = pi5  & ~n4435;
  assign n4437 = pi5  & ~n4436;
  assign n4438 = ~n4435 & ~n4436;
  assign n4439 = ~n4437 & ~n4438;
  assign n4440 = n4428 & ~n4439;
  assign n4441 = ~n4428 & n4439;
  assign n4442 = ~n4440 & ~n4441;
  assign n4443 = ~n4231 & n4442;
  assign n4444 = ~n4231 & ~n4443;
  assign n4445 = ~n4440 & ~n4443;
  assign n4446 = ~n4441 & n4445;
  assign n4447 = ~n4444 & ~n4446;
  assign n4448 = ~n4207 & ~n4209;
  assign n4449 = ~pi97  & ~pi98 ;
  assign n4450 = pi97  & pi98 ;
  assign n4451 = ~n4449 & ~n4450;
  assign n4452 = ~n4448 & n4451;
  assign n4453 = n4448 & ~n4451;
  assign n4454 = ~n4452 & ~n4453;
  assign n4455 = n262 & n4454;
  assign n4456 = pi96  & n288;
  assign n4457 = pi98  & n267;
  assign n4458 = pi97  & n269;
  assign n4459 = ~n4457 & ~n4458;
  assign n4460 = ~n4456 & n4459;
  assign n4461 = ~n4455 & n4460;
  assign n4462 = pi2  & ~n4461;
  assign n4463 = pi2  & ~n4462;
  assign n4464 = ~n4461 & ~n4462;
  assign n4465 = ~n4463 & ~n4464;
  assign n4466 = ~n4447 & n4465;
  assign n4467 = n4447 & ~n4465;
  assign n4468 = ~n4466 & ~n4467;
  assign n4469 = ~n4229 & ~n4468;
  assign n4470 = n4229 & n4468;
  assign po34  = ~n4469 & ~n4470;
  assign n4472 = ~n4447 & ~n4465;
  assign n4473 = ~n4469 & ~n4472;
  assign n4474 = n687 & n2801;
  assign n4475 = pi88  & n763;
  assign n4476 = pi90  & n685;
  assign n4477 = pi89  & n680;
  assign n4478 = ~n4476 & ~n4477;
  assign n4479 = ~n4475 & n4478;
  assign n4480 = ~n4474 & n4479;
  assign n4481 = pi11  & ~n4480;
  assign n4482 = pi11  & ~n4481;
  assign n4483 = ~n4480 & ~n4481;
  assign n4484 = ~n4482 & ~n4483;
  assign n4485 = ~n4382 & ~n4389;
  assign n4486 = ~n4363 & ~n4369;
  assign n4487 = ~n4305 & ~n4311;
  assign n4488 = n809 & n2523;
  assign n4489 = pi73  & n2667;
  assign n4490 = pi75  & n2521;
  assign n4491 = pi74  & n2516;
  assign n4492 = ~n4490 & ~n4491;
  assign n4493 = ~n4489 & n4492;
  assign n4494 = ~n4488 & n4493;
  assign n4495 = pi26  & ~n4494;
  assign n4496 = pi26  & ~n4495;
  assign n4497 = ~n4494 & ~n4495;
  assign n4498 = ~n4496 & ~n4497;
  assign n4499 = ~n4289 & ~n4291;
  assign n4500 = ~n4283 & ~n4285;
  assign n4501 = n286 & n4271;
  assign n4502 = n4027 & n4263;
  assign n4503 = ~n4268 & n4502;
  assign n4504 = pi64  & n4503;
  assign n4505 = pi66  & n4269;
  assign n4506 = pi65  & n4264;
  assign n4507 = ~n4505 & ~n4506;
  assign n4508 = ~n4501 & n4507;
  assign n4509 = ~n4504 & n4508;
  assign n4510 = pi35  & ~n4509;
  assign n4511 = pi35  & ~n4510;
  assign n4512 = ~n4509 & ~n4510;
  assign n4513 = ~n4511 & ~n4512;
  assign n4514 = ~n4279 & n4513;
  assign n4515 = n4279 & ~n4513;
  assign n4516 = ~n4514 & ~n4515;
  assign n4517 = n401 & n3622;
  assign n4518 = pi67  & n3814;
  assign n4519 = pi69  & n3620;
  assign n4520 = pi68  & n3615;
  assign n4521 = ~n4519 & ~n4520;
  assign n4522 = ~n4518 & n4521;
  assign n4523 = ~n4517 & n4522;
  assign n4524 = pi32  & ~n4523;
  assign n4525 = pi32  & ~n4524;
  assign n4526 = ~n4523 & ~n4524;
  assign n4527 = ~n4525 & ~n4526;
  assign n4528 = n4516 & ~n4527;
  assign n4529 = ~n4516 & n4527;
  assign n4530 = ~n4528 & ~n4529;
  assign n4531 = ~n4500 & n4530;
  assign n4532 = ~n4500 & ~n4531;
  assign n4533 = ~n4528 & ~n4531;
  assign n4534 = ~n4529 & n4533;
  assign n4535 = ~n4532 & ~n4534;
  assign n4536 = n576 & n3034;
  assign n4537 = pi70  & n3225;
  assign n4538 = pi72  & n3032;
  assign n4539 = pi71  & n3027;
  assign n4540 = ~n4538 & ~n4539;
  assign n4541 = ~n4537 & n4540;
  assign n4542 = ~n4536 & n4541;
  assign n4543 = pi29  & ~n4542;
  assign n4544 = pi29  & ~n4543;
  assign n4545 = ~n4542 & ~n4543;
  assign n4546 = ~n4544 & ~n4545;
  assign n4547 = ~n4535 & ~n4546;
  assign n4548 = ~n4535 & ~n4547;
  assign n4549 = ~n4546 & ~n4547;
  assign n4550 = ~n4548 & ~n4549;
  assign n4551 = ~n4499 & ~n4550;
  assign n4552 = n4499 & n4550;
  assign n4553 = ~n4551 & ~n4552;
  assign n4554 = ~n4498 & n4553;
  assign n4555 = ~n4498 & ~n4554;
  assign n4556 = n4553 & ~n4554;
  assign n4557 = ~n4555 & ~n4556;
  assign n4558 = ~n4487 & ~n4557;
  assign n4559 = ~n4487 & ~n4558;
  assign n4560 = ~n4557 & ~n4558;
  assign n4561 = ~n4559 & ~n4560;
  assign n4562 = n1025 & n2043;
  assign n4563 = pi76  & n2180;
  assign n4564 = pi78  & n2041;
  assign n4565 = pi77  & n2036;
  assign n4566 = ~n4564 & ~n4565;
  assign n4567 = ~n4563 & n4566;
  assign n4568 = ~n4562 & n4567;
  assign n4569 = pi23  & ~n4568;
  assign n4570 = pi23  & ~n4569;
  assign n4571 = ~n4568 & ~n4569;
  assign n4572 = ~n4570 & ~n4571;
  assign n4573 = n4561 & n4572;
  assign n4574 = ~n4561 & ~n4572;
  assign n4575 = ~n4573 & ~n4574;
  assign n4576 = ~n4329 & n4575;
  assign n4577 = n4329 & ~n4575;
  assign n4578 = ~n4576 & ~n4577;
  assign n4579 = n1434 & n1611;
  assign n4580 = pi79  & n1745;
  assign n4581 = pi81  & n1609;
  assign n4582 = pi80  & n1604;
  assign n4583 = ~n4581 & ~n4582;
  assign n4584 = ~n4580 & n4583;
  assign n4585 = ~n4579 & n4584;
  assign n4586 = pi20  & ~n4585;
  assign n4587 = pi20  & ~n4586;
  assign n4588 = ~n4585 & ~n4586;
  assign n4589 = ~n4587 & ~n4588;
  assign n4590 = n4578 & ~n4589;
  assign n4591 = n4578 & ~n4590;
  assign n4592 = ~n4589 & ~n4590;
  assign n4593 = ~n4591 & ~n4592;
  assign n4594 = ~n4343 & ~n4350;
  assign n4595 = n4593 & n4594;
  assign n4596 = ~n4593 & ~n4594;
  assign n4597 = ~n4595 & ~n4596;
  assign n4598 = n1297 & n1834;
  assign n4599 = pi82  & n1366;
  assign n4600 = pi84  & n1295;
  assign n4601 = pi83  & n1290;
  assign n4602 = ~n4600 & ~n4601;
  assign n4603 = ~n4599 & n4602;
  assign n4604 = ~n4598 & n4603;
  assign n4605 = pi17  & ~n4604;
  assign n4606 = pi17  & ~n4605;
  assign n4607 = ~n4604 & ~n4605;
  assign n4608 = ~n4606 & ~n4607;
  assign n4609 = n4597 & ~n4608;
  assign n4610 = ~n4597 & n4608;
  assign n4611 = ~n4609 & ~n4610;
  assign n4612 = ~n4486 & n4611;
  assign n4613 = ~n4486 & ~n4612;
  assign n4614 = ~n4609 & ~n4612;
  assign n4615 = ~n4610 & n4614;
  assign n4616 = ~n4613 & ~n4615;
  assign n4617 = n938 & n2288;
  assign n4618 = pi85  & n1052;
  assign n4619 = pi87  & n936;
  assign n4620 = pi86  & n931;
  assign n4621 = ~n4619 & ~n4620;
  assign n4622 = ~n4618 & n4621;
  assign n4623 = ~n4617 & n4622;
  assign n4624 = pi14  & ~n4623;
  assign n4625 = pi14  & ~n4624;
  assign n4626 = ~n4623 & ~n4624;
  assign n4627 = ~n4625 & ~n4626;
  assign n4628 = n4616 & n4627;
  assign n4629 = ~n4616 & ~n4627;
  assign n4630 = ~n4628 & ~n4629;
  assign n4631 = ~n4485 & n4630;
  assign n4632 = n4485 & ~n4630;
  assign n4633 = ~n4631 & ~n4632;
  assign n4634 = n4484 & ~n4633;
  assign n4635 = ~n4484 & n4633;
  assign n4636 = ~n4634 & ~n4635;
  assign n4637 = ~n4407 & n4636;
  assign n4638 = n4407 & ~n4636;
  assign n4639 = ~n4637 & ~n4638;
  assign n4640 = n498 & n3371;
  assign n4641 = pi91  & n537;
  assign n4642 = pi93  & n496;
  assign n4643 = pi92  & n491;
  assign n4644 = ~n4642 & ~n4643;
  assign n4645 = ~n4641 & n4644;
  assign n4646 = ~n4640 & n4645;
  assign n4647 = pi8  & ~n4646;
  assign n4648 = pi8  & ~n4647;
  assign n4649 = ~n4646 & ~n4647;
  assign n4650 = ~n4648 & ~n4649;
  assign n4651 = n4639 & ~n4650;
  assign n4652 = n4639 & ~n4651;
  assign n4653 = ~n4650 & ~n4651;
  assign n4654 = ~n4652 & ~n4653;
  assign n4655 = ~n4421 & ~n4427;
  assign n4656 = n4654 & n4655;
  assign n4657 = ~n4654 & ~n4655;
  assign n4658 = ~n4656 & ~n4657;
  assign n4659 = n342 & n4001;
  assign n4660 = pi94  & n380;
  assign n4661 = pi96  & n340;
  assign n4662 = pi95  & n335;
  assign n4663 = ~n4661 & ~n4662;
  assign n4664 = ~n4660 & n4663;
  assign n4665 = ~n4659 & n4664;
  assign n4666 = pi5  & ~n4665;
  assign n4667 = pi5  & ~n4666;
  assign n4668 = ~n4665 & ~n4666;
  assign n4669 = ~n4667 & ~n4668;
  assign n4670 = n4658 & ~n4669;
  assign n4671 = ~n4658 & n4669;
  assign n4672 = ~n4670 & ~n4671;
  assign n4673 = ~n4445 & n4672;
  assign n4674 = ~n4445 & ~n4673;
  assign n4675 = ~n4670 & ~n4673;
  assign n4676 = ~n4671 & n4675;
  assign n4677 = ~n4674 & ~n4676;
  assign n4678 = ~n4450 & ~n4452;
  assign n4679 = ~pi98  & ~pi99 ;
  assign n4680 = pi98  & pi99 ;
  assign n4681 = ~n4679 & ~n4680;
  assign n4682 = ~n4678 & n4681;
  assign n4683 = n4678 & ~n4681;
  assign n4684 = ~n4682 & ~n4683;
  assign n4685 = n262 & n4684;
  assign n4686 = pi97  & n288;
  assign n4687 = pi99  & n267;
  assign n4688 = pi98  & n269;
  assign n4689 = ~n4687 & ~n4688;
  assign n4690 = ~n4686 & n4689;
  assign n4691 = ~n4685 & n4690;
  assign n4692 = pi2  & ~n4691;
  assign n4693 = pi2  & ~n4692;
  assign n4694 = ~n4691 & ~n4692;
  assign n4695 = ~n4693 & ~n4694;
  assign n4696 = ~n4677 & n4695;
  assign n4697 = n4677 & ~n4695;
  assign n4698 = ~n4696 & ~n4697;
  assign n4699 = ~n4473 & ~n4698;
  assign n4700 = n4473 & n4698;
  assign po35  = ~n4699 & ~n4700;
  assign n4702 = n342 & n4211;
  assign n4703 = pi95  & n380;
  assign n4704 = pi97  & n340;
  assign n4705 = pi96  & n335;
  assign n4706 = ~n4704 & ~n4705;
  assign n4707 = ~n4703 & n4706;
  assign n4708 = ~n4702 & n4707;
  assign n4709 = pi5  & ~n4708;
  assign n4710 = pi5  & ~n4709;
  assign n4711 = ~n4708 & ~n4709;
  assign n4712 = ~n4710 & ~n4711;
  assign n4713 = ~n4651 & ~n4657;
  assign n4714 = ~n4635 & ~n4637;
  assign n4715 = ~n4629 & ~n4631;
  assign n4716 = ~n4590 & ~n4596;
  assign n4717 = ~n4574 & ~n4576;
  assign n4718 = ~n4547 & ~n4551;
  assign n4719 = pi35  & ~pi36 ;
  assign n4720 = ~pi35  & pi36 ;
  assign n4721 = ~n4719 & ~n4720;
  assign n4722 = pi64  & ~n4721;
  assign n4723 = ~n4515 & n4722;
  assign n4724 = n4515 & ~n4722;
  assign n4725 = ~n4723 & ~n4724;
  assign n4726 = n309 & n4271;
  assign n4727 = pi65  & n4503;
  assign n4728 = pi67  & n4269;
  assign n4729 = pi66  & n4264;
  assign n4730 = ~n4728 & ~n4729;
  assign n4731 = ~n4727 & n4730;
  assign n4732 = ~n4726 & n4731;
  assign n4733 = pi35  & ~n4732;
  assign n4734 = pi35  & ~n4733;
  assign n4735 = ~n4732 & ~n4733;
  assign n4736 = ~n4734 & ~n4735;
  assign n4737 = ~n4725 & ~n4736;
  assign n4738 = n4725 & n4736;
  assign n4739 = ~n4737 & ~n4738;
  assign n4740 = n450 & n3622;
  assign n4741 = pi68  & n3814;
  assign n4742 = pi70  & n3620;
  assign n4743 = pi69  & n3615;
  assign n4744 = ~n4742 & ~n4743;
  assign n4745 = ~n4741 & n4744;
  assign n4746 = ~n4740 & n4745;
  assign n4747 = pi32  & ~n4746;
  assign n4748 = pi32  & ~n4747;
  assign n4749 = ~n4746 & ~n4747;
  assign n4750 = ~n4748 & ~n4749;
  assign n4751 = n4739 & ~n4750;
  assign n4752 = n4739 & ~n4751;
  assign n4753 = ~n4750 & ~n4751;
  assign n4754 = ~n4752 & ~n4753;
  assign n4755 = ~n4533 & n4754;
  assign n4756 = n4533 & ~n4754;
  assign n4757 = ~n4755 & ~n4756;
  assign n4758 = n642 & n3034;
  assign n4759 = pi71  & n3225;
  assign n4760 = pi73  & n3032;
  assign n4761 = pi72  & n3027;
  assign n4762 = ~n4760 & ~n4761;
  assign n4763 = ~n4759 & n4762;
  assign n4764 = ~n4758 & n4763;
  assign n4765 = pi29  & ~n4764;
  assign n4766 = pi29  & ~n4765;
  assign n4767 = ~n4764 & ~n4765;
  assign n4768 = ~n4766 & ~n4767;
  assign n4769 = ~n4757 & ~n4768;
  assign n4770 = n4757 & n4768;
  assign n4771 = ~n4769 & ~n4770;
  assign n4772 = n4718 & ~n4771;
  assign n4773 = ~n4718 & n4771;
  assign n4774 = ~n4772 & ~n4773;
  assign n4775 = n891 & n2523;
  assign n4776 = pi74  & n2667;
  assign n4777 = pi76  & n2521;
  assign n4778 = pi75  & n2516;
  assign n4779 = ~n4777 & ~n4778;
  assign n4780 = ~n4776 & n4779;
  assign n4781 = ~n4775 & n4780;
  assign n4782 = pi26  & ~n4781;
  assign n4783 = pi26  & ~n4782;
  assign n4784 = ~n4781 & ~n4782;
  assign n4785 = ~n4783 & ~n4784;
  assign n4786 = ~n4774 & n4785;
  assign n4787 = n4774 & ~n4785;
  assign n4788 = ~n4786 & ~n4787;
  assign n4789 = ~n4554 & ~n4558;
  assign n4790 = n4788 & ~n4789;
  assign n4791 = ~n4788 & n4789;
  assign n4792 = ~n4790 & ~n4791;
  assign n4793 = n1122 & n2043;
  assign n4794 = pi77  & n2180;
  assign n4795 = pi79  & n2041;
  assign n4796 = pi78  & n2036;
  assign n4797 = ~n4795 & ~n4796;
  assign n4798 = ~n4794 & n4797;
  assign n4799 = ~n4793 & n4798;
  assign n4800 = pi23  & ~n4799;
  assign n4801 = pi23  & ~n4800;
  assign n4802 = ~n4799 & ~n4800;
  assign n4803 = ~n4801 & ~n4802;
  assign n4804 = n4792 & ~n4803;
  assign n4805 = n4792 & ~n4804;
  assign n4806 = ~n4803 & ~n4804;
  assign n4807 = ~n4805 & ~n4806;
  assign n4808 = ~n4717 & n4807;
  assign n4809 = n4717 & ~n4807;
  assign n4810 = ~n4808 & ~n4809;
  assign n4811 = n1554 & n1611;
  assign n4812 = pi80  & n1745;
  assign n4813 = pi82  & n1609;
  assign n4814 = pi81  & n1604;
  assign n4815 = ~n4813 & ~n4814;
  assign n4816 = ~n4812 & n4815;
  assign n4817 = ~n4811 & n4816;
  assign n4818 = pi20  & ~n4817;
  assign n4819 = pi20  & ~n4818;
  assign n4820 = ~n4817 & ~n4818;
  assign n4821 = ~n4819 & ~n4820;
  assign n4822 = ~n4810 & ~n4821;
  assign n4823 = n4810 & n4821;
  assign n4824 = ~n4822 & ~n4823;
  assign n4825 = n4716 & ~n4824;
  assign n4826 = ~n4716 & n4824;
  assign n4827 = ~n4825 & ~n4826;
  assign n4828 = n1297 & n1972;
  assign n4829 = pi83  & n1366;
  assign n4830 = pi85  & n1295;
  assign n4831 = pi84  & n1290;
  assign n4832 = ~n4830 & ~n4831;
  assign n4833 = ~n4829 & n4832;
  assign n4834 = ~n4828 & n4833;
  assign n4835 = pi17  & ~n4834;
  assign n4836 = pi17  & ~n4835;
  assign n4837 = ~n4834 & ~n4835;
  assign n4838 = ~n4836 & ~n4837;
  assign n4839 = n4827 & ~n4838;
  assign n4840 = n4827 & ~n4839;
  assign n4841 = ~n4838 & ~n4839;
  assign n4842 = ~n4840 & ~n4841;
  assign n4843 = ~n4614 & n4842;
  assign n4844 = n4614 & ~n4842;
  assign n4845 = ~n4843 & ~n4844;
  assign n4846 = n938 & n2446;
  assign n4847 = pi86  & n1052;
  assign n4848 = pi88  & n936;
  assign n4849 = pi87  & n931;
  assign n4850 = ~n4848 & ~n4849;
  assign n4851 = ~n4847 & n4850;
  assign n4852 = ~n4846 & n4851;
  assign n4853 = pi14  & ~n4852;
  assign n4854 = pi14  & ~n4853;
  assign n4855 = ~n4852 & ~n4853;
  assign n4856 = ~n4854 & ~n4855;
  assign n4857 = n4845 & n4856;
  assign n4858 = ~n4845 & ~n4856;
  assign n4859 = ~n4857 & ~n4858;
  assign n4860 = ~n4715 & n4859;
  assign n4861 = n4715 & ~n4859;
  assign n4862 = ~n4860 & ~n4861;
  assign n4863 = n687 & n2978;
  assign n4864 = pi89  & n763;
  assign n4865 = pi91  & n685;
  assign n4866 = pi90  & n680;
  assign n4867 = ~n4865 & ~n4866;
  assign n4868 = ~n4864 & n4867;
  assign n4869 = ~n4863 & n4868;
  assign n4870 = pi11  & ~n4869;
  assign n4871 = pi11  & ~n4870;
  assign n4872 = ~n4869 & ~n4870;
  assign n4873 = ~n4871 & ~n4872;
  assign n4874 = n4862 & ~n4873;
  assign n4875 = n4862 & ~n4874;
  assign n4876 = ~n4873 & ~n4874;
  assign n4877 = ~n4875 & ~n4876;
  assign n4878 = ~n4714 & n4877;
  assign n4879 = n4714 & ~n4877;
  assign n4880 = ~n4878 & ~n4879;
  assign n4881 = n498 & n3565;
  assign n4882 = pi92  & n537;
  assign n4883 = pi94  & n496;
  assign n4884 = pi93  & n491;
  assign n4885 = ~n4883 & ~n4884;
  assign n4886 = ~n4882 & n4885;
  assign n4887 = ~n4881 & n4886;
  assign n4888 = pi8  & ~n4887;
  assign n4889 = pi8  & ~n4888;
  assign n4890 = ~n4887 & ~n4888;
  assign n4891 = ~n4889 & ~n4890;
  assign n4892 = n4880 & n4891;
  assign n4893 = ~n4880 & ~n4891;
  assign n4894 = ~n4892 & ~n4893;
  assign n4895 = ~n4713 & n4894;
  assign n4896 = n4713 & ~n4894;
  assign n4897 = ~n4895 & ~n4896;
  assign n4898 = ~n4712 & n4897;
  assign n4899 = n4712 & ~n4897;
  assign n4900 = ~n4898 & ~n4899;
  assign n4901 = ~n4675 & n4900;
  assign n4902 = n4675 & ~n4900;
  assign n4903 = ~n4901 & ~n4902;
  assign n4904 = ~n4680 & ~n4682;
  assign n4905 = ~pi99  & ~pi100 ;
  assign n4906 = pi99  & pi100 ;
  assign n4907 = ~n4905 & ~n4906;
  assign n4908 = ~n4904 & n4907;
  assign n4909 = n4904 & ~n4907;
  assign n4910 = ~n4908 & ~n4909;
  assign n4911 = n262 & n4910;
  assign n4912 = pi98  & n288;
  assign n4913 = pi100  & n267;
  assign n4914 = pi99  & n269;
  assign n4915 = ~n4913 & ~n4914;
  assign n4916 = ~n4912 & n4915;
  assign n4917 = ~n4911 & n4916;
  assign n4918 = pi2  & ~n4917;
  assign n4919 = pi2  & ~n4918;
  assign n4920 = ~n4917 & ~n4918;
  assign n4921 = ~n4919 & ~n4920;
  assign n4922 = n4903 & ~n4921;
  assign n4923 = n4903 & ~n4922;
  assign n4924 = ~n4921 & ~n4922;
  assign n4925 = ~n4923 & ~n4924;
  assign n4926 = ~n4677 & ~n4695;
  assign n4927 = ~n4699 & ~n4926;
  assign n4928 = ~n4925 & ~n4927;
  assign n4929 = n4925 & n4927;
  assign po36  = ~n4928 & ~n4929;
  assign n4931 = ~n4922 & ~n4928;
  assign n4932 = ~n4893 & ~n4895;
  assign n4933 = n498 & n3784;
  assign n4934 = pi93  & n537;
  assign n4935 = pi95  & n496;
  assign n4936 = pi94  & n491;
  assign n4937 = ~n4935 & ~n4936;
  assign n4938 = ~n4934 & n4937;
  assign n4939 = ~n4933 & n4938;
  assign n4940 = pi8  & ~n4939;
  assign n4941 = pi8  & ~n4940;
  assign n4942 = ~n4939 & ~n4940;
  assign n4943 = ~n4941 & ~n4942;
  assign n4944 = ~n4714 & ~n4877;
  assign n4945 = ~n4874 & ~n4944;
  assign n4946 = ~n4858 & ~n4860;
  assign n4947 = ~n4787 & ~n4790;
  assign n4948 = n999 & n2523;
  assign n4949 = pi75  & n2667;
  assign n4950 = pi77  & n2521;
  assign n4951 = pi76  & n2516;
  assign n4952 = ~n4950 & ~n4951;
  assign n4953 = ~n4949 & n4952;
  assign n4954 = ~n4948 & n4953;
  assign n4955 = pi26  & ~n4954;
  assign n4956 = pi26  & ~n4955;
  assign n4957 = ~n4954 & ~n4955;
  assign n4958 = ~n4956 & ~n4957;
  assign n4959 = ~n4769 & ~n4773;
  assign n4960 = n729 & n3034;
  assign n4961 = pi72  & n3225;
  assign n4962 = pi74  & n3032;
  assign n4963 = pi73  & n3027;
  assign n4964 = ~n4962 & ~n4963;
  assign n4965 = ~n4961 & n4964;
  assign n4966 = ~n4960 & n4965;
  assign n4967 = pi29  & ~n4966;
  assign n4968 = pi29  & ~n4967;
  assign n4969 = ~n4966 & ~n4967;
  assign n4970 = ~n4968 & ~n4969;
  assign n4971 = ~n4533 & ~n4754;
  assign n4972 = ~n4751 & ~n4971;
  assign n4973 = n475 & n3622;
  assign n4974 = pi69  & n3814;
  assign n4975 = pi71  & n3620;
  assign n4976 = pi70  & n3615;
  assign n4977 = ~n4975 & ~n4976;
  assign n4978 = ~n4974 & n4977;
  assign n4979 = ~n4973 & n4978;
  assign n4980 = pi32  & ~n4979;
  assign n4981 = pi32  & ~n4980;
  assign n4982 = ~n4979 & ~n4980;
  assign n4983 = ~n4981 & ~n4982;
  assign n4984 = n4515 & n4722;
  assign n4985 = ~n4737 & ~n4984;
  assign n4986 = n359 & n4271;
  assign n4987 = pi66  & n4503;
  assign n4988 = pi68  & n4269;
  assign n4989 = pi67  & n4264;
  assign n4990 = ~n4988 & ~n4989;
  assign n4991 = ~n4987 & n4990;
  assign n4992 = ~n4986 & n4991;
  assign n4993 = pi35  & ~n4992;
  assign n4994 = pi35  & ~n4993;
  assign n4995 = ~n4992 & ~n4993;
  assign n4996 = ~n4994 & ~n4995;
  assign n4997 = pi38  & ~n4722;
  assign n4998 = ~pi36  & pi37 ;
  assign n4999 = pi36  & ~pi37 ;
  assign n5000 = ~n4998 & ~n4999;
  assign n5001 = n4721 & ~n5000;
  assign n5002 = pi64  & n5001;
  assign n5003 = ~pi37  & pi38 ;
  assign n5004 = pi37  & ~pi38 ;
  assign n5005 = ~n5003 & ~n5004;
  assign n5006 = ~n4721 & n5005;
  assign n5007 = pi65  & n5006;
  assign n5008 = ~n4721 & ~n5005;
  assign n5009 = ~n265 & n5008;
  assign n5010 = ~n5002 & ~n5007;
  assign n5011 = ~n5009 & n5010;
  assign n5012 = pi38  & ~n5011;
  assign n5013 = pi38  & ~n5012;
  assign n5014 = ~n5011 & ~n5012;
  assign n5015 = ~n5013 & ~n5014;
  assign n5016 = n4997 & ~n5015;
  assign n5017 = ~n4997 & n5015;
  assign n5018 = ~n5016 & ~n5017;
  assign n5019 = n4996 & ~n5018;
  assign n5020 = ~n4996 & n5018;
  assign n5021 = ~n5019 & ~n5020;
  assign n5022 = ~n4985 & n5021;
  assign n5023 = n4985 & ~n5021;
  assign n5024 = ~n5022 & ~n5023;
  assign n5025 = n4983 & ~n5024;
  assign n5026 = ~n4983 & n5024;
  assign n5027 = ~n5025 & ~n5026;
  assign n5028 = ~n4972 & n5027;
  assign n5029 = n4972 & ~n5027;
  assign n5030 = ~n5028 & ~n5029;
  assign n5031 = n4970 & ~n5030;
  assign n5032 = ~n4970 & n5030;
  assign n5033 = ~n5031 & ~n5032;
  assign n5034 = ~n4959 & n5033;
  assign n5035 = n4959 & ~n5033;
  assign n5036 = ~n5034 & ~n5035;
  assign n5037 = n4958 & ~n5036;
  assign n5038 = ~n4958 & n5036;
  assign n5039 = ~n5037 & ~n5038;
  assign n5040 = ~n4947 & n5039;
  assign n5041 = n4947 & ~n5039;
  assign n5042 = ~n5040 & ~n5041;
  assign n5043 = n1225 & n2043;
  assign n5044 = pi78  & n2180;
  assign n5045 = pi80  & n2041;
  assign n5046 = pi79  & n2036;
  assign n5047 = ~n5045 & ~n5046;
  assign n5048 = ~n5044 & n5047;
  assign n5049 = ~n5043 & n5048;
  assign n5050 = pi23  & ~n5049;
  assign n5051 = pi23  & ~n5050;
  assign n5052 = ~n5049 & ~n5050;
  assign n5053 = ~n5051 & ~n5052;
  assign n5054 = n5042 & ~n5053;
  assign n5055 = n5042 & ~n5054;
  assign n5056 = ~n5053 & ~n5054;
  assign n5057 = ~n5055 & ~n5056;
  assign n5058 = ~n4717 & ~n4807;
  assign n5059 = ~n4804 & ~n5058;
  assign n5060 = n5057 & n5059;
  assign n5061 = ~n5057 & ~n5059;
  assign n5062 = ~n5060 & ~n5061;
  assign n5063 = n1611 & n1696;
  assign n5064 = pi81  & n1745;
  assign n5065 = pi83  & n1609;
  assign n5066 = pi82  & n1604;
  assign n5067 = ~n5065 & ~n5066;
  assign n5068 = ~n5064 & n5067;
  assign n5069 = ~n5063 & n5068;
  assign n5070 = pi20  & ~n5069;
  assign n5071 = pi20  & ~n5070;
  assign n5072 = ~n5069 & ~n5070;
  assign n5073 = ~n5071 & ~n5072;
  assign n5074 = n5062 & ~n5073;
  assign n5075 = n5062 & ~n5074;
  assign n5076 = ~n5073 & ~n5074;
  assign n5077 = ~n5075 & ~n5076;
  assign n5078 = ~n4822 & ~n4826;
  assign n5079 = n5077 & n5078;
  assign n5080 = ~n5077 & ~n5078;
  assign n5081 = ~n5079 & ~n5080;
  assign n5082 = n1297 & n2133;
  assign n5083 = pi84  & n1366;
  assign n5084 = pi86  & n1295;
  assign n5085 = pi85  & n1290;
  assign n5086 = ~n5084 & ~n5085;
  assign n5087 = ~n5083 & n5086;
  assign n5088 = ~n5082 & n5087;
  assign n5089 = pi17  & ~n5088;
  assign n5090 = pi17  & ~n5089;
  assign n5091 = ~n5088 & ~n5089;
  assign n5092 = ~n5090 & ~n5091;
  assign n5093 = n5081 & ~n5092;
  assign n5094 = n5081 & ~n5093;
  assign n5095 = ~n5092 & ~n5093;
  assign n5096 = ~n5094 & ~n5095;
  assign n5097 = ~n4614 & ~n4842;
  assign n5098 = ~n4839 & ~n5097;
  assign n5099 = n5096 & n5098;
  assign n5100 = ~n5096 & ~n5098;
  assign n5101 = ~n5099 & ~n5100;
  assign n5102 = n938 & n2473;
  assign n5103 = pi87  & n1052;
  assign n5104 = pi89  & n936;
  assign n5105 = pi88  & n931;
  assign n5106 = ~n5104 & ~n5105;
  assign n5107 = ~n5103 & n5106;
  assign n5108 = ~n5102 & n5107;
  assign n5109 = pi14  & ~n5108;
  assign n5110 = pi14  & ~n5109;
  assign n5111 = ~n5108 & ~n5109;
  assign n5112 = ~n5110 & ~n5111;
  assign n5113 = n5101 & ~n5112;
  assign n5114 = ~n5101 & n5112;
  assign n5115 = ~n5113 & ~n5114;
  assign n5116 = ~n4946 & n5115;
  assign n5117 = ~n4946 & ~n5116;
  assign n5118 = ~n5113 & ~n5116;
  assign n5119 = ~n5114 & n5118;
  assign n5120 = ~n5117 & ~n5119;
  assign n5121 = n687 & n3177;
  assign n5122 = pi90  & n763;
  assign n5123 = pi92  & n685;
  assign n5124 = pi91  & n680;
  assign n5125 = ~n5123 & ~n5124;
  assign n5126 = ~n5122 & n5125;
  assign n5127 = ~n5121 & n5126;
  assign n5128 = pi11  & ~n5127;
  assign n5129 = pi11  & ~n5128;
  assign n5130 = ~n5127 & ~n5128;
  assign n5131 = ~n5129 & ~n5130;
  assign n5132 = n5120 & n5131;
  assign n5133 = ~n5120 & ~n5131;
  assign n5134 = ~n5132 & ~n5133;
  assign n5135 = ~n4945 & n5134;
  assign n5136 = n4945 & ~n5134;
  assign n5137 = ~n5135 & ~n5136;
  assign n5138 = n4943 & ~n5137;
  assign n5139 = ~n4943 & n5137;
  assign n5140 = ~n5138 & ~n5139;
  assign n5141 = ~n4932 & n5140;
  assign n5142 = n4932 & ~n5140;
  assign n5143 = ~n5141 & ~n5142;
  assign n5144 = n342 & n4454;
  assign n5145 = pi96  & n380;
  assign n5146 = pi98  & n340;
  assign n5147 = pi97  & n335;
  assign n5148 = ~n5146 & ~n5147;
  assign n5149 = ~n5145 & n5148;
  assign n5150 = ~n5144 & n5149;
  assign n5151 = pi5  & ~n5150;
  assign n5152 = pi5  & ~n5151;
  assign n5153 = ~n5150 & ~n5151;
  assign n5154 = ~n5152 & ~n5153;
  assign n5155 = n5143 & ~n5154;
  assign n5156 = n5143 & ~n5155;
  assign n5157 = ~n5154 & ~n5155;
  assign n5158 = ~n5156 & ~n5157;
  assign n5159 = ~n4898 & ~n4901;
  assign n5160 = n5158 & n5159;
  assign n5161 = ~n5158 & ~n5159;
  assign n5162 = ~n5160 & ~n5161;
  assign n5163 = ~n4906 & ~n4908;
  assign n5164 = ~pi100  & ~pi101 ;
  assign n5165 = pi100  & pi101 ;
  assign n5166 = ~n5164 & ~n5165;
  assign n5167 = ~n5163 & n5166;
  assign n5168 = n5163 & ~n5166;
  assign n5169 = ~n5167 & ~n5168;
  assign n5170 = n262 & n5169;
  assign n5171 = pi99  & n288;
  assign n5172 = pi101  & n267;
  assign n5173 = pi100  & n269;
  assign n5174 = ~n5172 & ~n5173;
  assign n5175 = ~n5171 & n5174;
  assign n5176 = ~n5170 & n5175;
  assign n5177 = pi2  & ~n5176;
  assign n5178 = pi2  & ~n5177;
  assign n5179 = ~n5176 & ~n5177;
  assign n5180 = ~n5178 & ~n5179;
  assign n5181 = ~n5162 & n5180;
  assign n5182 = n5162 & ~n5180;
  assign n5183 = ~n5181 & ~n5182;
  assign n5184 = ~n4931 & n5183;
  assign n5185 = n4931 & ~n5183;
  assign po37  = ~n5184 & ~n5185;
  assign n5187 = ~n5155 & ~n5161;
  assign n5188 = n342 & n4684;
  assign n5189 = pi97  & n380;
  assign n5190 = pi99  & n340;
  assign n5191 = pi98  & n335;
  assign n5192 = ~n5190 & ~n5191;
  assign n5193 = ~n5189 & n5192;
  assign n5194 = ~n5188 & n5193;
  assign n5195 = pi5  & ~n5194;
  assign n5196 = pi5  & ~n5195;
  assign n5197 = ~n5194 & ~n5195;
  assign n5198 = ~n5196 & ~n5197;
  assign n5199 = ~n5139 & ~n5141;
  assign n5200 = n498 & n4001;
  assign n5201 = pi94  & n537;
  assign n5202 = pi96  & n496;
  assign n5203 = pi95  & n491;
  assign n5204 = ~n5202 & ~n5203;
  assign n5205 = ~n5201 & n5204;
  assign n5206 = ~n5200 & n5205;
  assign n5207 = pi8  & ~n5206;
  assign n5208 = pi8  & ~n5207;
  assign n5209 = ~n5206 & ~n5207;
  assign n5210 = ~n5208 & ~n5209;
  assign n5211 = ~n5133 & ~n5135;
  assign n5212 = n687 & n3371;
  assign n5213 = pi91  & n763;
  assign n5214 = pi93  & n685;
  assign n5215 = pi92  & n680;
  assign n5216 = ~n5214 & ~n5215;
  assign n5217 = ~n5213 & n5216;
  assign n5218 = ~n5212 & n5217;
  assign n5219 = pi11  & ~n5218;
  assign n5220 = pi11  & ~n5219;
  assign n5221 = ~n5218 & ~n5219;
  assign n5222 = ~n5220 & ~n5221;
  assign n5223 = ~n5093 & ~n5100;
  assign n5224 = ~n5038 & ~n5040;
  assign n5225 = ~n5032 & ~n5034;
  assign n5226 = n809 & n3034;
  assign n5227 = pi73  & n3225;
  assign n5228 = pi75  & n3032;
  assign n5229 = pi74  & n3027;
  assign n5230 = ~n5228 & ~n5229;
  assign n5231 = ~n5227 & n5230;
  assign n5232 = ~n5226 & n5231;
  assign n5233 = pi29  & ~n5232;
  assign n5234 = pi29  & ~n5233;
  assign n5235 = ~n5232 & ~n5233;
  assign n5236 = ~n5234 & ~n5235;
  assign n5237 = ~n5026 & ~n5028;
  assign n5238 = ~n5020 & ~n5022;
  assign n5239 = n286 & n5008;
  assign n5240 = n4721 & n5000;
  assign n5241 = ~n5005 & n5240;
  assign n5242 = pi64  & n5241;
  assign n5243 = pi66  & n5006;
  assign n5244 = pi65  & n5001;
  assign n5245 = ~n5243 & ~n5244;
  assign n5246 = ~n5239 & n5245;
  assign n5247 = ~n5242 & n5246;
  assign n5248 = pi38  & ~n5247;
  assign n5249 = pi38  & ~n5248;
  assign n5250 = ~n5247 & ~n5248;
  assign n5251 = ~n5249 & ~n5250;
  assign n5252 = ~n5016 & n5251;
  assign n5253 = n5016 & ~n5251;
  assign n5254 = ~n5252 & ~n5253;
  assign n5255 = n401 & n4271;
  assign n5256 = pi67  & n4503;
  assign n5257 = pi69  & n4269;
  assign n5258 = pi68  & n4264;
  assign n5259 = ~n5257 & ~n5258;
  assign n5260 = ~n5256 & n5259;
  assign n5261 = ~n5255 & n5260;
  assign n5262 = pi35  & ~n5261;
  assign n5263 = pi35  & ~n5262;
  assign n5264 = ~n5261 & ~n5262;
  assign n5265 = ~n5263 & ~n5264;
  assign n5266 = n5254 & ~n5265;
  assign n5267 = n5254 & ~n5266;
  assign n5268 = ~n5265 & ~n5266;
  assign n5269 = ~n5267 & ~n5268;
  assign n5270 = ~n5238 & n5269;
  assign n5271 = n5238 & ~n5269;
  assign n5272 = ~n5270 & ~n5271;
  assign n5273 = n576 & n3622;
  assign n5274 = pi70  & n3814;
  assign n5275 = pi72  & n3620;
  assign n5276 = pi71  & n3615;
  assign n5277 = ~n5275 & ~n5276;
  assign n5278 = ~n5274 & n5277;
  assign n5279 = ~n5273 & n5278;
  assign n5280 = pi32  & ~n5279;
  assign n5281 = pi32  & ~n5280;
  assign n5282 = ~n5279 & ~n5280;
  assign n5283 = ~n5281 & ~n5282;
  assign n5284 = ~n5272 & ~n5283;
  assign n5285 = n5272 & n5283;
  assign n5286 = ~n5284 & ~n5285;
  assign n5287 = ~n5237 & n5286;
  assign n5288 = n5237 & ~n5286;
  assign n5289 = ~n5287 & ~n5288;
  assign n5290 = ~n5236 & n5289;
  assign n5291 = ~n5236 & ~n5290;
  assign n5292 = n5289 & ~n5290;
  assign n5293 = ~n5291 & ~n5292;
  assign n5294 = ~n5225 & ~n5293;
  assign n5295 = ~n5225 & ~n5294;
  assign n5296 = ~n5293 & ~n5294;
  assign n5297 = ~n5295 & ~n5296;
  assign n5298 = n1025 & n2523;
  assign n5299 = pi76  & n2667;
  assign n5300 = pi78  & n2521;
  assign n5301 = pi77  & n2516;
  assign n5302 = ~n5300 & ~n5301;
  assign n5303 = ~n5299 & n5302;
  assign n5304 = ~n5298 & n5303;
  assign n5305 = pi26  & ~n5304;
  assign n5306 = pi26  & ~n5305;
  assign n5307 = ~n5304 & ~n5305;
  assign n5308 = ~n5306 & ~n5307;
  assign n5309 = n5297 & n5308;
  assign n5310 = ~n5297 & ~n5308;
  assign n5311 = ~n5309 & ~n5310;
  assign n5312 = ~n5224 & n5311;
  assign n5313 = n5224 & ~n5311;
  assign n5314 = ~n5312 & ~n5313;
  assign n5315 = n1434 & n2043;
  assign n5316 = pi79  & n2180;
  assign n5317 = pi81  & n2041;
  assign n5318 = pi80  & n2036;
  assign n5319 = ~n5317 & ~n5318;
  assign n5320 = ~n5316 & n5319;
  assign n5321 = ~n5315 & n5320;
  assign n5322 = pi23  & ~n5321;
  assign n5323 = pi23  & ~n5322;
  assign n5324 = ~n5321 & ~n5322;
  assign n5325 = ~n5323 & ~n5324;
  assign n5326 = n5314 & ~n5325;
  assign n5327 = n5314 & ~n5326;
  assign n5328 = ~n5325 & ~n5326;
  assign n5329 = ~n5327 & ~n5328;
  assign n5330 = ~n5054 & ~n5061;
  assign n5331 = n5329 & n5330;
  assign n5332 = ~n5329 & ~n5330;
  assign n5333 = ~n5331 & ~n5332;
  assign n5334 = n1611 & n1834;
  assign n5335 = pi82  & n1745;
  assign n5336 = pi84  & n1609;
  assign n5337 = pi83  & n1604;
  assign n5338 = ~n5336 & ~n5337;
  assign n5339 = ~n5335 & n5338;
  assign n5340 = ~n5334 & n5339;
  assign n5341 = pi20  & ~n5340;
  assign n5342 = pi20  & ~n5341;
  assign n5343 = ~n5340 & ~n5341;
  assign n5344 = ~n5342 & ~n5343;
  assign n5345 = n5333 & ~n5344;
  assign n5346 = n5333 & ~n5345;
  assign n5347 = ~n5344 & ~n5345;
  assign n5348 = ~n5346 & ~n5347;
  assign n5349 = ~n5074 & ~n5080;
  assign n5350 = n5348 & n5349;
  assign n5351 = ~n5348 & ~n5349;
  assign n5352 = ~n5350 & ~n5351;
  assign n5353 = n1297 & n2288;
  assign n5354 = pi85  & n1366;
  assign n5355 = pi87  & n1295;
  assign n5356 = pi86  & n1290;
  assign n5357 = ~n5355 & ~n5356;
  assign n5358 = ~n5354 & n5357;
  assign n5359 = ~n5353 & n5358;
  assign n5360 = pi17  & ~n5359;
  assign n5361 = pi17  & ~n5360;
  assign n5362 = ~n5359 & ~n5360;
  assign n5363 = ~n5361 & ~n5362;
  assign n5364 = n5352 & ~n5363;
  assign n5365 = ~n5352 & n5363;
  assign n5366 = ~n5364 & ~n5365;
  assign n5367 = ~n5223 & n5366;
  assign n5368 = ~n5223 & ~n5367;
  assign n5369 = ~n5364 & ~n5367;
  assign n5370 = ~n5365 & n5369;
  assign n5371 = ~n5368 & ~n5370;
  assign n5372 = n938 & n2801;
  assign n5373 = pi88  & n1052;
  assign n5374 = pi90  & n936;
  assign n5375 = pi89  & n931;
  assign n5376 = ~n5374 & ~n5375;
  assign n5377 = ~n5373 & n5376;
  assign n5378 = ~n5372 & n5377;
  assign n5379 = pi14  & ~n5378;
  assign n5380 = pi14  & ~n5379;
  assign n5381 = ~n5378 & ~n5379;
  assign n5382 = ~n5380 & ~n5381;
  assign n5383 = n5371 & n5382;
  assign n5384 = ~n5371 & ~n5382;
  assign n5385 = ~n5383 & ~n5384;
  assign n5386 = ~n5118 & n5385;
  assign n5387 = n5118 & ~n5385;
  assign n5388 = ~n5386 & ~n5387;
  assign n5389 = n5222 & ~n5388;
  assign n5390 = ~n5222 & n5388;
  assign n5391 = ~n5389 & ~n5390;
  assign n5392 = ~n5211 & n5391;
  assign n5393 = n5211 & ~n5391;
  assign n5394 = ~n5392 & ~n5393;
  assign n5395 = n5210 & ~n5394;
  assign n5396 = ~n5210 & n5394;
  assign n5397 = ~n5395 & ~n5396;
  assign n5398 = ~n5199 & n5397;
  assign n5399 = n5199 & ~n5397;
  assign n5400 = ~n5398 & ~n5399;
  assign n5401 = n5198 & ~n5400;
  assign n5402 = ~n5198 & n5400;
  assign n5403 = ~n5401 & ~n5402;
  assign n5404 = ~n5187 & n5403;
  assign n5405 = n5187 & ~n5403;
  assign n5406 = ~n5404 & ~n5405;
  assign n5407 = ~n5165 & ~n5167;
  assign n5408 = ~pi101  & ~pi102 ;
  assign n5409 = pi101  & pi102 ;
  assign n5410 = ~n5408 & ~n5409;
  assign n5411 = ~n5407 & n5410;
  assign n5412 = n5407 & ~n5410;
  assign n5413 = ~n5411 & ~n5412;
  assign n5414 = n262 & n5413;
  assign n5415 = pi100  & n288;
  assign n5416 = pi102  & n267;
  assign n5417 = pi101  & n269;
  assign n5418 = ~n5416 & ~n5417;
  assign n5419 = ~n5415 & n5418;
  assign n5420 = ~n5414 & n5419;
  assign n5421 = pi2  & ~n5420;
  assign n5422 = pi2  & ~n5421;
  assign n5423 = ~n5420 & ~n5421;
  assign n5424 = ~n5422 & ~n5423;
  assign n5425 = n5406 & ~n5424;
  assign n5426 = n5406 & ~n5425;
  assign n5427 = ~n5424 & ~n5425;
  assign n5428 = ~n5426 & ~n5427;
  assign n5429 = ~n5182 & ~n5184;
  assign n5430 = ~n5428 & ~n5429;
  assign n5431 = n5428 & n5429;
  assign po38  = ~n5430 & ~n5431;
  assign n5433 = ~n5402 & ~n5404;
  assign n5434 = ~n5396 & ~n5398;
  assign n5435 = ~n5390 & ~n5392;
  assign n5436 = ~n5384 & ~n5386;
  assign n5437 = ~n5326 & ~n5332;
  assign n5438 = ~n5310 & ~n5312;
  assign n5439 = pi38  & ~pi39 ;
  assign n5440 = ~pi38  & pi39 ;
  assign n5441 = ~n5439 & ~n5440;
  assign n5442 = pi64  & ~n5441;
  assign n5443 = ~n5253 & n5442;
  assign n5444 = n5253 & ~n5442;
  assign n5445 = ~n5443 & ~n5444;
  assign n5446 = n309 & n5008;
  assign n5447 = pi65  & n5241;
  assign n5448 = pi67  & n5006;
  assign n5449 = pi66  & n5001;
  assign n5450 = ~n5448 & ~n5449;
  assign n5451 = ~n5447 & n5450;
  assign n5452 = ~n5446 & n5451;
  assign n5453 = pi38  & ~n5452;
  assign n5454 = pi38  & ~n5453;
  assign n5455 = ~n5452 & ~n5453;
  assign n5456 = ~n5454 & ~n5455;
  assign n5457 = ~n5445 & ~n5456;
  assign n5458 = n5445 & n5456;
  assign n5459 = ~n5457 & ~n5458;
  assign n5460 = n450 & n4271;
  assign n5461 = pi68  & n4503;
  assign n5462 = pi70  & n4269;
  assign n5463 = pi69  & n4264;
  assign n5464 = ~n5462 & ~n5463;
  assign n5465 = ~n5461 & n5464;
  assign n5466 = ~n5460 & n5465;
  assign n5467 = pi35  & ~n5466;
  assign n5468 = pi35  & ~n5467;
  assign n5469 = ~n5466 & ~n5467;
  assign n5470 = ~n5468 & ~n5469;
  assign n5471 = n5459 & ~n5470;
  assign n5472 = n5459 & ~n5471;
  assign n5473 = ~n5470 & ~n5471;
  assign n5474 = ~n5472 & ~n5473;
  assign n5475 = ~n5238 & ~n5269;
  assign n5476 = ~n5266 & ~n5475;
  assign n5477 = n5474 & n5476;
  assign n5478 = ~n5474 & ~n5476;
  assign n5479 = ~n5477 & ~n5478;
  assign n5480 = n642 & n3622;
  assign n5481 = pi71  & n3814;
  assign n5482 = pi73  & n3620;
  assign n5483 = pi72  & n3615;
  assign n5484 = ~n5482 & ~n5483;
  assign n5485 = ~n5481 & n5484;
  assign n5486 = ~n5480 & n5485;
  assign n5487 = pi32  & ~n5486;
  assign n5488 = pi32  & ~n5487;
  assign n5489 = ~n5486 & ~n5487;
  assign n5490 = ~n5488 & ~n5489;
  assign n5491 = n5479 & ~n5490;
  assign n5492 = n5479 & ~n5491;
  assign n5493 = ~n5490 & ~n5491;
  assign n5494 = ~n5492 & ~n5493;
  assign n5495 = ~n5284 & ~n5287;
  assign n5496 = n5494 & n5495;
  assign n5497 = ~n5494 & ~n5495;
  assign n5498 = ~n5496 & ~n5497;
  assign n5499 = n891 & n3034;
  assign n5500 = pi74  & n3225;
  assign n5501 = pi76  & n3032;
  assign n5502 = pi75  & n3027;
  assign n5503 = ~n5501 & ~n5502;
  assign n5504 = ~n5500 & n5503;
  assign n5505 = ~n5499 & n5504;
  assign n5506 = pi29  & ~n5505;
  assign n5507 = pi29  & ~n5506;
  assign n5508 = ~n5505 & ~n5506;
  assign n5509 = ~n5507 & ~n5508;
  assign n5510 = ~n5498 & n5509;
  assign n5511 = n5498 & ~n5509;
  assign n5512 = ~n5510 & ~n5511;
  assign n5513 = ~n5290 & ~n5294;
  assign n5514 = n5512 & ~n5513;
  assign n5515 = ~n5512 & n5513;
  assign n5516 = ~n5514 & ~n5515;
  assign n5517 = n1122 & n2523;
  assign n5518 = pi77  & n2667;
  assign n5519 = pi79  & n2521;
  assign n5520 = pi78  & n2516;
  assign n5521 = ~n5519 & ~n5520;
  assign n5522 = ~n5518 & n5521;
  assign n5523 = ~n5517 & n5522;
  assign n5524 = pi26  & ~n5523;
  assign n5525 = pi26  & ~n5524;
  assign n5526 = ~n5523 & ~n5524;
  assign n5527 = ~n5525 & ~n5526;
  assign n5528 = n5516 & ~n5527;
  assign n5529 = n5516 & ~n5528;
  assign n5530 = ~n5527 & ~n5528;
  assign n5531 = ~n5529 & ~n5530;
  assign n5532 = ~n5438 & n5531;
  assign n5533 = n5438 & ~n5531;
  assign n5534 = ~n5532 & ~n5533;
  assign n5535 = n1554 & n2043;
  assign n5536 = pi80  & n2180;
  assign n5537 = pi82  & n2041;
  assign n5538 = pi81  & n2036;
  assign n5539 = ~n5537 & ~n5538;
  assign n5540 = ~n5536 & n5539;
  assign n5541 = ~n5535 & n5540;
  assign n5542 = pi23  & ~n5541;
  assign n5543 = pi23  & ~n5542;
  assign n5544 = ~n5541 & ~n5542;
  assign n5545 = ~n5543 & ~n5544;
  assign n5546 = ~n5534 & ~n5545;
  assign n5547 = n5534 & n5545;
  assign n5548 = ~n5546 & ~n5547;
  assign n5549 = n5437 & ~n5548;
  assign n5550 = ~n5437 & n5548;
  assign n5551 = ~n5549 & ~n5550;
  assign n5552 = n1611 & n1972;
  assign n5553 = pi83  & n1745;
  assign n5554 = pi85  & n1609;
  assign n5555 = pi84  & n1604;
  assign n5556 = ~n5554 & ~n5555;
  assign n5557 = ~n5553 & n5556;
  assign n5558 = ~n5552 & n5557;
  assign n5559 = pi20  & ~n5558;
  assign n5560 = pi20  & ~n5559;
  assign n5561 = ~n5558 & ~n5559;
  assign n5562 = ~n5560 & ~n5561;
  assign n5563 = n5551 & ~n5562;
  assign n5564 = n5551 & ~n5563;
  assign n5565 = ~n5562 & ~n5563;
  assign n5566 = ~n5564 & ~n5565;
  assign n5567 = ~n5345 & ~n5351;
  assign n5568 = n5566 & n5567;
  assign n5569 = ~n5566 & ~n5567;
  assign n5570 = ~n5568 & ~n5569;
  assign n5571 = n1297 & n2446;
  assign n5572 = pi86  & n1366;
  assign n5573 = pi88  & n1295;
  assign n5574 = pi87  & n1290;
  assign n5575 = ~n5573 & ~n5574;
  assign n5576 = ~n5572 & n5575;
  assign n5577 = ~n5571 & n5576;
  assign n5578 = pi17  & ~n5577;
  assign n5579 = pi17  & ~n5578;
  assign n5580 = ~n5577 & ~n5578;
  assign n5581 = ~n5579 & ~n5580;
  assign n5582 = ~n5570 & n5581;
  assign n5583 = n5570 & ~n5581;
  assign n5584 = ~n5582 & ~n5583;
  assign n5585 = ~n5369 & n5584;
  assign n5586 = n5369 & ~n5584;
  assign n5587 = ~n5585 & ~n5586;
  assign n5588 = n938 & n2978;
  assign n5589 = pi89  & n1052;
  assign n5590 = pi91  & n936;
  assign n5591 = pi90  & n931;
  assign n5592 = ~n5590 & ~n5591;
  assign n5593 = ~n5589 & n5592;
  assign n5594 = ~n5588 & n5593;
  assign n5595 = pi14  & ~n5594;
  assign n5596 = pi14  & ~n5595;
  assign n5597 = ~n5594 & ~n5595;
  assign n5598 = ~n5596 & ~n5597;
  assign n5599 = n5587 & ~n5598;
  assign n5600 = n5587 & ~n5599;
  assign n5601 = ~n5598 & ~n5599;
  assign n5602 = ~n5600 & ~n5601;
  assign n5603 = ~n5436 & n5602;
  assign n5604 = n5436 & ~n5602;
  assign n5605 = ~n5603 & ~n5604;
  assign n5606 = n687 & n3565;
  assign n5607 = pi92  & n763;
  assign n5608 = pi94  & n685;
  assign n5609 = pi93  & n680;
  assign n5610 = ~n5608 & ~n5609;
  assign n5611 = ~n5607 & n5610;
  assign n5612 = ~n5606 & n5611;
  assign n5613 = pi11  & ~n5612;
  assign n5614 = pi11  & ~n5613;
  assign n5615 = ~n5612 & ~n5613;
  assign n5616 = ~n5614 & ~n5615;
  assign n5617 = ~n5605 & ~n5616;
  assign n5618 = n5605 & n5616;
  assign n5619 = ~n5617 & ~n5618;
  assign n5620 = ~n5435 & n5619;
  assign n5621 = n5435 & ~n5619;
  assign n5622 = ~n5620 & ~n5621;
  assign n5623 = n498 & n4211;
  assign n5624 = pi95  & n537;
  assign n5625 = pi97  & n496;
  assign n5626 = pi96  & n491;
  assign n5627 = ~n5625 & ~n5626;
  assign n5628 = ~n5624 & n5627;
  assign n5629 = ~n5623 & n5628;
  assign n5630 = pi8  & ~n5629;
  assign n5631 = pi8  & ~n5630;
  assign n5632 = ~n5629 & ~n5630;
  assign n5633 = ~n5631 & ~n5632;
  assign n5634 = n5622 & ~n5633;
  assign n5635 = n5622 & ~n5634;
  assign n5636 = ~n5633 & ~n5634;
  assign n5637 = ~n5635 & ~n5636;
  assign n5638 = ~n5434 & n5637;
  assign n5639 = n5434 & ~n5637;
  assign n5640 = ~n5638 & ~n5639;
  assign n5641 = n342 & n4910;
  assign n5642 = pi98  & n380;
  assign n5643 = pi100  & n340;
  assign n5644 = pi99  & n335;
  assign n5645 = ~n5643 & ~n5644;
  assign n5646 = ~n5642 & n5645;
  assign n5647 = ~n5641 & n5646;
  assign n5648 = pi5  & ~n5647;
  assign n5649 = pi5  & ~n5648;
  assign n5650 = ~n5647 & ~n5648;
  assign n5651 = ~n5649 & ~n5650;
  assign n5652 = n5640 & n5651;
  assign n5653 = ~n5640 & ~n5651;
  assign n5654 = ~n5652 & ~n5653;
  assign n5655 = ~n5433 & n5654;
  assign n5656 = n5433 & ~n5654;
  assign n5657 = ~n5655 & ~n5656;
  assign n5658 = ~n5409 & ~n5411;
  assign n5659 = ~pi102  & ~pi103 ;
  assign n5660 = pi102  & pi103 ;
  assign n5661 = ~n5659 & ~n5660;
  assign n5662 = ~n5658 & n5661;
  assign n5663 = n5658 & ~n5661;
  assign n5664 = ~n5662 & ~n5663;
  assign n5665 = n262 & n5664;
  assign n5666 = pi101  & n288;
  assign n5667 = pi103  & n267;
  assign n5668 = pi102  & n269;
  assign n5669 = ~n5667 & ~n5668;
  assign n5670 = ~n5666 & n5669;
  assign n5671 = ~n5665 & n5670;
  assign n5672 = pi2  & ~n5671;
  assign n5673 = pi2  & ~n5672;
  assign n5674 = ~n5671 & ~n5672;
  assign n5675 = ~n5673 & ~n5674;
  assign n5676 = n5657 & ~n5675;
  assign n5677 = n5657 & ~n5676;
  assign n5678 = ~n5675 & ~n5676;
  assign n5679 = ~n5677 & ~n5678;
  assign n5680 = ~n5425 & ~n5430;
  assign n5681 = ~n5679 & ~n5680;
  assign n5682 = n5679 & n5680;
  assign po39  = ~n5681 & ~n5682;
  assign n5684 = ~n5676 & ~n5681;
  assign n5685 = ~n5653 & ~n5655;
  assign n5686 = ~n5434 & ~n5637;
  assign n5687 = ~n5634 & ~n5686;
  assign n5688 = n498 & n4454;
  assign n5689 = pi96  & n537;
  assign n5690 = pi98  & n496;
  assign n5691 = pi97  & n491;
  assign n5692 = ~n5690 & ~n5691;
  assign n5693 = ~n5689 & n5692;
  assign n5694 = ~n5688 & n5693;
  assign n5695 = pi8  & ~n5694;
  assign n5696 = pi8  & ~n5695;
  assign n5697 = ~n5694 & ~n5695;
  assign n5698 = ~n5696 & ~n5697;
  assign n5699 = ~n5617 & ~n5620;
  assign n5700 = ~n5436 & ~n5602;
  assign n5701 = ~n5599 & ~n5700;
  assign n5702 = n938 & n3177;
  assign n5703 = pi90  & n1052;
  assign n5704 = pi92  & n936;
  assign n5705 = pi91  & n931;
  assign n5706 = ~n5704 & ~n5705;
  assign n5707 = ~n5703 & n5706;
  assign n5708 = ~n5702 & n5707;
  assign n5709 = pi14  & ~n5708;
  assign n5710 = pi14  & ~n5709;
  assign n5711 = ~n5708 & ~n5709;
  assign n5712 = ~n5710 & ~n5711;
  assign n5713 = ~n5511 & ~n5514;
  assign n5714 = ~n5491 & ~n5497;
  assign n5715 = n5253 & n5442;
  assign n5716 = ~n5457 & ~n5715;
  assign n5717 = n359 & n5008;
  assign n5718 = pi66  & n5241;
  assign n5719 = pi68  & n5006;
  assign n5720 = pi67  & n5001;
  assign n5721 = ~n5719 & ~n5720;
  assign n5722 = ~n5718 & n5721;
  assign n5723 = ~n5717 & n5722;
  assign n5724 = pi38  & ~n5723;
  assign n5725 = pi38  & ~n5724;
  assign n5726 = ~n5723 & ~n5724;
  assign n5727 = ~n5725 & ~n5726;
  assign n5728 = pi41  & ~n5442;
  assign n5729 = ~pi39  & pi40 ;
  assign n5730 = pi39  & ~pi40 ;
  assign n5731 = ~n5729 & ~n5730;
  assign n5732 = n5441 & ~n5731;
  assign n5733 = pi64  & n5732;
  assign n5734 = ~pi40  & pi41 ;
  assign n5735 = pi40  & ~pi41 ;
  assign n5736 = ~n5734 & ~n5735;
  assign n5737 = ~n5441 & n5736;
  assign n5738 = pi65  & n5737;
  assign n5739 = ~n5441 & ~n5736;
  assign n5740 = ~n265 & n5739;
  assign n5741 = ~n5733 & ~n5738;
  assign n5742 = ~n5740 & n5741;
  assign n5743 = pi41  & ~n5742;
  assign n5744 = pi41  & ~n5743;
  assign n5745 = ~n5742 & ~n5743;
  assign n5746 = ~n5744 & ~n5745;
  assign n5747 = n5728 & ~n5746;
  assign n5748 = ~n5728 & n5746;
  assign n5749 = ~n5747 & ~n5748;
  assign n5750 = n5727 & ~n5749;
  assign n5751 = ~n5727 & n5749;
  assign n5752 = ~n5750 & ~n5751;
  assign n5753 = ~n5716 & n5752;
  assign n5754 = n5716 & ~n5752;
  assign n5755 = ~n5753 & ~n5754;
  assign n5756 = n475 & n4271;
  assign n5757 = pi69  & n4503;
  assign n5758 = pi71  & n4269;
  assign n5759 = pi70  & n4264;
  assign n5760 = ~n5758 & ~n5759;
  assign n5761 = ~n5757 & n5760;
  assign n5762 = ~n5756 & n5761;
  assign n5763 = pi35  & ~n5762;
  assign n5764 = pi35  & ~n5763;
  assign n5765 = ~n5762 & ~n5763;
  assign n5766 = ~n5764 & ~n5765;
  assign n5767 = n5755 & ~n5766;
  assign n5768 = n5755 & ~n5767;
  assign n5769 = ~n5766 & ~n5767;
  assign n5770 = ~n5768 & ~n5769;
  assign n5771 = ~n5471 & ~n5478;
  assign n5772 = n5770 & n5771;
  assign n5773 = ~n5770 & ~n5771;
  assign n5774 = ~n5772 & ~n5773;
  assign n5775 = n729 & n3622;
  assign n5776 = pi72  & n3814;
  assign n5777 = pi74  & n3620;
  assign n5778 = pi73  & n3615;
  assign n5779 = ~n5777 & ~n5778;
  assign n5780 = ~n5776 & n5779;
  assign n5781 = ~n5775 & n5780;
  assign n5782 = pi32  & ~n5781;
  assign n5783 = pi32  & ~n5782;
  assign n5784 = ~n5781 & ~n5782;
  assign n5785 = ~n5783 & ~n5784;
  assign n5786 = n5774 & ~n5785;
  assign n5787 = ~n5774 & n5785;
  assign n5788 = ~n5786 & ~n5787;
  assign n5789 = ~n5714 & n5788;
  assign n5790 = ~n5714 & ~n5789;
  assign n5791 = ~n5786 & ~n5789;
  assign n5792 = ~n5787 & n5791;
  assign n5793 = ~n5790 & ~n5792;
  assign n5794 = n999 & n3034;
  assign n5795 = pi75  & n3225;
  assign n5796 = pi77  & n3032;
  assign n5797 = pi76  & n3027;
  assign n5798 = ~n5796 & ~n5797;
  assign n5799 = ~n5795 & n5798;
  assign n5800 = ~n5794 & n5799;
  assign n5801 = pi29  & ~n5800;
  assign n5802 = pi29  & ~n5801;
  assign n5803 = ~n5800 & ~n5801;
  assign n5804 = ~n5802 & ~n5803;
  assign n5805 = n5793 & n5804;
  assign n5806 = ~n5793 & ~n5804;
  assign n5807 = ~n5805 & ~n5806;
  assign n5808 = ~n5713 & n5807;
  assign n5809 = n5713 & ~n5807;
  assign n5810 = ~n5808 & ~n5809;
  assign n5811 = n1225 & n2523;
  assign n5812 = pi78  & n2667;
  assign n5813 = pi80  & n2521;
  assign n5814 = pi79  & n2516;
  assign n5815 = ~n5813 & ~n5814;
  assign n5816 = ~n5812 & n5815;
  assign n5817 = ~n5811 & n5816;
  assign n5818 = pi26  & ~n5817;
  assign n5819 = pi26  & ~n5818;
  assign n5820 = ~n5817 & ~n5818;
  assign n5821 = ~n5819 & ~n5820;
  assign n5822 = n5810 & ~n5821;
  assign n5823 = n5810 & ~n5822;
  assign n5824 = ~n5821 & ~n5822;
  assign n5825 = ~n5823 & ~n5824;
  assign n5826 = ~n5438 & ~n5531;
  assign n5827 = ~n5528 & ~n5826;
  assign n5828 = n5825 & n5827;
  assign n5829 = ~n5825 & ~n5827;
  assign n5830 = ~n5828 & ~n5829;
  assign n5831 = n1696 & n2043;
  assign n5832 = pi81  & n2180;
  assign n5833 = pi83  & n2041;
  assign n5834 = pi82  & n2036;
  assign n5835 = ~n5833 & ~n5834;
  assign n5836 = ~n5832 & n5835;
  assign n5837 = ~n5831 & n5836;
  assign n5838 = pi23  & ~n5837;
  assign n5839 = pi23  & ~n5838;
  assign n5840 = ~n5837 & ~n5838;
  assign n5841 = ~n5839 & ~n5840;
  assign n5842 = n5830 & ~n5841;
  assign n5843 = n5830 & ~n5842;
  assign n5844 = ~n5841 & ~n5842;
  assign n5845 = ~n5843 & ~n5844;
  assign n5846 = ~n5546 & ~n5550;
  assign n5847 = n5845 & n5846;
  assign n5848 = ~n5845 & ~n5846;
  assign n5849 = ~n5847 & ~n5848;
  assign n5850 = n1611 & n2133;
  assign n5851 = pi84  & n1745;
  assign n5852 = pi86  & n1609;
  assign n5853 = pi85  & n1604;
  assign n5854 = ~n5852 & ~n5853;
  assign n5855 = ~n5851 & n5854;
  assign n5856 = ~n5850 & n5855;
  assign n5857 = pi20  & ~n5856;
  assign n5858 = pi20  & ~n5857;
  assign n5859 = ~n5856 & ~n5857;
  assign n5860 = ~n5858 & ~n5859;
  assign n5861 = n5849 & ~n5860;
  assign n5862 = n5849 & ~n5861;
  assign n5863 = ~n5860 & ~n5861;
  assign n5864 = ~n5862 & ~n5863;
  assign n5865 = ~n5563 & ~n5569;
  assign n5866 = n5864 & n5865;
  assign n5867 = ~n5864 & ~n5865;
  assign n5868 = ~n5866 & ~n5867;
  assign n5869 = n1297 & n2473;
  assign n5870 = pi87  & n1366;
  assign n5871 = pi89  & n1295;
  assign n5872 = pi88  & n1290;
  assign n5873 = ~n5871 & ~n5872;
  assign n5874 = ~n5870 & n5873;
  assign n5875 = ~n5869 & n5874;
  assign n5876 = pi17  & ~n5875;
  assign n5877 = pi17  & ~n5876;
  assign n5878 = ~n5875 & ~n5876;
  assign n5879 = ~n5877 & ~n5878;
  assign n5880 = n5868 & ~n5879;
  assign n5881 = n5868 & ~n5880;
  assign n5882 = ~n5879 & ~n5880;
  assign n5883 = ~n5881 & ~n5882;
  assign n5884 = ~n5583 & ~n5585;
  assign n5885 = ~n5883 & ~n5884;
  assign n5886 = n5883 & n5884;
  assign n5887 = ~n5885 & ~n5886;
  assign n5888 = ~n5712 & n5887;
  assign n5889 = ~n5712 & ~n5888;
  assign n5890 = n5887 & ~n5888;
  assign n5891 = ~n5889 & ~n5890;
  assign n5892 = ~n5701 & ~n5891;
  assign n5893 = ~n5701 & ~n5892;
  assign n5894 = ~n5891 & ~n5892;
  assign n5895 = ~n5893 & ~n5894;
  assign n5896 = n687 & n3784;
  assign n5897 = pi93  & n763;
  assign n5898 = pi95  & n685;
  assign n5899 = pi94  & n680;
  assign n5900 = ~n5898 & ~n5899;
  assign n5901 = ~n5897 & n5900;
  assign n5902 = ~n5896 & n5901;
  assign n5903 = pi11  & ~n5902;
  assign n5904 = pi11  & ~n5903;
  assign n5905 = ~n5902 & ~n5903;
  assign n5906 = ~n5904 & ~n5905;
  assign n5907 = n5895 & n5906;
  assign n5908 = ~n5895 & ~n5906;
  assign n5909 = ~n5907 & ~n5908;
  assign n5910 = ~n5699 & n5909;
  assign n5911 = n5699 & ~n5909;
  assign n5912 = ~n5910 & ~n5911;
  assign n5913 = n5698 & ~n5912;
  assign n5914 = ~n5698 & n5912;
  assign n5915 = ~n5913 & ~n5914;
  assign n5916 = ~n5687 & n5915;
  assign n5917 = n5687 & ~n5915;
  assign n5918 = ~n5916 & ~n5917;
  assign n5919 = n342 & n5169;
  assign n5920 = pi99  & n380;
  assign n5921 = pi101  & n340;
  assign n5922 = pi100  & n335;
  assign n5923 = ~n5921 & ~n5922;
  assign n5924 = ~n5920 & n5923;
  assign n5925 = ~n5919 & n5924;
  assign n5926 = pi5  & ~n5925;
  assign n5927 = pi5  & ~n5926;
  assign n5928 = ~n5925 & ~n5926;
  assign n5929 = ~n5927 & ~n5928;
  assign n5930 = n5918 & ~n5929;
  assign n5931 = n5918 & ~n5930;
  assign n5932 = ~n5929 & ~n5930;
  assign n5933 = ~n5931 & ~n5932;
  assign n5934 = ~n5685 & n5933;
  assign n5935 = n5685 & ~n5933;
  assign n5936 = ~n5934 & ~n5935;
  assign n5937 = ~n5660 & ~n5662;
  assign n5938 = ~pi103  & ~pi104 ;
  assign n5939 = pi103  & pi104 ;
  assign n5940 = ~n5938 & ~n5939;
  assign n5941 = ~n5937 & n5940;
  assign n5942 = n5937 & ~n5940;
  assign n5943 = ~n5941 & ~n5942;
  assign n5944 = n262 & n5943;
  assign n5945 = pi102  & n288;
  assign n5946 = pi104  & n267;
  assign n5947 = pi103  & n269;
  assign n5948 = ~n5946 & ~n5947;
  assign n5949 = ~n5945 & n5948;
  assign n5950 = ~n5944 & n5949;
  assign n5951 = pi2  & ~n5950;
  assign n5952 = pi2  & ~n5951;
  assign n5953 = ~n5950 & ~n5951;
  assign n5954 = ~n5952 & ~n5953;
  assign n5955 = ~n5936 & ~n5954;
  assign n5956 = n5936 & n5954;
  assign n5957 = ~n5955 & ~n5956;
  assign n5958 = ~n5684 & n5957;
  assign n5959 = n5684 & ~n5957;
  assign po40  = ~n5958 & ~n5959;
  assign n5961 = ~n5955 & ~n5958;
  assign n5962 = ~n5685 & ~n5933;
  assign n5963 = ~n5930 & ~n5962;
  assign n5964 = ~n5914 & ~n5916;
  assign n5965 = ~n5908 & ~n5910;
  assign n5966 = n687 & n4001;
  assign n5967 = pi94  & n763;
  assign n5968 = pi96  & n685;
  assign n5969 = pi95  & n680;
  assign n5970 = ~n5968 & ~n5969;
  assign n5971 = ~n5967 & n5970;
  assign n5972 = ~n5966 & n5971;
  assign n5973 = pi11  & ~n5972;
  assign n5974 = pi11  & ~n5973;
  assign n5975 = ~n5972 & ~n5973;
  assign n5976 = ~n5974 & ~n5975;
  assign n5977 = ~n5888 & ~n5892;
  assign n5978 = n938 & n3371;
  assign n5979 = pi91  & n1052;
  assign n5980 = pi93  & n936;
  assign n5981 = pi92  & n931;
  assign n5982 = ~n5980 & ~n5981;
  assign n5983 = ~n5979 & n5982;
  assign n5984 = ~n5978 & n5983;
  assign n5985 = pi14  & ~n5984;
  assign n5986 = pi14  & ~n5985;
  assign n5987 = ~n5984 & ~n5985;
  assign n5988 = ~n5986 & ~n5987;
  assign n5989 = ~n5880 & ~n5885;
  assign n5990 = ~n5861 & ~n5867;
  assign n5991 = ~n5822 & ~n5829;
  assign n5992 = n1434 & n2523;
  assign n5993 = pi79  & n2667;
  assign n5994 = pi81  & n2521;
  assign n5995 = pi80  & n2516;
  assign n5996 = ~n5994 & ~n5995;
  assign n5997 = ~n5993 & n5996;
  assign n5998 = ~n5992 & n5997;
  assign n5999 = pi26  & ~n5998;
  assign n6000 = pi26  & ~n5999;
  assign n6001 = ~n5998 & ~n5999;
  assign n6002 = ~n6000 & ~n6001;
  assign n6003 = ~n5806 & ~n5808;
  assign n6004 = n1025 & n3034;
  assign n6005 = pi76  & n3225;
  assign n6006 = pi78  & n3032;
  assign n6007 = pi77  & n3027;
  assign n6008 = ~n6006 & ~n6007;
  assign n6009 = ~n6005 & n6008;
  assign n6010 = ~n6004 & n6009;
  assign n6011 = pi29  & ~n6010;
  assign n6012 = pi29  & ~n6011;
  assign n6013 = ~n6010 & ~n6011;
  assign n6014 = ~n6012 & ~n6013;
  assign n6015 = ~n5767 & ~n5773;
  assign n6016 = n576 & n4271;
  assign n6017 = pi70  & n4503;
  assign n6018 = pi72  & n4269;
  assign n6019 = pi71  & n4264;
  assign n6020 = ~n6018 & ~n6019;
  assign n6021 = ~n6017 & n6020;
  assign n6022 = ~n6016 & n6021;
  assign n6023 = pi35  & ~n6022;
  assign n6024 = pi35  & ~n6023;
  assign n6025 = ~n6022 & ~n6023;
  assign n6026 = ~n6024 & ~n6025;
  assign n6027 = ~n5751 & ~n5753;
  assign n6028 = n286 & n5739;
  assign n6029 = n5441 & n5731;
  assign n6030 = ~n5736 & n6029;
  assign n6031 = pi64  & n6030;
  assign n6032 = pi66  & n5737;
  assign n6033 = pi65  & n5732;
  assign n6034 = ~n6032 & ~n6033;
  assign n6035 = ~n6028 & n6034;
  assign n6036 = ~n6031 & n6035;
  assign n6037 = pi41  & ~n6036;
  assign n6038 = pi41  & ~n6037;
  assign n6039 = ~n6036 & ~n6037;
  assign n6040 = ~n6038 & ~n6039;
  assign n6041 = ~n5747 & n6040;
  assign n6042 = n5747 & ~n6040;
  assign n6043 = ~n6041 & ~n6042;
  assign n6044 = n401 & n5008;
  assign n6045 = pi67  & n5241;
  assign n6046 = pi69  & n5006;
  assign n6047 = pi68  & n5001;
  assign n6048 = ~n6046 & ~n6047;
  assign n6049 = ~n6045 & n6048;
  assign n6050 = ~n6044 & n6049;
  assign n6051 = pi38  & ~n6050;
  assign n6052 = pi38  & ~n6051;
  assign n6053 = ~n6050 & ~n6051;
  assign n6054 = ~n6052 & ~n6053;
  assign n6055 = n6043 & ~n6054;
  assign n6056 = n6043 & ~n6055;
  assign n6057 = ~n6054 & ~n6055;
  assign n6058 = ~n6056 & ~n6057;
  assign n6059 = ~n6027 & ~n6058;
  assign n6060 = n6027 & n6058;
  assign n6061 = ~n6059 & ~n6060;
  assign n6062 = ~n6026 & n6061;
  assign n6063 = ~n6026 & ~n6062;
  assign n6064 = n6061 & ~n6062;
  assign n6065 = ~n6063 & ~n6064;
  assign n6066 = ~n6015 & ~n6065;
  assign n6067 = ~n6015 & ~n6066;
  assign n6068 = ~n6065 & ~n6066;
  assign n6069 = ~n6067 & ~n6068;
  assign n6070 = n809 & n3622;
  assign n6071 = pi73  & n3814;
  assign n6072 = pi75  & n3620;
  assign n6073 = pi74  & n3615;
  assign n6074 = ~n6072 & ~n6073;
  assign n6075 = ~n6071 & n6074;
  assign n6076 = ~n6070 & n6075;
  assign n6077 = pi32  & ~n6076;
  assign n6078 = pi32  & ~n6077;
  assign n6079 = ~n6076 & ~n6077;
  assign n6080 = ~n6078 & ~n6079;
  assign n6081 = n6069 & n6080;
  assign n6082 = ~n6069 & ~n6080;
  assign n6083 = ~n6081 & ~n6082;
  assign n6084 = ~n5791 & n6083;
  assign n6085 = n5791 & ~n6083;
  assign n6086 = ~n6084 & ~n6085;
  assign n6087 = n6014 & ~n6086;
  assign n6088 = ~n6014 & n6086;
  assign n6089 = ~n6087 & ~n6088;
  assign n6090 = ~n6003 & n6089;
  assign n6091 = n6003 & ~n6089;
  assign n6092 = ~n6090 & ~n6091;
  assign n6093 = n6002 & ~n6092;
  assign n6094 = ~n6002 & n6092;
  assign n6095 = ~n6093 & ~n6094;
  assign n6096 = ~n5991 & n6095;
  assign n6097 = n5991 & ~n6095;
  assign n6098 = ~n6096 & ~n6097;
  assign n6099 = n1834 & n2043;
  assign n6100 = pi82  & n2180;
  assign n6101 = pi84  & n2041;
  assign n6102 = pi83  & n2036;
  assign n6103 = ~n6101 & ~n6102;
  assign n6104 = ~n6100 & n6103;
  assign n6105 = ~n6099 & n6104;
  assign n6106 = pi23  & ~n6105;
  assign n6107 = pi23  & ~n6106;
  assign n6108 = ~n6105 & ~n6106;
  assign n6109 = ~n6107 & ~n6108;
  assign n6110 = n6098 & ~n6109;
  assign n6111 = n6098 & ~n6110;
  assign n6112 = ~n6109 & ~n6110;
  assign n6113 = ~n6111 & ~n6112;
  assign n6114 = ~n5842 & ~n5848;
  assign n6115 = n6113 & n6114;
  assign n6116 = ~n6113 & ~n6114;
  assign n6117 = ~n6115 & ~n6116;
  assign n6118 = n1611 & n2288;
  assign n6119 = pi85  & n1745;
  assign n6120 = pi87  & n1609;
  assign n6121 = pi86  & n1604;
  assign n6122 = ~n6120 & ~n6121;
  assign n6123 = ~n6119 & n6122;
  assign n6124 = ~n6118 & n6123;
  assign n6125 = pi20  & ~n6124;
  assign n6126 = pi20  & ~n6125;
  assign n6127 = ~n6124 & ~n6125;
  assign n6128 = ~n6126 & ~n6127;
  assign n6129 = n6117 & ~n6128;
  assign n6130 = ~n6117 & n6128;
  assign n6131 = ~n6129 & ~n6130;
  assign n6132 = ~n5990 & n6131;
  assign n6133 = ~n5990 & ~n6132;
  assign n6134 = ~n6129 & ~n6132;
  assign n6135 = ~n6130 & n6134;
  assign n6136 = ~n6133 & ~n6135;
  assign n6137 = n1297 & n2801;
  assign n6138 = pi88  & n1366;
  assign n6139 = pi90  & n1295;
  assign n6140 = pi89  & n1290;
  assign n6141 = ~n6139 & ~n6140;
  assign n6142 = ~n6138 & n6141;
  assign n6143 = ~n6137 & n6142;
  assign n6144 = pi17  & ~n6143;
  assign n6145 = pi17  & ~n6144;
  assign n6146 = ~n6143 & ~n6144;
  assign n6147 = ~n6145 & ~n6146;
  assign n6148 = n6136 & n6147;
  assign n6149 = ~n6136 & ~n6147;
  assign n6150 = ~n6148 & ~n6149;
  assign n6151 = ~n5989 & n6150;
  assign n6152 = n5989 & ~n6150;
  assign n6153 = ~n6151 & ~n6152;
  assign n6154 = n5988 & ~n6153;
  assign n6155 = ~n5988 & n6153;
  assign n6156 = ~n6154 & ~n6155;
  assign n6157 = ~n5977 & n6156;
  assign n6158 = n5977 & ~n6156;
  assign n6159 = ~n6157 & ~n6158;
  assign n6160 = n5976 & ~n6159;
  assign n6161 = ~n5976 & n6159;
  assign n6162 = ~n6160 & ~n6161;
  assign n6163 = ~n5965 & n6162;
  assign n6164 = n5965 & ~n6162;
  assign n6165 = ~n6163 & ~n6164;
  assign n6166 = n498 & n4684;
  assign n6167 = pi97  & n537;
  assign n6168 = pi99  & n496;
  assign n6169 = pi98  & n491;
  assign n6170 = ~n6168 & ~n6169;
  assign n6171 = ~n6167 & n6170;
  assign n6172 = ~n6166 & n6171;
  assign n6173 = pi8  & ~n6172;
  assign n6174 = pi8  & ~n6173;
  assign n6175 = ~n6172 & ~n6173;
  assign n6176 = ~n6174 & ~n6175;
  assign n6177 = n6165 & ~n6176;
  assign n6178 = n6165 & ~n6177;
  assign n6179 = ~n6176 & ~n6177;
  assign n6180 = ~n6178 & ~n6179;
  assign n6181 = ~n5964 & n6180;
  assign n6182 = n5964 & ~n6180;
  assign n6183 = ~n6181 & ~n6182;
  assign n6184 = n342 & n5413;
  assign n6185 = pi100  & n380;
  assign n6186 = pi102  & n340;
  assign n6187 = pi101  & n335;
  assign n6188 = ~n6186 & ~n6187;
  assign n6189 = ~n6185 & n6188;
  assign n6190 = ~n6184 & n6189;
  assign n6191 = pi5  & ~n6190;
  assign n6192 = pi5  & ~n6191;
  assign n6193 = ~n6190 & ~n6191;
  assign n6194 = ~n6192 & ~n6193;
  assign n6195 = ~n6183 & ~n6194;
  assign n6196 = n6183 & n6194;
  assign n6197 = ~n6195 & ~n6196;
  assign n6198 = n5963 & ~n6197;
  assign n6199 = ~n5963 & n6197;
  assign n6200 = ~n6198 & ~n6199;
  assign n6201 = ~n5939 & ~n5941;
  assign n6202 = ~pi104  & ~pi105 ;
  assign n6203 = pi104  & pi105 ;
  assign n6204 = ~n6202 & ~n6203;
  assign n6205 = ~n6201 & n6204;
  assign n6206 = n6201 & ~n6204;
  assign n6207 = ~n6205 & ~n6206;
  assign n6208 = n262 & n6207;
  assign n6209 = pi103  & n288;
  assign n6210 = pi105  & n267;
  assign n6211 = pi104  & n269;
  assign n6212 = ~n6210 & ~n6211;
  assign n6213 = ~n6209 & n6212;
  assign n6214 = ~n6208 & n6213;
  assign n6215 = pi2  & ~n6214;
  assign n6216 = pi2  & ~n6215;
  assign n6217 = ~n6214 & ~n6215;
  assign n6218 = ~n6216 & ~n6217;
  assign n6219 = ~n6200 & n6218;
  assign n6220 = n6200 & ~n6218;
  assign n6221 = ~n6219 & ~n6220;
  assign n6222 = ~n5961 & n6221;
  assign n6223 = n5961 & ~n6221;
  assign po41  = ~n6222 & ~n6223;
  assign n6225 = ~n6195 & ~n6199;
  assign n6226 = n342 & n5664;
  assign n6227 = pi101  & n380;
  assign n6228 = pi103  & n340;
  assign n6229 = pi102  & n335;
  assign n6230 = ~n6228 & ~n6229;
  assign n6231 = ~n6227 & n6230;
  assign n6232 = ~n6226 & n6231;
  assign n6233 = pi5  & ~n6232;
  assign n6234 = pi5  & ~n6233;
  assign n6235 = ~n6232 & ~n6233;
  assign n6236 = ~n6234 & ~n6235;
  assign n6237 = ~n5964 & ~n6180;
  assign n6238 = ~n6177 & ~n6237;
  assign n6239 = ~n6161 & ~n6163;
  assign n6240 = ~n6155 & ~n6157;
  assign n6241 = ~n6149 & ~n6151;
  assign n6242 = ~n6094 & ~n6096;
  assign n6243 = ~n6088 & ~n6090;
  assign n6244 = ~n6082 & ~n6084;
  assign n6245 = n891 & n3622;
  assign n6246 = pi74  & n3814;
  assign n6247 = pi76  & n3620;
  assign n6248 = pi75  & n3615;
  assign n6249 = ~n6247 & ~n6248;
  assign n6250 = ~n6246 & n6249;
  assign n6251 = ~n6245 & n6250;
  assign n6252 = pi32  & ~n6251;
  assign n6253 = pi32  & ~n6252;
  assign n6254 = ~n6251 & ~n6252;
  assign n6255 = ~n6253 & ~n6254;
  assign n6256 = ~n6062 & ~n6066;
  assign n6257 = pi41  & ~pi42 ;
  assign n6258 = ~pi41  & pi42 ;
  assign n6259 = ~n6257 & ~n6258;
  assign n6260 = pi64  & ~n6259;
  assign n6261 = ~n6042 & n6260;
  assign n6262 = n6042 & ~n6260;
  assign n6263 = ~n6261 & ~n6262;
  assign n6264 = n309 & n5739;
  assign n6265 = pi65  & n6030;
  assign n6266 = pi67  & n5737;
  assign n6267 = pi66  & n5732;
  assign n6268 = ~n6266 & ~n6267;
  assign n6269 = ~n6265 & n6268;
  assign n6270 = ~n6264 & n6269;
  assign n6271 = pi41  & ~n6270;
  assign n6272 = pi41  & ~n6271;
  assign n6273 = ~n6270 & ~n6271;
  assign n6274 = ~n6272 & ~n6273;
  assign n6275 = ~n6263 & ~n6274;
  assign n6276 = n6263 & n6274;
  assign n6277 = ~n6275 & ~n6276;
  assign n6278 = n450 & n5008;
  assign n6279 = pi68  & n5241;
  assign n6280 = pi70  & n5006;
  assign n6281 = pi69  & n5001;
  assign n6282 = ~n6280 & ~n6281;
  assign n6283 = ~n6279 & n6282;
  assign n6284 = ~n6278 & n6283;
  assign n6285 = pi38  & ~n6284;
  assign n6286 = pi38  & ~n6285;
  assign n6287 = ~n6284 & ~n6285;
  assign n6288 = ~n6286 & ~n6287;
  assign n6289 = n6277 & ~n6288;
  assign n6290 = n6277 & ~n6289;
  assign n6291 = ~n6288 & ~n6289;
  assign n6292 = ~n6290 & ~n6291;
  assign n6293 = ~n6055 & ~n6059;
  assign n6294 = n6292 & n6293;
  assign n6295 = ~n6292 & ~n6293;
  assign n6296 = ~n6294 & ~n6295;
  assign n6297 = n642 & n4271;
  assign n6298 = pi71  & n4503;
  assign n6299 = pi73  & n4269;
  assign n6300 = pi72  & n4264;
  assign n6301 = ~n6299 & ~n6300;
  assign n6302 = ~n6298 & n6301;
  assign n6303 = ~n6297 & n6302;
  assign n6304 = pi35  & ~n6303;
  assign n6305 = pi35  & ~n6304;
  assign n6306 = ~n6303 & ~n6304;
  assign n6307 = ~n6305 & ~n6306;
  assign n6308 = ~n6296 & n6307;
  assign n6309 = n6296 & ~n6307;
  assign n6310 = ~n6308 & ~n6309;
  assign n6311 = ~n6256 & n6310;
  assign n6312 = n6256 & ~n6310;
  assign n6313 = ~n6311 & ~n6312;
  assign n6314 = ~n6255 & n6313;
  assign n6315 = ~n6255 & ~n6314;
  assign n6316 = n6313 & ~n6314;
  assign n6317 = ~n6315 & ~n6316;
  assign n6318 = ~n6244 & ~n6317;
  assign n6319 = ~n6244 & ~n6318;
  assign n6320 = ~n6317 & ~n6318;
  assign n6321 = ~n6319 & ~n6320;
  assign n6322 = n1122 & n3034;
  assign n6323 = pi77  & n3225;
  assign n6324 = pi79  & n3032;
  assign n6325 = pi78  & n3027;
  assign n6326 = ~n6324 & ~n6325;
  assign n6327 = ~n6323 & n6326;
  assign n6328 = ~n6322 & n6327;
  assign n6329 = pi29  & ~n6328;
  assign n6330 = pi29  & ~n6329;
  assign n6331 = ~n6328 & ~n6329;
  assign n6332 = ~n6330 & ~n6331;
  assign n6333 = ~n6321 & ~n6332;
  assign n6334 = ~n6321 & ~n6333;
  assign n6335 = ~n6332 & ~n6333;
  assign n6336 = ~n6334 & ~n6335;
  assign n6337 = ~n6243 & n6336;
  assign n6338 = n6243 & ~n6336;
  assign n6339 = ~n6337 & ~n6338;
  assign n6340 = n1554 & n2523;
  assign n6341 = pi80  & n2667;
  assign n6342 = pi82  & n2521;
  assign n6343 = pi81  & n2516;
  assign n6344 = ~n6342 & ~n6343;
  assign n6345 = ~n6341 & n6344;
  assign n6346 = ~n6340 & n6345;
  assign n6347 = pi26  & ~n6346;
  assign n6348 = pi26  & ~n6347;
  assign n6349 = ~n6346 & ~n6347;
  assign n6350 = ~n6348 & ~n6349;
  assign n6351 = ~n6339 & ~n6350;
  assign n6352 = n6339 & n6350;
  assign n6353 = ~n6351 & ~n6352;
  assign n6354 = ~n6242 & n6353;
  assign n6355 = n6242 & ~n6353;
  assign n6356 = ~n6354 & ~n6355;
  assign n6357 = n1972 & n2043;
  assign n6358 = pi83  & n2180;
  assign n6359 = pi85  & n2041;
  assign n6360 = pi84  & n2036;
  assign n6361 = ~n6359 & ~n6360;
  assign n6362 = ~n6358 & n6361;
  assign n6363 = ~n6357 & n6362;
  assign n6364 = pi23  & ~n6363;
  assign n6365 = pi23  & ~n6364;
  assign n6366 = ~n6363 & ~n6364;
  assign n6367 = ~n6365 & ~n6366;
  assign n6368 = n6356 & ~n6367;
  assign n6369 = n6356 & ~n6368;
  assign n6370 = ~n6367 & ~n6368;
  assign n6371 = ~n6369 & ~n6370;
  assign n6372 = ~n6110 & ~n6116;
  assign n6373 = n6371 & n6372;
  assign n6374 = ~n6371 & ~n6372;
  assign n6375 = ~n6373 & ~n6374;
  assign n6376 = n1611 & n2446;
  assign n6377 = pi86  & n1745;
  assign n6378 = pi88  & n1609;
  assign n6379 = pi87  & n1604;
  assign n6380 = ~n6378 & ~n6379;
  assign n6381 = ~n6377 & n6380;
  assign n6382 = ~n6376 & n6381;
  assign n6383 = pi20  & ~n6382;
  assign n6384 = pi20  & ~n6383;
  assign n6385 = ~n6382 & ~n6383;
  assign n6386 = ~n6384 & ~n6385;
  assign n6387 = ~n6375 & n6386;
  assign n6388 = n6375 & ~n6386;
  assign n6389 = ~n6387 & ~n6388;
  assign n6390 = ~n6134 & n6389;
  assign n6391 = n6134 & ~n6389;
  assign n6392 = ~n6390 & ~n6391;
  assign n6393 = n1297 & n2978;
  assign n6394 = pi89  & n1366;
  assign n6395 = pi91  & n1295;
  assign n6396 = pi90  & n1290;
  assign n6397 = ~n6395 & ~n6396;
  assign n6398 = ~n6394 & n6397;
  assign n6399 = ~n6393 & n6398;
  assign n6400 = pi17  & ~n6399;
  assign n6401 = pi17  & ~n6400;
  assign n6402 = ~n6399 & ~n6400;
  assign n6403 = ~n6401 & ~n6402;
  assign n6404 = n6392 & ~n6403;
  assign n6405 = n6392 & ~n6404;
  assign n6406 = ~n6403 & ~n6404;
  assign n6407 = ~n6405 & ~n6406;
  assign n6408 = ~n6241 & n6407;
  assign n6409 = n6241 & ~n6407;
  assign n6410 = ~n6408 & ~n6409;
  assign n6411 = n938 & n3565;
  assign n6412 = pi92  & n1052;
  assign n6413 = pi94  & n936;
  assign n6414 = pi93  & n931;
  assign n6415 = ~n6413 & ~n6414;
  assign n6416 = ~n6412 & n6415;
  assign n6417 = ~n6411 & n6416;
  assign n6418 = pi14  & ~n6417;
  assign n6419 = pi14  & ~n6418;
  assign n6420 = ~n6417 & ~n6418;
  assign n6421 = ~n6419 & ~n6420;
  assign n6422 = ~n6410 & ~n6421;
  assign n6423 = n6410 & n6421;
  assign n6424 = ~n6422 & ~n6423;
  assign n6425 = ~n6240 & n6424;
  assign n6426 = n6240 & ~n6424;
  assign n6427 = ~n6425 & ~n6426;
  assign n6428 = n687 & n4211;
  assign n6429 = pi95  & n763;
  assign n6430 = pi97  & n685;
  assign n6431 = pi96  & n680;
  assign n6432 = ~n6430 & ~n6431;
  assign n6433 = ~n6429 & n6432;
  assign n6434 = ~n6428 & n6433;
  assign n6435 = pi11  & ~n6434;
  assign n6436 = pi11  & ~n6435;
  assign n6437 = ~n6434 & ~n6435;
  assign n6438 = ~n6436 & ~n6437;
  assign n6439 = n6427 & ~n6438;
  assign n6440 = n6427 & ~n6439;
  assign n6441 = ~n6438 & ~n6439;
  assign n6442 = ~n6440 & ~n6441;
  assign n6443 = ~n6239 & n6442;
  assign n6444 = n6239 & ~n6442;
  assign n6445 = ~n6443 & ~n6444;
  assign n6446 = n498 & n4910;
  assign n6447 = pi98  & n537;
  assign n6448 = pi100  & n496;
  assign n6449 = pi99  & n491;
  assign n6450 = ~n6448 & ~n6449;
  assign n6451 = ~n6447 & n6450;
  assign n6452 = ~n6446 & n6451;
  assign n6453 = pi8  & ~n6452;
  assign n6454 = pi8  & ~n6453;
  assign n6455 = ~n6452 & ~n6453;
  assign n6456 = ~n6454 & ~n6455;
  assign n6457 = n6445 & n6456;
  assign n6458 = ~n6445 & ~n6456;
  assign n6459 = ~n6457 & ~n6458;
  assign n6460 = ~n6238 & n6459;
  assign n6461 = n6238 & ~n6459;
  assign n6462 = ~n6460 & ~n6461;
  assign n6463 = ~n6236 & n6462;
  assign n6464 = ~n6236 & ~n6463;
  assign n6465 = n6462 & ~n6463;
  assign n6466 = ~n6464 & ~n6465;
  assign n6467 = ~n6225 & ~n6466;
  assign n6468 = ~n6225 & ~n6467;
  assign n6469 = ~n6466 & ~n6467;
  assign n6470 = ~n6468 & ~n6469;
  assign n6471 = ~n6203 & ~n6205;
  assign n6472 = ~pi105  & ~pi106 ;
  assign n6473 = pi105  & pi106 ;
  assign n6474 = ~n6472 & ~n6473;
  assign n6475 = ~n6471 & n6474;
  assign n6476 = n6471 & ~n6474;
  assign n6477 = ~n6475 & ~n6476;
  assign n6478 = n262 & n6477;
  assign n6479 = pi104  & n288;
  assign n6480 = pi106  & n267;
  assign n6481 = pi105  & n269;
  assign n6482 = ~n6480 & ~n6481;
  assign n6483 = ~n6479 & n6482;
  assign n6484 = ~n6478 & n6483;
  assign n6485 = pi2  & ~n6484;
  assign n6486 = pi2  & ~n6485;
  assign n6487 = ~n6484 & ~n6485;
  assign n6488 = ~n6486 & ~n6487;
  assign n6489 = ~n6470 & ~n6488;
  assign n6490 = ~n6470 & ~n6489;
  assign n6491 = ~n6488 & ~n6489;
  assign n6492 = ~n6490 & ~n6491;
  assign n6493 = ~n6220 & ~n6222;
  assign n6494 = ~n6492 & ~n6493;
  assign n6495 = n6492 & n6493;
  assign po42  = ~n6494 & ~n6495;
  assign n6497 = ~n6463 & ~n6467;
  assign n6498 = ~n6458 & ~n6460;
  assign n6499 = ~n6422 & ~n6425;
  assign n6500 = ~n6241 & ~n6407;
  assign n6501 = ~n6404 & ~n6500;
  assign n6502 = n1297 & n3177;
  assign n6503 = pi90  & n1366;
  assign n6504 = pi92  & n1295;
  assign n6505 = pi91  & n1290;
  assign n6506 = ~n6504 & ~n6505;
  assign n6507 = ~n6503 & n6506;
  assign n6508 = ~n6502 & n6507;
  assign n6509 = pi17  & ~n6508;
  assign n6510 = pi17  & ~n6509;
  assign n6511 = ~n6508 & ~n6509;
  assign n6512 = ~n6510 & ~n6511;
  assign n6513 = ~n6314 & ~n6318;
  assign n6514 = ~n6309 & ~n6311;
  assign n6515 = n6042 & n6260;
  assign n6516 = ~n6275 & ~n6515;
  assign n6517 = n359 & n5739;
  assign n6518 = pi66  & n6030;
  assign n6519 = pi68  & n5737;
  assign n6520 = pi67  & n5732;
  assign n6521 = ~n6519 & ~n6520;
  assign n6522 = ~n6518 & n6521;
  assign n6523 = ~n6517 & n6522;
  assign n6524 = pi41  & ~n6523;
  assign n6525 = pi41  & ~n6524;
  assign n6526 = ~n6523 & ~n6524;
  assign n6527 = ~n6525 & ~n6526;
  assign n6528 = pi44  & ~n6260;
  assign n6529 = ~pi42  & pi43 ;
  assign n6530 = pi42  & ~pi43 ;
  assign n6531 = ~n6529 & ~n6530;
  assign n6532 = n6259 & ~n6531;
  assign n6533 = pi64  & n6532;
  assign n6534 = ~pi43  & pi44 ;
  assign n6535 = pi43  & ~pi44 ;
  assign n6536 = ~n6534 & ~n6535;
  assign n6537 = ~n6259 & n6536;
  assign n6538 = pi65  & n6537;
  assign n6539 = ~n6259 & ~n6536;
  assign n6540 = ~n265 & n6539;
  assign n6541 = ~n6533 & ~n6538;
  assign n6542 = ~n6540 & n6541;
  assign n6543 = pi44  & ~n6542;
  assign n6544 = pi44  & ~n6543;
  assign n6545 = ~n6542 & ~n6543;
  assign n6546 = ~n6544 & ~n6545;
  assign n6547 = n6528 & ~n6546;
  assign n6548 = ~n6528 & n6546;
  assign n6549 = ~n6547 & ~n6548;
  assign n6550 = n6527 & ~n6549;
  assign n6551 = ~n6527 & n6549;
  assign n6552 = ~n6550 & ~n6551;
  assign n6553 = ~n6516 & n6552;
  assign n6554 = n6516 & ~n6552;
  assign n6555 = ~n6553 & ~n6554;
  assign n6556 = n475 & n5008;
  assign n6557 = pi69  & n5241;
  assign n6558 = pi71  & n5006;
  assign n6559 = pi70  & n5001;
  assign n6560 = ~n6558 & ~n6559;
  assign n6561 = ~n6557 & n6560;
  assign n6562 = ~n6556 & n6561;
  assign n6563 = pi38  & ~n6562;
  assign n6564 = pi38  & ~n6563;
  assign n6565 = ~n6562 & ~n6563;
  assign n6566 = ~n6564 & ~n6565;
  assign n6567 = n6555 & ~n6566;
  assign n6568 = n6555 & ~n6567;
  assign n6569 = ~n6566 & ~n6567;
  assign n6570 = ~n6568 & ~n6569;
  assign n6571 = ~n6289 & ~n6295;
  assign n6572 = n6570 & n6571;
  assign n6573 = ~n6570 & ~n6571;
  assign n6574 = ~n6572 & ~n6573;
  assign n6575 = n729 & n4271;
  assign n6576 = pi72  & n4503;
  assign n6577 = pi74  & n4269;
  assign n6578 = pi73  & n4264;
  assign n6579 = ~n6577 & ~n6578;
  assign n6580 = ~n6576 & n6579;
  assign n6581 = ~n6575 & n6580;
  assign n6582 = pi35  & ~n6581;
  assign n6583 = pi35  & ~n6582;
  assign n6584 = ~n6581 & ~n6582;
  assign n6585 = ~n6583 & ~n6584;
  assign n6586 = n6574 & ~n6585;
  assign n6587 = ~n6574 & n6585;
  assign n6588 = ~n6586 & ~n6587;
  assign n6589 = ~n6514 & n6588;
  assign n6590 = ~n6514 & ~n6589;
  assign n6591 = ~n6586 & ~n6589;
  assign n6592 = ~n6587 & n6591;
  assign n6593 = ~n6590 & ~n6592;
  assign n6594 = n999 & n3622;
  assign n6595 = pi75  & n3814;
  assign n6596 = pi77  & n3620;
  assign n6597 = pi76  & n3615;
  assign n6598 = ~n6596 & ~n6597;
  assign n6599 = ~n6595 & n6598;
  assign n6600 = ~n6594 & n6599;
  assign n6601 = pi32  & ~n6600;
  assign n6602 = pi32  & ~n6601;
  assign n6603 = ~n6600 & ~n6601;
  assign n6604 = ~n6602 & ~n6603;
  assign n6605 = n6593 & n6604;
  assign n6606 = ~n6593 & ~n6604;
  assign n6607 = ~n6605 & ~n6606;
  assign n6608 = ~n6513 & n6607;
  assign n6609 = n6513 & ~n6607;
  assign n6610 = ~n6608 & ~n6609;
  assign n6611 = n1225 & n3034;
  assign n6612 = pi78  & n3225;
  assign n6613 = pi80  & n3032;
  assign n6614 = pi79  & n3027;
  assign n6615 = ~n6613 & ~n6614;
  assign n6616 = ~n6612 & n6615;
  assign n6617 = ~n6611 & n6616;
  assign n6618 = pi29  & ~n6617;
  assign n6619 = pi29  & ~n6618;
  assign n6620 = ~n6617 & ~n6618;
  assign n6621 = ~n6619 & ~n6620;
  assign n6622 = n6610 & ~n6621;
  assign n6623 = n6610 & ~n6622;
  assign n6624 = ~n6621 & ~n6622;
  assign n6625 = ~n6623 & ~n6624;
  assign n6626 = ~n6243 & ~n6336;
  assign n6627 = ~n6333 & ~n6626;
  assign n6628 = n6625 & n6627;
  assign n6629 = ~n6625 & ~n6627;
  assign n6630 = ~n6628 & ~n6629;
  assign n6631 = n1696 & n2523;
  assign n6632 = pi81  & n2667;
  assign n6633 = pi83  & n2521;
  assign n6634 = pi82  & n2516;
  assign n6635 = ~n6633 & ~n6634;
  assign n6636 = ~n6632 & n6635;
  assign n6637 = ~n6631 & n6636;
  assign n6638 = pi26  & ~n6637;
  assign n6639 = pi26  & ~n6638;
  assign n6640 = ~n6637 & ~n6638;
  assign n6641 = ~n6639 & ~n6640;
  assign n6642 = n6630 & ~n6641;
  assign n6643 = n6630 & ~n6642;
  assign n6644 = ~n6641 & ~n6642;
  assign n6645 = ~n6643 & ~n6644;
  assign n6646 = ~n6351 & ~n6354;
  assign n6647 = n6645 & n6646;
  assign n6648 = ~n6645 & ~n6646;
  assign n6649 = ~n6647 & ~n6648;
  assign n6650 = n2043 & n2133;
  assign n6651 = pi84  & n2180;
  assign n6652 = pi86  & n2041;
  assign n6653 = pi85  & n2036;
  assign n6654 = ~n6652 & ~n6653;
  assign n6655 = ~n6651 & n6654;
  assign n6656 = ~n6650 & n6655;
  assign n6657 = pi23  & ~n6656;
  assign n6658 = pi23  & ~n6657;
  assign n6659 = ~n6656 & ~n6657;
  assign n6660 = ~n6658 & ~n6659;
  assign n6661 = n6649 & ~n6660;
  assign n6662 = n6649 & ~n6661;
  assign n6663 = ~n6660 & ~n6661;
  assign n6664 = ~n6662 & ~n6663;
  assign n6665 = ~n6368 & ~n6374;
  assign n6666 = n6664 & n6665;
  assign n6667 = ~n6664 & ~n6665;
  assign n6668 = ~n6666 & ~n6667;
  assign n6669 = n1611 & n2473;
  assign n6670 = pi87  & n1745;
  assign n6671 = pi89  & n1609;
  assign n6672 = pi88  & n1604;
  assign n6673 = ~n6671 & ~n6672;
  assign n6674 = ~n6670 & n6673;
  assign n6675 = ~n6669 & n6674;
  assign n6676 = pi20  & ~n6675;
  assign n6677 = pi20  & ~n6676;
  assign n6678 = ~n6675 & ~n6676;
  assign n6679 = ~n6677 & ~n6678;
  assign n6680 = n6668 & ~n6679;
  assign n6681 = n6668 & ~n6680;
  assign n6682 = ~n6679 & ~n6680;
  assign n6683 = ~n6681 & ~n6682;
  assign n6684 = ~n6388 & ~n6390;
  assign n6685 = ~n6683 & ~n6684;
  assign n6686 = n6683 & n6684;
  assign n6687 = ~n6685 & ~n6686;
  assign n6688 = ~n6512 & n6687;
  assign n6689 = ~n6512 & ~n6688;
  assign n6690 = n6687 & ~n6688;
  assign n6691 = ~n6689 & ~n6690;
  assign n6692 = ~n6501 & ~n6691;
  assign n6693 = ~n6501 & ~n6692;
  assign n6694 = ~n6691 & ~n6692;
  assign n6695 = ~n6693 & ~n6694;
  assign n6696 = n938 & n3784;
  assign n6697 = pi93  & n1052;
  assign n6698 = pi95  & n936;
  assign n6699 = pi94  & n931;
  assign n6700 = ~n6698 & ~n6699;
  assign n6701 = ~n6697 & n6700;
  assign n6702 = ~n6696 & n6701;
  assign n6703 = pi14  & ~n6702;
  assign n6704 = pi14  & ~n6703;
  assign n6705 = ~n6702 & ~n6703;
  assign n6706 = ~n6704 & ~n6705;
  assign n6707 = n6695 & n6706;
  assign n6708 = ~n6695 & ~n6706;
  assign n6709 = ~n6707 & ~n6708;
  assign n6710 = ~n6499 & n6709;
  assign n6711 = n6499 & ~n6709;
  assign n6712 = ~n6710 & ~n6711;
  assign n6713 = n687 & n4454;
  assign n6714 = pi96  & n763;
  assign n6715 = pi98  & n685;
  assign n6716 = pi97  & n680;
  assign n6717 = ~n6715 & ~n6716;
  assign n6718 = ~n6714 & n6717;
  assign n6719 = ~n6713 & n6718;
  assign n6720 = pi11  & ~n6719;
  assign n6721 = pi11  & ~n6720;
  assign n6722 = ~n6719 & ~n6720;
  assign n6723 = ~n6721 & ~n6722;
  assign n6724 = n6712 & ~n6723;
  assign n6725 = n6712 & ~n6724;
  assign n6726 = ~n6723 & ~n6724;
  assign n6727 = ~n6725 & ~n6726;
  assign n6728 = ~n6239 & ~n6442;
  assign n6729 = ~n6439 & ~n6728;
  assign n6730 = n6727 & n6729;
  assign n6731 = ~n6727 & ~n6729;
  assign n6732 = ~n6730 & ~n6731;
  assign n6733 = n498 & n5169;
  assign n6734 = pi99  & n537;
  assign n6735 = pi101  & n496;
  assign n6736 = pi100  & n491;
  assign n6737 = ~n6735 & ~n6736;
  assign n6738 = ~n6734 & n6737;
  assign n6739 = ~n6733 & n6738;
  assign n6740 = pi8  & ~n6739;
  assign n6741 = pi8  & ~n6740;
  assign n6742 = ~n6739 & ~n6740;
  assign n6743 = ~n6741 & ~n6742;
  assign n6744 = n6732 & ~n6743;
  assign n6745 = ~n6732 & n6743;
  assign n6746 = ~n6744 & ~n6745;
  assign n6747 = ~n6498 & n6746;
  assign n6748 = ~n6498 & ~n6747;
  assign n6749 = ~n6744 & ~n6747;
  assign n6750 = ~n6745 & n6749;
  assign n6751 = ~n6748 & ~n6750;
  assign n6752 = n342 & n5943;
  assign n6753 = pi102  & n380;
  assign n6754 = pi104  & n340;
  assign n6755 = pi103  & n335;
  assign n6756 = ~n6754 & ~n6755;
  assign n6757 = ~n6753 & n6756;
  assign n6758 = ~n6752 & n6757;
  assign n6759 = pi5  & ~n6758;
  assign n6760 = pi5  & ~n6759;
  assign n6761 = ~n6758 & ~n6759;
  assign n6762 = ~n6760 & ~n6761;
  assign n6763 = n6751 & n6762;
  assign n6764 = ~n6751 & ~n6762;
  assign n6765 = ~n6763 & ~n6764;
  assign n6766 = ~n6497 & n6765;
  assign n6767 = n6497 & ~n6765;
  assign n6768 = ~n6766 & ~n6767;
  assign n6769 = ~n6473 & ~n6475;
  assign n6770 = ~pi106  & ~pi107 ;
  assign n6771 = pi106  & pi107 ;
  assign n6772 = ~n6770 & ~n6771;
  assign n6773 = ~n6769 & n6772;
  assign n6774 = n6769 & ~n6772;
  assign n6775 = ~n6773 & ~n6774;
  assign n6776 = n262 & n6775;
  assign n6777 = pi105  & n288;
  assign n6778 = pi107  & n267;
  assign n6779 = pi106  & n269;
  assign n6780 = ~n6778 & ~n6779;
  assign n6781 = ~n6777 & n6780;
  assign n6782 = ~n6776 & n6781;
  assign n6783 = pi2  & ~n6782;
  assign n6784 = pi2  & ~n6783;
  assign n6785 = ~n6782 & ~n6783;
  assign n6786 = ~n6784 & ~n6785;
  assign n6787 = n6768 & ~n6786;
  assign n6788 = n6768 & ~n6787;
  assign n6789 = ~n6786 & ~n6787;
  assign n6790 = ~n6788 & ~n6789;
  assign n6791 = ~n6489 & ~n6494;
  assign n6792 = ~n6790 & ~n6791;
  assign n6793 = n6790 & n6791;
  assign po43  = ~n6792 & ~n6793;
  assign n6795 = ~n6787 & ~n6792;
  assign n6796 = ~n6764 & ~n6766;
  assign n6797 = n342 & n6207;
  assign n6798 = pi103  & n380;
  assign n6799 = pi105  & n340;
  assign n6800 = pi104  & n335;
  assign n6801 = ~n6799 & ~n6800;
  assign n6802 = ~n6798 & n6801;
  assign n6803 = ~n6797 & n6802;
  assign n6804 = pi5  & ~n6803;
  assign n6805 = pi5  & ~n6804;
  assign n6806 = ~n6803 & ~n6804;
  assign n6807 = ~n6805 & ~n6806;
  assign n6808 = ~n6708 & ~n6710;
  assign n6809 = n938 & n4001;
  assign n6810 = pi94  & n1052;
  assign n6811 = pi96  & n936;
  assign n6812 = pi95  & n931;
  assign n6813 = ~n6811 & ~n6812;
  assign n6814 = ~n6810 & n6813;
  assign n6815 = ~n6809 & n6814;
  assign n6816 = pi14  & ~n6815;
  assign n6817 = pi14  & ~n6816;
  assign n6818 = ~n6815 & ~n6816;
  assign n6819 = ~n6817 & ~n6818;
  assign n6820 = ~n6688 & ~n6692;
  assign n6821 = n1297 & n3371;
  assign n6822 = pi91  & n1366;
  assign n6823 = pi93  & n1295;
  assign n6824 = pi92  & n1290;
  assign n6825 = ~n6823 & ~n6824;
  assign n6826 = ~n6822 & n6825;
  assign n6827 = ~n6821 & n6826;
  assign n6828 = pi17  & ~n6827;
  assign n6829 = pi17  & ~n6828;
  assign n6830 = ~n6827 & ~n6828;
  assign n6831 = ~n6829 & ~n6830;
  assign n6832 = ~n6680 & ~n6685;
  assign n6833 = ~n6661 & ~n6667;
  assign n6834 = ~n6622 & ~n6629;
  assign n6835 = n1434 & n3034;
  assign n6836 = pi79  & n3225;
  assign n6837 = pi81  & n3032;
  assign n6838 = pi80  & n3027;
  assign n6839 = ~n6837 & ~n6838;
  assign n6840 = ~n6836 & n6839;
  assign n6841 = ~n6835 & n6840;
  assign n6842 = pi29  & ~n6841;
  assign n6843 = pi29  & ~n6842;
  assign n6844 = ~n6841 & ~n6842;
  assign n6845 = ~n6843 & ~n6844;
  assign n6846 = ~n6606 & ~n6608;
  assign n6847 = n1025 & n3622;
  assign n6848 = pi76  & n3814;
  assign n6849 = pi78  & n3620;
  assign n6850 = pi77  & n3615;
  assign n6851 = ~n6849 & ~n6850;
  assign n6852 = ~n6848 & n6851;
  assign n6853 = ~n6847 & n6852;
  assign n6854 = pi32  & ~n6853;
  assign n6855 = pi32  & ~n6854;
  assign n6856 = ~n6853 & ~n6854;
  assign n6857 = ~n6855 & ~n6856;
  assign n6858 = ~n6567 & ~n6573;
  assign n6859 = n576 & n5008;
  assign n6860 = pi70  & n5241;
  assign n6861 = pi72  & n5006;
  assign n6862 = pi71  & n5001;
  assign n6863 = ~n6861 & ~n6862;
  assign n6864 = ~n6860 & n6863;
  assign n6865 = ~n6859 & n6864;
  assign n6866 = pi38  & ~n6865;
  assign n6867 = pi38  & ~n6866;
  assign n6868 = ~n6865 & ~n6866;
  assign n6869 = ~n6867 & ~n6868;
  assign n6870 = ~n6551 & ~n6553;
  assign n6871 = n286 & n6539;
  assign n6872 = n6259 & n6531;
  assign n6873 = ~n6536 & n6872;
  assign n6874 = pi64  & n6873;
  assign n6875 = pi66  & n6537;
  assign n6876 = pi65  & n6532;
  assign n6877 = ~n6875 & ~n6876;
  assign n6878 = ~n6871 & n6877;
  assign n6879 = ~n6874 & n6878;
  assign n6880 = pi44  & ~n6879;
  assign n6881 = pi44  & ~n6880;
  assign n6882 = ~n6879 & ~n6880;
  assign n6883 = ~n6881 & ~n6882;
  assign n6884 = ~n6547 & n6883;
  assign n6885 = n6547 & ~n6883;
  assign n6886 = ~n6884 & ~n6885;
  assign n6887 = n401 & n5739;
  assign n6888 = pi67  & n6030;
  assign n6889 = pi69  & n5737;
  assign n6890 = pi68  & n5732;
  assign n6891 = ~n6889 & ~n6890;
  assign n6892 = ~n6888 & n6891;
  assign n6893 = ~n6887 & n6892;
  assign n6894 = pi41  & ~n6893;
  assign n6895 = pi41  & ~n6894;
  assign n6896 = ~n6893 & ~n6894;
  assign n6897 = ~n6895 & ~n6896;
  assign n6898 = n6886 & ~n6897;
  assign n6899 = n6886 & ~n6898;
  assign n6900 = ~n6897 & ~n6898;
  assign n6901 = ~n6899 & ~n6900;
  assign n6902 = ~n6870 & ~n6901;
  assign n6903 = n6870 & n6901;
  assign n6904 = ~n6902 & ~n6903;
  assign n6905 = ~n6869 & n6904;
  assign n6906 = ~n6869 & ~n6905;
  assign n6907 = n6904 & ~n6905;
  assign n6908 = ~n6906 & ~n6907;
  assign n6909 = ~n6858 & ~n6908;
  assign n6910 = ~n6858 & ~n6909;
  assign n6911 = ~n6908 & ~n6909;
  assign n6912 = ~n6910 & ~n6911;
  assign n6913 = n809 & n4271;
  assign n6914 = pi73  & n4503;
  assign n6915 = pi75  & n4269;
  assign n6916 = pi74  & n4264;
  assign n6917 = ~n6915 & ~n6916;
  assign n6918 = ~n6914 & n6917;
  assign n6919 = ~n6913 & n6918;
  assign n6920 = pi35  & ~n6919;
  assign n6921 = pi35  & ~n6920;
  assign n6922 = ~n6919 & ~n6920;
  assign n6923 = ~n6921 & ~n6922;
  assign n6924 = n6912 & n6923;
  assign n6925 = ~n6912 & ~n6923;
  assign n6926 = ~n6924 & ~n6925;
  assign n6927 = ~n6591 & n6926;
  assign n6928 = n6591 & ~n6926;
  assign n6929 = ~n6927 & ~n6928;
  assign n6930 = n6857 & ~n6929;
  assign n6931 = ~n6857 & n6929;
  assign n6932 = ~n6930 & ~n6931;
  assign n6933 = ~n6846 & n6932;
  assign n6934 = n6846 & ~n6932;
  assign n6935 = ~n6933 & ~n6934;
  assign n6936 = n6845 & ~n6935;
  assign n6937 = ~n6845 & n6935;
  assign n6938 = ~n6936 & ~n6937;
  assign n6939 = ~n6834 & n6938;
  assign n6940 = n6834 & ~n6938;
  assign n6941 = ~n6939 & ~n6940;
  assign n6942 = n1834 & n2523;
  assign n6943 = pi82  & n2667;
  assign n6944 = pi84  & n2521;
  assign n6945 = pi83  & n2516;
  assign n6946 = ~n6944 & ~n6945;
  assign n6947 = ~n6943 & n6946;
  assign n6948 = ~n6942 & n6947;
  assign n6949 = pi26  & ~n6948;
  assign n6950 = pi26  & ~n6949;
  assign n6951 = ~n6948 & ~n6949;
  assign n6952 = ~n6950 & ~n6951;
  assign n6953 = n6941 & ~n6952;
  assign n6954 = n6941 & ~n6953;
  assign n6955 = ~n6952 & ~n6953;
  assign n6956 = ~n6954 & ~n6955;
  assign n6957 = ~n6642 & ~n6648;
  assign n6958 = n6956 & n6957;
  assign n6959 = ~n6956 & ~n6957;
  assign n6960 = ~n6958 & ~n6959;
  assign n6961 = n2043 & n2288;
  assign n6962 = pi85  & n2180;
  assign n6963 = pi87  & n2041;
  assign n6964 = pi86  & n2036;
  assign n6965 = ~n6963 & ~n6964;
  assign n6966 = ~n6962 & n6965;
  assign n6967 = ~n6961 & n6966;
  assign n6968 = pi23  & ~n6967;
  assign n6969 = pi23  & ~n6968;
  assign n6970 = ~n6967 & ~n6968;
  assign n6971 = ~n6969 & ~n6970;
  assign n6972 = n6960 & ~n6971;
  assign n6973 = ~n6960 & n6971;
  assign n6974 = ~n6972 & ~n6973;
  assign n6975 = ~n6833 & n6974;
  assign n6976 = ~n6833 & ~n6975;
  assign n6977 = ~n6972 & ~n6975;
  assign n6978 = ~n6973 & n6977;
  assign n6979 = ~n6976 & ~n6978;
  assign n6980 = n1611 & n2801;
  assign n6981 = pi88  & n1745;
  assign n6982 = pi90  & n1609;
  assign n6983 = pi89  & n1604;
  assign n6984 = ~n6982 & ~n6983;
  assign n6985 = ~n6981 & n6984;
  assign n6986 = ~n6980 & n6985;
  assign n6987 = pi20  & ~n6986;
  assign n6988 = pi20  & ~n6987;
  assign n6989 = ~n6986 & ~n6987;
  assign n6990 = ~n6988 & ~n6989;
  assign n6991 = n6979 & n6990;
  assign n6992 = ~n6979 & ~n6990;
  assign n6993 = ~n6991 & ~n6992;
  assign n6994 = ~n6832 & n6993;
  assign n6995 = n6832 & ~n6993;
  assign n6996 = ~n6994 & ~n6995;
  assign n6997 = n6831 & ~n6996;
  assign n6998 = ~n6831 & n6996;
  assign n6999 = ~n6997 & ~n6998;
  assign n7000 = ~n6820 & n6999;
  assign n7001 = n6820 & ~n6999;
  assign n7002 = ~n7000 & ~n7001;
  assign n7003 = n6819 & ~n7002;
  assign n7004 = ~n6819 & n7002;
  assign n7005 = ~n7003 & ~n7004;
  assign n7006 = ~n6808 & n7005;
  assign n7007 = n6808 & ~n7005;
  assign n7008 = ~n7006 & ~n7007;
  assign n7009 = n687 & n4684;
  assign n7010 = pi97  & n763;
  assign n7011 = pi99  & n685;
  assign n7012 = pi98  & n680;
  assign n7013 = ~n7011 & ~n7012;
  assign n7014 = ~n7010 & n7013;
  assign n7015 = ~n7009 & n7014;
  assign n7016 = pi11  & ~n7015;
  assign n7017 = pi11  & ~n7016;
  assign n7018 = ~n7015 & ~n7016;
  assign n7019 = ~n7017 & ~n7018;
  assign n7020 = n7008 & ~n7019;
  assign n7021 = n7008 & ~n7020;
  assign n7022 = ~n7019 & ~n7020;
  assign n7023 = ~n7021 & ~n7022;
  assign n7024 = ~n6724 & ~n6731;
  assign n7025 = n7023 & n7024;
  assign n7026 = ~n7023 & ~n7024;
  assign n7027 = ~n7025 & ~n7026;
  assign n7028 = n498 & n5413;
  assign n7029 = pi100  & n537;
  assign n7030 = pi102  & n496;
  assign n7031 = pi101  & n491;
  assign n7032 = ~n7030 & ~n7031;
  assign n7033 = ~n7029 & n7032;
  assign n7034 = ~n7028 & n7033;
  assign n7035 = pi8  & ~n7034;
  assign n7036 = pi8  & ~n7035;
  assign n7037 = ~n7034 & ~n7035;
  assign n7038 = ~n7036 & ~n7037;
  assign n7039 = n7027 & ~n7038;
  assign n7040 = n7027 & ~n7039;
  assign n7041 = ~n7038 & ~n7039;
  assign n7042 = ~n7040 & ~n7041;
  assign n7043 = ~n6749 & ~n7042;
  assign n7044 = n6749 & n7042;
  assign n7045 = ~n7043 & ~n7044;
  assign n7046 = ~n6807 & n7045;
  assign n7047 = ~n6807 & ~n7046;
  assign n7048 = n7045 & ~n7046;
  assign n7049 = ~n7047 & ~n7048;
  assign n7050 = ~n6796 & ~n7049;
  assign n7051 = ~n6796 & ~n7050;
  assign n7052 = ~n7049 & ~n7050;
  assign n7053 = ~n7051 & ~n7052;
  assign n7054 = ~n6771 & ~n6773;
  assign n7055 = ~pi107  & ~pi108 ;
  assign n7056 = pi107  & pi108 ;
  assign n7057 = ~n7055 & ~n7056;
  assign n7058 = ~n7054 & n7057;
  assign n7059 = n7054 & ~n7057;
  assign n7060 = ~n7058 & ~n7059;
  assign n7061 = n262 & n7060;
  assign n7062 = pi106  & n288;
  assign n7063 = pi108  & n267;
  assign n7064 = pi107  & n269;
  assign n7065 = ~n7063 & ~n7064;
  assign n7066 = ~n7062 & n7065;
  assign n7067 = ~n7061 & n7066;
  assign n7068 = pi2  & ~n7067;
  assign n7069 = pi2  & ~n7068;
  assign n7070 = ~n7067 & ~n7068;
  assign n7071 = ~n7069 & ~n7070;
  assign n7072 = ~n7053 & n7071;
  assign n7073 = n7053 & ~n7071;
  assign n7074 = ~n7072 & ~n7073;
  assign n7075 = ~n6795 & ~n7074;
  assign n7076 = n6795 & n7074;
  assign po44  = ~n7075 & ~n7076;
  assign n7078 = ~n7053 & ~n7071;
  assign n7079 = ~n7075 & ~n7078;
  assign n7080 = ~n7020 & ~n7026;
  assign n7081 = ~n7004 & ~n7006;
  assign n7082 = ~n6998 & ~n7000;
  assign n7083 = ~n6992 & ~n6994;
  assign n7084 = ~n6937 & ~n6939;
  assign n7085 = ~n6931 & ~n6933;
  assign n7086 = ~n6925 & ~n6927;
  assign n7087 = n891 & n4271;
  assign n7088 = pi74  & n4503;
  assign n7089 = pi76  & n4269;
  assign n7090 = pi75  & n4264;
  assign n7091 = ~n7089 & ~n7090;
  assign n7092 = ~n7088 & n7091;
  assign n7093 = ~n7087 & n7092;
  assign n7094 = pi35  & ~n7093;
  assign n7095 = pi35  & ~n7094;
  assign n7096 = ~n7093 & ~n7094;
  assign n7097 = ~n7095 & ~n7096;
  assign n7098 = ~n6905 & ~n6909;
  assign n7099 = pi44  & ~pi45 ;
  assign n7100 = ~pi44  & pi45 ;
  assign n7101 = ~n7099 & ~n7100;
  assign n7102 = pi64  & ~n7101;
  assign n7103 = ~n6885 & n7102;
  assign n7104 = n6885 & ~n7102;
  assign n7105 = ~n7103 & ~n7104;
  assign n7106 = n309 & n6539;
  assign n7107 = pi65  & n6873;
  assign n7108 = pi67  & n6537;
  assign n7109 = pi66  & n6532;
  assign n7110 = ~n7108 & ~n7109;
  assign n7111 = ~n7107 & n7110;
  assign n7112 = ~n7106 & n7111;
  assign n7113 = pi44  & ~n7112;
  assign n7114 = pi44  & ~n7113;
  assign n7115 = ~n7112 & ~n7113;
  assign n7116 = ~n7114 & ~n7115;
  assign n7117 = ~n7105 & ~n7116;
  assign n7118 = n7105 & n7116;
  assign n7119 = ~n7117 & ~n7118;
  assign n7120 = n450 & n5739;
  assign n7121 = pi68  & n6030;
  assign n7122 = pi70  & n5737;
  assign n7123 = pi69  & n5732;
  assign n7124 = ~n7122 & ~n7123;
  assign n7125 = ~n7121 & n7124;
  assign n7126 = ~n7120 & n7125;
  assign n7127 = pi41  & ~n7126;
  assign n7128 = pi41  & ~n7127;
  assign n7129 = ~n7126 & ~n7127;
  assign n7130 = ~n7128 & ~n7129;
  assign n7131 = n7119 & ~n7130;
  assign n7132 = n7119 & ~n7131;
  assign n7133 = ~n7130 & ~n7131;
  assign n7134 = ~n7132 & ~n7133;
  assign n7135 = ~n6898 & ~n6902;
  assign n7136 = n7134 & n7135;
  assign n7137 = ~n7134 & ~n7135;
  assign n7138 = ~n7136 & ~n7137;
  assign n7139 = n642 & n5008;
  assign n7140 = pi71  & n5241;
  assign n7141 = pi73  & n5006;
  assign n7142 = pi72  & n5001;
  assign n7143 = ~n7141 & ~n7142;
  assign n7144 = ~n7140 & n7143;
  assign n7145 = ~n7139 & n7144;
  assign n7146 = pi38  & ~n7145;
  assign n7147 = pi38  & ~n7146;
  assign n7148 = ~n7145 & ~n7146;
  assign n7149 = ~n7147 & ~n7148;
  assign n7150 = ~n7138 & n7149;
  assign n7151 = n7138 & ~n7149;
  assign n7152 = ~n7150 & ~n7151;
  assign n7153 = ~n7098 & n7152;
  assign n7154 = n7098 & ~n7152;
  assign n7155 = ~n7153 & ~n7154;
  assign n7156 = ~n7097 & n7155;
  assign n7157 = ~n7097 & ~n7156;
  assign n7158 = n7155 & ~n7156;
  assign n7159 = ~n7157 & ~n7158;
  assign n7160 = ~n7086 & ~n7159;
  assign n7161 = ~n7086 & ~n7160;
  assign n7162 = ~n7159 & ~n7160;
  assign n7163 = ~n7161 & ~n7162;
  assign n7164 = n1122 & n3622;
  assign n7165 = pi77  & n3814;
  assign n7166 = pi79  & n3620;
  assign n7167 = pi78  & n3615;
  assign n7168 = ~n7166 & ~n7167;
  assign n7169 = ~n7165 & n7168;
  assign n7170 = ~n7164 & n7169;
  assign n7171 = pi32  & ~n7170;
  assign n7172 = pi32  & ~n7171;
  assign n7173 = ~n7170 & ~n7171;
  assign n7174 = ~n7172 & ~n7173;
  assign n7175 = ~n7163 & ~n7174;
  assign n7176 = ~n7163 & ~n7175;
  assign n7177 = ~n7174 & ~n7175;
  assign n7178 = ~n7176 & ~n7177;
  assign n7179 = ~n7085 & n7178;
  assign n7180 = n7085 & ~n7178;
  assign n7181 = ~n7179 & ~n7180;
  assign n7182 = n1554 & n3034;
  assign n7183 = pi80  & n3225;
  assign n7184 = pi82  & n3032;
  assign n7185 = pi81  & n3027;
  assign n7186 = ~n7184 & ~n7185;
  assign n7187 = ~n7183 & n7186;
  assign n7188 = ~n7182 & n7187;
  assign n7189 = pi29  & ~n7188;
  assign n7190 = pi29  & ~n7189;
  assign n7191 = ~n7188 & ~n7189;
  assign n7192 = ~n7190 & ~n7191;
  assign n7193 = ~n7181 & ~n7192;
  assign n7194 = n7181 & n7192;
  assign n7195 = ~n7193 & ~n7194;
  assign n7196 = ~n7084 & n7195;
  assign n7197 = n7084 & ~n7195;
  assign n7198 = ~n7196 & ~n7197;
  assign n7199 = n1972 & n2523;
  assign n7200 = pi83  & n2667;
  assign n7201 = pi85  & n2521;
  assign n7202 = pi84  & n2516;
  assign n7203 = ~n7201 & ~n7202;
  assign n7204 = ~n7200 & n7203;
  assign n7205 = ~n7199 & n7204;
  assign n7206 = pi26  & ~n7205;
  assign n7207 = pi26  & ~n7206;
  assign n7208 = ~n7205 & ~n7206;
  assign n7209 = ~n7207 & ~n7208;
  assign n7210 = n7198 & ~n7209;
  assign n7211 = n7198 & ~n7210;
  assign n7212 = ~n7209 & ~n7210;
  assign n7213 = ~n7211 & ~n7212;
  assign n7214 = ~n6953 & ~n6959;
  assign n7215 = n7213 & n7214;
  assign n7216 = ~n7213 & ~n7214;
  assign n7217 = ~n7215 & ~n7216;
  assign n7218 = n2043 & n2446;
  assign n7219 = pi86  & n2180;
  assign n7220 = pi88  & n2041;
  assign n7221 = pi87  & n2036;
  assign n7222 = ~n7220 & ~n7221;
  assign n7223 = ~n7219 & n7222;
  assign n7224 = ~n7218 & n7223;
  assign n7225 = pi23  & ~n7224;
  assign n7226 = pi23  & ~n7225;
  assign n7227 = ~n7224 & ~n7225;
  assign n7228 = ~n7226 & ~n7227;
  assign n7229 = ~n7217 & n7228;
  assign n7230 = n7217 & ~n7228;
  assign n7231 = ~n7229 & ~n7230;
  assign n7232 = ~n6977 & n7231;
  assign n7233 = n6977 & ~n7231;
  assign n7234 = ~n7232 & ~n7233;
  assign n7235 = n1611 & n2978;
  assign n7236 = pi89  & n1745;
  assign n7237 = pi91  & n1609;
  assign n7238 = pi90  & n1604;
  assign n7239 = ~n7237 & ~n7238;
  assign n7240 = ~n7236 & n7239;
  assign n7241 = ~n7235 & n7240;
  assign n7242 = pi20  & ~n7241;
  assign n7243 = pi20  & ~n7242;
  assign n7244 = ~n7241 & ~n7242;
  assign n7245 = ~n7243 & ~n7244;
  assign n7246 = n7234 & ~n7245;
  assign n7247 = n7234 & ~n7246;
  assign n7248 = ~n7245 & ~n7246;
  assign n7249 = ~n7247 & ~n7248;
  assign n7250 = ~n7083 & n7249;
  assign n7251 = n7083 & ~n7249;
  assign n7252 = ~n7250 & ~n7251;
  assign n7253 = n1297 & n3565;
  assign n7254 = pi92  & n1366;
  assign n7255 = pi94  & n1295;
  assign n7256 = pi93  & n1290;
  assign n7257 = ~n7255 & ~n7256;
  assign n7258 = ~n7254 & n7257;
  assign n7259 = ~n7253 & n7258;
  assign n7260 = pi17  & ~n7259;
  assign n7261 = pi17  & ~n7260;
  assign n7262 = ~n7259 & ~n7260;
  assign n7263 = ~n7261 & ~n7262;
  assign n7264 = ~n7252 & ~n7263;
  assign n7265 = n7252 & n7263;
  assign n7266 = ~n7264 & ~n7265;
  assign n7267 = ~n7082 & n7266;
  assign n7268 = n7082 & ~n7266;
  assign n7269 = ~n7267 & ~n7268;
  assign n7270 = n938 & n4211;
  assign n7271 = pi95  & n1052;
  assign n7272 = pi97  & n936;
  assign n7273 = pi96  & n931;
  assign n7274 = ~n7272 & ~n7273;
  assign n7275 = ~n7271 & n7274;
  assign n7276 = ~n7270 & n7275;
  assign n7277 = pi14  & ~n7276;
  assign n7278 = pi14  & ~n7277;
  assign n7279 = ~n7276 & ~n7277;
  assign n7280 = ~n7278 & ~n7279;
  assign n7281 = n7269 & ~n7280;
  assign n7282 = n7269 & ~n7281;
  assign n7283 = ~n7280 & ~n7281;
  assign n7284 = ~n7282 & ~n7283;
  assign n7285 = ~n7081 & n7284;
  assign n7286 = n7081 & ~n7284;
  assign n7287 = ~n7285 & ~n7286;
  assign n7288 = n687 & n4910;
  assign n7289 = pi98  & n763;
  assign n7290 = pi100  & n685;
  assign n7291 = pi99  & n680;
  assign n7292 = ~n7290 & ~n7291;
  assign n7293 = ~n7289 & n7292;
  assign n7294 = ~n7288 & n7293;
  assign n7295 = pi11  & ~n7294;
  assign n7296 = pi11  & ~n7295;
  assign n7297 = ~n7294 & ~n7295;
  assign n7298 = ~n7296 & ~n7297;
  assign n7299 = ~n7287 & ~n7298;
  assign n7300 = n7287 & n7298;
  assign n7301 = ~n7299 & ~n7300;
  assign n7302 = n7080 & ~n7301;
  assign n7303 = ~n7080 & n7301;
  assign n7304 = ~n7302 & ~n7303;
  assign n7305 = n498 & n5664;
  assign n7306 = pi101  & n537;
  assign n7307 = pi103  & n496;
  assign n7308 = pi102  & n491;
  assign n7309 = ~n7307 & ~n7308;
  assign n7310 = ~n7306 & n7309;
  assign n7311 = ~n7305 & n7310;
  assign n7312 = pi8  & ~n7311;
  assign n7313 = pi8  & ~n7312;
  assign n7314 = ~n7311 & ~n7312;
  assign n7315 = ~n7313 & ~n7314;
  assign n7316 = n7304 & ~n7315;
  assign n7317 = n7304 & ~n7316;
  assign n7318 = ~n7315 & ~n7316;
  assign n7319 = ~n7317 & ~n7318;
  assign n7320 = ~n7039 & ~n7043;
  assign n7321 = n7319 & n7320;
  assign n7322 = ~n7319 & ~n7320;
  assign n7323 = ~n7321 & ~n7322;
  assign n7324 = n342 & n6477;
  assign n7325 = pi104  & n380;
  assign n7326 = pi106  & n340;
  assign n7327 = pi105  & n335;
  assign n7328 = ~n7326 & ~n7327;
  assign n7329 = ~n7325 & n7328;
  assign n7330 = ~n7324 & n7329;
  assign n7331 = pi5  & ~n7330;
  assign n7332 = pi5  & ~n7331;
  assign n7333 = ~n7330 & ~n7331;
  assign n7334 = ~n7332 & ~n7333;
  assign n7335 = n7323 & ~n7334;
  assign n7336 = n7323 & ~n7335;
  assign n7337 = ~n7334 & ~n7335;
  assign n7338 = ~n7336 & ~n7337;
  assign n7339 = ~n7046 & ~n7050;
  assign n7340 = n7338 & n7339;
  assign n7341 = ~n7338 & ~n7339;
  assign n7342 = ~n7340 & ~n7341;
  assign n7343 = ~n7056 & ~n7058;
  assign n7344 = ~pi108  & ~pi109 ;
  assign n7345 = pi108  & pi109 ;
  assign n7346 = ~n7344 & ~n7345;
  assign n7347 = ~n7343 & n7346;
  assign n7348 = n7343 & ~n7346;
  assign n7349 = ~n7347 & ~n7348;
  assign n7350 = n262 & n7349;
  assign n7351 = pi107  & n288;
  assign n7352 = pi109  & n267;
  assign n7353 = pi108  & n269;
  assign n7354 = ~n7352 & ~n7353;
  assign n7355 = ~n7351 & n7354;
  assign n7356 = ~n7350 & n7355;
  assign n7357 = pi2  & ~n7356;
  assign n7358 = pi2  & ~n7357;
  assign n7359 = ~n7356 & ~n7357;
  assign n7360 = ~n7358 & ~n7359;
  assign n7361 = ~n7342 & n7360;
  assign n7362 = n7342 & ~n7360;
  assign n7363 = ~n7361 & ~n7362;
  assign n7364 = ~n7079 & n7363;
  assign n7365 = n7079 & ~n7363;
  assign po45  = ~n7364 & ~n7365;
  assign n7367 = ~n7316 & ~n7322;
  assign n7368 = ~n7264 & ~n7267;
  assign n7369 = ~n7083 & ~n7249;
  assign n7370 = ~n7246 & ~n7369;
  assign n7371 = n1611 & n3177;
  assign n7372 = pi90  & n1745;
  assign n7373 = pi92  & n1609;
  assign n7374 = pi91  & n1604;
  assign n7375 = ~n7373 & ~n7374;
  assign n7376 = ~n7372 & n7375;
  assign n7377 = ~n7371 & n7376;
  assign n7378 = pi20  & ~n7377;
  assign n7379 = pi20  & ~n7378;
  assign n7380 = ~n7377 & ~n7378;
  assign n7381 = ~n7379 & ~n7380;
  assign n7382 = ~n7156 & ~n7160;
  assign n7383 = ~n7151 & ~n7153;
  assign n7384 = n6885 & n7102;
  assign n7385 = ~n7117 & ~n7384;
  assign n7386 = n359 & n6539;
  assign n7387 = pi66  & n6873;
  assign n7388 = pi68  & n6537;
  assign n7389 = pi67  & n6532;
  assign n7390 = ~n7388 & ~n7389;
  assign n7391 = ~n7387 & n7390;
  assign n7392 = ~n7386 & n7391;
  assign n7393 = pi44  & ~n7392;
  assign n7394 = pi44  & ~n7393;
  assign n7395 = ~n7392 & ~n7393;
  assign n7396 = ~n7394 & ~n7395;
  assign n7397 = pi47  & ~n7102;
  assign n7398 = ~pi45  & pi46 ;
  assign n7399 = pi45  & ~pi46 ;
  assign n7400 = ~n7398 & ~n7399;
  assign n7401 = n7101 & ~n7400;
  assign n7402 = pi64  & n7401;
  assign n7403 = ~pi46  & pi47 ;
  assign n7404 = pi46  & ~pi47 ;
  assign n7405 = ~n7403 & ~n7404;
  assign n7406 = ~n7101 & n7405;
  assign n7407 = pi65  & n7406;
  assign n7408 = ~n7101 & ~n7405;
  assign n7409 = ~n265 & n7408;
  assign n7410 = ~n7402 & ~n7407;
  assign n7411 = ~n7409 & n7410;
  assign n7412 = pi47  & ~n7411;
  assign n7413 = pi47  & ~n7412;
  assign n7414 = ~n7411 & ~n7412;
  assign n7415 = ~n7413 & ~n7414;
  assign n7416 = n7397 & ~n7415;
  assign n7417 = ~n7397 & n7415;
  assign n7418 = ~n7416 & ~n7417;
  assign n7419 = n7396 & ~n7418;
  assign n7420 = ~n7396 & n7418;
  assign n7421 = ~n7419 & ~n7420;
  assign n7422 = ~n7385 & n7421;
  assign n7423 = n7385 & ~n7421;
  assign n7424 = ~n7422 & ~n7423;
  assign n7425 = n475 & n5739;
  assign n7426 = pi69  & n6030;
  assign n7427 = pi71  & n5737;
  assign n7428 = pi70  & n5732;
  assign n7429 = ~n7427 & ~n7428;
  assign n7430 = ~n7426 & n7429;
  assign n7431 = ~n7425 & n7430;
  assign n7432 = pi41  & ~n7431;
  assign n7433 = pi41  & ~n7432;
  assign n7434 = ~n7431 & ~n7432;
  assign n7435 = ~n7433 & ~n7434;
  assign n7436 = n7424 & ~n7435;
  assign n7437 = n7424 & ~n7436;
  assign n7438 = ~n7435 & ~n7436;
  assign n7439 = ~n7437 & ~n7438;
  assign n7440 = ~n7131 & ~n7137;
  assign n7441 = n7439 & n7440;
  assign n7442 = ~n7439 & ~n7440;
  assign n7443 = ~n7441 & ~n7442;
  assign n7444 = n729 & n5008;
  assign n7445 = pi72  & n5241;
  assign n7446 = pi74  & n5006;
  assign n7447 = pi73  & n5001;
  assign n7448 = ~n7446 & ~n7447;
  assign n7449 = ~n7445 & n7448;
  assign n7450 = ~n7444 & n7449;
  assign n7451 = pi38  & ~n7450;
  assign n7452 = pi38  & ~n7451;
  assign n7453 = ~n7450 & ~n7451;
  assign n7454 = ~n7452 & ~n7453;
  assign n7455 = n7443 & ~n7454;
  assign n7456 = ~n7443 & n7454;
  assign n7457 = ~n7455 & ~n7456;
  assign n7458 = ~n7383 & n7457;
  assign n7459 = ~n7383 & ~n7458;
  assign n7460 = ~n7455 & ~n7458;
  assign n7461 = ~n7456 & n7460;
  assign n7462 = ~n7459 & ~n7461;
  assign n7463 = n999 & n4271;
  assign n7464 = pi75  & n4503;
  assign n7465 = pi77  & n4269;
  assign n7466 = pi76  & n4264;
  assign n7467 = ~n7465 & ~n7466;
  assign n7468 = ~n7464 & n7467;
  assign n7469 = ~n7463 & n7468;
  assign n7470 = pi35  & ~n7469;
  assign n7471 = pi35  & ~n7470;
  assign n7472 = ~n7469 & ~n7470;
  assign n7473 = ~n7471 & ~n7472;
  assign n7474 = n7462 & n7473;
  assign n7475 = ~n7462 & ~n7473;
  assign n7476 = ~n7474 & ~n7475;
  assign n7477 = ~n7382 & n7476;
  assign n7478 = n7382 & ~n7476;
  assign n7479 = ~n7477 & ~n7478;
  assign n7480 = n1225 & n3622;
  assign n7481 = pi78  & n3814;
  assign n7482 = pi80  & n3620;
  assign n7483 = pi79  & n3615;
  assign n7484 = ~n7482 & ~n7483;
  assign n7485 = ~n7481 & n7484;
  assign n7486 = ~n7480 & n7485;
  assign n7487 = pi32  & ~n7486;
  assign n7488 = pi32  & ~n7487;
  assign n7489 = ~n7486 & ~n7487;
  assign n7490 = ~n7488 & ~n7489;
  assign n7491 = n7479 & ~n7490;
  assign n7492 = n7479 & ~n7491;
  assign n7493 = ~n7490 & ~n7491;
  assign n7494 = ~n7492 & ~n7493;
  assign n7495 = ~n7085 & ~n7178;
  assign n7496 = ~n7175 & ~n7495;
  assign n7497 = n7494 & n7496;
  assign n7498 = ~n7494 & ~n7496;
  assign n7499 = ~n7497 & ~n7498;
  assign n7500 = n1696 & n3034;
  assign n7501 = pi81  & n3225;
  assign n7502 = pi83  & n3032;
  assign n7503 = pi82  & n3027;
  assign n7504 = ~n7502 & ~n7503;
  assign n7505 = ~n7501 & n7504;
  assign n7506 = ~n7500 & n7505;
  assign n7507 = pi29  & ~n7506;
  assign n7508 = pi29  & ~n7507;
  assign n7509 = ~n7506 & ~n7507;
  assign n7510 = ~n7508 & ~n7509;
  assign n7511 = n7499 & ~n7510;
  assign n7512 = n7499 & ~n7511;
  assign n7513 = ~n7510 & ~n7511;
  assign n7514 = ~n7512 & ~n7513;
  assign n7515 = ~n7193 & ~n7196;
  assign n7516 = n7514 & n7515;
  assign n7517 = ~n7514 & ~n7515;
  assign n7518 = ~n7516 & ~n7517;
  assign n7519 = n2133 & n2523;
  assign n7520 = pi84  & n2667;
  assign n7521 = pi86  & n2521;
  assign n7522 = pi85  & n2516;
  assign n7523 = ~n7521 & ~n7522;
  assign n7524 = ~n7520 & n7523;
  assign n7525 = ~n7519 & n7524;
  assign n7526 = pi26  & ~n7525;
  assign n7527 = pi26  & ~n7526;
  assign n7528 = ~n7525 & ~n7526;
  assign n7529 = ~n7527 & ~n7528;
  assign n7530 = n7518 & ~n7529;
  assign n7531 = n7518 & ~n7530;
  assign n7532 = ~n7529 & ~n7530;
  assign n7533 = ~n7531 & ~n7532;
  assign n7534 = ~n7210 & ~n7216;
  assign n7535 = n7533 & n7534;
  assign n7536 = ~n7533 & ~n7534;
  assign n7537 = ~n7535 & ~n7536;
  assign n7538 = n2043 & n2473;
  assign n7539 = pi87  & n2180;
  assign n7540 = pi89  & n2041;
  assign n7541 = pi88  & n2036;
  assign n7542 = ~n7540 & ~n7541;
  assign n7543 = ~n7539 & n7542;
  assign n7544 = ~n7538 & n7543;
  assign n7545 = pi23  & ~n7544;
  assign n7546 = pi23  & ~n7545;
  assign n7547 = ~n7544 & ~n7545;
  assign n7548 = ~n7546 & ~n7547;
  assign n7549 = n7537 & ~n7548;
  assign n7550 = n7537 & ~n7549;
  assign n7551 = ~n7548 & ~n7549;
  assign n7552 = ~n7550 & ~n7551;
  assign n7553 = ~n7230 & ~n7232;
  assign n7554 = ~n7552 & ~n7553;
  assign n7555 = n7552 & n7553;
  assign n7556 = ~n7554 & ~n7555;
  assign n7557 = ~n7381 & n7556;
  assign n7558 = ~n7381 & ~n7557;
  assign n7559 = n7556 & ~n7557;
  assign n7560 = ~n7558 & ~n7559;
  assign n7561 = ~n7370 & ~n7560;
  assign n7562 = ~n7370 & ~n7561;
  assign n7563 = ~n7560 & ~n7561;
  assign n7564 = ~n7562 & ~n7563;
  assign n7565 = n1297 & n3784;
  assign n7566 = pi93  & n1366;
  assign n7567 = pi95  & n1295;
  assign n7568 = pi94  & n1290;
  assign n7569 = ~n7567 & ~n7568;
  assign n7570 = ~n7566 & n7569;
  assign n7571 = ~n7565 & n7570;
  assign n7572 = pi17  & ~n7571;
  assign n7573 = pi17  & ~n7572;
  assign n7574 = ~n7571 & ~n7572;
  assign n7575 = ~n7573 & ~n7574;
  assign n7576 = n7564 & n7575;
  assign n7577 = ~n7564 & ~n7575;
  assign n7578 = ~n7576 & ~n7577;
  assign n7579 = ~n7368 & n7578;
  assign n7580 = n7368 & ~n7578;
  assign n7581 = ~n7579 & ~n7580;
  assign n7582 = n938 & n4454;
  assign n7583 = pi96  & n1052;
  assign n7584 = pi98  & n936;
  assign n7585 = pi97  & n931;
  assign n7586 = ~n7584 & ~n7585;
  assign n7587 = ~n7583 & n7586;
  assign n7588 = ~n7582 & n7587;
  assign n7589 = pi14  & ~n7588;
  assign n7590 = pi14  & ~n7589;
  assign n7591 = ~n7588 & ~n7589;
  assign n7592 = ~n7590 & ~n7591;
  assign n7593 = n7581 & ~n7592;
  assign n7594 = n7581 & ~n7593;
  assign n7595 = ~n7592 & ~n7593;
  assign n7596 = ~n7594 & ~n7595;
  assign n7597 = ~n7081 & ~n7284;
  assign n7598 = ~n7281 & ~n7597;
  assign n7599 = n7596 & n7598;
  assign n7600 = ~n7596 & ~n7598;
  assign n7601 = ~n7599 & ~n7600;
  assign n7602 = n687 & n5169;
  assign n7603 = pi99  & n763;
  assign n7604 = pi101  & n685;
  assign n7605 = pi100  & n680;
  assign n7606 = ~n7604 & ~n7605;
  assign n7607 = ~n7603 & n7606;
  assign n7608 = ~n7602 & n7607;
  assign n7609 = pi11  & ~n7608;
  assign n7610 = pi11  & ~n7609;
  assign n7611 = ~n7608 & ~n7609;
  assign n7612 = ~n7610 & ~n7611;
  assign n7613 = n7601 & ~n7612;
  assign n7614 = n7601 & ~n7613;
  assign n7615 = ~n7612 & ~n7613;
  assign n7616 = ~n7614 & ~n7615;
  assign n7617 = ~n7299 & ~n7303;
  assign n7618 = n7616 & n7617;
  assign n7619 = ~n7616 & ~n7617;
  assign n7620 = ~n7618 & ~n7619;
  assign n7621 = n498 & n5943;
  assign n7622 = pi102  & n537;
  assign n7623 = pi104  & n496;
  assign n7624 = pi103  & n491;
  assign n7625 = ~n7623 & ~n7624;
  assign n7626 = ~n7622 & n7625;
  assign n7627 = ~n7621 & n7626;
  assign n7628 = pi8  & ~n7627;
  assign n7629 = pi8  & ~n7628;
  assign n7630 = ~n7627 & ~n7628;
  assign n7631 = ~n7629 & ~n7630;
  assign n7632 = n7620 & ~n7631;
  assign n7633 = ~n7620 & n7631;
  assign n7634 = ~n7632 & ~n7633;
  assign n7635 = ~n7367 & n7634;
  assign n7636 = ~n7367 & ~n7635;
  assign n7637 = ~n7632 & ~n7635;
  assign n7638 = ~n7633 & n7637;
  assign n7639 = ~n7636 & ~n7638;
  assign n7640 = n342 & n6775;
  assign n7641 = pi105  & n380;
  assign n7642 = pi107  & n340;
  assign n7643 = pi106  & n335;
  assign n7644 = ~n7642 & ~n7643;
  assign n7645 = ~n7641 & n7644;
  assign n7646 = ~n7640 & n7645;
  assign n7647 = pi5  & ~n7646;
  assign n7648 = pi5  & ~n7647;
  assign n7649 = ~n7646 & ~n7647;
  assign n7650 = ~n7648 & ~n7649;
  assign n7651 = ~n7639 & ~n7650;
  assign n7652 = ~n7639 & ~n7651;
  assign n7653 = ~n7650 & ~n7651;
  assign n7654 = ~n7652 & ~n7653;
  assign n7655 = ~n7335 & ~n7341;
  assign n7656 = n7654 & n7655;
  assign n7657 = ~n7654 & ~n7655;
  assign n7658 = ~n7656 & ~n7657;
  assign n7659 = ~n7345 & ~n7347;
  assign n7660 = ~pi109  & ~pi110 ;
  assign n7661 = pi109  & pi110 ;
  assign n7662 = ~n7660 & ~n7661;
  assign n7663 = ~n7659 & n7662;
  assign n7664 = n7659 & ~n7662;
  assign n7665 = ~n7663 & ~n7664;
  assign n7666 = n262 & n7665;
  assign n7667 = pi108  & n288;
  assign n7668 = pi110  & n267;
  assign n7669 = pi109  & n269;
  assign n7670 = ~n7668 & ~n7669;
  assign n7671 = ~n7667 & n7670;
  assign n7672 = ~n7666 & n7671;
  assign n7673 = pi2  & ~n7672;
  assign n7674 = pi2  & ~n7673;
  assign n7675 = ~n7672 & ~n7673;
  assign n7676 = ~n7674 & ~n7675;
  assign n7677 = n7658 & ~n7676;
  assign n7678 = n7658 & ~n7677;
  assign n7679 = ~n7676 & ~n7677;
  assign n7680 = ~n7678 & ~n7679;
  assign n7681 = ~n7362 & ~n7364;
  assign n7682 = ~n7680 & ~n7681;
  assign n7683 = n7680 & n7681;
  assign po46  = ~n7682 & ~n7683;
  assign n7685 = ~n7651 & ~n7657;
  assign n7686 = ~n7577 & ~n7579;
  assign n7687 = n1297 & n4001;
  assign n7688 = pi94  & n1366;
  assign n7689 = pi96  & n1295;
  assign n7690 = pi95  & n1290;
  assign n7691 = ~n7689 & ~n7690;
  assign n7692 = ~n7688 & n7691;
  assign n7693 = ~n7687 & n7692;
  assign n7694 = pi17  & ~n7693;
  assign n7695 = pi17  & ~n7694;
  assign n7696 = ~n7693 & ~n7694;
  assign n7697 = ~n7695 & ~n7696;
  assign n7698 = ~n7557 & ~n7561;
  assign n7699 = n1611 & n3371;
  assign n7700 = pi91  & n1745;
  assign n7701 = pi93  & n1609;
  assign n7702 = pi92  & n1604;
  assign n7703 = ~n7701 & ~n7702;
  assign n7704 = ~n7700 & n7703;
  assign n7705 = ~n7699 & n7704;
  assign n7706 = pi20  & ~n7705;
  assign n7707 = pi20  & ~n7706;
  assign n7708 = ~n7705 & ~n7706;
  assign n7709 = ~n7707 & ~n7708;
  assign n7710 = ~n7549 & ~n7554;
  assign n7711 = ~n7530 & ~n7536;
  assign n7712 = ~n7491 & ~n7498;
  assign n7713 = n1434 & n3622;
  assign n7714 = pi79  & n3814;
  assign n7715 = pi81  & n3620;
  assign n7716 = pi80  & n3615;
  assign n7717 = ~n7715 & ~n7716;
  assign n7718 = ~n7714 & n7717;
  assign n7719 = ~n7713 & n7718;
  assign n7720 = pi32  & ~n7719;
  assign n7721 = pi32  & ~n7720;
  assign n7722 = ~n7719 & ~n7720;
  assign n7723 = ~n7721 & ~n7722;
  assign n7724 = ~n7475 & ~n7477;
  assign n7725 = ~n7436 & ~n7442;
  assign n7726 = n576 & n5739;
  assign n7727 = pi70  & n6030;
  assign n7728 = pi72  & n5737;
  assign n7729 = pi71  & n5732;
  assign n7730 = ~n7728 & ~n7729;
  assign n7731 = ~n7727 & n7730;
  assign n7732 = ~n7726 & n7731;
  assign n7733 = pi41  & ~n7732;
  assign n7734 = pi41  & ~n7733;
  assign n7735 = ~n7732 & ~n7733;
  assign n7736 = ~n7734 & ~n7735;
  assign n7737 = ~n7420 & ~n7422;
  assign n7738 = n286 & n7408;
  assign n7739 = n7101 & n7400;
  assign n7740 = ~n7405 & n7739;
  assign n7741 = pi64  & n7740;
  assign n7742 = pi66  & n7406;
  assign n7743 = pi65  & n7401;
  assign n7744 = ~n7742 & ~n7743;
  assign n7745 = ~n7738 & n7744;
  assign n7746 = ~n7741 & n7745;
  assign n7747 = pi47  & ~n7746;
  assign n7748 = pi47  & ~n7747;
  assign n7749 = ~n7746 & ~n7747;
  assign n7750 = ~n7748 & ~n7749;
  assign n7751 = ~n7416 & n7750;
  assign n7752 = n7416 & ~n7750;
  assign n7753 = ~n7751 & ~n7752;
  assign n7754 = n401 & n6539;
  assign n7755 = pi67  & n6873;
  assign n7756 = pi69  & n6537;
  assign n7757 = pi68  & n6532;
  assign n7758 = ~n7756 & ~n7757;
  assign n7759 = ~n7755 & n7758;
  assign n7760 = ~n7754 & n7759;
  assign n7761 = pi44  & ~n7760;
  assign n7762 = pi44  & ~n7761;
  assign n7763 = ~n7760 & ~n7761;
  assign n7764 = ~n7762 & ~n7763;
  assign n7765 = n7753 & ~n7764;
  assign n7766 = n7753 & ~n7765;
  assign n7767 = ~n7764 & ~n7765;
  assign n7768 = ~n7766 & ~n7767;
  assign n7769 = ~n7737 & ~n7768;
  assign n7770 = n7737 & n7768;
  assign n7771 = ~n7769 & ~n7770;
  assign n7772 = ~n7736 & n7771;
  assign n7773 = ~n7736 & ~n7772;
  assign n7774 = n7771 & ~n7772;
  assign n7775 = ~n7773 & ~n7774;
  assign n7776 = ~n7725 & ~n7775;
  assign n7777 = ~n7725 & ~n7776;
  assign n7778 = ~n7775 & ~n7776;
  assign n7779 = ~n7777 & ~n7778;
  assign n7780 = n809 & n5008;
  assign n7781 = pi73  & n5241;
  assign n7782 = pi75  & n5006;
  assign n7783 = pi74  & n5001;
  assign n7784 = ~n7782 & ~n7783;
  assign n7785 = ~n7781 & n7784;
  assign n7786 = ~n7780 & n7785;
  assign n7787 = pi38  & ~n7786;
  assign n7788 = pi38  & ~n7787;
  assign n7789 = ~n7786 & ~n7787;
  assign n7790 = ~n7788 & ~n7789;
  assign n7791 = n7779 & n7790;
  assign n7792 = ~n7779 & ~n7790;
  assign n7793 = ~n7791 & ~n7792;
  assign n7794 = ~n7460 & n7793;
  assign n7795 = n7460 & ~n7793;
  assign n7796 = ~n7794 & ~n7795;
  assign n7797 = n1025 & n4271;
  assign n7798 = pi76  & n4503;
  assign n7799 = pi78  & n4269;
  assign n7800 = pi77  & n4264;
  assign n7801 = ~n7799 & ~n7800;
  assign n7802 = ~n7798 & n7801;
  assign n7803 = ~n7797 & n7802;
  assign n7804 = pi35  & ~n7803;
  assign n7805 = pi35  & ~n7804;
  assign n7806 = ~n7803 & ~n7804;
  assign n7807 = ~n7805 & ~n7806;
  assign n7808 = n7796 & ~n7807;
  assign n7809 = n7796 & ~n7808;
  assign n7810 = ~n7807 & ~n7808;
  assign n7811 = ~n7809 & ~n7810;
  assign n7812 = ~n7724 & ~n7811;
  assign n7813 = n7724 & n7811;
  assign n7814 = ~n7812 & ~n7813;
  assign n7815 = ~n7723 & n7814;
  assign n7816 = ~n7723 & ~n7815;
  assign n7817 = n7814 & ~n7815;
  assign n7818 = ~n7816 & ~n7817;
  assign n7819 = ~n7712 & ~n7818;
  assign n7820 = ~n7712 & ~n7819;
  assign n7821 = ~n7818 & ~n7819;
  assign n7822 = ~n7820 & ~n7821;
  assign n7823 = n1834 & n3034;
  assign n7824 = pi82  & n3225;
  assign n7825 = pi84  & n3032;
  assign n7826 = pi83  & n3027;
  assign n7827 = ~n7825 & ~n7826;
  assign n7828 = ~n7824 & n7827;
  assign n7829 = ~n7823 & n7828;
  assign n7830 = pi29  & ~n7829;
  assign n7831 = pi29  & ~n7830;
  assign n7832 = ~n7829 & ~n7830;
  assign n7833 = ~n7831 & ~n7832;
  assign n7834 = ~n7822 & ~n7833;
  assign n7835 = ~n7822 & ~n7834;
  assign n7836 = ~n7833 & ~n7834;
  assign n7837 = ~n7835 & ~n7836;
  assign n7838 = ~n7511 & ~n7517;
  assign n7839 = n7837 & n7838;
  assign n7840 = ~n7837 & ~n7838;
  assign n7841 = ~n7839 & ~n7840;
  assign n7842 = n2288 & n2523;
  assign n7843 = pi85  & n2667;
  assign n7844 = pi87  & n2521;
  assign n7845 = pi86  & n2516;
  assign n7846 = ~n7844 & ~n7845;
  assign n7847 = ~n7843 & n7846;
  assign n7848 = ~n7842 & n7847;
  assign n7849 = pi26  & ~n7848;
  assign n7850 = pi26  & ~n7849;
  assign n7851 = ~n7848 & ~n7849;
  assign n7852 = ~n7850 & ~n7851;
  assign n7853 = n7841 & ~n7852;
  assign n7854 = ~n7841 & n7852;
  assign n7855 = ~n7853 & ~n7854;
  assign n7856 = ~n7711 & n7855;
  assign n7857 = ~n7711 & ~n7856;
  assign n7858 = ~n7853 & ~n7856;
  assign n7859 = ~n7854 & n7858;
  assign n7860 = ~n7857 & ~n7859;
  assign n7861 = n2043 & n2801;
  assign n7862 = pi88  & n2180;
  assign n7863 = pi90  & n2041;
  assign n7864 = pi89  & n2036;
  assign n7865 = ~n7863 & ~n7864;
  assign n7866 = ~n7862 & n7865;
  assign n7867 = ~n7861 & n7866;
  assign n7868 = pi23  & ~n7867;
  assign n7869 = pi23  & ~n7868;
  assign n7870 = ~n7867 & ~n7868;
  assign n7871 = ~n7869 & ~n7870;
  assign n7872 = n7860 & n7871;
  assign n7873 = ~n7860 & ~n7871;
  assign n7874 = ~n7872 & ~n7873;
  assign n7875 = ~n7710 & n7874;
  assign n7876 = n7710 & ~n7874;
  assign n7877 = ~n7875 & ~n7876;
  assign n7878 = n7709 & ~n7877;
  assign n7879 = ~n7709 & n7877;
  assign n7880 = ~n7878 & ~n7879;
  assign n7881 = ~n7698 & n7880;
  assign n7882 = n7698 & ~n7880;
  assign n7883 = ~n7881 & ~n7882;
  assign n7884 = n7697 & ~n7883;
  assign n7885 = ~n7697 & n7883;
  assign n7886 = ~n7884 & ~n7885;
  assign n7887 = ~n7686 & n7886;
  assign n7888 = n7686 & ~n7886;
  assign n7889 = ~n7887 & ~n7888;
  assign n7890 = n938 & n4684;
  assign n7891 = pi97  & n1052;
  assign n7892 = pi99  & n936;
  assign n7893 = pi98  & n931;
  assign n7894 = ~n7892 & ~n7893;
  assign n7895 = ~n7891 & n7894;
  assign n7896 = ~n7890 & n7895;
  assign n7897 = pi14  & ~n7896;
  assign n7898 = pi14  & ~n7897;
  assign n7899 = ~n7896 & ~n7897;
  assign n7900 = ~n7898 & ~n7899;
  assign n7901 = n7889 & ~n7900;
  assign n7902 = n7889 & ~n7901;
  assign n7903 = ~n7900 & ~n7901;
  assign n7904 = ~n7902 & ~n7903;
  assign n7905 = ~n7593 & ~n7600;
  assign n7906 = n7904 & n7905;
  assign n7907 = ~n7904 & ~n7905;
  assign n7908 = ~n7906 & ~n7907;
  assign n7909 = n687 & n5413;
  assign n7910 = pi100  & n763;
  assign n7911 = pi102  & n685;
  assign n7912 = pi101  & n680;
  assign n7913 = ~n7911 & ~n7912;
  assign n7914 = ~n7910 & n7913;
  assign n7915 = ~n7909 & n7914;
  assign n7916 = pi11  & ~n7915;
  assign n7917 = pi11  & ~n7916;
  assign n7918 = ~n7915 & ~n7916;
  assign n7919 = ~n7917 & ~n7918;
  assign n7920 = n7908 & ~n7919;
  assign n7921 = n7908 & ~n7920;
  assign n7922 = ~n7919 & ~n7920;
  assign n7923 = ~n7921 & ~n7922;
  assign n7924 = ~n7613 & ~n7619;
  assign n7925 = n7923 & n7924;
  assign n7926 = ~n7923 & ~n7924;
  assign n7927 = ~n7925 & ~n7926;
  assign n7928 = n498 & n6207;
  assign n7929 = pi103  & n537;
  assign n7930 = pi105  & n496;
  assign n7931 = pi104  & n491;
  assign n7932 = ~n7930 & ~n7931;
  assign n7933 = ~n7929 & n7932;
  assign n7934 = ~n7928 & n7933;
  assign n7935 = pi8  & ~n7934;
  assign n7936 = pi8  & ~n7935;
  assign n7937 = ~n7934 & ~n7935;
  assign n7938 = ~n7936 & ~n7937;
  assign n7939 = n7927 & ~n7938;
  assign n7940 = ~n7927 & n7938;
  assign n7941 = ~n7939 & ~n7940;
  assign n7942 = ~n7637 & n7941;
  assign n7943 = ~n7637 & ~n7942;
  assign n7944 = ~n7939 & ~n7942;
  assign n7945 = ~n7940 & n7944;
  assign n7946 = ~n7943 & ~n7945;
  assign n7947 = n342 & n7060;
  assign n7948 = pi106  & n380;
  assign n7949 = pi108  & n340;
  assign n7950 = pi107  & n335;
  assign n7951 = ~n7949 & ~n7950;
  assign n7952 = ~n7948 & n7951;
  assign n7953 = ~n7947 & n7952;
  assign n7954 = pi5  & ~n7953;
  assign n7955 = pi5  & ~n7954;
  assign n7956 = ~n7953 & ~n7954;
  assign n7957 = ~n7955 & ~n7956;
  assign n7958 = n7946 & n7957;
  assign n7959 = ~n7946 & ~n7957;
  assign n7960 = ~n7958 & ~n7959;
  assign n7961 = ~n7685 & n7960;
  assign n7962 = n7685 & ~n7960;
  assign n7963 = ~n7961 & ~n7962;
  assign n7964 = ~n7661 & ~n7663;
  assign n7965 = ~pi110  & ~pi111 ;
  assign n7966 = pi110  & pi111 ;
  assign n7967 = ~n7965 & ~n7966;
  assign n7968 = ~n7964 & n7967;
  assign n7969 = n7964 & ~n7967;
  assign n7970 = ~n7968 & ~n7969;
  assign n7971 = n262 & n7970;
  assign n7972 = pi109  & n288;
  assign n7973 = pi111  & n267;
  assign n7974 = pi110  & n269;
  assign n7975 = ~n7973 & ~n7974;
  assign n7976 = ~n7972 & n7975;
  assign n7977 = ~n7971 & n7976;
  assign n7978 = pi2  & ~n7977;
  assign n7979 = pi2  & ~n7978;
  assign n7980 = ~n7977 & ~n7978;
  assign n7981 = ~n7979 & ~n7980;
  assign n7982 = n7963 & ~n7981;
  assign n7983 = n7963 & ~n7982;
  assign n7984 = ~n7981 & ~n7982;
  assign n7985 = ~n7983 & ~n7984;
  assign n7986 = ~n7677 & ~n7682;
  assign n7987 = ~n7985 & ~n7986;
  assign n7988 = n7985 & n7986;
  assign po47  = ~n7987 & ~n7988;
  assign n7990 = ~n7982 & ~n7987;
  assign n7991 = ~n7966 & ~n7968;
  assign n7992 = ~pi111  & ~pi112 ;
  assign n7993 = pi111  & pi112 ;
  assign n7994 = ~n7992 & ~n7993;
  assign n7995 = ~n7991 & n7994;
  assign n7996 = n7991 & ~n7994;
  assign n7997 = ~n7995 & ~n7996;
  assign n7998 = n262 & n7997;
  assign n7999 = pi110  & n288;
  assign n8000 = pi112  & n267;
  assign n8001 = pi111  & n269;
  assign n8002 = ~n8000 & ~n8001;
  assign n8003 = ~n7999 & n8002;
  assign n8004 = ~n7998 & n8003;
  assign n8005 = pi2  & ~n8004;
  assign n8006 = pi2  & ~n8005;
  assign n8007 = ~n8004 & ~n8005;
  assign n8008 = ~n8006 & ~n8007;
  assign n8009 = ~n7959 & ~n7961;
  assign n8010 = ~n7901 & ~n7907;
  assign n8011 = ~n7885 & ~n7887;
  assign n8012 = ~n7879 & ~n7881;
  assign n8013 = ~n7873 & ~n7875;
  assign n8014 = ~n7808 & ~n7812;
  assign n8015 = n1122 & n4271;
  assign n8016 = pi77  & n4503;
  assign n8017 = pi79  & n4269;
  assign n8018 = pi78  & n4264;
  assign n8019 = ~n8017 & ~n8018;
  assign n8020 = ~n8016 & n8019;
  assign n8021 = ~n8015 & n8020;
  assign n8022 = pi35  & ~n8021;
  assign n8023 = pi35  & ~n8022;
  assign n8024 = ~n8021 & ~n8022;
  assign n8025 = ~n8023 & ~n8024;
  assign n8026 = ~n7792 & ~n7794;
  assign n8027 = n891 & n5008;
  assign n8028 = pi74  & n5241;
  assign n8029 = pi76  & n5006;
  assign n8030 = pi75  & n5001;
  assign n8031 = ~n8029 & ~n8030;
  assign n8032 = ~n8028 & n8031;
  assign n8033 = ~n8027 & n8032;
  assign n8034 = pi38  & ~n8033;
  assign n8035 = pi38  & ~n8034;
  assign n8036 = ~n8033 & ~n8034;
  assign n8037 = ~n8035 & ~n8036;
  assign n8038 = ~n7772 & ~n7776;
  assign n8039 = pi47  & ~pi48 ;
  assign n8040 = ~pi47  & pi48 ;
  assign n8041 = ~n8039 & ~n8040;
  assign n8042 = pi64  & ~n8041;
  assign n8043 = ~n7752 & n8042;
  assign n8044 = n7752 & ~n8042;
  assign n8045 = ~n8043 & ~n8044;
  assign n8046 = n309 & n7408;
  assign n8047 = pi65  & n7740;
  assign n8048 = pi67  & n7406;
  assign n8049 = pi66  & n7401;
  assign n8050 = ~n8048 & ~n8049;
  assign n8051 = ~n8047 & n8050;
  assign n8052 = ~n8046 & n8051;
  assign n8053 = pi47  & ~n8052;
  assign n8054 = pi47  & ~n8053;
  assign n8055 = ~n8052 & ~n8053;
  assign n8056 = ~n8054 & ~n8055;
  assign n8057 = ~n8045 & ~n8056;
  assign n8058 = n8045 & n8056;
  assign n8059 = ~n8057 & ~n8058;
  assign n8060 = n450 & n6539;
  assign n8061 = pi68  & n6873;
  assign n8062 = pi70  & n6537;
  assign n8063 = pi69  & n6532;
  assign n8064 = ~n8062 & ~n8063;
  assign n8065 = ~n8061 & n8064;
  assign n8066 = ~n8060 & n8065;
  assign n8067 = pi44  & ~n8066;
  assign n8068 = pi44  & ~n8067;
  assign n8069 = ~n8066 & ~n8067;
  assign n8070 = ~n8068 & ~n8069;
  assign n8071 = n8059 & ~n8070;
  assign n8072 = n8059 & ~n8071;
  assign n8073 = ~n8070 & ~n8071;
  assign n8074 = ~n8072 & ~n8073;
  assign n8075 = ~n7765 & ~n7769;
  assign n8076 = n8074 & n8075;
  assign n8077 = ~n8074 & ~n8075;
  assign n8078 = ~n8076 & ~n8077;
  assign n8079 = n642 & n5739;
  assign n8080 = pi71  & n6030;
  assign n8081 = pi73  & n5737;
  assign n8082 = pi72  & n5732;
  assign n8083 = ~n8081 & ~n8082;
  assign n8084 = ~n8080 & n8083;
  assign n8085 = ~n8079 & n8084;
  assign n8086 = pi41  & ~n8085;
  assign n8087 = pi41  & ~n8086;
  assign n8088 = ~n8085 & ~n8086;
  assign n8089 = ~n8087 & ~n8088;
  assign n8090 = ~n8078 & n8089;
  assign n8091 = n8078 & ~n8089;
  assign n8092 = ~n8090 & ~n8091;
  assign n8093 = ~n8038 & n8092;
  assign n8094 = n8038 & ~n8092;
  assign n8095 = ~n8093 & ~n8094;
  assign n8096 = ~n8037 & n8095;
  assign n8097 = ~n8037 & ~n8096;
  assign n8098 = n8095 & ~n8096;
  assign n8099 = ~n8097 & ~n8098;
  assign n8100 = ~n8026 & ~n8099;
  assign n8101 = n8026 & n8099;
  assign n8102 = ~n8100 & ~n8101;
  assign n8103 = ~n8025 & n8102;
  assign n8104 = n8025 & ~n8102;
  assign n8105 = ~n8103 & ~n8104;
  assign n8106 = ~n8014 & n8105;
  assign n8107 = n8014 & ~n8105;
  assign n8108 = ~n8106 & ~n8107;
  assign n8109 = n1554 & n3622;
  assign n8110 = pi80  & n3814;
  assign n8111 = pi82  & n3620;
  assign n8112 = pi81  & n3615;
  assign n8113 = ~n8111 & ~n8112;
  assign n8114 = ~n8110 & n8113;
  assign n8115 = ~n8109 & n8114;
  assign n8116 = pi32  & ~n8115;
  assign n8117 = pi32  & ~n8116;
  assign n8118 = ~n8115 & ~n8116;
  assign n8119 = ~n8117 & ~n8118;
  assign n8120 = n8108 & ~n8119;
  assign n8121 = n8108 & ~n8120;
  assign n8122 = ~n8119 & ~n8120;
  assign n8123 = ~n8121 & ~n8122;
  assign n8124 = ~n7815 & ~n7819;
  assign n8125 = n8123 & n8124;
  assign n8126 = ~n8123 & ~n8124;
  assign n8127 = ~n8125 & ~n8126;
  assign n8128 = n1972 & n3034;
  assign n8129 = pi83  & n3225;
  assign n8130 = pi85  & n3032;
  assign n8131 = pi84  & n3027;
  assign n8132 = ~n8130 & ~n8131;
  assign n8133 = ~n8129 & n8132;
  assign n8134 = ~n8128 & n8133;
  assign n8135 = pi29  & ~n8134;
  assign n8136 = pi29  & ~n8135;
  assign n8137 = ~n8134 & ~n8135;
  assign n8138 = ~n8136 & ~n8137;
  assign n8139 = n8127 & ~n8138;
  assign n8140 = n8127 & ~n8139;
  assign n8141 = ~n8138 & ~n8139;
  assign n8142 = ~n8140 & ~n8141;
  assign n8143 = ~n7834 & ~n7840;
  assign n8144 = n8142 & n8143;
  assign n8145 = ~n8142 & ~n8143;
  assign n8146 = ~n8144 & ~n8145;
  assign n8147 = n2446 & n2523;
  assign n8148 = pi86  & n2667;
  assign n8149 = pi88  & n2521;
  assign n8150 = pi87  & n2516;
  assign n8151 = ~n8149 & ~n8150;
  assign n8152 = ~n8148 & n8151;
  assign n8153 = ~n8147 & n8152;
  assign n8154 = pi26  & ~n8153;
  assign n8155 = pi26  & ~n8154;
  assign n8156 = ~n8153 & ~n8154;
  assign n8157 = ~n8155 & ~n8156;
  assign n8158 = ~n8146 & n8157;
  assign n8159 = n8146 & ~n8157;
  assign n8160 = ~n8158 & ~n8159;
  assign n8161 = ~n7858 & n8160;
  assign n8162 = n7858 & ~n8160;
  assign n8163 = ~n8161 & ~n8162;
  assign n8164 = n2043 & n2978;
  assign n8165 = pi89  & n2180;
  assign n8166 = pi91  & n2041;
  assign n8167 = pi90  & n2036;
  assign n8168 = ~n8166 & ~n8167;
  assign n8169 = ~n8165 & n8168;
  assign n8170 = ~n8164 & n8169;
  assign n8171 = pi23  & ~n8170;
  assign n8172 = pi23  & ~n8171;
  assign n8173 = ~n8170 & ~n8171;
  assign n8174 = ~n8172 & ~n8173;
  assign n8175 = n8163 & ~n8174;
  assign n8176 = n8163 & ~n8175;
  assign n8177 = ~n8174 & ~n8175;
  assign n8178 = ~n8176 & ~n8177;
  assign n8179 = ~n8013 & n8178;
  assign n8180 = n8013 & ~n8178;
  assign n8181 = ~n8179 & ~n8180;
  assign n8182 = n1611 & n3565;
  assign n8183 = pi92  & n1745;
  assign n8184 = pi94  & n1609;
  assign n8185 = pi93  & n1604;
  assign n8186 = ~n8184 & ~n8185;
  assign n8187 = ~n8183 & n8186;
  assign n8188 = ~n8182 & n8187;
  assign n8189 = pi20  & ~n8188;
  assign n8190 = pi20  & ~n8189;
  assign n8191 = ~n8188 & ~n8189;
  assign n8192 = ~n8190 & ~n8191;
  assign n8193 = ~n8181 & ~n8192;
  assign n8194 = n8181 & n8192;
  assign n8195 = ~n8193 & ~n8194;
  assign n8196 = ~n8012 & n8195;
  assign n8197 = n8012 & ~n8195;
  assign n8198 = ~n8196 & ~n8197;
  assign n8199 = n1297 & n4211;
  assign n8200 = pi95  & n1366;
  assign n8201 = pi97  & n1295;
  assign n8202 = pi96  & n1290;
  assign n8203 = ~n8201 & ~n8202;
  assign n8204 = ~n8200 & n8203;
  assign n8205 = ~n8199 & n8204;
  assign n8206 = pi17  & ~n8205;
  assign n8207 = pi17  & ~n8206;
  assign n8208 = ~n8205 & ~n8206;
  assign n8209 = ~n8207 & ~n8208;
  assign n8210 = n8198 & ~n8209;
  assign n8211 = n8198 & ~n8210;
  assign n8212 = ~n8209 & ~n8210;
  assign n8213 = ~n8211 & ~n8212;
  assign n8214 = ~n8011 & n8213;
  assign n8215 = n8011 & ~n8213;
  assign n8216 = ~n8214 & ~n8215;
  assign n8217 = n938 & n4910;
  assign n8218 = pi98  & n1052;
  assign n8219 = pi100  & n936;
  assign n8220 = pi99  & n931;
  assign n8221 = ~n8219 & ~n8220;
  assign n8222 = ~n8218 & n8221;
  assign n8223 = ~n8217 & n8222;
  assign n8224 = pi14  & ~n8223;
  assign n8225 = pi14  & ~n8224;
  assign n8226 = ~n8223 & ~n8224;
  assign n8227 = ~n8225 & ~n8226;
  assign n8228 = ~n8216 & ~n8227;
  assign n8229 = n8216 & n8227;
  assign n8230 = ~n8228 & ~n8229;
  assign n8231 = n8010 & ~n8230;
  assign n8232 = ~n8010 & n8230;
  assign n8233 = ~n8231 & ~n8232;
  assign n8234 = n687 & n5664;
  assign n8235 = pi101  & n763;
  assign n8236 = pi103  & n685;
  assign n8237 = pi102  & n680;
  assign n8238 = ~n8236 & ~n8237;
  assign n8239 = ~n8235 & n8238;
  assign n8240 = ~n8234 & n8239;
  assign n8241 = pi11  & ~n8240;
  assign n8242 = pi11  & ~n8241;
  assign n8243 = ~n8240 & ~n8241;
  assign n8244 = ~n8242 & ~n8243;
  assign n8245 = n8233 & ~n8244;
  assign n8246 = n8233 & ~n8245;
  assign n8247 = ~n8244 & ~n8245;
  assign n8248 = ~n8246 & ~n8247;
  assign n8249 = ~n7920 & ~n7926;
  assign n8250 = n8248 & n8249;
  assign n8251 = ~n8248 & ~n8249;
  assign n8252 = ~n8250 & ~n8251;
  assign n8253 = n498 & n6477;
  assign n8254 = pi104  & n537;
  assign n8255 = pi106  & n496;
  assign n8256 = pi105  & n491;
  assign n8257 = ~n8255 & ~n8256;
  assign n8258 = ~n8254 & n8257;
  assign n8259 = ~n8253 & n8258;
  assign n8260 = pi8  & ~n8259;
  assign n8261 = pi8  & ~n8260;
  assign n8262 = ~n8259 & ~n8260;
  assign n8263 = ~n8261 & ~n8262;
  assign n8264 = n8252 & ~n8263;
  assign n8265 = n8252 & ~n8264;
  assign n8266 = ~n8263 & ~n8264;
  assign n8267 = ~n8265 & ~n8266;
  assign n8268 = ~n7944 & n8267;
  assign n8269 = n7944 & ~n8267;
  assign n8270 = ~n8268 & ~n8269;
  assign n8271 = n342 & n7349;
  assign n8272 = pi107  & n380;
  assign n8273 = pi109  & n340;
  assign n8274 = pi108  & n335;
  assign n8275 = ~n8273 & ~n8274;
  assign n8276 = ~n8272 & n8275;
  assign n8277 = ~n8271 & n8276;
  assign n8278 = pi5  & ~n8277;
  assign n8279 = pi5  & ~n8278;
  assign n8280 = ~n8277 & ~n8278;
  assign n8281 = ~n8279 & ~n8280;
  assign n8282 = ~n8270 & ~n8281;
  assign n8283 = n8270 & n8281;
  assign n8284 = ~n8282 & ~n8283;
  assign n8285 = ~n8009 & n8284;
  assign n8286 = n8009 & ~n8284;
  assign n8287 = ~n8285 & ~n8286;
  assign n8288 = n8008 & ~n8287;
  assign n8289 = ~n8008 & n8287;
  assign n8290 = ~n8288 & ~n8289;
  assign n8291 = ~n7990 & n8290;
  assign n8292 = n7990 & ~n8290;
  assign po48  = ~n8291 & ~n8292;
  assign n8294 = ~n8289 & ~n8291;
  assign n8295 = ~n8013 & ~n8178;
  assign n8296 = ~n8175 & ~n8295;
  assign n8297 = n2043 & n3177;
  assign n8298 = pi90  & n2180;
  assign n8299 = pi92  & n2041;
  assign n8300 = pi91  & n2036;
  assign n8301 = ~n8299 & ~n8300;
  assign n8302 = ~n8298 & n8301;
  assign n8303 = ~n8297 & n8302;
  assign n8304 = pi23  & ~n8303;
  assign n8305 = pi23  & ~n8304;
  assign n8306 = ~n8303 & ~n8304;
  assign n8307 = ~n8305 & ~n8306;
  assign n8308 = ~n8096 & ~n8100;
  assign n8309 = ~n8091 & ~n8093;
  assign n8310 = n7752 & n8042;
  assign n8311 = ~n8057 & ~n8310;
  assign n8312 = n359 & n7408;
  assign n8313 = pi66  & n7740;
  assign n8314 = pi68  & n7406;
  assign n8315 = pi67  & n7401;
  assign n8316 = ~n8314 & ~n8315;
  assign n8317 = ~n8313 & n8316;
  assign n8318 = ~n8312 & n8317;
  assign n8319 = pi47  & ~n8318;
  assign n8320 = pi47  & ~n8319;
  assign n8321 = ~n8318 & ~n8319;
  assign n8322 = ~n8320 & ~n8321;
  assign n8323 = pi50  & ~n8042;
  assign n8324 = ~pi48  & pi49 ;
  assign n8325 = pi48  & ~pi49 ;
  assign n8326 = ~n8324 & ~n8325;
  assign n8327 = n8041 & ~n8326;
  assign n8328 = pi64  & n8327;
  assign n8329 = ~pi49  & pi50 ;
  assign n8330 = pi49  & ~pi50 ;
  assign n8331 = ~n8329 & ~n8330;
  assign n8332 = ~n8041 & n8331;
  assign n8333 = pi65  & n8332;
  assign n8334 = ~n8041 & ~n8331;
  assign n8335 = ~n265 & n8334;
  assign n8336 = ~n8328 & ~n8333;
  assign n8337 = ~n8335 & n8336;
  assign n8338 = pi50  & ~n8337;
  assign n8339 = pi50  & ~n8338;
  assign n8340 = ~n8337 & ~n8338;
  assign n8341 = ~n8339 & ~n8340;
  assign n8342 = n8323 & ~n8341;
  assign n8343 = ~n8323 & n8341;
  assign n8344 = ~n8342 & ~n8343;
  assign n8345 = n8322 & ~n8344;
  assign n8346 = ~n8322 & n8344;
  assign n8347 = ~n8345 & ~n8346;
  assign n8348 = ~n8311 & n8347;
  assign n8349 = n8311 & ~n8347;
  assign n8350 = ~n8348 & ~n8349;
  assign n8351 = n475 & n6539;
  assign n8352 = pi69  & n6873;
  assign n8353 = pi71  & n6537;
  assign n8354 = pi70  & n6532;
  assign n8355 = ~n8353 & ~n8354;
  assign n8356 = ~n8352 & n8355;
  assign n8357 = ~n8351 & n8356;
  assign n8358 = pi44  & ~n8357;
  assign n8359 = pi44  & ~n8358;
  assign n8360 = ~n8357 & ~n8358;
  assign n8361 = ~n8359 & ~n8360;
  assign n8362 = n8350 & ~n8361;
  assign n8363 = n8350 & ~n8362;
  assign n8364 = ~n8361 & ~n8362;
  assign n8365 = ~n8363 & ~n8364;
  assign n8366 = ~n8071 & ~n8077;
  assign n8367 = n8365 & n8366;
  assign n8368 = ~n8365 & ~n8366;
  assign n8369 = ~n8367 & ~n8368;
  assign n8370 = n729 & n5739;
  assign n8371 = pi72  & n6030;
  assign n8372 = pi74  & n5737;
  assign n8373 = pi73  & n5732;
  assign n8374 = ~n8372 & ~n8373;
  assign n8375 = ~n8371 & n8374;
  assign n8376 = ~n8370 & n8375;
  assign n8377 = pi41  & ~n8376;
  assign n8378 = pi41  & ~n8377;
  assign n8379 = ~n8376 & ~n8377;
  assign n8380 = ~n8378 & ~n8379;
  assign n8381 = n8369 & ~n8380;
  assign n8382 = ~n8369 & n8380;
  assign n8383 = ~n8381 & ~n8382;
  assign n8384 = ~n8309 & n8383;
  assign n8385 = ~n8309 & ~n8384;
  assign n8386 = ~n8381 & ~n8384;
  assign n8387 = ~n8382 & n8386;
  assign n8388 = ~n8385 & ~n8387;
  assign n8389 = n999 & n5008;
  assign n8390 = pi75  & n5241;
  assign n8391 = pi77  & n5006;
  assign n8392 = pi76  & n5001;
  assign n8393 = ~n8391 & ~n8392;
  assign n8394 = ~n8390 & n8393;
  assign n8395 = ~n8389 & n8394;
  assign n8396 = pi38  & ~n8395;
  assign n8397 = pi38  & ~n8396;
  assign n8398 = ~n8395 & ~n8396;
  assign n8399 = ~n8397 & ~n8398;
  assign n8400 = n8388 & n8399;
  assign n8401 = ~n8388 & ~n8399;
  assign n8402 = ~n8400 & ~n8401;
  assign n8403 = ~n8308 & n8402;
  assign n8404 = n8308 & ~n8402;
  assign n8405 = ~n8403 & ~n8404;
  assign n8406 = n1225 & n4271;
  assign n8407 = pi78  & n4503;
  assign n8408 = pi80  & n4269;
  assign n8409 = pi79  & n4264;
  assign n8410 = ~n8408 & ~n8409;
  assign n8411 = ~n8407 & n8410;
  assign n8412 = ~n8406 & n8411;
  assign n8413 = pi35  & ~n8412;
  assign n8414 = pi35  & ~n8413;
  assign n8415 = ~n8412 & ~n8413;
  assign n8416 = ~n8414 & ~n8415;
  assign n8417 = n8405 & ~n8416;
  assign n8418 = n8405 & ~n8417;
  assign n8419 = ~n8416 & ~n8417;
  assign n8420 = ~n8418 & ~n8419;
  assign n8421 = ~n8103 & ~n8106;
  assign n8422 = n8420 & n8421;
  assign n8423 = ~n8420 & ~n8421;
  assign n8424 = ~n8422 & ~n8423;
  assign n8425 = n1696 & n3622;
  assign n8426 = pi81  & n3814;
  assign n8427 = pi83  & n3620;
  assign n8428 = pi82  & n3615;
  assign n8429 = ~n8427 & ~n8428;
  assign n8430 = ~n8426 & n8429;
  assign n8431 = ~n8425 & n8430;
  assign n8432 = pi32  & ~n8431;
  assign n8433 = pi32  & ~n8432;
  assign n8434 = ~n8431 & ~n8432;
  assign n8435 = ~n8433 & ~n8434;
  assign n8436 = n8424 & ~n8435;
  assign n8437 = n8424 & ~n8436;
  assign n8438 = ~n8435 & ~n8436;
  assign n8439 = ~n8437 & ~n8438;
  assign n8440 = ~n8120 & ~n8126;
  assign n8441 = n8439 & n8440;
  assign n8442 = ~n8439 & ~n8440;
  assign n8443 = ~n8441 & ~n8442;
  assign n8444 = n2133 & n3034;
  assign n8445 = pi84  & n3225;
  assign n8446 = pi86  & n3032;
  assign n8447 = pi85  & n3027;
  assign n8448 = ~n8446 & ~n8447;
  assign n8449 = ~n8445 & n8448;
  assign n8450 = ~n8444 & n8449;
  assign n8451 = pi29  & ~n8450;
  assign n8452 = pi29  & ~n8451;
  assign n8453 = ~n8450 & ~n8451;
  assign n8454 = ~n8452 & ~n8453;
  assign n8455 = n8443 & ~n8454;
  assign n8456 = n8443 & ~n8455;
  assign n8457 = ~n8454 & ~n8455;
  assign n8458 = ~n8456 & ~n8457;
  assign n8459 = ~n8139 & ~n8145;
  assign n8460 = n8458 & n8459;
  assign n8461 = ~n8458 & ~n8459;
  assign n8462 = ~n8460 & ~n8461;
  assign n8463 = n2473 & n2523;
  assign n8464 = pi87  & n2667;
  assign n8465 = pi89  & n2521;
  assign n8466 = pi88  & n2516;
  assign n8467 = ~n8465 & ~n8466;
  assign n8468 = ~n8464 & n8467;
  assign n8469 = ~n8463 & n8468;
  assign n8470 = pi26  & ~n8469;
  assign n8471 = pi26  & ~n8470;
  assign n8472 = ~n8469 & ~n8470;
  assign n8473 = ~n8471 & ~n8472;
  assign n8474 = n8462 & ~n8473;
  assign n8475 = n8462 & ~n8474;
  assign n8476 = ~n8473 & ~n8474;
  assign n8477 = ~n8475 & ~n8476;
  assign n8478 = ~n8159 & ~n8161;
  assign n8479 = ~n8477 & ~n8478;
  assign n8480 = n8477 & n8478;
  assign n8481 = ~n8479 & ~n8480;
  assign n8482 = ~n8307 & n8481;
  assign n8483 = ~n8307 & ~n8482;
  assign n8484 = n8481 & ~n8482;
  assign n8485 = ~n8483 & ~n8484;
  assign n8486 = ~n8296 & ~n8485;
  assign n8487 = ~n8296 & ~n8486;
  assign n8488 = ~n8485 & ~n8486;
  assign n8489 = ~n8487 & ~n8488;
  assign n8490 = n1611 & n3784;
  assign n8491 = pi93  & n1745;
  assign n8492 = pi95  & n1609;
  assign n8493 = pi94  & n1604;
  assign n8494 = ~n8492 & ~n8493;
  assign n8495 = ~n8491 & n8494;
  assign n8496 = ~n8490 & n8495;
  assign n8497 = pi20  & ~n8496;
  assign n8498 = pi20  & ~n8497;
  assign n8499 = ~n8496 & ~n8497;
  assign n8500 = ~n8498 & ~n8499;
  assign n8501 = ~n8489 & ~n8500;
  assign n8502 = ~n8489 & ~n8501;
  assign n8503 = ~n8500 & ~n8501;
  assign n8504 = ~n8502 & ~n8503;
  assign n8505 = ~n8193 & ~n8196;
  assign n8506 = n8504 & n8505;
  assign n8507 = ~n8504 & ~n8505;
  assign n8508 = ~n8506 & ~n8507;
  assign n8509 = n1297 & n4454;
  assign n8510 = pi96  & n1366;
  assign n8511 = pi98  & n1295;
  assign n8512 = pi97  & n1290;
  assign n8513 = ~n8511 & ~n8512;
  assign n8514 = ~n8510 & n8513;
  assign n8515 = ~n8509 & n8514;
  assign n8516 = pi17  & ~n8515;
  assign n8517 = pi17  & ~n8516;
  assign n8518 = ~n8515 & ~n8516;
  assign n8519 = ~n8517 & ~n8518;
  assign n8520 = n8508 & ~n8519;
  assign n8521 = n8508 & ~n8520;
  assign n8522 = ~n8519 & ~n8520;
  assign n8523 = ~n8521 & ~n8522;
  assign n8524 = ~n8011 & ~n8213;
  assign n8525 = ~n8210 & ~n8524;
  assign n8526 = n8523 & n8525;
  assign n8527 = ~n8523 & ~n8525;
  assign n8528 = ~n8526 & ~n8527;
  assign n8529 = n938 & n5169;
  assign n8530 = pi99  & n1052;
  assign n8531 = pi101  & n936;
  assign n8532 = pi100  & n931;
  assign n8533 = ~n8531 & ~n8532;
  assign n8534 = ~n8530 & n8533;
  assign n8535 = ~n8529 & n8534;
  assign n8536 = pi14  & ~n8535;
  assign n8537 = pi14  & ~n8536;
  assign n8538 = ~n8535 & ~n8536;
  assign n8539 = ~n8537 & ~n8538;
  assign n8540 = n8528 & ~n8539;
  assign n8541 = n8528 & ~n8540;
  assign n8542 = ~n8539 & ~n8540;
  assign n8543 = ~n8541 & ~n8542;
  assign n8544 = ~n8228 & ~n8232;
  assign n8545 = n8543 & n8544;
  assign n8546 = ~n8543 & ~n8544;
  assign n8547 = ~n8545 & ~n8546;
  assign n8548 = n687 & n5943;
  assign n8549 = pi102  & n763;
  assign n8550 = pi104  & n685;
  assign n8551 = pi103  & n680;
  assign n8552 = ~n8550 & ~n8551;
  assign n8553 = ~n8549 & n8552;
  assign n8554 = ~n8548 & n8553;
  assign n8555 = pi11  & ~n8554;
  assign n8556 = pi11  & ~n8555;
  assign n8557 = ~n8554 & ~n8555;
  assign n8558 = ~n8556 & ~n8557;
  assign n8559 = n8547 & ~n8558;
  assign n8560 = n8547 & ~n8559;
  assign n8561 = ~n8558 & ~n8559;
  assign n8562 = ~n8560 & ~n8561;
  assign n8563 = ~n8245 & ~n8251;
  assign n8564 = n8562 & n8563;
  assign n8565 = ~n8562 & ~n8563;
  assign n8566 = ~n8564 & ~n8565;
  assign n8567 = n498 & n6775;
  assign n8568 = pi105  & n537;
  assign n8569 = pi107  & n496;
  assign n8570 = pi106  & n491;
  assign n8571 = ~n8569 & ~n8570;
  assign n8572 = ~n8568 & n8571;
  assign n8573 = ~n8567 & n8572;
  assign n8574 = pi8  & ~n8573;
  assign n8575 = pi8  & ~n8574;
  assign n8576 = ~n8573 & ~n8574;
  assign n8577 = ~n8575 & ~n8576;
  assign n8578 = n8566 & ~n8577;
  assign n8579 = n8566 & ~n8578;
  assign n8580 = ~n8577 & ~n8578;
  assign n8581 = ~n8579 & ~n8580;
  assign n8582 = ~n7944 & ~n8267;
  assign n8583 = ~n8264 & ~n8582;
  assign n8584 = n8581 & n8583;
  assign n8585 = ~n8581 & ~n8583;
  assign n8586 = ~n8584 & ~n8585;
  assign n8587 = n342 & n7665;
  assign n8588 = pi108  & n380;
  assign n8589 = pi110  & n340;
  assign n8590 = pi109  & n335;
  assign n8591 = ~n8589 & ~n8590;
  assign n8592 = ~n8588 & n8591;
  assign n8593 = ~n8587 & n8592;
  assign n8594 = pi5  & ~n8593;
  assign n8595 = pi5  & ~n8594;
  assign n8596 = ~n8593 & ~n8594;
  assign n8597 = ~n8595 & ~n8596;
  assign n8598 = n8586 & ~n8597;
  assign n8599 = n8586 & ~n8598;
  assign n8600 = ~n8597 & ~n8598;
  assign n8601 = ~n8599 & ~n8600;
  assign n8602 = ~n8282 & ~n8285;
  assign n8603 = n8601 & n8602;
  assign n8604 = ~n8601 & ~n8602;
  assign n8605 = ~n8603 & ~n8604;
  assign n8606 = ~n7993 & ~n7995;
  assign n8607 = ~pi112  & ~pi113 ;
  assign n8608 = pi112  & pi113 ;
  assign n8609 = ~n8607 & ~n8608;
  assign n8610 = ~n8606 & n8609;
  assign n8611 = n8606 & ~n8609;
  assign n8612 = ~n8610 & ~n8611;
  assign n8613 = n262 & n8612;
  assign n8614 = pi111  & n288;
  assign n8615 = pi113  & n267;
  assign n8616 = pi112  & n269;
  assign n8617 = ~n8615 & ~n8616;
  assign n8618 = ~n8614 & n8617;
  assign n8619 = ~n8613 & n8618;
  assign n8620 = pi2  & ~n8619;
  assign n8621 = pi2  & ~n8620;
  assign n8622 = ~n8619 & ~n8620;
  assign n8623 = ~n8621 & ~n8622;
  assign n8624 = ~n8605 & n8623;
  assign n8625 = n8605 & ~n8623;
  assign n8626 = ~n8624 & ~n8625;
  assign n8627 = ~n8294 & n8626;
  assign n8628 = n8294 & ~n8626;
  assign po49  = ~n8627 & ~n8628;
  assign n8630 = ~n8578 & ~n8585;
  assign n8631 = ~n8501 & ~n8507;
  assign n8632 = n1611 & n4001;
  assign n8633 = pi94  & n1745;
  assign n8634 = pi96  & n1609;
  assign n8635 = pi95  & n1604;
  assign n8636 = ~n8634 & ~n8635;
  assign n8637 = ~n8633 & n8636;
  assign n8638 = ~n8632 & n8637;
  assign n8639 = pi20  & ~n8638;
  assign n8640 = pi20  & ~n8639;
  assign n8641 = ~n8638 & ~n8639;
  assign n8642 = ~n8640 & ~n8641;
  assign n8643 = ~n8482 & ~n8486;
  assign n8644 = n2043 & n3371;
  assign n8645 = pi91  & n2180;
  assign n8646 = pi93  & n2041;
  assign n8647 = pi92  & n2036;
  assign n8648 = ~n8646 & ~n8647;
  assign n8649 = ~n8645 & n8648;
  assign n8650 = ~n8644 & n8649;
  assign n8651 = pi23  & ~n8650;
  assign n8652 = pi23  & ~n8651;
  assign n8653 = ~n8650 & ~n8651;
  assign n8654 = ~n8652 & ~n8653;
  assign n8655 = ~n8474 & ~n8479;
  assign n8656 = ~n8455 & ~n8461;
  assign n8657 = ~n8417 & ~n8423;
  assign n8658 = n1434 & n4271;
  assign n8659 = pi79  & n4503;
  assign n8660 = pi81  & n4269;
  assign n8661 = pi80  & n4264;
  assign n8662 = ~n8660 & ~n8661;
  assign n8663 = ~n8659 & n8662;
  assign n8664 = ~n8658 & n8663;
  assign n8665 = pi35  & ~n8664;
  assign n8666 = pi35  & ~n8665;
  assign n8667 = ~n8664 & ~n8665;
  assign n8668 = ~n8666 & ~n8667;
  assign n8669 = ~n8401 & ~n8403;
  assign n8670 = ~n8362 & ~n8368;
  assign n8671 = n576 & n6539;
  assign n8672 = pi70  & n6873;
  assign n8673 = pi72  & n6537;
  assign n8674 = pi71  & n6532;
  assign n8675 = ~n8673 & ~n8674;
  assign n8676 = ~n8672 & n8675;
  assign n8677 = ~n8671 & n8676;
  assign n8678 = pi44  & ~n8677;
  assign n8679 = pi44  & ~n8678;
  assign n8680 = ~n8677 & ~n8678;
  assign n8681 = ~n8679 & ~n8680;
  assign n8682 = ~n8346 & ~n8348;
  assign n8683 = n286 & n8334;
  assign n8684 = n8041 & n8326;
  assign n8685 = ~n8331 & n8684;
  assign n8686 = pi64  & n8685;
  assign n8687 = pi66  & n8332;
  assign n8688 = pi65  & n8327;
  assign n8689 = ~n8687 & ~n8688;
  assign n8690 = ~n8683 & n8689;
  assign n8691 = ~n8686 & n8690;
  assign n8692 = pi50  & ~n8691;
  assign n8693 = pi50  & ~n8692;
  assign n8694 = ~n8691 & ~n8692;
  assign n8695 = ~n8693 & ~n8694;
  assign n8696 = ~n8342 & n8695;
  assign n8697 = n8342 & ~n8695;
  assign n8698 = ~n8696 & ~n8697;
  assign n8699 = n401 & n7408;
  assign n8700 = pi67  & n7740;
  assign n8701 = pi69  & n7406;
  assign n8702 = pi68  & n7401;
  assign n8703 = ~n8701 & ~n8702;
  assign n8704 = ~n8700 & n8703;
  assign n8705 = ~n8699 & n8704;
  assign n8706 = pi47  & ~n8705;
  assign n8707 = pi47  & ~n8706;
  assign n8708 = ~n8705 & ~n8706;
  assign n8709 = ~n8707 & ~n8708;
  assign n8710 = n8698 & ~n8709;
  assign n8711 = n8698 & ~n8710;
  assign n8712 = ~n8709 & ~n8710;
  assign n8713 = ~n8711 & ~n8712;
  assign n8714 = ~n8682 & ~n8713;
  assign n8715 = n8682 & n8713;
  assign n8716 = ~n8714 & ~n8715;
  assign n8717 = ~n8681 & n8716;
  assign n8718 = ~n8681 & ~n8717;
  assign n8719 = n8716 & ~n8717;
  assign n8720 = ~n8718 & ~n8719;
  assign n8721 = ~n8670 & ~n8720;
  assign n8722 = ~n8670 & ~n8721;
  assign n8723 = ~n8720 & ~n8721;
  assign n8724 = ~n8722 & ~n8723;
  assign n8725 = n809 & n5739;
  assign n8726 = pi73  & n6030;
  assign n8727 = pi75  & n5737;
  assign n8728 = pi74  & n5732;
  assign n8729 = ~n8727 & ~n8728;
  assign n8730 = ~n8726 & n8729;
  assign n8731 = ~n8725 & n8730;
  assign n8732 = pi41  & ~n8731;
  assign n8733 = pi41  & ~n8732;
  assign n8734 = ~n8731 & ~n8732;
  assign n8735 = ~n8733 & ~n8734;
  assign n8736 = n8724 & n8735;
  assign n8737 = ~n8724 & ~n8735;
  assign n8738 = ~n8736 & ~n8737;
  assign n8739 = ~n8386 & n8738;
  assign n8740 = n8386 & ~n8738;
  assign n8741 = ~n8739 & ~n8740;
  assign n8742 = n1025 & n5008;
  assign n8743 = pi76  & n5241;
  assign n8744 = pi78  & n5006;
  assign n8745 = pi77  & n5001;
  assign n8746 = ~n8744 & ~n8745;
  assign n8747 = ~n8743 & n8746;
  assign n8748 = ~n8742 & n8747;
  assign n8749 = pi38  & ~n8748;
  assign n8750 = pi38  & ~n8749;
  assign n8751 = ~n8748 & ~n8749;
  assign n8752 = ~n8750 & ~n8751;
  assign n8753 = n8741 & ~n8752;
  assign n8754 = n8741 & ~n8753;
  assign n8755 = ~n8752 & ~n8753;
  assign n8756 = ~n8754 & ~n8755;
  assign n8757 = ~n8669 & ~n8756;
  assign n8758 = n8669 & n8756;
  assign n8759 = ~n8757 & ~n8758;
  assign n8760 = ~n8668 & n8759;
  assign n8761 = ~n8668 & ~n8760;
  assign n8762 = n8759 & ~n8760;
  assign n8763 = ~n8761 & ~n8762;
  assign n8764 = ~n8657 & ~n8763;
  assign n8765 = ~n8657 & ~n8764;
  assign n8766 = ~n8763 & ~n8764;
  assign n8767 = ~n8765 & ~n8766;
  assign n8768 = n1834 & n3622;
  assign n8769 = pi82  & n3814;
  assign n8770 = pi84  & n3620;
  assign n8771 = pi83  & n3615;
  assign n8772 = ~n8770 & ~n8771;
  assign n8773 = ~n8769 & n8772;
  assign n8774 = ~n8768 & n8773;
  assign n8775 = pi32  & ~n8774;
  assign n8776 = pi32  & ~n8775;
  assign n8777 = ~n8774 & ~n8775;
  assign n8778 = ~n8776 & ~n8777;
  assign n8779 = ~n8767 & ~n8778;
  assign n8780 = ~n8767 & ~n8779;
  assign n8781 = ~n8778 & ~n8779;
  assign n8782 = ~n8780 & ~n8781;
  assign n8783 = ~n8436 & ~n8442;
  assign n8784 = n8782 & n8783;
  assign n8785 = ~n8782 & ~n8783;
  assign n8786 = ~n8784 & ~n8785;
  assign n8787 = n2288 & n3034;
  assign n8788 = pi85  & n3225;
  assign n8789 = pi87  & n3032;
  assign n8790 = pi86  & n3027;
  assign n8791 = ~n8789 & ~n8790;
  assign n8792 = ~n8788 & n8791;
  assign n8793 = ~n8787 & n8792;
  assign n8794 = pi29  & ~n8793;
  assign n8795 = pi29  & ~n8794;
  assign n8796 = ~n8793 & ~n8794;
  assign n8797 = ~n8795 & ~n8796;
  assign n8798 = n8786 & ~n8797;
  assign n8799 = ~n8786 & n8797;
  assign n8800 = ~n8798 & ~n8799;
  assign n8801 = ~n8656 & n8800;
  assign n8802 = ~n8656 & ~n8801;
  assign n8803 = ~n8798 & ~n8801;
  assign n8804 = ~n8799 & n8803;
  assign n8805 = ~n8802 & ~n8804;
  assign n8806 = n2523 & n2801;
  assign n8807 = pi88  & n2667;
  assign n8808 = pi90  & n2521;
  assign n8809 = pi89  & n2516;
  assign n8810 = ~n8808 & ~n8809;
  assign n8811 = ~n8807 & n8810;
  assign n8812 = ~n8806 & n8811;
  assign n8813 = pi26  & ~n8812;
  assign n8814 = pi26  & ~n8813;
  assign n8815 = ~n8812 & ~n8813;
  assign n8816 = ~n8814 & ~n8815;
  assign n8817 = n8805 & n8816;
  assign n8818 = ~n8805 & ~n8816;
  assign n8819 = ~n8817 & ~n8818;
  assign n8820 = ~n8655 & n8819;
  assign n8821 = n8655 & ~n8819;
  assign n8822 = ~n8820 & ~n8821;
  assign n8823 = n8654 & ~n8822;
  assign n8824 = ~n8654 & n8822;
  assign n8825 = ~n8823 & ~n8824;
  assign n8826 = ~n8643 & n8825;
  assign n8827 = n8643 & ~n8825;
  assign n8828 = ~n8826 & ~n8827;
  assign n8829 = n8642 & ~n8828;
  assign n8830 = ~n8642 & n8828;
  assign n8831 = ~n8829 & ~n8830;
  assign n8832 = ~n8631 & n8831;
  assign n8833 = n8631 & ~n8831;
  assign n8834 = ~n8832 & ~n8833;
  assign n8835 = n1297 & n4684;
  assign n8836 = pi97  & n1366;
  assign n8837 = pi99  & n1295;
  assign n8838 = pi98  & n1290;
  assign n8839 = ~n8837 & ~n8838;
  assign n8840 = ~n8836 & n8839;
  assign n8841 = ~n8835 & n8840;
  assign n8842 = pi17  & ~n8841;
  assign n8843 = pi17  & ~n8842;
  assign n8844 = ~n8841 & ~n8842;
  assign n8845 = ~n8843 & ~n8844;
  assign n8846 = n8834 & ~n8845;
  assign n8847 = n8834 & ~n8846;
  assign n8848 = ~n8845 & ~n8846;
  assign n8849 = ~n8847 & ~n8848;
  assign n8850 = ~n8520 & ~n8527;
  assign n8851 = n8849 & n8850;
  assign n8852 = ~n8849 & ~n8850;
  assign n8853 = ~n8851 & ~n8852;
  assign n8854 = n938 & n5413;
  assign n8855 = pi100  & n1052;
  assign n8856 = pi102  & n936;
  assign n8857 = pi101  & n931;
  assign n8858 = ~n8856 & ~n8857;
  assign n8859 = ~n8855 & n8858;
  assign n8860 = ~n8854 & n8859;
  assign n8861 = pi14  & ~n8860;
  assign n8862 = pi14  & ~n8861;
  assign n8863 = ~n8860 & ~n8861;
  assign n8864 = ~n8862 & ~n8863;
  assign n8865 = n8853 & ~n8864;
  assign n8866 = n8853 & ~n8865;
  assign n8867 = ~n8864 & ~n8865;
  assign n8868 = ~n8866 & ~n8867;
  assign n8869 = ~n8540 & ~n8546;
  assign n8870 = n8868 & n8869;
  assign n8871 = ~n8868 & ~n8869;
  assign n8872 = ~n8870 & ~n8871;
  assign n8873 = n687 & n6207;
  assign n8874 = pi103  & n763;
  assign n8875 = pi105  & n685;
  assign n8876 = pi104  & n680;
  assign n8877 = ~n8875 & ~n8876;
  assign n8878 = ~n8874 & n8877;
  assign n8879 = ~n8873 & n8878;
  assign n8880 = pi11  & ~n8879;
  assign n8881 = pi11  & ~n8880;
  assign n8882 = ~n8879 & ~n8880;
  assign n8883 = ~n8881 & ~n8882;
  assign n8884 = n8872 & ~n8883;
  assign n8885 = n8872 & ~n8884;
  assign n8886 = ~n8883 & ~n8884;
  assign n8887 = ~n8885 & ~n8886;
  assign n8888 = ~n8559 & ~n8565;
  assign n8889 = n8887 & n8888;
  assign n8890 = ~n8887 & ~n8888;
  assign n8891 = ~n8889 & ~n8890;
  assign n8892 = n498 & n7060;
  assign n8893 = pi106  & n537;
  assign n8894 = pi108  & n496;
  assign n8895 = pi107  & n491;
  assign n8896 = ~n8894 & ~n8895;
  assign n8897 = ~n8893 & n8896;
  assign n8898 = ~n8892 & n8897;
  assign n8899 = pi8  & ~n8898;
  assign n8900 = pi8  & ~n8899;
  assign n8901 = ~n8898 & ~n8899;
  assign n8902 = ~n8900 & ~n8901;
  assign n8903 = n8891 & ~n8902;
  assign n8904 = ~n8891 & n8902;
  assign n8905 = ~n8903 & ~n8904;
  assign n8906 = ~n8630 & n8905;
  assign n8907 = ~n8630 & ~n8906;
  assign n8908 = ~n8903 & ~n8906;
  assign n8909 = ~n8904 & n8908;
  assign n8910 = ~n8907 & ~n8909;
  assign n8911 = n342 & n7970;
  assign n8912 = pi109  & n380;
  assign n8913 = pi111  & n340;
  assign n8914 = pi110  & n335;
  assign n8915 = ~n8913 & ~n8914;
  assign n8916 = ~n8912 & n8915;
  assign n8917 = ~n8911 & n8916;
  assign n8918 = pi5  & ~n8917;
  assign n8919 = pi5  & ~n8918;
  assign n8920 = ~n8917 & ~n8918;
  assign n8921 = ~n8919 & ~n8920;
  assign n8922 = ~n8910 & ~n8921;
  assign n8923 = ~n8910 & ~n8922;
  assign n8924 = ~n8921 & ~n8922;
  assign n8925 = ~n8923 & ~n8924;
  assign n8926 = ~n8598 & ~n8604;
  assign n8927 = n8925 & n8926;
  assign n8928 = ~n8925 & ~n8926;
  assign n8929 = ~n8927 & ~n8928;
  assign n8930 = ~n8608 & ~n8610;
  assign n8931 = ~pi113  & ~pi114 ;
  assign n8932 = pi113  & pi114 ;
  assign n8933 = ~n8931 & ~n8932;
  assign n8934 = ~n8930 & n8933;
  assign n8935 = n8930 & ~n8933;
  assign n8936 = ~n8934 & ~n8935;
  assign n8937 = n262 & n8936;
  assign n8938 = pi112  & n288;
  assign n8939 = pi114  & n267;
  assign n8940 = pi113  & n269;
  assign n8941 = ~n8939 & ~n8940;
  assign n8942 = ~n8938 & n8941;
  assign n8943 = ~n8937 & n8942;
  assign n8944 = pi2  & ~n8943;
  assign n8945 = pi2  & ~n8944;
  assign n8946 = ~n8943 & ~n8944;
  assign n8947 = ~n8945 & ~n8946;
  assign n8948 = n8929 & ~n8947;
  assign n8949 = n8929 & ~n8948;
  assign n8950 = ~n8947 & ~n8948;
  assign n8951 = ~n8949 & ~n8950;
  assign n8952 = ~n8625 & ~n8627;
  assign n8953 = ~n8951 & ~n8952;
  assign n8954 = n8951 & n8952;
  assign po50  = ~n8953 & ~n8954;
  assign n8956 = ~n8948 & ~n8953;
  assign n8957 = ~n8932 & ~n8934;
  assign n8958 = ~pi114  & ~pi115 ;
  assign n8959 = pi114  & pi115 ;
  assign n8960 = ~n8958 & ~n8959;
  assign n8961 = ~n8957 & n8960;
  assign n8962 = n8957 & ~n8960;
  assign n8963 = ~n8961 & ~n8962;
  assign n8964 = n262 & n8963;
  assign n8965 = pi113  & n288;
  assign n8966 = pi115  & n267;
  assign n8967 = pi114  & n269;
  assign n8968 = ~n8966 & ~n8967;
  assign n8969 = ~n8965 & n8968;
  assign n8970 = ~n8964 & n8969;
  assign n8971 = pi2  & ~n8970;
  assign n8972 = pi2  & ~n8971;
  assign n8973 = ~n8970 & ~n8971;
  assign n8974 = ~n8972 & ~n8973;
  assign n8975 = ~n8922 & ~n8928;
  assign n8976 = ~n8846 & ~n8852;
  assign n8977 = ~n8830 & ~n8832;
  assign n8978 = ~n8824 & ~n8826;
  assign n8979 = ~n8818 & ~n8820;
  assign n8980 = ~n8760 & ~n8764;
  assign n8981 = n1554 & n4271;
  assign n8982 = pi80  & n4503;
  assign n8983 = pi82  & n4269;
  assign n8984 = pi81  & n4264;
  assign n8985 = ~n8983 & ~n8984;
  assign n8986 = ~n8982 & n8985;
  assign n8987 = ~n8981 & n8986;
  assign n8988 = pi35  & ~n8987;
  assign n8989 = pi35  & ~n8988;
  assign n8990 = ~n8987 & ~n8988;
  assign n8991 = ~n8989 & ~n8990;
  assign n8992 = ~n8753 & ~n8757;
  assign n8993 = n1122 & n5008;
  assign n8994 = pi77  & n5241;
  assign n8995 = pi79  & n5006;
  assign n8996 = pi78  & n5001;
  assign n8997 = ~n8995 & ~n8996;
  assign n8998 = ~n8994 & n8997;
  assign n8999 = ~n8993 & n8998;
  assign n9000 = pi38  & ~n8999;
  assign n9001 = pi38  & ~n9000;
  assign n9002 = ~n8999 & ~n9000;
  assign n9003 = ~n9001 & ~n9002;
  assign n9004 = ~n8737 & ~n8739;
  assign n9005 = n891 & n5739;
  assign n9006 = pi74  & n6030;
  assign n9007 = pi76  & n5737;
  assign n9008 = pi75  & n5732;
  assign n9009 = ~n9007 & ~n9008;
  assign n9010 = ~n9006 & n9009;
  assign n9011 = ~n9005 & n9010;
  assign n9012 = pi41  & ~n9011;
  assign n9013 = pi41  & ~n9012;
  assign n9014 = ~n9011 & ~n9012;
  assign n9015 = ~n9013 & ~n9014;
  assign n9016 = ~n8717 & ~n8721;
  assign n9017 = pi50  & ~pi51 ;
  assign n9018 = ~pi50  & pi51 ;
  assign n9019 = ~n9017 & ~n9018;
  assign n9020 = pi64  & ~n9019;
  assign n9021 = ~n8697 & n9020;
  assign n9022 = n8697 & ~n9020;
  assign n9023 = ~n9021 & ~n9022;
  assign n9024 = n309 & n8334;
  assign n9025 = pi65  & n8685;
  assign n9026 = pi67  & n8332;
  assign n9027 = pi66  & n8327;
  assign n9028 = ~n9026 & ~n9027;
  assign n9029 = ~n9025 & n9028;
  assign n9030 = ~n9024 & n9029;
  assign n9031 = pi50  & ~n9030;
  assign n9032 = pi50  & ~n9031;
  assign n9033 = ~n9030 & ~n9031;
  assign n9034 = ~n9032 & ~n9033;
  assign n9035 = ~n9023 & ~n9034;
  assign n9036 = n9023 & n9034;
  assign n9037 = ~n9035 & ~n9036;
  assign n9038 = n450 & n7408;
  assign n9039 = pi68  & n7740;
  assign n9040 = pi70  & n7406;
  assign n9041 = pi69  & n7401;
  assign n9042 = ~n9040 & ~n9041;
  assign n9043 = ~n9039 & n9042;
  assign n9044 = ~n9038 & n9043;
  assign n9045 = pi47  & ~n9044;
  assign n9046 = pi47  & ~n9045;
  assign n9047 = ~n9044 & ~n9045;
  assign n9048 = ~n9046 & ~n9047;
  assign n9049 = n9037 & ~n9048;
  assign n9050 = n9037 & ~n9049;
  assign n9051 = ~n9048 & ~n9049;
  assign n9052 = ~n9050 & ~n9051;
  assign n9053 = ~n8710 & ~n8714;
  assign n9054 = n9052 & n9053;
  assign n9055 = ~n9052 & ~n9053;
  assign n9056 = ~n9054 & ~n9055;
  assign n9057 = n642 & n6539;
  assign n9058 = pi71  & n6873;
  assign n9059 = pi73  & n6537;
  assign n9060 = pi72  & n6532;
  assign n9061 = ~n9059 & ~n9060;
  assign n9062 = ~n9058 & n9061;
  assign n9063 = ~n9057 & n9062;
  assign n9064 = pi44  & ~n9063;
  assign n9065 = pi44  & ~n9064;
  assign n9066 = ~n9063 & ~n9064;
  assign n9067 = ~n9065 & ~n9066;
  assign n9068 = ~n9056 & n9067;
  assign n9069 = n9056 & ~n9067;
  assign n9070 = ~n9068 & ~n9069;
  assign n9071 = ~n9016 & n9070;
  assign n9072 = n9016 & ~n9070;
  assign n9073 = ~n9071 & ~n9072;
  assign n9074 = ~n9015 & n9073;
  assign n9075 = ~n9015 & ~n9074;
  assign n9076 = n9073 & ~n9074;
  assign n9077 = ~n9075 & ~n9076;
  assign n9078 = ~n9004 & ~n9077;
  assign n9079 = n9004 & n9077;
  assign n9080 = ~n9078 & ~n9079;
  assign n9081 = ~n9003 & n9080;
  assign n9082 = n9003 & ~n9080;
  assign n9083 = ~n9081 & ~n9082;
  assign n9084 = ~n8992 & n9083;
  assign n9085 = n8992 & ~n9083;
  assign n9086 = ~n9084 & ~n9085;
  assign n9087 = ~n8991 & n9086;
  assign n9088 = n8991 & ~n9086;
  assign n9089 = ~n9087 & ~n9088;
  assign n9090 = ~n8980 & n9089;
  assign n9091 = n8980 & ~n9089;
  assign n9092 = ~n9090 & ~n9091;
  assign n9093 = n1972 & n3622;
  assign n9094 = pi83  & n3814;
  assign n9095 = pi85  & n3620;
  assign n9096 = pi84  & n3615;
  assign n9097 = ~n9095 & ~n9096;
  assign n9098 = ~n9094 & n9097;
  assign n9099 = ~n9093 & n9098;
  assign n9100 = pi32  & ~n9099;
  assign n9101 = pi32  & ~n9100;
  assign n9102 = ~n9099 & ~n9100;
  assign n9103 = ~n9101 & ~n9102;
  assign n9104 = n9092 & ~n9103;
  assign n9105 = n9092 & ~n9104;
  assign n9106 = ~n9103 & ~n9104;
  assign n9107 = ~n9105 & ~n9106;
  assign n9108 = ~n8779 & ~n8785;
  assign n9109 = n9107 & n9108;
  assign n9110 = ~n9107 & ~n9108;
  assign n9111 = ~n9109 & ~n9110;
  assign n9112 = n2446 & n3034;
  assign n9113 = pi86  & n3225;
  assign n9114 = pi88  & n3032;
  assign n9115 = pi87  & n3027;
  assign n9116 = ~n9114 & ~n9115;
  assign n9117 = ~n9113 & n9116;
  assign n9118 = ~n9112 & n9117;
  assign n9119 = pi29  & ~n9118;
  assign n9120 = pi29  & ~n9119;
  assign n9121 = ~n9118 & ~n9119;
  assign n9122 = ~n9120 & ~n9121;
  assign n9123 = ~n9111 & n9122;
  assign n9124 = n9111 & ~n9122;
  assign n9125 = ~n9123 & ~n9124;
  assign n9126 = ~n8803 & n9125;
  assign n9127 = n8803 & ~n9125;
  assign n9128 = ~n9126 & ~n9127;
  assign n9129 = n2523 & n2978;
  assign n9130 = pi89  & n2667;
  assign n9131 = pi91  & n2521;
  assign n9132 = pi90  & n2516;
  assign n9133 = ~n9131 & ~n9132;
  assign n9134 = ~n9130 & n9133;
  assign n9135 = ~n9129 & n9134;
  assign n9136 = pi26  & ~n9135;
  assign n9137 = pi26  & ~n9136;
  assign n9138 = ~n9135 & ~n9136;
  assign n9139 = ~n9137 & ~n9138;
  assign n9140 = n9128 & ~n9139;
  assign n9141 = n9128 & ~n9140;
  assign n9142 = ~n9139 & ~n9140;
  assign n9143 = ~n9141 & ~n9142;
  assign n9144 = ~n8979 & n9143;
  assign n9145 = n8979 & ~n9143;
  assign n9146 = ~n9144 & ~n9145;
  assign n9147 = n2043 & n3565;
  assign n9148 = pi92  & n2180;
  assign n9149 = pi94  & n2041;
  assign n9150 = pi93  & n2036;
  assign n9151 = ~n9149 & ~n9150;
  assign n9152 = ~n9148 & n9151;
  assign n9153 = ~n9147 & n9152;
  assign n9154 = pi23  & ~n9153;
  assign n9155 = pi23  & ~n9154;
  assign n9156 = ~n9153 & ~n9154;
  assign n9157 = ~n9155 & ~n9156;
  assign n9158 = ~n9146 & ~n9157;
  assign n9159 = n9146 & n9157;
  assign n9160 = ~n9158 & ~n9159;
  assign n9161 = ~n8978 & n9160;
  assign n9162 = n8978 & ~n9160;
  assign n9163 = ~n9161 & ~n9162;
  assign n9164 = n1611 & n4211;
  assign n9165 = pi95  & n1745;
  assign n9166 = pi97  & n1609;
  assign n9167 = pi96  & n1604;
  assign n9168 = ~n9166 & ~n9167;
  assign n9169 = ~n9165 & n9168;
  assign n9170 = ~n9164 & n9169;
  assign n9171 = pi20  & ~n9170;
  assign n9172 = pi20  & ~n9171;
  assign n9173 = ~n9170 & ~n9171;
  assign n9174 = ~n9172 & ~n9173;
  assign n9175 = n9163 & ~n9174;
  assign n9176 = n9163 & ~n9175;
  assign n9177 = ~n9174 & ~n9175;
  assign n9178 = ~n9176 & ~n9177;
  assign n9179 = ~n8977 & n9178;
  assign n9180 = n8977 & ~n9178;
  assign n9181 = ~n9179 & ~n9180;
  assign n9182 = n1297 & n4910;
  assign n9183 = pi98  & n1366;
  assign n9184 = pi100  & n1295;
  assign n9185 = pi99  & n1290;
  assign n9186 = ~n9184 & ~n9185;
  assign n9187 = ~n9183 & n9186;
  assign n9188 = ~n9182 & n9187;
  assign n9189 = pi17  & ~n9188;
  assign n9190 = pi17  & ~n9189;
  assign n9191 = ~n9188 & ~n9189;
  assign n9192 = ~n9190 & ~n9191;
  assign n9193 = ~n9181 & ~n9192;
  assign n9194 = n9181 & n9192;
  assign n9195 = ~n9193 & ~n9194;
  assign n9196 = n8976 & ~n9195;
  assign n9197 = ~n8976 & n9195;
  assign n9198 = ~n9196 & ~n9197;
  assign n9199 = n938 & n5664;
  assign n9200 = pi101  & n1052;
  assign n9201 = pi103  & n936;
  assign n9202 = pi102  & n931;
  assign n9203 = ~n9201 & ~n9202;
  assign n9204 = ~n9200 & n9203;
  assign n9205 = ~n9199 & n9204;
  assign n9206 = pi14  & ~n9205;
  assign n9207 = pi14  & ~n9206;
  assign n9208 = ~n9205 & ~n9206;
  assign n9209 = ~n9207 & ~n9208;
  assign n9210 = n9198 & ~n9209;
  assign n9211 = n9198 & ~n9210;
  assign n9212 = ~n9209 & ~n9210;
  assign n9213 = ~n9211 & ~n9212;
  assign n9214 = ~n8865 & ~n8871;
  assign n9215 = n9213 & n9214;
  assign n9216 = ~n9213 & ~n9214;
  assign n9217 = ~n9215 & ~n9216;
  assign n9218 = n687 & n6477;
  assign n9219 = pi104  & n763;
  assign n9220 = pi106  & n685;
  assign n9221 = pi105  & n680;
  assign n9222 = ~n9220 & ~n9221;
  assign n9223 = ~n9219 & n9222;
  assign n9224 = ~n9218 & n9223;
  assign n9225 = pi11  & ~n9224;
  assign n9226 = pi11  & ~n9225;
  assign n9227 = ~n9224 & ~n9225;
  assign n9228 = ~n9226 & ~n9227;
  assign n9229 = ~n9217 & n9228;
  assign n9230 = n9217 & ~n9228;
  assign n9231 = ~n9229 & ~n9230;
  assign n9232 = ~n8884 & ~n8890;
  assign n9233 = n9231 & ~n9232;
  assign n9234 = ~n9231 & n9232;
  assign n9235 = ~n9233 & ~n9234;
  assign n9236 = n498 & n7349;
  assign n9237 = pi107  & n537;
  assign n9238 = pi109  & n496;
  assign n9239 = pi108  & n491;
  assign n9240 = ~n9238 & ~n9239;
  assign n9241 = ~n9237 & n9240;
  assign n9242 = ~n9236 & n9241;
  assign n9243 = pi8  & ~n9242;
  assign n9244 = pi8  & ~n9243;
  assign n9245 = ~n9242 & ~n9243;
  assign n9246 = ~n9244 & ~n9245;
  assign n9247 = n9235 & ~n9246;
  assign n9248 = n9235 & ~n9247;
  assign n9249 = ~n9246 & ~n9247;
  assign n9250 = ~n9248 & ~n9249;
  assign n9251 = ~n8908 & n9250;
  assign n9252 = n8908 & ~n9250;
  assign n9253 = ~n9251 & ~n9252;
  assign n9254 = n342 & n7997;
  assign n9255 = pi110  & n380;
  assign n9256 = pi112  & n340;
  assign n9257 = pi111  & n335;
  assign n9258 = ~n9256 & ~n9257;
  assign n9259 = ~n9255 & n9258;
  assign n9260 = ~n9254 & n9259;
  assign n9261 = pi5  & ~n9260;
  assign n9262 = pi5  & ~n9261;
  assign n9263 = ~n9260 & ~n9261;
  assign n9264 = ~n9262 & ~n9263;
  assign n9265 = n9253 & n9264;
  assign n9266 = ~n9253 & ~n9264;
  assign n9267 = ~n9265 & ~n9266;
  assign n9268 = ~n8975 & n9267;
  assign n9269 = n8975 & ~n9267;
  assign n9270 = ~n9268 & ~n9269;
  assign n9271 = ~n8974 & n9270;
  assign n9272 = n8974 & ~n9270;
  assign n9273 = ~n9271 & ~n9272;
  assign n9274 = ~n8956 & n9273;
  assign n9275 = n8956 & ~n9273;
  assign po51  = ~n9274 & ~n9275;
  assign n9277 = ~n9271 & ~n9274;
  assign n9278 = ~n9266 & ~n9268;
  assign n9279 = ~n9230 & ~n9233;
  assign n9280 = ~n8979 & ~n9143;
  assign n9281 = ~n9140 & ~n9280;
  assign n9282 = ~n9124 & ~n9126;
  assign n9283 = ~n9087 & ~n9090;
  assign n9284 = ~n9074 & ~n9078;
  assign n9285 = ~n9069 & ~n9071;
  assign n9286 = n8697 & n9020;
  assign n9287 = ~n9035 & ~n9286;
  assign n9288 = n359 & n8334;
  assign n9289 = pi66  & n8685;
  assign n9290 = pi68  & n8332;
  assign n9291 = pi67  & n8327;
  assign n9292 = ~n9290 & ~n9291;
  assign n9293 = ~n9289 & n9292;
  assign n9294 = ~n9288 & n9293;
  assign n9295 = pi50  & ~n9294;
  assign n9296 = pi50  & ~n9295;
  assign n9297 = ~n9294 & ~n9295;
  assign n9298 = ~n9296 & ~n9297;
  assign n9299 = pi53  & ~n9020;
  assign n9300 = ~pi51  & pi52 ;
  assign n9301 = pi51  & ~pi52 ;
  assign n9302 = ~n9300 & ~n9301;
  assign n9303 = n9019 & ~n9302;
  assign n9304 = pi64  & n9303;
  assign n9305 = ~pi52  & pi53 ;
  assign n9306 = pi52  & ~pi53 ;
  assign n9307 = ~n9305 & ~n9306;
  assign n9308 = ~n9019 & n9307;
  assign n9309 = pi65  & n9308;
  assign n9310 = ~n9019 & ~n9307;
  assign n9311 = ~n265 & n9310;
  assign n9312 = ~n9304 & ~n9309;
  assign n9313 = ~n9311 & n9312;
  assign n9314 = pi53  & ~n9313;
  assign n9315 = pi53  & ~n9314;
  assign n9316 = ~n9313 & ~n9314;
  assign n9317 = ~n9315 & ~n9316;
  assign n9318 = n9299 & ~n9317;
  assign n9319 = ~n9299 & n9317;
  assign n9320 = ~n9318 & ~n9319;
  assign n9321 = n9298 & ~n9320;
  assign n9322 = ~n9298 & n9320;
  assign n9323 = ~n9321 & ~n9322;
  assign n9324 = ~n9287 & n9323;
  assign n9325 = n9287 & ~n9323;
  assign n9326 = ~n9324 & ~n9325;
  assign n9327 = n475 & n7408;
  assign n9328 = pi69  & n7740;
  assign n9329 = pi71  & n7406;
  assign n9330 = pi70  & n7401;
  assign n9331 = ~n9329 & ~n9330;
  assign n9332 = ~n9328 & n9331;
  assign n9333 = ~n9327 & n9332;
  assign n9334 = pi47  & ~n9333;
  assign n9335 = pi47  & ~n9334;
  assign n9336 = ~n9333 & ~n9334;
  assign n9337 = ~n9335 & ~n9336;
  assign n9338 = n9326 & ~n9337;
  assign n9339 = n9326 & ~n9338;
  assign n9340 = ~n9337 & ~n9338;
  assign n9341 = ~n9339 & ~n9340;
  assign n9342 = ~n9049 & ~n9055;
  assign n9343 = n9341 & n9342;
  assign n9344 = ~n9341 & ~n9342;
  assign n9345 = ~n9343 & ~n9344;
  assign n9346 = n729 & n6539;
  assign n9347 = pi72  & n6873;
  assign n9348 = pi74  & n6537;
  assign n9349 = pi73  & n6532;
  assign n9350 = ~n9348 & ~n9349;
  assign n9351 = ~n9347 & n9350;
  assign n9352 = ~n9346 & n9351;
  assign n9353 = pi44  & ~n9352;
  assign n9354 = pi44  & ~n9353;
  assign n9355 = ~n9352 & ~n9353;
  assign n9356 = ~n9354 & ~n9355;
  assign n9357 = n9345 & ~n9356;
  assign n9358 = ~n9345 & n9356;
  assign n9359 = ~n9357 & ~n9358;
  assign n9360 = ~n9285 & n9359;
  assign n9361 = ~n9285 & ~n9360;
  assign n9362 = ~n9357 & ~n9360;
  assign n9363 = ~n9358 & n9362;
  assign n9364 = ~n9361 & ~n9363;
  assign n9365 = n999 & n5739;
  assign n9366 = pi75  & n6030;
  assign n9367 = pi77  & n5737;
  assign n9368 = pi76  & n5732;
  assign n9369 = ~n9367 & ~n9368;
  assign n9370 = ~n9366 & n9369;
  assign n9371 = ~n9365 & n9370;
  assign n9372 = pi41  & ~n9371;
  assign n9373 = pi41  & ~n9372;
  assign n9374 = ~n9371 & ~n9372;
  assign n9375 = ~n9373 & ~n9374;
  assign n9376 = n9364 & n9375;
  assign n9377 = ~n9364 & ~n9375;
  assign n9378 = ~n9376 & ~n9377;
  assign n9379 = ~n9284 & n9378;
  assign n9380 = n9284 & ~n9378;
  assign n9381 = ~n9379 & ~n9380;
  assign n9382 = n1225 & n5008;
  assign n9383 = pi78  & n5241;
  assign n9384 = pi80  & n5006;
  assign n9385 = pi79  & n5001;
  assign n9386 = ~n9384 & ~n9385;
  assign n9387 = ~n9383 & n9386;
  assign n9388 = ~n9382 & n9387;
  assign n9389 = pi38  & ~n9388;
  assign n9390 = pi38  & ~n9389;
  assign n9391 = ~n9388 & ~n9389;
  assign n9392 = ~n9390 & ~n9391;
  assign n9393 = n9381 & ~n9392;
  assign n9394 = n9381 & ~n9393;
  assign n9395 = ~n9392 & ~n9393;
  assign n9396 = ~n9394 & ~n9395;
  assign n9397 = ~n9081 & ~n9084;
  assign n9398 = n9396 & n9397;
  assign n9399 = ~n9396 & ~n9397;
  assign n9400 = ~n9398 & ~n9399;
  assign n9401 = n1696 & n4271;
  assign n9402 = pi81  & n4503;
  assign n9403 = pi83  & n4269;
  assign n9404 = pi82  & n4264;
  assign n9405 = ~n9403 & ~n9404;
  assign n9406 = ~n9402 & n9405;
  assign n9407 = ~n9401 & n9406;
  assign n9408 = pi35  & ~n9407;
  assign n9409 = pi35  & ~n9408;
  assign n9410 = ~n9407 & ~n9408;
  assign n9411 = ~n9409 & ~n9410;
  assign n9412 = n9400 & ~n9411;
  assign n9413 = ~n9400 & n9411;
  assign n9414 = ~n9412 & ~n9413;
  assign n9415 = ~n9283 & n9414;
  assign n9416 = ~n9283 & ~n9415;
  assign n9417 = ~n9412 & ~n9415;
  assign n9418 = ~n9413 & n9417;
  assign n9419 = ~n9416 & ~n9418;
  assign n9420 = n2133 & n3622;
  assign n9421 = pi84  & n3814;
  assign n9422 = pi86  & n3620;
  assign n9423 = pi85  & n3615;
  assign n9424 = ~n9422 & ~n9423;
  assign n9425 = ~n9421 & n9424;
  assign n9426 = ~n9420 & n9425;
  assign n9427 = pi32  & ~n9426;
  assign n9428 = pi32  & ~n9427;
  assign n9429 = ~n9426 & ~n9427;
  assign n9430 = ~n9428 & ~n9429;
  assign n9431 = ~n9419 & ~n9430;
  assign n9432 = ~n9419 & ~n9431;
  assign n9433 = ~n9430 & ~n9431;
  assign n9434 = ~n9432 & ~n9433;
  assign n9435 = ~n9104 & ~n9110;
  assign n9436 = n9434 & n9435;
  assign n9437 = ~n9434 & ~n9435;
  assign n9438 = ~n9436 & ~n9437;
  assign n9439 = n2473 & n3034;
  assign n9440 = pi87  & n3225;
  assign n9441 = pi89  & n3032;
  assign n9442 = pi88  & n3027;
  assign n9443 = ~n9441 & ~n9442;
  assign n9444 = ~n9440 & n9443;
  assign n9445 = ~n9439 & n9444;
  assign n9446 = pi29  & ~n9445;
  assign n9447 = pi29  & ~n9446;
  assign n9448 = ~n9445 & ~n9446;
  assign n9449 = ~n9447 & ~n9448;
  assign n9450 = n9438 & ~n9449;
  assign n9451 = n9438 & ~n9450;
  assign n9452 = ~n9449 & ~n9450;
  assign n9453 = ~n9451 & ~n9452;
  assign n9454 = ~n9282 & n9453;
  assign n9455 = n9282 & ~n9453;
  assign n9456 = ~n9454 & ~n9455;
  assign n9457 = n2523 & n3177;
  assign n9458 = pi90  & n2667;
  assign n9459 = pi92  & n2521;
  assign n9460 = pi91  & n2516;
  assign n9461 = ~n9459 & ~n9460;
  assign n9462 = ~n9458 & n9461;
  assign n9463 = ~n9457 & n9462;
  assign n9464 = pi26  & ~n9463;
  assign n9465 = pi26  & ~n9464;
  assign n9466 = ~n9463 & ~n9464;
  assign n9467 = ~n9465 & ~n9466;
  assign n9468 = ~n9456 & ~n9467;
  assign n9469 = n9456 & n9467;
  assign n9470 = ~n9468 & ~n9469;
  assign n9471 = n9281 & ~n9470;
  assign n9472 = ~n9281 & n9470;
  assign n9473 = ~n9471 & ~n9472;
  assign n9474 = n2043 & n3784;
  assign n9475 = pi93  & n2180;
  assign n9476 = pi95  & n2041;
  assign n9477 = pi94  & n2036;
  assign n9478 = ~n9476 & ~n9477;
  assign n9479 = ~n9475 & n9478;
  assign n9480 = ~n9474 & n9479;
  assign n9481 = pi23  & ~n9480;
  assign n9482 = pi23  & ~n9481;
  assign n9483 = ~n9480 & ~n9481;
  assign n9484 = ~n9482 & ~n9483;
  assign n9485 = n9473 & ~n9484;
  assign n9486 = n9473 & ~n9485;
  assign n9487 = ~n9484 & ~n9485;
  assign n9488 = ~n9486 & ~n9487;
  assign n9489 = ~n9158 & ~n9161;
  assign n9490 = n9488 & n9489;
  assign n9491 = ~n9488 & ~n9489;
  assign n9492 = ~n9490 & ~n9491;
  assign n9493 = n1611 & n4454;
  assign n9494 = pi96  & n1745;
  assign n9495 = pi98  & n1609;
  assign n9496 = pi97  & n1604;
  assign n9497 = ~n9495 & ~n9496;
  assign n9498 = ~n9494 & n9497;
  assign n9499 = ~n9493 & n9498;
  assign n9500 = pi20  & ~n9499;
  assign n9501 = pi20  & ~n9500;
  assign n9502 = ~n9499 & ~n9500;
  assign n9503 = ~n9501 & ~n9502;
  assign n9504 = n9492 & ~n9503;
  assign n9505 = n9492 & ~n9504;
  assign n9506 = ~n9503 & ~n9504;
  assign n9507 = ~n9505 & ~n9506;
  assign n9508 = ~n8977 & ~n9178;
  assign n9509 = ~n9175 & ~n9508;
  assign n9510 = n9507 & n9509;
  assign n9511 = ~n9507 & ~n9509;
  assign n9512 = ~n9510 & ~n9511;
  assign n9513 = n1297 & n5169;
  assign n9514 = pi99  & n1366;
  assign n9515 = pi101  & n1295;
  assign n9516 = pi100  & n1290;
  assign n9517 = ~n9515 & ~n9516;
  assign n9518 = ~n9514 & n9517;
  assign n9519 = ~n9513 & n9518;
  assign n9520 = pi17  & ~n9519;
  assign n9521 = pi17  & ~n9520;
  assign n9522 = ~n9519 & ~n9520;
  assign n9523 = ~n9521 & ~n9522;
  assign n9524 = n9512 & ~n9523;
  assign n9525 = n9512 & ~n9524;
  assign n9526 = ~n9523 & ~n9524;
  assign n9527 = ~n9525 & ~n9526;
  assign n9528 = ~n9193 & ~n9197;
  assign n9529 = n9527 & n9528;
  assign n9530 = ~n9527 & ~n9528;
  assign n9531 = ~n9529 & ~n9530;
  assign n9532 = n938 & n5943;
  assign n9533 = pi102  & n1052;
  assign n9534 = pi104  & n936;
  assign n9535 = pi103  & n931;
  assign n9536 = ~n9534 & ~n9535;
  assign n9537 = ~n9533 & n9536;
  assign n9538 = ~n9532 & n9537;
  assign n9539 = pi14  & ~n9538;
  assign n9540 = pi14  & ~n9539;
  assign n9541 = ~n9538 & ~n9539;
  assign n9542 = ~n9540 & ~n9541;
  assign n9543 = n9531 & ~n9542;
  assign n9544 = n9531 & ~n9543;
  assign n9545 = ~n9542 & ~n9543;
  assign n9546 = ~n9544 & ~n9545;
  assign n9547 = ~n9210 & ~n9216;
  assign n9548 = n9546 & n9547;
  assign n9549 = ~n9546 & ~n9547;
  assign n9550 = ~n9548 & ~n9549;
  assign n9551 = n687 & n6775;
  assign n9552 = pi105  & n763;
  assign n9553 = pi107  & n685;
  assign n9554 = pi106  & n680;
  assign n9555 = ~n9553 & ~n9554;
  assign n9556 = ~n9552 & n9555;
  assign n9557 = ~n9551 & n9556;
  assign n9558 = pi11  & ~n9557;
  assign n9559 = pi11  & ~n9558;
  assign n9560 = ~n9557 & ~n9558;
  assign n9561 = ~n9559 & ~n9560;
  assign n9562 = n9550 & ~n9561;
  assign n9563 = ~n9550 & n9561;
  assign n9564 = ~n9562 & ~n9563;
  assign n9565 = ~n9279 & n9564;
  assign n9566 = ~n9279 & ~n9565;
  assign n9567 = ~n9562 & ~n9565;
  assign n9568 = ~n9563 & n9567;
  assign n9569 = ~n9566 & ~n9568;
  assign n9570 = n498 & n7665;
  assign n9571 = pi108  & n537;
  assign n9572 = pi110  & n496;
  assign n9573 = pi109  & n491;
  assign n9574 = ~n9572 & ~n9573;
  assign n9575 = ~n9571 & n9574;
  assign n9576 = ~n9570 & n9575;
  assign n9577 = pi8  & ~n9576;
  assign n9578 = pi8  & ~n9577;
  assign n9579 = ~n9576 & ~n9577;
  assign n9580 = ~n9578 & ~n9579;
  assign n9581 = ~n9569 & ~n9580;
  assign n9582 = ~n9569 & ~n9581;
  assign n9583 = ~n9580 & ~n9581;
  assign n9584 = ~n9582 & ~n9583;
  assign n9585 = ~n8908 & ~n9250;
  assign n9586 = ~n9247 & ~n9585;
  assign n9587 = n9584 & n9586;
  assign n9588 = ~n9584 & ~n9586;
  assign n9589 = ~n9587 & ~n9588;
  assign n9590 = n342 & n8612;
  assign n9591 = pi111  & n380;
  assign n9592 = pi113  & n340;
  assign n9593 = pi112  & n335;
  assign n9594 = ~n9592 & ~n9593;
  assign n9595 = ~n9591 & n9594;
  assign n9596 = ~n9590 & n9595;
  assign n9597 = pi5  & ~n9596;
  assign n9598 = pi5  & ~n9597;
  assign n9599 = ~n9596 & ~n9597;
  assign n9600 = ~n9598 & ~n9599;
  assign n9601 = n9589 & ~n9600;
  assign n9602 = n9589 & ~n9601;
  assign n9603 = ~n9600 & ~n9601;
  assign n9604 = ~n9602 & ~n9603;
  assign n9605 = ~n9278 & n9604;
  assign n9606 = n9278 & ~n9604;
  assign n9607 = ~n9605 & ~n9606;
  assign n9608 = ~n8959 & ~n8961;
  assign n9609 = ~pi115  & ~pi116 ;
  assign n9610 = pi115  & pi116 ;
  assign n9611 = ~n9609 & ~n9610;
  assign n9612 = ~n9608 & n9611;
  assign n9613 = n9608 & ~n9611;
  assign n9614 = ~n9612 & ~n9613;
  assign n9615 = n262 & n9614;
  assign n9616 = pi114  & n288;
  assign n9617 = pi116  & n267;
  assign n9618 = pi115  & n269;
  assign n9619 = ~n9617 & ~n9618;
  assign n9620 = ~n9616 & n9619;
  assign n9621 = ~n9615 & n9620;
  assign n9622 = pi2  & ~n9621;
  assign n9623 = pi2  & ~n9622;
  assign n9624 = ~n9621 & ~n9622;
  assign n9625 = ~n9623 & ~n9624;
  assign n9626 = ~n9607 & ~n9625;
  assign n9627 = n9607 & n9625;
  assign n9628 = ~n9626 & ~n9627;
  assign n9629 = ~n9277 & n9628;
  assign n9630 = n9277 & ~n9628;
  assign po52  = ~n9629 & ~n9630;
  assign n9632 = ~n9626 & ~n9629;
  assign n9633 = ~n9278 & ~n9604;
  assign n9634 = ~n9601 & ~n9633;
  assign n9635 = ~n9485 & ~n9491;
  assign n9636 = n2043 & n4001;
  assign n9637 = pi94  & n2180;
  assign n9638 = pi96  & n2041;
  assign n9639 = pi95  & n2036;
  assign n9640 = ~n9638 & ~n9639;
  assign n9641 = ~n9637 & n9640;
  assign n9642 = ~n9636 & n9641;
  assign n9643 = pi23  & ~n9642;
  assign n9644 = pi23  & ~n9643;
  assign n9645 = ~n9642 & ~n9643;
  assign n9646 = ~n9644 & ~n9645;
  assign n9647 = ~n9468 & ~n9472;
  assign n9648 = n2523 & n3371;
  assign n9649 = pi91  & n2667;
  assign n9650 = pi93  & n2521;
  assign n9651 = pi92  & n2516;
  assign n9652 = ~n9650 & ~n9651;
  assign n9653 = ~n9649 & n9652;
  assign n9654 = ~n9648 & n9653;
  assign n9655 = pi26  & ~n9654;
  assign n9656 = pi26  & ~n9655;
  assign n9657 = ~n9654 & ~n9655;
  assign n9658 = ~n9656 & ~n9657;
  assign n9659 = ~n9282 & ~n9453;
  assign n9660 = ~n9450 & ~n9659;
  assign n9661 = ~n9431 & ~n9437;
  assign n9662 = n2288 & n3622;
  assign n9663 = pi85  & n3814;
  assign n9664 = pi87  & n3620;
  assign n9665 = pi86  & n3615;
  assign n9666 = ~n9664 & ~n9665;
  assign n9667 = ~n9663 & n9666;
  assign n9668 = ~n9662 & n9667;
  assign n9669 = pi32  & ~n9668;
  assign n9670 = pi32  & ~n9669;
  assign n9671 = ~n9668 & ~n9669;
  assign n9672 = ~n9670 & ~n9671;
  assign n9673 = ~n9393 & ~n9399;
  assign n9674 = n1434 & n5008;
  assign n9675 = pi79  & n5241;
  assign n9676 = pi81  & n5006;
  assign n9677 = pi80  & n5001;
  assign n9678 = ~n9676 & ~n9677;
  assign n9679 = ~n9675 & n9678;
  assign n9680 = ~n9674 & n9679;
  assign n9681 = pi38  & ~n9680;
  assign n9682 = pi38  & ~n9681;
  assign n9683 = ~n9680 & ~n9681;
  assign n9684 = ~n9682 & ~n9683;
  assign n9685 = ~n9377 & ~n9379;
  assign n9686 = n809 & n6539;
  assign n9687 = pi73  & n6873;
  assign n9688 = pi75  & n6537;
  assign n9689 = pi74  & n6532;
  assign n9690 = ~n9688 & ~n9689;
  assign n9691 = ~n9687 & n9690;
  assign n9692 = ~n9686 & n9691;
  assign n9693 = pi44  & ~n9692;
  assign n9694 = pi44  & ~n9693;
  assign n9695 = ~n9692 & ~n9693;
  assign n9696 = ~n9694 & ~n9695;
  assign n9697 = ~n9338 & ~n9344;
  assign n9698 = ~n9322 & ~n9324;
  assign n9699 = n286 & n9310;
  assign n9700 = n9019 & n9302;
  assign n9701 = ~n9307 & n9700;
  assign n9702 = pi64  & n9701;
  assign n9703 = pi66  & n9308;
  assign n9704 = pi65  & n9303;
  assign n9705 = ~n9703 & ~n9704;
  assign n9706 = ~n9699 & n9705;
  assign n9707 = ~n9702 & n9706;
  assign n9708 = pi53  & ~n9707;
  assign n9709 = pi53  & ~n9708;
  assign n9710 = ~n9707 & ~n9708;
  assign n9711 = ~n9709 & ~n9710;
  assign n9712 = ~n9318 & n9711;
  assign n9713 = n9318 & ~n9711;
  assign n9714 = ~n9712 & ~n9713;
  assign n9715 = n401 & n8334;
  assign n9716 = pi67  & n8685;
  assign n9717 = pi69  & n8332;
  assign n9718 = pi68  & n8327;
  assign n9719 = ~n9717 & ~n9718;
  assign n9720 = ~n9716 & n9719;
  assign n9721 = ~n9715 & n9720;
  assign n9722 = pi50  & ~n9721;
  assign n9723 = pi50  & ~n9722;
  assign n9724 = ~n9721 & ~n9722;
  assign n9725 = ~n9723 & ~n9724;
  assign n9726 = n9714 & ~n9725;
  assign n9727 = ~n9714 & n9725;
  assign n9728 = ~n9726 & ~n9727;
  assign n9729 = ~n9698 & n9728;
  assign n9730 = ~n9698 & ~n9729;
  assign n9731 = ~n9726 & ~n9729;
  assign n9732 = ~n9727 & n9731;
  assign n9733 = ~n9730 & ~n9732;
  assign n9734 = n576 & n7408;
  assign n9735 = pi70  & n7740;
  assign n9736 = pi72  & n7406;
  assign n9737 = pi71  & n7401;
  assign n9738 = ~n9736 & ~n9737;
  assign n9739 = ~n9735 & n9738;
  assign n9740 = ~n9734 & n9739;
  assign n9741 = pi47  & ~n9740;
  assign n9742 = pi47  & ~n9741;
  assign n9743 = ~n9740 & ~n9741;
  assign n9744 = ~n9742 & ~n9743;
  assign n9745 = n9733 & n9744;
  assign n9746 = ~n9733 & ~n9744;
  assign n9747 = ~n9745 & ~n9746;
  assign n9748 = ~n9697 & n9747;
  assign n9749 = n9697 & ~n9747;
  assign n9750 = ~n9748 & ~n9749;
  assign n9751 = n9696 & ~n9750;
  assign n9752 = ~n9696 & n9750;
  assign n9753 = ~n9751 & ~n9752;
  assign n9754 = ~n9362 & n9753;
  assign n9755 = n9362 & ~n9753;
  assign n9756 = ~n9754 & ~n9755;
  assign n9757 = n1025 & n5739;
  assign n9758 = pi76  & n6030;
  assign n9759 = pi78  & n5737;
  assign n9760 = pi77  & n5732;
  assign n9761 = ~n9759 & ~n9760;
  assign n9762 = ~n9758 & n9761;
  assign n9763 = ~n9757 & n9762;
  assign n9764 = pi41  & ~n9763;
  assign n9765 = pi41  & ~n9764;
  assign n9766 = ~n9763 & ~n9764;
  assign n9767 = ~n9765 & ~n9766;
  assign n9768 = n9756 & ~n9767;
  assign n9769 = n9756 & ~n9768;
  assign n9770 = ~n9767 & ~n9768;
  assign n9771 = ~n9769 & ~n9770;
  assign n9772 = ~n9685 & ~n9771;
  assign n9773 = n9685 & n9771;
  assign n9774 = ~n9772 & ~n9773;
  assign n9775 = ~n9684 & n9774;
  assign n9776 = ~n9684 & ~n9775;
  assign n9777 = n9774 & ~n9775;
  assign n9778 = ~n9776 & ~n9777;
  assign n9779 = ~n9673 & ~n9778;
  assign n9780 = ~n9673 & ~n9779;
  assign n9781 = ~n9778 & ~n9779;
  assign n9782 = ~n9780 & ~n9781;
  assign n9783 = n1834 & n4271;
  assign n9784 = pi82  & n4503;
  assign n9785 = pi84  & n4269;
  assign n9786 = pi83  & n4264;
  assign n9787 = ~n9785 & ~n9786;
  assign n9788 = ~n9784 & n9787;
  assign n9789 = ~n9783 & n9788;
  assign n9790 = pi35  & ~n9789;
  assign n9791 = pi35  & ~n9790;
  assign n9792 = ~n9789 & ~n9790;
  assign n9793 = ~n9791 & ~n9792;
  assign n9794 = ~n9782 & ~n9793;
  assign n9795 = ~n9782 & ~n9794;
  assign n9796 = ~n9793 & ~n9794;
  assign n9797 = ~n9795 & ~n9796;
  assign n9798 = ~n9417 & ~n9797;
  assign n9799 = n9417 & n9797;
  assign n9800 = ~n9798 & ~n9799;
  assign n9801 = ~n9672 & n9800;
  assign n9802 = ~n9672 & ~n9801;
  assign n9803 = n9800 & ~n9801;
  assign n9804 = ~n9802 & ~n9803;
  assign n9805 = ~n9661 & ~n9804;
  assign n9806 = ~n9661 & ~n9805;
  assign n9807 = ~n9804 & ~n9805;
  assign n9808 = ~n9806 & ~n9807;
  assign n9809 = n2801 & n3034;
  assign n9810 = pi88  & n3225;
  assign n9811 = pi90  & n3032;
  assign n9812 = pi89  & n3027;
  assign n9813 = ~n9811 & ~n9812;
  assign n9814 = ~n9810 & n9813;
  assign n9815 = ~n9809 & n9814;
  assign n9816 = pi29  & ~n9815;
  assign n9817 = pi29  & ~n9816;
  assign n9818 = ~n9815 & ~n9816;
  assign n9819 = ~n9817 & ~n9818;
  assign n9820 = n9808 & n9819;
  assign n9821 = ~n9808 & ~n9819;
  assign n9822 = ~n9820 & ~n9821;
  assign n9823 = ~n9660 & n9822;
  assign n9824 = n9660 & ~n9822;
  assign n9825 = ~n9823 & ~n9824;
  assign n9826 = n9658 & ~n9825;
  assign n9827 = ~n9658 & n9825;
  assign n9828 = ~n9826 & ~n9827;
  assign n9829 = ~n9647 & n9828;
  assign n9830 = n9647 & ~n9828;
  assign n9831 = ~n9829 & ~n9830;
  assign n9832 = n9646 & ~n9831;
  assign n9833 = ~n9646 & n9831;
  assign n9834 = ~n9832 & ~n9833;
  assign n9835 = ~n9635 & n9834;
  assign n9836 = n9635 & ~n9834;
  assign n9837 = ~n9835 & ~n9836;
  assign n9838 = n1611 & n4684;
  assign n9839 = pi97  & n1745;
  assign n9840 = pi99  & n1609;
  assign n9841 = pi98  & n1604;
  assign n9842 = ~n9840 & ~n9841;
  assign n9843 = ~n9839 & n9842;
  assign n9844 = ~n9838 & n9843;
  assign n9845 = pi20  & ~n9844;
  assign n9846 = pi20  & ~n9845;
  assign n9847 = ~n9844 & ~n9845;
  assign n9848 = ~n9846 & ~n9847;
  assign n9849 = n9837 & ~n9848;
  assign n9850 = n9837 & ~n9849;
  assign n9851 = ~n9848 & ~n9849;
  assign n9852 = ~n9850 & ~n9851;
  assign n9853 = ~n9504 & ~n9511;
  assign n9854 = n9852 & n9853;
  assign n9855 = ~n9852 & ~n9853;
  assign n9856 = ~n9854 & ~n9855;
  assign n9857 = n1297 & n5413;
  assign n9858 = pi100  & n1366;
  assign n9859 = pi102  & n1295;
  assign n9860 = pi101  & n1290;
  assign n9861 = ~n9859 & ~n9860;
  assign n9862 = ~n9858 & n9861;
  assign n9863 = ~n9857 & n9862;
  assign n9864 = pi17  & ~n9863;
  assign n9865 = pi17  & ~n9864;
  assign n9866 = ~n9863 & ~n9864;
  assign n9867 = ~n9865 & ~n9866;
  assign n9868 = n9856 & ~n9867;
  assign n9869 = n9856 & ~n9868;
  assign n9870 = ~n9867 & ~n9868;
  assign n9871 = ~n9869 & ~n9870;
  assign n9872 = ~n9524 & ~n9530;
  assign n9873 = n9871 & n9872;
  assign n9874 = ~n9871 & ~n9872;
  assign n9875 = ~n9873 & ~n9874;
  assign n9876 = n938 & n6207;
  assign n9877 = pi103  & n1052;
  assign n9878 = pi105  & n936;
  assign n9879 = pi104  & n931;
  assign n9880 = ~n9878 & ~n9879;
  assign n9881 = ~n9877 & n9880;
  assign n9882 = ~n9876 & n9881;
  assign n9883 = pi14  & ~n9882;
  assign n9884 = pi14  & ~n9883;
  assign n9885 = ~n9882 & ~n9883;
  assign n9886 = ~n9884 & ~n9885;
  assign n9887 = n9875 & ~n9886;
  assign n9888 = n9875 & ~n9887;
  assign n9889 = ~n9886 & ~n9887;
  assign n9890 = ~n9888 & ~n9889;
  assign n9891 = ~n9543 & ~n9549;
  assign n9892 = n9890 & n9891;
  assign n9893 = ~n9890 & ~n9891;
  assign n9894 = ~n9892 & ~n9893;
  assign n9895 = n687 & n7060;
  assign n9896 = pi106  & n763;
  assign n9897 = pi108  & n685;
  assign n9898 = pi107  & n680;
  assign n9899 = ~n9897 & ~n9898;
  assign n9900 = ~n9896 & n9899;
  assign n9901 = ~n9895 & n9900;
  assign n9902 = pi11  & ~n9901;
  assign n9903 = pi11  & ~n9902;
  assign n9904 = ~n9901 & ~n9902;
  assign n9905 = ~n9903 & ~n9904;
  assign n9906 = n9894 & ~n9905;
  assign n9907 = ~n9894 & n9905;
  assign n9908 = ~n9906 & ~n9907;
  assign n9909 = ~n9567 & n9908;
  assign n9910 = ~n9567 & ~n9909;
  assign n9911 = ~n9906 & ~n9909;
  assign n9912 = ~n9907 & n9911;
  assign n9913 = ~n9910 & ~n9912;
  assign n9914 = n498 & n7970;
  assign n9915 = pi109  & n537;
  assign n9916 = pi111  & n496;
  assign n9917 = pi110  & n491;
  assign n9918 = ~n9916 & ~n9917;
  assign n9919 = ~n9915 & n9918;
  assign n9920 = ~n9914 & n9919;
  assign n9921 = pi8  & ~n9920;
  assign n9922 = pi8  & ~n9921;
  assign n9923 = ~n9920 & ~n9921;
  assign n9924 = ~n9922 & ~n9923;
  assign n9925 = ~n9913 & ~n9924;
  assign n9926 = ~n9913 & ~n9925;
  assign n9927 = ~n9924 & ~n9925;
  assign n9928 = ~n9926 & ~n9927;
  assign n9929 = ~n9581 & ~n9588;
  assign n9930 = n9928 & n9929;
  assign n9931 = ~n9928 & ~n9929;
  assign n9932 = ~n9930 & ~n9931;
  assign n9933 = n342 & n8936;
  assign n9934 = pi112  & n380;
  assign n9935 = pi114  & n340;
  assign n9936 = pi113  & n335;
  assign n9937 = ~n9935 & ~n9936;
  assign n9938 = ~n9934 & n9937;
  assign n9939 = ~n9933 & n9938;
  assign n9940 = pi5  & ~n9939;
  assign n9941 = pi5  & ~n9940;
  assign n9942 = ~n9939 & ~n9940;
  assign n9943 = ~n9941 & ~n9942;
  assign n9944 = n9932 & ~n9943;
  assign n9945 = ~n9932 & n9943;
  assign n9946 = ~n9944 & ~n9945;
  assign n9947 = ~n9634 & n9946;
  assign n9948 = ~n9634 & ~n9947;
  assign n9949 = ~n9944 & ~n9947;
  assign n9950 = ~n9945 & n9949;
  assign n9951 = ~n9948 & ~n9950;
  assign n9952 = ~n9610 & ~n9612;
  assign n9953 = ~pi116  & ~pi117 ;
  assign n9954 = pi116  & pi117 ;
  assign n9955 = ~n9953 & ~n9954;
  assign n9956 = ~n9952 & n9955;
  assign n9957 = n9952 & ~n9955;
  assign n9958 = ~n9956 & ~n9957;
  assign n9959 = n262 & n9958;
  assign n9960 = pi115  & n288;
  assign n9961 = pi117  & n267;
  assign n9962 = pi116  & n269;
  assign n9963 = ~n9961 & ~n9962;
  assign n9964 = ~n9960 & n9963;
  assign n9965 = ~n9959 & n9964;
  assign n9966 = pi2  & ~n9965;
  assign n9967 = pi2  & ~n9966;
  assign n9968 = ~n9965 & ~n9966;
  assign n9969 = ~n9967 & ~n9968;
  assign n9970 = ~n9951 & n9969;
  assign n9971 = n9951 & ~n9969;
  assign n9972 = ~n9970 & ~n9971;
  assign n9973 = ~n9632 & ~n9972;
  assign n9974 = n9632 & n9972;
  assign po53  = ~n9973 & ~n9974;
  assign n9976 = ~n9951 & ~n9969;
  assign n9977 = ~n9973 & ~n9976;
  assign n9978 = ~n9954 & ~n9956;
  assign n9979 = ~pi117  & ~pi118 ;
  assign n9980 = pi117  & pi118 ;
  assign n9981 = ~n9979 & ~n9980;
  assign n9982 = ~n9978 & n9981;
  assign n9983 = n9978 & ~n9981;
  assign n9984 = ~n9982 & ~n9983;
  assign n9985 = n262 & n9984;
  assign n9986 = pi116  & n288;
  assign n9987 = pi118  & n267;
  assign n9988 = pi117  & n269;
  assign n9989 = ~n9987 & ~n9988;
  assign n9990 = ~n9986 & n9989;
  assign n9991 = ~n9985 & n9990;
  assign n9992 = pi2  & ~n9991;
  assign n9993 = pi2  & ~n9992;
  assign n9994 = ~n9991 & ~n9992;
  assign n9995 = ~n9993 & ~n9994;
  assign n9996 = n687 & n7349;
  assign n9997 = pi107  & n763;
  assign n9998 = pi109  & n685;
  assign n9999 = pi108  & n680;
  assign n10000 = ~n9998 & ~n9999;
  assign n10001 = ~n9997 & n10000;
  assign n10002 = ~n9996 & n10001;
  assign n10003 = pi11  & ~n10002;
  assign n10004 = pi11  & ~n10003;
  assign n10005 = ~n10002 & ~n10003;
  assign n10006 = ~n10004 & ~n10005;
  assign n10007 = ~n9887 & ~n9893;
  assign n10008 = ~n9849 & ~n9855;
  assign n10009 = ~n9833 & ~n9835;
  assign n10010 = ~n9827 & ~n9829;
  assign n10011 = n2523 & n3565;
  assign n10012 = pi92  & n2667;
  assign n10013 = pi94  & n2521;
  assign n10014 = pi93  & n2516;
  assign n10015 = ~n10013 & ~n10014;
  assign n10016 = ~n10012 & n10015;
  assign n10017 = ~n10011 & n10016;
  assign n10018 = pi26  & ~n10017;
  assign n10019 = pi26  & ~n10018;
  assign n10020 = ~n10017 & ~n10018;
  assign n10021 = ~n10019 & ~n10020;
  assign n10022 = ~n9821 & ~n9823;
  assign n10023 = n2978 & n3034;
  assign n10024 = pi89  & n3225;
  assign n10025 = pi91  & n3032;
  assign n10026 = pi90  & n3027;
  assign n10027 = ~n10025 & ~n10026;
  assign n10028 = ~n10024 & n10027;
  assign n10029 = ~n10023 & n10028;
  assign n10030 = pi29  & ~n10029;
  assign n10031 = pi29  & ~n10030;
  assign n10032 = ~n10029 & ~n10030;
  assign n10033 = ~n10031 & ~n10032;
  assign n10034 = ~n9801 & ~n9805;
  assign n10035 = n2446 & n3622;
  assign n10036 = pi86  & n3814;
  assign n10037 = pi88  & n3620;
  assign n10038 = pi87  & n3615;
  assign n10039 = ~n10037 & ~n10038;
  assign n10040 = ~n10036 & n10039;
  assign n10041 = ~n10035 & n10040;
  assign n10042 = pi32  & ~n10041;
  assign n10043 = pi32  & ~n10042;
  assign n10044 = ~n10041 & ~n10042;
  assign n10045 = ~n10043 & ~n10044;
  assign n10046 = ~n9794 & ~n9798;
  assign n10047 = n1972 & n4271;
  assign n10048 = pi83  & n4503;
  assign n10049 = pi85  & n4269;
  assign n10050 = pi84  & n4264;
  assign n10051 = ~n10049 & ~n10050;
  assign n10052 = ~n10048 & n10051;
  assign n10053 = ~n10047 & n10052;
  assign n10054 = pi35  & ~n10053;
  assign n10055 = pi35  & ~n10054;
  assign n10056 = ~n10053 & ~n10054;
  assign n10057 = ~n10055 & ~n10056;
  assign n10058 = ~n9775 & ~n9779;
  assign n10059 = n1554 & n5008;
  assign n10060 = pi80  & n5241;
  assign n10061 = pi82  & n5006;
  assign n10062 = pi81  & n5001;
  assign n10063 = ~n10061 & ~n10062;
  assign n10064 = ~n10060 & n10063;
  assign n10065 = ~n10059 & n10064;
  assign n10066 = pi38  & ~n10065;
  assign n10067 = pi38  & ~n10066;
  assign n10068 = ~n10065 & ~n10066;
  assign n10069 = ~n10067 & ~n10068;
  assign n10070 = ~n9768 & ~n9772;
  assign n10071 = n1122 & n5739;
  assign n10072 = pi77  & n6030;
  assign n10073 = pi79  & n5737;
  assign n10074 = pi78  & n5732;
  assign n10075 = ~n10073 & ~n10074;
  assign n10076 = ~n10072 & n10075;
  assign n10077 = ~n10071 & n10076;
  assign n10078 = pi41  & ~n10077;
  assign n10079 = pi41  & ~n10078;
  assign n10080 = ~n10077 & ~n10078;
  assign n10081 = ~n10079 & ~n10080;
  assign n10082 = ~n9752 & ~n9754;
  assign n10083 = n891 & n6539;
  assign n10084 = pi74  & n6873;
  assign n10085 = pi76  & n6537;
  assign n10086 = pi75  & n6532;
  assign n10087 = ~n10085 & ~n10086;
  assign n10088 = ~n10084 & n10087;
  assign n10089 = ~n10083 & n10088;
  assign n10090 = pi44  & ~n10089;
  assign n10091 = pi44  & ~n10090;
  assign n10092 = ~n10089 & ~n10090;
  assign n10093 = ~n10091 & ~n10092;
  assign n10094 = ~n9746 & ~n9748;
  assign n10095 = n642 & n7408;
  assign n10096 = pi71  & n7740;
  assign n10097 = pi73  & n7406;
  assign n10098 = pi72  & n7401;
  assign n10099 = ~n10097 & ~n10098;
  assign n10100 = ~n10096 & n10099;
  assign n10101 = ~n10095 & n10100;
  assign n10102 = pi47  & ~n10101;
  assign n10103 = pi47  & ~n10102;
  assign n10104 = ~n10101 & ~n10102;
  assign n10105 = ~n10103 & ~n10104;
  assign n10106 = pi53  & ~pi54 ;
  assign n10107 = ~pi53  & pi54 ;
  assign n10108 = ~n10106 & ~n10107;
  assign n10109 = pi64  & ~n10108;
  assign n10110 = ~n9713 & n10109;
  assign n10111 = n9713 & ~n10109;
  assign n10112 = ~n10110 & ~n10111;
  assign n10113 = n309 & n9310;
  assign n10114 = pi65  & n9701;
  assign n10115 = pi67  & n9308;
  assign n10116 = pi66  & n9303;
  assign n10117 = ~n10115 & ~n10116;
  assign n10118 = ~n10114 & n10117;
  assign n10119 = ~n10113 & n10118;
  assign n10120 = pi53  & ~n10119;
  assign n10121 = pi53  & ~n10120;
  assign n10122 = ~n10119 & ~n10120;
  assign n10123 = ~n10121 & ~n10122;
  assign n10124 = ~n10112 & ~n10123;
  assign n10125 = n10112 & n10123;
  assign n10126 = ~n10124 & ~n10125;
  assign n10127 = n450 & n8334;
  assign n10128 = pi68  & n8685;
  assign n10129 = pi70  & n8332;
  assign n10130 = pi69  & n8327;
  assign n10131 = ~n10129 & ~n10130;
  assign n10132 = ~n10128 & n10131;
  assign n10133 = ~n10127 & n10132;
  assign n10134 = pi50  & ~n10133;
  assign n10135 = pi50  & ~n10134;
  assign n10136 = ~n10133 & ~n10134;
  assign n10137 = ~n10135 & ~n10136;
  assign n10138 = n10126 & ~n10137;
  assign n10139 = n10126 & ~n10138;
  assign n10140 = ~n10137 & ~n10138;
  assign n10141 = ~n10139 & ~n10140;
  assign n10142 = ~n9731 & ~n10141;
  assign n10143 = n9731 & n10141;
  assign n10144 = ~n10142 & ~n10143;
  assign n10145 = ~n10105 & n10144;
  assign n10146 = ~n10105 & ~n10145;
  assign n10147 = n10144 & ~n10145;
  assign n10148 = ~n10146 & ~n10147;
  assign n10149 = ~n10094 & ~n10148;
  assign n10150 = n10094 & n10148;
  assign n10151 = ~n10149 & ~n10150;
  assign n10152 = ~n10093 & n10151;
  assign n10153 = ~n10093 & ~n10152;
  assign n10154 = n10151 & ~n10152;
  assign n10155 = ~n10153 & ~n10154;
  assign n10156 = ~n10082 & ~n10155;
  assign n10157 = n10082 & n10155;
  assign n10158 = ~n10156 & ~n10157;
  assign n10159 = ~n10081 & n10158;
  assign n10160 = n10081 & ~n10158;
  assign n10161 = ~n10159 & ~n10160;
  assign n10162 = ~n10070 & n10161;
  assign n10163 = n10070 & ~n10161;
  assign n10164 = ~n10162 & ~n10163;
  assign n10165 = ~n10069 & n10164;
  assign n10166 = ~n10069 & ~n10165;
  assign n10167 = n10164 & ~n10165;
  assign n10168 = ~n10166 & ~n10167;
  assign n10169 = ~n10058 & ~n10168;
  assign n10170 = n10058 & n10168;
  assign n10171 = ~n10169 & ~n10170;
  assign n10172 = ~n10057 & n10171;
  assign n10173 = n10057 & ~n10171;
  assign n10174 = ~n10172 & ~n10173;
  assign n10175 = ~n10046 & n10174;
  assign n10176 = n10046 & ~n10174;
  assign n10177 = ~n10175 & ~n10176;
  assign n10178 = ~n10045 & n10177;
  assign n10179 = n10045 & ~n10177;
  assign n10180 = ~n10178 & ~n10179;
  assign n10181 = ~n10034 & n10180;
  assign n10182 = n10034 & ~n10180;
  assign n10183 = ~n10181 & ~n10182;
  assign n10184 = ~n10033 & n10183;
  assign n10185 = n10033 & ~n10183;
  assign n10186 = ~n10184 & ~n10185;
  assign n10187 = ~n10022 & n10186;
  assign n10188 = n10022 & ~n10186;
  assign n10189 = ~n10187 & ~n10188;
  assign n10190 = ~n10021 & n10189;
  assign n10191 = n10021 & ~n10189;
  assign n10192 = ~n10190 & ~n10191;
  assign n10193 = ~n10010 & n10192;
  assign n10194 = n10010 & ~n10192;
  assign n10195 = ~n10193 & ~n10194;
  assign n10196 = n2043 & n4211;
  assign n10197 = pi95  & n2180;
  assign n10198 = pi97  & n2041;
  assign n10199 = pi96  & n2036;
  assign n10200 = ~n10198 & ~n10199;
  assign n10201 = ~n10197 & n10200;
  assign n10202 = ~n10196 & n10201;
  assign n10203 = pi23  & ~n10202;
  assign n10204 = pi23  & ~n10203;
  assign n10205 = ~n10202 & ~n10203;
  assign n10206 = ~n10204 & ~n10205;
  assign n10207 = n10195 & ~n10206;
  assign n10208 = n10195 & ~n10207;
  assign n10209 = ~n10206 & ~n10207;
  assign n10210 = ~n10208 & ~n10209;
  assign n10211 = ~n10009 & n10210;
  assign n10212 = n10009 & ~n10210;
  assign n10213 = ~n10211 & ~n10212;
  assign n10214 = n1611 & n4910;
  assign n10215 = pi98  & n1745;
  assign n10216 = pi100  & n1609;
  assign n10217 = pi99  & n1604;
  assign n10218 = ~n10216 & ~n10217;
  assign n10219 = ~n10215 & n10218;
  assign n10220 = ~n10214 & n10219;
  assign n10221 = pi20  & ~n10220;
  assign n10222 = pi20  & ~n10221;
  assign n10223 = ~n10220 & ~n10221;
  assign n10224 = ~n10222 & ~n10223;
  assign n10225 = ~n10213 & ~n10224;
  assign n10226 = n10213 & n10224;
  assign n10227 = ~n10225 & ~n10226;
  assign n10228 = n10008 & ~n10227;
  assign n10229 = ~n10008 & n10227;
  assign n10230 = ~n10228 & ~n10229;
  assign n10231 = n1297 & n5664;
  assign n10232 = pi101  & n1366;
  assign n10233 = pi103  & n1295;
  assign n10234 = pi102  & n1290;
  assign n10235 = ~n10233 & ~n10234;
  assign n10236 = ~n10232 & n10235;
  assign n10237 = ~n10231 & n10236;
  assign n10238 = pi17  & ~n10237;
  assign n10239 = pi17  & ~n10238;
  assign n10240 = ~n10237 & ~n10238;
  assign n10241 = ~n10239 & ~n10240;
  assign n10242 = n10230 & ~n10241;
  assign n10243 = n10230 & ~n10242;
  assign n10244 = ~n10241 & ~n10242;
  assign n10245 = ~n10243 & ~n10244;
  assign n10246 = ~n9868 & ~n9874;
  assign n10247 = n10245 & n10246;
  assign n10248 = ~n10245 & ~n10246;
  assign n10249 = ~n10247 & ~n10248;
  assign n10250 = n938 & n6477;
  assign n10251 = pi104  & n1052;
  assign n10252 = pi106  & n936;
  assign n10253 = pi105  & n931;
  assign n10254 = ~n10252 & ~n10253;
  assign n10255 = ~n10251 & n10254;
  assign n10256 = ~n10250 & n10255;
  assign n10257 = pi14  & ~n10256;
  assign n10258 = pi14  & ~n10257;
  assign n10259 = ~n10256 & ~n10257;
  assign n10260 = ~n10258 & ~n10259;
  assign n10261 = ~n10249 & n10260;
  assign n10262 = n10249 & ~n10260;
  assign n10263 = ~n10261 & ~n10262;
  assign n10264 = ~n10007 & n10263;
  assign n10265 = n10007 & ~n10263;
  assign n10266 = ~n10264 & ~n10265;
  assign n10267 = ~n10006 & n10266;
  assign n10268 = ~n10006 & ~n10267;
  assign n10269 = n10266 & ~n10267;
  assign n10270 = ~n10268 & ~n10269;
  assign n10271 = ~n9911 & ~n10270;
  assign n10272 = ~n9911 & ~n10271;
  assign n10273 = ~n10270 & ~n10271;
  assign n10274 = ~n10272 & ~n10273;
  assign n10275 = n498 & n7997;
  assign n10276 = pi110  & n537;
  assign n10277 = pi112  & n496;
  assign n10278 = pi111  & n491;
  assign n10279 = ~n10277 & ~n10278;
  assign n10280 = ~n10276 & n10279;
  assign n10281 = ~n10275 & n10280;
  assign n10282 = pi8  & ~n10281;
  assign n10283 = pi8  & ~n10282;
  assign n10284 = ~n10281 & ~n10282;
  assign n10285 = ~n10283 & ~n10284;
  assign n10286 = ~n10274 & ~n10285;
  assign n10287 = ~n10274 & ~n10286;
  assign n10288 = ~n10285 & ~n10286;
  assign n10289 = ~n10287 & ~n10288;
  assign n10290 = ~n9925 & ~n9931;
  assign n10291 = n10289 & n10290;
  assign n10292 = ~n10289 & ~n10290;
  assign n10293 = ~n10291 & ~n10292;
  assign n10294 = n342 & n8963;
  assign n10295 = pi113  & n380;
  assign n10296 = pi115  & n340;
  assign n10297 = pi114  & n335;
  assign n10298 = ~n10296 & ~n10297;
  assign n10299 = ~n10295 & n10298;
  assign n10300 = ~n10294 & n10299;
  assign n10301 = pi5  & ~n10300;
  assign n10302 = pi5  & ~n10301;
  assign n10303 = ~n10300 & ~n10301;
  assign n10304 = ~n10302 & ~n10303;
  assign n10305 = ~n10293 & n10304;
  assign n10306 = n10293 & ~n10304;
  assign n10307 = ~n10305 & ~n10306;
  assign n10308 = ~n9949 & n10307;
  assign n10309 = n9949 & ~n10307;
  assign n10310 = ~n10308 & ~n10309;
  assign n10311 = ~n9995 & n10310;
  assign n10312 = n9995 & ~n10310;
  assign n10313 = ~n10311 & ~n10312;
  assign n10314 = ~n9977 & n10313;
  assign n10315 = n9977 & ~n10313;
  assign po54  = ~n10314 & ~n10315;
  assign n10317 = ~n10311 & ~n10314;
  assign n10318 = ~n10306 & ~n10308;
  assign n10319 = ~n10286 & ~n10292;
  assign n10320 = n498 & n8612;
  assign n10321 = pi111  & n537;
  assign n10322 = pi113  & n496;
  assign n10323 = pi112  & n491;
  assign n10324 = ~n10322 & ~n10323;
  assign n10325 = ~n10321 & n10324;
  assign n10326 = ~n10320 & n10325;
  assign n10327 = pi8  & ~n10326;
  assign n10328 = pi8  & ~n10327;
  assign n10329 = ~n10326 & ~n10327;
  assign n10330 = ~n10328 & ~n10329;
  assign n10331 = ~n10267 & ~n10271;
  assign n10332 = ~n10262 & ~n10264;
  assign n10333 = ~n10165 & ~n10169;
  assign n10334 = ~n10152 & ~n10156;
  assign n10335 = n999 & n6539;
  assign n10336 = pi75  & n6873;
  assign n10337 = pi77  & n6537;
  assign n10338 = pi76  & n6532;
  assign n10339 = ~n10337 & ~n10338;
  assign n10340 = ~n10336 & n10339;
  assign n10341 = ~n10335 & n10340;
  assign n10342 = pi44  & ~n10341;
  assign n10343 = pi44  & ~n10342;
  assign n10344 = ~n10341 & ~n10342;
  assign n10345 = ~n10343 & ~n10344;
  assign n10346 = ~n10145 & ~n10149;
  assign n10347 = n729 & n7408;
  assign n10348 = pi72  & n7740;
  assign n10349 = pi74  & n7406;
  assign n10350 = pi73  & n7401;
  assign n10351 = ~n10349 & ~n10350;
  assign n10352 = ~n10348 & n10351;
  assign n10353 = ~n10347 & n10352;
  assign n10354 = pi47  & ~n10353;
  assign n10355 = pi47  & ~n10354;
  assign n10356 = ~n10353 & ~n10354;
  assign n10357 = ~n10355 & ~n10356;
  assign n10358 = ~n10138 & ~n10142;
  assign n10359 = n475 & n8334;
  assign n10360 = pi69  & n8685;
  assign n10361 = pi71  & n8332;
  assign n10362 = pi70  & n8327;
  assign n10363 = ~n10361 & ~n10362;
  assign n10364 = ~n10360 & n10363;
  assign n10365 = ~n10359 & n10364;
  assign n10366 = pi50  & ~n10365;
  assign n10367 = pi50  & ~n10366;
  assign n10368 = ~n10365 & ~n10366;
  assign n10369 = ~n10367 & ~n10368;
  assign n10370 = n9713 & n10109;
  assign n10371 = ~n10124 & ~n10370;
  assign n10372 = n359 & n9310;
  assign n10373 = pi66  & n9701;
  assign n10374 = pi68  & n9308;
  assign n10375 = pi67  & n9303;
  assign n10376 = ~n10374 & ~n10375;
  assign n10377 = ~n10373 & n10376;
  assign n10378 = ~n10372 & n10377;
  assign n10379 = pi53  & ~n10378;
  assign n10380 = pi53  & ~n10379;
  assign n10381 = ~n10378 & ~n10379;
  assign n10382 = ~n10380 & ~n10381;
  assign n10383 = pi56  & ~n10109;
  assign n10384 = ~pi54  & pi55 ;
  assign n10385 = pi54  & ~pi55 ;
  assign n10386 = ~n10384 & ~n10385;
  assign n10387 = n10108 & ~n10386;
  assign n10388 = pi64  & n10387;
  assign n10389 = ~pi55  & pi56 ;
  assign n10390 = pi55  & ~pi56 ;
  assign n10391 = ~n10389 & ~n10390;
  assign n10392 = ~n10108 & n10391;
  assign n10393 = pi65  & n10392;
  assign n10394 = ~n10108 & ~n10391;
  assign n10395 = ~n265 & n10394;
  assign n10396 = ~n10388 & ~n10393;
  assign n10397 = ~n10395 & n10396;
  assign n10398 = pi56  & ~n10397;
  assign n10399 = pi56  & ~n10398;
  assign n10400 = ~n10397 & ~n10398;
  assign n10401 = ~n10399 & ~n10400;
  assign n10402 = n10383 & ~n10401;
  assign n10403 = ~n10383 & n10401;
  assign n10404 = ~n10402 & ~n10403;
  assign n10405 = n10382 & ~n10404;
  assign n10406 = ~n10382 & n10404;
  assign n10407 = ~n10405 & ~n10406;
  assign n10408 = ~n10371 & n10407;
  assign n10409 = n10371 & ~n10407;
  assign n10410 = ~n10408 & ~n10409;
  assign n10411 = n10369 & ~n10410;
  assign n10412 = ~n10369 & n10410;
  assign n10413 = ~n10411 & ~n10412;
  assign n10414 = ~n10358 & n10413;
  assign n10415 = n10358 & ~n10413;
  assign n10416 = ~n10414 & ~n10415;
  assign n10417 = n10357 & ~n10416;
  assign n10418 = ~n10357 & n10416;
  assign n10419 = ~n10417 & ~n10418;
  assign n10420 = ~n10346 & n10419;
  assign n10421 = n10346 & ~n10419;
  assign n10422 = ~n10420 & ~n10421;
  assign n10423 = n10345 & ~n10422;
  assign n10424 = ~n10345 & n10422;
  assign n10425 = ~n10423 & ~n10424;
  assign n10426 = ~n10334 & n10425;
  assign n10427 = n10334 & ~n10425;
  assign n10428 = ~n10426 & ~n10427;
  assign n10429 = n1225 & n5739;
  assign n10430 = pi78  & n6030;
  assign n10431 = pi80  & n5737;
  assign n10432 = pi79  & n5732;
  assign n10433 = ~n10431 & ~n10432;
  assign n10434 = ~n10430 & n10433;
  assign n10435 = ~n10429 & n10434;
  assign n10436 = pi41  & ~n10435;
  assign n10437 = pi41  & ~n10436;
  assign n10438 = ~n10435 & ~n10436;
  assign n10439 = ~n10437 & ~n10438;
  assign n10440 = n10428 & ~n10439;
  assign n10441 = n10428 & ~n10440;
  assign n10442 = ~n10439 & ~n10440;
  assign n10443 = ~n10441 & ~n10442;
  assign n10444 = ~n10159 & ~n10162;
  assign n10445 = n10443 & n10444;
  assign n10446 = ~n10443 & ~n10444;
  assign n10447 = ~n10445 & ~n10446;
  assign n10448 = n1696 & n5008;
  assign n10449 = pi81  & n5241;
  assign n10450 = pi83  & n5006;
  assign n10451 = pi82  & n5001;
  assign n10452 = ~n10450 & ~n10451;
  assign n10453 = ~n10449 & n10452;
  assign n10454 = ~n10448 & n10453;
  assign n10455 = pi38  & ~n10454;
  assign n10456 = pi38  & ~n10455;
  assign n10457 = ~n10454 & ~n10455;
  assign n10458 = ~n10456 & ~n10457;
  assign n10459 = n10447 & ~n10458;
  assign n10460 = ~n10447 & n10458;
  assign n10461 = ~n10459 & ~n10460;
  assign n10462 = ~n10333 & n10461;
  assign n10463 = ~n10333 & ~n10462;
  assign n10464 = ~n10459 & ~n10462;
  assign n10465 = ~n10460 & n10464;
  assign n10466 = ~n10463 & ~n10465;
  assign n10467 = n2133 & n4271;
  assign n10468 = pi84  & n4503;
  assign n10469 = pi86  & n4269;
  assign n10470 = pi85  & n4264;
  assign n10471 = ~n10469 & ~n10470;
  assign n10472 = ~n10468 & n10471;
  assign n10473 = ~n10467 & n10472;
  assign n10474 = pi35  & ~n10473;
  assign n10475 = pi35  & ~n10474;
  assign n10476 = ~n10473 & ~n10474;
  assign n10477 = ~n10475 & ~n10476;
  assign n10478 = ~n10466 & ~n10477;
  assign n10479 = ~n10466 & ~n10478;
  assign n10480 = ~n10477 & ~n10478;
  assign n10481 = ~n10479 & ~n10480;
  assign n10482 = ~n10172 & ~n10175;
  assign n10483 = n10481 & n10482;
  assign n10484 = ~n10481 & ~n10482;
  assign n10485 = ~n10483 & ~n10484;
  assign n10486 = n2473 & n3622;
  assign n10487 = pi87  & n3814;
  assign n10488 = pi89  & n3620;
  assign n10489 = pi88  & n3615;
  assign n10490 = ~n10488 & ~n10489;
  assign n10491 = ~n10487 & n10490;
  assign n10492 = ~n10486 & n10491;
  assign n10493 = pi32  & ~n10492;
  assign n10494 = pi32  & ~n10493;
  assign n10495 = ~n10492 & ~n10493;
  assign n10496 = ~n10494 & ~n10495;
  assign n10497 = n10485 & ~n10496;
  assign n10498 = n10485 & ~n10497;
  assign n10499 = ~n10496 & ~n10497;
  assign n10500 = ~n10498 & ~n10499;
  assign n10501 = ~n10178 & ~n10181;
  assign n10502 = n10500 & n10501;
  assign n10503 = ~n10500 & ~n10501;
  assign n10504 = ~n10502 & ~n10503;
  assign n10505 = n3034 & n3177;
  assign n10506 = pi90  & n3225;
  assign n10507 = pi92  & n3032;
  assign n10508 = pi91  & n3027;
  assign n10509 = ~n10507 & ~n10508;
  assign n10510 = ~n10506 & n10509;
  assign n10511 = ~n10505 & n10510;
  assign n10512 = pi29  & ~n10511;
  assign n10513 = pi29  & ~n10512;
  assign n10514 = ~n10511 & ~n10512;
  assign n10515 = ~n10513 & ~n10514;
  assign n10516 = n10504 & ~n10515;
  assign n10517 = n10504 & ~n10516;
  assign n10518 = ~n10515 & ~n10516;
  assign n10519 = ~n10517 & ~n10518;
  assign n10520 = ~n10184 & ~n10187;
  assign n10521 = n10519 & n10520;
  assign n10522 = ~n10519 & ~n10520;
  assign n10523 = ~n10521 & ~n10522;
  assign n10524 = n2523 & n3784;
  assign n10525 = pi93  & n2667;
  assign n10526 = pi95  & n2521;
  assign n10527 = pi94  & n2516;
  assign n10528 = ~n10526 & ~n10527;
  assign n10529 = ~n10525 & n10528;
  assign n10530 = ~n10524 & n10529;
  assign n10531 = pi26  & ~n10530;
  assign n10532 = pi26  & ~n10531;
  assign n10533 = ~n10530 & ~n10531;
  assign n10534 = ~n10532 & ~n10533;
  assign n10535 = n10523 & ~n10534;
  assign n10536 = n10523 & ~n10535;
  assign n10537 = ~n10534 & ~n10535;
  assign n10538 = ~n10536 & ~n10537;
  assign n10539 = ~n10190 & ~n10193;
  assign n10540 = n10538 & n10539;
  assign n10541 = ~n10538 & ~n10539;
  assign n10542 = ~n10540 & ~n10541;
  assign n10543 = n2043 & n4454;
  assign n10544 = pi96  & n2180;
  assign n10545 = pi98  & n2041;
  assign n10546 = pi97  & n2036;
  assign n10547 = ~n10545 & ~n10546;
  assign n10548 = ~n10544 & n10547;
  assign n10549 = ~n10543 & n10548;
  assign n10550 = pi23  & ~n10549;
  assign n10551 = pi23  & ~n10550;
  assign n10552 = ~n10549 & ~n10550;
  assign n10553 = ~n10551 & ~n10552;
  assign n10554 = n10542 & ~n10553;
  assign n10555 = n10542 & ~n10554;
  assign n10556 = ~n10553 & ~n10554;
  assign n10557 = ~n10555 & ~n10556;
  assign n10558 = ~n10009 & ~n10210;
  assign n10559 = ~n10207 & ~n10558;
  assign n10560 = n10557 & n10559;
  assign n10561 = ~n10557 & ~n10559;
  assign n10562 = ~n10560 & ~n10561;
  assign n10563 = n1611 & n5169;
  assign n10564 = pi99  & n1745;
  assign n10565 = pi101  & n1609;
  assign n10566 = pi100  & n1604;
  assign n10567 = ~n10565 & ~n10566;
  assign n10568 = ~n10564 & n10567;
  assign n10569 = ~n10563 & n10568;
  assign n10570 = pi20  & ~n10569;
  assign n10571 = pi20  & ~n10570;
  assign n10572 = ~n10569 & ~n10570;
  assign n10573 = ~n10571 & ~n10572;
  assign n10574 = n10562 & ~n10573;
  assign n10575 = n10562 & ~n10574;
  assign n10576 = ~n10573 & ~n10574;
  assign n10577 = ~n10575 & ~n10576;
  assign n10578 = ~n10225 & ~n10229;
  assign n10579 = n10577 & n10578;
  assign n10580 = ~n10577 & ~n10578;
  assign n10581 = ~n10579 & ~n10580;
  assign n10582 = n1297 & n5943;
  assign n10583 = pi102  & n1366;
  assign n10584 = pi104  & n1295;
  assign n10585 = pi103  & n1290;
  assign n10586 = ~n10584 & ~n10585;
  assign n10587 = ~n10583 & n10586;
  assign n10588 = ~n10582 & n10587;
  assign n10589 = pi17  & ~n10588;
  assign n10590 = pi17  & ~n10589;
  assign n10591 = ~n10588 & ~n10589;
  assign n10592 = ~n10590 & ~n10591;
  assign n10593 = n10581 & ~n10592;
  assign n10594 = n10581 & ~n10593;
  assign n10595 = ~n10592 & ~n10593;
  assign n10596 = ~n10594 & ~n10595;
  assign n10597 = ~n10242 & ~n10248;
  assign n10598 = n10596 & n10597;
  assign n10599 = ~n10596 & ~n10597;
  assign n10600 = ~n10598 & ~n10599;
  assign n10601 = n938 & n6775;
  assign n10602 = pi105  & n1052;
  assign n10603 = pi107  & n936;
  assign n10604 = pi106  & n931;
  assign n10605 = ~n10603 & ~n10604;
  assign n10606 = ~n10602 & n10605;
  assign n10607 = ~n10601 & n10606;
  assign n10608 = pi14  & ~n10607;
  assign n10609 = pi14  & ~n10608;
  assign n10610 = ~n10607 & ~n10608;
  assign n10611 = ~n10609 & ~n10610;
  assign n10612 = n10600 & ~n10611;
  assign n10613 = ~n10600 & n10611;
  assign n10614 = ~n10612 & ~n10613;
  assign n10615 = ~n10332 & n10614;
  assign n10616 = ~n10332 & ~n10615;
  assign n10617 = ~n10612 & ~n10615;
  assign n10618 = ~n10613 & n10617;
  assign n10619 = ~n10616 & ~n10618;
  assign n10620 = n687 & n7665;
  assign n10621 = pi108  & n763;
  assign n10622 = pi110  & n685;
  assign n10623 = pi109  & n680;
  assign n10624 = ~n10622 & ~n10623;
  assign n10625 = ~n10621 & n10624;
  assign n10626 = ~n10620 & n10625;
  assign n10627 = pi11  & ~n10626;
  assign n10628 = pi11  & ~n10627;
  assign n10629 = ~n10626 & ~n10627;
  assign n10630 = ~n10628 & ~n10629;
  assign n10631 = n10619 & n10630;
  assign n10632 = ~n10619 & ~n10630;
  assign n10633 = ~n10631 & ~n10632;
  assign n10634 = ~n10331 & n10633;
  assign n10635 = n10331 & ~n10633;
  assign n10636 = ~n10634 & ~n10635;
  assign n10637 = n10330 & ~n10636;
  assign n10638 = ~n10330 & n10636;
  assign n10639 = ~n10637 & ~n10638;
  assign n10640 = ~n10319 & n10639;
  assign n10641 = n10319 & ~n10639;
  assign n10642 = ~n10640 & ~n10641;
  assign n10643 = n342 & n9614;
  assign n10644 = pi114  & n380;
  assign n10645 = pi116  & n340;
  assign n10646 = pi115  & n335;
  assign n10647 = ~n10645 & ~n10646;
  assign n10648 = ~n10644 & n10647;
  assign n10649 = ~n10643 & n10648;
  assign n10650 = pi5  & ~n10649;
  assign n10651 = pi5  & ~n10650;
  assign n10652 = ~n10649 & ~n10650;
  assign n10653 = ~n10651 & ~n10652;
  assign n10654 = n10642 & ~n10653;
  assign n10655 = n10642 & ~n10654;
  assign n10656 = ~n10653 & ~n10654;
  assign n10657 = ~n10655 & ~n10656;
  assign n10658 = ~n10318 & n10657;
  assign n10659 = n10318 & ~n10657;
  assign n10660 = ~n10658 & ~n10659;
  assign n10661 = ~n9980 & ~n9982;
  assign n10662 = ~pi118  & ~pi119 ;
  assign n10663 = pi118  & pi119 ;
  assign n10664 = ~n10662 & ~n10663;
  assign n10665 = ~n10661 & n10664;
  assign n10666 = n10661 & ~n10664;
  assign n10667 = ~n10665 & ~n10666;
  assign n10668 = n262 & n10667;
  assign n10669 = pi117  & n288;
  assign n10670 = pi119  & n267;
  assign n10671 = pi118  & n269;
  assign n10672 = ~n10670 & ~n10671;
  assign n10673 = ~n10669 & n10672;
  assign n10674 = ~n10668 & n10673;
  assign n10675 = pi2  & ~n10674;
  assign n10676 = pi2  & ~n10675;
  assign n10677 = ~n10674 & ~n10675;
  assign n10678 = ~n10676 & ~n10677;
  assign n10679 = ~n10660 & ~n10678;
  assign n10680 = n10660 & n10678;
  assign n10681 = ~n10679 & ~n10680;
  assign n10682 = ~n10317 & n10681;
  assign n10683 = n10317 & ~n10681;
  assign po55  = ~n10682 & ~n10683;
  assign n10685 = ~n10318 & ~n10657;
  assign n10686 = ~n10654 & ~n10685;
  assign n10687 = ~n10638 & ~n10640;
  assign n10688 = n498 & n8936;
  assign n10689 = pi112  & n537;
  assign n10690 = pi114  & n496;
  assign n10691 = pi113  & n491;
  assign n10692 = ~n10690 & ~n10691;
  assign n10693 = ~n10689 & n10692;
  assign n10694 = ~n10688 & n10693;
  assign n10695 = pi8  & ~n10694;
  assign n10696 = pi8  & ~n10695;
  assign n10697 = ~n10694 & ~n10695;
  assign n10698 = ~n10696 & ~n10697;
  assign n10699 = ~n10632 & ~n10634;
  assign n10700 = ~n10535 & ~n10541;
  assign n10701 = n2523 & n4001;
  assign n10702 = pi94  & n2667;
  assign n10703 = pi96  & n2521;
  assign n10704 = pi95  & n2516;
  assign n10705 = ~n10703 & ~n10704;
  assign n10706 = ~n10702 & n10705;
  assign n10707 = ~n10701 & n10706;
  assign n10708 = pi26  & ~n10707;
  assign n10709 = pi26  & ~n10708;
  assign n10710 = ~n10707 & ~n10708;
  assign n10711 = ~n10709 & ~n10710;
  assign n10712 = ~n10516 & ~n10522;
  assign n10713 = ~n10497 & ~n10503;
  assign n10714 = ~n10478 & ~n10484;
  assign n10715 = ~n10440 & ~n10446;
  assign n10716 = n1434 & n5739;
  assign n10717 = pi79  & n6030;
  assign n10718 = pi81  & n5737;
  assign n10719 = pi80  & n5732;
  assign n10720 = ~n10718 & ~n10719;
  assign n10721 = ~n10717 & n10720;
  assign n10722 = ~n10716 & n10721;
  assign n10723 = pi41  & ~n10722;
  assign n10724 = pi41  & ~n10723;
  assign n10725 = ~n10722 & ~n10723;
  assign n10726 = ~n10724 & ~n10725;
  assign n10727 = ~n10424 & ~n10426;
  assign n10728 = ~n10418 & ~n10420;
  assign n10729 = n809 & n7408;
  assign n10730 = pi73  & n7740;
  assign n10731 = pi75  & n7406;
  assign n10732 = pi74  & n7401;
  assign n10733 = ~n10731 & ~n10732;
  assign n10734 = ~n10730 & n10733;
  assign n10735 = ~n10729 & n10734;
  assign n10736 = pi47  & ~n10735;
  assign n10737 = pi47  & ~n10736;
  assign n10738 = ~n10735 & ~n10736;
  assign n10739 = ~n10737 & ~n10738;
  assign n10740 = ~n10412 & ~n10414;
  assign n10741 = ~n10406 & ~n10408;
  assign n10742 = n286 & n10394;
  assign n10743 = n10108 & n10386;
  assign n10744 = ~n10391 & n10743;
  assign n10745 = pi64  & n10744;
  assign n10746 = pi66  & n10392;
  assign n10747 = pi65  & n10387;
  assign n10748 = ~n10746 & ~n10747;
  assign n10749 = ~n10742 & n10748;
  assign n10750 = ~n10745 & n10749;
  assign n10751 = pi56  & ~n10750;
  assign n10752 = pi56  & ~n10751;
  assign n10753 = ~n10750 & ~n10751;
  assign n10754 = ~n10752 & ~n10753;
  assign n10755 = ~n10402 & n10754;
  assign n10756 = n10402 & ~n10754;
  assign n10757 = ~n10755 & ~n10756;
  assign n10758 = n401 & n9310;
  assign n10759 = pi67  & n9701;
  assign n10760 = pi69  & n9308;
  assign n10761 = pi68  & n9303;
  assign n10762 = ~n10760 & ~n10761;
  assign n10763 = ~n10759 & n10762;
  assign n10764 = ~n10758 & n10763;
  assign n10765 = pi53  & ~n10764;
  assign n10766 = pi53  & ~n10765;
  assign n10767 = ~n10764 & ~n10765;
  assign n10768 = ~n10766 & ~n10767;
  assign n10769 = n10757 & ~n10768;
  assign n10770 = ~n10757 & n10768;
  assign n10771 = ~n10769 & ~n10770;
  assign n10772 = ~n10741 & n10771;
  assign n10773 = ~n10741 & ~n10772;
  assign n10774 = ~n10769 & ~n10772;
  assign n10775 = ~n10770 & n10774;
  assign n10776 = ~n10773 & ~n10775;
  assign n10777 = n576 & n8334;
  assign n10778 = pi70  & n8685;
  assign n10779 = pi72  & n8332;
  assign n10780 = pi71  & n8327;
  assign n10781 = ~n10779 & ~n10780;
  assign n10782 = ~n10778 & n10781;
  assign n10783 = ~n10777 & n10782;
  assign n10784 = pi50  & ~n10783;
  assign n10785 = pi50  & ~n10784;
  assign n10786 = ~n10783 & ~n10784;
  assign n10787 = ~n10785 & ~n10786;
  assign n10788 = n10776 & n10787;
  assign n10789 = ~n10776 & ~n10787;
  assign n10790 = ~n10788 & ~n10789;
  assign n10791 = ~n10740 & n10790;
  assign n10792 = n10740 & ~n10790;
  assign n10793 = ~n10791 & ~n10792;
  assign n10794 = n10739 & ~n10793;
  assign n10795 = ~n10739 & n10793;
  assign n10796 = ~n10794 & ~n10795;
  assign n10797 = ~n10728 & n10796;
  assign n10798 = n10728 & ~n10796;
  assign n10799 = ~n10797 & ~n10798;
  assign n10800 = n1025 & n6539;
  assign n10801 = pi76  & n6873;
  assign n10802 = pi78  & n6537;
  assign n10803 = pi77  & n6532;
  assign n10804 = ~n10802 & ~n10803;
  assign n10805 = ~n10801 & n10804;
  assign n10806 = ~n10800 & n10805;
  assign n10807 = pi44  & ~n10806;
  assign n10808 = pi44  & ~n10807;
  assign n10809 = ~n10806 & ~n10807;
  assign n10810 = ~n10808 & ~n10809;
  assign n10811 = n10799 & ~n10810;
  assign n10812 = n10799 & ~n10811;
  assign n10813 = ~n10810 & ~n10811;
  assign n10814 = ~n10812 & ~n10813;
  assign n10815 = ~n10727 & ~n10814;
  assign n10816 = n10727 & n10814;
  assign n10817 = ~n10815 & ~n10816;
  assign n10818 = ~n10726 & n10817;
  assign n10819 = ~n10726 & ~n10818;
  assign n10820 = n10817 & ~n10818;
  assign n10821 = ~n10819 & ~n10820;
  assign n10822 = ~n10715 & ~n10821;
  assign n10823 = ~n10715 & ~n10822;
  assign n10824 = ~n10821 & ~n10822;
  assign n10825 = ~n10823 & ~n10824;
  assign n10826 = n1834 & n5008;
  assign n10827 = pi82  & n5241;
  assign n10828 = pi84  & n5006;
  assign n10829 = pi83  & n5001;
  assign n10830 = ~n10828 & ~n10829;
  assign n10831 = ~n10827 & n10830;
  assign n10832 = ~n10826 & n10831;
  assign n10833 = pi38  & ~n10832;
  assign n10834 = pi38  & ~n10833;
  assign n10835 = ~n10832 & ~n10833;
  assign n10836 = ~n10834 & ~n10835;
  assign n10837 = ~n10825 & ~n10836;
  assign n10838 = ~n10825 & ~n10837;
  assign n10839 = ~n10836 & ~n10837;
  assign n10840 = ~n10838 & ~n10839;
  assign n10841 = ~n10464 & n10840;
  assign n10842 = n10464 & ~n10840;
  assign n10843 = ~n10841 & ~n10842;
  assign n10844 = n2288 & n4271;
  assign n10845 = pi85  & n4503;
  assign n10846 = pi87  & n4269;
  assign n10847 = pi86  & n4264;
  assign n10848 = ~n10846 & ~n10847;
  assign n10849 = ~n10845 & n10848;
  assign n10850 = ~n10844 & n10849;
  assign n10851 = pi35  & ~n10850;
  assign n10852 = pi35  & ~n10851;
  assign n10853 = ~n10850 & ~n10851;
  assign n10854 = ~n10852 & ~n10853;
  assign n10855 = ~n10843 & ~n10854;
  assign n10856 = n10843 & n10854;
  assign n10857 = ~n10855 & ~n10856;
  assign n10858 = n10714 & ~n10857;
  assign n10859 = ~n10714 & n10857;
  assign n10860 = ~n10858 & ~n10859;
  assign n10861 = n2801 & n3622;
  assign n10862 = pi88  & n3814;
  assign n10863 = pi90  & n3620;
  assign n10864 = pi89  & n3615;
  assign n10865 = ~n10863 & ~n10864;
  assign n10866 = ~n10862 & n10865;
  assign n10867 = ~n10861 & n10866;
  assign n10868 = pi32  & ~n10867;
  assign n10869 = pi32  & ~n10868;
  assign n10870 = ~n10867 & ~n10868;
  assign n10871 = ~n10869 & ~n10870;
  assign n10872 = n10860 & ~n10871;
  assign n10873 = ~n10860 & n10871;
  assign n10874 = ~n10872 & ~n10873;
  assign n10875 = ~n10713 & n10874;
  assign n10876 = ~n10713 & ~n10875;
  assign n10877 = ~n10872 & ~n10875;
  assign n10878 = ~n10873 & n10877;
  assign n10879 = ~n10876 & ~n10878;
  assign n10880 = n3034 & n3371;
  assign n10881 = pi91  & n3225;
  assign n10882 = pi93  & n3032;
  assign n10883 = pi92  & n3027;
  assign n10884 = ~n10882 & ~n10883;
  assign n10885 = ~n10881 & n10884;
  assign n10886 = ~n10880 & n10885;
  assign n10887 = pi29  & ~n10886;
  assign n10888 = pi29  & ~n10887;
  assign n10889 = ~n10886 & ~n10887;
  assign n10890 = ~n10888 & ~n10889;
  assign n10891 = n10879 & n10890;
  assign n10892 = ~n10879 & ~n10890;
  assign n10893 = ~n10891 & ~n10892;
  assign n10894 = ~n10712 & n10893;
  assign n10895 = n10712 & ~n10893;
  assign n10896 = ~n10894 & ~n10895;
  assign n10897 = n10711 & ~n10896;
  assign n10898 = ~n10711 & n10896;
  assign n10899 = ~n10897 & ~n10898;
  assign n10900 = ~n10700 & n10899;
  assign n10901 = n10700 & ~n10899;
  assign n10902 = ~n10900 & ~n10901;
  assign n10903 = n2043 & n4684;
  assign n10904 = pi97  & n2180;
  assign n10905 = pi99  & n2041;
  assign n10906 = pi98  & n2036;
  assign n10907 = ~n10905 & ~n10906;
  assign n10908 = ~n10904 & n10907;
  assign n10909 = ~n10903 & n10908;
  assign n10910 = pi23  & ~n10909;
  assign n10911 = pi23  & ~n10910;
  assign n10912 = ~n10909 & ~n10910;
  assign n10913 = ~n10911 & ~n10912;
  assign n10914 = n10902 & ~n10913;
  assign n10915 = n10902 & ~n10914;
  assign n10916 = ~n10913 & ~n10914;
  assign n10917 = ~n10915 & ~n10916;
  assign n10918 = ~n10554 & ~n10561;
  assign n10919 = n10917 & n10918;
  assign n10920 = ~n10917 & ~n10918;
  assign n10921 = ~n10919 & ~n10920;
  assign n10922 = n1611 & n5413;
  assign n10923 = pi100  & n1745;
  assign n10924 = pi102  & n1609;
  assign n10925 = pi101  & n1604;
  assign n10926 = ~n10924 & ~n10925;
  assign n10927 = ~n10923 & n10926;
  assign n10928 = ~n10922 & n10927;
  assign n10929 = pi20  & ~n10928;
  assign n10930 = pi20  & ~n10929;
  assign n10931 = ~n10928 & ~n10929;
  assign n10932 = ~n10930 & ~n10931;
  assign n10933 = n10921 & ~n10932;
  assign n10934 = n10921 & ~n10933;
  assign n10935 = ~n10932 & ~n10933;
  assign n10936 = ~n10934 & ~n10935;
  assign n10937 = ~n10574 & ~n10580;
  assign n10938 = n10936 & n10937;
  assign n10939 = ~n10936 & ~n10937;
  assign n10940 = ~n10938 & ~n10939;
  assign n10941 = n1297 & n6207;
  assign n10942 = pi103  & n1366;
  assign n10943 = pi105  & n1295;
  assign n10944 = pi104  & n1290;
  assign n10945 = ~n10943 & ~n10944;
  assign n10946 = ~n10942 & n10945;
  assign n10947 = ~n10941 & n10946;
  assign n10948 = pi17  & ~n10947;
  assign n10949 = pi17  & ~n10948;
  assign n10950 = ~n10947 & ~n10948;
  assign n10951 = ~n10949 & ~n10950;
  assign n10952 = n10940 & ~n10951;
  assign n10953 = n10940 & ~n10952;
  assign n10954 = ~n10951 & ~n10952;
  assign n10955 = ~n10953 & ~n10954;
  assign n10956 = ~n10593 & ~n10599;
  assign n10957 = n10955 & n10956;
  assign n10958 = ~n10955 & ~n10956;
  assign n10959 = ~n10957 & ~n10958;
  assign n10960 = n938 & n7060;
  assign n10961 = pi106  & n1052;
  assign n10962 = pi108  & n936;
  assign n10963 = pi107  & n931;
  assign n10964 = ~n10962 & ~n10963;
  assign n10965 = ~n10961 & n10964;
  assign n10966 = ~n10960 & n10965;
  assign n10967 = pi14  & ~n10966;
  assign n10968 = pi14  & ~n10967;
  assign n10969 = ~n10966 & ~n10967;
  assign n10970 = ~n10968 & ~n10969;
  assign n10971 = n10959 & ~n10970;
  assign n10972 = ~n10959 & n10970;
  assign n10973 = ~n10971 & ~n10972;
  assign n10974 = ~n10617 & n10973;
  assign n10975 = ~n10617 & ~n10974;
  assign n10976 = ~n10971 & ~n10974;
  assign n10977 = ~n10972 & n10976;
  assign n10978 = ~n10975 & ~n10977;
  assign n10979 = n687 & n7970;
  assign n10980 = pi109  & n763;
  assign n10981 = pi111  & n685;
  assign n10982 = pi110  & n680;
  assign n10983 = ~n10981 & ~n10982;
  assign n10984 = ~n10980 & n10983;
  assign n10985 = ~n10979 & n10984;
  assign n10986 = pi11  & ~n10985;
  assign n10987 = pi11  & ~n10986;
  assign n10988 = ~n10985 & ~n10986;
  assign n10989 = ~n10987 & ~n10988;
  assign n10990 = ~n10978 & ~n10989;
  assign n10991 = ~n10978 & ~n10990;
  assign n10992 = ~n10989 & ~n10990;
  assign n10993 = ~n10991 & ~n10992;
  assign n10994 = ~n10699 & ~n10993;
  assign n10995 = n10699 & n10993;
  assign n10996 = ~n10994 & ~n10995;
  assign n10997 = ~n10698 & n10996;
  assign n10998 = ~n10698 & ~n10997;
  assign n10999 = n10996 & ~n10997;
  assign n11000 = ~n10998 & ~n10999;
  assign n11001 = ~n10687 & ~n11000;
  assign n11002 = ~n10687 & ~n11001;
  assign n11003 = ~n11000 & ~n11001;
  assign n11004 = ~n11002 & ~n11003;
  assign n11005 = n342 & n9958;
  assign n11006 = pi115  & n380;
  assign n11007 = pi117  & n340;
  assign n11008 = pi116  & n335;
  assign n11009 = ~n11007 & ~n11008;
  assign n11010 = ~n11006 & n11009;
  assign n11011 = ~n11005 & n11010;
  assign n11012 = pi5  & ~n11011;
  assign n11013 = pi5  & ~n11012;
  assign n11014 = ~n11011 & ~n11012;
  assign n11015 = ~n11013 & ~n11014;
  assign n11016 = n11004 & n11015;
  assign n11017 = ~n11004 & ~n11015;
  assign n11018 = ~n11016 & ~n11017;
  assign n11019 = ~n10686 & n11018;
  assign n11020 = n10686 & ~n11018;
  assign n11021 = ~n11019 & ~n11020;
  assign n11022 = ~n10663 & ~n10665;
  assign n11023 = ~pi119  & ~pi120 ;
  assign n11024 = pi119  & pi120 ;
  assign n11025 = ~n11023 & ~n11024;
  assign n11026 = ~n11022 & n11025;
  assign n11027 = n11022 & ~n11025;
  assign n11028 = ~n11026 & ~n11027;
  assign n11029 = n262 & n11028;
  assign n11030 = pi118  & n288;
  assign n11031 = pi120  & n267;
  assign n11032 = pi119  & n269;
  assign n11033 = ~n11031 & ~n11032;
  assign n11034 = ~n11030 & n11033;
  assign n11035 = ~n11029 & n11034;
  assign n11036 = pi2  & ~n11035;
  assign n11037 = pi2  & ~n11036;
  assign n11038 = ~n11035 & ~n11036;
  assign n11039 = ~n11037 & ~n11038;
  assign n11040 = n11021 & ~n11039;
  assign n11041 = n11021 & ~n11040;
  assign n11042 = ~n11039 & ~n11040;
  assign n11043 = ~n11041 & ~n11042;
  assign n11044 = ~n10679 & ~n10682;
  assign n11045 = ~n11043 & ~n11044;
  assign n11046 = n11043 & n11044;
  assign po56  = ~n11045 & ~n11046;
  assign n11048 = ~n11017 & ~n11019;
  assign n11049 = n342 & n9984;
  assign n11050 = pi116  & n380;
  assign n11051 = pi118  & n340;
  assign n11052 = pi117  & n335;
  assign n11053 = ~n11051 & ~n11052;
  assign n11054 = ~n11050 & n11053;
  assign n11055 = ~n11049 & n11054;
  assign n11056 = pi5  & ~n11055;
  assign n11057 = pi5  & ~n11056;
  assign n11058 = ~n11055 & ~n11056;
  assign n11059 = ~n11057 & ~n11058;
  assign n11060 = ~n10997 & ~n11001;
  assign n11061 = n498 & n8963;
  assign n11062 = pi113  & n537;
  assign n11063 = pi115  & n496;
  assign n11064 = pi114  & n491;
  assign n11065 = ~n11063 & ~n11064;
  assign n11066 = ~n11062 & n11065;
  assign n11067 = ~n11061 & n11066;
  assign n11068 = pi8  & ~n11067;
  assign n11069 = pi8  & ~n11068;
  assign n11070 = ~n11067 & ~n11068;
  assign n11071 = ~n11069 & ~n11070;
  assign n11072 = ~n10990 & ~n10994;
  assign n11073 = n687 & n7997;
  assign n11074 = pi110  & n763;
  assign n11075 = pi112  & n685;
  assign n11076 = pi111  & n680;
  assign n11077 = ~n11075 & ~n11076;
  assign n11078 = ~n11074 & n11077;
  assign n11079 = ~n11073 & n11078;
  assign n11080 = pi11  & ~n11079;
  assign n11081 = pi11  & ~n11080;
  assign n11082 = ~n11079 & ~n11080;
  assign n11083 = ~n11081 & ~n11082;
  assign n11084 = n938 & n7349;
  assign n11085 = pi107  & n1052;
  assign n11086 = pi109  & n936;
  assign n11087 = pi108  & n931;
  assign n11088 = ~n11086 & ~n11087;
  assign n11089 = ~n11085 & n11088;
  assign n11090 = ~n11084 & n11089;
  assign n11091 = pi14  & ~n11090;
  assign n11092 = pi14  & ~n11091;
  assign n11093 = ~n11090 & ~n11091;
  assign n11094 = ~n11092 & ~n11093;
  assign n11095 = ~n10952 & ~n10958;
  assign n11096 = ~n10914 & ~n10920;
  assign n11097 = ~n10898 & ~n10900;
  assign n11098 = ~n10892 & ~n10894;
  assign n11099 = n3034 & n3565;
  assign n11100 = pi92  & n3225;
  assign n11101 = pi94  & n3032;
  assign n11102 = pi93  & n3027;
  assign n11103 = ~n11101 & ~n11102;
  assign n11104 = ~n11100 & n11103;
  assign n11105 = ~n11099 & n11104;
  assign n11106 = pi29  & ~n11105;
  assign n11107 = pi29  & ~n11106;
  assign n11108 = ~n11105 & ~n11106;
  assign n11109 = ~n11107 & ~n11108;
  assign n11110 = ~n10464 & ~n10840;
  assign n11111 = ~n10837 & ~n11110;
  assign n11112 = n1972 & n5008;
  assign n11113 = pi83  & n5241;
  assign n11114 = pi85  & n5006;
  assign n11115 = pi84  & n5001;
  assign n11116 = ~n11114 & ~n11115;
  assign n11117 = ~n11113 & n11116;
  assign n11118 = ~n11112 & n11117;
  assign n11119 = pi38  & ~n11118;
  assign n11120 = pi38  & ~n11119;
  assign n11121 = ~n11118 & ~n11119;
  assign n11122 = ~n11120 & ~n11121;
  assign n11123 = ~n10818 & ~n10822;
  assign n11124 = n1554 & n5739;
  assign n11125 = pi80  & n6030;
  assign n11126 = pi82  & n5737;
  assign n11127 = pi81  & n5732;
  assign n11128 = ~n11126 & ~n11127;
  assign n11129 = ~n11125 & n11128;
  assign n11130 = ~n11124 & n11129;
  assign n11131 = pi41  & ~n11130;
  assign n11132 = pi41  & ~n11131;
  assign n11133 = ~n11130 & ~n11131;
  assign n11134 = ~n11132 & ~n11133;
  assign n11135 = ~n10811 & ~n10815;
  assign n11136 = n1122 & n6539;
  assign n11137 = pi77  & n6873;
  assign n11138 = pi79  & n6537;
  assign n11139 = pi78  & n6532;
  assign n11140 = ~n11138 & ~n11139;
  assign n11141 = ~n11137 & n11140;
  assign n11142 = ~n11136 & n11141;
  assign n11143 = pi44  & ~n11142;
  assign n11144 = pi44  & ~n11143;
  assign n11145 = ~n11142 & ~n11143;
  assign n11146 = ~n11144 & ~n11145;
  assign n11147 = ~n10795 & ~n10797;
  assign n11148 = n891 & n7408;
  assign n11149 = pi74  & n7740;
  assign n11150 = pi76  & n7406;
  assign n11151 = pi75  & n7401;
  assign n11152 = ~n11150 & ~n11151;
  assign n11153 = ~n11149 & n11152;
  assign n11154 = ~n11148 & n11153;
  assign n11155 = pi47  & ~n11154;
  assign n11156 = pi47  & ~n11155;
  assign n11157 = ~n11154 & ~n11155;
  assign n11158 = ~n11156 & ~n11157;
  assign n11159 = ~n10789 & ~n10791;
  assign n11160 = pi56  & ~pi57 ;
  assign n11161 = ~pi56  & pi57 ;
  assign n11162 = ~n11160 & ~n11161;
  assign n11163 = pi64  & ~n11162;
  assign n11164 = ~n10756 & n11163;
  assign n11165 = n10756 & ~n11163;
  assign n11166 = ~n11164 & ~n11165;
  assign n11167 = n309 & n10394;
  assign n11168 = pi65  & n10744;
  assign n11169 = pi67  & n10392;
  assign n11170 = pi66  & n10387;
  assign n11171 = ~n11169 & ~n11170;
  assign n11172 = ~n11168 & n11171;
  assign n11173 = ~n11167 & n11172;
  assign n11174 = pi56  & ~n11173;
  assign n11175 = pi56  & ~n11174;
  assign n11176 = ~n11173 & ~n11174;
  assign n11177 = ~n11175 & ~n11176;
  assign n11178 = ~n11166 & ~n11177;
  assign n11179 = n11166 & n11177;
  assign n11180 = ~n11178 & ~n11179;
  assign n11181 = n450 & n9310;
  assign n11182 = pi68  & n9701;
  assign n11183 = pi70  & n9308;
  assign n11184 = pi69  & n9303;
  assign n11185 = ~n11183 & ~n11184;
  assign n11186 = ~n11182 & n11185;
  assign n11187 = ~n11181 & n11186;
  assign n11188 = pi53  & ~n11187;
  assign n11189 = pi53  & ~n11188;
  assign n11190 = ~n11187 & ~n11188;
  assign n11191 = ~n11189 & ~n11190;
  assign n11192 = n11180 & ~n11191;
  assign n11193 = n11180 & ~n11192;
  assign n11194 = ~n11191 & ~n11192;
  assign n11195 = ~n11193 & ~n11194;
  assign n11196 = ~n10774 & n11195;
  assign n11197 = n10774 & ~n11195;
  assign n11198 = ~n11196 & ~n11197;
  assign n11199 = n642 & n8334;
  assign n11200 = pi71  & n8685;
  assign n11201 = pi73  & n8332;
  assign n11202 = pi72  & n8327;
  assign n11203 = ~n11201 & ~n11202;
  assign n11204 = ~n11200 & n11203;
  assign n11205 = ~n11199 & n11204;
  assign n11206 = pi50  & ~n11205;
  assign n11207 = pi50  & ~n11206;
  assign n11208 = ~n11205 & ~n11206;
  assign n11209 = ~n11207 & ~n11208;
  assign n11210 = ~n11198 & ~n11209;
  assign n11211 = n11198 & n11209;
  assign n11212 = ~n11210 & ~n11211;
  assign n11213 = ~n11159 & n11212;
  assign n11214 = n11159 & ~n11212;
  assign n11215 = ~n11213 & ~n11214;
  assign n11216 = n11158 & ~n11215;
  assign n11217 = ~n11158 & n11215;
  assign n11218 = ~n11216 & ~n11217;
  assign n11219 = ~n11147 & n11218;
  assign n11220 = n11147 & ~n11218;
  assign n11221 = ~n11219 & ~n11220;
  assign n11222 = ~n11146 & n11221;
  assign n11223 = n11146 & ~n11221;
  assign n11224 = ~n11222 & ~n11223;
  assign n11225 = ~n11135 & n11224;
  assign n11226 = n11135 & ~n11224;
  assign n11227 = ~n11225 & ~n11226;
  assign n11228 = ~n11134 & n11227;
  assign n11229 = ~n11134 & ~n11228;
  assign n11230 = n11227 & ~n11228;
  assign n11231 = ~n11229 & ~n11230;
  assign n11232 = ~n11123 & ~n11231;
  assign n11233 = n11123 & n11231;
  assign n11234 = ~n11232 & ~n11233;
  assign n11235 = ~n11122 & n11234;
  assign n11236 = n11122 & ~n11234;
  assign n11237 = ~n11235 & ~n11236;
  assign n11238 = ~n11111 & n11237;
  assign n11239 = n11111 & ~n11237;
  assign n11240 = ~n11238 & ~n11239;
  assign n11241 = n2446 & n4271;
  assign n11242 = pi86  & n4503;
  assign n11243 = pi88  & n4269;
  assign n11244 = pi87  & n4264;
  assign n11245 = ~n11243 & ~n11244;
  assign n11246 = ~n11242 & n11245;
  assign n11247 = ~n11241 & n11246;
  assign n11248 = pi35  & ~n11247;
  assign n11249 = pi35  & ~n11248;
  assign n11250 = ~n11247 & ~n11248;
  assign n11251 = ~n11249 & ~n11250;
  assign n11252 = n11240 & ~n11251;
  assign n11253 = n11240 & ~n11252;
  assign n11254 = ~n11251 & ~n11252;
  assign n11255 = ~n11253 & ~n11254;
  assign n11256 = ~n10855 & ~n10859;
  assign n11257 = n11255 & n11256;
  assign n11258 = ~n11255 & ~n11256;
  assign n11259 = ~n11257 & ~n11258;
  assign n11260 = n2978 & n3622;
  assign n11261 = pi89  & n3814;
  assign n11262 = pi91  & n3620;
  assign n11263 = pi90  & n3615;
  assign n11264 = ~n11262 & ~n11263;
  assign n11265 = ~n11261 & n11264;
  assign n11266 = ~n11260 & n11265;
  assign n11267 = pi32  & ~n11266;
  assign n11268 = pi32  & ~n11267;
  assign n11269 = ~n11266 & ~n11267;
  assign n11270 = ~n11268 & ~n11269;
  assign n11271 = ~n11259 & n11270;
  assign n11272 = n11259 & ~n11270;
  assign n11273 = ~n11271 & ~n11272;
  assign n11274 = ~n10877 & n11273;
  assign n11275 = n10877 & ~n11273;
  assign n11276 = ~n11274 & ~n11275;
  assign n11277 = ~n11109 & n11276;
  assign n11278 = n11109 & ~n11276;
  assign n11279 = ~n11277 & ~n11278;
  assign n11280 = ~n11098 & n11279;
  assign n11281 = n11098 & ~n11279;
  assign n11282 = ~n11280 & ~n11281;
  assign n11283 = n2523 & n4211;
  assign n11284 = pi95  & n2667;
  assign n11285 = pi97  & n2521;
  assign n11286 = pi96  & n2516;
  assign n11287 = ~n11285 & ~n11286;
  assign n11288 = ~n11284 & n11287;
  assign n11289 = ~n11283 & n11288;
  assign n11290 = pi26  & ~n11289;
  assign n11291 = pi26  & ~n11290;
  assign n11292 = ~n11289 & ~n11290;
  assign n11293 = ~n11291 & ~n11292;
  assign n11294 = n11282 & ~n11293;
  assign n11295 = n11282 & ~n11294;
  assign n11296 = ~n11293 & ~n11294;
  assign n11297 = ~n11295 & ~n11296;
  assign n11298 = ~n11097 & n11297;
  assign n11299 = n11097 & ~n11297;
  assign n11300 = ~n11298 & ~n11299;
  assign n11301 = n2043 & n4910;
  assign n11302 = pi98  & n2180;
  assign n11303 = pi100  & n2041;
  assign n11304 = pi99  & n2036;
  assign n11305 = ~n11303 & ~n11304;
  assign n11306 = ~n11302 & n11305;
  assign n11307 = ~n11301 & n11306;
  assign n11308 = pi23  & ~n11307;
  assign n11309 = pi23  & ~n11308;
  assign n11310 = ~n11307 & ~n11308;
  assign n11311 = ~n11309 & ~n11310;
  assign n11312 = ~n11300 & ~n11311;
  assign n11313 = n11300 & n11311;
  assign n11314 = ~n11312 & ~n11313;
  assign n11315 = n11096 & ~n11314;
  assign n11316 = ~n11096 & n11314;
  assign n11317 = ~n11315 & ~n11316;
  assign n11318 = n1611 & n5664;
  assign n11319 = pi101  & n1745;
  assign n11320 = pi103  & n1609;
  assign n11321 = pi102  & n1604;
  assign n11322 = ~n11320 & ~n11321;
  assign n11323 = ~n11319 & n11322;
  assign n11324 = ~n11318 & n11323;
  assign n11325 = pi20  & ~n11324;
  assign n11326 = pi20  & ~n11325;
  assign n11327 = ~n11324 & ~n11325;
  assign n11328 = ~n11326 & ~n11327;
  assign n11329 = n11317 & ~n11328;
  assign n11330 = n11317 & ~n11329;
  assign n11331 = ~n11328 & ~n11329;
  assign n11332 = ~n11330 & ~n11331;
  assign n11333 = ~n10933 & ~n10939;
  assign n11334 = n11332 & n11333;
  assign n11335 = ~n11332 & ~n11333;
  assign n11336 = ~n11334 & ~n11335;
  assign n11337 = n1297 & n6477;
  assign n11338 = pi104  & n1366;
  assign n11339 = pi106  & n1295;
  assign n11340 = pi105  & n1290;
  assign n11341 = ~n11339 & ~n11340;
  assign n11342 = ~n11338 & n11341;
  assign n11343 = ~n11337 & n11342;
  assign n11344 = pi17  & ~n11343;
  assign n11345 = pi17  & ~n11344;
  assign n11346 = ~n11343 & ~n11344;
  assign n11347 = ~n11345 & ~n11346;
  assign n11348 = ~n11336 & n11347;
  assign n11349 = n11336 & ~n11347;
  assign n11350 = ~n11348 & ~n11349;
  assign n11351 = ~n11095 & n11350;
  assign n11352 = n11095 & ~n11350;
  assign n11353 = ~n11351 & ~n11352;
  assign n11354 = ~n11094 & n11353;
  assign n11355 = ~n11094 & ~n11354;
  assign n11356 = n11353 & ~n11354;
  assign n11357 = ~n11355 & ~n11356;
  assign n11358 = ~n10976 & ~n11357;
  assign n11359 = n10976 & n11357;
  assign n11360 = ~n11358 & ~n11359;
  assign n11361 = ~n11083 & n11360;
  assign n11362 = ~n11083 & ~n11361;
  assign n11363 = n11360 & ~n11361;
  assign n11364 = ~n11362 & ~n11363;
  assign n11365 = ~n11072 & ~n11364;
  assign n11366 = n11072 & n11364;
  assign n11367 = ~n11365 & ~n11366;
  assign n11368 = ~n11071 & n11367;
  assign n11369 = ~n11071 & ~n11368;
  assign n11370 = n11367 & ~n11368;
  assign n11371 = ~n11369 & ~n11370;
  assign n11372 = ~n11060 & ~n11371;
  assign n11373 = n11060 & n11371;
  assign n11374 = ~n11372 & ~n11373;
  assign n11375 = ~n11059 & n11374;
  assign n11376 = ~n11059 & ~n11375;
  assign n11377 = n11374 & ~n11375;
  assign n11378 = ~n11376 & ~n11377;
  assign n11379 = ~n11048 & ~n11378;
  assign n11380 = ~n11048 & ~n11379;
  assign n11381 = ~n11378 & ~n11379;
  assign n11382 = ~n11380 & ~n11381;
  assign n11383 = ~n11024 & ~n11026;
  assign n11384 = ~pi120  & ~pi121 ;
  assign n11385 = pi120  & pi121 ;
  assign n11386 = ~n11384 & ~n11385;
  assign n11387 = ~n11383 & n11386;
  assign n11388 = n11383 & ~n11386;
  assign n11389 = ~n11387 & ~n11388;
  assign n11390 = n262 & n11389;
  assign n11391 = pi119  & n288;
  assign n11392 = pi121  & n267;
  assign n11393 = pi120  & n269;
  assign n11394 = ~n11392 & ~n11393;
  assign n11395 = ~n11391 & n11394;
  assign n11396 = ~n11390 & n11395;
  assign n11397 = pi2  & ~n11396;
  assign n11398 = pi2  & ~n11397;
  assign n11399 = ~n11396 & ~n11397;
  assign n11400 = ~n11398 & ~n11399;
  assign n11401 = ~n11382 & ~n11400;
  assign n11402 = ~n11382 & ~n11401;
  assign n11403 = ~n11400 & ~n11401;
  assign n11404 = ~n11402 & ~n11403;
  assign n11405 = ~n11040 & ~n11045;
  assign n11406 = ~n11404 & ~n11405;
  assign n11407 = n11404 & n11405;
  assign po57  = ~n11406 & ~n11407;
  assign n11409 = ~n11375 & ~n11379;
  assign n11410 = n342 & n10667;
  assign n11411 = pi117  & n380;
  assign n11412 = pi119  & n340;
  assign n11413 = pi118  & n335;
  assign n11414 = ~n11412 & ~n11413;
  assign n11415 = ~n11411 & n11414;
  assign n11416 = ~n11410 & n11415;
  assign n11417 = pi5  & ~n11416;
  assign n11418 = pi5  & ~n11417;
  assign n11419 = ~n11416 & ~n11417;
  assign n11420 = ~n11418 & ~n11419;
  assign n11421 = ~n11368 & ~n11372;
  assign n11422 = n498 & n9614;
  assign n11423 = pi114  & n537;
  assign n11424 = pi116  & n496;
  assign n11425 = pi115  & n491;
  assign n11426 = ~n11424 & ~n11425;
  assign n11427 = ~n11423 & n11426;
  assign n11428 = ~n11422 & n11427;
  assign n11429 = pi8  & ~n11428;
  assign n11430 = pi8  & ~n11429;
  assign n11431 = ~n11428 & ~n11429;
  assign n11432 = ~n11430 & ~n11431;
  assign n11433 = ~n11361 & ~n11365;
  assign n11434 = n687 & n8612;
  assign n11435 = pi111  & n763;
  assign n11436 = pi113  & n685;
  assign n11437 = pi112  & n680;
  assign n11438 = ~n11436 & ~n11437;
  assign n11439 = ~n11435 & n11438;
  assign n11440 = ~n11434 & n11439;
  assign n11441 = pi11  & ~n11440;
  assign n11442 = pi11  & ~n11441;
  assign n11443 = ~n11440 & ~n11441;
  assign n11444 = ~n11442 & ~n11443;
  assign n11445 = ~n11354 & ~n11358;
  assign n11446 = ~n11349 & ~n11351;
  assign n11447 = ~n11277 & ~n11280;
  assign n11448 = ~n11272 & ~n11274;
  assign n11449 = ~n11228 & ~n11232;
  assign n11450 = ~n11217 & ~n11219;
  assign n11451 = ~n10774 & ~n11195;
  assign n11452 = ~n11192 & ~n11451;
  assign n11453 = n475 & n9310;
  assign n11454 = pi69  & n9701;
  assign n11455 = pi71  & n9308;
  assign n11456 = pi70  & n9303;
  assign n11457 = ~n11455 & ~n11456;
  assign n11458 = ~n11454 & n11457;
  assign n11459 = ~n11453 & n11458;
  assign n11460 = pi53  & ~n11459;
  assign n11461 = pi53  & ~n11460;
  assign n11462 = ~n11459 & ~n11460;
  assign n11463 = ~n11461 & ~n11462;
  assign n11464 = n10756 & n11163;
  assign n11465 = ~n11178 & ~n11464;
  assign n11466 = n359 & n10394;
  assign n11467 = pi66  & n10744;
  assign n11468 = pi68  & n10392;
  assign n11469 = pi67  & n10387;
  assign n11470 = ~n11468 & ~n11469;
  assign n11471 = ~n11467 & n11470;
  assign n11472 = ~n11466 & n11471;
  assign n11473 = pi56  & ~n11472;
  assign n11474 = pi56  & ~n11473;
  assign n11475 = ~n11472 & ~n11473;
  assign n11476 = ~n11474 & ~n11475;
  assign n11477 = pi59  & ~n11163;
  assign n11478 = ~pi57  & pi58 ;
  assign n11479 = pi57  & ~pi58 ;
  assign n11480 = ~n11478 & ~n11479;
  assign n11481 = n11162 & ~n11480;
  assign n11482 = pi64  & n11481;
  assign n11483 = ~pi58  & pi59 ;
  assign n11484 = pi58  & ~pi59 ;
  assign n11485 = ~n11483 & ~n11484;
  assign n11486 = ~n11162 & n11485;
  assign n11487 = pi65  & n11486;
  assign n11488 = ~n11162 & ~n11485;
  assign n11489 = ~n265 & n11488;
  assign n11490 = ~n11482 & ~n11487;
  assign n11491 = ~n11489 & n11490;
  assign n11492 = pi59  & ~n11491;
  assign n11493 = pi59  & ~n11492;
  assign n11494 = ~n11491 & ~n11492;
  assign n11495 = ~n11493 & ~n11494;
  assign n11496 = n11477 & ~n11495;
  assign n11497 = ~n11477 & n11495;
  assign n11498 = ~n11496 & ~n11497;
  assign n11499 = n11476 & ~n11498;
  assign n11500 = ~n11476 & n11498;
  assign n11501 = ~n11499 & ~n11500;
  assign n11502 = ~n11465 & n11501;
  assign n11503 = n11465 & ~n11501;
  assign n11504 = ~n11502 & ~n11503;
  assign n11505 = n11463 & ~n11504;
  assign n11506 = ~n11463 & n11504;
  assign n11507 = ~n11505 & ~n11506;
  assign n11508 = ~n11452 & n11507;
  assign n11509 = n11452 & ~n11507;
  assign n11510 = ~n11508 & ~n11509;
  assign n11511 = n729 & n8334;
  assign n11512 = pi72  & n8685;
  assign n11513 = pi74  & n8332;
  assign n11514 = pi73  & n8327;
  assign n11515 = ~n11513 & ~n11514;
  assign n11516 = ~n11512 & n11515;
  assign n11517 = ~n11511 & n11516;
  assign n11518 = pi50  & ~n11517;
  assign n11519 = pi50  & ~n11518;
  assign n11520 = ~n11517 & ~n11518;
  assign n11521 = ~n11519 & ~n11520;
  assign n11522 = n11510 & ~n11521;
  assign n11523 = n11510 & ~n11522;
  assign n11524 = ~n11521 & ~n11522;
  assign n11525 = ~n11523 & ~n11524;
  assign n11526 = ~n11210 & ~n11213;
  assign n11527 = n11525 & n11526;
  assign n11528 = ~n11525 & ~n11526;
  assign n11529 = ~n11527 & ~n11528;
  assign n11530 = n999 & n7408;
  assign n11531 = pi75  & n7740;
  assign n11532 = pi77  & n7406;
  assign n11533 = pi76  & n7401;
  assign n11534 = ~n11532 & ~n11533;
  assign n11535 = ~n11531 & n11534;
  assign n11536 = ~n11530 & n11535;
  assign n11537 = pi47  & ~n11536;
  assign n11538 = pi47  & ~n11537;
  assign n11539 = ~n11536 & ~n11537;
  assign n11540 = ~n11538 & ~n11539;
  assign n11541 = n11529 & ~n11540;
  assign n11542 = ~n11529 & n11540;
  assign n11543 = ~n11541 & ~n11542;
  assign n11544 = ~n11450 & n11543;
  assign n11545 = ~n11450 & ~n11544;
  assign n11546 = ~n11541 & ~n11544;
  assign n11547 = ~n11542 & n11546;
  assign n11548 = ~n11545 & ~n11547;
  assign n11549 = n1225 & n6539;
  assign n11550 = pi78  & n6873;
  assign n11551 = pi80  & n6537;
  assign n11552 = pi79  & n6532;
  assign n11553 = ~n11551 & ~n11552;
  assign n11554 = ~n11550 & n11553;
  assign n11555 = ~n11549 & n11554;
  assign n11556 = pi44  & ~n11555;
  assign n11557 = pi44  & ~n11556;
  assign n11558 = ~n11555 & ~n11556;
  assign n11559 = ~n11557 & ~n11558;
  assign n11560 = ~n11548 & ~n11559;
  assign n11561 = ~n11548 & ~n11560;
  assign n11562 = ~n11559 & ~n11560;
  assign n11563 = ~n11561 & ~n11562;
  assign n11564 = ~n11222 & ~n11225;
  assign n11565 = n11563 & n11564;
  assign n11566 = ~n11563 & ~n11564;
  assign n11567 = ~n11565 & ~n11566;
  assign n11568 = n1696 & n5739;
  assign n11569 = pi81  & n6030;
  assign n11570 = pi83  & n5737;
  assign n11571 = pi82  & n5732;
  assign n11572 = ~n11570 & ~n11571;
  assign n11573 = ~n11569 & n11572;
  assign n11574 = ~n11568 & n11573;
  assign n11575 = pi41  & ~n11574;
  assign n11576 = pi41  & ~n11575;
  assign n11577 = ~n11574 & ~n11575;
  assign n11578 = ~n11576 & ~n11577;
  assign n11579 = n11567 & ~n11578;
  assign n11580 = ~n11567 & n11578;
  assign n11581 = ~n11579 & ~n11580;
  assign n11582 = ~n11449 & n11581;
  assign n11583 = ~n11449 & ~n11582;
  assign n11584 = ~n11579 & ~n11582;
  assign n11585 = ~n11580 & n11584;
  assign n11586 = ~n11583 & ~n11585;
  assign n11587 = n2133 & n5008;
  assign n11588 = pi84  & n5241;
  assign n11589 = pi86  & n5006;
  assign n11590 = pi85  & n5001;
  assign n11591 = ~n11589 & ~n11590;
  assign n11592 = ~n11588 & n11591;
  assign n11593 = ~n11587 & n11592;
  assign n11594 = pi38  & ~n11593;
  assign n11595 = pi38  & ~n11594;
  assign n11596 = ~n11593 & ~n11594;
  assign n11597 = ~n11595 & ~n11596;
  assign n11598 = ~n11586 & ~n11597;
  assign n11599 = ~n11586 & ~n11598;
  assign n11600 = ~n11597 & ~n11598;
  assign n11601 = ~n11599 & ~n11600;
  assign n11602 = ~n11235 & ~n11238;
  assign n11603 = n11601 & n11602;
  assign n11604 = ~n11601 & ~n11602;
  assign n11605 = ~n11603 & ~n11604;
  assign n11606 = n2473 & n4271;
  assign n11607 = pi87  & n4503;
  assign n11608 = pi89  & n4269;
  assign n11609 = pi88  & n4264;
  assign n11610 = ~n11608 & ~n11609;
  assign n11611 = ~n11607 & n11610;
  assign n11612 = ~n11606 & n11611;
  assign n11613 = pi35  & ~n11612;
  assign n11614 = pi35  & ~n11613;
  assign n11615 = ~n11612 & ~n11613;
  assign n11616 = ~n11614 & ~n11615;
  assign n11617 = n11605 & ~n11616;
  assign n11618 = n11605 & ~n11617;
  assign n11619 = ~n11616 & ~n11617;
  assign n11620 = ~n11618 & ~n11619;
  assign n11621 = ~n11252 & ~n11258;
  assign n11622 = n11620 & n11621;
  assign n11623 = ~n11620 & ~n11621;
  assign n11624 = ~n11622 & ~n11623;
  assign n11625 = n3177 & n3622;
  assign n11626 = pi90  & n3814;
  assign n11627 = pi92  & n3620;
  assign n11628 = pi91  & n3615;
  assign n11629 = ~n11627 & ~n11628;
  assign n11630 = ~n11626 & n11629;
  assign n11631 = ~n11625 & n11630;
  assign n11632 = pi32  & ~n11631;
  assign n11633 = pi32  & ~n11632;
  assign n11634 = ~n11631 & ~n11632;
  assign n11635 = ~n11633 & ~n11634;
  assign n11636 = n11624 & ~n11635;
  assign n11637 = n11624 & ~n11636;
  assign n11638 = ~n11635 & ~n11636;
  assign n11639 = ~n11637 & ~n11638;
  assign n11640 = ~n11448 & n11639;
  assign n11641 = n11448 & ~n11639;
  assign n11642 = ~n11640 & ~n11641;
  assign n11643 = n3034 & n3784;
  assign n11644 = pi93  & n3225;
  assign n11645 = pi95  & n3032;
  assign n11646 = pi94  & n3027;
  assign n11647 = ~n11645 & ~n11646;
  assign n11648 = ~n11644 & n11647;
  assign n11649 = ~n11643 & n11648;
  assign n11650 = pi29  & ~n11649;
  assign n11651 = pi29  & ~n11650;
  assign n11652 = ~n11649 & ~n11650;
  assign n11653 = ~n11651 & ~n11652;
  assign n11654 = ~n11642 & ~n11653;
  assign n11655 = n11642 & n11653;
  assign n11656 = ~n11654 & ~n11655;
  assign n11657 = n11447 & ~n11656;
  assign n11658 = ~n11447 & n11656;
  assign n11659 = ~n11657 & ~n11658;
  assign n11660 = n2523 & n4454;
  assign n11661 = pi96  & n2667;
  assign n11662 = pi98  & n2521;
  assign n11663 = pi97  & n2516;
  assign n11664 = ~n11662 & ~n11663;
  assign n11665 = ~n11661 & n11664;
  assign n11666 = ~n11660 & n11665;
  assign n11667 = pi26  & ~n11666;
  assign n11668 = pi26  & ~n11667;
  assign n11669 = ~n11666 & ~n11667;
  assign n11670 = ~n11668 & ~n11669;
  assign n11671 = n11659 & ~n11670;
  assign n11672 = n11659 & ~n11671;
  assign n11673 = ~n11670 & ~n11671;
  assign n11674 = ~n11672 & ~n11673;
  assign n11675 = ~n11097 & ~n11297;
  assign n11676 = ~n11294 & ~n11675;
  assign n11677 = n11674 & n11676;
  assign n11678 = ~n11674 & ~n11676;
  assign n11679 = ~n11677 & ~n11678;
  assign n11680 = n2043 & n5169;
  assign n11681 = pi99  & n2180;
  assign n11682 = pi101  & n2041;
  assign n11683 = pi100  & n2036;
  assign n11684 = ~n11682 & ~n11683;
  assign n11685 = ~n11681 & n11684;
  assign n11686 = ~n11680 & n11685;
  assign n11687 = pi23  & ~n11686;
  assign n11688 = pi23  & ~n11687;
  assign n11689 = ~n11686 & ~n11687;
  assign n11690 = ~n11688 & ~n11689;
  assign n11691 = n11679 & ~n11690;
  assign n11692 = n11679 & ~n11691;
  assign n11693 = ~n11690 & ~n11691;
  assign n11694 = ~n11692 & ~n11693;
  assign n11695 = ~n11312 & ~n11316;
  assign n11696 = n11694 & n11695;
  assign n11697 = ~n11694 & ~n11695;
  assign n11698 = ~n11696 & ~n11697;
  assign n11699 = n1611 & n5943;
  assign n11700 = pi102  & n1745;
  assign n11701 = pi104  & n1609;
  assign n11702 = pi103  & n1604;
  assign n11703 = ~n11701 & ~n11702;
  assign n11704 = ~n11700 & n11703;
  assign n11705 = ~n11699 & n11704;
  assign n11706 = pi20  & ~n11705;
  assign n11707 = pi20  & ~n11706;
  assign n11708 = ~n11705 & ~n11706;
  assign n11709 = ~n11707 & ~n11708;
  assign n11710 = n11698 & ~n11709;
  assign n11711 = n11698 & ~n11710;
  assign n11712 = ~n11709 & ~n11710;
  assign n11713 = ~n11711 & ~n11712;
  assign n11714 = ~n11329 & ~n11335;
  assign n11715 = n11713 & n11714;
  assign n11716 = ~n11713 & ~n11714;
  assign n11717 = ~n11715 & ~n11716;
  assign n11718 = n1297 & n6775;
  assign n11719 = pi105  & n1366;
  assign n11720 = pi107  & n1295;
  assign n11721 = pi106  & n1290;
  assign n11722 = ~n11720 & ~n11721;
  assign n11723 = ~n11719 & n11722;
  assign n11724 = ~n11718 & n11723;
  assign n11725 = pi17  & ~n11724;
  assign n11726 = pi17  & ~n11725;
  assign n11727 = ~n11724 & ~n11725;
  assign n11728 = ~n11726 & ~n11727;
  assign n11729 = n11717 & ~n11728;
  assign n11730 = ~n11717 & n11728;
  assign n11731 = ~n11729 & ~n11730;
  assign n11732 = ~n11446 & n11731;
  assign n11733 = ~n11446 & ~n11732;
  assign n11734 = ~n11729 & ~n11732;
  assign n11735 = ~n11730 & n11734;
  assign n11736 = ~n11733 & ~n11735;
  assign n11737 = n938 & n7665;
  assign n11738 = pi108  & n1052;
  assign n11739 = pi110  & n936;
  assign n11740 = pi109  & n931;
  assign n11741 = ~n11739 & ~n11740;
  assign n11742 = ~n11738 & n11741;
  assign n11743 = ~n11737 & n11742;
  assign n11744 = pi14  & ~n11743;
  assign n11745 = pi14  & ~n11744;
  assign n11746 = ~n11743 & ~n11744;
  assign n11747 = ~n11745 & ~n11746;
  assign n11748 = n11736 & n11747;
  assign n11749 = ~n11736 & ~n11747;
  assign n11750 = ~n11748 & ~n11749;
  assign n11751 = ~n11445 & n11750;
  assign n11752 = n11445 & ~n11750;
  assign n11753 = ~n11751 & ~n11752;
  assign n11754 = n11444 & ~n11753;
  assign n11755 = ~n11444 & n11753;
  assign n11756 = ~n11754 & ~n11755;
  assign n11757 = ~n11433 & n11756;
  assign n11758 = n11433 & ~n11756;
  assign n11759 = ~n11757 & ~n11758;
  assign n11760 = n11432 & ~n11759;
  assign n11761 = ~n11432 & n11759;
  assign n11762 = ~n11760 & ~n11761;
  assign n11763 = ~n11421 & n11762;
  assign n11764 = n11421 & ~n11762;
  assign n11765 = ~n11763 & ~n11764;
  assign n11766 = n11420 & ~n11765;
  assign n11767 = ~n11420 & n11765;
  assign n11768 = ~n11766 & ~n11767;
  assign n11769 = ~n11409 & n11768;
  assign n11770 = n11409 & ~n11768;
  assign n11771 = ~n11769 & ~n11770;
  assign n11772 = ~n11385 & ~n11387;
  assign n11773 = ~pi121  & ~pi122 ;
  assign n11774 = pi121  & pi122 ;
  assign n11775 = ~n11773 & ~n11774;
  assign n11776 = ~n11772 & n11775;
  assign n11777 = n11772 & ~n11775;
  assign n11778 = ~n11776 & ~n11777;
  assign n11779 = n262 & n11778;
  assign n11780 = pi120  & n288;
  assign n11781 = pi122  & n267;
  assign n11782 = pi121  & n269;
  assign n11783 = ~n11781 & ~n11782;
  assign n11784 = ~n11780 & n11783;
  assign n11785 = ~n11779 & n11784;
  assign n11786 = pi2  & ~n11785;
  assign n11787 = pi2  & ~n11786;
  assign n11788 = ~n11785 & ~n11786;
  assign n11789 = ~n11787 & ~n11788;
  assign n11790 = n11771 & ~n11789;
  assign n11791 = n11771 & ~n11790;
  assign n11792 = ~n11789 & ~n11790;
  assign n11793 = ~n11791 & ~n11792;
  assign n11794 = ~n11401 & ~n11406;
  assign n11795 = ~n11793 & ~n11794;
  assign n11796 = n11793 & n11794;
  assign po58  = ~n11795 & ~n11796;
  assign n11798 = ~n11790 & ~n11795;
  assign n11799 = ~n11767 & ~n11769;
  assign n11800 = ~n11761 & ~n11763;
  assign n11801 = n498 & n9958;
  assign n11802 = pi115  & n537;
  assign n11803 = pi117  & n496;
  assign n11804 = pi116  & n491;
  assign n11805 = ~n11803 & ~n11804;
  assign n11806 = ~n11802 & n11805;
  assign n11807 = ~n11801 & n11806;
  assign n11808 = pi8  & ~n11807;
  assign n11809 = pi8  & ~n11808;
  assign n11810 = ~n11807 & ~n11808;
  assign n11811 = ~n11809 & ~n11810;
  assign n11812 = ~n11755 & ~n11757;
  assign n11813 = ~n11749 & ~n11751;
  assign n11814 = ~n11710 & ~n11716;
  assign n11815 = ~n11654 & ~n11658;
  assign n11816 = ~n11448 & ~n11639;
  assign n11817 = ~n11636 & ~n11816;
  assign n11818 = ~n11598 & ~n11604;
  assign n11819 = ~n11560 & ~n11566;
  assign n11820 = n1434 & n6539;
  assign n11821 = pi79  & n6873;
  assign n11822 = pi81  & n6537;
  assign n11823 = pi80  & n6532;
  assign n11824 = ~n11822 & ~n11823;
  assign n11825 = ~n11821 & n11824;
  assign n11826 = ~n11820 & n11825;
  assign n11827 = pi44  & ~n11826;
  assign n11828 = pi44  & ~n11827;
  assign n11829 = ~n11826 & ~n11827;
  assign n11830 = ~n11828 & ~n11829;
  assign n11831 = ~n11522 & ~n11528;
  assign n11832 = n809 & n8334;
  assign n11833 = pi73  & n8685;
  assign n11834 = pi75  & n8332;
  assign n11835 = pi74  & n8327;
  assign n11836 = ~n11834 & ~n11835;
  assign n11837 = ~n11833 & n11836;
  assign n11838 = ~n11832 & n11837;
  assign n11839 = pi50  & ~n11838;
  assign n11840 = pi50  & ~n11839;
  assign n11841 = ~n11838 & ~n11839;
  assign n11842 = ~n11840 & ~n11841;
  assign n11843 = ~n11506 & ~n11508;
  assign n11844 = ~n11500 & ~n11502;
  assign n11845 = n286 & n11488;
  assign n11846 = n11162 & n11480;
  assign n11847 = ~n11485 & n11846;
  assign n11848 = pi64  & n11847;
  assign n11849 = pi66  & n11486;
  assign n11850 = pi65  & n11481;
  assign n11851 = ~n11849 & ~n11850;
  assign n11852 = ~n11845 & n11851;
  assign n11853 = ~n11848 & n11852;
  assign n11854 = pi59  & ~n11853;
  assign n11855 = pi59  & ~n11854;
  assign n11856 = ~n11853 & ~n11854;
  assign n11857 = ~n11855 & ~n11856;
  assign n11858 = ~n11496 & n11857;
  assign n11859 = n11496 & ~n11857;
  assign n11860 = ~n11858 & ~n11859;
  assign n11861 = n401 & n10394;
  assign n11862 = pi67  & n10744;
  assign n11863 = pi69  & n10392;
  assign n11864 = pi68  & n10387;
  assign n11865 = ~n11863 & ~n11864;
  assign n11866 = ~n11862 & n11865;
  assign n11867 = ~n11861 & n11866;
  assign n11868 = pi56  & ~n11867;
  assign n11869 = pi56  & ~n11868;
  assign n11870 = ~n11867 & ~n11868;
  assign n11871 = ~n11869 & ~n11870;
  assign n11872 = n11860 & ~n11871;
  assign n11873 = ~n11860 & n11871;
  assign n11874 = ~n11872 & ~n11873;
  assign n11875 = ~n11844 & n11874;
  assign n11876 = ~n11844 & ~n11875;
  assign n11877 = ~n11872 & ~n11875;
  assign n11878 = ~n11873 & n11877;
  assign n11879 = ~n11876 & ~n11878;
  assign n11880 = n576 & n9310;
  assign n11881 = pi70  & n9701;
  assign n11882 = pi72  & n9308;
  assign n11883 = pi71  & n9303;
  assign n11884 = ~n11882 & ~n11883;
  assign n11885 = ~n11881 & n11884;
  assign n11886 = ~n11880 & n11885;
  assign n11887 = pi53  & ~n11886;
  assign n11888 = pi53  & ~n11887;
  assign n11889 = ~n11886 & ~n11887;
  assign n11890 = ~n11888 & ~n11889;
  assign n11891 = n11879 & n11890;
  assign n11892 = ~n11879 & ~n11890;
  assign n11893 = ~n11891 & ~n11892;
  assign n11894 = ~n11843 & n11893;
  assign n11895 = n11843 & ~n11893;
  assign n11896 = ~n11894 & ~n11895;
  assign n11897 = n11842 & ~n11896;
  assign n11898 = ~n11842 & n11896;
  assign n11899 = ~n11897 & ~n11898;
  assign n11900 = ~n11831 & n11899;
  assign n11901 = n11831 & ~n11899;
  assign n11902 = ~n11900 & ~n11901;
  assign n11903 = n1025 & n7408;
  assign n11904 = pi76  & n7740;
  assign n11905 = pi78  & n7406;
  assign n11906 = pi77  & n7401;
  assign n11907 = ~n11905 & ~n11906;
  assign n11908 = ~n11904 & n11907;
  assign n11909 = ~n11903 & n11908;
  assign n11910 = pi47  & ~n11909;
  assign n11911 = pi47  & ~n11910;
  assign n11912 = ~n11909 & ~n11910;
  assign n11913 = ~n11911 & ~n11912;
  assign n11914 = n11902 & ~n11913;
  assign n11915 = n11902 & ~n11914;
  assign n11916 = ~n11913 & ~n11914;
  assign n11917 = ~n11915 & ~n11916;
  assign n11918 = ~n11546 & ~n11917;
  assign n11919 = n11546 & n11917;
  assign n11920 = ~n11918 & ~n11919;
  assign n11921 = ~n11830 & n11920;
  assign n11922 = ~n11830 & ~n11921;
  assign n11923 = n11920 & ~n11921;
  assign n11924 = ~n11922 & ~n11923;
  assign n11925 = ~n11819 & ~n11924;
  assign n11926 = ~n11819 & ~n11925;
  assign n11927 = ~n11924 & ~n11925;
  assign n11928 = ~n11926 & ~n11927;
  assign n11929 = n1834 & n5739;
  assign n11930 = pi82  & n6030;
  assign n11931 = pi84  & n5737;
  assign n11932 = pi83  & n5732;
  assign n11933 = ~n11931 & ~n11932;
  assign n11934 = ~n11930 & n11933;
  assign n11935 = ~n11929 & n11934;
  assign n11936 = pi41  & ~n11935;
  assign n11937 = pi41  & ~n11936;
  assign n11938 = ~n11935 & ~n11936;
  assign n11939 = ~n11937 & ~n11938;
  assign n11940 = ~n11928 & ~n11939;
  assign n11941 = ~n11928 & ~n11940;
  assign n11942 = ~n11939 & ~n11940;
  assign n11943 = ~n11941 & ~n11942;
  assign n11944 = ~n11584 & n11943;
  assign n11945 = n11584 & ~n11943;
  assign n11946 = ~n11944 & ~n11945;
  assign n11947 = n2288 & n5008;
  assign n11948 = pi85  & n5241;
  assign n11949 = pi87  & n5006;
  assign n11950 = pi86  & n5001;
  assign n11951 = ~n11949 & ~n11950;
  assign n11952 = ~n11948 & n11951;
  assign n11953 = ~n11947 & n11952;
  assign n11954 = pi38  & ~n11953;
  assign n11955 = pi38  & ~n11954;
  assign n11956 = ~n11953 & ~n11954;
  assign n11957 = ~n11955 & ~n11956;
  assign n11958 = ~n11946 & ~n11957;
  assign n11959 = n11946 & n11957;
  assign n11960 = ~n11958 & ~n11959;
  assign n11961 = n11818 & ~n11960;
  assign n11962 = ~n11818 & n11960;
  assign n11963 = ~n11961 & ~n11962;
  assign n11964 = n2801 & n4271;
  assign n11965 = pi88  & n4503;
  assign n11966 = pi90  & n4269;
  assign n11967 = pi89  & n4264;
  assign n11968 = ~n11966 & ~n11967;
  assign n11969 = ~n11965 & n11968;
  assign n11970 = ~n11964 & n11969;
  assign n11971 = pi35  & ~n11970;
  assign n11972 = pi35  & ~n11971;
  assign n11973 = ~n11970 & ~n11971;
  assign n11974 = ~n11972 & ~n11973;
  assign n11975 = n11963 & ~n11974;
  assign n11976 = n11963 & ~n11975;
  assign n11977 = ~n11974 & ~n11975;
  assign n11978 = ~n11976 & ~n11977;
  assign n11979 = ~n11617 & ~n11623;
  assign n11980 = n11978 & n11979;
  assign n11981 = ~n11978 & ~n11979;
  assign n11982 = ~n11980 & ~n11981;
  assign n11983 = n3371 & n3622;
  assign n11984 = pi91  & n3814;
  assign n11985 = pi93  & n3620;
  assign n11986 = pi92  & n3615;
  assign n11987 = ~n11985 & ~n11986;
  assign n11988 = ~n11984 & n11987;
  assign n11989 = ~n11983 & n11988;
  assign n11990 = pi32  & ~n11989;
  assign n11991 = pi32  & ~n11990;
  assign n11992 = ~n11989 & ~n11990;
  assign n11993 = ~n11991 & ~n11992;
  assign n11994 = n11982 & ~n11993;
  assign n11995 = ~n11982 & n11993;
  assign n11996 = ~n11994 & ~n11995;
  assign n11997 = ~n11817 & n11996;
  assign n11998 = ~n11817 & ~n11997;
  assign n11999 = ~n11994 & ~n11997;
  assign n12000 = ~n11995 & n11999;
  assign n12001 = ~n11998 & ~n12000;
  assign n12002 = n3034 & n4001;
  assign n12003 = pi94  & n3225;
  assign n12004 = pi96  & n3032;
  assign n12005 = pi95  & n3027;
  assign n12006 = ~n12004 & ~n12005;
  assign n12007 = ~n12003 & n12006;
  assign n12008 = ~n12002 & n12007;
  assign n12009 = pi29  & ~n12008;
  assign n12010 = pi29  & ~n12009;
  assign n12011 = ~n12008 & ~n12009;
  assign n12012 = ~n12010 & ~n12011;
  assign n12013 = n12001 & n12012;
  assign n12014 = ~n12001 & ~n12012;
  assign n12015 = ~n12013 & ~n12014;
  assign n12016 = ~n11815 & n12015;
  assign n12017 = n11815 & ~n12015;
  assign n12018 = ~n12016 & ~n12017;
  assign n12019 = n2523 & n4684;
  assign n12020 = pi97  & n2667;
  assign n12021 = pi99  & n2521;
  assign n12022 = pi98  & n2516;
  assign n12023 = ~n12021 & ~n12022;
  assign n12024 = ~n12020 & n12023;
  assign n12025 = ~n12019 & n12024;
  assign n12026 = pi26  & ~n12025;
  assign n12027 = pi26  & ~n12026;
  assign n12028 = ~n12025 & ~n12026;
  assign n12029 = ~n12027 & ~n12028;
  assign n12030 = n12018 & ~n12029;
  assign n12031 = n12018 & ~n12030;
  assign n12032 = ~n12029 & ~n12030;
  assign n12033 = ~n12031 & ~n12032;
  assign n12034 = ~n11671 & ~n11678;
  assign n12035 = n12033 & n12034;
  assign n12036 = ~n12033 & ~n12034;
  assign n12037 = ~n12035 & ~n12036;
  assign n12038 = n2043 & n5413;
  assign n12039 = pi100  & n2180;
  assign n12040 = pi102  & n2041;
  assign n12041 = pi101  & n2036;
  assign n12042 = ~n12040 & ~n12041;
  assign n12043 = ~n12039 & n12042;
  assign n12044 = ~n12038 & n12043;
  assign n12045 = pi23  & ~n12044;
  assign n12046 = pi23  & ~n12045;
  assign n12047 = ~n12044 & ~n12045;
  assign n12048 = ~n12046 & ~n12047;
  assign n12049 = n12037 & ~n12048;
  assign n12050 = n12037 & ~n12049;
  assign n12051 = ~n12048 & ~n12049;
  assign n12052 = ~n12050 & ~n12051;
  assign n12053 = ~n11691 & ~n11697;
  assign n12054 = n12052 & n12053;
  assign n12055 = ~n12052 & ~n12053;
  assign n12056 = ~n12054 & ~n12055;
  assign n12057 = n1611 & n6207;
  assign n12058 = pi103  & n1745;
  assign n12059 = pi105  & n1609;
  assign n12060 = pi104  & n1604;
  assign n12061 = ~n12059 & ~n12060;
  assign n12062 = ~n12058 & n12061;
  assign n12063 = ~n12057 & n12062;
  assign n12064 = pi20  & ~n12063;
  assign n12065 = pi20  & ~n12064;
  assign n12066 = ~n12063 & ~n12064;
  assign n12067 = ~n12065 & ~n12066;
  assign n12068 = n12056 & ~n12067;
  assign n12069 = ~n12056 & n12067;
  assign n12070 = ~n12068 & ~n12069;
  assign n12071 = ~n11814 & n12070;
  assign n12072 = ~n11814 & ~n12071;
  assign n12073 = ~n12068 & ~n12071;
  assign n12074 = ~n12069 & n12073;
  assign n12075 = ~n12072 & ~n12074;
  assign n12076 = n1297 & n7060;
  assign n12077 = pi106  & n1366;
  assign n12078 = pi108  & n1295;
  assign n12079 = pi107  & n1290;
  assign n12080 = ~n12078 & ~n12079;
  assign n12081 = ~n12077 & n12080;
  assign n12082 = ~n12076 & n12081;
  assign n12083 = pi17  & ~n12082;
  assign n12084 = pi17  & ~n12083;
  assign n12085 = ~n12082 & ~n12083;
  assign n12086 = ~n12084 & ~n12085;
  assign n12087 = ~n12075 & ~n12086;
  assign n12088 = ~n12075 & ~n12087;
  assign n12089 = ~n12086 & ~n12087;
  assign n12090 = ~n12088 & ~n12089;
  assign n12091 = ~n11734 & n12090;
  assign n12092 = n11734 & ~n12090;
  assign n12093 = ~n12091 & ~n12092;
  assign n12094 = n938 & n7970;
  assign n12095 = pi109  & n1052;
  assign n12096 = pi111  & n936;
  assign n12097 = pi110  & n931;
  assign n12098 = ~n12096 & ~n12097;
  assign n12099 = ~n12095 & n12098;
  assign n12100 = ~n12094 & n12099;
  assign n12101 = pi14  & ~n12100;
  assign n12102 = pi14  & ~n12101;
  assign n12103 = ~n12100 & ~n12101;
  assign n12104 = ~n12102 & ~n12103;
  assign n12105 = ~n12093 & ~n12104;
  assign n12106 = n12093 & n12104;
  assign n12107 = ~n12105 & ~n12106;
  assign n12108 = ~n11813 & n12107;
  assign n12109 = n11813 & ~n12107;
  assign n12110 = ~n12108 & ~n12109;
  assign n12111 = n687 & n8936;
  assign n12112 = pi112  & n763;
  assign n12113 = pi114  & n685;
  assign n12114 = pi113  & n680;
  assign n12115 = ~n12113 & ~n12114;
  assign n12116 = ~n12112 & n12115;
  assign n12117 = ~n12111 & n12116;
  assign n12118 = pi11  & ~n12117;
  assign n12119 = pi11  & ~n12118;
  assign n12120 = ~n12117 & ~n12118;
  assign n12121 = ~n12119 & ~n12120;
  assign n12122 = n12110 & ~n12121;
  assign n12123 = n12110 & ~n12122;
  assign n12124 = ~n12121 & ~n12122;
  assign n12125 = ~n12123 & ~n12124;
  assign n12126 = ~n11812 & ~n12125;
  assign n12127 = n11812 & n12125;
  assign n12128 = ~n12126 & ~n12127;
  assign n12129 = ~n11811 & n12128;
  assign n12130 = ~n11811 & ~n12129;
  assign n12131 = n12128 & ~n12129;
  assign n12132 = ~n12130 & ~n12131;
  assign n12133 = ~n11800 & ~n12132;
  assign n12134 = ~n11800 & ~n12133;
  assign n12135 = ~n12132 & ~n12133;
  assign n12136 = ~n12134 & ~n12135;
  assign n12137 = n342 & n11028;
  assign n12138 = pi118  & n380;
  assign n12139 = pi120  & n340;
  assign n12140 = pi119  & n335;
  assign n12141 = ~n12139 & ~n12140;
  assign n12142 = ~n12138 & n12141;
  assign n12143 = ~n12137 & n12142;
  assign n12144 = pi5  & ~n12143;
  assign n12145 = pi5  & ~n12144;
  assign n12146 = ~n12143 & ~n12144;
  assign n12147 = ~n12145 & ~n12146;
  assign n12148 = ~n12136 & ~n12147;
  assign n12149 = ~n12136 & ~n12148;
  assign n12150 = ~n12147 & ~n12148;
  assign n12151 = ~n12149 & ~n12150;
  assign n12152 = ~n11774 & ~n11776;
  assign n12153 = ~pi122  & ~pi123 ;
  assign n12154 = pi122  & pi123 ;
  assign n12155 = ~n12153 & ~n12154;
  assign n12156 = ~n12152 & n12155;
  assign n12157 = n12152 & ~n12155;
  assign n12158 = ~n12156 & ~n12157;
  assign n12159 = n262 & n12158;
  assign n12160 = pi121  & n288;
  assign n12161 = pi123  & n267;
  assign n12162 = pi122  & n269;
  assign n12163 = ~n12161 & ~n12162;
  assign n12164 = ~n12160 & n12163;
  assign n12165 = ~n12159 & n12164;
  assign n12166 = pi2  & ~n12165;
  assign n12167 = pi2  & ~n12166;
  assign n12168 = ~n12165 & ~n12166;
  assign n12169 = ~n12167 & ~n12168;
  assign n12170 = ~n12151 & n12169;
  assign n12171 = n12151 & ~n12169;
  assign n12172 = ~n12170 & ~n12171;
  assign n12173 = ~n11799 & ~n12172;
  assign n12174 = ~n11799 & ~n12173;
  assign n12175 = ~n12172 & ~n12173;
  assign n12176 = ~n12174 & ~n12175;
  assign n12177 = ~n11798 & ~n12176;
  assign n12178 = n11798 & n12176;
  assign po59  = ~n12177 & ~n12178;
  assign n12180 = ~n12173 & ~n12177;
  assign n12181 = ~n12151 & ~n12169;
  assign n12182 = ~n12148 & ~n12181;
  assign n12183 = ~n12154 & ~n12156;
  assign n12184 = ~pi123  & ~pi124 ;
  assign n12185 = pi123  & pi124 ;
  assign n12186 = ~n12184 & ~n12185;
  assign n12187 = ~n12183 & n12186;
  assign n12188 = n12183 & ~n12186;
  assign n12189 = ~n12187 & ~n12188;
  assign n12190 = n262 & n12189;
  assign n12191 = pi122  & n288;
  assign n12192 = pi124  & n267;
  assign n12193 = pi123  & n269;
  assign n12194 = ~n12192 & ~n12193;
  assign n12195 = ~n12191 & n12194;
  assign n12196 = ~n12190 & n12195;
  assign n12197 = pi2  & ~n12196;
  assign n12198 = pi2  & ~n12197;
  assign n12199 = ~n12196 & ~n12197;
  assign n12200 = ~n12198 & ~n12199;
  assign n12201 = n342 & n11389;
  assign n12202 = pi119  & n380;
  assign n12203 = pi121  & n340;
  assign n12204 = pi120  & n335;
  assign n12205 = ~n12203 & ~n12204;
  assign n12206 = ~n12202 & n12205;
  assign n12207 = ~n12201 & n12206;
  assign n12208 = pi5  & ~n12207;
  assign n12209 = pi5  & ~n12208;
  assign n12210 = ~n12207 & ~n12208;
  assign n12211 = ~n12209 & ~n12210;
  assign n12212 = ~n12129 & ~n12133;
  assign n12213 = n498 & n9984;
  assign n12214 = pi116  & n537;
  assign n12215 = pi118  & n496;
  assign n12216 = pi117  & n491;
  assign n12217 = ~n12215 & ~n12216;
  assign n12218 = ~n12214 & n12217;
  assign n12219 = ~n12213 & n12218;
  assign n12220 = pi8  & ~n12219;
  assign n12221 = pi8  & ~n12220;
  assign n12222 = ~n12219 & ~n12220;
  assign n12223 = ~n12221 & ~n12222;
  assign n12224 = ~n12122 & ~n12126;
  assign n12225 = n687 & n8963;
  assign n12226 = pi113  & n763;
  assign n12227 = pi115  & n685;
  assign n12228 = pi114  & n680;
  assign n12229 = ~n12227 & ~n12228;
  assign n12230 = ~n12226 & n12229;
  assign n12231 = ~n12225 & n12230;
  assign n12232 = pi11  & ~n12231;
  assign n12233 = pi11  & ~n12232;
  assign n12234 = ~n12231 & ~n12232;
  assign n12235 = ~n12233 & ~n12234;
  assign n12236 = ~n12105 & ~n12108;
  assign n12237 = n938 & n7997;
  assign n12238 = pi110  & n1052;
  assign n12239 = pi112  & n936;
  assign n12240 = pi111  & n931;
  assign n12241 = ~n12239 & ~n12240;
  assign n12242 = ~n12238 & n12241;
  assign n12243 = ~n12237 & n12242;
  assign n12244 = pi14  & ~n12243;
  assign n12245 = pi14  & ~n12244;
  assign n12246 = ~n12243 & ~n12244;
  assign n12247 = ~n12245 & ~n12246;
  assign n12248 = ~n11734 & ~n12090;
  assign n12249 = ~n12087 & ~n12248;
  assign n12250 = n1297 & n7349;
  assign n12251 = pi107  & n1366;
  assign n12252 = pi109  & n1295;
  assign n12253 = pi108  & n1290;
  assign n12254 = ~n12252 & ~n12253;
  assign n12255 = ~n12251 & n12254;
  assign n12256 = ~n12250 & n12255;
  assign n12257 = pi17  & ~n12256;
  assign n12258 = pi17  & ~n12257;
  assign n12259 = ~n12256 & ~n12257;
  assign n12260 = ~n12258 & ~n12259;
  assign n12261 = ~n12030 & ~n12036;
  assign n12262 = ~n12014 & ~n12016;
  assign n12263 = ~n11584 & ~n11943;
  assign n12264 = ~n11940 & ~n12263;
  assign n12265 = n1972 & n5739;
  assign n12266 = pi83  & n6030;
  assign n12267 = pi85  & n5737;
  assign n12268 = pi84  & n5732;
  assign n12269 = ~n12267 & ~n12268;
  assign n12270 = ~n12266 & n12269;
  assign n12271 = ~n12265 & n12270;
  assign n12272 = pi41  & ~n12271;
  assign n12273 = pi41  & ~n12272;
  assign n12274 = ~n12271 & ~n12272;
  assign n12275 = ~n12273 & ~n12274;
  assign n12276 = ~n11921 & ~n11925;
  assign n12277 = n1554 & n6539;
  assign n12278 = pi80  & n6873;
  assign n12279 = pi82  & n6537;
  assign n12280 = pi81  & n6532;
  assign n12281 = ~n12279 & ~n12280;
  assign n12282 = ~n12278 & n12281;
  assign n12283 = ~n12277 & n12282;
  assign n12284 = pi44  & ~n12283;
  assign n12285 = pi44  & ~n12284;
  assign n12286 = ~n12283 & ~n12284;
  assign n12287 = ~n12285 & ~n12286;
  assign n12288 = ~n11914 & ~n11918;
  assign n12289 = n1122 & n7408;
  assign n12290 = pi77  & n7740;
  assign n12291 = pi79  & n7406;
  assign n12292 = pi78  & n7401;
  assign n12293 = ~n12291 & ~n12292;
  assign n12294 = ~n12290 & n12293;
  assign n12295 = ~n12289 & n12294;
  assign n12296 = pi47  & ~n12295;
  assign n12297 = pi47  & ~n12296;
  assign n12298 = ~n12295 & ~n12296;
  assign n12299 = ~n12297 & ~n12298;
  assign n12300 = ~n11898 & ~n11900;
  assign n12301 = n891 & n8334;
  assign n12302 = pi74  & n8685;
  assign n12303 = pi76  & n8332;
  assign n12304 = pi75  & n8327;
  assign n12305 = ~n12303 & ~n12304;
  assign n12306 = ~n12302 & n12305;
  assign n12307 = ~n12301 & n12306;
  assign n12308 = pi50  & ~n12307;
  assign n12309 = pi50  & ~n12308;
  assign n12310 = ~n12307 & ~n12308;
  assign n12311 = ~n12309 & ~n12310;
  assign n12312 = ~n11892 & ~n11894;
  assign n12313 = pi59  & ~pi60 ;
  assign n12314 = ~pi59  & pi60 ;
  assign n12315 = ~n12313 & ~n12314;
  assign n12316 = pi64  & ~n12315;
  assign n12317 = ~n11859 & n12316;
  assign n12318 = n11859 & ~n12316;
  assign n12319 = ~n12317 & ~n12318;
  assign n12320 = n309 & n11488;
  assign n12321 = pi65  & n11847;
  assign n12322 = pi67  & n11486;
  assign n12323 = pi66  & n11481;
  assign n12324 = ~n12322 & ~n12323;
  assign n12325 = ~n12321 & n12324;
  assign n12326 = ~n12320 & n12325;
  assign n12327 = pi59  & ~n12326;
  assign n12328 = pi59  & ~n12327;
  assign n12329 = ~n12326 & ~n12327;
  assign n12330 = ~n12328 & ~n12329;
  assign n12331 = ~n12319 & ~n12330;
  assign n12332 = n12319 & n12330;
  assign n12333 = ~n12331 & ~n12332;
  assign n12334 = n450 & n10394;
  assign n12335 = pi68  & n10744;
  assign n12336 = pi70  & n10392;
  assign n12337 = pi69  & n10387;
  assign n12338 = ~n12336 & ~n12337;
  assign n12339 = ~n12335 & n12338;
  assign n12340 = ~n12334 & n12339;
  assign n12341 = pi56  & ~n12340;
  assign n12342 = pi56  & ~n12341;
  assign n12343 = ~n12340 & ~n12341;
  assign n12344 = ~n12342 & ~n12343;
  assign n12345 = n12333 & ~n12344;
  assign n12346 = n12333 & ~n12345;
  assign n12347 = ~n12344 & ~n12345;
  assign n12348 = ~n12346 & ~n12347;
  assign n12349 = ~n11877 & n12348;
  assign n12350 = n11877 & ~n12348;
  assign n12351 = ~n12349 & ~n12350;
  assign n12352 = n642 & n9310;
  assign n12353 = pi71  & n9701;
  assign n12354 = pi73  & n9308;
  assign n12355 = pi72  & n9303;
  assign n12356 = ~n12354 & ~n12355;
  assign n12357 = ~n12353 & n12356;
  assign n12358 = ~n12352 & n12357;
  assign n12359 = pi53  & ~n12358;
  assign n12360 = pi53  & ~n12359;
  assign n12361 = ~n12358 & ~n12359;
  assign n12362 = ~n12360 & ~n12361;
  assign n12363 = ~n12351 & ~n12362;
  assign n12364 = n12351 & n12362;
  assign n12365 = ~n12363 & ~n12364;
  assign n12366 = ~n12312 & n12365;
  assign n12367 = n12312 & ~n12365;
  assign n12368 = ~n12366 & ~n12367;
  assign n12369 = n12311 & ~n12368;
  assign n12370 = ~n12311 & n12368;
  assign n12371 = ~n12369 & ~n12370;
  assign n12372 = ~n12300 & n12371;
  assign n12373 = n12300 & ~n12371;
  assign n12374 = ~n12372 & ~n12373;
  assign n12375 = ~n12299 & n12374;
  assign n12376 = n12299 & ~n12374;
  assign n12377 = ~n12375 & ~n12376;
  assign n12378 = ~n12288 & n12377;
  assign n12379 = n12288 & ~n12377;
  assign n12380 = ~n12378 & ~n12379;
  assign n12381 = ~n12287 & n12380;
  assign n12382 = ~n12287 & ~n12381;
  assign n12383 = n12380 & ~n12381;
  assign n12384 = ~n12382 & ~n12383;
  assign n12385 = ~n12276 & ~n12384;
  assign n12386 = n12276 & n12384;
  assign n12387 = ~n12385 & ~n12386;
  assign n12388 = ~n12275 & n12387;
  assign n12389 = n12275 & ~n12387;
  assign n12390 = ~n12388 & ~n12389;
  assign n12391 = ~n12264 & n12390;
  assign n12392 = n12264 & ~n12390;
  assign n12393 = ~n12391 & ~n12392;
  assign n12394 = n2446 & n5008;
  assign n12395 = pi86  & n5241;
  assign n12396 = pi88  & n5006;
  assign n12397 = pi87  & n5001;
  assign n12398 = ~n12396 & ~n12397;
  assign n12399 = ~n12395 & n12398;
  assign n12400 = ~n12394 & n12399;
  assign n12401 = pi38  & ~n12400;
  assign n12402 = pi38  & ~n12401;
  assign n12403 = ~n12400 & ~n12401;
  assign n12404 = ~n12402 & ~n12403;
  assign n12405 = n12393 & ~n12404;
  assign n12406 = n12393 & ~n12405;
  assign n12407 = ~n12404 & ~n12405;
  assign n12408 = ~n12406 & ~n12407;
  assign n12409 = ~n11958 & ~n11962;
  assign n12410 = n12408 & n12409;
  assign n12411 = ~n12408 & ~n12409;
  assign n12412 = ~n12410 & ~n12411;
  assign n12413 = n2978 & n4271;
  assign n12414 = pi89  & n4503;
  assign n12415 = pi91  & n4269;
  assign n12416 = pi90  & n4264;
  assign n12417 = ~n12415 & ~n12416;
  assign n12418 = ~n12414 & n12417;
  assign n12419 = ~n12413 & n12418;
  assign n12420 = pi35  & ~n12419;
  assign n12421 = pi35  & ~n12420;
  assign n12422 = ~n12419 & ~n12420;
  assign n12423 = ~n12421 & ~n12422;
  assign n12424 = n12412 & ~n12423;
  assign n12425 = n12412 & ~n12424;
  assign n12426 = ~n12423 & ~n12424;
  assign n12427 = ~n12425 & ~n12426;
  assign n12428 = ~n11975 & ~n11981;
  assign n12429 = n12427 & n12428;
  assign n12430 = ~n12427 & ~n12428;
  assign n12431 = ~n12429 & ~n12430;
  assign n12432 = n3565 & n3622;
  assign n12433 = pi92  & n3814;
  assign n12434 = pi94  & n3620;
  assign n12435 = pi93  & n3615;
  assign n12436 = ~n12434 & ~n12435;
  assign n12437 = ~n12433 & n12436;
  assign n12438 = ~n12432 & n12437;
  assign n12439 = pi32  & ~n12438;
  assign n12440 = pi32  & ~n12439;
  assign n12441 = ~n12438 & ~n12439;
  assign n12442 = ~n12440 & ~n12441;
  assign n12443 = ~n12431 & n12442;
  assign n12444 = n12431 & ~n12442;
  assign n12445 = ~n12443 & ~n12444;
  assign n12446 = ~n11999 & n12445;
  assign n12447 = n11999 & ~n12445;
  assign n12448 = ~n12446 & ~n12447;
  assign n12449 = n3034 & n4211;
  assign n12450 = pi95  & n3225;
  assign n12451 = pi97  & n3032;
  assign n12452 = pi96  & n3027;
  assign n12453 = ~n12451 & ~n12452;
  assign n12454 = ~n12450 & n12453;
  assign n12455 = ~n12449 & n12454;
  assign n12456 = pi29  & ~n12455;
  assign n12457 = pi29  & ~n12456;
  assign n12458 = ~n12455 & ~n12456;
  assign n12459 = ~n12457 & ~n12458;
  assign n12460 = n12448 & ~n12459;
  assign n12461 = n12448 & ~n12460;
  assign n12462 = ~n12459 & ~n12460;
  assign n12463 = ~n12461 & ~n12462;
  assign n12464 = ~n12262 & n12463;
  assign n12465 = n12262 & ~n12463;
  assign n12466 = ~n12464 & ~n12465;
  assign n12467 = n2523 & n4910;
  assign n12468 = pi98  & n2667;
  assign n12469 = pi100  & n2521;
  assign n12470 = pi99  & n2516;
  assign n12471 = ~n12469 & ~n12470;
  assign n12472 = ~n12468 & n12471;
  assign n12473 = ~n12467 & n12472;
  assign n12474 = pi26  & ~n12473;
  assign n12475 = pi26  & ~n12474;
  assign n12476 = ~n12473 & ~n12474;
  assign n12477 = ~n12475 & ~n12476;
  assign n12478 = ~n12466 & ~n12477;
  assign n12479 = n12466 & n12477;
  assign n12480 = ~n12478 & ~n12479;
  assign n12481 = n12261 & ~n12480;
  assign n12482 = ~n12261 & n12480;
  assign n12483 = ~n12481 & ~n12482;
  assign n12484 = n2043 & n5664;
  assign n12485 = pi101  & n2180;
  assign n12486 = pi103  & n2041;
  assign n12487 = pi102  & n2036;
  assign n12488 = ~n12486 & ~n12487;
  assign n12489 = ~n12485 & n12488;
  assign n12490 = ~n12484 & n12489;
  assign n12491 = pi23  & ~n12490;
  assign n12492 = pi23  & ~n12491;
  assign n12493 = ~n12490 & ~n12491;
  assign n12494 = ~n12492 & ~n12493;
  assign n12495 = n12483 & ~n12494;
  assign n12496 = n12483 & ~n12495;
  assign n12497 = ~n12494 & ~n12495;
  assign n12498 = ~n12496 & ~n12497;
  assign n12499 = ~n12049 & ~n12055;
  assign n12500 = n12498 & n12499;
  assign n12501 = ~n12498 & ~n12499;
  assign n12502 = ~n12500 & ~n12501;
  assign n12503 = n1611 & n6477;
  assign n12504 = pi104  & n1745;
  assign n12505 = pi106  & n1609;
  assign n12506 = pi105  & n1604;
  assign n12507 = ~n12505 & ~n12506;
  assign n12508 = ~n12504 & n12507;
  assign n12509 = ~n12503 & n12508;
  assign n12510 = pi20  & ~n12509;
  assign n12511 = pi20  & ~n12510;
  assign n12512 = ~n12509 & ~n12510;
  assign n12513 = ~n12511 & ~n12512;
  assign n12514 = ~n12502 & n12513;
  assign n12515 = n12502 & ~n12513;
  assign n12516 = ~n12514 & ~n12515;
  assign n12517 = ~n12073 & n12516;
  assign n12518 = n12073 & ~n12516;
  assign n12519 = ~n12517 & ~n12518;
  assign n12520 = ~n12260 & n12519;
  assign n12521 = ~n12260 & ~n12520;
  assign n12522 = n12519 & ~n12520;
  assign n12523 = ~n12521 & ~n12522;
  assign n12524 = ~n12249 & ~n12523;
  assign n12525 = n12249 & n12523;
  assign n12526 = ~n12524 & ~n12525;
  assign n12527 = ~n12247 & n12526;
  assign n12528 = ~n12247 & ~n12527;
  assign n12529 = n12526 & ~n12527;
  assign n12530 = ~n12528 & ~n12529;
  assign n12531 = ~n12236 & ~n12530;
  assign n12532 = n12236 & n12530;
  assign n12533 = ~n12531 & ~n12532;
  assign n12534 = ~n12235 & n12533;
  assign n12535 = ~n12235 & ~n12534;
  assign n12536 = n12533 & ~n12534;
  assign n12537 = ~n12535 & ~n12536;
  assign n12538 = ~n12224 & ~n12537;
  assign n12539 = n12224 & n12537;
  assign n12540 = ~n12538 & ~n12539;
  assign n12541 = ~n12223 & n12540;
  assign n12542 = n12223 & ~n12540;
  assign n12543 = ~n12541 & ~n12542;
  assign n12544 = ~n12212 & n12543;
  assign n12545 = n12212 & ~n12543;
  assign n12546 = ~n12544 & ~n12545;
  assign n12547 = ~n12211 & n12546;
  assign n12548 = n12211 & ~n12546;
  assign n12549 = ~n12547 & ~n12548;
  assign n12550 = ~n12200 & n12549;
  assign n12551 = n12200 & ~n12549;
  assign n12552 = ~n12550 & ~n12551;
  assign n12553 = ~n12182 & n12552;
  assign n12554 = n12182 & ~n12552;
  assign n12555 = ~n12553 & ~n12554;
  assign n12556 = ~n12180 & n12555;
  assign n12557 = n12180 & ~n12555;
  assign po60  = ~n12556 & ~n12557;
  assign n12559 = ~n12534 & ~n12538;
  assign n12560 = n687 & n9614;
  assign n12561 = pi114  & n763;
  assign n12562 = pi116  & n685;
  assign n12563 = pi115  & n680;
  assign n12564 = ~n12562 & ~n12563;
  assign n12565 = ~n12561 & n12564;
  assign n12566 = ~n12560 & n12565;
  assign n12567 = pi11  & ~n12566;
  assign n12568 = pi11  & ~n12567;
  assign n12569 = ~n12566 & ~n12567;
  assign n12570 = ~n12568 & ~n12569;
  assign n12571 = ~n12527 & ~n12531;
  assign n12572 = n938 & n8612;
  assign n12573 = pi111  & n1052;
  assign n12574 = pi113  & n936;
  assign n12575 = pi112  & n931;
  assign n12576 = ~n12574 & ~n12575;
  assign n12577 = ~n12573 & n12576;
  assign n12578 = ~n12572 & n12577;
  assign n12579 = pi14  & ~n12578;
  assign n12580 = pi14  & ~n12579;
  assign n12581 = ~n12578 & ~n12579;
  assign n12582 = ~n12580 & ~n12581;
  assign n12583 = ~n12520 & ~n12524;
  assign n12584 = ~n12515 & ~n12517;
  assign n12585 = ~n12262 & ~n12463;
  assign n12586 = ~n12460 & ~n12585;
  assign n12587 = ~n12444 & ~n12446;
  assign n12588 = ~n12381 & ~n12385;
  assign n12589 = ~n12370 & ~n12372;
  assign n12590 = ~n11877 & ~n12348;
  assign n12591 = ~n12345 & ~n12590;
  assign n12592 = n475 & n10394;
  assign n12593 = pi69  & n10744;
  assign n12594 = pi71  & n10392;
  assign n12595 = pi70  & n10387;
  assign n12596 = ~n12594 & ~n12595;
  assign n12597 = ~n12593 & n12596;
  assign n12598 = ~n12592 & n12597;
  assign n12599 = pi56  & ~n12598;
  assign n12600 = pi56  & ~n12599;
  assign n12601 = ~n12598 & ~n12599;
  assign n12602 = ~n12600 & ~n12601;
  assign n12603 = n11859 & n12316;
  assign n12604 = ~n12331 & ~n12603;
  assign n12605 = n359 & n11488;
  assign n12606 = pi66  & n11847;
  assign n12607 = pi68  & n11486;
  assign n12608 = pi67  & n11481;
  assign n12609 = ~n12607 & ~n12608;
  assign n12610 = ~n12606 & n12609;
  assign n12611 = ~n12605 & n12610;
  assign n12612 = pi59  & ~n12611;
  assign n12613 = pi59  & ~n12612;
  assign n12614 = ~n12611 & ~n12612;
  assign n12615 = ~n12613 & ~n12614;
  assign n12616 = pi62  & ~n12316;
  assign n12617 = ~pi60  & pi61 ;
  assign n12618 = pi60  & ~pi61 ;
  assign n12619 = ~n12617 & ~n12618;
  assign n12620 = n12315 & ~n12619;
  assign n12621 = pi64  & n12620;
  assign n12622 = ~pi61  & pi62 ;
  assign n12623 = pi61  & ~pi62 ;
  assign n12624 = ~n12622 & ~n12623;
  assign n12625 = ~n12315 & n12624;
  assign n12626 = pi65  & n12625;
  assign n12627 = ~n12315 & ~n12624;
  assign n12628 = ~n265 & n12627;
  assign n12629 = ~n12621 & ~n12626;
  assign n12630 = ~n12628 & n12629;
  assign n12631 = pi62  & ~n12630;
  assign n12632 = pi62  & ~n12631;
  assign n12633 = ~n12630 & ~n12631;
  assign n12634 = ~n12632 & ~n12633;
  assign n12635 = n12616 & ~n12634;
  assign n12636 = ~n12616 & n12634;
  assign n12637 = ~n12635 & ~n12636;
  assign n12638 = n12615 & ~n12637;
  assign n12639 = ~n12615 & n12637;
  assign n12640 = ~n12638 & ~n12639;
  assign n12641 = ~n12604 & n12640;
  assign n12642 = n12604 & ~n12640;
  assign n12643 = ~n12641 & ~n12642;
  assign n12644 = n12602 & ~n12643;
  assign n12645 = ~n12602 & n12643;
  assign n12646 = ~n12644 & ~n12645;
  assign n12647 = ~n12591 & n12646;
  assign n12648 = n12591 & ~n12646;
  assign n12649 = ~n12647 & ~n12648;
  assign n12650 = n729 & n9310;
  assign n12651 = pi72  & n9701;
  assign n12652 = pi74  & n9308;
  assign n12653 = pi73  & n9303;
  assign n12654 = ~n12652 & ~n12653;
  assign n12655 = ~n12651 & n12654;
  assign n12656 = ~n12650 & n12655;
  assign n12657 = pi53  & ~n12656;
  assign n12658 = pi53  & ~n12657;
  assign n12659 = ~n12656 & ~n12657;
  assign n12660 = ~n12658 & ~n12659;
  assign n12661 = n12649 & ~n12660;
  assign n12662 = n12649 & ~n12661;
  assign n12663 = ~n12660 & ~n12661;
  assign n12664 = ~n12662 & ~n12663;
  assign n12665 = ~n12363 & ~n12366;
  assign n12666 = n12664 & n12665;
  assign n12667 = ~n12664 & ~n12665;
  assign n12668 = ~n12666 & ~n12667;
  assign n12669 = n999 & n8334;
  assign n12670 = pi75  & n8685;
  assign n12671 = pi77  & n8332;
  assign n12672 = pi76  & n8327;
  assign n12673 = ~n12671 & ~n12672;
  assign n12674 = ~n12670 & n12673;
  assign n12675 = ~n12669 & n12674;
  assign n12676 = pi50  & ~n12675;
  assign n12677 = pi50  & ~n12676;
  assign n12678 = ~n12675 & ~n12676;
  assign n12679 = ~n12677 & ~n12678;
  assign n12680 = n12668 & ~n12679;
  assign n12681 = ~n12668 & n12679;
  assign n12682 = ~n12680 & ~n12681;
  assign n12683 = ~n12589 & n12682;
  assign n12684 = ~n12589 & ~n12683;
  assign n12685 = ~n12680 & ~n12683;
  assign n12686 = ~n12681 & n12685;
  assign n12687 = ~n12684 & ~n12686;
  assign n12688 = n1225 & n7408;
  assign n12689 = pi78  & n7740;
  assign n12690 = pi80  & n7406;
  assign n12691 = pi79  & n7401;
  assign n12692 = ~n12690 & ~n12691;
  assign n12693 = ~n12689 & n12692;
  assign n12694 = ~n12688 & n12693;
  assign n12695 = pi47  & ~n12694;
  assign n12696 = pi47  & ~n12695;
  assign n12697 = ~n12694 & ~n12695;
  assign n12698 = ~n12696 & ~n12697;
  assign n12699 = ~n12687 & ~n12698;
  assign n12700 = ~n12687 & ~n12699;
  assign n12701 = ~n12698 & ~n12699;
  assign n12702 = ~n12700 & ~n12701;
  assign n12703 = ~n12375 & ~n12378;
  assign n12704 = n12702 & n12703;
  assign n12705 = ~n12702 & ~n12703;
  assign n12706 = ~n12704 & ~n12705;
  assign n12707 = n1696 & n6539;
  assign n12708 = pi81  & n6873;
  assign n12709 = pi83  & n6537;
  assign n12710 = pi82  & n6532;
  assign n12711 = ~n12709 & ~n12710;
  assign n12712 = ~n12708 & n12711;
  assign n12713 = ~n12707 & n12712;
  assign n12714 = pi44  & ~n12713;
  assign n12715 = pi44  & ~n12714;
  assign n12716 = ~n12713 & ~n12714;
  assign n12717 = ~n12715 & ~n12716;
  assign n12718 = n12706 & ~n12717;
  assign n12719 = ~n12706 & n12717;
  assign n12720 = ~n12718 & ~n12719;
  assign n12721 = ~n12588 & n12720;
  assign n12722 = ~n12588 & ~n12721;
  assign n12723 = ~n12718 & ~n12721;
  assign n12724 = ~n12719 & n12723;
  assign n12725 = ~n12722 & ~n12724;
  assign n12726 = n2133 & n5739;
  assign n12727 = pi84  & n6030;
  assign n12728 = pi86  & n5737;
  assign n12729 = pi85  & n5732;
  assign n12730 = ~n12728 & ~n12729;
  assign n12731 = ~n12727 & n12730;
  assign n12732 = ~n12726 & n12731;
  assign n12733 = pi41  & ~n12732;
  assign n12734 = pi41  & ~n12733;
  assign n12735 = ~n12732 & ~n12733;
  assign n12736 = ~n12734 & ~n12735;
  assign n12737 = ~n12725 & ~n12736;
  assign n12738 = ~n12725 & ~n12737;
  assign n12739 = ~n12736 & ~n12737;
  assign n12740 = ~n12738 & ~n12739;
  assign n12741 = ~n12388 & ~n12391;
  assign n12742 = n12740 & n12741;
  assign n12743 = ~n12740 & ~n12741;
  assign n12744 = ~n12742 & ~n12743;
  assign n12745 = n2473 & n5008;
  assign n12746 = pi87  & n5241;
  assign n12747 = pi89  & n5006;
  assign n12748 = pi88  & n5001;
  assign n12749 = ~n12747 & ~n12748;
  assign n12750 = ~n12746 & n12749;
  assign n12751 = ~n12745 & n12750;
  assign n12752 = pi38  & ~n12751;
  assign n12753 = pi38  & ~n12752;
  assign n12754 = ~n12751 & ~n12752;
  assign n12755 = ~n12753 & ~n12754;
  assign n12756 = n12744 & ~n12755;
  assign n12757 = n12744 & ~n12756;
  assign n12758 = ~n12755 & ~n12756;
  assign n12759 = ~n12757 & ~n12758;
  assign n12760 = ~n12405 & ~n12411;
  assign n12761 = n12759 & n12760;
  assign n12762 = ~n12759 & ~n12760;
  assign n12763 = ~n12761 & ~n12762;
  assign n12764 = n3177 & n4271;
  assign n12765 = pi90  & n4503;
  assign n12766 = pi92  & n4269;
  assign n12767 = pi91  & n4264;
  assign n12768 = ~n12766 & ~n12767;
  assign n12769 = ~n12765 & n12768;
  assign n12770 = ~n12764 & n12769;
  assign n12771 = pi35  & ~n12770;
  assign n12772 = pi35  & ~n12771;
  assign n12773 = ~n12770 & ~n12771;
  assign n12774 = ~n12772 & ~n12773;
  assign n12775 = n12763 & ~n12774;
  assign n12776 = n12763 & ~n12775;
  assign n12777 = ~n12774 & ~n12775;
  assign n12778 = ~n12776 & ~n12777;
  assign n12779 = ~n12424 & ~n12430;
  assign n12780 = n12778 & n12779;
  assign n12781 = ~n12778 & ~n12779;
  assign n12782 = ~n12780 & ~n12781;
  assign n12783 = n3622 & n3784;
  assign n12784 = pi93  & n3814;
  assign n12785 = pi95  & n3620;
  assign n12786 = pi94  & n3615;
  assign n12787 = ~n12785 & ~n12786;
  assign n12788 = ~n12784 & n12787;
  assign n12789 = ~n12783 & n12788;
  assign n12790 = pi32  & ~n12789;
  assign n12791 = pi32  & ~n12790;
  assign n12792 = ~n12789 & ~n12790;
  assign n12793 = ~n12791 & ~n12792;
  assign n12794 = n12782 & ~n12793;
  assign n12795 = n12782 & ~n12794;
  assign n12796 = ~n12793 & ~n12794;
  assign n12797 = ~n12795 & ~n12796;
  assign n12798 = ~n12587 & n12797;
  assign n12799 = n12587 & ~n12797;
  assign n12800 = ~n12798 & ~n12799;
  assign n12801 = n3034 & n4454;
  assign n12802 = pi96  & n3225;
  assign n12803 = pi98  & n3032;
  assign n12804 = pi97  & n3027;
  assign n12805 = ~n12803 & ~n12804;
  assign n12806 = ~n12802 & n12805;
  assign n12807 = ~n12801 & n12806;
  assign n12808 = pi29  & ~n12807;
  assign n12809 = pi29  & ~n12808;
  assign n12810 = ~n12807 & ~n12808;
  assign n12811 = ~n12809 & ~n12810;
  assign n12812 = ~n12800 & ~n12811;
  assign n12813 = n12800 & n12811;
  assign n12814 = ~n12812 & ~n12813;
  assign n12815 = n12586 & ~n12814;
  assign n12816 = ~n12586 & n12814;
  assign n12817 = ~n12815 & ~n12816;
  assign n12818 = n2523 & n5169;
  assign n12819 = pi99  & n2667;
  assign n12820 = pi101  & n2521;
  assign n12821 = pi100  & n2516;
  assign n12822 = ~n12820 & ~n12821;
  assign n12823 = ~n12819 & n12822;
  assign n12824 = ~n12818 & n12823;
  assign n12825 = pi26  & ~n12824;
  assign n12826 = pi26  & ~n12825;
  assign n12827 = ~n12824 & ~n12825;
  assign n12828 = ~n12826 & ~n12827;
  assign n12829 = n12817 & ~n12828;
  assign n12830 = n12817 & ~n12829;
  assign n12831 = ~n12828 & ~n12829;
  assign n12832 = ~n12830 & ~n12831;
  assign n12833 = ~n12478 & ~n12482;
  assign n12834 = n12832 & n12833;
  assign n12835 = ~n12832 & ~n12833;
  assign n12836 = ~n12834 & ~n12835;
  assign n12837 = n2043 & n5943;
  assign n12838 = pi102  & n2180;
  assign n12839 = pi104  & n2041;
  assign n12840 = pi103  & n2036;
  assign n12841 = ~n12839 & ~n12840;
  assign n12842 = ~n12838 & n12841;
  assign n12843 = ~n12837 & n12842;
  assign n12844 = pi23  & ~n12843;
  assign n12845 = pi23  & ~n12844;
  assign n12846 = ~n12843 & ~n12844;
  assign n12847 = ~n12845 & ~n12846;
  assign n12848 = n12836 & ~n12847;
  assign n12849 = n12836 & ~n12848;
  assign n12850 = ~n12847 & ~n12848;
  assign n12851 = ~n12849 & ~n12850;
  assign n12852 = ~n12495 & ~n12501;
  assign n12853 = n12851 & n12852;
  assign n12854 = ~n12851 & ~n12852;
  assign n12855 = ~n12853 & ~n12854;
  assign n12856 = n1611 & n6775;
  assign n12857 = pi105  & n1745;
  assign n12858 = pi107  & n1609;
  assign n12859 = pi106  & n1604;
  assign n12860 = ~n12858 & ~n12859;
  assign n12861 = ~n12857 & n12860;
  assign n12862 = ~n12856 & n12861;
  assign n12863 = pi20  & ~n12862;
  assign n12864 = pi20  & ~n12863;
  assign n12865 = ~n12862 & ~n12863;
  assign n12866 = ~n12864 & ~n12865;
  assign n12867 = n12855 & ~n12866;
  assign n12868 = ~n12855 & n12866;
  assign n12869 = ~n12867 & ~n12868;
  assign n12870 = ~n12584 & n12869;
  assign n12871 = ~n12584 & ~n12870;
  assign n12872 = ~n12867 & ~n12870;
  assign n12873 = ~n12868 & n12872;
  assign n12874 = ~n12871 & ~n12873;
  assign n12875 = n1297 & n7665;
  assign n12876 = pi108  & n1366;
  assign n12877 = pi110  & n1295;
  assign n12878 = pi109  & n1290;
  assign n12879 = ~n12877 & ~n12878;
  assign n12880 = ~n12876 & n12879;
  assign n12881 = ~n12875 & n12880;
  assign n12882 = pi17  & ~n12881;
  assign n12883 = pi17  & ~n12882;
  assign n12884 = ~n12881 & ~n12882;
  assign n12885 = ~n12883 & ~n12884;
  assign n12886 = n12874 & n12885;
  assign n12887 = ~n12874 & ~n12885;
  assign n12888 = ~n12886 & ~n12887;
  assign n12889 = ~n12583 & n12888;
  assign n12890 = n12583 & ~n12888;
  assign n12891 = ~n12889 & ~n12890;
  assign n12892 = n12582 & ~n12891;
  assign n12893 = ~n12582 & n12891;
  assign n12894 = ~n12892 & ~n12893;
  assign n12895 = ~n12571 & n12894;
  assign n12896 = n12571 & ~n12894;
  assign n12897 = ~n12895 & ~n12896;
  assign n12898 = n12570 & ~n12897;
  assign n12899 = ~n12570 & n12897;
  assign n12900 = ~n12898 & ~n12899;
  assign n12901 = ~n12559 & n12900;
  assign n12902 = n12559 & ~n12900;
  assign n12903 = ~n12901 & ~n12902;
  assign n12904 = n498 & n10667;
  assign n12905 = pi117  & n537;
  assign n12906 = pi119  & n496;
  assign n12907 = pi118  & n491;
  assign n12908 = ~n12906 & ~n12907;
  assign n12909 = ~n12905 & n12908;
  assign n12910 = ~n12904 & n12909;
  assign n12911 = pi8  & ~n12910;
  assign n12912 = pi8  & ~n12911;
  assign n12913 = ~n12910 & ~n12911;
  assign n12914 = ~n12912 & ~n12913;
  assign n12915 = n12903 & ~n12914;
  assign n12916 = n12903 & ~n12915;
  assign n12917 = ~n12914 & ~n12915;
  assign n12918 = ~n12916 & ~n12917;
  assign n12919 = ~n12541 & ~n12544;
  assign n12920 = n12918 & n12919;
  assign n12921 = ~n12918 & ~n12919;
  assign n12922 = ~n12920 & ~n12921;
  assign n12923 = n342 & n11778;
  assign n12924 = pi120  & n380;
  assign n12925 = pi122  & n340;
  assign n12926 = pi121  & n335;
  assign n12927 = ~n12925 & ~n12926;
  assign n12928 = ~n12924 & n12927;
  assign n12929 = ~n12923 & n12928;
  assign n12930 = pi5  & ~n12929;
  assign n12931 = pi5  & ~n12930;
  assign n12932 = ~n12929 & ~n12930;
  assign n12933 = ~n12931 & ~n12932;
  assign n12934 = ~n12922 & n12933;
  assign n12935 = n12922 & ~n12933;
  assign n12936 = ~n12934 & ~n12935;
  assign n12937 = ~n12185 & ~n12187;
  assign n12938 = ~pi124  & ~pi125 ;
  assign n12939 = pi124  & pi125 ;
  assign n12940 = ~n12938 & ~n12939;
  assign n12941 = ~n12937 & n12940;
  assign n12942 = n12937 & ~n12940;
  assign n12943 = ~n12941 & ~n12942;
  assign n12944 = n262 & n12943;
  assign n12945 = pi123  & n288;
  assign n12946 = pi125  & n267;
  assign n12947 = pi124  & n269;
  assign n12948 = ~n12946 & ~n12947;
  assign n12949 = ~n12945 & n12948;
  assign n12950 = ~n12944 & n12949;
  assign n12951 = pi2  & ~n12950;
  assign n12952 = pi2  & ~n12951;
  assign n12953 = ~n12950 & ~n12951;
  assign n12954 = ~n12952 & ~n12953;
  assign n12955 = n12936 & ~n12954;
  assign n12956 = n12936 & ~n12955;
  assign n12957 = ~n12954 & ~n12955;
  assign n12958 = ~n12956 & ~n12957;
  assign n12959 = ~n12547 & ~n12550;
  assign n12960 = n12958 & n12959;
  assign n12961 = ~n12958 & ~n12959;
  assign n12962 = ~n12960 & ~n12961;
  assign n12963 = ~n12553 & ~n12556;
  assign n12964 = n12962 & ~n12963;
  assign n12965 = ~n12962 & n12963;
  assign po61  = ~n12964 & ~n12965;
  assign n12967 = ~n12961 & ~n12964;
  assign n12968 = ~n12935 & ~n12955;
  assign n12969 = ~n12899 & ~n12901;
  assign n12970 = ~n12893 & ~n12895;
  assign n12971 = ~n12887 & ~n12889;
  assign n12972 = ~n12848 & ~n12854;
  assign n12973 = ~n12587 & ~n12797;
  assign n12974 = ~n12794 & ~n12973;
  assign n12975 = ~n12737 & ~n12743;
  assign n12976 = ~n12699 & ~n12705;
  assign n12977 = n1434 & n7408;
  assign n12978 = pi79  & n7740;
  assign n12979 = pi81  & n7406;
  assign n12980 = pi80  & n7401;
  assign n12981 = ~n12979 & ~n12980;
  assign n12982 = ~n12978 & n12981;
  assign n12983 = ~n12977 & n12982;
  assign n12984 = pi47  & ~n12983;
  assign n12985 = pi47  & ~n12984;
  assign n12986 = ~n12983 & ~n12984;
  assign n12987 = ~n12985 & ~n12986;
  assign n12988 = ~n12661 & ~n12667;
  assign n12989 = n809 & n9310;
  assign n12990 = pi73  & n9701;
  assign n12991 = pi75  & n9308;
  assign n12992 = pi74  & n9303;
  assign n12993 = ~n12991 & ~n12992;
  assign n12994 = ~n12990 & n12993;
  assign n12995 = ~n12989 & n12994;
  assign n12996 = pi53  & ~n12995;
  assign n12997 = pi53  & ~n12996;
  assign n12998 = ~n12995 & ~n12996;
  assign n12999 = ~n12997 & ~n12998;
  assign n13000 = ~n12645 & ~n12647;
  assign n13001 = ~n12639 & ~n12641;
  assign n13002 = n286 & n12627;
  assign n13003 = n12315 & n12619;
  assign n13004 = ~n12624 & n13003;
  assign n13005 = pi64  & n13004;
  assign n13006 = pi66  & n12625;
  assign n13007 = pi65  & n12620;
  assign n13008 = ~n13006 & ~n13007;
  assign n13009 = ~n13002 & n13008;
  assign n13010 = ~n13005 & n13009;
  assign n13011 = pi62  & ~n13010;
  assign n13012 = pi62  & ~n13011;
  assign n13013 = ~n13010 & ~n13011;
  assign n13014 = ~n13012 & ~n13013;
  assign n13015 = ~n12635 & n13014;
  assign n13016 = n12635 & ~n13014;
  assign n13017 = ~n13015 & ~n13016;
  assign n13018 = n401 & n11488;
  assign n13019 = pi67  & n11847;
  assign n13020 = pi69  & n11486;
  assign n13021 = pi68  & n11481;
  assign n13022 = ~n13020 & ~n13021;
  assign n13023 = ~n13019 & n13022;
  assign n13024 = ~n13018 & n13023;
  assign n13025 = pi59  & ~n13024;
  assign n13026 = pi59  & ~n13025;
  assign n13027 = ~n13024 & ~n13025;
  assign n13028 = ~n13026 & ~n13027;
  assign n13029 = n13017 & ~n13028;
  assign n13030 = ~n13017 & n13028;
  assign n13031 = ~n13029 & ~n13030;
  assign n13032 = ~n13001 & n13031;
  assign n13033 = ~n13001 & ~n13032;
  assign n13034 = ~n13029 & ~n13032;
  assign n13035 = ~n13030 & n13034;
  assign n13036 = ~n13033 & ~n13035;
  assign n13037 = n576 & n10394;
  assign n13038 = pi70  & n10744;
  assign n13039 = pi72  & n10392;
  assign n13040 = pi71  & n10387;
  assign n13041 = ~n13039 & ~n13040;
  assign n13042 = ~n13038 & n13041;
  assign n13043 = ~n13037 & n13042;
  assign n13044 = pi56  & ~n13043;
  assign n13045 = pi56  & ~n13044;
  assign n13046 = ~n13043 & ~n13044;
  assign n13047 = ~n13045 & ~n13046;
  assign n13048 = n13036 & n13047;
  assign n13049 = ~n13036 & ~n13047;
  assign n13050 = ~n13048 & ~n13049;
  assign n13051 = ~n13000 & n13050;
  assign n13052 = n13000 & ~n13050;
  assign n13053 = ~n13051 & ~n13052;
  assign n13054 = n12999 & ~n13053;
  assign n13055 = ~n12999 & n13053;
  assign n13056 = ~n13054 & ~n13055;
  assign n13057 = ~n12988 & n13056;
  assign n13058 = n12988 & ~n13056;
  assign n13059 = ~n13057 & ~n13058;
  assign n13060 = n1025 & n8334;
  assign n13061 = pi76  & n8685;
  assign n13062 = pi78  & n8332;
  assign n13063 = pi77  & n8327;
  assign n13064 = ~n13062 & ~n13063;
  assign n13065 = ~n13061 & n13064;
  assign n13066 = ~n13060 & n13065;
  assign n13067 = pi50  & ~n13066;
  assign n13068 = pi50  & ~n13067;
  assign n13069 = ~n13066 & ~n13067;
  assign n13070 = ~n13068 & ~n13069;
  assign n13071 = n13059 & ~n13070;
  assign n13072 = n13059 & ~n13071;
  assign n13073 = ~n13070 & ~n13071;
  assign n13074 = ~n13072 & ~n13073;
  assign n13075 = ~n12685 & ~n13074;
  assign n13076 = n12685 & n13074;
  assign n13077 = ~n13075 & ~n13076;
  assign n13078 = ~n12987 & n13077;
  assign n13079 = ~n12987 & ~n13078;
  assign n13080 = n13077 & ~n13078;
  assign n13081 = ~n13079 & ~n13080;
  assign n13082 = ~n12976 & ~n13081;
  assign n13083 = ~n12976 & ~n13082;
  assign n13084 = ~n13081 & ~n13082;
  assign n13085 = ~n13083 & ~n13084;
  assign n13086 = n1834 & n6539;
  assign n13087 = pi82  & n6873;
  assign n13088 = pi84  & n6537;
  assign n13089 = pi83  & n6532;
  assign n13090 = ~n13088 & ~n13089;
  assign n13091 = ~n13087 & n13090;
  assign n13092 = ~n13086 & n13091;
  assign n13093 = pi44  & ~n13092;
  assign n13094 = pi44  & ~n13093;
  assign n13095 = ~n13092 & ~n13093;
  assign n13096 = ~n13094 & ~n13095;
  assign n13097 = ~n13085 & ~n13096;
  assign n13098 = ~n13085 & ~n13097;
  assign n13099 = ~n13096 & ~n13097;
  assign n13100 = ~n13098 & ~n13099;
  assign n13101 = ~n12723 & n13100;
  assign n13102 = n12723 & ~n13100;
  assign n13103 = ~n13101 & ~n13102;
  assign n13104 = n2288 & n5739;
  assign n13105 = pi85  & n6030;
  assign n13106 = pi87  & n5737;
  assign n13107 = pi86  & n5732;
  assign n13108 = ~n13106 & ~n13107;
  assign n13109 = ~n13105 & n13108;
  assign n13110 = ~n13104 & n13109;
  assign n13111 = pi41  & ~n13110;
  assign n13112 = pi41  & ~n13111;
  assign n13113 = ~n13110 & ~n13111;
  assign n13114 = ~n13112 & ~n13113;
  assign n13115 = ~n13103 & ~n13114;
  assign n13116 = n13103 & n13114;
  assign n13117 = ~n13115 & ~n13116;
  assign n13118 = n12975 & ~n13117;
  assign n13119 = ~n12975 & n13117;
  assign n13120 = ~n13118 & ~n13119;
  assign n13121 = n2801 & n5008;
  assign n13122 = pi88  & n5241;
  assign n13123 = pi90  & n5006;
  assign n13124 = pi89  & n5001;
  assign n13125 = ~n13123 & ~n13124;
  assign n13126 = ~n13122 & n13125;
  assign n13127 = ~n13121 & n13126;
  assign n13128 = pi38  & ~n13127;
  assign n13129 = pi38  & ~n13128;
  assign n13130 = ~n13127 & ~n13128;
  assign n13131 = ~n13129 & ~n13130;
  assign n13132 = n13120 & ~n13131;
  assign n13133 = n13120 & ~n13132;
  assign n13134 = ~n13131 & ~n13132;
  assign n13135 = ~n13133 & ~n13134;
  assign n13136 = ~n12756 & ~n12762;
  assign n13137 = n13135 & n13136;
  assign n13138 = ~n13135 & ~n13136;
  assign n13139 = ~n13137 & ~n13138;
  assign n13140 = n3371 & n4271;
  assign n13141 = pi91  & n4503;
  assign n13142 = pi93  & n4269;
  assign n13143 = pi92  & n4264;
  assign n13144 = ~n13142 & ~n13143;
  assign n13145 = ~n13141 & n13144;
  assign n13146 = ~n13140 & n13145;
  assign n13147 = pi35  & ~n13146;
  assign n13148 = pi35  & ~n13147;
  assign n13149 = ~n13146 & ~n13147;
  assign n13150 = ~n13148 & ~n13149;
  assign n13151 = n13139 & ~n13150;
  assign n13152 = n13139 & ~n13151;
  assign n13153 = ~n13150 & ~n13151;
  assign n13154 = ~n13152 & ~n13153;
  assign n13155 = ~n12775 & ~n12781;
  assign n13156 = n13154 & n13155;
  assign n13157 = ~n13154 & ~n13155;
  assign n13158 = ~n13156 & ~n13157;
  assign n13159 = n3622 & n4001;
  assign n13160 = pi94  & n3814;
  assign n13161 = pi96  & n3620;
  assign n13162 = pi95  & n3615;
  assign n13163 = ~n13161 & ~n13162;
  assign n13164 = ~n13160 & n13163;
  assign n13165 = ~n13159 & n13164;
  assign n13166 = pi32  & ~n13165;
  assign n13167 = pi32  & ~n13166;
  assign n13168 = ~n13165 & ~n13166;
  assign n13169 = ~n13167 & ~n13168;
  assign n13170 = n13158 & ~n13169;
  assign n13171 = ~n13158 & n13169;
  assign n13172 = ~n13170 & ~n13171;
  assign n13173 = ~n12974 & n13172;
  assign n13174 = ~n12974 & ~n13173;
  assign n13175 = ~n13170 & ~n13173;
  assign n13176 = ~n13171 & n13175;
  assign n13177 = ~n13174 & ~n13176;
  assign n13178 = n3034 & n4684;
  assign n13179 = pi97  & n3225;
  assign n13180 = pi99  & n3032;
  assign n13181 = pi98  & n3027;
  assign n13182 = ~n13180 & ~n13181;
  assign n13183 = ~n13179 & n13182;
  assign n13184 = ~n13178 & n13183;
  assign n13185 = pi29  & ~n13184;
  assign n13186 = pi29  & ~n13185;
  assign n13187 = ~n13184 & ~n13185;
  assign n13188 = ~n13186 & ~n13187;
  assign n13189 = ~n13177 & ~n13188;
  assign n13190 = ~n13177 & ~n13189;
  assign n13191 = ~n13188 & ~n13189;
  assign n13192 = ~n13190 & ~n13191;
  assign n13193 = ~n12812 & ~n12816;
  assign n13194 = n13192 & n13193;
  assign n13195 = ~n13192 & ~n13193;
  assign n13196 = ~n13194 & ~n13195;
  assign n13197 = n2523 & n5413;
  assign n13198 = pi100  & n2667;
  assign n13199 = pi102  & n2521;
  assign n13200 = pi101  & n2516;
  assign n13201 = ~n13199 & ~n13200;
  assign n13202 = ~n13198 & n13201;
  assign n13203 = ~n13197 & n13202;
  assign n13204 = pi26  & ~n13203;
  assign n13205 = pi26  & ~n13204;
  assign n13206 = ~n13203 & ~n13204;
  assign n13207 = ~n13205 & ~n13206;
  assign n13208 = n13196 & ~n13207;
  assign n13209 = n13196 & ~n13208;
  assign n13210 = ~n13207 & ~n13208;
  assign n13211 = ~n13209 & ~n13210;
  assign n13212 = ~n12829 & ~n12835;
  assign n13213 = n13211 & n13212;
  assign n13214 = ~n13211 & ~n13212;
  assign n13215 = ~n13213 & ~n13214;
  assign n13216 = n2043 & n6207;
  assign n13217 = pi103  & n2180;
  assign n13218 = pi105  & n2041;
  assign n13219 = pi104  & n2036;
  assign n13220 = ~n13218 & ~n13219;
  assign n13221 = ~n13217 & n13220;
  assign n13222 = ~n13216 & n13221;
  assign n13223 = pi23  & ~n13222;
  assign n13224 = pi23  & ~n13223;
  assign n13225 = ~n13222 & ~n13223;
  assign n13226 = ~n13224 & ~n13225;
  assign n13227 = n13215 & ~n13226;
  assign n13228 = ~n13215 & n13226;
  assign n13229 = ~n13227 & ~n13228;
  assign n13230 = ~n12972 & n13229;
  assign n13231 = ~n12972 & ~n13230;
  assign n13232 = ~n13227 & ~n13230;
  assign n13233 = ~n13228 & n13232;
  assign n13234 = ~n13231 & ~n13233;
  assign n13235 = n1611 & n7060;
  assign n13236 = pi106  & n1745;
  assign n13237 = pi108  & n1609;
  assign n13238 = pi107  & n1604;
  assign n13239 = ~n13237 & ~n13238;
  assign n13240 = ~n13236 & n13239;
  assign n13241 = ~n13235 & n13240;
  assign n13242 = pi20  & ~n13241;
  assign n13243 = pi20  & ~n13242;
  assign n13244 = ~n13241 & ~n13242;
  assign n13245 = ~n13243 & ~n13244;
  assign n13246 = ~n13234 & ~n13245;
  assign n13247 = ~n13234 & ~n13246;
  assign n13248 = ~n13245 & ~n13246;
  assign n13249 = ~n13247 & ~n13248;
  assign n13250 = ~n12872 & n13249;
  assign n13251 = n12872 & ~n13249;
  assign n13252 = ~n13250 & ~n13251;
  assign n13253 = n1297 & n7970;
  assign n13254 = pi109  & n1366;
  assign n13255 = pi111  & n1295;
  assign n13256 = pi110  & n1290;
  assign n13257 = ~n13255 & ~n13256;
  assign n13258 = ~n13254 & n13257;
  assign n13259 = ~n13253 & n13258;
  assign n13260 = pi17  & ~n13259;
  assign n13261 = pi17  & ~n13260;
  assign n13262 = ~n13259 & ~n13260;
  assign n13263 = ~n13261 & ~n13262;
  assign n13264 = ~n13252 & ~n13263;
  assign n13265 = n13252 & n13263;
  assign n13266 = ~n13264 & ~n13265;
  assign n13267 = ~n12971 & n13266;
  assign n13268 = n12971 & ~n13266;
  assign n13269 = ~n13267 & ~n13268;
  assign n13270 = n938 & n8936;
  assign n13271 = pi112  & n1052;
  assign n13272 = pi114  & n936;
  assign n13273 = pi113  & n931;
  assign n13274 = ~n13272 & ~n13273;
  assign n13275 = ~n13271 & n13274;
  assign n13276 = ~n13270 & n13275;
  assign n13277 = pi14  & ~n13276;
  assign n13278 = pi14  & ~n13277;
  assign n13279 = ~n13276 & ~n13277;
  assign n13280 = ~n13278 & ~n13279;
  assign n13281 = n13269 & ~n13280;
  assign n13282 = n13269 & ~n13281;
  assign n13283 = ~n13280 & ~n13281;
  assign n13284 = ~n13282 & ~n13283;
  assign n13285 = ~n12970 & n13284;
  assign n13286 = n12970 & ~n13284;
  assign n13287 = ~n13285 & ~n13286;
  assign n13288 = n687 & n9958;
  assign n13289 = pi115  & n763;
  assign n13290 = pi117  & n685;
  assign n13291 = pi116  & n680;
  assign n13292 = ~n13290 & ~n13291;
  assign n13293 = ~n13289 & n13292;
  assign n13294 = ~n13288 & n13293;
  assign n13295 = pi11  & ~n13294;
  assign n13296 = pi11  & ~n13295;
  assign n13297 = ~n13294 & ~n13295;
  assign n13298 = ~n13296 & ~n13297;
  assign n13299 = ~n13287 & ~n13298;
  assign n13300 = n13287 & n13298;
  assign n13301 = ~n13299 & ~n13300;
  assign n13302 = ~n12969 & n13301;
  assign n13303 = n12969 & ~n13301;
  assign n13304 = ~n13302 & ~n13303;
  assign n13305 = n498 & n11028;
  assign n13306 = pi118  & n537;
  assign n13307 = pi120  & n496;
  assign n13308 = pi119  & n491;
  assign n13309 = ~n13307 & ~n13308;
  assign n13310 = ~n13306 & n13309;
  assign n13311 = ~n13305 & n13310;
  assign n13312 = pi8  & ~n13311;
  assign n13313 = pi8  & ~n13312;
  assign n13314 = ~n13311 & ~n13312;
  assign n13315 = ~n13313 & ~n13314;
  assign n13316 = ~n13304 & n13315;
  assign n13317 = n13304 & ~n13315;
  assign n13318 = ~n13316 & ~n13317;
  assign n13319 = n342 & n12158;
  assign n13320 = pi121  & n380;
  assign n13321 = pi123  & n340;
  assign n13322 = pi122  & n335;
  assign n13323 = ~n13321 & ~n13322;
  assign n13324 = ~n13320 & n13323;
  assign n13325 = ~n13319 & n13324;
  assign n13326 = pi5  & ~n13325;
  assign n13327 = pi5  & ~n13326;
  assign n13328 = ~n13325 & ~n13326;
  assign n13329 = ~n13327 & ~n13328;
  assign n13330 = n13318 & ~n13329;
  assign n13331 = n13318 & ~n13330;
  assign n13332 = ~n13329 & ~n13330;
  assign n13333 = ~n13331 & ~n13332;
  assign n13334 = ~n12915 & ~n12921;
  assign n13335 = n13333 & n13334;
  assign n13336 = ~n13333 & ~n13334;
  assign n13337 = ~n13335 & ~n13336;
  assign n13338 = ~n12939 & ~n12941;
  assign n13339 = ~pi125  & ~pi126 ;
  assign n13340 = pi125  & pi126 ;
  assign n13341 = ~n13339 & ~n13340;
  assign n13342 = ~n13338 & n13341;
  assign n13343 = n13338 & ~n13341;
  assign n13344 = ~n13342 & ~n13343;
  assign n13345 = n262 & n13344;
  assign n13346 = pi124  & n288;
  assign n13347 = pi126  & n267;
  assign n13348 = pi125  & n269;
  assign n13349 = ~n13347 & ~n13348;
  assign n13350 = ~n13346 & n13349;
  assign n13351 = ~n13345 & n13350;
  assign n13352 = pi2  & ~n13351;
  assign n13353 = pi2  & ~n13352;
  assign n13354 = ~n13351 & ~n13352;
  assign n13355 = ~n13353 & ~n13354;
  assign n13356 = ~n13337 & n13355;
  assign n13357 = n13337 & ~n13355;
  assign n13358 = ~n13356 & ~n13357;
  assign n13359 = ~n12968 & n13358;
  assign n13360 = n12968 & ~n13358;
  assign n13361 = ~n13359 & ~n13360;
  assign n13362 = ~n12967 & n13361;
  assign n13363 = n12967 & ~n13361;
  assign po62  = ~n13362 & ~n13363;
  assign n13365 = ~n12970 & ~n13284;
  assign n13366 = ~n13281 & ~n13365;
  assign n13367 = n938 & n8963;
  assign n13368 = pi113  & n1052;
  assign n13369 = pi115  & n936;
  assign n13370 = pi114  & n931;
  assign n13371 = ~n13369 & ~n13370;
  assign n13372 = ~n13368 & n13371;
  assign n13373 = ~n13367 & n13372;
  assign n13374 = pi14  & ~n13373;
  assign n13375 = pi14  & ~n13374;
  assign n13376 = ~n13373 & ~n13374;
  assign n13377 = ~n13375 & ~n13376;
  assign n13378 = ~n13264 & ~n13267;
  assign n13379 = n1297 & n7997;
  assign n13380 = pi110  & n1366;
  assign n13381 = pi112  & n1295;
  assign n13382 = pi111  & n1290;
  assign n13383 = ~n13381 & ~n13382;
  assign n13384 = ~n13380 & n13383;
  assign n13385 = ~n13379 & n13384;
  assign n13386 = pi17  & ~n13385;
  assign n13387 = pi17  & ~n13386;
  assign n13388 = ~n13385 & ~n13386;
  assign n13389 = ~n13387 & ~n13388;
  assign n13390 = ~n12872 & ~n13249;
  assign n13391 = ~n13246 & ~n13390;
  assign n13392 = n1611 & n7349;
  assign n13393 = pi107  & n1745;
  assign n13394 = pi109  & n1609;
  assign n13395 = pi108  & n1604;
  assign n13396 = ~n13394 & ~n13395;
  assign n13397 = ~n13393 & n13396;
  assign n13398 = ~n13392 & n13397;
  assign n13399 = pi20  & ~n13398;
  assign n13400 = pi20  & ~n13399;
  assign n13401 = ~n13398 & ~n13399;
  assign n13402 = ~n13400 & ~n13401;
  assign n13403 = n2043 & n6477;
  assign n13404 = pi104  & n2180;
  assign n13405 = pi106  & n2041;
  assign n13406 = pi105  & n2036;
  assign n13407 = ~n13405 & ~n13406;
  assign n13408 = ~n13404 & n13407;
  assign n13409 = ~n13403 & n13408;
  assign n13410 = pi23  & ~n13409;
  assign n13411 = pi23  & ~n13410;
  assign n13412 = ~n13409 & ~n13410;
  assign n13413 = ~n13411 & ~n13412;
  assign n13414 = ~n13208 & ~n13214;
  assign n13415 = ~n13189 & ~n13195;
  assign n13416 = ~n12723 & ~n13100;
  assign n13417 = ~n13097 & ~n13416;
  assign n13418 = n1972 & n6539;
  assign n13419 = pi83  & n6873;
  assign n13420 = pi85  & n6537;
  assign n13421 = pi84  & n6532;
  assign n13422 = ~n13420 & ~n13421;
  assign n13423 = ~n13419 & n13422;
  assign n13424 = ~n13418 & n13423;
  assign n13425 = pi44  & ~n13424;
  assign n13426 = pi44  & ~n13425;
  assign n13427 = ~n13424 & ~n13425;
  assign n13428 = ~n13426 & ~n13427;
  assign n13429 = ~n13078 & ~n13082;
  assign n13430 = ~n13055 & ~n13057;
  assign n13431 = ~n13049 & ~n13051;
  assign n13432 = pi62  & ~pi63 ;
  assign n13433 = ~pi62  & pi63 ;
  assign n13434 = ~n13432 & ~n13433;
  assign n13435 = pi64  & ~n13434;
  assign n13436 = n13016 & n13435;
  assign n13437 = n13016 & ~n13436;
  assign n13438 = n13435 & ~n13436;
  assign n13439 = ~n13437 & ~n13438;
  assign n13440 = n309 & n12627;
  assign n13441 = pi65  & n13004;
  assign n13442 = pi67  & n12625;
  assign n13443 = pi66  & n12620;
  assign n13444 = ~n13442 & ~n13443;
  assign n13445 = ~n13441 & n13444;
  assign n13446 = ~n13440 & n13445;
  assign n13447 = pi62  & ~n13446;
  assign n13448 = pi62  & ~n13447;
  assign n13449 = ~n13446 & ~n13447;
  assign n13450 = ~n13448 & ~n13449;
  assign n13451 = ~n13439 & ~n13450;
  assign n13452 = ~n13439 & ~n13451;
  assign n13453 = ~n13450 & ~n13451;
  assign n13454 = ~n13452 & ~n13453;
  assign n13455 = n450 & n11488;
  assign n13456 = pi68  & n11847;
  assign n13457 = pi70  & n11486;
  assign n13458 = pi69  & n11481;
  assign n13459 = ~n13457 & ~n13458;
  assign n13460 = ~n13456 & n13459;
  assign n13461 = ~n13455 & n13460;
  assign n13462 = pi59  & ~n13461;
  assign n13463 = pi59  & ~n13462;
  assign n13464 = ~n13461 & ~n13462;
  assign n13465 = ~n13463 & ~n13464;
  assign n13466 = n13454 & n13465;
  assign n13467 = ~n13454 & ~n13465;
  assign n13468 = ~n13466 & ~n13467;
  assign n13469 = ~n13034 & n13468;
  assign n13470 = n13034 & ~n13468;
  assign n13471 = ~n13469 & ~n13470;
  assign n13472 = n642 & n10394;
  assign n13473 = pi71  & n10744;
  assign n13474 = pi73  & n10392;
  assign n13475 = pi72  & n10387;
  assign n13476 = ~n13474 & ~n13475;
  assign n13477 = ~n13473 & n13476;
  assign n13478 = ~n13472 & n13477;
  assign n13479 = pi56  & ~n13478;
  assign n13480 = pi56  & ~n13479;
  assign n13481 = ~n13478 & ~n13479;
  assign n13482 = ~n13480 & ~n13481;
  assign n13483 = n13471 & ~n13482;
  assign n13484 = n13471 & ~n13483;
  assign n13485 = ~n13482 & ~n13483;
  assign n13486 = ~n13484 & ~n13485;
  assign n13487 = ~n13431 & n13486;
  assign n13488 = n13431 & ~n13486;
  assign n13489 = ~n13487 & ~n13488;
  assign n13490 = n891 & n9310;
  assign n13491 = pi74  & n9701;
  assign n13492 = pi76  & n9308;
  assign n13493 = pi75  & n9303;
  assign n13494 = ~n13492 & ~n13493;
  assign n13495 = ~n13491 & n13494;
  assign n13496 = ~n13490 & n13495;
  assign n13497 = pi53  & ~n13496;
  assign n13498 = pi53  & ~n13497;
  assign n13499 = ~n13496 & ~n13497;
  assign n13500 = ~n13498 & ~n13499;
  assign n13501 = n13489 & n13500;
  assign n13502 = ~n13489 & ~n13500;
  assign n13503 = ~n13501 & ~n13502;
  assign n13504 = ~n13430 & n13503;
  assign n13505 = n13430 & ~n13503;
  assign n13506 = ~n13504 & ~n13505;
  assign n13507 = n1122 & n8334;
  assign n13508 = pi77  & n8685;
  assign n13509 = pi79  & n8332;
  assign n13510 = pi78  & n8327;
  assign n13511 = ~n13509 & ~n13510;
  assign n13512 = ~n13508 & n13511;
  assign n13513 = ~n13507 & n13512;
  assign n13514 = pi50  & ~n13513;
  assign n13515 = pi50  & ~n13514;
  assign n13516 = ~n13513 & ~n13514;
  assign n13517 = ~n13515 & ~n13516;
  assign n13518 = n13506 & ~n13517;
  assign n13519 = n13506 & ~n13518;
  assign n13520 = ~n13517 & ~n13518;
  assign n13521 = ~n13519 & ~n13520;
  assign n13522 = ~n13071 & ~n13075;
  assign n13523 = n13521 & n13522;
  assign n13524 = ~n13521 & ~n13522;
  assign n13525 = ~n13523 & ~n13524;
  assign n13526 = n1554 & n7408;
  assign n13527 = pi80  & n7740;
  assign n13528 = pi82  & n7406;
  assign n13529 = pi81  & n7401;
  assign n13530 = ~n13528 & ~n13529;
  assign n13531 = ~n13527 & n13530;
  assign n13532 = ~n13526 & n13531;
  assign n13533 = pi47  & ~n13532;
  assign n13534 = pi47  & ~n13533;
  assign n13535 = ~n13532 & ~n13533;
  assign n13536 = ~n13534 & ~n13535;
  assign n13537 = ~n13525 & n13536;
  assign n13538 = n13525 & ~n13536;
  assign n13539 = ~n13537 & ~n13538;
  assign n13540 = ~n13429 & n13539;
  assign n13541 = n13429 & ~n13539;
  assign n13542 = ~n13540 & ~n13541;
  assign n13543 = ~n13428 & n13542;
  assign n13544 = n13428 & ~n13542;
  assign n13545 = ~n13543 & ~n13544;
  assign n13546 = ~n13417 & n13545;
  assign n13547 = n13417 & ~n13545;
  assign n13548 = ~n13546 & ~n13547;
  assign n13549 = n2446 & n5739;
  assign n13550 = pi86  & n6030;
  assign n13551 = pi88  & n5737;
  assign n13552 = pi87  & n5732;
  assign n13553 = ~n13551 & ~n13552;
  assign n13554 = ~n13550 & n13553;
  assign n13555 = ~n13549 & n13554;
  assign n13556 = pi41  & ~n13555;
  assign n13557 = pi41  & ~n13556;
  assign n13558 = ~n13555 & ~n13556;
  assign n13559 = ~n13557 & ~n13558;
  assign n13560 = n13548 & ~n13559;
  assign n13561 = n13548 & ~n13560;
  assign n13562 = ~n13559 & ~n13560;
  assign n13563 = ~n13561 & ~n13562;
  assign n13564 = ~n13115 & ~n13119;
  assign n13565 = n13563 & n13564;
  assign n13566 = ~n13563 & ~n13564;
  assign n13567 = ~n13565 & ~n13566;
  assign n13568 = n2978 & n5008;
  assign n13569 = pi89  & n5241;
  assign n13570 = pi91  & n5006;
  assign n13571 = pi90  & n5001;
  assign n13572 = ~n13570 & ~n13571;
  assign n13573 = ~n13569 & n13572;
  assign n13574 = ~n13568 & n13573;
  assign n13575 = pi38  & ~n13574;
  assign n13576 = pi38  & ~n13575;
  assign n13577 = ~n13574 & ~n13575;
  assign n13578 = ~n13576 & ~n13577;
  assign n13579 = n13567 & ~n13578;
  assign n13580 = n13567 & ~n13579;
  assign n13581 = ~n13578 & ~n13579;
  assign n13582 = ~n13580 & ~n13581;
  assign n13583 = ~n13132 & ~n13138;
  assign n13584 = n13582 & n13583;
  assign n13585 = ~n13582 & ~n13583;
  assign n13586 = ~n13584 & ~n13585;
  assign n13587 = n3565 & n4271;
  assign n13588 = pi92  & n4503;
  assign n13589 = pi94  & n4269;
  assign n13590 = pi93  & n4264;
  assign n13591 = ~n13589 & ~n13590;
  assign n13592 = ~n13588 & n13591;
  assign n13593 = ~n13587 & n13592;
  assign n13594 = pi35  & ~n13593;
  assign n13595 = pi35  & ~n13594;
  assign n13596 = ~n13593 & ~n13594;
  assign n13597 = ~n13595 & ~n13596;
  assign n13598 = ~n13586 & n13597;
  assign n13599 = n13586 & ~n13597;
  assign n13600 = ~n13598 & ~n13599;
  assign n13601 = ~n13151 & ~n13157;
  assign n13602 = n13600 & ~n13601;
  assign n13603 = ~n13600 & n13601;
  assign n13604 = ~n13602 & ~n13603;
  assign n13605 = n3622 & n4211;
  assign n13606 = pi95  & n3814;
  assign n13607 = pi97  & n3620;
  assign n13608 = pi96  & n3615;
  assign n13609 = ~n13607 & ~n13608;
  assign n13610 = ~n13606 & n13609;
  assign n13611 = ~n13605 & n13610;
  assign n13612 = pi32  & ~n13611;
  assign n13613 = pi32  & ~n13612;
  assign n13614 = ~n13611 & ~n13612;
  assign n13615 = ~n13613 & ~n13614;
  assign n13616 = n13604 & ~n13615;
  assign n13617 = n13604 & ~n13616;
  assign n13618 = ~n13615 & ~n13616;
  assign n13619 = ~n13617 & ~n13618;
  assign n13620 = ~n13175 & n13619;
  assign n13621 = n13175 & ~n13619;
  assign n13622 = ~n13620 & ~n13621;
  assign n13623 = n3034 & n4910;
  assign n13624 = pi98  & n3225;
  assign n13625 = pi100  & n3032;
  assign n13626 = pi99  & n3027;
  assign n13627 = ~n13625 & ~n13626;
  assign n13628 = ~n13624 & n13627;
  assign n13629 = ~n13623 & n13628;
  assign n13630 = pi29  & ~n13629;
  assign n13631 = pi29  & ~n13630;
  assign n13632 = ~n13629 & ~n13630;
  assign n13633 = ~n13631 & ~n13632;
  assign n13634 = ~n13622 & ~n13633;
  assign n13635 = n13622 & n13633;
  assign n13636 = ~n13634 & ~n13635;
  assign n13637 = n13415 & ~n13636;
  assign n13638 = ~n13415 & n13636;
  assign n13639 = ~n13637 & ~n13638;
  assign n13640 = n2523 & n5664;
  assign n13641 = pi101  & n2667;
  assign n13642 = pi103  & n2521;
  assign n13643 = pi102  & n2516;
  assign n13644 = ~n13642 & ~n13643;
  assign n13645 = ~n13641 & n13644;
  assign n13646 = ~n13640 & n13645;
  assign n13647 = pi26  & ~n13646;
  assign n13648 = pi26  & ~n13647;
  assign n13649 = ~n13646 & ~n13647;
  assign n13650 = ~n13648 & ~n13649;
  assign n13651 = ~n13639 & n13650;
  assign n13652 = n13639 & ~n13650;
  assign n13653 = ~n13651 & ~n13652;
  assign n13654 = ~n13414 & n13653;
  assign n13655 = n13414 & ~n13653;
  assign n13656 = ~n13654 & ~n13655;
  assign n13657 = ~n13413 & n13656;
  assign n13658 = ~n13413 & ~n13657;
  assign n13659 = n13656 & ~n13657;
  assign n13660 = ~n13658 & ~n13659;
  assign n13661 = ~n13232 & ~n13660;
  assign n13662 = n13232 & n13660;
  assign n13663 = ~n13661 & ~n13662;
  assign n13664 = ~n13402 & n13663;
  assign n13665 = ~n13402 & ~n13664;
  assign n13666 = n13663 & ~n13664;
  assign n13667 = ~n13665 & ~n13666;
  assign n13668 = ~n13391 & ~n13667;
  assign n13669 = n13391 & n13667;
  assign n13670 = ~n13668 & ~n13669;
  assign n13671 = ~n13389 & n13670;
  assign n13672 = ~n13389 & ~n13671;
  assign n13673 = n13670 & ~n13671;
  assign n13674 = ~n13672 & ~n13673;
  assign n13675 = ~n13378 & ~n13674;
  assign n13676 = n13378 & n13674;
  assign n13677 = ~n13675 & ~n13676;
  assign n13678 = ~n13377 & n13677;
  assign n13679 = n13377 & ~n13677;
  assign n13680 = ~n13678 & ~n13679;
  assign n13681 = ~n13366 & n13680;
  assign n13682 = n13366 & ~n13680;
  assign n13683 = ~n13681 & ~n13682;
  assign n13684 = n687 & n9984;
  assign n13685 = pi116  & n763;
  assign n13686 = pi118  & n685;
  assign n13687 = pi117  & n680;
  assign n13688 = ~n13686 & ~n13687;
  assign n13689 = ~n13685 & n13688;
  assign n13690 = ~n13684 & n13689;
  assign n13691 = pi11  & ~n13690;
  assign n13692 = pi11  & ~n13691;
  assign n13693 = ~n13690 & ~n13691;
  assign n13694 = ~n13692 & ~n13693;
  assign n13695 = n13683 & ~n13694;
  assign n13696 = n13683 & ~n13695;
  assign n13697 = ~n13694 & ~n13695;
  assign n13698 = ~n13696 & ~n13697;
  assign n13699 = ~n13299 & ~n13302;
  assign n13700 = n13698 & n13699;
  assign n13701 = ~n13698 & ~n13699;
  assign n13702 = ~n13700 & ~n13701;
  assign n13703 = n498 & n11389;
  assign n13704 = pi119  & n537;
  assign n13705 = pi121  & n496;
  assign n13706 = pi120  & n491;
  assign n13707 = ~n13705 & ~n13706;
  assign n13708 = ~n13704 & n13707;
  assign n13709 = ~n13703 & n13708;
  assign n13710 = pi8  & ~n13709;
  assign n13711 = pi8  & ~n13710;
  assign n13712 = ~n13709 & ~n13710;
  assign n13713 = ~n13711 & ~n13712;
  assign n13714 = n13702 & ~n13713;
  assign n13715 = n13702 & ~n13714;
  assign n13716 = ~n13713 & ~n13714;
  assign n13717 = ~n13715 & ~n13716;
  assign n13718 = n342 & n12189;
  assign n13719 = pi122  & n380;
  assign n13720 = pi124  & n340;
  assign n13721 = pi123  & n335;
  assign n13722 = ~n13720 & ~n13721;
  assign n13723 = ~n13719 & n13722;
  assign n13724 = ~n13718 & n13723;
  assign n13725 = pi5  & ~n13724;
  assign n13726 = pi5  & ~n13725;
  assign n13727 = ~n13724 & ~n13725;
  assign n13728 = ~n13726 & ~n13727;
  assign n13729 = ~n13717 & n13728;
  assign n13730 = n13717 & ~n13728;
  assign n13731 = ~n13729 & ~n13730;
  assign n13732 = ~n13317 & ~n13330;
  assign n13733 = n13731 & n13732;
  assign n13734 = ~n13731 & ~n13732;
  assign n13735 = ~n13733 & ~n13734;
  assign n13736 = ~n13340 & ~n13342;
  assign n13737 = pi126  & ~pi127 ;
  assign n13738 = ~pi126  & pi127 ;
  assign n13739 = ~n13737 & ~n13738;
  assign n13740 = ~n13736 & ~n13739;
  assign n13741 = n13736 & n13739;
  assign n13742 = ~n13740 & ~n13741;
  assign n13743 = n262 & n13742;
  assign n13744 = pi125  & n288;
  assign n13745 = pi127  & n267;
  assign n13746 = pi126  & n269;
  assign n13747 = ~n13745 & ~n13746;
  assign n13748 = ~n13744 & n13747;
  assign n13749 = ~n13743 & n13748;
  assign n13750 = pi2  & ~n13749;
  assign n13751 = pi2  & ~n13750;
  assign n13752 = ~n13749 & ~n13750;
  assign n13753 = ~n13751 & ~n13752;
  assign n13754 = n13735 & ~n13753;
  assign n13755 = n13735 & ~n13754;
  assign n13756 = ~n13753 & ~n13754;
  assign n13757 = ~n13755 & ~n13756;
  assign n13758 = ~n13336 & ~n13357;
  assign n13759 = ~n13757 & ~n13758;
  assign n13760 = ~n13757 & ~n13759;
  assign n13761 = ~n13758 & ~n13759;
  assign n13762 = ~n13760 & ~n13761;
  assign n13763 = ~n13359 & ~n13362;
  assign n13764 = ~n13762 & ~n13763;
  assign n13765 = n13762 & n13763;
  assign po63  = ~n13764 & ~n13765;
  assign n13767 = ~n13759 & ~n13764;
  assign n13768 = ~n13734 & ~n13754;
  assign n13769 = ~pi126  & ~n13740;
  assign n13770 = pi127  & ~n13769;
  assign n13771 = pi127  & ~n13770;
  assign n13772 = ~n13736 & n13737;
  assign n13773 = ~n13771 & ~n13772;
  assign n13774 = n262 & ~n13773;
  assign n13775 = pi126  & n288;
  assign n13776 = pi127  & n269;
  assign n13777 = ~n13775 & ~n13776;
  assign n13778 = ~n13774 & n13777;
  assign n13779 = pi2  & ~n13778;
  assign n13780 = pi2  & ~n13779;
  assign n13781 = ~n13778 & ~n13779;
  assign n13782 = ~n13780 & ~n13781;
  assign n13783 = ~n13717 & ~n13728;
  assign n13784 = ~n13714 & ~n13783;
  assign n13785 = ~n13695 & ~n13701;
  assign n13786 = n687 & n10667;
  assign n13787 = pi117  & n763;
  assign n13788 = pi119  & n685;
  assign n13789 = pi118  & n680;
  assign n13790 = ~n13788 & ~n13789;
  assign n13791 = ~n13787 & n13790;
  assign n13792 = ~n13786 & n13791;
  assign n13793 = pi11  & ~n13792;
  assign n13794 = pi11  & ~n13793;
  assign n13795 = ~n13792 & ~n13793;
  assign n13796 = ~n13794 & ~n13795;
  assign n13797 = ~n13678 & ~n13681;
  assign n13798 = n938 & n9614;
  assign n13799 = pi114  & n1052;
  assign n13800 = pi116  & n936;
  assign n13801 = pi115  & n931;
  assign n13802 = ~n13800 & ~n13801;
  assign n13803 = ~n13799 & n13802;
  assign n13804 = ~n13798 & n13803;
  assign n13805 = pi14  & ~n13804;
  assign n13806 = pi14  & ~n13805;
  assign n13807 = ~n13804 & ~n13805;
  assign n13808 = ~n13806 & ~n13807;
  assign n13809 = ~n13671 & ~n13675;
  assign n13810 = n1297 & n8612;
  assign n13811 = pi111  & n1366;
  assign n13812 = pi113  & n1295;
  assign n13813 = pi112  & n1290;
  assign n13814 = ~n13812 & ~n13813;
  assign n13815 = ~n13811 & n13814;
  assign n13816 = ~n13810 & n13815;
  assign n13817 = pi17  & ~n13816;
  assign n13818 = pi17  & ~n13817;
  assign n13819 = ~n13816 & ~n13817;
  assign n13820 = ~n13818 & ~n13819;
  assign n13821 = ~n13664 & ~n13668;
  assign n13822 = n1611 & n7665;
  assign n13823 = pi108  & n1745;
  assign n13824 = pi110  & n1609;
  assign n13825 = pi109  & n1604;
  assign n13826 = ~n13824 & ~n13825;
  assign n13827 = ~n13823 & n13826;
  assign n13828 = ~n13822 & n13827;
  assign n13829 = pi20  & ~n13828;
  assign n13830 = pi20  & ~n13829;
  assign n13831 = ~n13828 & ~n13829;
  assign n13832 = ~n13830 & ~n13831;
  assign n13833 = ~n13657 & ~n13661;
  assign n13834 = ~n13467 & ~n13469;
  assign n13835 = pi63  & n13434;
  assign n13836 = pi64  & n13835;
  assign n13837 = pi65  & ~n13434;
  assign n13838 = ~n13836 & ~n13837;
  assign n13839 = n359 & n12627;
  assign n13840 = pi66  & n13004;
  assign n13841 = pi68  & n12625;
  assign n13842 = pi67  & n12620;
  assign n13843 = ~n13841 & ~n13842;
  assign n13844 = ~n13840 & n13843;
  assign n13845 = ~n13839 & n13844;
  assign n13846 = pi62  & ~n13845;
  assign n13847 = pi62  & ~n13846;
  assign n13848 = ~n13845 & ~n13846;
  assign n13849 = ~n13847 & ~n13848;
  assign n13850 = ~n13838 & ~n13849;
  assign n13851 = ~n13838 & ~n13850;
  assign n13852 = ~n13849 & ~n13850;
  assign n13853 = ~n13851 & ~n13852;
  assign n13854 = ~n13436 & ~n13451;
  assign n13855 = n13853 & n13854;
  assign n13856 = ~n13853 & ~n13854;
  assign n13857 = ~n13855 & ~n13856;
  assign n13858 = n475 & n11488;
  assign n13859 = pi69  & n11847;
  assign n13860 = pi71  & n11486;
  assign n13861 = pi70  & n11481;
  assign n13862 = ~n13860 & ~n13861;
  assign n13863 = ~n13859 & n13862;
  assign n13864 = ~n13858 & n13863;
  assign n13865 = pi59  & ~n13864;
  assign n13866 = pi59  & ~n13865;
  assign n13867 = ~n13864 & ~n13865;
  assign n13868 = ~n13866 & ~n13867;
  assign n13869 = ~n13857 & n13868;
  assign n13870 = n13857 & ~n13868;
  assign n13871 = ~n13869 & ~n13870;
  assign n13872 = ~n13834 & n13871;
  assign n13873 = n13834 & ~n13871;
  assign n13874 = ~n13872 & ~n13873;
  assign n13875 = n729 & n10394;
  assign n13876 = pi72  & n10744;
  assign n13877 = pi74  & n10392;
  assign n13878 = pi73  & n10387;
  assign n13879 = ~n13877 & ~n13878;
  assign n13880 = ~n13876 & n13879;
  assign n13881 = ~n13875 & n13880;
  assign n13882 = pi56  & ~n13881;
  assign n13883 = pi56  & ~n13882;
  assign n13884 = ~n13881 & ~n13882;
  assign n13885 = ~n13883 & ~n13884;
  assign n13886 = n13874 & ~n13885;
  assign n13887 = n13874 & ~n13886;
  assign n13888 = ~n13885 & ~n13886;
  assign n13889 = ~n13887 & ~n13888;
  assign n13890 = ~n13431 & ~n13486;
  assign n13891 = ~n13483 & ~n13890;
  assign n13892 = n13889 & n13891;
  assign n13893 = ~n13889 & ~n13891;
  assign n13894 = ~n13892 & ~n13893;
  assign n13895 = n999 & n9310;
  assign n13896 = pi75  & n9701;
  assign n13897 = pi77  & n9308;
  assign n13898 = pi76  & n9303;
  assign n13899 = ~n13897 & ~n13898;
  assign n13900 = ~n13896 & n13899;
  assign n13901 = ~n13895 & n13900;
  assign n13902 = pi53  & ~n13901;
  assign n13903 = pi53  & ~n13902;
  assign n13904 = ~n13901 & ~n13902;
  assign n13905 = ~n13903 & ~n13904;
  assign n13906 = ~n13894 & n13905;
  assign n13907 = n13894 & ~n13905;
  assign n13908 = ~n13906 & ~n13907;
  assign n13909 = ~n13502 & ~n13504;
  assign n13910 = n13908 & ~n13909;
  assign n13911 = ~n13908 & n13909;
  assign n13912 = ~n13910 & ~n13911;
  assign n13913 = n1225 & n8334;
  assign n13914 = pi78  & n8685;
  assign n13915 = pi80  & n8332;
  assign n13916 = pi79  & n8327;
  assign n13917 = ~n13915 & ~n13916;
  assign n13918 = ~n13914 & n13917;
  assign n13919 = ~n13913 & n13918;
  assign n13920 = pi50  & ~n13919;
  assign n13921 = pi50  & ~n13920;
  assign n13922 = ~n13919 & ~n13920;
  assign n13923 = ~n13921 & ~n13922;
  assign n13924 = n13912 & ~n13923;
  assign n13925 = n13912 & ~n13924;
  assign n13926 = ~n13923 & ~n13924;
  assign n13927 = ~n13925 & ~n13926;
  assign n13928 = ~n13518 & ~n13524;
  assign n13929 = n13927 & n13928;
  assign n13930 = ~n13927 & ~n13928;
  assign n13931 = ~n13929 & ~n13930;
  assign n13932 = n1696 & n7408;
  assign n13933 = pi81  & n7740;
  assign n13934 = pi83  & n7406;
  assign n13935 = pi82  & n7401;
  assign n13936 = ~n13934 & ~n13935;
  assign n13937 = ~n13933 & n13936;
  assign n13938 = ~n13932 & n13937;
  assign n13939 = pi47  & ~n13938;
  assign n13940 = pi47  & ~n13939;
  assign n13941 = ~n13938 & ~n13939;
  assign n13942 = ~n13940 & ~n13941;
  assign n13943 = ~n13931 & n13942;
  assign n13944 = n13931 & ~n13942;
  assign n13945 = ~n13943 & ~n13944;
  assign n13946 = ~n13538 & ~n13540;
  assign n13947 = n13945 & ~n13946;
  assign n13948 = ~n13945 & n13946;
  assign n13949 = ~n13947 & ~n13948;
  assign n13950 = n2133 & n6539;
  assign n13951 = pi84  & n6873;
  assign n13952 = pi86  & n6537;
  assign n13953 = pi85  & n6532;
  assign n13954 = ~n13952 & ~n13953;
  assign n13955 = ~n13951 & n13954;
  assign n13956 = ~n13950 & n13955;
  assign n13957 = pi44  & ~n13956;
  assign n13958 = pi44  & ~n13957;
  assign n13959 = ~n13956 & ~n13957;
  assign n13960 = ~n13958 & ~n13959;
  assign n13961 = n13949 & ~n13960;
  assign n13962 = n13949 & ~n13961;
  assign n13963 = ~n13960 & ~n13961;
  assign n13964 = ~n13962 & ~n13963;
  assign n13965 = ~n13543 & ~n13546;
  assign n13966 = n13964 & n13965;
  assign n13967 = ~n13964 & ~n13965;
  assign n13968 = ~n13966 & ~n13967;
  assign n13969 = n2473 & n5739;
  assign n13970 = pi87  & n6030;
  assign n13971 = pi89  & n5737;
  assign n13972 = pi88  & n5732;
  assign n13973 = ~n13971 & ~n13972;
  assign n13974 = ~n13970 & n13973;
  assign n13975 = ~n13969 & n13974;
  assign n13976 = pi41  & ~n13975;
  assign n13977 = pi41  & ~n13976;
  assign n13978 = ~n13975 & ~n13976;
  assign n13979 = ~n13977 & ~n13978;
  assign n13980 = n13968 & ~n13979;
  assign n13981 = n13968 & ~n13980;
  assign n13982 = ~n13979 & ~n13980;
  assign n13983 = ~n13981 & ~n13982;
  assign n13984 = ~n13560 & ~n13566;
  assign n13985 = n13983 & n13984;
  assign n13986 = ~n13983 & ~n13984;
  assign n13987 = ~n13985 & ~n13986;
  assign n13988 = n3177 & n5008;
  assign n13989 = pi90  & n5241;
  assign n13990 = pi92  & n5006;
  assign n13991 = pi91  & n5001;
  assign n13992 = ~n13990 & ~n13991;
  assign n13993 = ~n13989 & n13992;
  assign n13994 = ~n13988 & n13993;
  assign n13995 = pi38  & ~n13994;
  assign n13996 = pi38  & ~n13995;
  assign n13997 = ~n13994 & ~n13995;
  assign n13998 = ~n13996 & ~n13997;
  assign n13999 = n13987 & ~n13998;
  assign n14000 = n13987 & ~n13999;
  assign n14001 = ~n13998 & ~n13999;
  assign n14002 = ~n14000 & ~n14001;
  assign n14003 = ~n13579 & ~n13585;
  assign n14004 = n14002 & n14003;
  assign n14005 = ~n14002 & ~n14003;
  assign n14006 = ~n14004 & ~n14005;
  assign n14007 = n3784 & n4271;
  assign n14008 = pi93  & n4503;
  assign n14009 = pi95  & n4269;
  assign n14010 = pi94  & n4264;
  assign n14011 = ~n14009 & ~n14010;
  assign n14012 = ~n14008 & n14011;
  assign n14013 = ~n14007 & n14012;
  assign n14014 = pi35  & ~n14013;
  assign n14015 = pi35  & ~n14014;
  assign n14016 = ~n14013 & ~n14014;
  assign n14017 = ~n14015 & ~n14016;
  assign n14018 = ~n14006 & n14017;
  assign n14019 = n14006 & ~n14017;
  assign n14020 = ~n14018 & ~n14019;
  assign n14021 = ~n13599 & ~n13602;
  assign n14022 = n14020 & ~n14021;
  assign n14023 = ~n14020 & n14021;
  assign n14024 = ~n14022 & ~n14023;
  assign n14025 = n3622 & n4454;
  assign n14026 = pi96  & n3814;
  assign n14027 = pi98  & n3620;
  assign n14028 = pi97  & n3615;
  assign n14029 = ~n14027 & ~n14028;
  assign n14030 = ~n14026 & n14029;
  assign n14031 = ~n14025 & n14030;
  assign n14032 = pi32  & ~n14031;
  assign n14033 = pi32  & ~n14032;
  assign n14034 = ~n14031 & ~n14032;
  assign n14035 = ~n14033 & ~n14034;
  assign n14036 = n14024 & ~n14035;
  assign n14037 = n14024 & ~n14036;
  assign n14038 = ~n14035 & ~n14036;
  assign n14039 = ~n14037 & ~n14038;
  assign n14040 = ~n13175 & ~n13619;
  assign n14041 = ~n13616 & ~n14040;
  assign n14042 = n14039 & n14041;
  assign n14043 = ~n14039 & ~n14041;
  assign n14044 = ~n14042 & ~n14043;
  assign n14045 = n3034 & n5169;
  assign n14046 = pi99  & n3225;
  assign n14047 = pi101  & n3032;
  assign n14048 = pi100  & n3027;
  assign n14049 = ~n14047 & ~n14048;
  assign n14050 = ~n14046 & n14049;
  assign n14051 = ~n14045 & n14050;
  assign n14052 = pi29  & ~n14051;
  assign n14053 = pi29  & ~n14052;
  assign n14054 = ~n14051 & ~n14052;
  assign n14055 = ~n14053 & ~n14054;
  assign n14056 = n14044 & ~n14055;
  assign n14057 = n14044 & ~n14056;
  assign n14058 = ~n14055 & ~n14056;
  assign n14059 = ~n14057 & ~n14058;
  assign n14060 = ~n13634 & ~n13638;
  assign n14061 = n14059 & n14060;
  assign n14062 = ~n14059 & ~n14060;
  assign n14063 = ~n14061 & ~n14062;
  assign n14064 = n2523 & n5943;
  assign n14065 = pi102  & n2667;
  assign n14066 = pi104  & n2521;
  assign n14067 = pi103  & n2516;
  assign n14068 = ~n14066 & ~n14067;
  assign n14069 = ~n14065 & n14068;
  assign n14070 = ~n14064 & n14069;
  assign n14071 = pi26  & ~n14070;
  assign n14072 = pi26  & ~n14071;
  assign n14073 = ~n14070 & ~n14071;
  assign n14074 = ~n14072 & ~n14073;
  assign n14075 = n14063 & ~n14074;
  assign n14076 = n14063 & ~n14075;
  assign n14077 = ~n14074 & ~n14075;
  assign n14078 = ~n14076 & ~n14077;
  assign n14079 = ~n13652 & ~n13654;
  assign n14080 = ~n14078 & ~n14079;
  assign n14081 = ~n14078 & ~n14080;
  assign n14082 = ~n14079 & ~n14080;
  assign n14083 = ~n14081 & ~n14082;
  assign n14084 = n2043 & n6775;
  assign n14085 = pi105  & n2180;
  assign n14086 = pi107  & n2041;
  assign n14087 = pi106  & n2036;
  assign n14088 = ~n14086 & ~n14087;
  assign n14089 = ~n14085 & n14088;
  assign n14090 = ~n14084 & n14089;
  assign n14091 = pi23  & ~n14090;
  assign n14092 = pi23  & ~n14091;
  assign n14093 = ~n14090 & ~n14091;
  assign n14094 = ~n14092 & ~n14093;
  assign n14095 = ~n14083 & n14094;
  assign n14096 = n14083 & ~n14094;
  assign n14097 = ~n14095 & ~n14096;
  assign n14098 = ~n13833 & ~n14097;
  assign n14099 = n13833 & n14097;
  assign n14100 = ~n14098 & ~n14099;
  assign n14101 = ~n13832 & n14100;
  assign n14102 = ~n13832 & ~n14101;
  assign n14103 = n14100 & ~n14101;
  assign n14104 = ~n14102 & ~n14103;
  assign n14105 = ~n13821 & ~n14104;
  assign n14106 = n13821 & n14104;
  assign n14107 = ~n14105 & ~n14106;
  assign n14108 = ~n13820 & n14107;
  assign n14109 = ~n13820 & ~n14108;
  assign n14110 = n14107 & ~n14108;
  assign n14111 = ~n14109 & ~n14110;
  assign n14112 = ~n13809 & ~n14111;
  assign n14113 = n13809 & n14111;
  assign n14114 = ~n14112 & ~n14113;
  assign n14115 = ~n13808 & n14114;
  assign n14116 = n13808 & ~n14114;
  assign n14117 = ~n14115 & ~n14116;
  assign n14118 = ~n13797 & n14117;
  assign n14119 = n13797 & ~n14117;
  assign n14120 = ~n14118 & ~n14119;
  assign n14121 = ~n13796 & n14120;
  assign n14122 = n13796 & ~n14120;
  assign n14123 = ~n14121 & ~n14122;
  assign n14124 = ~n13785 & n14123;
  assign n14125 = n13785 & ~n14123;
  assign n14126 = ~n14124 & ~n14125;
  assign n14127 = n498 & n11778;
  assign n14128 = pi120  & n537;
  assign n14129 = pi122  & n496;
  assign n14130 = pi121  & n491;
  assign n14131 = ~n14129 & ~n14130;
  assign n14132 = ~n14128 & n14131;
  assign n14133 = ~n14127 & n14132;
  assign n14134 = pi8  & ~n14133;
  assign n14135 = pi8  & ~n14134;
  assign n14136 = ~n14133 & ~n14134;
  assign n14137 = ~n14135 & ~n14136;
  assign n14138 = n14126 & ~n14137;
  assign n14139 = n14126 & ~n14138;
  assign n14140 = ~n14137 & ~n14138;
  assign n14141 = ~n14139 & ~n14140;
  assign n14142 = n342 & n12943;
  assign n14143 = pi123  & n380;
  assign n14144 = pi125  & n340;
  assign n14145 = pi124  & n335;
  assign n14146 = ~n14144 & ~n14145;
  assign n14147 = ~n14143 & n14146;
  assign n14148 = ~n14142 & n14147;
  assign n14149 = pi5  & ~n14148;
  assign n14150 = pi5  & ~n14149;
  assign n14151 = ~n14148 & ~n14149;
  assign n14152 = ~n14150 & ~n14151;
  assign n14153 = ~n14141 & n14152;
  assign n14154 = n14141 & ~n14152;
  assign n14155 = ~n14153 & ~n14154;
  assign n14156 = ~n13784 & ~n14155;
  assign n14157 = n13784 & n14155;
  assign n14158 = ~n14156 & ~n14157;
  assign n14159 = ~n13782 & n14158;
  assign n14160 = n13782 & ~n14158;
  assign n14161 = ~n14159 & ~n14160;
  assign n14162 = ~n13768 & n14161;
  assign n14163 = n13768 & ~n14161;
  assign n14164 = ~n14162 & ~n14163;
  assign n14165 = ~n13767 & n14164;
  assign n14166 = n13767 & ~n14164;
  assign po64  = ~n14165 & ~n14166;
  assign n14168 = ~n14108 & ~n14112;
  assign n14169 = ~n14101 & ~n14105;
  assign n14170 = n1611 & n7970;
  assign n14171 = pi109  & n1745;
  assign n14172 = pi111  & n1609;
  assign n14173 = pi110  & n1604;
  assign n14174 = ~n14172 & ~n14173;
  assign n14175 = ~n14171 & n14174;
  assign n14176 = ~n14170 & n14175;
  assign n14177 = pi20  & ~n14176;
  assign n14178 = pi20  & ~n14177;
  assign n14179 = ~n14176 & ~n14177;
  assign n14180 = ~n14178 & ~n14179;
  assign n14181 = ~n14075 & ~n14080;
  assign n14182 = ~n14019 & ~n14022;
  assign n14183 = ~n13961 & ~n13967;
  assign n14184 = ~n13944 & ~n13947;
  assign n14185 = ~n13924 & ~n13930;
  assign n14186 = ~n13907 & ~n13910;
  assign n14187 = ~n13886 & ~n13893;
  assign n14188 = ~n13870 & ~n13872;
  assign n14189 = pi65  & n13835;
  assign n14190 = pi66  & ~n13434;
  assign n14191 = ~n14189 & ~n14190;
  assign n14192 = n401 & n12627;
  assign n14193 = pi67  & n13004;
  assign n14194 = pi69  & n12625;
  assign n14195 = pi68  & n12620;
  assign n14196 = ~n14194 & ~n14195;
  assign n14197 = ~n14193 & n14196;
  assign n14198 = ~n14192 & n14197;
  assign n14199 = pi62  & ~n14198;
  assign n14200 = pi62  & ~n14199;
  assign n14201 = ~n14198 & ~n14199;
  assign n14202 = ~n14200 & ~n14201;
  assign n14203 = ~n14191 & ~n14202;
  assign n14204 = ~n14191 & ~n14203;
  assign n14205 = ~n14202 & ~n14203;
  assign n14206 = ~n14204 & ~n14205;
  assign n14207 = ~n13850 & ~n13856;
  assign n14208 = n14206 & n14207;
  assign n14209 = ~n14206 & ~n14207;
  assign n14210 = ~n14208 & ~n14209;
  assign n14211 = n576 & n11488;
  assign n14212 = pi70  & n11847;
  assign n14213 = pi72  & n11486;
  assign n14214 = pi71  & n11481;
  assign n14215 = ~n14213 & ~n14214;
  assign n14216 = ~n14212 & n14215;
  assign n14217 = ~n14211 & n14216;
  assign n14218 = pi59  & ~n14217;
  assign n14219 = pi59  & ~n14218;
  assign n14220 = ~n14217 & ~n14218;
  assign n14221 = ~n14219 & ~n14220;
  assign n14222 = n14210 & ~n14221;
  assign n14223 = ~n14210 & n14221;
  assign n14224 = ~n14222 & ~n14223;
  assign n14225 = ~n14188 & n14224;
  assign n14226 = ~n14188 & ~n14225;
  assign n14227 = ~n14222 & ~n14225;
  assign n14228 = ~n14223 & n14227;
  assign n14229 = ~n14226 & ~n14228;
  assign n14230 = n809 & n10394;
  assign n14231 = pi73  & n10744;
  assign n14232 = pi75  & n10392;
  assign n14233 = pi74  & n10387;
  assign n14234 = ~n14232 & ~n14233;
  assign n14235 = ~n14231 & n14234;
  assign n14236 = ~n14230 & n14235;
  assign n14237 = pi56  & ~n14236;
  assign n14238 = pi56  & ~n14237;
  assign n14239 = ~n14236 & ~n14237;
  assign n14240 = ~n14238 & ~n14239;
  assign n14241 = n14229 & n14240;
  assign n14242 = ~n14229 & ~n14240;
  assign n14243 = ~n14241 & ~n14242;
  assign n14244 = ~n14187 & n14243;
  assign n14245 = n14187 & ~n14243;
  assign n14246 = ~n14244 & ~n14245;
  assign n14247 = n1025 & n9310;
  assign n14248 = pi76  & n9701;
  assign n14249 = pi78  & n9308;
  assign n14250 = pi77  & n9303;
  assign n14251 = ~n14249 & ~n14250;
  assign n14252 = ~n14248 & n14251;
  assign n14253 = ~n14247 & n14252;
  assign n14254 = pi53  & ~n14253;
  assign n14255 = pi53  & ~n14254;
  assign n14256 = ~n14253 & ~n14254;
  assign n14257 = ~n14255 & ~n14256;
  assign n14258 = n14246 & ~n14257;
  assign n14259 = n14246 & ~n14258;
  assign n14260 = ~n14257 & ~n14258;
  assign n14261 = ~n14259 & ~n14260;
  assign n14262 = ~n14186 & n14261;
  assign n14263 = n14186 & ~n14261;
  assign n14264 = ~n14262 & ~n14263;
  assign n14265 = n1434 & n8334;
  assign n14266 = pi79  & n8685;
  assign n14267 = pi81  & n8332;
  assign n14268 = pi80  & n8327;
  assign n14269 = ~n14267 & ~n14268;
  assign n14270 = ~n14266 & n14269;
  assign n14271 = ~n14265 & n14270;
  assign n14272 = pi50  & ~n14271;
  assign n14273 = pi50  & ~n14272;
  assign n14274 = ~n14271 & ~n14272;
  assign n14275 = ~n14273 & ~n14274;
  assign n14276 = ~n14264 & ~n14275;
  assign n14277 = n14264 & n14275;
  assign n14278 = ~n14276 & ~n14277;
  assign n14279 = n14185 & ~n14278;
  assign n14280 = ~n14185 & n14278;
  assign n14281 = ~n14279 & ~n14280;
  assign n14282 = n1834 & n7408;
  assign n14283 = pi82  & n7740;
  assign n14284 = pi84  & n7406;
  assign n14285 = pi83  & n7401;
  assign n14286 = ~n14284 & ~n14285;
  assign n14287 = ~n14283 & n14286;
  assign n14288 = ~n14282 & n14287;
  assign n14289 = pi47  & ~n14288;
  assign n14290 = pi47  & ~n14289;
  assign n14291 = ~n14288 & ~n14289;
  assign n14292 = ~n14290 & ~n14291;
  assign n14293 = n14281 & ~n14292;
  assign n14294 = n14281 & ~n14293;
  assign n14295 = ~n14292 & ~n14293;
  assign n14296 = ~n14294 & ~n14295;
  assign n14297 = ~n14184 & n14296;
  assign n14298 = n14184 & ~n14296;
  assign n14299 = ~n14297 & ~n14298;
  assign n14300 = n2288 & n6539;
  assign n14301 = pi85  & n6873;
  assign n14302 = pi87  & n6537;
  assign n14303 = pi86  & n6532;
  assign n14304 = ~n14302 & ~n14303;
  assign n14305 = ~n14301 & n14304;
  assign n14306 = ~n14300 & n14305;
  assign n14307 = pi44  & ~n14306;
  assign n14308 = pi44  & ~n14307;
  assign n14309 = ~n14306 & ~n14307;
  assign n14310 = ~n14308 & ~n14309;
  assign n14311 = ~n14299 & ~n14310;
  assign n14312 = n14299 & n14310;
  assign n14313 = ~n14311 & ~n14312;
  assign n14314 = n14183 & ~n14313;
  assign n14315 = ~n14183 & n14313;
  assign n14316 = ~n14314 & ~n14315;
  assign n14317 = n2801 & n5739;
  assign n14318 = pi88  & n6030;
  assign n14319 = pi90  & n5737;
  assign n14320 = pi89  & n5732;
  assign n14321 = ~n14319 & ~n14320;
  assign n14322 = ~n14318 & n14321;
  assign n14323 = ~n14317 & n14322;
  assign n14324 = pi41  & ~n14323;
  assign n14325 = pi41  & ~n14324;
  assign n14326 = ~n14323 & ~n14324;
  assign n14327 = ~n14325 & ~n14326;
  assign n14328 = n14316 & ~n14327;
  assign n14329 = n14316 & ~n14328;
  assign n14330 = ~n14327 & ~n14328;
  assign n14331 = ~n14329 & ~n14330;
  assign n14332 = ~n13980 & ~n13986;
  assign n14333 = n14331 & n14332;
  assign n14334 = ~n14331 & ~n14332;
  assign n14335 = ~n14333 & ~n14334;
  assign n14336 = n3371 & n5008;
  assign n14337 = pi91  & n5241;
  assign n14338 = pi93  & n5006;
  assign n14339 = pi92  & n5001;
  assign n14340 = ~n14338 & ~n14339;
  assign n14341 = ~n14337 & n14340;
  assign n14342 = ~n14336 & n14341;
  assign n14343 = pi38  & ~n14342;
  assign n14344 = pi38  & ~n14343;
  assign n14345 = ~n14342 & ~n14343;
  assign n14346 = ~n14344 & ~n14345;
  assign n14347 = n14335 & ~n14346;
  assign n14348 = n14335 & ~n14347;
  assign n14349 = ~n14346 & ~n14347;
  assign n14350 = ~n14348 & ~n14349;
  assign n14351 = ~n13999 & ~n14005;
  assign n14352 = n14350 & n14351;
  assign n14353 = ~n14350 & ~n14351;
  assign n14354 = ~n14352 & ~n14353;
  assign n14355 = n4001 & n4271;
  assign n14356 = pi94  & n4503;
  assign n14357 = pi96  & n4269;
  assign n14358 = pi95  & n4264;
  assign n14359 = ~n14357 & ~n14358;
  assign n14360 = ~n14356 & n14359;
  assign n14361 = ~n14355 & n14360;
  assign n14362 = pi35  & ~n14361;
  assign n14363 = pi35  & ~n14362;
  assign n14364 = ~n14361 & ~n14362;
  assign n14365 = ~n14363 & ~n14364;
  assign n14366 = n14354 & ~n14365;
  assign n14367 = ~n14354 & n14365;
  assign n14368 = ~n14366 & ~n14367;
  assign n14369 = ~n14182 & n14368;
  assign n14370 = ~n14182 & ~n14369;
  assign n14371 = ~n14366 & ~n14369;
  assign n14372 = ~n14367 & n14371;
  assign n14373 = ~n14370 & ~n14372;
  assign n14374 = n3622 & n4684;
  assign n14375 = pi97  & n3814;
  assign n14376 = pi99  & n3620;
  assign n14377 = pi98  & n3615;
  assign n14378 = ~n14376 & ~n14377;
  assign n14379 = ~n14375 & n14378;
  assign n14380 = ~n14374 & n14379;
  assign n14381 = pi32  & ~n14380;
  assign n14382 = pi32  & ~n14381;
  assign n14383 = ~n14380 & ~n14381;
  assign n14384 = ~n14382 & ~n14383;
  assign n14385 = ~n14373 & ~n14384;
  assign n14386 = ~n14373 & ~n14385;
  assign n14387 = ~n14384 & ~n14385;
  assign n14388 = ~n14386 & ~n14387;
  assign n14389 = ~n14036 & ~n14043;
  assign n14390 = n14388 & n14389;
  assign n14391 = ~n14388 & ~n14389;
  assign n14392 = ~n14390 & ~n14391;
  assign n14393 = n3034 & n5413;
  assign n14394 = pi100  & n3225;
  assign n14395 = pi102  & n3032;
  assign n14396 = pi101  & n3027;
  assign n14397 = ~n14395 & ~n14396;
  assign n14398 = ~n14394 & n14397;
  assign n14399 = ~n14393 & n14398;
  assign n14400 = pi29  & ~n14399;
  assign n14401 = pi29  & ~n14400;
  assign n14402 = ~n14399 & ~n14400;
  assign n14403 = ~n14401 & ~n14402;
  assign n14404 = n14392 & ~n14403;
  assign n14405 = n14392 & ~n14404;
  assign n14406 = ~n14403 & ~n14404;
  assign n14407 = ~n14405 & ~n14406;
  assign n14408 = ~n14056 & ~n14062;
  assign n14409 = n14407 & n14408;
  assign n14410 = ~n14407 & ~n14408;
  assign n14411 = ~n14409 & ~n14410;
  assign n14412 = n2523 & n6207;
  assign n14413 = pi103  & n2667;
  assign n14414 = pi105  & n2521;
  assign n14415 = pi104  & n2516;
  assign n14416 = ~n14414 & ~n14415;
  assign n14417 = ~n14413 & n14416;
  assign n14418 = ~n14412 & n14417;
  assign n14419 = pi26  & ~n14418;
  assign n14420 = pi26  & ~n14419;
  assign n14421 = ~n14418 & ~n14419;
  assign n14422 = ~n14420 & ~n14421;
  assign n14423 = n14411 & ~n14422;
  assign n14424 = ~n14411 & n14422;
  assign n14425 = ~n14423 & ~n14424;
  assign n14426 = ~n14181 & n14425;
  assign n14427 = ~n14181 & ~n14426;
  assign n14428 = ~n14423 & ~n14426;
  assign n14429 = ~n14424 & n14428;
  assign n14430 = ~n14427 & ~n14429;
  assign n14431 = n2043 & n7060;
  assign n14432 = pi106  & n2180;
  assign n14433 = pi108  & n2041;
  assign n14434 = pi107  & n2036;
  assign n14435 = ~n14433 & ~n14434;
  assign n14436 = ~n14432 & n14435;
  assign n14437 = ~n14431 & n14436;
  assign n14438 = pi23  & ~n14437;
  assign n14439 = pi23  & ~n14438;
  assign n14440 = ~n14437 & ~n14438;
  assign n14441 = ~n14439 & ~n14440;
  assign n14442 = ~n14430 & ~n14441;
  assign n14443 = ~n14430 & ~n14442;
  assign n14444 = ~n14441 & ~n14442;
  assign n14445 = ~n14443 & ~n14444;
  assign n14446 = ~n14083 & ~n14094;
  assign n14447 = ~n14098 & ~n14446;
  assign n14448 = ~n14445 & ~n14447;
  assign n14449 = n14445 & n14447;
  assign n14450 = ~n14448 & ~n14449;
  assign n14451 = ~n14180 & n14450;
  assign n14452 = ~n14180 & ~n14451;
  assign n14453 = n14450 & ~n14451;
  assign n14454 = ~n14452 & ~n14453;
  assign n14455 = ~n14169 & ~n14454;
  assign n14456 = ~n14169 & ~n14455;
  assign n14457 = ~n14454 & ~n14455;
  assign n14458 = ~n14456 & ~n14457;
  assign n14459 = n1297 & n8936;
  assign n14460 = pi112  & n1366;
  assign n14461 = pi114  & n1295;
  assign n14462 = pi113  & n1290;
  assign n14463 = ~n14461 & ~n14462;
  assign n14464 = ~n14460 & n14463;
  assign n14465 = ~n14459 & n14464;
  assign n14466 = pi17  & ~n14465;
  assign n14467 = pi17  & ~n14466;
  assign n14468 = ~n14465 & ~n14466;
  assign n14469 = ~n14467 & ~n14468;
  assign n14470 = n14458 & n14469;
  assign n14471 = ~n14458 & ~n14469;
  assign n14472 = ~n14470 & ~n14471;
  assign n14473 = ~n14168 & n14472;
  assign n14474 = n14168 & ~n14472;
  assign n14475 = ~n14473 & ~n14474;
  assign n14476 = n938 & n9958;
  assign n14477 = pi115  & n1052;
  assign n14478 = pi117  & n936;
  assign n14479 = pi116  & n931;
  assign n14480 = ~n14478 & ~n14479;
  assign n14481 = ~n14477 & n14480;
  assign n14482 = ~n14476 & n14481;
  assign n14483 = pi14  & ~n14482;
  assign n14484 = pi14  & ~n14483;
  assign n14485 = ~n14482 & ~n14483;
  assign n14486 = ~n14484 & ~n14485;
  assign n14487 = n14475 & ~n14486;
  assign n14488 = n14475 & ~n14487;
  assign n14489 = ~n14486 & ~n14487;
  assign n14490 = ~n14488 & ~n14489;
  assign n14491 = ~n14115 & ~n14118;
  assign n14492 = n14490 & n14491;
  assign n14493 = ~n14490 & ~n14491;
  assign n14494 = ~n14492 & ~n14493;
  assign n14495 = n687 & n11028;
  assign n14496 = pi118  & n763;
  assign n14497 = pi120  & n685;
  assign n14498 = pi119  & n680;
  assign n14499 = ~n14497 & ~n14498;
  assign n14500 = ~n14496 & n14499;
  assign n14501 = ~n14495 & n14500;
  assign n14502 = pi11  & ~n14501;
  assign n14503 = pi11  & ~n14502;
  assign n14504 = ~n14501 & ~n14502;
  assign n14505 = ~n14503 & ~n14504;
  assign n14506 = ~n14494 & n14505;
  assign n14507 = n14494 & ~n14505;
  assign n14508 = ~n14506 & ~n14507;
  assign n14509 = n498 & n12158;
  assign n14510 = pi121  & n537;
  assign n14511 = pi123  & n496;
  assign n14512 = pi122  & n491;
  assign n14513 = ~n14511 & ~n14512;
  assign n14514 = ~n14510 & n14513;
  assign n14515 = ~n14509 & n14514;
  assign n14516 = pi8  & ~n14515;
  assign n14517 = pi8  & ~n14516;
  assign n14518 = ~n14515 & ~n14516;
  assign n14519 = ~n14517 & ~n14518;
  assign n14520 = n14508 & ~n14519;
  assign n14521 = n14508 & ~n14520;
  assign n14522 = ~n14519 & ~n14520;
  assign n14523 = ~n14521 & ~n14522;
  assign n14524 = ~n14121 & ~n14124;
  assign n14525 = n14523 & n14524;
  assign n14526 = ~n14523 & ~n14524;
  assign n14527 = ~n14525 & ~n14526;
  assign n14528 = n342 & n13344;
  assign n14529 = pi124  & n380;
  assign n14530 = pi126  & n340;
  assign n14531 = pi125  & n335;
  assign n14532 = ~n14530 & ~n14531;
  assign n14533 = ~n14529 & n14532;
  assign n14534 = ~n14528 & n14533;
  assign n14535 = pi5  & ~n14534;
  assign n14536 = pi5  & ~n14535;
  assign n14537 = ~n14534 & ~n14535;
  assign n14538 = ~n14536 & ~n14537;
  assign n14539 = n14527 & ~n14538;
  assign n14540 = n14527 & ~n14539;
  assign n14541 = ~n14538 & ~n14539;
  assign n14542 = ~n14540 & ~n14541;
  assign n14543 = ~n14141 & ~n14152;
  assign n14544 = ~n14138 & ~n14543;
  assign n14545 = n262 & n13770;
  assign n14546 = ~pi2  & ~n14545;
  assign n14547 = pi127  & n288;
  assign n14548 = ~n14545 & ~n14547;
  assign n14549 = pi2  & ~n14548;
  assign n14550 = ~n14546 & ~n14549;
  assign n14551 = ~n14544 & n14550;
  assign n14552 = n14544 & ~n14550;
  assign n14553 = ~n14551 & ~n14552;
  assign n14554 = ~n14542 & n14553;
  assign n14555 = ~n14542 & ~n14554;
  assign n14556 = n14553 & ~n14554;
  assign n14557 = ~n14555 & ~n14556;
  assign n14558 = ~n14156 & ~n14159;
  assign n14559 = n14557 & n14558;
  assign n14560 = ~n14557 & ~n14558;
  assign n14561 = ~n14559 & ~n14560;
  assign n14562 = ~n14162 & ~n14165;
  assign n14563 = n14561 & ~n14562;
  assign n14564 = ~n14561 & n14562;
  assign po65  = ~n14563 & ~n14564;
  assign n14566 = ~n14526 & ~n14539;
  assign n14567 = n342 & n13742;
  assign n14568 = pi125  & n380;
  assign n14569 = pi127  & n340;
  assign n14570 = pi126  & n335;
  assign n14571 = ~n14569 & ~n14570;
  assign n14572 = ~n14568 & n14571;
  assign n14573 = ~n14567 & n14572;
  assign n14574 = pi5  & ~n14573;
  assign n14575 = pi5  & ~n14574;
  assign n14576 = ~n14573 & ~n14574;
  assign n14577 = ~n14575 & ~n14576;
  assign n14578 = ~n14566 & ~n14577;
  assign n14579 = ~n14566 & ~n14578;
  assign n14580 = ~n14577 & ~n14578;
  assign n14581 = ~n14579 & ~n14580;
  assign n14582 = n687 & n11389;
  assign n14583 = pi119  & n763;
  assign n14584 = pi121  & n685;
  assign n14585 = pi120  & n680;
  assign n14586 = ~n14584 & ~n14585;
  assign n14587 = ~n14583 & n14586;
  assign n14588 = ~n14582 & n14587;
  assign n14589 = pi11  & ~n14588;
  assign n14590 = pi11  & ~n14589;
  assign n14591 = ~n14588 & ~n14589;
  assign n14592 = ~n14590 & ~n14591;
  assign n14593 = ~n14487 & ~n14493;
  assign n14594 = n14592 & n14593;
  assign n14595 = ~n14592 & ~n14593;
  assign n14596 = ~n14594 & ~n14595;
  assign n14597 = n1297 & n8963;
  assign n14598 = pi113  & n1366;
  assign n14599 = pi115  & n1295;
  assign n14600 = pi114  & n1290;
  assign n14601 = ~n14599 & ~n14600;
  assign n14602 = ~n14598 & n14601;
  assign n14603 = ~n14597 & n14602;
  assign n14604 = pi17  & ~n14603;
  assign n14605 = pi17  & ~n14604;
  assign n14606 = ~n14603 & ~n14604;
  assign n14607 = ~n14605 & ~n14606;
  assign n14608 = ~n14451 & ~n14455;
  assign n14609 = n14607 & n14608;
  assign n14610 = ~n14607 & ~n14608;
  assign n14611 = ~n14609 & ~n14610;
  assign n14612 = n1611 & n7997;
  assign n14613 = pi110  & n1745;
  assign n14614 = pi112  & n1609;
  assign n14615 = pi111  & n1604;
  assign n14616 = ~n14614 & ~n14615;
  assign n14617 = ~n14613 & n14616;
  assign n14618 = ~n14612 & n14617;
  assign n14619 = pi20  & ~n14618;
  assign n14620 = pi20  & ~n14619;
  assign n14621 = ~n14618 & ~n14619;
  assign n14622 = ~n14620 & ~n14621;
  assign n14623 = ~n14442 & ~n14448;
  assign n14624 = n14622 & n14623;
  assign n14625 = ~n14622 & ~n14623;
  assign n14626 = ~n14624 & ~n14625;
  assign n14627 = n2043 & n7349;
  assign n14628 = pi107  & n2180;
  assign n14629 = pi109  & n2041;
  assign n14630 = pi108  & n2036;
  assign n14631 = ~n14629 & ~n14630;
  assign n14632 = ~n14628 & n14631;
  assign n14633 = ~n14627 & n14632;
  assign n14634 = pi23  & ~n14633;
  assign n14635 = pi23  & ~n14634;
  assign n14636 = ~n14633 & ~n14634;
  assign n14637 = ~n14635 & ~n14636;
  assign n14638 = ~n14428 & n14637;
  assign n14639 = n14428 & ~n14637;
  assign n14640 = ~n14638 & ~n14639;
  assign n14641 = n2523 & n6477;
  assign n14642 = pi104  & n2667;
  assign n14643 = pi106  & n2521;
  assign n14644 = pi105  & n2516;
  assign n14645 = ~n14643 & ~n14644;
  assign n14646 = ~n14642 & n14645;
  assign n14647 = ~n14641 & n14646;
  assign n14648 = pi26  & ~n14647;
  assign n14649 = pi26  & ~n14648;
  assign n14650 = ~n14647 & ~n14648;
  assign n14651 = ~n14649 & ~n14650;
  assign n14652 = ~n14404 & ~n14410;
  assign n14653 = n14651 & n14652;
  assign n14654 = ~n14651 & ~n14652;
  assign n14655 = ~n14653 & ~n14654;
  assign n14656 = ~n14385 & ~n14391;
  assign n14657 = pi101  & n3225;
  assign n14658 = pi103  & n3032;
  assign n14659 = pi102  & n3027;
  assign n14660 = ~n14658 & ~n14659;
  assign n14661 = ~n14657 & n14660;
  assign n14662 = ~n3034 & n14661;
  assign n14663 = ~n5664 & n14661;
  assign n14664 = ~n14662 & ~n14663;
  assign n14665 = pi29  & ~n14664;
  assign n14666 = ~pi29  & n14664;
  assign n14667 = ~n14665 & ~n14666;
  assign n14668 = ~n14656 & ~n14667;
  assign n14669 = n14656 & n14667;
  assign n14670 = ~n14668 & ~n14669;
  assign n14671 = ~n14242 & ~n14244;
  assign n14672 = ~n14203 & ~n14209;
  assign n14673 = pi66  & n13835;
  assign n14674 = pi67  & ~n13434;
  assign n14675 = ~n14673 & ~n14674;
  assign n14676 = pi2  & ~n14675;
  assign n14677 = ~pi2  & n14675;
  assign n14678 = ~n14676 & ~n14677;
  assign n14679 = pi68  & n13004;
  assign n14680 = pi70  & n12625;
  assign n14681 = pi69  & n12620;
  assign n14682 = ~n14680 & ~n14681;
  assign n14683 = ~n14679 & n14682;
  assign n14684 = ~n12627 & n14683;
  assign n14685 = ~n450 & n14683;
  assign n14686 = ~n14684 & ~n14685;
  assign n14687 = pi62  & ~n14686;
  assign n14688 = ~pi62  & n14686;
  assign n14689 = ~n14687 & ~n14688;
  assign n14690 = n14678 & ~n14689;
  assign n14691 = ~n14678 & n14689;
  assign n14692 = ~n14690 & ~n14691;
  assign n14693 = ~n14672 & n14692;
  assign n14694 = n14672 & ~n14692;
  assign n14695 = ~n14693 & ~n14694;
  assign n14696 = n642 & n11488;
  assign n14697 = pi71  & n11847;
  assign n14698 = pi73  & n11486;
  assign n14699 = pi72  & n11481;
  assign n14700 = ~n14698 & ~n14699;
  assign n14701 = ~n14697 & n14700;
  assign n14702 = ~n14696 & n14701;
  assign n14703 = pi59  & ~n14702;
  assign n14704 = pi59  & ~n14703;
  assign n14705 = ~n14702 & ~n14703;
  assign n14706 = ~n14704 & ~n14705;
  assign n14707 = n14695 & ~n14706;
  assign n14708 = n14695 & ~n14707;
  assign n14709 = ~n14706 & ~n14707;
  assign n14710 = ~n14708 & ~n14709;
  assign n14711 = ~n14227 & n14710;
  assign n14712 = n14227 & ~n14710;
  assign n14713 = ~n14711 & ~n14712;
  assign n14714 = n891 & n10394;
  assign n14715 = pi74  & n10744;
  assign n14716 = pi76  & n10392;
  assign n14717 = pi75  & n10387;
  assign n14718 = ~n14716 & ~n14717;
  assign n14719 = ~n14715 & n14718;
  assign n14720 = ~n14714 & n14719;
  assign n14721 = pi56  & ~n14720;
  assign n14722 = pi56  & ~n14721;
  assign n14723 = ~n14720 & ~n14721;
  assign n14724 = ~n14722 & ~n14723;
  assign n14725 = n14713 & n14724;
  assign n14726 = ~n14713 & ~n14724;
  assign n14727 = ~n14725 & ~n14726;
  assign n14728 = ~n14671 & n14727;
  assign n14729 = n14671 & ~n14727;
  assign n14730 = ~n14728 & ~n14729;
  assign n14731 = n1122 & n9310;
  assign n14732 = pi77  & n9701;
  assign n14733 = pi79  & n9308;
  assign n14734 = pi78  & n9303;
  assign n14735 = ~n14733 & ~n14734;
  assign n14736 = ~n14732 & n14735;
  assign n14737 = ~n14731 & n14736;
  assign n14738 = pi53  & ~n14737;
  assign n14739 = pi53  & ~n14738;
  assign n14740 = ~n14737 & ~n14738;
  assign n14741 = ~n14739 & ~n14740;
  assign n14742 = n14730 & ~n14741;
  assign n14743 = n14730 & ~n14742;
  assign n14744 = ~n14741 & ~n14742;
  assign n14745 = ~n14743 & ~n14744;
  assign n14746 = ~n14186 & ~n14261;
  assign n14747 = ~n14258 & ~n14746;
  assign n14748 = n14745 & n14747;
  assign n14749 = ~n14745 & ~n14747;
  assign n14750 = ~n14748 & ~n14749;
  assign n14751 = n1554 & n8334;
  assign n14752 = pi80  & n8685;
  assign n14753 = pi82  & n8332;
  assign n14754 = pi81  & n8327;
  assign n14755 = ~n14753 & ~n14754;
  assign n14756 = ~n14752 & n14755;
  assign n14757 = ~n14751 & n14756;
  assign n14758 = pi50  & ~n14757;
  assign n14759 = pi50  & ~n14758;
  assign n14760 = ~n14757 & ~n14758;
  assign n14761 = ~n14759 & ~n14760;
  assign n14762 = n14750 & ~n14761;
  assign n14763 = n14750 & ~n14762;
  assign n14764 = ~n14761 & ~n14762;
  assign n14765 = ~n14763 & ~n14764;
  assign n14766 = ~n14276 & ~n14280;
  assign n14767 = n14765 & n14766;
  assign n14768 = ~n14765 & ~n14766;
  assign n14769 = ~n14767 & ~n14768;
  assign n14770 = n1972 & n7408;
  assign n14771 = pi83  & n7740;
  assign n14772 = pi85  & n7406;
  assign n14773 = pi84  & n7401;
  assign n14774 = ~n14772 & ~n14773;
  assign n14775 = ~n14771 & n14774;
  assign n14776 = ~n14770 & n14775;
  assign n14777 = pi47  & ~n14776;
  assign n14778 = pi47  & ~n14777;
  assign n14779 = ~n14776 & ~n14777;
  assign n14780 = ~n14778 & ~n14779;
  assign n14781 = ~n14769 & n14780;
  assign n14782 = n14769 & ~n14780;
  assign n14783 = ~n14781 & ~n14782;
  assign n14784 = ~n14184 & ~n14296;
  assign n14785 = ~n14293 & ~n14784;
  assign n14786 = n14783 & ~n14785;
  assign n14787 = ~n14783 & n14785;
  assign n14788 = ~n14786 & ~n14787;
  assign n14789 = n2446 & n6539;
  assign n14790 = pi86  & n6873;
  assign n14791 = pi88  & n6537;
  assign n14792 = pi87  & n6532;
  assign n14793 = ~n14791 & ~n14792;
  assign n14794 = ~n14790 & n14793;
  assign n14795 = ~n14789 & n14794;
  assign n14796 = pi44  & ~n14795;
  assign n14797 = pi44  & ~n14796;
  assign n14798 = ~n14795 & ~n14796;
  assign n14799 = ~n14797 & ~n14798;
  assign n14800 = n14788 & ~n14799;
  assign n14801 = n14788 & ~n14800;
  assign n14802 = ~n14799 & ~n14800;
  assign n14803 = ~n14801 & ~n14802;
  assign n14804 = ~n14311 & ~n14315;
  assign n14805 = n14803 & n14804;
  assign n14806 = ~n14803 & ~n14804;
  assign n14807 = ~n14805 & ~n14806;
  assign n14808 = n2978 & n5739;
  assign n14809 = pi89  & n6030;
  assign n14810 = pi91  & n5737;
  assign n14811 = pi90  & n5732;
  assign n14812 = ~n14810 & ~n14811;
  assign n14813 = ~n14809 & n14812;
  assign n14814 = ~n14808 & n14813;
  assign n14815 = pi41  & ~n14814;
  assign n14816 = pi41  & ~n14815;
  assign n14817 = ~n14814 & ~n14815;
  assign n14818 = ~n14816 & ~n14817;
  assign n14819 = n14807 & ~n14818;
  assign n14820 = n14807 & ~n14819;
  assign n14821 = ~n14818 & ~n14819;
  assign n14822 = ~n14820 & ~n14821;
  assign n14823 = ~n14328 & ~n14334;
  assign n14824 = n14822 & n14823;
  assign n14825 = ~n14822 & ~n14823;
  assign n14826 = ~n14824 & ~n14825;
  assign n14827 = n3565 & n5008;
  assign n14828 = pi92  & n5241;
  assign n14829 = pi94  & n5006;
  assign n14830 = pi93  & n5001;
  assign n14831 = ~n14829 & ~n14830;
  assign n14832 = ~n14828 & n14831;
  assign n14833 = ~n14827 & n14832;
  assign n14834 = pi38  & ~n14833;
  assign n14835 = pi38  & ~n14834;
  assign n14836 = ~n14833 & ~n14834;
  assign n14837 = ~n14835 & ~n14836;
  assign n14838 = ~n14826 & n14837;
  assign n14839 = n14826 & ~n14837;
  assign n14840 = ~n14838 & ~n14839;
  assign n14841 = ~n14347 & ~n14353;
  assign n14842 = n14840 & ~n14841;
  assign n14843 = ~n14840 & n14841;
  assign n14844 = ~n14842 & ~n14843;
  assign n14845 = n4211 & n4271;
  assign n14846 = pi95  & n4503;
  assign n14847 = pi97  & n4269;
  assign n14848 = pi96  & n4264;
  assign n14849 = ~n14847 & ~n14848;
  assign n14850 = ~n14846 & n14849;
  assign n14851 = ~n14845 & n14850;
  assign n14852 = pi35  & ~n14851;
  assign n14853 = pi35  & ~n14852;
  assign n14854 = ~n14851 & ~n14852;
  assign n14855 = ~n14853 & ~n14854;
  assign n14856 = n14844 & ~n14855;
  assign n14857 = n14844 & ~n14856;
  assign n14858 = ~n14855 & ~n14856;
  assign n14859 = ~n14857 & ~n14858;
  assign n14860 = pi98  & n3814;
  assign n14861 = pi100  & n3620;
  assign n14862 = pi99  & n3615;
  assign n14863 = ~n14861 & ~n14862;
  assign n14864 = ~n14860 & n14863;
  assign n14865 = ~n3622 & n14864;
  assign n14866 = ~n4910 & n14864;
  assign n14867 = ~n14865 & ~n14866;
  assign n14868 = pi32  & ~n14867;
  assign n14869 = ~pi32  & n14867;
  assign n14870 = ~n14868 & ~n14869;
  assign n14871 = ~n14371 & ~n14870;
  assign n14872 = ~n14371 & ~n14871;
  assign n14873 = ~n14870 & ~n14871;
  assign n14874 = ~n14872 & ~n14873;
  assign n14875 = ~n14859 & ~n14874;
  assign n14876 = ~n14859 & ~n14875;
  assign n14877 = ~n14874 & ~n14875;
  assign n14878 = ~n14876 & ~n14877;
  assign n14879 = n14670 & ~n14878;
  assign n14880 = n14670 & ~n14879;
  assign n14881 = ~n14878 & ~n14879;
  assign n14882 = ~n14880 & ~n14881;
  assign n14883 = n14655 & ~n14882;
  assign n14884 = ~n14655 & n14882;
  assign n14885 = ~n14883 & ~n14884;
  assign n14886 = ~n14640 & n14885;
  assign n14887 = ~n14640 & ~n14886;
  assign n14888 = n14885 & ~n14886;
  assign n14889 = ~n14887 & ~n14888;
  assign n14890 = n14626 & ~n14889;
  assign n14891 = ~n14626 & n14889;
  assign n14892 = ~n14890 & ~n14891;
  assign n14893 = n14611 & n14892;
  assign n14894 = n14611 & ~n14893;
  assign n14895 = n14892 & ~n14893;
  assign n14896 = ~n14894 & ~n14895;
  assign n14897 = ~n14471 & ~n14473;
  assign n14898 = pi116  & n1052;
  assign n14899 = pi118  & n936;
  assign n14900 = pi117  & n931;
  assign n14901 = ~n14899 & ~n14900;
  assign n14902 = ~n14898 & n14901;
  assign n14903 = ~n938 & n14902;
  assign n14904 = ~n9984 & n14902;
  assign n14905 = ~n14903 & ~n14904;
  assign n14906 = pi14  & ~n14905;
  assign n14907 = ~pi14  & n14905;
  assign n14908 = ~n14906 & ~n14907;
  assign n14909 = ~n14897 & ~n14908;
  assign n14910 = ~n14897 & ~n14909;
  assign n14911 = ~n14908 & ~n14909;
  assign n14912 = ~n14910 & ~n14911;
  assign n14913 = ~n14896 & ~n14912;
  assign n14914 = ~n14896 & ~n14913;
  assign n14915 = ~n14912 & ~n14913;
  assign n14916 = ~n14914 & ~n14915;
  assign n14917 = n14596 & ~n14916;
  assign n14918 = n14596 & ~n14917;
  assign n14919 = ~n14916 & ~n14917;
  assign n14920 = ~n14918 & ~n14919;
  assign n14921 = n498 & n12189;
  assign n14922 = pi122  & n537;
  assign n14923 = pi124  & n496;
  assign n14924 = pi123  & n491;
  assign n14925 = ~n14923 & ~n14924;
  assign n14926 = ~n14922 & n14925;
  assign n14927 = ~n14921 & n14926;
  assign n14928 = pi8  & ~n14927;
  assign n14929 = pi8  & ~n14928;
  assign n14930 = ~n14927 & ~n14928;
  assign n14931 = ~n14929 & ~n14930;
  assign n14932 = ~n14507 & ~n14520;
  assign n14933 = ~n14931 & ~n14932;
  assign n14934 = ~n14931 & ~n14933;
  assign n14935 = ~n14932 & ~n14933;
  assign n14936 = ~n14934 & ~n14935;
  assign n14937 = ~n14920 & ~n14936;
  assign n14938 = ~n14920 & ~n14937;
  assign n14939 = ~n14936 & ~n14937;
  assign n14940 = ~n14938 & ~n14939;
  assign n14941 = ~n14581 & ~n14940;
  assign n14942 = ~n14581 & ~n14941;
  assign n14943 = ~n14940 & ~n14941;
  assign n14944 = ~n14942 & ~n14943;
  assign n14945 = ~n14551 & ~n14554;
  assign n14946 = n14944 & n14945;
  assign n14947 = ~n14944 & ~n14945;
  assign n14948 = ~n14946 & ~n14947;
  assign n14949 = ~n14560 & ~n14563;
  assign n14950 = n14948 & ~n14949;
  assign n14951 = ~n14948 & n14949;
  assign po66  = ~n14950 & ~n14951;
  assign n14953 = ~n14947 & ~n14950;
  assign n14954 = ~n14578 & ~n14941;
  assign n14955 = n938 & n10667;
  assign n14956 = pi117  & n1052;
  assign n14957 = pi119  & n936;
  assign n14958 = pi118  & n931;
  assign n14959 = ~n14957 & ~n14958;
  assign n14960 = ~n14956 & n14959;
  assign n14961 = ~n14955 & n14960;
  assign n14962 = pi14  & ~n14961;
  assign n14963 = pi14  & ~n14962;
  assign n14964 = ~n14961 & ~n14962;
  assign n14965 = ~n14963 & ~n14964;
  assign n14966 = ~n14610 & ~n14893;
  assign n14967 = n14965 & n14966;
  assign n14968 = ~n14965 & ~n14966;
  assign n14969 = ~n14967 & ~n14968;
  assign n14970 = n1611 & n8612;
  assign n14971 = pi111  & n1745;
  assign n14972 = pi113  & n1609;
  assign n14973 = pi112  & n1604;
  assign n14974 = ~n14972 & ~n14973;
  assign n14975 = ~n14971 & n14974;
  assign n14976 = ~n14970 & n14975;
  assign n14977 = pi20  & ~n14976;
  assign n14978 = pi20  & ~n14977;
  assign n14979 = ~n14976 & ~n14977;
  assign n14980 = ~n14978 & ~n14979;
  assign n14981 = ~n14428 & ~n14637;
  assign n14982 = ~n14886 & ~n14981;
  assign n14983 = n14980 & n14982;
  assign n14984 = ~n14980 & ~n14982;
  assign n14985 = ~n14983 & ~n14984;
  assign n14986 = n2523 & n6775;
  assign n14987 = pi105  & n2667;
  assign n14988 = pi107  & n2521;
  assign n14989 = pi106  & n2516;
  assign n14990 = ~n14988 & ~n14989;
  assign n14991 = ~n14987 & n14990;
  assign n14992 = ~n14986 & n14991;
  assign n14993 = pi26  & ~n14992;
  assign n14994 = pi26  & ~n14993;
  assign n14995 = ~n14992 & ~n14993;
  assign n14996 = ~n14994 & ~n14995;
  assign n14997 = ~n14668 & ~n14879;
  assign n14998 = n14996 & n14997;
  assign n14999 = ~n14996 & ~n14997;
  assign n15000 = ~n14998 & ~n14999;
  assign n15001 = ~n14842 & ~n14856;
  assign n15002 = pi99  & n3814;
  assign n15003 = pi101  & n3620;
  assign n15004 = pi100  & n3615;
  assign n15005 = ~n15003 & ~n15004;
  assign n15006 = ~n15002 & n15005;
  assign n15007 = ~n3622 & n15006;
  assign n15008 = ~n5169 & n15006;
  assign n15009 = ~n15007 & ~n15008;
  assign n15010 = pi32  & ~n15009;
  assign n15011 = ~pi32  & n15009;
  assign n15012 = ~n15010 & ~n15011;
  assign n15013 = ~n15001 & ~n15012;
  assign n15014 = n15001 & n15012;
  assign n15015 = ~n15013 & ~n15014;
  assign n15016 = n4271 & n4454;
  assign n15017 = pi96  & n4503;
  assign n15018 = pi98  & n4269;
  assign n15019 = pi97  & n4264;
  assign n15020 = ~n15018 & ~n15019;
  assign n15021 = ~n15017 & n15020;
  assign n15022 = ~n15016 & n15021;
  assign n15023 = pi35  & ~n15022;
  assign n15024 = pi35  & ~n15023;
  assign n15025 = ~n15022 & ~n15023;
  assign n15026 = ~n15024 & ~n15025;
  assign n15027 = ~n14825 & ~n14839;
  assign n15028 = n475 & n12627;
  assign n15029 = pi69  & n13004;
  assign n15030 = pi71  & n12625;
  assign n15031 = pi70  & n12620;
  assign n15032 = ~n15030 & ~n15031;
  assign n15033 = ~n15029 & n15032;
  assign n15034 = ~n15028 & n15033;
  assign n15035 = pi62  & ~n15034;
  assign n15036 = pi62  & ~n15035;
  assign n15037 = ~n15034 & ~n15035;
  assign n15038 = ~n15036 & ~n15037;
  assign n15039 = pi67  & n13835;
  assign n15040 = pi68  & ~n13434;
  assign n15041 = ~n15039 & ~n15040;
  assign n15042 = pi2  & ~n15041;
  assign n15043 = pi2  & ~n15042;
  assign n15044 = ~n15041 & ~n15042;
  assign n15045 = ~n15043 & ~n15044;
  assign n15046 = ~n15038 & ~n15045;
  assign n15047 = ~n15038 & ~n15046;
  assign n15048 = ~n15045 & ~n15046;
  assign n15049 = ~n15047 & ~n15048;
  assign n15050 = ~n14676 & ~n14690;
  assign n15051 = n15049 & n15050;
  assign n15052 = ~n15049 & ~n15050;
  assign n15053 = ~n15051 & ~n15052;
  assign n15054 = n729 & n11488;
  assign n15055 = pi72  & n11847;
  assign n15056 = pi74  & n11486;
  assign n15057 = pi73  & n11481;
  assign n15058 = ~n15056 & ~n15057;
  assign n15059 = ~n15055 & n15058;
  assign n15060 = ~n15054 & n15059;
  assign n15061 = pi59  & ~n15060;
  assign n15062 = pi59  & ~n15061;
  assign n15063 = ~n15060 & ~n15061;
  assign n15064 = ~n15062 & ~n15063;
  assign n15065 = n15053 & ~n15064;
  assign n15066 = n15053 & ~n15065;
  assign n15067 = ~n15064 & ~n15065;
  assign n15068 = ~n15066 & ~n15067;
  assign n15069 = ~n14693 & ~n14707;
  assign n15070 = n15068 & n15069;
  assign n15071 = ~n15068 & ~n15069;
  assign n15072 = ~n15070 & ~n15071;
  assign n15073 = n999 & n10394;
  assign n15074 = pi75  & n10744;
  assign n15075 = pi77  & n10392;
  assign n15076 = pi76  & n10387;
  assign n15077 = ~n15075 & ~n15076;
  assign n15078 = ~n15074 & n15077;
  assign n15079 = ~n15073 & n15078;
  assign n15080 = pi56  & ~n15079;
  assign n15081 = pi56  & ~n15080;
  assign n15082 = ~n15079 & ~n15080;
  assign n15083 = ~n15081 & ~n15082;
  assign n15084 = ~n15072 & n15083;
  assign n15085 = n15072 & ~n15083;
  assign n15086 = ~n15084 & ~n15085;
  assign n15087 = ~n14227 & ~n14710;
  assign n15088 = ~n14726 & ~n15087;
  assign n15089 = n15086 & ~n15088;
  assign n15090 = ~n15086 & n15088;
  assign n15091 = ~n15089 & ~n15090;
  assign n15092 = n1225 & n9310;
  assign n15093 = pi78  & n9701;
  assign n15094 = pi80  & n9308;
  assign n15095 = pi79  & n9303;
  assign n15096 = ~n15094 & ~n15095;
  assign n15097 = ~n15093 & n15096;
  assign n15098 = ~n15092 & n15097;
  assign n15099 = pi53  & ~n15098;
  assign n15100 = pi53  & ~n15099;
  assign n15101 = ~n15098 & ~n15099;
  assign n15102 = ~n15100 & ~n15101;
  assign n15103 = n15091 & ~n15102;
  assign n15104 = n15091 & ~n15103;
  assign n15105 = ~n15102 & ~n15103;
  assign n15106 = ~n15104 & ~n15105;
  assign n15107 = ~n14728 & ~n14742;
  assign n15108 = n15106 & n15107;
  assign n15109 = ~n15106 & ~n15107;
  assign n15110 = ~n15108 & ~n15109;
  assign n15111 = n1696 & n8334;
  assign n15112 = pi81  & n8685;
  assign n15113 = pi83  & n8332;
  assign n15114 = pi82  & n8327;
  assign n15115 = ~n15113 & ~n15114;
  assign n15116 = ~n15112 & n15115;
  assign n15117 = ~n15111 & n15116;
  assign n15118 = pi50  & ~n15117;
  assign n15119 = pi50  & ~n15118;
  assign n15120 = ~n15117 & ~n15118;
  assign n15121 = ~n15119 & ~n15120;
  assign n15122 = n15110 & ~n15121;
  assign n15123 = n15110 & ~n15122;
  assign n15124 = ~n15121 & ~n15122;
  assign n15125 = ~n15123 & ~n15124;
  assign n15126 = ~n14749 & ~n14762;
  assign n15127 = n15125 & n15126;
  assign n15128 = ~n15125 & ~n15126;
  assign n15129 = ~n15127 & ~n15128;
  assign n15130 = n2133 & n7408;
  assign n15131 = pi84  & n7740;
  assign n15132 = pi86  & n7406;
  assign n15133 = pi85  & n7401;
  assign n15134 = ~n15132 & ~n15133;
  assign n15135 = ~n15131 & n15134;
  assign n15136 = ~n15130 & n15135;
  assign n15137 = pi47  & ~n15136;
  assign n15138 = pi47  & ~n15137;
  assign n15139 = ~n15136 & ~n15137;
  assign n15140 = ~n15138 & ~n15139;
  assign n15141 = n15129 & ~n15140;
  assign n15142 = n15129 & ~n15141;
  assign n15143 = ~n15140 & ~n15141;
  assign n15144 = ~n15142 & ~n15143;
  assign n15145 = ~n14768 & ~n14782;
  assign n15146 = ~n15144 & ~n15145;
  assign n15147 = ~n15144 & ~n15146;
  assign n15148 = ~n15145 & ~n15146;
  assign n15149 = ~n15147 & ~n15148;
  assign n15150 = n2473 & n6539;
  assign n15151 = pi87  & n6873;
  assign n15152 = pi89  & n6537;
  assign n15153 = pi88  & n6532;
  assign n15154 = ~n15152 & ~n15153;
  assign n15155 = ~n15151 & n15154;
  assign n15156 = ~n15150 & n15155;
  assign n15157 = pi44  & ~n15156;
  assign n15158 = pi44  & ~n15157;
  assign n15159 = ~n15156 & ~n15157;
  assign n15160 = ~n15158 & ~n15159;
  assign n15161 = ~n15149 & ~n15160;
  assign n15162 = ~n15149 & ~n15161;
  assign n15163 = ~n15160 & ~n15161;
  assign n15164 = ~n15162 & ~n15163;
  assign n15165 = ~n14786 & ~n14800;
  assign n15166 = n15164 & n15165;
  assign n15167 = ~n15164 & ~n15165;
  assign n15168 = ~n15166 & ~n15167;
  assign n15169 = n3177 & n5739;
  assign n15170 = pi90  & n6030;
  assign n15171 = pi92  & n5737;
  assign n15172 = pi91  & n5732;
  assign n15173 = ~n15171 & ~n15172;
  assign n15174 = ~n15170 & n15173;
  assign n15175 = ~n15169 & n15174;
  assign n15176 = pi41  & ~n15175;
  assign n15177 = pi41  & ~n15176;
  assign n15178 = ~n15175 & ~n15176;
  assign n15179 = ~n15177 & ~n15178;
  assign n15180 = n15168 & ~n15179;
  assign n15181 = n15168 & ~n15180;
  assign n15182 = ~n15179 & ~n15180;
  assign n15183 = ~n15181 & ~n15182;
  assign n15184 = ~n14806 & ~n14819;
  assign n15185 = n15183 & n15184;
  assign n15186 = ~n15183 & ~n15184;
  assign n15187 = ~n15185 & ~n15186;
  assign n15188 = n3784 & n5008;
  assign n15189 = pi93  & n5241;
  assign n15190 = pi95  & n5006;
  assign n15191 = pi94  & n5001;
  assign n15192 = ~n15190 & ~n15191;
  assign n15193 = ~n15189 & n15192;
  assign n15194 = ~n15188 & n15193;
  assign n15195 = pi38  & ~n15194;
  assign n15196 = pi38  & ~n15195;
  assign n15197 = ~n15194 & ~n15195;
  assign n15198 = ~n15196 & ~n15197;
  assign n15199 = ~n15187 & n15198;
  assign n15200 = n15187 & ~n15198;
  assign n15201 = ~n15199 & ~n15200;
  assign n15202 = ~n15027 & n15201;
  assign n15203 = ~n15027 & ~n15202;
  assign n15204 = n15201 & ~n15202;
  assign n15205 = ~n15203 & ~n15204;
  assign n15206 = ~n15026 & ~n15205;
  assign n15207 = ~n15026 & ~n15206;
  assign n15208 = ~n15205 & ~n15206;
  assign n15209 = ~n15207 & ~n15208;
  assign n15210 = ~n15015 & n15209;
  assign n15211 = n15015 & ~n15209;
  assign n15212 = ~n15210 & ~n15211;
  assign n15213 = ~n14871 & ~n14875;
  assign n15214 = pi102  & n3225;
  assign n15215 = pi104  & n3032;
  assign n15216 = pi103  & n3027;
  assign n15217 = ~n15215 & ~n15216;
  assign n15218 = ~n15214 & n15217;
  assign n15219 = ~n3034 & n15218;
  assign n15220 = ~n5943 & n15218;
  assign n15221 = ~n15219 & ~n15220;
  assign n15222 = pi29  & ~n15221;
  assign n15223 = ~pi29  & n15221;
  assign n15224 = ~n15222 & ~n15223;
  assign n15225 = ~n15213 & ~n15224;
  assign n15226 = ~n15213 & ~n15225;
  assign n15227 = ~n15224 & ~n15225;
  assign n15228 = ~n15226 & ~n15227;
  assign n15229 = n15212 & ~n15228;
  assign n15230 = n15212 & ~n15229;
  assign n15231 = ~n15228 & ~n15229;
  assign n15232 = ~n15230 & ~n15231;
  assign n15233 = n15000 & ~n15232;
  assign n15234 = n15000 & ~n15233;
  assign n15235 = ~n15232 & ~n15233;
  assign n15236 = ~n15234 & ~n15235;
  assign n15237 = n2043 & n7665;
  assign n15238 = pi108  & n2180;
  assign n15239 = pi110  & n2041;
  assign n15240 = pi109  & n2036;
  assign n15241 = ~n15239 & ~n15240;
  assign n15242 = ~n15238 & n15241;
  assign n15243 = ~n15237 & n15242;
  assign n15244 = pi23  & ~n15243;
  assign n15245 = pi23  & ~n15244;
  assign n15246 = ~n15243 & ~n15244;
  assign n15247 = ~n15245 & ~n15246;
  assign n15248 = ~n14654 & ~n14883;
  assign n15249 = ~n15247 & ~n15248;
  assign n15250 = ~n15247 & ~n15249;
  assign n15251 = ~n15248 & ~n15249;
  assign n15252 = ~n15250 & ~n15251;
  assign n15253 = ~n15236 & n15252;
  assign n15254 = n15236 & ~n15252;
  assign n15255 = ~n15253 & ~n15254;
  assign n15256 = n14985 & ~n15255;
  assign n15257 = n14985 & ~n15256;
  assign n15258 = ~n15255 & ~n15256;
  assign n15259 = ~n15257 & ~n15258;
  assign n15260 = n1297 & n9614;
  assign n15261 = pi114  & n1366;
  assign n15262 = pi116  & n1295;
  assign n15263 = pi115  & n1290;
  assign n15264 = ~n15262 & ~n15263;
  assign n15265 = ~n15261 & n15264;
  assign n15266 = ~n15260 & n15265;
  assign n15267 = pi17  & ~n15266;
  assign n15268 = pi17  & ~n15267;
  assign n15269 = ~n15266 & ~n15267;
  assign n15270 = ~n15268 & ~n15269;
  assign n15271 = ~n14625 & ~n14890;
  assign n15272 = ~n15270 & ~n15271;
  assign n15273 = ~n15270 & ~n15272;
  assign n15274 = ~n15271 & ~n15272;
  assign n15275 = ~n15273 & ~n15274;
  assign n15276 = ~n15259 & n15275;
  assign n15277 = n15259 & ~n15275;
  assign n15278 = ~n15276 & ~n15277;
  assign n15279 = n14969 & ~n15278;
  assign n15280 = n14969 & ~n15279;
  assign n15281 = ~n15278 & ~n15279;
  assign n15282 = ~n15280 & ~n15281;
  assign n15283 = ~n14909 & ~n14913;
  assign n15284 = pi120  & n763;
  assign n15285 = pi122  & n685;
  assign n15286 = pi121  & n680;
  assign n15287 = ~n15285 & ~n15286;
  assign n15288 = ~n15284 & n15287;
  assign n15289 = ~n687 & n15288;
  assign n15290 = ~n11778 & n15288;
  assign n15291 = ~n15289 & ~n15290;
  assign n15292 = pi11  & ~n15291;
  assign n15293 = ~pi11  & n15291;
  assign n15294 = ~n15292 & ~n15293;
  assign n15295 = ~n15283 & ~n15294;
  assign n15296 = ~n15283 & ~n15295;
  assign n15297 = ~n15294 & ~n15295;
  assign n15298 = ~n15296 & ~n15297;
  assign n15299 = ~n15282 & ~n15298;
  assign n15300 = ~n15282 & ~n15299;
  assign n15301 = ~n15298 & ~n15299;
  assign n15302 = ~n15300 & ~n15301;
  assign n15303 = ~n14595 & ~n14917;
  assign n15304 = pi123  & n537;
  assign n15305 = pi125  & n496;
  assign n15306 = pi124  & n491;
  assign n15307 = ~n15305 & ~n15306;
  assign n15308 = ~n15304 & n15307;
  assign n15309 = ~n498 & n15308;
  assign n15310 = ~n12943 & n15308;
  assign n15311 = ~n15309 & ~n15310;
  assign n15312 = pi8  & ~n15311;
  assign n15313 = ~pi8  & n15311;
  assign n15314 = ~n15312 & ~n15313;
  assign n15315 = ~n15303 & ~n15314;
  assign n15316 = ~n15303 & ~n15315;
  assign n15317 = ~n15314 & ~n15315;
  assign n15318 = ~n15316 & ~n15317;
  assign n15319 = ~n15302 & ~n15318;
  assign n15320 = ~n15302 & ~n15319;
  assign n15321 = ~n15318 & ~n15319;
  assign n15322 = ~n15320 & ~n15321;
  assign n15323 = ~n14933 & ~n14937;
  assign n15324 = pi126  & n380;
  assign n15325 = pi127  & n335;
  assign n15326 = ~n15324 & ~n15325;
  assign n15327 = ~n342 & n15326;
  assign n15328 = n13773 & n15326;
  assign n15329 = ~n15327 & ~n15328;
  assign n15330 = pi5  & ~n15329;
  assign n15331 = ~pi5  & n15329;
  assign n15332 = ~n15330 & ~n15331;
  assign n15333 = ~n15323 & ~n15332;
  assign n15334 = ~n15323 & ~n15333;
  assign n15335 = ~n15332 & ~n15333;
  assign n15336 = ~n15334 & ~n15335;
  assign n15337 = ~n15322 & ~n15336;
  assign n15338 = n15322 & n15336;
  assign n15339 = ~n15337 & ~n15338;
  assign n15340 = ~n14954 & n15339;
  assign n15341 = ~n14954 & ~n15340;
  assign n15342 = n15339 & ~n15340;
  assign n15343 = ~n15341 & ~n15342;
  assign n15344 = ~n14953 & ~n15343;
  assign n15345 = n14953 & n15343;
  assign po67  = ~n15344 & ~n15345;
  assign n15347 = ~n15340 & ~n15344;
  assign n15348 = ~n15333 & ~n15337;
  assign n15349 = ~n15315 & ~n15319;
  assign n15350 = pi127  & n380;
  assign n15351 = n342 & n13770;
  assign n15352 = ~n15350 & ~n15351;
  assign n15353 = pi5  & ~n15352;
  assign n15354 = pi5  & ~n15353;
  assign n15355 = ~n15352 & ~n15353;
  assign n15356 = ~n15354 & ~n15355;
  assign n15357 = ~n15349 & ~n15356;
  assign n15358 = ~n15349 & ~n15357;
  assign n15359 = ~n15356 & ~n15357;
  assign n15360 = ~n15358 & ~n15359;
  assign n15361 = n687 & n12158;
  assign n15362 = pi121  & n763;
  assign n15363 = pi123  & n685;
  assign n15364 = pi122  & n680;
  assign n15365 = ~n15363 & ~n15364;
  assign n15366 = ~n15362 & n15365;
  assign n15367 = ~n15361 & n15366;
  assign n15368 = pi11  & ~n15367;
  assign n15369 = pi11  & ~n15368;
  assign n15370 = ~n15367 & ~n15368;
  assign n15371 = ~n15369 & ~n15370;
  assign n15372 = ~n14968 & ~n15279;
  assign n15373 = n15371 & n15372;
  assign n15374 = ~n15371 & ~n15372;
  assign n15375 = ~n15373 & ~n15374;
  assign n15376 = n938 & n11028;
  assign n15377 = pi118  & n1052;
  assign n15378 = pi120  & n936;
  assign n15379 = pi119  & n931;
  assign n15380 = ~n15378 & ~n15379;
  assign n15381 = ~n15377 & n15380;
  assign n15382 = ~n15376 & n15381;
  assign n15383 = pi14  & ~n15382;
  assign n15384 = pi14  & ~n15383;
  assign n15385 = ~n15382 & ~n15383;
  assign n15386 = ~n15384 & ~n15385;
  assign n15387 = ~n15259 & ~n15275;
  assign n15388 = ~n15272 & ~n15387;
  assign n15389 = ~n15386 & ~n15388;
  assign n15390 = ~n15386 & ~n15389;
  assign n15391 = ~n15388 & ~n15389;
  assign n15392 = ~n15390 & ~n15391;
  assign n15393 = ~n14984 & ~n15256;
  assign n15394 = pi115  & n1366;
  assign n15395 = pi117  & n1295;
  assign n15396 = pi116  & n1290;
  assign n15397 = ~n15395 & ~n15396;
  assign n15398 = ~n15394 & n15397;
  assign n15399 = ~n1297 & n15398;
  assign n15400 = ~n9958 & n15398;
  assign n15401 = ~n15399 & ~n15400;
  assign n15402 = pi17  & ~n15401;
  assign n15403 = ~pi17  & n15401;
  assign n15404 = ~n15402 & ~n15403;
  assign n15405 = ~n15393 & ~n15404;
  assign n15406 = n15393 & n15404;
  assign n15407 = ~n15405 & ~n15406;
  assign n15408 = n1611 & n8936;
  assign n15409 = pi112  & n1745;
  assign n15410 = pi114  & n1609;
  assign n15411 = pi113  & n1604;
  assign n15412 = ~n15410 & ~n15411;
  assign n15413 = ~n15409 & n15412;
  assign n15414 = ~n15408 & n15413;
  assign n15415 = pi20  & ~n15414;
  assign n15416 = pi20  & ~n15415;
  assign n15417 = ~n15414 & ~n15415;
  assign n15418 = ~n15416 & ~n15417;
  assign n15419 = ~n15236 & ~n15252;
  assign n15420 = ~n15249 & ~n15419;
  assign n15421 = ~n15418 & ~n15420;
  assign n15422 = ~n15418 & ~n15421;
  assign n15423 = ~n15420 & ~n15421;
  assign n15424 = ~n15422 & ~n15423;
  assign n15425 = n2043 & n7970;
  assign n15426 = pi109  & n2180;
  assign n15427 = pi111  & n2041;
  assign n15428 = pi110  & n2036;
  assign n15429 = ~n15427 & ~n15428;
  assign n15430 = ~n15426 & n15429;
  assign n15431 = ~n15425 & n15430;
  assign n15432 = pi23  & ~n15431;
  assign n15433 = pi23  & ~n15432;
  assign n15434 = ~n15431 & ~n15432;
  assign n15435 = ~n15433 & ~n15434;
  assign n15436 = ~n14999 & ~n15233;
  assign n15437 = n15435 & n15436;
  assign n15438 = ~n15435 & ~n15436;
  assign n15439 = ~n15437 & ~n15438;
  assign n15440 = n3034 & n6207;
  assign n15441 = pi103  & n3225;
  assign n15442 = pi105  & n3032;
  assign n15443 = pi104  & n3027;
  assign n15444 = ~n15442 & ~n15443;
  assign n15445 = ~n15441 & n15444;
  assign n15446 = ~n15440 & n15445;
  assign n15447 = pi29  & ~n15446;
  assign n15448 = pi29  & ~n15447;
  assign n15449 = ~n15446 & ~n15447;
  assign n15450 = ~n15448 & ~n15449;
  assign n15451 = ~n15013 & ~n15211;
  assign n15452 = n15450 & n15451;
  assign n15453 = ~n15450 & ~n15451;
  assign n15454 = ~n15452 & ~n15453;
  assign n15455 = n576 & n12627;
  assign n15456 = pi70  & n13004;
  assign n15457 = pi72  & n12625;
  assign n15458 = pi71  & n12620;
  assign n15459 = ~n15457 & ~n15458;
  assign n15460 = ~n15456 & n15459;
  assign n15461 = ~n15455 & n15460;
  assign n15462 = pi62  & ~n15461;
  assign n15463 = pi62  & ~n15462;
  assign n15464 = ~n15461 & ~n15462;
  assign n15465 = ~n15463 & ~n15464;
  assign n15466 = pi68  & n13835;
  assign n15467 = pi69  & ~n13434;
  assign n15468 = ~n15466 & ~n15467;
  assign n15469 = pi2  & ~n15468;
  assign n15470 = pi2  & ~n15469;
  assign n15471 = ~n15468 & ~n15469;
  assign n15472 = ~n15470 & ~n15471;
  assign n15473 = ~n15465 & ~n15472;
  assign n15474 = ~n15465 & ~n15473;
  assign n15475 = ~n15472 & ~n15473;
  assign n15476 = ~n15474 & ~n15475;
  assign n15477 = ~n15042 & ~n15046;
  assign n15478 = n15476 & n15477;
  assign n15479 = ~n15476 & ~n15477;
  assign n15480 = ~n15478 & ~n15479;
  assign n15481 = n809 & n11488;
  assign n15482 = pi73  & n11847;
  assign n15483 = pi75  & n11486;
  assign n15484 = pi74  & n11481;
  assign n15485 = ~n15483 & ~n15484;
  assign n15486 = ~n15482 & n15485;
  assign n15487 = ~n15481 & n15486;
  assign n15488 = pi59  & ~n15487;
  assign n15489 = pi59  & ~n15488;
  assign n15490 = ~n15487 & ~n15488;
  assign n15491 = ~n15489 & ~n15490;
  assign n15492 = ~n15480 & n15491;
  assign n15493 = n15480 & ~n15491;
  assign n15494 = ~n15492 & ~n15493;
  assign n15495 = ~n15052 & ~n15065;
  assign n15496 = n15494 & ~n15495;
  assign n15497 = ~n15494 & n15495;
  assign n15498 = ~n15496 & ~n15497;
  assign n15499 = n1025 & n10394;
  assign n15500 = pi76  & n10744;
  assign n15501 = pi78  & n10392;
  assign n15502 = pi77  & n10387;
  assign n15503 = ~n15501 & ~n15502;
  assign n15504 = ~n15500 & n15503;
  assign n15505 = ~n15499 & n15504;
  assign n15506 = pi56  & ~n15505;
  assign n15507 = pi56  & ~n15506;
  assign n15508 = ~n15505 & ~n15506;
  assign n15509 = ~n15507 & ~n15508;
  assign n15510 = n15498 & ~n15509;
  assign n15511 = n15498 & ~n15510;
  assign n15512 = ~n15509 & ~n15510;
  assign n15513 = ~n15511 & ~n15512;
  assign n15514 = ~n15071 & ~n15085;
  assign n15515 = ~n15513 & ~n15514;
  assign n15516 = ~n15513 & ~n15515;
  assign n15517 = ~n15514 & ~n15515;
  assign n15518 = ~n15516 & ~n15517;
  assign n15519 = n1434 & n9310;
  assign n15520 = pi79  & n9701;
  assign n15521 = pi81  & n9308;
  assign n15522 = pi80  & n9303;
  assign n15523 = ~n15521 & ~n15522;
  assign n15524 = ~n15520 & n15523;
  assign n15525 = ~n15519 & n15524;
  assign n15526 = pi53  & ~n15525;
  assign n15527 = pi53  & ~n15526;
  assign n15528 = ~n15525 & ~n15526;
  assign n15529 = ~n15527 & ~n15528;
  assign n15530 = ~n15518 & ~n15529;
  assign n15531 = ~n15518 & ~n15530;
  assign n15532 = ~n15529 & ~n15530;
  assign n15533 = ~n15531 & ~n15532;
  assign n15534 = ~n15089 & ~n15103;
  assign n15535 = n15533 & n15534;
  assign n15536 = ~n15533 & ~n15534;
  assign n15537 = ~n15535 & ~n15536;
  assign n15538 = n1834 & n8334;
  assign n15539 = pi82  & n8685;
  assign n15540 = pi84  & n8332;
  assign n15541 = pi83  & n8327;
  assign n15542 = ~n15540 & ~n15541;
  assign n15543 = ~n15539 & n15542;
  assign n15544 = ~n15538 & n15543;
  assign n15545 = pi50  & ~n15544;
  assign n15546 = pi50  & ~n15545;
  assign n15547 = ~n15544 & ~n15545;
  assign n15548 = ~n15546 & ~n15547;
  assign n15549 = ~n15537 & n15548;
  assign n15550 = n15537 & ~n15548;
  assign n15551 = ~n15549 & ~n15550;
  assign n15552 = ~n15109 & ~n15122;
  assign n15553 = n15551 & ~n15552;
  assign n15554 = ~n15551 & n15552;
  assign n15555 = ~n15553 & ~n15554;
  assign n15556 = n2288 & n7408;
  assign n15557 = pi85  & n7740;
  assign n15558 = pi87  & n7406;
  assign n15559 = pi86  & n7401;
  assign n15560 = ~n15558 & ~n15559;
  assign n15561 = ~n15557 & n15560;
  assign n15562 = ~n15556 & n15561;
  assign n15563 = pi47  & ~n15562;
  assign n15564 = pi47  & ~n15563;
  assign n15565 = ~n15562 & ~n15563;
  assign n15566 = ~n15564 & ~n15565;
  assign n15567 = n15555 & ~n15566;
  assign n15568 = n15555 & ~n15567;
  assign n15569 = ~n15566 & ~n15567;
  assign n15570 = ~n15568 & ~n15569;
  assign n15571 = ~n15128 & ~n15141;
  assign n15572 = n15570 & n15571;
  assign n15573 = ~n15570 & ~n15571;
  assign n15574 = ~n15572 & ~n15573;
  assign n15575 = n2801 & n6539;
  assign n15576 = pi88  & n6873;
  assign n15577 = pi90  & n6537;
  assign n15578 = pi89  & n6532;
  assign n15579 = ~n15577 & ~n15578;
  assign n15580 = ~n15576 & n15579;
  assign n15581 = ~n15575 & n15580;
  assign n15582 = pi44  & ~n15581;
  assign n15583 = pi44  & ~n15582;
  assign n15584 = ~n15581 & ~n15582;
  assign n15585 = ~n15583 & ~n15584;
  assign n15586 = n15574 & ~n15585;
  assign n15587 = n15574 & ~n15586;
  assign n15588 = ~n15585 & ~n15586;
  assign n15589 = ~n15587 & ~n15588;
  assign n15590 = ~n15146 & ~n15161;
  assign n15591 = n15589 & n15590;
  assign n15592 = ~n15589 & ~n15590;
  assign n15593 = ~n15591 & ~n15592;
  assign n15594 = n3371 & n5739;
  assign n15595 = pi91  & n6030;
  assign n15596 = pi93  & n5737;
  assign n15597 = pi92  & n5732;
  assign n15598 = ~n15596 & ~n15597;
  assign n15599 = ~n15595 & n15598;
  assign n15600 = ~n15594 & n15599;
  assign n15601 = pi41  & ~n15600;
  assign n15602 = pi41  & ~n15601;
  assign n15603 = ~n15600 & ~n15601;
  assign n15604 = ~n15602 & ~n15603;
  assign n15605 = n15593 & ~n15604;
  assign n15606 = n15593 & ~n15605;
  assign n15607 = ~n15604 & ~n15605;
  assign n15608 = ~n15606 & ~n15607;
  assign n15609 = ~n15167 & ~n15180;
  assign n15610 = n15608 & n15609;
  assign n15611 = ~n15608 & ~n15609;
  assign n15612 = ~n15610 & ~n15611;
  assign n15613 = n4001 & n5008;
  assign n15614 = pi94  & n5241;
  assign n15615 = pi96  & n5006;
  assign n15616 = pi95  & n5001;
  assign n15617 = ~n15615 & ~n15616;
  assign n15618 = ~n15614 & n15617;
  assign n15619 = ~n15613 & n15618;
  assign n15620 = pi38  & ~n15619;
  assign n15621 = pi38  & ~n15620;
  assign n15622 = ~n15619 & ~n15620;
  assign n15623 = ~n15621 & ~n15622;
  assign n15624 = ~n15612 & n15623;
  assign n15625 = n15612 & ~n15623;
  assign n15626 = ~n15624 & ~n15625;
  assign n15627 = ~n15186 & ~n15200;
  assign n15628 = n15626 & ~n15627;
  assign n15629 = ~n15626 & n15627;
  assign n15630 = ~n15628 & ~n15629;
  assign n15631 = n4271 & n4684;
  assign n15632 = pi97  & n4503;
  assign n15633 = pi99  & n4269;
  assign n15634 = pi98  & n4264;
  assign n15635 = ~n15633 & ~n15634;
  assign n15636 = ~n15632 & n15635;
  assign n15637 = ~n15631 & n15636;
  assign n15638 = pi35  & ~n15637;
  assign n15639 = pi35  & ~n15638;
  assign n15640 = ~n15637 & ~n15638;
  assign n15641 = ~n15639 & ~n15640;
  assign n15642 = n15630 & ~n15641;
  assign n15643 = n15630 & ~n15642;
  assign n15644 = ~n15641 & ~n15642;
  assign n15645 = ~n15643 & ~n15644;
  assign n15646 = ~n15202 & ~n15206;
  assign n15647 = pi100  & n3814;
  assign n15648 = pi102  & n3620;
  assign n15649 = pi101  & n3615;
  assign n15650 = ~n15648 & ~n15649;
  assign n15651 = ~n15647 & n15650;
  assign n15652 = ~n3622 & n15651;
  assign n15653 = ~n5413 & n15651;
  assign n15654 = ~n15652 & ~n15653;
  assign n15655 = pi32  & ~n15654;
  assign n15656 = ~pi32  & n15654;
  assign n15657 = ~n15655 & ~n15656;
  assign n15658 = ~n15646 & ~n15657;
  assign n15659 = n15646 & n15657;
  assign n15660 = ~n15658 & ~n15659;
  assign n15661 = ~n15645 & n15660;
  assign n15662 = ~n15645 & ~n15661;
  assign n15663 = n15660 & ~n15661;
  assign n15664 = ~n15662 & ~n15663;
  assign n15665 = n15454 & ~n15664;
  assign n15666 = n15454 & ~n15665;
  assign n15667 = ~n15664 & ~n15665;
  assign n15668 = ~n15666 & ~n15667;
  assign n15669 = ~n15225 & ~n15229;
  assign n15670 = pi106  & n2667;
  assign n15671 = pi108  & n2521;
  assign n15672 = pi107  & n2516;
  assign n15673 = ~n15671 & ~n15672;
  assign n15674 = ~n15670 & n15673;
  assign n15675 = ~n2523 & n15674;
  assign n15676 = ~n7060 & n15674;
  assign n15677 = ~n15675 & ~n15676;
  assign n15678 = pi26  & ~n15677;
  assign n15679 = ~pi26  & n15677;
  assign n15680 = ~n15678 & ~n15679;
  assign n15681 = ~n15669 & ~n15680;
  assign n15682 = ~n15669 & ~n15681;
  assign n15683 = ~n15680 & ~n15681;
  assign n15684 = ~n15682 & ~n15683;
  assign n15685 = ~n15668 & ~n15684;
  assign n15686 = ~n15668 & ~n15685;
  assign n15687 = ~n15684 & ~n15685;
  assign n15688 = ~n15686 & ~n15687;
  assign n15689 = n15439 & ~n15688;
  assign n15690 = n15439 & ~n15689;
  assign n15691 = ~n15688 & ~n15689;
  assign n15692 = ~n15690 & ~n15691;
  assign n15693 = ~n15424 & n15692;
  assign n15694 = n15424 & ~n15692;
  assign n15695 = ~n15693 & ~n15694;
  assign n15696 = n15407 & ~n15695;
  assign n15697 = n15407 & ~n15696;
  assign n15698 = ~n15695 & ~n15696;
  assign n15699 = ~n15697 & ~n15698;
  assign n15700 = ~n15392 & n15699;
  assign n15701 = n15392 & ~n15699;
  assign n15702 = ~n15700 & ~n15701;
  assign n15703 = n15375 & ~n15702;
  assign n15704 = n15375 & ~n15703;
  assign n15705 = ~n15702 & ~n15703;
  assign n15706 = ~n15704 & ~n15705;
  assign n15707 = ~n15295 & ~n15299;
  assign n15708 = pi124  & n537;
  assign n15709 = pi126  & n496;
  assign n15710 = pi125  & n491;
  assign n15711 = ~n15709 & ~n15710;
  assign n15712 = ~n15708 & n15711;
  assign n15713 = ~n498 & n15712;
  assign n15714 = ~n13344 & n15712;
  assign n15715 = ~n15713 & ~n15714;
  assign n15716 = pi8  & ~n15715;
  assign n15717 = ~pi8  & n15715;
  assign n15718 = ~n15716 & ~n15717;
  assign n15719 = ~n15707 & ~n15718;
  assign n15720 = ~n15707 & ~n15719;
  assign n15721 = ~n15718 & ~n15719;
  assign n15722 = ~n15720 & ~n15721;
  assign n15723 = ~n15706 & ~n15722;
  assign n15724 = n15706 & n15722;
  assign n15725 = ~n15723 & ~n15724;
  assign n15726 = ~n15360 & n15725;
  assign n15727 = n15360 & ~n15725;
  assign n15728 = ~n15726 & ~n15727;
  assign n15729 = ~n15348 & n15728;
  assign n15730 = ~n15348 & ~n15729;
  assign n15731 = n15728 & ~n15729;
  assign n15732 = ~n15730 & ~n15731;
  assign n15733 = ~n15347 & ~n15732;
  assign n15734 = n15347 & n15732;
  assign po68  = ~n15733 & ~n15734;
  assign n15736 = ~n15729 & ~n15733;
  assign n15737 = ~n15357 & ~n15726;
  assign n15738 = ~n15719 & ~n15723;
  assign n15739 = n498 & n13742;
  assign n15740 = pi125  & n537;
  assign n15741 = pi127  & n496;
  assign n15742 = pi126  & n491;
  assign n15743 = ~n15741 & ~n15742;
  assign n15744 = ~n15740 & n15743;
  assign n15745 = ~n15739 & n15744;
  assign n15746 = pi8  & ~n15745;
  assign n15747 = pi8  & ~n15746;
  assign n15748 = ~n15745 & ~n15746;
  assign n15749 = ~n15747 & ~n15748;
  assign n15750 = ~n15738 & ~n15749;
  assign n15751 = ~n15738 & ~n15750;
  assign n15752 = ~n15749 & ~n15750;
  assign n15753 = ~n15751 & ~n15752;
  assign n15754 = n687 & n12189;
  assign n15755 = pi122  & n763;
  assign n15756 = pi124  & n685;
  assign n15757 = pi123  & n680;
  assign n15758 = ~n15756 & ~n15757;
  assign n15759 = ~n15755 & n15758;
  assign n15760 = ~n15754 & n15759;
  assign n15761 = pi11  & ~n15760;
  assign n15762 = pi11  & ~n15761;
  assign n15763 = ~n15760 & ~n15761;
  assign n15764 = ~n15762 & ~n15763;
  assign n15765 = ~n15374 & ~n15703;
  assign n15766 = n15764 & n15765;
  assign n15767 = ~n15764 & ~n15765;
  assign n15768 = ~n15766 & ~n15767;
  assign n15769 = ~n15405 & ~n15696;
  assign n15770 = n1297 & n9984;
  assign n15771 = pi116  & n1366;
  assign n15772 = pi118  & n1295;
  assign n15773 = pi117  & n1290;
  assign n15774 = ~n15772 & ~n15773;
  assign n15775 = ~n15771 & n15774;
  assign n15776 = ~n15770 & n15775;
  assign n15777 = pi17  & ~n15776;
  assign n15778 = pi17  & ~n15777;
  assign n15779 = ~n15776 & ~n15777;
  assign n15780 = ~n15778 & ~n15779;
  assign n15781 = ~n15769 & ~n15780;
  assign n15782 = ~n15769 & ~n15781;
  assign n15783 = ~n15780 & ~n15781;
  assign n15784 = ~n15782 & ~n15783;
  assign n15785 = n2043 & n7997;
  assign n15786 = pi110  & n2180;
  assign n15787 = pi112  & n2041;
  assign n15788 = pi111  & n2036;
  assign n15789 = ~n15787 & ~n15788;
  assign n15790 = ~n15786 & n15789;
  assign n15791 = ~n15785 & n15790;
  assign n15792 = pi23  & ~n15791;
  assign n15793 = pi23  & ~n15792;
  assign n15794 = ~n15791 & ~n15792;
  assign n15795 = ~n15793 & ~n15794;
  assign n15796 = ~n15438 & ~n15689;
  assign n15797 = n15795 & n15796;
  assign n15798 = ~n15795 & ~n15796;
  assign n15799 = ~n15797 & ~n15798;
  assign n15800 = ~n15681 & ~n15685;
  assign n15801 = n2523 & n7349;
  assign n15802 = pi107  & n2667;
  assign n15803 = pi109  & n2521;
  assign n15804 = pi108  & n2516;
  assign n15805 = ~n15803 & ~n15804;
  assign n15806 = ~n15802 & n15805;
  assign n15807 = ~n15801 & n15806;
  assign n15808 = pi26  & ~n15807;
  assign n15809 = pi26  & ~n15808;
  assign n15810 = ~n15807 & ~n15808;
  assign n15811 = ~n15809 & ~n15810;
  assign n15812 = ~n15800 & ~n15811;
  assign n15813 = ~n15800 & ~n15812;
  assign n15814 = ~n15811 & ~n15812;
  assign n15815 = ~n15813 & ~n15814;
  assign n15816 = n3034 & n6477;
  assign n15817 = pi104  & n3225;
  assign n15818 = pi106  & n3032;
  assign n15819 = pi105  & n3027;
  assign n15820 = ~n15818 & ~n15819;
  assign n15821 = ~n15817 & n15820;
  assign n15822 = ~n15816 & n15821;
  assign n15823 = pi29  & ~n15822;
  assign n15824 = pi29  & ~n15823;
  assign n15825 = ~n15822 & ~n15823;
  assign n15826 = ~n15824 & ~n15825;
  assign n15827 = ~n15453 & ~n15665;
  assign n15828 = n15826 & n15827;
  assign n15829 = ~n15826 & ~n15827;
  assign n15830 = ~n15828 & ~n15829;
  assign n15831 = ~n15628 & ~n15642;
  assign n15832 = ~n15611 & ~n15625;
  assign n15833 = ~n15592 & ~n15605;
  assign n15834 = ~n15553 & ~n15567;
  assign n15835 = ~n15536 & ~n15550;
  assign n15836 = ~n15479 & ~n15493;
  assign n15837 = n891 & n11488;
  assign n15838 = pi74  & n11847;
  assign n15839 = pi76  & n11486;
  assign n15840 = pi75  & n11481;
  assign n15841 = ~n15839 & ~n15840;
  assign n15842 = ~n15838 & n15841;
  assign n15843 = ~n15837 & n15842;
  assign n15844 = pi59  & ~n15843;
  assign n15845 = pi59  & ~n15844;
  assign n15846 = ~n15843 & ~n15844;
  assign n15847 = ~n15845 & ~n15846;
  assign n15848 = ~n15469 & ~n15473;
  assign n15849 = pi69  & n13835;
  assign n15850 = pi70  & ~n13434;
  assign n15851 = ~n15849 & ~n15850;
  assign n15852 = pi2  & ~pi5 ;
  assign n15853 = ~pi2  & pi5 ;
  assign n15854 = ~n15852 & ~n15853;
  assign n15855 = ~n15851 & ~n15854;
  assign n15856 = n15851 & n15854;
  assign n15857 = ~n15855 & ~n15856;
  assign n15858 = n15848 & ~n15857;
  assign n15859 = ~n15848 & n15857;
  assign n15860 = ~n15858 & ~n15859;
  assign n15861 = n642 & n12627;
  assign n15862 = pi71  & n13004;
  assign n15863 = pi73  & n12625;
  assign n15864 = pi72  & n12620;
  assign n15865 = ~n15863 & ~n15864;
  assign n15866 = ~n15862 & n15865;
  assign n15867 = ~n15861 & n15866;
  assign n15868 = pi62  & ~n15867;
  assign n15869 = pi62  & ~n15868;
  assign n15870 = ~n15867 & ~n15868;
  assign n15871 = ~n15869 & ~n15870;
  assign n15872 = ~n15860 & n15871;
  assign n15873 = n15860 & ~n15871;
  assign n15874 = ~n15872 & ~n15873;
  assign n15875 = ~n15847 & n15874;
  assign n15876 = ~n15847 & ~n15875;
  assign n15877 = n15874 & ~n15875;
  assign n15878 = ~n15876 & ~n15877;
  assign n15879 = ~n15836 & ~n15878;
  assign n15880 = ~n15836 & ~n15879;
  assign n15881 = ~n15878 & ~n15879;
  assign n15882 = ~n15880 & ~n15881;
  assign n15883 = n1122 & n10394;
  assign n15884 = pi77  & n10744;
  assign n15885 = pi79  & n10392;
  assign n15886 = pi78  & n10387;
  assign n15887 = ~n15885 & ~n15886;
  assign n15888 = ~n15884 & n15887;
  assign n15889 = ~n15883 & n15888;
  assign n15890 = pi56  & ~n15889;
  assign n15891 = pi56  & ~n15890;
  assign n15892 = ~n15889 & ~n15890;
  assign n15893 = ~n15891 & ~n15892;
  assign n15894 = ~n15882 & ~n15893;
  assign n15895 = ~n15882 & ~n15894;
  assign n15896 = ~n15893 & ~n15894;
  assign n15897 = ~n15895 & ~n15896;
  assign n15898 = ~n15496 & ~n15510;
  assign n15899 = n15897 & n15898;
  assign n15900 = ~n15897 & ~n15898;
  assign n15901 = ~n15899 & ~n15900;
  assign n15902 = n1554 & n9310;
  assign n15903 = pi80  & n9701;
  assign n15904 = pi82  & n9308;
  assign n15905 = pi81  & n9303;
  assign n15906 = ~n15904 & ~n15905;
  assign n15907 = ~n15903 & n15906;
  assign n15908 = ~n15902 & n15907;
  assign n15909 = pi53  & ~n15908;
  assign n15910 = pi53  & ~n15909;
  assign n15911 = ~n15908 & ~n15909;
  assign n15912 = ~n15910 & ~n15911;
  assign n15913 = n15901 & ~n15912;
  assign n15914 = n15901 & ~n15913;
  assign n15915 = ~n15912 & ~n15913;
  assign n15916 = ~n15914 & ~n15915;
  assign n15917 = ~n15515 & ~n15530;
  assign n15918 = n15916 & n15917;
  assign n15919 = ~n15916 & ~n15917;
  assign n15920 = ~n15918 & ~n15919;
  assign n15921 = n1972 & n8334;
  assign n15922 = pi83  & n8685;
  assign n15923 = pi85  & n8332;
  assign n15924 = pi84  & n8327;
  assign n15925 = ~n15923 & ~n15924;
  assign n15926 = ~n15922 & n15925;
  assign n15927 = ~n15921 & n15926;
  assign n15928 = pi50  & ~n15927;
  assign n15929 = pi50  & ~n15928;
  assign n15930 = ~n15927 & ~n15928;
  assign n15931 = ~n15929 & ~n15930;
  assign n15932 = n15920 & ~n15931;
  assign n15933 = n15920 & ~n15932;
  assign n15934 = ~n15931 & ~n15932;
  assign n15935 = ~n15933 & ~n15934;
  assign n15936 = ~n15835 & n15935;
  assign n15937 = n15835 & ~n15935;
  assign n15938 = ~n15936 & ~n15937;
  assign n15939 = n2446 & n7408;
  assign n15940 = pi86  & n7740;
  assign n15941 = pi88  & n7406;
  assign n15942 = pi87  & n7401;
  assign n15943 = ~n15941 & ~n15942;
  assign n15944 = ~n15940 & n15943;
  assign n15945 = ~n15939 & n15944;
  assign n15946 = pi47  & ~n15945;
  assign n15947 = pi47  & ~n15946;
  assign n15948 = ~n15945 & ~n15946;
  assign n15949 = ~n15947 & ~n15948;
  assign n15950 = ~n15938 & ~n15949;
  assign n15951 = n15938 & n15949;
  assign n15952 = ~n15950 & ~n15951;
  assign n15953 = n15834 & ~n15952;
  assign n15954 = ~n15834 & n15952;
  assign n15955 = ~n15953 & ~n15954;
  assign n15956 = n2978 & n6539;
  assign n15957 = pi89  & n6873;
  assign n15958 = pi91  & n6537;
  assign n15959 = pi90  & n6532;
  assign n15960 = ~n15958 & ~n15959;
  assign n15961 = ~n15957 & n15960;
  assign n15962 = ~n15956 & n15961;
  assign n15963 = pi44  & ~n15962;
  assign n15964 = pi44  & ~n15963;
  assign n15965 = ~n15962 & ~n15963;
  assign n15966 = ~n15964 & ~n15965;
  assign n15967 = n15955 & ~n15966;
  assign n15968 = n15955 & ~n15967;
  assign n15969 = ~n15966 & ~n15967;
  assign n15970 = ~n15968 & ~n15969;
  assign n15971 = ~n15573 & ~n15586;
  assign n15972 = n15970 & n15971;
  assign n15973 = ~n15970 & ~n15971;
  assign n15974 = ~n15972 & ~n15973;
  assign n15975 = n3565 & n5739;
  assign n15976 = pi92  & n6030;
  assign n15977 = pi94  & n5737;
  assign n15978 = pi93  & n5732;
  assign n15979 = ~n15977 & ~n15978;
  assign n15980 = ~n15976 & n15979;
  assign n15981 = ~n15975 & n15980;
  assign n15982 = pi41  & ~n15981;
  assign n15983 = pi41  & ~n15982;
  assign n15984 = ~n15981 & ~n15982;
  assign n15985 = ~n15983 & ~n15984;
  assign n15986 = ~n15974 & n15985;
  assign n15987 = n15974 & ~n15985;
  assign n15988 = ~n15833 & ~n15986;
  assign n15989 = ~n15987 & n15988;
  assign n15990 = ~n15833 & ~n15989;
  assign n15991 = ~n15987 & ~n15989;
  assign n15992 = ~n15986 & n15991;
  assign n15993 = ~n15990 & ~n15992;
  assign n15994 = n4211 & n5008;
  assign n15995 = pi95  & n5241;
  assign n15996 = pi97  & n5006;
  assign n15997 = pi96  & n5001;
  assign n15998 = ~n15996 & ~n15997;
  assign n15999 = ~n15995 & n15998;
  assign n16000 = ~n15994 & n15999;
  assign n16001 = pi38  & ~n16000;
  assign n16002 = pi38  & ~n16001;
  assign n16003 = ~n16000 & ~n16001;
  assign n16004 = ~n16002 & ~n16003;
  assign n16005 = ~n15993 & ~n16004;
  assign n16006 = ~n15993 & ~n16005;
  assign n16007 = ~n16004 & ~n16005;
  assign n16008 = ~n16006 & ~n16007;
  assign n16009 = ~n15832 & n16008;
  assign n16010 = n15832 & ~n16008;
  assign n16011 = ~n16009 & ~n16010;
  assign n16012 = n4271 & n4910;
  assign n16013 = pi98  & n4503;
  assign n16014 = pi100  & n4269;
  assign n16015 = pi99  & n4264;
  assign n16016 = ~n16014 & ~n16015;
  assign n16017 = ~n16013 & n16016;
  assign n16018 = ~n16012 & n16017;
  assign n16019 = pi35  & ~n16018;
  assign n16020 = pi35  & ~n16019;
  assign n16021 = ~n16018 & ~n16019;
  assign n16022 = ~n16020 & ~n16021;
  assign n16023 = ~n16011 & ~n16022;
  assign n16024 = n16011 & n16022;
  assign n16025 = ~n16023 & ~n16024;
  assign n16026 = n15831 & ~n16025;
  assign n16027 = ~n15831 & n16025;
  assign n16028 = ~n16026 & ~n16027;
  assign n16029 = n3622 & n5664;
  assign n16030 = pi101  & n3814;
  assign n16031 = pi103  & n3620;
  assign n16032 = pi102  & n3615;
  assign n16033 = ~n16031 & ~n16032;
  assign n16034 = ~n16030 & n16033;
  assign n16035 = ~n16029 & n16034;
  assign n16036 = pi32  & ~n16035;
  assign n16037 = pi32  & ~n16036;
  assign n16038 = ~n16035 & ~n16036;
  assign n16039 = ~n16037 & ~n16038;
  assign n16040 = ~n15658 & ~n15661;
  assign n16041 = n16039 & n16040;
  assign n16042 = ~n16039 & ~n16040;
  assign n16043 = ~n16041 & ~n16042;
  assign n16044 = n16028 & n16043;
  assign n16045 = ~n16028 & ~n16043;
  assign n16046 = ~n16044 & ~n16045;
  assign n16047 = n15830 & n16046;
  assign n16048 = ~n15830 & ~n16046;
  assign n16049 = ~n16047 & ~n16048;
  assign n16050 = ~n15815 & ~n16049;
  assign n16051 = n15815 & n16049;
  assign n16052 = ~n16050 & ~n16051;
  assign n16053 = n15799 & ~n16052;
  assign n16054 = n15799 & ~n16053;
  assign n16055 = ~n16052 & ~n16053;
  assign n16056 = ~n16054 & ~n16055;
  assign n16057 = n1611 & n8963;
  assign n16058 = pi113  & n1745;
  assign n16059 = pi115  & n1609;
  assign n16060 = pi114  & n1604;
  assign n16061 = ~n16059 & ~n16060;
  assign n16062 = ~n16058 & n16061;
  assign n16063 = ~n16057 & n16062;
  assign n16064 = pi20  & ~n16063;
  assign n16065 = pi20  & ~n16064;
  assign n16066 = ~n16063 & ~n16064;
  assign n16067 = ~n16065 & ~n16066;
  assign n16068 = ~n15424 & ~n15692;
  assign n16069 = ~n15421 & ~n16068;
  assign n16070 = ~n16067 & ~n16069;
  assign n16071 = n16067 & n16069;
  assign n16072 = ~n16070 & ~n16071;
  assign n16073 = ~n16056 & n16072;
  assign n16074 = ~n16056 & ~n16073;
  assign n16075 = n16072 & ~n16073;
  assign n16076 = ~n16074 & ~n16075;
  assign n16077 = ~n15784 & ~n16076;
  assign n16078 = ~n15784 & ~n16077;
  assign n16079 = ~n16076 & ~n16077;
  assign n16080 = ~n16078 & ~n16079;
  assign n16081 = n938 & n11389;
  assign n16082 = pi119  & n1052;
  assign n16083 = pi121  & n936;
  assign n16084 = pi120  & n931;
  assign n16085 = ~n16083 & ~n16084;
  assign n16086 = ~n16082 & n16085;
  assign n16087 = ~n16081 & n16086;
  assign n16088 = pi14  & ~n16087;
  assign n16089 = pi14  & ~n16088;
  assign n16090 = ~n16087 & ~n16088;
  assign n16091 = ~n16089 & ~n16090;
  assign n16092 = ~n15392 & ~n15699;
  assign n16093 = ~n15389 & ~n16092;
  assign n16094 = ~n16091 & ~n16093;
  assign n16095 = n16091 & n16093;
  assign n16096 = ~n16094 & ~n16095;
  assign n16097 = ~n16080 & n16096;
  assign n16098 = ~n16080 & ~n16097;
  assign n16099 = n16096 & ~n16097;
  assign n16100 = ~n16098 & ~n16099;
  assign n16101 = n15768 & ~n16100;
  assign n16102 = n15768 & ~n16101;
  assign n16103 = ~n16100 & ~n16101;
  assign n16104 = ~n16102 & ~n16103;
  assign n16105 = ~n15753 & n16104;
  assign n16106 = n15753 & ~n16104;
  assign n16107 = ~n16105 & ~n16106;
  assign n16108 = ~n15737 & ~n16107;
  assign n16109 = n15737 & n16107;
  assign n16110 = ~n16108 & ~n16109;
  assign n16111 = ~n15736 & n16110;
  assign n16112 = n15736 & ~n16110;
  assign po69  = ~n16111 & ~n16112;
  assign n16114 = ~n15767 & ~n16101;
  assign n16115 = pi126  & n537;
  assign n16116 = pi127  & n491;
  assign n16117 = ~n16115 & ~n16116;
  assign n16118 = ~n498 & n16117;
  assign n16119 = n13773 & n16117;
  assign n16120 = ~n16118 & ~n16119;
  assign n16121 = pi8  & ~n16120;
  assign n16122 = ~pi8  & n16120;
  assign n16123 = ~n16121 & ~n16122;
  assign n16124 = ~n16114 & ~n16123;
  assign n16125 = n16114 & n16123;
  assign n16126 = ~n16124 & ~n16125;
  assign n16127 = n687 & n12943;
  assign n16128 = pi123  & n763;
  assign n16129 = pi125  & n685;
  assign n16130 = pi124  & n680;
  assign n16131 = ~n16129 & ~n16130;
  assign n16132 = ~n16128 & n16131;
  assign n16133 = ~n16127 & n16132;
  assign n16134 = pi11  & ~n16133;
  assign n16135 = pi11  & ~n16134;
  assign n16136 = ~n16133 & ~n16134;
  assign n16137 = ~n16135 & ~n16136;
  assign n16138 = ~n16094 & ~n16097;
  assign n16139 = n16137 & n16138;
  assign n16140 = ~n16137 & ~n16138;
  assign n16141 = ~n16139 & ~n16140;
  assign n16142 = ~n15781 & ~n16077;
  assign n16143 = pi120  & n1052;
  assign n16144 = pi122  & n936;
  assign n16145 = pi121  & n931;
  assign n16146 = ~n16144 & ~n16145;
  assign n16147 = ~n16143 & n16146;
  assign n16148 = ~n938 & n16147;
  assign n16149 = ~n11778 & n16147;
  assign n16150 = ~n16148 & ~n16149;
  assign n16151 = pi14  & ~n16150;
  assign n16152 = ~pi14  & n16150;
  assign n16153 = ~n16151 & ~n16152;
  assign n16154 = ~n16142 & ~n16153;
  assign n16155 = n16142 & n16153;
  assign n16156 = ~n16154 & ~n16155;
  assign n16157 = n1297 & n10667;
  assign n16158 = pi117  & n1366;
  assign n16159 = pi119  & n1295;
  assign n16160 = pi118  & n1290;
  assign n16161 = ~n16159 & ~n16160;
  assign n16162 = ~n16158 & n16161;
  assign n16163 = ~n16157 & n16162;
  assign n16164 = pi17  & ~n16163;
  assign n16165 = pi17  & ~n16164;
  assign n16166 = ~n16163 & ~n16164;
  assign n16167 = ~n16165 & ~n16166;
  assign n16168 = ~n16070 & ~n16073;
  assign n16169 = n16167 & n16168;
  assign n16170 = ~n16167 & ~n16168;
  assign n16171 = ~n16169 & ~n16170;
  assign n16172 = n1611 & n9614;
  assign n16173 = pi114  & n1745;
  assign n16174 = pi116  & n1609;
  assign n16175 = pi115  & n1604;
  assign n16176 = ~n16174 & ~n16175;
  assign n16177 = ~n16173 & n16176;
  assign n16178 = ~n16172 & n16177;
  assign n16179 = pi20  & ~n16178;
  assign n16180 = pi20  & ~n16179;
  assign n16181 = ~n16178 & ~n16179;
  assign n16182 = ~n16180 & ~n16181;
  assign n16183 = ~n15798 & ~n16053;
  assign n16184 = n16182 & n16183;
  assign n16185 = ~n16182 & ~n16183;
  assign n16186 = ~n16184 & ~n16185;
  assign n16187 = n2043 & n8612;
  assign n16188 = pi111  & n2180;
  assign n16189 = pi113  & n2041;
  assign n16190 = pi112  & n2036;
  assign n16191 = ~n16189 & ~n16190;
  assign n16192 = ~n16188 & n16191;
  assign n16193 = ~n16187 & n16192;
  assign n16194 = pi23  & ~n16193;
  assign n16195 = pi23  & ~n16194;
  assign n16196 = ~n16193 & ~n16194;
  assign n16197 = ~n16195 & ~n16196;
  assign n16198 = ~n15815 & n16049;
  assign n16199 = ~n15812 & ~n16198;
  assign n16200 = ~n16197 & ~n16199;
  assign n16201 = ~n16197 & ~n16200;
  assign n16202 = ~n16199 & ~n16200;
  assign n16203 = ~n16201 & ~n16202;
  assign n16204 = ~n15829 & ~n16047;
  assign n16205 = pi108  & n2667;
  assign n16206 = pi110  & n2521;
  assign n16207 = pi109  & n2516;
  assign n16208 = ~n16206 & ~n16207;
  assign n16209 = ~n16205 & n16208;
  assign n16210 = ~n2523 & n16209;
  assign n16211 = ~n7665 & n16209;
  assign n16212 = ~n16210 & ~n16211;
  assign n16213 = pi26  & ~n16212;
  assign n16214 = ~pi26  & n16212;
  assign n16215 = ~n16213 & ~n16214;
  assign n16216 = ~n16204 & ~n16215;
  assign n16217 = n16204 & n16215;
  assign n16218 = ~n16216 & ~n16217;
  assign n16219 = n3034 & n6775;
  assign n16220 = pi105  & n3225;
  assign n16221 = pi107  & n3032;
  assign n16222 = pi106  & n3027;
  assign n16223 = ~n16221 & ~n16222;
  assign n16224 = ~n16220 & n16223;
  assign n16225 = ~n16219 & n16224;
  assign n16226 = pi29  & ~n16225;
  assign n16227 = pi29  & ~n16226;
  assign n16228 = ~n16225 & ~n16226;
  assign n16229 = ~n16227 & ~n16228;
  assign n16230 = ~n16042 & ~n16044;
  assign n16231 = ~n16229 & ~n16230;
  assign n16232 = ~n16229 & ~n16231;
  assign n16233 = ~n16230 & ~n16231;
  assign n16234 = ~n16232 & ~n16233;
  assign n16235 = n3622 & n5943;
  assign n16236 = pi102  & n3814;
  assign n16237 = pi104  & n3620;
  assign n16238 = pi103  & n3615;
  assign n16239 = ~n16237 & ~n16238;
  assign n16240 = ~n16236 & n16239;
  assign n16241 = ~n16235 & n16240;
  assign n16242 = pi32  & ~n16241;
  assign n16243 = pi32  & ~n16242;
  assign n16244 = ~n16241 & ~n16242;
  assign n16245 = ~n16243 & ~n16244;
  assign n16246 = ~n16023 & ~n16027;
  assign n16247 = n16245 & n16246;
  assign n16248 = ~n16245 & ~n16246;
  assign n16249 = ~n16247 & ~n16248;
  assign n16250 = n4271 & n5169;
  assign n16251 = pi99  & n4503;
  assign n16252 = pi101  & n4269;
  assign n16253 = pi100  & n4264;
  assign n16254 = ~n16252 & ~n16253;
  assign n16255 = ~n16251 & n16254;
  assign n16256 = ~n16250 & n16255;
  assign n16257 = pi35  & ~n16256;
  assign n16258 = pi35  & ~n16257;
  assign n16259 = ~n16256 & ~n16257;
  assign n16260 = ~n16258 & ~n16259;
  assign n16261 = ~n15832 & ~n16008;
  assign n16262 = ~n16005 & ~n16261;
  assign n16263 = n4454 & n5008;
  assign n16264 = pi96  & n5241;
  assign n16265 = pi98  & n5006;
  assign n16266 = pi97  & n5001;
  assign n16267 = ~n16265 & ~n16266;
  assign n16268 = ~n16264 & n16267;
  assign n16269 = ~n16263 & n16268;
  assign n16270 = pi38  & ~n16269;
  assign n16271 = pi38  & ~n16270;
  assign n16272 = ~n16269 & ~n16270;
  assign n16273 = ~n16271 & ~n16272;
  assign n16274 = ~n15859 & ~n15873;
  assign n16275 = ~pi2  & ~pi5 ;
  assign n16276 = ~n15855 & ~n16275;
  assign n16277 = pi70  & n13835;
  assign n16278 = pi71  & ~n13434;
  assign n16279 = ~n16277 & ~n16278;
  assign n16280 = ~n16276 & n16279;
  assign n16281 = n16276 & ~n16279;
  assign n16282 = ~n16280 & ~n16281;
  assign n16283 = pi72  & n13004;
  assign n16284 = pi74  & n12625;
  assign n16285 = pi73  & n12620;
  assign n16286 = ~n16284 & ~n16285;
  assign n16287 = ~n16283 & n16286;
  assign n16288 = ~n12627 & n16287;
  assign n16289 = ~n729 & n16287;
  assign n16290 = ~n16288 & ~n16289;
  assign n16291 = pi62  & ~n16290;
  assign n16292 = ~pi62  & n16290;
  assign n16293 = ~n16291 & ~n16292;
  assign n16294 = n16282 & ~n16293;
  assign n16295 = ~n16282 & n16293;
  assign n16296 = ~n16294 & ~n16295;
  assign n16297 = ~n16274 & n16296;
  assign n16298 = n16274 & ~n16296;
  assign n16299 = ~n16297 & ~n16298;
  assign n16300 = n999 & n11488;
  assign n16301 = pi75  & n11847;
  assign n16302 = pi77  & n11486;
  assign n16303 = pi76  & n11481;
  assign n16304 = ~n16302 & ~n16303;
  assign n16305 = ~n16301 & n16304;
  assign n16306 = ~n16300 & n16305;
  assign n16307 = pi59  & ~n16306;
  assign n16308 = pi59  & ~n16307;
  assign n16309 = ~n16306 & ~n16307;
  assign n16310 = ~n16308 & ~n16309;
  assign n16311 = n16299 & ~n16310;
  assign n16312 = n16299 & ~n16311;
  assign n16313 = ~n16310 & ~n16311;
  assign n16314 = ~n16312 & ~n16313;
  assign n16315 = ~n15875 & ~n15879;
  assign n16316 = n16314 & n16315;
  assign n16317 = ~n16314 & ~n16315;
  assign n16318 = ~n16316 & ~n16317;
  assign n16319 = n1225 & n10394;
  assign n16320 = pi78  & n10744;
  assign n16321 = pi80  & n10392;
  assign n16322 = pi79  & n10387;
  assign n16323 = ~n16321 & ~n16322;
  assign n16324 = ~n16320 & n16323;
  assign n16325 = ~n16319 & n16324;
  assign n16326 = pi56  & ~n16325;
  assign n16327 = pi56  & ~n16326;
  assign n16328 = ~n16325 & ~n16326;
  assign n16329 = ~n16327 & ~n16328;
  assign n16330 = n16318 & ~n16329;
  assign n16331 = n16318 & ~n16330;
  assign n16332 = ~n16329 & ~n16330;
  assign n16333 = ~n16331 & ~n16332;
  assign n16334 = ~n15894 & ~n15900;
  assign n16335 = n16333 & n16334;
  assign n16336 = ~n16333 & ~n16334;
  assign n16337 = ~n16335 & ~n16336;
  assign n16338 = n1696 & n9310;
  assign n16339 = pi81  & n9701;
  assign n16340 = pi83  & n9308;
  assign n16341 = pi82  & n9303;
  assign n16342 = ~n16340 & ~n16341;
  assign n16343 = ~n16339 & n16342;
  assign n16344 = ~n16338 & n16343;
  assign n16345 = pi53  & ~n16344;
  assign n16346 = pi53  & ~n16345;
  assign n16347 = ~n16344 & ~n16345;
  assign n16348 = ~n16346 & ~n16347;
  assign n16349 = n16337 & ~n16348;
  assign n16350 = n16337 & ~n16349;
  assign n16351 = ~n16348 & ~n16349;
  assign n16352 = ~n16350 & ~n16351;
  assign n16353 = ~n15913 & ~n15919;
  assign n16354 = n16352 & n16353;
  assign n16355 = ~n16352 & ~n16353;
  assign n16356 = ~n16354 & ~n16355;
  assign n16357 = n2133 & n8334;
  assign n16358 = pi84  & n8685;
  assign n16359 = pi86  & n8332;
  assign n16360 = pi85  & n8327;
  assign n16361 = ~n16359 & ~n16360;
  assign n16362 = ~n16358 & n16361;
  assign n16363 = ~n16357 & n16362;
  assign n16364 = pi50  & ~n16363;
  assign n16365 = pi50  & ~n16364;
  assign n16366 = ~n16363 & ~n16364;
  assign n16367 = ~n16365 & ~n16366;
  assign n16368 = n16356 & ~n16367;
  assign n16369 = n16356 & ~n16368;
  assign n16370 = ~n16367 & ~n16368;
  assign n16371 = ~n16369 & ~n16370;
  assign n16372 = ~n15835 & ~n15935;
  assign n16373 = ~n15932 & ~n16372;
  assign n16374 = n16371 & n16373;
  assign n16375 = ~n16371 & ~n16373;
  assign n16376 = ~n16374 & ~n16375;
  assign n16377 = n2473 & n7408;
  assign n16378 = pi87  & n7740;
  assign n16379 = pi89  & n7406;
  assign n16380 = pi88  & n7401;
  assign n16381 = ~n16379 & ~n16380;
  assign n16382 = ~n16378 & n16381;
  assign n16383 = ~n16377 & n16382;
  assign n16384 = pi47  & ~n16383;
  assign n16385 = pi47  & ~n16384;
  assign n16386 = ~n16383 & ~n16384;
  assign n16387 = ~n16385 & ~n16386;
  assign n16388 = n16376 & ~n16387;
  assign n16389 = n16376 & ~n16388;
  assign n16390 = ~n16387 & ~n16388;
  assign n16391 = ~n16389 & ~n16390;
  assign n16392 = ~n15950 & ~n15954;
  assign n16393 = n16391 & n16392;
  assign n16394 = ~n16391 & ~n16392;
  assign n16395 = ~n16393 & ~n16394;
  assign n16396 = n3177 & n6539;
  assign n16397 = pi90  & n6873;
  assign n16398 = pi92  & n6537;
  assign n16399 = pi91  & n6532;
  assign n16400 = ~n16398 & ~n16399;
  assign n16401 = ~n16397 & n16400;
  assign n16402 = ~n16396 & n16401;
  assign n16403 = pi44  & ~n16402;
  assign n16404 = pi44  & ~n16403;
  assign n16405 = ~n16402 & ~n16403;
  assign n16406 = ~n16404 & ~n16405;
  assign n16407 = n16395 & ~n16406;
  assign n16408 = n16395 & ~n16407;
  assign n16409 = ~n16406 & ~n16407;
  assign n16410 = ~n16408 & ~n16409;
  assign n16411 = ~n15967 & ~n15973;
  assign n16412 = n16410 & n16411;
  assign n16413 = ~n16410 & ~n16411;
  assign n16414 = ~n16412 & ~n16413;
  assign n16415 = n3784 & n5739;
  assign n16416 = pi93  & n6030;
  assign n16417 = pi95  & n5737;
  assign n16418 = pi94  & n5732;
  assign n16419 = ~n16417 & ~n16418;
  assign n16420 = ~n16416 & n16419;
  assign n16421 = ~n16415 & n16420;
  assign n16422 = pi41  & ~n16421;
  assign n16423 = pi41  & ~n16422;
  assign n16424 = ~n16421 & ~n16422;
  assign n16425 = ~n16423 & ~n16424;
  assign n16426 = ~n16414 & n16425;
  assign n16427 = n16414 & ~n16425;
  assign n16428 = ~n16426 & ~n16427;
  assign n16429 = ~n15991 & n16428;
  assign n16430 = n15991 & ~n16428;
  assign n16431 = ~n16429 & ~n16430;
  assign n16432 = ~n16273 & n16431;
  assign n16433 = n16273 & ~n16431;
  assign n16434 = ~n16432 & ~n16433;
  assign n16435 = ~n16262 & n16434;
  assign n16436 = n16262 & ~n16434;
  assign n16437 = ~n16435 & ~n16436;
  assign n16438 = ~n16260 & n16437;
  assign n16439 = ~n16260 & ~n16438;
  assign n16440 = n16437 & ~n16438;
  assign n16441 = ~n16439 & ~n16440;
  assign n16442 = n16249 & ~n16441;
  assign n16443 = n16249 & ~n16442;
  assign n16444 = ~n16441 & ~n16442;
  assign n16445 = ~n16443 & ~n16444;
  assign n16446 = ~n16234 & n16445;
  assign n16447 = n16234 & ~n16445;
  assign n16448 = ~n16446 & ~n16447;
  assign n16449 = n16218 & ~n16448;
  assign n16450 = n16218 & ~n16449;
  assign n16451 = ~n16448 & ~n16449;
  assign n16452 = ~n16450 & ~n16451;
  assign n16453 = ~n16203 & n16452;
  assign n16454 = n16203 & ~n16452;
  assign n16455 = ~n16453 & ~n16454;
  assign n16456 = n16186 & ~n16455;
  assign n16457 = n16186 & ~n16456;
  assign n16458 = ~n16455 & ~n16456;
  assign n16459 = ~n16457 & ~n16458;
  assign n16460 = n16171 & ~n16459;
  assign n16461 = ~n16171 & n16459;
  assign n16462 = ~n16460 & ~n16461;
  assign n16463 = n16156 & n16462;
  assign n16464 = n16156 & ~n16463;
  assign n16465 = n16462 & ~n16463;
  assign n16466 = ~n16464 & ~n16465;
  assign n16467 = n16141 & ~n16466;
  assign n16468 = ~n16141 & n16466;
  assign n16469 = ~n16467 & ~n16468;
  assign n16470 = n16126 & n16469;
  assign n16471 = n16126 & ~n16470;
  assign n16472 = n16469 & ~n16470;
  assign n16473 = ~n16471 & ~n16472;
  assign n16474 = ~n15753 & ~n16104;
  assign n16475 = ~n15750 & ~n16474;
  assign n16476 = ~n16473 & ~n16475;
  assign n16477 = ~n16473 & ~n16476;
  assign n16478 = ~n16475 & ~n16476;
  assign n16479 = ~n16477 & ~n16478;
  assign n16480 = ~n16108 & ~n16111;
  assign n16481 = ~n16479 & ~n16480;
  assign n16482 = n16479 & n16480;
  assign po70  = ~n16481 & ~n16482;
  assign n16484 = ~n16476 & ~n16481;
  assign n16485 = ~n16124 & ~n16470;
  assign n16486 = ~n16140 & ~n16467;
  assign n16487 = pi127  & n537;
  assign n16488 = n498 & n13770;
  assign n16489 = ~n16487 & ~n16488;
  assign n16490 = pi8  & ~n16489;
  assign n16491 = pi8  & ~n16490;
  assign n16492 = ~n16489 & ~n16490;
  assign n16493 = ~n16491 & ~n16492;
  assign n16494 = ~n16486 & ~n16493;
  assign n16495 = ~n16486 & ~n16494;
  assign n16496 = ~n16493 & ~n16494;
  assign n16497 = ~n16495 & ~n16496;
  assign n16498 = n1297 & n11028;
  assign n16499 = pi118  & n1366;
  assign n16500 = pi120  & n1295;
  assign n16501 = pi119  & n1290;
  assign n16502 = ~n16500 & ~n16501;
  assign n16503 = ~n16499 & n16502;
  assign n16504 = ~n16498 & n16503;
  assign n16505 = pi17  & ~n16504;
  assign n16506 = pi17  & ~n16505;
  assign n16507 = ~n16504 & ~n16505;
  assign n16508 = ~n16506 & ~n16507;
  assign n16509 = ~n16185 & ~n16456;
  assign n16510 = n16508 & n16509;
  assign n16511 = ~n16508 & ~n16509;
  assign n16512 = ~n16510 & ~n16511;
  assign n16513 = n2043 & n8936;
  assign n16514 = pi112  & n2180;
  assign n16515 = pi114  & n2041;
  assign n16516 = pi113  & n2036;
  assign n16517 = ~n16515 & ~n16516;
  assign n16518 = ~n16514 & n16517;
  assign n16519 = ~n16513 & n16518;
  assign n16520 = pi23  & ~n16519;
  assign n16521 = pi23  & ~n16520;
  assign n16522 = ~n16519 & ~n16520;
  assign n16523 = ~n16521 & ~n16522;
  assign n16524 = ~n16216 & ~n16449;
  assign n16525 = n16523 & n16524;
  assign n16526 = ~n16523 & ~n16524;
  assign n16527 = ~n16525 & ~n16526;
  assign n16528 = n2523 & n7970;
  assign n16529 = pi109  & n2667;
  assign n16530 = pi111  & n2521;
  assign n16531 = pi110  & n2516;
  assign n16532 = ~n16530 & ~n16531;
  assign n16533 = ~n16529 & n16532;
  assign n16534 = ~n16528 & n16533;
  assign n16535 = pi26  & ~n16534;
  assign n16536 = pi26  & ~n16535;
  assign n16537 = ~n16534 & ~n16535;
  assign n16538 = ~n16536 & ~n16537;
  assign n16539 = ~n16234 & ~n16445;
  assign n16540 = ~n16231 & ~n16539;
  assign n16541 = ~n16538 & ~n16540;
  assign n16542 = ~n16538 & ~n16541;
  assign n16543 = ~n16540 & ~n16541;
  assign n16544 = ~n16542 & ~n16543;
  assign n16545 = n3622 & n6207;
  assign n16546 = pi103  & n3814;
  assign n16547 = pi105  & n3620;
  assign n16548 = pi104  & n3615;
  assign n16549 = ~n16547 & ~n16548;
  assign n16550 = ~n16546 & n16549;
  assign n16551 = ~n16545 & n16550;
  assign n16552 = pi32  & ~n16551;
  assign n16553 = pi32  & ~n16552;
  assign n16554 = ~n16551 & ~n16552;
  assign n16555 = ~n16553 & ~n16554;
  assign n16556 = ~n16435 & ~n16438;
  assign n16557 = n16555 & n16556;
  assign n16558 = ~n16555 & ~n16556;
  assign n16559 = ~n16557 & ~n16558;
  assign n16560 = ~n16355 & ~n16368;
  assign n16561 = n2288 & n8334;
  assign n16562 = pi85  & n8685;
  assign n16563 = pi87  & n8332;
  assign n16564 = pi86  & n8327;
  assign n16565 = ~n16563 & ~n16564;
  assign n16566 = ~n16562 & n16565;
  assign n16567 = ~n16561 & n16566;
  assign n16568 = pi50  & ~n16567;
  assign n16569 = pi50  & ~n16568;
  assign n16570 = ~n16567 & ~n16568;
  assign n16571 = ~n16569 & ~n16570;
  assign n16572 = ~n16336 & ~n16349;
  assign n16573 = ~n16297 & ~n16311;
  assign n16574 = ~n16280 & ~n16294;
  assign n16575 = pi71  & n13835;
  assign n16576 = pi72  & ~n13434;
  assign n16577 = ~n16575 & ~n16576;
  assign n16578 = n16279 & ~n16577;
  assign n16579 = ~n16279 & n16577;
  assign n16580 = ~n16578 & ~n16579;
  assign n16581 = ~n16574 & n16580;
  assign n16582 = ~n16574 & ~n16581;
  assign n16583 = ~n16579 & ~n16581;
  assign n16584 = ~n16578 & n16583;
  assign n16585 = ~n16582 & ~n16584;
  assign n16586 = n809 & n12627;
  assign n16587 = pi73  & n13004;
  assign n16588 = pi75  & n12625;
  assign n16589 = pi74  & n12620;
  assign n16590 = ~n16588 & ~n16589;
  assign n16591 = ~n16587 & n16590;
  assign n16592 = ~n16586 & n16591;
  assign n16593 = pi62  & ~n16592;
  assign n16594 = pi62  & ~n16593;
  assign n16595 = ~n16592 & ~n16593;
  assign n16596 = ~n16594 & ~n16595;
  assign n16597 = ~n16585 & n16596;
  assign n16598 = n16585 & ~n16596;
  assign n16599 = ~n16597 & ~n16598;
  assign n16600 = n1025 & n11488;
  assign n16601 = pi76  & n11847;
  assign n16602 = pi78  & n11486;
  assign n16603 = pi77  & n11481;
  assign n16604 = ~n16602 & ~n16603;
  assign n16605 = ~n16601 & n16604;
  assign n16606 = ~n16600 & n16605;
  assign n16607 = pi59  & ~n16606;
  assign n16608 = pi59  & ~n16607;
  assign n16609 = ~n16606 & ~n16607;
  assign n16610 = ~n16608 & ~n16609;
  assign n16611 = ~n16599 & ~n16610;
  assign n16612 = n16599 & n16610;
  assign n16613 = ~n16611 & ~n16612;
  assign n16614 = n16573 & ~n16613;
  assign n16615 = ~n16573 & n16613;
  assign n16616 = ~n16614 & ~n16615;
  assign n16617 = n1434 & n10394;
  assign n16618 = pi79  & n10744;
  assign n16619 = pi81  & n10392;
  assign n16620 = pi80  & n10387;
  assign n16621 = ~n16619 & ~n16620;
  assign n16622 = ~n16618 & n16621;
  assign n16623 = ~n16617 & n16622;
  assign n16624 = pi56  & ~n16623;
  assign n16625 = pi56  & ~n16624;
  assign n16626 = ~n16623 & ~n16624;
  assign n16627 = ~n16625 & ~n16626;
  assign n16628 = n16616 & ~n16627;
  assign n16629 = n16616 & ~n16628;
  assign n16630 = ~n16627 & ~n16628;
  assign n16631 = ~n16629 & ~n16630;
  assign n16632 = ~n16317 & ~n16330;
  assign n16633 = n16631 & n16632;
  assign n16634 = ~n16631 & ~n16632;
  assign n16635 = ~n16633 & ~n16634;
  assign n16636 = n1834 & n9310;
  assign n16637 = pi82  & n9701;
  assign n16638 = pi84  & n9308;
  assign n16639 = pi83  & n9303;
  assign n16640 = ~n16638 & ~n16639;
  assign n16641 = ~n16637 & n16640;
  assign n16642 = ~n16636 & n16641;
  assign n16643 = pi53  & ~n16642;
  assign n16644 = pi53  & ~n16643;
  assign n16645 = ~n16642 & ~n16643;
  assign n16646 = ~n16644 & ~n16645;
  assign n16647 = ~n16635 & n16646;
  assign n16648 = n16635 & ~n16646;
  assign n16649 = ~n16647 & ~n16648;
  assign n16650 = ~n16572 & n16649;
  assign n16651 = ~n16572 & ~n16650;
  assign n16652 = n16649 & ~n16650;
  assign n16653 = ~n16651 & ~n16652;
  assign n16654 = ~n16571 & ~n16653;
  assign n16655 = n16571 & n16653;
  assign n16656 = ~n16654 & ~n16655;
  assign n16657 = ~n16560 & n16656;
  assign n16658 = n16560 & ~n16656;
  assign n16659 = ~n16657 & ~n16658;
  assign n16660 = n2801 & n7408;
  assign n16661 = pi88  & n7740;
  assign n16662 = pi90  & n7406;
  assign n16663 = pi89  & n7401;
  assign n16664 = ~n16662 & ~n16663;
  assign n16665 = ~n16661 & n16664;
  assign n16666 = ~n16660 & n16665;
  assign n16667 = pi47  & ~n16666;
  assign n16668 = pi47  & ~n16667;
  assign n16669 = ~n16666 & ~n16667;
  assign n16670 = ~n16668 & ~n16669;
  assign n16671 = n16659 & ~n16670;
  assign n16672 = n16659 & ~n16671;
  assign n16673 = ~n16670 & ~n16671;
  assign n16674 = ~n16672 & ~n16673;
  assign n16675 = ~n16375 & ~n16388;
  assign n16676 = n16674 & n16675;
  assign n16677 = ~n16674 & ~n16675;
  assign n16678 = ~n16676 & ~n16677;
  assign n16679 = n3371 & n6539;
  assign n16680 = pi91  & n6873;
  assign n16681 = pi93  & n6537;
  assign n16682 = pi92  & n6532;
  assign n16683 = ~n16681 & ~n16682;
  assign n16684 = ~n16680 & n16683;
  assign n16685 = ~n16679 & n16684;
  assign n16686 = pi44  & ~n16685;
  assign n16687 = pi44  & ~n16686;
  assign n16688 = ~n16685 & ~n16686;
  assign n16689 = ~n16687 & ~n16688;
  assign n16690 = n16678 & ~n16689;
  assign n16691 = n16678 & ~n16690;
  assign n16692 = ~n16689 & ~n16690;
  assign n16693 = ~n16691 & ~n16692;
  assign n16694 = ~n16394 & ~n16407;
  assign n16695 = n16693 & n16694;
  assign n16696 = ~n16693 & ~n16694;
  assign n16697 = ~n16695 & ~n16696;
  assign n16698 = n4001 & n5739;
  assign n16699 = pi94  & n6030;
  assign n16700 = pi96  & n5737;
  assign n16701 = pi95  & n5732;
  assign n16702 = ~n16700 & ~n16701;
  assign n16703 = ~n16699 & n16702;
  assign n16704 = ~n16698 & n16703;
  assign n16705 = pi41  & ~n16704;
  assign n16706 = pi41  & ~n16705;
  assign n16707 = ~n16704 & ~n16705;
  assign n16708 = ~n16706 & ~n16707;
  assign n16709 = ~n16697 & n16708;
  assign n16710 = n16697 & ~n16708;
  assign n16711 = ~n16709 & ~n16710;
  assign n16712 = ~n16413 & ~n16427;
  assign n16713 = n16711 & ~n16712;
  assign n16714 = ~n16711 & n16712;
  assign n16715 = ~n16713 & ~n16714;
  assign n16716 = n4684 & n5008;
  assign n16717 = pi97  & n5241;
  assign n16718 = pi99  & n5006;
  assign n16719 = pi98  & n5001;
  assign n16720 = ~n16718 & ~n16719;
  assign n16721 = ~n16717 & n16720;
  assign n16722 = ~n16716 & n16721;
  assign n16723 = pi38  & ~n16722;
  assign n16724 = pi38  & ~n16723;
  assign n16725 = ~n16722 & ~n16723;
  assign n16726 = ~n16724 & ~n16725;
  assign n16727 = n16715 & ~n16726;
  assign n16728 = n16715 & ~n16727;
  assign n16729 = ~n16726 & ~n16727;
  assign n16730 = ~n16728 & ~n16729;
  assign n16731 = ~n16429 & ~n16432;
  assign n16732 = n16730 & n16731;
  assign n16733 = ~n16730 & ~n16731;
  assign n16734 = ~n16732 & ~n16733;
  assign n16735 = n4271 & n5413;
  assign n16736 = pi100  & n4503;
  assign n16737 = pi102  & n4269;
  assign n16738 = pi101  & n4264;
  assign n16739 = ~n16737 & ~n16738;
  assign n16740 = ~n16736 & n16739;
  assign n16741 = ~n16735 & n16740;
  assign n16742 = pi35  & ~n16741;
  assign n16743 = pi35  & ~n16742;
  assign n16744 = ~n16741 & ~n16742;
  assign n16745 = ~n16743 & ~n16744;
  assign n16746 = n16734 & ~n16745;
  assign n16747 = ~n16734 & n16745;
  assign n16748 = ~n16746 & ~n16747;
  assign n16749 = n16559 & n16748;
  assign n16750 = n16559 & ~n16749;
  assign n16751 = n16748 & ~n16749;
  assign n16752 = ~n16750 & ~n16751;
  assign n16753 = ~n16248 & ~n16442;
  assign n16754 = pi106  & n3225;
  assign n16755 = pi108  & n3032;
  assign n16756 = pi107  & n3027;
  assign n16757 = ~n16755 & ~n16756;
  assign n16758 = ~n16754 & n16757;
  assign n16759 = ~n3034 & n16758;
  assign n16760 = ~n7060 & n16758;
  assign n16761 = ~n16759 & ~n16760;
  assign n16762 = pi29  & ~n16761;
  assign n16763 = ~pi29  & n16761;
  assign n16764 = ~n16762 & ~n16763;
  assign n16765 = ~n16753 & ~n16764;
  assign n16766 = ~n16753 & ~n16765;
  assign n16767 = ~n16764 & ~n16765;
  assign n16768 = ~n16766 & ~n16767;
  assign n16769 = ~n16752 & ~n16768;
  assign n16770 = ~n16752 & ~n16769;
  assign n16771 = ~n16768 & ~n16769;
  assign n16772 = ~n16770 & ~n16771;
  assign n16773 = ~n16544 & ~n16772;
  assign n16774 = ~n16544 & ~n16773;
  assign n16775 = ~n16772 & ~n16773;
  assign n16776 = ~n16774 & ~n16775;
  assign n16777 = ~n16527 & n16776;
  assign n16778 = n16527 & ~n16776;
  assign n16779 = ~n16777 & ~n16778;
  assign n16780 = ~n16203 & ~n16452;
  assign n16781 = ~n16200 & ~n16780;
  assign n16782 = pi115  & n1745;
  assign n16783 = pi117  & n1609;
  assign n16784 = pi116  & n1604;
  assign n16785 = ~n16783 & ~n16784;
  assign n16786 = ~n16782 & n16785;
  assign n16787 = ~n1611 & n16786;
  assign n16788 = ~n9958 & n16786;
  assign n16789 = ~n16787 & ~n16788;
  assign n16790 = pi20  & ~n16789;
  assign n16791 = ~pi20  & n16789;
  assign n16792 = ~n16790 & ~n16791;
  assign n16793 = ~n16781 & ~n16792;
  assign n16794 = ~n16781 & ~n16793;
  assign n16795 = ~n16792 & ~n16793;
  assign n16796 = ~n16794 & ~n16795;
  assign n16797 = n16779 & ~n16796;
  assign n16798 = n16779 & ~n16797;
  assign n16799 = ~n16796 & ~n16797;
  assign n16800 = ~n16798 & ~n16799;
  assign n16801 = n16512 & ~n16800;
  assign n16802 = n16512 & ~n16801;
  assign n16803 = ~n16800 & ~n16801;
  assign n16804 = ~n16802 & ~n16803;
  assign n16805 = n938 & n12158;
  assign n16806 = pi121  & n1052;
  assign n16807 = pi123  & n936;
  assign n16808 = pi122  & n931;
  assign n16809 = ~n16807 & ~n16808;
  assign n16810 = ~n16806 & n16809;
  assign n16811 = ~n16805 & n16810;
  assign n16812 = pi14  & ~n16811;
  assign n16813 = pi14  & ~n16812;
  assign n16814 = ~n16811 & ~n16812;
  assign n16815 = ~n16813 & ~n16814;
  assign n16816 = ~n16170 & ~n16460;
  assign n16817 = ~n16815 & ~n16816;
  assign n16818 = ~n16815 & ~n16817;
  assign n16819 = ~n16816 & ~n16817;
  assign n16820 = ~n16818 & ~n16819;
  assign n16821 = ~n16804 & n16820;
  assign n16822 = n16804 & ~n16820;
  assign n16823 = ~n16821 & ~n16822;
  assign n16824 = ~n16154 & ~n16463;
  assign n16825 = pi124  & n763;
  assign n16826 = pi126  & n685;
  assign n16827 = pi125  & n680;
  assign n16828 = ~n16826 & ~n16827;
  assign n16829 = ~n16825 & n16828;
  assign n16830 = ~n687 & n16829;
  assign n16831 = ~n13344 & n16829;
  assign n16832 = ~n16830 & ~n16831;
  assign n16833 = pi11  & ~n16832;
  assign n16834 = ~pi11  & n16832;
  assign n16835 = ~n16833 & ~n16834;
  assign n16836 = ~n16824 & ~n16835;
  assign n16837 = ~n16824 & ~n16836;
  assign n16838 = ~n16835 & ~n16836;
  assign n16839 = ~n16837 & ~n16838;
  assign n16840 = ~n16823 & ~n16839;
  assign n16841 = n16823 & n16839;
  assign n16842 = ~n16840 & ~n16841;
  assign n16843 = ~n16497 & n16842;
  assign n16844 = n16497 & ~n16842;
  assign n16845 = ~n16843 & ~n16844;
  assign n16846 = ~n16485 & n16845;
  assign n16847 = ~n16485 & ~n16846;
  assign n16848 = n16845 & ~n16846;
  assign n16849 = ~n16847 & ~n16848;
  assign n16850 = ~n16484 & ~n16849;
  assign n16851 = n16484 & n16849;
  assign po71  = ~n16850 & ~n16851;
  assign n16853 = ~n16846 & ~n16850;
  assign n16854 = ~n16494 & ~n16843;
  assign n16855 = ~n16836 & ~n16840;
  assign n16856 = n687 & n13742;
  assign n16857 = pi125  & n763;
  assign n16858 = pi127  & n685;
  assign n16859 = pi126  & n680;
  assign n16860 = ~n16858 & ~n16859;
  assign n16861 = ~n16857 & n16860;
  assign n16862 = ~n16856 & n16861;
  assign n16863 = pi11  & ~n16862;
  assign n16864 = pi11  & ~n16863;
  assign n16865 = ~n16862 & ~n16863;
  assign n16866 = ~n16864 & ~n16865;
  assign n16867 = ~n16855 & ~n16866;
  assign n16868 = ~n16855 & ~n16867;
  assign n16869 = ~n16866 & ~n16867;
  assign n16870 = ~n16868 & ~n16869;
  assign n16871 = ~n16804 & ~n16820;
  assign n16872 = ~n16817 & ~n16871;
  assign n16873 = n938 & n12189;
  assign n16874 = pi122  & n1052;
  assign n16875 = pi124  & n936;
  assign n16876 = pi123  & n931;
  assign n16877 = ~n16875 & ~n16876;
  assign n16878 = ~n16874 & n16877;
  assign n16879 = ~n16873 & n16878;
  assign n16880 = pi14  & ~n16879;
  assign n16881 = pi14  & ~n16880;
  assign n16882 = ~n16879 & ~n16880;
  assign n16883 = ~n16881 & ~n16882;
  assign n16884 = ~n16872 & n16883;
  assign n16885 = n16872 & ~n16883;
  assign n16886 = ~n16884 & ~n16885;
  assign n16887 = n1297 & n11389;
  assign n16888 = pi119  & n1366;
  assign n16889 = pi121  & n1295;
  assign n16890 = pi120  & n1290;
  assign n16891 = ~n16889 & ~n16890;
  assign n16892 = ~n16888 & n16891;
  assign n16893 = ~n16887 & n16892;
  assign n16894 = pi17  & ~n16893;
  assign n16895 = pi17  & ~n16894;
  assign n16896 = ~n16893 & ~n16894;
  assign n16897 = ~n16895 & ~n16896;
  assign n16898 = ~n16511 & ~n16801;
  assign n16899 = n16897 & n16898;
  assign n16900 = ~n16897 & ~n16898;
  assign n16901 = ~n16899 & ~n16900;
  assign n16902 = ~n16793 & ~n16797;
  assign n16903 = n1611 & n9984;
  assign n16904 = pi116  & n1745;
  assign n16905 = pi118  & n1609;
  assign n16906 = pi117  & n1604;
  assign n16907 = ~n16905 & ~n16906;
  assign n16908 = ~n16904 & n16907;
  assign n16909 = ~n16903 & n16908;
  assign n16910 = pi20  & ~n16909;
  assign n16911 = pi20  & ~n16910;
  assign n16912 = ~n16909 & ~n16910;
  assign n16913 = ~n16911 & ~n16912;
  assign n16914 = ~n16902 & ~n16913;
  assign n16915 = ~n16902 & ~n16914;
  assign n16916 = ~n16913 & ~n16914;
  assign n16917 = ~n16915 & ~n16916;
  assign n16918 = n2523 & n7997;
  assign n16919 = pi110  & n2667;
  assign n16920 = pi112  & n2521;
  assign n16921 = pi111  & n2516;
  assign n16922 = ~n16920 & ~n16921;
  assign n16923 = ~n16919 & n16922;
  assign n16924 = ~n16918 & n16923;
  assign n16925 = pi26  & ~n16924;
  assign n16926 = pi26  & ~n16925;
  assign n16927 = ~n16924 & ~n16925;
  assign n16928 = ~n16926 & ~n16927;
  assign n16929 = ~n16541 & ~n16773;
  assign n16930 = n16928 & n16929;
  assign n16931 = ~n16928 & ~n16929;
  assign n16932 = ~n16930 & ~n16931;
  assign n16933 = ~n16765 & ~n16769;
  assign n16934 = n3034 & n7349;
  assign n16935 = pi107  & n3225;
  assign n16936 = pi109  & n3032;
  assign n16937 = pi108  & n3027;
  assign n16938 = ~n16936 & ~n16937;
  assign n16939 = ~n16935 & n16938;
  assign n16940 = ~n16934 & n16939;
  assign n16941 = pi29  & ~n16940;
  assign n16942 = pi29  & ~n16941;
  assign n16943 = ~n16940 & ~n16941;
  assign n16944 = ~n16942 & ~n16943;
  assign n16945 = ~n16933 & ~n16944;
  assign n16946 = ~n16933 & ~n16945;
  assign n16947 = ~n16944 & ~n16945;
  assign n16948 = ~n16946 & ~n16947;
  assign n16949 = ~n16558 & ~n16749;
  assign n16950 = n3622 & n6477;
  assign n16951 = pi104  & n3814;
  assign n16952 = pi106  & n3620;
  assign n16953 = pi105  & n3615;
  assign n16954 = ~n16952 & ~n16953;
  assign n16955 = ~n16951 & n16954;
  assign n16956 = ~n16950 & n16955;
  assign n16957 = pi32  & ~n16956;
  assign n16958 = pi32  & ~n16957;
  assign n16959 = ~n16956 & ~n16957;
  assign n16960 = ~n16958 & ~n16959;
  assign n16961 = ~n16949 & ~n16960;
  assign n16962 = ~n16949 & ~n16961;
  assign n16963 = ~n16960 & ~n16961;
  assign n16964 = ~n16962 & ~n16963;
  assign n16965 = ~n16713 & ~n16727;
  assign n16966 = ~n16696 & ~n16710;
  assign n16967 = ~n16677 & ~n16690;
  assign n16968 = ~n16650 & ~n16654;
  assign n16969 = n2446 & n8334;
  assign n16970 = pi86  & n8685;
  assign n16971 = pi88  & n8332;
  assign n16972 = pi87  & n8327;
  assign n16973 = ~n16971 & ~n16972;
  assign n16974 = ~n16970 & n16973;
  assign n16975 = ~n16969 & n16974;
  assign n16976 = pi50  & ~n16975;
  assign n16977 = pi50  & ~n16976;
  assign n16978 = ~n16975 & ~n16976;
  assign n16979 = ~n16977 & ~n16978;
  assign n16980 = ~n16585 & ~n16596;
  assign n16981 = ~n16611 & ~n16980;
  assign n16982 = n891 & n12627;
  assign n16983 = pi74  & n13004;
  assign n16984 = pi76  & n12625;
  assign n16985 = pi75  & n12620;
  assign n16986 = ~n16984 & ~n16985;
  assign n16987 = ~n16983 & n16986;
  assign n16988 = ~n16982 & n16987;
  assign n16989 = pi62  & ~n16988;
  assign n16990 = pi62  & ~n16989;
  assign n16991 = ~n16988 & ~n16989;
  assign n16992 = ~n16990 & ~n16991;
  assign n16993 = pi72  & n13835;
  assign n16994 = pi73  & ~n13434;
  assign n16995 = ~n16993 & ~n16994;
  assign n16996 = pi8  & ~n16577;
  assign n16997 = ~pi8  & n16577;
  assign n16998 = ~n16996 & ~n16997;
  assign n16999 = ~n16995 & ~n16998;
  assign n17000 = n16995 & n16998;
  assign n17001 = ~n16999 & ~n17000;
  assign n17002 = ~n16583 & n17001;
  assign n17003 = n16583 & ~n17001;
  assign n17004 = ~n17002 & ~n17003;
  assign n17005 = n16992 & n17004;
  assign n17006 = ~n16992 & ~n17004;
  assign n17007 = ~n17005 & ~n17006;
  assign n17008 = n1122 & n11488;
  assign n17009 = pi77  & n11847;
  assign n17010 = pi79  & n11486;
  assign n17011 = pi78  & n11481;
  assign n17012 = ~n17010 & ~n17011;
  assign n17013 = ~n17009 & n17012;
  assign n17014 = ~n17008 & n17013;
  assign n17015 = pi59  & ~n17014;
  assign n17016 = pi59  & ~n17015;
  assign n17017 = ~n17014 & ~n17015;
  assign n17018 = ~n17016 & ~n17017;
  assign n17019 = ~n17007 & ~n17018;
  assign n17020 = n17007 & n17018;
  assign n17021 = ~n17019 & ~n17020;
  assign n17022 = ~n16981 & n17021;
  assign n17023 = n16981 & ~n17021;
  assign n17024 = ~n17022 & ~n17023;
  assign n17025 = n1554 & n10394;
  assign n17026 = pi80  & n10744;
  assign n17027 = pi82  & n10392;
  assign n17028 = pi81  & n10387;
  assign n17029 = ~n17027 & ~n17028;
  assign n17030 = ~n17026 & n17029;
  assign n17031 = ~n17025 & n17030;
  assign n17032 = pi56  & ~n17031;
  assign n17033 = pi56  & ~n17032;
  assign n17034 = ~n17031 & ~n17032;
  assign n17035 = ~n17033 & ~n17034;
  assign n17036 = n17024 & ~n17035;
  assign n17037 = n17024 & ~n17036;
  assign n17038 = ~n17035 & ~n17036;
  assign n17039 = ~n17037 & ~n17038;
  assign n17040 = ~n16615 & ~n16628;
  assign n17041 = n17039 & n17040;
  assign n17042 = ~n17039 & ~n17040;
  assign n17043 = ~n17041 & ~n17042;
  assign n17044 = n1972 & n9310;
  assign n17045 = pi83  & n9701;
  assign n17046 = pi85  & n9308;
  assign n17047 = pi84  & n9303;
  assign n17048 = ~n17046 & ~n17047;
  assign n17049 = ~n17045 & n17048;
  assign n17050 = ~n17044 & n17049;
  assign n17051 = pi53  & ~n17050;
  assign n17052 = pi53  & ~n17051;
  assign n17053 = ~n17050 & ~n17051;
  assign n17054 = ~n17052 & ~n17053;
  assign n17055 = n17043 & ~n17054;
  assign n17056 = n17043 & ~n17055;
  assign n17057 = ~n17054 & ~n17055;
  assign n17058 = ~n17056 & ~n17057;
  assign n17059 = ~n16634 & ~n16648;
  assign n17060 = ~n17058 & ~n17059;
  assign n17061 = n17058 & n17059;
  assign n17062 = ~n17060 & ~n17061;
  assign n17063 = ~n16979 & n17062;
  assign n17064 = ~n16979 & ~n17063;
  assign n17065 = n17062 & ~n17063;
  assign n17066 = ~n17064 & ~n17065;
  assign n17067 = ~n16968 & ~n17066;
  assign n17068 = ~n16968 & ~n17067;
  assign n17069 = ~n17066 & ~n17067;
  assign n17070 = ~n17068 & ~n17069;
  assign n17071 = n2978 & n7408;
  assign n17072 = pi89  & n7740;
  assign n17073 = pi91  & n7406;
  assign n17074 = pi90  & n7401;
  assign n17075 = ~n17073 & ~n17074;
  assign n17076 = ~n17072 & n17075;
  assign n17077 = ~n17071 & n17076;
  assign n17078 = pi47  & ~n17077;
  assign n17079 = pi47  & ~n17078;
  assign n17080 = ~n17077 & ~n17078;
  assign n17081 = ~n17079 & ~n17080;
  assign n17082 = ~n17070 & ~n17081;
  assign n17083 = ~n17070 & ~n17082;
  assign n17084 = ~n17081 & ~n17082;
  assign n17085 = ~n17083 & ~n17084;
  assign n17086 = ~n16657 & ~n16671;
  assign n17087 = n17085 & n17086;
  assign n17088 = ~n17085 & ~n17086;
  assign n17089 = ~n17087 & ~n17088;
  assign n17090 = n3565 & n6539;
  assign n17091 = pi92  & n6873;
  assign n17092 = pi94  & n6537;
  assign n17093 = pi93  & n6532;
  assign n17094 = ~n17092 & ~n17093;
  assign n17095 = ~n17091 & n17094;
  assign n17096 = ~n17090 & n17095;
  assign n17097 = pi44  & ~n17096;
  assign n17098 = pi44  & ~n17097;
  assign n17099 = ~n17096 & ~n17097;
  assign n17100 = ~n17098 & ~n17099;
  assign n17101 = ~n17089 & n17100;
  assign n17102 = n17089 & ~n17100;
  assign n17103 = ~n16967 & ~n17101;
  assign n17104 = ~n17102 & n17103;
  assign n17105 = ~n16967 & ~n17104;
  assign n17106 = ~n17102 & ~n17104;
  assign n17107 = ~n17101 & n17106;
  assign n17108 = ~n17105 & ~n17107;
  assign n17109 = n4211 & n5739;
  assign n17110 = pi95  & n6030;
  assign n17111 = pi97  & n5737;
  assign n17112 = pi96  & n5732;
  assign n17113 = ~n17111 & ~n17112;
  assign n17114 = ~n17110 & n17113;
  assign n17115 = ~n17109 & n17114;
  assign n17116 = pi41  & ~n17115;
  assign n17117 = pi41  & ~n17116;
  assign n17118 = ~n17115 & ~n17116;
  assign n17119 = ~n17117 & ~n17118;
  assign n17120 = ~n17108 & ~n17119;
  assign n17121 = ~n17108 & ~n17120;
  assign n17122 = ~n17119 & ~n17120;
  assign n17123 = ~n17121 & ~n17122;
  assign n17124 = ~n16966 & n17123;
  assign n17125 = n16966 & ~n17123;
  assign n17126 = ~n17124 & ~n17125;
  assign n17127 = n4910 & n5008;
  assign n17128 = pi98  & n5241;
  assign n17129 = pi100  & n5006;
  assign n17130 = pi99  & n5001;
  assign n17131 = ~n17129 & ~n17130;
  assign n17132 = ~n17128 & n17131;
  assign n17133 = ~n17127 & n17132;
  assign n17134 = pi38  & ~n17133;
  assign n17135 = pi38  & ~n17134;
  assign n17136 = ~n17133 & ~n17134;
  assign n17137 = ~n17135 & ~n17136;
  assign n17138 = ~n17126 & ~n17137;
  assign n17139 = n17126 & n17137;
  assign n17140 = ~n17138 & ~n17139;
  assign n17141 = n16965 & ~n17140;
  assign n17142 = ~n16965 & n17140;
  assign n17143 = ~n17141 & ~n17142;
  assign n17144 = n4271 & n5664;
  assign n17145 = pi101  & n4503;
  assign n17146 = pi103  & n4269;
  assign n17147 = pi102  & n4264;
  assign n17148 = ~n17146 & ~n17147;
  assign n17149 = ~n17145 & n17148;
  assign n17150 = ~n17144 & n17149;
  assign n17151 = pi35  & ~n17150;
  assign n17152 = pi35  & ~n17151;
  assign n17153 = ~n17150 & ~n17151;
  assign n17154 = ~n17152 & ~n17153;
  assign n17155 = n17143 & ~n17154;
  assign n17156 = n17143 & ~n17155;
  assign n17157 = ~n17154 & ~n17155;
  assign n17158 = ~n17156 & ~n17157;
  assign n17159 = ~n16733 & ~n16746;
  assign n17160 = ~n17158 & ~n17159;
  assign n17161 = ~n17158 & ~n17160;
  assign n17162 = ~n17159 & ~n17160;
  assign n17163 = ~n17161 & ~n17162;
  assign n17164 = ~n16964 & ~n17163;
  assign n17165 = ~n16964 & ~n17164;
  assign n17166 = ~n17163 & ~n17164;
  assign n17167 = ~n17165 & ~n17166;
  assign n17168 = ~n16948 & n17167;
  assign n17169 = n16948 & ~n17167;
  assign n17170 = ~n17168 & ~n17169;
  assign n17171 = n16932 & ~n17170;
  assign n17172 = n16932 & ~n17171;
  assign n17173 = ~n17170 & ~n17171;
  assign n17174 = ~n17172 & ~n17173;
  assign n17175 = n2043 & n8963;
  assign n17176 = pi113  & n2180;
  assign n17177 = pi115  & n2041;
  assign n17178 = pi114  & n2036;
  assign n17179 = ~n17177 & ~n17178;
  assign n17180 = ~n17176 & n17179;
  assign n17181 = ~n17175 & n17180;
  assign n17182 = pi23  & ~n17181;
  assign n17183 = pi23  & ~n17182;
  assign n17184 = ~n17181 & ~n17182;
  assign n17185 = ~n17183 & ~n17184;
  assign n17186 = ~n16526 & ~n16778;
  assign n17187 = ~n17185 & ~n17186;
  assign n17188 = n17185 & n17186;
  assign n17189 = ~n17187 & ~n17188;
  assign n17190 = ~n17174 & n17189;
  assign n17191 = ~n17174 & ~n17190;
  assign n17192 = n17189 & ~n17190;
  assign n17193 = ~n17191 & ~n17192;
  assign n17194 = ~n16917 & ~n17193;
  assign n17195 = ~n16917 & ~n17194;
  assign n17196 = ~n17193 & ~n17194;
  assign n17197 = ~n17195 & ~n17196;
  assign n17198 = n16901 & ~n17197;
  assign n17199 = ~n16901 & n17197;
  assign n17200 = ~n17198 & ~n17199;
  assign n17201 = ~n16886 & n17200;
  assign n17202 = ~n16886 & ~n17201;
  assign n17203 = n17200 & ~n17201;
  assign n17204 = ~n17202 & ~n17203;
  assign n17205 = ~n16870 & n17204;
  assign n17206 = n16870 & ~n17204;
  assign n17207 = ~n17205 & ~n17206;
  assign n17208 = ~n16854 & ~n17207;
  assign n17209 = ~n16854 & ~n17208;
  assign n17210 = ~n17207 & ~n17208;
  assign n17211 = ~n17209 & ~n17210;
  assign n17212 = ~n16853 & ~n17211;
  assign n17213 = n16853 & n17211;
  assign po72  = ~n17212 & ~n17213;
  assign n17215 = ~n17208 & ~n17212;
  assign n17216 = ~n16870 & ~n17204;
  assign n17217 = ~n16867 & ~n17216;
  assign n17218 = n938 & n12943;
  assign n17219 = pi123  & n1052;
  assign n17220 = pi125  & n936;
  assign n17221 = pi124  & n931;
  assign n17222 = ~n17220 & ~n17221;
  assign n17223 = ~n17219 & n17222;
  assign n17224 = ~n17218 & n17223;
  assign n17225 = pi14  & ~n17224;
  assign n17226 = pi14  & ~n17225;
  assign n17227 = ~n17224 & ~n17225;
  assign n17228 = ~n17226 & ~n17227;
  assign n17229 = ~n16900 & ~n17198;
  assign n17230 = ~n17228 & ~n17229;
  assign n17231 = ~n17228 & ~n17230;
  assign n17232 = ~n17229 & ~n17230;
  assign n17233 = ~n17231 & ~n17232;
  assign n17234 = n1611 & n10667;
  assign n17235 = pi117  & n1745;
  assign n17236 = pi119  & n1609;
  assign n17237 = pi118  & n1604;
  assign n17238 = ~n17236 & ~n17237;
  assign n17239 = ~n17235 & n17238;
  assign n17240 = ~n17234 & n17239;
  assign n17241 = pi20  & ~n17240;
  assign n17242 = pi20  & ~n17241;
  assign n17243 = ~n17240 & ~n17241;
  assign n17244 = ~n17242 & ~n17243;
  assign n17245 = ~n17187 & ~n17190;
  assign n17246 = n17244 & n17245;
  assign n17247 = ~n17244 & ~n17245;
  assign n17248 = ~n17246 & ~n17247;
  assign n17249 = n2043 & n9614;
  assign n17250 = pi114  & n2180;
  assign n17251 = pi116  & n2041;
  assign n17252 = pi115  & n2036;
  assign n17253 = ~n17251 & ~n17252;
  assign n17254 = ~n17250 & n17253;
  assign n17255 = ~n17249 & n17254;
  assign n17256 = pi23  & ~n17255;
  assign n17257 = pi23  & ~n17256;
  assign n17258 = ~n17255 & ~n17256;
  assign n17259 = ~n17257 & ~n17258;
  assign n17260 = ~n16931 & ~n17171;
  assign n17261 = n17259 & n17260;
  assign n17262 = ~n17259 & ~n17260;
  assign n17263 = ~n17261 & ~n17262;
  assign n17264 = n2523 & n8612;
  assign n17265 = pi111  & n2667;
  assign n17266 = pi113  & n2521;
  assign n17267 = pi112  & n2516;
  assign n17268 = ~n17266 & ~n17267;
  assign n17269 = ~n17265 & n17268;
  assign n17270 = ~n17264 & n17269;
  assign n17271 = pi26  & ~n17270;
  assign n17272 = pi26  & ~n17271;
  assign n17273 = ~n17270 & ~n17271;
  assign n17274 = ~n17272 & ~n17273;
  assign n17275 = ~n16948 & ~n17167;
  assign n17276 = ~n16945 & ~n17275;
  assign n17277 = ~n17274 & ~n17276;
  assign n17278 = ~n17274 & ~n17277;
  assign n17279 = ~n17276 & ~n17277;
  assign n17280 = ~n17278 & ~n17279;
  assign n17281 = n3622 & n6775;
  assign n17282 = pi105  & n3814;
  assign n17283 = pi107  & n3620;
  assign n17284 = pi106  & n3615;
  assign n17285 = ~n17283 & ~n17284;
  assign n17286 = ~n17282 & n17285;
  assign n17287 = ~n17281 & n17286;
  assign n17288 = pi32  & ~n17287;
  assign n17289 = pi32  & ~n17288;
  assign n17290 = ~n17287 & ~n17288;
  assign n17291 = ~n17289 & ~n17290;
  assign n17292 = ~n17155 & ~n17160;
  assign n17293 = n17291 & n17292;
  assign n17294 = ~n17291 & ~n17292;
  assign n17295 = ~n17293 & ~n17294;
  assign n17296 = n4271 & n5943;
  assign n17297 = pi102  & n4503;
  assign n17298 = pi104  & n4269;
  assign n17299 = pi103  & n4264;
  assign n17300 = ~n17298 & ~n17299;
  assign n17301 = ~n17297 & n17300;
  assign n17302 = ~n17296 & n17301;
  assign n17303 = pi35  & ~n17302;
  assign n17304 = pi35  & ~n17303;
  assign n17305 = ~n17302 & ~n17303;
  assign n17306 = ~n17304 & ~n17305;
  assign n17307 = ~n17138 & ~n17142;
  assign n17308 = n5008 & n5169;
  assign n17309 = pi99  & n5241;
  assign n17310 = pi101  & n5006;
  assign n17311 = pi100  & n5001;
  assign n17312 = ~n17310 & ~n17311;
  assign n17313 = ~n17309 & n17312;
  assign n17314 = ~n17308 & n17313;
  assign n17315 = pi38  & ~n17314;
  assign n17316 = pi38  & ~n17315;
  assign n17317 = ~n17314 & ~n17315;
  assign n17318 = ~n17316 & ~n17317;
  assign n17319 = ~n16966 & ~n17123;
  assign n17320 = ~n17120 & ~n17319;
  assign n17321 = n4454 & n5739;
  assign n17322 = pi96  & n6030;
  assign n17323 = pi98  & n5737;
  assign n17324 = pi97  & n5732;
  assign n17325 = ~n17323 & ~n17324;
  assign n17326 = ~n17322 & n17325;
  assign n17327 = ~n17321 & n17326;
  assign n17328 = pi41  & ~n17327;
  assign n17329 = pi41  & ~n17328;
  assign n17330 = ~n17327 & ~n17328;
  assign n17331 = ~n17329 & ~n17330;
  assign n17332 = n999 & n12627;
  assign n17333 = pi75  & n13004;
  assign n17334 = pi77  & n12625;
  assign n17335 = pi76  & n12620;
  assign n17336 = ~n17334 & ~n17335;
  assign n17337 = ~n17333 & n17336;
  assign n17338 = ~n17332 & n17337;
  assign n17339 = pi62  & ~n17338;
  assign n17340 = pi62  & ~n17339;
  assign n17341 = ~n17338 & ~n17339;
  assign n17342 = ~n17340 & ~n17341;
  assign n17343 = pi73  & n13835;
  assign n17344 = pi74  & ~n13434;
  assign n17345 = ~n17343 & ~n17344;
  assign n17346 = ~pi8  & ~n16577;
  assign n17347 = ~n16999 & ~n17346;
  assign n17348 = n17345 & ~n17347;
  assign n17349 = n17345 & ~n17348;
  assign n17350 = ~n17347 & ~n17348;
  assign n17351 = ~n17349 & ~n17350;
  assign n17352 = ~n17342 & ~n17351;
  assign n17353 = ~n17342 & ~n17352;
  assign n17354 = ~n17351 & ~n17352;
  assign n17355 = ~n17353 & ~n17354;
  assign n17356 = ~n17003 & ~n17005;
  assign n17357 = ~n17355 & n17356;
  assign n17358 = ~n17355 & ~n17357;
  assign n17359 = n17356 & ~n17357;
  assign n17360 = ~n17358 & ~n17359;
  assign n17361 = n1225 & n11488;
  assign n17362 = pi78  & n11847;
  assign n17363 = pi80  & n11486;
  assign n17364 = pi79  & n11481;
  assign n17365 = ~n17363 & ~n17364;
  assign n17366 = ~n17362 & n17365;
  assign n17367 = ~n17361 & n17366;
  assign n17368 = pi59  & ~n17367;
  assign n17369 = pi59  & ~n17368;
  assign n17370 = ~n17367 & ~n17368;
  assign n17371 = ~n17369 & ~n17370;
  assign n17372 = ~n17360 & ~n17371;
  assign n17373 = ~n17360 & ~n17372;
  assign n17374 = ~n17371 & ~n17372;
  assign n17375 = ~n17373 & ~n17374;
  assign n17376 = ~n17019 & ~n17022;
  assign n17377 = n17375 & n17376;
  assign n17378 = ~n17375 & ~n17376;
  assign n17379 = ~n17377 & ~n17378;
  assign n17380 = n1696 & n10394;
  assign n17381 = pi81  & n10744;
  assign n17382 = pi83  & n10392;
  assign n17383 = pi82  & n10387;
  assign n17384 = ~n17382 & ~n17383;
  assign n17385 = ~n17381 & n17384;
  assign n17386 = ~n17380 & n17385;
  assign n17387 = pi56  & ~n17386;
  assign n17388 = pi56  & ~n17387;
  assign n17389 = ~n17386 & ~n17387;
  assign n17390 = ~n17388 & ~n17389;
  assign n17391 = n17379 & ~n17390;
  assign n17392 = n17379 & ~n17391;
  assign n17393 = ~n17390 & ~n17391;
  assign n17394 = ~n17392 & ~n17393;
  assign n17395 = ~n17036 & ~n17042;
  assign n17396 = n17394 & n17395;
  assign n17397 = ~n17394 & ~n17395;
  assign n17398 = ~n17396 & ~n17397;
  assign n17399 = n2133 & n9310;
  assign n17400 = pi84  & n9701;
  assign n17401 = pi86  & n9308;
  assign n17402 = pi85  & n9303;
  assign n17403 = ~n17401 & ~n17402;
  assign n17404 = ~n17400 & n17403;
  assign n17405 = ~n17399 & n17404;
  assign n17406 = pi53  & ~n17405;
  assign n17407 = pi53  & ~n17406;
  assign n17408 = ~n17405 & ~n17406;
  assign n17409 = ~n17407 & ~n17408;
  assign n17410 = n17398 & ~n17409;
  assign n17411 = n17398 & ~n17410;
  assign n17412 = ~n17409 & ~n17410;
  assign n17413 = ~n17411 & ~n17412;
  assign n17414 = ~n17055 & ~n17060;
  assign n17415 = n17413 & n17414;
  assign n17416 = ~n17413 & ~n17414;
  assign n17417 = ~n17415 & ~n17416;
  assign n17418 = n2473 & n8334;
  assign n17419 = pi87  & n8685;
  assign n17420 = pi89  & n8332;
  assign n17421 = pi88  & n8327;
  assign n17422 = ~n17420 & ~n17421;
  assign n17423 = ~n17419 & n17422;
  assign n17424 = ~n17418 & n17423;
  assign n17425 = pi50  & ~n17424;
  assign n17426 = pi50  & ~n17425;
  assign n17427 = ~n17424 & ~n17425;
  assign n17428 = ~n17426 & ~n17427;
  assign n17429 = n17417 & ~n17428;
  assign n17430 = n17417 & ~n17429;
  assign n17431 = ~n17428 & ~n17429;
  assign n17432 = ~n17430 & ~n17431;
  assign n17433 = ~n17063 & ~n17067;
  assign n17434 = n17432 & n17433;
  assign n17435 = ~n17432 & ~n17433;
  assign n17436 = ~n17434 & ~n17435;
  assign n17437 = n3177 & n7408;
  assign n17438 = pi90  & n7740;
  assign n17439 = pi92  & n7406;
  assign n17440 = pi91  & n7401;
  assign n17441 = ~n17439 & ~n17440;
  assign n17442 = ~n17438 & n17441;
  assign n17443 = ~n17437 & n17442;
  assign n17444 = pi47  & ~n17443;
  assign n17445 = pi47  & ~n17444;
  assign n17446 = ~n17443 & ~n17444;
  assign n17447 = ~n17445 & ~n17446;
  assign n17448 = n17436 & ~n17447;
  assign n17449 = n17436 & ~n17448;
  assign n17450 = ~n17447 & ~n17448;
  assign n17451 = ~n17449 & ~n17450;
  assign n17452 = ~n17082 & ~n17088;
  assign n17453 = n17451 & n17452;
  assign n17454 = ~n17451 & ~n17452;
  assign n17455 = ~n17453 & ~n17454;
  assign n17456 = n3784 & n6539;
  assign n17457 = pi93  & n6873;
  assign n17458 = pi95  & n6537;
  assign n17459 = pi94  & n6532;
  assign n17460 = ~n17458 & ~n17459;
  assign n17461 = ~n17457 & n17460;
  assign n17462 = ~n17456 & n17461;
  assign n17463 = pi44  & ~n17462;
  assign n17464 = pi44  & ~n17463;
  assign n17465 = ~n17462 & ~n17463;
  assign n17466 = ~n17464 & ~n17465;
  assign n17467 = ~n17455 & n17466;
  assign n17468 = n17455 & ~n17466;
  assign n17469 = ~n17467 & ~n17468;
  assign n17470 = ~n17106 & n17469;
  assign n17471 = n17106 & ~n17469;
  assign n17472 = ~n17470 & ~n17471;
  assign n17473 = ~n17331 & n17472;
  assign n17474 = n17331 & ~n17472;
  assign n17475 = ~n17473 & ~n17474;
  assign n17476 = ~n17320 & n17475;
  assign n17477 = ~n17320 & ~n17476;
  assign n17478 = n17475 & ~n17476;
  assign n17479 = ~n17477 & ~n17478;
  assign n17480 = ~n17318 & ~n17479;
  assign n17481 = n17318 & n17479;
  assign n17482 = ~n17480 & ~n17481;
  assign n17483 = ~n17307 & n17482;
  assign n17484 = ~n17307 & ~n17483;
  assign n17485 = n17482 & ~n17483;
  assign n17486 = ~n17484 & ~n17485;
  assign n17487 = ~n17306 & ~n17486;
  assign n17488 = ~n17306 & ~n17487;
  assign n17489 = ~n17486 & ~n17487;
  assign n17490 = ~n17488 & ~n17489;
  assign n17491 = n17295 & ~n17490;
  assign n17492 = n17295 & ~n17491;
  assign n17493 = ~n17490 & ~n17491;
  assign n17494 = ~n17492 & ~n17493;
  assign n17495 = ~n16961 & ~n17164;
  assign n17496 = pi108  & n3225;
  assign n17497 = pi110  & n3032;
  assign n17498 = pi109  & n3027;
  assign n17499 = ~n17497 & ~n17498;
  assign n17500 = ~n17496 & n17499;
  assign n17501 = ~n3034 & n17500;
  assign n17502 = ~n7665 & n17500;
  assign n17503 = ~n17501 & ~n17502;
  assign n17504 = pi29  & ~n17503;
  assign n17505 = ~pi29  & n17503;
  assign n17506 = ~n17504 & ~n17505;
  assign n17507 = ~n17495 & ~n17506;
  assign n17508 = ~n17495 & ~n17507;
  assign n17509 = ~n17506 & ~n17507;
  assign n17510 = ~n17508 & ~n17509;
  assign n17511 = ~n17494 & ~n17510;
  assign n17512 = ~n17494 & ~n17511;
  assign n17513 = ~n17510 & ~n17511;
  assign n17514 = ~n17512 & ~n17513;
  assign n17515 = ~n17280 & ~n17514;
  assign n17516 = ~n17280 & ~n17515;
  assign n17517 = ~n17514 & ~n17515;
  assign n17518 = ~n17516 & ~n17517;
  assign n17519 = n17263 & ~n17518;
  assign n17520 = ~n17263 & n17518;
  assign n17521 = ~n17519 & ~n17520;
  assign n17522 = n17248 & n17521;
  assign n17523 = n17248 & ~n17522;
  assign n17524 = n17521 & ~n17522;
  assign n17525 = ~n17523 & ~n17524;
  assign n17526 = ~n16914 & ~n17194;
  assign n17527 = pi120  & n1366;
  assign n17528 = pi122  & n1295;
  assign n17529 = pi121  & n1290;
  assign n17530 = ~n17528 & ~n17529;
  assign n17531 = ~n17527 & n17530;
  assign n17532 = ~n1297 & n17531;
  assign n17533 = ~n11778 & n17531;
  assign n17534 = ~n17532 & ~n17533;
  assign n17535 = pi17  & ~n17534;
  assign n17536 = ~pi17  & n17534;
  assign n17537 = ~n17535 & ~n17536;
  assign n17538 = ~n17526 & ~n17537;
  assign n17539 = ~n17526 & ~n17538;
  assign n17540 = ~n17537 & ~n17538;
  assign n17541 = ~n17539 & ~n17540;
  assign n17542 = ~n17525 & ~n17541;
  assign n17543 = ~n17525 & ~n17542;
  assign n17544 = ~n17541 & ~n17542;
  assign n17545 = ~n17543 & ~n17544;
  assign n17546 = ~n17233 & ~n17545;
  assign n17547 = ~n17233 & ~n17546;
  assign n17548 = ~n17545 & ~n17546;
  assign n17549 = ~n17547 & ~n17548;
  assign n17550 = ~n16872 & ~n16883;
  assign n17551 = ~n17201 & ~n17550;
  assign n17552 = pi126  & n763;
  assign n17553 = pi127  & n680;
  assign n17554 = ~n17552 & ~n17553;
  assign n17555 = ~n687 & n17554;
  assign n17556 = n13773 & n17554;
  assign n17557 = ~n17555 & ~n17556;
  assign n17558 = pi11  & ~n17557;
  assign n17559 = ~pi11  & n17557;
  assign n17560 = ~n17558 & ~n17559;
  assign n17561 = ~n17551 & ~n17560;
  assign n17562 = ~n17551 & ~n17561;
  assign n17563 = ~n17560 & ~n17561;
  assign n17564 = ~n17562 & ~n17563;
  assign n17565 = ~n17549 & ~n17564;
  assign n17566 = n17549 & n17564;
  assign n17567 = ~n17565 & ~n17566;
  assign n17568 = ~n17217 & n17567;
  assign n17569 = ~n17217 & ~n17568;
  assign n17570 = n17567 & ~n17568;
  assign n17571 = ~n17569 & ~n17570;
  assign n17572 = ~n17215 & ~n17571;
  assign n17573 = n17215 & n17571;
  assign po73  = ~n17572 & ~n17573;
  assign n17575 = ~n17568 & ~n17572;
  assign n17576 = ~n17561 & ~n17565;
  assign n17577 = ~n17230 & ~n17546;
  assign n17578 = pi127  & n763;
  assign n17579 = n687 & n13770;
  assign n17580 = ~n17578 & ~n17579;
  assign n17581 = pi11  & ~n17580;
  assign n17582 = pi11  & ~n17581;
  assign n17583 = ~n17580 & ~n17581;
  assign n17584 = ~n17582 & ~n17583;
  assign n17585 = ~n17577 & ~n17584;
  assign n17586 = ~n17577 & ~n17585;
  assign n17587 = ~n17584 & ~n17585;
  assign n17588 = ~n17586 & ~n17587;
  assign n17589 = ~n17538 & ~n17542;
  assign n17590 = pi124  & n1052;
  assign n17591 = pi126  & n936;
  assign n17592 = pi125  & n931;
  assign n17593 = ~n17591 & ~n17592;
  assign n17594 = ~n17590 & n17593;
  assign n17595 = ~n938 & n17594;
  assign n17596 = ~n13344 & n17594;
  assign n17597 = ~n17595 & ~n17596;
  assign n17598 = pi14  & ~n17597;
  assign n17599 = ~pi14  & n17597;
  assign n17600 = ~n17598 & ~n17599;
  assign n17601 = ~n17589 & ~n17600;
  assign n17602 = n17589 & n17600;
  assign n17603 = ~n17601 & ~n17602;
  assign n17604 = n1297 & n12158;
  assign n17605 = pi121  & n1366;
  assign n17606 = pi123  & n1295;
  assign n17607 = pi122  & n1290;
  assign n17608 = ~n17606 & ~n17607;
  assign n17609 = ~n17605 & n17608;
  assign n17610 = ~n17604 & n17609;
  assign n17611 = pi17  & ~n17610;
  assign n17612 = pi17  & ~n17611;
  assign n17613 = ~n17610 & ~n17611;
  assign n17614 = ~n17612 & ~n17613;
  assign n17615 = ~n17247 & ~n17522;
  assign n17616 = n17614 & n17615;
  assign n17617 = ~n17614 & ~n17615;
  assign n17618 = ~n17616 & ~n17617;
  assign n17619 = n1611 & n11028;
  assign n17620 = pi118  & n1745;
  assign n17621 = pi120  & n1609;
  assign n17622 = pi119  & n1604;
  assign n17623 = ~n17621 & ~n17622;
  assign n17624 = ~n17620 & n17623;
  assign n17625 = ~n17619 & n17624;
  assign n17626 = pi20  & ~n17625;
  assign n17627 = pi20  & ~n17626;
  assign n17628 = ~n17625 & ~n17626;
  assign n17629 = ~n17627 & ~n17628;
  assign n17630 = ~n17262 & ~n17519;
  assign n17631 = ~n17629 & ~n17630;
  assign n17632 = ~n17629 & ~n17631;
  assign n17633 = ~n17630 & ~n17631;
  assign n17634 = ~n17632 & ~n17633;
  assign n17635 = ~n17507 & ~n17511;
  assign n17636 = pi112  & n2667;
  assign n17637 = pi114  & n2521;
  assign n17638 = pi113  & n2516;
  assign n17639 = ~n17637 & ~n17638;
  assign n17640 = ~n17636 & n17639;
  assign n17641 = ~n2523 & n17640;
  assign n17642 = ~n8936 & n17640;
  assign n17643 = ~n17641 & ~n17642;
  assign n17644 = pi26  & ~n17643;
  assign n17645 = ~pi26  & n17643;
  assign n17646 = ~n17644 & ~n17645;
  assign n17647 = ~n17635 & ~n17646;
  assign n17648 = n17635 & n17646;
  assign n17649 = ~n17647 & ~n17648;
  assign n17650 = n3034 & n7970;
  assign n17651 = pi109  & n3225;
  assign n17652 = pi111  & n3032;
  assign n17653 = pi110  & n3027;
  assign n17654 = ~n17652 & ~n17653;
  assign n17655 = ~n17651 & n17654;
  assign n17656 = ~n17650 & n17655;
  assign n17657 = pi29  & ~n17656;
  assign n17658 = pi29  & ~n17657;
  assign n17659 = ~n17656 & ~n17657;
  assign n17660 = ~n17658 & ~n17659;
  assign n17661 = ~n17294 & ~n17491;
  assign n17662 = n17660 & n17661;
  assign n17663 = ~n17660 & ~n17661;
  assign n17664 = ~n17662 & ~n17663;
  assign n17665 = ~n17483 & ~n17487;
  assign n17666 = pi106  & n3814;
  assign n17667 = pi108  & n3620;
  assign n17668 = pi107  & n3615;
  assign n17669 = ~n17667 & ~n17668;
  assign n17670 = ~n17666 & n17669;
  assign n17671 = ~n3622 & n17670;
  assign n17672 = ~n7060 & n17670;
  assign n17673 = ~n17671 & ~n17672;
  assign n17674 = pi32  & ~n17673;
  assign n17675 = ~pi32  & n17673;
  assign n17676 = ~n17674 & ~n17675;
  assign n17677 = ~n17665 & ~n17676;
  assign n17678 = n17665 & n17676;
  assign n17679 = ~n17677 & ~n17678;
  assign n17680 = n4271 & n6207;
  assign n17681 = pi103  & n4503;
  assign n17682 = pi105  & n4269;
  assign n17683 = pi104  & n4264;
  assign n17684 = ~n17682 & ~n17683;
  assign n17685 = ~n17681 & n17684;
  assign n17686 = ~n17680 & n17685;
  assign n17687 = pi35  & ~n17686;
  assign n17688 = pi35  & ~n17687;
  assign n17689 = ~n17686 & ~n17687;
  assign n17690 = ~n17688 & ~n17689;
  assign n17691 = ~n17476 & ~n17480;
  assign n17692 = ~n17416 & ~n17429;
  assign n17693 = n2801 & n8334;
  assign n17694 = pi88  & n8685;
  assign n17695 = pi90  & n8332;
  assign n17696 = pi89  & n8327;
  assign n17697 = ~n17695 & ~n17696;
  assign n17698 = ~n17694 & n17697;
  assign n17699 = ~n17693 & n17698;
  assign n17700 = pi50  & ~n17699;
  assign n17701 = pi50  & ~n17700;
  assign n17702 = ~n17699 & ~n17700;
  assign n17703 = ~n17701 & ~n17702;
  assign n17704 = ~n17397 & ~n17410;
  assign n17705 = n2288 & n9310;
  assign n17706 = pi85  & n9701;
  assign n17707 = pi87  & n9308;
  assign n17708 = pi86  & n9303;
  assign n17709 = ~n17707 & ~n17708;
  assign n17710 = ~n17706 & n17709;
  assign n17711 = ~n17705 & n17710;
  assign n17712 = pi53  & ~n17711;
  assign n17713 = pi53  & ~n17712;
  assign n17714 = ~n17711 & ~n17712;
  assign n17715 = ~n17713 & ~n17714;
  assign n17716 = ~n17378 & ~n17391;
  assign n17717 = ~n17348 & ~n17352;
  assign n17718 = pi74  & n13835;
  assign n17719 = pi75  & ~n13434;
  assign n17720 = ~n17718 & ~n17719;
  assign n17721 = n17345 & ~n17720;
  assign n17722 = n17345 & ~n17721;
  assign n17723 = ~n17720 & ~n17721;
  assign n17724 = ~n17722 & ~n17723;
  assign n17725 = ~n17717 & ~n17724;
  assign n17726 = ~n17717 & ~n17725;
  assign n17727 = ~n17724 & ~n17725;
  assign n17728 = ~n17726 & ~n17727;
  assign n17729 = n1025 & n12627;
  assign n17730 = pi76  & n13004;
  assign n17731 = pi78  & n12625;
  assign n17732 = pi77  & n12620;
  assign n17733 = ~n17731 & ~n17732;
  assign n17734 = ~n17730 & n17733;
  assign n17735 = ~n17729 & n17734;
  assign n17736 = pi62  & ~n17735;
  assign n17737 = pi62  & ~n17736;
  assign n17738 = ~n17735 & ~n17736;
  assign n17739 = ~n17737 & ~n17738;
  assign n17740 = ~n17728 & ~n17739;
  assign n17741 = ~n17728 & ~n17740;
  assign n17742 = ~n17739 & ~n17740;
  assign n17743 = ~n17741 & ~n17742;
  assign n17744 = n1434 & n11488;
  assign n17745 = pi79  & n11847;
  assign n17746 = pi81  & n11486;
  assign n17747 = pi80  & n11481;
  assign n17748 = ~n17746 & ~n17747;
  assign n17749 = ~n17745 & n17748;
  assign n17750 = ~n17744 & n17749;
  assign n17751 = pi59  & ~n17750;
  assign n17752 = pi59  & ~n17751;
  assign n17753 = ~n17750 & ~n17751;
  assign n17754 = ~n17752 & ~n17753;
  assign n17755 = ~n17743 & ~n17754;
  assign n17756 = ~n17743 & ~n17755;
  assign n17757 = ~n17754 & ~n17755;
  assign n17758 = ~n17756 & ~n17757;
  assign n17759 = ~n17357 & ~n17372;
  assign n17760 = n17758 & n17759;
  assign n17761 = ~n17758 & ~n17759;
  assign n17762 = ~n17760 & ~n17761;
  assign n17763 = n1834 & n10394;
  assign n17764 = pi82  & n10744;
  assign n17765 = pi84  & n10392;
  assign n17766 = pi83  & n10387;
  assign n17767 = ~n17765 & ~n17766;
  assign n17768 = ~n17764 & n17767;
  assign n17769 = ~n17763 & n17768;
  assign n17770 = pi56  & ~n17769;
  assign n17771 = pi56  & ~n17770;
  assign n17772 = ~n17769 & ~n17770;
  assign n17773 = ~n17771 & ~n17772;
  assign n17774 = ~n17762 & n17773;
  assign n17775 = n17762 & ~n17773;
  assign n17776 = ~n17774 & ~n17775;
  assign n17777 = ~n17716 & n17776;
  assign n17778 = ~n17716 & ~n17777;
  assign n17779 = n17776 & ~n17777;
  assign n17780 = ~n17778 & ~n17779;
  assign n17781 = ~n17715 & ~n17780;
  assign n17782 = n17715 & n17780;
  assign n17783 = ~n17781 & ~n17782;
  assign n17784 = ~n17704 & n17783;
  assign n17785 = n17704 & ~n17783;
  assign n17786 = ~n17784 & ~n17785;
  assign n17787 = ~n17703 & n17786;
  assign n17788 = n17703 & ~n17786;
  assign n17789 = ~n17787 & ~n17788;
  assign n17790 = ~n17692 & n17789;
  assign n17791 = n17692 & ~n17789;
  assign n17792 = ~n17790 & ~n17791;
  assign n17793 = n3371 & n7408;
  assign n17794 = pi91  & n7740;
  assign n17795 = pi93  & n7406;
  assign n17796 = pi92  & n7401;
  assign n17797 = ~n17795 & ~n17796;
  assign n17798 = ~n17794 & n17797;
  assign n17799 = ~n17793 & n17798;
  assign n17800 = pi47  & ~n17799;
  assign n17801 = pi47  & ~n17800;
  assign n17802 = ~n17799 & ~n17800;
  assign n17803 = ~n17801 & ~n17802;
  assign n17804 = n17792 & ~n17803;
  assign n17805 = n17792 & ~n17804;
  assign n17806 = ~n17803 & ~n17804;
  assign n17807 = ~n17805 & ~n17806;
  assign n17808 = ~n17435 & ~n17448;
  assign n17809 = n17807 & n17808;
  assign n17810 = ~n17807 & ~n17808;
  assign n17811 = ~n17809 & ~n17810;
  assign n17812 = n4001 & n6539;
  assign n17813 = pi94  & n6873;
  assign n17814 = pi96  & n6537;
  assign n17815 = pi95  & n6532;
  assign n17816 = ~n17814 & ~n17815;
  assign n17817 = ~n17813 & n17816;
  assign n17818 = ~n17812 & n17817;
  assign n17819 = pi44  & ~n17818;
  assign n17820 = pi44  & ~n17819;
  assign n17821 = ~n17818 & ~n17819;
  assign n17822 = ~n17820 & ~n17821;
  assign n17823 = ~n17811 & n17822;
  assign n17824 = n17811 & ~n17822;
  assign n17825 = ~n17823 & ~n17824;
  assign n17826 = ~n17454 & ~n17468;
  assign n17827 = n17825 & ~n17826;
  assign n17828 = ~n17825 & n17826;
  assign n17829 = ~n17827 & ~n17828;
  assign n17830 = n4684 & n5739;
  assign n17831 = pi97  & n6030;
  assign n17832 = pi99  & n5737;
  assign n17833 = pi98  & n5732;
  assign n17834 = ~n17832 & ~n17833;
  assign n17835 = ~n17831 & n17834;
  assign n17836 = ~n17830 & n17835;
  assign n17837 = pi41  & ~n17836;
  assign n17838 = pi41  & ~n17837;
  assign n17839 = ~n17836 & ~n17837;
  assign n17840 = ~n17838 & ~n17839;
  assign n17841 = n17829 & ~n17840;
  assign n17842 = n17829 & ~n17841;
  assign n17843 = ~n17840 & ~n17841;
  assign n17844 = ~n17842 & ~n17843;
  assign n17845 = ~n17470 & ~n17473;
  assign n17846 = n17844 & n17845;
  assign n17847 = ~n17844 & ~n17845;
  assign n17848 = ~n17846 & ~n17847;
  assign n17849 = n5008 & n5413;
  assign n17850 = pi100  & n5241;
  assign n17851 = pi102  & n5006;
  assign n17852 = pi101  & n5001;
  assign n17853 = ~n17851 & ~n17852;
  assign n17854 = ~n17850 & n17853;
  assign n17855 = ~n17849 & n17854;
  assign n17856 = pi38  & ~n17855;
  assign n17857 = pi38  & ~n17856;
  assign n17858 = ~n17855 & ~n17856;
  assign n17859 = ~n17857 & ~n17858;
  assign n17860 = ~n17848 & n17859;
  assign n17861 = n17848 & ~n17859;
  assign n17862 = ~n17860 & ~n17861;
  assign n17863 = ~n17691 & n17862;
  assign n17864 = n17691 & ~n17862;
  assign n17865 = ~n17863 & ~n17864;
  assign n17866 = ~n17690 & n17865;
  assign n17867 = ~n17690 & ~n17866;
  assign n17868 = n17865 & ~n17866;
  assign n17869 = ~n17867 & ~n17868;
  assign n17870 = n17679 & ~n17869;
  assign n17871 = n17679 & ~n17870;
  assign n17872 = ~n17869 & ~n17870;
  assign n17873 = ~n17871 & ~n17872;
  assign n17874 = n17664 & ~n17873;
  assign n17875 = ~n17664 & n17873;
  assign n17876 = ~n17874 & ~n17875;
  assign n17877 = n17649 & n17876;
  assign n17878 = n17649 & ~n17877;
  assign n17879 = n17876 & ~n17877;
  assign n17880 = ~n17878 & ~n17879;
  assign n17881 = ~n17277 & ~n17515;
  assign n17882 = pi115  & n2180;
  assign n17883 = pi117  & n2041;
  assign n17884 = pi116  & n2036;
  assign n17885 = ~n17883 & ~n17884;
  assign n17886 = ~n17882 & n17885;
  assign n17887 = ~n2043 & n17886;
  assign n17888 = ~n9958 & n17886;
  assign n17889 = ~n17887 & ~n17888;
  assign n17890 = pi23  & ~n17889;
  assign n17891 = ~pi23  & n17889;
  assign n17892 = ~n17890 & ~n17891;
  assign n17893 = ~n17881 & ~n17892;
  assign n17894 = ~n17881 & ~n17893;
  assign n17895 = ~n17892 & ~n17893;
  assign n17896 = ~n17894 & ~n17895;
  assign n17897 = ~n17880 & ~n17896;
  assign n17898 = ~n17880 & ~n17897;
  assign n17899 = ~n17896 & ~n17897;
  assign n17900 = ~n17898 & ~n17899;
  assign n17901 = ~n17634 & ~n17900;
  assign n17902 = ~n17634 & ~n17901;
  assign n17903 = ~n17900 & ~n17901;
  assign n17904 = ~n17902 & ~n17903;
  assign n17905 = n17618 & ~n17904;
  assign n17906 = ~n17618 & n17904;
  assign n17907 = ~n17905 & ~n17906;
  assign n17908 = n17603 & n17907;
  assign n17909 = n17603 & ~n17908;
  assign n17910 = n17907 & ~n17908;
  assign n17911 = ~n17909 & ~n17910;
  assign n17912 = ~n17588 & n17911;
  assign n17913 = n17588 & ~n17911;
  assign n17914 = ~n17912 & ~n17913;
  assign n17915 = ~n17576 & ~n17914;
  assign n17916 = ~n17576 & ~n17915;
  assign n17917 = ~n17914 & ~n17915;
  assign n17918 = ~n17916 & ~n17917;
  assign n17919 = ~n17575 & ~n17918;
  assign n17920 = n17575 & n17918;
  assign po74  = ~n17919 & ~n17920;
  assign n17922 = ~n17915 & ~n17919;
  assign n17923 = ~n17588 & ~n17911;
  assign n17924 = ~n17585 & ~n17923;
  assign n17925 = ~n17601 & ~n17908;
  assign n17926 = n938 & n13742;
  assign n17927 = pi125  & n1052;
  assign n17928 = pi127  & n936;
  assign n17929 = pi126  & n931;
  assign n17930 = ~n17928 & ~n17929;
  assign n17931 = ~n17927 & n17930;
  assign n17932 = ~n17926 & n17931;
  assign n17933 = pi14  & ~n17932;
  assign n17934 = pi14  & ~n17933;
  assign n17935 = ~n17932 & ~n17933;
  assign n17936 = ~n17934 & ~n17935;
  assign n17937 = ~n17925 & ~n17936;
  assign n17938 = ~n17925 & ~n17937;
  assign n17939 = ~n17936 & ~n17937;
  assign n17940 = ~n17938 & ~n17939;
  assign n17941 = ~n17617 & ~n17905;
  assign n17942 = n1297 & n12189;
  assign n17943 = pi122  & n1366;
  assign n17944 = pi124  & n1295;
  assign n17945 = pi123  & n1290;
  assign n17946 = ~n17944 & ~n17945;
  assign n17947 = ~n17943 & n17946;
  assign n17948 = ~n17942 & n17947;
  assign n17949 = pi17  & ~n17948;
  assign n17950 = pi17  & ~n17949;
  assign n17951 = ~n17948 & ~n17949;
  assign n17952 = ~n17950 & ~n17951;
  assign n17953 = ~n17941 & n17952;
  assign n17954 = n17941 & ~n17952;
  assign n17955 = ~n17953 & ~n17954;
  assign n17956 = n1611 & n11389;
  assign n17957 = pi119  & n1745;
  assign n17958 = pi121  & n1609;
  assign n17959 = pi120  & n1604;
  assign n17960 = ~n17958 & ~n17959;
  assign n17961 = ~n17957 & n17960;
  assign n17962 = ~n17956 & n17961;
  assign n17963 = pi20  & ~n17962;
  assign n17964 = pi20  & ~n17963;
  assign n17965 = ~n17962 & ~n17963;
  assign n17966 = ~n17964 & ~n17965;
  assign n17967 = ~n17631 & ~n17901;
  assign n17968 = n17966 & n17967;
  assign n17969 = ~n17966 & ~n17967;
  assign n17970 = ~n17968 & ~n17969;
  assign n17971 = ~n17893 & ~n17897;
  assign n17972 = n2043 & n9984;
  assign n17973 = pi116  & n2180;
  assign n17974 = pi118  & n2041;
  assign n17975 = pi117  & n2036;
  assign n17976 = ~n17974 & ~n17975;
  assign n17977 = ~n17973 & n17976;
  assign n17978 = ~n17972 & n17977;
  assign n17979 = pi23  & ~n17978;
  assign n17980 = pi23  & ~n17979;
  assign n17981 = ~n17978 & ~n17979;
  assign n17982 = ~n17980 & ~n17981;
  assign n17983 = ~n17971 & ~n17982;
  assign n17984 = ~n17971 & ~n17983;
  assign n17985 = ~n17982 & ~n17983;
  assign n17986 = ~n17984 & ~n17985;
  assign n17987 = n2523 & n8963;
  assign n17988 = pi113  & n2667;
  assign n17989 = pi115  & n2521;
  assign n17990 = pi114  & n2516;
  assign n17991 = ~n17989 & ~n17990;
  assign n17992 = ~n17988 & n17991;
  assign n17993 = ~n17987 & n17992;
  assign n17994 = pi26  & ~n17993;
  assign n17995 = pi26  & ~n17994;
  assign n17996 = ~n17993 & ~n17994;
  assign n17997 = ~n17995 & ~n17996;
  assign n17998 = ~n17647 & ~n17877;
  assign n17999 = n17997 & n17998;
  assign n18000 = ~n17997 & ~n17998;
  assign n18001 = ~n17999 & ~n18000;
  assign n18002 = ~n17663 & ~n17874;
  assign n18003 = n3034 & n7997;
  assign n18004 = pi110  & n3225;
  assign n18005 = pi112  & n3032;
  assign n18006 = pi111  & n3027;
  assign n18007 = ~n18005 & ~n18006;
  assign n18008 = ~n18004 & n18007;
  assign n18009 = ~n18003 & n18008;
  assign n18010 = pi29  & ~n18009;
  assign n18011 = pi29  & ~n18010;
  assign n18012 = ~n18009 & ~n18010;
  assign n18013 = ~n18011 & ~n18012;
  assign n18014 = ~n18002 & n18013;
  assign n18015 = n18002 & ~n18013;
  assign n18016 = ~n18014 & ~n18015;
  assign n18017 = ~n17863 & ~n17866;
  assign n18018 = ~n17847 & ~n17861;
  assign n18019 = ~n17827 & ~n17841;
  assign n18020 = ~n17810 & ~n17824;
  assign n18021 = ~n17790 & ~n17804;
  assign n18022 = ~n17777 & ~n17781;
  assign n18023 = n2446 & n9310;
  assign n18024 = pi86  & n9701;
  assign n18025 = pi88  & n9308;
  assign n18026 = pi87  & n9303;
  assign n18027 = ~n18025 & ~n18026;
  assign n18028 = ~n18024 & n18027;
  assign n18029 = ~n18023 & n18028;
  assign n18030 = pi53  & ~n18029;
  assign n18031 = pi53  & ~n18030;
  assign n18032 = ~n18029 & ~n18030;
  assign n18033 = ~n18031 & ~n18032;
  assign n18034 = ~n17721 & ~n17725;
  assign n18035 = n1122 & n12627;
  assign n18036 = pi77  & n13004;
  assign n18037 = pi79  & n12625;
  assign n18038 = pi78  & n12620;
  assign n18039 = ~n18037 & ~n18038;
  assign n18040 = ~n18036 & n18039;
  assign n18041 = ~n18035 & n18040;
  assign n18042 = pi62  & ~n18041;
  assign n18043 = pi62  & ~n18042;
  assign n18044 = ~n18041 & ~n18042;
  assign n18045 = ~n18043 & ~n18044;
  assign n18046 = pi75  & n13835;
  assign n18047 = pi76  & ~n13434;
  assign n18048 = ~n18046 & ~n18047;
  assign n18049 = pi11  & ~n17345;
  assign n18050 = ~pi11  & n17345;
  assign n18051 = ~n18049 & ~n18050;
  assign n18052 = ~n18048 & ~n18051;
  assign n18053 = n18048 & n18051;
  assign n18054 = ~n18052 & ~n18053;
  assign n18055 = ~n18045 & n18054;
  assign n18056 = ~n18045 & ~n18055;
  assign n18057 = n18054 & ~n18055;
  assign n18058 = ~n18056 & ~n18057;
  assign n18059 = ~n18034 & ~n18058;
  assign n18060 = ~n18034 & ~n18059;
  assign n18061 = ~n18058 & ~n18059;
  assign n18062 = ~n18060 & ~n18061;
  assign n18063 = n1554 & n11488;
  assign n18064 = pi80  & n11847;
  assign n18065 = pi82  & n11486;
  assign n18066 = pi81  & n11481;
  assign n18067 = ~n18065 & ~n18066;
  assign n18068 = ~n18064 & n18067;
  assign n18069 = ~n18063 & n18068;
  assign n18070 = pi59  & ~n18069;
  assign n18071 = pi59  & ~n18070;
  assign n18072 = ~n18069 & ~n18070;
  assign n18073 = ~n18071 & ~n18072;
  assign n18074 = ~n18062 & ~n18073;
  assign n18075 = ~n18062 & ~n18074;
  assign n18076 = ~n18073 & ~n18074;
  assign n18077 = ~n18075 & ~n18076;
  assign n18078 = ~n17740 & ~n17755;
  assign n18079 = n18077 & n18078;
  assign n18080 = ~n18077 & ~n18078;
  assign n18081 = ~n18079 & ~n18080;
  assign n18082 = n1972 & n10394;
  assign n18083 = pi83  & n10744;
  assign n18084 = pi85  & n10392;
  assign n18085 = pi84  & n10387;
  assign n18086 = ~n18084 & ~n18085;
  assign n18087 = ~n18083 & n18086;
  assign n18088 = ~n18082 & n18087;
  assign n18089 = pi56  & ~n18088;
  assign n18090 = pi56  & ~n18089;
  assign n18091 = ~n18088 & ~n18089;
  assign n18092 = ~n18090 & ~n18091;
  assign n18093 = n18081 & ~n18092;
  assign n18094 = n18081 & ~n18093;
  assign n18095 = ~n18092 & ~n18093;
  assign n18096 = ~n18094 & ~n18095;
  assign n18097 = ~n17761 & ~n17775;
  assign n18098 = ~n18096 & ~n18097;
  assign n18099 = n18096 & n18097;
  assign n18100 = ~n18098 & ~n18099;
  assign n18101 = ~n18033 & n18100;
  assign n18102 = ~n18033 & ~n18101;
  assign n18103 = n18100 & ~n18101;
  assign n18104 = ~n18102 & ~n18103;
  assign n18105 = ~n18022 & ~n18104;
  assign n18106 = ~n18022 & ~n18105;
  assign n18107 = ~n18104 & ~n18105;
  assign n18108 = ~n18106 & ~n18107;
  assign n18109 = n2978 & n8334;
  assign n18110 = pi89  & n8685;
  assign n18111 = pi91  & n8332;
  assign n18112 = pi90  & n8327;
  assign n18113 = ~n18111 & ~n18112;
  assign n18114 = ~n18110 & n18113;
  assign n18115 = ~n18109 & n18114;
  assign n18116 = pi50  & ~n18115;
  assign n18117 = pi50  & ~n18116;
  assign n18118 = ~n18115 & ~n18116;
  assign n18119 = ~n18117 & ~n18118;
  assign n18120 = ~n18108 & ~n18119;
  assign n18121 = ~n18108 & ~n18120;
  assign n18122 = ~n18119 & ~n18120;
  assign n18123 = ~n18121 & ~n18122;
  assign n18124 = ~n17784 & ~n17787;
  assign n18125 = n18123 & n18124;
  assign n18126 = ~n18123 & ~n18124;
  assign n18127 = ~n18125 & ~n18126;
  assign n18128 = n3565 & n7408;
  assign n18129 = pi92  & n7740;
  assign n18130 = pi94  & n7406;
  assign n18131 = pi93  & n7401;
  assign n18132 = ~n18130 & ~n18131;
  assign n18133 = ~n18129 & n18132;
  assign n18134 = ~n18128 & n18133;
  assign n18135 = pi47  & ~n18134;
  assign n18136 = pi47  & ~n18135;
  assign n18137 = ~n18134 & ~n18135;
  assign n18138 = ~n18136 & ~n18137;
  assign n18139 = ~n18127 & n18138;
  assign n18140 = n18127 & ~n18138;
  assign n18141 = ~n18021 & ~n18139;
  assign n18142 = ~n18140 & n18141;
  assign n18143 = ~n18021 & ~n18142;
  assign n18144 = ~n18140 & ~n18142;
  assign n18145 = ~n18139 & n18144;
  assign n18146 = ~n18143 & ~n18145;
  assign n18147 = n4211 & n6539;
  assign n18148 = pi95  & n6873;
  assign n18149 = pi97  & n6537;
  assign n18150 = pi96  & n6532;
  assign n18151 = ~n18149 & ~n18150;
  assign n18152 = ~n18148 & n18151;
  assign n18153 = ~n18147 & n18152;
  assign n18154 = pi44  & ~n18153;
  assign n18155 = pi44  & ~n18154;
  assign n18156 = ~n18153 & ~n18154;
  assign n18157 = ~n18155 & ~n18156;
  assign n18158 = ~n18146 & ~n18157;
  assign n18159 = ~n18146 & ~n18158;
  assign n18160 = ~n18157 & ~n18158;
  assign n18161 = ~n18159 & ~n18160;
  assign n18162 = ~n18020 & n18161;
  assign n18163 = n18020 & ~n18161;
  assign n18164 = ~n18162 & ~n18163;
  assign n18165 = n4910 & n5739;
  assign n18166 = pi98  & n6030;
  assign n18167 = pi100  & n5737;
  assign n18168 = pi99  & n5732;
  assign n18169 = ~n18167 & ~n18168;
  assign n18170 = ~n18166 & n18169;
  assign n18171 = ~n18165 & n18170;
  assign n18172 = pi41  & ~n18171;
  assign n18173 = pi41  & ~n18172;
  assign n18174 = ~n18171 & ~n18172;
  assign n18175 = ~n18173 & ~n18174;
  assign n18176 = ~n18164 & ~n18175;
  assign n18177 = n18164 & n18175;
  assign n18178 = ~n18176 & ~n18177;
  assign n18179 = n18019 & ~n18178;
  assign n18180 = ~n18019 & n18178;
  assign n18181 = ~n18179 & ~n18180;
  assign n18182 = n5008 & n5664;
  assign n18183 = pi101  & n5241;
  assign n18184 = pi103  & n5006;
  assign n18185 = pi102  & n5001;
  assign n18186 = ~n18184 & ~n18185;
  assign n18187 = ~n18183 & n18186;
  assign n18188 = ~n18182 & n18187;
  assign n18189 = pi38  & ~n18188;
  assign n18190 = pi38  & ~n18189;
  assign n18191 = ~n18188 & ~n18189;
  assign n18192 = ~n18190 & ~n18191;
  assign n18193 = n18181 & ~n18192;
  assign n18194 = n18181 & ~n18193;
  assign n18195 = ~n18192 & ~n18193;
  assign n18196 = ~n18194 & ~n18195;
  assign n18197 = ~n18018 & n18196;
  assign n18198 = n18018 & ~n18196;
  assign n18199 = ~n18197 & ~n18198;
  assign n18200 = n4271 & n6477;
  assign n18201 = pi104  & n4503;
  assign n18202 = pi106  & n4269;
  assign n18203 = pi105  & n4264;
  assign n18204 = ~n18202 & ~n18203;
  assign n18205 = ~n18201 & n18204;
  assign n18206 = ~n18200 & n18205;
  assign n18207 = pi35  & ~n18206;
  assign n18208 = pi35  & ~n18207;
  assign n18209 = ~n18206 & ~n18207;
  assign n18210 = ~n18208 & ~n18209;
  assign n18211 = ~n18199 & ~n18210;
  assign n18212 = n18199 & n18210;
  assign n18213 = ~n18211 & ~n18212;
  assign n18214 = n18017 & ~n18213;
  assign n18215 = ~n18017 & n18213;
  assign n18216 = ~n18214 & ~n18215;
  assign n18217 = ~n17677 & ~n17870;
  assign n18218 = n3622 & n7349;
  assign n18219 = pi107  & n3814;
  assign n18220 = pi109  & n3620;
  assign n18221 = pi108  & n3615;
  assign n18222 = ~n18220 & ~n18221;
  assign n18223 = ~n18219 & n18222;
  assign n18224 = ~n18218 & n18223;
  assign n18225 = pi32  & ~n18224;
  assign n18226 = pi32  & ~n18225;
  assign n18227 = ~n18224 & ~n18225;
  assign n18228 = ~n18226 & ~n18227;
  assign n18229 = ~n18217 & ~n18228;
  assign n18230 = ~n18217 & ~n18229;
  assign n18231 = ~n18228 & ~n18229;
  assign n18232 = ~n18230 & ~n18231;
  assign n18233 = n18216 & ~n18232;
  assign n18234 = ~n18216 & n18232;
  assign n18235 = ~n18233 & ~n18234;
  assign n18236 = ~n18016 & n18235;
  assign n18237 = ~n18016 & ~n18236;
  assign n18238 = n18235 & ~n18236;
  assign n18239 = ~n18237 & ~n18238;
  assign n18240 = n18001 & ~n18239;
  assign n18241 = ~n18001 & n18239;
  assign n18242 = ~n18240 & ~n18241;
  assign n18243 = ~n17986 & n18242;
  assign n18244 = ~n17986 & ~n18243;
  assign n18245 = n18242 & ~n18243;
  assign n18246 = ~n18244 & ~n18245;
  assign n18247 = n17970 & ~n18246;
  assign n18248 = ~n17970 & n18246;
  assign n18249 = ~n18247 & ~n18248;
  assign n18250 = ~n17955 & n18249;
  assign n18251 = ~n17955 & ~n18250;
  assign n18252 = n18249 & ~n18250;
  assign n18253 = ~n18251 & ~n18252;
  assign n18254 = ~n17940 & n18253;
  assign n18255 = n17940 & ~n18253;
  assign n18256 = ~n18254 & ~n18255;
  assign n18257 = ~n17924 & ~n18256;
  assign n18258 = ~n17924 & ~n18257;
  assign n18259 = ~n18256 & ~n18257;
  assign n18260 = ~n18258 & ~n18259;
  assign n18261 = ~n17922 & ~n18260;
  assign n18262 = n17922 & n18260;
  assign po75  = ~n18261 & ~n18262;
  assign n18264 = ~n18257 & ~n18261;
  assign n18265 = ~n17940 & ~n18253;
  assign n18266 = ~n17937 & ~n18265;
  assign n18267 = n1297 & n12943;
  assign n18268 = pi123  & n1366;
  assign n18269 = pi125  & n1295;
  assign n18270 = pi124  & n1290;
  assign n18271 = ~n18269 & ~n18270;
  assign n18272 = ~n18268 & n18271;
  assign n18273 = ~n18267 & n18272;
  assign n18274 = pi17  & ~n18273;
  assign n18275 = pi17  & ~n18274;
  assign n18276 = ~n18273 & ~n18274;
  assign n18277 = ~n18275 & ~n18276;
  assign n18278 = ~n17969 & ~n18247;
  assign n18279 = ~n18277 & ~n18278;
  assign n18280 = ~n18277 & ~n18279;
  assign n18281 = ~n18278 & ~n18279;
  assign n18282 = ~n18280 & ~n18281;
  assign n18283 = n2043 & n10667;
  assign n18284 = pi117  & n2180;
  assign n18285 = pi119  & n2041;
  assign n18286 = pi118  & n2036;
  assign n18287 = ~n18285 & ~n18286;
  assign n18288 = ~n18284 & n18287;
  assign n18289 = ~n18283 & n18288;
  assign n18290 = pi23  & ~n18289;
  assign n18291 = pi23  & ~n18290;
  assign n18292 = ~n18289 & ~n18290;
  assign n18293 = ~n18291 & ~n18292;
  assign n18294 = ~n18000 & ~n18240;
  assign n18295 = ~n18293 & ~n18294;
  assign n18296 = ~n18293 & ~n18295;
  assign n18297 = ~n18294 & ~n18295;
  assign n18298 = ~n18296 & ~n18297;
  assign n18299 = n3034 & n8612;
  assign n18300 = pi111  & n3225;
  assign n18301 = pi113  & n3032;
  assign n18302 = pi112  & n3027;
  assign n18303 = ~n18301 & ~n18302;
  assign n18304 = ~n18300 & n18303;
  assign n18305 = ~n18299 & n18304;
  assign n18306 = pi29  & ~n18305;
  assign n18307 = pi29  & ~n18306;
  assign n18308 = ~n18305 & ~n18306;
  assign n18309 = ~n18307 & ~n18308;
  assign n18310 = ~n18229 & ~n18233;
  assign n18311 = ~n18309 & ~n18310;
  assign n18312 = ~n18309 & ~n18311;
  assign n18313 = ~n18310 & ~n18311;
  assign n18314 = ~n18312 & ~n18313;
  assign n18315 = ~n18018 & ~n18196;
  assign n18316 = ~n18193 & ~n18315;
  assign n18317 = n5008 & n5943;
  assign n18318 = pi102  & n5241;
  assign n18319 = pi104  & n5006;
  assign n18320 = pi103  & n5001;
  assign n18321 = ~n18319 & ~n18320;
  assign n18322 = ~n18318 & n18321;
  assign n18323 = ~n18317 & n18322;
  assign n18324 = pi38  & ~n18323;
  assign n18325 = pi38  & ~n18324;
  assign n18326 = ~n18323 & ~n18324;
  assign n18327 = ~n18325 & ~n18326;
  assign n18328 = ~n18176 & ~n18180;
  assign n18329 = n5169 & n5739;
  assign n18330 = pi99  & n6030;
  assign n18331 = pi101  & n5737;
  assign n18332 = pi100  & n5732;
  assign n18333 = ~n18331 & ~n18332;
  assign n18334 = ~n18330 & n18333;
  assign n18335 = ~n18329 & n18334;
  assign n18336 = pi41  & ~n18335;
  assign n18337 = pi41  & ~n18336;
  assign n18338 = ~n18335 & ~n18336;
  assign n18339 = ~n18337 & ~n18338;
  assign n18340 = ~n18020 & ~n18161;
  assign n18341 = ~n18158 & ~n18340;
  assign n18342 = n4454 & n6539;
  assign n18343 = pi96  & n6873;
  assign n18344 = pi98  & n6537;
  assign n18345 = pi97  & n6532;
  assign n18346 = ~n18344 & ~n18345;
  assign n18347 = ~n18343 & n18346;
  assign n18348 = ~n18342 & n18347;
  assign n18349 = pi44  & ~n18348;
  assign n18350 = pi44  & ~n18349;
  assign n18351 = ~n18348 & ~n18349;
  assign n18352 = ~n18350 & ~n18351;
  assign n18353 = n3784 & n7408;
  assign n18354 = pi93  & n7740;
  assign n18355 = pi95  & n7406;
  assign n18356 = pi94  & n7401;
  assign n18357 = ~n18355 & ~n18356;
  assign n18358 = ~n18354 & n18357;
  assign n18359 = ~n18353 & n18358;
  assign n18360 = pi47  & ~n18359;
  assign n18361 = pi47  & ~n18360;
  assign n18362 = ~n18359 & ~n18360;
  assign n18363 = ~n18361 & ~n18362;
  assign n18364 = ~n18120 & ~n18126;
  assign n18365 = pi76  & n13835;
  assign n18366 = pi77  & ~n13434;
  assign n18367 = ~n18365 & ~n18366;
  assign n18368 = ~pi11  & ~n17345;
  assign n18369 = ~n18052 & ~n18368;
  assign n18370 = n18367 & ~n18369;
  assign n18371 = n18367 & ~n18370;
  assign n18372 = ~n18369 & ~n18370;
  assign n18373 = ~n18371 & ~n18372;
  assign n18374 = n1225 & n12627;
  assign n18375 = pi78  & n13004;
  assign n18376 = pi80  & n12625;
  assign n18377 = pi79  & n12620;
  assign n18378 = ~n18376 & ~n18377;
  assign n18379 = ~n18375 & n18378;
  assign n18380 = ~n18374 & n18379;
  assign n18381 = pi62  & ~n18380;
  assign n18382 = pi62  & ~n18381;
  assign n18383 = ~n18380 & ~n18381;
  assign n18384 = ~n18382 & ~n18383;
  assign n18385 = ~n18373 & n18384;
  assign n18386 = n18373 & ~n18384;
  assign n18387 = ~n18385 & ~n18386;
  assign n18388 = ~n18055 & ~n18059;
  assign n18389 = n18387 & n18388;
  assign n18390 = ~n18387 & ~n18388;
  assign n18391 = ~n18389 & ~n18390;
  assign n18392 = n1696 & n11488;
  assign n18393 = pi81  & n11847;
  assign n18394 = pi83  & n11486;
  assign n18395 = pi82  & n11481;
  assign n18396 = ~n18394 & ~n18395;
  assign n18397 = ~n18393 & n18396;
  assign n18398 = ~n18392 & n18397;
  assign n18399 = pi59  & ~n18398;
  assign n18400 = pi59  & ~n18399;
  assign n18401 = ~n18398 & ~n18399;
  assign n18402 = ~n18400 & ~n18401;
  assign n18403 = n18391 & ~n18402;
  assign n18404 = n18391 & ~n18403;
  assign n18405 = ~n18402 & ~n18403;
  assign n18406 = ~n18404 & ~n18405;
  assign n18407 = ~n18074 & ~n18080;
  assign n18408 = n18406 & n18407;
  assign n18409 = ~n18406 & ~n18407;
  assign n18410 = ~n18408 & ~n18409;
  assign n18411 = n2133 & n10394;
  assign n18412 = pi84  & n10744;
  assign n18413 = pi86  & n10392;
  assign n18414 = pi85  & n10387;
  assign n18415 = ~n18413 & ~n18414;
  assign n18416 = ~n18412 & n18415;
  assign n18417 = ~n18411 & n18416;
  assign n18418 = pi56  & ~n18417;
  assign n18419 = pi56  & ~n18418;
  assign n18420 = ~n18417 & ~n18418;
  assign n18421 = ~n18419 & ~n18420;
  assign n18422 = n18410 & ~n18421;
  assign n18423 = n18410 & ~n18422;
  assign n18424 = ~n18421 & ~n18422;
  assign n18425 = ~n18423 & ~n18424;
  assign n18426 = ~n18093 & ~n18098;
  assign n18427 = n18425 & n18426;
  assign n18428 = ~n18425 & ~n18426;
  assign n18429 = ~n18427 & ~n18428;
  assign n18430 = n2473 & n9310;
  assign n18431 = pi87  & n9701;
  assign n18432 = pi89  & n9308;
  assign n18433 = pi88  & n9303;
  assign n18434 = ~n18432 & ~n18433;
  assign n18435 = ~n18431 & n18434;
  assign n18436 = ~n18430 & n18435;
  assign n18437 = pi53  & ~n18436;
  assign n18438 = pi53  & ~n18437;
  assign n18439 = ~n18436 & ~n18437;
  assign n18440 = ~n18438 & ~n18439;
  assign n18441 = n18429 & ~n18440;
  assign n18442 = n18429 & ~n18441;
  assign n18443 = ~n18440 & ~n18441;
  assign n18444 = ~n18442 & ~n18443;
  assign n18445 = ~n18101 & ~n18105;
  assign n18446 = n18444 & n18445;
  assign n18447 = ~n18444 & ~n18445;
  assign n18448 = ~n18446 & ~n18447;
  assign n18449 = n3177 & n8334;
  assign n18450 = pi90  & n8685;
  assign n18451 = pi92  & n8332;
  assign n18452 = pi91  & n8327;
  assign n18453 = ~n18451 & ~n18452;
  assign n18454 = ~n18450 & n18453;
  assign n18455 = ~n18449 & n18454;
  assign n18456 = pi50  & ~n18455;
  assign n18457 = pi50  & ~n18456;
  assign n18458 = ~n18455 & ~n18456;
  assign n18459 = ~n18457 & ~n18458;
  assign n18460 = ~n18448 & n18459;
  assign n18461 = n18448 & ~n18459;
  assign n18462 = ~n18460 & ~n18461;
  assign n18463 = ~n18364 & n18462;
  assign n18464 = ~n18364 & ~n18463;
  assign n18465 = n18462 & ~n18463;
  assign n18466 = ~n18464 & ~n18465;
  assign n18467 = ~n18363 & ~n18466;
  assign n18468 = n18363 & n18466;
  assign n18469 = ~n18467 & ~n18468;
  assign n18470 = ~n18144 & n18469;
  assign n18471 = n18144 & ~n18469;
  assign n18472 = ~n18470 & ~n18471;
  assign n18473 = ~n18352 & n18472;
  assign n18474 = n18352 & ~n18472;
  assign n18475 = ~n18473 & ~n18474;
  assign n18476 = ~n18341 & n18475;
  assign n18477 = ~n18341 & ~n18476;
  assign n18478 = n18475 & ~n18476;
  assign n18479 = ~n18477 & ~n18478;
  assign n18480 = ~n18339 & ~n18479;
  assign n18481 = n18339 & n18479;
  assign n18482 = ~n18480 & ~n18481;
  assign n18483 = ~n18328 & n18482;
  assign n18484 = ~n18328 & ~n18483;
  assign n18485 = n18482 & ~n18483;
  assign n18486 = ~n18484 & ~n18485;
  assign n18487 = ~n18327 & ~n18486;
  assign n18488 = n18327 & n18486;
  assign n18489 = ~n18487 & ~n18488;
  assign n18490 = ~n18316 & n18489;
  assign n18491 = n18316 & ~n18489;
  assign n18492 = ~n18490 & ~n18491;
  assign n18493 = n4271 & n6775;
  assign n18494 = pi105  & n4503;
  assign n18495 = pi107  & n4269;
  assign n18496 = pi106  & n4264;
  assign n18497 = ~n18495 & ~n18496;
  assign n18498 = ~n18494 & n18497;
  assign n18499 = ~n18493 & n18498;
  assign n18500 = pi35  & ~n18499;
  assign n18501 = pi35  & ~n18500;
  assign n18502 = ~n18499 & ~n18500;
  assign n18503 = ~n18501 & ~n18502;
  assign n18504 = n18492 & ~n18503;
  assign n18505 = n18492 & ~n18504;
  assign n18506 = ~n18503 & ~n18504;
  assign n18507 = ~n18505 & ~n18506;
  assign n18508 = ~n18211 & ~n18215;
  assign n18509 = pi108  & n3814;
  assign n18510 = pi110  & n3620;
  assign n18511 = pi109  & n3615;
  assign n18512 = ~n18510 & ~n18511;
  assign n18513 = ~n18509 & n18512;
  assign n18514 = ~n3622 & n18513;
  assign n18515 = ~n7665 & n18513;
  assign n18516 = ~n18514 & ~n18515;
  assign n18517 = pi32  & ~n18516;
  assign n18518 = ~pi32  & n18516;
  assign n18519 = ~n18517 & ~n18518;
  assign n18520 = ~n18508 & ~n18519;
  assign n18521 = ~n18508 & ~n18520;
  assign n18522 = ~n18519 & ~n18520;
  assign n18523 = ~n18521 & ~n18522;
  assign n18524 = ~n18507 & ~n18523;
  assign n18525 = ~n18507 & ~n18524;
  assign n18526 = ~n18523 & ~n18524;
  assign n18527 = ~n18525 & ~n18526;
  assign n18528 = ~n18314 & ~n18527;
  assign n18529 = ~n18314 & ~n18528;
  assign n18530 = ~n18527 & ~n18528;
  assign n18531 = ~n18529 & ~n18530;
  assign n18532 = ~n18002 & ~n18013;
  assign n18533 = ~n18236 & ~n18532;
  assign n18534 = pi114  & n2667;
  assign n18535 = pi116  & n2521;
  assign n18536 = pi115  & n2516;
  assign n18537 = ~n18535 & ~n18536;
  assign n18538 = ~n18534 & n18537;
  assign n18539 = ~n2523 & n18538;
  assign n18540 = ~n9614 & n18538;
  assign n18541 = ~n18539 & ~n18540;
  assign n18542 = pi26  & ~n18541;
  assign n18543 = ~pi26  & n18541;
  assign n18544 = ~n18542 & ~n18543;
  assign n18545 = ~n18533 & ~n18544;
  assign n18546 = n18533 & n18544;
  assign n18547 = ~n18545 & ~n18546;
  assign n18548 = ~n18531 & n18547;
  assign n18549 = ~n18531 & ~n18548;
  assign n18550 = n18547 & ~n18548;
  assign n18551 = ~n18549 & ~n18550;
  assign n18552 = ~n18298 & ~n18551;
  assign n18553 = ~n18298 & ~n18552;
  assign n18554 = ~n18551 & ~n18552;
  assign n18555 = ~n18553 & ~n18554;
  assign n18556 = ~n17983 & ~n18243;
  assign n18557 = pi120  & n1745;
  assign n18558 = pi122  & n1609;
  assign n18559 = pi121  & n1604;
  assign n18560 = ~n18558 & ~n18559;
  assign n18561 = ~n18557 & n18560;
  assign n18562 = ~n1611 & n18561;
  assign n18563 = ~n11778 & n18561;
  assign n18564 = ~n18562 & ~n18563;
  assign n18565 = pi20  & ~n18564;
  assign n18566 = ~pi20  & n18564;
  assign n18567 = ~n18565 & ~n18566;
  assign n18568 = ~n18556 & ~n18567;
  assign n18569 = ~n18556 & ~n18568;
  assign n18570 = ~n18567 & ~n18568;
  assign n18571 = ~n18569 & ~n18570;
  assign n18572 = ~n18555 & ~n18571;
  assign n18573 = ~n18555 & ~n18572;
  assign n18574 = ~n18571 & ~n18572;
  assign n18575 = ~n18573 & ~n18574;
  assign n18576 = ~n18282 & ~n18575;
  assign n18577 = ~n18282 & ~n18576;
  assign n18578 = ~n18575 & ~n18576;
  assign n18579 = ~n18577 & ~n18578;
  assign n18580 = ~n17941 & ~n17952;
  assign n18581 = ~n18250 & ~n18580;
  assign n18582 = pi126  & n1052;
  assign n18583 = pi127  & n931;
  assign n18584 = ~n18582 & ~n18583;
  assign n18585 = ~n938 & n18584;
  assign n18586 = n13773 & n18584;
  assign n18587 = ~n18585 & ~n18586;
  assign n18588 = pi14  & ~n18587;
  assign n18589 = ~pi14  & n18587;
  assign n18590 = ~n18588 & ~n18589;
  assign n18591 = ~n18581 & ~n18590;
  assign n18592 = ~n18581 & ~n18591;
  assign n18593 = ~n18590 & ~n18591;
  assign n18594 = ~n18592 & ~n18593;
  assign n18595 = ~n18579 & ~n18594;
  assign n18596 = n18579 & n18594;
  assign n18597 = ~n18595 & ~n18596;
  assign n18598 = ~n18266 & n18597;
  assign n18599 = ~n18266 & ~n18598;
  assign n18600 = n18597 & ~n18598;
  assign n18601 = ~n18599 & ~n18600;
  assign n18602 = ~n18264 & ~n18601;
  assign n18603 = n18264 & n18601;
  assign po76  = ~n18602 & ~n18603;
  assign n18605 = ~n18598 & ~n18602;
  assign n18606 = ~n18591 & ~n18595;
  assign n18607 = ~n18279 & ~n18576;
  assign n18608 = pi127  & n1052;
  assign n18609 = n938 & n13770;
  assign n18610 = ~n18608 & ~n18609;
  assign n18611 = pi14  & ~n18610;
  assign n18612 = pi14  & ~n18611;
  assign n18613 = ~n18610 & ~n18611;
  assign n18614 = ~n18612 & ~n18613;
  assign n18615 = ~n18607 & ~n18614;
  assign n18616 = ~n18607 & ~n18615;
  assign n18617 = ~n18614 & ~n18615;
  assign n18618 = ~n18616 & ~n18617;
  assign n18619 = n1611 & n12158;
  assign n18620 = pi121  & n1745;
  assign n18621 = pi123  & n1609;
  assign n18622 = pi122  & n1604;
  assign n18623 = ~n18621 & ~n18622;
  assign n18624 = ~n18620 & n18623;
  assign n18625 = ~n18619 & n18624;
  assign n18626 = pi20  & ~n18625;
  assign n18627 = pi20  & ~n18626;
  assign n18628 = ~n18625 & ~n18626;
  assign n18629 = ~n18627 & ~n18628;
  assign n18630 = ~n18295 & ~n18552;
  assign n18631 = n18629 & n18630;
  assign n18632 = ~n18629 & ~n18630;
  assign n18633 = ~n18631 & ~n18632;
  assign n18634 = n2043 & n11028;
  assign n18635 = pi118  & n2180;
  assign n18636 = pi120  & n2041;
  assign n18637 = pi119  & n2036;
  assign n18638 = ~n18636 & ~n18637;
  assign n18639 = ~n18635 & n18638;
  assign n18640 = ~n18634 & n18639;
  assign n18641 = pi23  & ~n18640;
  assign n18642 = pi23  & ~n18641;
  assign n18643 = ~n18640 & ~n18641;
  assign n18644 = ~n18642 & ~n18643;
  assign n18645 = ~n18545 & ~n18548;
  assign n18646 = n18644 & n18645;
  assign n18647 = ~n18644 & ~n18645;
  assign n18648 = ~n18646 & ~n18647;
  assign n18649 = n2523 & n9958;
  assign n18650 = pi115  & n2667;
  assign n18651 = pi117  & n2521;
  assign n18652 = pi116  & n2516;
  assign n18653 = ~n18651 & ~n18652;
  assign n18654 = ~n18650 & n18653;
  assign n18655 = ~n18649 & n18654;
  assign n18656 = pi26  & ~n18655;
  assign n18657 = pi26  & ~n18656;
  assign n18658 = ~n18655 & ~n18656;
  assign n18659 = ~n18657 & ~n18658;
  assign n18660 = ~n18311 & ~n18528;
  assign n18661 = n18659 & n18660;
  assign n18662 = ~n18659 & ~n18660;
  assign n18663 = ~n18661 & ~n18662;
  assign n18664 = ~n18490 & ~n18504;
  assign n18665 = pi109  & n3814;
  assign n18666 = pi111  & n3620;
  assign n18667 = pi110  & n3615;
  assign n18668 = ~n18666 & ~n18667;
  assign n18669 = ~n18665 & n18668;
  assign n18670 = ~n3622 & n18669;
  assign n18671 = ~n7970 & n18669;
  assign n18672 = ~n18670 & ~n18671;
  assign n18673 = pi32  & ~n18672;
  assign n18674 = ~pi32  & n18672;
  assign n18675 = ~n18673 & ~n18674;
  assign n18676 = ~n18664 & ~n18675;
  assign n18677 = n18664 & n18675;
  assign n18678 = ~n18676 & ~n18677;
  assign n18679 = n4271 & n7060;
  assign n18680 = pi106  & n4503;
  assign n18681 = pi108  & n4269;
  assign n18682 = pi107  & n4264;
  assign n18683 = ~n18681 & ~n18682;
  assign n18684 = ~n18680 & n18683;
  assign n18685 = ~n18679 & n18684;
  assign n18686 = pi35  & ~n18685;
  assign n18687 = pi35  & ~n18686;
  assign n18688 = ~n18685 & ~n18686;
  assign n18689 = ~n18687 & ~n18688;
  assign n18690 = ~n18483 & ~n18487;
  assign n18691 = n5008 & n6207;
  assign n18692 = pi103  & n5241;
  assign n18693 = pi105  & n5006;
  assign n18694 = pi104  & n5001;
  assign n18695 = ~n18693 & ~n18694;
  assign n18696 = ~n18692 & n18695;
  assign n18697 = ~n18691 & n18696;
  assign n18698 = pi38  & ~n18697;
  assign n18699 = pi38  & ~n18698;
  assign n18700 = ~n18697 & ~n18698;
  assign n18701 = ~n18699 & ~n18700;
  assign n18702 = ~n18476 & ~n18480;
  assign n18703 = ~n18463 & ~n18467;
  assign n18704 = ~n18428 & ~n18441;
  assign n18705 = n2801 & n9310;
  assign n18706 = pi88  & n9701;
  assign n18707 = pi90  & n9308;
  assign n18708 = pi89  & n9303;
  assign n18709 = ~n18707 & ~n18708;
  assign n18710 = ~n18706 & n18709;
  assign n18711 = ~n18705 & n18710;
  assign n18712 = pi53  & ~n18711;
  assign n18713 = pi53  & ~n18712;
  assign n18714 = ~n18711 & ~n18712;
  assign n18715 = ~n18713 & ~n18714;
  assign n18716 = ~n18409 & ~n18422;
  assign n18717 = ~n18373 & ~n18384;
  assign n18718 = ~n18370 & ~n18717;
  assign n18719 = pi77  & n13835;
  assign n18720 = pi78  & ~n13434;
  assign n18721 = ~n18719 & ~n18720;
  assign n18722 = n18367 & ~n18721;
  assign n18723 = ~n18367 & n18721;
  assign n18724 = ~n18722 & ~n18723;
  assign n18725 = pi79  & n13004;
  assign n18726 = pi81  & n12625;
  assign n18727 = pi80  & n12620;
  assign n18728 = ~n18726 & ~n18727;
  assign n18729 = ~n18725 & n18728;
  assign n18730 = ~n12627 & n18729;
  assign n18731 = ~n1434 & n18729;
  assign n18732 = ~n18730 & ~n18731;
  assign n18733 = pi62  & ~n18732;
  assign n18734 = ~pi62  & n18732;
  assign n18735 = ~n18733 & ~n18734;
  assign n18736 = n18724 & ~n18735;
  assign n18737 = ~n18724 & n18735;
  assign n18738 = ~n18736 & ~n18737;
  assign n18739 = ~n18718 & n18738;
  assign n18740 = n18718 & ~n18738;
  assign n18741 = ~n18739 & ~n18740;
  assign n18742 = n1834 & n11488;
  assign n18743 = pi82  & n11847;
  assign n18744 = pi84  & n11486;
  assign n18745 = pi83  & n11481;
  assign n18746 = ~n18744 & ~n18745;
  assign n18747 = ~n18743 & n18746;
  assign n18748 = ~n18742 & n18747;
  assign n18749 = pi59  & ~n18748;
  assign n18750 = pi59  & ~n18749;
  assign n18751 = ~n18748 & ~n18749;
  assign n18752 = ~n18750 & ~n18751;
  assign n18753 = n18741 & ~n18752;
  assign n18754 = n18741 & ~n18753;
  assign n18755 = ~n18752 & ~n18753;
  assign n18756 = ~n18754 & ~n18755;
  assign n18757 = ~n18390 & ~n18403;
  assign n18758 = n18756 & n18757;
  assign n18759 = ~n18756 & ~n18757;
  assign n18760 = ~n18758 & ~n18759;
  assign n18761 = n2288 & n10394;
  assign n18762 = pi85  & n10744;
  assign n18763 = pi87  & n10392;
  assign n18764 = pi86  & n10387;
  assign n18765 = ~n18763 & ~n18764;
  assign n18766 = ~n18762 & n18765;
  assign n18767 = ~n18761 & n18766;
  assign n18768 = pi56  & ~n18767;
  assign n18769 = pi56  & ~n18768;
  assign n18770 = ~n18767 & ~n18768;
  assign n18771 = ~n18769 & ~n18770;
  assign n18772 = ~n18760 & n18771;
  assign n18773 = n18760 & ~n18771;
  assign n18774 = ~n18772 & ~n18773;
  assign n18775 = ~n18716 & n18774;
  assign n18776 = n18716 & ~n18774;
  assign n18777 = ~n18775 & ~n18776;
  assign n18778 = ~n18715 & n18777;
  assign n18779 = n18715 & ~n18777;
  assign n18780 = ~n18778 & ~n18779;
  assign n18781 = ~n18704 & n18780;
  assign n18782 = n18704 & ~n18780;
  assign n18783 = ~n18781 & ~n18782;
  assign n18784 = n3371 & n8334;
  assign n18785 = pi91  & n8685;
  assign n18786 = pi93  & n8332;
  assign n18787 = pi92  & n8327;
  assign n18788 = ~n18786 & ~n18787;
  assign n18789 = ~n18785 & n18788;
  assign n18790 = ~n18784 & n18789;
  assign n18791 = pi50  & ~n18790;
  assign n18792 = pi50  & ~n18791;
  assign n18793 = ~n18790 & ~n18791;
  assign n18794 = ~n18792 & ~n18793;
  assign n18795 = n18783 & ~n18794;
  assign n18796 = n18783 & ~n18795;
  assign n18797 = ~n18794 & ~n18795;
  assign n18798 = ~n18796 & ~n18797;
  assign n18799 = ~n18447 & ~n18461;
  assign n18800 = ~n18798 & ~n18799;
  assign n18801 = ~n18798 & ~n18800;
  assign n18802 = ~n18799 & ~n18800;
  assign n18803 = ~n18801 & ~n18802;
  assign n18804 = n4001 & n7408;
  assign n18805 = pi94  & n7740;
  assign n18806 = pi96  & n7406;
  assign n18807 = pi95  & n7401;
  assign n18808 = ~n18806 & ~n18807;
  assign n18809 = ~n18805 & n18808;
  assign n18810 = ~n18804 & n18809;
  assign n18811 = pi47  & ~n18810;
  assign n18812 = pi47  & ~n18811;
  assign n18813 = ~n18810 & ~n18811;
  assign n18814 = ~n18812 & ~n18813;
  assign n18815 = ~n18803 & n18814;
  assign n18816 = n18803 & ~n18814;
  assign n18817 = ~n18815 & ~n18816;
  assign n18818 = n18703 & n18817;
  assign n18819 = ~n18703 & ~n18817;
  assign n18820 = ~n18818 & ~n18819;
  assign n18821 = n4684 & n6539;
  assign n18822 = pi97  & n6873;
  assign n18823 = pi99  & n6537;
  assign n18824 = pi98  & n6532;
  assign n18825 = ~n18823 & ~n18824;
  assign n18826 = ~n18822 & n18825;
  assign n18827 = ~n18821 & n18826;
  assign n18828 = pi44  & ~n18827;
  assign n18829 = pi44  & ~n18828;
  assign n18830 = ~n18827 & ~n18828;
  assign n18831 = ~n18829 & ~n18830;
  assign n18832 = n18820 & ~n18831;
  assign n18833 = n18820 & ~n18832;
  assign n18834 = ~n18831 & ~n18832;
  assign n18835 = ~n18833 & ~n18834;
  assign n18836 = ~n18470 & ~n18473;
  assign n18837 = n18835 & n18836;
  assign n18838 = ~n18835 & ~n18836;
  assign n18839 = ~n18837 & ~n18838;
  assign n18840 = n5413 & n5739;
  assign n18841 = pi100  & n6030;
  assign n18842 = pi102  & n5737;
  assign n18843 = pi101  & n5732;
  assign n18844 = ~n18842 & ~n18843;
  assign n18845 = ~n18841 & n18844;
  assign n18846 = ~n18840 & n18845;
  assign n18847 = pi41  & ~n18846;
  assign n18848 = pi41  & ~n18847;
  assign n18849 = ~n18846 & ~n18847;
  assign n18850 = ~n18848 & ~n18849;
  assign n18851 = ~n18839 & n18850;
  assign n18852 = n18839 & ~n18850;
  assign n18853 = ~n18851 & ~n18852;
  assign n18854 = ~n18702 & n18853;
  assign n18855 = n18702 & ~n18853;
  assign n18856 = ~n18854 & ~n18855;
  assign n18857 = ~n18701 & n18856;
  assign n18858 = n18701 & ~n18856;
  assign n18859 = ~n18857 & ~n18858;
  assign n18860 = ~n18690 & n18859;
  assign n18861 = n18690 & ~n18859;
  assign n18862 = ~n18860 & ~n18861;
  assign n18863 = ~n18689 & n18862;
  assign n18864 = ~n18689 & ~n18863;
  assign n18865 = n18862 & ~n18863;
  assign n18866 = ~n18864 & ~n18865;
  assign n18867 = n18678 & ~n18866;
  assign n18868 = n18678 & ~n18867;
  assign n18869 = ~n18866 & ~n18867;
  assign n18870 = ~n18868 & ~n18869;
  assign n18871 = ~n18520 & ~n18524;
  assign n18872 = pi112  & n3225;
  assign n18873 = pi114  & n3032;
  assign n18874 = pi113  & n3027;
  assign n18875 = ~n18873 & ~n18874;
  assign n18876 = ~n18872 & n18875;
  assign n18877 = ~n3034 & n18876;
  assign n18878 = ~n8936 & n18876;
  assign n18879 = ~n18877 & ~n18878;
  assign n18880 = pi29  & ~n18879;
  assign n18881 = ~pi29  & n18879;
  assign n18882 = ~n18880 & ~n18881;
  assign n18883 = ~n18871 & ~n18882;
  assign n18884 = n18871 & n18882;
  assign n18885 = ~n18883 & ~n18884;
  assign n18886 = ~n18870 & n18885;
  assign n18887 = ~n18870 & ~n18886;
  assign n18888 = n18885 & ~n18886;
  assign n18889 = ~n18887 & ~n18888;
  assign n18890 = n18663 & ~n18889;
  assign n18891 = n18663 & ~n18890;
  assign n18892 = ~n18889 & ~n18890;
  assign n18893 = ~n18891 & ~n18892;
  assign n18894 = n18648 & ~n18893;
  assign n18895 = ~n18648 & n18893;
  assign n18896 = ~n18894 & ~n18895;
  assign n18897 = n18633 & n18896;
  assign n18898 = n18633 & ~n18897;
  assign n18899 = n18896 & ~n18897;
  assign n18900 = ~n18898 & ~n18899;
  assign n18901 = ~n18568 & ~n18572;
  assign n18902 = pi124  & n1366;
  assign n18903 = pi126  & n1295;
  assign n18904 = pi125  & n1290;
  assign n18905 = ~n18903 & ~n18904;
  assign n18906 = ~n18902 & n18905;
  assign n18907 = ~n1297 & n18906;
  assign n18908 = ~n13344 & n18906;
  assign n18909 = ~n18907 & ~n18908;
  assign n18910 = pi17  & ~n18909;
  assign n18911 = ~pi17  & n18909;
  assign n18912 = ~n18910 & ~n18911;
  assign n18913 = ~n18901 & ~n18912;
  assign n18914 = ~n18901 & ~n18913;
  assign n18915 = ~n18912 & ~n18913;
  assign n18916 = ~n18914 & ~n18915;
  assign n18917 = ~n18900 & ~n18916;
  assign n18918 = n18900 & n18916;
  assign n18919 = ~n18917 & ~n18918;
  assign n18920 = ~n18618 & n18919;
  assign n18921 = n18618 & ~n18919;
  assign n18922 = ~n18920 & ~n18921;
  assign n18923 = ~n18606 & n18922;
  assign n18924 = n18606 & ~n18922;
  assign n18925 = ~n18923 & ~n18924;
  assign n18926 = ~n18605 & n18925;
  assign n18927 = n18605 & ~n18925;
  assign po77  = ~n18926 & ~n18927;
  assign n18929 = ~n18913 & ~n18917;
  assign n18930 = n1297 & n13742;
  assign n18931 = pi125  & n1366;
  assign n18932 = pi127  & n1295;
  assign n18933 = pi126  & n1290;
  assign n18934 = ~n18932 & ~n18933;
  assign n18935 = ~n18931 & n18934;
  assign n18936 = ~n18930 & n18935;
  assign n18937 = pi17  & ~n18936;
  assign n18938 = pi17  & ~n18937;
  assign n18939 = ~n18936 & ~n18937;
  assign n18940 = ~n18938 & ~n18939;
  assign n18941 = ~n18929 & ~n18940;
  assign n18942 = ~n18929 & ~n18941;
  assign n18943 = ~n18940 & ~n18941;
  assign n18944 = ~n18942 & ~n18943;
  assign n18945 = n1611 & n12189;
  assign n18946 = pi122  & n1745;
  assign n18947 = pi124  & n1609;
  assign n18948 = pi123  & n1604;
  assign n18949 = ~n18947 & ~n18948;
  assign n18950 = ~n18946 & n18949;
  assign n18951 = ~n18945 & n18950;
  assign n18952 = pi20  & ~n18951;
  assign n18953 = pi20  & ~n18952;
  assign n18954 = ~n18951 & ~n18952;
  assign n18955 = ~n18953 & ~n18954;
  assign n18956 = ~n18632 & ~n18897;
  assign n18957 = n18955 & n18956;
  assign n18958 = ~n18955 & ~n18956;
  assign n18959 = ~n18957 & ~n18958;
  assign n18960 = ~n18647 & ~n18894;
  assign n18961 = n2043 & n11389;
  assign n18962 = pi119  & n2180;
  assign n18963 = pi121  & n2041;
  assign n18964 = pi120  & n2036;
  assign n18965 = ~n18963 & ~n18964;
  assign n18966 = ~n18962 & n18965;
  assign n18967 = ~n18961 & n18966;
  assign n18968 = pi23  & ~n18967;
  assign n18969 = pi23  & ~n18968;
  assign n18970 = ~n18967 & ~n18968;
  assign n18971 = ~n18969 & ~n18970;
  assign n18972 = ~n18960 & n18971;
  assign n18973 = n18960 & ~n18971;
  assign n18974 = ~n18972 & ~n18973;
  assign n18975 = n2523 & n9984;
  assign n18976 = pi116  & n2667;
  assign n18977 = pi118  & n2521;
  assign n18978 = pi117  & n2516;
  assign n18979 = ~n18977 & ~n18978;
  assign n18980 = ~n18976 & n18979;
  assign n18981 = ~n18975 & n18980;
  assign n18982 = pi26  & ~n18981;
  assign n18983 = pi26  & ~n18982;
  assign n18984 = ~n18981 & ~n18982;
  assign n18985 = ~n18983 & ~n18984;
  assign n18986 = ~n18662 & ~n18890;
  assign n18987 = n18985 & n18986;
  assign n18988 = ~n18985 & ~n18986;
  assign n18989 = ~n18987 & ~n18988;
  assign n18990 = n3034 & n8963;
  assign n18991 = pi113  & n3225;
  assign n18992 = pi115  & n3032;
  assign n18993 = pi114  & n3027;
  assign n18994 = ~n18992 & ~n18993;
  assign n18995 = ~n18991 & n18994;
  assign n18996 = ~n18990 & n18995;
  assign n18997 = pi29  & ~n18996;
  assign n18998 = pi29  & ~n18997;
  assign n18999 = ~n18996 & ~n18997;
  assign n19000 = ~n18998 & ~n18999;
  assign n19001 = ~n18883 & ~n18886;
  assign n19002 = n19000 & n19001;
  assign n19003 = ~n19000 & ~n19001;
  assign n19004 = ~n19002 & ~n19003;
  assign n19005 = ~n18854 & ~n18857;
  assign n19006 = ~n18838 & ~n18852;
  assign n19007 = ~n18819 & ~n18832;
  assign n19008 = ~n18803 & ~n18814;
  assign n19009 = ~n18800 & ~n19008;
  assign n19010 = ~n18759 & ~n18773;
  assign n19011 = pi78  & n13835;
  assign n19012 = pi79  & ~n13434;
  assign n19013 = ~n19011 & ~n19012;
  assign n19014 = ~pi14  & ~n19013;
  assign n19015 = ~pi14  & ~n19014;
  assign n19016 = ~n19013 & ~n19014;
  assign n19017 = ~n19015 & ~n19016;
  assign n19018 = ~n18367 & ~n19017;
  assign n19019 = ~n18367 & ~n19018;
  assign n19020 = ~n19017 & ~n19018;
  assign n19021 = ~n19019 & ~n19020;
  assign n19022 = n1554 & n12627;
  assign n19023 = pi80  & n13004;
  assign n19024 = pi82  & n12625;
  assign n19025 = pi81  & n12620;
  assign n19026 = ~n19024 & ~n19025;
  assign n19027 = ~n19023 & n19026;
  assign n19028 = ~n19022 & n19027;
  assign n19029 = pi62  & ~n19028;
  assign n19030 = pi62  & ~n19029;
  assign n19031 = ~n19028 & ~n19029;
  assign n19032 = ~n19030 & ~n19031;
  assign n19033 = ~n19021 & ~n19032;
  assign n19034 = ~n19021 & ~n19033;
  assign n19035 = ~n19032 & ~n19033;
  assign n19036 = ~n19034 & ~n19035;
  assign n19037 = ~n18722 & ~n18736;
  assign n19038 = n19036 & n19037;
  assign n19039 = ~n19036 & ~n19037;
  assign n19040 = ~n19038 & ~n19039;
  assign n19041 = n1972 & n11488;
  assign n19042 = pi83  & n11847;
  assign n19043 = pi85  & n11486;
  assign n19044 = pi84  & n11481;
  assign n19045 = ~n19043 & ~n19044;
  assign n19046 = ~n19042 & n19045;
  assign n19047 = ~n19041 & n19046;
  assign n19048 = pi59  & ~n19047;
  assign n19049 = pi59  & ~n19048;
  assign n19050 = ~n19047 & ~n19048;
  assign n19051 = ~n19049 & ~n19050;
  assign n19052 = n19040 & ~n19051;
  assign n19053 = n19040 & ~n19052;
  assign n19054 = ~n19051 & ~n19052;
  assign n19055 = ~n19053 & ~n19054;
  assign n19056 = ~n18739 & ~n18753;
  assign n19057 = n19055 & n19056;
  assign n19058 = ~n19055 & ~n19056;
  assign n19059 = ~n19057 & ~n19058;
  assign n19060 = n2446 & n10394;
  assign n19061 = pi86  & n10744;
  assign n19062 = pi88  & n10392;
  assign n19063 = pi87  & n10387;
  assign n19064 = ~n19062 & ~n19063;
  assign n19065 = ~n19061 & n19064;
  assign n19066 = ~n19060 & n19065;
  assign n19067 = pi56  & ~n19066;
  assign n19068 = pi56  & ~n19067;
  assign n19069 = ~n19066 & ~n19067;
  assign n19070 = ~n19068 & ~n19069;
  assign n19071 = ~n19059 & n19070;
  assign n19072 = n19059 & ~n19070;
  assign n19073 = ~n19010 & ~n19071;
  assign n19074 = ~n19072 & n19073;
  assign n19075 = ~n19010 & ~n19074;
  assign n19076 = ~n19072 & ~n19074;
  assign n19077 = ~n19071 & n19076;
  assign n19078 = ~n19075 & ~n19077;
  assign n19079 = n2978 & n9310;
  assign n19080 = pi89  & n9701;
  assign n19081 = pi91  & n9308;
  assign n19082 = pi90  & n9303;
  assign n19083 = ~n19081 & ~n19082;
  assign n19084 = ~n19080 & n19083;
  assign n19085 = ~n19079 & n19084;
  assign n19086 = pi53  & ~n19085;
  assign n19087 = pi53  & ~n19086;
  assign n19088 = ~n19085 & ~n19086;
  assign n19089 = ~n19087 & ~n19088;
  assign n19090 = ~n19078 & ~n19089;
  assign n19091 = ~n19078 & ~n19090;
  assign n19092 = ~n19089 & ~n19090;
  assign n19093 = ~n19091 & ~n19092;
  assign n19094 = ~n18775 & ~n18778;
  assign n19095 = n19093 & n19094;
  assign n19096 = ~n19093 & ~n19094;
  assign n19097 = ~n19095 & ~n19096;
  assign n19098 = n3565 & n8334;
  assign n19099 = pi92  & n8685;
  assign n19100 = pi94  & n8332;
  assign n19101 = pi93  & n8327;
  assign n19102 = ~n19100 & ~n19101;
  assign n19103 = ~n19099 & n19102;
  assign n19104 = ~n19098 & n19103;
  assign n19105 = pi50  & ~n19104;
  assign n19106 = pi50  & ~n19105;
  assign n19107 = ~n19104 & ~n19105;
  assign n19108 = ~n19106 & ~n19107;
  assign n19109 = n19097 & ~n19108;
  assign n19110 = n19097 & ~n19109;
  assign n19111 = ~n19108 & ~n19109;
  assign n19112 = ~n19110 & ~n19111;
  assign n19113 = ~n18781 & ~n18795;
  assign n19114 = n19112 & n19113;
  assign n19115 = ~n19112 & ~n19113;
  assign n19116 = ~n19114 & ~n19115;
  assign n19117 = n4211 & n7408;
  assign n19118 = pi95  & n7740;
  assign n19119 = pi97  & n7406;
  assign n19120 = pi96  & n7401;
  assign n19121 = ~n19119 & ~n19120;
  assign n19122 = ~n19118 & n19121;
  assign n19123 = ~n19117 & n19122;
  assign n19124 = pi47  & ~n19123;
  assign n19125 = pi47  & ~n19124;
  assign n19126 = ~n19123 & ~n19124;
  assign n19127 = ~n19125 & ~n19126;
  assign n19128 = n19116 & ~n19127;
  assign n19129 = n19116 & ~n19128;
  assign n19130 = ~n19127 & ~n19128;
  assign n19131 = ~n19129 & ~n19130;
  assign n19132 = ~n19009 & n19131;
  assign n19133 = n19009 & ~n19131;
  assign n19134 = ~n19132 & ~n19133;
  assign n19135 = n4910 & n6539;
  assign n19136 = pi98  & n6873;
  assign n19137 = pi100  & n6537;
  assign n19138 = pi99  & n6532;
  assign n19139 = ~n19137 & ~n19138;
  assign n19140 = ~n19136 & n19139;
  assign n19141 = ~n19135 & n19140;
  assign n19142 = pi44  & ~n19141;
  assign n19143 = pi44  & ~n19142;
  assign n19144 = ~n19141 & ~n19142;
  assign n19145 = ~n19143 & ~n19144;
  assign n19146 = ~n19134 & ~n19145;
  assign n19147 = n19134 & n19145;
  assign n19148 = ~n19146 & ~n19147;
  assign n19149 = n19007 & ~n19148;
  assign n19150 = ~n19007 & n19148;
  assign n19151 = ~n19149 & ~n19150;
  assign n19152 = n5664 & n5739;
  assign n19153 = pi101  & n6030;
  assign n19154 = pi103  & n5737;
  assign n19155 = pi102  & n5732;
  assign n19156 = ~n19154 & ~n19155;
  assign n19157 = ~n19153 & n19156;
  assign n19158 = ~n19152 & n19157;
  assign n19159 = pi41  & ~n19158;
  assign n19160 = pi41  & ~n19159;
  assign n19161 = ~n19158 & ~n19159;
  assign n19162 = ~n19160 & ~n19161;
  assign n19163 = n19151 & ~n19162;
  assign n19164 = n19151 & ~n19163;
  assign n19165 = ~n19162 & ~n19163;
  assign n19166 = ~n19164 & ~n19165;
  assign n19167 = ~n19006 & n19166;
  assign n19168 = n19006 & ~n19166;
  assign n19169 = ~n19167 & ~n19168;
  assign n19170 = n5008 & n6477;
  assign n19171 = pi104  & n5241;
  assign n19172 = pi106  & n5006;
  assign n19173 = pi105  & n5001;
  assign n19174 = ~n19172 & ~n19173;
  assign n19175 = ~n19171 & n19174;
  assign n19176 = ~n19170 & n19175;
  assign n19177 = pi38  & ~n19176;
  assign n19178 = pi38  & ~n19177;
  assign n19179 = ~n19176 & ~n19177;
  assign n19180 = ~n19178 & ~n19179;
  assign n19181 = ~n19169 & ~n19180;
  assign n19182 = n19169 & n19180;
  assign n19183 = ~n19181 & ~n19182;
  assign n19184 = n19005 & ~n19183;
  assign n19185 = ~n19005 & n19183;
  assign n19186 = ~n19184 & ~n19185;
  assign n19187 = n4271 & n7349;
  assign n19188 = pi107  & n4503;
  assign n19189 = pi109  & n4269;
  assign n19190 = pi108  & n4264;
  assign n19191 = ~n19189 & ~n19190;
  assign n19192 = ~n19188 & n19191;
  assign n19193 = ~n19187 & n19192;
  assign n19194 = pi35  & ~n19193;
  assign n19195 = pi35  & ~n19194;
  assign n19196 = ~n19193 & ~n19194;
  assign n19197 = ~n19195 & ~n19196;
  assign n19198 = n19186 & ~n19197;
  assign n19199 = n19186 & ~n19198;
  assign n19200 = ~n19197 & ~n19198;
  assign n19201 = ~n19199 & ~n19200;
  assign n19202 = ~n18860 & ~n18863;
  assign n19203 = n19201 & n19202;
  assign n19204 = ~n19201 & ~n19202;
  assign n19205 = ~n19203 & ~n19204;
  assign n19206 = ~n18676 & ~n18867;
  assign n19207 = n3622 & n7997;
  assign n19208 = pi110  & n3814;
  assign n19209 = pi112  & n3620;
  assign n19210 = pi111  & n3615;
  assign n19211 = ~n19209 & ~n19210;
  assign n19212 = ~n19208 & n19211;
  assign n19213 = ~n19207 & n19212;
  assign n19214 = pi32  & ~n19213;
  assign n19215 = pi32  & ~n19214;
  assign n19216 = ~n19213 & ~n19214;
  assign n19217 = ~n19215 & ~n19216;
  assign n19218 = ~n19206 & ~n19217;
  assign n19219 = ~n19206 & ~n19218;
  assign n19220 = ~n19217 & ~n19218;
  assign n19221 = ~n19219 & ~n19220;
  assign n19222 = n19205 & ~n19221;
  assign n19223 = ~n19205 & n19221;
  assign n19224 = ~n19222 & ~n19223;
  assign n19225 = n19004 & n19224;
  assign n19226 = n19004 & ~n19225;
  assign n19227 = n19224 & ~n19225;
  assign n19228 = ~n19226 & ~n19227;
  assign n19229 = n18989 & ~n19228;
  assign n19230 = ~n18989 & n19228;
  assign n19231 = ~n19229 & ~n19230;
  assign n19232 = ~n18974 & n19231;
  assign n19233 = ~n18974 & ~n19232;
  assign n19234 = n19231 & ~n19232;
  assign n19235 = ~n19233 & ~n19234;
  assign n19236 = n18959 & ~n19235;
  assign n19237 = ~n18959 & n19235;
  assign n19238 = ~n19236 & ~n19237;
  assign n19239 = ~n18944 & n19238;
  assign n19240 = ~n18944 & ~n19239;
  assign n19241 = n19238 & ~n19239;
  assign n19242 = ~n19240 & ~n19241;
  assign n19243 = ~n18615 & ~n18920;
  assign n19244 = n19242 & n19243;
  assign n19245 = ~n19242 & ~n19243;
  assign n19246 = ~n19244 & ~n19245;
  assign n19247 = ~n18923 & ~n18926;
  assign n19248 = n19246 & ~n19247;
  assign n19249 = ~n19246 & n19247;
  assign po78  = ~n19248 & ~n19249;
  assign n19251 = ~n18958 & ~n19236;
  assign n19252 = pi126  & n1366;
  assign n19253 = pi127  & n1290;
  assign n19254 = ~n19252 & ~n19253;
  assign n19255 = ~n1297 & n19254;
  assign n19256 = n13773 & n19254;
  assign n19257 = ~n19255 & ~n19256;
  assign n19258 = pi17  & ~n19257;
  assign n19259 = ~pi17  & n19257;
  assign n19260 = ~n19258 & ~n19259;
  assign n19261 = ~n19251 & ~n19260;
  assign n19262 = n19251 & n19260;
  assign n19263 = ~n19261 & ~n19262;
  assign n19264 = n1611 & n12943;
  assign n19265 = pi123  & n1745;
  assign n19266 = pi125  & n1609;
  assign n19267 = pi124  & n1604;
  assign n19268 = ~n19266 & ~n19267;
  assign n19269 = ~n19265 & n19268;
  assign n19270 = ~n19264 & n19269;
  assign n19271 = pi20  & ~n19270;
  assign n19272 = pi20  & ~n19271;
  assign n19273 = ~n19270 & ~n19271;
  assign n19274 = ~n19272 & ~n19273;
  assign n19275 = ~n18960 & ~n18971;
  assign n19276 = ~n19232 & ~n19275;
  assign n19277 = n19274 & n19276;
  assign n19278 = ~n19274 & ~n19276;
  assign n19279 = ~n19277 & ~n19278;
  assign n19280 = ~n18988 & ~n19229;
  assign n19281 = pi120  & n2180;
  assign n19282 = pi122  & n2041;
  assign n19283 = pi121  & n2036;
  assign n19284 = ~n19282 & ~n19283;
  assign n19285 = ~n19281 & n19284;
  assign n19286 = ~n2043 & n19285;
  assign n19287 = ~n11778 & n19285;
  assign n19288 = ~n19286 & ~n19287;
  assign n19289 = pi23  & ~n19288;
  assign n19290 = ~pi23  & n19288;
  assign n19291 = ~n19289 & ~n19290;
  assign n19292 = ~n19280 & ~n19291;
  assign n19293 = n19280 & n19291;
  assign n19294 = ~n19292 & ~n19293;
  assign n19295 = n2523 & n10667;
  assign n19296 = pi117  & n2667;
  assign n19297 = pi119  & n2521;
  assign n19298 = pi118  & n2516;
  assign n19299 = ~n19297 & ~n19298;
  assign n19300 = ~n19296 & n19299;
  assign n19301 = ~n19295 & n19300;
  assign n19302 = pi26  & ~n19301;
  assign n19303 = pi26  & ~n19302;
  assign n19304 = ~n19301 & ~n19302;
  assign n19305 = ~n19303 & ~n19304;
  assign n19306 = ~n19003 & ~n19225;
  assign n19307 = n19305 & n19306;
  assign n19308 = ~n19305 & ~n19306;
  assign n19309 = ~n19307 & ~n19308;
  assign n19310 = n3034 & n9614;
  assign n19311 = pi114  & n3225;
  assign n19312 = pi116  & n3032;
  assign n19313 = pi115  & n3027;
  assign n19314 = ~n19312 & ~n19313;
  assign n19315 = ~n19311 & n19314;
  assign n19316 = ~n19310 & n19315;
  assign n19317 = pi29  & ~n19316;
  assign n19318 = pi29  & ~n19317;
  assign n19319 = ~n19316 & ~n19317;
  assign n19320 = ~n19318 & ~n19319;
  assign n19321 = ~n19218 & ~n19222;
  assign n19322 = ~n19320 & ~n19321;
  assign n19323 = ~n19320 & ~n19322;
  assign n19324 = ~n19321 & ~n19322;
  assign n19325 = ~n19323 & ~n19324;
  assign n19326 = n3622 & n8612;
  assign n19327 = pi111  & n3814;
  assign n19328 = pi113  & n3620;
  assign n19329 = pi112  & n3615;
  assign n19330 = ~n19328 & ~n19329;
  assign n19331 = ~n19327 & n19330;
  assign n19332 = ~n19326 & n19331;
  assign n19333 = pi32  & ~n19332;
  assign n19334 = pi32  & ~n19333;
  assign n19335 = ~n19332 & ~n19333;
  assign n19336 = ~n19334 & ~n19335;
  assign n19337 = ~n19198 & ~n19204;
  assign n19338 = n19336 & n19337;
  assign n19339 = ~n19336 & ~n19337;
  assign n19340 = ~n19338 & ~n19339;
  assign n19341 = ~n19006 & ~n19166;
  assign n19342 = ~n19163 & ~n19341;
  assign n19343 = n5739 & n5943;
  assign n19344 = pi102  & n6030;
  assign n19345 = pi104  & n5737;
  assign n19346 = pi103  & n5732;
  assign n19347 = ~n19345 & ~n19346;
  assign n19348 = ~n19344 & n19347;
  assign n19349 = ~n19343 & n19348;
  assign n19350 = pi41  & ~n19349;
  assign n19351 = pi41  & ~n19350;
  assign n19352 = ~n19349 & ~n19350;
  assign n19353 = ~n19351 & ~n19352;
  assign n19354 = ~n19146 & ~n19150;
  assign n19355 = n5169 & n6539;
  assign n19356 = pi99  & n6873;
  assign n19357 = pi101  & n6537;
  assign n19358 = pi100  & n6532;
  assign n19359 = ~n19357 & ~n19358;
  assign n19360 = ~n19356 & n19359;
  assign n19361 = ~n19355 & n19360;
  assign n19362 = pi44  & ~n19361;
  assign n19363 = pi44  & ~n19362;
  assign n19364 = ~n19361 & ~n19362;
  assign n19365 = ~n19363 & ~n19364;
  assign n19366 = ~n19009 & ~n19131;
  assign n19367 = ~n19128 & ~n19366;
  assign n19368 = ~n19033 & ~n19039;
  assign n19369 = pi79  & n13835;
  assign n19370 = pi80  & ~n13434;
  assign n19371 = ~n19369 & ~n19370;
  assign n19372 = ~n19014 & ~n19018;
  assign n19373 = ~n19371 & n19372;
  assign n19374 = n19371 & ~n19372;
  assign n19375 = ~n19373 & ~n19374;
  assign n19376 = pi81  & n13004;
  assign n19377 = pi83  & n12625;
  assign n19378 = pi82  & n12620;
  assign n19379 = ~n19377 & ~n19378;
  assign n19380 = ~n19376 & n19379;
  assign n19381 = ~n12627 & n19380;
  assign n19382 = ~n1696 & n19380;
  assign n19383 = ~n19381 & ~n19382;
  assign n19384 = pi62  & ~n19383;
  assign n19385 = ~pi62  & n19383;
  assign n19386 = ~n19384 & ~n19385;
  assign n19387 = n19375 & ~n19386;
  assign n19388 = ~n19375 & n19386;
  assign n19389 = ~n19387 & ~n19388;
  assign n19390 = ~n19368 & n19389;
  assign n19391 = n19368 & ~n19389;
  assign n19392 = ~n19390 & ~n19391;
  assign n19393 = n2133 & n11488;
  assign n19394 = pi84  & n11847;
  assign n19395 = pi86  & n11486;
  assign n19396 = pi85  & n11481;
  assign n19397 = ~n19395 & ~n19396;
  assign n19398 = ~n19394 & n19397;
  assign n19399 = ~n19393 & n19398;
  assign n19400 = pi59  & ~n19399;
  assign n19401 = pi59  & ~n19400;
  assign n19402 = ~n19399 & ~n19400;
  assign n19403 = ~n19401 & ~n19402;
  assign n19404 = n19392 & ~n19403;
  assign n19405 = n19392 & ~n19404;
  assign n19406 = ~n19403 & ~n19404;
  assign n19407 = ~n19405 & ~n19406;
  assign n19408 = ~n19052 & ~n19058;
  assign n19409 = n19407 & n19408;
  assign n19410 = ~n19407 & ~n19408;
  assign n19411 = ~n19409 & ~n19410;
  assign n19412 = n2473 & n10394;
  assign n19413 = pi87  & n10744;
  assign n19414 = pi89  & n10392;
  assign n19415 = pi88  & n10387;
  assign n19416 = ~n19414 & ~n19415;
  assign n19417 = ~n19413 & n19416;
  assign n19418 = ~n19412 & n19417;
  assign n19419 = pi56  & ~n19418;
  assign n19420 = pi56  & ~n19419;
  assign n19421 = ~n19418 & ~n19419;
  assign n19422 = ~n19420 & ~n19421;
  assign n19423 = n19411 & ~n19422;
  assign n19424 = n19411 & ~n19423;
  assign n19425 = ~n19422 & ~n19423;
  assign n19426 = ~n19424 & ~n19425;
  assign n19427 = ~n19076 & n19426;
  assign n19428 = n19076 & ~n19426;
  assign n19429 = ~n19427 & ~n19428;
  assign n19430 = n3177 & n9310;
  assign n19431 = pi90  & n9701;
  assign n19432 = pi92  & n9308;
  assign n19433 = pi91  & n9303;
  assign n19434 = ~n19432 & ~n19433;
  assign n19435 = ~n19431 & n19434;
  assign n19436 = ~n19430 & n19435;
  assign n19437 = pi53  & ~n19436;
  assign n19438 = pi53  & ~n19437;
  assign n19439 = ~n19436 & ~n19437;
  assign n19440 = ~n19438 & ~n19439;
  assign n19441 = n19429 & n19440;
  assign n19442 = ~n19429 & ~n19440;
  assign n19443 = ~n19441 & ~n19442;
  assign n19444 = ~n19090 & ~n19096;
  assign n19445 = n19443 & ~n19444;
  assign n19446 = ~n19443 & n19444;
  assign n19447 = ~n19445 & ~n19446;
  assign n19448 = n3784 & n8334;
  assign n19449 = pi93  & n8685;
  assign n19450 = pi95  & n8332;
  assign n19451 = pi94  & n8327;
  assign n19452 = ~n19450 & ~n19451;
  assign n19453 = ~n19449 & n19452;
  assign n19454 = ~n19448 & n19453;
  assign n19455 = pi50  & ~n19454;
  assign n19456 = pi50  & ~n19455;
  assign n19457 = ~n19454 & ~n19455;
  assign n19458 = ~n19456 & ~n19457;
  assign n19459 = n19447 & ~n19458;
  assign n19460 = n19447 & ~n19459;
  assign n19461 = ~n19458 & ~n19459;
  assign n19462 = ~n19460 & ~n19461;
  assign n19463 = ~n19109 & ~n19115;
  assign n19464 = n19462 & n19463;
  assign n19465 = ~n19462 & ~n19463;
  assign n19466 = ~n19464 & ~n19465;
  assign n19467 = n4454 & n7408;
  assign n19468 = pi96  & n7740;
  assign n19469 = pi98  & n7406;
  assign n19470 = pi97  & n7401;
  assign n19471 = ~n19469 & ~n19470;
  assign n19472 = ~n19468 & n19471;
  assign n19473 = ~n19467 & n19472;
  assign n19474 = pi47  & ~n19473;
  assign n19475 = pi47  & ~n19474;
  assign n19476 = ~n19473 & ~n19474;
  assign n19477 = ~n19475 & ~n19476;
  assign n19478 = ~n19466 & n19477;
  assign n19479 = n19466 & ~n19477;
  assign n19480 = ~n19478 & ~n19479;
  assign n19481 = ~n19367 & n19480;
  assign n19482 = ~n19367 & ~n19481;
  assign n19483 = n19480 & ~n19481;
  assign n19484 = ~n19482 & ~n19483;
  assign n19485 = ~n19365 & ~n19484;
  assign n19486 = n19365 & n19484;
  assign n19487 = ~n19485 & ~n19486;
  assign n19488 = ~n19354 & n19487;
  assign n19489 = ~n19354 & ~n19488;
  assign n19490 = n19487 & ~n19488;
  assign n19491 = ~n19489 & ~n19490;
  assign n19492 = ~n19353 & ~n19491;
  assign n19493 = n19353 & n19491;
  assign n19494 = ~n19492 & ~n19493;
  assign n19495 = ~n19342 & n19494;
  assign n19496 = n19342 & ~n19494;
  assign n19497 = ~n19495 & ~n19496;
  assign n19498 = n5008 & n6775;
  assign n19499 = pi105  & n5241;
  assign n19500 = pi107  & n5006;
  assign n19501 = pi106  & n5001;
  assign n19502 = ~n19500 & ~n19501;
  assign n19503 = ~n19499 & n19502;
  assign n19504 = ~n19498 & n19503;
  assign n19505 = pi38  & ~n19504;
  assign n19506 = pi38  & ~n19505;
  assign n19507 = ~n19504 & ~n19505;
  assign n19508 = ~n19506 & ~n19507;
  assign n19509 = n19497 & ~n19508;
  assign n19510 = n19497 & ~n19509;
  assign n19511 = ~n19508 & ~n19509;
  assign n19512 = ~n19510 & ~n19511;
  assign n19513 = ~n19181 & ~n19185;
  assign n19514 = n19512 & n19513;
  assign n19515 = ~n19512 & ~n19513;
  assign n19516 = ~n19514 & ~n19515;
  assign n19517 = n4271 & n7665;
  assign n19518 = pi108  & n4503;
  assign n19519 = pi110  & n4269;
  assign n19520 = pi109  & n4264;
  assign n19521 = ~n19519 & ~n19520;
  assign n19522 = ~n19518 & n19521;
  assign n19523 = ~n19517 & n19522;
  assign n19524 = pi35  & ~n19523;
  assign n19525 = pi35  & ~n19524;
  assign n19526 = ~n19523 & ~n19524;
  assign n19527 = ~n19525 & ~n19526;
  assign n19528 = n19516 & ~n19527;
  assign n19529 = n19516 & ~n19528;
  assign n19530 = ~n19527 & ~n19528;
  assign n19531 = ~n19529 & ~n19530;
  assign n19532 = n19340 & ~n19531;
  assign n19533 = ~n19340 & n19531;
  assign n19534 = ~n19532 & ~n19533;
  assign n19535 = ~n19325 & n19534;
  assign n19536 = ~n19325 & ~n19535;
  assign n19537 = n19534 & ~n19535;
  assign n19538 = ~n19536 & ~n19537;
  assign n19539 = n19309 & ~n19538;
  assign n19540 = ~n19309 & n19538;
  assign n19541 = ~n19539 & ~n19540;
  assign n19542 = n19294 & n19541;
  assign n19543 = n19294 & ~n19542;
  assign n19544 = n19541 & ~n19542;
  assign n19545 = ~n19543 & ~n19544;
  assign n19546 = n19279 & ~n19545;
  assign n19547 = ~n19279 & n19545;
  assign n19548 = ~n19546 & ~n19547;
  assign n19549 = n19263 & n19548;
  assign n19550 = n19263 & ~n19549;
  assign n19551 = n19548 & ~n19549;
  assign n19552 = ~n19550 & ~n19551;
  assign n19553 = ~n18941 & ~n19239;
  assign n19554 = n19552 & n19553;
  assign n19555 = ~n19552 & ~n19553;
  assign n19556 = ~n19554 & ~n19555;
  assign n19557 = ~n19245 & ~n19248;
  assign n19558 = n19556 & ~n19557;
  assign n19559 = ~n19556 & n19557;
  assign po79  = ~n19558 & ~n19559;
  assign n19561 = ~n19555 & ~n19558;
  assign n19562 = ~n19261 & ~n19549;
  assign n19563 = ~n19278 & ~n19546;
  assign n19564 = pi127  & n1366;
  assign n19565 = n1297 & n13770;
  assign n19566 = ~n19564 & ~n19565;
  assign n19567 = pi17  & ~n19566;
  assign n19568 = pi17  & ~n19567;
  assign n19569 = ~n19566 & ~n19567;
  assign n19570 = ~n19568 & ~n19569;
  assign n19571 = ~n19563 & ~n19570;
  assign n19572 = ~n19563 & ~n19571;
  assign n19573 = ~n19570 & ~n19571;
  assign n19574 = ~n19572 & ~n19573;
  assign n19575 = n1611 & n13344;
  assign n19576 = pi124  & n1745;
  assign n19577 = pi126  & n1609;
  assign n19578 = pi125  & n1604;
  assign n19579 = ~n19577 & ~n19578;
  assign n19580 = ~n19576 & n19579;
  assign n19581 = ~n19575 & n19580;
  assign n19582 = pi20  & ~n19581;
  assign n19583 = pi20  & ~n19582;
  assign n19584 = ~n19581 & ~n19582;
  assign n19585 = ~n19583 & ~n19584;
  assign n19586 = ~n19292 & ~n19542;
  assign n19587 = n19585 & n19586;
  assign n19588 = ~n19585 & ~n19586;
  assign n19589 = ~n19587 & ~n19588;
  assign n19590 = n2043 & n12158;
  assign n19591 = pi121  & n2180;
  assign n19592 = pi123  & n2041;
  assign n19593 = pi122  & n2036;
  assign n19594 = ~n19592 & ~n19593;
  assign n19595 = ~n19591 & n19594;
  assign n19596 = ~n19590 & n19595;
  assign n19597 = pi23  & ~n19596;
  assign n19598 = pi23  & ~n19597;
  assign n19599 = ~n19596 & ~n19597;
  assign n19600 = ~n19598 & ~n19599;
  assign n19601 = ~n19308 & ~n19539;
  assign n19602 = ~n19600 & ~n19601;
  assign n19603 = ~n19600 & ~n19602;
  assign n19604 = ~n19601 & ~n19602;
  assign n19605 = ~n19603 & ~n19604;
  assign n19606 = n2523 & n11028;
  assign n19607 = pi118  & n2667;
  assign n19608 = pi120  & n2521;
  assign n19609 = pi119  & n2516;
  assign n19610 = ~n19608 & ~n19609;
  assign n19611 = ~n19607 & n19610;
  assign n19612 = ~n19606 & n19611;
  assign n19613 = pi26  & ~n19612;
  assign n19614 = pi26  & ~n19613;
  assign n19615 = ~n19612 & ~n19613;
  assign n19616 = ~n19614 & ~n19615;
  assign n19617 = ~n19322 & ~n19535;
  assign n19618 = n19616 & n19617;
  assign n19619 = ~n19616 & ~n19617;
  assign n19620 = ~n19618 & ~n19619;
  assign n19621 = n3034 & n9958;
  assign n19622 = pi115  & n3225;
  assign n19623 = pi117  & n3032;
  assign n19624 = pi116  & n3027;
  assign n19625 = ~n19623 & ~n19624;
  assign n19626 = ~n19622 & n19625;
  assign n19627 = ~n19621 & n19626;
  assign n19628 = pi29  & ~n19627;
  assign n19629 = pi29  & ~n19628;
  assign n19630 = ~n19627 & ~n19628;
  assign n19631 = ~n19629 & ~n19630;
  assign n19632 = ~n19339 & ~n19532;
  assign n19633 = ~n19631 & ~n19632;
  assign n19634 = ~n19631 & ~n19633;
  assign n19635 = ~n19632 & ~n19633;
  assign n19636 = ~n19634 & ~n19635;
  assign n19637 = n3622 & n8936;
  assign n19638 = pi112  & n3814;
  assign n19639 = pi114  & n3620;
  assign n19640 = pi113  & n3615;
  assign n19641 = ~n19639 & ~n19640;
  assign n19642 = ~n19638 & n19641;
  assign n19643 = ~n19637 & n19642;
  assign n19644 = pi32  & ~n19643;
  assign n19645 = pi32  & ~n19644;
  assign n19646 = ~n19643 & ~n19644;
  assign n19647 = ~n19645 & ~n19646;
  assign n19648 = ~n19515 & ~n19528;
  assign n19649 = n19647 & n19648;
  assign n19650 = ~n19647 & ~n19648;
  assign n19651 = ~n19649 & ~n19650;
  assign n19652 = ~n19495 & ~n19509;
  assign n19653 = n5008 & n7060;
  assign n19654 = pi106  & n5241;
  assign n19655 = pi108  & n5006;
  assign n19656 = pi107  & n5001;
  assign n19657 = ~n19655 & ~n19656;
  assign n19658 = ~n19654 & n19657;
  assign n19659 = ~n19653 & n19658;
  assign n19660 = pi38  & ~n19659;
  assign n19661 = pi38  & ~n19660;
  assign n19662 = ~n19659 & ~n19660;
  assign n19663 = ~n19661 & ~n19662;
  assign n19664 = ~n19488 & ~n19492;
  assign n19665 = n5739 & n6207;
  assign n19666 = pi103  & n6030;
  assign n19667 = pi105  & n5737;
  assign n19668 = pi104  & n5732;
  assign n19669 = ~n19667 & ~n19668;
  assign n19670 = ~n19666 & n19669;
  assign n19671 = ~n19665 & n19670;
  assign n19672 = pi41  & ~n19671;
  assign n19673 = pi41  & ~n19672;
  assign n19674 = ~n19671 & ~n19672;
  assign n19675 = ~n19673 & ~n19674;
  assign n19676 = ~n19481 & ~n19485;
  assign n19677 = ~n19410 & ~n19423;
  assign n19678 = n2801 & n10394;
  assign n19679 = pi88  & n10744;
  assign n19680 = pi90  & n10392;
  assign n19681 = pi89  & n10387;
  assign n19682 = ~n19680 & ~n19681;
  assign n19683 = ~n19679 & n19682;
  assign n19684 = ~n19678 & n19683;
  assign n19685 = pi56  & ~n19684;
  assign n19686 = pi56  & ~n19685;
  assign n19687 = ~n19684 & ~n19685;
  assign n19688 = ~n19686 & ~n19687;
  assign n19689 = ~n19390 & ~n19404;
  assign n19690 = n1834 & n12627;
  assign n19691 = pi82  & n13004;
  assign n19692 = pi84  & n12625;
  assign n19693 = pi83  & n12620;
  assign n19694 = ~n19692 & ~n19693;
  assign n19695 = ~n19691 & n19694;
  assign n19696 = ~n19690 & n19695;
  assign n19697 = pi62  & ~n19696;
  assign n19698 = pi62  & ~n19697;
  assign n19699 = ~n19696 & ~n19697;
  assign n19700 = ~n19698 & ~n19699;
  assign n19701 = pi80  & n13835;
  assign n19702 = pi81  & ~n13434;
  assign n19703 = ~n19701 & ~n19702;
  assign n19704 = n19371 & ~n19703;
  assign n19705 = ~n19371 & n19703;
  assign n19706 = ~n19704 & ~n19705;
  assign n19707 = ~n19700 & n19706;
  assign n19708 = ~n19700 & ~n19707;
  assign n19709 = ~n19705 & ~n19707;
  assign n19710 = ~n19704 & n19709;
  assign n19711 = ~n19708 & ~n19710;
  assign n19712 = ~n19374 & ~n19387;
  assign n19713 = n19711 & n19712;
  assign n19714 = ~n19711 & ~n19712;
  assign n19715 = ~n19713 & ~n19714;
  assign n19716 = n2288 & n11488;
  assign n19717 = pi85  & n11847;
  assign n19718 = pi87  & n11486;
  assign n19719 = pi86  & n11481;
  assign n19720 = ~n19718 & ~n19719;
  assign n19721 = ~n19717 & n19720;
  assign n19722 = ~n19716 & n19721;
  assign n19723 = pi59  & ~n19722;
  assign n19724 = pi59  & ~n19723;
  assign n19725 = ~n19722 & ~n19723;
  assign n19726 = ~n19724 & ~n19725;
  assign n19727 = ~n19715 & n19726;
  assign n19728 = n19715 & ~n19726;
  assign n19729 = ~n19727 & ~n19728;
  assign n19730 = ~n19689 & n19729;
  assign n19731 = n19689 & ~n19729;
  assign n19732 = ~n19730 & ~n19731;
  assign n19733 = ~n19688 & n19732;
  assign n19734 = n19688 & ~n19732;
  assign n19735 = ~n19733 & ~n19734;
  assign n19736 = ~n19677 & n19735;
  assign n19737 = n19677 & ~n19735;
  assign n19738 = ~n19736 & ~n19737;
  assign n19739 = n3371 & n9310;
  assign n19740 = pi91  & n9701;
  assign n19741 = pi93  & n9308;
  assign n19742 = pi92  & n9303;
  assign n19743 = ~n19741 & ~n19742;
  assign n19744 = ~n19740 & n19743;
  assign n19745 = ~n19739 & n19744;
  assign n19746 = pi53  & ~n19745;
  assign n19747 = pi53  & ~n19746;
  assign n19748 = ~n19745 & ~n19746;
  assign n19749 = ~n19747 & ~n19748;
  assign n19750 = n19738 & ~n19749;
  assign n19751 = n19738 & ~n19750;
  assign n19752 = ~n19749 & ~n19750;
  assign n19753 = ~n19751 & ~n19752;
  assign n19754 = ~n19076 & ~n19426;
  assign n19755 = ~n19442 & ~n19754;
  assign n19756 = ~n19753 & ~n19755;
  assign n19757 = ~n19753 & ~n19756;
  assign n19758 = ~n19755 & ~n19756;
  assign n19759 = ~n19757 & ~n19758;
  assign n19760 = n4001 & n8334;
  assign n19761 = pi94  & n8685;
  assign n19762 = pi96  & n8332;
  assign n19763 = pi95  & n8327;
  assign n19764 = ~n19762 & ~n19763;
  assign n19765 = ~n19761 & n19764;
  assign n19766 = ~n19760 & n19765;
  assign n19767 = pi50  & ~n19766;
  assign n19768 = pi50  & ~n19767;
  assign n19769 = ~n19766 & ~n19767;
  assign n19770 = ~n19768 & ~n19769;
  assign n19771 = ~n19759 & n19770;
  assign n19772 = n19759 & ~n19770;
  assign n19773 = ~n19771 & ~n19772;
  assign n19774 = ~n19445 & ~n19459;
  assign n19775 = n19773 & n19774;
  assign n19776 = ~n19773 & ~n19774;
  assign n19777 = ~n19775 & ~n19776;
  assign n19778 = n4684 & n7408;
  assign n19779 = pi97  & n7740;
  assign n19780 = pi99  & n7406;
  assign n19781 = pi98  & n7401;
  assign n19782 = ~n19780 & ~n19781;
  assign n19783 = ~n19779 & n19782;
  assign n19784 = ~n19778 & n19783;
  assign n19785 = pi47  & ~n19784;
  assign n19786 = pi47  & ~n19785;
  assign n19787 = ~n19784 & ~n19785;
  assign n19788 = ~n19786 & ~n19787;
  assign n19789 = n19777 & ~n19788;
  assign n19790 = n19777 & ~n19789;
  assign n19791 = ~n19788 & ~n19789;
  assign n19792 = ~n19790 & ~n19791;
  assign n19793 = ~n19465 & ~n19479;
  assign n19794 = ~n19792 & ~n19793;
  assign n19795 = ~n19792 & ~n19794;
  assign n19796 = ~n19793 & ~n19794;
  assign n19797 = ~n19795 & ~n19796;
  assign n19798 = n5413 & n6539;
  assign n19799 = pi100  & n6873;
  assign n19800 = pi102  & n6537;
  assign n19801 = pi101  & n6532;
  assign n19802 = ~n19800 & ~n19801;
  assign n19803 = ~n19799 & n19802;
  assign n19804 = ~n19798 & n19803;
  assign n19805 = pi44  & ~n19804;
  assign n19806 = pi44  & ~n19805;
  assign n19807 = ~n19804 & ~n19805;
  assign n19808 = ~n19806 & ~n19807;
  assign n19809 = ~n19797 & n19808;
  assign n19810 = n19797 & ~n19808;
  assign n19811 = ~n19809 & ~n19810;
  assign n19812 = ~n19676 & ~n19811;
  assign n19813 = n19676 & n19811;
  assign n19814 = ~n19812 & ~n19813;
  assign n19815 = ~n19675 & n19814;
  assign n19816 = n19675 & ~n19814;
  assign n19817 = ~n19815 & ~n19816;
  assign n19818 = ~n19664 & n19817;
  assign n19819 = n19664 & ~n19817;
  assign n19820 = ~n19818 & ~n19819;
  assign n19821 = ~n19663 & n19820;
  assign n19822 = n19663 & ~n19820;
  assign n19823 = ~n19821 & ~n19822;
  assign n19824 = ~n19652 & n19823;
  assign n19825 = n19652 & ~n19823;
  assign n19826 = ~n19824 & ~n19825;
  assign n19827 = n4271 & n7970;
  assign n19828 = pi109  & n4503;
  assign n19829 = pi111  & n4269;
  assign n19830 = pi110  & n4264;
  assign n19831 = ~n19829 & ~n19830;
  assign n19832 = ~n19828 & n19831;
  assign n19833 = ~n19827 & n19832;
  assign n19834 = pi35  & ~n19833;
  assign n19835 = pi35  & ~n19834;
  assign n19836 = ~n19833 & ~n19834;
  assign n19837 = ~n19835 & ~n19836;
  assign n19838 = n19826 & ~n19837;
  assign n19839 = n19826 & ~n19838;
  assign n19840 = ~n19837 & ~n19838;
  assign n19841 = ~n19839 & ~n19840;
  assign n19842 = n19651 & ~n19841;
  assign n19843 = ~n19651 & n19841;
  assign n19844 = ~n19842 & ~n19843;
  assign n19845 = ~n19636 & n19844;
  assign n19846 = ~n19636 & ~n19845;
  assign n19847 = n19844 & ~n19845;
  assign n19848 = ~n19846 & ~n19847;
  assign n19849 = n19620 & ~n19848;
  assign n19850 = ~n19620 & n19848;
  assign n19851 = ~n19849 & ~n19850;
  assign n19852 = ~n19605 & n19851;
  assign n19853 = ~n19605 & ~n19852;
  assign n19854 = n19851 & ~n19852;
  assign n19855 = ~n19853 & ~n19854;
  assign n19856 = ~n19589 & n19855;
  assign n19857 = n19589 & ~n19855;
  assign n19858 = ~n19856 & ~n19857;
  assign n19859 = ~n19574 & n19858;
  assign n19860 = n19574 & ~n19858;
  assign n19861 = ~n19859 & ~n19860;
  assign n19862 = ~n19562 & n19861;
  assign n19863 = ~n19562 & ~n19862;
  assign n19864 = n19861 & ~n19862;
  assign n19865 = ~n19863 & ~n19864;
  assign n19866 = ~n19561 & ~n19865;
  assign n19867 = n19561 & n19865;
  assign po80  = ~n19866 & ~n19867;
  assign n19869 = ~n19862 & ~n19866;
  assign n19870 = ~n19571 & ~n19859;
  assign n19871 = ~n19588 & ~n19857;
  assign n19872 = n1611 & n13742;
  assign n19873 = pi125  & n1745;
  assign n19874 = pi127  & n1609;
  assign n19875 = pi126  & n1604;
  assign n19876 = ~n19874 & ~n19875;
  assign n19877 = ~n19873 & n19876;
  assign n19878 = ~n19872 & n19877;
  assign n19879 = pi20  & ~n19878;
  assign n19880 = pi20  & ~n19879;
  assign n19881 = ~n19878 & ~n19879;
  assign n19882 = ~n19880 & ~n19881;
  assign n19883 = ~n19871 & ~n19882;
  assign n19884 = ~n19871 & ~n19883;
  assign n19885 = ~n19882 & ~n19883;
  assign n19886 = ~n19884 & ~n19885;
  assign n19887 = n2043 & n12189;
  assign n19888 = pi122  & n2180;
  assign n19889 = pi124  & n2041;
  assign n19890 = pi123  & n2036;
  assign n19891 = ~n19889 & ~n19890;
  assign n19892 = ~n19888 & n19891;
  assign n19893 = ~n19887 & n19892;
  assign n19894 = pi23  & ~n19893;
  assign n19895 = pi23  & ~n19894;
  assign n19896 = ~n19893 & ~n19894;
  assign n19897 = ~n19895 & ~n19896;
  assign n19898 = ~n19602 & ~n19852;
  assign n19899 = n19897 & n19898;
  assign n19900 = ~n19897 & ~n19898;
  assign n19901 = ~n19899 & ~n19900;
  assign n19902 = n3034 & n9984;
  assign n19903 = pi116  & n3225;
  assign n19904 = pi118  & n3032;
  assign n19905 = pi117  & n3027;
  assign n19906 = ~n19904 & ~n19905;
  assign n19907 = ~n19903 & n19906;
  assign n19908 = ~n19902 & n19907;
  assign n19909 = pi29  & ~n19908;
  assign n19910 = pi29  & ~n19909;
  assign n19911 = ~n19908 & ~n19909;
  assign n19912 = ~n19910 & ~n19911;
  assign n19913 = ~n19633 & ~n19845;
  assign n19914 = n19912 & n19913;
  assign n19915 = ~n19912 & ~n19913;
  assign n19916 = ~n19914 & ~n19915;
  assign n19917 = ~n19812 & ~n19815;
  assign n19918 = ~n19797 & ~n19808;
  assign n19919 = ~n19794 & ~n19918;
  assign n19920 = ~n19776 & ~n19789;
  assign n19921 = ~n19714 & ~n19728;
  assign n19922 = n1972 & n12627;
  assign n19923 = pi83  & n13004;
  assign n19924 = pi85  & n12625;
  assign n19925 = pi84  & n12620;
  assign n19926 = ~n19924 & ~n19925;
  assign n19927 = ~n19923 & n19926;
  assign n19928 = ~n19922 & n19927;
  assign n19929 = pi62  & ~n19928;
  assign n19930 = pi62  & ~n19929;
  assign n19931 = ~n19928 & ~n19929;
  assign n19932 = ~n19930 & ~n19931;
  assign n19933 = pi81  & n13835;
  assign n19934 = pi82  & ~n13434;
  assign n19935 = ~n19933 & ~n19934;
  assign n19936 = ~pi17  & ~n19935;
  assign n19937 = pi17  & n19935;
  assign n19938 = ~n19936 & ~n19937;
  assign n19939 = ~n19703 & n19938;
  assign n19940 = n19703 & ~n19938;
  assign n19941 = ~n19939 & ~n19940;
  assign n19942 = ~n19932 & n19941;
  assign n19943 = ~n19932 & ~n19942;
  assign n19944 = n19941 & ~n19942;
  assign n19945 = ~n19943 & ~n19944;
  assign n19946 = ~n19709 & ~n19945;
  assign n19947 = ~n19709 & ~n19946;
  assign n19948 = ~n19945 & ~n19946;
  assign n19949 = ~n19947 & ~n19948;
  assign n19950 = n2446 & n11488;
  assign n19951 = pi86  & n11847;
  assign n19952 = pi88  & n11486;
  assign n19953 = pi87  & n11481;
  assign n19954 = ~n19952 & ~n19953;
  assign n19955 = ~n19951 & n19954;
  assign n19956 = ~n19950 & n19955;
  assign n19957 = pi59  & ~n19956;
  assign n19958 = pi59  & ~n19957;
  assign n19959 = ~n19956 & ~n19957;
  assign n19960 = ~n19958 & ~n19959;
  assign n19961 = n19949 & n19960;
  assign n19962 = ~n19949 & ~n19960;
  assign n19963 = ~n19961 & ~n19962;
  assign n19964 = ~n19921 & n19963;
  assign n19965 = n19921 & ~n19963;
  assign n19966 = ~n19964 & ~n19965;
  assign n19967 = n2978 & n10394;
  assign n19968 = pi89  & n10744;
  assign n19969 = pi91  & n10392;
  assign n19970 = pi90  & n10387;
  assign n19971 = ~n19969 & ~n19970;
  assign n19972 = ~n19968 & n19971;
  assign n19973 = ~n19967 & n19972;
  assign n19974 = pi56  & ~n19973;
  assign n19975 = pi56  & ~n19974;
  assign n19976 = ~n19973 & ~n19974;
  assign n19977 = ~n19975 & ~n19976;
  assign n19978 = n19966 & ~n19977;
  assign n19979 = n19966 & ~n19978;
  assign n19980 = ~n19977 & ~n19978;
  assign n19981 = ~n19979 & ~n19980;
  assign n19982 = ~n19730 & ~n19733;
  assign n19983 = n19981 & n19982;
  assign n19984 = ~n19981 & ~n19982;
  assign n19985 = ~n19983 & ~n19984;
  assign n19986 = n3565 & n9310;
  assign n19987 = pi92  & n9701;
  assign n19988 = pi94  & n9308;
  assign n19989 = pi93  & n9303;
  assign n19990 = ~n19988 & ~n19989;
  assign n19991 = ~n19987 & n19990;
  assign n19992 = ~n19986 & n19991;
  assign n19993 = pi53  & ~n19992;
  assign n19994 = pi53  & ~n19993;
  assign n19995 = ~n19992 & ~n19993;
  assign n19996 = ~n19994 & ~n19995;
  assign n19997 = n19985 & ~n19996;
  assign n19998 = n19985 & ~n19997;
  assign n19999 = ~n19996 & ~n19997;
  assign n20000 = ~n19998 & ~n19999;
  assign n20001 = ~n19736 & ~n19750;
  assign n20002 = n20000 & n20001;
  assign n20003 = ~n20000 & ~n20001;
  assign n20004 = ~n20002 & ~n20003;
  assign n20005 = n4211 & n8334;
  assign n20006 = pi95  & n8685;
  assign n20007 = pi97  & n8332;
  assign n20008 = pi96  & n8327;
  assign n20009 = ~n20007 & ~n20008;
  assign n20010 = ~n20006 & n20009;
  assign n20011 = ~n20005 & n20010;
  assign n20012 = pi50  & ~n20011;
  assign n20013 = pi50  & ~n20012;
  assign n20014 = ~n20011 & ~n20012;
  assign n20015 = ~n20013 & ~n20014;
  assign n20016 = ~n19759 & ~n19770;
  assign n20017 = ~n19756 & ~n20016;
  assign n20018 = ~n20015 & ~n20017;
  assign n20019 = n20015 & n20017;
  assign n20020 = ~n20018 & ~n20019;
  assign n20021 = ~n20004 & n20020;
  assign n20022 = n20004 & ~n20020;
  assign n20023 = ~n20021 & ~n20022;
  assign n20024 = n4910 & n7408;
  assign n20025 = pi98  & n7740;
  assign n20026 = pi100  & n7406;
  assign n20027 = pi99  & n7401;
  assign n20028 = ~n20026 & ~n20027;
  assign n20029 = ~n20025 & n20028;
  assign n20030 = ~n20024 & n20029;
  assign n20031 = pi47  & ~n20030;
  assign n20032 = pi47  & ~n20031;
  assign n20033 = ~n20030 & ~n20031;
  assign n20034 = ~n20032 & ~n20033;
  assign n20035 = ~n20023 & ~n20034;
  assign n20036 = n20023 & n20034;
  assign n20037 = ~n20035 & ~n20036;
  assign n20038 = n19920 & ~n20037;
  assign n20039 = ~n19920 & n20037;
  assign n20040 = ~n20038 & ~n20039;
  assign n20041 = n5664 & n6539;
  assign n20042 = pi101  & n6873;
  assign n20043 = pi103  & n6537;
  assign n20044 = pi102  & n6532;
  assign n20045 = ~n20043 & ~n20044;
  assign n20046 = ~n20042 & n20045;
  assign n20047 = ~n20041 & n20046;
  assign n20048 = pi44  & ~n20047;
  assign n20049 = pi44  & ~n20048;
  assign n20050 = ~n20047 & ~n20048;
  assign n20051 = ~n20049 & ~n20050;
  assign n20052 = n20040 & ~n20051;
  assign n20053 = n20040 & ~n20052;
  assign n20054 = ~n20051 & ~n20052;
  assign n20055 = ~n20053 & ~n20054;
  assign n20056 = ~n19919 & n20055;
  assign n20057 = n19919 & ~n20055;
  assign n20058 = ~n20056 & ~n20057;
  assign n20059 = n5739 & n6477;
  assign n20060 = pi104  & n6030;
  assign n20061 = pi106  & n5737;
  assign n20062 = pi105  & n5732;
  assign n20063 = ~n20061 & ~n20062;
  assign n20064 = ~n20060 & n20063;
  assign n20065 = ~n20059 & n20064;
  assign n20066 = pi41  & ~n20065;
  assign n20067 = pi41  & ~n20066;
  assign n20068 = ~n20065 & ~n20066;
  assign n20069 = ~n20067 & ~n20068;
  assign n20070 = ~n20058 & ~n20069;
  assign n20071 = n20058 & n20069;
  assign n20072 = ~n20070 & ~n20071;
  assign n20073 = n19917 & ~n20072;
  assign n20074 = ~n19917 & n20072;
  assign n20075 = ~n20073 & ~n20074;
  assign n20076 = n5008 & n7349;
  assign n20077 = pi107  & n5241;
  assign n20078 = pi109  & n5006;
  assign n20079 = pi108  & n5001;
  assign n20080 = ~n20078 & ~n20079;
  assign n20081 = ~n20077 & n20080;
  assign n20082 = ~n20076 & n20081;
  assign n20083 = pi38  & ~n20082;
  assign n20084 = pi38  & ~n20083;
  assign n20085 = ~n20082 & ~n20083;
  assign n20086 = ~n20084 & ~n20085;
  assign n20087 = n20075 & ~n20086;
  assign n20088 = n20075 & ~n20087;
  assign n20089 = ~n20086 & ~n20087;
  assign n20090 = ~n20088 & ~n20089;
  assign n20091 = ~n19818 & ~n19821;
  assign n20092 = n20090 & n20091;
  assign n20093 = ~n20090 & ~n20091;
  assign n20094 = ~n20092 & ~n20093;
  assign n20095 = n4271 & n7997;
  assign n20096 = pi110  & n4503;
  assign n20097 = pi112  & n4269;
  assign n20098 = pi111  & n4264;
  assign n20099 = ~n20097 & ~n20098;
  assign n20100 = ~n20096 & n20099;
  assign n20101 = ~n20095 & n20100;
  assign n20102 = pi35  & ~n20101;
  assign n20103 = pi35  & ~n20102;
  assign n20104 = ~n20101 & ~n20102;
  assign n20105 = ~n20103 & ~n20104;
  assign n20106 = n20094 & ~n20105;
  assign n20107 = n20094 & ~n20106;
  assign n20108 = ~n20105 & ~n20106;
  assign n20109 = ~n20107 & ~n20108;
  assign n20110 = ~n19824 & ~n19838;
  assign n20111 = n20109 & n20110;
  assign n20112 = ~n20109 & ~n20110;
  assign n20113 = ~n20111 & ~n20112;
  assign n20114 = n3622 & n8963;
  assign n20115 = pi113  & n3814;
  assign n20116 = pi115  & n3620;
  assign n20117 = pi114  & n3615;
  assign n20118 = ~n20116 & ~n20117;
  assign n20119 = ~n20115 & n20118;
  assign n20120 = ~n20114 & n20119;
  assign n20121 = pi32  & ~n20120;
  assign n20122 = pi32  & ~n20121;
  assign n20123 = ~n20120 & ~n20121;
  assign n20124 = ~n20122 & ~n20123;
  assign n20125 = ~n19650 & ~n19842;
  assign n20126 = ~n20124 & ~n20125;
  assign n20127 = n20124 & n20125;
  assign n20128 = ~n20126 & ~n20127;
  assign n20129 = n20113 & n20128;
  assign n20130 = n20113 & ~n20129;
  assign n20131 = n20128 & ~n20129;
  assign n20132 = ~n20130 & ~n20131;
  assign n20133 = n19916 & ~n20132;
  assign n20134 = n19916 & ~n20133;
  assign n20135 = ~n20132 & ~n20133;
  assign n20136 = ~n20134 & ~n20135;
  assign n20137 = n2523 & n11389;
  assign n20138 = pi119  & n2667;
  assign n20139 = pi121  & n2521;
  assign n20140 = pi120  & n2516;
  assign n20141 = ~n20139 & ~n20140;
  assign n20142 = ~n20138 & n20141;
  assign n20143 = ~n20137 & n20142;
  assign n20144 = pi26  & ~n20143;
  assign n20145 = pi26  & ~n20144;
  assign n20146 = ~n20143 & ~n20144;
  assign n20147 = ~n20145 & ~n20146;
  assign n20148 = ~n19619 & ~n19849;
  assign n20149 = ~n20147 & ~n20148;
  assign n20150 = n20147 & n20148;
  assign n20151 = ~n20149 & ~n20150;
  assign n20152 = ~n20136 & n20151;
  assign n20153 = ~n20136 & ~n20152;
  assign n20154 = n20151 & ~n20152;
  assign n20155 = ~n20153 & ~n20154;
  assign n20156 = n19901 & ~n20155;
  assign n20157 = n19901 & ~n20156;
  assign n20158 = ~n20155 & ~n20156;
  assign n20159 = ~n20157 & ~n20158;
  assign n20160 = ~n19886 & n20159;
  assign n20161 = n19886 & ~n20159;
  assign n20162 = ~n20160 & ~n20161;
  assign n20163 = ~n19870 & ~n20162;
  assign n20164 = ~n19870 & ~n20163;
  assign n20165 = ~n20162 & ~n20163;
  assign n20166 = ~n20164 & ~n20165;
  assign n20167 = ~n19869 & ~n20166;
  assign n20168 = n19869 & n20166;
  assign po81  = ~n20167 & ~n20168;
  assign n20170 = ~n20163 & ~n20167;
  assign n20171 = ~n19886 & ~n20159;
  assign n20172 = ~n19883 & ~n20171;
  assign n20173 = n2043 & n12943;
  assign n20174 = pi123  & n2180;
  assign n20175 = pi125  & n2041;
  assign n20176 = pi124  & n2036;
  assign n20177 = ~n20175 & ~n20176;
  assign n20178 = ~n20174 & n20177;
  assign n20179 = ~n20173 & n20178;
  assign n20180 = pi23  & ~n20179;
  assign n20181 = pi23  & ~n20180;
  assign n20182 = ~n20179 & ~n20180;
  assign n20183 = ~n20181 & ~n20182;
  assign n20184 = ~n20149 & ~n20152;
  assign n20185 = n20183 & n20184;
  assign n20186 = ~n20183 & ~n20184;
  assign n20187 = ~n20185 & ~n20186;
  assign n20188 = n2523 & n11778;
  assign n20189 = pi120  & n2667;
  assign n20190 = pi122  & n2521;
  assign n20191 = pi121  & n2516;
  assign n20192 = ~n20190 & ~n20191;
  assign n20193 = ~n20189 & n20192;
  assign n20194 = ~n20188 & n20193;
  assign n20195 = pi26  & ~n20194;
  assign n20196 = pi26  & ~n20195;
  assign n20197 = ~n20194 & ~n20195;
  assign n20198 = ~n20196 & ~n20197;
  assign n20199 = ~n19915 & ~n20133;
  assign n20200 = n20198 & n20199;
  assign n20201 = ~n20198 & ~n20199;
  assign n20202 = ~n20200 & ~n20201;
  assign n20203 = n3034 & n10667;
  assign n20204 = pi117  & n3225;
  assign n20205 = pi119  & n3032;
  assign n20206 = pi118  & n3027;
  assign n20207 = ~n20205 & ~n20206;
  assign n20208 = ~n20204 & n20207;
  assign n20209 = ~n20203 & n20208;
  assign n20210 = pi29  & ~n20209;
  assign n20211 = pi29  & ~n20210;
  assign n20212 = ~n20209 & ~n20210;
  assign n20213 = ~n20211 & ~n20212;
  assign n20214 = ~n20126 & ~n20129;
  assign n20215 = n20213 & n20214;
  assign n20216 = ~n20213 & ~n20214;
  assign n20217 = ~n20215 & ~n20216;
  assign n20218 = n3622 & n9614;
  assign n20219 = pi114  & n3814;
  assign n20220 = pi116  & n3620;
  assign n20221 = pi115  & n3615;
  assign n20222 = ~n20220 & ~n20221;
  assign n20223 = ~n20219 & n20222;
  assign n20224 = ~n20218 & n20223;
  assign n20225 = pi32  & ~n20224;
  assign n20226 = pi32  & ~n20225;
  assign n20227 = ~n20224 & ~n20225;
  assign n20228 = ~n20226 & ~n20227;
  assign n20229 = ~n20106 & ~n20112;
  assign n20230 = n20228 & n20229;
  assign n20231 = ~n20228 & ~n20229;
  assign n20232 = ~n20230 & ~n20231;
  assign n20233 = ~n19919 & ~n20055;
  assign n20234 = ~n20052 & ~n20233;
  assign n20235 = n5943 & n6539;
  assign n20236 = pi102  & n6873;
  assign n20237 = pi104  & n6537;
  assign n20238 = pi103  & n6532;
  assign n20239 = ~n20237 & ~n20238;
  assign n20240 = ~n20236 & n20239;
  assign n20241 = ~n20235 & n20240;
  assign n20242 = pi44  & ~n20241;
  assign n20243 = pi44  & ~n20242;
  assign n20244 = ~n20241 & ~n20242;
  assign n20245 = ~n20243 & ~n20244;
  assign n20246 = ~n20035 & ~n20039;
  assign n20247 = ~n19962 & ~n19964;
  assign n20248 = pi82  & n13835;
  assign n20249 = pi83  & ~n13434;
  assign n20250 = ~n20248 & ~n20249;
  assign n20251 = ~n19936 & ~n19939;
  assign n20252 = ~n20250 & n20251;
  assign n20253 = n20250 & ~n20251;
  assign n20254 = ~n20252 & ~n20253;
  assign n20255 = n2133 & n12627;
  assign n20256 = pi84  & n13004;
  assign n20257 = pi86  & n12625;
  assign n20258 = pi85  & n12620;
  assign n20259 = ~n20257 & ~n20258;
  assign n20260 = ~n20256 & n20259;
  assign n20261 = ~n20255 & n20260;
  assign n20262 = pi62  & ~n20261;
  assign n20263 = pi62  & ~n20262;
  assign n20264 = ~n20261 & ~n20262;
  assign n20265 = ~n20263 & ~n20264;
  assign n20266 = ~n20254 & n20265;
  assign n20267 = n20254 & ~n20265;
  assign n20268 = ~n20266 & ~n20267;
  assign n20269 = ~n19942 & ~n19946;
  assign n20270 = n20268 & ~n20269;
  assign n20271 = ~n20268 & n20269;
  assign n20272 = ~n20270 & ~n20271;
  assign n20273 = n2473 & n11488;
  assign n20274 = pi87  & n11847;
  assign n20275 = pi89  & n11486;
  assign n20276 = pi88  & n11481;
  assign n20277 = ~n20275 & ~n20276;
  assign n20278 = ~n20274 & n20277;
  assign n20279 = ~n20273 & n20278;
  assign n20280 = pi59  & ~n20279;
  assign n20281 = pi59  & ~n20280;
  assign n20282 = ~n20279 & ~n20280;
  assign n20283 = ~n20281 & ~n20282;
  assign n20284 = n20272 & ~n20283;
  assign n20285 = n20272 & ~n20284;
  assign n20286 = ~n20283 & ~n20284;
  assign n20287 = ~n20285 & ~n20286;
  assign n20288 = ~n20247 & n20287;
  assign n20289 = n20247 & ~n20287;
  assign n20290 = ~n20288 & ~n20289;
  assign n20291 = n3177 & n10394;
  assign n20292 = pi90  & n10744;
  assign n20293 = pi92  & n10392;
  assign n20294 = pi91  & n10387;
  assign n20295 = ~n20293 & ~n20294;
  assign n20296 = ~n20292 & n20295;
  assign n20297 = ~n20291 & n20296;
  assign n20298 = pi56  & ~n20297;
  assign n20299 = pi56  & ~n20298;
  assign n20300 = ~n20297 & ~n20298;
  assign n20301 = ~n20299 & ~n20300;
  assign n20302 = n20290 & n20301;
  assign n20303 = ~n20290 & ~n20301;
  assign n20304 = ~n20302 & ~n20303;
  assign n20305 = ~n19978 & ~n19984;
  assign n20306 = n20304 & ~n20305;
  assign n20307 = ~n20304 & n20305;
  assign n20308 = ~n20306 & ~n20307;
  assign n20309 = n3784 & n9310;
  assign n20310 = pi93  & n9701;
  assign n20311 = pi95  & n9308;
  assign n20312 = pi94  & n9303;
  assign n20313 = ~n20311 & ~n20312;
  assign n20314 = ~n20310 & n20313;
  assign n20315 = ~n20309 & n20314;
  assign n20316 = pi53  & ~n20315;
  assign n20317 = pi53  & ~n20316;
  assign n20318 = ~n20315 & ~n20316;
  assign n20319 = ~n20317 & ~n20318;
  assign n20320 = n20308 & ~n20319;
  assign n20321 = n20308 & ~n20320;
  assign n20322 = ~n20319 & ~n20320;
  assign n20323 = ~n20321 & ~n20322;
  assign n20324 = ~n19997 & ~n20003;
  assign n20325 = n20323 & n20324;
  assign n20326 = ~n20323 & ~n20324;
  assign n20327 = ~n20325 & ~n20326;
  assign n20328 = n4454 & n8334;
  assign n20329 = pi96  & n8685;
  assign n20330 = pi98  & n8332;
  assign n20331 = pi97  & n8327;
  assign n20332 = ~n20330 & ~n20331;
  assign n20333 = ~n20329 & n20332;
  assign n20334 = ~n20328 & n20333;
  assign n20335 = pi50  & ~n20334;
  assign n20336 = pi50  & ~n20335;
  assign n20337 = ~n20334 & ~n20335;
  assign n20338 = ~n20336 & ~n20337;
  assign n20339 = n20327 & ~n20338;
  assign n20340 = n20327 & ~n20339;
  assign n20341 = ~n20338 & ~n20339;
  assign n20342 = ~n20340 & ~n20341;
  assign n20343 = ~n20019 & ~n20021;
  assign n20344 = n20342 & ~n20343;
  assign n20345 = ~n20342 & n20343;
  assign n20346 = ~n20344 & ~n20345;
  assign n20347 = n5169 & n7408;
  assign n20348 = pi99  & n7740;
  assign n20349 = pi101  & n7406;
  assign n20350 = pi100  & n7401;
  assign n20351 = ~n20349 & ~n20350;
  assign n20352 = ~n20348 & n20351;
  assign n20353 = ~n20347 & n20352;
  assign n20354 = pi47  & ~n20353;
  assign n20355 = pi47  & ~n20354;
  assign n20356 = ~n20353 & ~n20354;
  assign n20357 = ~n20355 & ~n20356;
  assign n20358 = ~n20346 & n20357;
  assign n20359 = n20346 & ~n20357;
  assign n20360 = ~n20358 & ~n20359;
  assign n20361 = ~n20246 & n20360;
  assign n20362 = ~n20246 & ~n20361;
  assign n20363 = n20360 & ~n20361;
  assign n20364 = ~n20362 & ~n20363;
  assign n20365 = ~n20245 & ~n20364;
  assign n20366 = n20245 & n20364;
  assign n20367 = ~n20365 & ~n20366;
  assign n20368 = ~n20234 & n20367;
  assign n20369 = n20234 & ~n20367;
  assign n20370 = ~n20368 & ~n20369;
  assign n20371 = n5739 & n6775;
  assign n20372 = pi105  & n6030;
  assign n20373 = pi107  & n5737;
  assign n20374 = pi106  & n5732;
  assign n20375 = ~n20373 & ~n20374;
  assign n20376 = ~n20372 & n20375;
  assign n20377 = ~n20371 & n20376;
  assign n20378 = pi41  & ~n20377;
  assign n20379 = pi41  & ~n20378;
  assign n20380 = ~n20377 & ~n20378;
  assign n20381 = ~n20379 & ~n20380;
  assign n20382 = n20370 & ~n20381;
  assign n20383 = n20370 & ~n20382;
  assign n20384 = ~n20381 & ~n20382;
  assign n20385 = ~n20383 & ~n20384;
  assign n20386 = ~n20070 & ~n20074;
  assign n20387 = n20385 & n20386;
  assign n20388 = ~n20385 & ~n20386;
  assign n20389 = ~n20387 & ~n20388;
  assign n20390 = n5008 & n7665;
  assign n20391 = pi108  & n5241;
  assign n20392 = pi110  & n5006;
  assign n20393 = pi109  & n5001;
  assign n20394 = ~n20392 & ~n20393;
  assign n20395 = ~n20391 & n20394;
  assign n20396 = ~n20390 & n20395;
  assign n20397 = pi38  & ~n20396;
  assign n20398 = pi38  & ~n20397;
  assign n20399 = ~n20396 & ~n20397;
  assign n20400 = ~n20398 & ~n20399;
  assign n20401 = n20389 & ~n20400;
  assign n20402 = n20389 & ~n20401;
  assign n20403 = ~n20400 & ~n20401;
  assign n20404 = ~n20402 & ~n20403;
  assign n20405 = ~n20087 & ~n20093;
  assign n20406 = n20404 & n20405;
  assign n20407 = ~n20404 & ~n20405;
  assign n20408 = ~n20406 & ~n20407;
  assign n20409 = n4271 & n8612;
  assign n20410 = pi111  & n4503;
  assign n20411 = pi113  & n4269;
  assign n20412 = pi112  & n4264;
  assign n20413 = ~n20411 & ~n20412;
  assign n20414 = ~n20410 & n20413;
  assign n20415 = ~n20409 & n20414;
  assign n20416 = pi35  & ~n20415;
  assign n20417 = pi35  & ~n20416;
  assign n20418 = ~n20415 & ~n20416;
  assign n20419 = ~n20417 & ~n20418;
  assign n20420 = n20408 & ~n20419;
  assign n20421 = n20408 & ~n20420;
  assign n20422 = ~n20419 & ~n20420;
  assign n20423 = ~n20421 & ~n20422;
  assign n20424 = n20232 & ~n20423;
  assign n20425 = ~n20232 & n20423;
  assign n20426 = ~n20424 & ~n20425;
  assign n20427 = n20217 & n20426;
  assign n20428 = n20217 & ~n20427;
  assign n20429 = n20426 & ~n20427;
  assign n20430 = ~n20428 & ~n20429;
  assign n20431 = n20202 & ~n20430;
  assign n20432 = ~n20202 & n20430;
  assign n20433 = ~n20431 & ~n20432;
  assign n20434 = n20187 & n20433;
  assign n20435 = n20187 & ~n20434;
  assign n20436 = n20433 & ~n20434;
  assign n20437 = ~n20435 & ~n20436;
  assign n20438 = ~n19900 & ~n20156;
  assign n20439 = pi126  & n1745;
  assign n20440 = pi127  & n1604;
  assign n20441 = ~n20439 & ~n20440;
  assign n20442 = ~n1611 & n20441;
  assign n20443 = n13773 & n20441;
  assign n20444 = ~n20442 & ~n20443;
  assign n20445 = pi20  & ~n20444;
  assign n20446 = ~pi20  & n20444;
  assign n20447 = ~n20445 & ~n20446;
  assign n20448 = ~n20438 & ~n20447;
  assign n20449 = ~n20438 & ~n20448;
  assign n20450 = ~n20447 & ~n20448;
  assign n20451 = ~n20449 & ~n20450;
  assign n20452 = ~n20437 & ~n20451;
  assign n20453 = n20437 & n20451;
  assign n20454 = ~n20452 & ~n20453;
  assign n20455 = ~n20172 & n20454;
  assign n20456 = ~n20172 & ~n20455;
  assign n20457 = n20454 & ~n20455;
  assign n20458 = ~n20456 & ~n20457;
  assign n20459 = ~n20170 & ~n20458;
  assign n20460 = n20170 & n20458;
  assign po82  = ~n20459 & ~n20460;
  assign n20462 = ~n20455 & ~n20459;
  assign n20463 = ~n20448 & ~n20452;
  assign n20464 = ~n20186 & ~n20434;
  assign n20465 = pi127  & n1745;
  assign n20466 = n1611 & n13770;
  assign n20467 = ~n20465 & ~n20466;
  assign n20468 = pi20  & ~n20467;
  assign n20469 = pi20  & ~n20468;
  assign n20470 = ~n20467 & ~n20468;
  assign n20471 = ~n20469 & ~n20470;
  assign n20472 = ~n20464 & ~n20471;
  assign n20473 = ~n20464 & ~n20472;
  assign n20474 = ~n20471 & ~n20472;
  assign n20475 = ~n20473 & ~n20474;
  assign n20476 = n2043 & n13344;
  assign n20477 = pi124  & n2180;
  assign n20478 = pi126  & n2041;
  assign n20479 = pi125  & n2036;
  assign n20480 = ~n20478 & ~n20479;
  assign n20481 = ~n20477 & n20480;
  assign n20482 = ~n20476 & n20481;
  assign n20483 = pi23  & ~n20482;
  assign n20484 = pi23  & ~n20483;
  assign n20485 = ~n20482 & ~n20483;
  assign n20486 = ~n20484 & ~n20485;
  assign n20487 = ~n20201 & ~n20431;
  assign n20488 = ~n20486 & ~n20487;
  assign n20489 = ~n20486 & ~n20488;
  assign n20490 = ~n20487 & ~n20488;
  assign n20491 = ~n20489 & ~n20490;
  assign n20492 = n2523 & n12158;
  assign n20493 = pi121  & n2667;
  assign n20494 = pi123  & n2521;
  assign n20495 = pi122  & n2516;
  assign n20496 = ~n20494 & ~n20495;
  assign n20497 = ~n20493 & n20496;
  assign n20498 = ~n20492 & n20497;
  assign n20499 = pi26  & ~n20498;
  assign n20500 = pi26  & ~n20499;
  assign n20501 = ~n20498 & ~n20499;
  assign n20502 = ~n20500 & ~n20501;
  assign n20503 = ~n20216 & ~n20427;
  assign n20504 = n20502 & n20503;
  assign n20505 = ~n20502 & ~n20503;
  assign n20506 = ~n20504 & ~n20505;
  assign n20507 = n3034 & n11028;
  assign n20508 = pi118  & n3225;
  assign n20509 = pi120  & n3032;
  assign n20510 = pi119  & n3027;
  assign n20511 = ~n20509 & ~n20510;
  assign n20512 = ~n20508 & n20511;
  assign n20513 = ~n20507 & n20512;
  assign n20514 = pi29  & ~n20513;
  assign n20515 = pi29  & ~n20514;
  assign n20516 = ~n20513 & ~n20514;
  assign n20517 = ~n20515 & ~n20516;
  assign n20518 = ~n20231 & ~n20424;
  assign n20519 = ~n20517 & ~n20518;
  assign n20520 = ~n20517 & ~n20519;
  assign n20521 = ~n20518 & ~n20519;
  assign n20522 = ~n20520 & ~n20521;
  assign n20523 = n3622 & n9958;
  assign n20524 = pi115  & n3814;
  assign n20525 = pi117  & n3620;
  assign n20526 = pi116  & n3615;
  assign n20527 = ~n20525 & ~n20526;
  assign n20528 = ~n20524 & n20527;
  assign n20529 = ~n20523 & n20528;
  assign n20530 = pi32  & ~n20529;
  assign n20531 = pi32  & ~n20530;
  assign n20532 = ~n20529 & ~n20530;
  assign n20533 = ~n20531 & ~n20532;
  assign n20534 = ~n20407 & ~n20420;
  assign n20535 = n20533 & n20534;
  assign n20536 = ~n20533 & ~n20534;
  assign n20537 = ~n20535 & ~n20536;
  assign n20538 = ~n20368 & ~n20382;
  assign n20539 = n5739 & n7060;
  assign n20540 = pi106  & n6030;
  assign n20541 = pi108  & n5737;
  assign n20542 = pi107  & n5732;
  assign n20543 = ~n20541 & ~n20542;
  assign n20544 = ~n20540 & n20543;
  assign n20545 = ~n20539 & n20544;
  assign n20546 = pi41  & ~n20545;
  assign n20547 = pi41  & ~n20546;
  assign n20548 = ~n20545 & ~n20546;
  assign n20549 = ~n20547 & ~n20548;
  assign n20550 = ~n20361 & ~n20365;
  assign n20551 = n6207 & n6539;
  assign n20552 = pi103  & n6873;
  assign n20553 = pi105  & n6537;
  assign n20554 = pi104  & n6532;
  assign n20555 = ~n20553 & ~n20554;
  assign n20556 = ~n20552 & n20555;
  assign n20557 = ~n20551 & n20556;
  assign n20558 = pi44  & ~n20557;
  assign n20559 = pi44  & ~n20558;
  assign n20560 = ~n20557 & ~n20558;
  assign n20561 = ~n20559 & ~n20560;
  assign n20562 = ~n20345 & ~n20359;
  assign n20563 = n5413 & n7408;
  assign n20564 = pi100  & n7740;
  assign n20565 = pi102  & n7406;
  assign n20566 = pi101  & n7401;
  assign n20567 = ~n20565 & ~n20566;
  assign n20568 = ~n20564 & n20567;
  assign n20569 = ~n20563 & n20568;
  assign n20570 = pi47  & ~n20569;
  assign n20571 = pi47  & ~n20570;
  assign n20572 = ~n20569 & ~n20570;
  assign n20573 = ~n20571 & ~n20572;
  assign n20574 = ~n20326 & ~n20339;
  assign n20575 = n4684 & n8334;
  assign n20576 = pi97  & n8685;
  assign n20577 = pi99  & n8332;
  assign n20578 = pi98  & n8327;
  assign n20579 = ~n20577 & ~n20578;
  assign n20580 = ~n20576 & n20579;
  assign n20581 = ~n20575 & n20580;
  assign n20582 = pi50  & ~n20581;
  assign n20583 = pi50  & ~n20582;
  assign n20584 = ~n20581 & ~n20582;
  assign n20585 = ~n20583 & ~n20584;
  assign n20586 = ~n20306 & ~n20320;
  assign n20587 = ~n20270 & ~n20284;
  assign n20588 = n2801 & n11488;
  assign n20589 = pi88  & n11847;
  assign n20590 = pi90  & n11486;
  assign n20591 = pi89  & n11481;
  assign n20592 = ~n20590 & ~n20591;
  assign n20593 = ~n20589 & n20592;
  assign n20594 = ~n20588 & n20593;
  assign n20595 = pi59  & ~n20594;
  assign n20596 = pi59  & ~n20595;
  assign n20597 = ~n20594 & ~n20595;
  assign n20598 = ~n20596 & ~n20597;
  assign n20599 = ~n20253 & ~n20267;
  assign n20600 = pi83  & n13835;
  assign n20601 = pi84  & ~n13434;
  assign n20602 = ~n20600 & ~n20601;
  assign n20603 = ~n20250 & n20602;
  assign n20604 = n20250 & ~n20602;
  assign n20605 = ~n20603 & ~n20604;
  assign n20606 = pi85  & n13004;
  assign n20607 = pi87  & n12625;
  assign n20608 = pi86  & n12620;
  assign n20609 = ~n20607 & ~n20608;
  assign n20610 = ~n20606 & n20609;
  assign n20611 = ~n12627 & n20610;
  assign n20612 = ~n2288 & n20610;
  assign n20613 = ~n20611 & ~n20612;
  assign n20614 = pi62  & ~n20613;
  assign n20615 = ~pi62  & n20613;
  assign n20616 = ~n20614 & ~n20615;
  assign n20617 = n20605 & ~n20616;
  assign n20618 = ~n20605 & n20616;
  assign n20619 = ~n20617 & ~n20618;
  assign n20620 = ~n20599 & n20619;
  assign n20621 = n20599 & ~n20619;
  assign n20622 = ~n20620 & ~n20621;
  assign n20623 = ~n20598 & n20622;
  assign n20624 = n20598 & ~n20622;
  assign n20625 = ~n20623 & ~n20624;
  assign n20626 = ~n20587 & n20625;
  assign n20627 = n20587 & ~n20625;
  assign n20628 = ~n20626 & ~n20627;
  assign n20629 = n3371 & n10394;
  assign n20630 = pi91  & n10744;
  assign n20631 = pi93  & n10392;
  assign n20632 = pi92  & n10387;
  assign n20633 = ~n20631 & ~n20632;
  assign n20634 = ~n20630 & n20633;
  assign n20635 = ~n20629 & n20634;
  assign n20636 = pi56  & ~n20635;
  assign n20637 = pi56  & ~n20636;
  assign n20638 = ~n20635 & ~n20636;
  assign n20639 = ~n20637 & ~n20638;
  assign n20640 = n20628 & ~n20639;
  assign n20641 = n20628 & ~n20640;
  assign n20642 = ~n20639 & ~n20640;
  assign n20643 = ~n20641 & ~n20642;
  assign n20644 = ~n20247 & ~n20287;
  assign n20645 = ~n20303 & ~n20644;
  assign n20646 = ~n20643 & ~n20645;
  assign n20647 = ~n20643 & ~n20646;
  assign n20648 = ~n20645 & ~n20646;
  assign n20649 = ~n20647 & ~n20648;
  assign n20650 = n4001 & n9310;
  assign n20651 = pi94  & n9701;
  assign n20652 = pi96  & n9308;
  assign n20653 = pi95  & n9303;
  assign n20654 = ~n20652 & ~n20653;
  assign n20655 = ~n20651 & n20654;
  assign n20656 = ~n20650 & n20655;
  assign n20657 = pi53  & ~n20656;
  assign n20658 = pi53  & ~n20657;
  assign n20659 = ~n20656 & ~n20657;
  assign n20660 = ~n20658 & ~n20659;
  assign n20661 = ~n20649 & n20660;
  assign n20662 = n20649 & ~n20660;
  assign n20663 = ~n20661 & ~n20662;
  assign n20664 = ~n20586 & ~n20663;
  assign n20665 = n20586 & n20663;
  assign n20666 = ~n20664 & ~n20665;
  assign n20667 = ~n20585 & n20666;
  assign n20668 = n20585 & ~n20666;
  assign n20669 = ~n20667 & ~n20668;
  assign n20670 = ~n20574 & n20669;
  assign n20671 = n20574 & ~n20669;
  assign n20672 = ~n20670 & ~n20671;
  assign n20673 = ~n20573 & n20672;
  assign n20674 = n20573 & ~n20672;
  assign n20675 = ~n20673 & ~n20674;
  assign n20676 = ~n20562 & n20675;
  assign n20677 = n20562 & ~n20675;
  assign n20678 = ~n20676 & ~n20677;
  assign n20679 = ~n20561 & n20678;
  assign n20680 = n20561 & ~n20678;
  assign n20681 = ~n20679 & ~n20680;
  assign n20682 = ~n20550 & n20681;
  assign n20683 = n20550 & ~n20681;
  assign n20684 = ~n20682 & ~n20683;
  assign n20685 = ~n20549 & n20684;
  assign n20686 = n20549 & ~n20684;
  assign n20687 = ~n20685 & ~n20686;
  assign n20688 = ~n20538 & n20687;
  assign n20689 = n20538 & ~n20687;
  assign n20690 = ~n20688 & ~n20689;
  assign n20691 = n5008 & n7970;
  assign n20692 = pi109  & n5241;
  assign n20693 = pi111  & n5006;
  assign n20694 = pi110  & n5001;
  assign n20695 = ~n20693 & ~n20694;
  assign n20696 = ~n20692 & n20695;
  assign n20697 = ~n20691 & n20696;
  assign n20698 = pi38  & ~n20697;
  assign n20699 = pi38  & ~n20698;
  assign n20700 = ~n20697 & ~n20698;
  assign n20701 = ~n20699 & ~n20700;
  assign n20702 = n20690 & ~n20701;
  assign n20703 = n20690 & ~n20702;
  assign n20704 = ~n20701 & ~n20702;
  assign n20705 = ~n20703 & ~n20704;
  assign n20706 = ~n20388 & ~n20401;
  assign n20707 = n20705 & n20706;
  assign n20708 = ~n20705 & ~n20706;
  assign n20709 = ~n20707 & ~n20708;
  assign n20710 = n4271 & n8936;
  assign n20711 = pi112  & n4503;
  assign n20712 = pi114  & n4269;
  assign n20713 = pi113  & n4264;
  assign n20714 = ~n20712 & ~n20713;
  assign n20715 = ~n20711 & n20714;
  assign n20716 = ~n20710 & n20715;
  assign n20717 = pi35  & ~n20716;
  assign n20718 = pi35  & ~n20717;
  assign n20719 = ~n20716 & ~n20717;
  assign n20720 = ~n20718 & ~n20719;
  assign n20721 = n20709 & ~n20720;
  assign n20722 = ~n20709 & n20720;
  assign n20723 = ~n20721 & ~n20722;
  assign n20724 = n20537 & n20723;
  assign n20725 = n20537 & ~n20724;
  assign n20726 = n20723 & ~n20724;
  assign n20727 = ~n20725 & ~n20726;
  assign n20728 = ~n20522 & n20727;
  assign n20729 = n20522 & ~n20727;
  assign n20730 = ~n20728 & ~n20729;
  assign n20731 = n20506 & ~n20730;
  assign n20732 = n20506 & ~n20731;
  assign n20733 = ~n20730 & ~n20731;
  assign n20734 = ~n20732 & ~n20733;
  assign n20735 = ~n20491 & n20734;
  assign n20736 = n20491 & ~n20734;
  assign n20737 = ~n20735 & ~n20736;
  assign n20738 = ~n20475 & ~n20737;
  assign n20739 = n20475 & n20737;
  assign n20740 = ~n20738 & ~n20739;
  assign n20741 = ~n20463 & n20740;
  assign n20742 = n20463 & ~n20740;
  assign n20743 = ~n20741 & ~n20742;
  assign n20744 = ~n20462 & n20743;
  assign n20745 = n20462 & ~n20743;
  assign po83  = ~n20744 & ~n20745;
  assign n20747 = ~n20491 & ~n20734;
  assign n20748 = ~n20488 & ~n20747;
  assign n20749 = n2043 & n13742;
  assign n20750 = pi125  & n2180;
  assign n20751 = pi127  & n2041;
  assign n20752 = pi126  & n2036;
  assign n20753 = ~n20751 & ~n20752;
  assign n20754 = ~n20750 & n20753;
  assign n20755 = ~n20749 & n20754;
  assign n20756 = pi23  & ~n20755;
  assign n20757 = pi23  & ~n20756;
  assign n20758 = ~n20755 & ~n20756;
  assign n20759 = ~n20757 & ~n20758;
  assign n20760 = ~n20748 & ~n20759;
  assign n20761 = ~n20748 & ~n20760;
  assign n20762 = ~n20759 & ~n20760;
  assign n20763 = ~n20761 & ~n20762;
  assign n20764 = n2523 & n12189;
  assign n20765 = pi122  & n2667;
  assign n20766 = pi124  & n2521;
  assign n20767 = pi123  & n2516;
  assign n20768 = ~n20766 & ~n20767;
  assign n20769 = ~n20765 & n20768;
  assign n20770 = ~n20764 & n20769;
  assign n20771 = pi26  & ~n20770;
  assign n20772 = pi26  & ~n20771;
  assign n20773 = ~n20770 & ~n20771;
  assign n20774 = ~n20772 & ~n20773;
  assign n20775 = ~n20505 & ~n20731;
  assign n20776 = n20774 & n20775;
  assign n20777 = ~n20774 & ~n20775;
  assign n20778 = ~n20776 & ~n20777;
  assign n20779 = ~n20522 & ~n20727;
  assign n20780 = ~n20519 & ~n20779;
  assign n20781 = n3034 & n11389;
  assign n20782 = pi119  & n3225;
  assign n20783 = pi121  & n3032;
  assign n20784 = pi120  & n3027;
  assign n20785 = ~n20783 & ~n20784;
  assign n20786 = ~n20782 & n20785;
  assign n20787 = ~n20781 & n20786;
  assign n20788 = pi29  & ~n20787;
  assign n20789 = pi29  & ~n20788;
  assign n20790 = ~n20787 & ~n20788;
  assign n20791 = ~n20789 & ~n20790;
  assign n20792 = ~n20780 & n20791;
  assign n20793 = n20780 & ~n20791;
  assign n20794 = ~n20792 & ~n20793;
  assign n20795 = n3622 & n9984;
  assign n20796 = pi116  & n3814;
  assign n20797 = pi118  & n3620;
  assign n20798 = pi117  & n3615;
  assign n20799 = ~n20797 & ~n20798;
  assign n20800 = ~n20796 & n20799;
  assign n20801 = ~n20795 & n20800;
  assign n20802 = pi32  & ~n20801;
  assign n20803 = pi32  & ~n20802;
  assign n20804 = ~n20801 & ~n20802;
  assign n20805 = ~n20803 & ~n20804;
  assign n20806 = ~n20536 & ~n20724;
  assign n20807 = n20805 & n20806;
  assign n20808 = ~n20805 & ~n20806;
  assign n20809 = ~n20807 & ~n20808;
  assign n20810 = ~n20708 & ~n20721;
  assign n20811 = ~n20664 & ~n20667;
  assign n20812 = pi84  & n13835;
  assign n20813 = pi85  & ~n13434;
  assign n20814 = ~n20812 & ~n20813;
  assign n20815 = ~pi20  & ~n20814;
  assign n20816 = pi20  & n20814;
  assign n20817 = ~n20815 & ~n20816;
  assign n20818 = ~n20602 & n20817;
  assign n20819 = n20602 & ~n20817;
  assign n20820 = ~n20818 & ~n20819;
  assign n20821 = n2446 & n12627;
  assign n20822 = pi86  & n13004;
  assign n20823 = pi88  & n12625;
  assign n20824 = pi87  & n12620;
  assign n20825 = ~n20823 & ~n20824;
  assign n20826 = ~n20822 & n20825;
  assign n20827 = ~n20821 & n20826;
  assign n20828 = pi62  & ~n20827;
  assign n20829 = pi62  & ~n20828;
  assign n20830 = ~n20827 & ~n20828;
  assign n20831 = ~n20829 & ~n20830;
  assign n20832 = n20820 & ~n20831;
  assign n20833 = n20820 & ~n20832;
  assign n20834 = ~n20831 & ~n20832;
  assign n20835 = ~n20833 & ~n20834;
  assign n20836 = ~n20603 & ~n20617;
  assign n20837 = ~n20835 & ~n20836;
  assign n20838 = ~n20835 & ~n20837;
  assign n20839 = ~n20836 & ~n20837;
  assign n20840 = ~n20838 & ~n20839;
  assign n20841 = n2978 & n11488;
  assign n20842 = pi89  & n11847;
  assign n20843 = pi91  & n11486;
  assign n20844 = pi90  & n11481;
  assign n20845 = ~n20843 & ~n20844;
  assign n20846 = ~n20842 & n20845;
  assign n20847 = ~n20841 & n20846;
  assign n20848 = pi59  & ~n20847;
  assign n20849 = pi59  & ~n20848;
  assign n20850 = ~n20847 & ~n20848;
  assign n20851 = ~n20849 & ~n20850;
  assign n20852 = ~n20840 & ~n20851;
  assign n20853 = ~n20840 & ~n20852;
  assign n20854 = ~n20851 & ~n20852;
  assign n20855 = ~n20853 & ~n20854;
  assign n20856 = ~n20620 & ~n20623;
  assign n20857 = n20855 & n20856;
  assign n20858 = ~n20855 & ~n20856;
  assign n20859 = ~n20857 & ~n20858;
  assign n20860 = n3565 & n10394;
  assign n20861 = pi92  & n10744;
  assign n20862 = pi94  & n10392;
  assign n20863 = pi93  & n10387;
  assign n20864 = ~n20862 & ~n20863;
  assign n20865 = ~n20861 & n20864;
  assign n20866 = ~n20860 & n20865;
  assign n20867 = pi56  & ~n20866;
  assign n20868 = pi56  & ~n20867;
  assign n20869 = ~n20866 & ~n20867;
  assign n20870 = ~n20868 & ~n20869;
  assign n20871 = n20859 & ~n20870;
  assign n20872 = n20859 & ~n20871;
  assign n20873 = ~n20870 & ~n20871;
  assign n20874 = ~n20872 & ~n20873;
  assign n20875 = ~n20626 & ~n20640;
  assign n20876 = n20874 & n20875;
  assign n20877 = ~n20874 & ~n20875;
  assign n20878 = ~n20876 & ~n20877;
  assign n20879 = n4211 & n9310;
  assign n20880 = pi95  & n9701;
  assign n20881 = pi97  & n9308;
  assign n20882 = pi96  & n9303;
  assign n20883 = ~n20881 & ~n20882;
  assign n20884 = ~n20880 & n20883;
  assign n20885 = ~n20879 & n20884;
  assign n20886 = pi53  & ~n20885;
  assign n20887 = pi53  & ~n20886;
  assign n20888 = ~n20885 & ~n20886;
  assign n20889 = ~n20887 & ~n20888;
  assign n20890 = ~n20649 & ~n20660;
  assign n20891 = ~n20646 & ~n20890;
  assign n20892 = ~n20889 & ~n20891;
  assign n20893 = n20889 & n20891;
  assign n20894 = ~n20892 & ~n20893;
  assign n20895 = ~n20878 & n20894;
  assign n20896 = n20878 & ~n20894;
  assign n20897 = ~n20895 & ~n20896;
  assign n20898 = n4910 & n8334;
  assign n20899 = pi98  & n8685;
  assign n20900 = pi100  & n8332;
  assign n20901 = pi99  & n8327;
  assign n20902 = ~n20900 & ~n20901;
  assign n20903 = ~n20899 & n20902;
  assign n20904 = ~n20898 & n20903;
  assign n20905 = pi50  & ~n20904;
  assign n20906 = pi50  & ~n20905;
  assign n20907 = ~n20904 & ~n20905;
  assign n20908 = ~n20906 & ~n20907;
  assign n20909 = ~n20897 & ~n20908;
  assign n20910 = n20897 & n20908;
  assign n20911 = ~n20909 & ~n20910;
  assign n20912 = n20811 & ~n20911;
  assign n20913 = ~n20811 & n20911;
  assign n20914 = ~n20912 & ~n20913;
  assign n20915 = n5664 & n7408;
  assign n20916 = pi101  & n7740;
  assign n20917 = pi103  & n7406;
  assign n20918 = pi102  & n7401;
  assign n20919 = ~n20917 & ~n20918;
  assign n20920 = ~n20916 & n20919;
  assign n20921 = ~n20915 & n20920;
  assign n20922 = pi47  & ~n20921;
  assign n20923 = pi47  & ~n20922;
  assign n20924 = ~n20921 & ~n20922;
  assign n20925 = ~n20923 & ~n20924;
  assign n20926 = n20914 & ~n20925;
  assign n20927 = n20914 & ~n20926;
  assign n20928 = ~n20925 & ~n20926;
  assign n20929 = ~n20927 & ~n20928;
  assign n20930 = ~n20670 & ~n20673;
  assign n20931 = n20929 & n20930;
  assign n20932 = ~n20929 & ~n20930;
  assign n20933 = ~n20931 & ~n20932;
  assign n20934 = n6477 & n6539;
  assign n20935 = pi104  & n6873;
  assign n20936 = pi106  & n6537;
  assign n20937 = pi105  & n6532;
  assign n20938 = ~n20936 & ~n20937;
  assign n20939 = ~n20935 & n20938;
  assign n20940 = ~n20934 & n20939;
  assign n20941 = pi44  & ~n20940;
  assign n20942 = pi44  & ~n20941;
  assign n20943 = ~n20940 & ~n20941;
  assign n20944 = ~n20942 & ~n20943;
  assign n20945 = n20933 & ~n20944;
  assign n20946 = n20933 & ~n20945;
  assign n20947 = ~n20944 & ~n20945;
  assign n20948 = ~n20946 & ~n20947;
  assign n20949 = ~n20676 & ~n20679;
  assign n20950 = n20948 & n20949;
  assign n20951 = ~n20948 & ~n20949;
  assign n20952 = ~n20950 & ~n20951;
  assign n20953 = n5739 & n7349;
  assign n20954 = pi107  & n6030;
  assign n20955 = pi109  & n5737;
  assign n20956 = pi108  & n5732;
  assign n20957 = ~n20955 & ~n20956;
  assign n20958 = ~n20954 & n20957;
  assign n20959 = ~n20953 & n20958;
  assign n20960 = pi41  & ~n20959;
  assign n20961 = pi41  & ~n20960;
  assign n20962 = ~n20959 & ~n20960;
  assign n20963 = ~n20961 & ~n20962;
  assign n20964 = n20952 & ~n20963;
  assign n20965 = n20952 & ~n20964;
  assign n20966 = ~n20963 & ~n20964;
  assign n20967 = ~n20965 & ~n20966;
  assign n20968 = ~n20682 & ~n20685;
  assign n20969 = n20967 & n20968;
  assign n20970 = ~n20967 & ~n20968;
  assign n20971 = ~n20969 & ~n20970;
  assign n20972 = n5008 & n7997;
  assign n20973 = pi110  & n5241;
  assign n20974 = pi112  & n5006;
  assign n20975 = pi111  & n5001;
  assign n20976 = ~n20974 & ~n20975;
  assign n20977 = ~n20973 & n20976;
  assign n20978 = ~n20972 & n20977;
  assign n20979 = pi38  & ~n20978;
  assign n20980 = pi38  & ~n20979;
  assign n20981 = ~n20978 & ~n20979;
  assign n20982 = ~n20980 & ~n20981;
  assign n20983 = n20971 & ~n20982;
  assign n20984 = n20971 & ~n20983;
  assign n20985 = ~n20982 & ~n20983;
  assign n20986 = ~n20984 & ~n20985;
  assign n20987 = ~n20688 & ~n20702;
  assign n20988 = n20986 & n20987;
  assign n20989 = ~n20986 & ~n20987;
  assign n20990 = ~n20988 & ~n20989;
  assign n20991 = n4271 & n8963;
  assign n20992 = pi113  & n4503;
  assign n20993 = pi115  & n4269;
  assign n20994 = pi114  & n4264;
  assign n20995 = ~n20993 & ~n20994;
  assign n20996 = ~n20992 & n20995;
  assign n20997 = ~n20991 & n20996;
  assign n20998 = pi35  & ~n20997;
  assign n20999 = pi35  & ~n20998;
  assign n21000 = ~n20997 & ~n20998;
  assign n21001 = ~n20999 & ~n21000;
  assign n21002 = ~n20990 & n21001;
  assign n21003 = n20990 & ~n21001;
  assign n21004 = ~n20810 & ~n21002;
  assign n21005 = ~n21003 & n21004;
  assign n21006 = ~n20810 & ~n21005;
  assign n21007 = ~n21003 & ~n21005;
  assign n21008 = ~n21002 & n21007;
  assign n21009 = ~n21006 & ~n21008;
  assign n21010 = n20809 & ~n21009;
  assign n21011 = ~n20809 & n21009;
  assign n21012 = ~n21010 & ~n21011;
  assign n21013 = ~n20794 & n21012;
  assign n21014 = ~n20794 & ~n21013;
  assign n21015 = n21012 & ~n21013;
  assign n21016 = ~n21014 & ~n21015;
  assign n21017 = n20778 & ~n21016;
  assign n21018 = ~n20778 & n21016;
  assign n21019 = ~n21017 & ~n21018;
  assign n21020 = ~n20763 & n21019;
  assign n21021 = ~n20763 & ~n21020;
  assign n21022 = n21019 & ~n21020;
  assign n21023 = ~n21021 & ~n21022;
  assign n21024 = ~n20472 & ~n20738;
  assign n21025 = n21023 & n21024;
  assign n21026 = ~n21023 & ~n21024;
  assign n21027 = ~n21025 & ~n21026;
  assign n21028 = ~n20741 & ~n20744;
  assign n21029 = n21027 & ~n21028;
  assign n21030 = ~n21027 & n21028;
  assign po84  = ~n21029 & ~n21030;
  assign n21032 = ~n20777 & ~n21017;
  assign n21033 = pi126  & n2180;
  assign n21034 = pi127  & n2036;
  assign n21035 = ~n21033 & ~n21034;
  assign n21036 = ~n2043 & n21035;
  assign n21037 = n13773 & n21035;
  assign n21038 = ~n21036 & ~n21037;
  assign n21039 = pi23  & ~n21038;
  assign n21040 = ~pi23  & n21038;
  assign n21041 = ~n21039 & ~n21040;
  assign n21042 = ~n21032 & ~n21041;
  assign n21043 = n21032 & n21041;
  assign n21044 = ~n21042 & ~n21043;
  assign n21045 = n2523 & n12943;
  assign n21046 = pi123  & n2667;
  assign n21047 = pi125  & n2521;
  assign n21048 = pi124  & n2516;
  assign n21049 = ~n21047 & ~n21048;
  assign n21050 = ~n21046 & n21049;
  assign n21051 = ~n21045 & n21050;
  assign n21052 = pi26  & ~n21051;
  assign n21053 = pi26  & ~n21052;
  assign n21054 = ~n21051 & ~n21052;
  assign n21055 = ~n21053 & ~n21054;
  assign n21056 = ~n20780 & ~n20791;
  assign n21057 = ~n21013 & ~n21056;
  assign n21058 = n21055 & n21057;
  assign n21059 = ~n21055 & ~n21057;
  assign n21060 = ~n21058 & ~n21059;
  assign n21061 = ~n20808 & ~n21010;
  assign n21062 = pi120  & n3225;
  assign n21063 = pi122  & n3032;
  assign n21064 = pi121  & n3027;
  assign n21065 = ~n21063 & ~n21064;
  assign n21066 = ~n21062 & n21065;
  assign n21067 = ~n3034 & n21066;
  assign n21068 = ~n11778 & n21066;
  assign n21069 = ~n21067 & ~n21068;
  assign n21070 = pi29  & ~n21069;
  assign n21071 = ~pi29  & n21069;
  assign n21072 = ~n21070 & ~n21071;
  assign n21073 = ~n21061 & ~n21072;
  assign n21074 = n21061 & n21072;
  assign n21075 = ~n21073 & ~n21074;
  assign n21076 = n3622 & n10667;
  assign n21077 = pi117  & n3814;
  assign n21078 = pi119  & n3620;
  assign n21079 = pi118  & n3615;
  assign n21080 = ~n21078 & ~n21079;
  assign n21081 = ~n21077 & n21080;
  assign n21082 = ~n21076 & n21081;
  assign n21083 = pi32  & ~n21082;
  assign n21084 = pi32  & ~n21083;
  assign n21085 = ~n21082 & ~n21083;
  assign n21086 = ~n21084 & ~n21085;
  assign n21087 = ~n21007 & n21086;
  assign n21088 = n21007 & ~n21086;
  assign n21089 = ~n21087 & ~n21088;
  assign n21090 = ~n20926 & ~n20932;
  assign n21091 = n5943 & n7408;
  assign n21092 = pi102  & n7740;
  assign n21093 = pi104  & n7406;
  assign n21094 = pi103  & n7401;
  assign n21095 = ~n21093 & ~n21094;
  assign n21096 = ~n21092 & n21095;
  assign n21097 = ~n21091 & n21096;
  assign n21098 = pi47  & ~n21097;
  assign n21099 = pi47  & ~n21098;
  assign n21100 = ~n21097 & ~n21098;
  assign n21101 = ~n21099 & ~n21100;
  assign n21102 = ~n20909 & ~n20913;
  assign n21103 = ~n20852 & ~n20858;
  assign n21104 = n3177 & n11488;
  assign n21105 = pi90  & n11847;
  assign n21106 = pi92  & n11486;
  assign n21107 = pi91  & n11481;
  assign n21108 = ~n21106 & ~n21107;
  assign n21109 = ~n21105 & n21108;
  assign n21110 = ~n21104 & n21109;
  assign n21111 = pi59  & ~n21110;
  assign n21112 = pi59  & ~n21111;
  assign n21113 = ~n21110 & ~n21111;
  assign n21114 = ~n21112 & ~n21113;
  assign n21115 = ~n20832 & ~n20837;
  assign n21116 = pi85  & n13835;
  assign n21117 = pi86  & ~n13434;
  assign n21118 = ~n21116 & ~n21117;
  assign n21119 = ~n20815 & ~n20818;
  assign n21120 = ~n21118 & n21119;
  assign n21121 = n21118 & ~n21119;
  assign n21122 = ~n21120 & ~n21121;
  assign n21123 = pi87  & n13004;
  assign n21124 = pi89  & n12625;
  assign n21125 = pi88  & n12620;
  assign n21126 = ~n21124 & ~n21125;
  assign n21127 = ~n21123 & n21126;
  assign n21128 = ~n12627 & n21127;
  assign n21129 = ~n2473 & n21127;
  assign n21130 = ~n21128 & ~n21129;
  assign n21131 = pi62  & ~n21130;
  assign n21132 = ~pi62  & n21130;
  assign n21133 = ~n21131 & ~n21132;
  assign n21134 = n21122 & ~n21133;
  assign n21135 = ~n21122 & n21133;
  assign n21136 = ~n21134 & ~n21135;
  assign n21137 = ~n21115 & n21136;
  assign n21138 = n21115 & ~n21136;
  assign n21139 = ~n21137 & ~n21138;
  assign n21140 = ~n21114 & n21139;
  assign n21141 = n21114 & ~n21139;
  assign n21142 = ~n21140 & ~n21141;
  assign n21143 = ~n21103 & n21142;
  assign n21144 = n21103 & ~n21142;
  assign n21145 = ~n21143 & ~n21144;
  assign n21146 = n3784 & n10394;
  assign n21147 = pi93  & n10744;
  assign n21148 = pi95  & n10392;
  assign n21149 = pi94  & n10387;
  assign n21150 = ~n21148 & ~n21149;
  assign n21151 = ~n21147 & n21150;
  assign n21152 = ~n21146 & n21151;
  assign n21153 = pi56  & ~n21152;
  assign n21154 = pi56  & ~n21153;
  assign n21155 = ~n21152 & ~n21153;
  assign n21156 = ~n21154 & ~n21155;
  assign n21157 = n21145 & ~n21156;
  assign n21158 = n21145 & ~n21157;
  assign n21159 = ~n21156 & ~n21157;
  assign n21160 = ~n21158 & ~n21159;
  assign n21161 = ~n20871 & ~n20877;
  assign n21162 = n21160 & n21161;
  assign n21163 = ~n21160 & ~n21161;
  assign n21164 = ~n21162 & ~n21163;
  assign n21165 = n4454 & n9310;
  assign n21166 = pi96  & n9701;
  assign n21167 = pi98  & n9308;
  assign n21168 = pi97  & n9303;
  assign n21169 = ~n21167 & ~n21168;
  assign n21170 = ~n21166 & n21169;
  assign n21171 = ~n21165 & n21170;
  assign n21172 = pi53  & ~n21171;
  assign n21173 = pi53  & ~n21172;
  assign n21174 = ~n21171 & ~n21172;
  assign n21175 = ~n21173 & ~n21174;
  assign n21176 = n21164 & ~n21175;
  assign n21177 = n21164 & ~n21176;
  assign n21178 = ~n21175 & ~n21176;
  assign n21179 = ~n21177 & ~n21178;
  assign n21180 = ~n20893 & ~n20895;
  assign n21181 = n21179 & ~n21180;
  assign n21182 = ~n21179 & n21180;
  assign n21183 = ~n21181 & ~n21182;
  assign n21184 = n5169 & n8334;
  assign n21185 = pi99  & n8685;
  assign n21186 = pi101  & n8332;
  assign n21187 = pi100  & n8327;
  assign n21188 = ~n21186 & ~n21187;
  assign n21189 = ~n21185 & n21188;
  assign n21190 = ~n21184 & n21189;
  assign n21191 = pi50  & ~n21190;
  assign n21192 = pi50  & ~n21191;
  assign n21193 = ~n21190 & ~n21191;
  assign n21194 = ~n21192 & ~n21193;
  assign n21195 = ~n21183 & n21194;
  assign n21196 = n21183 & ~n21194;
  assign n21197 = ~n21195 & ~n21196;
  assign n21198 = ~n21102 & n21197;
  assign n21199 = ~n21102 & ~n21198;
  assign n21200 = n21197 & ~n21198;
  assign n21201 = ~n21199 & ~n21200;
  assign n21202 = ~n21101 & ~n21201;
  assign n21203 = n21101 & n21201;
  assign n21204 = ~n21202 & ~n21203;
  assign n21205 = ~n21090 & n21204;
  assign n21206 = n21090 & ~n21204;
  assign n21207 = ~n21205 & ~n21206;
  assign n21208 = n6539 & n6775;
  assign n21209 = pi105  & n6873;
  assign n21210 = pi107  & n6537;
  assign n21211 = pi106  & n6532;
  assign n21212 = ~n21210 & ~n21211;
  assign n21213 = ~n21209 & n21212;
  assign n21214 = ~n21208 & n21213;
  assign n21215 = pi44  & ~n21214;
  assign n21216 = pi44  & ~n21215;
  assign n21217 = ~n21214 & ~n21215;
  assign n21218 = ~n21216 & ~n21217;
  assign n21219 = n21207 & ~n21218;
  assign n21220 = n21207 & ~n21219;
  assign n21221 = ~n21218 & ~n21219;
  assign n21222 = ~n21220 & ~n21221;
  assign n21223 = ~n20945 & ~n20951;
  assign n21224 = n21222 & n21223;
  assign n21225 = ~n21222 & ~n21223;
  assign n21226 = ~n21224 & ~n21225;
  assign n21227 = n5739 & n7665;
  assign n21228 = pi108  & n6030;
  assign n21229 = pi110  & n5737;
  assign n21230 = pi109  & n5732;
  assign n21231 = ~n21229 & ~n21230;
  assign n21232 = ~n21228 & n21231;
  assign n21233 = ~n21227 & n21232;
  assign n21234 = pi41  & ~n21233;
  assign n21235 = pi41  & ~n21234;
  assign n21236 = ~n21233 & ~n21234;
  assign n21237 = ~n21235 & ~n21236;
  assign n21238 = n21226 & ~n21237;
  assign n21239 = n21226 & ~n21238;
  assign n21240 = ~n21237 & ~n21238;
  assign n21241 = ~n21239 & ~n21240;
  assign n21242 = ~n20964 & ~n20970;
  assign n21243 = n21241 & n21242;
  assign n21244 = ~n21241 & ~n21242;
  assign n21245 = ~n21243 & ~n21244;
  assign n21246 = n5008 & n8612;
  assign n21247 = pi111  & n5241;
  assign n21248 = pi113  & n5006;
  assign n21249 = pi112  & n5001;
  assign n21250 = ~n21248 & ~n21249;
  assign n21251 = ~n21247 & n21250;
  assign n21252 = ~n21246 & n21251;
  assign n21253 = pi38  & ~n21252;
  assign n21254 = pi38  & ~n21253;
  assign n21255 = ~n21252 & ~n21253;
  assign n21256 = ~n21254 & ~n21255;
  assign n21257 = n21245 & ~n21256;
  assign n21258 = n21245 & ~n21257;
  assign n21259 = ~n21256 & ~n21257;
  assign n21260 = ~n21258 & ~n21259;
  assign n21261 = ~n20983 & ~n20989;
  assign n21262 = n21260 & n21261;
  assign n21263 = ~n21260 & ~n21261;
  assign n21264 = ~n21262 & ~n21263;
  assign n21265 = n4271 & n9614;
  assign n21266 = pi114  & n4503;
  assign n21267 = pi116  & n4269;
  assign n21268 = pi115  & n4264;
  assign n21269 = ~n21267 & ~n21268;
  assign n21270 = ~n21266 & n21269;
  assign n21271 = ~n21265 & n21270;
  assign n21272 = pi35  & ~n21271;
  assign n21273 = pi35  & ~n21272;
  assign n21274 = ~n21271 & ~n21272;
  assign n21275 = ~n21273 & ~n21274;
  assign n21276 = n21264 & ~n21275;
  assign n21277 = n21264 & ~n21276;
  assign n21278 = ~n21275 & ~n21276;
  assign n21279 = ~n21277 & ~n21278;
  assign n21280 = ~n21089 & ~n21279;
  assign n21281 = n21089 & n21279;
  assign n21282 = ~n21280 & ~n21281;
  assign n21283 = n21075 & n21282;
  assign n21284 = n21075 & ~n21283;
  assign n21285 = n21282 & ~n21283;
  assign n21286 = ~n21284 & ~n21285;
  assign n21287 = n21060 & ~n21286;
  assign n21288 = ~n21060 & n21286;
  assign n21289 = ~n21287 & ~n21288;
  assign n21290 = n21044 & n21289;
  assign n21291 = n21044 & ~n21290;
  assign n21292 = n21289 & ~n21290;
  assign n21293 = ~n21291 & ~n21292;
  assign n21294 = ~n20760 & ~n21020;
  assign n21295 = n21293 & n21294;
  assign n21296 = ~n21293 & ~n21294;
  assign n21297 = ~n21295 & ~n21296;
  assign n21298 = ~n21026 & ~n21029;
  assign n21299 = n21297 & ~n21298;
  assign n21300 = ~n21297 & n21298;
  assign po85  = ~n21299 & ~n21300;
  assign n21302 = ~n21296 & ~n21299;
  assign n21303 = ~n21042 & ~n21290;
  assign n21304 = ~n21059 & ~n21287;
  assign n21305 = pi127  & n2180;
  assign n21306 = n2043 & n13770;
  assign n21307 = ~n21305 & ~n21306;
  assign n21308 = pi23  & ~n21307;
  assign n21309 = pi23  & ~n21308;
  assign n21310 = ~n21307 & ~n21308;
  assign n21311 = ~n21309 & ~n21310;
  assign n21312 = ~n21304 & ~n21311;
  assign n21313 = ~n21304 & ~n21312;
  assign n21314 = ~n21311 & ~n21312;
  assign n21315 = ~n21313 & ~n21314;
  assign n21316 = n2523 & n13344;
  assign n21317 = pi124  & n2667;
  assign n21318 = pi126  & n2521;
  assign n21319 = pi125  & n2516;
  assign n21320 = ~n21318 & ~n21319;
  assign n21321 = ~n21317 & n21320;
  assign n21322 = ~n21316 & n21321;
  assign n21323 = pi26  & ~n21322;
  assign n21324 = pi26  & ~n21323;
  assign n21325 = ~n21322 & ~n21323;
  assign n21326 = ~n21324 & ~n21325;
  assign n21327 = ~n21073 & ~n21283;
  assign n21328 = n21326 & n21327;
  assign n21329 = ~n21326 & ~n21327;
  assign n21330 = ~n21328 & ~n21329;
  assign n21331 = n3034 & n12158;
  assign n21332 = pi121  & n3225;
  assign n21333 = pi123  & n3032;
  assign n21334 = pi122  & n3027;
  assign n21335 = ~n21333 & ~n21334;
  assign n21336 = ~n21332 & n21335;
  assign n21337 = ~n21331 & n21336;
  assign n21338 = pi29  & ~n21337;
  assign n21339 = pi29  & ~n21338;
  assign n21340 = ~n21337 & ~n21338;
  assign n21341 = ~n21339 & ~n21340;
  assign n21342 = ~n21007 & ~n21086;
  assign n21343 = ~n21280 & ~n21342;
  assign n21344 = ~n21341 & ~n21343;
  assign n21345 = ~n21341 & ~n21344;
  assign n21346 = ~n21343 & ~n21344;
  assign n21347 = ~n21345 & ~n21346;
  assign n21348 = n3622 & n11028;
  assign n21349 = pi118  & n3814;
  assign n21350 = pi120  & n3620;
  assign n21351 = pi119  & n3615;
  assign n21352 = ~n21350 & ~n21351;
  assign n21353 = ~n21349 & n21352;
  assign n21354 = ~n21348 & n21353;
  assign n21355 = pi32  & ~n21354;
  assign n21356 = pi32  & ~n21355;
  assign n21357 = ~n21354 & ~n21355;
  assign n21358 = ~n21356 & ~n21357;
  assign n21359 = ~n21263 & ~n21276;
  assign n21360 = n21358 & n21359;
  assign n21361 = ~n21358 & ~n21359;
  assign n21362 = ~n21360 & ~n21361;
  assign n21363 = n4271 & n9958;
  assign n21364 = pi115  & n4503;
  assign n21365 = pi117  & n4269;
  assign n21366 = pi116  & n4264;
  assign n21367 = ~n21365 & ~n21366;
  assign n21368 = ~n21364 & n21367;
  assign n21369 = ~n21363 & n21368;
  assign n21370 = pi35  & ~n21369;
  assign n21371 = pi35  & ~n21370;
  assign n21372 = ~n21369 & ~n21370;
  assign n21373 = ~n21371 & ~n21372;
  assign n21374 = ~n21244 & ~n21257;
  assign n21375 = ~n21205 & ~n21219;
  assign n21376 = n6539 & n7060;
  assign n21377 = pi106  & n6873;
  assign n21378 = pi108  & n6537;
  assign n21379 = pi107  & n6532;
  assign n21380 = ~n21378 & ~n21379;
  assign n21381 = ~n21377 & n21380;
  assign n21382 = ~n21376 & n21381;
  assign n21383 = pi44  & ~n21382;
  assign n21384 = pi44  & ~n21383;
  assign n21385 = ~n21382 & ~n21383;
  assign n21386 = ~n21384 & ~n21385;
  assign n21387 = ~n21198 & ~n21202;
  assign n21388 = ~n21163 & ~n21176;
  assign n21389 = n4684 & n9310;
  assign n21390 = pi97  & n9701;
  assign n21391 = pi99  & n9308;
  assign n21392 = pi98  & n9303;
  assign n21393 = ~n21391 & ~n21392;
  assign n21394 = ~n21390 & n21393;
  assign n21395 = ~n21389 & n21394;
  assign n21396 = pi53  & ~n21395;
  assign n21397 = pi53  & ~n21396;
  assign n21398 = ~n21395 & ~n21396;
  assign n21399 = ~n21397 & ~n21398;
  assign n21400 = ~n21143 & ~n21157;
  assign n21401 = ~n21121 & ~n21134;
  assign n21402 = pi86  & n13835;
  assign n21403 = pi87  & ~n13434;
  assign n21404 = ~n21402 & ~n21403;
  assign n21405 = ~n21118 & n21404;
  assign n21406 = n21118 & ~n21404;
  assign n21407 = ~n21405 & ~n21406;
  assign n21408 = pi88  & n13004;
  assign n21409 = pi90  & n12625;
  assign n21410 = pi89  & n12620;
  assign n21411 = ~n21409 & ~n21410;
  assign n21412 = ~n21408 & n21411;
  assign n21413 = ~n12627 & n21412;
  assign n21414 = ~n2801 & n21412;
  assign n21415 = ~n21413 & ~n21414;
  assign n21416 = pi62  & ~n21415;
  assign n21417 = ~pi62  & n21415;
  assign n21418 = ~n21416 & ~n21417;
  assign n21419 = n21407 & ~n21418;
  assign n21420 = ~n21407 & n21418;
  assign n21421 = ~n21419 & ~n21420;
  assign n21422 = ~n21401 & n21421;
  assign n21423 = n21401 & ~n21421;
  assign n21424 = ~n21422 & ~n21423;
  assign n21425 = n3371 & n11488;
  assign n21426 = pi91  & n11847;
  assign n21427 = pi93  & n11486;
  assign n21428 = pi92  & n11481;
  assign n21429 = ~n21427 & ~n21428;
  assign n21430 = ~n21426 & n21429;
  assign n21431 = ~n21425 & n21430;
  assign n21432 = pi59  & ~n21431;
  assign n21433 = pi59  & ~n21432;
  assign n21434 = ~n21431 & ~n21432;
  assign n21435 = ~n21433 & ~n21434;
  assign n21436 = n21424 & ~n21435;
  assign n21437 = n21424 & ~n21436;
  assign n21438 = ~n21435 & ~n21436;
  assign n21439 = ~n21437 & ~n21438;
  assign n21440 = ~n21137 & ~n21140;
  assign n21441 = n21439 & n21440;
  assign n21442 = ~n21439 & ~n21440;
  assign n21443 = ~n21441 & ~n21442;
  assign n21444 = n4001 & n10394;
  assign n21445 = pi94  & n10744;
  assign n21446 = pi96  & n10392;
  assign n21447 = pi95  & n10387;
  assign n21448 = ~n21446 & ~n21447;
  assign n21449 = ~n21445 & n21448;
  assign n21450 = ~n21444 & n21449;
  assign n21451 = pi56  & ~n21450;
  assign n21452 = pi56  & ~n21451;
  assign n21453 = ~n21450 & ~n21451;
  assign n21454 = ~n21452 & ~n21453;
  assign n21455 = ~n21443 & n21454;
  assign n21456 = n21443 & ~n21454;
  assign n21457 = ~n21455 & ~n21456;
  assign n21458 = ~n21400 & n21457;
  assign n21459 = n21400 & ~n21457;
  assign n21460 = ~n21458 & ~n21459;
  assign n21461 = ~n21399 & n21460;
  assign n21462 = n21399 & ~n21460;
  assign n21463 = ~n21461 & ~n21462;
  assign n21464 = ~n21388 & n21463;
  assign n21465 = n21388 & ~n21463;
  assign n21466 = ~n21464 & ~n21465;
  assign n21467 = n5413 & n8334;
  assign n21468 = pi100  & n8685;
  assign n21469 = pi102  & n8332;
  assign n21470 = pi101  & n8327;
  assign n21471 = ~n21469 & ~n21470;
  assign n21472 = ~n21468 & n21471;
  assign n21473 = ~n21467 & n21472;
  assign n21474 = pi50  & ~n21473;
  assign n21475 = pi50  & ~n21474;
  assign n21476 = ~n21473 & ~n21474;
  assign n21477 = ~n21475 & ~n21476;
  assign n21478 = n21466 & ~n21477;
  assign n21479 = n21466 & ~n21478;
  assign n21480 = ~n21477 & ~n21478;
  assign n21481 = ~n21479 & ~n21480;
  assign n21482 = ~n21182 & ~n21196;
  assign n21483 = ~n21481 & ~n21482;
  assign n21484 = ~n21481 & ~n21483;
  assign n21485 = ~n21482 & ~n21483;
  assign n21486 = ~n21484 & ~n21485;
  assign n21487 = n6207 & n7408;
  assign n21488 = pi103  & n7740;
  assign n21489 = pi105  & n7406;
  assign n21490 = pi104  & n7401;
  assign n21491 = ~n21489 & ~n21490;
  assign n21492 = ~n21488 & n21491;
  assign n21493 = ~n21487 & n21492;
  assign n21494 = pi47  & ~n21493;
  assign n21495 = pi47  & ~n21494;
  assign n21496 = ~n21493 & ~n21494;
  assign n21497 = ~n21495 & ~n21496;
  assign n21498 = ~n21486 & n21497;
  assign n21499 = n21486 & ~n21497;
  assign n21500 = ~n21498 & ~n21499;
  assign n21501 = ~n21387 & ~n21500;
  assign n21502 = n21387 & n21500;
  assign n21503 = ~n21501 & ~n21502;
  assign n21504 = ~n21386 & n21503;
  assign n21505 = n21386 & ~n21503;
  assign n21506 = ~n21504 & ~n21505;
  assign n21507 = ~n21375 & n21506;
  assign n21508 = n21375 & ~n21506;
  assign n21509 = ~n21507 & ~n21508;
  assign n21510 = n5739 & n7970;
  assign n21511 = pi109  & n6030;
  assign n21512 = pi111  & n5737;
  assign n21513 = pi110  & n5732;
  assign n21514 = ~n21512 & ~n21513;
  assign n21515 = ~n21511 & n21514;
  assign n21516 = ~n21510 & n21515;
  assign n21517 = pi41  & ~n21516;
  assign n21518 = pi41  & ~n21517;
  assign n21519 = ~n21516 & ~n21517;
  assign n21520 = ~n21518 & ~n21519;
  assign n21521 = n21509 & ~n21520;
  assign n21522 = n21509 & ~n21521;
  assign n21523 = ~n21520 & ~n21521;
  assign n21524 = ~n21522 & ~n21523;
  assign n21525 = ~n21225 & ~n21238;
  assign n21526 = n21524 & n21525;
  assign n21527 = ~n21524 & ~n21525;
  assign n21528 = ~n21526 & ~n21527;
  assign n21529 = n5008 & n8936;
  assign n21530 = pi112  & n5241;
  assign n21531 = pi114  & n5006;
  assign n21532 = pi113  & n5001;
  assign n21533 = ~n21531 & ~n21532;
  assign n21534 = ~n21530 & n21533;
  assign n21535 = ~n21529 & n21534;
  assign n21536 = pi38  & ~n21535;
  assign n21537 = pi38  & ~n21536;
  assign n21538 = ~n21535 & ~n21536;
  assign n21539 = ~n21537 & ~n21538;
  assign n21540 = ~n21528 & n21539;
  assign n21541 = n21528 & ~n21539;
  assign n21542 = ~n21540 & ~n21541;
  assign n21543 = ~n21374 & n21542;
  assign n21544 = ~n21374 & ~n21543;
  assign n21545 = n21542 & ~n21543;
  assign n21546 = ~n21544 & ~n21545;
  assign n21547 = ~n21373 & ~n21546;
  assign n21548 = ~n21373 & ~n21547;
  assign n21549 = ~n21546 & ~n21547;
  assign n21550 = ~n21548 & ~n21549;
  assign n21551 = n21362 & ~n21550;
  assign n21552 = n21362 & ~n21551;
  assign n21553 = ~n21550 & ~n21551;
  assign n21554 = ~n21552 & ~n21553;
  assign n21555 = ~n21347 & n21554;
  assign n21556 = n21347 & ~n21554;
  assign n21557 = ~n21555 & ~n21556;
  assign n21558 = n21330 & ~n21557;
  assign n21559 = n21330 & ~n21558;
  assign n21560 = ~n21557 & ~n21558;
  assign n21561 = ~n21559 & ~n21560;
  assign n21562 = ~n21315 & n21561;
  assign n21563 = n21315 & ~n21561;
  assign n21564 = ~n21562 & ~n21563;
  assign n21565 = ~n21303 & ~n21564;
  assign n21566 = ~n21303 & ~n21565;
  assign n21567 = ~n21564 & ~n21565;
  assign n21568 = ~n21566 & ~n21567;
  assign n21569 = ~n21302 & ~n21568;
  assign n21570 = n21302 & n21568;
  assign po86  = ~n21569 & ~n21570;
  assign n21572 = ~n21565 & ~n21569;
  assign n21573 = ~n21315 & ~n21561;
  assign n21574 = ~n21312 & ~n21573;
  assign n21575 = ~n21329 & ~n21558;
  assign n21576 = n2523 & n13742;
  assign n21577 = pi125  & n2667;
  assign n21578 = pi127  & n2521;
  assign n21579 = pi126  & n2516;
  assign n21580 = ~n21578 & ~n21579;
  assign n21581 = ~n21577 & n21580;
  assign n21582 = ~n21576 & n21581;
  assign n21583 = pi26  & ~n21582;
  assign n21584 = pi26  & ~n21583;
  assign n21585 = ~n21582 & ~n21583;
  assign n21586 = ~n21584 & ~n21585;
  assign n21587 = ~n21575 & ~n21586;
  assign n21588 = ~n21575 & ~n21587;
  assign n21589 = ~n21586 & ~n21587;
  assign n21590 = ~n21588 & ~n21589;
  assign n21591 = ~n21347 & ~n21554;
  assign n21592 = ~n21344 & ~n21591;
  assign n21593 = n3034 & n12189;
  assign n21594 = pi122  & n3225;
  assign n21595 = pi124  & n3032;
  assign n21596 = pi123  & n3027;
  assign n21597 = ~n21595 & ~n21596;
  assign n21598 = ~n21594 & n21597;
  assign n21599 = ~n21593 & n21598;
  assign n21600 = pi29  & ~n21599;
  assign n21601 = pi29  & ~n21600;
  assign n21602 = ~n21599 & ~n21600;
  assign n21603 = ~n21601 & ~n21602;
  assign n21604 = ~n21592 & n21603;
  assign n21605 = n21592 & ~n21603;
  assign n21606 = ~n21604 & ~n21605;
  assign n21607 = n3622 & n11389;
  assign n21608 = pi119  & n3814;
  assign n21609 = pi121  & n3620;
  assign n21610 = pi120  & n3615;
  assign n21611 = ~n21609 & ~n21610;
  assign n21612 = ~n21608 & n21611;
  assign n21613 = ~n21607 & n21612;
  assign n21614 = pi32  & ~n21613;
  assign n21615 = pi32  & ~n21614;
  assign n21616 = ~n21613 & ~n21614;
  assign n21617 = ~n21615 & ~n21616;
  assign n21618 = ~n21361 & ~n21551;
  assign n21619 = n21617 & n21618;
  assign n21620 = ~n21617 & ~n21618;
  assign n21621 = ~n21619 & ~n21620;
  assign n21622 = ~n21543 & ~n21547;
  assign n21623 = ~n21527 & ~n21541;
  assign n21624 = ~n21501 & ~n21504;
  assign n21625 = ~n21486 & ~n21497;
  assign n21626 = ~n21483 & ~n21625;
  assign n21627 = ~n21422 & ~n21436;
  assign n21628 = ~n21405 & ~n21419;
  assign n21629 = pi87  & n13835;
  assign n21630 = pi88  & ~n13434;
  assign n21631 = ~n21629 & ~n21630;
  assign n21632 = ~pi23  & ~n21631;
  assign n21633 = pi23  & n21631;
  assign n21634 = ~n21632 & ~n21633;
  assign n21635 = ~n21404 & n21634;
  assign n21636 = n21404 & ~n21634;
  assign n21637 = ~n21635 & ~n21636;
  assign n21638 = n2978 & n12627;
  assign n21639 = pi89  & n13004;
  assign n21640 = pi91  & n12625;
  assign n21641 = pi90  & n12620;
  assign n21642 = ~n21640 & ~n21641;
  assign n21643 = ~n21639 & n21642;
  assign n21644 = ~n21638 & n21643;
  assign n21645 = pi62  & ~n21644;
  assign n21646 = pi62  & ~n21645;
  assign n21647 = ~n21644 & ~n21645;
  assign n21648 = ~n21646 & ~n21647;
  assign n21649 = n21637 & ~n21648;
  assign n21650 = n21637 & ~n21649;
  assign n21651 = ~n21648 & ~n21649;
  assign n21652 = ~n21650 & ~n21651;
  assign n21653 = ~n21628 & n21652;
  assign n21654 = n21628 & ~n21652;
  assign n21655 = ~n21653 & ~n21654;
  assign n21656 = n3565 & n11488;
  assign n21657 = pi92  & n11847;
  assign n21658 = pi94  & n11486;
  assign n21659 = pi93  & n11481;
  assign n21660 = ~n21658 & ~n21659;
  assign n21661 = ~n21657 & n21660;
  assign n21662 = ~n21656 & n21661;
  assign n21663 = pi59  & ~n21662;
  assign n21664 = pi59  & ~n21663;
  assign n21665 = ~n21662 & ~n21663;
  assign n21666 = ~n21664 & ~n21665;
  assign n21667 = ~n21655 & ~n21666;
  assign n21668 = n21655 & n21666;
  assign n21669 = ~n21667 & ~n21668;
  assign n21670 = n21627 & ~n21669;
  assign n21671 = ~n21627 & n21669;
  assign n21672 = ~n21670 & ~n21671;
  assign n21673 = n4211 & n10394;
  assign n21674 = pi95  & n10744;
  assign n21675 = pi97  & n10392;
  assign n21676 = pi96  & n10387;
  assign n21677 = ~n21675 & ~n21676;
  assign n21678 = ~n21674 & n21677;
  assign n21679 = ~n21673 & n21678;
  assign n21680 = pi56  & ~n21679;
  assign n21681 = pi56  & ~n21680;
  assign n21682 = ~n21679 & ~n21680;
  assign n21683 = ~n21681 & ~n21682;
  assign n21684 = ~n21442 & ~n21456;
  assign n21685 = ~n21683 & ~n21684;
  assign n21686 = n21683 & n21684;
  assign n21687 = ~n21685 & ~n21686;
  assign n21688 = n21672 & n21687;
  assign n21689 = ~n21672 & ~n21687;
  assign n21690 = ~n21688 & ~n21689;
  assign n21691 = n4910 & n9310;
  assign n21692 = pi98  & n9701;
  assign n21693 = pi100  & n9308;
  assign n21694 = pi99  & n9303;
  assign n21695 = ~n21693 & ~n21694;
  assign n21696 = ~n21692 & n21695;
  assign n21697 = ~n21691 & n21696;
  assign n21698 = pi53  & ~n21697;
  assign n21699 = pi53  & ~n21698;
  assign n21700 = ~n21697 & ~n21698;
  assign n21701 = ~n21699 & ~n21700;
  assign n21702 = n21690 & ~n21701;
  assign n21703 = n21690 & ~n21702;
  assign n21704 = ~n21701 & ~n21702;
  assign n21705 = ~n21703 & ~n21704;
  assign n21706 = ~n21458 & ~n21461;
  assign n21707 = n21705 & n21706;
  assign n21708 = ~n21705 & ~n21706;
  assign n21709 = ~n21707 & ~n21708;
  assign n21710 = n5664 & n8334;
  assign n21711 = pi101  & n8685;
  assign n21712 = pi103  & n8332;
  assign n21713 = pi102  & n8327;
  assign n21714 = ~n21712 & ~n21713;
  assign n21715 = ~n21711 & n21714;
  assign n21716 = ~n21710 & n21715;
  assign n21717 = pi50  & ~n21716;
  assign n21718 = pi50  & ~n21717;
  assign n21719 = ~n21716 & ~n21717;
  assign n21720 = ~n21718 & ~n21719;
  assign n21721 = n21709 & ~n21720;
  assign n21722 = n21709 & ~n21721;
  assign n21723 = ~n21720 & ~n21721;
  assign n21724 = ~n21722 & ~n21723;
  assign n21725 = ~n21464 & ~n21478;
  assign n21726 = n21724 & n21725;
  assign n21727 = ~n21724 & ~n21725;
  assign n21728 = ~n21726 & ~n21727;
  assign n21729 = n6477 & n7408;
  assign n21730 = pi104  & n7740;
  assign n21731 = pi106  & n7406;
  assign n21732 = pi105  & n7401;
  assign n21733 = ~n21731 & ~n21732;
  assign n21734 = ~n21730 & n21733;
  assign n21735 = ~n21729 & n21734;
  assign n21736 = pi47  & ~n21735;
  assign n21737 = pi47  & ~n21736;
  assign n21738 = ~n21735 & ~n21736;
  assign n21739 = ~n21737 & ~n21738;
  assign n21740 = n21728 & ~n21739;
  assign n21741 = n21728 & ~n21740;
  assign n21742 = ~n21739 & ~n21740;
  assign n21743 = ~n21741 & ~n21742;
  assign n21744 = ~n21626 & n21743;
  assign n21745 = n21626 & ~n21743;
  assign n21746 = ~n21744 & ~n21745;
  assign n21747 = n6539 & n7349;
  assign n21748 = pi107  & n6873;
  assign n21749 = pi109  & n6537;
  assign n21750 = pi108  & n6532;
  assign n21751 = ~n21749 & ~n21750;
  assign n21752 = ~n21748 & n21751;
  assign n21753 = ~n21747 & n21752;
  assign n21754 = pi44  & ~n21753;
  assign n21755 = pi44  & ~n21754;
  assign n21756 = ~n21753 & ~n21754;
  assign n21757 = ~n21755 & ~n21756;
  assign n21758 = ~n21746 & ~n21757;
  assign n21759 = n21746 & n21757;
  assign n21760 = ~n21758 & ~n21759;
  assign n21761 = n21624 & ~n21760;
  assign n21762 = ~n21624 & n21760;
  assign n21763 = ~n21761 & ~n21762;
  assign n21764 = n5739 & n7997;
  assign n21765 = pi110  & n6030;
  assign n21766 = pi112  & n5737;
  assign n21767 = pi111  & n5732;
  assign n21768 = ~n21766 & ~n21767;
  assign n21769 = ~n21765 & n21768;
  assign n21770 = ~n21764 & n21769;
  assign n21771 = pi41  & ~n21770;
  assign n21772 = pi41  & ~n21771;
  assign n21773 = ~n21770 & ~n21771;
  assign n21774 = ~n21772 & ~n21773;
  assign n21775 = n21763 & ~n21774;
  assign n21776 = n21763 & ~n21775;
  assign n21777 = ~n21774 & ~n21775;
  assign n21778 = ~n21776 & ~n21777;
  assign n21779 = ~n21507 & ~n21521;
  assign n21780 = n21778 & n21779;
  assign n21781 = ~n21778 & ~n21779;
  assign n21782 = ~n21780 & ~n21781;
  assign n21783 = n5008 & n8963;
  assign n21784 = pi113  & n5241;
  assign n21785 = pi115  & n5006;
  assign n21786 = pi114  & n5001;
  assign n21787 = ~n21785 & ~n21786;
  assign n21788 = ~n21784 & n21787;
  assign n21789 = ~n21783 & n21788;
  assign n21790 = pi38  & ~n21789;
  assign n21791 = pi38  & ~n21790;
  assign n21792 = ~n21789 & ~n21790;
  assign n21793 = ~n21791 & ~n21792;
  assign n21794 = ~n21782 & n21793;
  assign n21795 = n21782 & ~n21793;
  assign n21796 = ~n21623 & ~n21794;
  assign n21797 = ~n21795 & n21796;
  assign n21798 = ~n21623 & ~n21797;
  assign n21799 = ~n21795 & ~n21797;
  assign n21800 = ~n21794 & n21799;
  assign n21801 = ~n21798 & ~n21800;
  assign n21802 = n4271 & n9984;
  assign n21803 = pi116  & n4503;
  assign n21804 = pi118  & n4269;
  assign n21805 = pi117  & n4264;
  assign n21806 = ~n21804 & ~n21805;
  assign n21807 = ~n21803 & n21806;
  assign n21808 = ~n21802 & n21807;
  assign n21809 = pi35  & ~n21808;
  assign n21810 = pi35  & ~n21809;
  assign n21811 = ~n21808 & ~n21809;
  assign n21812 = ~n21810 & ~n21811;
  assign n21813 = n21801 & n21812;
  assign n21814 = ~n21801 & ~n21812;
  assign n21815 = ~n21813 & ~n21814;
  assign n21816 = ~n21622 & n21815;
  assign n21817 = n21622 & ~n21815;
  assign n21818 = ~n21816 & ~n21817;
  assign n21819 = n21621 & n21818;
  assign n21820 = ~n21621 & ~n21818;
  assign n21821 = ~n21819 & ~n21820;
  assign n21822 = ~n21606 & n21821;
  assign n21823 = ~n21606 & ~n21822;
  assign n21824 = n21821 & ~n21822;
  assign n21825 = ~n21823 & ~n21824;
  assign n21826 = ~n21590 & n21825;
  assign n21827 = n21590 & ~n21825;
  assign n21828 = ~n21826 & ~n21827;
  assign n21829 = ~n21574 & ~n21828;
  assign n21830 = ~n21574 & ~n21829;
  assign n21831 = ~n21828 & ~n21829;
  assign n21832 = ~n21830 & ~n21831;
  assign n21833 = ~n21572 & ~n21832;
  assign n21834 = n21572 & n21832;
  assign po87  = ~n21833 & ~n21834;
  assign n21836 = ~n21829 & ~n21833;
  assign n21837 = ~n21590 & ~n21825;
  assign n21838 = ~n21587 & ~n21837;
  assign n21839 = n3034 & n12943;
  assign n21840 = pi123  & n3225;
  assign n21841 = pi125  & n3032;
  assign n21842 = pi124  & n3027;
  assign n21843 = ~n21841 & ~n21842;
  assign n21844 = ~n21840 & n21843;
  assign n21845 = ~n21839 & n21844;
  assign n21846 = pi29  & ~n21845;
  assign n21847 = pi29  & ~n21846;
  assign n21848 = ~n21845 & ~n21846;
  assign n21849 = ~n21847 & ~n21848;
  assign n21850 = ~n21620 & ~n21819;
  assign n21851 = ~n21849 & ~n21850;
  assign n21852 = ~n21849 & ~n21851;
  assign n21853 = ~n21850 & ~n21851;
  assign n21854 = ~n21852 & ~n21853;
  assign n21855 = ~n21814 & ~n21816;
  assign n21856 = pi120  & n3814;
  assign n21857 = pi122  & n3620;
  assign n21858 = pi121  & n3615;
  assign n21859 = ~n21857 & ~n21858;
  assign n21860 = ~n21856 & n21859;
  assign n21861 = ~n3622 & n21860;
  assign n21862 = ~n11778 & n21860;
  assign n21863 = ~n21861 & ~n21862;
  assign n21864 = pi32  & ~n21863;
  assign n21865 = ~pi32  & n21863;
  assign n21866 = ~n21864 & ~n21865;
  assign n21867 = ~n21855 & ~n21866;
  assign n21868 = n21855 & n21866;
  assign n21869 = ~n21867 & ~n21868;
  assign n21870 = ~n21721 & ~n21727;
  assign n21871 = n5943 & n8334;
  assign n21872 = pi102  & n8685;
  assign n21873 = pi104  & n8332;
  assign n21874 = pi103  & n8327;
  assign n21875 = ~n21873 & ~n21874;
  assign n21876 = ~n21872 & n21875;
  assign n21877 = ~n21871 & n21876;
  assign n21878 = pi50  & ~n21877;
  assign n21879 = pi50  & ~n21878;
  assign n21880 = ~n21877 & ~n21878;
  assign n21881 = ~n21879 & ~n21880;
  assign n21882 = ~n21702 & ~n21708;
  assign n21883 = ~n21628 & ~n21652;
  assign n21884 = ~n21649 & ~n21883;
  assign n21885 = pi88  & n13835;
  assign n21886 = pi89  & ~n13434;
  assign n21887 = ~n21885 & ~n21886;
  assign n21888 = ~n21632 & ~n21635;
  assign n21889 = ~n21887 & n21888;
  assign n21890 = n21887 & ~n21888;
  assign n21891 = ~n21889 & ~n21890;
  assign n21892 = pi90  & n13004;
  assign n21893 = pi92  & n12625;
  assign n21894 = pi91  & n12620;
  assign n21895 = ~n21893 & ~n21894;
  assign n21896 = ~n21892 & n21895;
  assign n21897 = ~n12627 & n21896;
  assign n21898 = ~n3177 & n21896;
  assign n21899 = ~n21897 & ~n21898;
  assign n21900 = pi62  & ~n21899;
  assign n21901 = ~pi62  & n21899;
  assign n21902 = ~n21900 & ~n21901;
  assign n21903 = n21891 & ~n21902;
  assign n21904 = ~n21891 & n21902;
  assign n21905 = ~n21903 & ~n21904;
  assign n21906 = ~n21884 & n21905;
  assign n21907 = n21884 & ~n21905;
  assign n21908 = ~n21906 & ~n21907;
  assign n21909 = n3784 & n11488;
  assign n21910 = pi93  & n11847;
  assign n21911 = pi95  & n11486;
  assign n21912 = pi94  & n11481;
  assign n21913 = ~n21911 & ~n21912;
  assign n21914 = ~n21910 & n21913;
  assign n21915 = ~n21909 & n21914;
  assign n21916 = pi59  & ~n21915;
  assign n21917 = pi59  & ~n21916;
  assign n21918 = ~n21915 & ~n21916;
  assign n21919 = ~n21917 & ~n21918;
  assign n21920 = n21908 & ~n21919;
  assign n21921 = n21908 & ~n21920;
  assign n21922 = ~n21919 & ~n21920;
  assign n21923 = ~n21921 & ~n21922;
  assign n21924 = ~n21667 & ~n21671;
  assign n21925 = n21923 & n21924;
  assign n21926 = ~n21923 & ~n21924;
  assign n21927 = ~n21925 & ~n21926;
  assign n21928 = n4454 & n10394;
  assign n21929 = pi96  & n10744;
  assign n21930 = pi98  & n10392;
  assign n21931 = pi97  & n10387;
  assign n21932 = ~n21930 & ~n21931;
  assign n21933 = ~n21929 & n21932;
  assign n21934 = ~n21928 & n21933;
  assign n21935 = pi56  & ~n21934;
  assign n21936 = pi56  & ~n21935;
  assign n21937 = ~n21934 & ~n21935;
  assign n21938 = ~n21936 & ~n21937;
  assign n21939 = n21927 & ~n21938;
  assign n21940 = n21927 & ~n21939;
  assign n21941 = ~n21938 & ~n21939;
  assign n21942 = ~n21940 & ~n21941;
  assign n21943 = ~n21685 & ~n21688;
  assign n21944 = n21942 & n21943;
  assign n21945 = ~n21942 & ~n21943;
  assign n21946 = ~n21944 & ~n21945;
  assign n21947 = n5169 & n9310;
  assign n21948 = pi99  & n9701;
  assign n21949 = pi101  & n9308;
  assign n21950 = pi100  & n9303;
  assign n21951 = ~n21949 & ~n21950;
  assign n21952 = ~n21948 & n21951;
  assign n21953 = ~n21947 & n21952;
  assign n21954 = pi53  & ~n21953;
  assign n21955 = pi53  & ~n21954;
  assign n21956 = ~n21953 & ~n21954;
  assign n21957 = ~n21955 & ~n21956;
  assign n21958 = ~n21946 & n21957;
  assign n21959 = n21946 & ~n21957;
  assign n21960 = ~n21958 & ~n21959;
  assign n21961 = ~n21882 & n21960;
  assign n21962 = ~n21882 & ~n21961;
  assign n21963 = n21960 & ~n21961;
  assign n21964 = ~n21962 & ~n21963;
  assign n21965 = ~n21881 & ~n21964;
  assign n21966 = n21881 & n21964;
  assign n21967 = ~n21965 & ~n21966;
  assign n21968 = ~n21870 & n21967;
  assign n21969 = n21870 & ~n21967;
  assign n21970 = ~n21968 & ~n21969;
  assign n21971 = n6775 & n7408;
  assign n21972 = pi105  & n7740;
  assign n21973 = pi107  & n7406;
  assign n21974 = pi106  & n7401;
  assign n21975 = ~n21973 & ~n21974;
  assign n21976 = ~n21972 & n21975;
  assign n21977 = ~n21971 & n21976;
  assign n21978 = pi47  & ~n21977;
  assign n21979 = pi47  & ~n21978;
  assign n21980 = ~n21977 & ~n21978;
  assign n21981 = ~n21979 & ~n21980;
  assign n21982 = n21970 & ~n21981;
  assign n21983 = n21970 & ~n21982;
  assign n21984 = ~n21981 & ~n21982;
  assign n21985 = ~n21983 & ~n21984;
  assign n21986 = ~n21626 & ~n21743;
  assign n21987 = ~n21740 & ~n21986;
  assign n21988 = n21985 & n21987;
  assign n21989 = ~n21985 & ~n21987;
  assign n21990 = ~n21988 & ~n21989;
  assign n21991 = n6539 & n7665;
  assign n21992 = pi108  & n6873;
  assign n21993 = pi110  & n6537;
  assign n21994 = pi109  & n6532;
  assign n21995 = ~n21993 & ~n21994;
  assign n21996 = ~n21992 & n21995;
  assign n21997 = ~n21991 & n21996;
  assign n21998 = pi44  & ~n21997;
  assign n21999 = pi44  & ~n21998;
  assign n22000 = ~n21997 & ~n21998;
  assign n22001 = ~n21999 & ~n22000;
  assign n22002 = n21990 & ~n22001;
  assign n22003 = n21990 & ~n22002;
  assign n22004 = ~n22001 & ~n22002;
  assign n22005 = ~n22003 & ~n22004;
  assign n22006 = ~n21758 & ~n21762;
  assign n22007 = n22005 & n22006;
  assign n22008 = ~n22005 & ~n22006;
  assign n22009 = ~n22007 & ~n22008;
  assign n22010 = n5739 & n8612;
  assign n22011 = pi111  & n6030;
  assign n22012 = pi113  & n5737;
  assign n22013 = pi112  & n5732;
  assign n22014 = ~n22012 & ~n22013;
  assign n22015 = ~n22011 & n22014;
  assign n22016 = ~n22010 & n22015;
  assign n22017 = pi41  & ~n22016;
  assign n22018 = pi41  & ~n22017;
  assign n22019 = ~n22016 & ~n22017;
  assign n22020 = ~n22018 & ~n22019;
  assign n22021 = n22009 & ~n22020;
  assign n22022 = n22009 & ~n22021;
  assign n22023 = ~n22020 & ~n22021;
  assign n22024 = ~n22022 & ~n22023;
  assign n22025 = ~n21775 & ~n21781;
  assign n22026 = n22024 & n22025;
  assign n22027 = ~n22024 & ~n22025;
  assign n22028 = ~n22026 & ~n22027;
  assign n22029 = n5008 & n9614;
  assign n22030 = pi114  & n5241;
  assign n22031 = pi116  & n5006;
  assign n22032 = pi115  & n5001;
  assign n22033 = ~n22031 & ~n22032;
  assign n22034 = ~n22030 & n22033;
  assign n22035 = ~n22029 & n22034;
  assign n22036 = pi38  & ~n22035;
  assign n22037 = pi38  & ~n22036;
  assign n22038 = ~n22035 & ~n22036;
  assign n22039 = ~n22037 & ~n22038;
  assign n22040 = n22028 & ~n22039;
  assign n22041 = n22028 & ~n22040;
  assign n22042 = ~n22039 & ~n22040;
  assign n22043 = ~n22041 & ~n22042;
  assign n22044 = ~n21799 & n22043;
  assign n22045 = n21799 & ~n22043;
  assign n22046 = ~n22044 & ~n22045;
  assign n22047 = n4271 & n10667;
  assign n22048 = pi117  & n4503;
  assign n22049 = pi119  & n4269;
  assign n22050 = pi118  & n4264;
  assign n22051 = ~n22049 & ~n22050;
  assign n22052 = ~n22048 & n22051;
  assign n22053 = ~n22047 & n22052;
  assign n22054 = pi35  & ~n22053;
  assign n22055 = pi35  & ~n22054;
  assign n22056 = ~n22053 & ~n22054;
  assign n22057 = ~n22055 & ~n22056;
  assign n22058 = ~n22046 & ~n22057;
  assign n22059 = n22046 & n22057;
  assign n22060 = ~n22058 & ~n22059;
  assign n22061 = n21869 & n22060;
  assign n22062 = ~n21869 & ~n22060;
  assign n22063 = ~n22061 & ~n22062;
  assign n22064 = ~n21854 & n22063;
  assign n22065 = ~n21854 & ~n22064;
  assign n22066 = n22063 & ~n22064;
  assign n22067 = ~n22065 & ~n22066;
  assign n22068 = ~n21592 & ~n21603;
  assign n22069 = ~n21822 & ~n22068;
  assign n22070 = pi126  & n2667;
  assign n22071 = pi127  & n2516;
  assign n22072 = ~n22070 & ~n22071;
  assign n22073 = ~n2523 & n22072;
  assign n22074 = n13773 & n22072;
  assign n22075 = ~n22073 & ~n22074;
  assign n22076 = pi26  & ~n22075;
  assign n22077 = ~pi26  & n22075;
  assign n22078 = ~n22076 & ~n22077;
  assign n22079 = ~n22069 & ~n22078;
  assign n22080 = ~n22069 & ~n22079;
  assign n22081 = ~n22078 & ~n22079;
  assign n22082 = ~n22080 & ~n22081;
  assign n22083 = ~n22067 & ~n22082;
  assign n22084 = n22067 & n22082;
  assign n22085 = ~n22083 & ~n22084;
  assign n22086 = ~n21838 & n22085;
  assign n22087 = ~n21838 & ~n22086;
  assign n22088 = n22085 & ~n22086;
  assign n22089 = ~n22087 & ~n22088;
  assign n22090 = ~n21836 & ~n22089;
  assign n22091 = n21836 & n22089;
  assign po88  = ~n22090 & ~n22091;
  assign n22093 = ~n22086 & ~n22090;
  assign n22094 = ~n22079 & ~n22083;
  assign n22095 = ~n21851 & ~n22064;
  assign n22096 = pi127  & n2667;
  assign n22097 = n2523 & n13770;
  assign n22098 = ~n22096 & ~n22097;
  assign n22099 = pi26  & ~n22098;
  assign n22100 = pi26  & ~n22099;
  assign n22101 = ~n22098 & ~n22099;
  assign n22102 = ~n22100 & ~n22101;
  assign n22103 = ~n22095 & ~n22102;
  assign n22104 = ~n22095 & ~n22103;
  assign n22105 = ~n22102 & ~n22103;
  assign n22106 = ~n22104 & ~n22105;
  assign n22107 = n3034 & n13344;
  assign n22108 = pi124  & n3225;
  assign n22109 = pi126  & n3032;
  assign n22110 = pi125  & n3027;
  assign n22111 = ~n22109 & ~n22110;
  assign n22112 = ~n22108 & n22111;
  assign n22113 = ~n22107 & n22112;
  assign n22114 = pi29  & ~n22113;
  assign n22115 = pi29  & ~n22114;
  assign n22116 = ~n22113 & ~n22114;
  assign n22117 = ~n22115 & ~n22116;
  assign n22118 = ~n21867 & ~n22061;
  assign n22119 = n22117 & n22118;
  assign n22120 = ~n22117 & ~n22118;
  assign n22121 = ~n22119 & ~n22120;
  assign n22122 = n3622 & n12158;
  assign n22123 = pi121  & n3814;
  assign n22124 = pi123  & n3620;
  assign n22125 = pi122  & n3615;
  assign n22126 = ~n22124 & ~n22125;
  assign n22127 = ~n22123 & n22126;
  assign n22128 = ~n22122 & n22127;
  assign n22129 = pi32  & ~n22128;
  assign n22130 = pi32  & ~n22129;
  assign n22131 = ~n22128 & ~n22129;
  assign n22132 = ~n22130 & ~n22131;
  assign n22133 = ~n21799 & ~n22043;
  assign n22134 = ~n22058 & ~n22133;
  assign n22135 = n22132 & n22134;
  assign n22136 = ~n22132 & ~n22134;
  assign n22137 = ~n22135 & ~n22136;
  assign n22138 = n4271 & n11028;
  assign n22139 = pi118  & n4503;
  assign n22140 = pi120  & n4269;
  assign n22141 = pi119  & n4264;
  assign n22142 = ~n22140 & ~n22141;
  assign n22143 = ~n22139 & n22142;
  assign n22144 = ~n22138 & n22143;
  assign n22145 = pi35  & ~n22144;
  assign n22146 = pi35  & ~n22145;
  assign n22147 = ~n22144 & ~n22145;
  assign n22148 = ~n22146 & ~n22147;
  assign n22149 = ~n22027 & ~n22040;
  assign n22150 = n5008 & n9958;
  assign n22151 = pi115  & n5241;
  assign n22152 = pi117  & n5006;
  assign n22153 = pi116  & n5001;
  assign n22154 = ~n22152 & ~n22153;
  assign n22155 = ~n22151 & n22154;
  assign n22156 = ~n22150 & n22155;
  assign n22157 = pi38  & ~n22156;
  assign n22158 = pi38  & ~n22157;
  assign n22159 = ~n22156 & ~n22157;
  assign n22160 = ~n22158 & ~n22159;
  assign n22161 = ~n22008 & ~n22021;
  assign n22162 = ~n21968 & ~n21982;
  assign n22163 = n7060 & n7408;
  assign n22164 = pi106  & n7740;
  assign n22165 = pi108  & n7406;
  assign n22166 = pi107  & n7401;
  assign n22167 = ~n22165 & ~n22166;
  assign n22168 = ~n22164 & n22167;
  assign n22169 = ~n22163 & n22168;
  assign n22170 = pi47  & ~n22169;
  assign n22171 = pi47  & ~n22170;
  assign n22172 = ~n22169 & ~n22170;
  assign n22173 = ~n22171 & ~n22172;
  assign n22174 = ~n21961 & ~n21965;
  assign n22175 = ~n21926 & ~n21939;
  assign n22176 = n4684 & n10394;
  assign n22177 = pi97  & n10744;
  assign n22178 = pi99  & n10392;
  assign n22179 = pi98  & n10387;
  assign n22180 = ~n22178 & ~n22179;
  assign n22181 = ~n22177 & n22180;
  assign n22182 = ~n22176 & n22181;
  assign n22183 = pi56  & ~n22182;
  assign n22184 = pi56  & ~n22183;
  assign n22185 = ~n22182 & ~n22183;
  assign n22186 = ~n22184 & ~n22185;
  assign n22187 = ~n21906 & ~n21920;
  assign n22188 = n4001 & n11488;
  assign n22189 = pi94  & n11847;
  assign n22190 = pi96  & n11486;
  assign n22191 = pi95  & n11481;
  assign n22192 = ~n22190 & ~n22191;
  assign n22193 = ~n22189 & n22192;
  assign n22194 = ~n22188 & n22193;
  assign n22195 = pi59  & ~n22194;
  assign n22196 = pi59  & ~n22195;
  assign n22197 = ~n22194 & ~n22195;
  assign n22198 = ~n22196 & ~n22197;
  assign n22199 = ~n21890 & ~n21903;
  assign n22200 = pi89  & n13835;
  assign n22201 = pi90  & ~n13434;
  assign n22202 = ~n22200 & ~n22201;
  assign n22203 = ~n21887 & n22202;
  assign n22204 = n21887 & ~n22202;
  assign n22205 = ~n22203 & ~n22204;
  assign n22206 = pi91  & n13004;
  assign n22207 = pi93  & n12625;
  assign n22208 = pi92  & n12620;
  assign n22209 = ~n22207 & ~n22208;
  assign n22210 = ~n22206 & n22209;
  assign n22211 = ~n12627 & n22210;
  assign n22212 = ~n3371 & n22210;
  assign n22213 = ~n22211 & ~n22212;
  assign n22214 = pi62  & ~n22213;
  assign n22215 = ~pi62  & n22213;
  assign n22216 = ~n22214 & ~n22215;
  assign n22217 = n22205 & ~n22216;
  assign n22218 = ~n22205 & n22216;
  assign n22219 = ~n22217 & ~n22218;
  assign n22220 = ~n22199 & n22219;
  assign n22221 = n22199 & ~n22219;
  assign n22222 = ~n22220 & ~n22221;
  assign n22223 = ~n22198 & n22222;
  assign n22224 = n22198 & ~n22222;
  assign n22225 = ~n22223 & ~n22224;
  assign n22226 = ~n22187 & n22225;
  assign n22227 = n22187 & ~n22225;
  assign n22228 = ~n22226 & ~n22227;
  assign n22229 = ~n22186 & n22228;
  assign n22230 = n22186 & ~n22228;
  assign n22231 = ~n22229 & ~n22230;
  assign n22232 = ~n22175 & n22231;
  assign n22233 = n22175 & ~n22231;
  assign n22234 = ~n22232 & ~n22233;
  assign n22235 = n5413 & n9310;
  assign n22236 = pi100  & n9701;
  assign n22237 = pi102  & n9308;
  assign n22238 = pi101  & n9303;
  assign n22239 = ~n22237 & ~n22238;
  assign n22240 = ~n22236 & n22239;
  assign n22241 = ~n22235 & n22240;
  assign n22242 = pi53  & ~n22241;
  assign n22243 = pi53  & ~n22242;
  assign n22244 = ~n22241 & ~n22242;
  assign n22245 = ~n22243 & ~n22244;
  assign n22246 = n22234 & ~n22245;
  assign n22247 = n22234 & ~n22246;
  assign n22248 = ~n22245 & ~n22246;
  assign n22249 = ~n22247 & ~n22248;
  assign n22250 = ~n21945 & ~n21959;
  assign n22251 = ~n22249 & ~n22250;
  assign n22252 = ~n22249 & ~n22251;
  assign n22253 = ~n22250 & ~n22251;
  assign n22254 = ~n22252 & ~n22253;
  assign n22255 = n6207 & n8334;
  assign n22256 = pi103  & n8685;
  assign n22257 = pi105  & n8332;
  assign n22258 = pi104  & n8327;
  assign n22259 = ~n22257 & ~n22258;
  assign n22260 = ~n22256 & n22259;
  assign n22261 = ~n22255 & n22260;
  assign n22262 = pi50  & ~n22261;
  assign n22263 = pi50  & ~n22262;
  assign n22264 = ~n22261 & ~n22262;
  assign n22265 = ~n22263 & ~n22264;
  assign n22266 = ~n22254 & n22265;
  assign n22267 = n22254 & ~n22265;
  assign n22268 = ~n22266 & ~n22267;
  assign n22269 = ~n22174 & ~n22268;
  assign n22270 = n22174 & n22268;
  assign n22271 = ~n22269 & ~n22270;
  assign n22272 = ~n22173 & n22271;
  assign n22273 = n22173 & ~n22271;
  assign n22274 = ~n22272 & ~n22273;
  assign n22275 = ~n22162 & n22274;
  assign n22276 = n22162 & ~n22274;
  assign n22277 = ~n22275 & ~n22276;
  assign n22278 = n6539 & n7970;
  assign n22279 = pi109  & n6873;
  assign n22280 = pi111  & n6537;
  assign n22281 = pi110  & n6532;
  assign n22282 = ~n22280 & ~n22281;
  assign n22283 = ~n22279 & n22282;
  assign n22284 = ~n22278 & n22283;
  assign n22285 = pi44  & ~n22284;
  assign n22286 = pi44  & ~n22285;
  assign n22287 = ~n22284 & ~n22285;
  assign n22288 = ~n22286 & ~n22287;
  assign n22289 = n22277 & ~n22288;
  assign n22290 = n22277 & ~n22289;
  assign n22291 = ~n22288 & ~n22289;
  assign n22292 = ~n22290 & ~n22291;
  assign n22293 = ~n21989 & ~n22002;
  assign n22294 = n22292 & n22293;
  assign n22295 = ~n22292 & ~n22293;
  assign n22296 = ~n22294 & ~n22295;
  assign n22297 = n5739 & n8936;
  assign n22298 = pi112  & n6030;
  assign n22299 = pi114  & n5737;
  assign n22300 = pi113  & n5732;
  assign n22301 = ~n22299 & ~n22300;
  assign n22302 = ~n22298 & n22301;
  assign n22303 = ~n22297 & n22302;
  assign n22304 = pi41  & ~n22303;
  assign n22305 = pi41  & ~n22304;
  assign n22306 = ~n22303 & ~n22304;
  assign n22307 = ~n22305 & ~n22306;
  assign n22308 = ~n22296 & n22307;
  assign n22309 = n22296 & ~n22307;
  assign n22310 = ~n22308 & ~n22309;
  assign n22311 = ~n22161 & n22310;
  assign n22312 = ~n22161 & ~n22311;
  assign n22313 = n22310 & ~n22311;
  assign n22314 = ~n22312 & ~n22313;
  assign n22315 = ~n22160 & ~n22314;
  assign n22316 = n22160 & n22314;
  assign n22317 = ~n22315 & ~n22316;
  assign n22318 = ~n22149 & n22317;
  assign n22319 = n22149 & ~n22317;
  assign n22320 = ~n22318 & ~n22319;
  assign n22321 = ~n22148 & n22320;
  assign n22322 = ~n22148 & ~n22321;
  assign n22323 = n22320 & ~n22321;
  assign n22324 = ~n22322 & ~n22323;
  assign n22325 = n22137 & ~n22324;
  assign n22326 = n22137 & ~n22325;
  assign n22327 = ~n22324 & ~n22325;
  assign n22328 = ~n22326 & ~n22327;
  assign n22329 = ~n22121 & n22328;
  assign n22330 = n22121 & ~n22328;
  assign n22331 = ~n22329 & ~n22330;
  assign n22332 = ~n22106 & n22331;
  assign n22333 = n22106 & ~n22331;
  assign n22334 = ~n22332 & ~n22333;
  assign n22335 = ~n22094 & n22334;
  assign n22336 = n22094 & ~n22334;
  assign n22337 = ~n22335 & ~n22336;
  assign n22338 = ~n22093 & n22337;
  assign n22339 = n22093 & ~n22337;
  assign po89  = ~n22338 & ~n22339;
  assign n22341 = ~n22103 & ~n22332;
  assign n22342 = ~n22120 & ~n22330;
  assign n22343 = n3034 & n13742;
  assign n22344 = pi125  & n3225;
  assign n22345 = pi127  & n3032;
  assign n22346 = pi126  & n3027;
  assign n22347 = ~n22345 & ~n22346;
  assign n22348 = ~n22344 & n22347;
  assign n22349 = ~n22343 & n22348;
  assign n22350 = pi29  & ~n22349;
  assign n22351 = pi29  & ~n22350;
  assign n22352 = ~n22349 & ~n22350;
  assign n22353 = ~n22351 & ~n22352;
  assign n22354 = ~n22342 & ~n22353;
  assign n22355 = ~n22342 & ~n22354;
  assign n22356 = ~n22353 & ~n22354;
  assign n22357 = ~n22355 & ~n22356;
  assign n22358 = ~n22311 & ~n22315;
  assign n22359 = ~n22295 & ~n22309;
  assign n22360 = ~n22269 & ~n22272;
  assign n22361 = ~n22254 & ~n22265;
  assign n22362 = ~n22251 & ~n22361;
  assign n22363 = n4211 & n11488;
  assign n22364 = pi95  & n11847;
  assign n22365 = pi97  & n11486;
  assign n22366 = pi96  & n11481;
  assign n22367 = ~n22365 & ~n22366;
  assign n22368 = ~n22364 & n22367;
  assign n22369 = ~n22363 & n22368;
  assign n22370 = pi59  & ~n22369;
  assign n22371 = pi59  & ~n22370;
  assign n22372 = ~n22369 & ~n22370;
  assign n22373 = ~n22371 & ~n22372;
  assign n22374 = ~n22220 & ~n22223;
  assign n22375 = n22373 & n22374;
  assign n22376 = ~n22373 & ~n22374;
  assign n22377 = ~n22375 & ~n22376;
  assign n22378 = ~n22203 & ~n22217;
  assign n22379 = pi90  & n13835;
  assign n22380 = pi91  & ~n13434;
  assign n22381 = ~n22379 & ~n22380;
  assign n22382 = ~pi26  & ~n22381;
  assign n22383 = pi26  & n22381;
  assign n22384 = ~n22382 & ~n22383;
  assign n22385 = ~n22202 & n22384;
  assign n22386 = n22202 & ~n22384;
  assign n22387 = ~n22385 & ~n22386;
  assign n22388 = ~n22378 & n22387;
  assign n22389 = n22378 & ~n22387;
  assign n22390 = ~n22388 & ~n22389;
  assign n22391 = n3565 & n12627;
  assign n22392 = pi92  & n13004;
  assign n22393 = pi94  & n12625;
  assign n22394 = pi93  & n12620;
  assign n22395 = ~n22393 & ~n22394;
  assign n22396 = ~n22392 & n22395;
  assign n22397 = ~n22391 & n22396;
  assign n22398 = pi62  & ~n22397;
  assign n22399 = pi62  & ~n22398;
  assign n22400 = ~n22397 & ~n22398;
  assign n22401 = ~n22399 & ~n22400;
  assign n22402 = n22390 & ~n22401;
  assign n22403 = n22390 & ~n22402;
  assign n22404 = ~n22401 & ~n22402;
  assign n22405 = ~n22403 & ~n22404;
  assign n22406 = ~n22377 & n22405;
  assign n22407 = n22377 & ~n22405;
  assign n22408 = ~n22406 & ~n22407;
  assign n22409 = n4910 & n10394;
  assign n22410 = pi98  & n10744;
  assign n22411 = pi100  & n10392;
  assign n22412 = pi99  & n10387;
  assign n22413 = ~n22411 & ~n22412;
  assign n22414 = ~n22410 & n22413;
  assign n22415 = ~n22409 & n22414;
  assign n22416 = pi56  & ~n22415;
  assign n22417 = pi56  & ~n22416;
  assign n22418 = ~n22415 & ~n22416;
  assign n22419 = ~n22417 & ~n22418;
  assign n22420 = n22408 & ~n22419;
  assign n22421 = n22408 & ~n22420;
  assign n22422 = ~n22419 & ~n22420;
  assign n22423 = ~n22421 & ~n22422;
  assign n22424 = ~n22226 & ~n22229;
  assign n22425 = n22423 & n22424;
  assign n22426 = ~n22423 & ~n22424;
  assign n22427 = ~n22425 & ~n22426;
  assign n22428 = n5664 & n9310;
  assign n22429 = pi101  & n9701;
  assign n22430 = pi103  & n9308;
  assign n22431 = pi102  & n9303;
  assign n22432 = ~n22430 & ~n22431;
  assign n22433 = ~n22429 & n22432;
  assign n22434 = ~n22428 & n22433;
  assign n22435 = pi53  & ~n22434;
  assign n22436 = pi53  & ~n22435;
  assign n22437 = ~n22434 & ~n22435;
  assign n22438 = ~n22436 & ~n22437;
  assign n22439 = n22427 & ~n22438;
  assign n22440 = n22427 & ~n22439;
  assign n22441 = ~n22438 & ~n22439;
  assign n22442 = ~n22440 & ~n22441;
  assign n22443 = ~n22232 & ~n22246;
  assign n22444 = n22442 & n22443;
  assign n22445 = ~n22442 & ~n22443;
  assign n22446 = ~n22444 & ~n22445;
  assign n22447 = n6477 & n8334;
  assign n22448 = pi104  & n8685;
  assign n22449 = pi106  & n8332;
  assign n22450 = pi105  & n8327;
  assign n22451 = ~n22449 & ~n22450;
  assign n22452 = ~n22448 & n22451;
  assign n22453 = ~n22447 & n22452;
  assign n22454 = pi50  & ~n22453;
  assign n22455 = pi50  & ~n22454;
  assign n22456 = ~n22453 & ~n22454;
  assign n22457 = ~n22455 & ~n22456;
  assign n22458 = n22446 & ~n22457;
  assign n22459 = n22446 & ~n22458;
  assign n22460 = ~n22457 & ~n22458;
  assign n22461 = ~n22459 & ~n22460;
  assign n22462 = ~n22362 & n22461;
  assign n22463 = n22362 & ~n22461;
  assign n22464 = ~n22462 & ~n22463;
  assign n22465 = n7349 & n7408;
  assign n22466 = pi107  & n7740;
  assign n22467 = pi109  & n7406;
  assign n22468 = pi108  & n7401;
  assign n22469 = ~n22467 & ~n22468;
  assign n22470 = ~n22466 & n22469;
  assign n22471 = ~n22465 & n22470;
  assign n22472 = pi47  & ~n22471;
  assign n22473 = pi47  & ~n22472;
  assign n22474 = ~n22471 & ~n22472;
  assign n22475 = ~n22473 & ~n22474;
  assign n22476 = ~n22464 & ~n22475;
  assign n22477 = n22464 & n22475;
  assign n22478 = ~n22476 & ~n22477;
  assign n22479 = n22360 & ~n22478;
  assign n22480 = ~n22360 & n22478;
  assign n22481 = ~n22479 & ~n22480;
  assign n22482 = n6539 & n7997;
  assign n22483 = pi110  & n6873;
  assign n22484 = pi112  & n6537;
  assign n22485 = pi111  & n6532;
  assign n22486 = ~n22484 & ~n22485;
  assign n22487 = ~n22483 & n22486;
  assign n22488 = ~n22482 & n22487;
  assign n22489 = pi44  & ~n22488;
  assign n22490 = pi44  & ~n22489;
  assign n22491 = ~n22488 & ~n22489;
  assign n22492 = ~n22490 & ~n22491;
  assign n22493 = n22481 & ~n22492;
  assign n22494 = n22481 & ~n22493;
  assign n22495 = ~n22492 & ~n22493;
  assign n22496 = ~n22494 & ~n22495;
  assign n22497 = ~n22275 & ~n22289;
  assign n22498 = n22496 & n22497;
  assign n22499 = ~n22496 & ~n22497;
  assign n22500 = ~n22498 & ~n22499;
  assign n22501 = n5739 & n8963;
  assign n22502 = pi113  & n6030;
  assign n22503 = pi115  & n5737;
  assign n22504 = pi114  & n5732;
  assign n22505 = ~n22503 & ~n22504;
  assign n22506 = ~n22502 & n22505;
  assign n22507 = ~n22501 & n22506;
  assign n22508 = pi41  & ~n22507;
  assign n22509 = pi41  & ~n22508;
  assign n22510 = ~n22507 & ~n22508;
  assign n22511 = ~n22509 & ~n22510;
  assign n22512 = ~n22500 & n22511;
  assign n22513 = n22500 & ~n22511;
  assign n22514 = ~n22359 & ~n22512;
  assign n22515 = ~n22513 & n22514;
  assign n22516 = ~n22359 & ~n22515;
  assign n22517 = ~n22513 & ~n22515;
  assign n22518 = ~n22512 & n22517;
  assign n22519 = ~n22516 & ~n22518;
  assign n22520 = n5008 & n9984;
  assign n22521 = pi116  & n5241;
  assign n22522 = pi118  & n5006;
  assign n22523 = pi117  & n5001;
  assign n22524 = ~n22522 & ~n22523;
  assign n22525 = ~n22521 & n22524;
  assign n22526 = ~n22520 & n22525;
  assign n22527 = pi38  & ~n22526;
  assign n22528 = pi38  & ~n22527;
  assign n22529 = ~n22526 & ~n22527;
  assign n22530 = ~n22528 & ~n22529;
  assign n22531 = n22519 & n22530;
  assign n22532 = ~n22519 & ~n22530;
  assign n22533 = ~n22531 & ~n22532;
  assign n22534 = ~n22358 & n22533;
  assign n22535 = n22358 & ~n22533;
  assign n22536 = ~n22534 & ~n22535;
  assign n22537 = n4271 & n11389;
  assign n22538 = pi119  & n4503;
  assign n22539 = pi121  & n4269;
  assign n22540 = pi120  & n4264;
  assign n22541 = ~n22539 & ~n22540;
  assign n22542 = ~n22538 & n22541;
  assign n22543 = ~n22537 & n22542;
  assign n22544 = pi35  & ~n22543;
  assign n22545 = pi35  & ~n22544;
  assign n22546 = ~n22543 & ~n22544;
  assign n22547 = ~n22545 & ~n22546;
  assign n22548 = n22536 & ~n22547;
  assign n22549 = n22536 & ~n22548;
  assign n22550 = ~n22547 & ~n22548;
  assign n22551 = ~n22549 & ~n22550;
  assign n22552 = ~n22318 & ~n22321;
  assign n22553 = n22551 & n22552;
  assign n22554 = ~n22551 & ~n22552;
  assign n22555 = ~n22553 & ~n22554;
  assign n22556 = n3622 & n12189;
  assign n22557 = pi122  & n3814;
  assign n22558 = pi124  & n3620;
  assign n22559 = pi123  & n3615;
  assign n22560 = ~n22558 & ~n22559;
  assign n22561 = ~n22557 & n22560;
  assign n22562 = ~n22556 & n22561;
  assign n22563 = pi32  & ~n22562;
  assign n22564 = pi32  & ~n22563;
  assign n22565 = ~n22562 & ~n22563;
  assign n22566 = ~n22564 & ~n22565;
  assign n22567 = ~n22136 & ~n22325;
  assign n22568 = n22566 & n22567;
  assign n22569 = ~n22566 & ~n22567;
  assign n22570 = ~n22568 & ~n22569;
  assign n22571 = n22555 & ~n22570;
  assign n22572 = ~n22555 & n22570;
  assign n22573 = ~n22571 & ~n22572;
  assign n22574 = ~n22357 & ~n22573;
  assign n22575 = n22357 & n22573;
  assign n22576 = ~n22574 & ~n22575;
  assign n22577 = n22341 & ~n22576;
  assign n22578 = ~n22341 & n22576;
  assign n22579 = ~n22577 & ~n22578;
  assign n22580 = ~n22335 & ~n22338;
  assign n22581 = n22579 & ~n22580;
  assign n22582 = ~n22579 & n22580;
  assign po90  = ~n22581 & ~n22582;
  assign n22584 = pi126  & n3225;
  assign n22585 = pi127  & n3027;
  assign n22586 = ~n22584 & ~n22585;
  assign n22587 = ~n3034 & n22586;
  assign n22588 = n13773 & n22586;
  assign n22589 = ~n22587 & ~n22588;
  assign n22590 = pi29  & ~n22589;
  assign n22591 = ~pi29  & n22589;
  assign n22592 = ~n22590 & ~n22591;
  assign n22593 = ~n22568 & ~n22572;
  assign n22594 = ~n22592 & n22593;
  assign n22595 = n22592 & ~n22593;
  assign n22596 = ~n22594 & ~n22595;
  assign n22597 = n3622 & n12943;
  assign n22598 = pi123  & n3814;
  assign n22599 = pi125  & n3620;
  assign n22600 = pi124  & n3615;
  assign n22601 = ~n22599 & ~n22600;
  assign n22602 = ~n22598 & n22601;
  assign n22603 = ~n22597 & n22602;
  assign n22604 = pi32  & ~n22603;
  assign n22605 = pi32  & ~n22604;
  assign n22606 = ~n22603 & ~n22604;
  assign n22607 = ~n22605 & ~n22606;
  assign n22608 = ~n22548 & ~n22554;
  assign n22609 = n22607 & n22608;
  assign n22610 = ~n22607 & ~n22608;
  assign n22611 = ~n22609 & ~n22610;
  assign n22612 = ~n22532 & ~n22534;
  assign n22613 = ~n22439 & ~n22445;
  assign n22614 = n5943 & n9310;
  assign n22615 = pi102  & n9701;
  assign n22616 = pi104  & n9308;
  assign n22617 = pi103  & n9303;
  assign n22618 = ~n22616 & ~n22617;
  assign n22619 = ~n22615 & n22618;
  assign n22620 = ~n22614 & n22619;
  assign n22621 = pi53  & ~n22620;
  assign n22622 = pi53  & ~n22621;
  assign n22623 = ~n22620 & ~n22621;
  assign n22624 = ~n22622 & ~n22623;
  assign n22625 = ~n22420 & ~n22426;
  assign n22626 = pi91  & n13835;
  assign n22627 = pi92  & ~n13434;
  assign n22628 = ~n22626 & ~n22627;
  assign n22629 = ~n22382 & ~n22385;
  assign n22630 = ~n22628 & n22629;
  assign n22631 = n22628 & ~n22629;
  assign n22632 = ~n22630 & ~n22631;
  assign n22633 = n3784 & n12627;
  assign n22634 = pi93  & n13004;
  assign n22635 = pi95  & n12625;
  assign n22636 = pi94  & n12620;
  assign n22637 = ~n22635 & ~n22636;
  assign n22638 = ~n22634 & n22637;
  assign n22639 = ~n22633 & n22638;
  assign n22640 = pi62  & ~n22639;
  assign n22641 = pi62  & ~n22640;
  assign n22642 = ~n22639 & ~n22640;
  assign n22643 = ~n22641 & ~n22642;
  assign n22644 = ~n22632 & n22643;
  assign n22645 = n22632 & ~n22643;
  assign n22646 = ~n22644 & ~n22645;
  assign n22647 = ~n22388 & ~n22402;
  assign n22648 = n22646 & ~n22647;
  assign n22649 = ~n22646 & n22647;
  assign n22650 = ~n22648 & ~n22649;
  assign n22651 = n4454 & n11488;
  assign n22652 = pi96  & n11847;
  assign n22653 = pi98  & n11486;
  assign n22654 = pi97  & n11481;
  assign n22655 = ~n22653 & ~n22654;
  assign n22656 = ~n22652 & n22655;
  assign n22657 = ~n22651 & n22656;
  assign n22658 = pi59  & ~n22657;
  assign n22659 = pi59  & ~n22658;
  assign n22660 = ~n22657 & ~n22658;
  assign n22661 = ~n22659 & ~n22660;
  assign n22662 = n22650 & ~n22661;
  assign n22663 = n22650 & ~n22662;
  assign n22664 = ~n22661 & ~n22662;
  assign n22665 = ~n22663 & ~n22664;
  assign n22666 = ~n22376 & ~n22407;
  assign n22667 = ~n22665 & ~n22666;
  assign n22668 = ~n22665 & ~n22667;
  assign n22669 = ~n22666 & ~n22667;
  assign n22670 = ~n22668 & ~n22669;
  assign n22671 = n5169 & n10394;
  assign n22672 = pi99  & n10744;
  assign n22673 = pi101  & n10392;
  assign n22674 = pi100  & n10387;
  assign n22675 = ~n22673 & ~n22674;
  assign n22676 = ~n22672 & n22675;
  assign n22677 = ~n22671 & n22676;
  assign n22678 = pi56  & ~n22677;
  assign n22679 = pi56  & ~n22678;
  assign n22680 = ~n22677 & ~n22678;
  assign n22681 = ~n22679 & ~n22680;
  assign n22682 = ~n22670 & n22681;
  assign n22683 = n22670 & ~n22681;
  assign n22684 = ~n22682 & ~n22683;
  assign n22685 = ~n22625 & ~n22684;
  assign n22686 = ~n22625 & ~n22685;
  assign n22687 = ~n22684 & ~n22685;
  assign n22688 = ~n22686 & ~n22687;
  assign n22689 = ~n22624 & ~n22688;
  assign n22690 = n22624 & n22688;
  assign n22691 = ~n22689 & ~n22690;
  assign n22692 = ~n22613 & n22691;
  assign n22693 = n22613 & ~n22691;
  assign n22694 = ~n22692 & ~n22693;
  assign n22695 = n6775 & n8334;
  assign n22696 = pi105  & n8685;
  assign n22697 = pi107  & n8332;
  assign n22698 = pi106  & n8327;
  assign n22699 = ~n22697 & ~n22698;
  assign n22700 = ~n22696 & n22699;
  assign n22701 = ~n22695 & n22700;
  assign n22702 = pi50  & ~n22701;
  assign n22703 = pi50  & ~n22702;
  assign n22704 = ~n22701 & ~n22702;
  assign n22705 = ~n22703 & ~n22704;
  assign n22706 = n22694 & ~n22705;
  assign n22707 = n22694 & ~n22706;
  assign n22708 = ~n22705 & ~n22706;
  assign n22709 = ~n22707 & ~n22708;
  assign n22710 = ~n22362 & ~n22461;
  assign n22711 = ~n22458 & ~n22710;
  assign n22712 = n22709 & n22711;
  assign n22713 = ~n22709 & ~n22711;
  assign n22714 = ~n22712 & ~n22713;
  assign n22715 = n7408 & n7665;
  assign n22716 = pi108  & n7740;
  assign n22717 = pi110  & n7406;
  assign n22718 = pi109  & n7401;
  assign n22719 = ~n22717 & ~n22718;
  assign n22720 = ~n22716 & n22719;
  assign n22721 = ~n22715 & n22720;
  assign n22722 = pi47  & ~n22721;
  assign n22723 = pi47  & ~n22722;
  assign n22724 = ~n22721 & ~n22722;
  assign n22725 = ~n22723 & ~n22724;
  assign n22726 = n22714 & ~n22725;
  assign n22727 = n22714 & ~n22726;
  assign n22728 = ~n22725 & ~n22726;
  assign n22729 = ~n22727 & ~n22728;
  assign n22730 = ~n22476 & ~n22480;
  assign n22731 = n22729 & n22730;
  assign n22732 = ~n22729 & ~n22730;
  assign n22733 = ~n22731 & ~n22732;
  assign n22734 = n6539 & n8612;
  assign n22735 = pi111  & n6873;
  assign n22736 = pi113  & n6537;
  assign n22737 = pi112  & n6532;
  assign n22738 = ~n22736 & ~n22737;
  assign n22739 = ~n22735 & n22738;
  assign n22740 = ~n22734 & n22739;
  assign n22741 = pi44  & ~n22740;
  assign n22742 = pi44  & ~n22741;
  assign n22743 = ~n22740 & ~n22741;
  assign n22744 = ~n22742 & ~n22743;
  assign n22745 = n22733 & ~n22744;
  assign n22746 = n22733 & ~n22745;
  assign n22747 = ~n22744 & ~n22745;
  assign n22748 = ~n22746 & ~n22747;
  assign n22749 = ~n22493 & ~n22499;
  assign n22750 = n22748 & n22749;
  assign n22751 = ~n22748 & ~n22749;
  assign n22752 = ~n22750 & ~n22751;
  assign n22753 = n5739 & n9614;
  assign n22754 = pi114  & n6030;
  assign n22755 = pi116  & n5737;
  assign n22756 = pi115  & n5732;
  assign n22757 = ~n22755 & ~n22756;
  assign n22758 = ~n22754 & n22757;
  assign n22759 = ~n22753 & n22758;
  assign n22760 = pi41  & ~n22759;
  assign n22761 = pi41  & ~n22760;
  assign n22762 = ~n22759 & ~n22760;
  assign n22763 = ~n22761 & ~n22762;
  assign n22764 = n22752 & ~n22763;
  assign n22765 = n22752 & ~n22764;
  assign n22766 = ~n22763 & ~n22764;
  assign n22767 = ~n22765 & ~n22766;
  assign n22768 = ~n22517 & n22767;
  assign n22769 = n22517 & ~n22767;
  assign n22770 = ~n22768 & ~n22769;
  assign n22771 = n5008 & n10667;
  assign n22772 = pi117  & n5241;
  assign n22773 = pi119  & n5006;
  assign n22774 = pi118  & n5001;
  assign n22775 = ~n22773 & ~n22774;
  assign n22776 = ~n22772 & n22775;
  assign n22777 = ~n22771 & n22776;
  assign n22778 = pi38  & ~n22777;
  assign n22779 = pi38  & ~n22778;
  assign n22780 = ~n22777 & ~n22778;
  assign n22781 = ~n22779 & ~n22780;
  assign n22782 = ~n22770 & ~n22781;
  assign n22783 = n22770 & n22781;
  assign n22784 = ~n22782 & ~n22783;
  assign n22785 = ~n22612 & n22784;
  assign n22786 = n22612 & ~n22784;
  assign n22787 = ~n22785 & ~n22786;
  assign n22788 = n4271 & n11778;
  assign n22789 = pi120  & n4503;
  assign n22790 = pi122  & n4269;
  assign n22791 = pi121  & n4264;
  assign n22792 = ~n22790 & ~n22791;
  assign n22793 = ~n22789 & n22792;
  assign n22794 = ~n22788 & n22793;
  assign n22795 = pi35  & ~n22794;
  assign n22796 = pi35  & ~n22795;
  assign n22797 = ~n22794 & ~n22795;
  assign n22798 = ~n22796 & ~n22797;
  assign n22799 = n22787 & ~n22798;
  assign n22800 = n22787 & ~n22799;
  assign n22801 = ~n22798 & ~n22799;
  assign n22802 = ~n22800 & ~n22801;
  assign n22803 = n22611 & ~n22802;
  assign n22804 = ~n22611 & n22802;
  assign n22805 = ~n22803 & ~n22804;
  assign n22806 = n22596 & n22805;
  assign n22807 = n22596 & ~n22806;
  assign n22808 = n22805 & ~n22806;
  assign n22809 = ~n22807 & ~n22808;
  assign n22810 = ~n22354 & ~n22574;
  assign n22811 = n22809 & n22810;
  assign n22812 = ~n22809 & ~n22810;
  assign n22813 = ~n22811 & ~n22812;
  assign n22814 = ~n22578 & ~n22581;
  assign n22815 = n22813 & ~n22814;
  assign n22816 = ~n22813 & n22814;
  assign po91  = ~n22815 & ~n22816;
  assign n22818 = ~n22812 & ~n22815;
  assign n22819 = ~n22594 & ~n22806;
  assign n22820 = ~n22610 & ~n22803;
  assign n22821 = pi127  & n3225;
  assign n22822 = n3034 & n13770;
  assign n22823 = ~n22821 & ~n22822;
  assign n22824 = pi29  & ~n22823;
  assign n22825 = pi29  & ~n22824;
  assign n22826 = ~n22823 & ~n22824;
  assign n22827 = ~n22825 & ~n22826;
  assign n22828 = ~n22820 & ~n22827;
  assign n22829 = ~n22820 & ~n22828;
  assign n22830 = ~n22827 & ~n22828;
  assign n22831 = ~n22829 & ~n22830;
  assign n22832 = n3622 & n13344;
  assign n22833 = pi124  & n3814;
  assign n22834 = pi126  & n3620;
  assign n22835 = pi125  & n3615;
  assign n22836 = ~n22834 & ~n22835;
  assign n22837 = ~n22833 & n22836;
  assign n22838 = ~n22832 & n22837;
  assign n22839 = pi32  & ~n22838;
  assign n22840 = pi32  & ~n22839;
  assign n22841 = ~n22838 & ~n22839;
  assign n22842 = ~n22840 & ~n22841;
  assign n22843 = ~n22785 & ~n22799;
  assign n22844 = n22842 & n22843;
  assign n22845 = ~n22842 & ~n22843;
  assign n22846 = ~n22844 & ~n22845;
  assign n22847 = ~n22517 & ~n22767;
  assign n22848 = ~n22782 & ~n22847;
  assign n22849 = n5008 & n11028;
  assign n22850 = pi118  & n5241;
  assign n22851 = pi120  & n5006;
  assign n22852 = pi119  & n5001;
  assign n22853 = ~n22851 & ~n22852;
  assign n22854 = ~n22850 & n22853;
  assign n22855 = ~n22849 & n22854;
  assign n22856 = pi38  & ~n22855;
  assign n22857 = pi38  & ~n22856;
  assign n22858 = ~n22855 & ~n22856;
  assign n22859 = ~n22857 & ~n22858;
  assign n22860 = ~n22751 & ~n22764;
  assign n22861 = n5739 & n9958;
  assign n22862 = pi115  & n6030;
  assign n22863 = pi117  & n5737;
  assign n22864 = pi116  & n5732;
  assign n22865 = ~n22863 & ~n22864;
  assign n22866 = ~n22862 & n22865;
  assign n22867 = ~n22861 & n22866;
  assign n22868 = pi41  & ~n22867;
  assign n22869 = pi41  & ~n22868;
  assign n22870 = ~n22867 & ~n22868;
  assign n22871 = ~n22869 & ~n22870;
  assign n22872 = ~n22732 & ~n22745;
  assign n22873 = ~n22692 & ~n22706;
  assign n22874 = n7060 & n8334;
  assign n22875 = pi106  & n8685;
  assign n22876 = pi108  & n8332;
  assign n22877 = pi107  & n8327;
  assign n22878 = ~n22876 & ~n22877;
  assign n22879 = ~n22875 & n22878;
  assign n22880 = ~n22874 & n22879;
  assign n22881 = pi50  & ~n22880;
  assign n22882 = pi50  & ~n22881;
  assign n22883 = ~n22880 & ~n22881;
  assign n22884 = ~n22882 & ~n22883;
  assign n22885 = ~n22685 & ~n22689;
  assign n22886 = ~n22648 & ~n22662;
  assign n22887 = n4684 & n11488;
  assign n22888 = pi97  & n11847;
  assign n22889 = pi99  & n11486;
  assign n22890 = pi98  & n11481;
  assign n22891 = ~n22889 & ~n22890;
  assign n22892 = ~n22888 & n22891;
  assign n22893 = ~n22887 & n22892;
  assign n22894 = pi59  & ~n22893;
  assign n22895 = pi59  & ~n22894;
  assign n22896 = ~n22893 & ~n22894;
  assign n22897 = ~n22895 & ~n22896;
  assign n22898 = ~n22631 & ~n22645;
  assign n22899 = pi92  & n13835;
  assign n22900 = pi93  & ~n13434;
  assign n22901 = ~n22899 & ~n22900;
  assign n22902 = n22628 & ~n22901;
  assign n22903 = ~n22628 & n22901;
  assign n22904 = ~n22902 & ~n22903;
  assign n22905 = ~n22898 & n22904;
  assign n22906 = ~n22898 & ~n22905;
  assign n22907 = ~n22903 & ~n22905;
  assign n22908 = ~n22902 & n22907;
  assign n22909 = ~n22906 & ~n22908;
  assign n22910 = n4001 & n12627;
  assign n22911 = pi94  & n13004;
  assign n22912 = pi96  & n12625;
  assign n22913 = pi95  & n12620;
  assign n22914 = ~n22912 & ~n22913;
  assign n22915 = ~n22911 & n22914;
  assign n22916 = ~n22910 & n22915;
  assign n22917 = pi62  & ~n22916;
  assign n22918 = pi62  & ~n22917;
  assign n22919 = ~n22916 & ~n22917;
  assign n22920 = ~n22918 & ~n22919;
  assign n22921 = ~n22909 & n22920;
  assign n22922 = n22909 & ~n22920;
  assign n22923 = ~n22921 & ~n22922;
  assign n22924 = ~n22897 & ~n22923;
  assign n22925 = n22897 & n22923;
  assign n22926 = ~n22924 & ~n22925;
  assign n22927 = ~n22886 & n22926;
  assign n22928 = n22886 & ~n22926;
  assign n22929 = ~n22927 & ~n22928;
  assign n22930 = n5413 & n10394;
  assign n22931 = pi100  & n10744;
  assign n22932 = pi102  & n10392;
  assign n22933 = pi101  & n10387;
  assign n22934 = ~n22932 & ~n22933;
  assign n22935 = ~n22931 & n22934;
  assign n22936 = ~n22930 & n22935;
  assign n22937 = pi56  & ~n22936;
  assign n22938 = pi56  & ~n22937;
  assign n22939 = ~n22936 & ~n22937;
  assign n22940 = ~n22938 & ~n22939;
  assign n22941 = n22929 & ~n22940;
  assign n22942 = n22929 & ~n22941;
  assign n22943 = ~n22940 & ~n22941;
  assign n22944 = ~n22942 & ~n22943;
  assign n22945 = ~n22670 & ~n22681;
  assign n22946 = ~n22667 & ~n22945;
  assign n22947 = ~n22944 & ~n22946;
  assign n22948 = ~n22944 & ~n22947;
  assign n22949 = ~n22946 & ~n22947;
  assign n22950 = ~n22948 & ~n22949;
  assign n22951 = n6207 & n9310;
  assign n22952 = pi103  & n9701;
  assign n22953 = pi105  & n9308;
  assign n22954 = pi104  & n9303;
  assign n22955 = ~n22953 & ~n22954;
  assign n22956 = ~n22952 & n22955;
  assign n22957 = ~n22951 & n22956;
  assign n22958 = pi53  & ~n22957;
  assign n22959 = pi53  & ~n22958;
  assign n22960 = ~n22957 & ~n22958;
  assign n22961 = ~n22959 & ~n22960;
  assign n22962 = ~n22950 & n22961;
  assign n22963 = n22950 & ~n22961;
  assign n22964 = ~n22962 & ~n22963;
  assign n22965 = ~n22885 & ~n22964;
  assign n22966 = n22885 & n22964;
  assign n22967 = ~n22965 & ~n22966;
  assign n22968 = ~n22884 & n22967;
  assign n22969 = n22884 & ~n22967;
  assign n22970 = ~n22968 & ~n22969;
  assign n22971 = ~n22873 & n22970;
  assign n22972 = n22873 & ~n22970;
  assign n22973 = ~n22971 & ~n22972;
  assign n22974 = n7408 & n7970;
  assign n22975 = pi109  & n7740;
  assign n22976 = pi111  & n7406;
  assign n22977 = pi110  & n7401;
  assign n22978 = ~n22976 & ~n22977;
  assign n22979 = ~n22975 & n22978;
  assign n22980 = ~n22974 & n22979;
  assign n22981 = pi47  & ~n22980;
  assign n22982 = pi47  & ~n22981;
  assign n22983 = ~n22980 & ~n22981;
  assign n22984 = ~n22982 & ~n22983;
  assign n22985 = n22973 & ~n22984;
  assign n22986 = n22973 & ~n22985;
  assign n22987 = ~n22984 & ~n22985;
  assign n22988 = ~n22986 & ~n22987;
  assign n22989 = ~n22713 & ~n22726;
  assign n22990 = n22988 & n22989;
  assign n22991 = ~n22988 & ~n22989;
  assign n22992 = ~n22990 & ~n22991;
  assign n22993 = n6539 & n8936;
  assign n22994 = pi112  & n6873;
  assign n22995 = pi114  & n6537;
  assign n22996 = pi113  & n6532;
  assign n22997 = ~n22995 & ~n22996;
  assign n22998 = ~n22994 & n22997;
  assign n22999 = ~n22993 & n22998;
  assign n23000 = pi44  & ~n22999;
  assign n23001 = pi44  & ~n23000;
  assign n23002 = ~n22999 & ~n23000;
  assign n23003 = ~n23001 & ~n23002;
  assign n23004 = ~n22992 & n23003;
  assign n23005 = n22992 & ~n23003;
  assign n23006 = ~n23004 & ~n23005;
  assign n23007 = ~n22872 & n23006;
  assign n23008 = ~n22872 & ~n23007;
  assign n23009 = n23006 & ~n23007;
  assign n23010 = ~n23008 & ~n23009;
  assign n23011 = ~n22871 & ~n23010;
  assign n23012 = n22871 & n23010;
  assign n23013 = ~n23011 & ~n23012;
  assign n23014 = ~n22860 & n23013;
  assign n23015 = n22860 & ~n23013;
  assign n23016 = ~n23014 & ~n23015;
  assign n23017 = ~n22859 & n23016;
  assign n23018 = n22859 & ~n23016;
  assign n23019 = ~n23017 & ~n23018;
  assign n23020 = ~n22848 & n23019;
  assign n23021 = n22848 & ~n23019;
  assign n23022 = ~n23020 & ~n23021;
  assign n23023 = n4271 & n12158;
  assign n23024 = pi121  & n4503;
  assign n23025 = pi123  & n4269;
  assign n23026 = pi122  & n4264;
  assign n23027 = ~n23025 & ~n23026;
  assign n23028 = ~n23024 & n23027;
  assign n23029 = ~n23023 & n23028;
  assign n23030 = pi35  & ~n23029;
  assign n23031 = pi35  & ~n23030;
  assign n23032 = ~n23029 & ~n23030;
  assign n23033 = ~n23031 & ~n23032;
  assign n23034 = n23022 & ~n23033;
  assign n23035 = n23022 & ~n23034;
  assign n23036 = ~n23033 & ~n23034;
  assign n23037 = ~n23035 & ~n23036;
  assign n23038 = ~n22846 & n23037;
  assign n23039 = n22846 & ~n23037;
  assign n23040 = ~n23038 & ~n23039;
  assign n23041 = ~n22831 & n23040;
  assign n23042 = n22831 & ~n23040;
  assign n23043 = ~n23041 & ~n23042;
  assign n23044 = ~n22819 & n23043;
  assign n23045 = ~n22819 & ~n23044;
  assign n23046 = n23043 & ~n23044;
  assign n23047 = ~n23045 & ~n23046;
  assign n23048 = ~n22818 & ~n23047;
  assign n23049 = n22818 & n23047;
  assign po92  = ~n23048 & ~n23049;
  assign n23051 = ~n23044 & ~n23048;
  assign n23052 = ~n22828 & ~n23041;
  assign n23053 = ~n23007 & ~n23011;
  assign n23054 = ~n22991 & ~n23005;
  assign n23055 = ~n22965 & ~n22968;
  assign n23056 = ~n22950 & ~n22961;
  assign n23057 = ~n22947 & ~n23056;
  assign n23058 = ~n22909 & ~n22920;
  assign n23059 = ~n22924 & ~n23058;
  assign n23060 = pi93  & n13835;
  assign n23061 = pi94  & ~n13434;
  assign n23062 = ~n23060 & ~n23061;
  assign n23063 = ~pi29  & ~n23062;
  assign n23064 = pi29  & n23062;
  assign n23065 = ~n23063 & ~n23064;
  assign n23066 = ~n22901 & n23065;
  assign n23067 = ~n22901 & ~n23066;
  assign n23068 = n23065 & ~n23066;
  assign n23069 = ~n23067 & ~n23068;
  assign n23070 = ~n22907 & ~n23069;
  assign n23071 = ~n22907 & ~n23070;
  assign n23072 = ~n23069 & ~n23070;
  assign n23073 = ~n23071 & ~n23072;
  assign n23074 = n4211 & n12627;
  assign n23075 = pi95  & n13004;
  assign n23076 = pi97  & n12625;
  assign n23077 = pi96  & n12620;
  assign n23078 = ~n23076 & ~n23077;
  assign n23079 = ~n23075 & n23078;
  assign n23080 = ~n23074 & n23079;
  assign n23081 = pi62  & ~n23080;
  assign n23082 = pi62  & ~n23081;
  assign n23083 = ~n23080 & ~n23081;
  assign n23084 = ~n23082 & ~n23083;
  assign n23085 = ~n23073 & n23084;
  assign n23086 = n23073 & ~n23084;
  assign n23087 = ~n23085 & ~n23086;
  assign n23088 = n4910 & n11488;
  assign n23089 = pi98  & n11847;
  assign n23090 = pi100  & n11486;
  assign n23091 = pi99  & n11481;
  assign n23092 = ~n23090 & ~n23091;
  assign n23093 = ~n23089 & n23092;
  assign n23094 = ~n23088 & n23093;
  assign n23095 = pi59  & ~n23094;
  assign n23096 = pi59  & ~n23095;
  assign n23097 = ~n23094 & ~n23095;
  assign n23098 = ~n23096 & ~n23097;
  assign n23099 = ~n23087 & ~n23098;
  assign n23100 = n23087 & n23098;
  assign n23101 = ~n23099 & ~n23100;
  assign n23102 = ~n23059 & n23101;
  assign n23103 = n23059 & ~n23101;
  assign n23104 = ~n23102 & ~n23103;
  assign n23105 = n5664 & n10394;
  assign n23106 = pi101  & n10744;
  assign n23107 = pi103  & n10392;
  assign n23108 = pi102  & n10387;
  assign n23109 = ~n23107 & ~n23108;
  assign n23110 = ~n23106 & n23109;
  assign n23111 = ~n23105 & n23110;
  assign n23112 = pi56  & ~n23111;
  assign n23113 = pi56  & ~n23112;
  assign n23114 = ~n23111 & ~n23112;
  assign n23115 = ~n23113 & ~n23114;
  assign n23116 = n23104 & ~n23115;
  assign n23117 = n23104 & ~n23116;
  assign n23118 = ~n23115 & ~n23116;
  assign n23119 = ~n23117 & ~n23118;
  assign n23120 = ~n22927 & ~n22941;
  assign n23121 = n23119 & n23120;
  assign n23122 = ~n23119 & ~n23120;
  assign n23123 = ~n23121 & ~n23122;
  assign n23124 = n6477 & n9310;
  assign n23125 = pi104  & n9701;
  assign n23126 = pi106  & n9308;
  assign n23127 = pi105  & n9303;
  assign n23128 = ~n23126 & ~n23127;
  assign n23129 = ~n23125 & n23128;
  assign n23130 = ~n23124 & n23129;
  assign n23131 = pi53  & ~n23130;
  assign n23132 = pi53  & ~n23131;
  assign n23133 = ~n23130 & ~n23131;
  assign n23134 = ~n23132 & ~n23133;
  assign n23135 = n23123 & ~n23134;
  assign n23136 = n23123 & ~n23135;
  assign n23137 = ~n23134 & ~n23135;
  assign n23138 = ~n23136 & ~n23137;
  assign n23139 = ~n23057 & n23138;
  assign n23140 = n23057 & ~n23138;
  assign n23141 = ~n23139 & ~n23140;
  assign n23142 = n7349 & n8334;
  assign n23143 = pi107  & n8685;
  assign n23144 = pi109  & n8332;
  assign n23145 = pi108  & n8327;
  assign n23146 = ~n23144 & ~n23145;
  assign n23147 = ~n23143 & n23146;
  assign n23148 = ~n23142 & n23147;
  assign n23149 = pi50  & ~n23148;
  assign n23150 = pi50  & ~n23149;
  assign n23151 = ~n23148 & ~n23149;
  assign n23152 = ~n23150 & ~n23151;
  assign n23153 = ~n23141 & ~n23152;
  assign n23154 = n23141 & n23152;
  assign n23155 = ~n23153 & ~n23154;
  assign n23156 = n23055 & ~n23155;
  assign n23157 = ~n23055 & n23155;
  assign n23158 = ~n23156 & ~n23157;
  assign n23159 = n7408 & n7997;
  assign n23160 = pi110  & n7740;
  assign n23161 = pi112  & n7406;
  assign n23162 = pi111  & n7401;
  assign n23163 = ~n23161 & ~n23162;
  assign n23164 = ~n23160 & n23163;
  assign n23165 = ~n23159 & n23164;
  assign n23166 = pi47  & ~n23165;
  assign n23167 = pi47  & ~n23166;
  assign n23168 = ~n23165 & ~n23166;
  assign n23169 = ~n23167 & ~n23168;
  assign n23170 = n23158 & ~n23169;
  assign n23171 = n23158 & ~n23170;
  assign n23172 = ~n23169 & ~n23170;
  assign n23173 = ~n23171 & ~n23172;
  assign n23174 = ~n22971 & ~n22985;
  assign n23175 = n23173 & n23174;
  assign n23176 = ~n23173 & ~n23174;
  assign n23177 = ~n23175 & ~n23176;
  assign n23178 = n6539 & n8963;
  assign n23179 = pi113  & n6873;
  assign n23180 = pi115  & n6537;
  assign n23181 = pi114  & n6532;
  assign n23182 = ~n23180 & ~n23181;
  assign n23183 = ~n23179 & n23182;
  assign n23184 = ~n23178 & n23183;
  assign n23185 = pi44  & ~n23184;
  assign n23186 = pi44  & ~n23185;
  assign n23187 = ~n23184 & ~n23185;
  assign n23188 = ~n23186 & ~n23187;
  assign n23189 = ~n23177 & n23188;
  assign n23190 = n23177 & ~n23188;
  assign n23191 = ~n23054 & ~n23189;
  assign n23192 = ~n23190 & n23191;
  assign n23193 = ~n23054 & ~n23192;
  assign n23194 = ~n23190 & ~n23192;
  assign n23195 = ~n23189 & n23194;
  assign n23196 = ~n23193 & ~n23195;
  assign n23197 = n5739 & n9984;
  assign n23198 = pi116  & n6030;
  assign n23199 = pi118  & n5737;
  assign n23200 = pi117  & n5732;
  assign n23201 = ~n23199 & ~n23200;
  assign n23202 = ~n23198 & n23201;
  assign n23203 = ~n23197 & n23202;
  assign n23204 = pi41  & ~n23203;
  assign n23205 = pi41  & ~n23204;
  assign n23206 = ~n23203 & ~n23204;
  assign n23207 = ~n23205 & ~n23206;
  assign n23208 = n23196 & n23207;
  assign n23209 = ~n23196 & ~n23207;
  assign n23210 = ~n23208 & ~n23209;
  assign n23211 = ~n23053 & n23210;
  assign n23212 = n23053 & ~n23210;
  assign n23213 = ~n23211 & ~n23212;
  assign n23214 = n5008 & n11389;
  assign n23215 = pi119  & n5241;
  assign n23216 = pi121  & n5006;
  assign n23217 = pi120  & n5001;
  assign n23218 = ~n23216 & ~n23217;
  assign n23219 = ~n23215 & n23218;
  assign n23220 = ~n23214 & n23219;
  assign n23221 = pi38  & ~n23220;
  assign n23222 = pi38  & ~n23221;
  assign n23223 = ~n23220 & ~n23221;
  assign n23224 = ~n23222 & ~n23223;
  assign n23225 = n23213 & ~n23224;
  assign n23226 = n23213 & ~n23225;
  assign n23227 = ~n23224 & ~n23225;
  assign n23228 = ~n23226 & ~n23227;
  assign n23229 = ~n23014 & ~n23017;
  assign n23230 = n23228 & n23229;
  assign n23231 = ~n23228 & ~n23229;
  assign n23232 = ~n23230 & ~n23231;
  assign n23233 = n4271 & n12189;
  assign n23234 = pi122  & n4503;
  assign n23235 = pi124  & n4269;
  assign n23236 = pi123  & n4264;
  assign n23237 = ~n23235 & ~n23236;
  assign n23238 = ~n23234 & n23237;
  assign n23239 = ~n23233 & n23238;
  assign n23240 = pi35  & ~n23239;
  assign n23241 = pi35  & ~n23240;
  assign n23242 = ~n23239 & ~n23240;
  assign n23243 = ~n23241 & ~n23242;
  assign n23244 = n23232 & ~n23243;
  assign n23245 = n23232 & ~n23244;
  assign n23246 = ~n23243 & ~n23244;
  assign n23247 = ~n23245 & ~n23246;
  assign n23248 = ~n23020 & ~n23034;
  assign n23249 = n23247 & n23248;
  assign n23250 = ~n23247 & ~n23248;
  assign n23251 = ~n23249 & ~n23250;
  assign n23252 = ~n22845 & ~n23039;
  assign n23253 = n3622 & n13742;
  assign n23254 = pi125  & n3814;
  assign n23255 = pi127  & n3620;
  assign n23256 = pi126  & n3615;
  assign n23257 = ~n23255 & ~n23256;
  assign n23258 = ~n23254 & n23257;
  assign n23259 = ~n23253 & n23258;
  assign n23260 = pi32  & ~n23259;
  assign n23261 = pi32  & ~n23260;
  assign n23262 = ~n23259 & ~n23260;
  assign n23263 = ~n23261 & ~n23262;
  assign n23264 = ~n23252 & ~n23263;
  assign n23265 = ~n23252 & ~n23264;
  assign n23266 = ~n23263 & ~n23264;
  assign n23267 = ~n23265 & ~n23266;
  assign n23268 = ~n23251 & n23267;
  assign n23269 = n23251 & ~n23267;
  assign n23270 = ~n23268 & ~n23269;
  assign n23271 = ~n23052 & n23270;
  assign n23272 = n23052 & ~n23270;
  assign n23273 = ~n23271 & ~n23272;
  assign n23274 = ~n23051 & n23273;
  assign n23275 = n23051 & ~n23273;
  assign po93  = ~n23274 & ~n23275;
  assign n23277 = ~n23244 & ~n23250;
  assign n23278 = pi126  & n3814;
  assign n23279 = pi127  & n3615;
  assign n23280 = ~n23278 & ~n23279;
  assign n23281 = ~n3622 & n23280;
  assign n23282 = n13773 & n23280;
  assign n23283 = ~n23281 & ~n23282;
  assign n23284 = pi32  & ~n23283;
  assign n23285 = ~pi32  & n23283;
  assign n23286 = ~n23284 & ~n23285;
  assign n23287 = ~n23277 & ~n23286;
  assign n23288 = n23277 & n23286;
  assign n23289 = ~n23287 & ~n23288;
  assign n23290 = ~n23209 & ~n23211;
  assign n23291 = ~n23116 & ~n23122;
  assign n23292 = n5943 & n10394;
  assign n23293 = pi102  & n10744;
  assign n23294 = pi104  & n10392;
  assign n23295 = pi103  & n10387;
  assign n23296 = ~n23294 & ~n23295;
  assign n23297 = ~n23293 & n23296;
  assign n23298 = ~n23292 & n23297;
  assign n23299 = pi56  & ~n23298;
  assign n23300 = pi56  & ~n23299;
  assign n23301 = ~n23298 & ~n23299;
  assign n23302 = ~n23300 & ~n23301;
  assign n23303 = ~n23099 & ~n23102;
  assign n23304 = n5169 & n11488;
  assign n23305 = pi99  & n11847;
  assign n23306 = pi101  & n11486;
  assign n23307 = pi100  & n11481;
  assign n23308 = ~n23306 & ~n23307;
  assign n23309 = ~n23305 & n23308;
  assign n23310 = ~n23304 & n23309;
  assign n23311 = pi59  & ~n23310;
  assign n23312 = pi59  & ~n23311;
  assign n23313 = ~n23310 & ~n23311;
  assign n23314 = ~n23312 & ~n23313;
  assign n23315 = ~n23073 & ~n23084;
  assign n23316 = ~n23070 & ~n23315;
  assign n23317 = pi94  & n13835;
  assign n23318 = pi95  & ~n13434;
  assign n23319 = ~n23317 & ~n23318;
  assign n23320 = ~n23063 & ~n23066;
  assign n23321 = ~n23319 & n23320;
  assign n23322 = n23319 & ~n23320;
  assign n23323 = ~n23321 & ~n23322;
  assign n23324 = n4454 & n12627;
  assign n23325 = pi96  & n13004;
  assign n23326 = pi98  & n12625;
  assign n23327 = pi97  & n12620;
  assign n23328 = ~n23326 & ~n23327;
  assign n23329 = ~n23325 & n23328;
  assign n23330 = ~n23324 & n23329;
  assign n23331 = pi62  & ~n23330;
  assign n23332 = pi62  & ~n23331;
  assign n23333 = ~n23330 & ~n23331;
  assign n23334 = ~n23332 & ~n23333;
  assign n23335 = ~n23323 & n23334;
  assign n23336 = n23323 & ~n23334;
  assign n23337 = ~n23335 & ~n23336;
  assign n23338 = ~n23316 & n23337;
  assign n23339 = ~n23316 & ~n23338;
  assign n23340 = n23337 & ~n23338;
  assign n23341 = ~n23339 & ~n23340;
  assign n23342 = ~n23314 & ~n23341;
  assign n23343 = n23314 & n23341;
  assign n23344 = ~n23342 & ~n23343;
  assign n23345 = ~n23303 & n23344;
  assign n23346 = ~n23303 & ~n23345;
  assign n23347 = n23344 & ~n23345;
  assign n23348 = ~n23346 & ~n23347;
  assign n23349 = ~n23302 & ~n23348;
  assign n23350 = n23302 & n23348;
  assign n23351 = ~n23349 & ~n23350;
  assign n23352 = ~n23291 & n23351;
  assign n23353 = n23291 & ~n23351;
  assign n23354 = ~n23352 & ~n23353;
  assign n23355 = n6775 & n9310;
  assign n23356 = pi105  & n9701;
  assign n23357 = pi107  & n9308;
  assign n23358 = pi106  & n9303;
  assign n23359 = ~n23357 & ~n23358;
  assign n23360 = ~n23356 & n23359;
  assign n23361 = ~n23355 & n23360;
  assign n23362 = pi53  & ~n23361;
  assign n23363 = pi53  & ~n23362;
  assign n23364 = ~n23361 & ~n23362;
  assign n23365 = ~n23363 & ~n23364;
  assign n23366 = n23354 & ~n23365;
  assign n23367 = n23354 & ~n23366;
  assign n23368 = ~n23365 & ~n23366;
  assign n23369 = ~n23367 & ~n23368;
  assign n23370 = ~n23057 & ~n23138;
  assign n23371 = ~n23135 & ~n23370;
  assign n23372 = n23369 & n23371;
  assign n23373 = ~n23369 & ~n23371;
  assign n23374 = ~n23372 & ~n23373;
  assign n23375 = n7665 & n8334;
  assign n23376 = pi108  & n8685;
  assign n23377 = pi110  & n8332;
  assign n23378 = pi109  & n8327;
  assign n23379 = ~n23377 & ~n23378;
  assign n23380 = ~n23376 & n23379;
  assign n23381 = ~n23375 & n23380;
  assign n23382 = pi50  & ~n23381;
  assign n23383 = pi50  & ~n23382;
  assign n23384 = ~n23381 & ~n23382;
  assign n23385 = ~n23383 & ~n23384;
  assign n23386 = n23374 & ~n23385;
  assign n23387 = n23374 & ~n23386;
  assign n23388 = ~n23385 & ~n23386;
  assign n23389 = ~n23387 & ~n23388;
  assign n23390 = ~n23153 & ~n23157;
  assign n23391 = n23389 & n23390;
  assign n23392 = ~n23389 & ~n23390;
  assign n23393 = ~n23391 & ~n23392;
  assign n23394 = n7408 & n8612;
  assign n23395 = pi111  & n7740;
  assign n23396 = pi113  & n7406;
  assign n23397 = pi112  & n7401;
  assign n23398 = ~n23396 & ~n23397;
  assign n23399 = ~n23395 & n23398;
  assign n23400 = ~n23394 & n23399;
  assign n23401 = pi47  & ~n23400;
  assign n23402 = pi47  & ~n23401;
  assign n23403 = ~n23400 & ~n23401;
  assign n23404 = ~n23402 & ~n23403;
  assign n23405 = n23393 & ~n23404;
  assign n23406 = n23393 & ~n23405;
  assign n23407 = ~n23404 & ~n23405;
  assign n23408 = ~n23406 & ~n23407;
  assign n23409 = ~n23170 & ~n23176;
  assign n23410 = n23408 & n23409;
  assign n23411 = ~n23408 & ~n23409;
  assign n23412 = ~n23410 & ~n23411;
  assign n23413 = n6539 & n9614;
  assign n23414 = pi114  & n6873;
  assign n23415 = pi116  & n6537;
  assign n23416 = pi115  & n6532;
  assign n23417 = ~n23415 & ~n23416;
  assign n23418 = ~n23414 & n23417;
  assign n23419 = ~n23413 & n23418;
  assign n23420 = pi44  & ~n23419;
  assign n23421 = pi44  & ~n23420;
  assign n23422 = ~n23419 & ~n23420;
  assign n23423 = ~n23421 & ~n23422;
  assign n23424 = n23412 & ~n23423;
  assign n23425 = n23412 & ~n23424;
  assign n23426 = ~n23423 & ~n23424;
  assign n23427 = ~n23425 & ~n23426;
  assign n23428 = ~n23194 & n23427;
  assign n23429 = n23194 & ~n23427;
  assign n23430 = ~n23428 & ~n23429;
  assign n23431 = n5739 & n10667;
  assign n23432 = pi117  & n6030;
  assign n23433 = pi119  & n5737;
  assign n23434 = pi118  & n5732;
  assign n23435 = ~n23433 & ~n23434;
  assign n23436 = ~n23432 & n23435;
  assign n23437 = ~n23431 & n23436;
  assign n23438 = pi41  & ~n23437;
  assign n23439 = pi41  & ~n23438;
  assign n23440 = ~n23437 & ~n23438;
  assign n23441 = ~n23439 & ~n23440;
  assign n23442 = ~n23430 & ~n23441;
  assign n23443 = n23430 & n23441;
  assign n23444 = ~n23442 & ~n23443;
  assign n23445 = ~n23290 & n23444;
  assign n23446 = n23290 & ~n23444;
  assign n23447 = ~n23445 & ~n23446;
  assign n23448 = n5008 & n11778;
  assign n23449 = pi120  & n5241;
  assign n23450 = pi122  & n5006;
  assign n23451 = pi121  & n5001;
  assign n23452 = ~n23450 & ~n23451;
  assign n23453 = ~n23449 & n23452;
  assign n23454 = ~n23448 & n23453;
  assign n23455 = pi38  & ~n23454;
  assign n23456 = pi38  & ~n23455;
  assign n23457 = ~n23454 & ~n23455;
  assign n23458 = ~n23456 & ~n23457;
  assign n23459 = n23447 & ~n23458;
  assign n23460 = n23447 & ~n23459;
  assign n23461 = ~n23458 & ~n23459;
  assign n23462 = ~n23460 & ~n23461;
  assign n23463 = ~n23225 & ~n23231;
  assign n23464 = n23462 & n23463;
  assign n23465 = ~n23462 & ~n23463;
  assign n23466 = ~n23464 & ~n23465;
  assign n23467 = n4271 & n12943;
  assign n23468 = pi123  & n4503;
  assign n23469 = pi125  & n4269;
  assign n23470 = pi124  & n4264;
  assign n23471 = ~n23469 & ~n23470;
  assign n23472 = ~n23468 & n23471;
  assign n23473 = ~n23467 & n23472;
  assign n23474 = pi35  & ~n23473;
  assign n23475 = pi35  & ~n23474;
  assign n23476 = ~n23473 & ~n23474;
  assign n23477 = ~n23475 & ~n23476;
  assign n23478 = n23466 & ~n23477;
  assign n23479 = ~n23466 & n23477;
  assign n23480 = ~n23478 & ~n23479;
  assign n23481 = n23289 & n23480;
  assign n23482 = n23289 & ~n23481;
  assign n23483 = n23480 & ~n23481;
  assign n23484 = ~n23482 & ~n23483;
  assign n23485 = ~n23264 & ~n23269;
  assign n23486 = ~n23484 & ~n23485;
  assign n23487 = ~n23484 & ~n23486;
  assign n23488 = ~n23485 & ~n23486;
  assign n23489 = ~n23487 & ~n23488;
  assign n23490 = ~n23271 & ~n23274;
  assign n23491 = ~n23489 & ~n23490;
  assign n23492 = n23489 & n23490;
  assign po94  = ~n23491 & ~n23492;
  assign n23494 = ~n23486 & ~n23491;
  assign n23495 = ~n23287 & ~n23481;
  assign n23496 = ~n23465 & ~n23478;
  assign n23497 = pi127  & n3814;
  assign n23498 = n3622 & n13770;
  assign n23499 = ~n23497 & ~n23498;
  assign n23500 = pi32  & ~n23499;
  assign n23501 = pi32  & ~n23500;
  assign n23502 = ~n23499 & ~n23500;
  assign n23503 = ~n23501 & ~n23502;
  assign n23504 = ~n23496 & ~n23503;
  assign n23505 = ~n23496 & ~n23504;
  assign n23506 = ~n23503 & ~n23504;
  assign n23507 = ~n23505 & ~n23506;
  assign n23508 = ~n23194 & ~n23427;
  assign n23509 = ~n23442 & ~n23508;
  assign n23510 = n5739 & n11028;
  assign n23511 = pi118  & n6030;
  assign n23512 = pi120  & n5737;
  assign n23513 = pi119  & n5732;
  assign n23514 = ~n23512 & ~n23513;
  assign n23515 = ~n23511 & n23514;
  assign n23516 = ~n23510 & n23515;
  assign n23517 = pi41  & ~n23516;
  assign n23518 = pi41  & ~n23517;
  assign n23519 = ~n23516 & ~n23517;
  assign n23520 = ~n23518 & ~n23519;
  assign n23521 = ~n23411 & ~n23424;
  assign n23522 = n6539 & n9958;
  assign n23523 = pi115  & n6873;
  assign n23524 = pi117  & n6537;
  assign n23525 = pi116  & n6532;
  assign n23526 = ~n23524 & ~n23525;
  assign n23527 = ~n23523 & n23526;
  assign n23528 = ~n23522 & n23527;
  assign n23529 = pi44  & ~n23528;
  assign n23530 = pi44  & ~n23529;
  assign n23531 = ~n23528 & ~n23529;
  assign n23532 = ~n23530 & ~n23531;
  assign n23533 = ~n23392 & ~n23405;
  assign n23534 = ~n23352 & ~n23366;
  assign n23535 = n7060 & n9310;
  assign n23536 = pi106  & n9701;
  assign n23537 = pi108  & n9308;
  assign n23538 = pi107  & n9303;
  assign n23539 = ~n23537 & ~n23538;
  assign n23540 = ~n23536 & n23539;
  assign n23541 = ~n23535 & n23540;
  assign n23542 = pi53  & ~n23541;
  assign n23543 = pi53  & ~n23542;
  assign n23544 = ~n23541 & ~n23542;
  assign n23545 = ~n23543 & ~n23544;
  assign n23546 = ~n23345 & ~n23349;
  assign n23547 = n6207 & n10394;
  assign n23548 = pi103  & n10744;
  assign n23549 = pi105  & n10392;
  assign n23550 = pi104  & n10387;
  assign n23551 = ~n23549 & ~n23550;
  assign n23552 = ~n23548 & n23551;
  assign n23553 = ~n23547 & n23552;
  assign n23554 = pi56  & ~n23553;
  assign n23555 = pi56  & ~n23554;
  assign n23556 = ~n23553 & ~n23554;
  assign n23557 = ~n23555 & ~n23556;
  assign n23558 = ~n23338 & ~n23342;
  assign n23559 = ~n23322 & ~n23336;
  assign n23560 = pi95  & n13835;
  assign n23561 = pi96  & ~n13434;
  assign n23562 = ~n23560 & ~n23561;
  assign n23563 = ~n23319 & n23562;
  assign n23564 = n23319 & ~n23562;
  assign n23565 = ~n23563 & ~n23564;
  assign n23566 = ~n23559 & n23565;
  assign n23567 = ~n23559 & ~n23566;
  assign n23568 = ~n23563 & ~n23566;
  assign n23569 = ~n23564 & n23568;
  assign n23570 = ~n23567 & ~n23569;
  assign n23571 = n4684 & n12627;
  assign n23572 = pi97  & n13004;
  assign n23573 = pi99  & n12625;
  assign n23574 = pi98  & n12620;
  assign n23575 = ~n23573 & ~n23574;
  assign n23576 = ~n23572 & n23575;
  assign n23577 = ~n23571 & n23576;
  assign n23578 = pi62  & ~n23577;
  assign n23579 = pi62  & ~n23578;
  assign n23580 = ~n23577 & ~n23578;
  assign n23581 = ~n23579 & ~n23580;
  assign n23582 = ~n23570 & ~n23581;
  assign n23583 = ~n23570 & ~n23582;
  assign n23584 = ~n23581 & ~n23582;
  assign n23585 = ~n23583 & ~n23584;
  assign n23586 = n5413 & n11488;
  assign n23587 = pi100  & n11847;
  assign n23588 = pi102  & n11486;
  assign n23589 = pi101  & n11481;
  assign n23590 = ~n23588 & ~n23589;
  assign n23591 = ~n23587 & n23590;
  assign n23592 = ~n23586 & n23591;
  assign n23593 = pi59  & ~n23592;
  assign n23594 = pi59  & ~n23593;
  assign n23595 = ~n23592 & ~n23593;
  assign n23596 = ~n23594 & ~n23595;
  assign n23597 = ~n23585 & n23596;
  assign n23598 = n23585 & ~n23596;
  assign n23599 = ~n23597 & ~n23598;
  assign n23600 = ~n23558 & ~n23599;
  assign n23601 = n23558 & n23599;
  assign n23602 = ~n23600 & ~n23601;
  assign n23603 = ~n23557 & n23602;
  assign n23604 = n23557 & ~n23602;
  assign n23605 = ~n23603 & ~n23604;
  assign n23606 = ~n23546 & n23605;
  assign n23607 = n23546 & ~n23605;
  assign n23608 = ~n23606 & ~n23607;
  assign n23609 = ~n23545 & n23608;
  assign n23610 = n23545 & ~n23608;
  assign n23611 = ~n23609 & ~n23610;
  assign n23612 = ~n23534 & n23611;
  assign n23613 = n23534 & ~n23611;
  assign n23614 = ~n23612 & ~n23613;
  assign n23615 = n7970 & n8334;
  assign n23616 = pi109  & n8685;
  assign n23617 = pi111  & n8332;
  assign n23618 = pi110  & n8327;
  assign n23619 = ~n23617 & ~n23618;
  assign n23620 = ~n23616 & n23619;
  assign n23621 = ~n23615 & n23620;
  assign n23622 = pi50  & ~n23621;
  assign n23623 = pi50  & ~n23622;
  assign n23624 = ~n23621 & ~n23622;
  assign n23625 = ~n23623 & ~n23624;
  assign n23626 = n23614 & ~n23625;
  assign n23627 = n23614 & ~n23626;
  assign n23628 = ~n23625 & ~n23626;
  assign n23629 = ~n23627 & ~n23628;
  assign n23630 = ~n23373 & ~n23386;
  assign n23631 = n23629 & n23630;
  assign n23632 = ~n23629 & ~n23630;
  assign n23633 = ~n23631 & ~n23632;
  assign n23634 = n7408 & n8936;
  assign n23635 = pi112  & n7740;
  assign n23636 = pi114  & n7406;
  assign n23637 = pi113  & n7401;
  assign n23638 = ~n23636 & ~n23637;
  assign n23639 = ~n23635 & n23638;
  assign n23640 = ~n23634 & n23639;
  assign n23641 = pi47  & ~n23640;
  assign n23642 = pi47  & ~n23641;
  assign n23643 = ~n23640 & ~n23641;
  assign n23644 = ~n23642 & ~n23643;
  assign n23645 = ~n23633 & n23644;
  assign n23646 = n23633 & ~n23644;
  assign n23647 = ~n23645 & ~n23646;
  assign n23648 = ~n23533 & n23647;
  assign n23649 = ~n23533 & ~n23648;
  assign n23650 = n23647 & ~n23648;
  assign n23651 = ~n23649 & ~n23650;
  assign n23652 = ~n23532 & ~n23651;
  assign n23653 = n23532 & n23651;
  assign n23654 = ~n23652 & ~n23653;
  assign n23655 = ~n23521 & n23654;
  assign n23656 = n23521 & ~n23654;
  assign n23657 = ~n23655 & ~n23656;
  assign n23658 = ~n23520 & n23657;
  assign n23659 = n23520 & ~n23657;
  assign n23660 = ~n23658 & ~n23659;
  assign n23661 = ~n23509 & n23660;
  assign n23662 = n23509 & ~n23660;
  assign n23663 = ~n23661 & ~n23662;
  assign n23664 = n5008 & n12158;
  assign n23665 = pi121  & n5241;
  assign n23666 = pi123  & n5006;
  assign n23667 = pi122  & n5001;
  assign n23668 = ~n23666 & ~n23667;
  assign n23669 = ~n23665 & n23668;
  assign n23670 = ~n23664 & n23669;
  assign n23671 = pi38  & ~n23670;
  assign n23672 = pi38  & ~n23671;
  assign n23673 = ~n23670 & ~n23671;
  assign n23674 = ~n23672 & ~n23673;
  assign n23675 = n23663 & ~n23674;
  assign n23676 = n23663 & ~n23675;
  assign n23677 = ~n23674 & ~n23675;
  assign n23678 = ~n23676 & ~n23677;
  assign n23679 = ~n23445 & ~n23459;
  assign n23680 = n23678 & n23679;
  assign n23681 = ~n23678 & ~n23679;
  assign n23682 = ~n23680 & ~n23681;
  assign n23683 = n4271 & n13344;
  assign n23684 = pi124  & n4503;
  assign n23685 = pi126  & n4269;
  assign n23686 = pi125  & n4264;
  assign n23687 = ~n23685 & ~n23686;
  assign n23688 = ~n23684 & n23687;
  assign n23689 = ~n23683 & n23688;
  assign n23690 = pi35  & ~n23689;
  assign n23691 = pi35  & ~n23690;
  assign n23692 = ~n23689 & ~n23690;
  assign n23693 = ~n23691 & ~n23692;
  assign n23694 = n23682 & ~n23693;
  assign n23695 = n23682 & ~n23694;
  assign n23696 = ~n23693 & ~n23694;
  assign n23697 = ~n23695 & ~n23696;
  assign n23698 = ~n23507 & n23697;
  assign n23699 = n23507 & ~n23697;
  assign n23700 = ~n23698 & ~n23699;
  assign n23701 = ~n23495 & ~n23700;
  assign n23702 = ~n23495 & ~n23701;
  assign n23703 = ~n23700 & ~n23701;
  assign n23704 = ~n23702 & ~n23703;
  assign n23705 = ~n23494 & ~n23704;
  assign n23706 = n23494 & n23704;
  assign po95  = ~n23705 & ~n23706;
  assign n23708 = ~n23701 & ~n23705;
  assign n23709 = ~n23507 & ~n23697;
  assign n23710 = ~n23504 & ~n23709;
  assign n23711 = ~n23648 & ~n23652;
  assign n23712 = ~n23632 & ~n23646;
  assign n23713 = ~n23585 & ~n23596;
  assign n23714 = ~n23582 & ~n23713;
  assign n23715 = pi96  & n13835;
  assign n23716 = pi97  & ~n13434;
  assign n23717 = ~n23715 & ~n23716;
  assign n23718 = ~pi32  & ~n23717;
  assign n23719 = pi32  & n23717;
  assign n23720 = ~n23718 & ~n23719;
  assign n23721 = ~n23562 & n23720;
  assign n23722 = ~n23562 & ~n23721;
  assign n23723 = n23720 & ~n23721;
  assign n23724 = ~n23722 & ~n23723;
  assign n23725 = ~n23568 & ~n23724;
  assign n23726 = ~n23568 & ~n23725;
  assign n23727 = ~n23724 & ~n23725;
  assign n23728 = ~n23726 & ~n23727;
  assign n23729 = n4910 & n12627;
  assign n23730 = pi98  & n13004;
  assign n23731 = pi100  & n12625;
  assign n23732 = pi99  & n12620;
  assign n23733 = ~n23731 & ~n23732;
  assign n23734 = ~n23730 & n23733;
  assign n23735 = ~n23729 & n23734;
  assign n23736 = pi62  & ~n23735;
  assign n23737 = pi62  & ~n23736;
  assign n23738 = ~n23735 & ~n23736;
  assign n23739 = ~n23737 & ~n23738;
  assign n23740 = ~n23728 & n23739;
  assign n23741 = n23728 & ~n23739;
  assign n23742 = ~n23740 & ~n23741;
  assign n23743 = n5664 & n11488;
  assign n23744 = pi101  & n11847;
  assign n23745 = pi103  & n11486;
  assign n23746 = pi102  & n11481;
  assign n23747 = ~n23745 & ~n23746;
  assign n23748 = ~n23744 & n23747;
  assign n23749 = ~n23743 & n23748;
  assign n23750 = pi59  & ~n23749;
  assign n23751 = pi59  & ~n23750;
  assign n23752 = ~n23749 & ~n23750;
  assign n23753 = ~n23751 & ~n23752;
  assign n23754 = ~n23742 & ~n23753;
  assign n23755 = n23742 & n23753;
  assign n23756 = ~n23754 & ~n23755;
  assign n23757 = ~n23714 & n23756;
  assign n23758 = n23714 & ~n23756;
  assign n23759 = ~n23757 & ~n23758;
  assign n23760 = n6477 & n10394;
  assign n23761 = pi104  & n10744;
  assign n23762 = pi106  & n10392;
  assign n23763 = pi105  & n10387;
  assign n23764 = ~n23762 & ~n23763;
  assign n23765 = ~n23761 & n23764;
  assign n23766 = ~n23760 & n23765;
  assign n23767 = pi56  & ~n23766;
  assign n23768 = pi56  & ~n23767;
  assign n23769 = ~n23766 & ~n23767;
  assign n23770 = ~n23768 & ~n23769;
  assign n23771 = n23759 & ~n23770;
  assign n23772 = n23759 & ~n23771;
  assign n23773 = ~n23770 & ~n23771;
  assign n23774 = ~n23772 & ~n23773;
  assign n23775 = ~n23600 & ~n23603;
  assign n23776 = n23774 & n23775;
  assign n23777 = ~n23774 & ~n23775;
  assign n23778 = ~n23776 & ~n23777;
  assign n23779 = n7349 & n9310;
  assign n23780 = pi107  & n9701;
  assign n23781 = pi109  & n9308;
  assign n23782 = pi108  & n9303;
  assign n23783 = ~n23781 & ~n23782;
  assign n23784 = ~n23780 & n23783;
  assign n23785 = ~n23779 & n23784;
  assign n23786 = pi53  & ~n23785;
  assign n23787 = pi53  & ~n23786;
  assign n23788 = ~n23785 & ~n23786;
  assign n23789 = ~n23787 & ~n23788;
  assign n23790 = n23778 & ~n23789;
  assign n23791 = n23778 & ~n23790;
  assign n23792 = ~n23789 & ~n23790;
  assign n23793 = ~n23791 & ~n23792;
  assign n23794 = ~n23606 & ~n23609;
  assign n23795 = n23793 & n23794;
  assign n23796 = ~n23793 & ~n23794;
  assign n23797 = ~n23795 & ~n23796;
  assign n23798 = n7997 & n8334;
  assign n23799 = pi110  & n8685;
  assign n23800 = pi112  & n8332;
  assign n23801 = pi111  & n8327;
  assign n23802 = ~n23800 & ~n23801;
  assign n23803 = ~n23799 & n23802;
  assign n23804 = ~n23798 & n23803;
  assign n23805 = pi50  & ~n23804;
  assign n23806 = pi50  & ~n23805;
  assign n23807 = ~n23804 & ~n23805;
  assign n23808 = ~n23806 & ~n23807;
  assign n23809 = n23797 & ~n23808;
  assign n23810 = n23797 & ~n23809;
  assign n23811 = ~n23808 & ~n23809;
  assign n23812 = ~n23810 & ~n23811;
  assign n23813 = ~n23612 & ~n23626;
  assign n23814 = n23812 & n23813;
  assign n23815 = ~n23812 & ~n23813;
  assign n23816 = ~n23814 & ~n23815;
  assign n23817 = n7408 & n8963;
  assign n23818 = pi113  & n7740;
  assign n23819 = pi115  & n7406;
  assign n23820 = pi114  & n7401;
  assign n23821 = ~n23819 & ~n23820;
  assign n23822 = ~n23818 & n23821;
  assign n23823 = ~n23817 & n23822;
  assign n23824 = pi47  & ~n23823;
  assign n23825 = pi47  & ~n23824;
  assign n23826 = ~n23823 & ~n23824;
  assign n23827 = ~n23825 & ~n23826;
  assign n23828 = ~n23816 & n23827;
  assign n23829 = n23816 & ~n23827;
  assign n23830 = ~n23712 & ~n23828;
  assign n23831 = ~n23829 & n23830;
  assign n23832 = ~n23712 & ~n23831;
  assign n23833 = ~n23829 & ~n23831;
  assign n23834 = ~n23828 & n23833;
  assign n23835 = ~n23832 & ~n23834;
  assign n23836 = n6539 & n9984;
  assign n23837 = pi116  & n6873;
  assign n23838 = pi118  & n6537;
  assign n23839 = pi117  & n6532;
  assign n23840 = ~n23838 & ~n23839;
  assign n23841 = ~n23837 & n23840;
  assign n23842 = ~n23836 & n23841;
  assign n23843 = pi44  & ~n23842;
  assign n23844 = pi44  & ~n23843;
  assign n23845 = ~n23842 & ~n23843;
  assign n23846 = ~n23844 & ~n23845;
  assign n23847 = n23835 & n23846;
  assign n23848 = ~n23835 & ~n23846;
  assign n23849 = ~n23847 & ~n23848;
  assign n23850 = ~n23711 & n23849;
  assign n23851 = n23711 & ~n23849;
  assign n23852 = ~n23850 & ~n23851;
  assign n23853 = n5739 & n11389;
  assign n23854 = pi119  & n6030;
  assign n23855 = pi121  & n5737;
  assign n23856 = pi120  & n5732;
  assign n23857 = ~n23855 & ~n23856;
  assign n23858 = ~n23854 & n23857;
  assign n23859 = ~n23853 & n23858;
  assign n23860 = pi41  & ~n23859;
  assign n23861 = pi41  & ~n23860;
  assign n23862 = ~n23859 & ~n23860;
  assign n23863 = ~n23861 & ~n23862;
  assign n23864 = n23852 & ~n23863;
  assign n23865 = n23852 & ~n23864;
  assign n23866 = ~n23863 & ~n23864;
  assign n23867 = ~n23865 & ~n23866;
  assign n23868 = ~n23655 & ~n23658;
  assign n23869 = n23867 & n23868;
  assign n23870 = ~n23867 & ~n23868;
  assign n23871 = ~n23869 & ~n23870;
  assign n23872 = n5008 & n12189;
  assign n23873 = pi122  & n5241;
  assign n23874 = pi124  & n5006;
  assign n23875 = pi123  & n5001;
  assign n23876 = ~n23874 & ~n23875;
  assign n23877 = ~n23873 & n23876;
  assign n23878 = ~n23872 & n23877;
  assign n23879 = pi38  & ~n23878;
  assign n23880 = pi38  & ~n23879;
  assign n23881 = ~n23878 & ~n23879;
  assign n23882 = ~n23880 & ~n23881;
  assign n23883 = n23871 & ~n23882;
  assign n23884 = n23871 & ~n23883;
  assign n23885 = ~n23882 & ~n23883;
  assign n23886 = ~n23884 & ~n23885;
  assign n23887 = ~n23661 & ~n23675;
  assign n23888 = n23886 & n23887;
  assign n23889 = ~n23886 & ~n23887;
  assign n23890 = ~n23888 & ~n23889;
  assign n23891 = ~n23681 & ~n23694;
  assign n23892 = n4271 & n13742;
  assign n23893 = pi125  & n4503;
  assign n23894 = pi127  & n4269;
  assign n23895 = pi126  & n4264;
  assign n23896 = ~n23894 & ~n23895;
  assign n23897 = ~n23893 & n23896;
  assign n23898 = ~n23892 & n23897;
  assign n23899 = pi35  & ~n23898;
  assign n23900 = pi35  & ~n23899;
  assign n23901 = ~n23898 & ~n23899;
  assign n23902 = ~n23900 & ~n23901;
  assign n23903 = ~n23891 & ~n23902;
  assign n23904 = ~n23891 & ~n23903;
  assign n23905 = ~n23902 & ~n23903;
  assign n23906 = ~n23904 & ~n23905;
  assign n23907 = ~n23890 & n23906;
  assign n23908 = n23890 & ~n23906;
  assign n23909 = ~n23907 & ~n23908;
  assign n23910 = ~n23710 & n23909;
  assign n23911 = n23710 & ~n23909;
  assign n23912 = ~n23910 & ~n23911;
  assign n23913 = ~n23708 & n23912;
  assign n23914 = n23708 & ~n23912;
  assign po96  = ~n23913 & ~n23914;
  assign n23916 = ~n23883 & ~n23889;
  assign n23917 = pi126  & n4503;
  assign n23918 = pi127  & n4264;
  assign n23919 = ~n23917 & ~n23918;
  assign n23920 = ~n4271 & n23919;
  assign n23921 = n13773 & n23919;
  assign n23922 = ~n23920 & ~n23921;
  assign n23923 = pi35  & ~n23922;
  assign n23924 = ~pi35  & n23922;
  assign n23925 = ~n23923 & ~n23924;
  assign n23926 = ~n23916 & ~n23925;
  assign n23927 = n23916 & n23925;
  assign n23928 = ~n23926 & ~n23927;
  assign n23929 = ~n23848 & ~n23850;
  assign n23930 = ~n23754 & ~n23757;
  assign n23931 = n5943 & n11488;
  assign n23932 = pi102  & n11847;
  assign n23933 = pi104  & n11486;
  assign n23934 = pi103  & n11481;
  assign n23935 = ~n23933 & ~n23934;
  assign n23936 = ~n23932 & n23935;
  assign n23937 = ~n23931 & n23936;
  assign n23938 = pi59  & ~n23937;
  assign n23939 = pi59  & ~n23938;
  assign n23940 = ~n23937 & ~n23938;
  assign n23941 = ~n23939 & ~n23940;
  assign n23942 = ~n23728 & ~n23739;
  assign n23943 = ~n23725 & ~n23942;
  assign n23944 = pi97  & n13835;
  assign n23945 = pi98  & ~n13434;
  assign n23946 = ~n23944 & ~n23945;
  assign n23947 = ~n23718 & ~n23721;
  assign n23948 = ~n23946 & n23947;
  assign n23949 = n23946 & ~n23947;
  assign n23950 = ~n23948 & ~n23949;
  assign n23951 = n5169 & n12627;
  assign n23952 = pi99  & n13004;
  assign n23953 = pi101  & n12625;
  assign n23954 = pi100  & n12620;
  assign n23955 = ~n23953 & ~n23954;
  assign n23956 = ~n23952 & n23955;
  assign n23957 = ~n23951 & n23956;
  assign n23958 = pi62  & ~n23957;
  assign n23959 = pi62  & ~n23958;
  assign n23960 = ~n23957 & ~n23958;
  assign n23961 = ~n23959 & ~n23960;
  assign n23962 = ~n23950 & n23961;
  assign n23963 = n23950 & ~n23961;
  assign n23964 = ~n23962 & ~n23963;
  assign n23965 = ~n23943 & n23964;
  assign n23966 = ~n23943 & ~n23965;
  assign n23967 = n23964 & ~n23965;
  assign n23968 = ~n23966 & ~n23967;
  assign n23969 = ~n23941 & ~n23968;
  assign n23970 = n23941 & n23968;
  assign n23971 = ~n23969 & ~n23970;
  assign n23972 = ~n23930 & n23971;
  assign n23973 = n23930 & ~n23971;
  assign n23974 = ~n23972 & ~n23973;
  assign n23975 = n6775 & n10394;
  assign n23976 = pi105  & n10744;
  assign n23977 = pi107  & n10392;
  assign n23978 = pi106  & n10387;
  assign n23979 = ~n23977 & ~n23978;
  assign n23980 = ~n23976 & n23979;
  assign n23981 = ~n23975 & n23980;
  assign n23982 = pi56  & ~n23981;
  assign n23983 = pi56  & ~n23982;
  assign n23984 = ~n23981 & ~n23982;
  assign n23985 = ~n23983 & ~n23984;
  assign n23986 = n23974 & ~n23985;
  assign n23987 = n23974 & ~n23986;
  assign n23988 = ~n23985 & ~n23986;
  assign n23989 = ~n23987 & ~n23988;
  assign n23990 = ~n23771 & ~n23777;
  assign n23991 = n23989 & n23990;
  assign n23992 = ~n23989 & ~n23990;
  assign n23993 = ~n23991 & ~n23992;
  assign n23994 = n7665 & n9310;
  assign n23995 = pi108  & n9701;
  assign n23996 = pi110  & n9308;
  assign n23997 = pi109  & n9303;
  assign n23998 = ~n23996 & ~n23997;
  assign n23999 = ~n23995 & n23998;
  assign n24000 = ~n23994 & n23999;
  assign n24001 = pi53  & ~n24000;
  assign n24002 = pi53  & ~n24001;
  assign n24003 = ~n24000 & ~n24001;
  assign n24004 = ~n24002 & ~n24003;
  assign n24005 = n23993 & ~n24004;
  assign n24006 = n23993 & ~n24005;
  assign n24007 = ~n24004 & ~n24005;
  assign n24008 = ~n24006 & ~n24007;
  assign n24009 = ~n23790 & ~n23796;
  assign n24010 = n24008 & n24009;
  assign n24011 = ~n24008 & ~n24009;
  assign n24012 = ~n24010 & ~n24011;
  assign n24013 = n8334 & n8612;
  assign n24014 = pi111  & n8685;
  assign n24015 = pi113  & n8332;
  assign n24016 = pi112  & n8327;
  assign n24017 = ~n24015 & ~n24016;
  assign n24018 = ~n24014 & n24017;
  assign n24019 = ~n24013 & n24018;
  assign n24020 = pi50  & ~n24019;
  assign n24021 = pi50  & ~n24020;
  assign n24022 = ~n24019 & ~n24020;
  assign n24023 = ~n24021 & ~n24022;
  assign n24024 = n24012 & ~n24023;
  assign n24025 = n24012 & ~n24024;
  assign n24026 = ~n24023 & ~n24024;
  assign n24027 = ~n24025 & ~n24026;
  assign n24028 = ~n23809 & ~n23815;
  assign n24029 = n24027 & n24028;
  assign n24030 = ~n24027 & ~n24028;
  assign n24031 = ~n24029 & ~n24030;
  assign n24032 = n7408 & n9614;
  assign n24033 = pi114  & n7740;
  assign n24034 = pi116  & n7406;
  assign n24035 = pi115  & n7401;
  assign n24036 = ~n24034 & ~n24035;
  assign n24037 = ~n24033 & n24036;
  assign n24038 = ~n24032 & n24037;
  assign n24039 = pi47  & ~n24038;
  assign n24040 = pi47  & ~n24039;
  assign n24041 = ~n24038 & ~n24039;
  assign n24042 = ~n24040 & ~n24041;
  assign n24043 = n24031 & ~n24042;
  assign n24044 = n24031 & ~n24043;
  assign n24045 = ~n24042 & ~n24043;
  assign n24046 = ~n24044 & ~n24045;
  assign n24047 = ~n23833 & n24046;
  assign n24048 = n23833 & ~n24046;
  assign n24049 = ~n24047 & ~n24048;
  assign n24050 = n6539 & n10667;
  assign n24051 = pi117  & n6873;
  assign n24052 = pi119  & n6537;
  assign n24053 = pi118  & n6532;
  assign n24054 = ~n24052 & ~n24053;
  assign n24055 = ~n24051 & n24054;
  assign n24056 = ~n24050 & n24055;
  assign n24057 = pi44  & ~n24056;
  assign n24058 = pi44  & ~n24057;
  assign n24059 = ~n24056 & ~n24057;
  assign n24060 = ~n24058 & ~n24059;
  assign n24061 = ~n24049 & ~n24060;
  assign n24062 = n24049 & n24060;
  assign n24063 = ~n24061 & ~n24062;
  assign n24064 = ~n23929 & n24063;
  assign n24065 = n23929 & ~n24063;
  assign n24066 = ~n24064 & ~n24065;
  assign n24067 = n5739 & n11778;
  assign n24068 = pi120  & n6030;
  assign n24069 = pi122  & n5737;
  assign n24070 = pi121  & n5732;
  assign n24071 = ~n24069 & ~n24070;
  assign n24072 = ~n24068 & n24071;
  assign n24073 = ~n24067 & n24072;
  assign n24074 = pi41  & ~n24073;
  assign n24075 = pi41  & ~n24074;
  assign n24076 = ~n24073 & ~n24074;
  assign n24077 = ~n24075 & ~n24076;
  assign n24078 = n24066 & ~n24077;
  assign n24079 = n24066 & ~n24078;
  assign n24080 = ~n24077 & ~n24078;
  assign n24081 = ~n24079 & ~n24080;
  assign n24082 = ~n23864 & ~n23870;
  assign n24083 = n24081 & n24082;
  assign n24084 = ~n24081 & ~n24082;
  assign n24085 = ~n24083 & ~n24084;
  assign n24086 = n5008 & n12943;
  assign n24087 = pi123  & n5241;
  assign n24088 = pi125  & n5006;
  assign n24089 = pi124  & n5001;
  assign n24090 = ~n24088 & ~n24089;
  assign n24091 = ~n24087 & n24090;
  assign n24092 = ~n24086 & n24091;
  assign n24093 = pi38  & ~n24092;
  assign n24094 = pi38  & ~n24093;
  assign n24095 = ~n24092 & ~n24093;
  assign n24096 = ~n24094 & ~n24095;
  assign n24097 = n24085 & ~n24096;
  assign n24098 = ~n24085 & n24096;
  assign n24099 = ~n24097 & ~n24098;
  assign n24100 = n23928 & n24099;
  assign n24101 = n23928 & ~n24100;
  assign n24102 = n24099 & ~n24100;
  assign n24103 = ~n24101 & ~n24102;
  assign n24104 = ~n23903 & ~n23908;
  assign n24105 = ~n24103 & ~n24104;
  assign n24106 = ~n24103 & ~n24105;
  assign n24107 = ~n24104 & ~n24105;
  assign n24108 = ~n24106 & ~n24107;
  assign n24109 = ~n23910 & ~n23913;
  assign n24110 = ~n24108 & ~n24109;
  assign n24111 = n24108 & n24109;
  assign po97  = ~n24110 & ~n24111;
  assign n24113 = ~n24105 & ~n24110;
  assign n24114 = ~n23926 & ~n24100;
  assign n24115 = ~n24084 & ~n24097;
  assign n24116 = pi127  & n4503;
  assign n24117 = n4271 & n13770;
  assign n24118 = ~n24116 & ~n24117;
  assign n24119 = pi35  & ~n24118;
  assign n24120 = pi35  & ~n24119;
  assign n24121 = ~n24118 & ~n24119;
  assign n24122 = ~n24120 & ~n24121;
  assign n24123 = ~n24115 & ~n24122;
  assign n24124 = ~n24115 & ~n24123;
  assign n24125 = ~n24122 & ~n24123;
  assign n24126 = ~n24124 & ~n24125;
  assign n24127 = ~n23833 & ~n24046;
  assign n24128 = ~n24061 & ~n24127;
  assign n24129 = n6539 & n11028;
  assign n24130 = pi118  & n6873;
  assign n24131 = pi120  & n6537;
  assign n24132 = pi119  & n6532;
  assign n24133 = ~n24131 & ~n24132;
  assign n24134 = ~n24130 & n24133;
  assign n24135 = ~n24129 & n24134;
  assign n24136 = pi44  & ~n24135;
  assign n24137 = pi44  & ~n24136;
  assign n24138 = ~n24135 & ~n24136;
  assign n24139 = ~n24137 & ~n24138;
  assign n24140 = ~n24030 & ~n24043;
  assign n24141 = n7408 & n9958;
  assign n24142 = pi115  & n7740;
  assign n24143 = pi117  & n7406;
  assign n24144 = pi116  & n7401;
  assign n24145 = ~n24143 & ~n24144;
  assign n24146 = ~n24142 & n24145;
  assign n24147 = ~n24141 & n24146;
  assign n24148 = pi47  & ~n24147;
  assign n24149 = pi47  & ~n24148;
  assign n24150 = ~n24147 & ~n24148;
  assign n24151 = ~n24149 & ~n24150;
  assign n24152 = ~n24011 & ~n24024;
  assign n24153 = ~n23972 & ~n23986;
  assign n24154 = n7060 & n10394;
  assign n24155 = pi106  & n10744;
  assign n24156 = pi108  & n10392;
  assign n24157 = pi107  & n10387;
  assign n24158 = ~n24156 & ~n24157;
  assign n24159 = ~n24155 & n24158;
  assign n24160 = ~n24154 & n24159;
  assign n24161 = pi56  & ~n24160;
  assign n24162 = pi56  & ~n24161;
  assign n24163 = ~n24160 & ~n24161;
  assign n24164 = ~n24162 & ~n24163;
  assign n24165 = ~n23965 & ~n23969;
  assign n24166 = ~n23949 & ~n23963;
  assign n24167 = pi98  & n13835;
  assign n24168 = pi99  & ~n13434;
  assign n24169 = ~n24167 & ~n24168;
  assign n24170 = ~n23946 & n24169;
  assign n24171 = n23946 & ~n24169;
  assign n24172 = ~n24170 & ~n24171;
  assign n24173 = ~n24166 & n24172;
  assign n24174 = ~n24166 & ~n24173;
  assign n24175 = ~n24170 & ~n24173;
  assign n24176 = ~n24171 & n24175;
  assign n24177 = ~n24174 & ~n24176;
  assign n24178 = n5413 & n12627;
  assign n24179 = pi100  & n13004;
  assign n24180 = pi102  & n12625;
  assign n24181 = pi101  & n12620;
  assign n24182 = ~n24180 & ~n24181;
  assign n24183 = ~n24179 & n24182;
  assign n24184 = ~n24178 & n24183;
  assign n24185 = pi62  & ~n24184;
  assign n24186 = pi62  & ~n24185;
  assign n24187 = ~n24184 & ~n24185;
  assign n24188 = ~n24186 & ~n24187;
  assign n24189 = ~n24177 & ~n24188;
  assign n24190 = ~n24177 & ~n24189;
  assign n24191 = ~n24188 & ~n24189;
  assign n24192 = ~n24190 & ~n24191;
  assign n24193 = n6207 & n11488;
  assign n24194 = pi103  & n11847;
  assign n24195 = pi105  & n11486;
  assign n24196 = pi104  & n11481;
  assign n24197 = ~n24195 & ~n24196;
  assign n24198 = ~n24194 & n24197;
  assign n24199 = ~n24193 & n24198;
  assign n24200 = pi59  & ~n24199;
  assign n24201 = pi59  & ~n24200;
  assign n24202 = ~n24199 & ~n24200;
  assign n24203 = ~n24201 & ~n24202;
  assign n24204 = ~n24192 & n24203;
  assign n24205 = n24192 & ~n24203;
  assign n24206 = ~n24204 & ~n24205;
  assign n24207 = ~n24165 & ~n24206;
  assign n24208 = n24165 & n24206;
  assign n24209 = ~n24207 & ~n24208;
  assign n24210 = ~n24164 & n24209;
  assign n24211 = n24164 & ~n24209;
  assign n24212 = ~n24210 & ~n24211;
  assign n24213 = ~n24153 & n24212;
  assign n24214 = n24153 & ~n24212;
  assign n24215 = ~n24213 & ~n24214;
  assign n24216 = n7970 & n9310;
  assign n24217 = pi109  & n9701;
  assign n24218 = pi111  & n9308;
  assign n24219 = pi110  & n9303;
  assign n24220 = ~n24218 & ~n24219;
  assign n24221 = ~n24217 & n24220;
  assign n24222 = ~n24216 & n24221;
  assign n24223 = pi53  & ~n24222;
  assign n24224 = pi53  & ~n24223;
  assign n24225 = ~n24222 & ~n24223;
  assign n24226 = ~n24224 & ~n24225;
  assign n24227 = n24215 & ~n24226;
  assign n24228 = n24215 & ~n24227;
  assign n24229 = ~n24226 & ~n24227;
  assign n24230 = ~n24228 & ~n24229;
  assign n24231 = ~n23992 & ~n24005;
  assign n24232 = n24230 & n24231;
  assign n24233 = ~n24230 & ~n24231;
  assign n24234 = ~n24232 & ~n24233;
  assign n24235 = n8334 & n8936;
  assign n24236 = pi112  & n8685;
  assign n24237 = pi114  & n8332;
  assign n24238 = pi113  & n8327;
  assign n24239 = ~n24237 & ~n24238;
  assign n24240 = ~n24236 & n24239;
  assign n24241 = ~n24235 & n24240;
  assign n24242 = pi50  & ~n24241;
  assign n24243 = pi50  & ~n24242;
  assign n24244 = ~n24241 & ~n24242;
  assign n24245 = ~n24243 & ~n24244;
  assign n24246 = ~n24234 & n24245;
  assign n24247 = n24234 & ~n24245;
  assign n24248 = ~n24246 & ~n24247;
  assign n24249 = ~n24152 & n24248;
  assign n24250 = ~n24152 & ~n24249;
  assign n24251 = n24248 & ~n24249;
  assign n24252 = ~n24250 & ~n24251;
  assign n24253 = ~n24151 & ~n24252;
  assign n24254 = n24151 & n24252;
  assign n24255 = ~n24253 & ~n24254;
  assign n24256 = ~n24140 & n24255;
  assign n24257 = n24140 & ~n24255;
  assign n24258 = ~n24256 & ~n24257;
  assign n24259 = ~n24139 & n24258;
  assign n24260 = n24139 & ~n24258;
  assign n24261 = ~n24259 & ~n24260;
  assign n24262 = ~n24128 & n24261;
  assign n24263 = n24128 & ~n24261;
  assign n24264 = ~n24262 & ~n24263;
  assign n24265 = n5739 & n12158;
  assign n24266 = pi121  & n6030;
  assign n24267 = pi123  & n5737;
  assign n24268 = pi122  & n5732;
  assign n24269 = ~n24267 & ~n24268;
  assign n24270 = ~n24266 & n24269;
  assign n24271 = ~n24265 & n24270;
  assign n24272 = pi41  & ~n24271;
  assign n24273 = pi41  & ~n24272;
  assign n24274 = ~n24271 & ~n24272;
  assign n24275 = ~n24273 & ~n24274;
  assign n24276 = n24264 & ~n24275;
  assign n24277 = n24264 & ~n24276;
  assign n24278 = ~n24275 & ~n24276;
  assign n24279 = ~n24277 & ~n24278;
  assign n24280 = ~n24064 & ~n24078;
  assign n24281 = n24279 & n24280;
  assign n24282 = ~n24279 & ~n24280;
  assign n24283 = ~n24281 & ~n24282;
  assign n24284 = n5008 & n13344;
  assign n24285 = pi124  & n5241;
  assign n24286 = pi126  & n5006;
  assign n24287 = pi125  & n5001;
  assign n24288 = ~n24286 & ~n24287;
  assign n24289 = ~n24285 & n24288;
  assign n24290 = ~n24284 & n24289;
  assign n24291 = pi38  & ~n24290;
  assign n24292 = pi38  & ~n24291;
  assign n24293 = ~n24290 & ~n24291;
  assign n24294 = ~n24292 & ~n24293;
  assign n24295 = n24283 & ~n24294;
  assign n24296 = n24283 & ~n24295;
  assign n24297 = ~n24294 & ~n24295;
  assign n24298 = ~n24296 & ~n24297;
  assign n24299 = ~n24126 & n24298;
  assign n24300 = n24126 & ~n24298;
  assign n24301 = ~n24299 & ~n24300;
  assign n24302 = ~n24114 & ~n24301;
  assign n24303 = n24114 & n24301;
  assign n24304 = ~n24302 & ~n24303;
  assign n24305 = ~n24113 & n24304;
  assign n24306 = n24113 & ~n24304;
  assign po98  = ~n24305 & ~n24306;
  assign n24308 = ~n24302 & ~n24305;
  assign n24309 = ~n24249 & ~n24253;
  assign n24310 = n7408 & n9984;
  assign n24311 = pi116  & n7740;
  assign n24312 = pi118  & n7406;
  assign n24313 = pi117  & n7401;
  assign n24314 = ~n24312 & ~n24313;
  assign n24315 = ~n24311 & n24314;
  assign n24316 = ~n24310 & n24315;
  assign n24317 = pi47  & ~n24316;
  assign n24318 = pi47  & ~n24317;
  assign n24319 = ~n24316 & ~n24317;
  assign n24320 = ~n24318 & ~n24319;
  assign n24321 = ~n24233 & ~n24247;
  assign n24322 = pi99  & n13835;
  assign n24323 = pi100  & ~n13434;
  assign n24324 = ~n24322 & ~n24323;
  assign n24325 = pi35  & ~n24169;
  assign n24326 = ~pi35  & n24169;
  assign n24327 = ~n24325 & ~n24326;
  assign n24328 = ~n24324 & ~n24327;
  assign n24329 = n24324 & n24327;
  assign n24330 = ~n24328 & ~n24329;
  assign n24331 = ~n24175 & n24330;
  assign n24332 = n24175 & ~n24330;
  assign n24333 = ~n24331 & ~n24332;
  assign n24334 = n5664 & n12627;
  assign n24335 = pi101  & n13004;
  assign n24336 = pi103  & n12625;
  assign n24337 = pi102  & n12620;
  assign n24338 = ~n24336 & ~n24337;
  assign n24339 = ~n24335 & n24338;
  assign n24340 = ~n24334 & n24339;
  assign n24341 = pi62  & ~n24340;
  assign n24342 = pi62  & ~n24341;
  assign n24343 = ~n24340 & ~n24341;
  assign n24344 = ~n24342 & ~n24343;
  assign n24345 = ~n24333 & n24344;
  assign n24346 = n24333 & ~n24344;
  assign n24347 = ~n24345 & ~n24346;
  assign n24348 = n6477 & n11488;
  assign n24349 = pi104  & n11847;
  assign n24350 = pi106  & n11486;
  assign n24351 = pi105  & n11481;
  assign n24352 = ~n24350 & ~n24351;
  assign n24353 = ~n24349 & n24352;
  assign n24354 = ~n24348 & n24353;
  assign n24355 = pi59  & ~n24354;
  assign n24356 = pi59  & ~n24355;
  assign n24357 = ~n24354 & ~n24355;
  assign n24358 = ~n24356 & ~n24357;
  assign n24359 = n24347 & ~n24358;
  assign n24360 = n24347 & ~n24359;
  assign n24361 = ~n24358 & ~n24359;
  assign n24362 = ~n24360 & ~n24361;
  assign n24363 = ~n24192 & ~n24203;
  assign n24364 = ~n24189 & ~n24363;
  assign n24365 = ~n24362 & ~n24364;
  assign n24366 = ~n24362 & ~n24365;
  assign n24367 = ~n24364 & ~n24365;
  assign n24368 = ~n24366 & ~n24367;
  assign n24369 = n7349 & n10394;
  assign n24370 = pi107  & n10744;
  assign n24371 = pi109  & n10392;
  assign n24372 = pi108  & n10387;
  assign n24373 = ~n24371 & ~n24372;
  assign n24374 = ~n24370 & n24373;
  assign n24375 = ~n24369 & n24374;
  assign n24376 = pi56  & ~n24375;
  assign n24377 = pi56  & ~n24376;
  assign n24378 = ~n24375 & ~n24376;
  assign n24379 = ~n24377 & ~n24378;
  assign n24380 = ~n24368 & ~n24379;
  assign n24381 = ~n24368 & ~n24380;
  assign n24382 = ~n24379 & ~n24380;
  assign n24383 = ~n24381 & ~n24382;
  assign n24384 = ~n24207 & ~n24210;
  assign n24385 = n24383 & n24384;
  assign n24386 = ~n24383 & ~n24384;
  assign n24387 = ~n24385 & ~n24386;
  assign n24388 = n7997 & n9310;
  assign n24389 = pi110  & n9701;
  assign n24390 = pi112  & n9308;
  assign n24391 = pi111  & n9303;
  assign n24392 = ~n24390 & ~n24391;
  assign n24393 = ~n24389 & n24392;
  assign n24394 = ~n24388 & n24393;
  assign n24395 = pi53  & ~n24394;
  assign n24396 = pi53  & ~n24395;
  assign n24397 = ~n24394 & ~n24395;
  assign n24398 = ~n24396 & ~n24397;
  assign n24399 = n24387 & ~n24398;
  assign n24400 = n24387 & ~n24399;
  assign n24401 = ~n24398 & ~n24399;
  assign n24402 = ~n24400 & ~n24401;
  assign n24403 = ~n24213 & ~n24227;
  assign n24404 = n24402 & n24403;
  assign n24405 = ~n24402 & ~n24403;
  assign n24406 = ~n24404 & ~n24405;
  assign n24407 = n8334 & n8963;
  assign n24408 = pi113  & n8685;
  assign n24409 = pi115  & n8332;
  assign n24410 = pi114  & n8327;
  assign n24411 = ~n24409 & ~n24410;
  assign n24412 = ~n24408 & n24411;
  assign n24413 = ~n24407 & n24412;
  assign n24414 = pi50  & ~n24413;
  assign n24415 = pi50  & ~n24414;
  assign n24416 = ~n24413 & ~n24414;
  assign n24417 = ~n24415 & ~n24416;
  assign n24418 = ~n24406 & n24417;
  assign n24419 = n24406 & ~n24417;
  assign n24420 = ~n24418 & ~n24419;
  assign n24421 = ~n24321 & n24420;
  assign n24422 = n24321 & ~n24420;
  assign n24423 = ~n24421 & ~n24422;
  assign n24424 = ~n24320 & n24423;
  assign n24425 = n24320 & ~n24423;
  assign n24426 = ~n24424 & ~n24425;
  assign n24427 = ~n24309 & n24426;
  assign n24428 = n24309 & ~n24426;
  assign n24429 = ~n24427 & ~n24428;
  assign n24430 = n6539 & n11389;
  assign n24431 = pi119  & n6873;
  assign n24432 = pi121  & n6537;
  assign n24433 = pi120  & n6532;
  assign n24434 = ~n24432 & ~n24433;
  assign n24435 = ~n24431 & n24434;
  assign n24436 = ~n24430 & n24435;
  assign n24437 = pi44  & ~n24436;
  assign n24438 = pi44  & ~n24437;
  assign n24439 = ~n24436 & ~n24437;
  assign n24440 = ~n24438 & ~n24439;
  assign n24441 = n24429 & ~n24440;
  assign n24442 = n24429 & ~n24441;
  assign n24443 = ~n24440 & ~n24441;
  assign n24444 = ~n24442 & ~n24443;
  assign n24445 = ~n24256 & ~n24259;
  assign n24446 = n24444 & n24445;
  assign n24447 = ~n24444 & ~n24445;
  assign n24448 = ~n24446 & ~n24447;
  assign n24449 = n5739 & n12189;
  assign n24450 = pi122  & n6030;
  assign n24451 = pi124  & n5737;
  assign n24452 = pi123  & n5732;
  assign n24453 = ~n24451 & ~n24452;
  assign n24454 = ~n24450 & n24453;
  assign n24455 = ~n24449 & n24454;
  assign n24456 = pi41  & ~n24455;
  assign n24457 = pi41  & ~n24456;
  assign n24458 = ~n24455 & ~n24456;
  assign n24459 = ~n24457 & ~n24458;
  assign n24460 = n24448 & ~n24459;
  assign n24461 = n24448 & ~n24460;
  assign n24462 = ~n24459 & ~n24460;
  assign n24463 = ~n24461 & ~n24462;
  assign n24464 = ~n24262 & ~n24276;
  assign n24465 = n24463 & n24464;
  assign n24466 = ~n24463 & ~n24464;
  assign n24467 = ~n24465 & ~n24466;
  assign n24468 = n5008 & n13742;
  assign n24469 = pi125  & n5241;
  assign n24470 = pi127  & n5006;
  assign n24471 = pi126  & n5001;
  assign n24472 = ~n24470 & ~n24471;
  assign n24473 = ~n24469 & n24472;
  assign n24474 = ~n24468 & n24473;
  assign n24475 = pi38  & ~n24474;
  assign n24476 = pi38  & ~n24475;
  assign n24477 = ~n24474 & ~n24475;
  assign n24478 = ~n24476 & ~n24477;
  assign n24479 = n24467 & ~n24478;
  assign n24480 = n24467 & ~n24479;
  assign n24481 = ~n24478 & ~n24479;
  assign n24482 = ~n24480 & ~n24481;
  assign n24483 = ~n24282 & ~n24295;
  assign n24484 = n24482 & n24483;
  assign n24485 = ~n24482 & ~n24483;
  assign n24486 = ~n24484 & ~n24485;
  assign n24487 = ~n24126 & ~n24298;
  assign n24488 = ~n24123 & ~n24487;
  assign n24489 = n24486 & ~n24488;
  assign n24490 = ~n24486 & n24488;
  assign n24491 = ~n24489 & ~n24490;
  assign n24492 = ~n24308 & n24491;
  assign n24493 = n24308 & ~n24491;
  assign po99  = ~n24492 & ~n24493;
  assign n24495 = ~n24460 & ~n24466;
  assign n24496 = pi126  & n5241;
  assign n24497 = pi127  & n5001;
  assign n24498 = ~n24496 & ~n24497;
  assign n24499 = ~n5008 & n24498;
  assign n24500 = n13773 & n24498;
  assign n24501 = ~n24499 & ~n24500;
  assign n24502 = pi38  & ~n24501;
  assign n24503 = ~pi38  & n24501;
  assign n24504 = ~n24502 & ~n24503;
  assign n24505 = ~n24495 & ~n24504;
  assign n24506 = n24495 & n24504;
  assign n24507 = ~n24505 & ~n24506;
  assign n24508 = n5943 & n12627;
  assign n24509 = pi102  & n13004;
  assign n24510 = pi104  & n12625;
  assign n24511 = pi103  & n12620;
  assign n24512 = ~n24510 & ~n24511;
  assign n24513 = ~n24509 & n24512;
  assign n24514 = ~n24508 & n24513;
  assign n24515 = pi62  & ~n24514;
  assign n24516 = pi62  & ~n24515;
  assign n24517 = ~n24514 & ~n24515;
  assign n24518 = ~n24516 & ~n24517;
  assign n24519 = pi100  & n13835;
  assign n24520 = pi101  & ~n13434;
  assign n24521 = ~n24519 & ~n24520;
  assign n24522 = ~pi35  & ~n24169;
  assign n24523 = ~n24328 & ~n24522;
  assign n24524 = n24521 & ~n24523;
  assign n24525 = n24521 & ~n24524;
  assign n24526 = ~n24523 & ~n24524;
  assign n24527 = ~n24525 & ~n24526;
  assign n24528 = ~n24518 & ~n24527;
  assign n24529 = ~n24518 & ~n24528;
  assign n24530 = ~n24527 & ~n24528;
  assign n24531 = ~n24529 & ~n24530;
  assign n24532 = ~n24331 & ~n24346;
  assign n24533 = n24531 & n24532;
  assign n24534 = ~n24531 & ~n24532;
  assign n24535 = ~n24533 & ~n24534;
  assign n24536 = n6775 & n11488;
  assign n24537 = pi105  & n11847;
  assign n24538 = pi107  & n11486;
  assign n24539 = pi106  & n11481;
  assign n24540 = ~n24538 & ~n24539;
  assign n24541 = ~n24537 & n24540;
  assign n24542 = ~n24536 & n24541;
  assign n24543 = pi59  & ~n24542;
  assign n24544 = pi59  & ~n24543;
  assign n24545 = ~n24542 & ~n24543;
  assign n24546 = ~n24544 & ~n24545;
  assign n24547 = n24535 & ~n24546;
  assign n24548 = n24535 & ~n24547;
  assign n24549 = ~n24546 & ~n24547;
  assign n24550 = ~n24548 & ~n24549;
  assign n24551 = ~n24359 & ~n24365;
  assign n24552 = n24550 & n24551;
  assign n24553 = ~n24550 & ~n24551;
  assign n24554 = ~n24552 & ~n24553;
  assign n24555 = n7665 & n10394;
  assign n24556 = pi108  & n10744;
  assign n24557 = pi110  & n10392;
  assign n24558 = pi109  & n10387;
  assign n24559 = ~n24557 & ~n24558;
  assign n24560 = ~n24556 & n24559;
  assign n24561 = ~n24555 & n24560;
  assign n24562 = pi56  & ~n24561;
  assign n24563 = pi56  & ~n24562;
  assign n24564 = ~n24561 & ~n24562;
  assign n24565 = ~n24563 & ~n24564;
  assign n24566 = n24554 & ~n24565;
  assign n24567 = n24554 & ~n24566;
  assign n24568 = ~n24565 & ~n24566;
  assign n24569 = ~n24567 & ~n24568;
  assign n24570 = ~n24380 & ~n24386;
  assign n24571 = n24569 & n24570;
  assign n24572 = ~n24569 & ~n24570;
  assign n24573 = ~n24571 & ~n24572;
  assign n24574 = n8612 & n9310;
  assign n24575 = pi111  & n9701;
  assign n24576 = pi113  & n9308;
  assign n24577 = pi112  & n9303;
  assign n24578 = ~n24576 & ~n24577;
  assign n24579 = ~n24575 & n24578;
  assign n24580 = ~n24574 & n24579;
  assign n24581 = pi53  & ~n24580;
  assign n24582 = pi53  & ~n24581;
  assign n24583 = ~n24580 & ~n24581;
  assign n24584 = ~n24582 & ~n24583;
  assign n24585 = n24573 & ~n24584;
  assign n24586 = n24573 & ~n24585;
  assign n24587 = ~n24584 & ~n24585;
  assign n24588 = ~n24586 & ~n24587;
  assign n24589 = ~n24399 & ~n24405;
  assign n24590 = n24588 & n24589;
  assign n24591 = ~n24588 & ~n24589;
  assign n24592 = ~n24590 & ~n24591;
  assign n24593 = n8334 & n9614;
  assign n24594 = pi114  & n8685;
  assign n24595 = pi116  & n8332;
  assign n24596 = pi115  & n8327;
  assign n24597 = ~n24595 & ~n24596;
  assign n24598 = ~n24594 & n24597;
  assign n24599 = ~n24593 & n24598;
  assign n24600 = pi50  & ~n24599;
  assign n24601 = pi50  & ~n24600;
  assign n24602 = ~n24599 & ~n24600;
  assign n24603 = ~n24601 & ~n24602;
  assign n24604 = n24592 & ~n24603;
  assign n24605 = n24592 & ~n24604;
  assign n24606 = ~n24603 & ~n24604;
  assign n24607 = ~n24605 & ~n24606;
  assign n24608 = ~n24419 & ~n24421;
  assign n24609 = ~n24607 & ~n24608;
  assign n24610 = ~n24607 & ~n24609;
  assign n24611 = ~n24608 & ~n24609;
  assign n24612 = ~n24610 & ~n24611;
  assign n24613 = n7408 & n10667;
  assign n24614 = pi117  & n7740;
  assign n24615 = pi119  & n7406;
  assign n24616 = pi118  & n7401;
  assign n24617 = ~n24615 & ~n24616;
  assign n24618 = ~n24614 & n24617;
  assign n24619 = ~n24613 & n24618;
  assign n24620 = pi47  & ~n24619;
  assign n24621 = pi47  & ~n24620;
  assign n24622 = ~n24619 & ~n24620;
  assign n24623 = ~n24621 & ~n24622;
  assign n24624 = ~n24612 & ~n24623;
  assign n24625 = ~n24612 & ~n24624;
  assign n24626 = ~n24623 & ~n24624;
  assign n24627 = ~n24625 & ~n24626;
  assign n24628 = ~n24424 & ~n24427;
  assign n24629 = n24627 & n24628;
  assign n24630 = ~n24627 & ~n24628;
  assign n24631 = ~n24629 & ~n24630;
  assign n24632 = n6539 & n11778;
  assign n24633 = pi120  & n6873;
  assign n24634 = pi122  & n6537;
  assign n24635 = pi121  & n6532;
  assign n24636 = ~n24634 & ~n24635;
  assign n24637 = ~n24633 & n24636;
  assign n24638 = ~n24632 & n24637;
  assign n24639 = pi44  & ~n24638;
  assign n24640 = pi44  & ~n24639;
  assign n24641 = ~n24638 & ~n24639;
  assign n24642 = ~n24640 & ~n24641;
  assign n24643 = n24631 & ~n24642;
  assign n24644 = n24631 & ~n24643;
  assign n24645 = ~n24642 & ~n24643;
  assign n24646 = ~n24644 & ~n24645;
  assign n24647 = ~n24441 & ~n24447;
  assign n24648 = n24646 & n24647;
  assign n24649 = ~n24646 & ~n24647;
  assign n24650 = ~n24648 & ~n24649;
  assign n24651 = n5739 & n12943;
  assign n24652 = pi123  & n6030;
  assign n24653 = pi125  & n5737;
  assign n24654 = pi124  & n5732;
  assign n24655 = ~n24653 & ~n24654;
  assign n24656 = ~n24652 & n24655;
  assign n24657 = ~n24651 & n24656;
  assign n24658 = pi41  & ~n24657;
  assign n24659 = pi41  & ~n24658;
  assign n24660 = ~n24657 & ~n24658;
  assign n24661 = ~n24659 & ~n24660;
  assign n24662 = n24650 & ~n24661;
  assign n24663 = ~n24650 & n24661;
  assign n24664 = ~n24662 & ~n24663;
  assign n24665 = n24507 & n24664;
  assign n24666 = n24507 & ~n24665;
  assign n24667 = n24664 & ~n24665;
  assign n24668 = ~n24666 & ~n24667;
  assign n24669 = ~n24479 & ~n24485;
  assign n24670 = n24668 & n24669;
  assign n24671 = ~n24668 & ~n24669;
  assign n24672 = ~n24670 & ~n24671;
  assign n24673 = ~n24489 & ~n24492;
  assign n24674 = n24672 & ~n24673;
  assign n24675 = ~n24672 & n24673;
  assign po100  = ~n24674 & ~n24675;
  assign n24677 = ~n24671 & ~n24674;
  assign n24678 = ~n24505 & ~n24665;
  assign n24679 = ~n24649 & ~n24662;
  assign n24680 = pi127  & n5241;
  assign n24681 = n5008 & n13770;
  assign n24682 = ~n24680 & ~n24681;
  assign n24683 = pi38  & ~n24682;
  assign n24684 = pi38  & ~n24683;
  assign n24685 = ~n24682 & ~n24683;
  assign n24686 = ~n24684 & ~n24685;
  assign n24687 = ~n24679 & ~n24686;
  assign n24688 = ~n24679 & ~n24687;
  assign n24689 = ~n24686 & ~n24687;
  assign n24690 = ~n24688 & ~n24689;
  assign n24691 = ~n24609 & ~n24624;
  assign n24692 = n7408 & n11028;
  assign n24693 = pi118  & n7740;
  assign n24694 = pi120  & n7406;
  assign n24695 = pi119  & n7401;
  assign n24696 = ~n24694 & ~n24695;
  assign n24697 = ~n24693 & n24696;
  assign n24698 = ~n24692 & n24697;
  assign n24699 = pi47  & ~n24698;
  assign n24700 = pi47  & ~n24699;
  assign n24701 = ~n24698 & ~n24699;
  assign n24702 = ~n24700 & ~n24701;
  assign n24703 = ~n24591 & ~n24604;
  assign n24704 = n8334 & n9958;
  assign n24705 = pi115  & n8685;
  assign n24706 = pi117  & n8332;
  assign n24707 = pi116  & n8327;
  assign n24708 = ~n24706 & ~n24707;
  assign n24709 = ~n24705 & n24708;
  assign n24710 = ~n24704 & n24709;
  assign n24711 = pi50  & ~n24710;
  assign n24712 = pi50  & ~n24711;
  assign n24713 = ~n24710 & ~n24711;
  assign n24714 = ~n24712 & ~n24713;
  assign n24715 = ~n24572 & ~n24585;
  assign n24716 = ~n24524 & ~n24528;
  assign n24717 = pi101  & n13835;
  assign n24718 = pi102  & ~n13434;
  assign n24719 = ~n24717 & ~n24718;
  assign n24720 = n24521 & ~n24719;
  assign n24721 = n24521 & ~n24720;
  assign n24722 = ~n24719 & ~n24720;
  assign n24723 = ~n24721 & ~n24722;
  assign n24724 = ~n24716 & ~n24723;
  assign n24725 = ~n24716 & ~n24724;
  assign n24726 = ~n24723 & ~n24724;
  assign n24727 = ~n24725 & ~n24726;
  assign n24728 = n6207 & n12627;
  assign n24729 = pi103  & n13004;
  assign n24730 = pi105  & n12625;
  assign n24731 = pi104  & n12620;
  assign n24732 = ~n24730 & ~n24731;
  assign n24733 = ~n24729 & n24732;
  assign n24734 = ~n24728 & n24733;
  assign n24735 = pi62  & ~n24734;
  assign n24736 = pi62  & ~n24735;
  assign n24737 = ~n24734 & ~n24735;
  assign n24738 = ~n24736 & ~n24737;
  assign n24739 = ~n24727 & ~n24738;
  assign n24740 = ~n24727 & ~n24739;
  assign n24741 = ~n24738 & ~n24739;
  assign n24742 = ~n24740 & ~n24741;
  assign n24743 = n7060 & n11488;
  assign n24744 = pi106  & n11847;
  assign n24745 = pi108  & n11486;
  assign n24746 = pi107  & n11481;
  assign n24747 = ~n24745 & ~n24746;
  assign n24748 = ~n24744 & n24747;
  assign n24749 = ~n24743 & n24748;
  assign n24750 = pi59  & ~n24749;
  assign n24751 = pi59  & ~n24750;
  assign n24752 = ~n24749 & ~n24750;
  assign n24753 = ~n24751 & ~n24752;
  assign n24754 = ~n24742 & n24753;
  assign n24755 = n24742 & ~n24753;
  assign n24756 = ~n24754 & ~n24755;
  assign n24757 = ~n24534 & ~n24547;
  assign n24758 = n24756 & n24757;
  assign n24759 = ~n24756 & ~n24757;
  assign n24760 = ~n24758 & ~n24759;
  assign n24761 = n7970 & n10394;
  assign n24762 = pi109  & n10744;
  assign n24763 = pi111  & n10392;
  assign n24764 = pi110  & n10387;
  assign n24765 = ~n24763 & ~n24764;
  assign n24766 = ~n24762 & n24765;
  assign n24767 = ~n24761 & n24766;
  assign n24768 = pi56  & ~n24767;
  assign n24769 = pi56  & ~n24768;
  assign n24770 = ~n24767 & ~n24768;
  assign n24771 = ~n24769 & ~n24770;
  assign n24772 = n24760 & ~n24771;
  assign n24773 = n24760 & ~n24772;
  assign n24774 = ~n24771 & ~n24772;
  assign n24775 = ~n24773 & ~n24774;
  assign n24776 = ~n24553 & ~n24566;
  assign n24777 = n24775 & n24776;
  assign n24778 = ~n24775 & ~n24776;
  assign n24779 = ~n24777 & ~n24778;
  assign n24780 = n8936 & n9310;
  assign n24781 = pi112  & n9701;
  assign n24782 = pi114  & n9308;
  assign n24783 = pi113  & n9303;
  assign n24784 = ~n24782 & ~n24783;
  assign n24785 = ~n24781 & n24784;
  assign n24786 = ~n24780 & n24785;
  assign n24787 = pi53  & ~n24786;
  assign n24788 = pi53  & ~n24787;
  assign n24789 = ~n24786 & ~n24787;
  assign n24790 = ~n24788 & ~n24789;
  assign n24791 = ~n24779 & n24790;
  assign n24792 = n24779 & ~n24790;
  assign n24793 = ~n24791 & ~n24792;
  assign n24794 = ~n24715 & n24793;
  assign n24795 = ~n24715 & ~n24794;
  assign n24796 = n24793 & ~n24794;
  assign n24797 = ~n24795 & ~n24796;
  assign n24798 = ~n24714 & ~n24797;
  assign n24799 = n24714 & n24797;
  assign n24800 = ~n24798 & ~n24799;
  assign n24801 = ~n24703 & n24800;
  assign n24802 = n24703 & ~n24800;
  assign n24803 = ~n24801 & ~n24802;
  assign n24804 = ~n24702 & n24803;
  assign n24805 = n24702 & ~n24803;
  assign n24806 = ~n24804 & ~n24805;
  assign n24807 = ~n24691 & n24806;
  assign n24808 = n24691 & ~n24806;
  assign n24809 = ~n24807 & ~n24808;
  assign n24810 = n6539 & n12158;
  assign n24811 = pi121  & n6873;
  assign n24812 = pi123  & n6537;
  assign n24813 = pi122  & n6532;
  assign n24814 = ~n24812 & ~n24813;
  assign n24815 = ~n24811 & n24814;
  assign n24816 = ~n24810 & n24815;
  assign n24817 = pi44  & ~n24816;
  assign n24818 = pi44  & ~n24817;
  assign n24819 = ~n24816 & ~n24817;
  assign n24820 = ~n24818 & ~n24819;
  assign n24821 = n24809 & ~n24820;
  assign n24822 = n24809 & ~n24821;
  assign n24823 = ~n24820 & ~n24821;
  assign n24824 = ~n24822 & ~n24823;
  assign n24825 = ~n24630 & ~n24643;
  assign n24826 = n24824 & n24825;
  assign n24827 = ~n24824 & ~n24825;
  assign n24828 = ~n24826 & ~n24827;
  assign n24829 = n5739 & n13344;
  assign n24830 = pi124  & n6030;
  assign n24831 = pi126  & n5737;
  assign n24832 = pi125  & n5732;
  assign n24833 = ~n24831 & ~n24832;
  assign n24834 = ~n24830 & n24833;
  assign n24835 = ~n24829 & n24834;
  assign n24836 = pi41  & ~n24835;
  assign n24837 = pi41  & ~n24836;
  assign n24838 = ~n24835 & ~n24836;
  assign n24839 = ~n24837 & ~n24838;
  assign n24840 = n24828 & ~n24839;
  assign n24841 = n24828 & ~n24840;
  assign n24842 = ~n24839 & ~n24840;
  assign n24843 = ~n24841 & ~n24842;
  assign n24844 = ~n24690 & n24843;
  assign n24845 = n24690 & ~n24843;
  assign n24846 = ~n24844 & ~n24845;
  assign n24847 = ~n24678 & ~n24846;
  assign n24848 = n24678 & n24846;
  assign n24849 = ~n24847 & ~n24848;
  assign n24850 = ~n24677 & n24849;
  assign n24851 = n24677 & ~n24849;
  assign po101  = ~n24850 & ~n24851;
  assign n24853 = ~n24847 & ~n24850;
  assign n24854 = ~n24794 & ~n24798;
  assign n24855 = n8334 & n9984;
  assign n24856 = pi116  & n8685;
  assign n24857 = pi118  & n8332;
  assign n24858 = pi117  & n8327;
  assign n24859 = ~n24857 & ~n24858;
  assign n24860 = ~n24856 & n24859;
  assign n24861 = ~n24855 & n24860;
  assign n24862 = pi50  & ~n24861;
  assign n24863 = pi50  & ~n24862;
  assign n24864 = ~n24861 & ~n24862;
  assign n24865 = ~n24863 & ~n24864;
  assign n24866 = ~n24778 & ~n24792;
  assign n24867 = ~n24720 & ~n24724;
  assign n24868 = pi102  & n13835;
  assign n24869 = pi103  & ~n13434;
  assign n24870 = ~n24868 & ~n24869;
  assign n24871 = pi38  & ~n24521;
  assign n24872 = ~pi38  & n24521;
  assign n24873 = ~n24871 & ~n24872;
  assign n24874 = ~n24870 & ~n24873;
  assign n24875 = n24870 & n24873;
  assign n24876 = ~n24874 & ~n24875;
  assign n24877 = ~n24867 & n24876;
  assign n24878 = n24867 & ~n24876;
  assign n24879 = ~n24877 & ~n24878;
  assign n24880 = n6477 & n12627;
  assign n24881 = pi104  & n13004;
  assign n24882 = pi106  & n12625;
  assign n24883 = pi105  & n12620;
  assign n24884 = ~n24882 & ~n24883;
  assign n24885 = ~n24881 & n24884;
  assign n24886 = ~n24880 & n24885;
  assign n24887 = pi62  & ~n24886;
  assign n24888 = pi62  & ~n24887;
  assign n24889 = ~n24886 & ~n24887;
  assign n24890 = ~n24888 & ~n24889;
  assign n24891 = n24879 & ~n24890;
  assign n24892 = n24879 & ~n24891;
  assign n24893 = ~n24890 & ~n24891;
  assign n24894 = ~n24892 & ~n24893;
  assign n24895 = n7349 & n11488;
  assign n24896 = pi107  & n11847;
  assign n24897 = pi109  & n11486;
  assign n24898 = pi108  & n11481;
  assign n24899 = ~n24897 & ~n24898;
  assign n24900 = ~n24896 & n24899;
  assign n24901 = ~n24895 & n24900;
  assign n24902 = pi59  & ~n24901;
  assign n24903 = pi59  & ~n24902;
  assign n24904 = ~n24901 & ~n24902;
  assign n24905 = ~n24903 & ~n24904;
  assign n24906 = ~n24894 & ~n24905;
  assign n24907 = ~n24894 & ~n24906;
  assign n24908 = ~n24905 & ~n24906;
  assign n24909 = ~n24907 & ~n24908;
  assign n24910 = ~n24742 & ~n24753;
  assign n24911 = ~n24739 & ~n24910;
  assign n24912 = ~n24909 & ~n24911;
  assign n24913 = ~n24909 & ~n24912;
  assign n24914 = ~n24911 & ~n24912;
  assign n24915 = ~n24913 & ~n24914;
  assign n24916 = n7997 & n10394;
  assign n24917 = pi110  & n10744;
  assign n24918 = pi112  & n10392;
  assign n24919 = pi111  & n10387;
  assign n24920 = ~n24918 & ~n24919;
  assign n24921 = ~n24917 & n24920;
  assign n24922 = ~n24916 & n24921;
  assign n24923 = pi56  & ~n24922;
  assign n24924 = pi56  & ~n24923;
  assign n24925 = ~n24922 & ~n24923;
  assign n24926 = ~n24924 & ~n24925;
  assign n24927 = ~n24915 & ~n24926;
  assign n24928 = ~n24915 & ~n24927;
  assign n24929 = ~n24926 & ~n24927;
  assign n24930 = ~n24928 & ~n24929;
  assign n24931 = ~n24759 & ~n24772;
  assign n24932 = n24930 & n24931;
  assign n24933 = ~n24930 & ~n24931;
  assign n24934 = ~n24932 & ~n24933;
  assign n24935 = n8963 & n9310;
  assign n24936 = pi113  & n9701;
  assign n24937 = pi115  & n9308;
  assign n24938 = pi114  & n9303;
  assign n24939 = ~n24937 & ~n24938;
  assign n24940 = ~n24936 & n24939;
  assign n24941 = ~n24935 & n24940;
  assign n24942 = pi53  & ~n24941;
  assign n24943 = pi53  & ~n24942;
  assign n24944 = ~n24941 & ~n24942;
  assign n24945 = ~n24943 & ~n24944;
  assign n24946 = ~n24934 & n24945;
  assign n24947 = n24934 & ~n24945;
  assign n24948 = ~n24946 & ~n24947;
  assign n24949 = ~n24866 & n24948;
  assign n24950 = n24866 & ~n24948;
  assign n24951 = ~n24949 & ~n24950;
  assign n24952 = ~n24865 & n24951;
  assign n24953 = n24865 & ~n24951;
  assign n24954 = ~n24952 & ~n24953;
  assign n24955 = ~n24854 & n24954;
  assign n24956 = n24854 & ~n24954;
  assign n24957 = ~n24955 & ~n24956;
  assign n24958 = n7408 & n11389;
  assign n24959 = pi119  & n7740;
  assign n24960 = pi121  & n7406;
  assign n24961 = pi120  & n7401;
  assign n24962 = ~n24960 & ~n24961;
  assign n24963 = ~n24959 & n24962;
  assign n24964 = ~n24958 & n24963;
  assign n24965 = pi47  & ~n24964;
  assign n24966 = pi47  & ~n24965;
  assign n24967 = ~n24964 & ~n24965;
  assign n24968 = ~n24966 & ~n24967;
  assign n24969 = n24957 & ~n24968;
  assign n24970 = n24957 & ~n24969;
  assign n24971 = ~n24968 & ~n24969;
  assign n24972 = ~n24970 & ~n24971;
  assign n24973 = ~n24801 & ~n24804;
  assign n24974 = n24972 & n24973;
  assign n24975 = ~n24972 & ~n24973;
  assign n24976 = ~n24974 & ~n24975;
  assign n24977 = n6539 & n12189;
  assign n24978 = pi122  & n6873;
  assign n24979 = pi124  & n6537;
  assign n24980 = pi123  & n6532;
  assign n24981 = ~n24979 & ~n24980;
  assign n24982 = ~n24978 & n24981;
  assign n24983 = ~n24977 & n24982;
  assign n24984 = pi44  & ~n24983;
  assign n24985 = pi44  & ~n24984;
  assign n24986 = ~n24983 & ~n24984;
  assign n24987 = ~n24985 & ~n24986;
  assign n24988 = n24976 & ~n24987;
  assign n24989 = n24976 & ~n24988;
  assign n24990 = ~n24987 & ~n24988;
  assign n24991 = ~n24989 & ~n24990;
  assign n24992 = ~n24807 & ~n24821;
  assign n24993 = n24991 & n24992;
  assign n24994 = ~n24991 & ~n24992;
  assign n24995 = ~n24993 & ~n24994;
  assign n24996 = n5739 & n13742;
  assign n24997 = pi125  & n6030;
  assign n24998 = pi127  & n5737;
  assign n24999 = pi126  & n5732;
  assign n25000 = ~n24998 & ~n24999;
  assign n25001 = ~n24997 & n25000;
  assign n25002 = ~n24996 & n25001;
  assign n25003 = pi41  & ~n25002;
  assign n25004 = pi41  & ~n25003;
  assign n25005 = ~n25002 & ~n25003;
  assign n25006 = ~n25004 & ~n25005;
  assign n25007 = n24995 & ~n25006;
  assign n25008 = n24995 & ~n25007;
  assign n25009 = ~n25006 & ~n25007;
  assign n25010 = ~n25008 & ~n25009;
  assign n25011 = ~n24827 & ~n24840;
  assign n25012 = n25010 & n25011;
  assign n25013 = ~n25010 & ~n25011;
  assign n25014 = ~n25012 & ~n25013;
  assign n25015 = ~n24690 & ~n24843;
  assign n25016 = ~n24687 & ~n25015;
  assign n25017 = n25014 & ~n25016;
  assign n25018 = ~n25014 & n25016;
  assign n25019 = ~n25017 & ~n25018;
  assign n25020 = ~n24853 & n25019;
  assign n25021 = n24853 & ~n25019;
  assign po102  = ~n25020 & ~n25021;
  assign n25023 = ~n24988 & ~n24994;
  assign n25024 = pi126  & n6030;
  assign n25025 = pi127  & n5732;
  assign n25026 = ~n25024 & ~n25025;
  assign n25027 = ~n5739 & n25026;
  assign n25028 = n13773 & n25026;
  assign n25029 = ~n25027 & ~n25028;
  assign n25030 = pi41  & ~n25029;
  assign n25031 = ~pi41  & n25029;
  assign n25032 = ~n25030 & ~n25031;
  assign n25033 = ~n25023 & ~n25032;
  assign n25034 = n25023 & n25032;
  assign n25035 = ~n25033 & ~n25034;
  assign n25036 = ~n24877 & ~n24891;
  assign n25037 = pi103  & n13835;
  assign n25038 = pi104  & ~n13434;
  assign n25039 = ~n25037 & ~n25038;
  assign n25040 = ~pi38  & ~n24521;
  assign n25041 = ~n24874 & ~n25040;
  assign n25042 = n25039 & ~n25041;
  assign n25043 = ~n25039 & n25041;
  assign n25044 = ~n25042 & ~n25043;
  assign n25045 = pi105  & n13004;
  assign n25046 = pi107  & n12625;
  assign n25047 = pi106  & n12620;
  assign n25048 = ~n25046 & ~n25047;
  assign n25049 = ~n25045 & n25048;
  assign n25050 = ~n12627 & n25049;
  assign n25051 = ~n6775 & n25049;
  assign n25052 = ~n25050 & ~n25051;
  assign n25053 = pi62  & ~n25052;
  assign n25054 = ~pi62  & n25052;
  assign n25055 = ~n25053 & ~n25054;
  assign n25056 = n25044 & ~n25055;
  assign n25057 = ~n25044 & n25055;
  assign n25058 = ~n25056 & ~n25057;
  assign n25059 = ~n25036 & n25058;
  assign n25060 = n25036 & ~n25058;
  assign n25061 = ~n25059 & ~n25060;
  assign n25062 = n7665 & n11488;
  assign n25063 = pi108  & n11847;
  assign n25064 = pi110  & n11486;
  assign n25065 = pi109  & n11481;
  assign n25066 = ~n25064 & ~n25065;
  assign n25067 = ~n25063 & n25066;
  assign n25068 = ~n25062 & n25067;
  assign n25069 = pi59  & ~n25068;
  assign n25070 = pi59  & ~n25069;
  assign n25071 = ~n25068 & ~n25069;
  assign n25072 = ~n25070 & ~n25071;
  assign n25073 = n25061 & ~n25072;
  assign n25074 = n25061 & ~n25073;
  assign n25075 = ~n25072 & ~n25073;
  assign n25076 = ~n25074 & ~n25075;
  assign n25077 = ~n24906 & ~n24912;
  assign n25078 = n25076 & n25077;
  assign n25079 = ~n25076 & ~n25077;
  assign n25080 = ~n25078 & ~n25079;
  assign n25081 = n8612 & n10394;
  assign n25082 = pi111  & n10744;
  assign n25083 = pi113  & n10392;
  assign n25084 = pi112  & n10387;
  assign n25085 = ~n25083 & ~n25084;
  assign n25086 = ~n25082 & n25085;
  assign n25087 = ~n25081 & n25086;
  assign n25088 = pi56  & ~n25087;
  assign n25089 = pi56  & ~n25088;
  assign n25090 = ~n25087 & ~n25088;
  assign n25091 = ~n25089 & ~n25090;
  assign n25092 = n25080 & ~n25091;
  assign n25093 = n25080 & ~n25092;
  assign n25094 = ~n25091 & ~n25092;
  assign n25095 = ~n25093 & ~n25094;
  assign n25096 = ~n24927 & ~n24933;
  assign n25097 = n25095 & n25096;
  assign n25098 = ~n25095 & ~n25096;
  assign n25099 = ~n25097 & ~n25098;
  assign n25100 = n9310 & n9614;
  assign n25101 = pi114  & n9701;
  assign n25102 = pi116  & n9308;
  assign n25103 = pi115  & n9303;
  assign n25104 = ~n25102 & ~n25103;
  assign n25105 = ~n25101 & n25104;
  assign n25106 = ~n25100 & n25105;
  assign n25107 = pi53  & ~n25106;
  assign n25108 = pi53  & ~n25107;
  assign n25109 = ~n25106 & ~n25107;
  assign n25110 = ~n25108 & ~n25109;
  assign n25111 = n25099 & ~n25110;
  assign n25112 = n25099 & ~n25111;
  assign n25113 = ~n25110 & ~n25111;
  assign n25114 = ~n25112 & ~n25113;
  assign n25115 = ~n24947 & ~n24949;
  assign n25116 = ~n25114 & ~n25115;
  assign n25117 = ~n25114 & ~n25116;
  assign n25118 = ~n25115 & ~n25116;
  assign n25119 = ~n25117 & ~n25118;
  assign n25120 = n8334 & n10667;
  assign n25121 = pi117  & n8685;
  assign n25122 = pi119  & n8332;
  assign n25123 = pi118  & n8327;
  assign n25124 = ~n25122 & ~n25123;
  assign n25125 = ~n25121 & n25124;
  assign n25126 = ~n25120 & n25125;
  assign n25127 = pi50  & ~n25126;
  assign n25128 = pi50  & ~n25127;
  assign n25129 = ~n25126 & ~n25127;
  assign n25130 = ~n25128 & ~n25129;
  assign n25131 = ~n25119 & ~n25130;
  assign n25132 = ~n25119 & ~n25131;
  assign n25133 = ~n25130 & ~n25131;
  assign n25134 = ~n25132 & ~n25133;
  assign n25135 = ~n24952 & ~n24955;
  assign n25136 = n25134 & n25135;
  assign n25137 = ~n25134 & ~n25135;
  assign n25138 = ~n25136 & ~n25137;
  assign n25139 = n7408 & n11778;
  assign n25140 = pi120  & n7740;
  assign n25141 = pi122  & n7406;
  assign n25142 = pi121  & n7401;
  assign n25143 = ~n25141 & ~n25142;
  assign n25144 = ~n25140 & n25143;
  assign n25145 = ~n25139 & n25144;
  assign n25146 = pi47  & ~n25145;
  assign n25147 = pi47  & ~n25146;
  assign n25148 = ~n25145 & ~n25146;
  assign n25149 = ~n25147 & ~n25148;
  assign n25150 = n25138 & ~n25149;
  assign n25151 = n25138 & ~n25150;
  assign n25152 = ~n25149 & ~n25150;
  assign n25153 = ~n25151 & ~n25152;
  assign n25154 = ~n24969 & ~n24975;
  assign n25155 = n25153 & n25154;
  assign n25156 = ~n25153 & ~n25154;
  assign n25157 = ~n25155 & ~n25156;
  assign n25158 = n6539 & n12943;
  assign n25159 = pi123  & n6873;
  assign n25160 = pi125  & n6537;
  assign n25161 = pi124  & n6532;
  assign n25162 = ~n25160 & ~n25161;
  assign n25163 = ~n25159 & n25162;
  assign n25164 = ~n25158 & n25163;
  assign n25165 = pi44  & ~n25164;
  assign n25166 = pi44  & ~n25165;
  assign n25167 = ~n25164 & ~n25165;
  assign n25168 = ~n25166 & ~n25167;
  assign n25169 = n25157 & ~n25168;
  assign n25170 = ~n25157 & n25168;
  assign n25171 = ~n25169 & ~n25170;
  assign n25172 = n25035 & n25171;
  assign n25173 = n25035 & ~n25172;
  assign n25174 = n25171 & ~n25172;
  assign n25175 = ~n25173 & ~n25174;
  assign n25176 = ~n25007 & ~n25013;
  assign n25177 = n25175 & n25176;
  assign n25178 = ~n25175 & ~n25176;
  assign n25179 = ~n25177 & ~n25178;
  assign n25180 = ~n25017 & ~n25020;
  assign n25181 = n25179 & ~n25180;
  assign n25182 = ~n25179 & n25180;
  assign po103  = ~n25181 & ~n25182;
  assign n25184 = ~n25178 & ~n25181;
  assign n25185 = ~n25033 & ~n25172;
  assign n25186 = ~n25156 & ~n25169;
  assign n25187 = pi127  & n6030;
  assign n25188 = n5739 & n13770;
  assign n25189 = ~n25187 & ~n25188;
  assign n25190 = pi41  & ~n25189;
  assign n25191 = pi41  & ~n25190;
  assign n25192 = ~n25189 & ~n25190;
  assign n25193 = ~n25191 & ~n25192;
  assign n25194 = ~n25186 & ~n25193;
  assign n25195 = ~n25186 & ~n25194;
  assign n25196 = ~n25193 & ~n25194;
  assign n25197 = ~n25195 & ~n25196;
  assign n25198 = ~n25116 & ~n25131;
  assign n25199 = n8334 & n11028;
  assign n25200 = pi118  & n8685;
  assign n25201 = pi120  & n8332;
  assign n25202 = pi119  & n8327;
  assign n25203 = ~n25201 & ~n25202;
  assign n25204 = ~n25200 & n25203;
  assign n25205 = ~n25199 & n25204;
  assign n25206 = pi50  & ~n25205;
  assign n25207 = pi50  & ~n25206;
  assign n25208 = ~n25205 & ~n25206;
  assign n25209 = ~n25207 & ~n25208;
  assign n25210 = ~n25098 & ~n25111;
  assign n25211 = n9310 & n9958;
  assign n25212 = pi115  & n9701;
  assign n25213 = pi117  & n9308;
  assign n25214 = pi116  & n9303;
  assign n25215 = ~n25213 & ~n25214;
  assign n25216 = ~n25212 & n25215;
  assign n25217 = ~n25211 & n25216;
  assign n25218 = pi53  & ~n25217;
  assign n25219 = pi53  & ~n25218;
  assign n25220 = ~n25217 & ~n25218;
  assign n25221 = ~n25219 & ~n25220;
  assign n25222 = ~n25079 & ~n25092;
  assign n25223 = ~n25059 & ~n25073;
  assign n25224 = ~n25042 & ~n25056;
  assign n25225 = pi104  & n13835;
  assign n25226 = pi105  & ~n13434;
  assign n25227 = ~n25225 & ~n25226;
  assign n25228 = n25039 & ~n25227;
  assign n25229 = n25039 & ~n25228;
  assign n25230 = ~n25227 & ~n25228;
  assign n25231 = ~n25229 & ~n25230;
  assign n25232 = ~n25224 & ~n25231;
  assign n25233 = ~n25224 & ~n25232;
  assign n25234 = ~n25231 & ~n25232;
  assign n25235 = ~n25233 & ~n25234;
  assign n25236 = n7060 & n12627;
  assign n25237 = pi106  & n13004;
  assign n25238 = pi108  & n12625;
  assign n25239 = pi107  & n12620;
  assign n25240 = ~n25238 & ~n25239;
  assign n25241 = ~n25237 & n25240;
  assign n25242 = ~n25236 & n25241;
  assign n25243 = pi62  & ~n25242;
  assign n25244 = pi62  & ~n25243;
  assign n25245 = ~n25242 & ~n25243;
  assign n25246 = ~n25244 & ~n25245;
  assign n25247 = ~n25235 & n25246;
  assign n25248 = n25235 & ~n25246;
  assign n25249 = ~n25247 & ~n25248;
  assign n25250 = n7970 & n11488;
  assign n25251 = pi109  & n11847;
  assign n25252 = pi111  & n11486;
  assign n25253 = pi110  & n11481;
  assign n25254 = ~n25252 & ~n25253;
  assign n25255 = ~n25251 & n25254;
  assign n25256 = ~n25250 & n25255;
  assign n25257 = pi59  & ~n25256;
  assign n25258 = pi59  & ~n25257;
  assign n25259 = ~n25256 & ~n25257;
  assign n25260 = ~n25258 & ~n25259;
  assign n25261 = ~n25249 & ~n25260;
  assign n25262 = n25249 & n25260;
  assign n25263 = ~n25261 & ~n25262;
  assign n25264 = n25223 & ~n25263;
  assign n25265 = ~n25223 & n25263;
  assign n25266 = ~n25264 & ~n25265;
  assign n25267 = n8936 & n10394;
  assign n25268 = pi112  & n10744;
  assign n25269 = pi114  & n10392;
  assign n25270 = pi113  & n10387;
  assign n25271 = ~n25269 & ~n25270;
  assign n25272 = ~n25268 & n25271;
  assign n25273 = ~n25267 & n25272;
  assign n25274 = pi56  & ~n25273;
  assign n25275 = pi56  & ~n25274;
  assign n25276 = ~n25273 & ~n25274;
  assign n25277 = ~n25275 & ~n25276;
  assign n25278 = ~n25266 & n25277;
  assign n25279 = n25266 & ~n25277;
  assign n25280 = ~n25278 & ~n25279;
  assign n25281 = ~n25222 & n25280;
  assign n25282 = ~n25222 & ~n25281;
  assign n25283 = n25280 & ~n25281;
  assign n25284 = ~n25282 & ~n25283;
  assign n25285 = ~n25221 & ~n25284;
  assign n25286 = n25221 & n25284;
  assign n25287 = ~n25285 & ~n25286;
  assign n25288 = ~n25210 & n25287;
  assign n25289 = ~n25210 & ~n25288;
  assign n25290 = n25287 & ~n25288;
  assign n25291 = ~n25289 & ~n25290;
  assign n25292 = ~n25209 & ~n25291;
  assign n25293 = n25209 & n25291;
  assign n25294 = ~n25292 & ~n25293;
  assign n25295 = ~n25198 & n25294;
  assign n25296 = n25198 & ~n25294;
  assign n25297 = ~n25295 & ~n25296;
  assign n25298 = n7408 & n12158;
  assign n25299 = pi121  & n7740;
  assign n25300 = pi123  & n7406;
  assign n25301 = pi122  & n7401;
  assign n25302 = ~n25300 & ~n25301;
  assign n25303 = ~n25299 & n25302;
  assign n25304 = ~n25298 & n25303;
  assign n25305 = pi47  & ~n25304;
  assign n25306 = pi47  & ~n25305;
  assign n25307 = ~n25304 & ~n25305;
  assign n25308 = ~n25306 & ~n25307;
  assign n25309 = n25297 & ~n25308;
  assign n25310 = n25297 & ~n25309;
  assign n25311 = ~n25308 & ~n25309;
  assign n25312 = ~n25310 & ~n25311;
  assign n25313 = ~n25137 & ~n25150;
  assign n25314 = n25312 & n25313;
  assign n25315 = ~n25312 & ~n25313;
  assign n25316 = ~n25314 & ~n25315;
  assign n25317 = n6539 & n13344;
  assign n25318 = pi124  & n6873;
  assign n25319 = pi126  & n6537;
  assign n25320 = pi125  & n6532;
  assign n25321 = ~n25319 & ~n25320;
  assign n25322 = ~n25318 & n25321;
  assign n25323 = ~n25317 & n25322;
  assign n25324 = pi44  & ~n25323;
  assign n25325 = pi44  & ~n25324;
  assign n25326 = ~n25323 & ~n25324;
  assign n25327 = ~n25325 & ~n25326;
  assign n25328 = n25316 & ~n25327;
  assign n25329 = n25316 & ~n25328;
  assign n25330 = ~n25327 & ~n25328;
  assign n25331 = ~n25329 & ~n25330;
  assign n25332 = ~n25197 & n25331;
  assign n25333 = n25197 & ~n25331;
  assign n25334 = ~n25332 & ~n25333;
  assign n25335 = ~n25185 & ~n25334;
  assign n25336 = n25185 & n25334;
  assign n25337 = ~n25335 & ~n25336;
  assign n25338 = ~n25184 & n25337;
  assign n25339 = n25184 & ~n25337;
  assign po104  = ~n25338 & ~n25339;
  assign n25341 = ~n25335 & ~n25338;
  assign n25342 = ~n25288 & ~n25292;
  assign n25343 = n8334 & n11389;
  assign n25344 = pi119  & n8685;
  assign n25345 = pi121  & n8332;
  assign n25346 = pi120  & n8327;
  assign n25347 = ~n25345 & ~n25346;
  assign n25348 = ~n25344 & n25347;
  assign n25349 = ~n25343 & n25348;
  assign n25350 = pi50  & ~n25349;
  assign n25351 = pi50  & ~n25350;
  assign n25352 = ~n25349 & ~n25350;
  assign n25353 = ~n25351 & ~n25352;
  assign n25354 = ~n25281 & ~n25285;
  assign n25355 = ~n25265 & ~n25279;
  assign n25356 = n8963 & n10394;
  assign n25357 = pi113  & n10744;
  assign n25358 = pi115  & n10392;
  assign n25359 = pi114  & n10387;
  assign n25360 = ~n25358 & ~n25359;
  assign n25361 = ~n25357 & n25360;
  assign n25362 = ~n25356 & n25361;
  assign n25363 = pi56  & ~n25362;
  assign n25364 = pi56  & ~n25363;
  assign n25365 = ~n25362 & ~n25363;
  assign n25366 = ~n25364 & ~n25365;
  assign n25367 = pi41  & ~n25039;
  assign n25368 = ~pi41  & n25039;
  assign n25369 = ~n25367 & ~n25368;
  assign n25370 = pi105  & n13835;
  assign n25371 = pi106  & ~n13434;
  assign n25372 = ~n25370 & ~n25371;
  assign n25373 = n25369 & n25372;
  assign n25374 = ~n25369 & ~n25372;
  assign n25375 = ~n25373 & ~n25374;
  assign n25376 = n7349 & n12627;
  assign n25377 = pi107  & n13004;
  assign n25378 = pi109  & n12625;
  assign n25379 = pi108  & n12620;
  assign n25380 = ~n25378 & ~n25379;
  assign n25381 = ~n25377 & n25380;
  assign n25382 = ~n25376 & n25381;
  assign n25383 = pi62  & ~n25382;
  assign n25384 = pi62  & ~n25383;
  assign n25385 = ~n25382 & ~n25383;
  assign n25386 = ~n25384 & ~n25385;
  assign n25387 = n25375 & ~n25386;
  assign n25388 = n25375 & ~n25387;
  assign n25389 = ~n25386 & ~n25387;
  assign n25390 = ~n25388 & ~n25389;
  assign n25391 = ~n25228 & ~n25232;
  assign n25392 = n25390 & n25391;
  assign n25393 = ~n25390 & ~n25391;
  assign n25394 = ~n25392 & ~n25393;
  assign n25395 = n7997 & n11488;
  assign n25396 = pi110  & n11847;
  assign n25397 = pi112  & n11486;
  assign n25398 = pi111  & n11481;
  assign n25399 = ~n25397 & ~n25398;
  assign n25400 = ~n25396 & n25399;
  assign n25401 = ~n25395 & n25400;
  assign n25402 = pi59  & ~n25401;
  assign n25403 = pi59  & ~n25402;
  assign n25404 = ~n25401 & ~n25402;
  assign n25405 = ~n25403 & ~n25404;
  assign n25406 = n25394 & ~n25405;
  assign n25407 = n25394 & ~n25406;
  assign n25408 = ~n25405 & ~n25406;
  assign n25409 = ~n25407 & ~n25408;
  assign n25410 = ~n25235 & ~n25246;
  assign n25411 = ~n25261 & ~n25410;
  assign n25412 = ~n25409 & ~n25411;
  assign n25413 = n25409 & n25411;
  assign n25414 = ~n25412 & ~n25413;
  assign n25415 = ~n25366 & n25414;
  assign n25416 = ~n25366 & ~n25415;
  assign n25417 = n25414 & ~n25415;
  assign n25418 = ~n25416 & ~n25417;
  assign n25419 = ~n25355 & ~n25418;
  assign n25420 = ~n25355 & ~n25419;
  assign n25421 = ~n25418 & ~n25419;
  assign n25422 = ~n25420 & ~n25421;
  assign n25423 = n9310 & n9984;
  assign n25424 = pi116  & n9701;
  assign n25425 = pi118  & n9308;
  assign n25426 = pi117  & n9303;
  assign n25427 = ~n25425 & ~n25426;
  assign n25428 = ~n25424 & n25427;
  assign n25429 = ~n25423 & n25428;
  assign n25430 = pi53  & ~n25429;
  assign n25431 = pi53  & ~n25430;
  assign n25432 = ~n25429 & ~n25430;
  assign n25433 = ~n25431 & ~n25432;
  assign n25434 = n25422 & n25433;
  assign n25435 = ~n25422 & ~n25433;
  assign n25436 = ~n25434 & ~n25435;
  assign n25437 = ~n25354 & n25436;
  assign n25438 = n25354 & ~n25436;
  assign n25439 = ~n25437 & ~n25438;
  assign n25440 = n25353 & ~n25439;
  assign n25441 = ~n25353 & n25439;
  assign n25442 = ~n25440 & ~n25441;
  assign n25443 = ~n25342 & n25442;
  assign n25444 = n25342 & ~n25442;
  assign n25445 = ~n25443 & ~n25444;
  assign n25446 = n7408 & n12189;
  assign n25447 = pi122  & n7740;
  assign n25448 = pi124  & n7406;
  assign n25449 = pi123  & n7401;
  assign n25450 = ~n25448 & ~n25449;
  assign n25451 = ~n25447 & n25450;
  assign n25452 = ~n25446 & n25451;
  assign n25453 = pi47  & ~n25452;
  assign n25454 = pi47  & ~n25453;
  assign n25455 = ~n25452 & ~n25453;
  assign n25456 = ~n25454 & ~n25455;
  assign n25457 = n25445 & ~n25456;
  assign n25458 = n25445 & ~n25457;
  assign n25459 = ~n25456 & ~n25457;
  assign n25460 = ~n25458 & ~n25459;
  assign n25461 = ~n25295 & ~n25309;
  assign n25462 = n25460 & n25461;
  assign n25463 = ~n25460 & ~n25461;
  assign n25464 = ~n25462 & ~n25463;
  assign n25465 = n6539 & n13742;
  assign n25466 = pi125  & n6873;
  assign n25467 = pi127  & n6537;
  assign n25468 = pi126  & n6532;
  assign n25469 = ~n25467 & ~n25468;
  assign n25470 = ~n25466 & n25469;
  assign n25471 = ~n25465 & n25470;
  assign n25472 = pi44  & ~n25471;
  assign n25473 = pi44  & ~n25472;
  assign n25474 = ~n25471 & ~n25472;
  assign n25475 = ~n25473 & ~n25474;
  assign n25476 = n25464 & ~n25475;
  assign n25477 = n25464 & ~n25476;
  assign n25478 = ~n25475 & ~n25476;
  assign n25479 = ~n25477 & ~n25478;
  assign n25480 = ~n25315 & ~n25328;
  assign n25481 = n25479 & n25480;
  assign n25482 = ~n25479 & ~n25480;
  assign n25483 = ~n25481 & ~n25482;
  assign n25484 = ~n25197 & ~n25331;
  assign n25485 = ~n25194 & ~n25484;
  assign n25486 = n25483 & ~n25485;
  assign n25487 = ~n25483 & n25485;
  assign n25488 = ~n25486 & ~n25487;
  assign n25489 = ~n25341 & n25488;
  assign n25490 = n25341 & ~n25488;
  assign po105  = ~n25489 & ~n25490;
  assign n25492 = ~n25457 & ~n25463;
  assign n25493 = pi126  & n6873;
  assign n25494 = pi127  & n6532;
  assign n25495 = ~n25493 & ~n25494;
  assign n25496 = ~n6539 & n25495;
  assign n25497 = n13773 & n25495;
  assign n25498 = ~n25496 & ~n25497;
  assign n25499 = pi44  & ~n25498;
  assign n25500 = ~pi44  & n25498;
  assign n25501 = ~n25499 & ~n25500;
  assign n25502 = ~n25492 & ~n25501;
  assign n25503 = n25492 & n25501;
  assign n25504 = ~n25502 & ~n25503;
  assign n25505 = n7408 & n12943;
  assign n25506 = pi123  & n7740;
  assign n25507 = pi125  & n7406;
  assign n25508 = pi124  & n7401;
  assign n25509 = ~n25507 & ~n25508;
  assign n25510 = ~n25506 & n25509;
  assign n25511 = ~n25505 & n25510;
  assign n25512 = pi47  & ~n25511;
  assign n25513 = pi47  & ~n25512;
  assign n25514 = ~n25511 & ~n25512;
  assign n25515 = ~n25513 & ~n25514;
  assign n25516 = ~n25441 & ~n25443;
  assign n25517 = ~n25435 & ~n25437;
  assign n25518 = ~n25387 & ~n25393;
  assign n25519 = pi106  & n13835;
  assign n25520 = pi107  & ~n13434;
  assign n25521 = ~n25519 & ~n25520;
  assign n25522 = ~pi41  & ~n25039;
  assign n25523 = ~n25374 & ~n25522;
  assign n25524 = n25521 & ~n25523;
  assign n25525 = n25521 & ~n25524;
  assign n25526 = ~n25523 & ~n25524;
  assign n25527 = ~n25525 & ~n25526;
  assign n25528 = pi108  & n13004;
  assign n25529 = pi110  & n12625;
  assign n25530 = pi109  & n12620;
  assign n25531 = ~n25529 & ~n25530;
  assign n25532 = ~n25528 & n25531;
  assign n25533 = ~n12627 & n25532;
  assign n25534 = ~n7665 & n25532;
  assign n25535 = ~n25533 & ~n25534;
  assign n25536 = pi62  & ~n25535;
  assign n25537 = ~pi62  & n25535;
  assign n25538 = ~n25536 & ~n25537;
  assign n25539 = ~n25527 & ~n25538;
  assign n25540 = n25527 & n25538;
  assign n25541 = ~n25539 & ~n25540;
  assign n25542 = ~n25518 & n25541;
  assign n25543 = n25518 & ~n25541;
  assign n25544 = ~n25542 & ~n25543;
  assign n25545 = n8612 & n11488;
  assign n25546 = pi111  & n11847;
  assign n25547 = pi113  & n11486;
  assign n25548 = pi112  & n11481;
  assign n25549 = ~n25547 & ~n25548;
  assign n25550 = ~n25546 & n25549;
  assign n25551 = ~n25545 & n25550;
  assign n25552 = pi59  & ~n25551;
  assign n25553 = pi59  & ~n25552;
  assign n25554 = ~n25551 & ~n25552;
  assign n25555 = ~n25553 & ~n25554;
  assign n25556 = n25544 & ~n25555;
  assign n25557 = n25544 & ~n25556;
  assign n25558 = ~n25555 & ~n25556;
  assign n25559 = ~n25557 & ~n25558;
  assign n25560 = ~n25406 & ~n25412;
  assign n25561 = n25559 & n25560;
  assign n25562 = ~n25559 & ~n25560;
  assign n25563 = ~n25561 & ~n25562;
  assign n25564 = n9614 & n10394;
  assign n25565 = pi114  & n10744;
  assign n25566 = pi116  & n10392;
  assign n25567 = pi115  & n10387;
  assign n25568 = ~n25566 & ~n25567;
  assign n25569 = ~n25565 & n25568;
  assign n25570 = ~n25564 & n25569;
  assign n25571 = pi56  & ~n25570;
  assign n25572 = pi56  & ~n25571;
  assign n25573 = ~n25570 & ~n25571;
  assign n25574 = ~n25572 & ~n25573;
  assign n25575 = n25563 & ~n25574;
  assign n25576 = n25563 & ~n25575;
  assign n25577 = ~n25574 & ~n25575;
  assign n25578 = ~n25576 & ~n25577;
  assign n25579 = ~n25415 & ~n25419;
  assign n25580 = n25578 & n25579;
  assign n25581 = ~n25578 & ~n25579;
  assign n25582 = ~n25580 & ~n25581;
  assign n25583 = n9310 & n10667;
  assign n25584 = pi117  & n9701;
  assign n25585 = pi119  & n9308;
  assign n25586 = pi118  & n9303;
  assign n25587 = ~n25585 & ~n25586;
  assign n25588 = ~n25584 & n25587;
  assign n25589 = ~n25583 & n25588;
  assign n25590 = pi53  & ~n25589;
  assign n25591 = pi53  & ~n25590;
  assign n25592 = ~n25589 & ~n25590;
  assign n25593 = ~n25591 & ~n25592;
  assign n25594 = n25582 & ~n25593;
  assign n25595 = n25582 & ~n25594;
  assign n25596 = ~n25593 & ~n25594;
  assign n25597 = ~n25595 & ~n25596;
  assign n25598 = ~n25517 & n25597;
  assign n25599 = n25517 & ~n25597;
  assign n25600 = ~n25598 & ~n25599;
  assign n25601 = n8334 & n11778;
  assign n25602 = pi120  & n8685;
  assign n25603 = pi122  & n8332;
  assign n25604 = pi121  & n8327;
  assign n25605 = ~n25603 & ~n25604;
  assign n25606 = ~n25602 & n25605;
  assign n25607 = ~n25601 & n25606;
  assign n25608 = pi50  & ~n25607;
  assign n25609 = pi50  & ~n25608;
  assign n25610 = ~n25607 & ~n25608;
  assign n25611 = ~n25609 & ~n25610;
  assign n25612 = n25600 & n25611;
  assign n25613 = ~n25600 & ~n25611;
  assign n25614 = ~n25612 & ~n25613;
  assign n25615 = ~n25516 & n25614;
  assign n25616 = ~n25516 & ~n25615;
  assign n25617 = n25614 & ~n25615;
  assign n25618 = ~n25616 & ~n25617;
  assign n25619 = ~n25515 & ~n25618;
  assign n25620 = ~n25515 & ~n25619;
  assign n25621 = ~n25618 & ~n25619;
  assign n25622 = ~n25620 & ~n25621;
  assign n25623 = n25504 & ~n25622;
  assign n25624 = n25504 & ~n25623;
  assign n25625 = ~n25622 & ~n25623;
  assign n25626 = ~n25624 & ~n25625;
  assign n25627 = ~n25476 & ~n25482;
  assign n25628 = n25626 & n25627;
  assign n25629 = ~n25626 & ~n25627;
  assign n25630 = ~n25628 & ~n25629;
  assign n25631 = ~n25486 & ~n25489;
  assign n25632 = n25630 & ~n25631;
  assign n25633 = ~n25630 & n25631;
  assign po106  = ~n25632 & ~n25633;
  assign n25635 = ~n25629 & ~n25632;
  assign n25636 = ~n25502 & ~n25623;
  assign n25637 = ~n25615 & ~n25619;
  assign n25638 = pi127  & n6873;
  assign n25639 = n6539 & n13770;
  assign n25640 = ~n25638 & ~n25639;
  assign n25641 = pi44  & ~n25640;
  assign n25642 = pi44  & ~n25641;
  assign n25643 = ~n25640 & ~n25641;
  assign n25644 = ~n25642 & ~n25643;
  assign n25645 = ~n25637 & ~n25644;
  assign n25646 = ~n25637 & ~n25645;
  assign n25647 = ~n25644 & ~n25645;
  assign n25648 = ~n25646 & ~n25647;
  assign n25649 = ~n25581 & ~n25594;
  assign n25650 = n9310 & n11028;
  assign n25651 = pi118  & n9701;
  assign n25652 = pi120  & n9308;
  assign n25653 = pi119  & n9303;
  assign n25654 = ~n25652 & ~n25653;
  assign n25655 = ~n25651 & n25654;
  assign n25656 = ~n25650 & n25655;
  assign n25657 = pi53  & ~n25656;
  assign n25658 = pi53  & ~n25657;
  assign n25659 = ~n25656 & ~n25657;
  assign n25660 = ~n25658 & ~n25659;
  assign n25661 = ~n25562 & ~n25575;
  assign n25662 = n9958 & n10394;
  assign n25663 = pi115  & n10744;
  assign n25664 = pi117  & n10392;
  assign n25665 = pi116  & n10387;
  assign n25666 = ~n25664 & ~n25665;
  assign n25667 = ~n25663 & n25666;
  assign n25668 = ~n25662 & n25667;
  assign n25669 = pi56  & ~n25668;
  assign n25670 = pi56  & ~n25669;
  assign n25671 = ~n25668 & ~n25669;
  assign n25672 = ~n25670 & ~n25671;
  assign n25673 = ~n25542 & ~n25556;
  assign n25674 = n8936 & n11488;
  assign n25675 = pi112  & n11847;
  assign n25676 = pi114  & n11486;
  assign n25677 = pi113  & n11481;
  assign n25678 = ~n25676 & ~n25677;
  assign n25679 = ~n25675 & n25678;
  assign n25680 = ~n25674 & n25679;
  assign n25681 = pi59  & ~n25680;
  assign n25682 = pi59  & ~n25681;
  assign n25683 = ~n25680 & ~n25681;
  assign n25684 = ~n25682 & ~n25683;
  assign n25685 = ~n25524 & ~n25539;
  assign n25686 = pi107  & n13835;
  assign n25687 = pi108  & ~n13434;
  assign n25688 = ~n25686 & ~n25687;
  assign n25689 = n25521 & ~n25688;
  assign n25690 = ~n25521 & n25688;
  assign n25691 = ~n25689 & ~n25690;
  assign n25692 = pi109  & n13004;
  assign n25693 = pi111  & n12625;
  assign n25694 = pi110  & n12620;
  assign n25695 = ~n25693 & ~n25694;
  assign n25696 = ~n25692 & n25695;
  assign n25697 = ~n12627 & n25696;
  assign n25698 = ~n7970 & n25696;
  assign n25699 = ~n25697 & ~n25698;
  assign n25700 = pi62  & ~n25699;
  assign n25701 = ~pi62  & n25699;
  assign n25702 = ~n25700 & ~n25701;
  assign n25703 = n25691 & ~n25702;
  assign n25704 = ~n25691 & n25702;
  assign n25705 = ~n25703 & ~n25704;
  assign n25706 = ~n25685 & n25705;
  assign n25707 = ~n25685 & ~n25706;
  assign n25708 = n25705 & ~n25706;
  assign n25709 = ~n25707 & ~n25708;
  assign n25710 = ~n25684 & ~n25709;
  assign n25711 = n25684 & n25709;
  assign n25712 = ~n25710 & ~n25711;
  assign n25713 = ~n25673 & n25712;
  assign n25714 = ~n25673 & ~n25713;
  assign n25715 = n25712 & ~n25713;
  assign n25716 = ~n25714 & ~n25715;
  assign n25717 = ~n25672 & ~n25716;
  assign n25718 = n25672 & n25716;
  assign n25719 = ~n25717 & ~n25718;
  assign n25720 = ~n25661 & n25719;
  assign n25721 = ~n25661 & ~n25720;
  assign n25722 = n25719 & ~n25720;
  assign n25723 = ~n25721 & ~n25722;
  assign n25724 = ~n25660 & ~n25723;
  assign n25725 = n25660 & n25723;
  assign n25726 = ~n25724 & ~n25725;
  assign n25727 = ~n25649 & n25726;
  assign n25728 = n25649 & ~n25726;
  assign n25729 = ~n25727 & ~n25728;
  assign n25730 = n8334 & n12158;
  assign n25731 = pi121  & n8685;
  assign n25732 = pi123  & n8332;
  assign n25733 = pi122  & n8327;
  assign n25734 = ~n25732 & ~n25733;
  assign n25735 = ~n25731 & n25734;
  assign n25736 = ~n25730 & n25735;
  assign n25737 = pi50  & ~n25736;
  assign n25738 = pi50  & ~n25737;
  assign n25739 = ~n25736 & ~n25737;
  assign n25740 = ~n25738 & ~n25739;
  assign n25741 = n25729 & ~n25740;
  assign n25742 = n25729 & ~n25741;
  assign n25743 = ~n25740 & ~n25741;
  assign n25744 = ~n25742 & ~n25743;
  assign n25745 = ~n25517 & ~n25597;
  assign n25746 = ~n25613 & ~n25745;
  assign n25747 = ~n25744 & ~n25746;
  assign n25748 = ~n25744 & ~n25747;
  assign n25749 = ~n25746 & ~n25747;
  assign n25750 = ~n25748 & ~n25749;
  assign n25751 = n7408 & n13344;
  assign n25752 = pi124  & n7740;
  assign n25753 = pi126  & n7406;
  assign n25754 = pi125  & n7401;
  assign n25755 = ~n25753 & ~n25754;
  assign n25756 = ~n25752 & n25755;
  assign n25757 = ~n25751 & n25756;
  assign n25758 = pi47  & ~n25757;
  assign n25759 = pi47  & ~n25758;
  assign n25760 = ~n25757 & ~n25758;
  assign n25761 = ~n25759 & ~n25760;
  assign n25762 = ~n25750 & ~n25761;
  assign n25763 = ~n25750 & ~n25762;
  assign n25764 = ~n25761 & ~n25762;
  assign n25765 = ~n25763 & ~n25764;
  assign n25766 = ~n25648 & n25765;
  assign n25767 = n25648 & ~n25765;
  assign n25768 = ~n25766 & ~n25767;
  assign n25769 = ~n25636 & ~n25768;
  assign n25770 = n25636 & n25768;
  assign n25771 = ~n25769 & ~n25770;
  assign n25772 = ~n25635 & n25771;
  assign n25773 = n25635 & ~n25771;
  assign po107  = ~n25772 & ~n25773;
  assign n25775 = ~n25769 & ~n25772;
  assign n25776 = ~n25727 & ~n25741;
  assign n25777 = n8334 & n12189;
  assign n25778 = pi122  & n8685;
  assign n25779 = pi124  & n8332;
  assign n25780 = pi123  & n8327;
  assign n25781 = ~n25779 & ~n25780;
  assign n25782 = ~n25778 & n25781;
  assign n25783 = ~n25777 & n25782;
  assign n25784 = pi50  & ~n25783;
  assign n25785 = pi50  & ~n25784;
  assign n25786 = ~n25783 & ~n25784;
  assign n25787 = ~n25785 & ~n25786;
  assign n25788 = ~n25720 & ~n25724;
  assign n25789 = n9310 & n11389;
  assign n25790 = pi119  & n9701;
  assign n25791 = pi121  & n9308;
  assign n25792 = pi120  & n9303;
  assign n25793 = ~n25791 & ~n25792;
  assign n25794 = ~n25790 & n25793;
  assign n25795 = ~n25789 & n25794;
  assign n25796 = pi53  & ~n25795;
  assign n25797 = pi53  & ~n25796;
  assign n25798 = ~n25795 & ~n25796;
  assign n25799 = ~n25797 & ~n25798;
  assign n25800 = ~n25713 & ~n25717;
  assign n25801 = n9984 & n10394;
  assign n25802 = pi116  & n10744;
  assign n25803 = pi118  & n10392;
  assign n25804 = pi117  & n10387;
  assign n25805 = ~n25803 & ~n25804;
  assign n25806 = ~n25802 & n25805;
  assign n25807 = ~n25801 & n25806;
  assign n25808 = pi56  & ~n25807;
  assign n25809 = pi56  & ~n25808;
  assign n25810 = ~n25807 & ~n25808;
  assign n25811 = ~n25809 & ~n25810;
  assign n25812 = ~n25706 & ~n25710;
  assign n25813 = ~n25689 & ~n25703;
  assign n25814 = pi108  & n13835;
  assign n25815 = pi109  & ~n13434;
  assign n25816 = ~n25814 & ~n25815;
  assign n25817 = ~pi44  & ~n25816;
  assign n25818 = pi44  & n25816;
  assign n25819 = ~n25817 & ~n25818;
  assign n25820 = ~n25521 & n25819;
  assign n25821 = ~n25521 & ~n25820;
  assign n25822 = n25819 & ~n25820;
  assign n25823 = ~n25821 & ~n25822;
  assign n25824 = ~n25813 & ~n25823;
  assign n25825 = ~n25813 & ~n25824;
  assign n25826 = ~n25823 & ~n25824;
  assign n25827 = ~n25825 & ~n25826;
  assign n25828 = n7997 & n12627;
  assign n25829 = pi110  & n13004;
  assign n25830 = pi112  & n12625;
  assign n25831 = pi111  & n12620;
  assign n25832 = ~n25830 & ~n25831;
  assign n25833 = ~n25829 & n25832;
  assign n25834 = ~n25828 & n25833;
  assign n25835 = pi62  & ~n25834;
  assign n25836 = pi62  & ~n25835;
  assign n25837 = ~n25834 & ~n25835;
  assign n25838 = ~n25836 & ~n25837;
  assign n25839 = ~n25827 & ~n25838;
  assign n25840 = ~n25827 & ~n25839;
  assign n25841 = ~n25838 & ~n25839;
  assign n25842 = ~n25840 & ~n25841;
  assign n25843 = n8963 & n11488;
  assign n25844 = pi113  & n11847;
  assign n25845 = pi115  & n11486;
  assign n25846 = pi114  & n11481;
  assign n25847 = ~n25845 & ~n25846;
  assign n25848 = ~n25844 & n25847;
  assign n25849 = ~n25843 & n25848;
  assign n25850 = pi59  & ~n25849;
  assign n25851 = pi59  & ~n25850;
  assign n25852 = ~n25849 & ~n25850;
  assign n25853 = ~n25851 & ~n25852;
  assign n25854 = n25842 & n25853;
  assign n25855 = ~n25842 & ~n25853;
  assign n25856 = ~n25854 & ~n25855;
  assign n25857 = ~n25812 & n25856;
  assign n25858 = n25812 & ~n25856;
  assign n25859 = ~n25857 & ~n25858;
  assign n25860 = n25811 & ~n25859;
  assign n25861 = ~n25811 & n25859;
  assign n25862 = ~n25860 & ~n25861;
  assign n25863 = ~n25800 & n25862;
  assign n25864 = n25800 & ~n25862;
  assign n25865 = ~n25863 & ~n25864;
  assign n25866 = n25799 & ~n25865;
  assign n25867 = ~n25799 & n25865;
  assign n25868 = ~n25866 & ~n25867;
  assign n25869 = ~n25788 & n25868;
  assign n25870 = n25788 & ~n25868;
  assign n25871 = ~n25869 & ~n25870;
  assign n25872 = n25787 & ~n25871;
  assign n25873 = ~n25787 & n25871;
  assign n25874 = ~n25872 & ~n25873;
  assign n25875 = ~n25776 & n25874;
  assign n25876 = n25776 & ~n25874;
  assign n25877 = ~n25875 & ~n25876;
  assign n25878 = n7408 & n13742;
  assign n25879 = pi125  & n7740;
  assign n25880 = pi127  & n7406;
  assign n25881 = pi126  & n7401;
  assign n25882 = ~n25880 & ~n25881;
  assign n25883 = ~n25879 & n25882;
  assign n25884 = ~n25878 & n25883;
  assign n25885 = pi47  & ~n25884;
  assign n25886 = pi47  & ~n25885;
  assign n25887 = ~n25884 & ~n25885;
  assign n25888 = ~n25886 & ~n25887;
  assign n25889 = n25877 & ~n25888;
  assign n25890 = n25877 & ~n25889;
  assign n25891 = ~n25888 & ~n25889;
  assign n25892 = ~n25890 & ~n25891;
  assign n25893 = ~n25747 & ~n25762;
  assign n25894 = n25892 & n25893;
  assign n25895 = ~n25892 & ~n25893;
  assign n25896 = ~n25894 & ~n25895;
  assign n25897 = ~n25648 & ~n25765;
  assign n25898 = ~n25645 & ~n25897;
  assign n25899 = n25896 & ~n25898;
  assign n25900 = ~n25896 & n25898;
  assign n25901 = ~n25899 & ~n25900;
  assign n25902 = ~n25775 & n25901;
  assign n25903 = n25775 & ~n25901;
  assign po108  = ~n25902 & ~n25903;
  assign n25905 = ~n25873 & ~n25875;
  assign n25906 = pi126  & n7740;
  assign n25907 = pi127  & n7401;
  assign n25908 = ~n25906 & ~n25907;
  assign n25909 = ~n7408 & n25908;
  assign n25910 = n13773 & n25908;
  assign n25911 = ~n25909 & ~n25910;
  assign n25912 = pi47  & ~n25911;
  assign n25913 = ~pi47  & n25911;
  assign n25914 = ~n25912 & ~n25913;
  assign n25915 = ~n25905 & ~n25914;
  assign n25916 = n25905 & n25914;
  assign n25917 = ~n25915 & ~n25916;
  assign n25918 = n8334 & n12943;
  assign n25919 = pi123  & n8685;
  assign n25920 = pi125  & n8332;
  assign n25921 = pi124  & n8327;
  assign n25922 = ~n25920 & ~n25921;
  assign n25923 = ~n25919 & n25922;
  assign n25924 = ~n25918 & n25923;
  assign n25925 = pi50  & ~n25924;
  assign n25926 = pi50  & ~n25925;
  assign n25927 = ~n25924 & ~n25925;
  assign n25928 = ~n25926 & ~n25927;
  assign n25929 = ~n25867 & ~n25869;
  assign n25930 = ~n25861 & ~n25863;
  assign n25931 = ~n25855 & ~n25857;
  assign n25932 = n9614 & n11488;
  assign n25933 = pi114  & n11847;
  assign n25934 = pi116  & n11486;
  assign n25935 = pi115  & n11481;
  assign n25936 = ~n25934 & ~n25935;
  assign n25937 = ~n25933 & n25936;
  assign n25938 = ~n25932 & n25937;
  assign n25939 = pi59  & ~n25938;
  assign n25940 = pi59  & ~n25939;
  assign n25941 = ~n25938 & ~n25939;
  assign n25942 = ~n25940 & ~n25941;
  assign n25943 = ~n25824 & ~n25839;
  assign n25944 = pi109  & n13835;
  assign n25945 = pi110  & ~n13434;
  assign n25946 = ~n25944 & ~n25945;
  assign n25947 = ~n25817 & ~n25820;
  assign n25948 = ~n25946 & n25947;
  assign n25949 = n25946 & ~n25947;
  assign n25950 = ~n25948 & ~n25949;
  assign n25951 = n8612 & n12627;
  assign n25952 = pi111  & n13004;
  assign n25953 = pi113  & n12625;
  assign n25954 = pi112  & n12620;
  assign n25955 = ~n25953 & ~n25954;
  assign n25956 = ~n25952 & n25955;
  assign n25957 = ~n25951 & n25956;
  assign n25958 = pi62  & ~n25957;
  assign n25959 = pi62  & ~n25958;
  assign n25960 = ~n25957 & ~n25958;
  assign n25961 = ~n25959 & ~n25960;
  assign n25962 = ~n25950 & n25961;
  assign n25963 = n25950 & ~n25961;
  assign n25964 = ~n25962 & ~n25963;
  assign n25965 = ~n25943 & n25964;
  assign n25966 = ~n25943 & ~n25965;
  assign n25967 = n25964 & ~n25965;
  assign n25968 = ~n25966 & ~n25967;
  assign n25969 = ~n25942 & ~n25968;
  assign n25970 = n25942 & n25968;
  assign n25971 = ~n25969 & ~n25970;
  assign n25972 = ~n25931 & n25971;
  assign n25973 = n25931 & ~n25971;
  assign n25974 = ~n25972 & ~n25973;
  assign n25975 = n10394 & n10667;
  assign n25976 = pi117  & n10744;
  assign n25977 = pi119  & n10392;
  assign n25978 = pi118  & n10387;
  assign n25979 = ~n25977 & ~n25978;
  assign n25980 = ~n25976 & n25979;
  assign n25981 = ~n25975 & n25980;
  assign n25982 = pi56  & ~n25981;
  assign n25983 = pi56  & ~n25982;
  assign n25984 = ~n25981 & ~n25982;
  assign n25985 = ~n25983 & ~n25984;
  assign n25986 = n25974 & ~n25985;
  assign n25987 = n25974 & ~n25986;
  assign n25988 = ~n25985 & ~n25986;
  assign n25989 = ~n25987 & ~n25988;
  assign n25990 = ~n25930 & n25989;
  assign n25991 = n25930 & ~n25989;
  assign n25992 = ~n25990 & ~n25991;
  assign n25993 = n9310 & n11778;
  assign n25994 = pi120  & n9701;
  assign n25995 = pi122  & n9308;
  assign n25996 = pi121  & n9303;
  assign n25997 = ~n25995 & ~n25996;
  assign n25998 = ~n25994 & n25997;
  assign n25999 = ~n25993 & n25998;
  assign n26000 = pi53  & ~n25999;
  assign n26001 = pi53  & ~n26000;
  assign n26002 = ~n25999 & ~n26000;
  assign n26003 = ~n26001 & ~n26002;
  assign n26004 = n25992 & n26003;
  assign n26005 = ~n25992 & ~n26003;
  assign n26006 = ~n26004 & ~n26005;
  assign n26007 = ~n25929 & n26006;
  assign n26008 = ~n25929 & ~n26007;
  assign n26009 = n26006 & ~n26007;
  assign n26010 = ~n26008 & ~n26009;
  assign n26011 = ~n25928 & ~n26010;
  assign n26012 = ~n25928 & ~n26011;
  assign n26013 = ~n26010 & ~n26011;
  assign n26014 = ~n26012 & ~n26013;
  assign n26015 = n25917 & ~n26014;
  assign n26016 = n25917 & ~n26015;
  assign n26017 = ~n26014 & ~n26015;
  assign n26018 = ~n26016 & ~n26017;
  assign n26019 = ~n25889 & ~n25895;
  assign n26020 = n26018 & n26019;
  assign n26021 = ~n26018 & ~n26019;
  assign n26022 = ~n26020 & ~n26021;
  assign n26023 = ~n25899 & ~n25902;
  assign n26024 = n26022 & ~n26023;
  assign n26025 = ~n26022 & n26023;
  assign po109  = ~n26024 & ~n26025;
  assign n26027 = ~n25972 & ~n25986;
  assign n26028 = n10394 & n11028;
  assign n26029 = pi118  & n10744;
  assign n26030 = pi120  & n10392;
  assign n26031 = pi119  & n10387;
  assign n26032 = ~n26030 & ~n26031;
  assign n26033 = ~n26029 & n26032;
  assign n26034 = ~n26028 & n26033;
  assign n26035 = pi56  & ~n26034;
  assign n26036 = pi56  & ~n26035;
  assign n26037 = ~n26034 & ~n26035;
  assign n26038 = ~n26036 & ~n26037;
  assign n26039 = ~n25965 & ~n25969;
  assign n26040 = n9958 & n11488;
  assign n26041 = pi115  & n11847;
  assign n26042 = pi117  & n11486;
  assign n26043 = pi116  & n11481;
  assign n26044 = ~n26042 & ~n26043;
  assign n26045 = ~n26041 & n26044;
  assign n26046 = ~n26040 & n26045;
  assign n26047 = pi59  & ~n26046;
  assign n26048 = pi59  & ~n26047;
  assign n26049 = ~n26046 & ~n26047;
  assign n26050 = ~n26048 & ~n26049;
  assign n26051 = ~n25949 & ~n25963;
  assign n26052 = pi110  & n13835;
  assign n26053 = pi111  & ~n13434;
  assign n26054 = ~n26052 & ~n26053;
  assign n26055 = n25946 & ~n26054;
  assign n26056 = ~n25946 & n26054;
  assign n26057 = ~n26055 & ~n26056;
  assign n26058 = ~n26051 & n26057;
  assign n26059 = ~n26051 & ~n26058;
  assign n26060 = ~n26056 & ~n26058;
  assign n26061 = ~n26055 & n26060;
  assign n26062 = ~n26059 & ~n26061;
  assign n26063 = n8936 & n12627;
  assign n26064 = pi112  & n13004;
  assign n26065 = pi114  & n12625;
  assign n26066 = pi113  & n12620;
  assign n26067 = ~n26065 & ~n26066;
  assign n26068 = ~n26064 & n26067;
  assign n26069 = ~n26063 & n26068;
  assign n26070 = pi62  & ~n26069;
  assign n26071 = pi62  & ~n26070;
  assign n26072 = ~n26069 & ~n26070;
  assign n26073 = ~n26071 & ~n26072;
  assign n26074 = ~n26062 & n26073;
  assign n26075 = n26062 & ~n26073;
  assign n26076 = ~n26074 & ~n26075;
  assign n26077 = ~n26050 & ~n26076;
  assign n26078 = n26050 & n26076;
  assign n26079 = ~n26077 & ~n26078;
  assign n26080 = ~n26039 & n26079;
  assign n26081 = ~n26039 & ~n26080;
  assign n26082 = n26079 & ~n26080;
  assign n26083 = ~n26081 & ~n26082;
  assign n26084 = ~n26038 & ~n26083;
  assign n26085 = n26038 & n26083;
  assign n26086 = ~n26084 & ~n26085;
  assign n26087 = ~n26027 & n26086;
  assign n26088 = n26027 & ~n26086;
  assign n26089 = ~n26087 & ~n26088;
  assign n26090 = n9310 & n12158;
  assign n26091 = pi121  & n9701;
  assign n26092 = pi123  & n9308;
  assign n26093 = pi122  & n9303;
  assign n26094 = ~n26092 & ~n26093;
  assign n26095 = ~n26091 & n26094;
  assign n26096 = ~n26090 & n26095;
  assign n26097 = pi53  & ~n26096;
  assign n26098 = pi53  & ~n26097;
  assign n26099 = ~n26096 & ~n26097;
  assign n26100 = ~n26098 & ~n26099;
  assign n26101 = n26089 & ~n26100;
  assign n26102 = n26089 & ~n26101;
  assign n26103 = ~n26100 & ~n26101;
  assign n26104 = ~n26102 & ~n26103;
  assign n26105 = ~n25930 & ~n25989;
  assign n26106 = ~n26005 & ~n26105;
  assign n26107 = ~n26104 & ~n26106;
  assign n26108 = ~n26104 & ~n26107;
  assign n26109 = ~n26106 & ~n26107;
  assign n26110 = ~n26108 & ~n26109;
  assign n26111 = n8334 & n13344;
  assign n26112 = pi124  & n8685;
  assign n26113 = pi126  & n8332;
  assign n26114 = pi125  & n8327;
  assign n26115 = ~n26113 & ~n26114;
  assign n26116 = ~n26112 & n26115;
  assign n26117 = ~n26111 & n26116;
  assign n26118 = pi50  & ~n26117;
  assign n26119 = pi50  & ~n26118;
  assign n26120 = ~n26117 & ~n26118;
  assign n26121 = ~n26119 & ~n26120;
  assign n26122 = ~n26110 & ~n26121;
  assign n26123 = ~n26110 & ~n26122;
  assign n26124 = ~n26121 & ~n26122;
  assign n26125 = ~n26123 & ~n26124;
  assign n26126 = ~n26007 & ~n26011;
  assign n26127 = pi127  & n7740;
  assign n26128 = ~n7408 & ~n26127;
  assign n26129 = ~n13770 & ~n26127;
  assign n26130 = ~n26128 & ~n26129;
  assign n26131 = pi47  & ~n26130;
  assign n26132 = ~pi47  & n26130;
  assign n26133 = ~n26131 & ~n26132;
  assign n26134 = ~n26126 & ~n26133;
  assign n26135 = n26126 & n26133;
  assign n26136 = ~n26134 & ~n26135;
  assign n26137 = ~n26125 & n26136;
  assign n26138 = ~n26125 & ~n26137;
  assign n26139 = n26136 & ~n26137;
  assign n26140 = ~n26138 & ~n26139;
  assign n26141 = ~n25915 & ~n26015;
  assign n26142 = n26140 & n26141;
  assign n26143 = ~n26140 & ~n26141;
  assign n26144 = ~n26142 & ~n26143;
  assign n26145 = ~n26021 & ~n26024;
  assign n26146 = n26144 & ~n26145;
  assign n26147 = ~n26144 & n26145;
  assign po110  = ~n26146 & ~n26147;
  assign n26149 = ~n26087 & ~n26101;
  assign n26150 = n9310 & n12189;
  assign n26151 = pi122  & n9701;
  assign n26152 = pi124  & n9308;
  assign n26153 = pi123  & n9303;
  assign n26154 = ~n26152 & ~n26153;
  assign n26155 = ~n26151 & n26154;
  assign n26156 = ~n26150 & n26155;
  assign n26157 = pi53  & ~n26156;
  assign n26158 = pi53  & ~n26157;
  assign n26159 = ~n26156 & ~n26157;
  assign n26160 = ~n26158 & ~n26159;
  assign n26161 = ~n26080 & ~n26084;
  assign n26162 = n10394 & n11389;
  assign n26163 = pi119  & n10744;
  assign n26164 = pi121  & n10392;
  assign n26165 = pi120  & n10387;
  assign n26166 = ~n26164 & ~n26165;
  assign n26167 = ~n26163 & n26166;
  assign n26168 = ~n26162 & n26167;
  assign n26169 = pi56  & ~n26168;
  assign n26170 = pi56  & ~n26169;
  assign n26171 = ~n26168 & ~n26169;
  assign n26172 = ~n26170 & ~n26171;
  assign n26173 = ~n26062 & ~n26073;
  assign n26174 = ~n26077 & ~n26173;
  assign n26175 = n8963 & n12627;
  assign n26176 = pi113  & n13004;
  assign n26177 = pi115  & n12625;
  assign n26178 = pi114  & n12620;
  assign n26179 = ~n26177 & ~n26178;
  assign n26180 = ~n26176 & n26179;
  assign n26181 = ~n26175 & n26180;
  assign n26182 = pi62  & ~n26181;
  assign n26183 = pi62  & ~n26182;
  assign n26184 = ~n26181 & ~n26182;
  assign n26185 = ~n26183 & ~n26184;
  assign n26186 = pi111  & n13835;
  assign n26187 = pi112  & ~n13434;
  assign n26188 = ~n26186 & ~n26187;
  assign n26189 = pi47  & ~n26054;
  assign n26190 = ~pi47  & n26054;
  assign n26191 = ~n26189 & ~n26190;
  assign n26192 = ~n26188 & ~n26191;
  assign n26193 = n26188 & n26191;
  assign n26194 = ~n26192 & ~n26193;
  assign n26195 = ~n26185 & n26194;
  assign n26196 = ~n26185 & ~n26195;
  assign n26197 = n26194 & ~n26195;
  assign n26198 = ~n26196 & ~n26197;
  assign n26199 = ~n26060 & ~n26198;
  assign n26200 = ~n26060 & ~n26199;
  assign n26201 = ~n26198 & ~n26199;
  assign n26202 = ~n26200 & ~n26201;
  assign n26203 = n9984 & n11488;
  assign n26204 = pi116  & n11847;
  assign n26205 = pi118  & n11486;
  assign n26206 = pi117  & n11481;
  assign n26207 = ~n26205 & ~n26206;
  assign n26208 = ~n26204 & n26207;
  assign n26209 = ~n26203 & n26208;
  assign n26210 = pi59  & ~n26209;
  assign n26211 = pi59  & ~n26210;
  assign n26212 = ~n26209 & ~n26210;
  assign n26213 = ~n26211 & ~n26212;
  assign n26214 = n26202 & n26213;
  assign n26215 = ~n26202 & ~n26213;
  assign n26216 = ~n26214 & ~n26215;
  assign n26217 = ~n26174 & n26216;
  assign n26218 = n26174 & ~n26216;
  assign n26219 = ~n26217 & ~n26218;
  assign n26220 = n26172 & ~n26219;
  assign n26221 = ~n26172 & n26219;
  assign n26222 = ~n26220 & ~n26221;
  assign n26223 = ~n26161 & n26222;
  assign n26224 = n26161 & ~n26222;
  assign n26225 = ~n26223 & ~n26224;
  assign n26226 = n26160 & ~n26225;
  assign n26227 = ~n26160 & n26225;
  assign n26228 = ~n26226 & ~n26227;
  assign n26229 = ~n26149 & n26228;
  assign n26230 = n26149 & ~n26228;
  assign n26231 = ~n26229 & ~n26230;
  assign n26232 = n8334 & n13742;
  assign n26233 = pi125  & n8685;
  assign n26234 = pi127  & n8332;
  assign n26235 = pi126  & n8327;
  assign n26236 = ~n26234 & ~n26235;
  assign n26237 = ~n26233 & n26236;
  assign n26238 = ~n26232 & n26237;
  assign n26239 = pi50  & ~n26238;
  assign n26240 = pi50  & ~n26239;
  assign n26241 = ~n26238 & ~n26239;
  assign n26242 = ~n26240 & ~n26241;
  assign n26243 = n26231 & ~n26242;
  assign n26244 = n26231 & ~n26243;
  assign n26245 = ~n26242 & ~n26243;
  assign n26246 = ~n26244 & ~n26245;
  assign n26247 = ~n26107 & ~n26122;
  assign n26248 = n26246 & n26247;
  assign n26249 = ~n26246 & ~n26247;
  assign n26250 = ~n26248 & ~n26249;
  assign n26251 = ~n26134 & ~n26137;
  assign n26252 = ~n26250 & n26251;
  assign n26253 = n26250 & ~n26251;
  assign n26254 = ~n26252 & ~n26253;
  assign n26255 = ~n26143 & ~n26146;
  assign n26256 = n26254 & ~n26255;
  assign n26257 = ~n26254 & n26255;
  assign po111  = ~n26256 & ~n26257;
  assign n26259 = ~n26227 & ~n26229;
  assign n26260 = n9310 & n12943;
  assign n26261 = pi123  & n9701;
  assign n26262 = pi125  & n9308;
  assign n26263 = pi124  & n9303;
  assign n26264 = ~n26262 & ~n26263;
  assign n26265 = ~n26261 & n26264;
  assign n26266 = ~n26260 & n26265;
  assign n26267 = pi53  & ~n26266;
  assign n26268 = pi53  & ~n26267;
  assign n26269 = ~n26266 & ~n26267;
  assign n26270 = ~n26268 & ~n26269;
  assign n26271 = ~n26221 & ~n26223;
  assign n26272 = n10394 & n11778;
  assign n26273 = pi120  & n10744;
  assign n26274 = pi122  & n10392;
  assign n26275 = pi121  & n10387;
  assign n26276 = ~n26274 & ~n26275;
  assign n26277 = ~n26273 & n26276;
  assign n26278 = ~n26272 & n26277;
  assign n26279 = pi56  & ~n26278;
  assign n26280 = pi56  & ~n26279;
  assign n26281 = ~n26278 & ~n26279;
  assign n26282 = ~n26280 & ~n26281;
  assign n26283 = ~n26215 & ~n26217;
  assign n26284 = n10667 & n11488;
  assign n26285 = pi117  & n11847;
  assign n26286 = pi119  & n11486;
  assign n26287 = pi118  & n11481;
  assign n26288 = ~n26286 & ~n26287;
  assign n26289 = ~n26285 & n26288;
  assign n26290 = ~n26284 & n26289;
  assign n26291 = pi59  & ~n26290;
  assign n26292 = pi59  & ~n26291;
  assign n26293 = ~n26290 & ~n26291;
  assign n26294 = ~n26292 & ~n26293;
  assign n26295 = ~n26195 & ~n26199;
  assign n26296 = pi112  & n13835;
  assign n26297 = pi113  & ~n13434;
  assign n26298 = ~n26296 & ~n26297;
  assign n26299 = ~pi47  & ~n26054;
  assign n26300 = ~n26192 & ~n26299;
  assign n26301 = n26298 & ~n26300;
  assign n26302 = ~n26298 & n26300;
  assign n26303 = ~n26301 & ~n26302;
  assign n26304 = pi114  & n13004;
  assign n26305 = pi116  & n12625;
  assign n26306 = pi115  & n12620;
  assign n26307 = ~n26305 & ~n26306;
  assign n26308 = ~n26304 & n26307;
  assign n26309 = ~n12627 & n26308;
  assign n26310 = ~n9614 & n26308;
  assign n26311 = ~n26309 & ~n26310;
  assign n26312 = pi62  & ~n26311;
  assign n26313 = ~pi62  & n26311;
  assign n26314 = ~n26312 & ~n26313;
  assign n26315 = n26303 & ~n26314;
  assign n26316 = ~n26303 & n26314;
  assign n26317 = ~n26315 & ~n26316;
  assign n26318 = ~n26295 & n26317;
  assign n26319 = ~n26295 & ~n26318;
  assign n26320 = n26317 & ~n26318;
  assign n26321 = ~n26319 & ~n26320;
  assign n26322 = ~n26294 & ~n26321;
  assign n26323 = n26294 & n26321;
  assign n26324 = ~n26322 & ~n26323;
  assign n26325 = ~n26283 & n26324;
  assign n26326 = n26283 & ~n26324;
  assign n26327 = ~n26325 & ~n26326;
  assign n26328 = ~n26282 & n26327;
  assign n26329 = n26282 & ~n26327;
  assign n26330 = ~n26328 & ~n26329;
  assign n26331 = ~n26271 & n26330;
  assign n26332 = ~n26271 & ~n26331;
  assign n26333 = n26330 & ~n26331;
  assign n26334 = ~n26332 & ~n26333;
  assign n26335 = ~n26270 & ~n26334;
  assign n26336 = n26270 & n26334;
  assign n26337 = ~n26335 & ~n26336;
  assign n26338 = ~n26259 & n26337;
  assign n26339 = n26259 & ~n26337;
  assign n26340 = ~n26338 & ~n26339;
  assign n26341 = n8334 & ~n13773;
  assign n26342 = pi126  & n8685;
  assign n26343 = pi127  & n8327;
  assign n26344 = ~n26342 & ~n26343;
  assign n26345 = ~n26341 & n26344;
  assign n26346 = pi50  & ~n26345;
  assign n26347 = pi50  & ~n26346;
  assign n26348 = ~n26345 & ~n26346;
  assign n26349 = ~n26347 & ~n26348;
  assign n26350 = n26340 & ~n26349;
  assign n26351 = n26340 & ~n26350;
  assign n26352 = ~n26349 & ~n26350;
  assign n26353 = ~n26351 & ~n26352;
  assign n26354 = ~n26243 & ~n26249;
  assign n26355 = n26353 & n26354;
  assign n26356 = ~n26353 & ~n26354;
  assign n26357 = ~n26355 & ~n26356;
  assign n26358 = ~n26253 & ~n26256;
  assign n26359 = n26357 & ~n26358;
  assign n26360 = ~n26357 & n26358;
  assign po112  = ~n26359 & ~n26360;
  assign n26362 = ~n26318 & ~n26322;
  assign n26363 = n9958 & n12627;
  assign n26364 = pi115  & n13004;
  assign n26365 = pi117  & n12625;
  assign n26366 = pi116  & n12620;
  assign n26367 = ~n26365 & ~n26366;
  assign n26368 = ~n26364 & n26367;
  assign n26369 = ~n26363 & n26368;
  assign n26370 = pi62  & ~n26369;
  assign n26371 = pi62  & ~n26370;
  assign n26372 = ~n26369 & ~n26370;
  assign n26373 = ~n26371 & ~n26372;
  assign n26374 = pi113  & n13835;
  assign n26375 = pi114  & ~n13434;
  assign n26376 = ~n26374 & ~n26375;
  assign n26377 = n26298 & ~n26376;
  assign n26378 = n26298 & ~n26377;
  assign n26379 = ~n26376 & ~n26377;
  assign n26380 = ~n26378 & ~n26379;
  assign n26381 = ~n26373 & ~n26380;
  assign n26382 = ~n26373 & ~n26381;
  assign n26383 = ~n26380 & ~n26381;
  assign n26384 = ~n26382 & ~n26383;
  assign n26385 = ~n26301 & ~n26315;
  assign n26386 = n26384 & n26385;
  assign n26387 = ~n26384 & ~n26385;
  assign n26388 = ~n26386 & ~n26387;
  assign n26389 = n11028 & n11488;
  assign n26390 = pi118  & n11847;
  assign n26391 = pi120  & n11486;
  assign n26392 = pi119  & n11481;
  assign n26393 = ~n26391 & ~n26392;
  assign n26394 = ~n26390 & n26393;
  assign n26395 = ~n26389 & n26394;
  assign n26396 = pi59  & ~n26395;
  assign n26397 = pi59  & ~n26396;
  assign n26398 = ~n26395 & ~n26396;
  assign n26399 = ~n26397 & ~n26398;
  assign n26400 = ~n26388 & n26399;
  assign n26401 = n26388 & ~n26399;
  assign n26402 = ~n26400 & ~n26401;
  assign n26403 = ~n26362 & n26402;
  assign n26404 = n26362 & ~n26402;
  assign n26405 = ~n26403 & ~n26404;
  assign n26406 = n10394 & n12158;
  assign n26407 = pi121  & n10744;
  assign n26408 = pi123  & n10392;
  assign n26409 = pi122  & n10387;
  assign n26410 = ~n26408 & ~n26409;
  assign n26411 = ~n26407 & n26410;
  assign n26412 = ~n26406 & n26411;
  assign n26413 = pi56  & ~n26412;
  assign n26414 = pi56  & ~n26413;
  assign n26415 = ~n26412 & ~n26413;
  assign n26416 = ~n26414 & ~n26415;
  assign n26417 = n26405 & ~n26416;
  assign n26418 = n26405 & ~n26417;
  assign n26419 = ~n26416 & ~n26417;
  assign n26420 = ~n26418 & ~n26419;
  assign n26421 = ~n26325 & ~n26328;
  assign n26422 = n26420 & n26421;
  assign n26423 = ~n26420 & ~n26421;
  assign n26424 = ~n26422 & ~n26423;
  assign n26425 = n9310 & n13344;
  assign n26426 = pi124  & n9701;
  assign n26427 = pi126  & n9308;
  assign n26428 = pi125  & n9303;
  assign n26429 = ~n26427 & ~n26428;
  assign n26430 = ~n26426 & n26429;
  assign n26431 = ~n26425 & n26430;
  assign n26432 = pi53  & ~n26431;
  assign n26433 = pi53  & ~n26432;
  assign n26434 = ~n26431 & ~n26432;
  assign n26435 = ~n26433 & ~n26434;
  assign n26436 = n26424 & ~n26435;
  assign n26437 = n26424 & ~n26436;
  assign n26438 = ~n26435 & ~n26436;
  assign n26439 = ~n26437 & ~n26438;
  assign n26440 = ~n26331 & ~n26335;
  assign n26441 = pi127  & n8685;
  assign n26442 = ~n8334 & ~n26441;
  assign n26443 = ~n13770 & ~n26441;
  assign n26444 = ~n26442 & ~n26443;
  assign n26445 = pi50  & ~n26444;
  assign n26446 = ~pi50  & n26444;
  assign n26447 = ~n26445 & ~n26446;
  assign n26448 = ~n26440 & ~n26447;
  assign n26449 = n26440 & n26447;
  assign n26450 = ~n26448 & ~n26449;
  assign n26451 = ~n26439 & n26450;
  assign n26452 = ~n26439 & ~n26451;
  assign n26453 = n26450 & ~n26451;
  assign n26454 = ~n26452 & ~n26453;
  assign n26455 = ~n26338 & ~n26350;
  assign n26456 = n26454 & n26455;
  assign n26457 = ~n26454 & ~n26455;
  assign n26458 = ~n26456 & ~n26457;
  assign n26459 = ~n26356 & ~n26359;
  assign n26460 = n26458 & ~n26459;
  assign n26461 = ~n26458 & n26459;
  assign po113  = ~n26460 & ~n26461;
  assign n26463 = ~n26403 & ~n26417;
  assign n26464 = n10394 & n12189;
  assign n26465 = pi122  & n10744;
  assign n26466 = pi124  & n10392;
  assign n26467 = pi123  & n10387;
  assign n26468 = ~n26466 & ~n26467;
  assign n26469 = ~n26465 & n26468;
  assign n26470 = ~n26464 & n26469;
  assign n26471 = pi56  & ~n26470;
  assign n26472 = pi56  & ~n26471;
  assign n26473 = ~n26470 & ~n26471;
  assign n26474 = ~n26472 & ~n26473;
  assign n26475 = ~n26387 & ~n26401;
  assign n26476 = n11389 & n11488;
  assign n26477 = pi119  & n11847;
  assign n26478 = pi121  & n11486;
  assign n26479 = pi120  & n11481;
  assign n26480 = ~n26478 & ~n26479;
  assign n26481 = ~n26477 & n26480;
  assign n26482 = ~n26476 & n26481;
  assign n26483 = pi59  & ~n26482;
  assign n26484 = pi59  & ~n26483;
  assign n26485 = ~n26482 & ~n26483;
  assign n26486 = ~n26484 & ~n26485;
  assign n26487 = n9984 & n12627;
  assign n26488 = pi116  & n13004;
  assign n26489 = pi118  & n12625;
  assign n26490 = pi117  & n12620;
  assign n26491 = ~n26489 & ~n26490;
  assign n26492 = ~n26488 & n26491;
  assign n26493 = ~n26487 & n26492;
  assign n26494 = pi62  & ~n26493;
  assign n26495 = pi62  & ~n26494;
  assign n26496 = ~n26493 & ~n26494;
  assign n26497 = ~n26495 & ~n26496;
  assign n26498 = ~n26377 & ~n26381;
  assign n26499 = pi114  & n13835;
  assign n26500 = pi115  & ~n13434;
  assign n26501 = ~n26499 & ~n26500;
  assign n26502 = ~pi50  & ~n26501;
  assign n26503 = pi50  & n26501;
  assign n26504 = ~n26502 & ~n26503;
  assign n26505 = ~n26298 & n26504;
  assign n26506 = n26298 & ~n26504;
  assign n26507 = ~n26505 & ~n26506;
  assign n26508 = ~n26498 & n26507;
  assign n26509 = ~n26498 & ~n26508;
  assign n26510 = n26507 & ~n26508;
  assign n26511 = ~n26509 & ~n26510;
  assign n26512 = ~n26497 & ~n26511;
  assign n26513 = n26497 & n26511;
  assign n26514 = ~n26512 & ~n26513;
  assign n26515 = ~n26486 & n26514;
  assign n26516 = ~n26486 & ~n26515;
  assign n26517 = n26514 & ~n26515;
  assign n26518 = ~n26516 & ~n26517;
  assign n26519 = ~n26475 & ~n26518;
  assign n26520 = n26475 & n26518;
  assign n26521 = ~n26519 & ~n26520;
  assign n26522 = ~n26474 & n26521;
  assign n26523 = n26474 & ~n26521;
  assign n26524 = ~n26522 & ~n26523;
  assign n26525 = ~n26463 & n26524;
  assign n26526 = n26463 & ~n26524;
  assign n26527 = ~n26525 & ~n26526;
  assign n26528 = n9310 & n13742;
  assign n26529 = pi125  & n9701;
  assign n26530 = pi127  & n9308;
  assign n26531 = pi126  & n9303;
  assign n26532 = ~n26530 & ~n26531;
  assign n26533 = ~n26529 & n26532;
  assign n26534 = ~n26528 & n26533;
  assign n26535 = pi53  & ~n26534;
  assign n26536 = pi53  & ~n26535;
  assign n26537 = ~n26534 & ~n26535;
  assign n26538 = ~n26536 & ~n26537;
  assign n26539 = n26527 & ~n26538;
  assign n26540 = n26527 & ~n26539;
  assign n26541 = ~n26538 & ~n26539;
  assign n26542 = ~n26540 & ~n26541;
  assign n26543 = ~n26423 & ~n26436;
  assign n26544 = n26542 & n26543;
  assign n26545 = ~n26542 & ~n26543;
  assign n26546 = ~n26544 & ~n26545;
  assign n26547 = ~n26448 & ~n26451;
  assign n26548 = ~n26546 & n26547;
  assign n26549 = n26546 & ~n26547;
  assign n26550 = ~n26548 & ~n26549;
  assign n26551 = ~n26457 & ~n26460;
  assign n26552 = n26550 & ~n26551;
  assign n26553 = ~n26550 & n26551;
  assign po114  = ~n26552 & ~n26553;
  assign n26555 = ~n26522 & ~n26525;
  assign n26556 = n10394 & n12943;
  assign n26557 = pi123  & n10744;
  assign n26558 = pi125  & n10392;
  assign n26559 = pi124  & n10387;
  assign n26560 = ~n26558 & ~n26559;
  assign n26561 = ~n26557 & n26560;
  assign n26562 = ~n26556 & n26561;
  assign n26563 = pi56  & ~n26562;
  assign n26564 = pi56  & ~n26563;
  assign n26565 = ~n26562 & ~n26563;
  assign n26566 = ~n26564 & ~n26565;
  assign n26567 = ~n26515 & ~n26519;
  assign n26568 = n11488 & n11778;
  assign n26569 = pi120  & n11847;
  assign n26570 = pi122  & n11486;
  assign n26571 = pi121  & n11481;
  assign n26572 = ~n26570 & ~n26571;
  assign n26573 = ~n26569 & n26572;
  assign n26574 = ~n26568 & n26573;
  assign n26575 = pi59  & ~n26574;
  assign n26576 = pi59  & ~n26575;
  assign n26577 = ~n26574 & ~n26575;
  assign n26578 = ~n26576 & ~n26577;
  assign n26579 = ~n26508 & ~n26512;
  assign n26580 = pi115  & n13835;
  assign n26581 = pi116  & ~n13434;
  assign n26582 = ~n26580 & ~n26581;
  assign n26583 = ~n26502 & ~n26505;
  assign n26584 = ~n26582 & n26583;
  assign n26585 = n26582 & ~n26583;
  assign n26586 = ~n26584 & ~n26585;
  assign n26587 = n10667 & n12627;
  assign n26588 = pi117  & n13004;
  assign n26589 = pi119  & n12625;
  assign n26590 = pi118  & n12620;
  assign n26591 = ~n26589 & ~n26590;
  assign n26592 = ~n26588 & n26591;
  assign n26593 = ~n26587 & n26592;
  assign n26594 = pi62  & ~n26593;
  assign n26595 = pi62  & ~n26594;
  assign n26596 = ~n26593 & ~n26594;
  assign n26597 = ~n26595 & ~n26596;
  assign n26598 = ~n26586 & n26597;
  assign n26599 = n26586 & ~n26597;
  assign n26600 = ~n26598 & ~n26599;
  assign n26601 = ~n26579 & n26600;
  assign n26602 = n26579 & ~n26600;
  assign n26603 = ~n26601 & ~n26602;
  assign n26604 = ~n26578 & n26603;
  assign n26605 = n26578 & ~n26603;
  assign n26606 = ~n26604 & ~n26605;
  assign n26607 = ~n26567 & n26606;
  assign n26608 = ~n26567 & ~n26607;
  assign n26609 = n26606 & ~n26607;
  assign n26610 = ~n26608 & ~n26609;
  assign n26611 = ~n26566 & ~n26610;
  assign n26612 = n26566 & n26610;
  assign n26613 = ~n26611 & ~n26612;
  assign n26614 = ~n26555 & n26613;
  assign n26615 = n26555 & ~n26613;
  assign n26616 = ~n26614 & ~n26615;
  assign n26617 = n9310 & ~n13773;
  assign n26618 = pi126  & n9701;
  assign n26619 = pi127  & n9303;
  assign n26620 = ~n26618 & ~n26619;
  assign n26621 = ~n26617 & n26620;
  assign n26622 = pi53  & ~n26621;
  assign n26623 = pi53  & ~n26622;
  assign n26624 = ~n26621 & ~n26622;
  assign n26625 = ~n26623 & ~n26624;
  assign n26626 = n26616 & ~n26625;
  assign n26627 = n26616 & ~n26626;
  assign n26628 = ~n26625 & ~n26626;
  assign n26629 = ~n26627 & ~n26628;
  assign n26630 = ~n26539 & ~n26545;
  assign n26631 = n26629 & n26630;
  assign n26632 = ~n26629 & ~n26630;
  assign n26633 = ~n26631 & ~n26632;
  assign n26634 = ~n26549 & ~n26552;
  assign n26635 = n26633 & ~n26634;
  assign n26636 = ~n26633 & n26634;
  assign po115  = ~n26635 & ~n26636;
  assign n26638 = ~n26601 & ~n26604;
  assign n26639 = ~n26585 & ~n26599;
  assign n26640 = pi116  & n13835;
  assign n26641 = pi117  & ~n13434;
  assign n26642 = ~n26640 & ~n26641;
  assign n26643 = n26582 & ~n26642;
  assign n26644 = ~n26582 & n26642;
  assign n26645 = ~n26643 & ~n26644;
  assign n26646 = ~n26639 & n26645;
  assign n26647 = ~n26639 & ~n26646;
  assign n26648 = ~n26644 & ~n26646;
  assign n26649 = ~n26643 & n26648;
  assign n26650 = ~n26647 & ~n26649;
  assign n26651 = n11028 & n12627;
  assign n26652 = pi118  & n13004;
  assign n26653 = pi120  & n12625;
  assign n26654 = pi119  & n12620;
  assign n26655 = ~n26653 & ~n26654;
  assign n26656 = ~n26652 & n26655;
  assign n26657 = ~n26651 & n26656;
  assign n26658 = pi62  & ~n26657;
  assign n26659 = pi62  & ~n26658;
  assign n26660 = ~n26657 & ~n26658;
  assign n26661 = ~n26659 & ~n26660;
  assign n26662 = ~n26650 & n26661;
  assign n26663 = n26650 & ~n26661;
  assign n26664 = ~n26662 & ~n26663;
  assign n26665 = n11488 & n12158;
  assign n26666 = pi121  & n11847;
  assign n26667 = pi123  & n11486;
  assign n26668 = pi122  & n11481;
  assign n26669 = ~n26667 & ~n26668;
  assign n26670 = ~n26666 & n26669;
  assign n26671 = ~n26665 & n26670;
  assign n26672 = pi59  & ~n26671;
  assign n26673 = pi59  & ~n26672;
  assign n26674 = ~n26671 & ~n26672;
  assign n26675 = ~n26673 & ~n26674;
  assign n26676 = ~n26664 & ~n26675;
  assign n26677 = n26664 & n26675;
  assign n26678 = ~n26676 & ~n26677;
  assign n26679 = n26638 & ~n26678;
  assign n26680 = ~n26638 & n26678;
  assign n26681 = ~n26679 & ~n26680;
  assign n26682 = n10394 & n13344;
  assign n26683 = pi124  & n10744;
  assign n26684 = pi126  & n10392;
  assign n26685 = pi125  & n10387;
  assign n26686 = ~n26684 & ~n26685;
  assign n26687 = ~n26683 & n26686;
  assign n26688 = ~n26682 & n26687;
  assign n26689 = pi56  & ~n26688;
  assign n26690 = pi56  & ~n26689;
  assign n26691 = ~n26688 & ~n26689;
  assign n26692 = ~n26690 & ~n26691;
  assign n26693 = n26681 & ~n26692;
  assign n26694 = n26681 & ~n26693;
  assign n26695 = ~n26692 & ~n26693;
  assign n26696 = ~n26694 & ~n26695;
  assign n26697 = ~n26607 & ~n26611;
  assign n26698 = pi127  & n9701;
  assign n26699 = ~n9310 & ~n26698;
  assign n26700 = ~n13770 & ~n26698;
  assign n26701 = ~n26699 & ~n26700;
  assign n26702 = pi53  & ~n26701;
  assign n26703 = ~pi53  & n26701;
  assign n26704 = ~n26702 & ~n26703;
  assign n26705 = ~n26697 & ~n26704;
  assign n26706 = n26697 & n26704;
  assign n26707 = ~n26705 & ~n26706;
  assign n26708 = ~n26696 & n26707;
  assign n26709 = ~n26696 & ~n26708;
  assign n26710 = n26707 & ~n26708;
  assign n26711 = ~n26709 & ~n26710;
  assign n26712 = ~n26614 & ~n26626;
  assign n26713 = n26711 & n26712;
  assign n26714 = ~n26711 & ~n26712;
  assign n26715 = ~n26713 & ~n26714;
  assign n26716 = ~n26632 & ~n26635;
  assign n26717 = n26715 & ~n26716;
  assign n26718 = ~n26715 & n26716;
  assign po116  = ~n26717 & ~n26718;
  assign n26720 = ~n26714 & ~n26717;
  assign n26721 = ~n26705 & ~n26708;
  assign n26722 = ~n26680 & ~n26693;
  assign n26723 = n10394 & n13742;
  assign n26724 = pi125  & n10744;
  assign n26725 = pi127  & n10392;
  assign n26726 = pi126  & n10387;
  assign n26727 = ~n26725 & ~n26726;
  assign n26728 = ~n26724 & n26727;
  assign n26729 = ~n26723 & n26728;
  assign n26730 = pi56  & ~n26729;
  assign n26731 = pi56  & ~n26730;
  assign n26732 = ~n26729 & ~n26730;
  assign n26733 = ~n26731 & ~n26732;
  assign n26734 = ~n26722 & ~n26733;
  assign n26735 = ~n26722 & ~n26734;
  assign n26736 = ~n26733 & ~n26734;
  assign n26737 = ~n26735 & ~n26736;
  assign n26738 = ~n26650 & ~n26661;
  assign n26739 = ~n26676 & ~n26738;
  assign n26740 = n11488 & n12189;
  assign n26741 = pi122  & n11847;
  assign n26742 = pi124  & n11486;
  assign n26743 = pi123  & n11481;
  assign n26744 = ~n26742 & ~n26743;
  assign n26745 = ~n26741 & n26744;
  assign n26746 = ~n26740 & n26745;
  assign n26747 = pi59  & ~n26746;
  assign n26748 = pi59  & ~n26747;
  assign n26749 = ~n26746 & ~n26747;
  assign n26750 = ~n26748 & ~n26749;
  assign n26751 = pi53  & ~n26642;
  assign n26752 = ~pi53  & n26642;
  assign n26753 = ~n26751 & ~n26752;
  assign n26754 = pi117  & n13835;
  assign n26755 = pi118  & ~n13434;
  assign n26756 = ~n26754 & ~n26755;
  assign n26757 = n26753 & n26756;
  assign n26758 = ~n26753 & ~n26756;
  assign n26759 = ~n26757 & ~n26758;
  assign n26760 = n11389 & n12627;
  assign n26761 = pi119  & n13004;
  assign n26762 = pi121  & n12625;
  assign n26763 = pi120  & n12620;
  assign n26764 = ~n26762 & ~n26763;
  assign n26765 = ~n26761 & n26764;
  assign n26766 = ~n26760 & n26765;
  assign n26767 = pi62  & ~n26766;
  assign n26768 = pi62  & ~n26767;
  assign n26769 = ~n26766 & ~n26767;
  assign n26770 = ~n26768 & ~n26769;
  assign n26771 = n26759 & ~n26770;
  assign n26772 = n26759 & ~n26771;
  assign n26773 = ~n26770 & ~n26771;
  assign n26774 = ~n26772 & ~n26773;
  assign n26775 = ~n26648 & ~n26774;
  assign n26776 = n26648 & n26774;
  assign n26777 = ~n26775 & ~n26776;
  assign n26778 = ~n26750 & n26777;
  assign n26779 = ~n26750 & ~n26778;
  assign n26780 = n26777 & ~n26778;
  assign n26781 = ~n26779 & ~n26780;
  assign n26782 = ~n26739 & ~n26781;
  assign n26783 = ~n26739 & ~n26782;
  assign n26784 = ~n26781 & ~n26782;
  assign n26785 = ~n26783 & ~n26784;
  assign n26786 = ~n26737 & n26785;
  assign n26787 = n26737 & ~n26785;
  assign n26788 = ~n26786 & ~n26787;
  assign n26789 = ~n26721 & ~n26788;
  assign n26790 = n26721 & n26788;
  assign n26791 = ~n26789 & ~n26790;
  assign n26792 = ~n26720 & n26791;
  assign n26793 = n26720 & ~n26791;
  assign po117  = ~n26792 & ~n26793;
  assign n26795 = ~n26778 & ~n26782;
  assign n26796 = n11488 & n12943;
  assign n26797 = pi123  & n11847;
  assign n26798 = pi125  & n11486;
  assign n26799 = pi124  & n11481;
  assign n26800 = ~n26798 & ~n26799;
  assign n26801 = ~n26797 & n26800;
  assign n26802 = ~n26796 & n26801;
  assign n26803 = pi59  & ~n26802;
  assign n26804 = pi59  & ~n26803;
  assign n26805 = ~n26802 & ~n26803;
  assign n26806 = ~n26804 & ~n26805;
  assign n26807 = ~n26771 & ~n26775;
  assign n26808 = pi118  & n13835;
  assign n26809 = pi119  & ~n13434;
  assign n26810 = ~n26808 & ~n26809;
  assign n26811 = ~pi53  & ~n26642;
  assign n26812 = ~n26758 & ~n26811;
  assign n26813 = n26810 & ~n26812;
  assign n26814 = ~n26810 & n26812;
  assign n26815 = ~n26813 & ~n26814;
  assign n26816 = pi120  & n13004;
  assign n26817 = pi122  & n12625;
  assign n26818 = pi121  & n12620;
  assign n26819 = ~n26817 & ~n26818;
  assign n26820 = ~n26816 & n26819;
  assign n26821 = ~n12627 & n26820;
  assign n26822 = ~n11778 & n26820;
  assign n26823 = ~n26821 & ~n26822;
  assign n26824 = pi62  & ~n26823;
  assign n26825 = ~pi62  & n26823;
  assign n26826 = ~n26824 & ~n26825;
  assign n26827 = n26815 & ~n26826;
  assign n26828 = ~n26815 & n26826;
  assign n26829 = ~n26827 & ~n26828;
  assign n26830 = ~n26807 & n26829;
  assign n26831 = ~n26807 & ~n26830;
  assign n26832 = n26829 & ~n26830;
  assign n26833 = ~n26831 & ~n26832;
  assign n26834 = ~n26806 & ~n26833;
  assign n26835 = n26806 & n26833;
  assign n26836 = ~n26834 & ~n26835;
  assign n26837 = ~n26795 & n26836;
  assign n26838 = n26795 & ~n26836;
  assign n26839 = ~n26837 & ~n26838;
  assign n26840 = n10394 & ~n13773;
  assign n26841 = pi126  & n10744;
  assign n26842 = pi127  & n10387;
  assign n26843 = ~n26841 & ~n26842;
  assign n26844 = ~n26840 & n26843;
  assign n26845 = pi56  & ~n26844;
  assign n26846 = pi56  & ~n26845;
  assign n26847 = ~n26844 & ~n26845;
  assign n26848 = ~n26846 & ~n26847;
  assign n26849 = n26839 & ~n26848;
  assign n26850 = n26839 & ~n26849;
  assign n26851 = ~n26848 & ~n26849;
  assign n26852 = ~n26850 & ~n26851;
  assign n26853 = ~n26737 & ~n26785;
  assign n26854 = ~n26734 & ~n26853;
  assign n26855 = ~n26852 & ~n26854;
  assign n26856 = ~n26852 & ~n26855;
  assign n26857 = ~n26854 & ~n26855;
  assign n26858 = ~n26856 & ~n26857;
  assign n26859 = ~n26789 & ~n26792;
  assign n26860 = ~n26858 & ~n26859;
  assign n26861 = n26858 & n26859;
  assign po118  = ~n26860 & ~n26861;
  assign n26863 = n12158 & n12627;
  assign n26864 = pi121  & n13004;
  assign n26865 = pi123  & n12625;
  assign n26866 = pi122  & n12620;
  assign n26867 = ~n26865 & ~n26866;
  assign n26868 = ~n26864 & n26867;
  assign n26869 = ~n26863 & n26868;
  assign n26870 = pi62  & ~n26869;
  assign n26871 = pi62  & ~n26870;
  assign n26872 = ~n26869 & ~n26870;
  assign n26873 = ~n26871 & ~n26872;
  assign n26874 = pi119  & n13835;
  assign n26875 = pi120  & ~n13434;
  assign n26876 = ~n26874 & ~n26875;
  assign n26877 = n26810 & ~n26876;
  assign n26878 = n26810 & ~n26877;
  assign n26879 = ~n26876 & ~n26877;
  assign n26880 = ~n26878 & ~n26879;
  assign n26881 = ~n26873 & ~n26880;
  assign n26882 = ~n26873 & ~n26881;
  assign n26883 = ~n26880 & ~n26881;
  assign n26884 = ~n26882 & ~n26883;
  assign n26885 = ~n26813 & ~n26827;
  assign n26886 = n26884 & n26885;
  assign n26887 = ~n26884 & ~n26885;
  assign n26888 = ~n26886 & ~n26887;
  assign n26889 = n11488 & n13344;
  assign n26890 = pi124  & n11847;
  assign n26891 = pi126  & n11486;
  assign n26892 = pi125  & n11481;
  assign n26893 = ~n26891 & ~n26892;
  assign n26894 = ~n26890 & n26893;
  assign n26895 = ~n26889 & n26894;
  assign n26896 = pi59  & ~n26895;
  assign n26897 = pi59  & ~n26896;
  assign n26898 = ~n26895 & ~n26896;
  assign n26899 = ~n26897 & ~n26898;
  assign n26900 = n26888 & ~n26899;
  assign n26901 = n26888 & ~n26900;
  assign n26902 = ~n26899 & ~n26900;
  assign n26903 = ~n26901 & ~n26902;
  assign n26904 = ~n26830 & ~n26834;
  assign n26905 = pi127  & n10744;
  assign n26906 = ~n10394 & ~n26905;
  assign n26907 = ~n13770 & ~n26905;
  assign n26908 = ~n26906 & ~n26907;
  assign n26909 = pi56  & ~n26908;
  assign n26910 = ~pi56  & n26908;
  assign n26911 = ~n26909 & ~n26910;
  assign n26912 = ~n26904 & ~n26911;
  assign n26913 = n26904 & n26911;
  assign n26914 = ~n26912 & ~n26913;
  assign n26915 = ~n26903 & n26914;
  assign n26916 = ~n26903 & ~n26915;
  assign n26917 = n26914 & ~n26915;
  assign n26918 = ~n26916 & ~n26917;
  assign n26919 = ~n26837 & ~n26849;
  assign n26920 = n26918 & n26919;
  assign n26921 = ~n26918 & ~n26919;
  assign n26922 = ~n26920 & ~n26921;
  assign n26923 = ~n26855 & ~n26860;
  assign n26924 = n26922 & ~n26923;
  assign n26925 = ~n26922 & n26923;
  assign po119  = ~n26924 & ~n26925;
  assign n26927 = ~n26887 & ~n26900;
  assign n26928 = n11488 & n13742;
  assign n26929 = pi125  & n11847;
  assign n26930 = pi127  & n11486;
  assign n26931 = pi126  & n11481;
  assign n26932 = ~n26930 & ~n26931;
  assign n26933 = ~n26929 & n26932;
  assign n26934 = ~n26928 & n26933;
  assign n26935 = pi59  & ~n26934;
  assign n26936 = pi59  & ~n26935;
  assign n26937 = ~n26934 & ~n26935;
  assign n26938 = ~n26936 & ~n26937;
  assign n26939 = ~n26927 & ~n26938;
  assign n26940 = ~n26927 & ~n26939;
  assign n26941 = ~n26938 & ~n26939;
  assign n26942 = ~n26940 & ~n26941;
  assign n26943 = pi120  & n13835;
  assign n26944 = pi121  & ~n13434;
  assign n26945 = ~n26943 & ~n26944;
  assign n26946 = ~pi56  & ~n26945;
  assign n26947 = ~pi56  & ~n26946;
  assign n26948 = ~n26945 & ~n26946;
  assign n26949 = ~n26947 & ~n26948;
  assign n26950 = ~n26810 & ~n26949;
  assign n26951 = ~n26810 & ~n26950;
  assign n26952 = ~n26949 & ~n26950;
  assign n26953 = ~n26951 & ~n26952;
  assign n26954 = ~n26877 & ~n26881;
  assign n26955 = n26953 & n26954;
  assign n26956 = ~n26953 & ~n26954;
  assign n26957 = ~n26955 & ~n26956;
  assign n26958 = n12189 & n12627;
  assign n26959 = pi122  & n13004;
  assign n26960 = pi124  & n12625;
  assign n26961 = pi123  & n12620;
  assign n26962 = ~n26960 & ~n26961;
  assign n26963 = ~n26959 & n26962;
  assign n26964 = ~n26958 & n26963;
  assign n26965 = pi62  & ~n26964;
  assign n26966 = pi62  & ~n26965;
  assign n26967 = ~n26964 & ~n26965;
  assign n26968 = ~n26966 & ~n26967;
  assign n26969 = n26957 & ~n26968;
  assign n26970 = ~n26957 & n26968;
  assign n26971 = ~n26969 & ~n26970;
  assign n26972 = ~n26942 & n26971;
  assign n26973 = ~n26942 & ~n26972;
  assign n26974 = n26971 & ~n26972;
  assign n26975 = ~n26973 & ~n26974;
  assign n26976 = ~n26912 & ~n26915;
  assign n26977 = n26975 & n26976;
  assign n26978 = ~n26975 & ~n26976;
  assign n26979 = ~n26977 & ~n26978;
  assign n26980 = ~n26921 & ~n26924;
  assign n26981 = n26979 & ~n26980;
  assign n26982 = ~n26979 & n26980;
  assign po120  = ~n26981 & ~n26982;
  assign n26984 = ~n26956 & ~n26969;
  assign n26985 = pi121  & n13835;
  assign n26986 = pi122  & ~n13434;
  assign n26987 = ~n26985 & ~n26986;
  assign n26988 = ~n26946 & ~n26950;
  assign n26989 = ~n26987 & n26988;
  assign n26990 = n26987 & ~n26988;
  assign n26991 = ~n26989 & ~n26990;
  assign n26992 = pi123  & n13004;
  assign n26993 = pi125  & n12625;
  assign n26994 = pi124  & n12620;
  assign n26995 = ~n26993 & ~n26994;
  assign n26996 = ~n26992 & n26995;
  assign n26997 = ~n12627 & n26996;
  assign n26998 = ~n12943 & n26996;
  assign n26999 = ~n26997 & ~n26998;
  assign n27000 = pi62  & ~n26999;
  assign n27001 = ~pi62  & n26999;
  assign n27002 = ~n27000 & ~n27001;
  assign n27003 = n26991 & ~n27002;
  assign n27004 = ~n26991 & n27002;
  assign n27005 = ~n27003 & ~n27004;
  assign n27006 = ~n26984 & n27005;
  assign n27007 = n26984 & ~n27005;
  assign n27008 = ~n27006 & ~n27007;
  assign n27009 = n11488 & ~n13773;
  assign n27010 = pi126  & n11847;
  assign n27011 = pi127  & n11481;
  assign n27012 = ~n27010 & ~n27011;
  assign n27013 = ~n27009 & n27012;
  assign n27014 = pi59  & ~n27013;
  assign n27015 = pi59  & ~n27014;
  assign n27016 = ~n27013 & ~n27014;
  assign n27017 = ~n27015 & ~n27016;
  assign n27018 = n27008 & ~n27017;
  assign n27019 = n27008 & ~n27018;
  assign n27020 = ~n27017 & ~n27018;
  assign n27021 = ~n27019 & ~n27020;
  assign n27022 = ~n26939 & ~n26972;
  assign n27023 = n27021 & n27022;
  assign n27024 = ~n27021 & ~n27022;
  assign n27025 = ~n27023 & ~n27024;
  assign n27026 = ~n26978 & ~n26981;
  assign n27027 = n27025 & ~n27026;
  assign n27028 = ~n27025 & n27026;
  assign po121  = ~n27027 & ~n27028;
  assign n27030 = ~n27024 & ~n27027;
  assign n27031 = ~n27006 & ~n27018;
  assign n27032 = ~n26990 & ~n27003;
  assign n27033 = pi122  & n13835;
  assign n27034 = pi123  & ~n13434;
  assign n27035 = ~n27033 & ~n27034;
  assign n27036 = n26987 & ~n27035;
  assign n27037 = ~n26987 & n27035;
  assign n27038 = ~n27036 & ~n27037;
  assign n27039 = ~n27032 & n27038;
  assign n27040 = ~n27032 & ~n27039;
  assign n27041 = ~n27037 & ~n27039;
  assign n27042 = ~n27036 & n27041;
  assign n27043 = ~n27040 & ~n27042;
  assign n27044 = n12627 & n13344;
  assign n27045 = pi124  & n13004;
  assign n27046 = pi126  & n12625;
  assign n27047 = pi125  & n12620;
  assign n27048 = ~n27046 & ~n27047;
  assign n27049 = ~n27045 & n27048;
  assign n27050 = ~n27044 & n27049;
  assign n27051 = pi62  & ~n27050;
  assign n27052 = pi62  & ~n27051;
  assign n27053 = ~n27050 & ~n27051;
  assign n27054 = ~n27052 & ~n27053;
  assign n27055 = pi127  & n11847;
  assign n27056 = n11488 & n13770;
  assign n27057 = ~n27055 & ~n27056;
  assign n27058 = pi59  & ~n27057;
  assign n27059 = pi59  & ~n27058;
  assign n27060 = ~n27057 & ~n27058;
  assign n27061 = ~n27059 & ~n27060;
  assign n27062 = ~n27054 & ~n27061;
  assign n27063 = ~n27054 & ~n27062;
  assign n27064 = ~n27061 & ~n27062;
  assign n27065 = ~n27063 & ~n27064;
  assign n27066 = ~n27043 & n27065;
  assign n27067 = n27043 & ~n27065;
  assign n27068 = ~n27066 & ~n27067;
  assign n27069 = ~n27031 & ~n27068;
  assign n27070 = ~n27031 & ~n27069;
  assign n27071 = ~n27068 & ~n27069;
  assign n27072 = ~n27070 & ~n27071;
  assign n27073 = ~n27030 & ~n27072;
  assign n27074 = n27030 & n27072;
  assign po122  = ~n27073 & ~n27074;
  assign n27076 = ~n27069 & ~n27073;
  assign n27077 = ~n27043 & ~n27065;
  assign n27078 = ~n27062 & ~n27077;
  assign n27079 = pi59  & ~n27035;
  assign n27080 = ~pi59  & n27035;
  assign n27081 = ~n27079 & ~n27080;
  assign n27082 = pi123  & n13835;
  assign n27083 = pi124  & ~n13434;
  assign n27084 = ~n27082 & ~n27083;
  assign n27085 = n27081 & n27084;
  assign n27086 = ~n27081 & ~n27084;
  assign n27087 = ~n27085 & ~n27086;
  assign n27088 = n12627 & n13742;
  assign n27089 = pi125  & n13004;
  assign n27090 = pi127  & n12625;
  assign n27091 = pi126  & n12620;
  assign n27092 = ~n27090 & ~n27091;
  assign n27093 = ~n27089 & n27092;
  assign n27094 = ~n27088 & n27093;
  assign n27095 = pi62  & ~n27094;
  assign n27096 = pi62  & ~n27095;
  assign n27097 = ~n27094 & ~n27095;
  assign n27098 = ~n27096 & ~n27097;
  assign n27099 = n27087 & ~n27098;
  assign n27100 = n27087 & ~n27099;
  assign n27101 = ~n27098 & ~n27099;
  assign n27102 = ~n27100 & ~n27101;
  assign n27103 = ~n27041 & ~n27102;
  assign n27104 = n27041 & n27102;
  assign n27105 = ~n27103 & ~n27104;
  assign n27106 = ~n27078 & n27105;
  assign n27107 = ~n27078 & ~n27106;
  assign n27108 = n27105 & ~n27106;
  assign n27109 = ~n27107 & ~n27108;
  assign n27110 = ~n27076 & ~n27109;
  assign n27111 = n27076 & n27109;
  assign po123  = ~n27110 & ~n27111;
  assign n27113 = ~n27106 & ~n27110;
  assign n27114 = ~n27099 & ~n27103;
  assign n27115 = pi124  & n13835;
  assign n27116 = pi125  & ~n13434;
  assign n27117 = ~n27115 & ~n27116;
  assign n27118 = ~pi59  & ~n27035;
  assign n27119 = ~n27086 & ~n27118;
  assign n27120 = n27117 & ~n27119;
  assign n27121 = ~n27117 & n27119;
  assign n27122 = ~n27120 & ~n27121;
  assign n27123 = pi126  & n13004;
  assign n27124 = pi127  & n12620;
  assign n27125 = ~n27123 & ~n27124;
  assign n27126 = ~n12627 & n27125;
  assign n27127 = n13773 & n27125;
  assign n27128 = ~n27126 & ~n27127;
  assign n27129 = pi62  & ~n27128;
  assign n27130 = ~pi62  & n27128;
  assign n27131 = ~n27129 & ~n27130;
  assign n27132 = n27122 & ~n27131;
  assign n27133 = ~n27122 & n27131;
  assign n27134 = ~n27132 & ~n27133;
  assign n27135 = ~n27114 & n27134;
  assign n27136 = ~n27114 & ~n27135;
  assign n27137 = n27134 & ~n27135;
  assign n27138 = ~n27136 & ~n27137;
  assign n27139 = ~n27113 & ~n27138;
  assign n27140 = n27113 & n27138;
  assign po124  = ~n27139 & ~n27140;
  assign n27142 = ~n27135 & ~n27139;
  assign n27143 = ~n27120 & ~n27132;
  assign n27144 = pi125  & n13835;
  assign n27145 = pi126  & ~n13434;
  assign n27146 = ~n27144 & ~n27145;
  assign n27147 = n27117 & ~n27146;
  assign n27148 = ~n27117 & n27146;
  assign n27149 = ~n27147 & ~n27148;
  assign n27150 = pi127  & n13004;
  assign n27151 = ~n12627 & ~n27150;
  assign n27152 = ~n13770 & ~n27150;
  assign n27153 = ~n27151 & ~n27152;
  assign n27154 = pi62  & ~n27153;
  assign n27155 = ~pi62  & n27153;
  assign n27156 = ~n27154 & ~n27155;
  assign n27157 = n27149 & ~n27156;
  assign n27158 = ~n27149 & n27156;
  assign n27159 = ~n27157 & ~n27158;
  assign n27160 = ~n27143 & n27159;
  assign n27161 = ~n27143 & ~n27160;
  assign n27162 = n27159 & ~n27160;
  assign n27163 = ~n27161 & ~n27162;
  assign n27164 = ~n27142 & ~n27163;
  assign n27165 = n27142 & n27163;
  assign po125  = ~n27164 & ~n27165;
  assign n27167 = ~n27160 & ~n27164;
  assign n27168 = ~n27147 & ~n27157;
  assign n27169 = pi126  & n13835;
  assign n27170 = pi127  & ~n13434;
  assign n27171 = ~n27169 & ~n27170;
  assign n27172 = ~pi62  & ~n27171;
  assign n27173 = pi62  & n27171;
  assign n27174 = ~n27172 & ~n27173;
  assign n27175 = ~n27117 & n27174;
  assign n27176 = n27117 & ~n27174;
  assign n27177 = ~n27175 & ~n27176;
  assign n27178 = ~n27168 & n27177;
  assign n27179 = n27168 & ~n27177;
  assign n27180 = ~n27178 & ~n27179;
  assign n27181 = ~n27167 & n27180;
  assign n27182 = n27167 & ~n27180;
  assign po126  = ~n27181 & ~n27182;
  assign n27184 = ~n27172 & ~n27175;
  assign n27185 = pi127  & n13835;
  assign n27186 = ~n27184 & n27185;
  assign n27187 = n27184 & ~n27185;
  assign n27188 = ~n27186 & ~n27187;
  assign n27189 = ~n27178 & ~n27181;
  assign n27190 = n27188 & n27189;
  assign n27191 = ~n27188 & ~n27189;
  assign po127  = ~n27190 & ~n27191;
endmodule
