module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 ,
    pi7 , pi8 , pi9 , pi10 , pi11 , pi12 ,
    pi13 , pi14 , pi15 , pi16 , pi17 , pi18 ,
    pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 ,
    pi31 , pi32 , pi33 , pi34 , pi35 , pi36 ,
    pi37 , pi38 , pi39 , pi40 , pi41 , pi42 ,
    pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 ,
    pi55 , pi56 , pi57 , pi58 , pi59 , pi60 ,
    pi61 , pi62 , pi63 , pi64 , pi65 , pi66 ,
    pi67 , pi68 , pi69 , pi70 , pi71 , pi72 ,
    pi73 , pi74 , pi75 , pi76 , pi77 , pi78 ,
    pi79 , pi80 , pi81 , pi82 , pi83 , pi84 ,
    pi85 , pi86 , pi87 , pi88 , pi89 , pi90 ,
    pi91 , pi92 , pi93 , pi94 , pi95 , pi96 ,
    pi97 , pi98 , pi99 , pi100 , pi101 , pi102 ,
    pi103 , pi104 , pi105 , pi106 , pi107 , pi108 ,
    pi109 , pi110 , pi111 , pi112 , pi113 , pi114 ,
    pi115 , pi116 , pi117 , pi118 , pi119 , pi120 ,
    pi121 , pi122 , pi123 , pi124 , pi125 , pi126 ,
    pi127 , pi128 , pi129 , pi130 , pi131 , pi132 , pi133 ,
    pi134 , pi135 , pi136 , pi137 , pi138 , pi139 ,
    pi140 , pi141 , pi142 , pi143 , pi144 , pi145 ,
    pi146 , pi147 , pi148 , pi149 , pi150 , pi151 ,
    pi152 , pi153 , pi154 , pi155 , pi156 , pi157 ,
    pi158 , pi159 , pi160 , pi161 , pi162 , pi163 ,
    pi164 , pi165 , pi166 , pi167 , pi168 , pi169 ,
    pi170 , pi171 , pi172 , pi173 , pi174 , pi175 ,
    pi176 , pi177 , pi178 , pi179 , pi180 , pi181 ,
    pi182 , pi183 , pi184 , pi185 , pi186 , pi187 ,
    pi188 , pi189 , pi190 , pi191 , pi192 , pi193 ,
    pi194 , pi195 , pi196 , pi197 , pi198 , pi199 ,
    pi200 , pi201 , pi202 , pi203 , pi204 , pi205 ,
    pi206 , pi207 , pi208 , pi209 , pi210 , pi211 ,
    pi212 , pi213 , pi214 , pi215 , pi216 , pi217 ,
    pi218 , pi219 , pi220 , pi221 , pi222 , pi223 ,
    pi224 , pi225 , pi226 , pi227 , pi228 , pi229 ,
    pi230 , pi231 , pi232 , pi233 , pi234 , pi235 ,
    pi236 , pi237 , pi238 , pi239 , pi240 , pi241 ,
    pi242 , pi243 , pi244 , pi245 , pi246 , pi247 ,
    pi248 , pi249 , pi250 , pi251 , pi252 , pi253 ,
    pi254 , pi255 , pi256 , pi257 , pi258 , pi259 ,
    pi260 , pi261 , pi262 , pi263 , pi264 , pi265 , pi266 ,
    pi267 , pi268 , pi269 , pi270 , pi271 , pi272 ,
    pi273 , pi274 , pi275 , pi276 , pi277 , pi278 ,
    pi279 , pi280 , pi281 , pi282 , pi283 , pi284 ,
    pi285 , pi286 , pi287 , pi288 , pi289 , pi290 ,
    pi291 , pi292 , pi293 , pi294 , pi295 , pi296 ,
    pi297 , pi298 , pi299 , pi300 , pi301 , pi302 ,
    pi303 , pi304 , pi305 , pi306 , pi307 , pi308 ,
    pi309 , pi310 , pi311 , pi312 , pi313 , pi314 ,
    pi315 , pi316 , pi317 , pi318 , pi319 , pi320 ,
    pi321 , pi322 , pi323 , pi324 , pi325 , pi326 ,
    pi327 , pi328 , pi329 , pi330 , pi331 , pi332 ,
    pi333 , pi334 , pi335 , pi336 , pi337 , pi338 ,
    pi339 , pi340 , pi341 , pi342 , pi343 , pi344 ,
    pi345 , pi346 , pi347 , pi348 , pi349 , pi350 ,
    pi351 , pi352 , pi353 , pi354 , pi355 , pi356 ,
    pi357 , pi358 , pi359 , pi360 , pi361 , pi362 ,
    pi363 , pi364 , pi365 , pi366 , pi367 , pi368 ,
    pi369 , pi370 , pi371 , pi372 , pi373 , pi374 ,
    pi375 , pi376 , pi377 , pi378 , pi379 , pi380 ,
    pi381 , pi382 , pi383 , pi384 , pi385 , pi386 ,
    pi387 , pi388 , pi389 , pi390 , pi391 , pi392 , pi393 ,
    pi394 , pi395 , pi396 , pi397 , pi398 , pi399 ,
    pi400 , pi401 , pi402 , pi403 , pi404 , pi405 ,
    pi406 , pi407 , pi408 , pi409 , pi410 , pi411 ,
    pi412 , pi413 , pi414 , pi415 , pi416 , pi417 ,
    pi418 , pi419 , pi420 , pi421 , pi422 , pi423 ,
    pi424 , pi425 , pi426 , pi427 , pi428 , pi429 ,
    pi430 , pi431 , pi432 , pi433 , pi434 , pi435 ,
    pi436 , pi437 , pi438 , pi439 , pi440 , pi441 ,
    pi442 , pi443 , pi444 , pi445 , pi446 , pi447 ,
    pi448 , pi449 , pi450 , pi451 , pi452 , pi453 ,
    pi454 , pi455 , pi456 , pi457 , pi458 , pi459 ,
    pi460 , pi461 , pi462 , pi463 , pi464 , pi465 ,
    pi466 , pi467 , pi468 , pi469 , pi470 , pi471 ,
    pi472 , pi473 , pi474 , pi475 , pi476 , pi477 ,
    pi478 , pi479 , pi480 , pi481 , pi482 , pi483 ,
    pi484 , pi485 , pi486 , pi487 , pi488 , pi489 ,
    pi490 , pi491 , pi492 , pi493 , pi494 , pi495 ,
    pi496 , pi497 , pi498 , pi499 , pi500 , pi501 ,
    pi502 , pi503 , pi504 , pi505 , pi506 , pi507 ,
    pi508 , pi509 , pi510 , pi511 ,
    po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 , po14 ,
    po15 , po16 , po17 , po18 , po19 ,
    po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 ,
    po30 , po31 , po32 , po33 , po34 ,
    po35 , po36 , po37 , po38 , po39 ,
    po40 , po41 , po42 , po43 , po44 ,
    po45 , po46 , po47 , po48 , po49 ,
    po50 , po51 , po52 , po53 , po54 ,
    po55 , po56 , po57 , po58 , po59 ,
    po60 , po61 , po62 , po63 , po64 ,
    po65 , po66 , po67 , po68 , po69 ,
    po70 , po71 , po72 , po73 , po74 ,
    po75 , po76 , po77 , po78 , po79 ,
    po80 , po81 , po82 , po83 , po84 ,
    po85 , po86 , po87 , po88 , po89 ,
    po90 , po91 , po92 , po93 , po94 ,
    po95 , po96 , po97 , po98 , po99 ,
    po100 , po101 , po102 , po103 ,
    po104 , po105 , po106 , po107 ,
    po108 , po109 , po110 , po111 ,
    po112 , po113 , po114 , po115 ,
    po116 , po117 , po118 , po119 ,
    po120 , po121 , po122 , po123 ,
    po124 , po125 , po126 , po127 ,
    po128 , po129   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 ,
    pi6 , pi7 , pi8 , pi9 , pi10 , pi11 ,
    pi12 , pi13 , pi14 , pi15 , pi16 , pi17 ,
    pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 ,
    pi30 , pi31 , pi32 , pi33 , pi34 , pi35 ,
    pi36 , pi37 , pi38 , pi39 , pi40 , pi41 ,
    pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 ,
    pi54 , pi55 , pi56 , pi57 , pi58 , pi59 ,
    pi60 , pi61 , pi62 , pi63 , pi64 , pi65 ,
    pi66 , pi67 , pi68 , pi69 , pi70 , pi71 ,
    pi72 , pi73 , pi74 , pi75 , pi76 , pi77 ,
    pi78 , pi79 , pi80 , pi81 , pi82 , pi83 ,
    pi84 , pi85 , pi86 , pi87 , pi88 , pi89 ,
    pi90 , pi91 , pi92 , pi93 , pi94 , pi95 ,
    pi96 , pi97 , pi98 , pi99 , pi100 , pi101 ,
    pi102 , pi103 , pi104 , pi105 , pi106 , pi107 ,
    pi108 , pi109 , pi110 , pi111 , pi112 , pi113 ,
    pi114 , pi115 , pi116 , pi117 , pi118 , pi119 ,
    pi120 , pi121 , pi122 , pi123 , pi124 , pi125 ,
    pi126 , pi127 , pi128 , pi129 , pi130 , pi131 ,
    pi132 , pi133 , pi134 , pi135 , pi136 , pi137 , pi138 ,
    pi139 , pi140 , pi141 , pi142 , pi143 , pi144 ,
    pi145 , pi146 , pi147 , pi148 , pi149 , pi150 ,
    pi151 , pi152 , pi153 , pi154 , pi155 , pi156 ,
    pi157 , pi158 , pi159 , pi160 , pi161 , pi162 ,
    pi163 , pi164 , pi165 , pi166 , pi167 , pi168 ,
    pi169 , pi170 , pi171 , pi172 , pi173 , pi174 ,
    pi175 , pi176 , pi177 , pi178 , pi179 , pi180 ,
    pi181 , pi182 , pi183 , pi184 , pi185 , pi186 ,
    pi187 , pi188 , pi189 , pi190 , pi191 , pi192 ,
    pi193 , pi194 , pi195 , pi196 , pi197 , pi198 ,
    pi199 , pi200 , pi201 , pi202 , pi203 , pi204 ,
    pi205 , pi206 , pi207 , pi208 , pi209 , pi210 ,
    pi211 , pi212 , pi213 , pi214 , pi215 , pi216 ,
    pi217 , pi218 , pi219 , pi220 , pi221 , pi222 ,
    pi223 , pi224 , pi225 , pi226 , pi227 , pi228 ,
    pi229 , pi230 , pi231 , pi232 , pi233 , pi234 ,
    pi235 , pi236 , pi237 , pi238 , pi239 , pi240 ,
    pi241 , pi242 , pi243 , pi244 , pi245 , pi246 ,
    pi247 , pi248 , pi249 , pi250 , pi251 , pi252 ,
    pi253 , pi254 , pi255 , pi256 , pi257 , pi258 ,
    pi259 , pi260 , pi261 , pi262 , pi263 , pi264 , pi265 ,
    pi266 , pi267 , pi268 , pi269 , pi270 , pi271 ,
    pi272 , pi273 , pi274 , pi275 , pi276 , pi277 ,
    pi278 , pi279 , pi280 , pi281 , pi282 , pi283 ,
    pi284 , pi285 , pi286 , pi287 , pi288 , pi289 ,
    pi290 , pi291 , pi292 , pi293 , pi294 , pi295 ,
    pi296 , pi297 , pi298 , pi299 , pi300 , pi301 ,
    pi302 , pi303 , pi304 , pi305 , pi306 , pi307 ,
    pi308 , pi309 , pi310 , pi311 , pi312 , pi313 ,
    pi314 , pi315 , pi316 , pi317 , pi318 , pi319 ,
    pi320 , pi321 , pi322 , pi323 , pi324 , pi325 ,
    pi326 , pi327 , pi328 , pi329 , pi330 , pi331 ,
    pi332 , pi333 , pi334 , pi335 , pi336 , pi337 ,
    pi338 , pi339 , pi340 , pi341 , pi342 , pi343 ,
    pi344 , pi345 , pi346 , pi347 , pi348 , pi349 ,
    pi350 , pi351 , pi352 , pi353 , pi354 , pi355 ,
    pi356 , pi357 , pi358 , pi359 , pi360 , pi361 ,
    pi362 , pi363 , pi364 , pi365 , pi366 , pi367 ,
    pi368 , pi369 , pi370 , pi371 , pi372 , pi373 ,
    pi374 , pi375 , pi376 , pi377 , pi378 , pi379 ,
    pi380 , pi381 , pi382 , pi383 , pi384 , pi385 ,
    pi386 , pi387 , pi388 , pi389 , pi390 , pi391 , pi392 ,
    pi393 , pi394 , pi395 , pi396 , pi397 , pi398 ,
    pi399 , pi400 , pi401 , pi402 , pi403 , pi404 ,
    pi405 , pi406 , pi407 , pi408 , pi409 , pi410 ,
    pi411 , pi412 , pi413 , pi414 , pi415 , pi416 ,
    pi417 , pi418 , pi419 , pi420 , pi421 , pi422 ,
    pi423 , pi424 , pi425 , pi426 , pi427 , pi428 ,
    pi429 , pi430 , pi431 , pi432 , pi433 , pi434 ,
    pi435 , pi436 , pi437 , pi438 , pi439 , pi440 ,
    pi441 , pi442 , pi443 , pi444 , pi445 , pi446 ,
    pi447 , pi448 , pi449 , pi450 , pi451 , pi452 ,
    pi453 , pi454 , pi455 , pi456 , pi457 , pi458 ,
    pi459 , pi460 , pi461 , pi462 , pi463 , pi464 ,
    pi465 , pi466 , pi467 , pi468 , pi469 , pi470 ,
    pi471 , pi472 , pi473 , pi474 , pi475 , pi476 ,
    pi477 , pi478 , pi479 , pi480 , pi481 , pi482 ,
    pi483 , pi484 , pi485 , pi486 , pi487 , pi488 ,
    pi489 , pi490 , pi491 , pi492 , pi493 , pi494 ,
    pi495 , pi496 , pi497 , pi498 , pi499 , pi500 ,
    pi501 , pi502 , pi503 , pi504 , pi505 , pi506 ,
    pi507 , pi508 , pi509 , pi510 , pi511 ;
  output po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 , po14 ,
    po15 , po16 , po17 , po18 , po19 ,
    po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 ,
    po30 , po31 , po32 , po33 , po34 ,
    po35 , po36 , po37 , po38 , po39 ,
    po40 , po41 , po42 , po43 , po44 ,
    po45 , po46 , po47 , po48 , po49 ,
    po50 , po51 , po52 , po53 , po54 ,
    po55 , po56 , po57 , po58 , po59 ,
    po60 , po61 , po62 , po63 , po64 ,
    po65 , po66 , po67 , po68 , po69 ,
    po70 , po71 , po72 , po73 , po74 ,
    po75 , po76 , po77 , po78 , po79 ,
    po80 , po81 , po82 , po83 , po84 ,
    po85 , po86 , po87 , po88 , po89 ,
    po90 , po91 , po92 , po93 , po94 ,
    po95 , po96 , po97 , po98 , po99 ,
    po100 , po101 , po102 , po103 ,
    po104 , po105 , po106 , po107 ,
    po108 , po109 , po110 , po111 ,
    po112 , po113 , po114 , po115 ,
    po116 , po117 , po118 , po119 ,
    po120 , po121 , po122 , po123 ,
    po124 , po125 , po126 , po127 ,
    po128 , po129 ;
  wire n643, n644, n645, n646, n647, n648, n649,
    n650, n651, n652, n653, n654, n655, n656,
    n657, n658, n659, n660, n661, n662, n663,
    n664, n665, n666, n667, n668, n669, n670,
    n671, n672, n673, n674, n675, n676, n677,
    n678, n679, n680, n681, n682, n683, n684,
    n685, n686, n687, n688, n689, n690, n691,
    n692, n693, n694, n695, n696, n697, n698,
    n699, n700, n701, n702, n703, n704, n705,
    n706, n707, n708, n709, n710, n711, n712,
    n713, n714, n715, n716, n717, n718, n719,
    n720, n721, n722, n723, n724, n725, n726,
    n727, n728, n729, n730, n731, n732, n733,
    n734, n735, n736, n737, n738, n739, n740,
    n741, n742, n743, n744, n745, n746, n747,
    n748, n749, n750, n751, n752, n753, n754,
    n755, n756, n757, n758, n759, n760, n761,
    n762, n763, n764, n765, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n775,
    n776, n777, n778, n779, n780, n781, n782,
    n783, n784, n785, n786, n787, n788, n789,
    n790, n791, n792, n793, n794, n795, n796,
    n797, n798, n799, n800, n801, n802, n803,
    n804, n805, n806, n807, n808, n809, n810,
    n811, n812, n813, n814, n815, n816, n817,
    n818, n819, n820, n821, n822, n823, n824,
    n825, n826, n827, n828, n829, n830, n831,
    n832, n833, n834, n835, n836, n837, n838,
    n839, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n851, n852,
    n853, n854, n855, n856, n857, n858, n859,
    n860, n861, n862, n863, n864, n865, n866,
    n867, n868, n869, n870, n871, n872, n873,
    n874, n875, n876, n877, n878, n879, n880,
    n881, n882, n883, n884, n885, n886, n887,
    n888, n889, n890, n891, n892, n893, n894,
    n895, n896, n897, n898, n899, n900, n901,
    n902, n903, n904, n905, n906, n907, n908,
    n909, n910, n911, n912, n913, n914, n915,
    n916, n917, n918, n919, n920, n921, n922,
    n923, n924, n925, n926, n927, n928, n929,
    n930, n931, n932, n933, n934, n935, n936,
    n937, n938, n939, n940, n941, n942, n943,
    n944, n945, n946, n947, n948, n949, n950,
    n951, n952, n953, n954, n955, n956, n957,
    n958, n959, n960, n961, n962, n963, n964,
    n965, n966, n967, n968, n969, n970, n971,
    n972, n973, n974, n975, n976, n977, n978,
    n979, n980, n981, n982, n983, n984, n985,
    n986, n987, n988, n989, n990, n991, n992,
    n993, n994, n995, n996, n997, n998, n999,
    n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011,
    n1012, n1013, n1014, n1015, n1016, n1017,
    n1018, n1019, n1020, n1021, n1022, n1023,
    n1024, n1025, n1026, n1027, n1028, n1029,
    n1030, n1031, n1032, n1033, n1034, n1035,
    n1036, n1037, n1038, n1039, n1040, n1041,
    n1042, n1043, n1044, n1045, n1046, n1047,
    n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059,
    n1060, n1061, n1062, n1063, n1064, n1065,
    n1066, n1067, n1068, n1069, n1070, n1071,
    n1072, n1073, n1074, n1075, n1076, n1077,
    n1078, n1079, n1080, n1081, n1082, n1083,
    n1084, n1085, n1086, n1087, n1088, n1089,
    n1090, n1091, n1092, n1093, n1094, n1095,
    n1096, n1097, n1098, n1099, n1100, n1101,
    n1102, n1103, n1104, n1105, n1106, n1107,
    n1108, n1109, n1110, n1111, n1112, n1113,
    n1114, n1115, n1116, n1117, n1118, n1119,
    n1120, n1121, n1122, n1123, n1124, n1125,
    n1126, n1127, n1128, n1129, n1130, n1131,
    n1132, n1133, n1134, n1135, n1136, n1137,
    n1138, n1139, n1140, n1141, n1142, n1143,
    n1144, n1145, n1146, n1147, n1148, n1149,
    n1150, n1151, n1152, n1153, n1154, n1155,
    n1156, n1157, n1158, n1159, n1160, n1161,
    n1162, n1163, n1164, n1165, n1166, n1167,
    n1168, n1169, n1170, n1171, n1172, n1173,
    n1174, n1175, n1176, n1177, n1178, n1179,
    n1180, n1181, n1182, n1183, n1184, n1185,
    n1186, n1187, n1188, n1189, n1190, n1191,
    n1192, n1193, n1194, n1195, n1196, n1197,
    n1198, n1199, n1200, n1201, n1202, n1203,
    n1204, n1205, n1206, n1207, n1208, n1209,
    n1210, n1211, n1212, n1213, n1214, n1215,
    n1216, n1217, n1218, n1219, n1220, n1221,
    n1222, n1223, n1224, n1225, n1226, n1227,
    n1228, n1229, n1230, n1231, n1232, n1233,
    n1234, n1235, n1236, n1237, n1238, n1239,
    n1240, n1241, n1242, n1243, n1244, n1245,
    n1246, n1247, n1248, n1249, n1250, n1251,
    n1252, n1253, n1254, n1255, n1256, n1257,
    n1258, n1259, n1260, n1261, n1262, n1263,
    n1264, n1265, n1266, n1267, n1268, n1269,
    n1270, n1271, n1272, n1273, n1274, n1275,
    n1276, n1277, n1278, n1279, n1280, n1281,
    n1282, n1283, n1284, n1285, n1286, n1287,
    n1288, n1289, n1290, n1291, n1292, n1293,
    n1294, n1295, n1296, n1297, n1298, n1299,
    n1300, n1301, n1302, n1303, n1304, n1305,
    n1306, n1307, n1308, n1309, n1310, n1311,
    n1312, n1313, n1314, n1315, n1316, n1317,
    n1318, n1319, n1320, n1321, n1322, n1323,
    n1324, n1325, n1326, n1327, n1328, n1329,
    n1330, n1331, n1332, n1333, n1334, n1335,
    n1336, n1337, n1338, n1339, n1340, n1341,
    n1342, n1343, n1344, n1345, n1346, n1347,
    n1348, n1349, n1350, n1351, n1352, n1353,
    n1354, n1355, n1356, n1357, n1358, n1359,
    n1360, n1361, n1362, n1363, n1364, n1365,
    n1366, n1367, n1368, n1369, n1370, n1371,
    n1372, n1373, n1374, n1375, n1376, n1377,
    n1378, n1379, n1380, n1381, n1382, n1383,
    n1384, n1385, n1386, n1387, n1388, n1389,
    n1390, n1391, n1392, n1393, n1394, n1395,
    n1396, n1397, n1398, n1399, n1400, n1401,
    n1402, n1403, n1404, n1405, n1406, n1407,
    n1408, n1409, n1410, n1411, n1412, n1413,
    n1414, n1415, n1416, n1417, n1418, n1419,
    n1420, n1421, n1422, n1423, n1424, n1425,
    n1426, n1427, n1428, n1429, n1430, n1431,
    n1432, n1433, n1434, n1435, n1436, n1437,
    n1438, n1439, n1440, n1441, n1442, n1443,
    n1444, n1445, n1446, n1447, n1448, n1449,
    n1450, n1451, n1452, n1453, n1454, n1455,
    n1456, n1457, n1458, n1459, n1460, n1461,
    n1462, n1463, n1464, n1465, n1466, n1467,
    n1468, n1469, n1470, n1471, n1472, n1473,
    n1474, n1475, n1476, n1477, n1478, n1479,
    n1480, n1481, n1482, n1483, n1484, n1485,
    n1486, n1487, n1488, n1489, n1490, n1491,
    n1492, n1493, n1494, n1495, n1496, n1497,
    n1498, n1499, n1500, n1501, n1502, n1503,
    n1504, n1505, n1506, n1507, n1508, n1509,
    n1510, n1511, n1512, n1513, n1514, n1515,
    n1516, n1517, n1518, n1519, n1520, n1521,
    n1522, n1523, n1524, n1525, n1526, n1527,
    n1528, n1529, n1530, n1531, n1532, n1533,
    n1534, n1535, n1536, n1537, n1538, n1539,
    n1540, n1541, n1542, n1543, n1544, n1545,
    n1546, n1547, n1548, n1549, n1550, n1551,
    n1552, n1553, n1554, n1555, n1556, n1557,
    n1558, n1559, n1560, n1561, n1562, n1563,
    n1564, n1565, n1566, n1567, n1568, n1569,
    n1570, n1571, n1572, n1573, n1574, n1575,
    n1576, n1577, n1578, n1579, n1580, n1581,
    n1582, n1583, n1584, n1585, n1586, n1587,
    n1588, n1589, n1590, n1591, n1592, n1593,
    n1594, n1595, n1596, n1597, n1598, n1599,
    n1600, n1601, n1602, n1603, n1604, n1605,
    n1606, n1607, n1608, n1609, n1610, n1611,
    n1612, n1613, n1614, n1615, n1616, n1617,
    n1618, n1619, n1620, n1621, n1622, n1623,
    n1624, n1625, n1626, n1627, n1628, n1629,
    n1630, n1631, n1632, n1633, n1634, n1635,
    n1636, n1637, n1638, n1639, n1640, n1641,
    n1642, n1643, n1644, n1645, n1646, n1647,
    n1648, n1649, n1650, n1651, n1652, n1653,
    n1654, n1655, n1656, n1657, n1658, n1659,
    n1660, n1661, n1662, n1663, n1664, n1665,
    n1666, n1667, n1668, n1669, n1670, n1671,
    n1672, n1673, n1674, n1675, n1676, n1677,
    n1678, n1679, n1680, n1681, n1682, n1683,
    n1684, n1685, n1686, n1687, n1688, n1689,
    n1690, n1691, n1692, n1693, n1694, n1695,
    n1696, n1697, n1698, n1699, n1700, n1701,
    n1702, n1703, n1704, n1705, n1706, n1707,
    n1708, n1709, n1710, n1711, n1712, n1713,
    n1714, n1715, n1716, n1717, n1718, n1719,
    n1720, n1721, n1722, n1723, n1724, n1725,
    n1726, n1727, n1728, n1729, n1730, n1731,
    n1732, n1733, n1734, n1735, n1736, n1737,
    n1738, n1739, n1740, n1741, n1742, n1743,
    n1744, n1745, n1746, n1747, n1748, n1749,
    n1750, n1751, n1752, n1753, n1754, n1755,
    n1756, n1757, n1758, n1759, n1760, n1761,
    n1762, n1763, n1764, n1765, n1766, n1767,
    n1768, n1769, n1770, n1771, n1772, n1773,
    n1774, n1775, n1776, n1777, n1778, n1779,
    n1780, n1781, n1782, n1783, n1784, n1785,
    n1786, n1787, n1788, n1789, n1790, n1791,
    n1792, n1793, n1794, n1795, n1796, n1797,
    n1798, n1799, n1800, n1801, n1802, n1803,
    n1804, n1805, n1806, n1807, n1808, n1809,
    n1810, n1811, n1812, n1813, n1814, n1815,
    n1816, n1817, n1818, n1819, n1820, n1821,
    n1822, n1823, n1824, n1825, n1826, n1827,
    n1828, n1829, n1830, n1831, n1832, n1833,
    n1834, n1835, n1836, n1837, n1838, n1839,
    n1840, n1841, n1842, n1843, n1844, n1845,
    n1846, n1847, n1848, n1849, n1850, n1851,
    n1852, n1853, n1854, n1855, n1856, n1857,
    n1858, n1859, n1860, n1861, n1862, n1863,
    n1864, n1865, n1866, n1867, n1868, n1869,
    n1870, n1871, n1872, n1873, n1874, n1875,
    n1876, n1877, n1878, n1879, n1880, n1881,
    n1882, n1883, n1884, n1885, n1886, n1887,
    n1888, n1889, n1890, n1891, n1892, n1893,
    n1894, n1895, n1896, n1897, n1898, n1899,
    n1900, n1901, n1902, n1903, n1904, n1905,
    n1906, n1907, n1908, n1909, n1910, n1911,
    n1912, n1913, n1914, n1915, n1916, n1917,
    n1918, n1919, n1920, n1921, n1922, n1923,
    n1924, n1925, n1926, n1927, n1928, n1929,
    n1930, n1931, n1932, n1933, n1934, n1935,
    n1936, n1937, n1938, n1939, n1940, n1941,
    n1942, n1943, n1944, n1945, n1946, n1947,
    n1948, n1949, n1950, n1951, n1952, n1953,
    n1954, n1955, n1956, n1957, n1958, n1959,
    n1960, n1961, n1962, n1963, n1964, n1965,
    n1966, n1967, n1968, n1969, n1970, n1971,
    n1972, n1973, n1974, n1975, n1976, n1977,
    n1978, n1979, n1980, n1981, n1982, n1983,
    n1984, n1985, n1986, n1987, n1988, n1989,
    n1990, n1991, n1992, n1993, n1994, n1995,
    n1996, n1997, n1998, n1999, n2000, n2001,
    n2002, n2003, n2004, n2005, n2006, n2007,
    n2008, n2009, n2010, n2011, n2012, n2013,
    n2014, n2015, n2016, n2017, n2018, n2019,
    n2020, n2021, n2022, n2023, n2024, n2025,
    n2026, n2027, n2028, n2029, n2030, n2031,
    n2032, n2033, n2034, n2035, n2036, n2037,
    n2038, n2039, n2040, n2041, n2042, n2043,
    n2044, n2045, n2046, n2047, n2048, n2049,
    n2050, n2051, n2052, n2053, n2054, n2055,
    n2056, n2057, n2058, n2059, n2060, n2061,
    n2062, n2063, n2064, n2065, n2066, n2067,
    n2068, n2069, n2070, n2071, n2072, n2073,
    n2074, n2075, n2076, n2077, n2078, n2079,
    n2080, n2081, n2082, n2083, n2084, n2085,
    n2086, n2087, n2088, n2089, n2090, n2091,
    n2092, n2093, n2094, n2095, n2096, n2097,
    n2098, n2099, n2100, n2101, n2102, n2103,
    n2104, n2105, n2106, n2107, n2108, n2109,
    n2110, n2111, n2112, n2113, n2114, n2115,
    n2116, n2117, n2118, n2119, n2120, n2121,
    n2122, n2123, n2124, n2125, n2126, n2127,
    n2128, n2129, n2130, n2131, n2132, n2133,
    n2134, n2135, n2136, n2137, n2138, n2139,
    n2140, n2141, n2142, n2143, n2144, n2145,
    n2146, n2147, n2148, n2149, n2150, n2151,
    n2152, n2153, n2154, n2155, n2156, n2157,
    n2158, n2159, n2160, n2161, n2162, n2163,
    n2164, n2165, n2166, n2167, n2168, n2169,
    n2170, n2171, n2172, n2173, n2174, n2175,
    n2176, n2177, n2178, n2179, n2180, n2181,
    n2182, n2183, n2184, n2185, n2186, n2187,
    n2188, n2189, n2190, n2191, n2192, n2193,
    n2194, n2195, n2196, n2197, n2198, n2199,
    n2200, n2201, n2202, n2203, n2204, n2205,
    n2206, n2207, n2208, n2209, n2210, n2211,
    n2212, n2213, n2214, n2215, n2216, n2217,
    n2218, n2219, n2220, n2221, n2222, n2223,
    n2224, n2225, n2226, n2227, n2228, n2229,
    n2230, n2231, n2232, n2233, n2234, n2235,
    n2236, n2237, n2238, n2239, n2240, n2241,
    n2242, n2243, n2244, n2245, n2246, n2247,
    n2248, n2249, n2250, n2251, n2252, n2253,
    n2254, n2255, n2256, n2257, n2258, n2259,
    n2260, n2261, n2262, n2263, n2264, n2265,
    n2266, n2267, n2268, n2269, n2270, n2271,
    n2272, n2273, n2274, n2275, n2276, n2277,
    n2278, n2279, n2280, n2281, n2282, n2283,
    n2284, n2285, n2286, n2287, n2288, n2289,
    n2290, n2291, n2292, n2293, n2294, n2295,
    n2296, n2297, n2298, n2299, n2300, n2301,
    n2302, n2303, n2304, n2305, n2306, n2307,
    n2308, n2309, n2310, n2311, n2312, n2313,
    n2314, n2315, n2316, n2317, n2318, n2319,
    n2320, n2321, n2322, n2323, n2324, n2325,
    n2326, n2327, n2328, n2329, n2330, n2331,
    n2332, n2333, n2334, n2335, n2336, n2337,
    n2338, n2339, n2340, n2341, n2342, n2343,
    n2344, n2345, n2346, n2347, n2348, n2349,
    n2350, n2351, n2352, n2353, n2354, n2355,
    n2356, n2357, n2358, n2359, n2360, n2361,
    n2362, n2363, n2364, n2365, n2366, n2367,
    n2368, n2369, n2370, n2371, n2372, n2373,
    n2374, n2375, n2376, n2377, n2378, n2379,
    n2380, n2381, n2382, n2383, n2384, n2385,
    n2386, n2387, n2388, n2389, n2390, n2391,
    n2392, n2393, n2394, n2395, n2396, n2397,
    n2398, n2399, n2400, n2401, n2402, n2403,
    n2404, n2405, n2406, n2407, n2408, n2409,
    n2410, n2411, n2412, n2413, n2414, n2415,
    n2416, n2417, n2418, n2419, n2420, n2421,
    n2422, n2423, n2424, n2425, n2426, n2427,
    n2428, n2429, n2430, n2431, n2432, n2433,
    n2434, n2435, n2436, n2437, n2438, n2439,
    n2440, n2441, n2442, n2443, n2444, n2445,
    n2446, n2447, n2448, n2449, n2450, n2451,
    n2452, n2453, n2454, n2455, n2456, n2457,
    n2458, n2459, n2460, n2461, n2462, n2463,
    n2464, n2465, n2466, n2467, n2468, n2469,
    n2470, n2471, n2472, n2473, n2474, n2475,
    n2476, n2477, n2478, n2479, n2480, n2481,
    n2482, n2483, n2484, n2485, n2486, n2487,
    n2488, n2489, n2490, n2491, n2492, n2493,
    n2494, n2495, n2496, n2497, n2498, n2499,
    n2500, n2501, n2502, n2503, n2504, n2505,
    n2506, n2507, n2508, n2509, n2510, n2511,
    n2512, n2513, n2514, n2515, n2516, n2517,
    n2518, n2519, n2520, n2521, n2522, n2523,
    n2524, n2525, n2526, n2527, n2528, n2529,
    n2530, n2531, n2532, n2533, n2534, n2535,
    n2536, n2537, n2538, n2539, n2540, n2541,
    n2542, n2543, n2544, n2545, n2546, n2547,
    n2548, n2549, n2550, n2551, n2552, n2553,
    n2554, n2555, n2556, n2557, n2558, n2559,
    n2560, n2561, n2562, n2563, n2564, n2565,
    n2566, n2567, n2568, n2569, n2570, n2571,
    n2572, n2573, n2574, n2575, n2576, n2577,
    n2578, n2579, n2580, n2581, n2582, n2583,
    n2584, n2585, n2586, n2587, n2588, n2589,
    n2590, n2591, n2592, n2593, n2594, n2595,
    n2596, n2597, n2598, n2599, n2600, n2601,
    n2602, n2603, n2604, n2605, n2606, n2607,
    n2608, n2609, n2610, n2611, n2612, n2613,
    n2614, n2615, n2616, n2617, n2618, n2619,
    n2620, n2621, n2622, n2623, n2624, n2625,
    n2626, n2627, n2628, n2629, n2630, n2631,
    n2632, n2633, n2634, n2635, n2636, n2637,
    n2638, n2639, n2640, n2641, n2642, n2643,
    n2644, n2645, n2646, n2647, n2648, n2649,
    n2650, n2651, n2652, n2653, n2654, n2655,
    n2656, n2657, n2658, n2659, n2660, n2661,
    n2662, n2663, n2664, n2665, n2666, n2667,
    n2668, n2669, n2670, n2671, n2672, n2673,
    n2674, n2675, n2676, n2677, n2678, n2679,
    n2680, n2681, n2682, n2683, n2684, n2685,
    n2686, n2687, n2688, n2689, n2690, n2691,
    n2692, n2693, n2694, n2695, n2696, n2697,
    n2698, n2699, n2700, n2701, n2702, n2703,
    n2704, n2705, n2706, n2707, n2708, n2709,
    n2710, n2711, n2712, n2713, n2714, n2715,
    n2716, n2717, n2718, n2719, n2720, n2721,
    n2722, n2723, n2724, n2725, n2726, n2727,
    n2728, n2729, n2730, n2731, n2732, n2733,
    n2734, n2735, n2736, n2737, n2738, n2739,
    n2740, n2741, n2742, n2743, n2744, n2745,
    n2746, n2747, n2748, n2749, n2750, n2751,
    n2752, n2753, n2754, n2755, n2756, n2757,
    n2758, n2759, n2760, n2761, n2762, n2763,
    n2764, n2765, n2766, n2767, n2768, n2769,
    n2770, n2771, n2772, n2773, n2774, n2775,
    n2776, n2777, n2778, n2779, n2780, n2781,
    n2782, n2783, n2784, n2785, n2786, n2787,
    n2788, n2789, n2790, n2791, n2792, n2793,
    n2794, n2795, n2796, n2797, n2798, n2799,
    n2800, n2801, n2802, n2803, n2804, n2805,
    n2806, n2807, n2808, n2809, n2810, n2811,
    n2812, n2813, n2814, n2815, n2816, n2817,
    n2818, n2819, n2820, n2821, n2822, n2823,
    n2824, n2825, n2826, n2827, n2828, n2829,
    n2830, n2831, n2832, n2833, n2834, n2835,
    n2836, n2837, n2838, n2839, n2840, n2841,
    n2842, n2843, n2844, n2845, n2846, n2847,
    n2848, n2849, n2850, n2851, n2852, n2853,
    n2854, n2855, n2856, n2857, n2858, n2859,
    n2860, n2861, n2862, n2863, n2864, n2865,
    n2866, n2867, n2868, n2869, n2870, n2871,
    n2872, n2873, n2874, n2875, n2876, n2877,
    n2878, n2879, n2880, n2881, n2882, n2883,
    n2884, n2885, n2886, n2887, n2888, n2889,
    n2890, n2891, n2892, n2893, n2894, n2895,
    n2896, n2897, n2898, n2899, n2900, n2901,
    n2902, n2903, n2904, n2905, n2906, n2907,
    n2908, n2909, n2910, n2911, n2912, n2913,
    n2914, n2915, n2916, n2917, n2918, n2919,
    n2920, n2921, n2922, n2923, n2924, n2925,
    n2926, n2927, n2928, n2929, n2930, n2931,
    n2932, n2933, n2934, n2935, n2936, n2937,
    n2938, n2939, n2940, n2941, n2942, n2943,
    n2944, n2945, n2946, n2947, n2948, n2949,
    n2950, n2951, n2952, n2953, n2954, n2955,
    n2956, n2957, n2958, n2959, n2960, n2961,
    n2962, n2963, n2964, n2965, n2966, n2967,
    n2968, n2969, n2970, n2971, n2972, n2973,
    n2974, n2975, n2976, n2977, n2978, n2979,
    n2980, n2981, n2982, n2983, n2984, n2985,
    n2986, n2987, n2988, n2989, n2990, n2991,
    n2992, n2993, n2994, n2995, n2996, n2997,
    n2998, n2999, n3000, n3001, n3002, n3003,
    n3004, n3005, n3006, n3007, n3008, n3009,
    n3010, n3011, n3012, n3013, n3014, n3015,
    n3016, n3017, n3018, n3019, n3020, n3021,
    n3022, n3023, n3024, n3025, n3026, n3027,
    n3028, n3029, n3030, n3031, n3032, n3033,
    n3034, n3035, n3036, n3037, n3038, n3039,
    n3040, n3041, n3042, n3043, n3044, n3045,
    n3046, n3047, n3048, n3049, n3050, n3051,
    n3052, n3053, n3054, n3055, n3056, n3057,
    n3058, n3059, n3060, n3061, n3062, n3063,
    n3064, n3065, n3066, n3067, n3068, n3069,
    n3070, n3071, n3072, n3073, n3074, n3075,
    n3076, n3077, n3078, n3079, n3080, n3081,
    n3082, n3083, n3084, n3085, n3086, n3087,
    n3088, n3089, n3090, n3091, n3092, n3093,
    n3094, n3095, n3096, n3097, n3098, n3099,
    n3100, n3101, n3102, n3103, n3104, n3105,
    n3106, n3107, n3108, n3109, n3110, n3111,
    n3112, n3113, n3114, n3115, n3117, n3118,
    n3120, n3121, n3123, n3124, n3126, n3127,
    n3129, n3130, n3132, n3133, n3135, n3136,
    n3138, n3139, n3141, n3142, n3144, n3145,
    n3147, n3148, n3150, n3151, n3153, n3154,
    n3156, n3157, n3159, n3160, n3162, n3163,
    n3165, n3166, n3168, n3169, n3171, n3172,
    n3174, n3175, n3177, n3178, n3180, n3181,
    n3183, n3184, n3186, n3187, n3189, n3190,
    n3192, n3193, n3195, n3196, n3198, n3199,
    n3201, n3202, n3204, n3205, n3207, n3208,
    n3210, n3211, n3213, n3214, n3216, n3217,
    n3219, n3220, n3222, n3223, n3225, n3226,
    n3228, n3229, n3231, n3232, n3234, n3235,
    n3237, n3238, n3240, n3241, n3243, n3244,
    n3246, n3247, n3249, n3250, n3252, n3253,
    n3255, n3256, n3258, n3259, n3261, n3262,
    n3264, n3265, n3267, n3268, n3270, n3271,
    n3273, n3274, n3276, n3277, n3279, n3280,
    n3282, n3283, n3285, n3286, n3288, n3289,
    n3291, n3292, n3294, n3295, n3297, n3298,
    n3300, n3301, n3303, n3304, n3306, n3307,
    n3309, n3310, n3312, n3313, n3315, n3316,
    n3318, n3319, n3321, n3322, n3324, n3325,
    n3327, n3328, n3330, n3331, n3333, n3334,
    n3336, n3337, n3339, n3340, n3342, n3343,
    n3345, n3346, n3348, n3349, n3351, n3352,
    n3354, n3355, n3357, n3358, n3360, n3361,
    n3363, n3364, n3366, n3367, n3369, n3370,
    n3372, n3373, n3375, n3376, n3378, n3379,
    n3381, n3382, n3384, n3385, n3387, n3388,
    n3390, n3391, n3393, n3394, n3396, n3397,
    n3399, n3400, n3402, n3403, n3405, n3406,
    n3408, n3409, n3411, n3412, n3414, n3415,
    n3417, n3418, n3420, n3421, n3423, n3424,
    n3426, n3427, n3429, n3430, n3432, n3433,
    n3435, n3436, n3438, n3439, n3441, n3442,
    n3444, n3445, n3447, n3448, n3450, n3451,
    n3453, n3454, n3456, n3457, n3459, n3460,
    n3462, n3463, n3465, n3466, n3468, n3469,
    n3471, n3472, n3474, n3475, n3477, n3478,
    n3480, n3481, n3483, n3484, n3486, n3487,
    n3489, n3490, n3492, n3493, n3495, n3496,
    n3499, n3500;
  assign n643 = ~pi383  & pi511 ;
  assign n644 = ~pi382  & pi510 ;
  assign n645 = ~pi381  & pi509 ;
  assign n646 = ~n644 & ~n645;
  assign n647 = pi380  & ~pi508 ;
  assign n648 = pi381  & ~pi509 ;
  assign n649 = ~n647 & ~n648;
  assign n650 = n646 & ~n649;
  assign n651 = pi382  & ~pi510 ;
  assign n652 = ~n650 & ~n651;
  assign n653 = ~pi377  & pi505 ;
  assign n654 = ~pi379  & pi507 ;
  assign n655 = ~pi378  & pi506 ;
  assign n656 = ~n654 & ~n655;
  assign n657 = ~pi375  & pi503 ;
  assign n658 = ~pi502  & ~n657;
  assign n659 = pi374  & ~n657;
  assign n660 = ~n658 & ~n659;
  assign n661 = ~pi369  & pi497 ;
  assign n662 = ~pi371  & pi499 ;
  assign n663 = ~pi370  & pi498 ;
  assign n664 = ~n662 & ~n663;
  assign n665 = ~pi367  & pi495 ;
  assign n666 = ~pi494  & ~n665;
  assign n667 = pi366  & ~n665;
  assign n668 = ~n666 & ~n667;
  assign n669 = ~pi361  & pi489 ;
  assign n670 = ~pi363  & pi491 ;
  assign n671 = ~pi362  & pi490 ;
  assign n672 = ~n670 & ~n671;
  assign n673 = ~pi359  & pi487 ;
  assign n674 = ~pi486  & ~n673;
  assign n675 = pi358  & ~n673;
  assign n676 = ~n674 & ~n675;
  assign n677 = ~pi353  & pi481 ;
  assign n678 = ~pi355  & pi483 ;
  assign n679 = ~pi354  & pi482 ;
  assign n680 = ~n678 & ~n679;
  assign n681 = ~pi351  & pi479 ;
  assign n682 = ~pi478  & ~n681;
  assign n683 = pi350  & ~n681;
  assign n684 = ~n682 & ~n683;
  assign n685 = ~pi345  & pi473 ;
  assign n686 = ~pi347  & pi475 ;
  assign n687 = ~pi346  & pi474 ;
  assign n688 = ~n686 & ~n687;
  assign n689 = ~pi343  & pi471 ;
  assign n690 = ~pi470  & ~n689;
  assign n691 = pi342  & ~n689;
  assign n692 = ~n690 & ~n691;
  assign n693 = ~pi337  & pi465 ;
  assign n694 = ~pi339  & pi467 ;
  assign n695 = ~pi338  & pi466 ;
  assign n696 = ~n694 & ~n695;
  assign n697 = ~pi335  & pi463 ;
  assign n698 = ~pi462  & ~n697;
  assign n699 = pi334  & ~n697;
  assign n700 = ~n698 & ~n699;
  assign n701 = ~pi329  & pi457 ;
  assign n702 = ~pi331  & pi459 ;
  assign n703 = ~pi330  & pi458 ;
  assign n704 = ~n702 & ~n703;
  assign n705 = ~pi327  & pi455 ;
  assign n706 = ~pi454  & ~n705;
  assign n707 = pi326  & ~n705;
  assign n708 = ~n706 & ~n707;
  assign n709 = ~pi321  & pi449 ;
  assign n710 = ~pi323  & pi451 ;
  assign n711 = ~pi322  & pi450 ;
  assign n712 = ~n710 & ~n711;
  assign n713 = pi315  & ~pi443 ;
  assign n714 = ~pi315  & pi443 ;
  assign n715 = ~pi314  & pi442 ;
  assign n716 = ~n714 & ~n715;
  assign n717 = pi314  & ~pi442 ;
  assign n718 = pi313  & ~pi441 ;
  assign n719 = ~pi313  & pi441 ;
  assign n720 = ~pi440  & ~n719;
  assign n721 = pi312  & n720;
  assign n722 = ~n718 & ~n721;
  assign n723 = ~n717 & n722;
  assign n724 = n716 & ~n723;
  assign n725 = ~n713 & ~n724;
  assign n726 = ~pi319  & pi447 ;
  assign n727 = ~pi446  & ~n726;
  assign n728 = pi318  & ~n726;
  assign n729 = ~n727 & ~n728;
  assign n730 = ~pi317  & pi445 ;
  assign n731 = ~pi316  & pi444 ;
  assign n732 = ~n730 & ~n731;
  assign n733 = ~n729 & n732;
  assign n734 = ~n725 & n733;
  assign n735 = ~pi446  & n728;
  assign n736 = pi319  & ~pi447 ;
  assign n737 = pi317  & ~pi445 ;
  assign n738 = ~pi444  & ~n730;
  assign n739 = pi316  & n738;
  assign n740 = ~n737 & ~n739;
  assign n741 = ~n729 & ~n740;
  assign n742 = ~pi312  & pi440 ;
  assign n743 = n733 & ~n742;
  assign n744 = pi311  & ~pi439 ;
  assign n745 = ~pi311  & pi439 ;
  assign n746 = ~pi310  & pi438 ;
  assign n747 = ~n745 & ~n746;
  assign n748 = pi310  & ~pi438 ;
  assign n749 = pi309  & ~pi437 ;
  assign n750 = ~pi309  & pi437 ;
  assign n751 = ~pi436  & ~n750;
  assign n752 = pi308  & n751;
  assign n753 = ~n749 & ~n752;
  assign n754 = ~n748 & n753;
  assign n755 = n747 & ~n754;
  assign n756 = pi307  & ~pi435 ;
  assign n757 = ~pi307  & pi435 ;
  assign n758 = ~pi306  & pi434 ;
  assign n759 = ~n757 & ~n758;
  assign n760 = pi306  & ~pi434 ;
  assign n761 = pi305  & ~pi433 ;
  assign n762 = ~pi305  & pi433 ;
  assign n763 = ~pi432  & ~n762;
  assign n764 = pi304  & n763;
  assign n765 = ~n761 & ~n764;
  assign n766 = ~n760 & n765;
  assign n767 = n759 & ~n766;
  assign n768 = ~n756 & ~n767;
  assign n769 = ~pi308  & pi436 ;
  assign n770 = n747 & ~n769;
  assign n771 = ~n750 & n770;
  assign n772 = ~n768 & n771;
  assign n773 = ~n755 & ~n772;
  assign n774 = ~pi304  & pi432 ;
  assign n775 = n759 & ~n774;
  assign n776 = pi299  & ~pi427 ;
  assign n777 = ~pi299  & pi427 ;
  assign n778 = ~pi298  & pi426 ;
  assign n779 = ~n777 & ~n778;
  assign n780 = pi298  & ~pi426 ;
  assign n781 = pi297  & ~pi425 ;
  assign n782 = ~pi297  & pi425 ;
  assign n783 = ~pi424  & ~n782;
  assign n784 = pi296  & n783;
  assign n785 = ~n781 & ~n784;
  assign n786 = ~n780 & n785;
  assign n787 = n779 & ~n786;
  assign n788 = ~n776 & ~n787;
  assign n789 = ~pi303  & pi431 ;
  assign n790 = ~pi430  & ~n789;
  assign n791 = pi302  & ~n789;
  assign n792 = ~n790 & ~n791;
  assign n793 = ~pi301  & pi429 ;
  assign n794 = ~pi300  & pi428 ;
  assign n795 = ~n793 & ~n794;
  assign n796 = ~n792 & n795;
  assign n797 = ~n788 & n796;
  assign n798 = ~pi430  & n791;
  assign n799 = pi303  & ~pi431 ;
  assign n800 = pi301  & ~pi429 ;
  assign n801 = ~pi428  & ~n793;
  assign n802 = pi300  & n801;
  assign n803 = ~n800 & ~n802;
  assign n804 = ~n792 & ~n803;
  assign n805 = ~pi296  & pi424 ;
  assign n806 = n796 & ~n805;
  assign n807 = ~pi295  & pi423 ;
  assign n808 = ~pi422  & ~n807;
  assign n809 = pi294  & ~n807;
  assign n810 = ~n808 & ~n809;
  assign n811 = ~pi293  & pi421 ;
  assign n812 = ~pi292  & pi420 ;
  assign n813 = ~n811 & ~n812;
  assign n814 = ~n810 & n813;
  assign n815 = pi287  & ~pi415 ;
  assign n816 = pi286  & ~pi414 ;
  assign n817 = ~pi286  & pi414 ;
  assign n818 = pi285  & ~pi413 ;
  assign n819 = ~pi285  & pi413 ;
  assign n820 = pi284  & ~pi412 ;
  assign n821 = ~pi284  & pi412 ;
  assign n822 = pi283  & ~pi411 ;
  assign n823 = ~pi283  & pi411 ;
  assign n824 = pi282  & ~pi410 ;
  assign n825 = ~pi282  & pi410 ;
  assign n826 = pi281  & ~pi409 ;
  assign n827 = ~pi281  & pi409 ;
  assign n828 = pi280  & ~pi408 ;
  assign n829 = ~pi280  & pi408 ;
  assign n830 = pi279  & ~pi407 ;
  assign n831 = ~pi279  & pi407 ;
  assign n832 = pi278  & ~pi406 ;
  assign n833 = ~pi278  & pi406 ;
  assign n834 = pi277  & ~pi405 ;
  assign n835 = ~pi277  & pi405 ;
  assign n836 = pi276  & ~pi404 ;
  assign n837 = ~pi276  & pi404 ;
  assign n838 = pi275  & ~pi403 ;
  assign n839 = ~pi275  & pi403 ;
  assign n840 = pi274  & ~pi402 ;
  assign n841 = ~pi274  & pi402 ;
  assign n842 = pi273  & ~pi401 ;
  assign n843 = ~pi273  & pi401 ;
  assign n844 = pi272  & ~pi400 ;
  assign n845 = ~pi272  & pi400 ;
  assign n846 = pi271  & ~pi399 ;
  assign n847 = ~pi271  & pi399 ;
  assign n848 = pi270  & ~pi398 ;
  assign n849 = ~pi270  & pi398 ;
  assign n850 = pi269  & ~pi397 ;
  assign n851 = ~pi269  & pi397 ;
  assign n852 = pi268  & ~pi396 ;
  assign n853 = ~pi268  & pi396 ;
  assign n854 = pi267  & ~pi395 ;
  assign n855 = ~pi267  & pi395 ;
  assign n856 = pi266  & ~pi394 ;
  assign n857 = ~pi266  & pi394 ;
  assign n858 = pi265  & ~pi393 ;
  assign n859 = ~pi265  & pi393 ;
  assign n860 = pi264  & ~pi392 ;
  assign n861 = ~pi264  & pi392 ;
  assign n862 = pi263  & ~pi391 ;
  assign n863 = ~pi263  & pi391 ;
  assign n864 = pi262  & ~pi390 ;
  assign n865 = ~pi262  & pi390 ;
  assign n866 = pi261  & ~pi389 ;
  assign n867 = ~pi261  & pi389 ;
  assign n868 = pi260  & ~pi388 ;
  assign n869 = ~pi260  & pi388 ;
  assign n870 = pi259  & ~pi387 ;
  assign n871 = ~pi259  & pi387 ;
  assign n872 = pi258  & ~pi386 ;
  assign n873 = ~pi258  & pi386 ;
  assign n874 = pi257  & ~pi385 ;
  assign n875 = pi256  & ~pi384 ;
  assign n876 = ~pi257  & pi385 ;
  assign n877 = n875 & ~n876;
  assign n878 = ~n874 & ~n877;
  assign n879 = ~n873 & ~n878;
  assign n880 = ~n872 & ~n879;
  assign n881 = ~n871 & ~n880;
  assign n882 = ~n870 & ~n881;
  assign n883 = ~n869 & ~n882;
  assign n884 = ~n868 & ~n883;
  assign n885 = ~n867 & ~n884;
  assign n886 = ~n866 & ~n885;
  assign n887 = ~n865 & ~n886;
  assign n888 = ~n864 & ~n887;
  assign n889 = ~n863 & ~n888;
  assign n890 = ~n862 & ~n889;
  assign n891 = ~n861 & ~n890;
  assign n892 = ~n860 & ~n891;
  assign n893 = ~n859 & ~n892;
  assign n894 = ~n858 & ~n893;
  assign n895 = ~n857 & ~n894;
  assign n896 = ~n856 & ~n895;
  assign n897 = ~n855 & ~n896;
  assign n898 = ~n854 & ~n897;
  assign n899 = ~n853 & ~n898;
  assign n900 = ~n852 & ~n899;
  assign n901 = ~n851 & ~n900;
  assign n902 = ~n850 & ~n901;
  assign n903 = ~n849 & ~n902;
  assign n904 = ~n848 & ~n903;
  assign n905 = ~n847 & ~n904;
  assign n906 = ~n846 & ~n905;
  assign n907 = ~n845 & ~n906;
  assign n908 = ~n844 & ~n907;
  assign n909 = ~n843 & ~n908;
  assign n910 = ~n842 & ~n909;
  assign n911 = ~n841 & ~n910;
  assign n912 = ~n840 & ~n911;
  assign n913 = ~n839 & ~n912;
  assign n914 = ~n838 & ~n913;
  assign n915 = ~n837 & ~n914;
  assign n916 = ~n836 & ~n915;
  assign n917 = ~n835 & ~n916;
  assign n918 = ~n834 & ~n917;
  assign n919 = ~n833 & ~n918;
  assign n920 = ~n832 & ~n919;
  assign n921 = ~n831 & ~n920;
  assign n922 = ~n830 & ~n921;
  assign n923 = ~n829 & ~n922;
  assign n924 = ~n828 & ~n923;
  assign n925 = ~n827 & ~n924;
  assign n926 = ~n826 & ~n925;
  assign n927 = ~n825 & ~n926;
  assign n928 = ~n824 & ~n927;
  assign n929 = ~n823 & ~n928;
  assign n930 = ~n822 & ~n929;
  assign n931 = ~n821 & ~n930;
  assign n932 = ~n820 & ~n931;
  assign n933 = ~n819 & ~n932;
  assign n934 = ~n818 & ~n933;
  assign n935 = ~n817 & ~n934;
  assign n936 = ~n816 & ~n935;
  assign n937 = ~n815 & n936;
  assign n938 = n814 & ~n937;
  assign n939 = ~pi289  & pi417 ;
  assign n940 = ~pi288  & pi416 ;
  assign n941 = ~pi291  & pi419 ;
  assign n942 = ~pi290  & pi418 ;
  assign n943 = ~n941 & ~n942;
  assign n944 = ~pi287  & pi415 ;
  assign n945 = n943 & ~n944;
  assign n946 = ~n940 & n945;
  assign n947 = ~n939 & n946;
  assign n948 = n938 & n947;
  assign n949 = pi291  & ~pi419 ;
  assign n950 = pi290  & ~pi418 ;
  assign n951 = pi289  & ~pi417 ;
  assign n952 = ~pi416  & ~n939;
  assign n953 = pi288  & n952;
  assign n954 = ~n951 & ~n953;
  assign n955 = ~n950 & n954;
  assign n956 = n943 & ~n955;
  assign n957 = ~n949 & ~n956;
  assign n958 = n814 & ~n957;
  assign n959 = pi295  & ~pi423 ;
  assign n960 = pi293  & ~pi421 ;
  assign n961 = ~pi420  & ~n811;
  assign n962 = pi292  & n961;
  assign n963 = ~n960 & ~n962;
  assign n964 = ~n810 & ~n963;
  assign n965 = ~n959 & ~n964;
  assign n966 = ~n958 & n965;
  assign n967 = ~n948 & n966;
  assign n968 = pi294  & n808;
  assign n969 = n967 & ~n968;
  assign n970 = n779 & ~n969;
  assign n971 = ~n782 & n970;
  assign n972 = n806 & n971;
  assign n973 = ~n804 & ~n972;
  assign n974 = ~n799 & n973;
  assign n975 = ~n798 & n974;
  assign n976 = ~n797 & n975;
  assign n977 = n771 & ~n976;
  assign n978 = ~n762 & n977;
  assign n979 = n775 & n978;
  assign n980 = n773 & ~n979;
  assign n981 = ~n744 & n980;
  assign n982 = n716 & ~n981;
  assign n983 = ~n719 & n982;
  assign n984 = n743 & n983;
  assign n985 = ~n741 & ~n984;
  assign n986 = ~n736 & n985;
  assign n987 = ~n735 & n986;
  assign n988 = ~n734 & n987;
  assign n989 = n712 & ~n988;
  assign n990 = ~n709 & n989;
  assign n991 = ~pi320  & pi448 ;
  assign n992 = n990 & ~n991;
  assign n993 = pi323  & ~pi451 ;
  assign n994 = pi322  & ~pi450 ;
  assign n995 = pi321  & ~pi449 ;
  assign n996 = ~pi448  & ~n709;
  assign n997 = pi320  & n996;
  assign n998 = ~n995 & ~n997;
  assign n999 = ~n994 & n998;
  assign n1000 = n712 & ~n999;
  assign n1001 = ~n993 & ~n1000;
  assign n1002 = ~n992 & n1001;
  assign n1003 = ~n708 & ~n1002;
  assign n1004 = ~pi325  & pi453 ;
  assign n1005 = ~pi324  & pi452 ;
  assign n1006 = ~n1004 & ~n1005;
  assign n1007 = n1003 & n1006;
  assign n1008 = ~pi454  & n707;
  assign n1009 = pi327  & ~pi455 ;
  assign n1010 = pi325  & ~pi453 ;
  assign n1011 = ~pi452  & ~n1004;
  assign n1012 = pi324  & n1011;
  assign n1013 = ~n1010 & ~n1012;
  assign n1014 = ~n708 & ~n1013;
  assign n1015 = ~n1009 & ~n1014;
  assign n1016 = ~n1008 & n1015;
  assign n1017 = ~n1007 & n1016;
  assign n1018 = n704 & ~n1017;
  assign n1019 = ~n701 & n1018;
  assign n1020 = ~pi328  & pi456 ;
  assign n1021 = n1019 & ~n1020;
  assign n1022 = pi331  & ~pi459 ;
  assign n1023 = pi330  & ~pi458 ;
  assign n1024 = pi329  & ~pi457 ;
  assign n1025 = ~pi456  & ~n701;
  assign n1026 = pi328  & n1025;
  assign n1027 = ~n1024 & ~n1026;
  assign n1028 = ~n1023 & n1027;
  assign n1029 = n704 & ~n1028;
  assign n1030 = ~n1022 & ~n1029;
  assign n1031 = ~n1021 & n1030;
  assign n1032 = ~n700 & ~n1031;
  assign n1033 = ~pi333  & pi461 ;
  assign n1034 = ~pi332  & pi460 ;
  assign n1035 = ~n1033 & ~n1034;
  assign n1036 = n1032 & n1035;
  assign n1037 = ~pi462  & n699;
  assign n1038 = pi335  & ~pi463 ;
  assign n1039 = pi333  & ~pi461 ;
  assign n1040 = ~pi460  & ~n1033;
  assign n1041 = pi332  & n1040;
  assign n1042 = ~n1039 & ~n1041;
  assign n1043 = ~n700 & ~n1042;
  assign n1044 = ~n1038 & ~n1043;
  assign n1045 = ~n1037 & n1044;
  assign n1046 = ~n1036 & n1045;
  assign n1047 = n696 & ~n1046;
  assign n1048 = ~n693 & n1047;
  assign n1049 = ~pi336  & pi464 ;
  assign n1050 = n1048 & ~n1049;
  assign n1051 = pi339  & ~pi467 ;
  assign n1052 = pi338  & ~pi466 ;
  assign n1053 = pi337  & ~pi465 ;
  assign n1054 = ~pi464  & ~n693;
  assign n1055 = pi336  & n1054;
  assign n1056 = ~n1053 & ~n1055;
  assign n1057 = ~n1052 & n1056;
  assign n1058 = n696 & ~n1057;
  assign n1059 = ~n1051 & ~n1058;
  assign n1060 = ~n1050 & n1059;
  assign n1061 = ~n692 & ~n1060;
  assign n1062 = ~pi341  & pi469 ;
  assign n1063 = ~pi340  & pi468 ;
  assign n1064 = ~n1062 & ~n1063;
  assign n1065 = n1061 & n1064;
  assign n1066 = ~pi470  & n691;
  assign n1067 = pi343  & ~pi471 ;
  assign n1068 = pi341  & ~pi469 ;
  assign n1069 = ~pi468  & ~n1062;
  assign n1070 = pi340  & n1069;
  assign n1071 = ~n1068 & ~n1070;
  assign n1072 = ~n692 & ~n1071;
  assign n1073 = ~n1067 & ~n1072;
  assign n1074 = ~n1066 & n1073;
  assign n1075 = ~n1065 & n1074;
  assign n1076 = n688 & ~n1075;
  assign n1077 = ~n685 & n1076;
  assign n1078 = ~pi344  & pi472 ;
  assign n1079 = n1077 & ~n1078;
  assign n1080 = pi347  & ~pi475 ;
  assign n1081 = pi346  & ~pi474 ;
  assign n1082 = pi345  & ~pi473 ;
  assign n1083 = ~pi472  & ~n685;
  assign n1084 = pi344  & n1083;
  assign n1085 = ~n1082 & ~n1084;
  assign n1086 = ~n1081 & n1085;
  assign n1087 = n688 & ~n1086;
  assign n1088 = ~n1080 & ~n1087;
  assign n1089 = ~n1079 & n1088;
  assign n1090 = ~n684 & ~n1089;
  assign n1091 = ~pi349  & pi477 ;
  assign n1092 = ~pi348  & pi476 ;
  assign n1093 = ~n1091 & ~n1092;
  assign n1094 = n1090 & n1093;
  assign n1095 = ~pi478  & n683;
  assign n1096 = pi351  & ~pi479 ;
  assign n1097 = pi349  & ~pi477 ;
  assign n1098 = ~pi476  & ~n1091;
  assign n1099 = pi348  & n1098;
  assign n1100 = ~n1097 & ~n1099;
  assign n1101 = ~n684 & ~n1100;
  assign n1102 = ~n1096 & ~n1101;
  assign n1103 = ~n1095 & n1102;
  assign n1104 = ~n1094 & n1103;
  assign n1105 = n680 & ~n1104;
  assign n1106 = ~n677 & n1105;
  assign n1107 = ~pi352  & pi480 ;
  assign n1108 = n1106 & ~n1107;
  assign n1109 = pi355  & ~pi483 ;
  assign n1110 = pi354  & ~pi482 ;
  assign n1111 = pi353  & ~pi481 ;
  assign n1112 = ~pi480  & ~n677;
  assign n1113 = pi352  & n1112;
  assign n1114 = ~n1111 & ~n1113;
  assign n1115 = ~n1110 & n1114;
  assign n1116 = n680 & ~n1115;
  assign n1117 = ~n1109 & ~n1116;
  assign n1118 = ~n1108 & n1117;
  assign n1119 = ~n676 & ~n1118;
  assign n1120 = ~pi357  & pi485 ;
  assign n1121 = ~pi356  & pi484 ;
  assign n1122 = ~n1120 & ~n1121;
  assign n1123 = n1119 & n1122;
  assign n1124 = ~pi486  & n675;
  assign n1125 = pi359  & ~pi487 ;
  assign n1126 = pi357  & ~pi485 ;
  assign n1127 = ~pi484  & ~n1120;
  assign n1128 = pi356  & n1127;
  assign n1129 = ~n1126 & ~n1128;
  assign n1130 = ~n676 & ~n1129;
  assign n1131 = ~n1125 & ~n1130;
  assign n1132 = ~n1124 & n1131;
  assign n1133 = ~n1123 & n1132;
  assign n1134 = n672 & ~n1133;
  assign n1135 = ~n669 & n1134;
  assign n1136 = ~pi360  & pi488 ;
  assign n1137 = n1135 & ~n1136;
  assign n1138 = pi363  & ~pi491 ;
  assign n1139 = pi362  & ~pi490 ;
  assign n1140 = pi361  & ~pi489 ;
  assign n1141 = ~pi488  & ~n669;
  assign n1142 = pi360  & n1141;
  assign n1143 = ~n1140 & ~n1142;
  assign n1144 = ~n1139 & n1143;
  assign n1145 = n672 & ~n1144;
  assign n1146 = ~n1138 & ~n1145;
  assign n1147 = ~n1137 & n1146;
  assign n1148 = ~n668 & ~n1147;
  assign n1149 = ~pi365  & pi493 ;
  assign n1150 = ~pi364  & pi492 ;
  assign n1151 = ~n1149 & ~n1150;
  assign n1152 = n1148 & n1151;
  assign n1153 = ~pi494  & n667;
  assign n1154 = pi367  & ~pi495 ;
  assign n1155 = pi365  & ~pi493 ;
  assign n1156 = ~pi492  & ~n1149;
  assign n1157 = pi364  & n1156;
  assign n1158 = ~n1155 & ~n1157;
  assign n1159 = ~n668 & ~n1158;
  assign n1160 = ~n1154 & ~n1159;
  assign n1161 = ~n1153 & n1160;
  assign n1162 = ~n1152 & n1161;
  assign n1163 = n664 & ~n1162;
  assign n1164 = ~n661 & n1163;
  assign n1165 = ~pi368  & pi496 ;
  assign n1166 = n1164 & ~n1165;
  assign n1167 = pi371  & ~pi499 ;
  assign n1168 = pi370  & ~pi498 ;
  assign n1169 = pi369  & ~pi497 ;
  assign n1170 = ~pi496  & ~n661;
  assign n1171 = pi368  & n1170;
  assign n1172 = ~n1169 & ~n1171;
  assign n1173 = ~n1168 & n1172;
  assign n1174 = n664 & ~n1173;
  assign n1175 = ~n1167 & ~n1174;
  assign n1176 = ~n1166 & n1175;
  assign n1177 = ~n660 & ~n1176;
  assign n1178 = ~pi373  & pi501 ;
  assign n1179 = ~pi372  & pi500 ;
  assign n1180 = ~n1178 & ~n1179;
  assign n1181 = n1177 & n1180;
  assign n1182 = ~pi502  & n659;
  assign n1183 = pi375  & ~pi503 ;
  assign n1184 = pi373  & ~pi501 ;
  assign n1185 = ~pi500  & ~n1178;
  assign n1186 = pi372  & n1185;
  assign n1187 = ~n1184 & ~n1186;
  assign n1188 = ~n660 & ~n1187;
  assign n1189 = ~n1183 & ~n1188;
  assign n1190 = ~n1182 & n1189;
  assign n1191 = ~n1181 & n1190;
  assign n1192 = n656 & ~n1191;
  assign n1193 = ~n653 & n1192;
  assign n1194 = ~pi376  & pi504 ;
  assign n1195 = n1193 & ~n1194;
  assign n1196 = pi379  & ~pi507 ;
  assign n1197 = pi378  & ~pi506 ;
  assign n1198 = pi377  & ~pi505 ;
  assign n1199 = ~pi504  & ~n653;
  assign n1200 = pi376  & n1199;
  assign n1201 = ~n1198 & ~n1200;
  assign n1202 = ~n1197 & n1201;
  assign n1203 = n656 & ~n1202;
  assign n1204 = ~n1196 & ~n1203;
  assign n1205 = ~n1195 & n1204;
  assign n1206 = n646 & ~n1205;
  assign n1207 = ~pi380  & pi508 ;
  assign n1208 = n1206 & ~n1207;
  assign n1209 = n652 & ~n1208;
  assign n1210 = pi383  & ~pi511 ;
  assign n1211 = ~n1209 & ~n1210;
  assign n1212 = ~n643 & ~n1211;
  assign n1213 = pi384  & n1212;
  assign n1214 = pi256  & ~n1212;
  assign n1215 = ~n1213 & ~n1214;
  assign n1216 = pi383  & pi511 ;
  assign n1217 = pi127  & pi255 ;
  assign n1218 = ~n1216 & n1217;
  assign n1219 = ~pi127  & pi255 ;
  assign n1220 = pi127  & ~pi255 ;
  assign n1221 = ~pi126  & pi254 ;
  assign n1222 = ~pi125  & pi253 ;
  assign n1223 = ~n1221 & ~n1222;
  assign n1224 = pi124  & ~pi252 ;
  assign n1225 = pi125  & ~pi253 ;
  assign n1226 = ~n1224 & ~n1225;
  assign n1227 = n1223 & ~n1226;
  assign n1228 = pi126  & ~pi254 ;
  assign n1229 = ~n1227 & ~n1228;
  assign n1230 = ~n1220 & ~n1229;
  assign n1231 = ~pi121  & pi249 ;
  assign n1232 = ~pi123  & pi251 ;
  assign n1233 = ~pi122  & pi250 ;
  assign n1234 = ~n1232 & ~n1233;
  assign n1235 = ~pi119  & pi247 ;
  assign n1236 = ~pi246  & ~n1235;
  assign n1237 = pi118  & ~n1235;
  assign n1238 = ~n1236 & ~n1237;
  assign n1239 = ~pi113  & pi241 ;
  assign n1240 = ~pi115  & pi243 ;
  assign n1241 = ~pi114  & pi242 ;
  assign n1242 = ~n1240 & ~n1241;
  assign n1243 = ~pi111  & pi239 ;
  assign n1244 = ~pi238  & ~n1243;
  assign n1245 = pi110  & ~n1243;
  assign n1246 = ~n1244 & ~n1245;
  assign n1247 = ~pi105  & pi233 ;
  assign n1248 = ~pi107  & pi235 ;
  assign n1249 = ~pi106  & pi234 ;
  assign n1250 = ~n1248 & ~n1249;
  assign n1251 = ~pi103  & pi231 ;
  assign n1252 = ~pi230  & ~n1251;
  assign n1253 = pi102  & ~n1251;
  assign n1254 = ~n1252 & ~n1253;
  assign n1255 = ~pi97  & pi225 ;
  assign n1256 = ~pi99  & pi227 ;
  assign n1257 = ~pi98  & pi226 ;
  assign n1258 = ~n1256 & ~n1257;
  assign n1259 = ~pi95  & pi223 ;
  assign n1260 = ~pi222  & ~n1259;
  assign n1261 = pi94  & ~n1259;
  assign n1262 = ~n1260 & ~n1261;
  assign n1263 = ~pi89  & pi217 ;
  assign n1264 = ~pi91  & pi219 ;
  assign n1265 = ~pi90  & pi218 ;
  assign n1266 = ~n1264 & ~n1265;
  assign n1267 = ~pi87  & pi215 ;
  assign n1268 = ~pi214  & ~n1267;
  assign n1269 = pi86  & ~n1267;
  assign n1270 = ~n1268 & ~n1269;
  assign n1271 = ~pi81  & pi209 ;
  assign n1272 = ~pi83  & pi211 ;
  assign n1273 = ~pi82  & pi210 ;
  assign n1274 = ~n1272 & ~n1273;
  assign n1275 = ~pi79  & pi207 ;
  assign n1276 = ~pi206  & ~n1275;
  assign n1277 = pi78  & ~n1275;
  assign n1278 = ~n1276 & ~n1277;
  assign n1279 = ~pi73  & pi201 ;
  assign n1280 = ~pi75  & pi203 ;
  assign n1281 = ~pi74  & pi202 ;
  assign n1282 = ~n1280 & ~n1281;
  assign n1283 = ~pi71  & pi199 ;
  assign n1284 = ~pi198  & ~n1283;
  assign n1285 = pi70  & ~n1283;
  assign n1286 = ~n1284 & ~n1285;
  assign n1287 = ~pi65  & pi193 ;
  assign n1288 = ~pi67  & pi195 ;
  assign n1289 = ~pi66  & pi194 ;
  assign n1290 = ~n1288 & ~n1289;
  assign n1291 = pi59  & ~pi187 ;
  assign n1292 = ~pi59  & pi187 ;
  assign n1293 = ~pi58  & pi186 ;
  assign n1294 = ~n1292 & ~n1293;
  assign n1295 = pi58  & ~pi186 ;
  assign n1296 = pi57  & ~pi185 ;
  assign n1297 = ~pi57  & pi185 ;
  assign n1298 = ~pi184  & ~n1297;
  assign n1299 = pi56  & n1298;
  assign n1300 = ~n1296 & ~n1299;
  assign n1301 = ~n1295 & n1300;
  assign n1302 = n1294 & ~n1301;
  assign n1303 = ~n1291 & ~n1302;
  assign n1304 = ~pi63  & pi191 ;
  assign n1305 = ~pi190  & ~n1304;
  assign n1306 = pi62  & ~n1304;
  assign n1307 = ~n1305 & ~n1306;
  assign n1308 = ~pi61  & pi189 ;
  assign n1309 = ~pi60  & pi188 ;
  assign n1310 = ~n1308 & ~n1309;
  assign n1311 = ~n1307 & n1310;
  assign n1312 = ~n1303 & n1311;
  assign n1313 = ~pi190  & n1306;
  assign n1314 = pi63  & ~pi191 ;
  assign n1315 = pi61  & ~pi189 ;
  assign n1316 = ~pi188  & ~n1308;
  assign n1317 = pi60  & n1316;
  assign n1318 = ~n1315 & ~n1317;
  assign n1319 = ~n1307 & ~n1318;
  assign n1320 = ~pi56  & pi184 ;
  assign n1321 = n1311 & ~n1320;
  assign n1322 = pi55  & ~pi183 ;
  assign n1323 = ~pi55  & pi183 ;
  assign n1324 = ~pi54  & pi182 ;
  assign n1325 = ~n1323 & ~n1324;
  assign n1326 = pi54  & ~pi182 ;
  assign n1327 = pi53  & ~pi181 ;
  assign n1328 = ~pi53  & pi181 ;
  assign n1329 = ~pi180  & ~n1328;
  assign n1330 = pi52  & n1329;
  assign n1331 = ~n1327 & ~n1330;
  assign n1332 = ~n1326 & n1331;
  assign n1333 = n1325 & ~n1332;
  assign n1334 = pi51  & ~pi179 ;
  assign n1335 = ~pi51  & pi179 ;
  assign n1336 = ~pi50  & pi178 ;
  assign n1337 = ~n1335 & ~n1336;
  assign n1338 = pi50  & ~pi178 ;
  assign n1339 = pi49  & ~pi177 ;
  assign n1340 = ~pi49  & pi177 ;
  assign n1341 = ~pi176  & ~n1340;
  assign n1342 = pi48  & n1341;
  assign n1343 = ~n1339 & ~n1342;
  assign n1344 = ~n1338 & n1343;
  assign n1345 = n1337 & ~n1344;
  assign n1346 = ~n1334 & ~n1345;
  assign n1347 = ~pi52  & pi180 ;
  assign n1348 = n1325 & ~n1347;
  assign n1349 = ~n1328 & n1348;
  assign n1350 = ~n1346 & n1349;
  assign n1351 = ~n1333 & ~n1350;
  assign n1352 = ~pi48  & pi176 ;
  assign n1353 = n1337 & ~n1352;
  assign n1354 = pi43  & ~pi171 ;
  assign n1355 = ~pi43  & pi171 ;
  assign n1356 = ~pi42  & pi170 ;
  assign n1357 = ~n1355 & ~n1356;
  assign n1358 = pi42  & ~pi170 ;
  assign n1359 = pi41  & ~pi169 ;
  assign n1360 = ~pi41  & pi169 ;
  assign n1361 = ~pi168  & ~n1360;
  assign n1362 = pi40  & n1361;
  assign n1363 = ~n1359 & ~n1362;
  assign n1364 = ~n1358 & n1363;
  assign n1365 = n1357 & ~n1364;
  assign n1366 = ~n1354 & ~n1365;
  assign n1367 = ~pi47  & pi175 ;
  assign n1368 = ~pi174  & ~n1367;
  assign n1369 = pi46  & ~n1367;
  assign n1370 = ~n1368 & ~n1369;
  assign n1371 = ~pi45  & pi173 ;
  assign n1372 = ~pi44  & pi172 ;
  assign n1373 = ~n1371 & ~n1372;
  assign n1374 = ~n1370 & n1373;
  assign n1375 = ~n1366 & n1374;
  assign n1376 = ~pi174  & n1369;
  assign n1377 = pi47  & ~pi175 ;
  assign n1378 = pi45  & ~pi173 ;
  assign n1379 = ~pi172  & ~n1371;
  assign n1380 = pi44  & n1379;
  assign n1381 = ~n1378 & ~n1380;
  assign n1382 = ~n1370 & ~n1381;
  assign n1383 = ~pi40  & pi168 ;
  assign n1384 = n1374 & ~n1383;
  assign n1385 = ~pi39  & pi167 ;
  assign n1386 = ~pi166  & ~n1385;
  assign n1387 = pi38  & ~n1385;
  assign n1388 = ~n1386 & ~n1387;
  assign n1389 = ~pi37  & pi165 ;
  assign n1390 = ~pi36  & pi164 ;
  assign n1391 = ~n1389 & ~n1390;
  assign n1392 = ~n1388 & n1391;
  assign n1393 = pi31  & ~pi159 ;
  assign n1394 = pi30  & ~pi158 ;
  assign n1395 = ~pi30  & pi158 ;
  assign n1396 = pi29  & ~pi157 ;
  assign n1397 = ~pi29  & pi157 ;
  assign n1398 = pi28  & ~pi156 ;
  assign n1399 = ~pi28  & pi156 ;
  assign n1400 = pi27  & ~pi155 ;
  assign n1401 = ~pi27  & pi155 ;
  assign n1402 = pi26  & ~pi154 ;
  assign n1403 = ~pi26  & pi154 ;
  assign n1404 = pi25  & ~pi153 ;
  assign n1405 = ~pi25  & pi153 ;
  assign n1406 = pi24  & ~pi152 ;
  assign n1407 = ~pi24  & pi152 ;
  assign n1408 = pi23  & ~pi151 ;
  assign n1409 = ~pi23  & pi151 ;
  assign n1410 = pi22  & ~pi150 ;
  assign n1411 = ~pi22  & pi150 ;
  assign n1412 = pi21  & ~pi149 ;
  assign n1413 = ~pi21  & pi149 ;
  assign n1414 = pi20  & ~pi148 ;
  assign n1415 = ~pi20  & pi148 ;
  assign n1416 = pi19  & ~pi147 ;
  assign n1417 = ~pi19  & pi147 ;
  assign n1418 = pi18  & ~pi146 ;
  assign n1419 = ~pi18  & pi146 ;
  assign n1420 = pi17  & ~pi145 ;
  assign n1421 = ~pi17  & pi145 ;
  assign n1422 = pi16  & ~pi144 ;
  assign n1423 = ~pi16  & pi144 ;
  assign n1424 = pi15  & ~pi143 ;
  assign n1425 = ~pi15  & pi143 ;
  assign n1426 = pi14  & ~pi142 ;
  assign n1427 = ~pi14  & pi142 ;
  assign n1428 = pi13  & ~pi141 ;
  assign n1429 = ~pi13  & pi141 ;
  assign n1430 = pi12  & ~pi140 ;
  assign n1431 = ~pi12  & pi140 ;
  assign n1432 = pi11  & ~pi139 ;
  assign n1433 = ~pi11  & pi139 ;
  assign n1434 = pi10  & ~pi138 ;
  assign n1435 = ~pi10  & pi138 ;
  assign n1436 = pi9  & ~pi137 ;
  assign n1437 = ~pi9  & pi137 ;
  assign n1438 = pi8  & ~pi136 ;
  assign n1439 = ~pi8  & pi136 ;
  assign n1440 = pi7  & ~pi135 ;
  assign n1441 = ~pi7  & pi135 ;
  assign n1442 = pi6  & ~pi134 ;
  assign n1443 = ~pi6  & pi134 ;
  assign n1444 = pi5  & ~pi133 ;
  assign n1445 = ~pi5  & pi133 ;
  assign n1446 = pi4  & ~pi132 ;
  assign n1447 = ~pi4  & pi132 ;
  assign n1448 = pi3  & ~pi131 ;
  assign n1449 = ~pi3  & pi131 ;
  assign n1450 = pi2  & ~pi130 ;
  assign n1451 = ~pi2  & pi130 ;
  assign n1452 = pi0  & ~pi128 ;
  assign n1453 = ~pi1  & pi129 ;
  assign n1454 = n1452 & ~n1453;
  assign n1455 = pi1  & ~pi129 ;
  assign n1456 = ~n1454 & ~n1455;
  assign n1457 = ~n1451 & ~n1456;
  assign n1458 = ~n1450 & ~n1457;
  assign n1459 = ~n1449 & ~n1458;
  assign n1460 = ~n1448 & ~n1459;
  assign n1461 = ~n1447 & ~n1460;
  assign n1462 = ~n1446 & ~n1461;
  assign n1463 = ~n1445 & ~n1462;
  assign n1464 = ~n1444 & ~n1463;
  assign n1465 = ~n1443 & ~n1464;
  assign n1466 = ~n1442 & ~n1465;
  assign n1467 = ~n1441 & ~n1466;
  assign n1468 = ~n1440 & ~n1467;
  assign n1469 = ~n1439 & ~n1468;
  assign n1470 = ~n1438 & ~n1469;
  assign n1471 = ~n1437 & ~n1470;
  assign n1472 = ~n1436 & ~n1471;
  assign n1473 = ~n1435 & ~n1472;
  assign n1474 = ~n1434 & ~n1473;
  assign n1475 = ~n1433 & ~n1474;
  assign n1476 = ~n1432 & ~n1475;
  assign n1477 = ~n1431 & ~n1476;
  assign n1478 = ~n1430 & ~n1477;
  assign n1479 = ~n1429 & ~n1478;
  assign n1480 = ~n1428 & ~n1479;
  assign n1481 = ~n1427 & ~n1480;
  assign n1482 = ~n1426 & ~n1481;
  assign n1483 = ~n1425 & ~n1482;
  assign n1484 = ~n1424 & ~n1483;
  assign n1485 = ~n1423 & ~n1484;
  assign n1486 = ~n1422 & ~n1485;
  assign n1487 = ~n1421 & ~n1486;
  assign n1488 = ~n1420 & ~n1487;
  assign n1489 = ~n1419 & ~n1488;
  assign n1490 = ~n1418 & ~n1489;
  assign n1491 = ~n1417 & ~n1490;
  assign n1492 = ~n1416 & ~n1491;
  assign n1493 = ~n1415 & ~n1492;
  assign n1494 = ~n1414 & ~n1493;
  assign n1495 = ~n1413 & ~n1494;
  assign n1496 = ~n1412 & ~n1495;
  assign n1497 = ~n1411 & ~n1496;
  assign n1498 = ~n1410 & ~n1497;
  assign n1499 = ~n1409 & ~n1498;
  assign n1500 = ~n1408 & ~n1499;
  assign n1501 = ~n1407 & ~n1500;
  assign n1502 = ~n1406 & ~n1501;
  assign n1503 = ~n1405 & ~n1502;
  assign n1504 = ~n1404 & ~n1503;
  assign n1505 = ~n1403 & ~n1504;
  assign n1506 = ~n1402 & ~n1505;
  assign n1507 = ~n1401 & ~n1506;
  assign n1508 = ~n1400 & ~n1507;
  assign n1509 = ~n1399 & ~n1508;
  assign n1510 = ~n1398 & ~n1509;
  assign n1511 = ~n1397 & ~n1510;
  assign n1512 = ~n1396 & ~n1511;
  assign n1513 = ~n1395 & ~n1512;
  assign n1514 = ~n1394 & ~n1513;
  assign n1515 = ~n1393 & n1514;
  assign n1516 = n1392 & ~n1515;
  assign n1517 = ~pi33  & pi161 ;
  assign n1518 = ~pi32  & pi160 ;
  assign n1519 = ~pi35  & pi163 ;
  assign n1520 = ~pi34  & pi162 ;
  assign n1521 = ~n1519 & ~n1520;
  assign n1522 = ~pi31  & pi159 ;
  assign n1523 = n1521 & ~n1522;
  assign n1524 = ~n1518 & n1523;
  assign n1525 = ~n1517 & n1524;
  assign n1526 = n1516 & n1525;
  assign n1527 = pi35  & ~pi163 ;
  assign n1528 = pi34  & ~pi162 ;
  assign n1529 = pi33  & ~pi161 ;
  assign n1530 = ~pi160  & ~n1517;
  assign n1531 = pi32  & n1530;
  assign n1532 = ~n1529 & ~n1531;
  assign n1533 = ~n1528 & n1532;
  assign n1534 = n1521 & ~n1533;
  assign n1535 = ~n1527 & ~n1534;
  assign n1536 = n1392 & ~n1535;
  assign n1537 = pi39  & ~pi167 ;
  assign n1538 = pi37  & ~pi165 ;
  assign n1539 = ~pi164  & ~n1389;
  assign n1540 = pi36  & n1539;
  assign n1541 = ~n1538 & ~n1540;
  assign n1542 = ~n1388 & ~n1541;
  assign n1543 = ~n1537 & ~n1542;
  assign n1544 = ~n1536 & n1543;
  assign n1545 = ~n1526 & n1544;
  assign n1546 = pi38  & n1386;
  assign n1547 = n1545 & ~n1546;
  assign n1548 = n1357 & ~n1547;
  assign n1549 = ~n1360 & n1548;
  assign n1550 = n1384 & n1549;
  assign n1551 = ~n1382 & ~n1550;
  assign n1552 = ~n1377 & n1551;
  assign n1553 = ~n1376 & n1552;
  assign n1554 = ~n1375 & n1553;
  assign n1555 = n1349 & ~n1554;
  assign n1556 = ~n1340 & n1555;
  assign n1557 = n1353 & n1556;
  assign n1558 = n1351 & ~n1557;
  assign n1559 = ~n1322 & n1558;
  assign n1560 = n1294 & ~n1559;
  assign n1561 = ~n1297 & n1560;
  assign n1562 = n1321 & n1561;
  assign n1563 = ~n1319 & ~n1562;
  assign n1564 = ~n1314 & n1563;
  assign n1565 = ~n1313 & n1564;
  assign n1566 = ~n1312 & n1565;
  assign n1567 = n1290 & ~n1566;
  assign n1568 = ~n1287 & n1567;
  assign n1569 = ~pi64  & pi192 ;
  assign n1570 = n1568 & ~n1569;
  assign n1571 = pi67  & ~pi195 ;
  assign n1572 = pi66  & ~pi194 ;
  assign n1573 = pi65  & ~pi193 ;
  assign n1574 = ~pi192  & ~n1287;
  assign n1575 = pi64  & n1574;
  assign n1576 = ~n1573 & ~n1575;
  assign n1577 = ~n1572 & n1576;
  assign n1578 = n1290 & ~n1577;
  assign n1579 = ~n1571 & ~n1578;
  assign n1580 = ~n1570 & n1579;
  assign n1581 = ~n1286 & ~n1580;
  assign n1582 = ~pi69  & pi197 ;
  assign n1583 = ~pi68  & pi196 ;
  assign n1584 = ~n1582 & ~n1583;
  assign n1585 = n1581 & n1584;
  assign n1586 = ~pi198  & n1285;
  assign n1587 = pi71  & ~pi199 ;
  assign n1588 = pi69  & ~pi197 ;
  assign n1589 = ~pi196  & ~n1582;
  assign n1590 = pi68  & n1589;
  assign n1591 = ~n1588 & ~n1590;
  assign n1592 = ~n1286 & ~n1591;
  assign n1593 = ~n1587 & ~n1592;
  assign n1594 = ~n1586 & n1593;
  assign n1595 = ~n1585 & n1594;
  assign n1596 = n1282 & ~n1595;
  assign n1597 = ~n1279 & n1596;
  assign n1598 = ~pi72  & pi200 ;
  assign n1599 = n1597 & ~n1598;
  assign n1600 = pi75  & ~pi203 ;
  assign n1601 = pi74  & ~pi202 ;
  assign n1602 = pi73  & ~pi201 ;
  assign n1603 = ~pi200  & ~n1279;
  assign n1604 = pi72  & n1603;
  assign n1605 = ~n1602 & ~n1604;
  assign n1606 = ~n1601 & n1605;
  assign n1607 = n1282 & ~n1606;
  assign n1608 = ~n1600 & ~n1607;
  assign n1609 = ~n1599 & n1608;
  assign n1610 = ~n1278 & ~n1609;
  assign n1611 = ~pi77  & pi205 ;
  assign n1612 = ~pi76  & pi204 ;
  assign n1613 = ~n1611 & ~n1612;
  assign n1614 = n1610 & n1613;
  assign n1615 = ~pi206  & n1277;
  assign n1616 = pi79  & ~pi207 ;
  assign n1617 = pi77  & ~pi205 ;
  assign n1618 = ~pi204  & ~n1611;
  assign n1619 = pi76  & n1618;
  assign n1620 = ~n1617 & ~n1619;
  assign n1621 = ~n1278 & ~n1620;
  assign n1622 = ~n1616 & ~n1621;
  assign n1623 = ~n1615 & n1622;
  assign n1624 = ~n1614 & n1623;
  assign n1625 = n1274 & ~n1624;
  assign n1626 = ~n1271 & n1625;
  assign n1627 = ~pi80  & pi208 ;
  assign n1628 = n1626 & ~n1627;
  assign n1629 = pi83  & ~pi211 ;
  assign n1630 = pi82  & ~pi210 ;
  assign n1631 = pi81  & ~pi209 ;
  assign n1632 = ~pi208  & ~n1271;
  assign n1633 = pi80  & n1632;
  assign n1634 = ~n1631 & ~n1633;
  assign n1635 = ~n1630 & n1634;
  assign n1636 = n1274 & ~n1635;
  assign n1637 = ~n1629 & ~n1636;
  assign n1638 = ~n1628 & n1637;
  assign n1639 = ~n1270 & ~n1638;
  assign n1640 = ~pi85  & pi213 ;
  assign n1641 = ~pi84  & pi212 ;
  assign n1642 = ~n1640 & ~n1641;
  assign n1643 = n1639 & n1642;
  assign n1644 = ~pi214  & n1269;
  assign n1645 = pi87  & ~pi215 ;
  assign n1646 = pi85  & ~pi213 ;
  assign n1647 = ~pi212  & ~n1640;
  assign n1648 = pi84  & n1647;
  assign n1649 = ~n1646 & ~n1648;
  assign n1650 = ~n1270 & ~n1649;
  assign n1651 = ~n1645 & ~n1650;
  assign n1652 = ~n1644 & n1651;
  assign n1653 = ~n1643 & n1652;
  assign n1654 = n1266 & ~n1653;
  assign n1655 = ~n1263 & n1654;
  assign n1656 = ~pi88  & pi216 ;
  assign n1657 = n1655 & ~n1656;
  assign n1658 = pi91  & ~pi219 ;
  assign n1659 = pi90  & ~pi218 ;
  assign n1660 = pi89  & ~pi217 ;
  assign n1661 = ~pi216  & ~n1263;
  assign n1662 = pi88  & n1661;
  assign n1663 = ~n1660 & ~n1662;
  assign n1664 = ~n1659 & n1663;
  assign n1665 = n1266 & ~n1664;
  assign n1666 = ~n1658 & ~n1665;
  assign n1667 = ~n1657 & n1666;
  assign n1668 = ~n1262 & ~n1667;
  assign n1669 = ~pi93  & pi221 ;
  assign n1670 = ~pi92  & pi220 ;
  assign n1671 = ~n1669 & ~n1670;
  assign n1672 = n1668 & n1671;
  assign n1673 = ~pi222  & n1261;
  assign n1674 = pi95  & ~pi223 ;
  assign n1675 = pi93  & ~pi221 ;
  assign n1676 = ~pi220  & ~n1669;
  assign n1677 = pi92  & n1676;
  assign n1678 = ~n1675 & ~n1677;
  assign n1679 = ~n1262 & ~n1678;
  assign n1680 = ~n1674 & ~n1679;
  assign n1681 = ~n1673 & n1680;
  assign n1682 = ~n1672 & n1681;
  assign n1683 = n1258 & ~n1682;
  assign n1684 = ~n1255 & n1683;
  assign n1685 = ~pi96  & pi224 ;
  assign n1686 = n1684 & ~n1685;
  assign n1687 = pi99  & ~pi227 ;
  assign n1688 = pi98  & ~pi226 ;
  assign n1689 = pi97  & ~pi225 ;
  assign n1690 = ~pi224  & ~n1255;
  assign n1691 = pi96  & n1690;
  assign n1692 = ~n1689 & ~n1691;
  assign n1693 = ~n1688 & n1692;
  assign n1694 = n1258 & ~n1693;
  assign n1695 = ~n1687 & ~n1694;
  assign n1696 = ~n1686 & n1695;
  assign n1697 = ~n1254 & ~n1696;
  assign n1698 = ~pi101  & pi229 ;
  assign n1699 = ~pi100  & pi228 ;
  assign n1700 = ~n1698 & ~n1699;
  assign n1701 = n1697 & n1700;
  assign n1702 = ~pi230  & n1253;
  assign n1703 = pi103  & ~pi231 ;
  assign n1704 = pi101  & ~pi229 ;
  assign n1705 = ~pi228  & ~n1698;
  assign n1706 = pi100  & n1705;
  assign n1707 = ~n1704 & ~n1706;
  assign n1708 = ~n1254 & ~n1707;
  assign n1709 = ~n1703 & ~n1708;
  assign n1710 = ~n1702 & n1709;
  assign n1711 = ~n1701 & n1710;
  assign n1712 = n1250 & ~n1711;
  assign n1713 = ~n1247 & n1712;
  assign n1714 = ~pi104  & pi232 ;
  assign n1715 = n1713 & ~n1714;
  assign n1716 = pi107  & ~pi235 ;
  assign n1717 = pi106  & ~pi234 ;
  assign n1718 = pi105  & ~pi233 ;
  assign n1719 = ~pi232  & ~n1247;
  assign n1720 = pi104  & n1719;
  assign n1721 = ~n1718 & ~n1720;
  assign n1722 = ~n1717 & n1721;
  assign n1723 = n1250 & ~n1722;
  assign n1724 = ~n1716 & ~n1723;
  assign n1725 = ~n1715 & n1724;
  assign n1726 = ~n1246 & ~n1725;
  assign n1727 = ~pi109  & pi237 ;
  assign n1728 = ~pi108  & pi236 ;
  assign n1729 = ~n1727 & ~n1728;
  assign n1730 = n1726 & n1729;
  assign n1731 = ~pi238  & n1245;
  assign n1732 = pi111  & ~pi239 ;
  assign n1733 = pi109  & ~pi237 ;
  assign n1734 = ~pi236  & ~n1727;
  assign n1735 = pi108  & n1734;
  assign n1736 = ~n1733 & ~n1735;
  assign n1737 = ~n1246 & ~n1736;
  assign n1738 = ~n1732 & ~n1737;
  assign n1739 = ~n1731 & n1738;
  assign n1740 = ~n1730 & n1739;
  assign n1741 = n1242 & ~n1740;
  assign n1742 = ~n1239 & n1741;
  assign n1743 = ~pi112  & pi240 ;
  assign n1744 = n1742 & ~n1743;
  assign n1745 = pi115  & ~pi243 ;
  assign n1746 = pi114  & ~pi242 ;
  assign n1747 = pi113  & ~pi241 ;
  assign n1748 = ~pi240  & ~n1239;
  assign n1749 = pi112  & n1748;
  assign n1750 = ~n1747 & ~n1749;
  assign n1751 = ~n1746 & n1750;
  assign n1752 = n1242 & ~n1751;
  assign n1753 = ~n1745 & ~n1752;
  assign n1754 = ~n1744 & n1753;
  assign n1755 = ~n1238 & ~n1754;
  assign n1756 = ~pi117  & pi245 ;
  assign n1757 = ~pi116  & pi244 ;
  assign n1758 = ~n1756 & ~n1757;
  assign n1759 = n1755 & n1758;
  assign n1760 = ~pi246  & n1237;
  assign n1761 = pi119  & ~pi247 ;
  assign n1762 = pi117  & ~pi245 ;
  assign n1763 = ~pi244  & ~n1756;
  assign n1764 = pi116  & n1763;
  assign n1765 = ~n1762 & ~n1764;
  assign n1766 = ~n1238 & ~n1765;
  assign n1767 = ~n1761 & ~n1766;
  assign n1768 = ~n1760 & n1767;
  assign n1769 = ~n1759 & n1768;
  assign n1770 = n1234 & ~n1769;
  assign n1771 = ~n1231 & n1770;
  assign n1772 = ~pi120  & pi248 ;
  assign n1773 = n1771 & ~n1772;
  assign n1774 = pi123  & ~pi251 ;
  assign n1775 = pi122  & ~pi250 ;
  assign n1776 = pi121  & ~pi249 ;
  assign n1777 = ~pi248  & ~n1231;
  assign n1778 = pi120  & n1777;
  assign n1779 = ~n1776 & ~n1778;
  assign n1780 = ~n1775 & n1779;
  assign n1781 = n1234 & ~n1780;
  assign n1782 = ~n1774 & ~n1781;
  assign n1783 = ~n1773 & n1782;
  assign n1784 = n1223 & ~n1783;
  assign n1785 = ~pi124  & pi252 ;
  assign n1786 = n1784 & ~n1785;
  assign n1787 = ~n1220 & n1786;
  assign n1788 = ~n1230 & ~n1787;
  assign n1789 = ~n1219 & n1788;
  assign n1790 = pi254  & n1789;
  assign n1791 = pi126  & ~n1789;
  assign n1792 = ~n1790 & ~n1791;
  assign n1793 = pi510  & n1212;
  assign n1794 = pi382  & ~n1212;
  assign n1795 = ~n1793 & ~n1794;
  assign n1796 = n1792 & ~n1795;
  assign n1797 = pi253  & n1789;
  assign n1798 = pi125  & ~n1789;
  assign n1799 = ~n1797 & ~n1798;
  assign n1800 = pi509  & n1212;
  assign n1801 = pi381  & ~n1212;
  assign n1802 = ~n1800 & ~n1801;
  assign n1803 = n1799 & ~n1802;
  assign n1804 = ~n1796 & ~n1803;
  assign n1805 = pi252  & n1789;
  assign n1806 = pi124  & ~n1789;
  assign n1807 = ~n1805 & ~n1806;
  assign n1808 = pi508  & n1212;
  assign n1809 = pi380  & ~n1212;
  assign n1810 = ~n1808 & ~n1809;
  assign n1811 = ~n1807 & n1810;
  assign n1812 = ~n1799 & n1802;
  assign n1813 = ~n1811 & ~n1812;
  assign n1814 = n1804 & ~n1813;
  assign n1815 = ~n1792 & n1795;
  assign n1816 = ~n1814 & ~n1815;
  assign n1817 = ~n1218 & ~n1816;
  assign n1818 = n1216 & ~n1217;
  assign n1819 = n1807 & ~n1810;
  assign n1820 = pi251  & n1789;
  assign n1821 = pi123  & ~n1789;
  assign n1822 = ~n1820 & ~n1821;
  assign n1823 = pi507  & n1212;
  assign n1824 = pi379  & ~n1212;
  assign n1825 = ~n1823 & ~n1824;
  assign n1826 = n1822 & ~n1825;
  assign n1827 = pi506  & n1212;
  assign n1828 = pi378  & ~n1212;
  assign n1829 = ~n1827 & ~n1828;
  assign n1830 = pi250  & n1789;
  assign n1831 = pi122  & ~n1789;
  assign n1832 = ~n1830 & ~n1831;
  assign n1833 = ~n1829 & n1832;
  assign n1834 = ~n1826 & ~n1833;
  assign n1835 = pi245  & n1789;
  assign n1836 = pi117  & ~n1789;
  assign n1837 = ~n1835 & ~n1836;
  assign n1838 = pi501  & n1212;
  assign n1839 = pi373  & ~n1212;
  assign n1840 = ~n1838 & ~n1839;
  assign n1841 = ~n1837 & n1840;
  assign n1842 = pi244  & n1789;
  assign n1843 = pi116  & ~n1789;
  assign n1844 = ~n1842 & ~n1843;
  assign n1845 = pi500  & n1212;
  assign n1846 = pi372  & ~n1212;
  assign n1847 = ~n1845 & ~n1846;
  assign n1848 = ~n1844 & n1847;
  assign n1849 = ~n1841 & ~n1848;
  assign n1850 = pi247  & n1789;
  assign n1851 = pi119  & ~n1789;
  assign n1852 = ~n1850 & ~n1851;
  assign n1853 = pi503  & n1212;
  assign n1854 = pi375  & ~n1212;
  assign n1855 = ~n1853 & ~n1854;
  assign n1856 = n1852 & ~n1855;
  assign n1857 = n1837 & ~n1840;
  assign n1858 = ~n1856 & ~n1857;
  assign n1859 = pi502  & n1212;
  assign n1860 = pi374  & ~n1212;
  assign n1861 = ~n1859 & ~n1860;
  assign n1862 = pi246  & n1789;
  assign n1863 = pi118  & ~n1789;
  assign n1864 = ~n1862 & ~n1863;
  assign n1865 = ~n1861 & n1864;
  assign n1866 = n1858 & ~n1865;
  assign n1867 = ~n1849 & n1866;
  assign n1868 = ~n1856 & ~n1864;
  assign n1869 = n1861 & n1868;
  assign n1870 = ~n1852 & n1855;
  assign n1871 = pi241  & n1789;
  assign n1872 = pi113  & ~n1789;
  assign n1873 = ~n1871 & ~n1872;
  assign n1874 = pi497  & n1212;
  assign n1875 = pi369  & ~n1212;
  assign n1876 = ~n1874 & ~n1875;
  assign n1877 = n1873 & ~n1876;
  assign n1878 = pi243  & n1789;
  assign n1879 = pi115  & ~n1789;
  assign n1880 = ~n1878 & ~n1879;
  assign n1881 = pi499  & n1212;
  assign n1882 = pi371  & ~n1212;
  assign n1883 = ~n1881 & ~n1882;
  assign n1884 = n1880 & ~n1883;
  assign n1885 = pi498  & n1212;
  assign n1886 = pi370  & ~n1212;
  assign n1887 = ~n1885 & ~n1886;
  assign n1888 = pi242  & n1789;
  assign n1889 = pi114  & ~n1789;
  assign n1890 = ~n1888 & ~n1889;
  assign n1891 = ~n1887 & n1890;
  assign n1892 = ~n1884 & ~n1891;
  assign n1893 = pi494  & n1212;
  assign n1894 = pi366  & ~n1212;
  assign n1895 = ~n1893 & ~n1894;
  assign n1896 = pi239  & n1789;
  assign n1897 = pi111  & ~n1789;
  assign n1898 = ~n1896 & ~n1897;
  assign n1899 = pi495  & n1212;
  assign n1900 = pi367  & ~n1212;
  assign n1901 = ~n1899 & ~n1900;
  assign n1902 = n1898 & ~n1901;
  assign n1903 = pi238  & n1789;
  assign n1904 = pi110  & ~n1789;
  assign n1905 = ~n1903 & ~n1904;
  assign n1906 = ~n1902 & ~n1905;
  assign n1907 = n1895 & n1906;
  assign n1908 = n1895 & ~n1902;
  assign n1909 = ~n1906 & ~n1908;
  assign n1910 = pi237  & n1789;
  assign n1911 = pi109  & ~n1789;
  assign n1912 = ~n1910 & ~n1911;
  assign n1913 = pi493  & n1212;
  assign n1914 = pi365  & ~n1212;
  assign n1915 = ~n1913 & ~n1914;
  assign n1916 = ~n1912 & n1915;
  assign n1917 = pi236  & n1789;
  assign n1918 = pi108  & ~n1789;
  assign n1919 = ~n1917 & ~n1918;
  assign n1920 = n1912 & ~n1915;
  assign n1921 = pi492  & n1212;
  assign n1922 = pi364  & ~n1212;
  assign n1923 = ~n1921 & ~n1922;
  assign n1924 = ~n1920 & n1923;
  assign n1925 = ~n1919 & n1924;
  assign n1926 = ~n1916 & ~n1925;
  assign n1927 = ~n1909 & ~n1926;
  assign n1928 = ~n1898 & n1901;
  assign n1929 = pi233  & n1789;
  assign n1930 = pi105  & ~n1789;
  assign n1931 = ~n1929 & ~n1930;
  assign n1932 = pi489  & n1212;
  assign n1933 = pi361  & ~n1212;
  assign n1934 = ~n1932 & ~n1933;
  assign n1935 = n1931 & ~n1934;
  assign n1936 = pi235  & n1789;
  assign n1937 = pi107  & ~n1789;
  assign n1938 = ~n1936 & ~n1937;
  assign n1939 = pi491  & n1212;
  assign n1940 = pi363  & ~n1212;
  assign n1941 = ~n1939 & ~n1940;
  assign n1942 = n1938 & ~n1941;
  assign n1943 = pi490  & n1212;
  assign n1944 = pi362  & ~n1212;
  assign n1945 = ~n1943 & ~n1944;
  assign n1946 = pi234  & n1789;
  assign n1947 = pi106  & ~n1789;
  assign n1948 = ~n1946 & ~n1947;
  assign n1949 = ~n1945 & n1948;
  assign n1950 = ~n1942 & ~n1949;
  assign n1951 = pi486  & n1212;
  assign n1952 = pi358  & ~n1212;
  assign n1953 = ~n1951 & ~n1952;
  assign n1954 = pi231  & n1789;
  assign n1955 = pi103  & ~n1789;
  assign n1956 = ~n1954 & ~n1955;
  assign n1957 = pi487  & n1212;
  assign n1958 = pi359  & ~n1212;
  assign n1959 = ~n1957 & ~n1958;
  assign n1960 = n1956 & ~n1959;
  assign n1961 = pi230  & n1789;
  assign n1962 = pi102  & ~n1789;
  assign n1963 = ~n1961 & ~n1962;
  assign n1964 = ~n1960 & ~n1963;
  assign n1965 = n1953 & n1964;
  assign n1966 = n1953 & ~n1960;
  assign n1967 = ~n1964 & ~n1966;
  assign n1968 = pi229  & n1789;
  assign n1969 = pi101  & ~n1789;
  assign n1970 = ~n1968 & ~n1969;
  assign n1971 = pi485  & n1212;
  assign n1972 = pi357  & ~n1212;
  assign n1973 = ~n1971 & ~n1972;
  assign n1974 = ~n1970 & n1973;
  assign n1975 = pi228  & n1789;
  assign n1976 = pi100  & ~n1789;
  assign n1977 = ~n1975 & ~n1976;
  assign n1978 = n1970 & ~n1973;
  assign n1979 = pi484  & n1212;
  assign n1980 = pi356  & ~n1212;
  assign n1981 = ~n1979 & ~n1980;
  assign n1982 = ~n1978 & n1981;
  assign n1983 = ~n1977 & n1982;
  assign n1984 = ~n1974 & ~n1983;
  assign n1985 = ~n1967 & ~n1984;
  assign n1986 = ~n1956 & n1959;
  assign n1987 = pi225  & n1789;
  assign n1988 = pi97  & ~n1789;
  assign n1989 = ~n1987 & ~n1988;
  assign n1990 = pi481  & n1212;
  assign n1991 = pi353  & ~n1212;
  assign n1992 = ~n1990 & ~n1991;
  assign n1993 = n1989 & ~n1992;
  assign n1994 = pi227  & n1789;
  assign n1995 = pi99  & ~n1789;
  assign n1996 = ~n1994 & ~n1995;
  assign n1997 = pi483  & n1212;
  assign n1998 = pi355  & ~n1212;
  assign n1999 = ~n1997 & ~n1998;
  assign n2000 = n1996 & ~n1999;
  assign n2001 = pi482  & n1212;
  assign n2002 = pi354  & ~n1212;
  assign n2003 = ~n2001 & ~n2002;
  assign n2004 = pi226  & n1789;
  assign n2005 = pi98  & ~n1789;
  assign n2006 = ~n2004 & ~n2005;
  assign n2007 = ~n2003 & n2006;
  assign n2008 = ~n2000 & ~n2007;
  assign n2009 = pi478  & n1212;
  assign n2010 = pi350  & ~n1212;
  assign n2011 = ~n2009 & ~n2010;
  assign n2012 = pi223  & n1789;
  assign n2013 = pi95  & ~n1789;
  assign n2014 = ~n2012 & ~n2013;
  assign n2015 = pi479  & n1212;
  assign n2016 = pi351  & ~n1212;
  assign n2017 = ~n2015 & ~n2016;
  assign n2018 = n2014 & ~n2017;
  assign n2019 = pi222  & n1789;
  assign n2020 = pi94  & ~n1789;
  assign n2021 = ~n2019 & ~n2020;
  assign n2022 = ~n2018 & ~n2021;
  assign n2023 = n2011 & n2022;
  assign n2024 = n2011 & ~n2018;
  assign n2025 = ~n2022 & ~n2024;
  assign n2026 = pi221  & n1789;
  assign n2027 = pi93  & ~n1789;
  assign n2028 = ~n2026 & ~n2027;
  assign n2029 = pi477  & n1212;
  assign n2030 = pi349  & ~n1212;
  assign n2031 = ~n2029 & ~n2030;
  assign n2032 = ~n2028 & n2031;
  assign n2033 = pi220  & n1789;
  assign n2034 = pi92  & ~n1789;
  assign n2035 = ~n2033 & ~n2034;
  assign n2036 = n2028 & ~n2031;
  assign n2037 = pi476  & n1212;
  assign n2038 = pi348  & ~n1212;
  assign n2039 = ~n2037 & ~n2038;
  assign n2040 = ~n2036 & n2039;
  assign n2041 = ~n2035 & n2040;
  assign n2042 = ~n2032 & ~n2041;
  assign n2043 = ~n2025 & ~n2042;
  assign n2044 = ~n2014 & n2017;
  assign n2045 = pi217  & n1789;
  assign n2046 = pi89  & ~n1789;
  assign n2047 = ~n2045 & ~n2046;
  assign n2048 = pi473  & n1212;
  assign n2049 = pi345  & ~n1212;
  assign n2050 = ~n2048 & ~n2049;
  assign n2051 = n2047 & ~n2050;
  assign n2052 = pi219  & n1789;
  assign n2053 = pi91  & ~n1789;
  assign n2054 = ~n2052 & ~n2053;
  assign n2055 = pi475  & n1212;
  assign n2056 = pi347  & ~n1212;
  assign n2057 = ~n2055 & ~n2056;
  assign n2058 = n2054 & ~n2057;
  assign n2059 = pi474  & n1212;
  assign n2060 = pi346  & ~n1212;
  assign n2061 = ~n2059 & ~n2060;
  assign n2062 = pi218  & n1789;
  assign n2063 = pi90  & ~n1789;
  assign n2064 = ~n2062 & ~n2063;
  assign n2065 = ~n2061 & n2064;
  assign n2066 = ~n2058 & ~n2065;
  assign n2067 = pi470  & n1212;
  assign n2068 = pi342  & ~n1212;
  assign n2069 = ~n2067 & ~n2068;
  assign n2070 = pi215  & n1789;
  assign n2071 = pi87  & ~n1789;
  assign n2072 = ~n2070 & ~n2071;
  assign n2073 = pi471  & n1212;
  assign n2074 = pi343  & ~n1212;
  assign n2075 = ~n2073 & ~n2074;
  assign n2076 = n2072 & ~n2075;
  assign n2077 = pi214  & n1789;
  assign n2078 = pi86  & ~n1789;
  assign n2079 = ~n2077 & ~n2078;
  assign n2080 = ~n2076 & ~n2079;
  assign n2081 = n2069 & n2080;
  assign n2082 = n2069 & ~n2076;
  assign n2083 = ~n2080 & ~n2082;
  assign n2084 = pi213  & n1789;
  assign n2085 = pi85  & ~n1789;
  assign n2086 = ~n2084 & ~n2085;
  assign n2087 = pi469  & n1212;
  assign n2088 = pi341  & ~n1212;
  assign n2089 = ~n2087 & ~n2088;
  assign n2090 = ~n2086 & n2089;
  assign n2091 = pi212  & n1789;
  assign n2092 = pi84  & ~n1789;
  assign n2093 = ~n2091 & ~n2092;
  assign n2094 = n2086 & ~n2089;
  assign n2095 = pi468  & n1212;
  assign n2096 = pi340  & ~n1212;
  assign n2097 = ~n2095 & ~n2096;
  assign n2098 = ~n2094 & n2097;
  assign n2099 = ~n2093 & n2098;
  assign n2100 = ~n2090 & ~n2099;
  assign n2101 = ~n2083 & ~n2100;
  assign n2102 = ~n2072 & n2075;
  assign n2103 = pi209  & n1789;
  assign n2104 = pi81  & ~n1789;
  assign n2105 = ~n2103 & ~n2104;
  assign n2106 = pi465  & n1212;
  assign n2107 = pi337  & ~n1212;
  assign n2108 = ~n2106 & ~n2107;
  assign n2109 = n2105 & ~n2108;
  assign n2110 = pi211  & n1789;
  assign n2111 = pi83  & ~n1789;
  assign n2112 = ~n2110 & ~n2111;
  assign n2113 = pi467  & n1212;
  assign n2114 = pi339  & ~n1212;
  assign n2115 = ~n2113 & ~n2114;
  assign n2116 = n2112 & ~n2115;
  assign n2117 = pi466  & n1212;
  assign n2118 = pi338  & ~n1212;
  assign n2119 = ~n2117 & ~n2118;
  assign n2120 = pi210  & n1789;
  assign n2121 = pi82  & ~n1789;
  assign n2122 = ~n2120 & ~n2121;
  assign n2123 = ~n2119 & n2122;
  assign n2124 = ~n2116 & ~n2123;
  assign n2125 = pi462  & n1212;
  assign n2126 = pi334  & ~n1212;
  assign n2127 = ~n2125 & ~n2126;
  assign n2128 = pi207  & n1789;
  assign n2129 = pi79  & ~n1789;
  assign n2130 = ~n2128 & ~n2129;
  assign n2131 = pi463  & n1212;
  assign n2132 = pi335  & ~n1212;
  assign n2133 = ~n2131 & ~n2132;
  assign n2134 = n2130 & ~n2133;
  assign n2135 = pi206  & n1789;
  assign n2136 = pi78  & ~n1789;
  assign n2137 = ~n2135 & ~n2136;
  assign n2138 = ~n2134 & ~n2137;
  assign n2139 = n2127 & n2138;
  assign n2140 = n2127 & ~n2134;
  assign n2141 = ~n2138 & ~n2140;
  assign n2142 = pi205  & n1789;
  assign n2143 = pi77  & ~n1789;
  assign n2144 = ~n2142 & ~n2143;
  assign n2145 = pi461  & n1212;
  assign n2146 = pi333  & ~n1212;
  assign n2147 = ~n2145 & ~n2146;
  assign n2148 = ~n2144 & n2147;
  assign n2149 = pi204  & n1789;
  assign n2150 = pi76  & ~n1789;
  assign n2151 = ~n2149 & ~n2150;
  assign n2152 = n2144 & ~n2147;
  assign n2153 = pi460  & n1212;
  assign n2154 = pi332  & ~n1212;
  assign n2155 = ~n2153 & ~n2154;
  assign n2156 = ~n2152 & n2155;
  assign n2157 = ~n2151 & n2156;
  assign n2158 = ~n2148 & ~n2157;
  assign n2159 = ~n2141 & ~n2158;
  assign n2160 = ~n2130 & n2133;
  assign n2161 = pi201  & n1789;
  assign n2162 = pi73  & ~n1789;
  assign n2163 = ~n2161 & ~n2162;
  assign n2164 = pi457  & n1212;
  assign n2165 = pi329  & ~n1212;
  assign n2166 = ~n2164 & ~n2165;
  assign n2167 = n2163 & ~n2166;
  assign n2168 = pi203  & n1789;
  assign n2169 = pi75  & ~n1789;
  assign n2170 = ~n2168 & ~n2169;
  assign n2171 = pi459  & n1212;
  assign n2172 = pi331  & ~n1212;
  assign n2173 = ~n2171 & ~n2172;
  assign n2174 = n2170 & ~n2173;
  assign n2175 = pi458  & n1212;
  assign n2176 = pi330  & ~n1212;
  assign n2177 = ~n2175 & ~n2176;
  assign n2178 = pi202  & n1789;
  assign n2179 = pi74  & ~n1789;
  assign n2180 = ~n2178 & ~n2179;
  assign n2181 = ~n2177 & n2180;
  assign n2182 = ~n2174 & ~n2181;
  assign n2183 = pi454  & n1212;
  assign n2184 = pi326  & ~n1212;
  assign n2185 = ~n2183 & ~n2184;
  assign n2186 = pi199  & n1789;
  assign n2187 = pi71  & ~n1789;
  assign n2188 = ~n2186 & ~n2187;
  assign n2189 = pi455  & n1212;
  assign n2190 = pi327  & ~n1212;
  assign n2191 = ~n2189 & ~n2190;
  assign n2192 = n2188 & ~n2191;
  assign n2193 = pi198  & n1789;
  assign n2194 = pi70  & ~n1789;
  assign n2195 = ~n2193 & ~n2194;
  assign n2196 = ~n2192 & ~n2195;
  assign n2197 = n2185 & n2196;
  assign n2198 = n2185 & ~n2192;
  assign n2199 = ~n2196 & ~n2198;
  assign n2200 = pi197  & n1789;
  assign n2201 = pi69  & ~n1789;
  assign n2202 = ~n2200 & ~n2201;
  assign n2203 = pi453  & n1212;
  assign n2204 = pi325  & ~n1212;
  assign n2205 = ~n2203 & ~n2204;
  assign n2206 = ~n2202 & n2205;
  assign n2207 = pi196  & n1789;
  assign n2208 = pi68  & ~n1789;
  assign n2209 = ~n2207 & ~n2208;
  assign n2210 = n2202 & ~n2205;
  assign n2211 = pi452  & n1212;
  assign n2212 = pi324  & ~n1212;
  assign n2213 = ~n2211 & ~n2212;
  assign n2214 = ~n2210 & n2213;
  assign n2215 = ~n2209 & n2214;
  assign n2216 = ~n2206 & ~n2215;
  assign n2217 = ~n2199 & ~n2216;
  assign n2218 = ~n2188 & n2191;
  assign n2219 = pi193  & n1789;
  assign n2220 = pi65  & ~n1789;
  assign n2221 = ~n2219 & ~n2220;
  assign n2222 = pi449  & n1212;
  assign n2223 = pi321  & ~n1212;
  assign n2224 = ~n2222 & ~n2223;
  assign n2225 = n2221 & ~n2224;
  assign n2226 = pi195  & n1789;
  assign n2227 = pi67  & ~n1789;
  assign n2228 = ~n2226 & ~n2227;
  assign n2229 = pi451  & n1212;
  assign n2230 = pi323  & ~n1212;
  assign n2231 = ~n2229 & ~n2230;
  assign n2232 = n2228 & ~n2231;
  assign n2233 = pi450  & n1212;
  assign n2234 = pi322  & ~n1212;
  assign n2235 = ~n2233 & ~n2234;
  assign n2236 = pi194  & n1789;
  assign n2237 = pi66  & ~n1789;
  assign n2238 = ~n2236 & ~n2237;
  assign n2239 = ~n2235 & n2238;
  assign n2240 = ~n2232 & ~n2239;
  assign n2241 = pi187  & n1789;
  assign n2242 = pi59  & ~n1789;
  assign n2243 = ~n2241 & ~n2242;
  assign n2244 = pi443  & n1212;
  assign n2245 = pi315  & ~n1212;
  assign n2246 = ~n2244 & ~n2245;
  assign n2247 = ~n2243 & n2246;
  assign n2248 = n2243 & ~n2246;
  assign n2249 = pi186  & n1789;
  assign n2250 = pi58  & ~n1789;
  assign n2251 = ~n2249 & ~n2250;
  assign n2252 = pi442  & n1212;
  assign n2253 = pi314  & ~n1212;
  assign n2254 = ~n2252 & ~n2253;
  assign n2255 = n2251 & ~n2254;
  assign n2256 = ~n2248 & ~n2255;
  assign n2257 = ~n2251 & n2254;
  assign n2258 = pi185  & n1789;
  assign n2259 = pi57  & ~n1789;
  assign n2260 = ~n2258 & ~n2259;
  assign n2261 = pi441  & n1212;
  assign n2262 = pi313  & ~n1212;
  assign n2263 = ~n2261 & ~n2262;
  assign n2264 = ~n2260 & n2263;
  assign n2265 = pi184  & n1789;
  assign n2266 = pi56  & ~n1789;
  assign n2267 = ~n2265 & ~n2266;
  assign n2268 = n2260 & ~n2263;
  assign n2269 = pi440  & n1212;
  assign n2270 = pi312  & ~n1212;
  assign n2271 = ~n2269 & ~n2270;
  assign n2272 = ~n2268 & n2271;
  assign n2273 = ~n2267 & n2272;
  assign n2274 = ~n2264 & ~n2273;
  assign n2275 = ~n2257 & n2274;
  assign n2276 = n2256 & ~n2275;
  assign n2277 = ~n2247 & ~n2276;
  assign n2278 = pi191  & n1789;
  assign n2279 = pi63  & ~n1789;
  assign n2280 = ~n2278 & ~n2279;
  assign n2281 = pi447  & n1212;
  assign n2282 = pi319  & ~n1212;
  assign n2283 = ~n2281 & ~n2282;
  assign n2284 = n2280 & ~n2283;
  assign n2285 = pi190  & n1789;
  assign n2286 = pi62  & ~n1789;
  assign n2287 = ~n2285 & ~n2286;
  assign n2288 = ~n2284 & ~n2287;
  assign n2289 = pi446  & n1212;
  assign n2290 = pi318  & ~n1212;
  assign n2291 = ~n2289 & ~n2290;
  assign n2292 = ~n2284 & n2291;
  assign n2293 = ~n2288 & ~n2292;
  assign n2294 = pi189  & n1789;
  assign n2295 = pi61  & ~n1789;
  assign n2296 = ~n2294 & ~n2295;
  assign n2297 = pi445  & n1212;
  assign n2298 = pi317  & ~n1212;
  assign n2299 = ~n2297 & ~n2298;
  assign n2300 = n2296 & ~n2299;
  assign n2301 = pi188  & n1789;
  assign n2302 = pi60  & ~n1789;
  assign n2303 = ~n2301 & ~n2302;
  assign n2304 = pi444  & n1212;
  assign n2305 = pi316  & ~n1212;
  assign n2306 = ~n2304 & ~n2305;
  assign n2307 = n2303 & ~n2306;
  assign n2308 = ~n2300 & ~n2307;
  assign n2309 = ~n2293 & n2308;
  assign n2310 = ~n2277 & n2309;
  assign n2311 = ~n2296 & n2299;
  assign n2312 = ~n2303 & n2306;
  assign n2313 = ~n2311 & ~n2312;
  assign n2314 = ~n2300 & ~n2313;
  assign n2315 = ~n2293 & n2314;
  assign n2316 = ~n2280 & n2283;
  assign n2317 = n2267 & ~n2271;
  assign n2318 = n2309 & ~n2317;
  assign n2319 = pi183  & n1789;
  assign n2320 = pi55  & ~n1789;
  assign n2321 = ~n2319 & ~n2320;
  assign n2322 = pi439  & n1212;
  assign n2323 = pi311  & ~n1212;
  assign n2324 = ~n2322 & ~n2323;
  assign n2325 = ~n2321 & n2324;
  assign n2326 = pi432  & n1212;
  assign n2327 = pi304  & ~n1212;
  assign n2328 = ~n2326 & ~n2327;
  assign n2329 = pi176  & n1789;
  assign n2330 = pi48  & ~n1789;
  assign n2331 = ~n2329 & ~n2330;
  assign n2332 = ~n2328 & n2331;
  assign n2333 = pi171  & n1789;
  assign n2334 = pi43  & ~n1789;
  assign n2335 = ~n2333 & ~n2334;
  assign n2336 = pi427  & n1212;
  assign n2337 = pi299  & ~n1212;
  assign n2338 = ~n2336 & ~n2337;
  assign n2339 = ~n2335 & n2338;
  assign n2340 = n2335 & ~n2338;
  assign n2341 = pi170  & n1789;
  assign n2342 = pi42  & ~n1789;
  assign n2343 = ~n2341 & ~n2342;
  assign n2344 = pi426  & n1212;
  assign n2345 = pi298  & ~n1212;
  assign n2346 = ~n2344 & ~n2345;
  assign n2347 = n2343 & ~n2346;
  assign n2348 = ~n2340 & ~n2347;
  assign n2349 = ~n2343 & n2346;
  assign n2350 = pi169  & n1789;
  assign n2351 = pi41  & ~n1789;
  assign n2352 = ~n2350 & ~n2351;
  assign n2353 = pi425  & n1212;
  assign n2354 = pi297  & ~n1212;
  assign n2355 = ~n2353 & ~n2354;
  assign n2356 = ~n2352 & n2355;
  assign n2357 = pi168  & n1789;
  assign n2358 = pi40  & ~n1789;
  assign n2359 = ~n2357 & ~n2358;
  assign n2360 = n2352 & ~n2355;
  assign n2361 = pi424  & n1212;
  assign n2362 = pi296  & ~n1212;
  assign n2363 = ~n2361 & ~n2362;
  assign n2364 = ~n2360 & n2363;
  assign n2365 = ~n2359 & n2364;
  assign n2366 = ~n2356 & ~n2365;
  assign n2367 = ~n2349 & n2366;
  assign n2368 = n2348 & ~n2367;
  assign n2369 = ~n2339 & ~n2368;
  assign n2370 = pi175  & n1789;
  assign n2371 = pi47  & ~n1789;
  assign n2372 = ~n2370 & ~n2371;
  assign n2373 = pi431  & n1212;
  assign n2374 = pi303  & ~n1212;
  assign n2375 = ~n2373 & ~n2374;
  assign n2376 = n2372 & ~n2375;
  assign n2377 = pi174  & n1789;
  assign n2378 = pi46  & ~n1789;
  assign n2379 = ~n2377 & ~n2378;
  assign n2380 = ~n2376 & ~n2379;
  assign n2381 = pi430  & n1212;
  assign n2382 = pi302  & ~n1212;
  assign n2383 = ~n2381 & ~n2382;
  assign n2384 = ~n2376 & n2383;
  assign n2385 = ~n2380 & ~n2384;
  assign n2386 = pi173  & n1789;
  assign n2387 = pi45  & ~n1789;
  assign n2388 = ~n2386 & ~n2387;
  assign n2389 = pi429  & n1212;
  assign n2390 = pi301  & ~n1212;
  assign n2391 = ~n2389 & ~n2390;
  assign n2392 = n2388 & ~n2391;
  assign n2393 = pi172  & n1789;
  assign n2394 = pi44  & ~n1789;
  assign n2395 = ~n2393 & ~n2394;
  assign n2396 = pi428  & n1212;
  assign n2397 = pi300  & ~n1212;
  assign n2398 = ~n2396 & ~n2397;
  assign n2399 = n2395 & ~n2398;
  assign n2400 = ~n2392 & ~n2399;
  assign n2401 = ~n2385 & n2400;
  assign n2402 = ~n2369 & n2401;
  assign n2403 = ~n2388 & n2391;
  assign n2404 = ~n2395 & n2398;
  assign n2405 = ~n2403 & ~n2404;
  assign n2406 = ~n2392 & ~n2405;
  assign n2407 = ~n2385 & n2406;
  assign n2408 = ~n2372 & n2375;
  assign n2409 = n2359 & ~n2363;
  assign n2410 = n2401 & ~n2409;
  assign n2411 = pi416  & n1212;
  assign n2412 = pi288  & ~n1212;
  assign n2413 = ~n2411 & ~n2412;
  assign n2414 = pi160  & n1789;
  assign n2415 = pi32  & ~n1789;
  assign n2416 = ~n2414 & ~n2415;
  assign n2417 = ~n2413 & n2416;
  assign n2418 = pi164  & n1789;
  assign n2419 = pi36  & ~n1789;
  assign n2420 = ~n2418 & ~n2419;
  assign n2421 = pi420  & n1212;
  assign n2422 = pi292  & ~n1212;
  assign n2423 = ~n2421 & ~n2422;
  assign n2424 = n2420 & ~n2423;
  assign n2425 = pi166  & n1789;
  assign n2426 = pi38  & ~n1789;
  assign n2427 = ~n2425 & ~n2426;
  assign n2428 = pi422  & n1212;
  assign n2429 = pi294  & ~n1212;
  assign n2430 = ~n2428 & ~n2429;
  assign n2431 = n2427 & ~n2430;
  assign n2432 = pi167  & n1789;
  assign n2433 = pi39  & ~n1789;
  assign n2434 = ~n2432 & ~n2433;
  assign n2435 = pi423  & n1212;
  assign n2436 = pi295  & ~n1212;
  assign n2437 = ~n2435 & ~n2436;
  assign n2438 = n2434 & ~n2437;
  assign n2439 = pi165  & n1789;
  assign n2440 = pi37  & ~n1789;
  assign n2441 = ~n2439 & ~n2440;
  assign n2442 = pi421  & n1212;
  assign n2443 = pi293  & ~n1212;
  assign n2444 = ~n2442 & ~n2443;
  assign n2445 = n2441 & ~n2444;
  assign n2446 = ~n2438 & ~n2445;
  assign n2447 = ~n2431 & n2446;
  assign n2448 = ~n2424 & n2447;
  assign n2449 = ~n2417 & n2448;
  assign n2450 = pi159  & n1789;
  assign n2451 = pi31  & ~n1789;
  assign n2452 = ~n2450 & ~n2451;
  assign n2453 = pi415  & n1212;
  assign n2454 = pi287  & ~n1212;
  assign n2455 = ~n2453 & ~n2454;
  assign n2456 = n2452 & ~n2455;
  assign n2457 = pi163  & n1789;
  assign n2458 = pi35  & ~n1789;
  assign n2459 = ~n2457 & ~n2458;
  assign n2460 = pi419  & n1212;
  assign n2461 = pi291  & ~n1212;
  assign n2462 = ~n2460 & ~n2461;
  assign n2463 = n2459 & ~n2462;
  assign n2464 = pi161  & n1789;
  assign n2465 = pi33  & ~n1789;
  assign n2466 = ~n2464 & ~n2465;
  assign n2467 = pi417  & n1212;
  assign n2468 = pi289  & ~n1212;
  assign n2469 = ~n2467 & ~n2468;
  assign n2470 = n2466 & ~n2469;
  assign n2471 = pi418  & n1212;
  assign n2472 = pi290  & ~n1212;
  assign n2473 = ~n2471 & ~n2472;
  assign n2474 = pi162  & n1789;
  assign n2475 = pi34  & ~n1789;
  assign n2476 = ~n2474 & ~n2475;
  assign n2477 = ~n2473 & n2476;
  assign n2478 = ~n2470 & ~n2477;
  assign n2479 = ~n2463 & n2478;
  assign n2480 = pi158  & n1789;
  assign n2481 = pi30  & ~n1789;
  assign n2482 = ~n2480 & ~n2481;
  assign n2483 = pi414  & n1212;
  assign n2484 = pi286  & ~n1212;
  assign n2485 = ~n2483 & ~n2484;
  assign n2486 = ~n2482 & n2485;
  assign n2487 = ~n2452 & n2455;
  assign n2488 = n2482 & ~n2485;
  assign n2489 = pi157  & n1789;
  assign n2490 = pi29  & ~n1789;
  assign n2491 = ~n2489 & ~n2490;
  assign n2492 = pi413  & n1212;
  assign n2493 = pi285  & ~n1212;
  assign n2494 = ~n2492 & ~n2493;
  assign n2495 = ~n2491 & n2494;
  assign n2496 = n2491 & ~n2494;
  assign n2497 = pi156  & n1789;
  assign n2498 = pi28  & ~n1789;
  assign n2499 = ~n2497 & ~n2498;
  assign n2500 = pi412  & n1212;
  assign n2501 = pi284  & ~n1212;
  assign n2502 = ~n2500 & ~n2501;
  assign n2503 = ~n2499 & n2502;
  assign n2504 = n2499 & ~n2502;
  assign n2505 = pi155  & n1789;
  assign n2506 = pi27  & ~n1789;
  assign n2507 = ~n2505 & ~n2506;
  assign n2508 = pi411  & n1212;
  assign n2509 = pi283  & ~n1212;
  assign n2510 = ~n2508 & ~n2509;
  assign n2511 = ~n2507 & n2510;
  assign n2512 = n2507 & ~n2510;
  assign n2513 = pi154  & n1789;
  assign n2514 = pi26  & ~n1789;
  assign n2515 = ~n2513 & ~n2514;
  assign n2516 = pi410  & n1212;
  assign n2517 = pi282  & ~n1212;
  assign n2518 = ~n2516 & ~n2517;
  assign n2519 = ~n2515 & n2518;
  assign n2520 = n2515 & ~n2518;
  assign n2521 = pi409  & n1212;
  assign n2522 = pi281  & ~n1212;
  assign n2523 = ~n2521 & ~n2522;
  assign n2524 = pi153  & n1789;
  assign n2525 = pi25  & ~n1789;
  assign n2526 = ~n2524 & ~n2525;
  assign n2527 = pi151  & n1789;
  assign n2528 = pi23  & ~n1789;
  assign n2529 = ~n2527 & ~n2528;
  assign n2530 = pi407  & n1212;
  assign n2531 = pi279  & ~n1212;
  assign n2532 = ~n2530 & ~n2531;
  assign n2533 = ~n2529 & n2532;
  assign n2534 = n2529 & ~n2532;
  assign n2535 = pi150  & n1789;
  assign n2536 = pi22  & ~n1789;
  assign n2537 = ~n2535 & ~n2536;
  assign n2538 = pi406  & n1212;
  assign n2539 = pi278  & ~n1212;
  assign n2540 = ~n2538 & ~n2539;
  assign n2541 = ~n2537 & n2540;
  assign n2542 = n2537 & ~n2540;
  assign n2543 = pi149  & n1789;
  assign n2544 = pi21  & ~n1789;
  assign n2545 = ~n2543 & ~n2544;
  assign n2546 = pi405  & n1212;
  assign n2547 = pi277  & ~n1212;
  assign n2548 = ~n2546 & ~n2547;
  assign n2549 = ~n2545 & n2548;
  assign n2550 = n2545 & ~n2548;
  assign n2551 = pi148  & n1789;
  assign n2552 = pi20  & ~n1789;
  assign n2553 = ~n2551 & ~n2552;
  assign n2554 = pi404  & n1212;
  assign n2555 = pi276  & ~n1212;
  assign n2556 = ~n2554 & ~n2555;
  assign n2557 = ~n2553 & n2556;
  assign n2558 = n2553 & ~n2556;
  assign n2559 = pi147  & n1789;
  assign n2560 = pi19  & ~n1789;
  assign n2561 = ~n2559 & ~n2560;
  assign n2562 = pi403  & n1212;
  assign n2563 = pi275  & ~n1212;
  assign n2564 = ~n2562 & ~n2563;
  assign n2565 = ~n2561 & n2564;
  assign n2566 = n2561 & ~n2564;
  assign n2567 = pi146  & n1789;
  assign n2568 = pi18  & ~n1789;
  assign n2569 = ~n2567 & ~n2568;
  assign n2570 = pi402  & n1212;
  assign n2571 = pi274  & ~n1212;
  assign n2572 = ~n2570 & ~n2571;
  assign n2573 = ~n2569 & n2572;
  assign n2574 = n2569 & ~n2572;
  assign n2575 = pi401  & n1212;
  assign n2576 = pi273  & ~n1212;
  assign n2577 = ~n2575 & ~n2576;
  assign n2578 = pi145  & n1789;
  assign n2579 = pi17  & ~n1789;
  assign n2580 = ~n2578 & ~n2579;
  assign n2581 = pi143  & n1789;
  assign n2582 = pi15  & ~n1789;
  assign n2583 = ~n2581 & ~n2582;
  assign n2584 = pi399  & n1212;
  assign n2585 = pi271  & ~n1212;
  assign n2586 = ~n2584 & ~n2585;
  assign n2587 = ~n2583 & n2586;
  assign n2588 = n2583 & ~n2586;
  assign n2589 = pi142  & n1789;
  assign n2590 = pi14  & ~n1789;
  assign n2591 = ~n2589 & ~n2590;
  assign n2592 = pi398  & n1212;
  assign n2593 = pi270  & ~n1212;
  assign n2594 = ~n2592 & ~n2593;
  assign n2595 = ~n2591 & n2594;
  assign n2596 = n2591 & ~n2594;
  assign n2597 = pi141  & n1789;
  assign n2598 = pi13  & ~n1789;
  assign n2599 = ~n2597 & ~n2598;
  assign n2600 = pi397  & n1212;
  assign n2601 = pi269  & ~n1212;
  assign n2602 = ~n2600 & ~n2601;
  assign n2603 = ~n2599 & n2602;
  assign n2604 = n2599 & ~n2602;
  assign n2605 = pi140  & n1789;
  assign n2606 = pi12  & ~n1789;
  assign n2607 = ~n2605 & ~n2606;
  assign n2608 = pi396  & n1212;
  assign n2609 = pi268  & ~n1212;
  assign n2610 = ~n2608 & ~n2609;
  assign n2611 = ~n2607 & n2610;
  assign n2612 = n2607 & ~n2610;
  assign n2613 = pi139  & n1789;
  assign n2614 = pi11  & ~n1789;
  assign n2615 = ~n2613 & ~n2614;
  assign n2616 = pi395  & n1212;
  assign n2617 = pi267  & ~n1212;
  assign n2618 = ~n2616 & ~n2617;
  assign n2619 = ~n2615 & n2618;
  assign n2620 = n2615 & ~n2618;
  assign n2621 = pi138  & n1789;
  assign n2622 = pi10  & ~n1789;
  assign n2623 = ~n2621 & ~n2622;
  assign n2624 = pi394  & n1212;
  assign n2625 = pi266  & ~n1212;
  assign n2626 = ~n2624 & ~n2625;
  assign n2627 = ~n2623 & n2626;
  assign n2628 = n2623 & ~n2626;
  assign n2629 = pi393  & n1212;
  assign n2630 = pi265  & ~n1212;
  assign n2631 = ~n2629 & ~n2630;
  assign n2632 = pi137  & n1789;
  assign n2633 = pi9  & ~n1789;
  assign n2634 = ~n2632 & ~n2633;
  assign n2635 = pi135  & n1789;
  assign n2636 = pi7  & ~n1789;
  assign n2637 = ~n2635 & ~n2636;
  assign n2638 = pi391  & n1212;
  assign n2639 = pi263  & ~n1212;
  assign n2640 = ~n2638 & ~n2639;
  assign n2641 = ~n2637 & n2640;
  assign n2642 = n2637 & ~n2640;
  assign n2643 = pi390  & n1212;
  assign n2644 = pi262  & ~n1212;
  assign n2645 = ~n2643 & ~n2644;
  assign n2646 = pi134  & n1789;
  assign n2647 = pi6  & ~n1789;
  assign n2648 = ~n2646 & ~n2647;
  assign n2649 = pi133  & n1789;
  assign n2650 = pi5  & ~n1789;
  assign n2651 = ~n2649 & ~n2650;
  assign n2652 = pi389  & n1212;
  assign n2653 = pi261  & ~n1212;
  assign n2654 = ~n2652 & ~n2653;
  assign n2655 = pi131  & n1789;
  assign n2656 = pi3  & ~n1789;
  assign n2657 = ~n2655 & ~n2656;
  assign n2658 = pi387  & n1212;
  assign n2659 = pi259  & ~n1212;
  assign n2660 = ~n2658 & ~n2659;
  assign n2661 = ~n2657 & n2660;
  assign n2662 = n2657 & ~n2660;
  assign n2663 = pi130  & n1789;
  assign n2664 = pi2  & ~n1789;
  assign n2665 = ~n2663 & ~n2664;
  assign n2666 = pi386  & n1212;
  assign n2667 = pi258  & ~n1212;
  assign n2668 = ~n2666 & ~n2667;
  assign n2669 = ~n2665 & n2668;
  assign n2670 = n2665 & ~n2668;
  assign n2671 = pi385  & n1212;
  assign n2672 = pi257  & ~n1212;
  assign n2673 = ~n2671 & ~n2672;
  assign n2674 = pi128  & n1789;
  assign n2675 = pi0  & ~n1789;
  assign n2676 = ~n2674 & ~n2675;
  assign n2677 = n1215 & ~n2676;
  assign n2678 = n2673 & n2677;
  assign n2679 = pi129  & n1789;
  assign n2680 = pi1  & ~n1789;
  assign n2681 = ~n2679 & ~n2680;
  assign n2682 = ~n2673 & ~n2677;
  assign n2683 = ~n2681 & ~n2682;
  assign n2684 = ~n2678 & ~n2683;
  assign n2685 = ~n2670 & ~n2684;
  assign n2686 = ~n2669 & ~n2685;
  assign n2687 = ~n2662 & ~n2686;
  assign n2688 = ~n2661 & ~n2687;
  assign n2689 = pi132  & n1789;
  assign n2690 = pi4  & ~n1789;
  assign n2691 = ~n2689 & ~n2690;
  assign n2692 = pi388  & n1212;
  assign n2693 = pi260  & ~n1212;
  assign n2694 = ~n2692 & ~n2693;
  assign n2695 = ~n2691 & n2694;
  assign n2696 = n2688 & ~n2695;
  assign n2697 = n2691 & ~n2694;
  assign n2698 = ~n2696 & ~n2697;
  assign n2699 = n2654 & n2698;
  assign n2700 = n2651 & ~n2699;
  assign n2701 = ~n2654 & ~n2698;
  assign n2702 = ~n2700 & ~n2701;
  assign n2703 = n2648 & ~n2702;
  assign n2704 = n2645 & ~n2703;
  assign n2705 = ~n2648 & n2702;
  assign n2706 = ~n2704 & ~n2705;
  assign n2707 = ~n2642 & ~n2706;
  assign n2708 = ~n2641 & ~n2707;
  assign n2709 = pi136  & n1789;
  assign n2710 = pi8  & ~n1789;
  assign n2711 = ~n2709 & ~n2710;
  assign n2712 = pi392  & n1212;
  assign n2713 = pi264  & ~n1212;
  assign n2714 = ~n2712 & ~n2713;
  assign n2715 = ~n2711 & n2714;
  assign n2716 = n2708 & ~n2715;
  assign n2717 = n2711 & ~n2714;
  assign n2718 = ~n2716 & ~n2717;
  assign n2719 = n2634 & ~n2718;
  assign n2720 = n2631 & ~n2719;
  assign n2721 = ~n2634 & n2718;
  assign n2722 = ~n2720 & ~n2721;
  assign n2723 = ~n2628 & ~n2722;
  assign n2724 = ~n2627 & ~n2723;
  assign n2725 = ~n2620 & ~n2724;
  assign n2726 = ~n2619 & ~n2725;
  assign n2727 = ~n2612 & ~n2726;
  assign n2728 = ~n2611 & ~n2727;
  assign n2729 = ~n2604 & ~n2728;
  assign n2730 = ~n2603 & ~n2729;
  assign n2731 = ~n2596 & ~n2730;
  assign n2732 = ~n2595 & ~n2731;
  assign n2733 = ~n2588 & ~n2732;
  assign n2734 = ~n2587 & ~n2733;
  assign n2735 = pi144  & n1789;
  assign n2736 = pi16  & ~n1789;
  assign n2737 = ~n2735 & ~n2736;
  assign n2738 = pi400  & n1212;
  assign n2739 = pi272  & ~n1212;
  assign n2740 = ~n2738 & ~n2739;
  assign n2741 = ~n2737 & n2740;
  assign n2742 = n2734 & ~n2741;
  assign n2743 = n2737 & ~n2740;
  assign n2744 = ~n2742 & ~n2743;
  assign n2745 = n2580 & ~n2744;
  assign n2746 = n2577 & ~n2745;
  assign n2747 = ~n2580 & n2744;
  assign n2748 = ~n2746 & ~n2747;
  assign n2749 = ~n2574 & ~n2748;
  assign n2750 = ~n2573 & ~n2749;
  assign n2751 = ~n2566 & ~n2750;
  assign n2752 = ~n2565 & ~n2751;
  assign n2753 = ~n2558 & ~n2752;
  assign n2754 = ~n2557 & ~n2753;
  assign n2755 = ~n2550 & ~n2754;
  assign n2756 = ~n2549 & ~n2755;
  assign n2757 = ~n2542 & ~n2756;
  assign n2758 = ~n2541 & ~n2757;
  assign n2759 = ~n2534 & ~n2758;
  assign n2760 = ~n2533 & ~n2759;
  assign n2761 = pi152  & n1789;
  assign n2762 = pi24  & ~n1789;
  assign n2763 = ~n2761 & ~n2762;
  assign n2764 = pi408  & n1212;
  assign n2765 = pi280  & ~n1212;
  assign n2766 = ~n2764 & ~n2765;
  assign n2767 = ~n2763 & n2766;
  assign n2768 = n2760 & ~n2767;
  assign n2769 = n2763 & ~n2766;
  assign n2770 = ~n2768 & ~n2769;
  assign n2771 = n2526 & ~n2770;
  assign n2772 = n2523 & ~n2771;
  assign n2773 = ~n2526 & n2770;
  assign n2774 = ~n2772 & ~n2773;
  assign n2775 = ~n2520 & ~n2774;
  assign n2776 = ~n2519 & ~n2775;
  assign n2777 = ~n2512 & ~n2776;
  assign n2778 = ~n2511 & ~n2777;
  assign n2779 = ~n2504 & ~n2778;
  assign n2780 = ~n2503 & ~n2779;
  assign n2781 = ~n2496 & ~n2780;
  assign n2782 = ~n2495 & ~n2781;
  assign n2783 = ~n2488 & ~n2782;
  assign n2784 = ~n2487 & ~n2783;
  assign n2785 = ~n2486 & n2784;
  assign n2786 = n2479 & ~n2785;
  assign n2787 = ~n2456 & n2786;
  assign n2788 = n2449 & n2787;
  assign n2789 = ~n2441 & n2444;
  assign n2790 = ~n2420 & n2423;
  assign n2791 = ~n2789 & ~n2790;
  assign n2792 = n2447 & ~n2791;
  assign n2793 = ~n2434 & n2437;
  assign n2794 = ~n2459 & n2462;
  assign n2795 = n2413 & ~n2416;
  assign n2796 = ~n2466 & n2469;
  assign n2797 = ~n2795 & ~n2796;
  assign n2798 = n2479 & ~n2797;
  assign n2799 = ~n2794 & ~n2798;
  assign n2800 = ~n2463 & n2473;
  assign n2801 = ~n2476 & n2800;
  assign n2802 = n2799 & ~n2801;
  assign n2803 = n2448 & ~n2802;
  assign n2804 = ~n2793 & ~n2803;
  assign n2805 = ~n2792 & n2804;
  assign n2806 = ~n2788 & n2805;
  assign n2807 = ~n2427 & n2430;
  assign n2808 = ~n2438 & n2807;
  assign n2809 = n2806 & ~n2808;
  assign n2810 = n2348 & ~n2809;
  assign n2811 = ~n2360 & n2810;
  assign n2812 = n2410 & n2811;
  assign n2813 = n2380 & n2383;
  assign n2814 = ~n2812 & ~n2813;
  assign n2815 = ~n2408 & n2814;
  assign n2816 = ~n2407 & n2815;
  assign n2817 = ~n2402 & n2816;
  assign n2818 = pi181  & n1789;
  assign n2819 = pi53  & ~n1789;
  assign n2820 = ~n2818 & ~n2819;
  assign n2821 = pi437  & n1212;
  assign n2822 = pi309  & ~n1212;
  assign n2823 = ~n2821 & ~n2822;
  assign n2824 = n2820 & ~n2823;
  assign n2825 = pi436  & n1212;
  assign n2826 = pi308  & ~n1212;
  assign n2827 = ~n2825 & ~n2826;
  assign n2828 = pi180  & n1789;
  assign n2829 = pi52  & ~n1789;
  assign n2830 = ~n2828 & ~n2829;
  assign n2831 = ~n2827 & n2830;
  assign n2832 = n2321 & ~n2324;
  assign n2833 = pi438  & n1212;
  assign n2834 = pi310  & ~n1212;
  assign n2835 = ~n2833 & ~n2834;
  assign n2836 = pi182  & n1789;
  assign n2837 = pi54  & ~n1789;
  assign n2838 = ~n2836 & ~n2837;
  assign n2839 = ~n2835 & n2838;
  assign n2840 = ~n2832 & ~n2839;
  assign n2841 = ~n2831 & n2840;
  assign n2842 = ~n2824 & n2841;
  assign n2843 = ~n2817 & n2842;
  assign n2844 = pi179  & n1789;
  assign n2845 = pi51  & ~n1789;
  assign n2846 = ~n2844 & ~n2845;
  assign n2847 = pi435  & n1212;
  assign n2848 = pi307  & ~n1212;
  assign n2849 = ~n2847 & ~n2848;
  assign n2850 = n2846 & ~n2849;
  assign n2851 = pi177  & n1789;
  assign n2852 = pi49  & ~n1789;
  assign n2853 = ~n2851 & ~n2852;
  assign n2854 = pi433  & n1212;
  assign n2855 = pi305  & ~n1212;
  assign n2856 = ~n2854 & ~n2855;
  assign n2857 = n2853 & ~n2856;
  assign n2858 = pi434  & n1212;
  assign n2859 = pi306  & ~n1212;
  assign n2860 = ~n2858 & ~n2859;
  assign n2861 = pi178  & n1789;
  assign n2862 = pi50  & ~n1789;
  assign n2863 = ~n2861 & ~n2862;
  assign n2864 = ~n2860 & n2863;
  assign n2865 = ~n2857 & ~n2864;
  assign n2866 = ~n2850 & n2865;
  assign n2867 = n2843 & n2866;
  assign n2868 = ~n2332 & n2867;
  assign n2869 = n2835 & ~n2838;
  assign n2870 = ~n2820 & n2823;
  assign n2871 = ~n2824 & ~n2830;
  assign n2872 = n2827 & n2871;
  assign n2873 = ~n2870 & ~n2872;
  assign n2874 = ~n2869 & n2873;
  assign n2875 = n2840 & ~n2874;
  assign n2876 = ~n2846 & n2849;
  assign n2877 = n2328 & ~n2331;
  assign n2878 = ~n2853 & n2856;
  assign n2879 = ~n2877 & ~n2878;
  assign n2880 = n2866 & ~n2879;
  assign n2881 = ~n2876 & ~n2880;
  assign n2882 = ~n2850 & n2860;
  assign n2883 = ~n2863 & n2882;
  assign n2884 = n2881 & ~n2883;
  assign n2885 = n2842 & ~n2884;
  assign n2886 = ~n2875 & ~n2885;
  assign n2887 = ~n2868 & n2886;
  assign n2888 = ~n2325 & n2887;
  assign n2889 = n2256 & ~n2888;
  assign n2890 = ~n2268 & n2889;
  assign n2891 = n2318 & n2890;
  assign n2892 = n2288 & n2291;
  assign n2893 = ~n2891 & ~n2892;
  assign n2894 = ~n2316 & n2893;
  assign n2895 = ~n2315 & n2894;
  assign n2896 = ~n2310 & n2895;
  assign n2897 = n2240 & ~n2896;
  assign n2898 = ~n2225 & n2897;
  assign n2899 = pi448  & n1212;
  assign n2900 = pi320  & ~n1212;
  assign n2901 = ~n2899 & ~n2900;
  assign n2902 = pi192  & n1789;
  assign n2903 = pi64  & ~n1789;
  assign n2904 = ~n2902 & ~n2903;
  assign n2905 = ~n2901 & n2904;
  assign n2906 = n2898 & ~n2905;
  assign n2907 = ~n2228 & n2231;
  assign n2908 = n2235 & ~n2238;
  assign n2909 = ~n2221 & n2224;
  assign n2910 = ~n2225 & ~n2904;
  assign n2911 = n2901 & n2910;
  assign n2912 = ~n2909 & ~n2911;
  assign n2913 = ~n2908 & n2912;
  assign n2914 = n2240 & ~n2913;
  assign n2915 = ~n2907 & ~n2914;
  assign n2916 = ~n2906 & n2915;
  assign n2917 = ~n2210 & ~n2916;
  assign n2918 = n2209 & ~n2213;
  assign n2919 = ~n2199 & ~n2918;
  assign n2920 = n2917 & n2919;
  assign n2921 = ~n2218 & ~n2920;
  assign n2922 = ~n2217 & n2921;
  assign n2923 = ~n2197 & n2922;
  assign n2924 = n2182 & ~n2923;
  assign n2925 = ~n2167 & n2924;
  assign n2926 = pi456  & n1212;
  assign n2927 = pi328  & ~n1212;
  assign n2928 = ~n2926 & ~n2927;
  assign n2929 = pi200  & n1789;
  assign n2930 = pi72  & ~n1789;
  assign n2931 = ~n2929 & ~n2930;
  assign n2932 = ~n2928 & n2931;
  assign n2933 = n2925 & ~n2932;
  assign n2934 = ~n2170 & n2173;
  assign n2935 = n2177 & ~n2180;
  assign n2936 = ~n2163 & n2166;
  assign n2937 = ~n2167 & ~n2931;
  assign n2938 = n2928 & n2937;
  assign n2939 = ~n2936 & ~n2938;
  assign n2940 = ~n2935 & n2939;
  assign n2941 = n2182 & ~n2940;
  assign n2942 = ~n2934 & ~n2941;
  assign n2943 = ~n2933 & n2942;
  assign n2944 = ~n2152 & ~n2943;
  assign n2945 = n2151 & ~n2155;
  assign n2946 = ~n2141 & ~n2945;
  assign n2947 = n2944 & n2946;
  assign n2948 = ~n2160 & ~n2947;
  assign n2949 = ~n2159 & n2948;
  assign n2950 = ~n2139 & n2949;
  assign n2951 = n2124 & ~n2950;
  assign n2952 = ~n2109 & n2951;
  assign n2953 = pi464  & n1212;
  assign n2954 = pi336  & ~n1212;
  assign n2955 = ~n2953 & ~n2954;
  assign n2956 = pi208  & n1789;
  assign n2957 = pi80  & ~n1789;
  assign n2958 = ~n2956 & ~n2957;
  assign n2959 = ~n2955 & n2958;
  assign n2960 = n2952 & ~n2959;
  assign n2961 = ~n2112 & n2115;
  assign n2962 = n2119 & ~n2122;
  assign n2963 = ~n2105 & n2108;
  assign n2964 = ~n2109 & ~n2958;
  assign n2965 = n2955 & n2964;
  assign n2966 = ~n2963 & ~n2965;
  assign n2967 = ~n2962 & n2966;
  assign n2968 = n2124 & ~n2967;
  assign n2969 = ~n2961 & ~n2968;
  assign n2970 = ~n2960 & n2969;
  assign n2971 = ~n2094 & ~n2970;
  assign n2972 = n2093 & ~n2097;
  assign n2973 = ~n2083 & ~n2972;
  assign n2974 = n2971 & n2973;
  assign n2975 = ~n2102 & ~n2974;
  assign n2976 = ~n2101 & n2975;
  assign n2977 = ~n2081 & n2976;
  assign n2978 = n2066 & ~n2977;
  assign n2979 = ~n2051 & n2978;
  assign n2980 = pi472  & n1212;
  assign n2981 = pi344  & ~n1212;
  assign n2982 = ~n2980 & ~n2981;
  assign n2983 = pi216  & n1789;
  assign n2984 = pi88  & ~n1789;
  assign n2985 = ~n2983 & ~n2984;
  assign n2986 = ~n2982 & n2985;
  assign n2987 = n2979 & ~n2986;
  assign n2988 = ~n2054 & n2057;
  assign n2989 = n2061 & ~n2064;
  assign n2990 = ~n2047 & n2050;
  assign n2991 = ~n2051 & ~n2985;
  assign n2992 = n2982 & n2991;
  assign n2993 = ~n2990 & ~n2992;
  assign n2994 = ~n2989 & n2993;
  assign n2995 = n2066 & ~n2994;
  assign n2996 = ~n2988 & ~n2995;
  assign n2997 = ~n2987 & n2996;
  assign n2998 = ~n2036 & ~n2997;
  assign n2999 = n2035 & ~n2039;
  assign n3000 = ~n2025 & ~n2999;
  assign n3001 = n2998 & n3000;
  assign n3002 = ~n2044 & ~n3001;
  assign n3003 = ~n2043 & n3002;
  assign n3004 = ~n2023 & n3003;
  assign n3005 = n2008 & ~n3004;
  assign n3006 = ~n1993 & n3005;
  assign n3007 = pi480  & n1212;
  assign n3008 = pi352  & ~n1212;
  assign n3009 = ~n3007 & ~n3008;
  assign n3010 = pi224  & n1789;
  assign n3011 = pi96  & ~n1789;
  assign n3012 = ~n3010 & ~n3011;
  assign n3013 = ~n3009 & n3012;
  assign n3014 = n3006 & ~n3013;
  assign n3015 = ~n1996 & n1999;
  assign n3016 = n2003 & ~n2006;
  assign n3017 = ~n1989 & n1992;
  assign n3018 = ~n1993 & ~n3012;
  assign n3019 = n3009 & n3018;
  assign n3020 = ~n3017 & ~n3019;
  assign n3021 = ~n3016 & n3020;
  assign n3022 = n2008 & ~n3021;
  assign n3023 = ~n3015 & ~n3022;
  assign n3024 = ~n3014 & n3023;
  assign n3025 = ~n1978 & ~n3024;
  assign n3026 = n1977 & ~n1981;
  assign n3027 = ~n1967 & ~n3026;
  assign n3028 = n3025 & n3027;
  assign n3029 = ~n1986 & ~n3028;
  assign n3030 = ~n1985 & n3029;
  assign n3031 = ~n1965 & n3030;
  assign n3032 = n1950 & ~n3031;
  assign n3033 = ~n1935 & n3032;
  assign n3034 = pi488  & n1212;
  assign n3035 = pi360  & ~n1212;
  assign n3036 = ~n3034 & ~n3035;
  assign n3037 = pi232  & n1789;
  assign n3038 = pi104  & ~n1789;
  assign n3039 = ~n3037 & ~n3038;
  assign n3040 = ~n3036 & n3039;
  assign n3041 = n3033 & ~n3040;
  assign n3042 = ~n1938 & n1941;
  assign n3043 = n1945 & ~n1948;
  assign n3044 = ~n1931 & n1934;
  assign n3045 = ~n1935 & ~n3039;
  assign n3046 = n3036 & n3045;
  assign n3047 = ~n3044 & ~n3046;
  assign n3048 = ~n3043 & n3047;
  assign n3049 = n1950 & ~n3048;
  assign n3050 = ~n3042 & ~n3049;
  assign n3051 = ~n3041 & n3050;
  assign n3052 = ~n1920 & ~n3051;
  assign n3053 = n1919 & ~n1923;
  assign n3054 = ~n1909 & ~n3053;
  assign n3055 = n3052 & n3054;
  assign n3056 = ~n1928 & ~n3055;
  assign n3057 = ~n1927 & n3056;
  assign n3058 = ~n1907 & n3057;
  assign n3059 = n1892 & ~n3058;
  assign n3060 = ~n1877 & n3059;
  assign n3061 = pi496  & n1212;
  assign n3062 = pi368  & ~n1212;
  assign n3063 = ~n3061 & ~n3062;
  assign n3064 = pi240  & n1789;
  assign n3065 = pi112  & ~n1789;
  assign n3066 = ~n3064 & ~n3065;
  assign n3067 = ~n3063 & n3066;
  assign n3068 = n3060 & ~n3067;
  assign n3069 = ~n1880 & n1883;
  assign n3070 = n1887 & ~n1890;
  assign n3071 = ~n1873 & n1876;
  assign n3072 = ~n1877 & ~n3066;
  assign n3073 = n3063 & n3072;
  assign n3074 = ~n3071 & ~n3073;
  assign n3075 = ~n3070 & n3074;
  assign n3076 = n1892 & ~n3075;
  assign n3077 = ~n3069 & ~n3076;
  assign n3078 = ~n3068 & n3077;
  assign n3079 = n1844 & ~n1847;
  assign n3080 = n1866 & ~n3079;
  assign n3081 = ~n3078 & n3080;
  assign n3082 = ~n1870 & ~n3081;
  assign n3083 = ~n1869 & n3082;
  assign n3084 = ~n1867 & n3083;
  assign n3085 = n1834 & ~n3084;
  assign n3086 = pi249  & n1789;
  assign n3087 = pi121  & ~n1789;
  assign n3088 = ~n3086 & ~n3087;
  assign n3089 = pi505  & n1212;
  assign n3090 = pi377  & ~n1212;
  assign n3091 = ~n3089 & ~n3090;
  assign n3092 = n3088 & ~n3091;
  assign n3093 = pi248  & n1789;
  assign n3094 = pi120  & ~n1789;
  assign n3095 = ~n3093 & ~n3094;
  assign n3096 = pi504  & n1212;
  assign n3097 = pi376  & ~n1212;
  assign n3098 = ~n3096 & ~n3097;
  assign n3099 = n3095 & ~n3098;
  assign n3100 = ~n3092 & ~n3099;
  assign n3101 = n3085 & n3100;
  assign n3102 = ~n1822 & n1825;
  assign n3103 = n1829 & ~n1832;
  assign n3104 = ~n3088 & n3091;
  assign n3105 = ~n3092 & n3098;
  assign n3106 = ~n3095 & n3105;
  assign n3107 = ~n3104 & ~n3106;
  assign n3108 = ~n3103 & n3107;
  assign n3109 = n1834 & ~n3108;
  assign n3110 = ~n3102 & ~n3109;
  assign n3111 = ~n3101 & n3110;
  assign n3112 = n1804 & ~n3111;
  assign n3113 = ~n1218 & n3112;
  assign n3114 = ~n1819 & n3113;
  assign n3115 = ~n1818 & ~n3114;
  assign po129  = ~n1817 & n3115;
  assign n3117 = ~n1215 & po129 ;
  assign n3118 = ~n2676 & ~po129 ;
  assign po0  = n3117 | n3118;
  assign n3120 = ~n2673 & po129 ;
  assign n3121 = ~n2681 & ~po129 ;
  assign po1  = n3120 | n3121;
  assign n3123 = ~n2668 & po129 ;
  assign n3124 = ~n2665 & ~po129 ;
  assign po2  = n3123 | n3124;
  assign n3126 = ~n2660 & po129 ;
  assign n3127 = ~n2657 & ~po129 ;
  assign po3  = n3126 | n3127;
  assign n3129 = ~n2694 & po129 ;
  assign n3130 = ~n2691 & ~po129 ;
  assign po4  = n3129 | n3130;
  assign n3132 = ~n2654 & po129 ;
  assign n3133 = ~n2651 & ~po129 ;
  assign po5  = n3132 | n3133;
  assign n3135 = ~n2645 & po129 ;
  assign n3136 = ~n2648 & ~po129 ;
  assign po6  = n3135 | n3136;
  assign n3138 = ~n2640 & po129 ;
  assign n3139 = ~n2637 & ~po129 ;
  assign po7  = n3138 | n3139;
  assign n3141 = ~n2714 & po129 ;
  assign n3142 = ~n2711 & ~po129 ;
  assign po8  = n3141 | n3142;
  assign n3144 = ~n2631 & po129 ;
  assign n3145 = ~n2634 & ~po129 ;
  assign po9  = n3144 | n3145;
  assign n3147 = ~n2626 & po129 ;
  assign n3148 = ~n2623 & ~po129 ;
  assign po10  = n3147 | n3148;
  assign n3150 = ~n2618 & po129 ;
  assign n3151 = ~n2615 & ~po129 ;
  assign po11  = n3150 | n3151;
  assign n3153 = ~n2610 & po129 ;
  assign n3154 = ~n2607 & ~po129 ;
  assign po12  = n3153 | n3154;
  assign n3156 = ~n2602 & po129 ;
  assign n3157 = ~n2599 & ~po129 ;
  assign po13  = n3156 | n3157;
  assign n3159 = ~n2594 & po129 ;
  assign n3160 = ~n2591 & ~po129 ;
  assign po14  = n3159 | n3160;
  assign n3162 = ~n2586 & po129 ;
  assign n3163 = ~n2583 & ~po129 ;
  assign po15  = n3162 | n3163;
  assign n3165 = ~n2740 & po129 ;
  assign n3166 = ~n2737 & ~po129 ;
  assign po16  = n3165 | n3166;
  assign n3168 = ~n2577 & po129 ;
  assign n3169 = ~n2580 & ~po129 ;
  assign po17  = n3168 | n3169;
  assign n3171 = ~n2572 & po129 ;
  assign n3172 = ~n2569 & ~po129 ;
  assign po18  = n3171 | n3172;
  assign n3174 = ~n2564 & po129 ;
  assign n3175 = ~n2561 & ~po129 ;
  assign po19  = n3174 | n3175;
  assign n3177 = ~n2556 & po129 ;
  assign n3178 = ~n2553 & ~po129 ;
  assign po20  = n3177 | n3178;
  assign n3180 = ~n2548 & po129 ;
  assign n3181 = ~n2545 & ~po129 ;
  assign po21  = n3180 | n3181;
  assign n3183 = ~n2540 & po129 ;
  assign n3184 = ~n2537 & ~po129 ;
  assign po22  = n3183 | n3184;
  assign n3186 = ~n2532 & po129 ;
  assign n3187 = ~n2529 & ~po129 ;
  assign po23  = n3186 | n3187;
  assign n3189 = ~n2766 & po129 ;
  assign n3190 = ~n2763 & ~po129 ;
  assign po24  = n3189 | n3190;
  assign n3192 = ~n2523 & po129 ;
  assign n3193 = ~n2526 & ~po129 ;
  assign po25  = n3192 | n3193;
  assign n3195 = ~n2518 & po129 ;
  assign n3196 = ~n2515 & ~po129 ;
  assign po26  = n3195 | n3196;
  assign n3198 = ~n2510 & po129 ;
  assign n3199 = ~n2507 & ~po129 ;
  assign po27  = n3198 | n3199;
  assign n3201 = ~n2502 & po129 ;
  assign n3202 = ~n2499 & ~po129 ;
  assign po28  = n3201 | n3202;
  assign n3204 = ~n2494 & po129 ;
  assign n3205 = ~n2491 & ~po129 ;
  assign po29  = n3204 | n3205;
  assign n3207 = ~n2485 & po129 ;
  assign n3208 = ~n2482 & ~po129 ;
  assign po30  = n3207 | n3208;
  assign n3210 = ~n2455 & po129 ;
  assign n3211 = ~n2452 & ~po129 ;
  assign po31  = n3210 | n3211;
  assign n3213 = ~n2413 & po129 ;
  assign n3214 = ~n2416 & ~po129 ;
  assign po32  = n3213 | n3214;
  assign n3216 = ~n2469 & po129 ;
  assign n3217 = ~n2466 & ~po129 ;
  assign po33  = n3216 | n3217;
  assign n3219 = ~n2473 & po129 ;
  assign n3220 = ~n2476 & ~po129 ;
  assign po34  = n3219 | n3220;
  assign n3222 = ~n2462 & po129 ;
  assign n3223 = ~n2459 & ~po129 ;
  assign po35  = n3222 | n3223;
  assign n3225 = ~n2423 & po129 ;
  assign n3226 = ~n2420 & ~po129 ;
  assign po36  = n3225 | n3226;
  assign n3228 = ~n2444 & po129 ;
  assign n3229 = ~n2441 & ~po129 ;
  assign po37  = n3228 | n3229;
  assign n3231 = ~n2430 & po129 ;
  assign n3232 = ~n2427 & ~po129 ;
  assign po38  = n3231 | n3232;
  assign n3234 = ~n2437 & po129 ;
  assign n3235 = ~n2434 & ~po129 ;
  assign po39  = n3234 | n3235;
  assign n3237 = ~n2363 & po129 ;
  assign n3238 = ~n2359 & ~po129 ;
  assign po40  = n3237 | n3238;
  assign n3240 = ~n2355 & po129 ;
  assign n3241 = ~n2352 & ~po129 ;
  assign po41  = n3240 | n3241;
  assign n3243 = ~n2346 & po129 ;
  assign n3244 = ~n2343 & ~po129 ;
  assign po42  = n3243 | n3244;
  assign n3246 = ~n2338 & po129 ;
  assign n3247 = ~n2335 & ~po129 ;
  assign po43  = n3246 | n3247;
  assign n3249 = ~n2398 & po129 ;
  assign n3250 = ~n2395 & ~po129 ;
  assign po44  = n3249 | n3250;
  assign n3252 = ~n2391 & po129 ;
  assign n3253 = ~n2388 & ~po129 ;
  assign po45  = n3252 | n3253;
  assign n3255 = ~n2383 & po129 ;
  assign n3256 = ~n2379 & ~po129 ;
  assign po46  = n3255 | n3256;
  assign n3258 = ~n2375 & po129 ;
  assign n3259 = ~n2372 & ~po129 ;
  assign po47  = n3258 | n3259;
  assign n3261 = ~n2328 & po129 ;
  assign n3262 = ~n2331 & ~po129 ;
  assign po48  = n3261 | n3262;
  assign n3264 = ~n2856 & po129 ;
  assign n3265 = ~n2853 & ~po129 ;
  assign po49  = n3264 | n3265;
  assign n3267 = ~n2860 & po129 ;
  assign n3268 = ~n2863 & ~po129 ;
  assign po50  = n3267 | n3268;
  assign n3270 = ~n2849 & po129 ;
  assign n3271 = ~n2846 & ~po129 ;
  assign po51  = n3270 | n3271;
  assign n3273 = ~n2827 & po129 ;
  assign n3274 = ~n2830 & ~po129 ;
  assign po52  = n3273 | n3274;
  assign n3276 = ~n2823 & po129 ;
  assign n3277 = ~n2820 & ~po129 ;
  assign po53  = n3276 | n3277;
  assign n3279 = ~n2835 & po129 ;
  assign n3280 = ~n2838 & ~po129 ;
  assign po54  = n3279 | n3280;
  assign n3282 = ~n2324 & po129 ;
  assign n3283 = ~n2321 & ~po129 ;
  assign po55  = n3282 | n3283;
  assign n3285 = ~n2271 & po129 ;
  assign n3286 = ~n2267 & ~po129 ;
  assign po56  = n3285 | n3286;
  assign n3288 = ~n2263 & po129 ;
  assign n3289 = ~n2260 & ~po129 ;
  assign po57  = n3288 | n3289;
  assign n3291 = ~n2254 & po129 ;
  assign n3292 = ~n2251 & ~po129 ;
  assign po58  = n3291 | n3292;
  assign n3294 = ~n2246 & po129 ;
  assign n3295 = ~n2243 & ~po129 ;
  assign po59  = n3294 | n3295;
  assign n3297 = ~n2306 & po129 ;
  assign n3298 = ~n2303 & ~po129 ;
  assign po60  = n3297 | n3298;
  assign n3300 = ~n2299 & po129 ;
  assign n3301 = ~n2296 & ~po129 ;
  assign po61  = n3300 | n3301;
  assign n3303 = ~n2291 & po129 ;
  assign n3304 = ~n2287 & ~po129 ;
  assign po62  = n3303 | n3304;
  assign n3306 = ~n2283 & po129 ;
  assign n3307 = ~n2280 & ~po129 ;
  assign po63  = n3306 | n3307;
  assign n3309 = ~n2901 & po129 ;
  assign n3310 = ~n2904 & ~po129 ;
  assign po64  = n3309 | n3310;
  assign n3312 = ~n2224 & po129 ;
  assign n3313 = ~n2221 & ~po129 ;
  assign po65  = n3312 | n3313;
  assign n3315 = ~n2235 & po129 ;
  assign n3316 = ~n2238 & ~po129 ;
  assign po66  = n3315 | n3316;
  assign n3318 = ~n2231 & po129 ;
  assign n3319 = ~n2228 & ~po129 ;
  assign po67  = n3318 | n3319;
  assign n3321 = ~n2213 & po129 ;
  assign n3322 = ~n2209 & ~po129 ;
  assign po68  = n3321 | n3322;
  assign n3324 = ~n2205 & po129 ;
  assign n3325 = ~n2202 & ~po129 ;
  assign po69  = n3324 | n3325;
  assign n3327 = ~n2185 & po129 ;
  assign n3328 = ~n2195 & ~po129 ;
  assign po70  = n3327 | n3328;
  assign n3330 = ~n2191 & po129 ;
  assign n3331 = ~n2188 & ~po129 ;
  assign po71  = n3330 | n3331;
  assign n3333 = ~n2928 & po129 ;
  assign n3334 = ~n2931 & ~po129 ;
  assign po72  = n3333 | n3334;
  assign n3336 = ~n2166 & po129 ;
  assign n3337 = ~n2163 & ~po129 ;
  assign po73  = n3336 | n3337;
  assign n3339 = ~n2177 & po129 ;
  assign n3340 = ~n2180 & ~po129 ;
  assign po74  = n3339 | n3340;
  assign n3342 = ~n2173 & po129 ;
  assign n3343 = ~n2170 & ~po129 ;
  assign po75  = n3342 | n3343;
  assign n3345 = ~n2155 & po129 ;
  assign n3346 = ~n2151 & ~po129 ;
  assign po76  = n3345 | n3346;
  assign n3348 = ~n2147 & po129 ;
  assign n3349 = ~n2144 & ~po129 ;
  assign po77  = n3348 | n3349;
  assign n3351 = ~n2127 & po129 ;
  assign n3352 = ~n2137 & ~po129 ;
  assign po78  = n3351 | n3352;
  assign n3354 = ~n2133 & po129 ;
  assign n3355 = ~n2130 & ~po129 ;
  assign po79  = n3354 | n3355;
  assign n3357 = ~n2955 & po129 ;
  assign n3358 = ~n2958 & ~po129 ;
  assign po80  = n3357 | n3358;
  assign n3360 = ~n2108 & po129 ;
  assign n3361 = ~n2105 & ~po129 ;
  assign po81  = n3360 | n3361;
  assign n3363 = ~n2119 & po129 ;
  assign n3364 = ~n2122 & ~po129 ;
  assign po82  = n3363 | n3364;
  assign n3366 = ~n2115 & po129 ;
  assign n3367 = ~n2112 & ~po129 ;
  assign po83  = n3366 | n3367;
  assign n3369 = ~n2097 & po129 ;
  assign n3370 = ~n2093 & ~po129 ;
  assign po84  = n3369 | n3370;
  assign n3372 = ~n2089 & po129 ;
  assign n3373 = ~n2086 & ~po129 ;
  assign po85  = n3372 | n3373;
  assign n3375 = ~n2069 & po129 ;
  assign n3376 = ~n2079 & ~po129 ;
  assign po86  = n3375 | n3376;
  assign n3378 = ~n2075 & po129 ;
  assign n3379 = ~n2072 & ~po129 ;
  assign po87  = n3378 | n3379;
  assign n3381 = ~n2982 & po129 ;
  assign n3382 = ~n2985 & ~po129 ;
  assign po88  = n3381 | n3382;
  assign n3384 = ~n2050 & po129 ;
  assign n3385 = ~n2047 & ~po129 ;
  assign po89  = n3384 | n3385;
  assign n3387 = ~n2061 & po129 ;
  assign n3388 = ~n2064 & ~po129 ;
  assign po90  = n3387 | n3388;
  assign n3390 = ~n2057 & po129 ;
  assign n3391 = ~n2054 & ~po129 ;
  assign po91  = n3390 | n3391;
  assign n3393 = ~n2039 & po129 ;
  assign n3394 = ~n2035 & ~po129 ;
  assign po92  = n3393 | n3394;
  assign n3396 = ~n2031 & po129 ;
  assign n3397 = ~n2028 & ~po129 ;
  assign po93  = n3396 | n3397;
  assign n3399 = ~n2011 & po129 ;
  assign n3400 = ~n2021 & ~po129 ;
  assign po94  = n3399 | n3400;
  assign n3402 = ~n2017 & po129 ;
  assign n3403 = ~n2014 & ~po129 ;
  assign po95  = n3402 | n3403;
  assign n3405 = ~n3009 & po129 ;
  assign n3406 = ~n3012 & ~po129 ;
  assign po96  = n3405 | n3406;
  assign n3408 = ~n1992 & po129 ;
  assign n3409 = ~n1989 & ~po129 ;
  assign po97  = n3408 | n3409;
  assign n3411 = ~n2003 & po129 ;
  assign n3412 = ~n2006 & ~po129 ;
  assign po98  = n3411 | n3412;
  assign n3414 = ~n1999 & po129 ;
  assign n3415 = ~n1996 & ~po129 ;
  assign po99  = n3414 | n3415;
  assign n3417 = ~n1981 & po129 ;
  assign n3418 = ~n1977 & ~po129 ;
  assign po100  = n3417 | n3418;
  assign n3420 = ~n1973 & po129 ;
  assign n3421 = ~n1970 & ~po129 ;
  assign po101  = n3420 | n3421;
  assign n3423 = ~n1953 & po129 ;
  assign n3424 = ~n1963 & ~po129 ;
  assign po102  = n3423 | n3424;
  assign n3426 = ~n1959 & po129 ;
  assign n3427 = ~n1956 & ~po129 ;
  assign po103  = n3426 | n3427;
  assign n3429 = ~n3036 & po129 ;
  assign n3430 = ~n3039 & ~po129 ;
  assign po104  = n3429 | n3430;
  assign n3432 = ~n1934 & po129 ;
  assign n3433 = ~n1931 & ~po129 ;
  assign po105  = n3432 | n3433;
  assign n3435 = ~n1945 & po129 ;
  assign n3436 = ~n1948 & ~po129 ;
  assign po106  = n3435 | n3436;
  assign n3438 = ~n1941 & po129 ;
  assign n3439 = ~n1938 & ~po129 ;
  assign po107  = n3438 | n3439;
  assign n3441 = ~n1923 & po129 ;
  assign n3442 = ~n1919 & ~po129 ;
  assign po108  = n3441 | n3442;
  assign n3444 = ~n1915 & po129 ;
  assign n3445 = ~n1912 & ~po129 ;
  assign po109  = n3444 | n3445;
  assign n3447 = ~n1895 & po129 ;
  assign n3448 = ~n1905 & ~po129 ;
  assign po110  = n3447 | n3448;
  assign n3450 = ~n1901 & po129 ;
  assign n3451 = ~n1898 & ~po129 ;
  assign po111  = n3450 | n3451;
  assign n3453 = ~n3063 & po129 ;
  assign n3454 = ~n3066 & ~po129 ;
  assign po112  = n3453 | n3454;
  assign n3456 = ~n1876 & po129 ;
  assign n3457 = ~n1873 & ~po129 ;
  assign po113  = n3456 | n3457;
  assign n3459 = ~n1887 & po129 ;
  assign n3460 = ~n1890 & ~po129 ;
  assign po114  = n3459 | n3460;
  assign n3462 = ~n1883 & po129 ;
  assign n3463 = ~n1880 & ~po129 ;
  assign po115  = n3462 | n3463;
  assign n3465 = ~n1847 & po129 ;
  assign n3466 = ~n1844 & ~po129 ;
  assign po116  = n3465 | n3466;
  assign n3468 = ~n1840 & po129 ;
  assign n3469 = ~n1837 & ~po129 ;
  assign po117  = n3468 | n3469;
  assign n3471 = ~n1861 & po129 ;
  assign n3472 = ~n1864 & ~po129 ;
  assign po118  = n3471 | n3472;
  assign n3474 = ~n1855 & po129 ;
  assign n3475 = ~n1852 & ~po129 ;
  assign po119  = n3474 | n3475;
  assign n3477 = ~n3098 & po129 ;
  assign n3478 = ~n3095 & ~po129 ;
  assign po120  = n3477 | n3478;
  assign n3480 = ~n3091 & po129 ;
  assign n3481 = ~n3088 & ~po129 ;
  assign po121  = n3480 | n3481;
  assign n3483 = ~n1829 & po129 ;
  assign n3484 = ~n1832 & ~po129 ;
  assign po122  = n3483 | n3484;
  assign n3486 = ~n1825 & po129 ;
  assign n3487 = ~n1822 & ~po129 ;
  assign po123  = n3486 | n3487;
  assign n3489 = ~n1810 & po129 ;
  assign n3490 = ~n1807 & ~po129 ;
  assign po124  = n3489 | n3490;
  assign n3492 = ~n1802 & po129 ;
  assign n3493 = ~n1799 & ~po129 ;
  assign po125  = n3492 | n3493;
  assign n3495 = ~n1795 & po129 ;
  assign n3496 = ~n1792 & ~po129 ;
  assign po126  = n3495 | n3496;
  assign po127  = n1216 & n1217;
  assign n3499 = n1789 & ~po129 ;
  assign n3500 = n1212 & po129 ;
  assign po128  = n3499 | n3500;
endmodule
