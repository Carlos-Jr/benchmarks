module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 , pi32 ,
    pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 , pi40 ,
    pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 , pi56 ,
    pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 , pi64 ,
    pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 , pi73 ,
    pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 , pi81 ,
    pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 , pi89 ,
    pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 , pi97 ,
    pi98 , pi99 , pi100 , pi101 , pi102 , pi103 , pi104 , pi105 ,
    pi106 , pi107 , pi108 , pi109 , pi110 , pi111 , pi112 , pi113 ,
    pi114 , pi115 , pi116 , pi117 , pi118 , pi119 , pi120 , pi121 ,
    pi122 , pi123 , pi124 , pi125 , pi126 , pi127 ,
    po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7 , po8 ,
    po9 , po10 , po11 , po12 , po13 , po14 , po15 , po16 ,
    po17 , po18 , po19 , po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 , po30 , po31 , po32 ,
    po33 , po34 , po35 , po36 , po37 , po38 , po39 , po40 ,
    po41 , po42 , po43 , po44 , po45 , po46 , po47 , po48 ,
    po49 , po50 , po51 , po52 , po53 , po54 , po55 , po56 ,
    po57 , po58 , po59 , po60 , po61 , po62 , po63 , po64 ,
    po65 , po66 , po67 , po68 , po69 , po70 , po71 , po72 ,
    po73 , po74 , po75 , po76 , po77 , po78 , po79 , po80 ,
    po81 , po82 , po83 , po84 , po85 , po86 , po87 , po88 ,
    po89 , po90 , po91 , po92 , po93 , po94 , po95 , po96 ,
    po97 , po98 , po99 , po100 , po101 , po102 , po103 ,
    po104 , po105 , po106 , po107 , po108 , po109 , po110 ,
    po111 , po112 , po113 , po114 , po115 , po116 , po117 ,
    po118 , po119 , po120 , po121 , po122 , po123 , po124 ,
    po125 , po126 , po127   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    pi32 , pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 ,
    pi56 , pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 ,
    pi64 , pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 ,
    pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 ,
    pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 ,
    pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 ,
    pi97 , pi98 , pi99 , pi100 , pi101 , pi102 , pi103 , pi104 ,
    pi105 , pi106 , pi107 , pi108 , pi109 , pi110 , pi111 , pi112 ,
    pi113 , pi114 , pi115 , pi116 , pi117 , pi118 , pi119 , pi120 ,
    pi121 , pi122 , pi123 , pi124 , pi125 , pi126 , pi127 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7 ,
    po8 , po9 , po10 , po11 , po12 , po13 , po14 , po15 ,
    po16 , po17 , po18 , po19 , po20 , po21 , po22 , po23 ,
    po24 , po25 , po26 , po27 , po28 , po29 , po30 , po31 ,
    po32 , po33 , po34 , po35 , po36 , po37 , po38 , po39 ,
    po40 , po41 , po42 , po43 , po44 , po45 , po46 , po47 ,
    po48 , po49 , po50 , po51 , po52 , po53 , po54 , po55 ,
    po56 , po57 , po58 , po59 , po60 , po61 , po62 , po63 ,
    po64 , po65 , po66 , po67 , po68 , po69 , po70 , po71 ,
    po72 , po73 , po74 , po75 , po76 , po77 , po78 , po79 ,
    po80 , po81 , po82 , po83 , po84 , po85 , po86 , po87 ,
    po88 , po89 , po90 , po91 , po92 , po93 , po94 , po95 ,
    po96 , po97 , po98 , po99 , po100 , po101 , po102 ,
    po103 , po104 , po105 , po106 , po107 , po108 , po109 ,
    po110 , po111 , po112 , po113 , po114 , po115 , po116 ,
    po117 , po118 , po119 , po120 , po121 , po122 , po123 ,
    po124 , po125 , po126 , po127 ;
  wire n258, n259, n260, n261, n262, n263, n264,
    n265, n266, n267, n268, n269, n270, n271,
    n272, n273, n274, n276, n277, n278, n279,
    n280, n281, n282, n283, n284, n285, n286,
    n287, n288, n289, n290, n291, n292, n293,
    n295, n296, n297, n298, n299, n300, n301,
    n302, n303, n304, n305, n306, n307, n308,
    n309, n310, n311, n312, n313, n314, n315,
    n316, n317, n318, n319, n320, n321, n322,
    n324, n325, n326, n327, n328, n329, n330,
    n331, n332, n333, n334, n335, n336, n337,
    n338, n339, n340, n341, n342, n343, n344,
    n345, n346, n347, n348, n349, n350, n351,
    n352, n353, n354, n355, n356, n357, n358,
    n359, n360, n361, n362, n363, n364, n366,
    n367, n368, n369, n370, n371, n372, n373,
    n374, n375, n376, n377, n378, n379, n380,
    n381, n382, n383, n384, n385, n386, n387,
    n388, n389, n390, n391, n392, n393, n394,
    n395, n396, n397, n398, n399, n400, n401,
    n402, n403, n405, n406, n407, n408, n409,
    n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423,
    n424, n425, n426, n427, n428, n429, n430,
    n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444,
    n445, n446, n447, n448, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487,
    n488, n489, n490, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501,
    n502, n503, n504, n505, n506, n507, n509,
    n510, n511, n512, n513, n514, n515, n516,
    n517, n518, n519, n520, n521, n522, n523,
    n524, n525, n526, n527, n528, n529, n530,
    n531, n532, n533, n534, n535, n536, n537,
    n538, n539, n540, n541, n542, n543, n544,
    n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n557, n558,
    n559, n560, n561, n562, n563, n565, n566,
    n567, n568, n569, n570, n571, n572, n573,
    n574, n575, n576, n577, n578, n579, n580,
    n581, n582, n583, n584, n585, n586, n587,
    n588, n589, n590, n591, n592, n593, n594,
    n595, n596, n597, n598, n599, n600, n601,
    n602, n603, n604, n605, n606, n607, n608,
    n609, n610, n611, n612, n613, n614, n615,
    n616, n617, n618, n619, n620, n621, n622,
    n623, n624, n625, n627, n628, n629, n630,
    n631, n632, n633, n634, n635, n636, n637,
    n638, n639, n640, n641, n642, n643, n644,
    n645, n646, n647, n648, n649, n650, n651,
    n652, n653, n654, n655, n656, n657, n658,
    n659, n660, n661, n662, n663, n664, n665,
    n666, n667, n668, n669, n670, n671, n672,
    n673, n674, n675, n676, n677, n678, n679,
    n680, n681, n682, n683, n684, n685, n686,
    n687, n688, n689, n690, n691, n692, n693,
    n694, n695, n696, n697, n698, n699, n700,
    n701, n703, n704, n705, n706, n707, n708,
    n709, n710, n711, n712, n713, n714, n715,
    n716, n717, n718, n719, n720, n721, n722,
    n723, n724, n725, n726, n727, n728, n729,
    n730, n731, n732, n733, n734, n735, n736,
    n737, n738, n739, n740, n741, n742, n743,
    n744, n745, n746, n747, n748, n749, n750,
    n751, n752, n753, n754, n755, n756, n757,
    n758, n759, n760, n761, n762, n763, n764,
    n765, n766, n767, n768, n769, n770, n771,
    n772, n773, n774, n776, n777, n778, n779,
    n780, n781, n782, n783, n784, n785, n786,
    n787, n788, n789, n790, n791, n792, n793,
    n794, n795, n796, n797, n798, n799, n800,
    n801, n802, n803, n804, n805, n806, n807,
    n808, n809, n810, n811, n812, n813, n814,
    n815, n816, n817, n818, n819, n820, n821,
    n822, n823, n824, n825, n826, n827, n828,
    n829, n830, n831, n832, n833, n834, n835,
    n836, n837, n838, n839, n840, n841, n842,
    n843, n844, n845, n846, n847, n848, n849,
    n850, n851, n852, n853, n855, n856, n857,
    n858, n859, n860, n861, n862, n863, n864,
    n865, n866, n867, n868, n869, n870, n871,
    n872, n873, n874, n875, n876, n877, n878,
    n879, n880, n881, n882, n883, n884, n885,
    n886, n887, n888, n889, n890, n891, n892,
    n893, n894, n895, n896, n897, n898, n899,
    n900, n901, n902, n903, n904, n905, n906,
    n907, n908, n909, n910, n911, n912, n913,
    n914, n915, n916, n917, n918, n919, n920,
    n921, n922, n923, n924, n925, n926, n927,
    n928, n929, n930, n931, n932, n933, n934,
    n935, n936, n937, n938, n939, n940, n941,
    n942, n943, n944, n945, n946, n948, n949,
    n950, n951, n952, n953, n954, n955, n956,
    n957, n958, n959, n960, n961, n962, n963,
    n964, n965, n966, n967, n968, n969, n970,
    n971, n972, n973, n974, n975, n976, n977,
    n978, n979, n980, n981, n982, n983, n984,
    n985, n986, n987, n988, n989, n990, n991,
    n992, n993, n994, n995, n996, n997, n998,
    n999, n1000, n1001, n1002, n1003, n1004,
    n1005, n1006, n1007, n1008, n1009, n1010,
    n1011, n1012, n1013, n1014, n1015, n1016,
    n1017, n1018, n1019, n1020, n1021, n1022,
    n1023, n1024, n1025, n1026, n1027, n1028,
    n1029, n1030, n1031, n1032, n1033, n1034,
    n1035, n1036, n1038, n1039, n1040, n1041,
    n1042, n1043, n1044, n1045, n1046, n1047,
    n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059,
    n1060, n1061, n1062, n1063, n1064, n1065,
    n1066, n1067, n1068, n1069, n1070, n1071,
    n1072, n1073, n1074, n1075, n1076, n1077,
    n1078, n1079, n1080, n1081, n1082, n1083,
    n1084, n1085, n1086, n1087, n1088, n1089,
    n1090, n1091, n1092, n1093, n1094, n1095,
    n1096, n1097, n1098, n1099, n1100, n1101,
    n1102, n1103, n1104, n1105, n1106, n1107,
    n1108, n1109, n1110, n1111, n1112, n1113,
    n1114, n1115, n1116, n1117, n1118, n1119,
    n1120, n1121, n1122, n1123, n1124, n1125,
    n1126, n1127, n1128, n1129, n1130, n1131,
    n1132, n1134, n1135, n1136, n1137, n1138,
    n1139, n1140, n1141, n1142, n1143, n1144,
    n1145, n1146, n1147, n1148, n1149, n1150,
    n1151, n1152, n1153, n1154, n1155, n1156,
    n1157, n1158, n1159, n1160, n1161, n1162,
    n1163, n1164, n1165, n1166, n1167, n1168,
    n1169, n1170, n1171, n1172, n1173, n1174,
    n1175, n1176, n1177, n1178, n1179, n1180,
    n1181, n1182, n1183, n1184, n1185, n1186,
    n1187, n1188, n1189, n1190, n1191, n1192,
    n1193, n1194, n1195, n1196, n1197, n1198,
    n1199, n1200, n1201, n1202, n1203, n1204,
    n1205, n1206, n1207, n1208, n1209, n1210,
    n1211, n1212, n1213, n1214, n1215, n1216,
    n1217, n1218, n1219, n1220, n1221, n1222,
    n1223, n1224, n1225, n1226, n1227, n1228,
    n1229, n1230, n1231, n1232, n1233, n1234,
    n1235, n1236, n1237, n1238, n1239, n1240,
    n1241, n1242, n1244, n1245, n1246, n1247,
    n1248, n1249, n1250, n1251, n1252, n1253,
    n1254, n1255, n1256, n1257, n1258, n1259,
    n1260, n1261, n1262, n1263, n1264, n1265,
    n1266, n1267, n1268, n1269, n1270, n1271,
    n1272, n1273, n1274, n1275, n1276, n1277,
    n1278, n1279, n1280, n1281, n1282, n1283,
    n1284, n1285, n1286, n1287, n1288, n1289,
    n1290, n1291, n1292, n1293, n1294, n1295,
    n1296, n1297, n1298, n1299, n1300, n1301,
    n1302, n1303, n1304, n1305, n1306, n1307,
    n1308, n1309, n1310, n1311, n1312, n1313,
    n1314, n1315, n1316, n1317, n1318, n1319,
    n1320, n1321, n1322, n1323, n1324, n1325,
    n1326, n1327, n1328, n1329, n1330, n1331,
    n1332, n1333, n1334, n1335, n1336, n1337,
    n1338, n1339, n1340, n1341, n1342, n1343,
    n1344, n1345, n1346, n1347, n1348, n1349,
    n1351, n1352, n1353, n1354, n1355, n1356,
    n1357, n1358, n1359, n1360, n1361, n1362,
    n1363, n1364, n1365, n1366, n1367, n1368,
    n1369, n1370, n1371, n1372, n1373, n1374,
    n1375, n1376, n1377, n1378, n1379, n1380,
    n1381, n1382, n1383, n1384, n1385, n1386,
    n1387, n1388, n1389, n1390, n1391, n1392,
    n1393, n1394, n1395, n1396, n1397, n1398,
    n1399, n1400, n1401, n1402, n1403, n1404,
    n1405, n1406, n1407, n1408, n1409, n1410,
    n1411, n1412, n1413, n1414, n1415, n1416,
    n1417, n1418, n1419, n1420, n1421, n1422,
    n1423, n1424, n1425, n1426, n1427, n1428,
    n1429, n1430, n1431, n1432, n1433, n1434,
    n1435, n1436, n1437, n1438, n1439, n1440,
    n1441, n1442, n1443, n1444, n1445, n1446,
    n1447, n1448, n1449, n1450, n1451, n1452,
    n1453, n1454, n1455, n1456, n1457, n1458,
    n1459, n1460, n1461, n1462, n1464, n1465,
    n1466, n1467, n1468, n1469, n1470, n1471,
    n1472, n1473, n1474, n1475, n1476, n1477,
    n1478, n1479, n1480, n1481, n1482, n1483,
    n1484, n1485, n1486, n1487, n1488, n1489,
    n1490, n1491, n1492, n1493, n1494, n1495,
    n1496, n1497, n1498, n1499, n1500, n1501,
    n1502, n1503, n1504, n1505, n1506, n1507,
    n1508, n1509, n1510, n1511, n1512, n1513,
    n1514, n1515, n1516, n1517, n1518, n1519,
    n1520, n1521, n1522, n1523, n1524, n1525,
    n1526, n1527, n1528, n1529, n1530, n1531,
    n1532, n1533, n1534, n1535, n1536, n1537,
    n1538, n1539, n1540, n1541, n1542, n1543,
    n1544, n1545, n1546, n1547, n1548, n1549,
    n1550, n1551, n1552, n1553, n1554, n1555,
    n1556, n1557, n1558, n1559, n1560, n1561,
    n1562, n1563, n1564, n1565, n1566, n1567,
    n1568, n1569, n1570, n1571, n1572, n1573,
    n1574, n1575, n1576, n1577, n1578, n1579,
    n1580, n1581, n1582, n1583, n1584, n1585,
    n1586, n1587, n1588, n1589, n1591, n1592,
    n1593, n1594, n1595, n1596, n1597, n1598,
    n1599, n1600, n1601, n1602, n1603, n1604,
    n1605, n1606, n1607, n1608, n1609, n1610,
    n1611, n1612, n1613, n1614, n1615, n1616,
    n1617, n1618, n1619, n1620, n1621, n1622,
    n1623, n1624, n1625, n1626, n1627, n1628,
    n1629, n1630, n1631, n1632, n1633, n1634,
    n1635, n1636, n1637, n1638, n1639, n1640,
    n1641, n1642, n1643, n1644, n1645, n1646,
    n1647, n1648, n1649, n1650, n1651, n1652,
    n1653, n1654, n1655, n1656, n1657, n1658,
    n1659, n1660, n1661, n1662, n1663, n1664,
    n1665, n1666, n1667, n1668, n1669, n1670,
    n1671, n1672, n1673, n1674, n1675, n1676,
    n1677, n1678, n1679, n1680, n1681, n1682,
    n1683, n1684, n1685, n1686, n1687, n1688,
    n1689, n1690, n1691, n1692, n1693, n1694,
    n1695, n1696, n1697, n1698, n1699, n1700,
    n1701, n1702, n1703, n1704, n1705, n1706,
    n1707, n1708, n1709, n1710, n1711, n1712,
    n1713, n1715, n1716, n1717, n1718, n1719,
    n1720, n1721, n1722, n1723, n1724, n1725,
    n1726, n1727, n1728, n1729, n1730, n1731,
    n1732, n1733, n1734, n1735, n1736, n1737,
    n1738, n1739, n1740, n1741, n1742, n1743,
    n1744, n1745, n1746, n1747, n1748, n1749,
    n1750, n1751, n1752, n1753, n1754, n1755,
    n1756, n1757, n1758, n1759, n1760, n1761,
    n1762, n1763, n1764, n1765, n1766, n1767,
    n1768, n1769, n1770, n1771, n1772, n1773,
    n1774, n1775, n1776, n1777, n1778, n1779,
    n1780, n1781, n1782, n1783, n1784, n1785,
    n1786, n1787, n1788, n1789, n1790, n1791,
    n1792, n1793, n1794, n1795, n1796, n1797,
    n1798, n1799, n1800, n1801, n1802, n1803,
    n1804, n1805, n1806, n1807, n1808, n1809,
    n1810, n1811, n1812, n1813, n1814, n1815,
    n1816, n1817, n1818, n1819, n1820, n1821,
    n1822, n1823, n1824, n1825, n1826, n1827,
    n1828, n1829, n1830, n1831, n1832, n1833,
    n1834, n1835, n1836, n1837, n1838, n1839,
    n1840, n1841, n1842, n1843, n1845, n1846,
    n1847, n1848, n1849, n1850, n1851, n1852,
    n1853, n1854, n1855, n1856, n1857, n1858,
    n1859, n1860, n1861, n1862, n1863, n1864,
    n1865, n1866, n1867, n1868, n1869, n1870,
    n1871, n1872, n1873, n1874, n1875, n1876,
    n1877, n1878, n1879, n1880, n1881, n1882,
    n1883, n1884, n1885, n1886, n1887, n1888,
    n1889, n1890, n1891, n1892, n1893, n1894,
    n1895, n1896, n1897, n1898, n1899, n1900,
    n1901, n1902, n1903, n1904, n1905, n1906,
    n1907, n1908, n1909, n1910, n1911, n1912,
    n1913, n1914, n1915, n1916, n1917, n1918,
    n1919, n1920, n1921, n1922, n1923, n1924,
    n1925, n1926, n1927, n1928, n1929, n1930,
    n1931, n1932, n1933, n1934, n1935, n1936,
    n1937, n1938, n1939, n1940, n1941, n1942,
    n1943, n1944, n1945, n1946, n1947, n1948,
    n1949, n1950, n1951, n1952, n1953, n1954,
    n1955, n1956, n1957, n1958, n1959, n1960,
    n1961, n1962, n1963, n1964, n1965, n1966,
    n1967, n1968, n1969, n1970, n1971, n1972,
    n1973, n1974, n1975, n1976, n1977, n1978,
    n1979, n1980, n1981, n1982, n1983, n1984,
    n1985, n1986, n1987, n1989, n1990, n1991,
    n1992, n1993, n1994, n1995, n1996, n1997,
    n1998, n1999, n2000, n2001, n2002, n2003,
    n2004, n2005, n2006, n2007, n2008, n2009,
    n2010, n2011, n2012, n2013, n2014, n2015,
    n2016, n2017, n2018, n2019, n2020, n2021,
    n2022, n2023, n2024, n2025, n2026, n2027,
    n2028, n2029, n2030, n2031, n2032, n2033,
    n2034, n2035, n2036, n2037, n2038, n2039,
    n2040, n2041, n2042, n2043, n2044, n2045,
    n2046, n2047, n2048, n2049, n2050, n2051,
    n2052, n2053, n2054, n2055, n2056, n2057,
    n2058, n2059, n2060, n2061, n2062, n2063,
    n2064, n2065, n2066, n2067, n2068, n2069,
    n2070, n2071, n2072, n2073, n2074, n2075,
    n2076, n2077, n2078, n2079, n2080, n2081,
    n2082, n2083, n2084, n2085, n2086, n2087,
    n2088, n2089, n2090, n2091, n2092, n2093,
    n2094, n2095, n2096, n2097, n2098, n2099,
    n2100, n2101, n2102, n2103, n2104, n2105,
    n2106, n2107, n2108, n2109, n2110, n2111,
    n2112, n2113, n2114, n2115, n2116, n2117,
    n2118, n2119, n2120, n2121, n2122, n2123,
    n2124, n2125, n2126, n2127, n2128, n2130,
    n2131, n2132, n2133, n2134, n2135, n2136,
    n2137, n2138, n2139, n2140, n2141, n2142,
    n2143, n2144, n2145, n2146, n2147, n2148,
    n2149, n2150, n2151, n2152, n2153, n2154,
    n2155, n2156, n2157, n2158, n2159, n2160,
    n2161, n2162, n2163, n2164, n2165, n2166,
    n2167, n2168, n2169, n2170, n2171, n2172,
    n2173, n2174, n2175, n2176, n2177, n2178,
    n2179, n2180, n2181, n2182, n2183, n2184,
    n2185, n2186, n2187, n2188, n2189, n2190,
    n2191, n2192, n2193, n2194, n2195, n2196,
    n2197, n2198, n2199, n2200, n2201, n2202,
    n2203, n2204, n2205, n2206, n2207, n2208,
    n2209, n2210, n2211, n2212, n2213, n2214,
    n2215, n2216, n2217, n2218, n2219, n2220,
    n2221, n2222, n2223, n2224, n2225, n2226,
    n2227, n2228, n2229, n2230, n2231, n2232,
    n2233, n2234, n2235, n2236, n2237, n2238,
    n2239, n2240, n2241, n2242, n2243, n2244,
    n2245, n2246, n2247, n2248, n2249, n2250,
    n2251, n2252, n2253, n2254, n2255, n2256,
    n2257, n2258, n2259, n2260, n2261, n2262,
    n2263, n2264, n2265, n2266, n2267, n2268,
    n2269, n2270, n2271, n2272, n2273, n2274,
    n2275, n2277, n2278, n2279, n2280, n2281,
    n2282, n2283, n2284, n2285, n2286, n2287,
    n2288, n2289, n2290, n2291, n2292, n2293,
    n2294, n2295, n2296, n2297, n2298, n2299,
    n2300, n2301, n2302, n2303, n2304, n2305,
    n2306, n2307, n2308, n2309, n2310, n2311,
    n2312, n2313, n2314, n2315, n2316, n2317,
    n2318, n2319, n2320, n2321, n2322, n2323,
    n2324, n2325, n2326, n2327, n2328, n2329,
    n2330, n2331, n2332, n2333, n2334, n2335,
    n2336, n2337, n2338, n2339, n2340, n2341,
    n2342, n2343, n2344, n2345, n2346, n2347,
    n2348, n2349, n2350, n2351, n2352, n2353,
    n2354, n2355, n2356, n2357, n2358, n2359,
    n2360, n2361, n2362, n2363, n2364, n2365,
    n2366, n2367, n2368, n2369, n2370, n2371,
    n2372, n2373, n2374, n2375, n2376, n2377,
    n2378, n2379, n2380, n2381, n2382, n2383,
    n2384, n2385, n2386, n2387, n2388, n2389,
    n2390, n2391, n2392, n2393, n2394, n2395,
    n2396, n2397, n2398, n2399, n2400, n2401,
    n2402, n2403, n2404, n2405, n2406, n2407,
    n2408, n2409, n2410, n2411, n2412, n2413,
    n2414, n2415, n2416, n2417, n2418, n2419,
    n2420, n2421, n2422, n2423, n2424, n2425,
    n2426, n2427, n2428, n2429, n2430, n2431,
    n2432, n2433, n2434, n2435, n2436, n2438,
    n2439, n2440, n2441, n2442, n2443, n2444,
    n2445, n2446, n2447, n2448, n2449, n2450,
    n2451, n2452, n2453, n2454, n2455, n2456,
    n2457, n2458, n2459, n2460, n2461, n2462,
    n2463, n2464, n2465, n2466, n2467, n2468,
    n2469, n2470, n2471, n2472, n2473, n2474,
    n2475, n2476, n2477, n2478, n2479, n2480,
    n2481, n2482, n2483, n2484, n2485, n2486,
    n2487, n2488, n2489, n2490, n2491, n2492,
    n2493, n2494, n2495, n2496, n2497, n2498,
    n2499, n2500, n2501, n2502, n2503, n2504,
    n2505, n2506, n2507, n2508, n2509, n2510,
    n2511, n2512, n2513, n2514, n2515, n2516,
    n2517, n2518, n2519, n2520, n2521, n2522,
    n2523, n2524, n2525, n2526, n2527, n2528,
    n2529, n2530, n2531, n2532, n2533, n2534,
    n2535, n2536, n2537, n2538, n2539, n2540,
    n2541, n2542, n2543, n2544, n2545, n2546,
    n2547, n2548, n2549, n2550, n2551, n2552,
    n2553, n2554, n2555, n2556, n2557, n2558,
    n2559, n2560, n2561, n2562, n2563, n2564,
    n2565, n2566, n2567, n2568, n2569, n2570,
    n2571, n2572, n2573, n2574, n2575, n2576,
    n2577, n2578, n2579, n2580, n2581, n2582,
    n2583, n2584, n2585, n2586, n2587, n2588,
    n2589, n2590, n2591, n2592, n2593, n2594,
    n2596, n2597, n2598, n2599, n2600, n2601,
    n2602, n2603, n2604, n2605, n2606, n2607,
    n2608, n2609, n2610, n2611, n2612, n2613,
    n2614, n2615, n2616, n2617, n2618, n2619,
    n2620, n2621, n2622, n2623, n2624, n2625,
    n2626, n2627, n2628, n2629, n2630, n2631,
    n2632, n2633, n2634, n2635, n2636, n2637,
    n2638, n2639, n2640, n2641, n2642, n2643,
    n2644, n2645, n2646, n2647, n2648, n2649,
    n2650, n2651, n2652, n2653, n2654, n2655,
    n2656, n2657, n2658, n2659, n2660, n2661,
    n2662, n2663, n2664, n2665, n2666, n2667,
    n2668, n2669, n2670, n2671, n2672, n2673,
    n2674, n2675, n2676, n2677, n2678, n2679,
    n2680, n2681, n2682, n2683, n2684, n2685,
    n2686, n2687, n2688, n2689, n2690, n2691,
    n2692, n2693, n2694, n2695, n2696, n2697,
    n2698, n2699, n2700, n2701, n2702, n2703,
    n2704, n2705, n2706, n2707, n2708, n2709,
    n2710, n2711, n2712, n2713, n2714, n2715,
    n2716, n2717, n2718, n2719, n2720, n2721,
    n2722, n2723, n2724, n2725, n2726, n2727,
    n2728, n2729, n2730, n2731, n2732, n2733,
    n2734, n2735, n2736, n2737, n2738, n2739,
    n2740, n2741, n2742, n2743, n2744, n2745,
    n2746, n2747, n2748, n2749, n2750, n2751,
    n2752, n2753, n2754, n2755, n2756, n2757,
    n2758, n2760, n2761, n2762, n2763, n2764,
    n2765, n2766, n2767, n2768, n2769, n2770,
    n2771, n2772, n2773, n2774, n2775, n2776,
    n2777, n2778, n2779, n2780, n2781, n2782,
    n2783, n2784, n2785, n2786, n2787, n2788,
    n2789, n2790, n2791, n2792, n2793, n2794,
    n2795, n2796, n2797, n2798, n2799, n2800,
    n2801, n2802, n2803, n2804, n2805, n2806,
    n2807, n2808, n2809, n2810, n2811, n2812,
    n2813, n2814, n2815, n2816, n2817, n2818,
    n2819, n2820, n2821, n2822, n2823, n2824,
    n2825, n2826, n2827, n2828, n2829, n2830,
    n2831, n2832, n2833, n2834, n2835, n2836,
    n2837, n2838, n2839, n2840, n2841, n2842,
    n2843, n2844, n2845, n2846, n2847, n2848,
    n2849, n2850, n2851, n2852, n2853, n2854,
    n2855, n2856, n2857, n2858, n2859, n2860,
    n2861, n2862, n2863, n2864, n2865, n2866,
    n2867, n2868, n2869, n2870, n2871, n2872,
    n2873, n2874, n2875, n2876, n2877, n2878,
    n2879, n2880, n2881, n2882, n2883, n2884,
    n2885, n2886, n2887, n2888, n2889, n2890,
    n2891, n2892, n2893, n2894, n2895, n2896,
    n2897, n2898, n2899, n2900, n2901, n2902,
    n2903, n2904, n2905, n2906, n2907, n2908,
    n2909, n2910, n2911, n2912, n2913, n2914,
    n2915, n2916, n2917, n2918, n2919, n2920,
    n2921, n2922, n2923, n2924, n2925, n2926,
    n2927, n2928, n2929, n2930, n2931, n2932,
    n2933, n2934, n2935, n2936, n2938, n2939,
    n2940, n2941, n2942, n2943, n2944, n2945,
    n2946, n2947, n2948, n2949, n2950, n2951,
    n2952, n2953, n2954, n2955, n2956, n2957,
    n2958, n2959, n2960, n2961, n2962, n2963,
    n2964, n2965, n2966, n2967, n2968, n2969,
    n2970, n2971, n2972, n2973, n2974, n2975,
    n2976, n2977, n2978, n2979, n2980, n2981,
    n2982, n2983, n2984, n2985, n2986, n2987,
    n2988, n2989, n2990, n2991, n2992, n2993,
    n2994, n2995, n2996, n2997, n2998, n2999,
    n3000, n3001, n3002, n3003, n3004, n3005,
    n3006, n3007, n3008, n3009, n3010, n3011,
    n3012, n3013, n3014, n3015, n3016, n3017,
    n3018, n3019, n3020, n3021, n3022, n3023,
    n3024, n3025, n3026, n3027, n3028, n3029,
    n3030, n3031, n3032, n3033, n3034, n3035,
    n3036, n3037, n3038, n3039, n3040, n3041,
    n3042, n3043, n3044, n3045, n3046, n3047,
    n3048, n3049, n3050, n3051, n3052, n3053,
    n3054, n3055, n3056, n3057, n3058, n3059,
    n3060, n3061, n3062, n3063, n3064, n3065,
    n3066, n3067, n3068, n3069, n3070, n3071,
    n3072, n3073, n3074, n3075, n3076, n3077,
    n3078, n3079, n3080, n3081, n3082, n3083,
    n3084, n3085, n3086, n3087, n3088, n3089,
    n3090, n3091, n3092, n3093, n3094, n3095,
    n3096, n3097, n3098, n3099, n3100, n3101,
    n3102, n3103, n3104, n3105, n3106, n3107,
    n3108, n3109, n3110, n3111, n3113, n3114,
    n3115, n3116, n3117, n3118, n3119, n3120,
    n3121, n3122, n3123, n3124, n3125, n3126,
    n3127, n3128, n3129, n3130, n3131, n3132,
    n3133, n3134, n3135, n3136, n3137, n3138,
    n3139, n3140, n3141, n3142, n3143, n3144,
    n3145, n3146, n3147, n3148, n3149, n3150,
    n3151, n3152, n3153, n3154, n3155, n3156,
    n3157, n3158, n3159, n3160, n3161, n3162,
    n3163, n3164, n3165, n3166, n3167, n3168,
    n3169, n3170, n3171, n3172, n3173, n3174,
    n3175, n3176, n3177, n3178, n3179, n3180,
    n3181, n3182, n3183, n3184, n3185, n3186,
    n3187, n3188, n3189, n3190, n3191, n3192,
    n3193, n3194, n3195, n3196, n3197, n3198,
    n3199, n3200, n3201, n3202, n3203, n3204,
    n3205, n3206, n3207, n3208, n3209, n3210,
    n3211, n3212, n3213, n3214, n3215, n3216,
    n3217, n3218, n3219, n3220, n3221, n3222,
    n3223, n3224, n3225, n3226, n3227, n3228,
    n3229, n3230, n3231, n3232, n3233, n3234,
    n3235, n3236, n3237, n3238, n3239, n3240,
    n3241, n3242, n3243, n3244, n3245, n3246,
    n3247, n3248, n3249, n3250, n3251, n3252,
    n3253, n3254, n3255, n3256, n3257, n3258,
    n3259, n3260, n3261, n3262, n3263, n3264,
    n3265, n3266, n3267, n3268, n3269, n3270,
    n3271, n3272, n3273, n3274, n3275, n3276,
    n3277, n3278, n3279, n3280, n3281, n3282,
    n3283, n3284, n3285, n3286, n3287, n3288,
    n3289, n3290, n3291, n3292, n3294, n3295,
    n3296, n3297, n3298, n3299, n3300, n3301,
    n3302, n3303, n3304, n3305, n3306, n3307,
    n3308, n3309, n3310, n3311, n3312, n3313,
    n3314, n3315, n3316, n3317, n3318, n3319,
    n3320, n3321, n3322, n3323, n3324, n3325,
    n3326, n3327, n3328, n3329, n3330, n3331,
    n3332, n3333, n3334, n3335, n3336, n3337,
    n3338, n3339, n3340, n3341, n3342, n3343,
    n3344, n3345, n3346, n3347, n3348, n3349,
    n3350, n3351, n3352, n3353, n3354, n3355,
    n3356, n3357, n3358, n3359, n3360, n3361,
    n3362, n3363, n3364, n3365, n3366, n3367,
    n3368, n3369, n3370, n3371, n3372, n3373,
    n3374, n3375, n3376, n3377, n3378, n3379,
    n3380, n3381, n3382, n3383, n3384, n3385,
    n3386, n3387, n3388, n3389, n3390, n3391,
    n3392, n3393, n3394, n3395, n3396, n3397,
    n3398, n3399, n3400, n3401, n3402, n3403,
    n3404, n3405, n3406, n3407, n3408, n3409,
    n3410, n3411, n3412, n3413, n3414, n3415,
    n3416, n3417, n3418, n3419, n3420, n3421,
    n3422, n3423, n3424, n3425, n3426, n3427,
    n3428, n3429, n3430, n3431, n3432, n3433,
    n3434, n3435, n3436, n3437, n3438, n3439,
    n3440, n3441, n3442, n3443, n3444, n3445,
    n3446, n3447, n3448, n3449, n3450, n3451,
    n3452, n3453, n3454, n3455, n3456, n3457,
    n3458, n3459, n3460, n3461, n3462, n3463,
    n3464, n3465, n3466, n3467, n3468, n3469,
    n3470, n3471, n3472, n3473, n3474, n3475,
    n3476, n3477, n3478, n3479, n3480, n3481,
    n3482, n3483, n3484, n3485, n3486, n3487,
    n3489, n3490, n3491, n3492, n3493, n3494,
    n3495, n3496, n3497, n3498, n3499, n3500,
    n3501, n3502, n3503, n3504, n3505, n3506,
    n3507, n3508, n3509, n3510, n3511, n3512,
    n3513, n3514, n3515, n3516, n3517, n3518,
    n3519, n3520, n3521, n3522, n3523, n3524,
    n3525, n3526, n3527, n3528, n3529, n3530,
    n3531, n3532, n3533, n3534, n3535, n3536,
    n3537, n3538, n3539, n3540, n3541, n3542,
    n3543, n3544, n3545, n3546, n3547, n3548,
    n3549, n3550, n3551, n3552, n3553, n3554,
    n3555, n3556, n3557, n3558, n3559, n3560,
    n3561, n3562, n3563, n3564, n3565, n3566,
    n3567, n3568, n3569, n3570, n3571, n3572,
    n3573, n3574, n3575, n3576, n3577, n3578,
    n3579, n3580, n3581, n3582, n3583, n3584,
    n3585, n3586, n3587, n3588, n3589, n3590,
    n3591, n3592, n3593, n3594, n3595, n3596,
    n3597, n3598, n3599, n3600, n3601, n3602,
    n3603, n3604, n3605, n3606, n3607, n3608,
    n3609, n3610, n3611, n3612, n3613, n3614,
    n3615, n3616, n3617, n3618, n3619, n3620,
    n3621, n3622, n3623, n3624, n3625, n3626,
    n3627, n3628, n3629, n3630, n3631, n3632,
    n3633, n3634, n3635, n3636, n3637, n3638,
    n3639, n3640, n3641, n3642, n3643, n3644,
    n3645, n3646, n3647, n3648, n3649, n3650,
    n3651, n3652, n3653, n3654, n3655, n3656,
    n3657, n3658, n3659, n3660, n3661, n3662,
    n3663, n3664, n3665, n3666, n3667, n3668,
    n3669, n3670, n3671, n3672, n3673, n3674,
    n3675, n3676, n3677, n3678, n3679, n3681,
    n3682, n3683, n3684, n3685, n3686, n3687,
    n3688, n3689, n3690, n3691, n3692, n3693,
    n3694, n3695, n3696, n3697, n3698, n3699,
    n3700, n3701, n3702, n3703, n3704, n3705,
    n3706, n3707, n3708, n3709, n3710, n3711,
    n3712, n3713, n3714, n3715, n3716, n3717,
    n3718, n3719, n3720, n3721, n3722, n3723,
    n3724, n3725, n3726, n3727, n3728, n3729,
    n3730, n3731, n3732, n3733, n3734, n3735,
    n3736, n3737, n3738, n3739, n3740, n3741,
    n3742, n3743, n3744, n3745, n3746, n3747,
    n3748, n3749, n3750, n3751, n3752, n3753,
    n3754, n3755, n3756, n3757, n3758, n3759,
    n3760, n3761, n3762, n3763, n3764, n3765,
    n3766, n3767, n3768, n3769, n3770, n3771,
    n3772, n3773, n3774, n3775, n3776, n3777,
    n3778, n3779, n3780, n3781, n3782, n3783,
    n3784, n3785, n3786, n3787, n3788, n3789,
    n3790, n3791, n3792, n3793, n3794, n3795,
    n3796, n3797, n3798, n3799, n3800, n3801,
    n3802, n3803, n3804, n3805, n3806, n3807,
    n3808, n3809, n3810, n3811, n3812, n3813,
    n3814, n3815, n3816, n3817, n3818, n3819,
    n3820, n3821, n3822, n3823, n3824, n3825,
    n3826, n3827, n3828, n3829, n3830, n3831,
    n3832, n3833, n3834, n3835, n3836, n3837,
    n3838, n3839, n3840, n3841, n3842, n3843,
    n3844, n3845, n3846, n3847, n3848, n3849,
    n3850, n3851, n3852, n3853, n3854, n3855,
    n3856, n3857, n3858, n3859, n3860, n3861,
    n3862, n3863, n3864, n3865, n3866, n3867,
    n3868, n3869, n3870, n3871, n3872, n3873,
    n3874, n3875, n3876, n3877, n3879, n3880,
    n3881, n3882, n3883, n3884, n3885, n3886,
    n3887, n3888, n3889, n3890, n3891, n3892,
    n3893, n3894, n3895, n3896, n3897, n3898,
    n3899, n3900, n3901, n3902, n3903, n3904,
    n3905, n3906, n3907, n3908, n3909, n3910,
    n3911, n3912, n3913, n3914, n3915, n3916,
    n3917, n3918, n3919, n3920, n3921, n3922,
    n3923, n3924, n3925, n3926, n3927, n3928,
    n3929, n3930, n3931, n3932, n3933, n3934,
    n3935, n3936, n3937, n3938, n3939, n3940,
    n3941, n3942, n3943, n3944, n3945, n3946,
    n3947, n3948, n3949, n3950, n3951, n3952,
    n3953, n3954, n3955, n3956, n3957, n3958,
    n3959, n3960, n3961, n3962, n3963, n3964,
    n3965, n3966, n3967, n3968, n3969, n3970,
    n3971, n3972, n3973, n3974, n3975, n3976,
    n3977, n3978, n3979, n3980, n3981, n3982,
    n3983, n3984, n3985, n3986, n3987, n3988,
    n3989, n3990, n3991, n3992, n3993, n3994,
    n3995, n3996, n3997, n3998, n3999, n4000,
    n4001, n4002, n4003, n4004, n4005, n4006,
    n4007, n4008, n4009, n4010, n4011, n4012,
    n4013, n4014, n4015, n4016, n4017, n4018,
    n4019, n4020, n4021, n4022, n4023, n4024,
    n4025, n4026, n4027, n4028, n4029, n4030,
    n4031, n4032, n4033, n4034, n4035, n4036,
    n4037, n4038, n4039, n4040, n4041, n4042,
    n4043, n4044, n4045, n4046, n4047, n4048,
    n4049, n4050, n4051, n4052, n4053, n4054,
    n4055, n4056, n4057, n4058, n4059, n4060,
    n4061, n4062, n4063, n4064, n4065, n4066,
    n4067, n4068, n4069, n4070, n4071, n4072,
    n4073, n4074, n4075, n4076, n4077, n4078,
    n4079, n4080, n4081, n4082, n4083, n4084,
    n4085, n4086, n4087, n4088, n4089, n4091,
    n4092, n4093, n4094, n4095, n4096, n4097,
    n4098, n4099, n4100, n4101, n4102, n4103,
    n4104, n4105, n4106, n4107, n4108, n4109,
    n4110, n4111, n4112, n4113, n4114, n4115,
    n4116, n4117, n4118, n4119, n4120, n4121,
    n4122, n4123, n4124, n4125, n4126, n4127,
    n4128, n4129, n4130, n4131, n4132, n4133,
    n4134, n4135, n4136, n4137, n4138, n4139,
    n4140, n4141, n4142, n4143, n4144, n4145,
    n4146, n4147, n4148, n4149, n4150, n4151,
    n4152, n4153, n4154, n4155, n4156, n4157,
    n4158, n4159, n4160, n4161, n4162, n4163,
    n4164, n4165, n4166, n4167, n4168, n4169,
    n4170, n4171, n4172, n4173, n4174, n4175,
    n4176, n4177, n4178, n4179, n4180, n4181,
    n4182, n4183, n4184, n4185, n4186, n4187,
    n4188, n4189, n4190, n4191, n4192, n4193,
    n4194, n4195, n4196, n4197, n4198, n4199,
    n4200, n4201, n4202, n4203, n4204, n4205,
    n4206, n4207, n4208, n4209, n4210, n4211,
    n4212, n4213, n4214, n4215, n4216, n4217,
    n4218, n4219, n4220, n4221, n4222, n4223,
    n4224, n4225, n4226, n4227, n4228, n4229,
    n4230, n4231, n4232, n4233, n4234, n4235,
    n4236, n4237, n4238, n4239, n4240, n4241,
    n4242, n4243, n4244, n4245, n4246, n4247,
    n4248, n4249, n4250, n4251, n4252, n4253,
    n4254, n4255, n4256, n4257, n4258, n4259,
    n4260, n4261, n4262, n4263, n4264, n4265,
    n4266, n4267, n4268, n4269, n4270, n4271,
    n4272, n4273, n4274, n4275, n4276, n4277,
    n4278, n4279, n4280, n4281, n4282, n4283,
    n4284, n4285, n4286, n4287, n4288, n4289,
    n4290, n4291, n4292, n4293, n4294, n4295,
    n4296, n4297, n4298, n4300, n4301, n4302,
    n4303, n4304, n4305, n4306, n4307, n4308,
    n4309, n4310, n4311, n4312, n4313, n4314,
    n4315, n4316, n4317, n4318, n4319, n4320,
    n4321, n4322, n4323, n4324, n4325, n4326,
    n4327, n4328, n4329, n4330, n4331, n4332,
    n4333, n4334, n4335, n4336, n4337, n4338,
    n4339, n4340, n4341, n4342, n4343, n4344,
    n4345, n4346, n4347, n4348, n4349, n4350,
    n4351, n4352, n4353, n4354, n4355, n4356,
    n4357, n4358, n4359, n4360, n4361, n4362,
    n4363, n4364, n4365, n4366, n4367, n4368,
    n4369, n4370, n4371, n4372, n4373, n4374,
    n4375, n4376, n4377, n4378, n4379, n4380,
    n4381, n4382, n4383, n4384, n4385, n4386,
    n4387, n4388, n4389, n4390, n4391, n4392,
    n4393, n4394, n4395, n4396, n4397, n4398,
    n4399, n4400, n4401, n4402, n4403, n4404,
    n4405, n4406, n4407, n4408, n4409, n4410,
    n4411, n4412, n4413, n4414, n4415, n4416,
    n4417, n4418, n4419, n4420, n4421, n4422,
    n4423, n4424, n4425, n4426, n4427, n4428,
    n4429, n4430, n4431, n4432, n4433, n4434,
    n4435, n4436, n4437, n4438, n4439, n4440,
    n4441, n4442, n4443, n4444, n4445, n4446,
    n4447, n4448, n4449, n4450, n4451, n4452,
    n4453, n4454, n4455, n4456, n4457, n4458,
    n4459, n4460, n4461, n4462, n4463, n4464,
    n4465, n4466, n4467, n4468, n4469, n4470,
    n4471, n4472, n4473, n4474, n4475, n4476,
    n4477, n4478, n4479, n4480, n4481, n4482,
    n4483, n4484, n4485, n4486, n4487, n4488,
    n4489, n4490, n4491, n4492, n4493, n4494,
    n4495, n4496, n4497, n4498, n4499, n4500,
    n4501, n4502, n4503, n4504, n4505, n4506,
    n4507, n4508, n4509, n4510, n4511, n4512,
    n4513, n4515, n4516, n4517, n4518, n4519,
    n4520, n4521, n4522, n4523, n4524, n4525,
    n4526, n4527, n4528, n4529, n4530, n4531,
    n4532, n4533, n4534, n4535, n4536, n4537,
    n4538, n4539, n4540, n4541, n4542, n4543,
    n4544, n4545, n4546, n4547, n4548, n4549,
    n4550, n4551, n4552, n4553, n4554, n4555,
    n4556, n4557, n4558, n4559, n4560, n4561,
    n4562, n4563, n4564, n4565, n4566, n4567,
    n4568, n4569, n4570, n4571, n4572, n4573,
    n4574, n4575, n4576, n4577, n4578, n4579,
    n4580, n4581, n4582, n4583, n4584, n4585,
    n4586, n4587, n4588, n4589, n4590, n4591,
    n4592, n4593, n4594, n4595, n4596, n4597,
    n4598, n4599, n4600, n4601, n4602, n4603,
    n4604, n4605, n4606, n4607, n4608, n4609,
    n4610, n4611, n4612, n4613, n4614, n4615,
    n4616, n4617, n4618, n4619, n4620, n4621,
    n4622, n4623, n4624, n4625, n4626, n4627,
    n4628, n4629, n4630, n4631, n4632, n4633,
    n4634, n4635, n4636, n4637, n4638, n4639,
    n4640, n4641, n4642, n4643, n4644, n4645,
    n4646, n4647, n4648, n4649, n4650, n4651,
    n4652, n4653, n4654, n4655, n4656, n4657,
    n4658, n4659, n4660, n4661, n4662, n4663,
    n4664, n4665, n4666, n4667, n4668, n4669,
    n4670, n4671, n4672, n4673, n4674, n4675,
    n4676, n4677, n4678, n4679, n4680, n4681,
    n4682, n4683, n4684, n4685, n4686, n4687,
    n4688, n4689, n4690, n4691, n4692, n4693,
    n4694, n4695, n4696, n4697, n4698, n4699,
    n4700, n4701, n4702, n4703, n4704, n4705,
    n4706, n4707, n4708, n4709, n4710, n4711,
    n4712, n4713, n4714, n4715, n4716, n4717,
    n4718, n4719, n4720, n4721, n4722, n4723,
    n4724, n4725, n4726, n4727, n4728, n4729,
    n4730, n4731, n4732, n4733, n4734, n4735,
    n4736, n4737, n4738, n4739, n4740, n4741,
    n4742, n4744, n4745, n4746, n4747, n4748,
    n4749, n4750, n4751, n4752, n4753, n4754,
    n4755, n4756, n4757, n4758, n4759, n4760,
    n4761, n4762, n4763, n4764, n4765, n4766,
    n4767, n4768, n4769, n4770, n4771, n4772,
    n4773, n4774, n4775, n4776, n4777, n4778,
    n4779, n4780, n4781, n4782, n4783, n4784,
    n4785, n4786, n4787, n4788, n4789, n4790,
    n4791, n4792, n4793, n4794, n4795, n4796,
    n4797, n4798, n4799, n4800, n4801, n4802,
    n4803, n4804, n4805, n4806, n4807, n4808,
    n4809, n4810, n4811, n4812, n4813, n4814,
    n4815, n4816, n4817, n4818, n4819, n4820,
    n4821, n4822, n4823, n4824, n4825, n4826,
    n4827, n4828, n4829, n4830, n4831, n4832,
    n4833, n4834, n4835, n4836, n4837, n4838,
    n4839, n4840, n4841, n4842, n4843, n4844,
    n4845, n4846, n4847, n4848, n4849, n4850,
    n4851, n4852, n4853, n4854, n4855, n4856,
    n4857, n4858, n4859, n4860, n4861, n4862,
    n4863, n4864, n4865, n4866, n4867, n4868,
    n4869, n4870, n4871, n4872, n4873, n4874,
    n4875, n4876, n4877, n4878, n4879, n4880,
    n4881, n4882, n4883, n4884, n4885, n4886,
    n4887, n4888, n4889, n4890, n4891, n4892,
    n4893, n4894, n4895, n4896, n4897, n4898,
    n4899, n4900, n4901, n4902, n4903, n4904,
    n4905, n4906, n4907, n4908, n4909, n4910,
    n4911, n4912, n4913, n4914, n4915, n4916,
    n4917, n4918, n4919, n4920, n4921, n4922,
    n4923, n4924, n4925, n4926, n4927, n4928,
    n4929, n4930, n4931, n4932, n4933, n4934,
    n4935, n4936, n4937, n4938, n4939, n4940,
    n4941, n4942, n4943, n4944, n4945, n4946,
    n4947, n4948, n4949, n4950, n4951, n4952,
    n4953, n4954, n4955, n4956, n4957, n4958,
    n4959, n4960, n4961, n4962, n4963, n4964,
    n4965, n4966, n4967, n4968, n4970, n4971,
    n4972, n4973, n4974, n4975, n4976, n4977,
    n4978, n4979, n4980, n4981, n4982, n4983,
    n4984, n4985, n4986, n4987, n4988, n4989,
    n4990, n4991, n4992, n4993, n4994, n4995,
    n4996, n4997, n4998, n4999, n5000, n5001,
    n5002, n5003, n5004, n5005, n5006, n5007,
    n5008, n5009, n5010, n5011, n5012, n5013,
    n5014, n5015, n5016, n5017, n5018, n5019,
    n5020, n5021, n5022, n5023, n5024, n5025,
    n5026, n5027, n5028, n5029, n5030, n5031,
    n5032, n5033, n5034, n5035, n5036, n5037,
    n5038, n5039, n5040, n5041, n5042, n5043,
    n5044, n5045, n5046, n5047, n5048, n5049,
    n5050, n5051, n5052, n5053, n5054, n5055,
    n5056, n5057, n5058, n5059, n5060, n5061,
    n5062, n5063, n5064, n5065, n5066, n5067,
    n5068, n5069, n5070, n5071, n5072, n5073,
    n5074, n5075, n5076, n5077, n5078, n5079,
    n5080, n5081, n5082, n5083, n5084, n5085,
    n5086, n5087, n5088, n5089, n5090, n5091,
    n5092, n5093, n5094, n5095, n5096, n5097,
    n5098, n5099, n5100, n5101, n5102, n5103,
    n5104, n5105, n5106, n5107, n5108, n5109,
    n5110, n5111, n5112, n5113, n5114, n5115,
    n5116, n5117, n5118, n5119, n5120, n5121,
    n5122, n5123, n5124, n5125, n5126, n5127,
    n5128, n5129, n5130, n5131, n5132, n5133,
    n5134, n5135, n5136, n5137, n5138, n5139,
    n5140, n5141, n5142, n5143, n5144, n5145,
    n5146, n5147, n5148, n5149, n5150, n5151,
    n5152, n5153, n5154, n5155, n5156, n5157,
    n5158, n5159, n5160, n5161, n5162, n5163,
    n5164, n5165, n5166, n5167, n5168, n5169,
    n5170, n5171, n5172, n5173, n5174, n5175,
    n5176, n5177, n5178, n5179, n5180, n5181,
    n5182, n5183, n5184, n5185, n5186, n5187,
    n5188, n5189, n5190, n5191, n5192, n5193,
    n5194, n5195, n5196, n5197, n5198, n5199,
    n5200, n5202, n5203, n5204, n5205, n5206,
    n5207, n5208, n5209, n5210, n5211, n5212,
    n5213, n5214, n5215, n5216, n5217, n5218,
    n5219, n5220, n5221, n5222, n5223, n5224,
    n5225, n5226, n5227, n5228, n5229, n5230,
    n5231, n5232, n5233, n5234, n5235, n5236,
    n5237, n5238, n5239, n5240, n5241, n5242,
    n5243, n5244, n5245, n5246, n5247, n5248,
    n5249, n5250, n5251, n5252, n5253, n5254,
    n5255, n5256, n5257, n5258, n5259, n5260,
    n5261, n5262, n5263, n5264, n5265, n5266,
    n5267, n5268, n5269, n5270, n5271, n5272,
    n5273, n5274, n5275, n5276, n5277, n5278,
    n5279, n5280, n5281, n5282, n5283, n5284,
    n5285, n5286, n5287, n5288, n5289, n5290,
    n5291, n5292, n5293, n5294, n5295, n5296,
    n5297, n5298, n5299, n5300, n5301, n5302,
    n5303, n5304, n5305, n5306, n5307, n5308,
    n5309, n5310, n5311, n5312, n5313, n5314,
    n5315, n5316, n5317, n5318, n5319, n5320,
    n5321, n5322, n5323, n5324, n5325, n5326,
    n5327, n5328, n5329, n5330, n5331, n5332,
    n5333, n5334, n5335, n5336, n5337, n5338,
    n5339, n5340, n5341, n5342, n5343, n5344,
    n5345, n5346, n5347, n5348, n5349, n5350,
    n5351, n5352, n5353, n5354, n5355, n5356,
    n5357, n5358, n5359, n5360, n5361, n5362,
    n5363, n5364, n5365, n5366, n5367, n5368,
    n5369, n5370, n5371, n5372, n5373, n5374,
    n5375, n5376, n5377, n5378, n5379, n5380,
    n5381, n5382, n5383, n5384, n5385, n5386,
    n5387, n5388, n5389, n5390, n5391, n5392,
    n5393, n5394, n5395, n5396, n5397, n5398,
    n5399, n5400, n5401, n5402, n5403, n5404,
    n5405, n5406, n5407, n5408, n5409, n5410,
    n5411, n5412, n5413, n5414, n5415, n5416,
    n5417, n5418, n5419, n5420, n5421, n5422,
    n5423, n5424, n5425, n5426, n5427, n5428,
    n5429, n5430, n5431, n5432, n5433, n5434,
    n5435, n5436, n5437, n5438, n5439, n5440,
    n5441, n5442, n5443, n5444, n5445, n5446,
    n5448, n5449, n5450, n5451, n5452, n5453,
    n5454, n5455, n5456, n5457, n5458, n5459,
    n5460, n5461, n5462, n5463, n5464, n5465,
    n5466, n5467, n5468, n5469, n5470, n5471,
    n5472, n5473, n5474, n5475, n5476, n5477,
    n5478, n5479, n5480, n5481, n5482, n5483,
    n5484, n5485, n5486, n5487, n5488, n5489,
    n5490, n5491, n5492, n5493, n5494, n5495,
    n5496, n5497, n5498, n5499, n5500, n5501,
    n5502, n5503, n5504, n5505, n5506, n5507,
    n5508, n5509, n5510, n5511, n5512, n5513,
    n5514, n5515, n5516, n5517, n5518, n5519,
    n5520, n5521, n5522, n5523, n5524, n5525,
    n5526, n5527, n5528, n5529, n5530, n5531,
    n5532, n5533, n5534, n5535, n5536, n5537,
    n5538, n5539, n5540, n5541, n5542, n5543,
    n5544, n5545, n5546, n5547, n5548, n5549,
    n5550, n5551, n5552, n5553, n5554, n5555,
    n5556, n5557, n5558, n5559, n5560, n5561,
    n5562, n5563, n5564, n5565, n5566, n5567,
    n5568, n5569, n5570, n5571, n5572, n5573,
    n5574, n5575, n5576, n5577, n5578, n5579,
    n5580, n5581, n5582, n5583, n5584, n5585,
    n5586, n5587, n5588, n5589, n5590, n5591,
    n5592, n5593, n5594, n5595, n5596, n5597,
    n5598, n5599, n5600, n5601, n5602, n5603,
    n5604, n5605, n5606, n5607, n5608, n5609,
    n5610, n5611, n5612, n5613, n5614, n5615,
    n5616, n5617, n5618, n5619, n5620, n5621,
    n5622, n5623, n5624, n5625, n5626, n5627,
    n5628, n5629, n5630, n5631, n5632, n5633,
    n5634, n5635, n5636, n5637, n5638, n5639,
    n5640, n5641, n5642, n5643, n5644, n5645,
    n5646, n5647, n5648, n5649, n5650, n5651,
    n5652, n5653, n5654, n5655, n5656, n5657,
    n5658, n5659, n5660, n5661, n5662, n5663,
    n5664, n5665, n5666, n5667, n5668, n5669,
    n5670, n5671, n5672, n5673, n5674, n5675,
    n5676, n5677, n5678, n5679, n5680, n5681,
    n5682, n5683, n5684, n5685, n5686, n5687,
    n5688, n5689, n5691, n5692, n5693, n5694,
    n5695, n5696, n5697, n5698, n5699, n5700,
    n5701, n5702, n5703, n5704, n5705, n5706,
    n5707, n5708, n5709, n5710, n5711, n5712,
    n5713, n5714, n5715, n5716, n5717, n5718,
    n5719, n5720, n5721, n5722, n5723, n5724,
    n5725, n5726, n5727, n5728, n5729, n5730,
    n5731, n5732, n5733, n5734, n5735, n5736,
    n5737, n5738, n5739, n5740, n5741, n5742,
    n5743, n5744, n5745, n5746, n5747, n5748,
    n5749, n5750, n5751, n5752, n5753, n5754,
    n5755, n5756, n5757, n5758, n5759, n5760,
    n5761, n5762, n5763, n5764, n5765, n5766,
    n5767, n5768, n5769, n5770, n5771, n5772,
    n5773, n5774, n5775, n5776, n5777, n5778,
    n5779, n5780, n5781, n5782, n5783, n5784,
    n5785, n5786, n5787, n5788, n5789, n5790,
    n5791, n5792, n5793, n5794, n5795, n5796,
    n5797, n5798, n5799, n5800, n5801, n5802,
    n5803, n5804, n5805, n5806, n5807, n5808,
    n5809, n5810, n5811, n5812, n5813, n5814,
    n5815, n5816, n5817, n5818, n5819, n5820,
    n5821, n5822, n5823, n5824, n5825, n5826,
    n5827, n5828, n5829, n5830, n5831, n5832,
    n5833, n5834, n5835, n5836, n5837, n5838,
    n5839, n5840, n5841, n5842, n5843, n5844,
    n5845, n5846, n5847, n5848, n5849, n5850,
    n5851, n5852, n5853, n5854, n5855, n5856,
    n5857, n5858, n5859, n5860, n5861, n5862,
    n5863, n5864, n5865, n5866, n5867, n5868,
    n5869, n5870, n5871, n5872, n5873, n5874,
    n5875, n5876, n5877, n5878, n5879, n5880,
    n5881, n5882, n5883, n5884, n5885, n5886,
    n5887, n5888, n5889, n5890, n5891, n5892,
    n5893, n5894, n5895, n5896, n5897, n5898,
    n5899, n5900, n5901, n5902, n5903, n5904,
    n5905, n5906, n5907, n5908, n5909, n5910,
    n5911, n5912, n5913, n5914, n5915, n5916,
    n5917, n5918, n5919, n5920, n5921, n5922,
    n5923, n5924, n5925, n5926, n5927, n5928,
    n5929, n5930, n5931, n5932, n5933, n5934,
    n5935, n5936, n5937, n5938, n5940, n5941,
    n5942, n5943, n5944, n5945, n5946, n5947,
    n5948, n5949, n5950, n5951, n5952, n5953,
    n5954, n5955, n5956, n5957, n5958, n5959,
    n5960, n5961, n5962, n5963, n5964, n5965,
    n5966, n5967, n5968, n5969, n5970, n5971,
    n5972, n5973, n5974, n5975, n5976, n5977,
    n5978, n5979, n5980, n5981, n5982, n5983,
    n5984, n5985, n5986, n5987, n5988, n5989,
    n5990, n5991, n5992, n5993, n5994, n5995,
    n5996, n5997, n5998, n5999, n6000, n6001,
    n6002, n6003, n6004, n6005, n6006, n6007,
    n6008, n6009, n6010, n6011, n6012, n6013,
    n6014, n6015, n6016, n6017, n6018, n6019,
    n6020, n6021, n6022, n6023, n6024, n6025,
    n6026, n6027, n6028, n6029, n6030, n6031,
    n6032, n6033, n6034, n6035, n6036, n6037,
    n6038, n6039, n6040, n6041, n6042, n6043,
    n6044, n6045, n6046, n6047, n6048, n6049,
    n6050, n6051, n6052, n6053, n6054, n6055,
    n6056, n6057, n6058, n6059, n6060, n6061,
    n6062, n6063, n6064, n6065, n6066, n6067,
    n6068, n6069, n6070, n6071, n6072, n6073,
    n6074, n6075, n6076, n6077, n6078, n6079,
    n6080, n6081, n6082, n6083, n6084, n6085,
    n6086, n6087, n6088, n6089, n6090, n6091,
    n6092, n6093, n6094, n6095, n6096, n6097,
    n6098, n6099, n6100, n6101, n6102, n6103,
    n6104, n6105, n6106, n6107, n6108, n6109,
    n6110, n6111, n6112, n6113, n6114, n6115,
    n6116, n6117, n6118, n6119, n6120, n6121,
    n6122, n6123, n6124, n6125, n6126, n6127,
    n6128, n6129, n6130, n6131, n6132, n6133,
    n6134, n6135, n6136, n6137, n6138, n6139,
    n6140, n6141, n6142, n6143, n6144, n6145,
    n6146, n6147, n6148, n6149, n6150, n6151,
    n6152, n6153, n6154, n6155, n6156, n6157,
    n6158, n6159, n6160, n6161, n6162, n6163,
    n6164, n6165, n6166, n6167, n6168, n6169,
    n6170, n6171, n6172, n6173, n6174, n6175,
    n6176, n6177, n6178, n6179, n6180, n6181,
    n6182, n6183, n6184, n6185, n6186, n6187,
    n6188, n6189, n6190, n6191, n6192, n6193,
    n6194, n6195, n6196, n6197, n6198, n6199,
    n6200, n6201, n6203, n6204, n6205, n6206,
    n6207, n6208, n6209, n6210, n6211, n6212,
    n6213, n6214, n6215, n6216, n6217, n6218,
    n6219, n6220, n6221, n6222, n6223, n6224,
    n6225, n6226, n6227, n6228, n6229, n6230,
    n6231, n6232, n6233, n6234, n6235, n6236,
    n6237, n6238, n6239, n6240, n6241, n6242,
    n6243, n6244, n6245, n6246, n6247, n6248,
    n6249, n6250, n6251, n6252, n6253, n6254,
    n6255, n6256, n6257, n6258, n6259, n6260,
    n6261, n6262, n6263, n6264, n6265, n6266,
    n6267, n6268, n6269, n6270, n6271, n6272,
    n6273, n6274, n6275, n6276, n6277, n6278,
    n6279, n6280, n6281, n6282, n6283, n6284,
    n6285, n6286, n6287, n6288, n6289, n6290,
    n6291, n6292, n6293, n6294, n6295, n6296,
    n6297, n6298, n6299, n6300, n6301, n6302,
    n6303, n6304, n6305, n6306, n6307, n6308,
    n6309, n6310, n6311, n6312, n6313, n6314,
    n6315, n6316, n6317, n6318, n6319, n6320,
    n6321, n6322, n6323, n6324, n6325, n6326,
    n6327, n6328, n6329, n6330, n6331, n6332,
    n6333, n6334, n6335, n6336, n6337, n6338,
    n6339, n6340, n6341, n6342, n6343, n6344,
    n6345, n6346, n6347, n6348, n6349, n6350,
    n6351, n6352, n6353, n6354, n6355, n6356,
    n6357, n6358, n6359, n6360, n6361, n6362,
    n6363, n6364, n6365, n6366, n6367, n6368,
    n6369, n6370, n6371, n6372, n6373, n6374,
    n6375, n6376, n6377, n6378, n6379, n6380,
    n6381, n6382, n6383, n6384, n6385, n6386,
    n6387, n6388, n6389, n6390, n6391, n6392,
    n6393, n6394, n6395, n6396, n6397, n6398,
    n6399, n6400, n6401, n6402, n6403, n6404,
    n6405, n6406, n6407, n6408, n6409, n6410,
    n6411, n6412, n6413, n6414, n6415, n6416,
    n6417, n6418, n6419, n6420, n6421, n6422,
    n6423, n6424, n6425, n6426, n6427, n6428,
    n6429, n6430, n6431, n6432, n6433, n6434,
    n6435, n6436, n6437, n6438, n6439, n6440,
    n6441, n6442, n6443, n6444, n6445, n6446,
    n6447, n6448, n6449, n6450, n6451, n6452,
    n6453, n6454, n6455, n6456, n6457, n6458,
    n6459, n6460, n6461, n6463, n6464, n6465,
    n6466, n6467, n6468, n6469, n6470, n6471,
    n6472, n6473, n6474, n6475, n6476, n6477,
    n6478, n6479, n6480, n6481, n6482, n6483,
    n6484, n6485, n6486, n6487, n6488, n6489,
    n6490, n6491, n6492, n6493, n6494, n6495,
    n6496, n6497, n6498, n6499, n6500, n6501,
    n6502, n6503, n6504, n6505, n6506, n6507,
    n6508, n6509, n6510, n6511, n6512, n6513,
    n6514, n6515, n6516, n6517, n6518, n6519,
    n6520, n6521, n6522, n6523, n6524, n6525,
    n6526, n6527, n6528, n6529, n6530, n6531,
    n6532, n6533, n6534, n6535, n6536, n6537,
    n6538, n6539, n6540, n6541, n6542, n6543,
    n6544, n6545, n6546, n6547, n6548, n6549,
    n6550, n6551, n6552, n6553, n6554, n6555,
    n6556, n6557, n6558, n6559, n6560, n6561,
    n6562, n6563, n6564, n6565, n6566, n6567,
    n6568, n6569, n6570, n6571, n6572, n6573,
    n6574, n6575, n6576, n6577, n6578, n6579,
    n6580, n6581, n6582, n6583, n6584, n6585,
    n6586, n6587, n6588, n6589, n6590, n6591,
    n6592, n6593, n6594, n6595, n6596, n6597,
    n6598, n6599, n6600, n6601, n6602, n6603,
    n6604, n6605, n6606, n6607, n6608, n6609,
    n6610, n6611, n6612, n6613, n6614, n6615,
    n6616, n6617, n6618, n6619, n6620, n6621,
    n6622, n6623, n6624, n6625, n6626, n6627,
    n6628, n6629, n6630, n6631, n6632, n6633,
    n6634, n6635, n6636, n6637, n6638, n6639,
    n6640, n6641, n6642, n6643, n6644, n6645,
    n6646, n6647, n6648, n6649, n6650, n6651,
    n6652, n6653, n6654, n6655, n6656, n6657,
    n6658, n6659, n6660, n6661, n6662, n6663,
    n6664, n6665, n6666, n6667, n6668, n6669,
    n6670, n6671, n6672, n6673, n6674, n6675,
    n6676, n6677, n6678, n6679, n6680, n6681,
    n6682, n6683, n6684, n6685, n6686, n6687,
    n6688, n6689, n6690, n6691, n6692, n6693,
    n6694, n6695, n6696, n6697, n6698, n6699,
    n6700, n6701, n6702, n6703, n6704, n6705,
    n6706, n6707, n6708, n6709, n6710, n6711,
    n6712, n6713, n6714, n6715, n6716, n6717,
    n6718, n6719, n6720, n6721, n6722, n6723,
    n6724, n6725, n6726, n6727, n6729, n6730,
    n6731, n6732, n6733, n6734, n6735, n6736,
    n6737, n6738, n6739, n6740, n6741, n6742,
    n6743, n6744, n6745, n6746, n6747, n6748,
    n6749, n6750, n6751, n6752, n6753, n6754,
    n6755, n6756, n6757, n6758, n6759, n6760,
    n6761, n6762, n6763, n6764, n6765, n6766,
    n6767, n6768, n6769, n6770, n6771, n6772,
    n6773, n6774, n6775, n6776, n6777, n6778,
    n6779, n6780, n6781, n6782, n6783, n6784,
    n6785, n6786, n6787, n6788, n6789, n6790,
    n6791, n6792, n6793, n6794, n6795, n6796,
    n6797, n6798, n6799, n6800, n6801, n6802,
    n6803, n6804, n6805, n6806, n6807, n6808,
    n6809, n6810, n6811, n6812, n6813, n6814,
    n6815, n6816, n6817, n6818, n6819, n6820,
    n6821, n6822, n6823, n6824, n6825, n6826,
    n6827, n6828, n6829, n6830, n6831, n6832,
    n6833, n6834, n6835, n6836, n6837, n6838,
    n6839, n6840, n6841, n6842, n6843, n6844,
    n6845, n6846, n6847, n6848, n6849, n6850,
    n6851, n6852, n6853, n6854, n6855, n6856,
    n6857, n6858, n6859, n6860, n6861, n6862,
    n6863, n6864, n6865, n6866, n6867, n6868,
    n6869, n6870, n6871, n6872, n6873, n6874,
    n6875, n6876, n6877, n6878, n6879, n6880,
    n6881, n6882, n6883, n6884, n6885, n6886,
    n6887, n6888, n6889, n6890, n6891, n6892,
    n6893, n6894, n6895, n6896, n6897, n6898,
    n6899, n6900, n6901, n6902, n6903, n6904,
    n6905, n6906, n6907, n6908, n6909, n6910,
    n6911, n6912, n6913, n6914, n6915, n6916,
    n6917, n6918, n6919, n6920, n6921, n6922,
    n6923, n6924, n6925, n6926, n6927, n6928,
    n6929, n6930, n6931, n6932, n6933, n6934,
    n6935, n6936, n6937, n6938, n6939, n6940,
    n6941, n6942, n6943, n6944, n6945, n6946,
    n6947, n6948, n6949, n6950, n6951, n6952,
    n6953, n6954, n6955, n6956, n6957, n6958,
    n6959, n6960, n6961, n6962, n6963, n6964,
    n6965, n6966, n6967, n6968, n6969, n6970,
    n6971, n6972, n6973, n6974, n6975, n6976,
    n6977, n6978, n6979, n6980, n6981, n6982,
    n6983, n6984, n6985, n6986, n6987, n6988,
    n6989, n6990, n6991, n6992, n6993, n6994,
    n6995, n6996, n6997, n6998, n6999, n7000,
    n7001, n7002, n7003, n7004, n7005, n7006,
    n7007, n7009, n7010, n7011, n7012, n7013,
    n7014, n7015, n7016, n7017, n7018, n7019,
    n7020, n7021, n7022, n7023, n7024, n7025,
    n7026, n7027, n7028, n7029, n7030, n7031,
    n7032, n7033, n7034, n7035, n7036, n7037,
    n7038, n7039, n7040, n7041, n7042, n7043,
    n7044, n7045, n7046, n7047, n7048, n7049,
    n7050, n7051, n7052, n7053, n7054, n7055,
    n7056, n7057, n7058, n7059, n7060, n7061,
    n7062, n7063, n7064, n7065, n7066, n7067,
    n7068, n7069, n7070, n7071, n7072, n7073,
    n7074, n7075, n7076, n7077, n7078, n7079,
    n7080, n7081, n7082, n7083, n7084, n7085,
    n7086, n7087, n7088, n7089, n7090, n7091,
    n7092, n7093, n7094, n7095, n7096, n7097,
    n7098, n7099, n7100, n7101, n7102, n7103,
    n7104, n7105, n7106, n7107, n7108, n7109,
    n7110, n7111, n7112, n7113, n7114, n7115,
    n7116, n7117, n7118, n7119, n7120, n7121,
    n7122, n7123, n7124, n7125, n7126, n7127,
    n7128, n7129, n7130, n7131, n7132, n7133,
    n7134, n7135, n7136, n7137, n7138, n7139,
    n7140, n7141, n7142, n7143, n7144, n7145,
    n7146, n7147, n7148, n7149, n7150, n7151,
    n7152, n7153, n7154, n7155, n7156, n7157,
    n7158, n7159, n7160, n7161, n7162, n7163,
    n7164, n7165, n7166, n7167, n7168, n7169,
    n7170, n7171, n7172, n7173, n7174, n7175,
    n7176, n7177, n7178, n7179, n7180, n7181,
    n7182, n7183, n7184, n7185, n7186, n7187,
    n7188, n7189, n7190, n7191, n7192, n7193,
    n7194, n7195, n7196, n7197, n7198, n7199,
    n7200, n7201, n7202, n7203, n7204, n7205,
    n7206, n7207, n7208, n7209, n7210, n7211,
    n7212, n7213, n7214, n7215, n7216, n7217,
    n7218, n7219, n7220, n7221, n7222, n7223,
    n7224, n7225, n7226, n7227, n7228, n7229,
    n7230, n7231, n7232, n7233, n7234, n7235,
    n7236, n7237, n7238, n7239, n7240, n7241,
    n7242, n7243, n7244, n7245, n7246, n7247,
    n7248, n7249, n7250, n7251, n7252, n7253,
    n7254, n7255, n7256, n7257, n7258, n7259,
    n7260, n7261, n7262, n7263, n7264, n7265,
    n7266, n7267, n7268, n7269, n7270, n7271,
    n7272, n7273, n7274, n7275, n7276, n7277,
    n7278, n7279, n7280, n7281, n7282, n7283,
    n7284, n7286, n7287, n7288, n7289, n7290,
    n7291, n7292, n7293, n7294, n7295, n7296,
    n7297, n7298, n7299, n7300, n7301, n7302,
    n7303, n7304, n7305, n7306, n7307, n7308,
    n7309, n7310, n7311, n7312, n7313, n7314,
    n7315, n7316, n7317, n7318, n7319, n7320,
    n7321, n7322, n7323, n7324, n7325, n7326,
    n7327, n7328, n7329, n7330, n7331, n7332,
    n7333, n7334, n7335, n7336, n7337, n7338,
    n7339, n7340, n7341, n7342, n7343, n7344,
    n7345, n7346, n7347, n7348, n7349, n7350,
    n7351, n7352, n7353, n7354, n7355, n7356,
    n7357, n7358, n7359, n7360, n7361, n7362,
    n7363, n7364, n7365, n7366, n7367, n7368,
    n7369, n7370, n7371, n7372, n7373, n7374,
    n7375, n7376, n7377, n7378, n7379, n7380,
    n7381, n7382, n7383, n7384, n7385, n7386,
    n7387, n7388, n7389, n7390, n7391, n7392,
    n7393, n7394, n7395, n7396, n7397, n7398,
    n7399, n7400, n7401, n7402, n7403, n7404,
    n7405, n7406, n7407, n7408, n7409, n7410,
    n7411, n7412, n7413, n7414, n7415, n7416,
    n7417, n7418, n7419, n7420, n7421, n7422,
    n7423, n7424, n7425, n7426, n7427, n7428,
    n7429, n7430, n7431, n7432, n7433, n7434,
    n7435, n7436, n7437, n7438, n7439, n7440,
    n7441, n7442, n7443, n7444, n7445, n7446,
    n7447, n7448, n7449, n7450, n7451, n7452,
    n7453, n7454, n7455, n7456, n7457, n7458,
    n7459, n7460, n7461, n7462, n7463, n7464,
    n7465, n7466, n7467, n7468, n7469, n7470,
    n7471, n7472, n7473, n7474, n7475, n7476,
    n7477, n7478, n7479, n7480, n7481, n7482,
    n7483, n7484, n7485, n7486, n7487, n7488,
    n7489, n7490, n7491, n7492, n7493, n7494,
    n7495, n7496, n7497, n7498, n7499, n7500,
    n7501, n7502, n7503, n7504, n7505, n7506,
    n7507, n7508, n7509, n7510, n7511, n7512,
    n7513, n7514, n7515, n7516, n7517, n7518,
    n7519, n7520, n7521, n7522, n7523, n7524,
    n7525, n7526, n7527, n7528, n7529, n7530,
    n7531, n7532, n7533, n7534, n7535, n7536,
    n7537, n7538, n7539, n7540, n7541, n7542,
    n7543, n7544, n7545, n7546, n7547, n7548,
    n7549, n7550, n7551, n7552, n7553, n7554,
    n7555, n7556, n7557, n7558, n7559, n7560,
    n7561, n7562, n7563, n7564, n7565, n7566,
    n7567, n7569, n7570, n7571, n7572, n7573,
    n7574, n7575, n7576, n7577, n7578, n7579,
    n7580, n7581, n7582, n7583, n7584, n7585,
    n7586, n7587, n7588, n7589, n7590, n7591,
    n7592, n7593, n7594, n7595, n7596, n7597,
    n7598, n7599, n7600, n7601, n7602, n7603,
    n7604, n7605, n7606, n7607, n7608, n7609,
    n7610, n7611, n7612, n7613, n7614, n7615,
    n7616, n7617, n7618, n7619, n7620, n7621,
    n7622, n7623, n7624, n7625, n7626, n7627,
    n7628, n7629, n7630, n7631, n7632, n7633,
    n7634, n7635, n7636, n7637, n7638, n7639,
    n7640, n7641, n7642, n7643, n7644, n7645,
    n7646, n7647, n7648, n7649, n7650, n7651,
    n7652, n7653, n7654, n7655, n7656, n7657,
    n7658, n7659, n7660, n7661, n7662, n7663,
    n7664, n7665, n7666, n7667, n7668, n7669,
    n7670, n7671, n7672, n7673, n7674, n7675,
    n7676, n7677, n7678, n7679, n7680, n7681,
    n7682, n7683, n7684, n7685, n7686, n7687,
    n7688, n7689, n7690, n7691, n7692, n7693,
    n7694, n7695, n7696, n7697, n7698, n7699,
    n7700, n7701, n7702, n7703, n7704, n7705,
    n7706, n7707, n7708, n7709, n7710, n7711,
    n7712, n7713, n7714, n7715, n7716, n7717,
    n7718, n7719, n7720, n7721, n7722, n7723,
    n7724, n7725, n7726, n7727, n7728, n7729,
    n7730, n7731, n7732, n7733, n7734, n7735,
    n7736, n7737, n7738, n7739, n7740, n7741,
    n7742, n7743, n7744, n7745, n7746, n7747,
    n7748, n7749, n7750, n7751, n7752, n7753,
    n7754, n7755, n7756, n7757, n7758, n7759,
    n7760, n7761, n7762, n7763, n7764, n7765,
    n7766, n7767, n7768, n7769, n7770, n7771,
    n7772, n7773, n7774, n7775, n7776, n7777,
    n7778, n7779, n7780, n7781, n7782, n7783,
    n7784, n7785, n7786, n7787, n7788, n7789,
    n7790, n7791, n7792, n7793, n7794, n7795,
    n7796, n7797, n7798, n7799, n7800, n7801,
    n7802, n7803, n7804, n7805, n7806, n7807,
    n7808, n7809, n7810, n7811, n7812, n7813,
    n7814, n7815, n7816, n7817, n7818, n7819,
    n7820, n7821, n7822, n7823, n7824, n7825,
    n7826, n7827, n7828, n7829, n7830, n7831,
    n7832, n7833, n7834, n7835, n7836, n7837,
    n7838, n7839, n7840, n7841, n7842, n7843,
    n7844, n7845, n7846, n7847, n7848, n7849,
    n7850, n7851, n7852, n7853, n7854, n7855,
    n7856, n7857, n7858, n7859, n7860, n7861,
    n7862, n7863, n7864, n7866, n7867, n7868,
    n7869, n7870, n7871, n7872, n7873, n7874,
    n7875, n7876, n7877, n7878, n7879, n7880,
    n7881, n7882, n7883, n7884, n7885, n7886,
    n7887, n7888, n7889, n7890, n7891, n7892,
    n7893, n7894, n7895, n7896, n7897, n7898,
    n7899, n7900, n7901, n7902, n7903, n7904,
    n7905, n7906, n7907, n7908, n7909, n7910,
    n7911, n7912, n7913, n7914, n7915, n7916,
    n7917, n7918, n7919, n7920, n7921, n7922,
    n7923, n7924, n7925, n7926, n7927, n7928,
    n7929, n7930, n7931, n7932, n7933, n7934,
    n7935, n7936, n7937, n7938, n7939, n7940,
    n7941, n7942, n7943, n7944, n7945, n7946,
    n7947, n7948, n7949, n7950, n7951, n7952,
    n7953, n7954, n7955, n7956, n7957, n7958,
    n7959, n7960, n7961, n7962, n7963, n7964,
    n7965, n7966, n7967, n7968, n7969, n7970,
    n7971, n7972, n7973, n7974, n7975, n7976,
    n7977, n7978, n7979, n7980, n7981, n7982,
    n7983, n7984, n7985, n7986, n7987, n7988,
    n7989, n7990, n7991, n7992, n7993, n7994,
    n7995, n7996, n7997, n7998, n7999, n8000,
    n8001, n8002, n8003, n8004, n8005, n8006,
    n8007, n8008, n8009, n8010, n8011, n8012,
    n8013, n8014, n8015, n8016, n8017, n8018,
    n8019, n8020, n8021, n8022, n8023, n8024,
    n8025, n8026, n8027, n8028, n8029, n8030,
    n8031, n8032, n8033, n8034, n8035, n8036,
    n8037, n8038, n8039, n8040, n8041, n8042,
    n8043, n8044, n8045, n8046, n8047, n8048,
    n8049, n8050, n8051, n8052, n8053, n8054,
    n8055, n8056, n8057, n8058, n8059, n8060,
    n8061, n8062, n8063, n8064, n8065, n8066,
    n8067, n8068, n8069, n8070, n8071, n8072,
    n8073, n8074, n8075, n8076, n8077, n8078,
    n8079, n8080, n8081, n8082, n8083, n8084,
    n8085, n8086, n8087, n8088, n8089, n8090,
    n8091, n8092, n8093, n8094, n8095, n8096,
    n8097, n8098, n8099, n8100, n8101, n8102,
    n8103, n8104, n8105, n8106, n8107, n8108,
    n8109, n8110, n8111, n8112, n8113, n8114,
    n8115, n8116, n8117, n8118, n8119, n8120,
    n8121, n8122, n8123, n8124, n8125, n8126,
    n8127, n8128, n8129, n8130, n8131, n8132,
    n8133, n8134, n8135, n8136, n8137, n8138,
    n8139, n8140, n8141, n8142, n8143, n8144,
    n8145, n8146, n8147, n8148, n8149, n8150,
    n8151, n8152, n8153, n8154, n8155, n8156,
    n8157, n8158, n8160, n8161, n8162, n8163,
    n8164, n8165, n8166, n8167, n8168, n8169,
    n8170, n8171, n8172, n8173, n8174, n8175,
    n8176, n8177, n8178, n8179, n8180, n8181,
    n8182, n8183, n8184, n8185, n8186, n8187,
    n8188, n8189, n8190, n8191, n8192, n8193,
    n8194, n8195, n8196, n8197, n8198, n8199,
    n8200, n8201, n8202, n8203, n8204, n8205,
    n8206, n8207, n8208, n8209, n8210, n8211,
    n8212, n8213, n8214, n8215, n8216, n8217,
    n8218, n8219, n8220, n8221, n8222, n8223,
    n8224, n8225, n8226, n8227, n8228, n8229,
    n8230, n8231, n8232, n8233, n8234, n8235,
    n8236, n8237, n8238, n8239, n8240, n8241,
    n8242, n8243, n8244, n8245, n8246, n8247,
    n8248, n8249, n8250, n8251, n8252, n8253,
    n8254, n8255, n8256, n8257, n8258, n8259,
    n8260, n8261, n8262, n8263, n8264, n8265,
    n8266, n8267, n8268, n8269, n8270, n8271,
    n8272, n8273, n8274, n8275, n8276, n8277,
    n8278, n8279, n8280, n8281, n8282, n8283,
    n8284, n8285, n8286, n8287, n8288, n8289,
    n8290, n8291, n8292, n8293, n8294, n8295,
    n8296, n8297, n8298, n8299, n8300, n8301,
    n8302, n8303, n8304, n8305, n8306, n8307,
    n8308, n8309, n8310, n8311, n8312, n8313,
    n8314, n8315, n8316, n8317, n8318, n8319,
    n8320, n8321, n8322, n8323, n8324, n8325,
    n8326, n8327, n8328, n8329, n8330, n8331,
    n8332, n8333, n8334, n8335, n8336, n8337,
    n8338, n8339, n8340, n8341, n8342, n8343,
    n8344, n8345, n8346, n8347, n8348, n8349,
    n8350, n8351, n8352, n8353, n8354, n8355,
    n8356, n8357, n8358, n8359, n8360, n8361,
    n8362, n8363, n8364, n8365, n8366, n8367,
    n8368, n8369, n8370, n8371, n8372, n8373,
    n8374, n8375, n8376, n8377, n8378, n8379,
    n8380, n8381, n8382, n8383, n8384, n8385,
    n8386, n8387, n8388, n8389, n8390, n8391,
    n8392, n8393, n8394, n8395, n8396, n8397,
    n8398, n8399, n8400, n8401, n8402, n8403,
    n8404, n8405, n8406, n8407, n8408, n8409,
    n8410, n8411, n8412, n8413, n8414, n8415,
    n8416, n8417, n8418, n8419, n8420, n8421,
    n8422, n8423, n8424, n8425, n8426, n8427,
    n8428, n8429, n8430, n8431, n8432, n8433,
    n8434, n8435, n8436, n8437, n8438, n8439,
    n8440, n8441, n8442, n8443, n8444, n8445,
    n8446, n8447, n8448, n8449, n8450, n8451,
    n8452, n8453, n8454, n8455, n8456, n8457,
    n8458, n8460, n8461, n8462, n8463, n8464,
    n8465, n8466, n8467, n8468, n8469, n8470,
    n8471, n8472, n8473, n8474, n8475, n8476,
    n8477, n8478, n8479, n8480, n8481, n8482,
    n8483, n8484, n8485, n8486, n8487, n8488,
    n8489, n8490, n8491, n8492, n8493, n8494,
    n8495, n8496, n8497, n8498, n8499, n8500,
    n8501, n8502, n8503, n8504, n8505, n8506,
    n8507, n8508, n8509, n8510, n8511, n8512,
    n8513, n8514, n8515, n8516, n8517, n8518,
    n8519, n8520, n8521, n8522, n8523, n8524,
    n8525, n8526, n8527, n8528, n8529, n8530,
    n8531, n8532, n8533, n8534, n8535, n8536,
    n8537, n8538, n8539, n8540, n8541, n8542,
    n8543, n8544, n8545, n8546, n8547, n8548,
    n8549, n8550, n8551, n8552, n8553, n8554,
    n8555, n8556, n8557, n8558, n8559, n8560,
    n8561, n8562, n8563, n8564, n8565, n8566,
    n8567, n8568, n8569, n8570, n8571, n8572,
    n8573, n8574, n8575, n8576, n8577, n8578,
    n8579, n8580, n8581, n8582, n8583, n8584,
    n8585, n8586, n8587, n8588, n8589, n8590,
    n8591, n8592, n8593, n8594, n8595, n8596,
    n8597, n8598, n8599, n8600, n8601, n8602,
    n8603, n8604, n8605, n8606, n8607, n8608,
    n8609, n8610, n8611, n8612, n8613, n8614,
    n8615, n8616, n8617, n8618, n8619, n8620,
    n8621, n8622, n8623, n8624, n8625, n8626,
    n8627, n8628, n8629, n8630, n8631, n8632,
    n8633, n8634, n8635, n8636, n8637, n8638,
    n8639, n8640, n8641, n8642, n8643, n8644,
    n8645, n8646, n8647, n8648, n8649, n8650,
    n8651, n8652, n8653, n8654, n8655, n8656,
    n8657, n8658, n8659, n8660, n8661, n8662,
    n8663, n8664, n8665, n8666, n8667, n8668,
    n8669, n8670, n8671, n8672, n8673, n8674,
    n8675, n8676, n8677, n8678, n8679, n8680,
    n8681, n8682, n8683, n8684, n8685, n8686,
    n8687, n8688, n8689, n8690, n8691, n8692,
    n8693, n8694, n8695, n8696, n8697, n8698,
    n8699, n8700, n8701, n8702, n8703, n8704,
    n8705, n8706, n8707, n8708, n8709, n8710,
    n8711, n8712, n8713, n8714, n8715, n8716,
    n8717, n8718, n8719, n8720, n8721, n8722,
    n8723, n8724, n8725, n8726, n8727, n8728,
    n8729, n8730, n8731, n8732, n8733, n8734,
    n8735, n8736, n8737, n8738, n8739, n8740,
    n8741, n8742, n8743, n8744, n8745, n8746,
    n8747, n8748, n8749, n8750, n8751, n8752,
    n8753, n8754, n8755, n8756, n8757, n8758,
    n8759, n8760, n8761, n8762, n8763, n8764,
    n8765, n8766, n8767, n8768, n8769, n8770,
    n8771, n8772, n8774, n8775, n8776, n8777,
    n8778, n8779, n8780, n8781, n8782, n8783,
    n8784, n8785, n8786, n8787, n8788, n8789,
    n8790, n8791, n8792, n8793, n8794, n8795,
    n8796, n8797, n8798, n8799, n8800, n8801,
    n8802, n8803, n8804, n8805, n8806, n8807,
    n8808, n8809, n8810, n8811, n8812, n8813,
    n8814, n8815, n8816, n8817, n8818, n8819,
    n8820, n8821, n8822, n8823, n8824, n8825,
    n8826, n8827, n8828, n8829, n8830, n8831,
    n8832, n8833, n8834, n8835, n8836, n8837,
    n8838, n8839, n8840, n8841, n8842, n8843,
    n8844, n8845, n8846, n8847, n8848, n8849,
    n8850, n8851, n8852, n8853, n8854, n8855,
    n8856, n8857, n8858, n8859, n8860, n8861,
    n8862, n8863, n8864, n8865, n8866, n8867,
    n8868, n8869, n8870, n8871, n8872, n8873,
    n8874, n8875, n8876, n8877, n8878, n8879,
    n8880, n8881, n8882, n8883, n8884, n8885,
    n8886, n8887, n8888, n8889, n8890, n8891,
    n8892, n8893, n8894, n8895, n8896, n8897,
    n8898, n8899, n8900, n8901, n8902, n8903,
    n8904, n8905, n8906, n8907, n8908, n8909,
    n8910, n8911, n8912, n8913, n8914, n8915,
    n8916, n8917, n8918, n8919, n8920, n8921,
    n8922, n8923, n8924, n8925, n8926, n8927,
    n8928, n8929, n8930, n8931, n8932, n8933,
    n8934, n8935, n8936, n8937, n8938, n8939,
    n8940, n8941, n8942, n8943, n8944, n8945,
    n8946, n8947, n8948, n8949, n8950, n8951,
    n8952, n8953, n8954, n8955, n8956, n8957,
    n8958, n8959, n8960, n8961, n8962, n8963,
    n8964, n8965, n8966, n8967, n8968, n8969,
    n8970, n8971, n8972, n8973, n8974, n8975,
    n8976, n8977, n8978, n8979, n8980, n8981,
    n8982, n8983, n8984, n8985, n8986, n8987,
    n8988, n8989, n8990, n8991, n8992, n8993,
    n8994, n8995, n8996, n8997, n8998, n8999,
    n9000, n9001, n9002, n9003, n9004, n9005,
    n9006, n9007, n9008, n9009, n9010, n9011,
    n9012, n9013, n9014, n9015, n9016, n9017,
    n9018, n9019, n9020, n9021, n9022, n9023,
    n9024, n9025, n9026, n9027, n9028, n9029,
    n9030, n9031, n9032, n9033, n9034, n9035,
    n9036, n9037, n9038, n9039, n9040, n9041,
    n9042, n9043, n9044, n9045, n9046, n9047,
    n9048, n9049, n9050, n9051, n9052, n9053,
    n9054, n9055, n9056, n9057, n9058, n9059,
    n9060, n9061, n9062, n9063, n9064, n9065,
    n9066, n9067, n9068, n9069, n9070, n9071,
    n9072, n9073, n9074, n9075, n9076, n9077,
    n9078, n9079, n9080, n9081, n9082, n9083,
    n9085, n9086, n9087, n9088, n9089, n9090,
    n9091, n9092, n9093, n9094, n9095, n9096,
    n9097, n9098, n9099, n9100, n9101, n9102,
    n9103, n9104, n9105, n9106, n9107, n9108,
    n9109, n9110, n9111, n9112, n9113, n9114,
    n9115, n9116, n9117, n9118, n9119, n9120,
    n9121, n9122, n9123, n9124, n9125, n9126,
    n9127, n9128, n9129, n9130, n9131, n9132,
    n9133, n9134, n9135, n9136, n9137, n9138,
    n9139, n9140, n9141, n9142, n9143, n9144,
    n9145, n9146, n9147, n9148, n9149, n9150,
    n9151, n9152, n9153, n9154, n9155, n9156,
    n9157, n9158, n9159, n9160, n9161, n9162,
    n9163, n9164, n9165, n9166, n9167, n9168,
    n9169, n9170, n9171, n9172, n9173, n9174,
    n9175, n9176, n9177, n9178, n9179, n9180,
    n9181, n9182, n9183, n9184, n9185, n9186,
    n9187, n9188, n9189, n9190, n9191, n9192,
    n9193, n9194, n9195, n9196, n9197, n9198,
    n9199, n9200, n9201, n9202, n9203, n9204,
    n9205, n9206, n9207, n9208, n9209, n9210,
    n9211, n9212, n9213, n9214, n9215, n9216,
    n9217, n9218, n9219, n9220, n9221, n9222,
    n9223, n9224, n9225, n9226, n9227, n9228,
    n9229, n9230, n9231, n9232, n9233, n9234,
    n9235, n9236, n9237, n9238, n9239, n9240,
    n9241, n9242, n9243, n9244, n9245, n9246,
    n9247, n9248, n9249, n9250, n9251, n9252,
    n9253, n9254, n9255, n9256, n9257, n9258,
    n9259, n9260, n9261, n9262, n9263, n9264,
    n9265, n9266, n9267, n9268, n9269, n9270,
    n9271, n9272, n9273, n9274, n9275, n9276,
    n9277, n9278, n9279, n9280, n9281, n9282,
    n9283, n9284, n9285, n9286, n9287, n9288,
    n9289, n9290, n9291, n9292, n9293, n9294,
    n9295, n9296, n9297, n9298, n9299, n9300,
    n9301, n9302, n9303, n9304, n9305, n9306,
    n9307, n9308, n9309, n9310, n9311, n9312,
    n9313, n9314, n9315, n9316, n9317, n9318,
    n9319, n9320, n9321, n9322, n9323, n9324,
    n9325, n9326, n9327, n9328, n9329, n9330,
    n9331, n9332, n9333, n9334, n9335, n9336,
    n9337, n9338, n9339, n9340, n9341, n9342,
    n9343, n9344, n9345, n9346, n9347, n9348,
    n9349, n9350, n9351, n9352, n9353, n9354,
    n9355, n9356, n9357, n9358, n9359, n9360,
    n9361, n9362, n9363, n9364, n9365, n9366,
    n9367, n9368, n9369, n9370, n9371, n9372,
    n9373, n9374, n9375, n9376, n9377, n9378,
    n9379, n9380, n9381, n9382, n9383, n9384,
    n9385, n9386, n9387, n9388, n9389, n9390,
    n9391, n9392, n9393, n9394, n9395, n9396,
    n9397, n9398, n9399, n9400, n9402, n9403,
    n9404, n9405, n9406, n9407, n9408, n9409,
    n9410, n9411, n9412, n9413, n9414, n9415,
    n9416, n9417, n9418, n9419, n9420, n9421,
    n9422, n9423, n9424, n9425, n9426, n9427,
    n9428, n9429, n9430, n9431, n9432, n9433,
    n9434, n9435, n9436, n9437, n9438, n9439,
    n9440, n9441, n9442, n9443, n9444, n9445,
    n9446, n9447, n9448, n9449, n9450, n9451,
    n9452, n9453, n9454, n9455, n9456, n9457,
    n9458, n9459, n9460, n9461, n9462, n9463,
    n9464, n9465, n9466, n9467, n9468, n9469,
    n9470, n9471, n9472, n9473, n9474, n9475,
    n9476, n9477, n9478, n9479, n9480, n9481,
    n9482, n9483, n9484, n9485, n9486, n9487,
    n9488, n9489, n9490, n9491, n9492, n9493,
    n9494, n9495, n9496, n9497, n9498, n9499,
    n9500, n9501, n9502, n9503, n9504, n9505,
    n9506, n9507, n9508, n9509, n9510, n9511,
    n9512, n9513, n9514, n9515, n9516, n9517,
    n9518, n9519, n9520, n9521, n9522, n9523,
    n9524, n9525, n9526, n9527, n9528, n9529,
    n9530, n9531, n9532, n9533, n9534, n9535,
    n9536, n9537, n9538, n9539, n9540, n9541,
    n9542, n9543, n9544, n9545, n9546, n9547,
    n9548, n9549, n9550, n9551, n9552, n9553,
    n9554, n9555, n9556, n9557, n9558, n9559,
    n9560, n9561, n9562, n9563, n9564, n9565,
    n9566, n9567, n9568, n9569, n9570, n9571,
    n9572, n9573, n9574, n9575, n9576, n9577,
    n9578, n9579, n9580, n9581, n9582, n9583,
    n9584, n9585, n9586, n9587, n9588, n9589,
    n9590, n9591, n9592, n9593, n9594, n9595,
    n9596, n9597, n9598, n9599, n9600, n9601,
    n9602, n9603, n9604, n9605, n9606, n9607,
    n9608, n9609, n9610, n9611, n9612, n9613,
    n9614, n9615, n9616, n9617, n9618, n9619,
    n9620, n9621, n9622, n9623, n9624, n9625,
    n9626, n9627, n9628, n9629, n9630, n9631,
    n9632, n9633, n9634, n9635, n9636, n9637,
    n9638, n9639, n9640, n9641, n9642, n9643,
    n9644, n9645, n9646, n9647, n9648, n9649,
    n9650, n9651, n9652, n9653, n9654, n9655,
    n9656, n9657, n9658, n9659, n9660, n9661,
    n9662, n9663, n9664, n9665, n9666, n9667,
    n9668, n9669, n9670, n9671, n9672, n9673,
    n9674, n9675, n9676, n9677, n9678, n9679,
    n9680, n9681, n9682, n9683, n9684, n9685,
    n9686, n9687, n9688, n9689, n9690, n9691,
    n9692, n9693, n9694, n9695, n9696, n9697,
    n9698, n9699, n9700, n9701, n9702, n9703,
    n9704, n9705, n9706, n9707, n9708, n9709,
    n9710, n9711, n9712, n9713, n9714, n9715,
    n9716, n9717, n9718, n9719, n9720, n9721,
    n9722, n9723, n9724, n9725, n9726, n9727,
    n9728, n9729, n9730, n9731, n9733, n9734,
    n9735, n9736, n9737, n9738, n9739, n9740,
    n9741, n9742, n9743, n9744, n9745, n9746,
    n9747, n9748, n9749, n9750, n9751, n9752,
    n9753, n9754, n9755, n9756, n9757, n9758,
    n9759, n9760, n9761, n9762, n9763, n9764,
    n9765, n9766, n9767, n9768, n9769, n9770,
    n9771, n9772, n9773, n9774, n9775, n9776,
    n9777, n9778, n9779, n9780, n9781, n9782,
    n9783, n9784, n9785, n9786, n9787, n9788,
    n9789, n9790, n9791, n9792, n9793, n9794,
    n9795, n9796, n9797, n9798, n9799, n9800,
    n9801, n9802, n9803, n9804, n9805, n9806,
    n9807, n9808, n9809, n9810, n9811, n9812,
    n9813, n9814, n9815, n9816, n9817, n9818,
    n9819, n9820, n9821, n9822, n9823, n9824,
    n9825, n9826, n9827, n9828, n9829, n9830,
    n9831, n9832, n9833, n9834, n9835, n9836,
    n9837, n9838, n9839, n9840, n9841, n9842,
    n9843, n9844, n9845, n9846, n9847, n9848,
    n9849, n9850, n9851, n9852, n9853, n9854,
    n9855, n9856, n9857, n9858, n9859, n9860,
    n9861, n9862, n9863, n9864, n9865, n9866,
    n9867, n9868, n9869, n9870, n9871, n9872,
    n9873, n9874, n9875, n9876, n9877, n9878,
    n9879, n9880, n9881, n9882, n9883, n9884,
    n9885, n9886, n9887, n9888, n9889, n9890,
    n9891, n9892, n9893, n9894, n9895, n9896,
    n9897, n9898, n9899, n9900, n9901, n9902,
    n9903, n9904, n9905, n9906, n9907, n9908,
    n9909, n9910, n9911, n9912, n9913, n9914,
    n9915, n9916, n9917, n9918, n9919, n9920,
    n9921, n9922, n9923, n9924, n9925, n9926,
    n9927, n9928, n9929, n9930, n9931, n9932,
    n9933, n9934, n9935, n9936, n9937, n9938,
    n9939, n9940, n9941, n9942, n9943, n9944,
    n9945, n9946, n9947, n9948, n9949, n9950,
    n9951, n9952, n9953, n9954, n9955, n9956,
    n9957, n9958, n9959, n9960, n9961, n9962,
    n9963, n9964, n9965, n9966, n9967, n9968,
    n9969, n9970, n9971, n9972, n9973, n9974,
    n9975, n9976, n9977, n9978, n9979, n9980,
    n9981, n9982, n9983, n9984, n9985, n9986,
    n9987, n9988, n9989, n9990, n9991, n9992,
    n9993, n9994, n9995, n9996, n9997, n9998,
    n9999, n10000, n10001, n10002, n10003, n10004,
    n10005, n10006, n10007, n10008, n10009, n10010,
    n10011, n10012, n10013, n10014, n10015, n10016,
    n10017, n10018, n10019, n10020, n10021, n10022,
    n10023, n10024, n10025, n10026, n10027, n10028,
    n10029, n10030, n10031, n10032, n10033, n10034,
    n10035, n10036, n10037, n10038, n10039, n10040,
    n10041, n10042, n10043, n10044, n10045, n10046,
    n10047, n10048, n10049, n10050, n10051, n10052,
    n10053, n10054, n10055, n10056, n10057, n10058,
    n10059, n10061, n10062, n10063, n10064, n10065,
    n10066, n10067, n10068, n10069, n10070, n10071,
    n10072, n10073, n10074, n10075, n10076, n10077,
    n10078, n10079, n10080, n10081, n10082, n10083,
    n10084, n10085, n10086, n10087, n10088, n10089,
    n10090, n10091, n10092, n10093, n10094, n10095,
    n10096, n10097, n10098, n10099, n10100, n10101,
    n10102, n10103, n10104, n10105, n10106, n10107,
    n10108, n10109, n10110, n10111, n10112, n10113,
    n10114, n10115, n10116, n10117, n10118, n10119,
    n10120, n10121, n10122, n10123, n10124, n10125,
    n10126, n10127, n10128, n10129, n10130, n10131,
    n10132, n10133, n10134, n10135, n10136, n10137,
    n10138, n10139, n10140, n10141, n10142, n10143,
    n10144, n10145, n10146, n10147, n10148, n10149,
    n10150, n10151, n10152, n10153, n10154, n10155,
    n10156, n10157, n10158, n10159, n10160, n10161,
    n10162, n10163, n10164, n10165, n10166, n10167,
    n10168, n10169, n10170, n10171, n10172, n10173,
    n10174, n10175, n10176, n10177, n10178, n10179,
    n10180, n10181, n10182, n10183, n10184, n10185,
    n10186, n10187, n10188, n10189, n10190, n10191,
    n10192, n10193, n10194, n10195, n10196, n10197,
    n10198, n10199, n10200, n10201, n10202, n10203,
    n10204, n10205, n10206, n10207, n10208, n10209,
    n10210, n10211, n10212, n10213, n10214, n10215,
    n10216, n10217, n10218, n10219, n10220, n10221,
    n10222, n10223, n10224, n10225, n10226, n10227,
    n10228, n10229, n10230, n10231, n10232, n10233,
    n10234, n10235, n10236, n10237, n10238, n10239,
    n10240, n10241, n10242, n10243, n10244, n10245,
    n10246, n10247, n10248, n10249, n10250, n10251,
    n10252, n10253, n10254, n10255, n10256, n10257,
    n10258, n10259, n10260, n10261, n10262, n10263,
    n10264, n10265, n10266, n10267, n10268, n10269,
    n10270, n10271, n10272, n10273, n10274, n10275,
    n10276, n10277, n10278, n10279, n10280, n10281,
    n10282, n10283, n10284, n10285, n10286, n10287,
    n10288, n10289, n10290, n10291, n10292, n10293,
    n10294, n10295, n10296, n10297, n10298, n10299,
    n10300, n10301, n10302, n10303, n10304, n10305,
    n10306, n10307, n10308, n10309, n10310, n10311,
    n10312, n10313, n10314, n10315, n10316, n10317,
    n10318, n10319, n10320, n10321, n10322, n10323,
    n10324, n10325, n10326, n10327, n10328, n10329,
    n10330, n10331, n10332, n10333, n10334, n10335,
    n10336, n10337, n10338, n10339, n10340, n10341,
    n10342, n10343, n10344, n10345, n10346, n10347,
    n10348, n10349, n10350, n10351, n10352, n10353,
    n10354, n10355, n10356, n10357, n10358, n10359,
    n10360, n10361, n10362, n10363, n10364, n10365,
    n10366, n10367, n10368, n10369, n10370, n10371,
    n10372, n10373, n10374, n10375, n10376, n10377,
    n10378, n10379, n10380, n10381, n10382, n10383,
    n10384, n10385, n10386, n10387, n10388, n10389,
    n10390, n10391, n10392, n10393, n10395, n10396,
    n10397, n10398, n10399, n10400, n10401, n10402,
    n10403, n10404, n10405, n10406, n10407, n10408,
    n10409, n10410, n10411, n10412, n10413, n10414,
    n10415, n10416, n10417, n10418, n10419, n10420,
    n10421, n10422, n10423, n10424, n10425, n10426,
    n10427, n10428, n10429, n10430, n10431, n10432,
    n10433, n10434, n10435, n10436, n10437, n10438,
    n10439, n10440, n10441, n10442, n10443, n10444,
    n10445, n10446, n10447, n10448, n10449, n10450,
    n10451, n10452, n10453, n10454, n10455, n10456,
    n10457, n10458, n10459, n10460, n10461, n10462,
    n10463, n10464, n10465, n10466, n10467, n10468,
    n10469, n10470, n10471, n10472, n10473, n10474,
    n10475, n10476, n10477, n10478, n10479, n10480,
    n10481, n10482, n10483, n10484, n10485, n10486,
    n10487, n10488, n10489, n10490, n10491, n10492,
    n10493, n10494, n10495, n10496, n10497, n10498,
    n10499, n10500, n10501, n10502, n10503, n10504,
    n10505, n10506, n10507, n10508, n10509, n10510,
    n10511, n10512, n10513, n10514, n10515, n10516,
    n10517, n10518, n10519, n10520, n10521, n10522,
    n10523, n10524, n10525, n10526, n10527, n10528,
    n10529, n10530, n10531, n10532, n10533, n10534,
    n10535, n10536, n10537, n10538, n10539, n10540,
    n10541, n10542, n10543, n10544, n10545, n10546,
    n10547, n10548, n10549, n10550, n10551, n10552,
    n10553, n10554, n10555, n10556, n10557, n10558,
    n10559, n10560, n10561, n10562, n10563, n10564,
    n10565, n10566, n10567, n10568, n10569, n10570,
    n10571, n10572, n10573, n10574, n10575, n10576,
    n10577, n10578, n10579, n10580, n10581, n10582,
    n10583, n10584, n10585, n10586, n10587, n10588,
    n10589, n10590, n10591, n10592, n10593, n10594,
    n10595, n10596, n10597, n10598, n10599, n10600,
    n10601, n10602, n10603, n10604, n10605, n10606,
    n10607, n10608, n10609, n10610, n10611, n10612,
    n10613, n10614, n10615, n10616, n10617, n10618,
    n10619, n10620, n10621, n10622, n10623, n10624,
    n10625, n10626, n10627, n10628, n10629, n10630,
    n10631, n10632, n10633, n10634, n10635, n10636,
    n10637, n10638, n10639, n10640, n10641, n10642,
    n10643, n10644, n10645, n10646, n10647, n10648,
    n10649, n10650, n10651, n10652, n10653, n10654,
    n10655, n10656, n10657, n10658, n10659, n10660,
    n10661, n10662, n10663, n10664, n10665, n10666,
    n10667, n10668, n10669, n10670, n10671, n10672,
    n10673, n10674, n10675, n10676, n10677, n10678,
    n10679, n10680, n10681, n10682, n10683, n10684,
    n10685, n10686, n10687, n10688, n10689, n10690,
    n10691, n10692, n10693, n10694, n10695, n10696,
    n10697, n10698, n10699, n10700, n10701, n10702,
    n10703, n10704, n10705, n10706, n10707, n10708,
    n10709, n10710, n10711, n10712, n10713, n10714,
    n10715, n10716, n10717, n10718, n10719, n10720,
    n10721, n10722, n10723, n10724, n10725, n10726,
    n10727, n10728, n10729, n10730, n10731, n10732,
    n10733, n10734, n10735, n10736, n10737, n10738,
    n10739, n10740, n10741, n10743, n10744, n10745,
    n10746, n10747, n10748, n10749, n10750, n10751,
    n10752, n10753, n10754, n10755, n10756, n10757,
    n10758, n10759, n10760, n10761, n10762, n10763,
    n10764, n10765, n10766, n10767, n10768, n10769,
    n10770, n10771, n10772, n10773, n10774, n10775,
    n10776, n10777, n10778, n10779, n10780, n10781,
    n10782, n10783, n10784, n10785, n10786, n10787,
    n10788, n10789, n10790, n10791, n10792, n10793,
    n10794, n10795, n10796, n10797, n10798, n10799,
    n10800, n10801, n10802, n10803, n10804, n10805,
    n10806, n10807, n10808, n10809, n10810, n10811,
    n10812, n10813, n10814, n10815, n10816, n10817,
    n10818, n10819, n10820, n10821, n10822, n10823,
    n10824, n10825, n10826, n10827, n10828, n10829,
    n10830, n10831, n10832, n10833, n10834, n10835,
    n10836, n10837, n10838, n10839, n10840, n10841,
    n10842, n10843, n10844, n10845, n10846, n10847,
    n10848, n10849, n10850, n10851, n10852, n10853,
    n10854, n10855, n10856, n10857, n10858, n10859,
    n10860, n10861, n10862, n10863, n10864, n10865,
    n10866, n10867, n10868, n10869, n10870, n10871,
    n10872, n10873, n10874, n10875, n10876, n10877,
    n10878, n10879, n10880, n10881, n10882, n10883,
    n10884, n10885, n10886, n10887, n10888, n10889,
    n10890, n10891, n10892, n10893, n10894, n10895,
    n10896, n10897, n10898, n10899, n10900, n10901,
    n10902, n10903, n10904, n10905, n10906, n10907,
    n10908, n10909, n10910, n10911, n10912, n10913,
    n10914, n10915, n10916, n10917, n10918, n10919,
    n10920, n10921, n10922, n10923, n10924, n10925,
    n10926, n10927, n10928, n10929, n10930, n10931,
    n10932, n10933, n10934, n10935, n10936, n10937,
    n10938, n10939, n10940, n10941, n10942, n10943,
    n10944, n10945, n10946, n10947, n10948, n10949,
    n10950, n10951, n10952, n10953, n10954, n10955,
    n10956, n10957, n10958, n10959, n10960, n10961,
    n10962, n10963, n10964, n10965, n10966, n10967,
    n10968, n10969, n10970, n10971, n10972, n10973,
    n10974, n10975, n10976, n10977, n10978, n10979,
    n10980, n10981, n10982, n10983, n10984, n10985,
    n10986, n10987, n10988, n10989, n10990, n10991,
    n10992, n10993, n10994, n10995, n10996, n10997,
    n10998, n10999, n11000, n11001, n11002, n11003,
    n11004, n11005, n11006, n11007, n11008, n11009,
    n11010, n11011, n11012, n11013, n11014, n11015,
    n11016, n11017, n11018, n11019, n11020, n11021,
    n11022, n11023, n11024, n11025, n11026, n11027,
    n11028, n11029, n11030, n11031, n11032, n11033,
    n11034, n11035, n11036, n11037, n11038, n11039,
    n11040, n11041, n11042, n11043, n11044, n11045,
    n11046, n11047, n11048, n11049, n11050, n11051,
    n11052, n11053, n11054, n11055, n11056, n11057,
    n11058, n11059, n11060, n11061, n11062, n11063,
    n11064, n11065, n11066, n11067, n11068, n11069,
    n11070, n11071, n11072, n11073, n11074, n11075,
    n11076, n11077, n11078, n11079, n11080, n11081,
    n11082, n11083, n11084, n11085, n11086, n11088,
    n11089, n11090, n11091, n11092, n11093, n11094,
    n11095, n11096, n11097, n11098, n11099, n11100,
    n11101, n11102, n11103, n11104, n11105, n11106,
    n11107, n11108, n11109, n11110, n11111, n11112,
    n11113, n11114, n11115, n11116, n11117, n11118,
    n11119, n11120, n11121, n11122, n11123, n11124,
    n11125, n11126, n11127, n11128, n11129, n11130,
    n11131, n11132, n11133, n11134, n11135, n11136,
    n11137, n11138, n11139, n11140, n11141, n11142,
    n11143, n11144, n11145, n11146, n11147, n11148,
    n11149, n11150, n11151, n11152, n11153, n11154,
    n11155, n11156, n11157, n11158, n11159, n11160,
    n11161, n11162, n11163, n11164, n11165, n11166,
    n11167, n11168, n11169, n11170, n11171, n11172,
    n11173, n11174, n11175, n11176, n11177, n11178,
    n11179, n11180, n11181, n11182, n11183, n11184,
    n11185, n11186, n11187, n11188, n11189, n11190,
    n11191, n11192, n11193, n11194, n11195, n11196,
    n11197, n11198, n11199, n11200, n11201, n11202,
    n11203, n11204, n11205, n11206, n11207, n11208,
    n11209, n11210, n11211, n11212, n11213, n11214,
    n11215, n11216, n11217, n11218, n11219, n11220,
    n11221, n11222, n11223, n11224, n11225, n11226,
    n11227, n11228, n11229, n11230, n11231, n11232,
    n11233, n11234, n11235, n11236, n11237, n11238,
    n11239, n11240, n11241, n11242, n11243, n11244,
    n11245, n11246, n11247, n11248, n11249, n11250,
    n11251, n11252, n11253, n11254, n11255, n11256,
    n11257, n11258, n11259, n11260, n11261, n11262,
    n11263, n11264, n11265, n11266, n11267, n11268,
    n11269, n11270, n11271, n11272, n11273, n11274,
    n11275, n11276, n11277, n11278, n11279, n11280,
    n11281, n11282, n11283, n11284, n11285, n11286,
    n11287, n11288, n11289, n11290, n11291, n11292,
    n11293, n11294, n11295, n11296, n11297, n11298,
    n11299, n11300, n11301, n11302, n11303, n11304,
    n11305, n11306, n11307, n11308, n11309, n11310,
    n11311, n11312, n11313, n11314, n11315, n11316,
    n11317, n11318, n11319, n11320, n11321, n11322,
    n11323, n11324, n11325, n11326, n11327, n11328,
    n11329, n11330, n11331, n11332, n11333, n11334,
    n11335, n11336, n11337, n11338, n11339, n11340,
    n11341, n11342, n11343, n11344, n11345, n11346,
    n11347, n11348, n11349, n11350, n11351, n11352,
    n11353, n11354, n11355, n11356, n11357, n11358,
    n11359, n11360, n11361, n11362, n11363, n11364,
    n11365, n11366, n11367, n11368, n11369, n11370,
    n11371, n11372, n11373, n11374, n11375, n11376,
    n11377, n11378, n11379, n11380, n11381, n11382,
    n11383, n11384, n11385, n11386, n11387, n11388,
    n11389, n11390, n11391, n11392, n11393, n11394,
    n11395, n11396, n11397, n11398, n11399, n11400,
    n11401, n11402, n11403, n11404, n11405, n11406,
    n11407, n11408, n11409, n11410, n11411, n11412,
    n11413, n11414, n11415, n11416, n11417, n11418,
    n11419, n11420, n11421, n11422, n11423, n11424,
    n11425, n11426, n11427, n11428, n11429, n11430,
    n11431, n11432, n11433, n11434, n11435, n11436,
    n11437, n11439, n11440, n11441, n11442, n11443,
    n11444, n11445, n11446, n11447, n11448, n11449,
    n11450, n11451, n11452, n11453, n11454, n11455,
    n11456, n11457, n11458, n11459, n11460, n11461,
    n11462, n11463, n11464, n11465, n11466, n11467,
    n11468, n11469, n11470, n11471, n11472, n11473,
    n11474, n11475, n11476, n11477, n11478, n11479,
    n11480, n11481, n11482, n11483, n11484, n11485,
    n11486, n11487, n11488, n11489, n11490, n11491,
    n11492, n11493, n11494, n11495, n11496, n11497,
    n11498, n11499, n11500, n11501, n11502, n11503,
    n11504, n11505, n11506, n11507, n11508, n11509,
    n11510, n11511, n11512, n11513, n11514, n11515,
    n11516, n11517, n11518, n11519, n11520, n11521,
    n11522, n11523, n11524, n11525, n11526, n11527,
    n11528, n11529, n11530, n11531, n11532, n11533,
    n11534, n11535, n11536, n11537, n11538, n11539,
    n11540, n11541, n11542, n11543, n11544, n11545,
    n11546, n11547, n11548, n11549, n11550, n11551,
    n11552, n11553, n11554, n11555, n11556, n11557,
    n11558, n11559, n11560, n11561, n11562, n11563,
    n11564, n11565, n11566, n11567, n11568, n11569,
    n11570, n11571, n11572, n11573, n11574, n11575,
    n11576, n11577, n11578, n11579, n11580, n11581,
    n11582, n11583, n11584, n11585, n11586, n11587,
    n11588, n11589, n11590, n11591, n11592, n11593,
    n11594, n11595, n11596, n11597, n11598, n11599,
    n11600, n11601, n11602, n11603, n11604, n11605,
    n11606, n11607, n11608, n11609, n11610, n11611,
    n11612, n11613, n11614, n11615, n11616, n11617,
    n11618, n11619, n11620, n11621, n11622, n11623,
    n11624, n11625, n11626, n11627, n11628, n11629,
    n11630, n11631, n11632, n11633, n11634, n11635,
    n11636, n11637, n11638, n11639, n11640, n11641,
    n11642, n11643, n11644, n11645, n11646, n11647,
    n11648, n11649, n11650, n11651, n11652, n11653,
    n11654, n11655, n11656, n11657, n11658, n11659,
    n11660, n11661, n11662, n11663, n11664, n11665,
    n11666, n11667, n11668, n11669, n11670, n11671,
    n11672, n11673, n11674, n11675, n11676, n11677,
    n11678, n11679, n11680, n11681, n11682, n11683,
    n11684, n11685, n11686, n11687, n11688, n11689,
    n11690, n11691, n11692, n11693, n11694, n11695,
    n11696, n11697, n11698, n11699, n11700, n11701,
    n11702, n11703, n11704, n11705, n11706, n11707,
    n11708, n11709, n11710, n11711, n11712, n11713,
    n11714, n11715, n11716, n11717, n11718, n11719,
    n11720, n11721, n11722, n11723, n11724, n11725,
    n11726, n11727, n11728, n11729, n11730, n11731,
    n11732, n11733, n11734, n11735, n11736, n11737,
    n11738, n11739, n11740, n11741, n11742, n11743,
    n11744, n11745, n11746, n11747, n11748, n11749,
    n11750, n11751, n11752, n11753, n11754, n11755,
    n11756, n11757, n11758, n11759, n11760, n11761,
    n11762, n11763, n11764, n11765, n11766, n11767,
    n11768, n11769, n11770, n11771, n11772, n11773,
    n11774, n11775, n11776, n11777, n11778, n11779,
    n11780, n11781, n11782, n11783, n11784, n11785,
    n11786, n11787, n11788, n11789, n11790, n11791,
    n11792, n11793, n11794, n11795, n11796, n11797,
    n11798, n11799, n11800, n11801, n11802, n11804,
    n11805, n11806, n11807, n11808, n11809, n11810,
    n11811, n11812, n11813, n11814, n11815, n11816,
    n11817, n11818, n11819, n11820, n11821, n11822,
    n11823, n11824, n11825, n11826, n11827, n11828,
    n11829, n11830, n11831, n11832, n11833, n11834,
    n11835, n11836, n11837, n11838, n11839, n11840,
    n11841, n11842, n11843, n11844, n11845, n11846,
    n11847, n11848, n11849, n11850, n11851, n11852,
    n11853, n11854, n11855, n11856, n11857, n11858,
    n11859, n11860, n11861, n11862, n11863, n11864,
    n11865, n11866, n11867, n11868, n11869, n11870,
    n11871, n11872, n11873, n11874, n11875, n11876,
    n11877, n11878, n11879, n11880, n11881, n11882,
    n11883, n11884, n11885, n11886, n11887, n11888,
    n11889, n11890, n11891, n11892, n11893, n11894,
    n11895, n11896, n11897, n11898, n11899, n11900,
    n11901, n11902, n11903, n11904, n11905, n11906,
    n11907, n11908, n11909, n11910, n11911, n11912,
    n11913, n11914, n11915, n11916, n11917, n11918,
    n11919, n11920, n11921, n11922, n11923, n11924,
    n11925, n11926, n11927, n11928, n11929, n11930,
    n11931, n11932, n11933, n11934, n11935, n11936,
    n11937, n11938, n11939, n11940, n11941, n11942,
    n11943, n11944, n11945, n11946, n11947, n11948,
    n11949, n11950, n11951, n11952, n11953, n11954,
    n11955, n11956, n11957, n11958, n11959, n11960,
    n11961, n11962, n11963, n11964, n11965, n11966,
    n11967, n11968, n11969, n11970, n11971, n11972,
    n11973, n11974, n11975, n11976, n11977, n11978,
    n11979, n11980, n11981, n11982, n11983, n11984,
    n11985, n11986, n11987, n11988, n11989, n11990,
    n11991, n11992, n11993, n11994, n11995, n11996,
    n11997, n11998, n11999, n12000, n12001, n12002,
    n12003, n12004, n12005, n12006, n12007, n12008,
    n12009, n12010, n12011, n12012, n12013, n12014,
    n12015, n12016, n12017, n12018, n12019, n12020,
    n12021, n12022, n12023, n12024, n12025, n12026,
    n12027, n12028, n12029, n12030, n12031, n12032,
    n12033, n12034, n12035, n12036, n12037, n12038,
    n12039, n12040, n12041, n12042, n12043, n12044,
    n12045, n12046, n12047, n12048, n12049, n12050,
    n12051, n12052, n12053, n12054, n12055, n12056,
    n12057, n12058, n12059, n12060, n12061, n12062,
    n12063, n12064, n12065, n12066, n12067, n12068,
    n12069, n12070, n12071, n12072, n12073, n12074,
    n12075, n12076, n12077, n12078, n12079, n12080,
    n12081, n12082, n12083, n12084, n12085, n12086,
    n12087, n12088, n12089, n12090, n12091, n12092,
    n12093, n12094, n12095, n12096, n12097, n12098,
    n12099, n12100, n12101, n12102, n12103, n12104,
    n12105, n12106, n12107, n12108, n12109, n12110,
    n12111, n12112, n12113, n12114, n12115, n12116,
    n12117, n12118, n12119, n12120, n12121, n12122,
    n12123, n12124, n12125, n12126, n12127, n12128,
    n12129, n12130, n12131, n12132, n12133, n12134,
    n12135, n12136, n12137, n12138, n12139, n12140,
    n12141, n12142, n12143, n12144, n12145, n12146,
    n12147, n12148, n12149, n12150, n12151, n12152,
    n12153, n12154, n12155, n12156, n12157, n12158,
    n12159, n12160, n12161, n12162, n12163, n12164,
    n12165, n12167, n12168, n12169, n12170, n12171,
    n12172, n12173, n12174, n12175, n12176, n12177,
    n12178, n12179, n12180, n12181, n12182, n12183,
    n12184, n12185, n12186, n12187, n12188, n12189,
    n12190, n12191, n12192, n12193, n12194, n12195,
    n12196, n12197, n12198, n12199, n12200, n12201,
    n12202, n12203, n12204, n12205, n12206, n12207,
    n12208, n12209, n12210, n12211, n12212, n12213,
    n12214, n12215, n12216, n12217, n12218, n12219,
    n12220, n12221, n12222, n12223, n12224, n12225,
    n12226, n12227, n12228, n12229, n12230, n12231,
    n12232, n12233, n12234, n12235, n12236, n12237,
    n12238, n12239, n12240, n12241, n12242, n12243,
    n12244, n12245, n12246, n12247, n12248, n12249,
    n12250, n12251, n12252, n12253, n12254, n12255,
    n12256, n12257, n12258, n12259, n12260, n12261,
    n12262, n12263, n12264, n12265, n12266, n12267,
    n12268, n12269, n12270, n12271, n12272, n12273,
    n12274, n12275, n12276, n12277, n12278, n12279,
    n12280, n12281, n12282, n12283, n12284, n12285,
    n12286, n12287, n12288, n12289, n12290, n12291,
    n12292, n12293, n12294, n12295, n12296, n12297,
    n12298, n12299, n12300, n12301, n12302, n12303,
    n12304, n12305, n12306, n12307, n12308, n12309,
    n12310, n12311, n12312, n12313, n12314, n12315,
    n12316, n12317, n12318, n12319, n12320, n12321,
    n12322, n12323, n12324, n12325, n12326, n12327,
    n12328, n12329, n12330, n12331, n12332, n12333,
    n12334, n12335, n12336, n12337, n12338, n12339,
    n12340, n12341, n12342, n12343, n12344, n12345,
    n12346, n12347, n12348, n12349, n12350, n12351,
    n12352, n12353, n12354, n12355, n12356, n12357,
    n12358, n12359, n12360, n12361, n12362, n12363,
    n12364, n12365, n12366, n12367, n12368, n12369,
    n12370, n12371, n12372, n12373, n12374, n12375,
    n12376, n12377, n12378, n12379, n12380, n12381,
    n12382, n12383, n12384, n12385, n12386, n12387,
    n12388, n12389, n12390, n12391, n12392, n12393,
    n12394, n12395, n12396, n12397, n12398, n12399,
    n12400, n12401, n12402, n12403, n12404, n12405,
    n12406, n12407, n12408, n12409, n12410, n12411,
    n12412, n12413, n12414, n12415, n12416, n12417,
    n12418, n12419, n12420, n12421, n12422, n12423,
    n12424, n12425, n12426, n12427, n12428, n12429,
    n12430, n12431, n12432, n12433, n12434, n12435,
    n12436, n12437, n12438, n12439, n12440, n12441,
    n12442, n12443, n12444, n12445, n12446, n12447,
    n12448, n12449, n12450, n12451, n12452, n12453,
    n12454, n12455, n12456, n12457, n12458, n12459,
    n12460, n12461, n12462, n12463, n12464, n12465,
    n12466, n12467, n12468, n12469, n12470, n12471,
    n12472, n12473, n12474, n12475, n12476, n12477,
    n12478, n12479, n12480, n12481, n12482, n12483,
    n12484, n12485, n12486, n12487, n12488, n12489,
    n12490, n12491, n12492, n12493, n12494, n12495,
    n12496, n12497, n12498, n12499, n12500, n12501,
    n12502, n12503, n12504, n12505, n12506, n12507,
    n12508, n12509, n12510, n12511, n12512, n12513,
    n12514, n12515, n12516, n12517, n12518, n12519,
    n12520, n12521, n12522, n12523, n12524, n12525,
    n12526, n12527, n12528, n12529, n12530, n12531,
    n12532, n12533, n12534, n12536, n12537, n12538,
    n12539, n12540, n12541, n12542, n12543, n12544,
    n12545, n12546, n12547, n12548, n12549, n12550,
    n12551, n12552, n12553, n12554, n12555, n12556,
    n12557, n12558, n12559, n12560, n12561, n12562,
    n12563, n12564, n12565, n12566, n12567, n12568,
    n12569, n12570, n12571, n12572, n12573, n12574,
    n12575, n12576, n12577, n12578, n12579, n12580,
    n12581, n12582, n12583, n12584, n12585, n12586,
    n12587, n12588, n12589, n12590, n12591, n12592,
    n12593, n12594, n12595, n12596, n12597, n12598,
    n12599, n12600, n12601, n12602, n12603, n12604,
    n12605, n12606, n12607, n12608, n12609, n12610,
    n12611, n12612, n12613, n12614, n12615, n12616,
    n12617, n12618, n12619, n12620, n12621, n12622,
    n12623, n12624, n12625, n12626, n12627, n12628,
    n12629, n12630, n12631, n12632, n12633, n12634,
    n12635, n12636, n12637, n12638, n12639, n12640,
    n12641, n12642, n12643, n12644, n12645, n12646,
    n12647, n12648, n12649, n12650, n12651, n12652,
    n12653, n12654, n12655, n12656, n12657, n12658,
    n12659, n12660, n12661, n12662, n12663, n12664,
    n12665, n12666, n12667, n12668, n12669, n12670,
    n12671, n12672, n12673, n12674, n12675, n12676,
    n12677, n12678, n12679, n12680, n12681, n12682,
    n12683, n12684, n12685, n12686, n12687, n12688,
    n12689, n12690, n12691, n12692, n12693, n12694,
    n12695, n12696, n12697, n12698, n12699, n12700,
    n12701, n12702, n12703, n12704, n12705, n12706,
    n12707, n12708, n12709, n12710, n12711, n12712,
    n12713, n12714, n12715, n12716, n12717, n12718,
    n12719, n12720, n12721, n12722, n12723, n12724,
    n12725, n12726, n12727, n12728, n12729, n12730,
    n12731, n12732, n12733, n12734, n12735, n12736,
    n12737, n12738, n12739, n12740, n12741, n12742,
    n12743, n12744, n12745, n12746, n12747, n12748,
    n12749, n12750, n12751, n12752, n12753, n12754,
    n12755, n12756, n12757, n12758, n12759, n12760,
    n12761, n12762, n12763, n12764, n12765, n12766,
    n12767, n12768, n12769, n12770, n12771, n12772,
    n12773, n12774, n12775, n12776, n12777, n12778,
    n12779, n12780, n12781, n12782, n12783, n12784,
    n12785, n12786, n12787, n12788, n12789, n12790,
    n12791, n12792, n12793, n12794, n12795, n12796,
    n12797, n12798, n12799, n12800, n12801, n12802,
    n12803, n12804, n12805, n12806, n12807, n12808,
    n12809, n12810, n12811, n12812, n12813, n12814,
    n12815, n12816, n12817, n12818, n12819, n12820,
    n12821, n12822, n12823, n12824, n12825, n12826,
    n12827, n12828, n12829, n12830, n12831, n12832,
    n12833, n12834, n12835, n12836, n12837, n12838,
    n12839, n12840, n12841, n12842, n12843, n12844,
    n12845, n12846, n12847, n12848, n12849, n12850,
    n12851, n12852, n12853, n12854, n12855, n12856,
    n12857, n12858, n12859, n12860, n12861, n12862,
    n12863, n12864, n12865, n12866, n12867, n12868,
    n12869, n12870, n12871, n12872, n12873, n12874,
    n12875, n12876, n12877, n12878, n12879, n12880,
    n12881, n12882, n12883, n12884, n12885, n12886,
    n12887, n12888, n12889, n12890, n12891, n12892,
    n12893, n12894, n12895, n12896, n12897, n12898,
    n12900, n12901, n12902, n12903, n12904, n12905,
    n12906, n12907, n12908, n12909, n12910, n12911,
    n12912, n12913, n12914, n12915, n12916, n12917,
    n12918, n12919, n12920, n12921, n12922, n12923,
    n12924, n12925, n12926, n12927, n12928, n12929,
    n12930, n12931, n12932, n12933, n12934, n12935,
    n12936, n12937, n12938, n12939, n12940, n12941,
    n12942, n12943, n12944, n12945, n12946, n12947,
    n12948, n12949, n12950, n12951, n12952, n12953,
    n12954, n12955, n12956, n12957, n12958, n12959,
    n12960, n12961, n12962, n12963, n12964, n12965,
    n12966, n12967, n12968, n12969, n12970, n12971,
    n12972, n12973, n12974, n12975, n12976, n12977,
    n12978, n12979, n12980, n12981, n12982, n12983,
    n12984, n12985, n12986, n12987, n12988, n12989,
    n12990, n12991, n12992, n12993, n12994, n12995,
    n12996, n12997, n12998, n12999, n13000, n13001,
    n13002, n13003, n13004, n13005, n13006, n13007,
    n13008, n13009, n13010, n13011, n13012, n13013,
    n13014, n13015, n13016, n13017, n13018, n13019,
    n13020, n13021, n13022, n13023, n13024, n13025,
    n13026, n13027, n13028, n13029, n13030, n13031,
    n13032, n13033, n13034, n13035, n13036, n13037,
    n13038, n13039, n13040, n13041, n13042, n13043,
    n13044, n13045, n13046, n13047, n13048, n13049,
    n13050, n13051, n13052, n13053, n13054, n13055,
    n13056, n13057, n13058, n13059, n13060, n13061,
    n13062, n13063, n13064, n13065, n13066, n13067,
    n13068, n13069, n13070, n13071, n13072, n13073,
    n13074, n13075, n13076, n13077, n13078, n13079,
    n13080, n13081, n13082, n13083, n13084, n13085,
    n13086, n13087, n13088, n13089, n13090, n13091,
    n13092, n13093, n13094, n13095, n13096, n13097,
    n13098, n13099, n13100, n13101, n13102, n13103,
    n13104, n13105, n13106, n13107, n13108, n13109,
    n13110, n13111, n13112, n13113, n13114, n13115,
    n13116, n13117, n13118, n13119, n13120, n13121,
    n13122, n13123, n13124, n13125, n13126, n13127,
    n13128, n13129, n13130, n13131, n13132, n13133,
    n13134, n13135, n13136, n13137, n13138, n13139,
    n13140, n13141, n13142, n13143, n13144, n13145,
    n13146, n13147, n13148, n13149, n13150, n13151,
    n13152, n13153, n13154, n13155, n13156, n13157,
    n13158, n13159, n13160, n13161, n13162, n13163,
    n13164, n13165, n13166, n13167, n13168, n13169,
    n13170, n13171, n13172, n13173, n13174, n13175,
    n13176, n13177, n13178, n13179, n13180, n13181,
    n13182, n13183, n13184, n13185, n13186, n13187,
    n13188, n13189, n13190, n13191, n13192, n13193,
    n13194, n13195, n13196, n13197, n13198, n13199,
    n13200, n13201, n13202, n13203, n13204, n13205,
    n13206, n13207, n13208, n13209, n13210, n13211,
    n13212, n13213, n13214, n13215, n13216, n13217,
    n13218, n13219, n13220, n13221, n13222, n13223,
    n13224, n13225, n13226, n13227, n13228, n13229,
    n13230, n13231, n13232, n13233, n13234, n13235,
    n13236, n13237, n13238, n13239, n13240, n13241,
    n13242, n13243, n13244, n13245, n13246, n13247,
    n13248, n13249, n13250, n13251, n13252, n13253,
    n13254, n13255, n13257, n13258, n13259, n13260,
    n13261, n13262, n13263, n13264, n13265, n13266,
    n13267, n13268, n13269, n13270, n13271, n13272,
    n13273, n13274, n13275, n13276, n13277, n13278,
    n13279, n13280, n13281, n13282, n13283, n13284,
    n13285, n13286, n13287, n13288, n13289, n13290,
    n13291, n13292, n13293, n13294, n13295, n13296,
    n13297, n13298, n13299, n13300, n13301, n13302,
    n13303, n13304, n13305, n13306, n13307, n13308,
    n13309, n13310, n13311, n13312, n13313, n13314,
    n13315, n13316, n13317, n13318, n13319, n13320,
    n13321, n13322, n13323, n13324, n13325, n13326,
    n13327, n13328, n13329, n13330, n13331, n13332,
    n13333, n13334, n13335, n13336, n13337, n13338,
    n13339, n13340, n13341, n13342, n13343, n13344,
    n13345, n13346, n13347, n13348, n13349, n13350,
    n13351, n13352, n13353, n13354, n13355, n13356,
    n13357, n13358, n13359, n13360, n13361, n13362,
    n13363, n13364, n13365, n13366, n13367, n13368,
    n13369, n13370, n13371, n13372, n13373, n13374,
    n13375, n13376, n13377, n13378, n13379, n13380,
    n13381, n13382, n13383, n13384, n13385, n13386,
    n13387, n13388, n13389, n13390, n13391, n13392,
    n13393, n13394, n13395, n13396, n13397, n13398,
    n13399, n13400, n13401, n13402, n13403, n13404,
    n13405, n13406, n13407, n13408, n13409, n13410,
    n13411, n13412, n13413, n13414, n13415, n13416,
    n13417, n13418, n13419, n13420, n13421, n13422,
    n13423, n13424, n13425, n13426, n13427, n13428,
    n13429, n13430, n13431, n13432, n13433, n13434,
    n13435, n13436, n13437, n13438, n13439, n13440,
    n13441, n13442, n13443, n13444, n13445, n13446,
    n13447, n13448, n13449, n13450, n13451, n13452,
    n13453, n13454, n13455, n13456, n13457, n13458,
    n13459, n13460, n13461, n13462, n13463, n13464,
    n13465, n13466, n13467, n13468, n13469, n13470,
    n13471, n13472, n13473, n13474, n13475, n13476,
    n13477, n13478, n13479, n13480, n13481, n13482,
    n13483, n13484, n13485, n13486, n13487, n13488,
    n13489, n13490, n13491, n13492, n13493, n13494,
    n13495, n13496, n13497, n13498, n13499, n13500,
    n13501, n13502, n13503, n13504, n13505, n13506,
    n13507, n13508, n13509, n13510, n13511, n13512,
    n13513, n13514, n13515, n13516, n13517, n13518,
    n13519, n13520, n13521, n13522, n13523, n13524,
    n13525, n13526, n13527, n13528, n13529, n13530,
    n13531, n13532, n13533, n13534, n13535, n13536,
    n13537, n13538, n13539, n13540, n13541, n13542,
    n13543, n13544, n13545, n13546, n13547, n13548,
    n13549, n13550, n13551, n13552, n13553, n13554,
    n13555, n13556, n13557, n13558, n13559, n13560,
    n13561, n13562, n13563, n13564, n13565, n13566,
    n13567, n13568, n13569, n13570, n13571, n13572,
    n13573, n13574, n13575, n13576, n13577, n13578,
    n13579, n13580, n13581, n13582, n13583, n13584,
    n13585, n13586, n13587, n13588, n13589, n13590,
    n13591, n13592, n13593, n13594, n13595, n13596,
    n13597, n13598, n13599, n13600, n13601, n13602,
    n13603, n13604, n13605, n13606, n13607, n13608,
    n13610, n13611, n13612, n13613, n13614, n13615,
    n13616, n13617, n13618, n13619, n13620, n13621,
    n13622, n13623, n13624, n13625, n13626, n13627,
    n13628, n13629, n13630, n13631, n13632, n13633,
    n13634, n13635, n13636, n13637, n13638, n13639,
    n13640, n13641, n13642, n13643, n13644, n13645,
    n13646, n13647, n13648, n13649, n13650, n13651,
    n13652, n13653, n13654, n13655, n13656, n13657,
    n13658, n13659, n13660, n13661, n13662, n13663,
    n13664, n13665, n13666, n13667, n13668, n13669,
    n13670, n13671, n13672, n13673, n13674, n13675,
    n13676, n13677, n13678, n13679, n13680, n13681,
    n13682, n13683, n13684, n13685, n13686, n13687,
    n13688, n13689, n13690, n13691, n13692, n13693,
    n13694, n13695, n13696, n13697, n13698, n13699,
    n13700, n13701, n13702, n13703, n13704, n13705,
    n13706, n13707, n13708, n13709, n13710, n13711,
    n13712, n13713, n13714, n13715, n13716, n13717,
    n13718, n13719, n13720, n13721, n13722, n13723,
    n13724, n13725, n13726, n13727, n13728, n13729,
    n13730, n13731, n13732, n13733, n13734, n13735,
    n13736, n13737, n13738, n13739, n13740, n13741,
    n13742, n13743, n13744, n13745, n13746, n13747,
    n13748, n13749, n13750, n13751, n13752, n13753,
    n13754, n13755, n13756, n13757, n13758, n13759,
    n13760, n13761, n13762, n13763, n13764, n13765,
    n13766, n13767, n13768, n13769, n13770, n13771,
    n13772, n13773, n13774, n13775, n13776, n13777,
    n13778, n13779, n13780, n13781, n13782, n13783,
    n13784, n13785, n13786, n13787, n13788, n13789,
    n13790, n13791, n13792, n13793, n13794, n13795,
    n13796, n13797, n13798, n13799, n13800, n13801,
    n13802, n13803, n13804, n13805, n13806, n13807,
    n13808, n13809, n13810, n13811, n13812, n13813,
    n13814, n13815, n13816, n13817, n13818, n13819,
    n13820, n13821, n13822, n13823, n13824, n13825,
    n13826, n13827, n13828, n13829, n13830, n13831,
    n13832, n13833, n13834, n13835, n13836, n13837,
    n13838, n13839, n13840, n13841, n13842, n13843,
    n13844, n13845, n13846, n13847, n13848, n13849,
    n13850, n13851, n13852, n13853, n13854, n13855,
    n13856, n13857, n13858, n13859, n13860, n13861,
    n13862, n13863, n13864, n13865, n13866, n13867,
    n13868, n13869, n13870, n13871, n13872, n13873,
    n13874, n13875, n13876, n13877, n13878, n13879,
    n13880, n13881, n13882, n13883, n13884, n13885,
    n13886, n13887, n13888, n13889, n13890, n13891,
    n13892, n13893, n13894, n13895, n13896, n13897,
    n13898, n13899, n13900, n13901, n13902, n13903,
    n13904, n13905, n13906, n13907, n13908, n13909,
    n13910, n13911, n13912, n13913, n13914, n13915,
    n13916, n13917, n13918, n13919, n13920, n13921,
    n13922, n13923, n13924, n13925, n13926, n13927,
    n13928, n13929, n13930, n13931, n13932, n13933,
    n13934, n13935, n13936, n13937, n13938, n13939,
    n13940, n13941, n13942, n13943, n13944, n13945,
    n13946, n13947, n13948, n13949, n13950, n13951,
    n13952, n13953, n13954, n13955, n13956, n13957,
    n13958, n13959, n13960, n13961, n13962, n13963,
    n13965, n13966, n13967, n13968, n13969, n13970,
    n13971, n13972, n13973, n13974, n13975, n13976,
    n13977, n13978, n13979, n13980, n13981, n13982,
    n13983, n13984, n13985, n13986, n13987, n13988,
    n13989, n13990, n13991, n13992, n13993, n13994,
    n13995, n13996, n13997, n13998, n13999, n14000,
    n14001, n14002, n14003, n14004, n14005, n14006,
    n14007, n14008, n14009, n14010, n14011, n14012,
    n14013, n14014, n14015, n14016, n14017, n14018,
    n14019, n14020, n14021, n14022, n14023, n14024,
    n14025, n14026, n14027, n14028, n14029, n14030,
    n14031, n14032, n14033, n14034, n14035, n14036,
    n14037, n14038, n14039, n14040, n14041, n14042,
    n14043, n14044, n14045, n14046, n14047, n14048,
    n14049, n14050, n14051, n14052, n14053, n14054,
    n14055, n14056, n14057, n14058, n14059, n14060,
    n14061, n14062, n14063, n14064, n14065, n14066,
    n14067, n14068, n14069, n14070, n14071, n14072,
    n14073, n14074, n14075, n14076, n14077, n14078,
    n14079, n14080, n14081, n14082, n14083, n14084,
    n14085, n14086, n14087, n14088, n14089, n14090,
    n14091, n14092, n14093, n14094, n14095, n14096,
    n14097, n14098, n14099, n14100, n14101, n14102,
    n14103, n14104, n14105, n14106, n14107, n14108,
    n14109, n14110, n14111, n14112, n14113, n14114,
    n14115, n14116, n14117, n14118, n14119, n14120,
    n14121, n14122, n14123, n14124, n14125, n14126,
    n14127, n14128, n14129, n14130, n14131, n14132,
    n14133, n14134, n14135, n14136, n14137, n14138,
    n14139, n14140, n14141, n14142, n14143, n14144,
    n14145, n14146, n14147, n14148, n14149, n14150,
    n14151, n14152, n14153, n14154, n14155, n14156,
    n14157, n14158, n14159, n14160, n14161, n14162,
    n14163, n14164, n14165, n14166, n14167, n14168,
    n14169, n14170, n14171, n14172, n14173, n14174,
    n14175, n14176, n14177, n14178, n14179, n14180,
    n14181, n14182, n14183, n14184, n14185, n14186,
    n14187, n14188, n14189, n14190, n14191, n14192,
    n14193, n14194, n14195, n14196, n14197, n14198,
    n14199, n14200, n14201, n14202, n14203, n14204,
    n14205, n14206, n14207, n14208, n14209, n14210,
    n14211, n14212, n14213, n14214, n14215, n14216,
    n14217, n14218, n14219, n14220, n14221, n14222,
    n14223, n14224, n14225, n14226, n14227, n14228,
    n14229, n14230, n14231, n14232, n14233, n14234,
    n14235, n14236, n14237, n14238, n14239, n14240,
    n14241, n14242, n14243, n14244, n14245, n14246,
    n14247, n14248, n14249, n14250, n14251, n14252,
    n14253, n14254, n14255, n14256, n14257, n14258,
    n14259, n14260, n14261, n14262, n14263, n14264,
    n14265, n14266, n14267, n14268, n14269, n14270,
    n14271, n14272, n14273, n14274, n14275, n14276,
    n14277, n14278, n14279, n14280, n14281, n14282,
    n14283, n14284, n14285, n14286, n14287, n14288,
    n14289, n14290, n14291, n14292, n14293, n14294,
    n14295, n14296, n14297, n14298, n14299, n14300,
    n14301, n14302, n14303, n14304, n14305, n14306,
    n14307, n14308, n14309, n14310, n14311, n14312,
    n14313, n14314, n14315, n14317, n14318, n14319,
    n14320, n14321, n14322, n14323, n14324, n14325,
    n14326, n14327, n14328, n14329, n14330, n14331,
    n14332, n14333, n14334, n14335, n14336, n14337,
    n14338, n14339, n14340, n14341, n14342, n14343,
    n14344, n14345, n14346, n14347, n14348, n14349,
    n14350, n14351, n14352, n14353, n14354, n14355,
    n14356, n14357, n14358, n14359, n14360, n14361,
    n14362, n14363, n14364, n14365, n14366, n14367,
    n14368, n14369, n14370, n14371, n14372, n14373,
    n14374, n14375, n14376, n14377, n14378, n14379,
    n14380, n14381, n14382, n14383, n14384, n14385,
    n14386, n14387, n14388, n14389, n14390, n14391,
    n14392, n14393, n14394, n14395, n14396, n14397,
    n14398, n14399, n14400, n14401, n14402, n14403,
    n14404, n14405, n14406, n14407, n14408, n14409,
    n14410, n14411, n14412, n14413, n14414, n14415,
    n14416, n14417, n14418, n14419, n14420, n14421,
    n14422, n14423, n14424, n14425, n14426, n14427,
    n14428, n14429, n14430, n14431, n14432, n14433,
    n14434, n14435, n14436, n14437, n14438, n14439,
    n14440, n14441, n14442, n14443, n14444, n14445,
    n14446, n14447, n14448, n14449, n14450, n14451,
    n14452, n14453, n14454, n14455, n14456, n14457,
    n14458, n14459, n14460, n14461, n14462, n14463,
    n14464, n14465, n14466, n14467, n14468, n14469,
    n14470, n14471, n14472, n14473, n14474, n14475,
    n14476, n14477, n14478, n14479, n14480, n14481,
    n14482, n14483, n14484, n14485, n14486, n14487,
    n14488, n14489, n14490, n14491, n14492, n14493,
    n14494, n14495, n14496, n14497, n14498, n14499,
    n14500, n14501, n14502, n14503, n14504, n14505,
    n14506, n14507, n14508, n14509, n14510, n14511,
    n14512, n14513, n14514, n14515, n14516, n14517,
    n14518, n14519, n14520, n14521, n14522, n14523,
    n14524, n14525, n14526, n14527, n14528, n14529,
    n14530, n14531, n14532, n14533, n14534, n14535,
    n14536, n14537, n14538, n14539, n14540, n14541,
    n14542, n14543, n14544, n14545, n14546, n14547,
    n14548, n14549, n14550, n14551, n14552, n14553,
    n14554, n14555, n14556, n14557, n14558, n14559,
    n14560, n14561, n14562, n14563, n14564, n14565,
    n14566, n14567, n14568, n14569, n14570, n14571,
    n14572, n14573, n14574, n14575, n14576, n14577,
    n14578, n14579, n14580, n14581, n14582, n14583,
    n14584, n14585, n14586, n14587, n14588, n14589,
    n14590, n14591, n14592, n14593, n14594, n14595,
    n14596, n14597, n14598, n14599, n14600, n14601,
    n14602, n14603, n14604, n14605, n14606, n14607,
    n14608, n14609, n14610, n14611, n14612, n14613,
    n14614, n14615, n14616, n14617, n14618, n14619,
    n14620, n14621, n14622, n14623, n14624, n14625,
    n14626, n14627, n14628, n14629, n14630, n14631,
    n14632, n14633, n14634, n14635, n14636, n14637,
    n14638, n14639, n14640, n14641, n14642, n14643,
    n14644, n14645, n14646, n14647, n14648, n14649,
    n14650, n14651, n14652, n14653, n14654, n14655,
    n14656, n14657, n14658, n14659, n14660, n14661,
    n14662, n14663, n14665, n14666, n14667, n14668,
    n14669, n14670, n14671, n14672, n14673, n14674,
    n14675, n14676, n14677, n14678, n14679, n14680,
    n14681, n14682, n14683, n14684, n14685, n14686,
    n14687, n14688, n14689, n14690, n14691, n14692,
    n14693, n14694, n14695, n14696, n14697, n14698,
    n14699, n14700, n14701, n14702, n14703, n14704,
    n14705, n14706, n14707, n14708, n14709, n14710,
    n14711, n14712, n14713, n14714, n14715, n14716,
    n14717, n14718, n14719, n14720, n14721, n14722,
    n14723, n14724, n14725, n14726, n14727, n14728,
    n14729, n14730, n14731, n14732, n14733, n14734,
    n14735, n14736, n14737, n14738, n14739, n14740,
    n14741, n14742, n14743, n14744, n14745, n14746,
    n14747, n14748, n14749, n14750, n14751, n14752,
    n14753, n14754, n14755, n14756, n14757, n14758,
    n14759, n14760, n14761, n14762, n14763, n14764,
    n14765, n14766, n14767, n14768, n14769, n14770,
    n14771, n14772, n14773, n14774, n14775, n14776,
    n14777, n14778, n14779, n14780, n14781, n14782,
    n14783, n14784, n14785, n14786, n14787, n14788,
    n14789, n14790, n14791, n14792, n14793, n14794,
    n14795, n14796, n14797, n14798, n14799, n14800,
    n14801, n14802, n14803, n14804, n14805, n14806,
    n14807, n14808, n14809, n14810, n14811, n14812,
    n14813, n14814, n14815, n14816, n14817, n14818,
    n14819, n14820, n14821, n14822, n14823, n14824,
    n14825, n14826, n14827, n14828, n14829, n14830,
    n14831, n14832, n14833, n14834, n14835, n14836,
    n14837, n14838, n14839, n14840, n14841, n14842,
    n14843, n14844, n14845, n14846, n14847, n14848,
    n14849, n14850, n14851, n14852, n14853, n14854,
    n14855, n14856, n14857, n14858, n14859, n14860,
    n14861, n14862, n14863, n14864, n14865, n14866,
    n14867, n14868, n14869, n14870, n14871, n14872,
    n14873, n14874, n14875, n14876, n14877, n14878,
    n14879, n14880, n14881, n14882, n14883, n14884,
    n14885, n14886, n14887, n14888, n14889, n14890,
    n14891, n14892, n14893, n14894, n14895, n14896,
    n14897, n14898, n14899, n14900, n14901, n14902,
    n14903, n14904, n14905, n14906, n14907, n14908,
    n14909, n14910, n14911, n14912, n14913, n14914,
    n14915, n14916, n14917, n14918, n14919, n14920,
    n14921, n14922, n14923, n14924, n14925, n14926,
    n14927, n14928, n14929, n14930, n14931, n14932,
    n14933, n14934, n14935, n14936, n14937, n14938,
    n14939, n14940, n14941, n14942, n14943, n14944,
    n14945, n14946, n14947, n14948, n14949, n14950,
    n14951, n14952, n14953, n14954, n14955, n14956,
    n14957, n14958, n14959, n14960, n14961, n14962,
    n14963, n14964, n14965, n14966, n14967, n14968,
    n14969, n14970, n14971, n14972, n14973, n14974,
    n14975, n14976, n14977, n14978, n14979, n14980,
    n14981, n14982, n14983, n14984, n14985, n14986,
    n14987, n14988, n14989, n14990, n14991, n14992,
    n14993, n14994, n14995, n14996, n14997, n14998,
    n15000, n15001, n15002, n15003, n15004, n15005,
    n15006, n15007, n15008, n15009, n15010, n15011,
    n15012, n15013, n15014, n15015, n15016, n15017,
    n15018, n15019, n15020, n15021, n15022, n15023,
    n15024, n15025, n15026, n15027, n15028, n15029,
    n15030, n15031, n15032, n15033, n15034, n15035,
    n15036, n15037, n15038, n15039, n15040, n15041,
    n15042, n15043, n15044, n15045, n15046, n15047,
    n15048, n15049, n15050, n15051, n15052, n15053,
    n15054, n15055, n15056, n15057, n15058, n15059,
    n15060, n15061, n15062, n15063, n15064, n15065,
    n15066, n15067, n15068, n15069, n15070, n15071,
    n15072, n15073, n15074, n15075, n15076, n15077,
    n15078, n15079, n15080, n15081, n15082, n15083,
    n15084, n15085, n15086, n15087, n15088, n15089,
    n15090, n15091, n15092, n15093, n15094, n15095,
    n15096, n15097, n15098, n15099, n15100, n15101,
    n15102, n15103, n15104, n15105, n15106, n15107,
    n15108, n15109, n15110, n15111, n15112, n15113,
    n15114, n15115, n15116, n15117, n15118, n15119,
    n15120, n15121, n15122, n15123, n15124, n15125,
    n15126, n15127, n15128, n15129, n15130, n15131,
    n15132, n15133, n15134, n15135, n15136, n15137,
    n15138, n15139, n15140, n15141, n15142, n15143,
    n15144, n15145, n15146, n15147, n15148, n15149,
    n15150, n15151, n15152, n15153, n15154, n15155,
    n15156, n15157, n15158, n15159, n15160, n15161,
    n15162, n15163, n15164, n15165, n15166, n15167,
    n15168, n15169, n15170, n15171, n15172, n15173,
    n15174, n15175, n15176, n15177, n15178, n15179,
    n15180, n15181, n15182, n15183, n15184, n15185,
    n15186, n15187, n15188, n15189, n15190, n15191,
    n15192, n15193, n15194, n15195, n15196, n15197,
    n15198, n15199, n15200, n15201, n15202, n15203,
    n15204, n15205, n15206, n15207, n15208, n15209,
    n15210, n15211, n15212, n15213, n15214, n15215,
    n15216, n15217, n15218, n15219, n15220, n15221,
    n15222, n15223, n15224, n15225, n15226, n15227,
    n15228, n15229, n15230, n15231, n15232, n15233,
    n15234, n15235, n15236, n15237, n15238, n15239,
    n15240, n15241, n15242, n15243, n15244, n15245,
    n15246, n15247, n15248, n15249, n15250, n15251,
    n15252, n15253, n15254, n15255, n15256, n15257,
    n15258, n15259, n15260, n15261, n15262, n15263,
    n15264, n15265, n15266, n15267, n15268, n15269,
    n15270, n15271, n15272, n15273, n15274, n15275,
    n15276, n15277, n15278, n15279, n15280, n15281,
    n15282, n15283, n15284, n15285, n15286, n15287,
    n15288, n15289, n15290, n15291, n15292, n15293,
    n15294, n15295, n15296, n15297, n15298, n15299,
    n15300, n15301, n15302, n15303, n15304, n15305,
    n15306, n15307, n15308, n15309, n15310, n15311,
    n15312, n15313, n15314, n15315, n15316, n15317,
    n15318, n15319, n15320, n15321, n15322, n15323,
    n15324, n15325, n15326, n15327, n15328, n15329,
    n15330, n15331, n15332, n15333, n15334, n15335,
    n15336, n15338, n15339, n15340, n15341, n15342,
    n15343, n15344, n15345, n15346, n15347, n15348,
    n15349, n15350, n15351, n15352, n15353, n15354,
    n15355, n15356, n15357, n15358, n15359, n15360,
    n15361, n15362, n15363, n15364, n15365, n15366,
    n15367, n15368, n15369, n15370, n15371, n15372,
    n15373, n15374, n15375, n15376, n15377, n15378,
    n15379, n15380, n15381, n15382, n15383, n15384,
    n15385, n15386, n15387, n15388, n15389, n15390,
    n15391, n15392, n15393, n15394, n15395, n15396,
    n15397, n15398, n15399, n15400, n15401, n15402,
    n15403, n15404, n15405, n15406, n15407, n15408,
    n15409, n15410, n15411, n15412, n15413, n15414,
    n15415, n15416, n15417, n15418, n15419, n15420,
    n15421, n15422, n15423, n15424, n15425, n15426,
    n15427, n15428, n15429, n15430, n15431, n15432,
    n15433, n15434, n15435, n15436, n15437, n15438,
    n15439, n15440, n15441, n15442, n15443, n15444,
    n15445, n15446, n15447, n15448, n15449, n15450,
    n15451, n15452, n15453, n15454, n15455, n15456,
    n15457, n15458, n15459, n15460, n15461, n15462,
    n15463, n15464, n15465, n15466, n15467, n15468,
    n15469, n15470, n15471, n15472, n15473, n15474,
    n15475, n15476, n15477, n15478, n15479, n15480,
    n15481, n15482, n15483, n15484, n15485, n15486,
    n15487, n15488, n15489, n15490, n15491, n15492,
    n15493, n15494, n15495, n15496, n15497, n15498,
    n15499, n15500, n15501, n15502, n15503, n15504,
    n15505, n15506, n15507, n15508, n15509, n15510,
    n15511, n15512, n15513, n15514, n15515, n15516,
    n15517, n15518, n15519, n15520, n15521, n15522,
    n15523, n15524, n15525, n15526, n15527, n15528,
    n15529, n15530, n15531, n15532, n15533, n15534,
    n15535, n15536, n15537, n15538, n15539, n15540,
    n15541, n15542, n15543, n15544, n15545, n15546,
    n15547, n15548, n15549, n15550, n15551, n15552,
    n15553, n15554, n15555, n15556, n15557, n15558,
    n15559, n15560, n15561, n15562, n15563, n15564,
    n15565, n15566, n15567, n15568, n15569, n15570,
    n15571, n15572, n15573, n15574, n15575, n15576,
    n15577, n15578, n15579, n15580, n15581, n15582,
    n15583, n15584, n15585, n15586, n15587, n15588,
    n15589, n15590, n15591, n15592, n15593, n15594,
    n15595, n15596, n15597, n15598, n15599, n15600,
    n15601, n15602, n15603, n15604, n15605, n15606,
    n15607, n15608, n15609, n15610, n15611, n15612,
    n15613, n15614, n15615, n15616, n15617, n15618,
    n15619, n15620, n15621, n15622, n15623, n15624,
    n15625, n15626, n15627, n15628, n15629, n15630,
    n15631, n15632, n15633, n15634, n15635, n15636,
    n15637, n15638, n15639, n15640, n15641, n15642,
    n15643, n15644, n15645, n15646, n15647, n15648,
    n15649, n15650, n15651, n15652, n15653, n15654,
    n15655, n15656, n15657, n15658, n15659, n15660,
    n15661, n15662, n15663, n15664, n15666, n15667,
    n15668, n15669, n15670, n15671, n15672, n15673,
    n15674, n15675, n15676, n15677, n15678, n15679,
    n15680, n15681, n15682, n15683, n15684, n15685,
    n15686, n15687, n15688, n15689, n15690, n15691,
    n15692, n15693, n15694, n15695, n15696, n15697,
    n15698, n15699, n15700, n15701, n15702, n15703,
    n15704, n15705, n15706, n15707, n15708, n15709,
    n15710, n15711, n15712, n15713, n15714, n15715,
    n15716, n15717, n15718, n15719, n15720, n15721,
    n15722, n15723, n15724, n15725, n15726, n15727,
    n15728, n15729, n15730, n15731, n15732, n15733,
    n15734, n15735, n15736, n15737, n15738, n15739,
    n15740, n15741, n15742, n15743, n15744, n15745,
    n15746, n15747, n15748, n15749, n15750, n15751,
    n15752, n15753, n15754, n15755, n15756, n15757,
    n15758, n15759, n15760, n15761, n15762, n15763,
    n15764, n15765, n15766, n15767, n15768, n15769,
    n15770, n15771, n15772, n15773, n15774, n15775,
    n15776, n15777, n15778, n15779, n15780, n15781,
    n15782, n15783, n15784, n15785, n15786, n15787,
    n15788, n15789, n15790, n15791, n15792, n15793,
    n15794, n15795, n15796, n15797, n15798, n15799,
    n15800, n15801, n15802, n15803, n15804, n15805,
    n15806, n15807, n15808, n15809, n15810, n15811,
    n15812, n15813, n15814, n15815, n15816, n15817,
    n15818, n15819, n15820, n15821, n15822, n15823,
    n15824, n15825, n15826, n15827, n15828, n15829,
    n15830, n15831, n15832, n15833, n15834, n15835,
    n15836, n15837, n15838, n15839, n15840, n15841,
    n15842, n15843, n15844, n15845, n15846, n15847,
    n15848, n15849, n15850, n15851, n15852, n15853,
    n15854, n15855, n15856, n15857, n15858, n15859,
    n15860, n15861, n15862, n15863, n15864, n15865,
    n15866, n15867, n15868, n15869, n15870, n15871,
    n15872, n15873, n15874, n15875, n15876, n15877,
    n15878, n15879, n15880, n15881, n15882, n15883,
    n15884, n15885, n15886, n15887, n15888, n15889,
    n15890, n15891, n15892, n15893, n15894, n15895,
    n15896, n15897, n15898, n15899, n15900, n15901,
    n15902, n15903, n15904, n15905, n15906, n15907,
    n15908, n15909, n15910, n15911, n15912, n15913,
    n15914, n15915, n15916, n15917, n15918, n15919,
    n15920, n15921, n15922, n15923, n15924, n15925,
    n15926, n15927, n15928, n15929, n15930, n15931,
    n15932, n15933, n15934, n15935, n15936, n15937,
    n15938, n15939, n15940, n15941, n15942, n15943,
    n15944, n15945, n15946, n15947, n15948, n15949,
    n15950, n15951, n15952, n15953, n15954, n15955,
    n15956, n15957, n15958, n15959, n15960, n15961,
    n15962, n15963, n15964, n15965, n15966, n15967,
    n15968, n15969, n15970, n15971, n15972, n15973,
    n15974, n15975, n15976, n15977, n15978, n15979,
    n15980, n15981, n15983, n15984, n15985, n15986,
    n15987, n15988, n15989, n15990, n15991, n15992,
    n15993, n15994, n15995, n15996, n15997, n15998,
    n15999, n16000, n16001, n16002, n16003, n16004,
    n16005, n16006, n16007, n16008, n16009, n16010,
    n16011, n16012, n16013, n16014, n16015, n16016,
    n16017, n16018, n16019, n16020, n16021, n16022,
    n16023, n16024, n16025, n16026, n16027, n16028,
    n16029, n16030, n16031, n16032, n16033, n16034,
    n16035, n16036, n16037, n16038, n16039, n16040,
    n16041, n16042, n16043, n16044, n16045, n16046,
    n16047, n16048, n16049, n16050, n16051, n16052,
    n16053, n16054, n16055, n16056, n16057, n16058,
    n16059, n16060, n16061, n16062, n16063, n16064,
    n16065, n16066, n16067, n16068, n16069, n16070,
    n16071, n16072, n16073, n16074, n16075, n16076,
    n16077, n16078, n16079, n16080, n16081, n16082,
    n16083, n16084, n16085, n16086, n16087, n16088,
    n16089, n16090, n16091, n16092, n16093, n16094,
    n16095, n16096, n16097, n16098, n16099, n16100,
    n16101, n16102, n16103, n16104, n16105, n16106,
    n16107, n16108, n16109, n16110, n16111, n16112,
    n16113, n16114, n16115, n16116, n16117, n16118,
    n16119, n16120, n16121, n16122, n16123, n16124,
    n16125, n16126, n16127, n16128, n16129, n16130,
    n16131, n16132, n16133, n16134, n16135, n16136,
    n16137, n16138, n16139, n16140, n16141, n16142,
    n16143, n16144, n16145, n16146, n16147, n16148,
    n16149, n16150, n16151, n16152, n16153, n16154,
    n16155, n16156, n16157, n16158, n16159, n16160,
    n16161, n16162, n16163, n16164, n16165, n16166,
    n16167, n16168, n16169, n16170, n16171, n16172,
    n16173, n16174, n16175, n16176, n16177, n16178,
    n16179, n16180, n16181, n16182, n16183, n16184,
    n16185, n16186, n16187, n16188, n16189, n16190,
    n16191, n16192, n16193, n16194, n16195, n16196,
    n16197, n16198, n16199, n16200, n16201, n16202,
    n16203, n16204, n16205, n16206, n16207, n16208,
    n16209, n16210, n16211, n16212, n16213, n16214,
    n16215, n16216, n16217, n16218, n16219, n16220,
    n16221, n16222, n16223, n16224, n16225, n16226,
    n16227, n16228, n16229, n16230, n16231, n16232,
    n16233, n16234, n16235, n16236, n16237, n16238,
    n16239, n16240, n16241, n16242, n16243, n16244,
    n16245, n16246, n16247, n16248, n16249, n16250,
    n16251, n16252, n16253, n16254, n16255, n16256,
    n16257, n16258, n16259, n16260, n16261, n16262,
    n16263, n16264, n16265, n16266, n16267, n16268,
    n16269, n16270, n16271, n16272, n16273, n16274,
    n16275, n16276, n16277, n16278, n16279, n16280,
    n16281, n16282, n16283, n16284, n16285, n16286,
    n16287, n16288, n16289, n16290, n16291, n16292,
    n16293, n16294, n16295, n16296, n16297, n16298,
    n16299, n16300, n16301, n16303, n16304, n16305,
    n16306, n16307, n16308, n16309, n16310, n16311,
    n16312, n16313, n16314, n16315, n16316, n16317,
    n16318, n16319, n16320, n16321, n16322, n16323,
    n16324, n16325, n16326, n16327, n16328, n16329,
    n16330, n16331, n16332, n16333, n16334, n16335,
    n16336, n16337, n16338, n16339, n16340, n16341,
    n16342, n16343, n16344, n16345, n16346, n16347,
    n16348, n16349, n16350, n16351, n16352, n16353,
    n16354, n16355, n16356, n16357, n16358, n16359,
    n16360, n16361, n16362, n16363, n16364, n16365,
    n16366, n16367, n16368, n16369, n16370, n16371,
    n16372, n16373, n16374, n16375, n16376, n16377,
    n16378, n16379, n16380, n16381, n16382, n16383,
    n16384, n16385, n16386, n16387, n16388, n16389,
    n16390, n16391, n16392, n16393, n16394, n16395,
    n16396, n16397, n16398, n16399, n16400, n16401,
    n16402, n16403, n16404, n16405, n16406, n16407,
    n16408, n16409, n16410, n16411, n16412, n16413,
    n16414, n16415, n16416, n16417, n16418, n16419,
    n16420, n16421, n16422, n16423, n16424, n16425,
    n16426, n16427, n16428, n16429, n16430, n16431,
    n16432, n16433, n16434, n16435, n16436, n16437,
    n16438, n16439, n16440, n16441, n16442, n16443,
    n16444, n16445, n16446, n16447, n16448, n16449,
    n16450, n16451, n16452, n16453, n16454, n16455,
    n16456, n16457, n16458, n16459, n16460, n16461,
    n16462, n16463, n16464, n16465, n16466, n16467,
    n16468, n16469, n16470, n16471, n16472, n16473,
    n16474, n16475, n16476, n16477, n16478, n16479,
    n16480, n16481, n16482, n16483, n16484, n16485,
    n16486, n16487, n16488, n16489, n16490, n16491,
    n16492, n16493, n16494, n16495, n16496, n16497,
    n16498, n16499, n16500, n16501, n16502, n16503,
    n16504, n16505, n16506, n16507, n16508, n16509,
    n16510, n16511, n16512, n16513, n16514, n16515,
    n16516, n16517, n16518, n16519, n16520, n16521,
    n16522, n16523, n16524, n16525, n16526, n16527,
    n16528, n16529, n16530, n16531, n16532, n16533,
    n16534, n16535, n16536, n16537, n16538, n16539,
    n16540, n16541, n16542, n16543, n16544, n16545,
    n16546, n16547, n16548, n16549, n16550, n16551,
    n16552, n16553, n16554, n16555, n16556, n16557,
    n16558, n16559, n16560, n16561, n16562, n16563,
    n16564, n16565, n16566, n16567, n16568, n16569,
    n16570, n16571, n16572, n16573, n16574, n16575,
    n16576, n16577, n16578, n16579, n16580, n16581,
    n16582, n16583, n16584, n16585, n16586, n16587,
    n16588, n16589, n16590, n16591, n16592, n16593,
    n16594, n16595, n16596, n16597, n16598, n16599,
    n16600, n16601, n16602, n16603, n16604, n16605,
    n16606, n16607, n16608, n16609, n16610, n16611,
    n16612, n16614, n16615, n16616, n16617, n16618,
    n16619, n16620, n16621, n16622, n16623, n16624,
    n16625, n16626, n16627, n16628, n16629, n16630,
    n16631, n16632, n16633, n16634, n16635, n16636,
    n16637, n16638, n16639, n16640, n16641, n16642,
    n16643, n16644, n16645, n16646, n16647, n16648,
    n16649, n16650, n16651, n16652, n16653, n16654,
    n16655, n16656, n16657, n16658, n16659, n16660,
    n16661, n16662, n16663, n16664, n16665, n16666,
    n16667, n16668, n16669, n16670, n16671, n16672,
    n16673, n16674, n16675, n16676, n16677, n16678,
    n16679, n16680, n16681, n16682, n16683, n16684,
    n16685, n16686, n16687, n16688, n16689, n16690,
    n16691, n16692, n16693, n16694, n16695, n16696,
    n16697, n16698, n16699, n16700, n16701, n16702,
    n16703, n16704, n16705, n16706, n16707, n16708,
    n16709, n16710, n16711, n16712, n16713, n16714,
    n16715, n16716, n16717, n16718, n16719, n16720,
    n16721, n16722, n16723, n16724, n16725, n16726,
    n16727, n16728, n16729, n16730, n16731, n16732,
    n16733, n16734, n16735, n16736, n16737, n16738,
    n16739, n16740, n16741, n16742, n16743, n16744,
    n16745, n16746, n16747, n16748, n16749, n16750,
    n16751, n16752, n16753, n16754, n16755, n16756,
    n16757, n16758, n16759, n16760, n16761, n16762,
    n16763, n16764, n16765, n16766, n16767, n16768,
    n16769, n16770, n16771, n16772, n16773, n16774,
    n16775, n16776, n16777, n16778, n16779, n16780,
    n16781, n16782, n16783, n16784, n16785, n16786,
    n16787, n16788, n16789, n16790, n16791, n16792,
    n16793, n16794, n16795, n16796, n16797, n16798,
    n16799, n16800, n16801, n16802, n16803, n16804,
    n16805, n16806, n16807, n16808, n16809, n16810,
    n16811, n16812, n16813, n16814, n16815, n16816,
    n16817, n16818, n16819, n16820, n16821, n16822,
    n16823, n16824, n16825, n16826, n16827, n16828,
    n16829, n16830, n16831, n16832, n16833, n16834,
    n16835, n16836, n16837, n16838, n16839, n16840,
    n16841, n16842, n16843, n16844, n16845, n16846,
    n16847, n16848, n16849, n16850, n16851, n16852,
    n16853, n16854, n16855, n16856, n16857, n16858,
    n16859, n16860, n16861, n16862, n16863, n16864,
    n16865, n16866, n16867, n16868, n16869, n16870,
    n16871, n16872, n16873, n16874, n16875, n16876,
    n16877, n16878, n16879, n16880, n16881, n16882,
    n16883, n16884, n16885, n16886, n16887, n16888,
    n16889, n16890, n16891, n16892, n16893, n16894,
    n16895, n16896, n16897, n16898, n16899, n16900,
    n16901, n16902, n16903, n16904, n16905, n16906,
    n16907, n16908, n16909, n16910, n16911, n16913,
    n16914, n16915, n16916, n16917, n16918, n16919,
    n16920, n16921, n16922, n16923, n16924, n16925,
    n16926, n16927, n16928, n16929, n16930, n16931,
    n16932, n16933, n16934, n16935, n16936, n16937,
    n16938, n16939, n16940, n16941, n16942, n16943,
    n16944, n16945, n16946, n16947, n16948, n16949,
    n16950, n16951, n16952, n16953, n16954, n16955,
    n16956, n16957, n16958, n16959, n16960, n16961,
    n16962, n16963, n16964, n16965, n16966, n16967,
    n16968, n16969, n16970, n16971, n16972, n16973,
    n16974, n16975, n16976, n16977, n16978, n16979,
    n16980, n16981, n16982, n16983, n16984, n16985,
    n16986, n16987, n16988, n16989, n16990, n16991,
    n16992, n16993, n16994, n16995, n16996, n16997,
    n16998, n16999, n17000, n17001, n17002, n17003,
    n17004, n17005, n17006, n17007, n17008, n17009,
    n17010, n17011, n17012, n17013, n17014, n17015,
    n17016, n17017, n17018, n17019, n17020, n17021,
    n17022, n17023, n17024, n17025, n17026, n17027,
    n17028, n17029, n17030, n17031, n17032, n17033,
    n17034, n17035, n17036, n17037, n17038, n17039,
    n17040, n17041, n17042, n17043, n17044, n17045,
    n17046, n17047, n17048, n17049, n17050, n17051,
    n17052, n17053, n17054, n17055, n17056, n17057,
    n17058, n17059, n17060, n17061, n17062, n17063,
    n17064, n17065, n17066, n17067, n17068, n17069,
    n17070, n17071, n17072, n17073, n17074, n17075,
    n17076, n17077, n17078, n17079, n17080, n17081,
    n17082, n17083, n17084, n17085, n17086, n17087,
    n17088, n17089, n17090, n17091, n17092, n17093,
    n17094, n17095, n17096, n17097, n17098, n17099,
    n17100, n17101, n17102, n17103, n17104, n17105,
    n17106, n17107, n17108, n17109, n17110, n17111,
    n17112, n17113, n17114, n17115, n17116, n17117,
    n17118, n17119, n17120, n17121, n17122, n17123,
    n17124, n17125, n17126, n17127, n17128, n17129,
    n17130, n17131, n17132, n17133, n17134, n17135,
    n17136, n17137, n17138, n17139, n17140, n17141,
    n17142, n17143, n17144, n17145, n17146, n17147,
    n17148, n17149, n17150, n17151, n17152, n17153,
    n17154, n17155, n17156, n17157, n17158, n17159,
    n17160, n17161, n17162, n17163, n17164, n17165,
    n17166, n17167, n17168, n17169, n17170, n17171,
    n17172, n17173, n17174, n17175, n17176, n17177,
    n17178, n17179, n17180, n17181, n17182, n17183,
    n17184, n17185, n17186, n17187, n17188, n17189,
    n17190, n17191, n17192, n17193, n17194, n17195,
    n17196, n17197, n17198, n17199, n17200, n17201,
    n17202, n17203, n17204, n17205, n17206, n17207,
    n17208, n17209, n17210, n17211, n17213, n17214,
    n17215, n17216, n17217, n17218, n17219, n17220,
    n17221, n17222, n17223, n17224, n17225, n17226,
    n17227, n17228, n17229, n17230, n17231, n17232,
    n17233, n17234, n17235, n17236, n17237, n17238,
    n17239, n17240, n17241, n17242, n17243, n17244,
    n17245, n17246, n17247, n17248, n17249, n17250,
    n17251, n17252, n17253, n17254, n17255, n17256,
    n17257, n17258, n17259, n17260, n17261, n17262,
    n17263, n17264, n17265, n17266, n17267, n17268,
    n17269, n17270, n17271, n17272, n17273, n17274,
    n17275, n17276, n17277, n17278, n17279, n17280,
    n17281, n17282, n17283, n17284, n17285, n17286,
    n17287, n17288, n17289, n17290, n17291, n17292,
    n17293, n17294, n17295, n17296, n17297, n17298,
    n17299, n17300, n17301, n17302, n17303, n17304,
    n17305, n17306, n17307, n17308, n17309, n17310,
    n17311, n17312, n17313, n17314, n17315, n17316,
    n17317, n17318, n17319, n17320, n17321, n17322,
    n17323, n17324, n17325, n17326, n17327, n17328,
    n17329, n17330, n17331, n17332, n17333, n17334,
    n17335, n17336, n17337, n17338, n17339, n17340,
    n17341, n17342, n17343, n17344, n17345, n17346,
    n17347, n17348, n17349, n17350, n17351, n17352,
    n17353, n17354, n17355, n17356, n17357, n17358,
    n17359, n17360, n17361, n17362, n17363, n17364,
    n17365, n17366, n17367, n17368, n17369, n17370,
    n17371, n17372, n17373, n17374, n17375, n17376,
    n17377, n17378, n17379, n17380, n17381, n17382,
    n17383, n17384, n17385, n17386, n17387, n17388,
    n17389, n17390, n17391, n17392, n17393, n17394,
    n17395, n17396, n17397, n17398, n17399, n17400,
    n17401, n17402, n17403, n17404, n17405, n17406,
    n17407, n17408, n17409, n17410, n17411, n17412,
    n17413, n17414, n17415, n17416, n17417, n17418,
    n17419, n17420, n17421, n17422, n17423, n17424,
    n17425, n17426, n17427, n17428, n17429, n17430,
    n17431, n17432, n17433, n17434, n17435, n17436,
    n17437, n17438, n17439, n17440, n17441, n17442,
    n17443, n17444, n17445, n17446, n17447, n17448,
    n17449, n17450, n17451, n17452, n17453, n17454,
    n17455, n17456, n17457, n17458, n17459, n17460,
    n17461, n17462, n17463, n17464, n17465, n17466,
    n17467, n17468, n17469, n17470, n17471, n17472,
    n17473, n17474, n17475, n17476, n17477, n17478,
    n17479, n17480, n17481, n17482, n17483, n17484,
    n17485, n17486, n17487, n17488, n17489, n17490,
    n17491, n17492, n17493, n17494, n17495, n17496,
    n17497, n17498, n17499, n17500, n17501, n17502,
    n17503, n17504, n17505, n17506, n17507, n17509,
    n17510, n17511, n17512, n17513, n17514, n17515,
    n17516, n17517, n17518, n17519, n17520, n17521,
    n17522, n17523, n17524, n17525, n17526, n17527,
    n17528, n17529, n17530, n17531, n17532, n17533,
    n17534, n17535, n17536, n17537, n17538, n17539,
    n17540, n17541, n17542, n17543, n17544, n17545,
    n17546, n17547, n17548, n17549, n17550, n17551,
    n17552, n17553, n17554, n17555, n17556, n17557,
    n17558, n17559, n17560, n17561, n17562, n17563,
    n17564, n17565, n17566, n17567, n17568, n17569,
    n17570, n17571, n17572, n17573, n17574, n17575,
    n17576, n17577, n17578, n17579, n17580, n17581,
    n17582, n17583, n17584, n17585, n17586, n17587,
    n17588, n17589, n17590, n17591, n17592, n17593,
    n17594, n17595, n17596, n17597, n17598, n17599,
    n17600, n17601, n17602, n17603, n17604, n17605,
    n17606, n17607, n17608, n17609, n17610, n17611,
    n17612, n17613, n17614, n17615, n17616, n17617,
    n17618, n17619, n17620, n17621, n17622, n17623,
    n17624, n17625, n17626, n17627, n17628, n17629,
    n17630, n17631, n17632, n17633, n17634, n17635,
    n17636, n17637, n17638, n17639, n17640, n17641,
    n17642, n17643, n17644, n17645, n17646, n17647,
    n17648, n17649, n17650, n17651, n17652, n17653,
    n17654, n17655, n17656, n17657, n17658, n17659,
    n17660, n17661, n17662, n17663, n17664, n17665,
    n17666, n17667, n17668, n17669, n17670, n17671,
    n17672, n17673, n17674, n17675, n17676, n17677,
    n17678, n17679, n17680, n17681, n17682, n17683,
    n17684, n17685, n17686, n17687, n17688, n17689,
    n17690, n17691, n17692, n17693, n17694, n17695,
    n17696, n17697, n17698, n17699, n17700, n17701,
    n17702, n17703, n17704, n17705, n17706, n17707,
    n17708, n17709, n17710, n17711, n17712, n17713,
    n17714, n17715, n17716, n17717, n17718, n17719,
    n17720, n17721, n17722, n17723, n17724, n17725,
    n17726, n17727, n17728, n17729, n17730, n17731,
    n17732, n17733, n17734, n17735, n17736, n17737,
    n17738, n17739, n17740, n17741, n17742, n17743,
    n17744, n17745, n17746, n17747, n17748, n17749,
    n17750, n17751, n17752, n17753, n17754, n17755,
    n17756, n17757, n17758, n17759, n17760, n17761,
    n17762, n17763, n17764, n17765, n17766, n17767,
    n17768, n17769, n17770, n17771, n17772, n17773,
    n17774, n17775, n17776, n17777, n17778, n17779,
    n17780, n17781, n17782, n17783, n17784, n17785,
    n17786, n17787, n17788, n17789, n17790, n17792,
    n17793, n17794, n17795, n17796, n17797, n17798,
    n17799, n17800, n17801, n17802, n17803, n17804,
    n17805, n17806, n17807, n17808, n17809, n17810,
    n17811, n17812, n17813, n17814, n17815, n17816,
    n17817, n17818, n17819, n17820, n17821, n17822,
    n17823, n17824, n17825, n17826, n17827, n17828,
    n17829, n17830, n17831, n17832, n17833, n17834,
    n17835, n17836, n17837, n17838, n17839, n17840,
    n17841, n17842, n17843, n17844, n17845, n17846,
    n17847, n17848, n17849, n17850, n17851, n17852,
    n17853, n17854, n17855, n17856, n17857, n17858,
    n17859, n17860, n17861, n17862, n17863, n17864,
    n17865, n17866, n17867, n17868, n17869, n17870,
    n17871, n17872, n17873, n17874, n17875, n17876,
    n17877, n17878, n17879, n17880, n17881, n17882,
    n17883, n17884, n17885, n17886, n17887, n17888,
    n17889, n17890, n17891, n17892, n17893, n17894,
    n17895, n17896, n17897, n17898, n17899, n17900,
    n17901, n17902, n17903, n17904, n17905, n17906,
    n17907, n17908, n17909, n17910, n17911, n17912,
    n17913, n17914, n17915, n17916, n17917, n17918,
    n17919, n17920, n17921, n17922, n17923, n17924,
    n17925, n17926, n17927, n17928, n17929, n17930,
    n17931, n17932, n17933, n17934, n17935, n17936,
    n17937, n17938, n17939, n17940, n17941, n17942,
    n17943, n17944, n17945, n17946, n17947, n17948,
    n17949, n17950, n17951, n17952, n17953, n17954,
    n17955, n17956, n17957, n17958, n17959, n17960,
    n17961, n17962, n17963, n17964, n17965, n17966,
    n17967, n17968, n17969, n17970, n17971, n17972,
    n17973, n17974, n17975, n17976, n17977, n17978,
    n17979, n17980, n17981, n17982, n17983, n17984,
    n17985, n17986, n17987, n17988, n17989, n17990,
    n17991, n17992, n17993, n17994, n17995, n17996,
    n17997, n17998, n17999, n18000, n18001, n18002,
    n18003, n18004, n18005, n18006, n18007, n18008,
    n18009, n18010, n18011, n18012, n18013, n18014,
    n18015, n18016, n18017, n18018, n18019, n18020,
    n18021, n18022, n18023, n18024, n18025, n18026,
    n18027, n18028, n18029, n18030, n18031, n18032,
    n18033, n18034, n18035, n18036, n18037, n18038,
    n18039, n18040, n18041, n18042, n18043, n18044,
    n18045, n18046, n18047, n18048, n18049, n18050,
    n18051, n18052, n18053, n18054, n18055, n18056,
    n18057, n18058, n18059, n18060, n18061, n18062,
    n18063, n18064, n18065, n18066, n18067, n18068,
    n18069, n18070, n18071, n18072, n18073, n18074,
    n18076, n18077, n18078, n18079, n18080, n18081,
    n18082, n18083, n18084, n18085, n18086, n18087,
    n18088, n18089, n18090, n18091, n18092, n18093,
    n18094, n18095, n18096, n18097, n18098, n18099,
    n18100, n18101, n18102, n18103, n18104, n18105,
    n18106, n18107, n18108, n18109, n18110, n18111,
    n18112, n18113, n18114, n18115, n18116, n18117,
    n18118, n18119, n18120, n18121, n18122, n18123,
    n18124, n18125, n18126, n18127, n18128, n18129,
    n18130, n18131, n18132, n18133, n18134, n18135,
    n18136, n18137, n18138, n18139, n18140, n18141,
    n18142, n18143, n18144, n18145, n18146, n18147,
    n18148, n18149, n18150, n18151, n18152, n18153,
    n18154, n18155, n18156, n18157, n18158, n18159,
    n18160, n18161, n18162, n18163, n18164, n18165,
    n18166, n18167, n18168, n18169, n18170, n18171,
    n18172, n18173, n18174, n18175, n18176, n18177,
    n18178, n18179, n18180, n18181, n18182, n18183,
    n18184, n18185, n18186, n18187, n18188, n18189,
    n18190, n18191, n18192, n18193, n18194, n18195,
    n18196, n18197, n18198, n18199, n18200, n18201,
    n18202, n18203, n18204, n18205, n18206, n18207,
    n18208, n18209, n18210, n18211, n18212, n18213,
    n18214, n18215, n18216, n18217, n18218, n18219,
    n18220, n18221, n18222, n18223, n18224, n18225,
    n18226, n18227, n18228, n18229, n18230, n18231,
    n18232, n18233, n18234, n18235, n18236, n18237,
    n18238, n18239, n18240, n18241, n18242, n18243,
    n18244, n18245, n18246, n18247, n18248, n18249,
    n18250, n18251, n18252, n18253, n18254, n18255,
    n18256, n18257, n18258, n18259, n18260, n18261,
    n18262, n18263, n18264, n18265, n18266, n18267,
    n18268, n18269, n18270, n18271, n18272, n18273,
    n18274, n18275, n18276, n18277, n18278, n18279,
    n18280, n18281, n18282, n18283, n18284, n18285,
    n18286, n18287, n18288, n18289, n18290, n18291,
    n18292, n18293, n18294, n18295, n18296, n18297,
    n18298, n18299, n18300, n18301, n18302, n18303,
    n18304, n18305, n18306, n18307, n18308, n18309,
    n18310, n18311, n18312, n18313, n18314, n18315,
    n18316, n18317, n18318, n18319, n18320, n18321,
    n18322, n18323, n18324, n18325, n18326, n18327,
    n18328, n18329, n18330, n18331, n18332, n18333,
    n18334, n18335, n18336, n18337, n18338, n18339,
    n18340, n18341, n18342, n18343, n18344, n18345,
    n18346, n18347, n18348, n18349, n18351, n18352,
    n18353, n18354, n18355, n18356, n18357, n18358,
    n18359, n18360, n18361, n18362, n18363, n18364,
    n18365, n18366, n18367, n18368, n18369, n18370,
    n18371, n18372, n18373, n18374, n18375, n18376,
    n18377, n18378, n18379, n18380, n18381, n18382,
    n18383, n18384, n18385, n18386, n18387, n18388,
    n18389, n18390, n18391, n18392, n18393, n18394,
    n18395, n18396, n18397, n18398, n18399, n18400,
    n18401, n18402, n18403, n18404, n18405, n18406,
    n18407, n18408, n18409, n18410, n18411, n18412,
    n18413, n18414, n18415, n18416, n18417, n18418,
    n18419, n18420, n18421, n18422, n18423, n18424,
    n18425, n18426, n18427, n18428, n18429, n18430,
    n18431, n18432, n18433, n18434, n18435, n18436,
    n18437, n18438, n18439, n18440, n18441, n18442,
    n18443, n18444, n18445, n18446, n18447, n18448,
    n18449, n18450, n18451, n18452, n18453, n18454,
    n18455, n18456, n18457, n18458, n18459, n18460,
    n18461, n18462, n18463, n18464, n18465, n18466,
    n18467, n18468, n18469, n18470, n18471, n18472,
    n18473, n18474, n18475, n18476, n18477, n18478,
    n18479, n18480, n18481, n18482, n18483, n18484,
    n18485, n18486, n18487, n18488, n18489, n18490,
    n18491, n18492, n18493, n18494, n18495, n18496,
    n18497, n18498, n18499, n18500, n18501, n18502,
    n18503, n18504, n18505, n18506, n18507, n18508,
    n18509, n18510, n18511, n18512, n18513, n18514,
    n18515, n18516, n18517, n18518, n18519, n18520,
    n18521, n18522, n18523, n18524, n18525, n18526,
    n18527, n18528, n18529, n18530, n18531, n18532,
    n18533, n18534, n18535, n18536, n18537, n18538,
    n18539, n18540, n18541, n18542, n18543, n18544,
    n18545, n18546, n18547, n18548, n18549, n18550,
    n18551, n18552, n18553, n18554, n18555, n18556,
    n18557, n18558, n18559, n18560, n18561, n18562,
    n18563, n18564, n18565, n18566, n18567, n18568,
    n18569, n18570, n18571, n18572, n18573, n18574,
    n18575, n18576, n18577, n18578, n18579, n18580,
    n18581, n18582, n18583, n18584, n18585, n18586,
    n18587, n18588, n18589, n18590, n18591, n18592,
    n18593, n18594, n18595, n18596, n18597, n18598,
    n18599, n18600, n18601, n18602, n18603, n18604,
    n18605, n18606, n18607, n18608, n18609, n18610,
    n18611, n18612, n18613, n18614, n18615, n18616,
    n18617, n18619, n18620, n18621, n18622, n18623,
    n18624, n18625, n18626, n18627, n18628, n18629,
    n18630, n18631, n18632, n18633, n18634, n18635,
    n18636, n18637, n18638, n18639, n18640, n18641,
    n18642, n18643, n18644, n18645, n18646, n18647,
    n18648, n18649, n18650, n18651, n18652, n18653,
    n18654, n18655, n18656, n18657, n18658, n18659,
    n18660, n18661, n18662, n18663, n18664, n18665,
    n18666, n18667, n18668, n18669, n18670, n18671,
    n18672, n18673, n18674, n18675, n18676, n18677,
    n18678, n18679, n18680, n18681, n18682, n18683,
    n18684, n18685, n18686, n18687, n18688, n18689,
    n18690, n18691, n18692, n18693, n18694, n18695,
    n18696, n18697, n18698, n18699, n18700, n18701,
    n18702, n18703, n18704, n18705, n18706, n18707,
    n18708, n18709, n18710, n18711, n18712, n18713,
    n18714, n18715, n18716, n18717, n18718, n18719,
    n18720, n18721, n18722, n18723, n18724, n18725,
    n18726, n18727, n18728, n18729, n18730, n18731,
    n18732, n18733, n18734, n18735, n18736, n18737,
    n18738, n18739, n18740, n18741, n18742, n18743,
    n18744, n18745, n18746, n18747, n18748, n18749,
    n18750, n18751, n18752, n18753, n18754, n18755,
    n18756, n18757, n18758, n18759, n18760, n18761,
    n18762, n18763, n18764, n18765, n18766, n18767,
    n18768, n18769, n18770, n18771, n18772, n18773,
    n18774, n18775, n18776, n18777, n18778, n18779,
    n18780, n18781, n18782, n18783, n18784, n18785,
    n18786, n18787, n18788, n18789, n18790, n18791,
    n18792, n18793, n18794, n18795, n18796, n18797,
    n18798, n18799, n18800, n18801, n18802, n18803,
    n18804, n18805, n18806, n18807, n18808, n18809,
    n18810, n18811, n18812, n18813, n18814, n18815,
    n18816, n18817, n18818, n18819, n18820, n18821,
    n18822, n18823, n18824, n18825, n18826, n18827,
    n18828, n18829, n18830, n18831, n18832, n18833,
    n18834, n18835, n18836, n18837, n18838, n18839,
    n18840, n18841, n18842, n18843, n18844, n18845,
    n18846, n18847, n18848, n18849, n18850, n18851,
    n18852, n18853, n18854, n18855, n18856, n18857,
    n18858, n18859, n18860, n18861, n18862, n18863,
    n18864, n18865, n18866, n18867, n18868, n18869,
    n18870, n18871, n18872, n18873, n18874, n18875,
    n18876, n18877, n18878, n18879, n18880, n18881,
    n18882, n18883, n18884, n18885, n18887, n18888,
    n18889, n18890, n18891, n18892, n18893, n18894,
    n18895, n18896, n18897, n18898, n18899, n18900,
    n18901, n18902, n18903, n18904, n18905, n18906,
    n18907, n18908, n18909, n18910, n18911, n18912,
    n18913, n18914, n18915, n18916, n18917, n18918,
    n18919, n18920, n18921, n18922, n18923, n18924,
    n18925, n18926, n18927, n18928, n18929, n18930,
    n18931, n18932, n18933, n18934, n18935, n18936,
    n18937, n18938, n18939, n18940, n18941, n18942,
    n18943, n18944, n18945, n18946, n18947, n18948,
    n18949, n18950, n18951, n18952, n18953, n18954,
    n18955, n18956, n18957, n18958, n18959, n18960,
    n18961, n18962, n18963, n18964, n18965, n18966,
    n18967, n18968, n18969, n18970, n18971, n18972,
    n18973, n18974, n18975, n18976, n18977, n18978,
    n18979, n18980, n18981, n18982, n18983, n18984,
    n18985, n18986, n18987, n18988, n18989, n18990,
    n18991, n18992, n18993, n18994, n18995, n18996,
    n18997, n18998, n18999, n19000, n19001, n19002,
    n19003, n19004, n19005, n19006, n19007, n19008,
    n19009, n19010, n19011, n19012, n19013, n19014,
    n19015, n19016, n19017, n19018, n19019, n19020,
    n19021, n19022, n19023, n19024, n19025, n19026,
    n19027, n19028, n19029, n19030, n19031, n19032,
    n19033, n19034, n19035, n19036, n19037, n19038,
    n19039, n19040, n19041, n19042, n19043, n19044,
    n19045, n19046, n19047, n19048, n19049, n19050,
    n19051, n19052, n19053, n19054, n19055, n19056,
    n19057, n19058, n19059, n19060, n19061, n19062,
    n19063, n19064, n19065, n19066, n19067, n19068,
    n19069, n19070, n19071, n19072, n19073, n19074,
    n19075, n19076, n19077, n19078, n19079, n19080,
    n19081, n19082, n19083, n19084, n19085, n19086,
    n19087, n19088, n19089, n19090, n19091, n19092,
    n19093, n19094, n19095, n19096, n19097, n19098,
    n19099, n19100, n19101, n19102, n19103, n19104,
    n19105, n19106, n19107, n19108, n19109, n19110,
    n19111, n19112, n19113, n19114, n19115, n19116,
    n19117, n19118, n19119, n19120, n19121, n19122,
    n19123, n19124, n19125, n19126, n19127, n19128,
    n19129, n19130, n19131, n19132, n19133, n19134,
    n19135, n19136, n19137, n19138, n19139, n19140,
    n19141, n19142, n19144, n19145, n19146, n19147,
    n19148, n19149, n19150, n19151, n19152, n19153,
    n19154, n19155, n19156, n19157, n19158, n19159,
    n19160, n19161, n19162, n19163, n19164, n19165,
    n19166, n19167, n19168, n19169, n19170, n19171,
    n19172, n19173, n19174, n19175, n19176, n19177,
    n19178, n19179, n19180, n19181, n19182, n19183,
    n19184, n19185, n19186, n19187, n19188, n19189,
    n19190, n19191, n19192, n19193, n19194, n19195,
    n19196, n19197, n19198, n19199, n19200, n19201,
    n19202, n19203, n19204, n19205, n19206, n19207,
    n19208, n19209, n19210, n19211, n19212, n19213,
    n19214, n19215, n19216, n19217, n19218, n19219,
    n19220, n19221, n19222, n19223, n19224, n19225,
    n19226, n19227, n19228, n19229, n19230, n19231,
    n19232, n19233, n19234, n19235, n19236, n19237,
    n19238, n19239, n19240, n19241, n19242, n19243,
    n19244, n19245, n19246, n19247, n19248, n19249,
    n19250, n19251, n19252, n19253, n19254, n19255,
    n19256, n19257, n19258, n19259, n19260, n19261,
    n19262, n19263, n19264, n19265, n19266, n19267,
    n19268, n19269, n19270, n19271, n19272, n19273,
    n19274, n19275, n19276, n19277, n19278, n19279,
    n19280, n19281, n19282, n19283, n19284, n19285,
    n19286, n19287, n19288, n19289, n19290, n19291,
    n19292, n19293, n19294, n19295, n19296, n19297,
    n19298, n19299, n19300, n19301, n19302, n19303,
    n19304, n19305, n19306, n19307, n19308, n19309,
    n19310, n19311, n19312, n19313, n19314, n19315,
    n19316, n19317, n19318, n19319, n19320, n19321,
    n19322, n19323, n19324, n19325, n19326, n19327,
    n19328, n19329, n19330, n19331, n19332, n19333,
    n19334, n19335, n19336, n19337, n19338, n19339,
    n19340, n19341, n19342, n19343, n19344, n19345,
    n19346, n19347, n19348, n19349, n19350, n19351,
    n19352, n19353, n19354, n19355, n19356, n19357,
    n19358, n19359, n19360, n19361, n19362, n19363,
    n19364, n19365, n19366, n19367, n19368, n19369,
    n19370, n19371, n19372, n19373, n19374, n19375,
    n19376, n19377, n19378, n19379, n19380, n19381,
    n19382, n19383, n19384, n19385, n19386, n19387,
    n19388, n19389, n19390, n19392, n19393, n19394,
    n19395, n19396, n19397, n19398, n19399, n19400,
    n19401, n19402, n19403, n19404, n19405, n19406,
    n19407, n19408, n19409, n19410, n19411, n19412,
    n19413, n19414, n19415, n19416, n19417, n19418,
    n19419, n19420, n19421, n19422, n19423, n19424,
    n19425, n19426, n19427, n19428, n19429, n19430,
    n19431, n19432, n19433, n19434, n19435, n19436,
    n19437, n19438, n19439, n19440, n19441, n19442,
    n19443, n19444, n19445, n19446, n19447, n19448,
    n19449, n19450, n19451, n19452, n19453, n19454,
    n19455, n19456, n19457, n19458, n19459, n19460,
    n19461, n19462, n19463, n19464, n19465, n19466,
    n19467, n19468, n19469, n19470, n19471, n19472,
    n19473, n19474, n19475, n19476, n19477, n19478,
    n19479, n19480, n19481, n19482, n19483, n19484,
    n19485, n19486, n19487, n19488, n19489, n19490,
    n19491, n19492, n19493, n19494, n19495, n19496,
    n19497, n19498, n19499, n19500, n19501, n19502,
    n19503, n19504, n19505, n19506, n19507, n19508,
    n19509, n19510, n19511, n19512, n19513, n19514,
    n19515, n19516, n19517, n19518, n19519, n19520,
    n19521, n19522, n19523, n19524, n19525, n19526,
    n19527, n19528, n19529, n19530, n19531, n19532,
    n19533, n19534, n19535, n19536, n19537, n19538,
    n19539, n19540, n19541, n19542, n19543, n19544,
    n19545, n19546, n19547, n19548, n19549, n19550,
    n19551, n19552, n19553, n19554, n19555, n19556,
    n19557, n19558, n19559, n19560, n19561, n19562,
    n19563, n19564, n19565, n19566, n19567, n19568,
    n19569, n19570, n19571, n19572, n19573, n19574,
    n19575, n19576, n19577, n19578, n19579, n19580,
    n19581, n19582, n19583, n19584, n19585, n19586,
    n19587, n19588, n19589, n19590, n19591, n19592,
    n19593, n19594, n19595, n19596, n19597, n19598,
    n19599, n19600, n19601, n19602, n19603, n19604,
    n19605, n19606, n19607, n19608, n19609, n19610,
    n19611, n19612, n19613, n19614, n19615, n19616,
    n19617, n19618, n19619, n19620, n19621, n19622,
    n19623, n19624, n19625, n19626, n19627, n19628,
    n19629, n19630, n19631, n19632, n19633, n19634,
    n19635, n19636, n19637, n19638, n19639, n19640,
    n19641, n19643, n19644, n19645, n19646, n19647,
    n19648, n19649, n19650, n19651, n19652, n19653,
    n19654, n19655, n19656, n19657, n19658, n19659,
    n19660, n19661, n19662, n19663, n19664, n19665,
    n19666, n19667, n19668, n19669, n19670, n19671,
    n19672, n19673, n19674, n19675, n19676, n19677,
    n19678, n19679, n19680, n19681, n19682, n19683,
    n19684, n19685, n19686, n19687, n19688, n19689,
    n19690, n19691, n19692, n19693, n19694, n19695,
    n19696, n19697, n19698, n19699, n19700, n19701,
    n19702, n19703, n19704, n19705, n19706, n19707,
    n19708, n19709, n19710, n19711, n19712, n19713,
    n19714, n19715, n19716, n19717, n19718, n19719,
    n19720, n19721, n19722, n19723, n19724, n19725,
    n19726, n19727, n19728, n19729, n19730, n19731,
    n19732, n19733, n19734, n19735, n19736, n19737,
    n19738, n19739, n19740, n19741, n19742, n19743,
    n19744, n19745, n19746, n19747, n19748, n19749,
    n19750, n19751, n19752, n19753, n19754, n19755,
    n19756, n19757, n19758, n19759, n19760, n19761,
    n19762, n19763, n19764, n19765, n19766, n19767,
    n19768, n19769, n19770, n19771, n19772, n19773,
    n19774, n19775, n19776, n19777, n19778, n19779,
    n19780, n19781, n19782, n19783, n19784, n19785,
    n19786, n19787, n19788, n19789, n19790, n19791,
    n19792, n19793, n19794, n19795, n19796, n19797,
    n19798, n19799, n19800, n19801, n19802, n19803,
    n19804, n19805, n19806, n19807, n19808, n19809,
    n19810, n19811, n19812, n19813, n19814, n19815,
    n19816, n19817, n19818, n19819, n19820, n19821,
    n19822, n19823, n19824, n19825, n19826, n19827,
    n19828, n19829, n19830, n19831, n19832, n19833,
    n19834, n19835, n19836, n19837, n19838, n19839,
    n19840, n19841, n19842, n19843, n19844, n19845,
    n19846, n19847, n19848, n19849, n19850, n19851,
    n19852, n19853, n19854, n19855, n19856, n19857,
    n19858, n19859, n19860, n19861, n19862, n19863,
    n19864, n19865, n19866, n19867, n19868, n19869,
    n19870, n19871, n19872, n19873, n19874, n19875,
    n19876, n19877, n19878, n19879, n19880, n19881,
    n19882, n19883, n19884, n19886, n19887, n19888,
    n19889, n19890, n19891, n19892, n19893, n19894,
    n19895, n19896, n19897, n19898, n19899, n19900,
    n19901, n19902, n19903, n19904, n19905, n19906,
    n19907, n19908, n19909, n19910, n19911, n19912,
    n19913, n19914, n19915, n19916, n19917, n19918,
    n19919, n19920, n19921, n19922, n19923, n19924,
    n19925, n19926, n19927, n19928, n19929, n19930,
    n19931, n19932, n19933, n19934, n19935, n19936,
    n19937, n19938, n19939, n19940, n19941, n19942,
    n19943, n19944, n19945, n19946, n19947, n19948,
    n19949, n19950, n19951, n19952, n19953, n19954,
    n19955, n19956, n19957, n19958, n19959, n19960,
    n19961, n19962, n19963, n19964, n19965, n19966,
    n19967, n19968, n19969, n19970, n19971, n19972,
    n19973, n19974, n19975, n19976, n19977, n19978,
    n19979, n19980, n19981, n19982, n19983, n19984,
    n19985, n19986, n19987, n19988, n19989, n19990,
    n19991, n19992, n19993, n19994, n19995, n19996,
    n19997, n19998, n19999, n20000, n20001, n20002,
    n20003, n20004, n20005, n20006, n20007, n20008,
    n20009, n20010, n20011, n20012, n20013, n20014,
    n20015, n20016, n20017, n20018, n20019, n20020,
    n20021, n20022, n20023, n20024, n20025, n20026,
    n20027, n20028, n20029, n20030, n20031, n20032,
    n20033, n20034, n20035, n20036, n20037, n20038,
    n20039, n20040, n20041, n20042, n20043, n20044,
    n20045, n20046, n20047, n20048, n20049, n20050,
    n20051, n20052, n20053, n20054, n20055, n20056,
    n20057, n20058, n20059, n20060, n20061, n20062,
    n20063, n20064, n20065, n20066, n20067, n20068,
    n20069, n20070, n20071, n20072, n20073, n20074,
    n20075, n20076, n20077, n20078, n20079, n20080,
    n20081, n20082, n20083, n20084, n20085, n20086,
    n20087, n20088, n20089, n20090, n20091, n20092,
    n20093, n20094, n20095, n20096, n20097, n20098,
    n20099, n20100, n20101, n20102, n20103, n20104,
    n20105, n20106, n20107, n20108, n20109, n20110,
    n20111, n20112, n20113, n20114, n20115, n20117,
    n20118, n20119, n20120, n20121, n20122, n20123,
    n20124, n20125, n20126, n20127, n20128, n20129,
    n20130, n20131, n20132, n20133, n20134, n20135,
    n20136, n20137, n20138, n20139, n20140, n20141,
    n20142, n20143, n20144, n20145, n20146, n20147,
    n20148, n20149, n20150, n20151, n20152, n20153,
    n20154, n20155, n20156, n20157, n20158, n20159,
    n20160, n20161, n20162, n20163, n20164, n20165,
    n20166, n20167, n20168, n20169, n20170, n20171,
    n20172, n20173, n20174, n20175, n20176, n20177,
    n20178, n20179, n20180, n20181, n20182, n20183,
    n20184, n20185, n20186, n20187, n20188, n20189,
    n20190, n20191, n20192, n20193, n20194, n20195,
    n20196, n20197, n20198, n20199, n20200, n20201,
    n20202, n20203, n20204, n20205, n20206, n20207,
    n20208, n20209, n20210, n20211, n20212, n20213,
    n20214, n20215, n20216, n20217, n20218, n20219,
    n20220, n20221, n20222, n20223, n20224, n20225,
    n20226, n20227, n20228, n20229, n20230, n20231,
    n20232, n20233, n20234, n20235, n20236, n20237,
    n20238, n20239, n20240, n20241, n20242, n20243,
    n20244, n20245, n20246, n20247, n20248, n20249,
    n20250, n20251, n20252, n20253, n20254, n20255,
    n20256, n20257, n20258, n20259, n20260, n20261,
    n20262, n20263, n20264, n20265, n20266, n20267,
    n20268, n20269, n20270, n20271, n20272, n20273,
    n20274, n20275, n20276, n20277, n20278, n20279,
    n20280, n20281, n20282, n20283, n20284, n20285,
    n20286, n20287, n20288, n20289, n20290, n20291,
    n20292, n20293, n20294, n20295, n20296, n20297,
    n20298, n20299, n20300, n20301, n20302, n20303,
    n20304, n20305, n20306, n20307, n20308, n20309,
    n20310, n20311, n20312, n20313, n20314, n20315,
    n20316, n20317, n20318, n20319, n20320, n20321,
    n20322, n20323, n20324, n20325, n20326, n20327,
    n20328, n20329, n20330, n20331, n20332, n20333,
    n20334, n20335, n20336, n20337, n20338, n20339,
    n20340, n20341, n20342, n20343, n20344, n20345,
    n20346, n20347, n20348, n20350, n20351, n20352,
    n20353, n20354, n20355, n20356, n20357, n20358,
    n20359, n20360, n20361, n20362, n20363, n20364,
    n20365, n20366, n20367, n20368, n20369, n20370,
    n20371, n20372, n20373, n20374, n20375, n20376,
    n20377, n20378, n20379, n20380, n20381, n20382,
    n20383, n20384, n20385, n20386, n20387, n20388,
    n20389, n20390, n20391, n20392, n20393, n20394,
    n20395, n20396, n20397, n20398, n20399, n20400,
    n20401, n20402, n20403, n20404, n20405, n20406,
    n20407, n20408, n20409, n20410, n20411, n20412,
    n20413, n20414, n20415, n20416, n20417, n20418,
    n20419, n20420, n20421, n20422, n20423, n20424,
    n20425, n20426, n20427, n20428, n20429, n20430,
    n20431, n20432, n20433, n20434, n20435, n20436,
    n20437, n20438, n20439, n20440, n20441, n20442,
    n20443, n20444, n20445, n20446, n20447, n20448,
    n20449, n20450, n20451, n20452, n20453, n20454,
    n20455, n20456, n20457, n20458, n20459, n20460,
    n20461, n20462, n20463, n20464, n20465, n20466,
    n20467, n20468, n20469, n20470, n20471, n20472,
    n20473, n20474, n20475, n20476, n20477, n20478,
    n20479, n20480, n20481, n20482, n20483, n20484,
    n20485, n20486, n20487, n20488, n20489, n20490,
    n20491, n20492, n20493, n20494, n20495, n20496,
    n20497, n20498, n20499, n20500, n20501, n20502,
    n20503, n20504, n20505, n20506, n20507, n20508,
    n20509, n20510, n20511, n20512, n20513, n20514,
    n20515, n20516, n20517, n20518, n20519, n20520,
    n20521, n20522, n20523, n20524, n20525, n20526,
    n20527, n20528, n20529, n20530, n20531, n20532,
    n20533, n20534, n20535, n20536, n20537, n20538,
    n20539, n20540, n20541, n20542, n20543, n20544,
    n20545, n20546, n20547, n20548, n20549, n20550,
    n20551, n20552, n20553, n20554, n20555, n20556,
    n20557, n20558, n20559, n20560, n20561, n20562,
    n20563, n20564, n20565, n20566, n20567, n20568,
    n20569, n20570, n20571, n20572, n20573, n20575,
    n20576, n20577, n20578, n20579, n20580, n20581,
    n20582, n20583, n20584, n20585, n20586, n20587,
    n20588, n20589, n20590, n20591, n20592, n20593,
    n20594, n20595, n20596, n20597, n20598, n20599,
    n20600, n20601, n20602, n20603, n20604, n20605,
    n20606, n20607, n20608, n20609, n20610, n20611,
    n20612, n20613, n20614, n20615, n20616, n20617,
    n20618, n20619, n20620, n20621, n20622, n20623,
    n20624, n20625, n20626, n20627, n20628, n20629,
    n20630, n20631, n20632, n20633, n20634, n20635,
    n20636, n20637, n20638, n20639, n20640, n20641,
    n20642, n20643, n20644, n20645, n20646, n20647,
    n20648, n20649, n20650, n20651, n20652, n20653,
    n20654, n20655, n20656, n20657, n20658, n20659,
    n20660, n20661, n20662, n20663, n20664, n20665,
    n20666, n20667, n20668, n20669, n20670, n20671,
    n20672, n20673, n20674, n20675, n20676, n20677,
    n20678, n20679, n20680, n20681, n20682, n20683,
    n20684, n20685, n20686, n20687, n20688, n20689,
    n20690, n20691, n20692, n20693, n20694, n20695,
    n20696, n20697, n20698, n20699, n20700, n20701,
    n20702, n20703, n20704, n20705, n20706, n20707,
    n20708, n20709, n20710, n20711, n20712, n20713,
    n20714, n20715, n20716, n20717, n20718, n20719,
    n20720, n20721, n20722, n20723, n20724, n20725,
    n20726, n20727, n20728, n20729, n20730, n20731,
    n20732, n20733, n20734, n20735, n20736, n20737,
    n20738, n20739, n20740, n20741, n20742, n20743,
    n20744, n20745, n20746, n20747, n20748, n20749,
    n20750, n20751, n20752, n20753, n20754, n20755,
    n20756, n20757, n20758, n20759, n20760, n20761,
    n20762, n20763, n20764, n20765, n20766, n20767,
    n20768, n20769, n20770, n20771, n20772, n20773,
    n20774, n20775, n20776, n20777, n20778, n20779,
    n20780, n20781, n20782, n20783, n20784, n20785,
    n20786, n20787, n20788, n20790, n20791, n20792,
    n20793, n20794, n20795, n20796, n20797, n20798,
    n20799, n20800, n20801, n20802, n20803, n20804,
    n20805, n20806, n20807, n20808, n20809, n20810,
    n20811, n20812, n20813, n20814, n20815, n20816,
    n20817, n20818, n20819, n20820, n20821, n20822,
    n20823, n20824, n20825, n20826, n20827, n20828,
    n20829, n20830, n20831, n20832, n20833, n20834,
    n20835, n20836, n20837, n20838, n20839, n20840,
    n20841, n20842, n20843, n20844, n20845, n20846,
    n20847, n20848, n20849, n20850, n20851, n20852,
    n20853, n20854, n20855, n20856, n20857, n20858,
    n20859, n20860, n20861, n20862, n20863, n20864,
    n20865, n20866, n20867, n20868, n20869, n20870,
    n20871, n20872, n20873, n20874, n20875, n20876,
    n20877, n20878, n20879, n20880, n20881, n20882,
    n20883, n20884, n20885, n20886, n20887, n20888,
    n20889, n20890, n20891, n20892, n20893, n20894,
    n20895, n20896, n20897, n20898, n20899, n20900,
    n20901, n20902, n20903, n20904, n20905, n20906,
    n20907, n20908, n20909, n20910, n20911, n20912,
    n20913, n20914, n20915, n20916, n20917, n20918,
    n20919, n20920, n20921, n20922, n20923, n20924,
    n20925, n20926, n20927, n20928, n20929, n20930,
    n20931, n20932, n20933, n20934, n20935, n20936,
    n20937, n20938, n20939, n20940, n20941, n20942,
    n20943, n20944, n20945, n20946, n20947, n20948,
    n20949, n20950, n20951, n20952, n20953, n20954,
    n20955, n20956, n20957, n20958, n20959, n20960,
    n20961, n20962, n20963, n20964, n20965, n20966,
    n20967, n20968, n20969, n20970, n20971, n20972,
    n20973, n20974, n20975, n20976, n20977, n20978,
    n20979, n20980, n20981, n20982, n20983, n20984,
    n20985, n20986, n20987, n20988, n20989, n20990,
    n20991, n20992, n20993, n20994, n20995, n20996,
    n20997, n20998, n20999, n21000, n21001, n21002,
    n21003, n21004, n21006, n21007, n21008, n21009,
    n21010, n21011, n21012, n21013, n21014, n21015,
    n21016, n21017, n21018, n21019, n21020, n21021,
    n21022, n21023, n21024, n21025, n21026, n21027,
    n21028, n21029, n21030, n21031, n21032, n21033,
    n21034, n21035, n21036, n21037, n21038, n21039,
    n21040, n21041, n21042, n21043, n21044, n21045,
    n21046, n21047, n21048, n21049, n21050, n21051,
    n21052, n21053, n21054, n21055, n21056, n21057,
    n21058, n21059, n21060, n21061, n21062, n21063,
    n21064, n21065, n21066, n21067, n21068, n21069,
    n21070, n21071, n21072, n21073, n21074, n21075,
    n21076, n21077, n21078, n21079, n21080, n21081,
    n21082, n21083, n21084, n21085, n21086, n21087,
    n21088, n21089, n21090, n21091, n21092, n21093,
    n21094, n21095, n21096, n21097, n21098, n21099,
    n21100, n21101, n21102, n21103, n21104, n21105,
    n21106, n21107, n21108, n21109, n21110, n21111,
    n21112, n21113, n21114, n21115, n21116, n21117,
    n21118, n21119, n21120, n21121, n21122, n21123,
    n21124, n21125, n21126, n21127, n21128, n21129,
    n21130, n21131, n21132, n21133, n21134, n21135,
    n21136, n21137, n21138, n21139, n21140, n21141,
    n21142, n21143, n21144, n21145, n21146, n21147,
    n21148, n21149, n21150, n21151, n21152, n21153,
    n21154, n21155, n21156, n21157, n21158, n21159,
    n21160, n21161, n21162, n21163, n21164, n21165,
    n21166, n21167, n21168, n21169, n21170, n21171,
    n21172, n21173, n21174, n21175, n21176, n21177,
    n21178, n21179, n21180, n21181, n21182, n21183,
    n21184, n21185, n21186, n21187, n21188, n21189,
    n21190, n21191, n21192, n21193, n21194, n21195,
    n21196, n21197, n21198, n21199, n21200, n21201,
    n21202, n21203, n21204, n21205, n21206, n21207,
    n21208, n21209, n21210, n21211, n21213, n21214,
    n21215, n21216, n21217, n21218, n21219, n21220,
    n21221, n21222, n21223, n21224, n21225, n21226,
    n21227, n21228, n21229, n21230, n21231, n21232,
    n21233, n21234, n21235, n21236, n21237, n21238,
    n21239, n21240, n21241, n21242, n21243, n21244,
    n21245, n21246, n21247, n21248, n21249, n21250,
    n21251, n21252, n21253, n21254, n21255, n21256,
    n21257, n21258, n21259, n21260, n21261, n21262,
    n21263, n21264, n21265, n21266, n21267, n21268,
    n21269, n21270, n21271, n21272, n21273, n21274,
    n21275, n21276, n21277, n21278, n21279, n21280,
    n21281, n21282, n21283, n21284, n21285, n21286,
    n21287, n21288, n21289, n21290, n21291, n21292,
    n21293, n21294, n21295, n21296, n21297, n21298,
    n21299, n21300, n21301, n21302, n21303, n21304,
    n21305, n21306, n21307, n21308, n21309, n21310,
    n21311, n21312, n21313, n21314, n21315, n21316,
    n21317, n21318, n21319, n21320, n21321, n21322,
    n21323, n21324, n21325, n21326, n21327, n21328,
    n21329, n21330, n21331, n21332, n21333, n21334,
    n21335, n21336, n21337, n21338, n21339, n21340,
    n21341, n21342, n21343, n21344, n21345, n21346,
    n21347, n21348, n21349, n21350, n21351, n21352,
    n21353, n21354, n21355, n21356, n21357, n21358,
    n21359, n21360, n21361, n21362, n21363, n21364,
    n21365, n21366, n21367, n21368, n21369, n21370,
    n21371, n21372, n21373, n21374, n21375, n21376,
    n21377, n21378, n21379, n21380, n21381, n21382,
    n21383, n21384, n21385, n21386, n21387, n21388,
    n21389, n21390, n21391, n21392, n21393, n21394,
    n21395, n21396, n21397, n21398, n21399, n21400,
    n21401, n21402, n21403, n21404, n21405, n21406,
    n21407, n21408, n21409, n21411, n21412, n21413,
    n21414, n21415, n21416, n21417, n21418, n21419,
    n21420, n21421, n21422, n21423, n21424, n21425,
    n21426, n21427, n21428, n21429, n21430, n21431,
    n21432, n21433, n21434, n21435, n21436, n21437,
    n21438, n21439, n21440, n21441, n21442, n21443,
    n21444, n21445, n21446, n21447, n21448, n21449,
    n21450, n21451, n21452, n21453, n21454, n21455,
    n21456, n21457, n21458, n21459, n21460, n21461,
    n21462, n21463, n21464, n21465, n21466, n21467,
    n21468, n21469, n21470, n21471, n21472, n21473,
    n21474, n21475, n21476, n21477, n21478, n21479,
    n21480, n21481, n21482, n21483, n21484, n21485,
    n21486, n21487, n21488, n21489, n21490, n21491,
    n21492, n21493, n21494, n21495, n21496, n21497,
    n21498, n21499, n21500, n21501, n21502, n21503,
    n21504, n21505, n21506, n21507, n21508, n21509,
    n21510, n21511, n21512, n21513, n21514, n21515,
    n21516, n21517, n21518, n21519, n21520, n21521,
    n21522, n21523, n21524, n21525, n21526, n21527,
    n21528, n21529, n21530, n21531, n21532, n21533,
    n21534, n21535, n21536, n21537, n21538, n21539,
    n21540, n21541, n21542, n21543, n21544, n21545,
    n21546, n21547, n21548, n21549, n21550, n21551,
    n21552, n21553, n21554, n21555, n21556, n21557,
    n21558, n21559, n21560, n21561, n21562, n21563,
    n21564, n21565, n21566, n21567, n21568, n21569,
    n21570, n21571, n21572, n21573, n21574, n21575,
    n21576, n21577, n21578, n21579, n21580, n21581,
    n21582, n21583, n21584, n21585, n21586, n21587,
    n21588, n21589, n21590, n21591, n21592, n21593,
    n21594, n21595, n21596, n21597, n21598, n21599,
    n21600, n21601, n21602, n21603, n21604, n21605,
    n21606, n21607, n21609, n21610, n21611, n21612,
    n21613, n21614, n21615, n21616, n21617, n21618,
    n21619, n21620, n21621, n21622, n21623, n21624,
    n21625, n21626, n21627, n21628, n21629, n21630,
    n21631, n21632, n21633, n21634, n21635, n21636,
    n21637, n21638, n21639, n21640, n21641, n21642,
    n21643, n21644, n21645, n21646, n21647, n21648,
    n21649, n21650, n21651, n21652, n21653, n21654,
    n21655, n21656, n21657, n21658, n21659, n21660,
    n21661, n21662, n21663, n21664, n21665, n21666,
    n21667, n21668, n21669, n21670, n21671, n21672,
    n21673, n21674, n21675, n21676, n21677, n21678,
    n21679, n21680, n21681, n21682, n21683, n21684,
    n21685, n21686, n21687, n21688, n21689, n21690,
    n21691, n21692, n21693, n21694, n21695, n21696,
    n21697, n21698, n21699, n21700, n21701, n21702,
    n21703, n21704, n21705, n21706, n21707, n21708,
    n21709, n21710, n21711, n21712, n21713, n21714,
    n21715, n21716, n21717, n21718, n21719, n21720,
    n21721, n21722, n21723, n21724, n21725, n21726,
    n21727, n21728, n21729, n21730, n21731, n21732,
    n21733, n21734, n21735, n21736, n21737, n21738,
    n21739, n21740, n21741, n21742, n21743, n21744,
    n21745, n21746, n21747, n21748, n21749, n21750,
    n21751, n21752, n21753, n21754, n21755, n21756,
    n21757, n21758, n21759, n21760, n21761, n21762,
    n21763, n21764, n21765, n21766, n21767, n21768,
    n21769, n21770, n21771, n21772, n21773, n21774,
    n21775, n21776, n21777, n21778, n21779, n21780,
    n21781, n21782, n21783, n21784, n21785, n21786,
    n21787, n21788, n21789, n21790, n21791, n21792,
    n21793, n21794, n21795, n21796, n21797, n21799,
    n21800, n21801, n21802, n21803, n21804, n21805,
    n21806, n21807, n21808, n21809, n21810, n21811,
    n21812, n21813, n21814, n21815, n21816, n21817,
    n21818, n21819, n21820, n21821, n21822, n21823,
    n21824, n21825, n21826, n21827, n21828, n21829,
    n21830, n21831, n21832, n21833, n21834, n21835,
    n21836, n21837, n21838, n21839, n21840, n21841,
    n21842, n21843, n21844, n21845, n21846, n21847,
    n21848, n21849, n21850, n21851, n21852, n21853,
    n21854, n21855, n21856, n21857, n21858, n21859,
    n21860, n21861, n21862, n21863, n21864, n21865,
    n21866, n21867, n21868, n21869, n21870, n21871,
    n21872, n21873, n21874, n21875, n21876, n21877,
    n21878, n21879, n21880, n21881, n21882, n21883,
    n21884, n21885, n21886, n21887, n21888, n21889,
    n21890, n21891, n21892, n21893, n21894, n21895,
    n21896, n21897, n21898, n21899, n21900, n21901,
    n21902, n21903, n21904, n21905, n21906, n21907,
    n21908, n21909, n21910, n21911, n21912, n21913,
    n21914, n21915, n21916, n21917, n21918, n21919,
    n21920, n21921, n21922, n21923, n21924, n21925,
    n21926, n21927, n21928, n21929, n21930, n21931,
    n21932, n21933, n21934, n21935, n21936, n21937,
    n21938, n21939, n21940, n21941, n21942, n21943,
    n21944, n21945, n21946, n21947, n21948, n21949,
    n21950, n21951, n21952, n21953, n21954, n21955,
    n21956, n21957, n21958, n21959, n21960, n21961,
    n21962, n21963, n21964, n21965, n21966, n21967,
    n21968, n21969, n21970, n21971, n21972, n21973,
    n21974, n21975, n21976, n21977, n21978, n21980,
    n21981, n21982, n21983, n21984, n21985, n21986,
    n21987, n21988, n21989, n21990, n21991, n21992,
    n21993, n21994, n21995, n21996, n21997, n21998,
    n21999, n22000, n22001, n22002, n22003, n22004,
    n22005, n22006, n22007, n22008, n22009, n22010,
    n22011, n22012, n22013, n22014, n22015, n22016,
    n22017, n22018, n22019, n22020, n22021, n22022,
    n22023, n22024, n22025, n22026, n22027, n22028,
    n22029, n22030, n22031, n22032, n22033, n22034,
    n22035, n22036, n22037, n22038, n22039, n22040,
    n22041, n22042, n22043, n22044, n22045, n22046,
    n22047, n22048, n22049, n22050, n22051, n22052,
    n22053, n22054, n22055, n22056, n22057, n22058,
    n22059, n22060, n22061, n22062, n22063, n22064,
    n22065, n22066, n22067, n22068, n22069, n22070,
    n22071, n22072, n22073, n22074, n22075, n22076,
    n22077, n22078, n22079, n22080, n22081, n22082,
    n22083, n22084, n22085, n22086, n22087, n22088,
    n22089, n22090, n22091, n22092, n22093, n22094,
    n22095, n22096, n22097, n22098, n22099, n22100,
    n22101, n22102, n22103, n22104, n22105, n22106,
    n22107, n22108, n22109, n22110, n22111, n22112,
    n22113, n22114, n22115, n22116, n22117, n22118,
    n22119, n22120, n22121, n22122, n22123, n22124,
    n22125, n22126, n22127, n22128, n22129, n22130,
    n22131, n22132, n22133, n22134, n22135, n22136,
    n22137, n22138, n22139, n22140, n22141, n22142,
    n22143, n22144, n22145, n22146, n22147, n22148,
    n22149, n22150, n22151, n22152, n22153, n22154,
    n22155, n22156, n22157, n22158, n22159, n22161,
    n22162, n22163, n22164, n22165, n22166, n22167,
    n22168, n22169, n22170, n22171, n22172, n22173,
    n22174, n22175, n22176, n22177, n22178, n22179,
    n22180, n22181, n22182, n22183, n22184, n22185,
    n22186, n22187, n22188, n22189, n22190, n22191,
    n22192, n22193, n22194, n22195, n22196, n22197,
    n22198, n22199, n22200, n22201, n22202, n22203,
    n22204, n22205, n22206, n22207, n22208, n22209,
    n22210, n22211, n22212, n22213, n22214, n22215,
    n22216, n22217, n22218, n22219, n22220, n22221,
    n22222, n22223, n22224, n22225, n22226, n22227,
    n22228, n22229, n22230, n22231, n22232, n22233,
    n22234, n22235, n22236, n22237, n22238, n22239,
    n22240, n22241, n22242, n22243, n22244, n22245,
    n22246, n22247, n22248, n22249, n22250, n22251,
    n22252, n22253, n22254, n22255, n22256, n22257,
    n22258, n22259, n22260, n22261, n22262, n22263,
    n22264, n22265, n22266, n22267, n22268, n22269,
    n22270, n22271, n22272, n22273, n22274, n22275,
    n22276, n22277, n22278, n22279, n22280, n22281,
    n22282, n22283, n22284, n22285, n22286, n22287,
    n22288, n22289, n22290, n22291, n22292, n22293,
    n22294, n22295, n22296, n22297, n22298, n22299,
    n22300, n22301, n22302, n22303, n22304, n22305,
    n22306, n22307, n22308, n22309, n22310, n22311,
    n22312, n22313, n22314, n22315, n22316, n22317,
    n22318, n22319, n22320, n22321, n22322, n22323,
    n22324, n22325, n22326, n22327, n22328, n22329,
    n22330, n22331, n22332, n22334, n22335, n22336,
    n22337, n22338, n22339, n22340, n22341, n22342,
    n22343, n22344, n22345, n22346, n22347, n22348,
    n22349, n22350, n22351, n22352, n22353, n22354,
    n22355, n22356, n22357, n22358, n22359, n22360,
    n22361, n22362, n22363, n22364, n22365, n22366,
    n22367, n22368, n22369, n22370, n22371, n22372,
    n22373, n22374, n22375, n22376, n22377, n22378,
    n22379, n22380, n22381, n22382, n22383, n22384,
    n22385, n22386, n22387, n22388, n22389, n22390,
    n22391, n22392, n22393, n22394, n22395, n22396,
    n22397, n22398, n22399, n22400, n22401, n22402,
    n22403, n22404, n22405, n22406, n22407, n22408,
    n22409, n22410, n22411, n22412, n22413, n22414,
    n22415, n22416, n22417, n22418, n22419, n22420,
    n22421, n22422, n22423, n22424, n22425, n22426,
    n22427, n22428, n22429, n22430, n22431, n22432,
    n22433, n22434, n22435, n22436, n22437, n22438,
    n22439, n22440, n22441, n22442, n22443, n22444,
    n22445, n22446, n22447, n22448, n22449, n22450,
    n22451, n22452, n22453, n22454, n22455, n22456,
    n22457, n22458, n22459, n22460, n22461, n22462,
    n22463, n22464, n22465, n22466, n22467, n22468,
    n22469, n22470, n22471, n22472, n22473, n22474,
    n22475, n22476, n22477, n22478, n22479, n22480,
    n22481, n22482, n22483, n22484, n22485, n22486,
    n22487, n22488, n22489, n22490, n22491, n22492,
    n22493, n22494, n22496, n22497, n22498, n22499,
    n22500, n22501, n22502, n22503, n22504, n22505,
    n22506, n22507, n22508, n22509, n22510, n22511,
    n22512, n22513, n22514, n22515, n22516, n22517,
    n22518, n22519, n22520, n22521, n22522, n22523,
    n22524, n22525, n22526, n22527, n22528, n22529,
    n22530, n22531, n22532, n22533, n22534, n22535,
    n22536, n22537, n22538, n22539, n22540, n22541,
    n22542, n22543, n22544, n22545, n22546, n22547,
    n22548, n22549, n22550, n22551, n22552, n22553,
    n22554, n22555, n22556, n22557, n22558, n22559,
    n22560, n22561, n22562, n22563, n22564, n22565,
    n22566, n22567, n22568, n22569, n22570, n22571,
    n22572, n22573, n22574, n22575, n22576, n22577,
    n22578, n22579, n22580, n22581, n22582, n22583,
    n22584, n22585, n22586, n22587, n22588, n22589,
    n22590, n22591, n22592, n22593, n22594, n22595,
    n22596, n22597, n22598, n22599, n22600, n22601,
    n22602, n22603, n22604, n22605, n22606, n22607,
    n22608, n22609, n22610, n22611, n22612, n22613,
    n22614, n22615, n22616, n22617, n22618, n22619,
    n22620, n22621, n22622, n22623, n22624, n22625,
    n22626, n22627, n22628, n22629, n22630, n22631,
    n22632, n22633, n22634, n22635, n22636, n22637,
    n22638, n22639, n22640, n22641, n22642, n22643,
    n22644, n22645, n22646, n22647, n22648, n22649,
    n22650, n22651, n22652, n22653, n22654, n22655,
    n22656, n22657, n22658, n22659, n22661, n22662,
    n22663, n22664, n22665, n22666, n22667, n22668,
    n22669, n22670, n22671, n22672, n22673, n22674,
    n22675, n22676, n22677, n22678, n22679, n22680,
    n22681, n22682, n22683, n22684, n22685, n22686,
    n22687, n22688, n22689, n22690, n22691, n22692,
    n22693, n22694, n22695, n22696, n22697, n22698,
    n22699, n22700, n22701, n22702, n22703, n22704,
    n22705, n22706, n22707, n22708, n22709, n22710,
    n22711, n22712, n22713, n22714, n22715, n22716,
    n22717, n22718, n22719, n22720, n22721, n22722,
    n22723, n22724, n22725, n22726, n22727, n22728,
    n22729, n22730, n22731, n22732, n22733, n22734,
    n22735, n22736, n22737, n22738, n22739, n22740,
    n22741, n22742, n22743, n22744, n22745, n22746,
    n22747, n22748, n22749, n22750, n22751, n22752,
    n22753, n22754, n22755, n22756, n22757, n22758,
    n22759, n22760, n22761, n22762, n22763, n22764,
    n22765, n22766, n22767, n22768, n22769, n22770,
    n22771, n22772, n22773, n22774, n22775, n22776,
    n22777, n22778, n22779, n22780, n22781, n22782,
    n22783, n22784, n22785, n22786, n22787, n22788,
    n22789, n22790, n22791, n22792, n22793, n22794,
    n22795, n22796, n22797, n22798, n22799, n22800,
    n22801, n22802, n22803, n22804, n22805, n22806,
    n22807, n22808, n22809, n22810, n22811, n22812,
    n22813, n22814, n22815, n22817, n22818, n22819,
    n22820, n22821, n22822, n22823, n22824, n22825,
    n22826, n22827, n22828, n22829, n22830, n22831,
    n22832, n22833, n22834, n22835, n22836, n22837,
    n22838, n22839, n22840, n22841, n22842, n22843,
    n22844, n22845, n22846, n22847, n22848, n22849,
    n22850, n22851, n22852, n22853, n22854, n22855,
    n22856, n22857, n22858, n22859, n22860, n22861,
    n22862, n22863, n22864, n22865, n22866, n22867,
    n22868, n22869, n22870, n22871, n22872, n22873,
    n22874, n22875, n22876, n22877, n22878, n22879,
    n22880, n22881, n22882, n22883, n22884, n22885,
    n22886, n22887, n22888, n22889, n22890, n22891,
    n22892, n22893, n22894, n22895, n22896, n22897,
    n22898, n22899, n22900, n22901, n22902, n22903,
    n22904, n22905, n22906, n22907, n22908, n22909,
    n22910, n22911, n22912, n22913, n22914, n22915,
    n22916, n22917, n22918, n22919, n22920, n22921,
    n22922, n22923, n22924, n22925, n22926, n22927,
    n22928, n22929, n22930, n22931, n22932, n22933,
    n22934, n22935, n22936, n22937, n22938, n22939,
    n22940, n22941, n22942, n22943, n22944, n22945,
    n22946, n22947, n22948, n22949, n22950, n22951,
    n22952, n22953, n22954, n22955, n22956, n22957,
    n22958, n22959, n22960, n22961, n22963, n22964,
    n22965, n22966, n22967, n22968, n22969, n22970,
    n22971, n22972, n22973, n22974, n22975, n22976,
    n22977, n22978, n22979, n22980, n22981, n22982,
    n22983, n22984, n22985, n22986, n22987, n22988,
    n22989, n22990, n22991, n22992, n22993, n22994,
    n22995, n22996, n22997, n22998, n22999, n23000,
    n23001, n23002, n23003, n23004, n23005, n23006,
    n23007, n23008, n23009, n23010, n23011, n23012,
    n23013, n23014, n23015, n23016, n23017, n23018,
    n23019, n23020, n23021, n23022, n23023, n23024,
    n23025, n23026, n23027, n23028, n23029, n23030,
    n23031, n23032, n23033, n23034, n23035, n23036,
    n23037, n23038, n23039, n23040, n23041, n23042,
    n23043, n23044, n23045, n23046, n23047, n23048,
    n23049, n23050, n23051, n23052, n23053, n23054,
    n23055, n23056, n23057, n23058, n23059, n23060,
    n23061, n23062, n23063, n23064, n23065, n23066,
    n23067, n23068, n23069, n23070, n23071, n23072,
    n23073, n23074, n23075, n23076, n23077, n23078,
    n23079, n23080, n23081, n23082, n23083, n23084,
    n23085, n23086, n23087, n23088, n23089, n23090,
    n23091, n23092, n23093, n23094, n23095, n23096,
    n23097, n23098, n23099, n23100, n23101, n23102,
    n23103, n23104, n23105, n23106, n23107, n23109,
    n23110, n23111, n23112, n23113, n23114, n23115,
    n23116, n23117, n23118, n23119, n23120, n23121,
    n23122, n23123, n23124, n23125, n23126, n23127,
    n23128, n23129, n23130, n23131, n23132, n23133,
    n23134, n23135, n23136, n23137, n23138, n23139,
    n23140, n23141, n23142, n23143, n23144, n23145,
    n23146, n23147, n23148, n23149, n23150, n23151,
    n23152, n23153, n23154, n23155, n23156, n23157,
    n23158, n23159, n23160, n23161, n23162, n23163,
    n23164, n23165, n23166, n23167, n23168, n23169,
    n23170, n23171, n23172, n23173, n23174, n23175,
    n23176, n23177, n23178, n23179, n23180, n23181,
    n23182, n23183, n23184, n23185, n23186, n23187,
    n23188, n23189, n23190, n23191, n23192, n23193,
    n23194, n23195, n23196, n23197, n23198, n23199,
    n23200, n23201, n23202, n23203, n23204, n23205,
    n23206, n23207, n23208, n23209, n23210, n23211,
    n23212, n23213, n23214, n23215, n23216, n23217,
    n23218, n23219, n23220, n23221, n23222, n23223,
    n23224, n23225, n23226, n23227, n23228, n23229,
    n23230, n23231, n23232, n23233, n23234, n23235,
    n23236, n23237, n23238, n23239, n23240, n23241,
    n23242, n23243, n23244, n23245, n23247, n23248,
    n23249, n23250, n23251, n23252, n23253, n23254,
    n23255, n23256, n23257, n23258, n23259, n23260,
    n23261, n23262, n23263, n23264, n23265, n23266,
    n23267, n23268, n23269, n23270, n23271, n23272,
    n23273, n23274, n23275, n23276, n23277, n23278,
    n23279, n23280, n23281, n23282, n23283, n23284,
    n23285, n23286, n23287, n23288, n23289, n23290,
    n23291, n23292, n23293, n23294, n23295, n23296,
    n23297, n23298, n23299, n23300, n23301, n23302,
    n23303, n23304, n23305, n23306, n23307, n23308,
    n23309, n23310, n23311, n23312, n23313, n23314,
    n23315, n23316, n23317, n23318, n23319, n23320,
    n23321, n23322, n23323, n23324, n23325, n23326,
    n23327, n23328, n23329, n23330, n23331, n23332,
    n23333, n23334, n23335, n23336, n23337, n23338,
    n23339, n23340, n23341, n23342, n23343, n23344,
    n23345, n23346, n23347, n23348, n23349, n23350,
    n23351, n23352, n23353, n23354, n23355, n23356,
    n23357, n23358, n23359, n23360, n23361, n23362,
    n23363, n23364, n23365, n23366, n23367, n23368,
    n23369, n23370, n23371, n23372, n23373, n23375,
    n23376, n23377, n23378, n23379, n23380, n23381,
    n23382, n23383, n23384, n23385, n23386, n23387,
    n23388, n23389, n23390, n23391, n23392, n23393,
    n23394, n23395, n23396, n23397, n23398, n23399,
    n23400, n23401, n23402, n23403, n23404, n23405,
    n23406, n23407, n23408, n23409, n23410, n23411,
    n23412, n23413, n23414, n23415, n23416, n23417,
    n23418, n23419, n23420, n23421, n23422, n23423,
    n23424, n23425, n23426, n23427, n23428, n23429,
    n23430, n23431, n23432, n23433, n23434, n23435,
    n23436, n23437, n23438, n23439, n23440, n23441,
    n23442, n23443, n23444, n23445, n23446, n23447,
    n23448, n23449, n23450, n23451, n23452, n23453,
    n23454, n23455, n23456, n23457, n23458, n23459,
    n23460, n23461, n23462, n23463, n23464, n23465,
    n23466, n23467, n23468, n23469, n23470, n23471,
    n23472, n23473, n23474, n23475, n23476, n23477,
    n23478, n23479, n23480, n23481, n23482, n23483,
    n23484, n23485, n23486, n23487, n23488, n23489,
    n23490, n23491, n23492, n23493, n23494, n23495,
    n23496, n23497, n23498, n23499, n23500, n23501,
    n23502, n23503, n23505, n23506, n23507, n23508,
    n23509, n23510, n23511, n23512, n23513, n23514,
    n23515, n23516, n23517, n23518, n23519, n23520,
    n23521, n23522, n23523, n23524, n23525, n23526,
    n23527, n23528, n23529, n23530, n23531, n23532,
    n23533, n23534, n23535, n23536, n23537, n23538,
    n23539, n23540, n23541, n23542, n23543, n23544,
    n23545, n23546, n23547, n23548, n23549, n23550,
    n23551, n23552, n23553, n23554, n23555, n23556,
    n23557, n23558, n23559, n23560, n23561, n23562,
    n23563, n23564, n23565, n23566, n23567, n23568,
    n23569, n23570, n23571, n23572, n23573, n23574,
    n23575, n23576, n23577, n23578, n23579, n23580,
    n23581, n23582, n23583, n23584, n23585, n23586,
    n23587, n23588, n23589, n23590, n23591, n23592,
    n23593, n23594, n23595, n23596, n23597, n23598,
    n23599, n23600, n23601, n23602, n23603, n23604,
    n23605, n23606, n23607, n23608, n23609, n23610,
    n23611, n23612, n23613, n23614, n23615, n23616,
    n23617, n23618, n23619, n23620, n23621, n23622,
    n23623, n23624, n23626, n23627, n23628, n23629,
    n23630, n23631, n23632, n23633, n23634, n23635,
    n23636, n23637, n23638, n23639, n23640, n23641,
    n23642, n23643, n23644, n23645, n23646, n23647,
    n23648, n23649, n23650, n23651, n23652, n23653,
    n23654, n23655, n23656, n23657, n23658, n23659,
    n23660, n23661, n23662, n23663, n23664, n23665,
    n23666, n23667, n23668, n23669, n23670, n23671,
    n23672, n23673, n23674, n23675, n23676, n23677,
    n23678, n23679, n23680, n23681, n23682, n23683,
    n23684, n23685, n23686, n23687, n23688, n23689,
    n23690, n23691, n23692, n23693, n23694, n23695,
    n23696, n23697, n23698, n23699, n23700, n23701,
    n23702, n23703, n23704, n23705, n23706, n23707,
    n23708, n23709, n23710, n23711, n23712, n23713,
    n23714, n23715, n23716, n23717, n23718, n23719,
    n23720, n23721, n23722, n23723, n23724, n23725,
    n23726, n23727, n23728, n23729, n23730, n23731,
    n23732, n23733, n23734, n23735, n23736, n23738,
    n23739, n23740, n23741, n23742, n23743, n23744,
    n23745, n23746, n23747, n23748, n23749, n23750,
    n23751, n23752, n23753, n23754, n23755, n23756,
    n23757, n23758, n23759, n23760, n23761, n23762,
    n23763, n23764, n23765, n23766, n23767, n23768,
    n23769, n23770, n23771, n23772, n23773, n23774,
    n23775, n23776, n23777, n23778, n23779, n23780,
    n23781, n23782, n23783, n23784, n23785, n23786,
    n23787, n23788, n23789, n23790, n23791, n23792,
    n23793, n23794, n23795, n23796, n23797, n23798,
    n23799, n23800, n23801, n23802, n23803, n23804,
    n23805, n23806, n23807, n23808, n23809, n23810,
    n23811, n23812, n23813, n23814, n23815, n23816,
    n23817, n23818, n23819, n23820, n23821, n23822,
    n23823, n23824, n23825, n23826, n23827, n23828,
    n23829, n23830, n23831, n23832, n23833, n23834,
    n23835, n23836, n23837, n23838, n23839, n23840,
    n23841, n23842, n23843, n23844, n23845, n23846,
    n23847, n23849, n23850, n23851, n23852, n23853,
    n23854, n23855, n23856, n23857, n23858, n23859,
    n23860, n23861, n23862, n23863, n23864, n23865,
    n23866, n23867, n23868, n23869, n23870, n23871,
    n23872, n23873, n23874, n23875, n23876, n23877,
    n23878, n23879, n23880, n23881, n23882, n23883,
    n23884, n23885, n23886, n23887, n23888, n23889,
    n23890, n23891, n23892, n23893, n23894, n23895,
    n23896, n23897, n23898, n23899, n23900, n23901,
    n23902, n23903, n23904, n23905, n23906, n23907,
    n23908, n23909, n23910, n23911, n23912, n23913,
    n23914, n23915, n23916, n23917, n23918, n23919,
    n23920, n23921, n23922, n23923, n23924, n23925,
    n23926, n23927, n23928, n23929, n23930, n23931,
    n23932, n23933, n23934, n23935, n23936, n23937,
    n23938, n23939, n23940, n23941, n23942, n23943,
    n23944, n23945, n23946, n23947, n23948, n23949,
    n23950, n23951, n23952, n23954, n23955, n23956,
    n23957, n23958, n23959, n23960, n23961, n23962,
    n23963, n23964, n23965, n23966, n23967, n23968,
    n23969, n23970, n23971, n23972, n23973, n23974,
    n23975, n23976, n23977, n23978, n23979, n23980,
    n23981, n23982, n23983, n23984, n23985, n23986,
    n23987, n23988, n23989, n23990, n23991, n23992,
    n23993, n23994, n23995, n23996, n23997, n23998,
    n23999, n24000, n24001, n24002, n24003, n24004,
    n24005, n24006, n24007, n24008, n24009, n24010,
    n24011, n24012, n24013, n24014, n24015, n24016,
    n24017, n24018, n24019, n24020, n24021, n24022,
    n24023, n24024, n24025, n24026, n24027, n24028,
    n24029, n24030, n24031, n24032, n24033, n24034,
    n24035, n24036, n24037, n24038, n24039, n24040,
    n24041, n24042, n24043, n24044, n24045, n24046,
    n24048, n24049, n24050, n24051, n24052, n24053,
    n24054, n24055, n24056, n24057, n24058, n24059,
    n24060, n24061, n24062, n24063, n24064, n24065,
    n24066, n24067, n24068, n24069, n24070, n24071,
    n24072, n24073, n24074, n24075, n24076, n24077,
    n24078, n24079, n24080, n24081, n24082, n24083,
    n24084, n24085, n24086, n24087, n24088, n24089,
    n24090, n24091, n24092, n24093, n24094, n24095,
    n24096, n24097, n24098, n24099, n24100, n24101,
    n24102, n24103, n24104, n24105, n24106, n24107,
    n24108, n24109, n24110, n24111, n24112, n24113,
    n24114, n24115, n24116, n24117, n24118, n24119,
    n24120, n24121, n24122, n24123, n24124, n24125,
    n24126, n24127, n24128, n24129, n24130, n24131,
    n24132, n24133, n24134, n24135, n24136, n24137,
    n24138, n24140, n24141, n24142, n24143, n24144,
    n24145, n24146, n24147, n24148, n24149, n24150,
    n24151, n24152, n24153, n24154, n24155, n24156,
    n24157, n24158, n24159, n24160, n24161, n24162,
    n24163, n24164, n24165, n24166, n24167, n24168,
    n24169, n24170, n24171, n24172, n24173, n24174,
    n24175, n24176, n24177, n24178, n24179, n24180,
    n24181, n24182, n24183, n24184, n24185, n24186,
    n24187, n24188, n24189, n24190, n24191, n24192,
    n24193, n24194, n24195, n24196, n24197, n24198,
    n24199, n24200, n24201, n24202, n24203, n24204,
    n24205, n24206, n24207, n24208, n24209, n24210,
    n24211, n24212, n24213, n24214, n24215, n24216,
    n24217, n24218, n24219, n24220, n24221, n24222,
    n24223, n24224, n24225, n24226, n24228, n24229,
    n24230, n24231, n24232, n24233, n24234, n24235,
    n24236, n24237, n24238, n24239, n24240, n24241,
    n24242, n24243, n24244, n24245, n24246, n24247,
    n24248, n24249, n24250, n24251, n24252, n24253,
    n24254, n24255, n24256, n24257, n24258, n24259,
    n24260, n24261, n24262, n24263, n24264, n24265,
    n24266, n24267, n24268, n24269, n24270, n24271,
    n24272, n24273, n24274, n24275, n24276, n24277,
    n24278, n24279, n24280, n24281, n24282, n24283,
    n24284, n24285, n24286, n24287, n24288, n24289,
    n24290, n24291, n24292, n24293, n24294, n24295,
    n24296, n24297, n24298, n24299, n24300, n24301,
    n24302, n24303, n24305, n24306, n24307, n24308,
    n24309, n24310, n24311, n24312, n24313, n24314,
    n24315, n24316, n24317, n24318, n24319, n24320,
    n24321, n24322, n24323, n24324, n24325, n24326,
    n24327, n24328, n24329, n24330, n24331, n24332,
    n24333, n24334, n24335, n24336, n24337, n24338,
    n24339, n24340, n24341, n24342, n24343, n24344,
    n24345, n24346, n24347, n24348, n24349, n24350,
    n24351, n24352, n24353, n24354, n24355, n24356,
    n24357, n24358, n24359, n24360, n24361, n24362,
    n24363, n24364, n24365, n24366, n24367, n24368,
    n24369, n24370, n24371, n24372, n24373, n24374,
    n24375, n24376, n24377, n24378, n24380, n24381,
    n24382, n24383, n24384, n24385, n24386, n24387,
    n24388, n24389, n24390, n24391, n24392, n24393,
    n24394, n24395, n24396, n24397, n24398, n24399,
    n24400, n24401, n24402, n24403, n24404, n24405,
    n24406, n24407, n24408, n24409, n24410, n24411,
    n24412, n24413, n24414, n24415, n24416, n24417,
    n24418, n24419, n24420, n24421, n24422, n24423,
    n24424, n24425, n24426, n24427, n24428, n24429,
    n24430, n24431, n24432, n24433, n24434, n24435,
    n24436, n24437, n24438, n24439, n24440, n24441,
    n24442, n24443, n24444, n24445, n24446, n24447,
    n24448, n24450, n24451, n24452, n24453, n24454,
    n24455, n24456, n24457, n24458, n24459, n24460,
    n24461, n24462, n24463, n24464, n24465, n24466,
    n24467, n24468, n24469, n24470, n24471, n24472,
    n24473, n24474, n24475, n24476, n24477, n24478,
    n24479, n24480, n24481, n24482, n24483, n24484,
    n24485, n24486, n24487, n24488, n24489, n24490,
    n24491, n24492, n24493, n24494, n24495, n24496,
    n24497, n24498, n24499, n24500, n24501, n24502,
    n24503, n24504, n24505, n24506, n24507, n24508,
    n24510, n24511, n24512, n24513, n24514, n24515,
    n24516, n24517, n24518, n24519, n24520, n24521,
    n24522, n24523, n24524, n24525, n24526, n24527,
    n24528, n24529, n24530, n24531, n24532, n24533,
    n24534, n24535, n24536, n24537, n24538, n24539,
    n24540, n24541, n24542, n24543, n24544, n24545,
    n24546, n24547, n24548, n24549, n24550, n24551,
    n24552, n24553, n24554, n24555, n24556, n24557,
    n24558, n24559, n24560, n24561, n24562, n24563,
    n24564, n24565, n24566, n24568, n24569, n24570,
    n24571, n24572, n24573, n24574, n24575, n24576,
    n24577, n24578, n24579, n24580, n24581, n24582,
    n24583, n24584, n24585, n24586, n24587, n24588,
    n24589, n24590, n24591, n24592, n24593, n24594,
    n24595, n24596, n24597, n24598, n24599, n24600,
    n24601, n24602, n24603, n24604, n24605, n24606,
    n24607, n24608, n24609, n24610, n24611, n24612,
    n24613, n24614, n24615, n24616, n24617, n24618,
    n24619, n24621, n24622, n24623, n24624, n24625,
    n24626, n24627, n24628, n24629, n24630, n24631,
    n24632, n24633, n24634, n24635, n24636, n24637,
    n24638, n24639, n24640, n24641, n24642, n24643,
    n24644, n24645, n24646, n24647, n24648, n24649,
    n24650, n24651, n24652, n24653, n24654, n24655,
    n24656, n24657, n24658, n24659, n24660, n24661,
    n24662, n24664, n24665, n24666, n24667, n24668,
    n24669, n24670, n24671, n24672, n24673, n24674,
    n24675, n24676, n24677, n24678, n24679, n24680,
    n24681, n24682, n24683, n24684, n24685, n24686,
    n24687, n24688, n24689, n24690, n24691, n24692,
    n24693, n24694, n24695, n24696, n24697, n24698,
    n24699, n24700, n24701, n24702, n24703, n24705,
    n24706, n24707, n24708, n24709, n24710, n24711,
    n24712, n24713, n24714, n24715, n24716, n24717,
    n24718, n24719, n24720, n24721, n24722, n24723,
    n24724, n24725, n24726, n24727, n24728, n24729,
    n24730, n24731, n24732, n24733, n24734, n24735,
    n24736, n24737, n24739, n24740, n24741, n24742,
    n24743, n24744, n24745, n24746, n24747, n24748,
    n24749, n24750, n24751, n24752, n24753, n24754,
    n24755, n24756, n24757, n24758, n24759, n24760,
    n24761, n24762, n24763, n24765, n24766, n24767,
    n24768, n24769, n24770, n24771, n24772, n24773,
    n24774, n24775, n24776, n24777, n24778, n24779,
    n24780, n24781, n24782, n24783, n24784, n24785,
    n24786, n24788, n24789, n24790, n24791, n24792,
    n24793, n24794, n24795, n24796, n24797, n24798,
    n24799, n24800, n24801, n24802, n24803, n24805,
    n24806, n24807, n24808, n24809, n24810, n24811;
  assign po0  = pi0  & pi64 ;
  assign n258 = pi2  & po0 ;
  assign n259 = ~pi1  & ~pi2 ;
  assign n260 = pi1  & pi2 ;
  assign n261 = ~n259 & ~n260;
  assign n262 = pi0  & n261;
  assign n263 = pi64  & pi65 ;
  assign n264 = ~pi64  & ~pi65 ;
  assign n265 = ~n263 & ~n264;
  assign n266 = n262 & n265;
  assign n267 = ~pi0  & pi1 ;
  assign n268 = pi64  & n267;
  assign n269 = pi0  & ~n261;
  assign n270 = pi65  & n269;
  assign n271 = ~n266 & ~n268;
  assign n272 = ~n270 & n271;
  assign n273 = n258 & ~n272;
  assign n274 = ~n258 & n272;
  assign po1  = ~n273 & ~n274;
  assign n276 = pi2  & ~po0 ;
  assign n277 = n272 & n276;
  assign n278 = pi2  & ~n277;
  assign n279 = pi66  & n269;
  assign n280 = pi65  & n267;
  assign n281 = ~pi0  & ~pi1 ;
  assign n282 = n261 & n281;
  assign n283 = pi64  & n282;
  assign n284 = ~pi64  & pi65 ;
  assign n285 = pi66  & ~n284;
  assign n286 = ~pi66  & n284;
  assign n287 = ~n285 & ~n286;
  assign n288 = n262 & ~n287;
  assign n289 = ~n279 & ~n280;
  assign n290 = ~n283 & ~n288;
  assign n291 = n289 & n290;
  assign n292 = ~n278 & n291;
  assign n293 = n278 & ~n291;
  assign po2  = ~n292 & ~n293;
  assign n295 = pi67  & n269;
  assign n296 = pi66  & n267;
  assign n297 = pi65  & n282;
  assign n298 = ~pi66  & ~pi67 ;
  assign n299 = pi66  & pi67 ;
  assign n300 = ~n298 & ~n299;
  assign n301 = ~pi64  & ~pi66 ;
  assign n302 = pi65  & ~n301;
  assign n303 = n300 & n302;
  assign n304 = ~n300 & ~n302;
  assign n305 = ~n303 & ~n304;
  assign n306 = n262 & n305;
  assign n307 = ~n295 & ~n296;
  assign n308 = ~n297 & n307;
  assign n309 = ~n306 & n308;
  assign n310 = pi2  & n309;
  assign n311 = ~pi2  & ~n309;
  assign n312 = ~n310 & ~n311;
  assign n313 = ~pi2  & ~pi3 ;
  assign n314 = pi2  & pi3 ;
  assign n315 = ~n313 & ~n314;
  assign n316 = pi64  & n315;
  assign n317 = ~n312 & n316;
  assign n318 = n312 & ~n316;
  assign n319 = ~n317 & ~n318;
  assign n320 = n277 & n291;
  assign n321 = n319 & n320;
  assign n322 = ~n319 & ~n320;
  assign po3  = ~n321 & ~n322;
  assign n324 = ~n317 & ~n321;
  assign n325 = pi68  & n269;
  assign n326 = pi67  & n267;
  assign n327 = pi66  & n282;
  assign n328 = ~n299 & ~n303;
  assign n329 = ~pi67  & ~pi68 ;
  assign n330 = pi67  & pi68 ;
  assign n331 = ~n329 & ~n330;
  assign n332 = ~n328 & n331;
  assign n333 = n328 & ~n331;
  assign n334 = ~n332 & ~n333;
  assign n335 = n262 & n334;
  assign n336 = ~n325 & ~n326;
  assign n337 = ~n327 & n336;
  assign n338 = ~n335 & n337;
  assign n339 = pi2  & n338;
  assign n340 = ~pi2  & ~n338;
  assign n341 = ~n339 & ~n340;
  assign n342 = pi5  & n316;
  assign n343 = ~pi4  & ~pi5 ;
  assign n344 = pi4  & pi5 ;
  assign n345 = ~n343 & ~n344;
  assign n346 = n315 & n345;
  assign n347 = n265 & n346;
  assign n348 = n315 & ~n345;
  assign n349 = pi65  & n348;
  assign n350 = ~pi3  & ~pi4 ;
  assign n351 = pi3  & pi4 ;
  assign n352 = ~n350 & ~n351;
  assign n353 = ~n315 & n352;
  assign n354 = pi64  & n353;
  assign n355 = ~n347 & ~n349;
  assign n356 = ~n354 & n355;
  assign n357 = n342 & ~n356;
  assign n358 = ~n342 & n356;
  assign n359 = ~n357 & ~n358;
  assign n360 = ~n341 & n359;
  assign n361 = n341 & ~n359;
  assign n362 = ~n360 & ~n361;
  assign n363 = ~n324 & n362;
  assign n364 = n324 & ~n362;
  assign po4  = ~n363 & ~n364;
  assign n366 = ~n360 & ~n363;
  assign n367 = pi69  & n269;
  assign n368 = pi68  & n267;
  assign n369 = pi67  & n282;
  assign n370 = ~n330 & ~n332;
  assign n371 = ~pi68  & ~pi69 ;
  assign n372 = pi68  & pi69 ;
  assign n373 = ~n371 & ~n372;
  assign n374 = ~n370 & n373;
  assign n375 = n370 & ~n373;
  assign n376 = ~n374 & ~n375;
  assign n377 = n262 & n376;
  assign n378 = ~n367 & ~n368;
  assign n379 = ~n369 & n378;
  assign n380 = ~n377 & n379;
  assign n381 = pi2  & n380;
  assign n382 = ~pi2  & ~n380;
  assign n383 = ~n381 & ~n382;
  assign n384 = pi5  & ~n316;
  assign n385 = n356 & n384;
  assign n386 = pi5  & ~n385;
  assign n387 = pi66  & n348;
  assign n388 = pi65  & n353;
  assign n389 = ~n287 & n346;
  assign n390 = ~n315 & n345;
  assign n391 = ~n352 & n390;
  assign n392 = pi64  & n391;
  assign n393 = ~n387 & ~n388;
  assign n394 = ~n389 & n393;
  assign n395 = ~n392 & n394;
  assign n396 = ~n386 & n395;
  assign n397 = n386 & ~n395;
  assign n398 = ~n396 & ~n397;
  assign n399 = ~n383 & n398;
  assign n400 = n383 & ~n398;
  assign n401 = ~n399 & ~n400;
  assign n402 = ~n366 & n401;
  assign n403 = n366 & ~n401;
  assign po5  = ~n402 & ~n403;
  assign n405 = ~n399 & ~n402;
  assign n406 = pi70  & n269;
  assign n407 = pi69  & n267;
  assign n408 = pi68  & n282;
  assign n409 = ~n372 & ~n374;
  assign n410 = ~pi69  & ~pi70 ;
  assign n411 = pi69  & pi70 ;
  assign n412 = ~n410 & ~n411;
  assign n413 = ~n409 & n412;
  assign n414 = n409 & ~n412;
  assign n415 = ~n413 & ~n414;
  assign n416 = n262 & n415;
  assign n417 = ~n406 & ~n407;
  assign n418 = ~n408 & n417;
  assign n419 = ~n416 & n418;
  assign n420 = pi2  & n419;
  assign n421 = ~pi2  & ~n419;
  assign n422 = ~n420 & ~n421;
  assign n423 = pi65  & n391;
  assign n424 = pi66  & n353;
  assign n425 = pi67  & n348;
  assign n426 = n305 & n346;
  assign n427 = ~n424 & ~n425;
  assign n428 = ~n423 & n427;
  assign n429 = ~n426 & n428;
  assign n430 = pi5  & n429;
  assign n431 = ~pi5  & ~n429;
  assign n432 = ~n430 & ~n431;
  assign n433 = ~pi5  & ~pi6 ;
  assign n434 = pi5  & pi6 ;
  assign n435 = ~n433 & ~n434;
  assign n436 = pi64  & n435;
  assign n437 = n385 & n395;
  assign n438 = n436 & n437;
  assign n439 = ~n436 & ~n437;
  assign n440 = ~n438 & ~n439;
  assign n441 = ~n432 & n440;
  assign n442 = n432 & ~n440;
  assign n443 = ~n441 & ~n442;
  assign n444 = ~n422 & n443;
  assign n445 = n422 & ~n443;
  assign n446 = ~n444 & ~n445;
  assign n447 = ~n405 & n446;
  assign n448 = n405 & ~n446;
  assign po6  = ~n447 & ~n448;
  assign n450 = ~n444 & ~n447;
  assign n451 = pi71  & n269;
  assign n452 = pi70  & n267;
  assign n453 = pi69  & n282;
  assign n454 = ~n411 & ~n413;
  assign n455 = ~pi70  & ~pi71 ;
  assign n456 = pi70  & pi71 ;
  assign n457 = ~n455 & ~n456;
  assign n458 = ~n454 & n457;
  assign n459 = n454 & ~n457;
  assign n460 = ~n458 & ~n459;
  assign n461 = n262 & n460;
  assign n462 = ~n451 & ~n452;
  assign n463 = ~n453 & n462;
  assign n464 = ~n461 & n463;
  assign n465 = pi2  & n464;
  assign n466 = ~pi2  & ~n464;
  assign n467 = ~n465 & ~n466;
  assign n468 = ~n438 & ~n441;
  assign n469 = pi66  & n391;
  assign n470 = pi67  & n353;
  assign n471 = pi68  & n348;
  assign n472 = n334 & n346;
  assign n473 = ~n470 & ~n471;
  assign n474 = ~n469 & n473;
  assign n475 = ~n472 & n474;
  assign n476 = pi5  & n475;
  assign n477 = ~pi5  & ~n475;
  assign n478 = ~n476 & ~n477;
  assign n479 = pi8  & n436;
  assign n480 = ~pi7  & ~pi8 ;
  assign n481 = pi7  & pi8 ;
  assign n482 = ~n480 & ~n481;
  assign n483 = n435 & n482;
  assign n484 = n265 & n483;
  assign n485 = n435 & ~n482;
  assign n486 = pi65  & n485;
  assign n487 = ~pi6  & ~pi7 ;
  assign n488 = pi6  & pi7 ;
  assign n489 = ~n487 & ~n488;
  assign n490 = ~n435 & n489;
  assign n491 = pi64  & n490;
  assign n492 = ~n484 & ~n486;
  assign n493 = ~n491 & n492;
  assign n494 = n479 & ~n493;
  assign n495 = ~n479 & n493;
  assign n496 = ~n494 & ~n495;
  assign n497 = ~n478 & n496;
  assign n498 = n478 & ~n496;
  assign n499 = ~n497 & ~n498;
  assign n500 = ~n468 & n499;
  assign n501 = n468 & ~n499;
  assign n502 = ~n500 & ~n501;
  assign n503 = ~n467 & n502;
  assign n504 = n467 & ~n502;
  assign n505 = ~n503 & ~n504;
  assign n506 = ~n450 & n505;
  assign n507 = n450 & ~n505;
  assign po7  = ~n506 & ~n507;
  assign n509 = ~n503 & ~n506;
  assign n510 = ~n497 & ~n500;
  assign n511 = pi67  & n391;
  assign n512 = pi68  & n353;
  assign n513 = pi69  & n348;
  assign n514 = n346 & n376;
  assign n515 = ~n512 & ~n513;
  assign n516 = ~n511 & n515;
  assign n517 = ~n514 & n516;
  assign n518 = pi5  & n517;
  assign n519 = ~pi5  & ~n517;
  assign n520 = ~n518 & ~n519;
  assign n521 = pi8  & ~n436;
  assign n522 = n493 & n521;
  assign n523 = pi8  & ~n522;
  assign n524 = ~n287 & n483;
  assign n525 = pi65  & n490;
  assign n526 = pi66  & n485;
  assign n527 = ~n435 & n482;
  assign n528 = ~n489 & n527;
  assign n529 = pi64  & n528;
  assign n530 = ~n524 & ~n525;
  assign n531 = ~n526 & n530;
  assign n532 = ~n529 & n531;
  assign n533 = ~n523 & n532;
  assign n534 = n523 & ~n532;
  assign n535 = ~n533 & ~n534;
  assign n536 = ~n520 & n535;
  assign n537 = n520 & ~n535;
  assign n538 = ~n536 & ~n537;
  assign n539 = n510 & ~n538;
  assign n540 = ~n510 & n538;
  assign n541 = ~n539 & ~n540;
  assign n542 = pi72  & n269;
  assign n543 = pi71  & n267;
  assign n544 = pi70  & n282;
  assign n545 = ~n456 & ~n458;
  assign n546 = ~pi71  & ~pi72 ;
  assign n547 = pi71  & pi72 ;
  assign n548 = ~n546 & ~n547;
  assign n549 = ~n545 & n548;
  assign n550 = n545 & ~n548;
  assign n551 = ~n549 & ~n550;
  assign n552 = n262 & n551;
  assign n553 = ~n542 & ~n543;
  assign n554 = ~n544 & n553;
  assign n555 = ~n552 & n554;
  assign n556 = pi2  & n555;
  assign n557 = ~pi2  & ~n555;
  assign n558 = ~n556 & ~n557;
  assign n559 = n541 & ~n558;
  assign n560 = ~n541 & n558;
  assign n561 = ~n559 & ~n560;
  assign n562 = ~n509 & n561;
  assign n563 = n509 & ~n561;
  assign po8  = ~n562 & ~n563;
  assign n565 = ~n559 & ~n562;
  assign n566 = ~n536 & ~n540;
  assign n567 = pi65  & n528;
  assign n568 = pi66  & n490;
  assign n569 = pi67  & n485;
  assign n570 = n305 & n483;
  assign n571 = ~n568 & ~n569;
  assign n572 = ~n567 & n571;
  assign n573 = ~n570 & n572;
  assign n574 = pi8  & n573;
  assign n575 = ~pi8  & ~n573;
  assign n576 = ~n574 & ~n575;
  assign n577 = ~pi8  & ~pi9 ;
  assign n578 = pi8  & pi9 ;
  assign n579 = ~n577 & ~n578;
  assign n580 = pi64  & n579;
  assign n581 = n522 & n532;
  assign n582 = n580 & n581;
  assign n583 = ~n580 & ~n581;
  assign n584 = ~n582 & ~n583;
  assign n585 = ~n576 & n584;
  assign n586 = n576 & ~n584;
  assign n587 = ~n585 & ~n586;
  assign n588 = pi68  & n391;
  assign n589 = pi69  & n353;
  assign n590 = pi70  & n348;
  assign n591 = n346 & n415;
  assign n592 = ~n589 & ~n590;
  assign n593 = ~n588 & n592;
  assign n594 = ~n591 & n593;
  assign n595 = pi5  & n594;
  assign n596 = ~pi5  & ~n594;
  assign n597 = ~n595 & ~n596;
  assign n598 = n587 & ~n597;
  assign n599 = ~n587 & n597;
  assign n600 = ~n598 & ~n599;
  assign n601 = n566 & ~n600;
  assign n602 = ~n566 & n600;
  assign n603 = ~n601 & ~n602;
  assign n604 = pi73  & n269;
  assign n605 = pi72  & n267;
  assign n606 = pi71  & n282;
  assign n607 = ~n547 & ~n549;
  assign n608 = ~pi72  & ~pi73 ;
  assign n609 = pi72  & pi73 ;
  assign n610 = ~n608 & ~n609;
  assign n611 = ~n607 & n610;
  assign n612 = n607 & ~n610;
  assign n613 = ~n611 & ~n612;
  assign n614 = n262 & n613;
  assign n615 = ~n604 & ~n605;
  assign n616 = ~n606 & n615;
  assign n617 = ~n614 & n616;
  assign n618 = pi2  & n617;
  assign n619 = ~pi2  & ~n617;
  assign n620 = ~n618 & ~n619;
  assign n621 = n603 & ~n620;
  assign n622 = ~n603 & n620;
  assign n623 = ~n621 & ~n622;
  assign n624 = ~n565 & n623;
  assign n625 = n565 & ~n623;
  assign po9  = ~n624 & ~n625;
  assign n627 = ~n621 & ~n624;
  assign n628 = ~n598 & ~n602;
  assign n629 = ~n582 & ~n585;
  assign n630 = pi66  & n528;
  assign n631 = pi67  & n490;
  assign n632 = pi68  & n485;
  assign n633 = n334 & n483;
  assign n634 = ~n631 & ~n632;
  assign n635 = ~n630 & n634;
  assign n636 = ~n633 & n635;
  assign n637 = pi8  & n636;
  assign n638 = ~pi8  & ~n636;
  assign n639 = ~n637 & ~n638;
  assign n640 = pi11  & n580;
  assign n641 = ~pi10  & ~pi11 ;
  assign n642 = pi10  & pi11 ;
  assign n643 = ~n641 & ~n642;
  assign n644 = n579 & n643;
  assign n645 = n265 & n644;
  assign n646 = n579 & ~n643;
  assign n647 = pi65  & n646;
  assign n648 = ~pi9  & ~pi10 ;
  assign n649 = pi9  & pi10 ;
  assign n650 = ~n648 & ~n649;
  assign n651 = ~n579 & n650;
  assign n652 = pi64  & n651;
  assign n653 = ~n645 & ~n647;
  assign n654 = ~n652 & n653;
  assign n655 = n640 & ~n654;
  assign n656 = ~n640 & n654;
  assign n657 = ~n655 & ~n656;
  assign n658 = n639 & ~n657;
  assign n659 = ~n639 & n657;
  assign n660 = ~n658 & ~n659;
  assign n661 = ~n629 & n660;
  assign n662 = n629 & ~n660;
  assign n663 = ~n661 & ~n662;
  assign n664 = pi69  & n391;
  assign n665 = pi70  & n353;
  assign n666 = pi71  & n348;
  assign n667 = n346 & n460;
  assign n668 = ~n665 & ~n666;
  assign n669 = ~n664 & n668;
  assign n670 = ~n667 & n669;
  assign n671 = pi5  & n670;
  assign n672 = ~pi5  & ~n670;
  assign n673 = ~n671 & ~n672;
  assign n674 = n663 & ~n673;
  assign n675 = ~n663 & n673;
  assign n676 = ~n674 & ~n675;
  assign n677 = n628 & ~n676;
  assign n678 = ~n628 & n676;
  assign n679 = ~n677 & ~n678;
  assign n680 = pi74  & n269;
  assign n681 = pi73  & n267;
  assign n682 = pi72  & n282;
  assign n683 = ~n609 & ~n611;
  assign n684 = ~pi73  & ~pi74 ;
  assign n685 = pi73  & pi74 ;
  assign n686 = ~n684 & ~n685;
  assign n687 = ~n683 & n686;
  assign n688 = n683 & ~n686;
  assign n689 = ~n687 & ~n688;
  assign n690 = n262 & n689;
  assign n691 = ~n680 & ~n681;
  assign n692 = ~n682 & n691;
  assign n693 = ~n690 & n692;
  assign n694 = pi2  & n693;
  assign n695 = ~pi2  & ~n693;
  assign n696 = ~n694 & ~n695;
  assign n697 = ~n679 & n696;
  assign n698 = n679 & ~n696;
  assign n699 = ~n697 & ~n698;
  assign n700 = ~n627 & n699;
  assign n701 = n627 & ~n699;
  assign po10  = ~n700 & ~n701;
  assign n703 = ~n698 & ~n700;
  assign n704 = pi75  & n269;
  assign n705 = pi74  & n267;
  assign n706 = pi73  & n282;
  assign n707 = ~n685 & ~n687;
  assign n708 = ~pi74  & ~pi75 ;
  assign n709 = pi74  & pi75 ;
  assign n710 = ~n708 & ~n709;
  assign n711 = ~n707 & n710;
  assign n712 = n707 & ~n710;
  assign n713 = ~n711 & ~n712;
  assign n714 = n262 & n713;
  assign n715 = ~n704 & ~n705;
  assign n716 = ~n706 & n715;
  assign n717 = ~n714 & n716;
  assign n718 = pi2  & n717;
  assign n719 = ~pi2  & ~n717;
  assign n720 = ~n718 & ~n719;
  assign n721 = ~n674 & ~n678;
  assign n722 = pi70  & n391;
  assign n723 = pi71  & n353;
  assign n724 = pi72  & n348;
  assign n725 = n346 & n551;
  assign n726 = ~n723 & ~n724;
  assign n727 = ~n722 & n726;
  assign n728 = ~n725 & n727;
  assign n729 = pi5  & n728;
  assign n730 = ~pi5  & ~n728;
  assign n731 = ~n729 & ~n730;
  assign n732 = ~n659 & ~n661;
  assign n733 = pi67  & n528;
  assign n734 = pi68  & n490;
  assign n735 = pi69  & n485;
  assign n736 = n376 & n483;
  assign n737 = ~n734 & ~n735;
  assign n738 = ~n733 & n737;
  assign n739 = ~n736 & n738;
  assign n740 = pi8  & n739;
  assign n741 = ~pi8  & ~n739;
  assign n742 = ~n740 & ~n741;
  assign n743 = pi11  & ~n580;
  assign n744 = n654 & n743;
  assign n745 = pi11  & ~n744;
  assign n746 = ~n287 & n644;
  assign n747 = pi65  & n651;
  assign n748 = pi66  & n646;
  assign n749 = ~n579 & n643;
  assign n750 = ~n650 & n749;
  assign n751 = pi64  & n750;
  assign n752 = ~n746 & ~n747;
  assign n753 = ~n748 & n752;
  assign n754 = ~n751 & n753;
  assign n755 = ~n745 & n754;
  assign n756 = n745 & ~n754;
  assign n757 = ~n755 & ~n756;
  assign n758 = ~n742 & n757;
  assign n759 = n742 & ~n757;
  assign n760 = ~n758 & ~n759;
  assign n761 = ~n732 & n760;
  assign n762 = n732 & ~n760;
  assign n763 = ~n761 & ~n762;
  assign n764 = ~n731 & n763;
  assign n765 = n731 & ~n763;
  assign n766 = ~n764 & ~n765;
  assign n767 = ~n721 & n766;
  assign n768 = n721 & ~n766;
  assign n769 = ~n767 & ~n768;
  assign n770 = ~n720 & n769;
  assign n771 = n720 & ~n769;
  assign n772 = ~n770 & ~n771;
  assign n773 = ~n703 & n772;
  assign n774 = n703 & ~n772;
  assign po11  = ~n773 & ~n774;
  assign n776 = ~n770 & ~n773;
  assign n777 = ~n758 & ~n761;
  assign n778 = pi65  & n750;
  assign n779 = pi66  & n651;
  assign n780 = pi67  & n646;
  assign n781 = n305 & n644;
  assign n782 = ~n779 & ~n780;
  assign n783 = ~n778 & n782;
  assign n784 = ~n781 & n783;
  assign n785 = pi11  & n784;
  assign n786 = ~pi11  & ~n784;
  assign n787 = ~n785 & ~n786;
  assign n788 = ~pi11  & ~pi12 ;
  assign n789 = pi11  & pi12 ;
  assign n790 = ~n788 & ~n789;
  assign n791 = pi64  & n790;
  assign n792 = n744 & n754;
  assign n793 = n791 & n792;
  assign n794 = ~n791 & ~n792;
  assign n795 = ~n793 & ~n794;
  assign n796 = ~n787 & n795;
  assign n797 = n787 & ~n795;
  assign n798 = ~n796 & ~n797;
  assign n799 = pi68  & n528;
  assign n800 = pi69  & n490;
  assign n801 = pi70  & n485;
  assign n802 = n415 & n483;
  assign n803 = ~n800 & ~n801;
  assign n804 = ~n799 & n803;
  assign n805 = ~n802 & n804;
  assign n806 = pi8  & n805;
  assign n807 = ~pi8  & ~n805;
  assign n808 = ~n806 & ~n807;
  assign n809 = n798 & ~n808;
  assign n810 = ~n798 & n808;
  assign n811 = ~n809 & ~n810;
  assign n812 = n777 & ~n811;
  assign n813 = ~n777 & n811;
  assign n814 = ~n812 & ~n813;
  assign n815 = pi71  & n391;
  assign n816 = pi72  & n353;
  assign n817 = pi73  & n348;
  assign n818 = n346 & n613;
  assign n819 = ~n816 & ~n817;
  assign n820 = ~n815 & n819;
  assign n821 = ~n818 & n820;
  assign n822 = pi5  & n821;
  assign n823 = ~pi5  & ~n821;
  assign n824 = ~n822 & ~n823;
  assign n825 = ~n814 & n824;
  assign n826 = n814 & ~n824;
  assign n827 = ~n825 & ~n826;
  assign n828 = ~n764 & ~n767;
  assign n829 = n827 & ~n828;
  assign n830 = ~n827 & n828;
  assign n831 = ~n829 & ~n830;
  assign n832 = pi76  & n269;
  assign n833 = pi75  & n267;
  assign n834 = pi74  & n282;
  assign n835 = ~n709 & ~n711;
  assign n836 = ~pi75  & ~pi76 ;
  assign n837 = pi75  & pi76 ;
  assign n838 = ~n836 & ~n837;
  assign n839 = ~n835 & n838;
  assign n840 = n835 & ~n838;
  assign n841 = ~n839 & ~n840;
  assign n842 = n262 & n841;
  assign n843 = ~n832 & ~n833;
  assign n844 = ~n834 & n843;
  assign n845 = ~n842 & n844;
  assign n846 = pi2  & n845;
  assign n847 = ~pi2  & ~n845;
  assign n848 = ~n846 & ~n847;
  assign n849 = n831 & ~n848;
  assign n850 = ~n831 & n848;
  assign n851 = ~n849 & ~n850;
  assign n852 = ~n776 & n851;
  assign n853 = n776 & ~n851;
  assign po12  = ~n852 & ~n853;
  assign n855 = ~n849 & ~n852;
  assign n856 = pi77  & n269;
  assign n857 = pi76  & n267;
  assign n858 = pi75  & n282;
  assign n859 = ~n837 & ~n839;
  assign n860 = ~pi76  & ~pi77 ;
  assign n861 = pi76  & pi77 ;
  assign n862 = ~n860 & ~n861;
  assign n863 = ~n859 & n862;
  assign n864 = n859 & ~n862;
  assign n865 = ~n863 & ~n864;
  assign n866 = n262 & n865;
  assign n867 = ~n856 & ~n857;
  assign n868 = ~n858 & n867;
  assign n869 = ~n866 & n868;
  assign n870 = pi2  & n869;
  assign n871 = ~pi2  & ~n869;
  assign n872 = ~n870 & ~n871;
  assign n873 = ~n826 & ~n829;
  assign n874 = ~n809 & ~n813;
  assign n875 = ~n793 & ~n796;
  assign n876 = pi66  & n750;
  assign n877 = pi67  & n651;
  assign n878 = pi68  & n646;
  assign n879 = n334 & n644;
  assign n880 = ~n877 & ~n878;
  assign n881 = ~n876 & n880;
  assign n882 = ~n879 & n881;
  assign n883 = pi11  & n882;
  assign n884 = ~pi11  & ~n882;
  assign n885 = ~n883 & ~n884;
  assign n886 = pi14  & n791;
  assign n887 = ~pi13  & ~pi14 ;
  assign n888 = pi13  & pi14 ;
  assign n889 = ~n887 & ~n888;
  assign n890 = n790 & n889;
  assign n891 = n265 & n890;
  assign n892 = n790 & ~n889;
  assign n893 = pi65  & n892;
  assign n894 = ~pi12  & ~pi13 ;
  assign n895 = pi12  & pi13 ;
  assign n896 = ~n894 & ~n895;
  assign n897 = ~n790 & n896;
  assign n898 = pi64  & n897;
  assign n899 = ~n891 & ~n893;
  assign n900 = ~n898 & n899;
  assign n901 = n886 & ~n900;
  assign n902 = ~n886 & n900;
  assign n903 = ~n901 & ~n902;
  assign n904 = n885 & ~n903;
  assign n905 = ~n885 & n903;
  assign n906 = ~n904 & ~n905;
  assign n907 = ~n875 & n906;
  assign n908 = n875 & ~n906;
  assign n909 = ~n907 & ~n908;
  assign n910 = pi69  & n528;
  assign n911 = pi70  & n490;
  assign n912 = pi71  & n485;
  assign n913 = n460 & n483;
  assign n914 = ~n911 & ~n912;
  assign n915 = ~n910 & n914;
  assign n916 = ~n913 & n915;
  assign n917 = pi8  & n916;
  assign n918 = ~pi8  & ~n916;
  assign n919 = ~n917 & ~n918;
  assign n920 = n909 & ~n919;
  assign n921 = ~n909 & n919;
  assign n922 = ~n920 & ~n921;
  assign n923 = n874 & ~n922;
  assign n924 = ~n874 & n922;
  assign n925 = ~n923 & ~n924;
  assign n926 = pi72  & n391;
  assign n927 = pi73  & n353;
  assign n928 = pi74  & n348;
  assign n929 = n346 & n689;
  assign n930 = ~n927 & ~n928;
  assign n931 = ~n926 & n930;
  assign n932 = ~n929 & n931;
  assign n933 = pi5  & n932;
  assign n934 = ~pi5  & ~n932;
  assign n935 = ~n933 & ~n934;
  assign n936 = n925 & ~n935;
  assign n937 = ~n925 & n935;
  assign n938 = ~n936 & ~n937;
  assign n939 = ~n873 & n938;
  assign n940 = n873 & ~n938;
  assign n941 = ~n939 & ~n940;
  assign n942 = ~n872 & n941;
  assign n943 = n872 & ~n941;
  assign n944 = ~n942 & ~n943;
  assign n945 = ~n855 & n944;
  assign n946 = n855 & ~n944;
  assign po13  = ~n945 & ~n946;
  assign n948 = ~n942 & ~n945;
  assign n949 = pi78  & n269;
  assign n950 = pi77  & n267;
  assign n951 = pi76  & n282;
  assign n952 = ~n861 & ~n863;
  assign n953 = ~pi77  & ~pi78 ;
  assign n954 = pi77  & pi78 ;
  assign n955 = ~n953 & ~n954;
  assign n956 = ~n952 & n955;
  assign n957 = n952 & ~n955;
  assign n958 = ~n956 & ~n957;
  assign n959 = n262 & n958;
  assign n960 = ~n949 & ~n950;
  assign n961 = ~n951 & n960;
  assign n962 = ~n959 & n961;
  assign n963 = pi2  & n962;
  assign n964 = ~pi2  & ~n962;
  assign n965 = ~n963 & ~n964;
  assign n966 = ~n936 & ~n939;
  assign n967 = pi73  & n391;
  assign n968 = pi74  & n353;
  assign n969 = pi75  & n348;
  assign n970 = n346 & n713;
  assign n971 = ~n968 & ~n969;
  assign n972 = ~n967 & n971;
  assign n973 = ~n970 & n972;
  assign n974 = pi5  & n973;
  assign n975 = ~pi5  & ~n973;
  assign n976 = ~n974 & ~n975;
  assign n977 = ~n920 & ~n924;
  assign n978 = pi70  & n528;
  assign n979 = pi71  & n490;
  assign n980 = pi72  & n485;
  assign n981 = n483 & n551;
  assign n982 = ~n979 & ~n980;
  assign n983 = ~n978 & n982;
  assign n984 = ~n981 & n983;
  assign n985 = pi8  & n984;
  assign n986 = ~pi8  & ~n984;
  assign n987 = ~n985 & ~n986;
  assign n988 = ~n905 & ~n907;
  assign n989 = pi67  & n750;
  assign n990 = pi68  & n651;
  assign n991 = pi69  & n646;
  assign n992 = n376 & n644;
  assign n993 = ~n990 & ~n991;
  assign n994 = ~n989 & n993;
  assign n995 = ~n992 & n994;
  assign n996 = pi11  & n995;
  assign n997 = ~pi11  & ~n995;
  assign n998 = ~n996 & ~n997;
  assign n999 = pi14  & ~n791;
  assign n1000 = n900 & n999;
  assign n1001 = pi14  & ~n1000;
  assign n1002 = ~n287 & n890;
  assign n1003 = pi65  & n897;
  assign n1004 = pi66  & n892;
  assign n1005 = ~n790 & n889;
  assign n1006 = ~n896 & n1005;
  assign n1007 = pi64  & n1006;
  assign n1008 = ~n1002 & ~n1003;
  assign n1009 = ~n1004 & n1008;
  assign n1010 = ~n1007 & n1009;
  assign n1011 = ~n1001 & n1010;
  assign n1012 = n1001 & ~n1010;
  assign n1013 = ~n1011 & ~n1012;
  assign n1014 = ~n998 & n1013;
  assign n1015 = n998 & ~n1013;
  assign n1016 = ~n1014 & ~n1015;
  assign n1017 = ~n988 & n1016;
  assign n1018 = n988 & ~n1016;
  assign n1019 = ~n1017 & ~n1018;
  assign n1020 = n987 & ~n1019;
  assign n1021 = ~n987 & n1019;
  assign n1022 = ~n1020 & ~n1021;
  assign n1023 = ~n977 & n1022;
  assign n1024 = n977 & ~n1022;
  assign n1025 = ~n1023 & ~n1024;
  assign n1026 = n976 & ~n1025;
  assign n1027 = ~n976 & n1025;
  assign n1028 = ~n1026 & ~n1027;
  assign n1029 = ~n966 & n1028;
  assign n1030 = n966 & ~n1028;
  assign n1031 = ~n1029 & ~n1030;
  assign n1032 = ~n965 & n1031;
  assign n1033 = n965 & ~n1031;
  assign n1034 = ~n1032 & ~n1033;
  assign n1035 = ~n948 & n1034;
  assign n1036 = n948 & ~n1034;
  assign po14  = ~n1035 & ~n1036;
  assign n1038 = ~n1032 & ~n1035;
  assign n1039 = pi79  & n269;
  assign n1040 = pi78  & n267;
  assign n1041 = pi77  & n282;
  assign n1042 = ~n954 & ~n956;
  assign n1043 = ~pi78  & ~pi79 ;
  assign n1044 = pi78  & pi79 ;
  assign n1045 = ~n1043 & ~n1044;
  assign n1046 = ~n1042 & n1045;
  assign n1047 = n1042 & ~n1045;
  assign n1048 = ~n1046 & ~n1047;
  assign n1049 = n262 & n1048;
  assign n1050 = ~n1039 & ~n1040;
  assign n1051 = ~n1041 & n1050;
  assign n1052 = ~n1049 & n1051;
  assign n1053 = pi2  & n1052;
  assign n1054 = ~pi2  & ~n1052;
  assign n1055 = ~n1053 & ~n1054;
  assign n1056 = ~n1027 & ~n1029;
  assign n1057 = pi74  & n391;
  assign n1058 = pi75  & n353;
  assign n1059 = pi76  & n348;
  assign n1060 = n346 & n841;
  assign n1061 = ~n1058 & ~n1059;
  assign n1062 = ~n1057 & n1061;
  assign n1063 = ~n1060 & n1062;
  assign n1064 = pi5  & n1063;
  assign n1065 = ~pi5  & ~n1063;
  assign n1066 = ~n1064 & ~n1065;
  assign n1067 = ~n1021 & ~n1023;
  assign n1068 = pi71  & n528;
  assign n1069 = pi72  & n490;
  assign n1070 = pi73  & n485;
  assign n1071 = n483 & n613;
  assign n1072 = ~n1069 & ~n1070;
  assign n1073 = ~n1068 & n1072;
  assign n1074 = ~n1071 & n1073;
  assign n1075 = pi8  & n1074;
  assign n1076 = ~pi8  & ~n1074;
  assign n1077 = ~n1075 & ~n1076;
  assign n1078 = ~n1014 & ~n1017;
  assign n1079 = pi65  & n1006;
  assign n1080 = pi66  & n897;
  assign n1081 = pi67  & n892;
  assign n1082 = n305 & n890;
  assign n1083 = ~n1080 & ~n1081;
  assign n1084 = ~n1079 & n1083;
  assign n1085 = ~n1082 & n1084;
  assign n1086 = pi14  & n1085;
  assign n1087 = ~pi14  & ~n1085;
  assign n1088 = ~n1086 & ~n1087;
  assign n1089 = ~pi14  & ~pi15 ;
  assign n1090 = pi14  & pi15 ;
  assign n1091 = ~n1089 & ~n1090;
  assign n1092 = pi64  & n1091;
  assign n1093 = n1000 & n1010;
  assign n1094 = n1092 & n1093;
  assign n1095 = ~n1092 & ~n1093;
  assign n1096 = ~n1094 & ~n1095;
  assign n1097 = ~n1088 & n1096;
  assign n1098 = n1088 & ~n1096;
  assign n1099 = ~n1097 & ~n1098;
  assign n1100 = pi68  & n750;
  assign n1101 = pi69  & n651;
  assign n1102 = pi70  & n646;
  assign n1103 = n415 & n644;
  assign n1104 = ~n1101 & ~n1102;
  assign n1105 = ~n1100 & n1104;
  assign n1106 = ~n1103 & n1105;
  assign n1107 = pi11  & n1106;
  assign n1108 = ~pi11  & ~n1106;
  assign n1109 = ~n1107 & ~n1108;
  assign n1110 = n1099 & ~n1109;
  assign n1111 = ~n1099 & n1109;
  assign n1112 = ~n1110 & ~n1111;
  assign n1113 = ~n1078 & n1112;
  assign n1114 = n1078 & ~n1112;
  assign n1115 = ~n1113 & ~n1114;
  assign n1116 = ~n1077 & n1115;
  assign n1117 = n1077 & ~n1115;
  assign n1118 = ~n1116 & ~n1117;
  assign n1119 = ~n1067 & n1118;
  assign n1120 = n1067 & ~n1118;
  assign n1121 = ~n1119 & ~n1120;
  assign n1122 = ~n1066 & n1121;
  assign n1123 = n1066 & ~n1121;
  assign n1124 = ~n1122 & ~n1123;
  assign n1125 = ~n1056 & n1124;
  assign n1126 = n1056 & ~n1124;
  assign n1127 = ~n1125 & ~n1126;
  assign n1128 = ~n1055 & n1127;
  assign n1129 = n1055 & ~n1127;
  assign n1130 = ~n1128 & ~n1129;
  assign n1131 = ~n1038 & n1130;
  assign n1132 = n1038 & ~n1130;
  assign po15  = ~n1131 & ~n1132;
  assign n1134 = ~n1128 & ~n1131;
  assign n1135 = pi80  & n269;
  assign n1136 = pi79  & n267;
  assign n1137 = pi78  & n282;
  assign n1138 = ~n1044 & ~n1046;
  assign n1139 = ~pi79  & ~pi80 ;
  assign n1140 = pi79  & pi80 ;
  assign n1141 = ~n1139 & ~n1140;
  assign n1142 = ~n1138 & n1141;
  assign n1143 = n1138 & ~n1141;
  assign n1144 = ~n1142 & ~n1143;
  assign n1145 = n262 & n1144;
  assign n1146 = ~n1135 & ~n1136;
  assign n1147 = ~n1137 & n1146;
  assign n1148 = ~n1145 & n1147;
  assign n1149 = pi2  & n1148;
  assign n1150 = ~pi2  & ~n1148;
  assign n1151 = ~n1149 & ~n1150;
  assign n1152 = ~n1122 & ~n1125;
  assign n1153 = pi75  & n391;
  assign n1154 = pi76  & n353;
  assign n1155 = pi77  & n348;
  assign n1156 = n346 & n865;
  assign n1157 = ~n1154 & ~n1155;
  assign n1158 = ~n1153 & n1157;
  assign n1159 = ~n1156 & n1158;
  assign n1160 = pi5  & n1159;
  assign n1161 = ~pi5  & ~n1159;
  assign n1162 = ~n1160 & ~n1161;
  assign n1163 = ~n1116 & ~n1119;
  assign n1164 = pi72  & n528;
  assign n1165 = pi73  & n490;
  assign n1166 = pi74  & n485;
  assign n1167 = n483 & n689;
  assign n1168 = ~n1165 & ~n1166;
  assign n1169 = ~n1164 & n1168;
  assign n1170 = ~n1167 & n1169;
  assign n1171 = pi8  & n1170;
  assign n1172 = ~pi8  & ~n1170;
  assign n1173 = ~n1171 & ~n1172;
  assign n1174 = ~n1110 & ~n1113;
  assign n1175 = pi69  & n750;
  assign n1176 = pi70  & n651;
  assign n1177 = pi71  & n646;
  assign n1178 = n460 & n644;
  assign n1179 = ~n1176 & ~n1177;
  assign n1180 = ~n1175 & n1179;
  assign n1181 = ~n1178 & n1180;
  assign n1182 = pi11  & n1181;
  assign n1183 = ~pi11  & ~n1181;
  assign n1184 = ~n1182 & ~n1183;
  assign n1185 = ~n1094 & ~n1097;
  assign n1186 = pi66  & n1006;
  assign n1187 = pi67  & n897;
  assign n1188 = pi68  & n892;
  assign n1189 = n334 & n890;
  assign n1190 = ~n1187 & ~n1188;
  assign n1191 = ~n1186 & n1190;
  assign n1192 = ~n1189 & n1191;
  assign n1193 = pi14  & n1192;
  assign n1194 = ~pi14  & ~n1192;
  assign n1195 = ~n1193 & ~n1194;
  assign n1196 = pi17  & n1092;
  assign n1197 = ~pi16  & ~pi17 ;
  assign n1198 = pi16  & pi17 ;
  assign n1199 = ~n1197 & ~n1198;
  assign n1200 = n1091 & n1199;
  assign n1201 = n265 & n1200;
  assign n1202 = n1091 & ~n1199;
  assign n1203 = pi65  & n1202;
  assign n1204 = ~pi15  & ~pi16 ;
  assign n1205 = pi15  & pi16 ;
  assign n1206 = ~n1204 & ~n1205;
  assign n1207 = ~n1091 & n1206;
  assign n1208 = pi64  & n1207;
  assign n1209 = ~n1201 & ~n1203;
  assign n1210 = ~n1208 & n1209;
  assign n1211 = n1196 & ~n1210;
  assign n1212 = ~n1196 & n1210;
  assign n1213 = ~n1211 & ~n1212;
  assign n1214 = n1195 & ~n1213;
  assign n1215 = ~n1195 & n1213;
  assign n1216 = ~n1214 & ~n1215;
  assign n1217 = ~n1185 & n1216;
  assign n1218 = n1185 & ~n1216;
  assign n1219 = ~n1217 & ~n1218;
  assign n1220 = n1184 & ~n1219;
  assign n1221 = ~n1184 & n1219;
  assign n1222 = ~n1220 & ~n1221;
  assign n1223 = ~n1174 & n1222;
  assign n1224 = n1174 & ~n1222;
  assign n1225 = ~n1223 & ~n1224;
  assign n1226 = n1173 & ~n1225;
  assign n1227 = ~n1173 & n1225;
  assign n1228 = ~n1226 & ~n1227;
  assign n1229 = ~n1163 & n1228;
  assign n1230 = n1163 & ~n1228;
  assign n1231 = ~n1229 & ~n1230;
  assign n1232 = n1162 & ~n1231;
  assign n1233 = ~n1162 & n1231;
  assign n1234 = ~n1232 & ~n1233;
  assign n1235 = ~n1152 & n1234;
  assign n1236 = n1152 & ~n1234;
  assign n1237 = ~n1235 & ~n1236;
  assign n1238 = ~n1151 & n1237;
  assign n1239 = n1151 & ~n1237;
  assign n1240 = ~n1238 & ~n1239;
  assign n1241 = ~n1134 & n1240;
  assign n1242 = n1134 & ~n1240;
  assign po16  = ~n1241 & ~n1242;
  assign n1244 = ~n1238 & ~n1241;
  assign n1245 = ~n1233 & ~n1235;
  assign n1246 = pi76  & n391;
  assign n1247 = pi77  & n353;
  assign n1248 = pi78  & n348;
  assign n1249 = n346 & n958;
  assign n1250 = ~n1247 & ~n1248;
  assign n1251 = ~n1246 & n1250;
  assign n1252 = ~n1249 & n1251;
  assign n1253 = pi5  & n1252;
  assign n1254 = ~pi5  & ~n1252;
  assign n1255 = ~n1253 & ~n1254;
  assign n1256 = ~n1227 & ~n1229;
  assign n1257 = pi73  & n528;
  assign n1258 = pi74  & n490;
  assign n1259 = pi75  & n485;
  assign n1260 = n483 & n713;
  assign n1261 = ~n1258 & ~n1259;
  assign n1262 = ~n1257 & n1261;
  assign n1263 = ~n1260 & n1262;
  assign n1264 = pi8  & n1263;
  assign n1265 = ~pi8  & ~n1263;
  assign n1266 = ~n1264 & ~n1265;
  assign n1267 = ~n1221 & ~n1223;
  assign n1268 = pi70  & n750;
  assign n1269 = pi71  & n651;
  assign n1270 = pi72  & n646;
  assign n1271 = n551 & n644;
  assign n1272 = ~n1269 & ~n1270;
  assign n1273 = ~n1268 & n1272;
  assign n1274 = ~n1271 & n1273;
  assign n1275 = pi11  & n1274;
  assign n1276 = ~pi11  & ~n1274;
  assign n1277 = ~n1275 & ~n1276;
  assign n1278 = ~n1215 & ~n1217;
  assign n1279 = pi67  & n1006;
  assign n1280 = pi68  & n897;
  assign n1281 = pi69  & n892;
  assign n1282 = n376 & n890;
  assign n1283 = ~n1280 & ~n1281;
  assign n1284 = ~n1279 & n1283;
  assign n1285 = ~n1282 & n1284;
  assign n1286 = pi14  & n1285;
  assign n1287 = ~pi14  & ~n1285;
  assign n1288 = ~n1286 & ~n1287;
  assign n1289 = pi17  & ~n1092;
  assign n1290 = n1210 & n1289;
  assign n1291 = pi17  & ~n1290;
  assign n1292 = ~n287 & n1200;
  assign n1293 = pi65  & n1207;
  assign n1294 = pi66  & n1202;
  assign n1295 = ~n1091 & n1199;
  assign n1296 = ~n1206 & n1295;
  assign n1297 = pi64  & n1296;
  assign n1298 = ~n1292 & ~n1293;
  assign n1299 = ~n1294 & n1298;
  assign n1300 = ~n1297 & n1299;
  assign n1301 = ~n1291 & n1300;
  assign n1302 = n1291 & ~n1300;
  assign n1303 = ~n1301 & ~n1302;
  assign n1304 = ~n1288 & n1303;
  assign n1305 = n1288 & ~n1303;
  assign n1306 = ~n1304 & ~n1305;
  assign n1307 = ~n1278 & n1306;
  assign n1308 = n1278 & ~n1306;
  assign n1309 = ~n1307 & ~n1308;
  assign n1310 = n1277 & ~n1309;
  assign n1311 = ~n1277 & n1309;
  assign n1312 = ~n1310 & ~n1311;
  assign n1313 = ~n1267 & n1312;
  assign n1314 = n1267 & ~n1312;
  assign n1315 = ~n1313 & ~n1314;
  assign n1316 = n1266 & ~n1315;
  assign n1317 = ~n1266 & n1315;
  assign n1318 = ~n1316 & ~n1317;
  assign n1319 = ~n1256 & n1318;
  assign n1320 = n1256 & ~n1318;
  assign n1321 = ~n1319 & ~n1320;
  assign n1322 = n1255 & ~n1321;
  assign n1323 = ~n1255 & n1321;
  assign n1324 = ~n1322 & ~n1323;
  assign n1325 = ~n1245 & n1324;
  assign n1326 = n1245 & ~n1324;
  assign n1327 = ~n1325 & ~n1326;
  assign n1328 = pi81  & n269;
  assign n1329 = pi80  & n267;
  assign n1330 = pi79  & n282;
  assign n1331 = ~n1140 & ~n1142;
  assign n1332 = ~pi80  & ~pi81 ;
  assign n1333 = pi80  & pi81 ;
  assign n1334 = ~n1332 & ~n1333;
  assign n1335 = ~n1331 & n1334;
  assign n1336 = n1331 & ~n1334;
  assign n1337 = ~n1335 & ~n1336;
  assign n1338 = n262 & n1337;
  assign n1339 = ~n1328 & ~n1329;
  assign n1340 = ~n1330 & n1339;
  assign n1341 = ~n1338 & n1340;
  assign n1342 = pi2  & n1341;
  assign n1343 = ~pi2  & ~n1341;
  assign n1344 = ~n1342 & ~n1343;
  assign n1345 = n1327 & ~n1344;
  assign n1346 = ~n1327 & n1344;
  assign n1347 = ~n1345 & ~n1346;
  assign n1348 = ~n1244 & n1347;
  assign n1349 = n1244 & ~n1347;
  assign po17  = ~n1348 & ~n1349;
  assign n1351 = ~n1345 & ~n1348;
  assign n1352 = ~n1323 & ~n1325;
  assign n1353 = pi77  & n391;
  assign n1354 = pi78  & n353;
  assign n1355 = pi79  & n348;
  assign n1356 = n346 & n1048;
  assign n1357 = ~n1354 & ~n1355;
  assign n1358 = ~n1353 & n1357;
  assign n1359 = ~n1356 & n1358;
  assign n1360 = pi5  & n1359;
  assign n1361 = ~pi5  & ~n1359;
  assign n1362 = ~n1360 & ~n1361;
  assign n1363 = ~n1317 & ~n1319;
  assign n1364 = pi74  & n528;
  assign n1365 = pi75  & n490;
  assign n1366 = pi76  & n485;
  assign n1367 = n483 & n841;
  assign n1368 = ~n1365 & ~n1366;
  assign n1369 = ~n1364 & n1368;
  assign n1370 = ~n1367 & n1369;
  assign n1371 = pi8  & n1370;
  assign n1372 = ~pi8  & ~n1370;
  assign n1373 = ~n1371 & ~n1372;
  assign n1374 = ~n1311 & ~n1313;
  assign n1375 = pi71  & n750;
  assign n1376 = pi72  & n651;
  assign n1377 = pi73  & n646;
  assign n1378 = n613 & n644;
  assign n1379 = ~n1376 & ~n1377;
  assign n1380 = ~n1375 & n1379;
  assign n1381 = ~n1378 & n1380;
  assign n1382 = pi11  & n1381;
  assign n1383 = ~pi11  & ~n1381;
  assign n1384 = ~n1382 & ~n1383;
  assign n1385 = ~n1304 & ~n1307;
  assign n1386 = pi65  & n1296;
  assign n1387 = pi66  & n1207;
  assign n1388 = pi67  & n1202;
  assign n1389 = n305 & n1200;
  assign n1390 = ~n1387 & ~n1388;
  assign n1391 = ~n1386 & n1390;
  assign n1392 = ~n1389 & n1391;
  assign n1393 = pi17  & n1392;
  assign n1394 = ~pi17  & ~n1392;
  assign n1395 = ~n1393 & ~n1394;
  assign n1396 = ~pi17  & ~pi18 ;
  assign n1397 = pi17  & pi18 ;
  assign n1398 = ~n1396 & ~n1397;
  assign n1399 = pi64  & n1398;
  assign n1400 = n1290 & n1300;
  assign n1401 = n1399 & n1400;
  assign n1402 = ~n1399 & ~n1400;
  assign n1403 = ~n1401 & ~n1402;
  assign n1404 = ~n1395 & n1403;
  assign n1405 = n1395 & ~n1403;
  assign n1406 = ~n1404 & ~n1405;
  assign n1407 = pi68  & n1006;
  assign n1408 = pi69  & n897;
  assign n1409 = pi70  & n892;
  assign n1410 = n415 & n890;
  assign n1411 = ~n1408 & ~n1409;
  assign n1412 = ~n1407 & n1411;
  assign n1413 = ~n1410 & n1412;
  assign n1414 = pi14  & n1413;
  assign n1415 = ~pi14  & ~n1413;
  assign n1416 = ~n1414 & ~n1415;
  assign n1417 = n1406 & ~n1416;
  assign n1418 = ~n1406 & n1416;
  assign n1419 = ~n1417 & ~n1418;
  assign n1420 = ~n1385 & n1419;
  assign n1421 = n1385 & ~n1419;
  assign n1422 = ~n1420 & ~n1421;
  assign n1423 = ~n1384 & n1422;
  assign n1424 = n1384 & ~n1422;
  assign n1425 = ~n1423 & ~n1424;
  assign n1426 = ~n1374 & n1425;
  assign n1427 = n1374 & ~n1425;
  assign n1428 = ~n1426 & ~n1427;
  assign n1429 = n1373 & ~n1428;
  assign n1430 = ~n1373 & n1428;
  assign n1431 = ~n1429 & ~n1430;
  assign n1432 = ~n1363 & n1431;
  assign n1433 = n1363 & ~n1431;
  assign n1434 = ~n1432 & ~n1433;
  assign n1435 = ~n1362 & n1434;
  assign n1436 = n1362 & ~n1434;
  assign n1437 = ~n1435 & ~n1436;
  assign n1438 = ~n1352 & n1437;
  assign n1439 = n1352 & ~n1437;
  assign n1440 = ~n1438 & ~n1439;
  assign n1441 = pi82  & n269;
  assign n1442 = pi81  & n267;
  assign n1443 = pi80  & n282;
  assign n1444 = ~n1333 & ~n1335;
  assign n1445 = ~pi81  & ~pi82 ;
  assign n1446 = pi81  & pi82 ;
  assign n1447 = ~n1445 & ~n1446;
  assign n1448 = ~n1444 & n1447;
  assign n1449 = n1444 & ~n1447;
  assign n1450 = ~n1448 & ~n1449;
  assign n1451 = n262 & n1450;
  assign n1452 = ~n1441 & ~n1442;
  assign n1453 = ~n1443 & n1452;
  assign n1454 = ~n1451 & n1453;
  assign n1455 = pi2  & n1454;
  assign n1456 = ~pi2  & ~n1454;
  assign n1457 = ~n1455 & ~n1456;
  assign n1458 = n1440 & ~n1457;
  assign n1459 = ~n1440 & n1457;
  assign n1460 = ~n1458 & ~n1459;
  assign n1461 = ~n1351 & n1460;
  assign n1462 = n1351 & ~n1460;
  assign po18  = ~n1461 & ~n1462;
  assign n1464 = ~n1458 & ~n1461;
  assign n1465 = ~n1435 & ~n1438;
  assign n1466 = ~n1423 & ~n1426;
  assign n1467 = ~n1417 & ~n1420;
  assign n1468 = pi69  & n1006;
  assign n1469 = pi70  & n897;
  assign n1470 = pi71  & n892;
  assign n1471 = n460 & n890;
  assign n1472 = ~n1469 & ~n1470;
  assign n1473 = ~n1468 & n1472;
  assign n1474 = ~n1471 & n1473;
  assign n1475 = pi14  & n1474;
  assign n1476 = ~pi14  & ~n1474;
  assign n1477 = ~n1475 & ~n1476;
  assign n1478 = ~n1401 & ~n1404;
  assign n1479 = pi66  & n1296;
  assign n1480 = pi67  & n1207;
  assign n1481 = pi68  & n1202;
  assign n1482 = n334 & n1200;
  assign n1483 = ~n1480 & ~n1481;
  assign n1484 = ~n1479 & n1483;
  assign n1485 = ~n1482 & n1484;
  assign n1486 = pi17  & n1485;
  assign n1487 = ~pi17  & ~n1485;
  assign n1488 = ~n1486 & ~n1487;
  assign n1489 = pi20  & n1399;
  assign n1490 = ~pi19  & ~pi20 ;
  assign n1491 = pi19  & pi20 ;
  assign n1492 = ~n1490 & ~n1491;
  assign n1493 = n1398 & n1492;
  assign n1494 = n265 & n1493;
  assign n1495 = n1398 & ~n1492;
  assign n1496 = pi65  & n1495;
  assign n1497 = ~pi18  & ~pi19 ;
  assign n1498 = pi18  & pi19 ;
  assign n1499 = ~n1497 & ~n1498;
  assign n1500 = ~n1398 & n1499;
  assign n1501 = pi64  & n1500;
  assign n1502 = ~n1494 & ~n1496;
  assign n1503 = ~n1501 & n1502;
  assign n1504 = n1489 & ~n1503;
  assign n1505 = ~n1489 & n1503;
  assign n1506 = ~n1504 & ~n1505;
  assign n1507 = ~n1488 & n1506;
  assign n1508 = n1488 & ~n1506;
  assign n1509 = ~n1507 & ~n1508;
  assign n1510 = ~n1478 & n1509;
  assign n1511 = n1478 & ~n1509;
  assign n1512 = ~n1510 & ~n1511;
  assign n1513 = ~n1477 & n1512;
  assign n1514 = n1477 & ~n1512;
  assign n1515 = ~n1513 & ~n1514;
  assign n1516 = ~n1467 & n1515;
  assign n1517 = n1467 & ~n1515;
  assign n1518 = ~n1516 & ~n1517;
  assign n1519 = pi72  & n750;
  assign n1520 = pi73  & n651;
  assign n1521 = pi74  & n646;
  assign n1522 = n644 & n689;
  assign n1523 = ~n1520 & ~n1521;
  assign n1524 = ~n1519 & n1523;
  assign n1525 = ~n1522 & n1524;
  assign n1526 = pi11  & n1525;
  assign n1527 = ~pi11  & ~n1525;
  assign n1528 = ~n1526 & ~n1527;
  assign n1529 = n1518 & ~n1528;
  assign n1530 = ~n1518 & n1528;
  assign n1531 = ~n1529 & ~n1530;
  assign n1532 = n1466 & ~n1531;
  assign n1533 = ~n1466 & n1531;
  assign n1534 = ~n1532 & ~n1533;
  assign n1535 = pi75  & n528;
  assign n1536 = pi76  & n490;
  assign n1537 = pi77  & n485;
  assign n1538 = n483 & n865;
  assign n1539 = ~n1536 & ~n1537;
  assign n1540 = ~n1535 & n1539;
  assign n1541 = ~n1538 & n1540;
  assign n1542 = pi8  & n1541;
  assign n1543 = ~pi8  & ~n1541;
  assign n1544 = ~n1542 & ~n1543;
  assign n1545 = ~n1534 & n1544;
  assign n1546 = n1534 & ~n1544;
  assign n1547 = ~n1545 & ~n1546;
  assign n1548 = ~n1430 & ~n1432;
  assign n1549 = n1547 & ~n1548;
  assign n1550 = ~n1547 & n1548;
  assign n1551 = ~n1549 & ~n1550;
  assign n1552 = pi78  & n391;
  assign n1553 = pi79  & n353;
  assign n1554 = pi80  & n348;
  assign n1555 = n346 & n1144;
  assign n1556 = ~n1553 & ~n1554;
  assign n1557 = ~n1552 & n1556;
  assign n1558 = ~n1555 & n1557;
  assign n1559 = pi5  & n1558;
  assign n1560 = ~pi5  & ~n1558;
  assign n1561 = ~n1559 & ~n1560;
  assign n1562 = n1551 & ~n1561;
  assign n1563 = ~n1551 & n1561;
  assign n1564 = ~n1562 & ~n1563;
  assign n1565 = n1465 & ~n1564;
  assign n1566 = ~n1465 & n1564;
  assign n1567 = ~n1565 & ~n1566;
  assign n1568 = pi83  & n269;
  assign n1569 = pi82  & n267;
  assign n1570 = pi81  & n282;
  assign n1571 = ~n1446 & ~n1448;
  assign n1572 = ~pi82  & ~pi83 ;
  assign n1573 = pi82  & pi83 ;
  assign n1574 = ~n1572 & ~n1573;
  assign n1575 = ~n1571 & n1574;
  assign n1576 = n1571 & ~n1574;
  assign n1577 = ~n1575 & ~n1576;
  assign n1578 = n262 & n1577;
  assign n1579 = ~n1568 & ~n1569;
  assign n1580 = ~n1570 & n1579;
  assign n1581 = ~n1578 & n1580;
  assign n1582 = pi2  & n1581;
  assign n1583 = ~pi2  & ~n1581;
  assign n1584 = ~n1582 & ~n1583;
  assign n1585 = n1567 & ~n1584;
  assign n1586 = ~n1567 & n1584;
  assign n1587 = ~n1585 & ~n1586;
  assign n1588 = ~n1464 & n1587;
  assign n1589 = n1464 & ~n1587;
  assign po19  = ~n1588 & ~n1589;
  assign n1591 = ~n1585 & ~n1588;
  assign n1592 = pi84  & n269;
  assign n1593 = pi83  & n267;
  assign n1594 = pi82  & n282;
  assign n1595 = ~n1573 & ~n1575;
  assign n1596 = ~pi83  & ~pi84 ;
  assign n1597 = pi83  & pi84 ;
  assign n1598 = ~n1596 & ~n1597;
  assign n1599 = ~n1595 & n1598;
  assign n1600 = n1595 & ~n1598;
  assign n1601 = ~n1599 & ~n1600;
  assign n1602 = n262 & n1601;
  assign n1603 = ~n1592 & ~n1593;
  assign n1604 = ~n1594 & n1603;
  assign n1605 = ~n1602 & n1604;
  assign n1606 = pi2  & n1605;
  assign n1607 = ~pi2  & ~n1605;
  assign n1608 = ~n1606 & ~n1607;
  assign n1609 = ~n1562 & ~n1566;
  assign n1610 = pi79  & n391;
  assign n1611 = pi80  & n353;
  assign n1612 = pi81  & n348;
  assign n1613 = n346 & n1337;
  assign n1614 = ~n1611 & ~n1612;
  assign n1615 = ~n1610 & n1614;
  assign n1616 = ~n1613 & n1615;
  assign n1617 = pi5  & n1616;
  assign n1618 = ~pi5  & ~n1616;
  assign n1619 = ~n1617 & ~n1618;
  assign n1620 = ~n1546 & ~n1549;
  assign n1621 = ~n1529 & ~n1533;
  assign n1622 = pi73  & n750;
  assign n1623 = pi74  & n651;
  assign n1624 = pi75  & n646;
  assign n1625 = n644 & n713;
  assign n1626 = ~n1623 & ~n1624;
  assign n1627 = ~n1622 & n1626;
  assign n1628 = ~n1625 & n1627;
  assign n1629 = pi11  & n1628;
  assign n1630 = ~pi11  & ~n1628;
  assign n1631 = ~n1629 & ~n1630;
  assign n1632 = ~n1513 & ~n1516;
  assign n1633 = pi70  & n1006;
  assign n1634 = pi71  & n897;
  assign n1635 = pi72  & n892;
  assign n1636 = n551 & n890;
  assign n1637 = ~n1634 & ~n1635;
  assign n1638 = ~n1633 & n1637;
  assign n1639 = ~n1636 & n1638;
  assign n1640 = pi14  & n1639;
  assign n1641 = ~pi14  & ~n1639;
  assign n1642 = ~n1640 & ~n1641;
  assign n1643 = ~n1507 & ~n1510;
  assign n1644 = pi67  & n1296;
  assign n1645 = pi68  & n1207;
  assign n1646 = pi69  & n1202;
  assign n1647 = n376 & n1200;
  assign n1648 = ~n1645 & ~n1646;
  assign n1649 = ~n1644 & n1648;
  assign n1650 = ~n1647 & n1649;
  assign n1651 = pi17  & n1650;
  assign n1652 = ~pi17  & ~n1650;
  assign n1653 = ~n1651 & ~n1652;
  assign n1654 = pi20  & ~n1399;
  assign n1655 = n1503 & n1654;
  assign n1656 = pi20  & ~n1655;
  assign n1657 = ~n287 & n1493;
  assign n1658 = pi65  & n1500;
  assign n1659 = pi66  & n1495;
  assign n1660 = ~n1398 & n1492;
  assign n1661 = ~n1499 & n1660;
  assign n1662 = pi64  & n1661;
  assign n1663 = ~n1657 & ~n1658;
  assign n1664 = ~n1659 & n1663;
  assign n1665 = ~n1662 & n1664;
  assign n1666 = ~n1656 & n1665;
  assign n1667 = n1656 & ~n1665;
  assign n1668 = ~n1666 & ~n1667;
  assign n1669 = ~n1653 & n1668;
  assign n1670 = n1653 & ~n1668;
  assign n1671 = ~n1669 & ~n1670;
  assign n1672 = ~n1643 & n1671;
  assign n1673 = n1643 & ~n1671;
  assign n1674 = ~n1672 & ~n1673;
  assign n1675 = n1642 & ~n1674;
  assign n1676 = ~n1642 & n1674;
  assign n1677 = ~n1675 & ~n1676;
  assign n1678 = ~n1632 & n1677;
  assign n1679 = n1632 & ~n1677;
  assign n1680 = ~n1678 & ~n1679;
  assign n1681 = n1631 & ~n1680;
  assign n1682 = ~n1631 & n1680;
  assign n1683 = ~n1681 & ~n1682;
  assign n1684 = ~n1621 & n1683;
  assign n1685 = n1621 & ~n1683;
  assign n1686 = ~n1684 & ~n1685;
  assign n1687 = pi76  & n528;
  assign n1688 = pi77  & n490;
  assign n1689 = pi78  & n485;
  assign n1690 = n483 & n958;
  assign n1691 = ~n1688 & ~n1689;
  assign n1692 = ~n1687 & n1691;
  assign n1693 = ~n1690 & n1692;
  assign n1694 = pi8  & n1693;
  assign n1695 = ~pi8  & ~n1693;
  assign n1696 = ~n1694 & ~n1695;
  assign n1697 = n1686 & ~n1696;
  assign n1698 = ~n1686 & n1696;
  assign n1699 = ~n1697 & ~n1698;
  assign n1700 = ~n1620 & n1699;
  assign n1701 = n1620 & ~n1699;
  assign n1702 = ~n1700 & ~n1701;
  assign n1703 = ~n1619 & n1702;
  assign n1704 = n1619 & ~n1702;
  assign n1705 = ~n1703 & ~n1704;
  assign n1706 = ~n1609 & n1705;
  assign n1707 = n1609 & ~n1705;
  assign n1708 = ~n1706 & ~n1707;
  assign n1709 = ~n1608 & n1708;
  assign n1710 = n1608 & ~n1708;
  assign n1711 = ~n1709 & ~n1710;
  assign n1712 = ~n1591 & n1711;
  assign n1713 = n1591 & ~n1711;
  assign po20  = ~n1712 & ~n1713;
  assign n1715 = ~n1709 & ~n1712;
  assign n1716 = ~n1703 & ~n1706;
  assign n1717 = ~n1697 & ~n1700;
  assign n1718 = pi77  & n528;
  assign n1719 = pi78  & n490;
  assign n1720 = pi79  & n485;
  assign n1721 = n483 & n1048;
  assign n1722 = ~n1719 & ~n1720;
  assign n1723 = ~n1718 & n1722;
  assign n1724 = ~n1721 & n1723;
  assign n1725 = pi8  & n1724;
  assign n1726 = ~pi8  & ~n1724;
  assign n1727 = ~n1725 & ~n1726;
  assign n1728 = ~n1682 & ~n1684;
  assign n1729 = pi74  & n750;
  assign n1730 = pi75  & n651;
  assign n1731 = pi76  & n646;
  assign n1732 = n644 & n841;
  assign n1733 = ~n1730 & ~n1731;
  assign n1734 = ~n1729 & n1733;
  assign n1735 = ~n1732 & n1734;
  assign n1736 = pi11  & n1735;
  assign n1737 = ~pi11  & ~n1735;
  assign n1738 = ~n1736 & ~n1737;
  assign n1739 = ~n1676 & ~n1678;
  assign n1740 = pi71  & n1006;
  assign n1741 = pi72  & n897;
  assign n1742 = pi73  & n892;
  assign n1743 = n613 & n890;
  assign n1744 = ~n1741 & ~n1742;
  assign n1745 = ~n1740 & n1744;
  assign n1746 = ~n1743 & n1745;
  assign n1747 = pi14  & n1746;
  assign n1748 = ~pi14  & ~n1746;
  assign n1749 = ~n1747 & ~n1748;
  assign n1750 = ~n1669 & ~n1672;
  assign n1751 = pi65  & n1661;
  assign n1752 = pi66  & n1500;
  assign n1753 = pi67  & n1495;
  assign n1754 = n305 & n1493;
  assign n1755 = ~n1752 & ~n1753;
  assign n1756 = ~n1751 & n1755;
  assign n1757 = ~n1754 & n1756;
  assign n1758 = pi20  & n1757;
  assign n1759 = ~pi20  & ~n1757;
  assign n1760 = ~n1758 & ~n1759;
  assign n1761 = ~pi20  & ~pi21 ;
  assign n1762 = pi20  & pi21 ;
  assign n1763 = ~n1761 & ~n1762;
  assign n1764 = pi64  & n1763;
  assign n1765 = n1655 & n1665;
  assign n1766 = n1764 & n1765;
  assign n1767 = ~n1764 & ~n1765;
  assign n1768 = ~n1766 & ~n1767;
  assign n1769 = ~n1760 & n1768;
  assign n1770 = n1760 & ~n1768;
  assign n1771 = ~n1769 & ~n1770;
  assign n1772 = pi68  & n1296;
  assign n1773 = pi69  & n1207;
  assign n1774 = pi70  & n1202;
  assign n1775 = n415 & n1200;
  assign n1776 = ~n1773 & ~n1774;
  assign n1777 = ~n1772 & n1776;
  assign n1778 = ~n1775 & n1777;
  assign n1779 = pi17  & n1778;
  assign n1780 = ~pi17  & ~n1778;
  assign n1781 = ~n1779 & ~n1780;
  assign n1782 = n1771 & ~n1781;
  assign n1783 = ~n1771 & n1781;
  assign n1784 = ~n1782 & ~n1783;
  assign n1785 = ~n1750 & n1784;
  assign n1786 = n1750 & ~n1784;
  assign n1787 = ~n1785 & ~n1786;
  assign n1788 = ~n1749 & n1787;
  assign n1789 = n1749 & ~n1787;
  assign n1790 = ~n1788 & ~n1789;
  assign n1791 = ~n1739 & n1790;
  assign n1792 = n1739 & ~n1790;
  assign n1793 = ~n1791 & ~n1792;
  assign n1794 = n1738 & ~n1793;
  assign n1795 = ~n1738 & n1793;
  assign n1796 = ~n1794 & ~n1795;
  assign n1797 = ~n1728 & n1796;
  assign n1798 = n1728 & ~n1796;
  assign n1799 = ~n1797 & ~n1798;
  assign n1800 = ~n1727 & n1799;
  assign n1801 = n1727 & ~n1799;
  assign n1802 = ~n1800 & ~n1801;
  assign n1803 = ~n1717 & n1802;
  assign n1804 = n1717 & ~n1802;
  assign n1805 = ~n1803 & ~n1804;
  assign n1806 = pi80  & n391;
  assign n1807 = pi81  & n353;
  assign n1808 = pi82  & n348;
  assign n1809 = n346 & n1450;
  assign n1810 = ~n1807 & ~n1808;
  assign n1811 = ~n1806 & n1810;
  assign n1812 = ~n1809 & n1811;
  assign n1813 = pi5  & n1812;
  assign n1814 = ~pi5  & ~n1812;
  assign n1815 = ~n1813 & ~n1814;
  assign n1816 = n1805 & ~n1815;
  assign n1817 = ~n1805 & n1815;
  assign n1818 = ~n1816 & ~n1817;
  assign n1819 = n1716 & ~n1818;
  assign n1820 = ~n1716 & n1818;
  assign n1821 = ~n1819 & ~n1820;
  assign n1822 = pi85  & n269;
  assign n1823 = pi84  & n267;
  assign n1824 = pi83  & n282;
  assign n1825 = ~n1597 & ~n1599;
  assign n1826 = ~pi84  & ~pi85 ;
  assign n1827 = pi84  & pi85 ;
  assign n1828 = ~n1826 & ~n1827;
  assign n1829 = ~n1825 & n1828;
  assign n1830 = n1825 & ~n1828;
  assign n1831 = ~n1829 & ~n1830;
  assign n1832 = n262 & n1831;
  assign n1833 = ~n1822 & ~n1823;
  assign n1834 = ~n1824 & n1833;
  assign n1835 = ~n1832 & n1834;
  assign n1836 = pi2  & n1835;
  assign n1837 = ~pi2  & ~n1835;
  assign n1838 = ~n1836 & ~n1837;
  assign n1839 = n1821 & ~n1838;
  assign n1840 = ~n1821 & n1838;
  assign n1841 = ~n1839 & ~n1840;
  assign n1842 = ~n1715 & n1841;
  assign n1843 = n1715 & ~n1841;
  assign po21  = ~n1842 & ~n1843;
  assign n1845 = ~n1839 & ~n1842;
  assign n1846 = ~n1816 & ~n1820;
  assign n1847 = ~n1800 & ~n1803;
  assign n1848 = pi78  & n528;
  assign n1849 = pi79  & n490;
  assign n1850 = pi80  & n485;
  assign n1851 = n483 & n1144;
  assign n1852 = ~n1849 & ~n1850;
  assign n1853 = ~n1848 & n1852;
  assign n1854 = ~n1851 & n1853;
  assign n1855 = pi8  & n1854;
  assign n1856 = ~pi8  & ~n1854;
  assign n1857 = ~n1855 & ~n1856;
  assign n1858 = ~n1795 & ~n1797;
  assign n1859 = ~n1788 & ~n1791;
  assign n1860 = ~n1782 & ~n1785;
  assign n1861 = pi69  & n1296;
  assign n1862 = pi70  & n1207;
  assign n1863 = pi71  & n1202;
  assign n1864 = n460 & n1200;
  assign n1865 = ~n1862 & ~n1863;
  assign n1866 = ~n1861 & n1865;
  assign n1867 = ~n1864 & n1866;
  assign n1868 = pi17  & n1867;
  assign n1869 = ~pi17  & ~n1867;
  assign n1870 = ~n1868 & ~n1869;
  assign n1871 = ~n1766 & ~n1769;
  assign n1872 = pi66  & n1661;
  assign n1873 = pi67  & n1500;
  assign n1874 = pi68  & n1495;
  assign n1875 = n334 & n1493;
  assign n1876 = ~n1873 & ~n1874;
  assign n1877 = ~n1872 & n1876;
  assign n1878 = ~n1875 & n1877;
  assign n1879 = pi20  & n1878;
  assign n1880 = ~pi20  & ~n1878;
  assign n1881 = ~n1879 & ~n1880;
  assign n1882 = pi23  & n1764;
  assign n1883 = ~pi22  & ~pi23 ;
  assign n1884 = pi22  & pi23 ;
  assign n1885 = ~n1883 & ~n1884;
  assign n1886 = n1763 & n1885;
  assign n1887 = n265 & n1886;
  assign n1888 = n1763 & ~n1885;
  assign n1889 = pi65  & n1888;
  assign n1890 = ~pi21  & ~pi22 ;
  assign n1891 = pi21  & pi22 ;
  assign n1892 = ~n1890 & ~n1891;
  assign n1893 = ~n1763 & n1892;
  assign n1894 = pi64  & n1893;
  assign n1895 = ~n1887 & ~n1889;
  assign n1896 = ~n1894 & n1895;
  assign n1897 = n1882 & ~n1896;
  assign n1898 = ~n1882 & n1896;
  assign n1899 = ~n1897 & ~n1898;
  assign n1900 = ~n1881 & n1899;
  assign n1901 = n1881 & ~n1899;
  assign n1902 = ~n1900 & ~n1901;
  assign n1903 = ~n1871 & n1902;
  assign n1904 = n1871 & ~n1902;
  assign n1905 = ~n1903 & ~n1904;
  assign n1906 = ~n1870 & n1905;
  assign n1907 = n1870 & ~n1905;
  assign n1908 = ~n1906 & ~n1907;
  assign n1909 = ~n1860 & n1908;
  assign n1910 = n1860 & ~n1908;
  assign n1911 = ~n1909 & ~n1910;
  assign n1912 = pi72  & n1006;
  assign n1913 = pi73  & n897;
  assign n1914 = pi74  & n892;
  assign n1915 = n689 & n890;
  assign n1916 = ~n1913 & ~n1914;
  assign n1917 = ~n1912 & n1916;
  assign n1918 = ~n1915 & n1917;
  assign n1919 = pi14  & n1918;
  assign n1920 = ~pi14  & ~n1918;
  assign n1921 = ~n1919 & ~n1920;
  assign n1922 = n1911 & ~n1921;
  assign n1923 = ~n1911 & n1921;
  assign n1924 = ~n1922 & ~n1923;
  assign n1925 = n1859 & ~n1924;
  assign n1926 = ~n1859 & n1924;
  assign n1927 = ~n1925 & ~n1926;
  assign n1928 = pi75  & n750;
  assign n1929 = pi76  & n651;
  assign n1930 = pi77  & n646;
  assign n1931 = n644 & n865;
  assign n1932 = ~n1929 & ~n1930;
  assign n1933 = ~n1928 & n1932;
  assign n1934 = ~n1931 & n1933;
  assign n1935 = pi11  & n1934;
  assign n1936 = ~pi11  & ~n1934;
  assign n1937 = ~n1935 & ~n1936;
  assign n1938 = ~n1927 & n1937;
  assign n1939 = n1927 & ~n1937;
  assign n1940 = ~n1938 & ~n1939;
  assign n1941 = ~n1858 & n1940;
  assign n1942 = n1858 & ~n1940;
  assign n1943 = ~n1941 & ~n1942;
  assign n1944 = ~n1857 & n1943;
  assign n1945 = n1857 & ~n1943;
  assign n1946 = ~n1944 & ~n1945;
  assign n1947 = ~n1847 & n1946;
  assign n1948 = n1847 & ~n1946;
  assign n1949 = ~n1947 & ~n1948;
  assign n1950 = pi81  & n391;
  assign n1951 = pi82  & n353;
  assign n1952 = pi83  & n348;
  assign n1953 = n346 & n1577;
  assign n1954 = ~n1951 & ~n1952;
  assign n1955 = ~n1950 & n1954;
  assign n1956 = ~n1953 & n1955;
  assign n1957 = pi5  & n1956;
  assign n1958 = ~pi5  & ~n1956;
  assign n1959 = ~n1957 & ~n1958;
  assign n1960 = n1949 & ~n1959;
  assign n1961 = ~n1949 & n1959;
  assign n1962 = ~n1960 & ~n1961;
  assign n1963 = n1846 & ~n1962;
  assign n1964 = ~n1846 & n1962;
  assign n1965 = ~n1963 & ~n1964;
  assign n1966 = pi86  & n269;
  assign n1967 = pi85  & n267;
  assign n1968 = pi84  & n282;
  assign n1969 = ~n1827 & ~n1829;
  assign n1970 = ~pi85  & ~pi86 ;
  assign n1971 = pi85  & pi86 ;
  assign n1972 = ~n1970 & ~n1971;
  assign n1973 = ~n1969 & n1972;
  assign n1974 = n1969 & ~n1972;
  assign n1975 = ~n1973 & ~n1974;
  assign n1976 = n262 & n1975;
  assign n1977 = ~n1966 & ~n1967;
  assign n1978 = ~n1968 & n1977;
  assign n1979 = ~n1976 & n1978;
  assign n1980 = pi2  & n1979;
  assign n1981 = ~pi2  & ~n1979;
  assign n1982 = ~n1980 & ~n1981;
  assign n1983 = ~n1965 & n1982;
  assign n1984 = n1965 & ~n1982;
  assign n1985 = ~n1983 & ~n1984;
  assign n1986 = ~n1845 & n1985;
  assign n1987 = n1845 & ~n1985;
  assign po22  = ~n1986 & ~n1987;
  assign n1989 = ~n1984 & ~n1986;
  assign n1990 = ~n1960 & ~n1964;
  assign n1991 = pi82  & n391;
  assign n1992 = pi83  & n353;
  assign n1993 = pi84  & n348;
  assign n1994 = n346 & n1601;
  assign n1995 = ~n1992 & ~n1993;
  assign n1996 = ~n1991 & n1995;
  assign n1997 = ~n1994 & n1996;
  assign n1998 = pi5  & n1997;
  assign n1999 = ~pi5  & ~n1997;
  assign n2000 = ~n1998 & ~n1999;
  assign n2001 = ~n1944 & ~n1947;
  assign n2002 = pi79  & n528;
  assign n2003 = pi80  & n490;
  assign n2004 = pi81  & n485;
  assign n2005 = n483 & n1337;
  assign n2006 = ~n2003 & ~n2004;
  assign n2007 = ~n2002 & n2006;
  assign n2008 = ~n2005 & n2007;
  assign n2009 = pi8  & n2008;
  assign n2010 = ~pi8  & ~n2008;
  assign n2011 = ~n2009 & ~n2010;
  assign n2012 = ~n1939 & ~n1941;
  assign n2013 = ~n1922 & ~n1926;
  assign n2014 = pi73  & n1006;
  assign n2015 = pi74  & n897;
  assign n2016 = pi75  & n892;
  assign n2017 = n713 & n890;
  assign n2018 = ~n2015 & ~n2016;
  assign n2019 = ~n2014 & n2018;
  assign n2020 = ~n2017 & n2019;
  assign n2021 = pi14  & n2020;
  assign n2022 = ~pi14  & ~n2020;
  assign n2023 = ~n2021 & ~n2022;
  assign n2024 = ~n1906 & ~n1909;
  assign n2025 = pi70  & n1296;
  assign n2026 = pi71  & n1207;
  assign n2027 = pi72  & n1202;
  assign n2028 = n551 & n1200;
  assign n2029 = ~n2026 & ~n2027;
  assign n2030 = ~n2025 & n2029;
  assign n2031 = ~n2028 & n2030;
  assign n2032 = pi17  & n2031;
  assign n2033 = ~pi17  & ~n2031;
  assign n2034 = ~n2032 & ~n2033;
  assign n2035 = ~n1900 & ~n1903;
  assign n2036 = pi67  & n1661;
  assign n2037 = pi68  & n1500;
  assign n2038 = pi69  & n1495;
  assign n2039 = n376 & n1493;
  assign n2040 = ~n2037 & ~n2038;
  assign n2041 = ~n2036 & n2040;
  assign n2042 = ~n2039 & n2041;
  assign n2043 = pi20  & n2042;
  assign n2044 = ~pi20  & ~n2042;
  assign n2045 = ~n2043 & ~n2044;
  assign n2046 = pi23  & ~n1764;
  assign n2047 = n1896 & n2046;
  assign n2048 = pi23  & ~n2047;
  assign n2049 = ~n287 & n1886;
  assign n2050 = pi65  & n1893;
  assign n2051 = pi66  & n1888;
  assign n2052 = ~n1763 & n1885;
  assign n2053 = ~n1892 & n2052;
  assign n2054 = pi64  & n2053;
  assign n2055 = ~n2049 & ~n2050;
  assign n2056 = ~n2051 & n2055;
  assign n2057 = ~n2054 & n2056;
  assign n2058 = ~n2048 & n2057;
  assign n2059 = n2048 & ~n2057;
  assign n2060 = ~n2058 & ~n2059;
  assign n2061 = ~n2045 & n2060;
  assign n2062 = n2045 & ~n2060;
  assign n2063 = ~n2061 & ~n2062;
  assign n2064 = ~n2035 & n2063;
  assign n2065 = n2035 & ~n2063;
  assign n2066 = ~n2064 & ~n2065;
  assign n2067 = n2034 & ~n2066;
  assign n2068 = ~n2034 & n2066;
  assign n2069 = ~n2067 & ~n2068;
  assign n2070 = ~n2024 & n2069;
  assign n2071 = n2024 & ~n2069;
  assign n2072 = ~n2070 & ~n2071;
  assign n2073 = n2023 & ~n2072;
  assign n2074 = ~n2023 & n2072;
  assign n2075 = ~n2073 & ~n2074;
  assign n2076 = ~n2013 & n2075;
  assign n2077 = n2013 & ~n2075;
  assign n2078 = ~n2076 & ~n2077;
  assign n2079 = pi76  & n750;
  assign n2080 = pi77  & n651;
  assign n2081 = pi78  & n646;
  assign n2082 = n644 & n958;
  assign n2083 = ~n2080 & ~n2081;
  assign n2084 = ~n2079 & n2083;
  assign n2085 = ~n2082 & n2084;
  assign n2086 = pi11  & n2085;
  assign n2087 = ~pi11  & ~n2085;
  assign n2088 = ~n2086 & ~n2087;
  assign n2089 = n2078 & ~n2088;
  assign n2090 = ~n2078 & n2088;
  assign n2091 = ~n2089 & ~n2090;
  assign n2092 = ~n2012 & n2091;
  assign n2093 = n2012 & ~n2091;
  assign n2094 = ~n2092 & ~n2093;
  assign n2095 = ~n2011 & n2094;
  assign n2096 = n2011 & ~n2094;
  assign n2097 = ~n2095 & ~n2096;
  assign n2098 = ~n2001 & n2097;
  assign n2099 = n2001 & ~n2097;
  assign n2100 = ~n2098 & ~n2099;
  assign n2101 = ~n2000 & n2100;
  assign n2102 = n2000 & ~n2100;
  assign n2103 = ~n2101 & ~n2102;
  assign n2104 = n1990 & ~n2103;
  assign n2105 = ~n1990 & n2103;
  assign n2106 = ~n2104 & ~n2105;
  assign n2107 = pi87  & n269;
  assign n2108 = pi86  & n267;
  assign n2109 = pi85  & n282;
  assign n2110 = ~n1971 & ~n1973;
  assign n2111 = ~pi86  & ~pi87 ;
  assign n2112 = pi86  & pi87 ;
  assign n2113 = ~n2111 & ~n2112;
  assign n2114 = ~n2110 & n2113;
  assign n2115 = n2110 & ~n2113;
  assign n2116 = ~n2114 & ~n2115;
  assign n2117 = n262 & n2116;
  assign n2118 = ~n2107 & ~n2108;
  assign n2119 = ~n2109 & n2118;
  assign n2120 = ~n2117 & n2119;
  assign n2121 = pi2  & n2120;
  assign n2122 = ~pi2  & ~n2120;
  assign n2123 = ~n2121 & ~n2122;
  assign n2124 = n2106 & ~n2123;
  assign n2125 = ~n2106 & n2123;
  assign n2126 = ~n2124 & ~n2125;
  assign n2127 = ~n1989 & n2126;
  assign n2128 = n1989 & ~n2126;
  assign po23  = ~n2127 & ~n2128;
  assign n2130 = ~n2124 & ~n2127;
  assign n2131 = pi88  & n269;
  assign n2132 = pi87  & n267;
  assign n2133 = pi86  & n282;
  assign n2134 = ~n2112 & ~n2114;
  assign n2135 = ~pi87  & ~pi88 ;
  assign n2136 = pi87  & pi88 ;
  assign n2137 = ~n2135 & ~n2136;
  assign n2138 = ~n2134 & n2137;
  assign n2139 = n2134 & ~n2137;
  assign n2140 = ~n2138 & ~n2139;
  assign n2141 = n262 & n2140;
  assign n2142 = ~n2131 & ~n2132;
  assign n2143 = ~n2133 & n2142;
  assign n2144 = ~n2141 & n2143;
  assign n2145 = pi2  & n2144;
  assign n2146 = ~pi2  & ~n2144;
  assign n2147 = ~n2145 & ~n2146;
  assign n2148 = ~n2101 & ~n2105;
  assign n2149 = pi83  & n391;
  assign n2150 = pi84  & n353;
  assign n2151 = pi85  & n348;
  assign n2152 = n346 & n1831;
  assign n2153 = ~n2150 & ~n2151;
  assign n2154 = ~n2149 & n2153;
  assign n2155 = ~n2152 & n2154;
  assign n2156 = pi5  & n2155;
  assign n2157 = ~pi5  & ~n2155;
  assign n2158 = ~n2156 & ~n2157;
  assign n2159 = ~n2095 & ~n2098;
  assign n2160 = ~n2089 & ~n2092;
  assign n2161 = ~n2074 & ~n2076;
  assign n2162 = pi74  & n1006;
  assign n2163 = pi75  & n897;
  assign n2164 = pi76  & n892;
  assign n2165 = n841 & n890;
  assign n2166 = ~n2163 & ~n2164;
  assign n2167 = ~n2162 & n2166;
  assign n2168 = ~n2165 & n2167;
  assign n2169 = pi14  & n2168;
  assign n2170 = ~pi14  & ~n2168;
  assign n2171 = ~n2169 & ~n2170;
  assign n2172 = ~n2068 & ~n2070;
  assign n2173 = pi71  & n1296;
  assign n2174 = pi72  & n1207;
  assign n2175 = pi73  & n1202;
  assign n2176 = n613 & n1200;
  assign n2177 = ~n2174 & ~n2175;
  assign n2178 = ~n2173 & n2177;
  assign n2179 = ~n2176 & n2178;
  assign n2180 = pi17  & n2179;
  assign n2181 = ~pi17  & ~n2179;
  assign n2182 = ~n2180 & ~n2181;
  assign n2183 = ~n2061 & ~n2064;
  assign n2184 = pi65  & n2053;
  assign n2185 = pi66  & n1893;
  assign n2186 = pi67  & n1888;
  assign n2187 = n305 & n1886;
  assign n2188 = ~n2185 & ~n2186;
  assign n2189 = ~n2184 & n2188;
  assign n2190 = ~n2187 & n2189;
  assign n2191 = pi23  & n2190;
  assign n2192 = ~pi23  & ~n2190;
  assign n2193 = ~n2191 & ~n2192;
  assign n2194 = ~pi23  & ~pi24 ;
  assign n2195 = pi23  & pi24 ;
  assign n2196 = ~n2194 & ~n2195;
  assign n2197 = pi64  & n2196;
  assign n2198 = n2047 & n2057;
  assign n2199 = n2197 & n2198;
  assign n2200 = ~n2197 & ~n2198;
  assign n2201 = ~n2199 & ~n2200;
  assign n2202 = ~n2193 & n2201;
  assign n2203 = n2193 & ~n2201;
  assign n2204 = ~n2202 & ~n2203;
  assign n2205 = pi68  & n1661;
  assign n2206 = pi69  & n1500;
  assign n2207 = pi70  & n1495;
  assign n2208 = n415 & n1493;
  assign n2209 = ~n2206 & ~n2207;
  assign n2210 = ~n2205 & n2209;
  assign n2211 = ~n2208 & n2210;
  assign n2212 = pi20  & n2211;
  assign n2213 = ~pi20  & ~n2211;
  assign n2214 = ~n2212 & ~n2213;
  assign n2215 = n2204 & ~n2214;
  assign n2216 = ~n2204 & n2214;
  assign n2217 = ~n2215 & ~n2216;
  assign n2218 = ~n2183 & n2217;
  assign n2219 = n2183 & ~n2217;
  assign n2220 = ~n2218 & ~n2219;
  assign n2221 = ~n2182 & n2220;
  assign n2222 = n2182 & ~n2220;
  assign n2223 = ~n2221 & ~n2222;
  assign n2224 = ~n2172 & n2223;
  assign n2225 = n2172 & ~n2223;
  assign n2226 = ~n2224 & ~n2225;
  assign n2227 = n2171 & ~n2226;
  assign n2228 = ~n2171 & n2226;
  assign n2229 = ~n2227 & ~n2228;
  assign n2230 = ~n2161 & n2229;
  assign n2231 = n2161 & ~n2229;
  assign n2232 = ~n2230 & ~n2231;
  assign n2233 = pi77  & n750;
  assign n2234 = pi78  & n651;
  assign n2235 = pi79  & n646;
  assign n2236 = n644 & n1048;
  assign n2237 = ~n2234 & ~n2235;
  assign n2238 = ~n2233 & n2237;
  assign n2239 = ~n2236 & n2238;
  assign n2240 = pi11  & n2239;
  assign n2241 = ~pi11  & ~n2239;
  assign n2242 = ~n2240 & ~n2241;
  assign n2243 = n2232 & ~n2242;
  assign n2244 = ~n2232 & n2242;
  assign n2245 = ~n2243 & ~n2244;
  assign n2246 = n2160 & ~n2245;
  assign n2247 = ~n2160 & n2245;
  assign n2248 = ~n2246 & ~n2247;
  assign n2249 = pi80  & n528;
  assign n2250 = pi81  & n490;
  assign n2251 = pi82  & n485;
  assign n2252 = n483 & n1450;
  assign n2253 = ~n2250 & ~n2251;
  assign n2254 = ~n2249 & n2253;
  assign n2255 = ~n2252 & n2254;
  assign n2256 = pi8  & n2255;
  assign n2257 = ~pi8  & ~n2255;
  assign n2258 = ~n2256 & ~n2257;
  assign n2259 = ~n2248 & n2258;
  assign n2260 = n2248 & ~n2258;
  assign n2261 = ~n2259 & ~n2260;
  assign n2262 = ~n2159 & n2261;
  assign n2263 = n2159 & ~n2261;
  assign n2264 = ~n2262 & ~n2263;
  assign n2265 = ~n2158 & n2264;
  assign n2266 = n2158 & ~n2264;
  assign n2267 = ~n2265 & ~n2266;
  assign n2268 = ~n2148 & n2267;
  assign n2269 = n2148 & ~n2267;
  assign n2270 = ~n2268 & ~n2269;
  assign n2271 = ~n2147 & n2270;
  assign n2272 = n2147 & ~n2270;
  assign n2273 = ~n2271 & ~n2272;
  assign n2274 = ~n2130 & n2273;
  assign n2275 = n2130 & ~n2273;
  assign po24  = ~n2274 & ~n2275;
  assign n2277 = ~n2271 & ~n2274;
  assign n2278 = pi89  & n269;
  assign n2279 = pi88  & n267;
  assign n2280 = pi87  & n282;
  assign n2281 = ~n2136 & ~n2138;
  assign n2282 = ~pi88  & ~pi89 ;
  assign n2283 = pi88  & pi89 ;
  assign n2284 = ~n2282 & ~n2283;
  assign n2285 = ~n2281 & n2284;
  assign n2286 = n2281 & ~n2284;
  assign n2287 = ~n2285 & ~n2286;
  assign n2288 = n262 & n2287;
  assign n2289 = ~n2278 & ~n2279;
  assign n2290 = ~n2280 & n2289;
  assign n2291 = ~n2288 & n2290;
  assign n2292 = pi2  & n2291;
  assign n2293 = ~pi2  & ~n2291;
  assign n2294 = ~n2292 & ~n2293;
  assign n2295 = ~n2265 & ~n2268;
  assign n2296 = pi84  & n391;
  assign n2297 = pi85  & n353;
  assign n2298 = pi86  & n348;
  assign n2299 = n346 & n1975;
  assign n2300 = ~n2297 & ~n2298;
  assign n2301 = ~n2296 & n2300;
  assign n2302 = ~n2299 & n2301;
  assign n2303 = pi5  & n2302;
  assign n2304 = ~pi5  & ~n2302;
  assign n2305 = ~n2303 & ~n2304;
  assign n2306 = ~n2260 & ~n2262;
  assign n2307 = ~n2243 & ~n2247;
  assign n2308 = ~n2221 & ~n2224;
  assign n2309 = ~n2215 & ~n2218;
  assign n2310 = pi69  & n1661;
  assign n2311 = pi70  & n1500;
  assign n2312 = pi71  & n1495;
  assign n2313 = n460 & n1493;
  assign n2314 = ~n2311 & ~n2312;
  assign n2315 = ~n2310 & n2314;
  assign n2316 = ~n2313 & n2315;
  assign n2317 = pi20  & n2316;
  assign n2318 = ~pi20  & ~n2316;
  assign n2319 = ~n2317 & ~n2318;
  assign n2320 = ~n2199 & ~n2202;
  assign n2321 = pi66  & n2053;
  assign n2322 = pi67  & n1893;
  assign n2323 = pi68  & n1888;
  assign n2324 = n334 & n1886;
  assign n2325 = ~n2322 & ~n2323;
  assign n2326 = ~n2321 & n2325;
  assign n2327 = ~n2324 & n2326;
  assign n2328 = pi23  & n2327;
  assign n2329 = ~pi23  & ~n2327;
  assign n2330 = ~n2328 & ~n2329;
  assign n2331 = pi26  & n2197;
  assign n2332 = ~pi25  & ~pi26 ;
  assign n2333 = pi25  & pi26 ;
  assign n2334 = ~n2332 & ~n2333;
  assign n2335 = n2196 & n2334;
  assign n2336 = n265 & n2335;
  assign n2337 = n2196 & ~n2334;
  assign n2338 = pi65  & n2337;
  assign n2339 = ~pi24  & ~pi25 ;
  assign n2340 = pi24  & pi25 ;
  assign n2341 = ~n2339 & ~n2340;
  assign n2342 = ~n2196 & n2341;
  assign n2343 = pi64  & n2342;
  assign n2344 = ~n2336 & ~n2338;
  assign n2345 = ~n2343 & n2344;
  assign n2346 = n2331 & ~n2345;
  assign n2347 = ~n2331 & n2345;
  assign n2348 = ~n2346 & ~n2347;
  assign n2349 = ~n2330 & n2348;
  assign n2350 = n2330 & ~n2348;
  assign n2351 = ~n2349 & ~n2350;
  assign n2352 = ~n2320 & n2351;
  assign n2353 = n2320 & ~n2351;
  assign n2354 = ~n2352 & ~n2353;
  assign n2355 = ~n2319 & n2354;
  assign n2356 = n2319 & ~n2354;
  assign n2357 = ~n2355 & ~n2356;
  assign n2358 = ~n2309 & n2357;
  assign n2359 = n2309 & ~n2357;
  assign n2360 = ~n2358 & ~n2359;
  assign n2361 = pi72  & n1296;
  assign n2362 = pi73  & n1207;
  assign n2363 = pi74  & n1202;
  assign n2364 = n689 & n1200;
  assign n2365 = ~n2362 & ~n2363;
  assign n2366 = ~n2361 & n2365;
  assign n2367 = ~n2364 & n2366;
  assign n2368 = pi17  & n2367;
  assign n2369 = ~pi17  & ~n2367;
  assign n2370 = ~n2368 & ~n2369;
  assign n2371 = n2360 & ~n2370;
  assign n2372 = ~n2360 & n2370;
  assign n2373 = ~n2371 & ~n2372;
  assign n2374 = n2308 & ~n2373;
  assign n2375 = ~n2308 & n2373;
  assign n2376 = ~n2374 & ~n2375;
  assign n2377 = pi75  & n1006;
  assign n2378 = pi76  & n897;
  assign n2379 = pi77  & n892;
  assign n2380 = n865 & n890;
  assign n2381 = ~n2378 & ~n2379;
  assign n2382 = ~n2377 & n2381;
  assign n2383 = ~n2380 & n2382;
  assign n2384 = pi14  & n2383;
  assign n2385 = ~pi14  & ~n2383;
  assign n2386 = ~n2384 & ~n2385;
  assign n2387 = ~n2376 & n2386;
  assign n2388 = n2376 & ~n2386;
  assign n2389 = ~n2387 & ~n2388;
  assign n2390 = ~n2228 & ~n2230;
  assign n2391 = n2389 & ~n2390;
  assign n2392 = ~n2389 & n2390;
  assign n2393 = ~n2391 & ~n2392;
  assign n2394 = pi78  & n750;
  assign n2395 = pi79  & n651;
  assign n2396 = pi80  & n646;
  assign n2397 = n644 & n1144;
  assign n2398 = ~n2395 & ~n2396;
  assign n2399 = ~n2394 & n2398;
  assign n2400 = ~n2397 & n2399;
  assign n2401 = pi11  & n2400;
  assign n2402 = ~pi11  & ~n2400;
  assign n2403 = ~n2401 & ~n2402;
  assign n2404 = n2393 & ~n2403;
  assign n2405 = ~n2393 & n2403;
  assign n2406 = ~n2404 & ~n2405;
  assign n2407 = n2307 & ~n2406;
  assign n2408 = ~n2307 & n2406;
  assign n2409 = ~n2407 & ~n2408;
  assign n2410 = pi81  & n528;
  assign n2411 = pi82  & n490;
  assign n2412 = pi83  & n485;
  assign n2413 = n483 & n1577;
  assign n2414 = ~n2411 & ~n2412;
  assign n2415 = ~n2410 & n2414;
  assign n2416 = ~n2413 & n2415;
  assign n2417 = pi8  & n2416;
  assign n2418 = ~pi8  & ~n2416;
  assign n2419 = ~n2417 & ~n2418;
  assign n2420 = n2409 & ~n2419;
  assign n2421 = ~n2409 & n2419;
  assign n2422 = ~n2420 & ~n2421;
  assign n2423 = ~n2306 & n2422;
  assign n2424 = n2306 & ~n2422;
  assign n2425 = ~n2423 & ~n2424;
  assign n2426 = ~n2305 & n2425;
  assign n2427 = n2305 & ~n2425;
  assign n2428 = ~n2426 & ~n2427;
  assign n2429 = ~n2295 & n2428;
  assign n2430 = n2295 & ~n2428;
  assign n2431 = ~n2429 & ~n2430;
  assign n2432 = ~n2294 & n2431;
  assign n2433 = n2294 & ~n2431;
  assign n2434 = ~n2432 & ~n2433;
  assign n2435 = ~n2277 & n2434;
  assign n2436 = n2277 & ~n2434;
  assign po25  = ~n2435 & ~n2436;
  assign n2438 = ~n2432 & ~n2435;
  assign n2439 = pi90  & n269;
  assign n2440 = pi89  & n267;
  assign n2441 = pi88  & n282;
  assign n2442 = ~n2283 & ~n2285;
  assign n2443 = ~pi89  & ~pi90 ;
  assign n2444 = pi89  & pi90 ;
  assign n2445 = ~n2443 & ~n2444;
  assign n2446 = ~n2442 & n2445;
  assign n2447 = n2442 & ~n2445;
  assign n2448 = ~n2446 & ~n2447;
  assign n2449 = n262 & n2448;
  assign n2450 = ~n2439 & ~n2440;
  assign n2451 = ~n2441 & n2450;
  assign n2452 = ~n2449 & n2451;
  assign n2453 = pi2  & n2452;
  assign n2454 = ~pi2  & ~n2452;
  assign n2455 = ~n2453 & ~n2454;
  assign n2456 = ~n2426 & ~n2429;
  assign n2457 = ~n2420 & ~n2423;
  assign n2458 = ~n2404 & ~n2408;
  assign n2459 = pi79  & n750;
  assign n2460 = pi80  & n651;
  assign n2461 = pi81  & n646;
  assign n2462 = n644 & n1337;
  assign n2463 = ~n2460 & ~n2461;
  assign n2464 = ~n2459 & n2463;
  assign n2465 = ~n2462 & n2464;
  assign n2466 = pi11  & n2465;
  assign n2467 = ~pi11  & ~n2465;
  assign n2468 = ~n2466 & ~n2467;
  assign n2469 = ~n2388 & ~n2391;
  assign n2470 = ~n2371 & ~n2375;
  assign n2471 = pi73  & n1296;
  assign n2472 = pi74  & n1207;
  assign n2473 = pi75  & n1202;
  assign n2474 = n713 & n1200;
  assign n2475 = ~n2472 & ~n2473;
  assign n2476 = ~n2471 & n2475;
  assign n2477 = ~n2474 & n2476;
  assign n2478 = pi17  & n2477;
  assign n2479 = ~pi17  & ~n2477;
  assign n2480 = ~n2478 & ~n2479;
  assign n2481 = ~n2355 & ~n2358;
  assign n2482 = pi70  & n1661;
  assign n2483 = pi71  & n1500;
  assign n2484 = pi72  & n1495;
  assign n2485 = n551 & n1493;
  assign n2486 = ~n2483 & ~n2484;
  assign n2487 = ~n2482 & n2486;
  assign n2488 = ~n2485 & n2487;
  assign n2489 = pi20  & n2488;
  assign n2490 = ~pi20  & ~n2488;
  assign n2491 = ~n2489 & ~n2490;
  assign n2492 = ~n2349 & ~n2352;
  assign n2493 = pi67  & n2053;
  assign n2494 = pi68  & n1893;
  assign n2495 = pi69  & n1888;
  assign n2496 = n376 & n1886;
  assign n2497 = ~n2494 & ~n2495;
  assign n2498 = ~n2493 & n2497;
  assign n2499 = ~n2496 & n2498;
  assign n2500 = pi23  & n2499;
  assign n2501 = ~pi23  & ~n2499;
  assign n2502 = ~n2500 & ~n2501;
  assign n2503 = pi26  & ~n2197;
  assign n2504 = n2345 & n2503;
  assign n2505 = pi26  & ~n2504;
  assign n2506 = ~n287 & n2335;
  assign n2507 = pi65  & n2342;
  assign n2508 = pi66  & n2337;
  assign n2509 = ~n2196 & n2334;
  assign n2510 = ~n2341 & n2509;
  assign n2511 = pi64  & n2510;
  assign n2512 = ~n2506 & ~n2507;
  assign n2513 = ~n2508 & n2512;
  assign n2514 = ~n2511 & n2513;
  assign n2515 = ~n2505 & n2514;
  assign n2516 = n2505 & ~n2514;
  assign n2517 = ~n2515 & ~n2516;
  assign n2518 = ~n2502 & n2517;
  assign n2519 = n2502 & ~n2517;
  assign n2520 = ~n2518 & ~n2519;
  assign n2521 = ~n2492 & n2520;
  assign n2522 = n2492 & ~n2520;
  assign n2523 = ~n2521 & ~n2522;
  assign n2524 = n2491 & ~n2523;
  assign n2525 = ~n2491 & n2523;
  assign n2526 = ~n2524 & ~n2525;
  assign n2527 = ~n2481 & n2526;
  assign n2528 = n2481 & ~n2526;
  assign n2529 = ~n2527 & ~n2528;
  assign n2530 = n2480 & ~n2529;
  assign n2531 = ~n2480 & n2529;
  assign n2532 = ~n2530 & ~n2531;
  assign n2533 = ~n2470 & n2532;
  assign n2534 = n2470 & ~n2532;
  assign n2535 = ~n2533 & ~n2534;
  assign n2536 = pi76  & n1006;
  assign n2537 = pi77  & n897;
  assign n2538 = pi78  & n892;
  assign n2539 = n890 & n958;
  assign n2540 = ~n2537 & ~n2538;
  assign n2541 = ~n2536 & n2540;
  assign n2542 = ~n2539 & n2541;
  assign n2543 = pi14  & n2542;
  assign n2544 = ~pi14  & ~n2542;
  assign n2545 = ~n2543 & ~n2544;
  assign n2546 = n2535 & ~n2545;
  assign n2547 = ~n2535 & n2545;
  assign n2548 = ~n2546 & ~n2547;
  assign n2549 = ~n2469 & n2548;
  assign n2550 = n2469 & ~n2548;
  assign n2551 = ~n2549 & ~n2550;
  assign n2552 = ~n2468 & n2551;
  assign n2553 = n2468 & ~n2551;
  assign n2554 = ~n2552 & ~n2553;
  assign n2555 = n2458 & ~n2554;
  assign n2556 = ~n2458 & n2554;
  assign n2557 = ~n2555 & ~n2556;
  assign n2558 = pi82  & n528;
  assign n2559 = pi83  & n490;
  assign n2560 = pi84  & n485;
  assign n2561 = n483 & n1601;
  assign n2562 = ~n2559 & ~n2560;
  assign n2563 = ~n2558 & n2562;
  assign n2564 = ~n2561 & n2563;
  assign n2565 = pi8  & n2564;
  assign n2566 = ~pi8  & ~n2564;
  assign n2567 = ~n2565 & ~n2566;
  assign n2568 = n2557 & ~n2567;
  assign n2569 = ~n2557 & n2567;
  assign n2570 = ~n2568 & ~n2569;
  assign n2571 = n2457 & ~n2570;
  assign n2572 = ~n2457 & n2570;
  assign n2573 = ~n2571 & ~n2572;
  assign n2574 = pi85  & n391;
  assign n2575 = pi86  & n353;
  assign n2576 = pi87  & n348;
  assign n2577 = n346 & n2116;
  assign n2578 = ~n2575 & ~n2576;
  assign n2579 = ~n2574 & n2578;
  assign n2580 = ~n2577 & n2579;
  assign n2581 = pi5  & n2580;
  assign n2582 = ~pi5  & ~n2580;
  assign n2583 = ~n2581 & ~n2582;
  assign n2584 = n2573 & ~n2583;
  assign n2585 = ~n2573 & n2583;
  assign n2586 = ~n2584 & ~n2585;
  assign n2587 = ~n2456 & n2586;
  assign n2588 = n2456 & ~n2586;
  assign n2589 = ~n2587 & ~n2588;
  assign n2590 = ~n2455 & n2589;
  assign n2591 = n2455 & ~n2589;
  assign n2592 = ~n2590 & ~n2591;
  assign n2593 = ~n2438 & n2592;
  assign n2594 = n2438 & ~n2592;
  assign po26  = ~n2593 & ~n2594;
  assign n2596 = ~n2590 & ~n2593;
  assign n2597 = ~n2584 & ~n2587;
  assign n2598 = ~n2552 & ~n2556;
  assign n2599 = ~n2546 & ~n2549;
  assign n2600 = ~n2531 & ~n2533;
  assign n2601 = pi74  & n1296;
  assign n2602 = pi75  & n1207;
  assign n2603 = pi76  & n1202;
  assign n2604 = n841 & n1200;
  assign n2605 = ~n2602 & ~n2603;
  assign n2606 = ~n2601 & n2605;
  assign n2607 = ~n2604 & n2606;
  assign n2608 = pi17  & n2607;
  assign n2609 = ~pi17  & ~n2607;
  assign n2610 = ~n2608 & ~n2609;
  assign n2611 = ~n2525 & ~n2527;
  assign n2612 = pi71  & n1661;
  assign n2613 = pi72  & n1500;
  assign n2614 = pi73  & n1495;
  assign n2615 = n613 & n1493;
  assign n2616 = ~n2613 & ~n2614;
  assign n2617 = ~n2612 & n2616;
  assign n2618 = ~n2615 & n2617;
  assign n2619 = pi20  & n2618;
  assign n2620 = ~pi20  & ~n2618;
  assign n2621 = ~n2619 & ~n2620;
  assign n2622 = ~n2518 & ~n2521;
  assign n2623 = pi65  & n2510;
  assign n2624 = pi66  & n2342;
  assign n2625 = pi67  & n2337;
  assign n2626 = n305 & n2335;
  assign n2627 = ~n2624 & ~n2625;
  assign n2628 = ~n2623 & n2627;
  assign n2629 = ~n2626 & n2628;
  assign n2630 = pi26  & n2629;
  assign n2631 = ~pi26  & ~n2629;
  assign n2632 = ~n2630 & ~n2631;
  assign n2633 = ~pi26  & ~pi27 ;
  assign n2634 = pi26  & pi27 ;
  assign n2635 = ~n2633 & ~n2634;
  assign n2636 = pi64  & n2635;
  assign n2637 = n2504 & n2514;
  assign n2638 = n2636 & n2637;
  assign n2639 = ~n2636 & ~n2637;
  assign n2640 = ~n2638 & ~n2639;
  assign n2641 = ~n2632 & n2640;
  assign n2642 = n2632 & ~n2640;
  assign n2643 = ~n2641 & ~n2642;
  assign n2644 = pi68  & n2053;
  assign n2645 = pi69  & n1893;
  assign n2646 = pi70  & n1888;
  assign n2647 = n415 & n1886;
  assign n2648 = ~n2645 & ~n2646;
  assign n2649 = ~n2644 & n2648;
  assign n2650 = ~n2647 & n2649;
  assign n2651 = pi23  & n2650;
  assign n2652 = ~pi23  & ~n2650;
  assign n2653 = ~n2651 & ~n2652;
  assign n2654 = n2643 & ~n2653;
  assign n2655 = ~n2643 & n2653;
  assign n2656 = ~n2654 & ~n2655;
  assign n2657 = ~n2622 & n2656;
  assign n2658 = n2622 & ~n2656;
  assign n2659 = ~n2657 & ~n2658;
  assign n2660 = ~n2621 & n2659;
  assign n2661 = n2621 & ~n2659;
  assign n2662 = ~n2660 & ~n2661;
  assign n2663 = ~n2611 & n2662;
  assign n2664 = n2611 & ~n2662;
  assign n2665 = ~n2663 & ~n2664;
  assign n2666 = n2610 & ~n2665;
  assign n2667 = ~n2610 & n2665;
  assign n2668 = ~n2666 & ~n2667;
  assign n2669 = ~n2600 & n2668;
  assign n2670 = n2600 & ~n2668;
  assign n2671 = ~n2669 & ~n2670;
  assign n2672 = pi77  & n1006;
  assign n2673 = pi78  & n897;
  assign n2674 = pi79  & n892;
  assign n2675 = n890 & n1048;
  assign n2676 = ~n2673 & ~n2674;
  assign n2677 = ~n2672 & n2676;
  assign n2678 = ~n2675 & n2677;
  assign n2679 = pi14  & n2678;
  assign n2680 = ~pi14  & ~n2678;
  assign n2681 = ~n2679 & ~n2680;
  assign n2682 = n2671 & ~n2681;
  assign n2683 = ~n2671 & n2681;
  assign n2684 = ~n2682 & ~n2683;
  assign n2685 = n2599 & ~n2684;
  assign n2686 = ~n2599 & n2684;
  assign n2687 = ~n2685 & ~n2686;
  assign n2688 = pi80  & n750;
  assign n2689 = pi81  & n651;
  assign n2690 = pi82  & n646;
  assign n2691 = n644 & n1450;
  assign n2692 = ~n2689 & ~n2690;
  assign n2693 = ~n2688 & n2692;
  assign n2694 = ~n2691 & n2693;
  assign n2695 = pi11  & n2694;
  assign n2696 = ~pi11  & ~n2694;
  assign n2697 = ~n2695 & ~n2696;
  assign n2698 = n2687 & ~n2697;
  assign n2699 = ~n2687 & n2697;
  assign n2700 = ~n2698 & ~n2699;
  assign n2701 = n2598 & ~n2700;
  assign n2702 = ~n2598 & n2700;
  assign n2703 = ~n2701 & ~n2702;
  assign n2704 = pi83  & n528;
  assign n2705 = pi84  & n490;
  assign n2706 = pi85  & n485;
  assign n2707 = n483 & n1831;
  assign n2708 = ~n2705 & ~n2706;
  assign n2709 = ~n2704 & n2708;
  assign n2710 = ~n2707 & n2709;
  assign n2711 = pi8  & n2710;
  assign n2712 = ~pi8  & ~n2710;
  assign n2713 = ~n2711 & ~n2712;
  assign n2714 = ~n2703 & n2713;
  assign n2715 = n2703 & ~n2713;
  assign n2716 = ~n2714 & ~n2715;
  assign n2717 = ~n2568 & ~n2572;
  assign n2718 = n2716 & ~n2717;
  assign n2719 = ~n2716 & n2717;
  assign n2720 = ~n2718 & ~n2719;
  assign n2721 = pi86  & n391;
  assign n2722 = pi87  & n353;
  assign n2723 = pi88  & n348;
  assign n2724 = n346 & n2140;
  assign n2725 = ~n2722 & ~n2723;
  assign n2726 = ~n2721 & n2725;
  assign n2727 = ~n2724 & n2726;
  assign n2728 = pi5  & n2727;
  assign n2729 = ~pi5  & ~n2727;
  assign n2730 = ~n2728 & ~n2729;
  assign n2731 = n2720 & ~n2730;
  assign n2732 = ~n2720 & n2730;
  assign n2733 = ~n2731 & ~n2732;
  assign n2734 = n2597 & ~n2733;
  assign n2735 = ~n2597 & n2733;
  assign n2736 = ~n2734 & ~n2735;
  assign n2737 = pi91  & n269;
  assign n2738 = pi90  & n267;
  assign n2739 = pi89  & n282;
  assign n2740 = ~n2444 & ~n2446;
  assign n2741 = ~pi90  & ~pi91 ;
  assign n2742 = pi90  & pi91 ;
  assign n2743 = ~n2741 & ~n2742;
  assign n2744 = ~n2740 & n2743;
  assign n2745 = n2740 & ~n2743;
  assign n2746 = ~n2744 & ~n2745;
  assign n2747 = n262 & n2746;
  assign n2748 = ~n2737 & ~n2738;
  assign n2749 = ~n2739 & n2748;
  assign n2750 = ~n2747 & n2749;
  assign n2751 = pi2  & n2750;
  assign n2752 = ~pi2  & ~n2750;
  assign n2753 = ~n2751 & ~n2752;
  assign n2754 = ~n2736 & n2753;
  assign n2755 = n2736 & ~n2753;
  assign n2756 = ~n2754 & ~n2755;
  assign n2757 = ~n2596 & n2756;
  assign n2758 = n2596 & ~n2756;
  assign po27  = ~n2757 & ~n2758;
  assign n2760 = ~n2755 & ~n2757;
  assign n2761 = ~n2731 & ~n2735;
  assign n2762 = ~n2698 & ~n2702;
  assign n2763 = ~n2682 & ~n2686;
  assign n2764 = pi78  & n1006;
  assign n2765 = pi79  & n897;
  assign n2766 = pi80  & n892;
  assign n2767 = n890 & n1144;
  assign n2768 = ~n2765 & ~n2766;
  assign n2769 = ~n2764 & n2768;
  assign n2770 = ~n2767 & n2769;
  assign n2771 = pi14  & n2770;
  assign n2772 = ~pi14  & ~n2770;
  assign n2773 = ~n2771 & ~n2772;
  assign n2774 = ~n2667 & ~n2669;
  assign n2775 = ~n2660 & ~n2663;
  assign n2776 = ~n2654 & ~n2657;
  assign n2777 = pi69  & n2053;
  assign n2778 = pi70  & n1893;
  assign n2779 = pi71  & n1888;
  assign n2780 = n460 & n1886;
  assign n2781 = ~n2778 & ~n2779;
  assign n2782 = ~n2777 & n2781;
  assign n2783 = ~n2780 & n2782;
  assign n2784 = pi23  & n2783;
  assign n2785 = ~pi23  & ~n2783;
  assign n2786 = ~n2784 & ~n2785;
  assign n2787 = ~n2638 & ~n2641;
  assign n2788 = pi66  & n2510;
  assign n2789 = pi67  & n2342;
  assign n2790 = pi68  & n2337;
  assign n2791 = n334 & n2335;
  assign n2792 = ~n2789 & ~n2790;
  assign n2793 = ~n2788 & n2792;
  assign n2794 = ~n2791 & n2793;
  assign n2795 = pi26  & n2794;
  assign n2796 = ~pi26  & ~n2794;
  assign n2797 = ~n2795 & ~n2796;
  assign n2798 = pi29  & n2636;
  assign n2799 = ~pi28  & ~pi29 ;
  assign n2800 = pi28  & pi29 ;
  assign n2801 = ~n2799 & ~n2800;
  assign n2802 = n2635 & n2801;
  assign n2803 = n265 & n2802;
  assign n2804 = n2635 & ~n2801;
  assign n2805 = pi65  & n2804;
  assign n2806 = ~pi27  & ~pi28 ;
  assign n2807 = pi27  & pi28 ;
  assign n2808 = ~n2806 & ~n2807;
  assign n2809 = ~n2635 & n2808;
  assign n2810 = pi64  & n2809;
  assign n2811 = ~n2803 & ~n2805;
  assign n2812 = ~n2810 & n2811;
  assign n2813 = n2798 & ~n2812;
  assign n2814 = ~n2798 & n2812;
  assign n2815 = ~n2813 & ~n2814;
  assign n2816 = ~n2797 & n2815;
  assign n2817 = n2797 & ~n2815;
  assign n2818 = ~n2816 & ~n2817;
  assign n2819 = ~n2787 & n2818;
  assign n2820 = n2787 & ~n2818;
  assign n2821 = ~n2819 & ~n2820;
  assign n2822 = ~n2786 & n2821;
  assign n2823 = n2786 & ~n2821;
  assign n2824 = ~n2822 & ~n2823;
  assign n2825 = ~n2776 & n2824;
  assign n2826 = n2776 & ~n2824;
  assign n2827 = ~n2825 & ~n2826;
  assign n2828 = pi72  & n1661;
  assign n2829 = pi73  & n1500;
  assign n2830 = pi74  & n1495;
  assign n2831 = n689 & n1493;
  assign n2832 = ~n2829 & ~n2830;
  assign n2833 = ~n2828 & n2832;
  assign n2834 = ~n2831 & n2833;
  assign n2835 = pi20  & n2834;
  assign n2836 = ~pi20  & ~n2834;
  assign n2837 = ~n2835 & ~n2836;
  assign n2838 = n2827 & ~n2837;
  assign n2839 = ~n2827 & n2837;
  assign n2840 = ~n2838 & ~n2839;
  assign n2841 = n2775 & ~n2840;
  assign n2842 = ~n2775 & n2840;
  assign n2843 = ~n2841 & ~n2842;
  assign n2844 = pi75  & n1296;
  assign n2845 = pi76  & n1207;
  assign n2846 = pi77  & n1202;
  assign n2847 = n865 & n1200;
  assign n2848 = ~n2845 & ~n2846;
  assign n2849 = ~n2844 & n2848;
  assign n2850 = ~n2847 & n2849;
  assign n2851 = pi17  & n2850;
  assign n2852 = ~pi17  & ~n2850;
  assign n2853 = ~n2851 & ~n2852;
  assign n2854 = n2843 & ~n2853;
  assign n2855 = ~n2843 & n2853;
  assign n2856 = ~n2854 & ~n2855;
  assign n2857 = ~n2774 & n2856;
  assign n2858 = n2774 & ~n2856;
  assign n2859 = ~n2857 & ~n2858;
  assign n2860 = ~n2773 & n2859;
  assign n2861 = n2773 & ~n2859;
  assign n2862 = ~n2860 & ~n2861;
  assign n2863 = n2763 & ~n2862;
  assign n2864 = ~n2763 & n2862;
  assign n2865 = ~n2863 & ~n2864;
  assign n2866 = pi81  & n750;
  assign n2867 = pi82  & n651;
  assign n2868 = pi83  & n646;
  assign n2869 = n644 & n1577;
  assign n2870 = ~n2867 & ~n2868;
  assign n2871 = ~n2866 & n2870;
  assign n2872 = ~n2869 & n2871;
  assign n2873 = pi11  & n2872;
  assign n2874 = ~pi11  & ~n2872;
  assign n2875 = ~n2873 & ~n2874;
  assign n2876 = n2865 & ~n2875;
  assign n2877 = ~n2865 & n2875;
  assign n2878 = ~n2876 & ~n2877;
  assign n2879 = n2762 & ~n2878;
  assign n2880 = ~n2762 & n2878;
  assign n2881 = ~n2879 & ~n2880;
  assign n2882 = pi84  & n528;
  assign n2883 = pi85  & n490;
  assign n2884 = pi86  & n485;
  assign n2885 = n483 & n1975;
  assign n2886 = ~n2883 & ~n2884;
  assign n2887 = ~n2882 & n2886;
  assign n2888 = ~n2885 & n2887;
  assign n2889 = pi8  & n2888;
  assign n2890 = ~pi8  & ~n2888;
  assign n2891 = ~n2889 & ~n2890;
  assign n2892 = ~n2881 & n2891;
  assign n2893 = n2881 & ~n2891;
  assign n2894 = ~n2892 & ~n2893;
  assign n2895 = ~n2715 & ~n2718;
  assign n2896 = n2894 & ~n2895;
  assign n2897 = ~n2894 & n2895;
  assign n2898 = ~n2896 & ~n2897;
  assign n2899 = pi87  & n391;
  assign n2900 = pi88  & n353;
  assign n2901 = pi89  & n348;
  assign n2902 = n346 & n2287;
  assign n2903 = ~n2900 & ~n2901;
  assign n2904 = ~n2899 & n2903;
  assign n2905 = ~n2902 & n2904;
  assign n2906 = pi5  & n2905;
  assign n2907 = ~pi5  & ~n2905;
  assign n2908 = ~n2906 & ~n2907;
  assign n2909 = n2898 & ~n2908;
  assign n2910 = ~n2898 & n2908;
  assign n2911 = ~n2909 & ~n2910;
  assign n2912 = n2761 & ~n2911;
  assign n2913 = ~n2761 & n2911;
  assign n2914 = ~n2912 & ~n2913;
  assign n2915 = pi92  & n269;
  assign n2916 = pi91  & n267;
  assign n2917 = pi90  & n282;
  assign n2918 = ~n2742 & ~n2744;
  assign n2919 = ~pi91  & ~pi92 ;
  assign n2920 = pi91  & pi92 ;
  assign n2921 = ~n2919 & ~n2920;
  assign n2922 = ~n2918 & n2921;
  assign n2923 = n2918 & ~n2921;
  assign n2924 = ~n2922 & ~n2923;
  assign n2925 = n262 & n2924;
  assign n2926 = ~n2915 & ~n2916;
  assign n2927 = ~n2917 & n2926;
  assign n2928 = ~n2925 & n2927;
  assign n2929 = pi2  & n2928;
  assign n2930 = ~pi2  & ~n2928;
  assign n2931 = ~n2929 & ~n2930;
  assign n2932 = ~n2914 & n2931;
  assign n2933 = n2914 & ~n2931;
  assign n2934 = ~n2932 & ~n2933;
  assign n2935 = ~n2760 & n2934;
  assign n2936 = n2760 & ~n2934;
  assign po28  = ~n2935 & ~n2936;
  assign n2938 = ~n2933 & ~n2935;
  assign n2939 = pi93  & n269;
  assign n2940 = pi92  & n267;
  assign n2941 = pi91  & n282;
  assign n2942 = ~n2920 & ~n2922;
  assign n2943 = ~pi92  & ~pi93 ;
  assign n2944 = pi92  & pi93 ;
  assign n2945 = ~n2943 & ~n2944;
  assign n2946 = ~n2942 & n2945;
  assign n2947 = n2942 & ~n2945;
  assign n2948 = ~n2946 & ~n2947;
  assign n2949 = n262 & n2948;
  assign n2950 = ~n2939 & ~n2940;
  assign n2951 = ~n2941 & n2950;
  assign n2952 = ~n2949 & n2951;
  assign n2953 = pi2  & n2952;
  assign n2954 = ~pi2  & ~n2952;
  assign n2955 = ~n2953 & ~n2954;
  assign n2956 = ~n2909 & ~n2913;
  assign n2957 = pi88  & n391;
  assign n2958 = pi89  & n353;
  assign n2959 = pi90  & n348;
  assign n2960 = n346 & n2448;
  assign n2961 = ~n2958 & ~n2959;
  assign n2962 = ~n2957 & n2961;
  assign n2963 = ~n2960 & n2962;
  assign n2964 = pi5  & n2963;
  assign n2965 = ~pi5  & ~n2963;
  assign n2966 = ~n2964 & ~n2965;
  assign n2967 = ~n2893 & ~n2896;
  assign n2968 = ~n2876 & ~n2880;
  assign n2969 = ~n2860 & ~n2864;
  assign n2970 = ~n2854 & ~n2857;
  assign n2971 = ~n2838 & ~n2842;
  assign n2972 = pi73  & n1661;
  assign n2973 = pi74  & n1500;
  assign n2974 = pi75  & n1495;
  assign n2975 = n713 & n1493;
  assign n2976 = ~n2973 & ~n2974;
  assign n2977 = ~n2972 & n2976;
  assign n2978 = ~n2975 & n2977;
  assign n2979 = pi20  & n2978;
  assign n2980 = ~pi20  & ~n2978;
  assign n2981 = ~n2979 & ~n2980;
  assign n2982 = ~n2822 & ~n2825;
  assign n2983 = pi70  & n2053;
  assign n2984 = pi71  & n1893;
  assign n2985 = pi72  & n1888;
  assign n2986 = n551 & n1886;
  assign n2987 = ~n2984 & ~n2985;
  assign n2988 = ~n2983 & n2987;
  assign n2989 = ~n2986 & n2988;
  assign n2990 = pi23  & n2989;
  assign n2991 = ~pi23  & ~n2989;
  assign n2992 = ~n2990 & ~n2991;
  assign n2993 = ~n2816 & ~n2819;
  assign n2994 = pi67  & n2510;
  assign n2995 = pi68  & n2342;
  assign n2996 = pi69  & n2337;
  assign n2997 = n376 & n2335;
  assign n2998 = ~n2995 & ~n2996;
  assign n2999 = ~n2994 & n2998;
  assign n3000 = ~n2997 & n2999;
  assign n3001 = pi26  & n3000;
  assign n3002 = ~pi26  & ~n3000;
  assign n3003 = ~n3001 & ~n3002;
  assign n3004 = pi29  & ~n2636;
  assign n3005 = n2812 & n3004;
  assign n3006 = pi29  & ~n3005;
  assign n3007 = ~n287 & n2802;
  assign n3008 = pi65  & n2809;
  assign n3009 = pi66  & n2804;
  assign n3010 = ~n2635 & n2801;
  assign n3011 = ~n2808 & n3010;
  assign n3012 = pi64  & n3011;
  assign n3013 = ~n3007 & ~n3008;
  assign n3014 = ~n3009 & n3013;
  assign n3015 = ~n3012 & n3014;
  assign n3016 = ~n3006 & n3015;
  assign n3017 = n3006 & ~n3015;
  assign n3018 = ~n3016 & ~n3017;
  assign n3019 = ~n3003 & n3018;
  assign n3020 = n3003 & ~n3018;
  assign n3021 = ~n3019 & ~n3020;
  assign n3022 = ~n2993 & n3021;
  assign n3023 = n2993 & ~n3021;
  assign n3024 = ~n3022 & ~n3023;
  assign n3025 = n2992 & ~n3024;
  assign n3026 = ~n2992 & n3024;
  assign n3027 = ~n3025 & ~n3026;
  assign n3028 = ~n2982 & n3027;
  assign n3029 = n2982 & ~n3027;
  assign n3030 = ~n3028 & ~n3029;
  assign n3031 = n2981 & ~n3030;
  assign n3032 = ~n2981 & n3030;
  assign n3033 = ~n3031 & ~n3032;
  assign n3034 = ~n2971 & n3033;
  assign n3035 = n2971 & ~n3033;
  assign n3036 = ~n3034 & ~n3035;
  assign n3037 = pi76  & n1296;
  assign n3038 = pi77  & n1207;
  assign n3039 = pi78  & n1202;
  assign n3040 = n958 & n1200;
  assign n3041 = ~n3038 & ~n3039;
  assign n3042 = ~n3037 & n3041;
  assign n3043 = ~n3040 & n3042;
  assign n3044 = pi17  & n3043;
  assign n3045 = ~pi17  & ~n3043;
  assign n3046 = ~n3044 & ~n3045;
  assign n3047 = n3036 & ~n3046;
  assign n3048 = ~n3036 & n3046;
  assign n3049 = ~n3047 & ~n3048;
  assign n3050 = n2970 & ~n3049;
  assign n3051 = ~n2970 & n3049;
  assign n3052 = ~n3050 & ~n3051;
  assign n3053 = pi79  & n1006;
  assign n3054 = pi80  & n897;
  assign n3055 = pi81  & n892;
  assign n3056 = n890 & n1337;
  assign n3057 = ~n3054 & ~n3055;
  assign n3058 = ~n3053 & n3057;
  assign n3059 = ~n3056 & n3058;
  assign n3060 = pi14  & n3059;
  assign n3061 = ~pi14  & ~n3059;
  assign n3062 = ~n3060 & ~n3061;
  assign n3063 = n3052 & ~n3062;
  assign n3064 = ~n3052 & n3062;
  assign n3065 = ~n3063 & ~n3064;
  assign n3066 = n2969 & ~n3065;
  assign n3067 = ~n2969 & n3065;
  assign n3068 = ~n3066 & ~n3067;
  assign n3069 = pi82  & n750;
  assign n3070 = pi83  & n651;
  assign n3071 = pi84  & n646;
  assign n3072 = n644 & n1601;
  assign n3073 = ~n3070 & ~n3071;
  assign n3074 = ~n3069 & n3073;
  assign n3075 = ~n3072 & n3074;
  assign n3076 = pi11  & n3075;
  assign n3077 = ~pi11  & ~n3075;
  assign n3078 = ~n3076 & ~n3077;
  assign n3079 = n3068 & ~n3078;
  assign n3080 = ~n3068 & n3078;
  assign n3081 = ~n3079 & ~n3080;
  assign n3082 = ~n2968 & n3081;
  assign n3083 = n2968 & ~n3081;
  assign n3084 = ~n3082 & ~n3083;
  assign n3085 = pi85  & n528;
  assign n3086 = pi86  & n490;
  assign n3087 = pi87  & n485;
  assign n3088 = n483 & n2116;
  assign n3089 = ~n3086 & ~n3087;
  assign n3090 = ~n3085 & n3089;
  assign n3091 = ~n3088 & n3090;
  assign n3092 = pi8  & n3091;
  assign n3093 = ~pi8  & ~n3091;
  assign n3094 = ~n3092 & ~n3093;
  assign n3095 = n3084 & ~n3094;
  assign n3096 = ~n3084 & n3094;
  assign n3097 = ~n3095 & ~n3096;
  assign n3098 = ~n2967 & n3097;
  assign n3099 = n2967 & ~n3097;
  assign n3100 = ~n3098 & ~n3099;
  assign n3101 = ~n2966 & n3100;
  assign n3102 = n2966 & ~n3100;
  assign n3103 = ~n3101 & ~n3102;
  assign n3104 = ~n2956 & n3103;
  assign n3105 = n2956 & ~n3103;
  assign n3106 = ~n3104 & ~n3105;
  assign n3107 = ~n2955 & n3106;
  assign n3108 = n2955 & ~n3106;
  assign n3109 = ~n3107 & ~n3108;
  assign n3110 = ~n2938 & n3109;
  assign n3111 = n2938 & ~n3109;
  assign po29  = ~n3110 & ~n3111;
  assign n3113 = ~n3107 & ~n3110;
  assign n3114 = ~n3101 & ~n3104;
  assign n3115 = ~n3095 & ~n3098;
  assign n3116 = pi86  & n528;
  assign n3117 = pi87  & n490;
  assign n3118 = pi88  & n485;
  assign n3119 = n483 & n2140;
  assign n3120 = ~n3117 & ~n3118;
  assign n3121 = ~n3116 & n3120;
  assign n3122 = ~n3119 & n3121;
  assign n3123 = pi8  & n3122;
  assign n3124 = ~pi8  & ~n3122;
  assign n3125 = ~n3123 & ~n3124;
  assign n3126 = ~n3079 & ~n3082;
  assign n3127 = ~n3063 & ~n3067;
  assign n3128 = ~n3047 & ~n3051;
  assign n3129 = ~n3032 & ~n3034;
  assign n3130 = pi74  & n1661;
  assign n3131 = pi75  & n1500;
  assign n3132 = pi76  & n1495;
  assign n3133 = n841 & n1493;
  assign n3134 = ~n3131 & ~n3132;
  assign n3135 = ~n3130 & n3134;
  assign n3136 = ~n3133 & n3135;
  assign n3137 = pi20  & n3136;
  assign n3138 = ~pi20  & ~n3136;
  assign n3139 = ~n3137 & ~n3138;
  assign n3140 = ~n3026 & ~n3028;
  assign n3141 = pi71  & n2053;
  assign n3142 = pi72  & n1893;
  assign n3143 = pi73  & n1888;
  assign n3144 = n613 & n1886;
  assign n3145 = ~n3142 & ~n3143;
  assign n3146 = ~n3141 & n3145;
  assign n3147 = ~n3144 & n3146;
  assign n3148 = pi23  & n3147;
  assign n3149 = ~pi23  & ~n3147;
  assign n3150 = ~n3148 & ~n3149;
  assign n3151 = ~n3019 & ~n3022;
  assign n3152 = pi65  & n3011;
  assign n3153 = pi66  & n2809;
  assign n3154 = pi67  & n2804;
  assign n3155 = n305 & n2802;
  assign n3156 = ~n3153 & ~n3154;
  assign n3157 = ~n3152 & n3156;
  assign n3158 = ~n3155 & n3157;
  assign n3159 = pi29  & n3158;
  assign n3160 = ~pi29  & ~n3158;
  assign n3161 = ~n3159 & ~n3160;
  assign n3162 = ~pi29  & ~pi30 ;
  assign n3163 = pi29  & pi30 ;
  assign n3164 = ~n3162 & ~n3163;
  assign n3165 = pi64  & n3164;
  assign n3166 = n3005 & n3015;
  assign n3167 = n3165 & n3166;
  assign n3168 = ~n3165 & ~n3166;
  assign n3169 = ~n3167 & ~n3168;
  assign n3170 = ~n3161 & n3169;
  assign n3171 = n3161 & ~n3169;
  assign n3172 = ~n3170 & ~n3171;
  assign n3173 = pi68  & n2510;
  assign n3174 = pi69  & n2342;
  assign n3175 = pi70  & n2337;
  assign n3176 = n415 & n2335;
  assign n3177 = ~n3174 & ~n3175;
  assign n3178 = ~n3173 & n3177;
  assign n3179 = ~n3176 & n3178;
  assign n3180 = pi26  & n3179;
  assign n3181 = ~pi26  & ~n3179;
  assign n3182 = ~n3180 & ~n3181;
  assign n3183 = n3172 & ~n3182;
  assign n3184 = ~n3172 & n3182;
  assign n3185 = ~n3183 & ~n3184;
  assign n3186 = ~n3151 & n3185;
  assign n3187 = n3151 & ~n3185;
  assign n3188 = ~n3186 & ~n3187;
  assign n3189 = ~n3150 & n3188;
  assign n3190 = n3150 & ~n3188;
  assign n3191 = ~n3189 & ~n3190;
  assign n3192 = ~n3140 & n3191;
  assign n3193 = n3140 & ~n3191;
  assign n3194 = ~n3192 & ~n3193;
  assign n3195 = n3139 & ~n3194;
  assign n3196 = ~n3139 & n3194;
  assign n3197 = ~n3195 & ~n3196;
  assign n3198 = ~n3129 & n3197;
  assign n3199 = n3129 & ~n3197;
  assign n3200 = ~n3198 & ~n3199;
  assign n3201 = pi77  & n1296;
  assign n3202 = pi78  & n1207;
  assign n3203 = pi79  & n1202;
  assign n3204 = n1048 & n1200;
  assign n3205 = ~n3202 & ~n3203;
  assign n3206 = ~n3201 & n3205;
  assign n3207 = ~n3204 & n3206;
  assign n3208 = pi17  & n3207;
  assign n3209 = ~pi17  & ~n3207;
  assign n3210 = ~n3208 & ~n3209;
  assign n3211 = n3200 & ~n3210;
  assign n3212 = ~n3200 & n3210;
  assign n3213 = ~n3211 & ~n3212;
  assign n3214 = n3128 & ~n3213;
  assign n3215 = ~n3128 & n3213;
  assign n3216 = ~n3214 & ~n3215;
  assign n3217 = pi80  & n1006;
  assign n3218 = pi81  & n897;
  assign n3219 = pi82  & n892;
  assign n3220 = n890 & n1450;
  assign n3221 = ~n3218 & ~n3219;
  assign n3222 = ~n3217 & n3221;
  assign n3223 = ~n3220 & n3222;
  assign n3224 = pi14  & n3223;
  assign n3225 = ~pi14  & ~n3223;
  assign n3226 = ~n3224 & ~n3225;
  assign n3227 = n3216 & ~n3226;
  assign n3228 = ~n3216 & n3226;
  assign n3229 = ~n3227 & ~n3228;
  assign n3230 = n3127 & ~n3229;
  assign n3231 = ~n3127 & n3229;
  assign n3232 = ~n3230 & ~n3231;
  assign n3233 = pi83  & n750;
  assign n3234 = pi84  & n651;
  assign n3235 = pi85  & n646;
  assign n3236 = n644 & n1831;
  assign n3237 = ~n3234 & ~n3235;
  assign n3238 = ~n3233 & n3237;
  assign n3239 = ~n3236 & n3238;
  assign n3240 = pi11  & n3239;
  assign n3241 = ~pi11  & ~n3239;
  assign n3242 = ~n3240 & ~n3241;
  assign n3243 = n3232 & ~n3242;
  assign n3244 = ~n3232 & n3242;
  assign n3245 = ~n3243 & ~n3244;
  assign n3246 = ~n3126 & n3245;
  assign n3247 = n3126 & ~n3245;
  assign n3248 = ~n3246 & ~n3247;
  assign n3249 = ~n3125 & n3248;
  assign n3250 = n3125 & ~n3248;
  assign n3251 = ~n3249 & ~n3250;
  assign n3252 = n3115 & ~n3251;
  assign n3253 = ~n3115 & n3251;
  assign n3254 = ~n3252 & ~n3253;
  assign n3255 = pi89  & n391;
  assign n3256 = pi90  & n353;
  assign n3257 = pi91  & n348;
  assign n3258 = n346 & n2746;
  assign n3259 = ~n3256 & ~n3257;
  assign n3260 = ~n3255 & n3259;
  assign n3261 = ~n3258 & n3260;
  assign n3262 = pi5  & n3261;
  assign n3263 = ~pi5  & ~n3261;
  assign n3264 = ~n3262 & ~n3263;
  assign n3265 = n3254 & ~n3264;
  assign n3266 = ~n3254 & n3264;
  assign n3267 = ~n3265 & ~n3266;
  assign n3268 = n3114 & ~n3267;
  assign n3269 = ~n3114 & n3267;
  assign n3270 = ~n3268 & ~n3269;
  assign n3271 = pi94  & n269;
  assign n3272 = pi93  & n267;
  assign n3273 = pi92  & n282;
  assign n3274 = ~n2944 & ~n2946;
  assign n3275 = ~pi93  & ~pi94 ;
  assign n3276 = pi93  & pi94 ;
  assign n3277 = ~n3275 & ~n3276;
  assign n3278 = ~n3274 & n3277;
  assign n3279 = n3274 & ~n3277;
  assign n3280 = ~n3278 & ~n3279;
  assign n3281 = n262 & n3280;
  assign n3282 = ~n3271 & ~n3272;
  assign n3283 = ~n3273 & n3282;
  assign n3284 = ~n3281 & n3283;
  assign n3285 = pi2  & n3284;
  assign n3286 = ~pi2  & ~n3284;
  assign n3287 = ~n3285 & ~n3286;
  assign n3288 = n3270 & ~n3287;
  assign n3289 = ~n3270 & n3287;
  assign n3290 = ~n3288 & ~n3289;
  assign n3291 = ~n3113 & n3290;
  assign n3292 = n3113 & ~n3290;
  assign po30  = ~n3291 & ~n3292;
  assign n3294 = ~n3288 & ~n3291;
  assign n3295 = ~n3265 & ~n3269;
  assign n3296 = ~n3249 & ~n3253;
  assign n3297 = ~n3243 & ~n3246;
  assign n3298 = ~n3227 & ~n3231;
  assign n3299 = ~n3211 & ~n3215;
  assign n3300 = ~n3189 & ~n3192;
  assign n3301 = ~n3183 & ~n3186;
  assign n3302 = pi69  & n2510;
  assign n3303 = pi70  & n2342;
  assign n3304 = pi71  & n2337;
  assign n3305 = n460 & n2335;
  assign n3306 = ~n3303 & ~n3304;
  assign n3307 = ~n3302 & n3306;
  assign n3308 = ~n3305 & n3307;
  assign n3309 = pi26  & n3308;
  assign n3310 = ~pi26  & ~n3308;
  assign n3311 = ~n3309 & ~n3310;
  assign n3312 = ~n3167 & ~n3170;
  assign n3313 = pi66  & n3011;
  assign n3314 = pi67  & n2809;
  assign n3315 = pi68  & n2804;
  assign n3316 = n334 & n2802;
  assign n3317 = ~n3314 & ~n3315;
  assign n3318 = ~n3313 & n3317;
  assign n3319 = ~n3316 & n3318;
  assign n3320 = pi29  & n3319;
  assign n3321 = ~pi29  & ~n3319;
  assign n3322 = ~n3320 & ~n3321;
  assign n3323 = pi32  & n3165;
  assign n3324 = ~pi31  & ~pi32 ;
  assign n3325 = pi31  & pi32 ;
  assign n3326 = ~n3324 & ~n3325;
  assign n3327 = n3164 & n3326;
  assign n3328 = n265 & n3327;
  assign n3329 = n3164 & ~n3326;
  assign n3330 = pi65  & n3329;
  assign n3331 = ~pi30  & ~pi31 ;
  assign n3332 = pi30  & pi31 ;
  assign n3333 = ~n3331 & ~n3332;
  assign n3334 = ~n3164 & n3333;
  assign n3335 = pi64  & n3334;
  assign n3336 = ~n3328 & ~n3330;
  assign n3337 = ~n3335 & n3336;
  assign n3338 = n3323 & ~n3337;
  assign n3339 = ~n3323 & n3337;
  assign n3340 = ~n3338 & ~n3339;
  assign n3341 = ~n3322 & n3340;
  assign n3342 = n3322 & ~n3340;
  assign n3343 = ~n3341 & ~n3342;
  assign n3344 = ~n3312 & n3343;
  assign n3345 = n3312 & ~n3343;
  assign n3346 = ~n3344 & ~n3345;
  assign n3347 = ~n3311 & n3346;
  assign n3348 = n3311 & ~n3346;
  assign n3349 = ~n3347 & ~n3348;
  assign n3350 = ~n3301 & n3349;
  assign n3351 = n3301 & ~n3349;
  assign n3352 = ~n3350 & ~n3351;
  assign n3353 = pi72  & n2053;
  assign n3354 = pi73  & n1893;
  assign n3355 = pi74  & n1888;
  assign n3356 = n689 & n1886;
  assign n3357 = ~n3354 & ~n3355;
  assign n3358 = ~n3353 & n3357;
  assign n3359 = ~n3356 & n3358;
  assign n3360 = pi23  & n3359;
  assign n3361 = ~pi23  & ~n3359;
  assign n3362 = ~n3360 & ~n3361;
  assign n3363 = n3352 & ~n3362;
  assign n3364 = ~n3352 & n3362;
  assign n3365 = ~n3363 & ~n3364;
  assign n3366 = n3300 & ~n3365;
  assign n3367 = ~n3300 & n3365;
  assign n3368 = ~n3366 & ~n3367;
  assign n3369 = pi75  & n1661;
  assign n3370 = pi76  & n1500;
  assign n3371 = pi77  & n1495;
  assign n3372 = n865 & n1493;
  assign n3373 = ~n3370 & ~n3371;
  assign n3374 = ~n3369 & n3373;
  assign n3375 = ~n3372 & n3374;
  assign n3376 = pi20  & n3375;
  assign n3377 = ~pi20  & ~n3375;
  assign n3378 = ~n3376 & ~n3377;
  assign n3379 = ~n3368 & n3378;
  assign n3380 = n3368 & ~n3378;
  assign n3381 = ~n3379 & ~n3380;
  assign n3382 = ~n3196 & ~n3198;
  assign n3383 = n3381 & ~n3382;
  assign n3384 = ~n3381 & n3382;
  assign n3385 = ~n3383 & ~n3384;
  assign n3386 = pi78  & n1296;
  assign n3387 = pi79  & n1207;
  assign n3388 = pi80  & n1202;
  assign n3389 = n1144 & n1200;
  assign n3390 = ~n3387 & ~n3388;
  assign n3391 = ~n3386 & n3390;
  assign n3392 = ~n3389 & n3391;
  assign n3393 = pi17  & n3392;
  assign n3394 = ~pi17  & ~n3392;
  assign n3395 = ~n3393 & ~n3394;
  assign n3396 = n3385 & ~n3395;
  assign n3397 = ~n3385 & n3395;
  assign n3398 = ~n3396 & ~n3397;
  assign n3399 = n3299 & ~n3398;
  assign n3400 = ~n3299 & n3398;
  assign n3401 = ~n3399 & ~n3400;
  assign n3402 = pi81  & n1006;
  assign n3403 = pi82  & n897;
  assign n3404 = pi83  & n892;
  assign n3405 = n890 & n1577;
  assign n3406 = ~n3403 & ~n3404;
  assign n3407 = ~n3402 & n3406;
  assign n3408 = ~n3405 & n3407;
  assign n3409 = pi14  & n3408;
  assign n3410 = ~pi14  & ~n3408;
  assign n3411 = ~n3409 & ~n3410;
  assign n3412 = n3401 & ~n3411;
  assign n3413 = ~n3401 & n3411;
  assign n3414 = ~n3412 & ~n3413;
  assign n3415 = n3298 & ~n3414;
  assign n3416 = ~n3298 & n3414;
  assign n3417 = ~n3415 & ~n3416;
  assign n3418 = pi84  & n750;
  assign n3419 = pi85  & n651;
  assign n3420 = pi86  & n646;
  assign n3421 = n644 & n1975;
  assign n3422 = ~n3419 & ~n3420;
  assign n3423 = ~n3418 & n3422;
  assign n3424 = ~n3421 & n3423;
  assign n3425 = pi11  & n3424;
  assign n3426 = ~pi11  & ~n3424;
  assign n3427 = ~n3425 & ~n3426;
  assign n3428 = n3417 & ~n3427;
  assign n3429 = ~n3417 & n3427;
  assign n3430 = ~n3428 & ~n3429;
  assign n3431 = n3297 & ~n3430;
  assign n3432 = ~n3297 & n3430;
  assign n3433 = ~n3431 & ~n3432;
  assign n3434 = pi87  & n528;
  assign n3435 = pi88  & n490;
  assign n3436 = pi89  & n485;
  assign n3437 = n483 & n2287;
  assign n3438 = ~n3435 & ~n3436;
  assign n3439 = ~n3434 & n3438;
  assign n3440 = ~n3437 & n3439;
  assign n3441 = pi8  & n3440;
  assign n3442 = ~pi8  & ~n3440;
  assign n3443 = ~n3441 & ~n3442;
  assign n3444 = n3433 & ~n3443;
  assign n3445 = ~n3433 & n3443;
  assign n3446 = ~n3444 & ~n3445;
  assign n3447 = n3296 & ~n3446;
  assign n3448 = ~n3296 & n3446;
  assign n3449 = ~n3447 & ~n3448;
  assign n3450 = pi90  & n391;
  assign n3451 = pi91  & n353;
  assign n3452 = pi92  & n348;
  assign n3453 = n346 & n2924;
  assign n3454 = ~n3451 & ~n3452;
  assign n3455 = ~n3450 & n3454;
  assign n3456 = ~n3453 & n3455;
  assign n3457 = pi5  & n3456;
  assign n3458 = ~pi5  & ~n3456;
  assign n3459 = ~n3457 & ~n3458;
  assign n3460 = n3449 & ~n3459;
  assign n3461 = ~n3449 & n3459;
  assign n3462 = ~n3460 & ~n3461;
  assign n3463 = n3295 & ~n3462;
  assign n3464 = ~n3295 & n3462;
  assign n3465 = ~n3463 & ~n3464;
  assign n3466 = pi95  & n269;
  assign n3467 = pi94  & n267;
  assign n3468 = pi93  & n282;
  assign n3469 = ~n3276 & ~n3278;
  assign n3470 = ~pi94  & ~pi95 ;
  assign n3471 = pi94  & pi95 ;
  assign n3472 = ~n3470 & ~n3471;
  assign n3473 = ~n3469 & n3472;
  assign n3474 = n3469 & ~n3472;
  assign n3475 = ~n3473 & ~n3474;
  assign n3476 = n262 & n3475;
  assign n3477 = ~n3466 & ~n3467;
  assign n3478 = ~n3468 & n3477;
  assign n3479 = ~n3476 & n3478;
  assign n3480 = pi2  & n3479;
  assign n3481 = ~pi2  & ~n3479;
  assign n3482 = ~n3480 & ~n3481;
  assign n3483 = n3465 & ~n3482;
  assign n3484 = ~n3465 & n3482;
  assign n3485 = ~n3483 & ~n3484;
  assign n3486 = ~n3294 & n3485;
  assign n3487 = n3294 & ~n3485;
  assign po31  = ~n3486 & ~n3487;
  assign n3489 = ~n3483 & ~n3486;
  assign n3490 = pi96  & n269;
  assign n3491 = pi95  & n267;
  assign n3492 = pi94  & n282;
  assign n3493 = ~n3471 & ~n3473;
  assign n3494 = ~pi95  & ~pi96 ;
  assign n3495 = pi95  & pi96 ;
  assign n3496 = ~n3494 & ~n3495;
  assign n3497 = ~n3493 & n3496;
  assign n3498 = n3493 & ~n3496;
  assign n3499 = ~n3497 & ~n3498;
  assign n3500 = n262 & n3499;
  assign n3501 = ~n3490 & ~n3491;
  assign n3502 = ~n3492 & n3501;
  assign n3503 = ~n3500 & n3502;
  assign n3504 = pi2  & n3503;
  assign n3505 = ~pi2  & ~n3503;
  assign n3506 = ~n3504 & ~n3505;
  assign n3507 = ~n3460 & ~n3464;
  assign n3508 = ~n3444 & ~n3448;
  assign n3509 = ~n3428 & ~n3432;
  assign n3510 = pi85  & n750;
  assign n3511 = pi86  & n651;
  assign n3512 = pi87  & n646;
  assign n3513 = n644 & n2116;
  assign n3514 = ~n3511 & ~n3512;
  assign n3515 = ~n3510 & n3514;
  assign n3516 = ~n3513 & n3515;
  assign n3517 = pi11  & n3516;
  assign n3518 = ~pi11  & ~n3516;
  assign n3519 = ~n3517 & ~n3518;
  assign n3520 = ~n3412 & ~n3416;
  assign n3521 = ~n3396 & ~n3400;
  assign n3522 = ~n3380 & ~n3383;
  assign n3523 = pi76  & n1661;
  assign n3524 = pi77  & n1500;
  assign n3525 = pi78  & n1495;
  assign n3526 = n958 & n1493;
  assign n3527 = ~n3524 & ~n3525;
  assign n3528 = ~n3523 & n3527;
  assign n3529 = ~n3526 & n3528;
  assign n3530 = pi20  & n3529;
  assign n3531 = ~pi20  & ~n3529;
  assign n3532 = ~n3530 & ~n3531;
  assign n3533 = ~n3363 & ~n3367;
  assign n3534 = ~n3347 & ~n3350;
  assign n3535 = ~n3341 & ~n3344;
  assign n3536 = pi67  & n3011;
  assign n3537 = pi68  & n2809;
  assign n3538 = pi69  & n2804;
  assign n3539 = n376 & n2802;
  assign n3540 = ~n3537 & ~n3538;
  assign n3541 = ~n3536 & n3540;
  assign n3542 = ~n3539 & n3541;
  assign n3543 = pi29  & n3542;
  assign n3544 = ~pi29  & ~n3542;
  assign n3545 = ~n3543 & ~n3544;
  assign n3546 = pi32  & ~n3165;
  assign n3547 = n3337 & n3546;
  assign n3548 = pi32  & ~n3547;
  assign n3549 = ~n287 & n3327;
  assign n3550 = pi65  & n3334;
  assign n3551 = pi66  & n3329;
  assign n3552 = ~n3164 & n3326;
  assign n3553 = ~n3333 & n3552;
  assign n3554 = pi64  & n3553;
  assign n3555 = ~n3549 & ~n3550;
  assign n3556 = ~n3551 & n3555;
  assign n3557 = ~n3554 & n3556;
  assign n3558 = ~n3548 & n3557;
  assign n3559 = n3548 & ~n3557;
  assign n3560 = ~n3558 & ~n3559;
  assign n3561 = ~n3545 & n3560;
  assign n3562 = n3545 & ~n3560;
  assign n3563 = ~n3561 & ~n3562;
  assign n3564 = ~n3535 & n3563;
  assign n3565 = n3535 & ~n3563;
  assign n3566 = ~n3564 & ~n3565;
  assign n3567 = pi70  & n2510;
  assign n3568 = pi71  & n2342;
  assign n3569 = pi72  & n2337;
  assign n3570 = n551 & n2335;
  assign n3571 = ~n3568 & ~n3569;
  assign n3572 = ~n3567 & n3571;
  assign n3573 = ~n3570 & n3572;
  assign n3574 = pi26  & n3573;
  assign n3575 = ~pi26  & ~n3573;
  assign n3576 = ~n3574 & ~n3575;
  assign n3577 = n3566 & ~n3576;
  assign n3578 = ~n3566 & n3576;
  assign n3579 = ~n3577 & ~n3578;
  assign n3580 = n3534 & ~n3579;
  assign n3581 = ~n3534 & n3579;
  assign n3582 = ~n3580 & ~n3581;
  assign n3583 = pi73  & n2053;
  assign n3584 = pi74  & n1893;
  assign n3585 = pi75  & n1888;
  assign n3586 = n713 & n1886;
  assign n3587 = ~n3584 & ~n3585;
  assign n3588 = ~n3583 & n3587;
  assign n3589 = ~n3586 & n3588;
  assign n3590 = pi23  & n3589;
  assign n3591 = ~pi23  & ~n3589;
  assign n3592 = ~n3590 & ~n3591;
  assign n3593 = n3582 & ~n3592;
  assign n3594 = ~n3582 & n3592;
  assign n3595 = ~n3593 & ~n3594;
  assign n3596 = ~n3533 & n3595;
  assign n3597 = n3533 & ~n3595;
  assign n3598 = ~n3596 & ~n3597;
  assign n3599 = n3532 & ~n3598;
  assign n3600 = ~n3532 & n3598;
  assign n3601 = ~n3599 & ~n3600;
  assign n3602 = ~n3522 & n3601;
  assign n3603 = n3522 & ~n3601;
  assign n3604 = ~n3602 & ~n3603;
  assign n3605 = pi79  & n1296;
  assign n3606 = pi80  & n1207;
  assign n3607 = pi81  & n1202;
  assign n3608 = n1200 & n1337;
  assign n3609 = ~n3606 & ~n3607;
  assign n3610 = ~n3605 & n3609;
  assign n3611 = ~n3608 & n3610;
  assign n3612 = pi17  & n3611;
  assign n3613 = ~pi17  & ~n3611;
  assign n3614 = ~n3612 & ~n3613;
  assign n3615 = n3604 & ~n3614;
  assign n3616 = ~n3604 & n3614;
  assign n3617 = ~n3615 & ~n3616;
  assign n3618 = n3521 & ~n3617;
  assign n3619 = ~n3521 & n3617;
  assign n3620 = ~n3618 & ~n3619;
  assign n3621 = pi82  & n1006;
  assign n3622 = pi83  & n897;
  assign n3623 = pi84  & n892;
  assign n3624 = n890 & n1601;
  assign n3625 = ~n3622 & ~n3623;
  assign n3626 = ~n3621 & n3625;
  assign n3627 = ~n3624 & n3626;
  assign n3628 = pi14  & n3627;
  assign n3629 = ~pi14  & ~n3627;
  assign n3630 = ~n3628 & ~n3629;
  assign n3631 = n3620 & ~n3630;
  assign n3632 = ~n3620 & n3630;
  assign n3633 = ~n3631 & ~n3632;
  assign n3634 = ~n3520 & n3633;
  assign n3635 = n3520 & ~n3633;
  assign n3636 = ~n3634 & ~n3635;
  assign n3637 = n3519 & ~n3636;
  assign n3638 = ~n3519 & n3636;
  assign n3639 = ~n3637 & ~n3638;
  assign n3640 = ~n3509 & n3639;
  assign n3641 = n3509 & ~n3639;
  assign n3642 = ~n3640 & ~n3641;
  assign n3643 = pi88  & n528;
  assign n3644 = pi89  & n490;
  assign n3645 = pi90  & n485;
  assign n3646 = n483 & n2448;
  assign n3647 = ~n3644 & ~n3645;
  assign n3648 = ~n3643 & n3647;
  assign n3649 = ~n3646 & n3648;
  assign n3650 = pi8  & n3649;
  assign n3651 = ~pi8  & ~n3649;
  assign n3652 = ~n3650 & ~n3651;
  assign n3653 = n3642 & ~n3652;
  assign n3654 = ~n3642 & n3652;
  assign n3655 = ~n3653 & ~n3654;
  assign n3656 = n3508 & ~n3655;
  assign n3657 = ~n3508 & n3655;
  assign n3658 = ~n3656 & ~n3657;
  assign n3659 = pi91  & n391;
  assign n3660 = pi92  & n353;
  assign n3661 = pi93  & n348;
  assign n3662 = n346 & n2948;
  assign n3663 = ~n3660 & ~n3661;
  assign n3664 = ~n3659 & n3663;
  assign n3665 = ~n3662 & n3664;
  assign n3666 = pi5  & n3665;
  assign n3667 = ~pi5  & ~n3665;
  assign n3668 = ~n3666 & ~n3667;
  assign n3669 = n3658 & ~n3668;
  assign n3670 = ~n3658 & n3668;
  assign n3671 = ~n3669 & ~n3670;
  assign n3672 = ~n3507 & n3671;
  assign n3673 = n3507 & ~n3671;
  assign n3674 = ~n3672 & ~n3673;
  assign n3675 = ~n3506 & n3674;
  assign n3676 = n3506 & ~n3674;
  assign n3677 = ~n3675 & ~n3676;
  assign n3678 = ~n3489 & n3677;
  assign n3679 = n3489 & ~n3677;
  assign po32  = ~n3678 & ~n3679;
  assign n3681 = ~n3675 & ~n3678;
  assign n3682 = pi97  & n269;
  assign n3683 = pi96  & n267;
  assign n3684 = pi95  & n282;
  assign n3685 = ~n3495 & ~n3497;
  assign n3686 = ~pi96  & ~pi97 ;
  assign n3687 = pi96  & pi97 ;
  assign n3688 = ~n3686 & ~n3687;
  assign n3689 = ~n3685 & n3688;
  assign n3690 = n3685 & ~n3688;
  assign n3691 = ~n3689 & ~n3690;
  assign n3692 = n262 & n3691;
  assign n3693 = ~n3682 & ~n3683;
  assign n3694 = ~n3684 & n3693;
  assign n3695 = ~n3692 & n3694;
  assign n3696 = pi2  & n3695;
  assign n3697 = ~pi2  & ~n3695;
  assign n3698 = ~n3696 & ~n3697;
  assign n3699 = ~n3669 & ~n3672;
  assign n3700 = ~n3653 & ~n3657;
  assign n3701 = ~n3638 & ~n3640;
  assign n3702 = pi86  & n750;
  assign n3703 = pi87  & n651;
  assign n3704 = pi88  & n646;
  assign n3705 = n644 & n2140;
  assign n3706 = ~n3703 & ~n3704;
  assign n3707 = ~n3702 & n3706;
  assign n3708 = ~n3705 & n3707;
  assign n3709 = pi11  & n3708;
  assign n3710 = ~pi11  & ~n3708;
  assign n3711 = ~n3709 & ~n3710;
  assign n3712 = ~n3631 & ~n3634;
  assign n3713 = ~n3615 & ~n3619;
  assign n3714 = pi80  & n1296;
  assign n3715 = pi81  & n1207;
  assign n3716 = pi82  & n1202;
  assign n3717 = n1200 & n1450;
  assign n3718 = ~n3715 & ~n3716;
  assign n3719 = ~n3714 & n3718;
  assign n3720 = ~n3717 & n3719;
  assign n3721 = pi17  & n3720;
  assign n3722 = ~pi17  & ~n3720;
  assign n3723 = ~n3721 & ~n3722;
  assign n3724 = ~n3600 & ~n3602;
  assign n3725 = ~n3593 & ~n3596;
  assign n3726 = ~n3577 & ~n3581;
  assign n3727 = pi71  & n2510;
  assign n3728 = pi72  & n2342;
  assign n3729 = pi73  & n2337;
  assign n3730 = n613 & n2335;
  assign n3731 = ~n3728 & ~n3729;
  assign n3732 = ~n3727 & n3731;
  assign n3733 = ~n3730 & n3732;
  assign n3734 = pi26  & n3733;
  assign n3735 = ~pi26  & ~n3733;
  assign n3736 = ~n3734 & ~n3735;
  assign n3737 = ~n3561 & ~n3564;
  assign n3738 = pi65  & n3553;
  assign n3739 = pi66  & n3334;
  assign n3740 = pi67  & n3329;
  assign n3741 = n305 & n3327;
  assign n3742 = ~n3739 & ~n3740;
  assign n3743 = ~n3738 & n3742;
  assign n3744 = ~n3741 & n3743;
  assign n3745 = pi32  & n3744;
  assign n3746 = ~pi32  & ~n3744;
  assign n3747 = ~n3745 & ~n3746;
  assign n3748 = ~pi32  & ~pi33 ;
  assign n3749 = pi32  & pi33 ;
  assign n3750 = ~n3748 & ~n3749;
  assign n3751 = pi64  & n3750;
  assign n3752 = n3547 & n3557;
  assign n3753 = n3751 & n3752;
  assign n3754 = ~n3751 & ~n3752;
  assign n3755 = ~n3753 & ~n3754;
  assign n3756 = ~n3747 & n3755;
  assign n3757 = n3747 & ~n3755;
  assign n3758 = ~n3756 & ~n3757;
  assign n3759 = pi68  & n3011;
  assign n3760 = pi69  & n2809;
  assign n3761 = pi70  & n2804;
  assign n3762 = n415 & n2802;
  assign n3763 = ~n3760 & ~n3761;
  assign n3764 = ~n3759 & n3763;
  assign n3765 = ~n3762 & n3764;
  assign n3766 = pi29  & n3765;
  assign n3767 = ~pi29  & ~n3765;
  assign n3768 = ~n3766 & ~n3767;
  assign n3769 = n3758 & ~n3768;
  assign n3770 = ~n3758 & n3768;
  assign n3771 = ~n3769 & ~n3770;
  assign n3772 = ~n3737 & n3771;
  assign n3773 = n3737 & ~n3771;
  assign n3774 = ~n3772 & ~n3773;
  assign n3775 = ~n3736 & n3774;
  assign n3776 = n3736 & ~n3774;
  assign n3777 = ~n3775 & ~n3776;
  assign n3778 = n3726 & ~n3777;
  assign n3779 = ~n3726 & n3777;
  assign n3780 = ~n3778 & ~n3779;
  assign n3781 = pi74  & n2053;
  assign n3782 = pi75  & n1893;
  assign n3783 = pi76  & n1888;
  assign n3784 = n841 & n1886;
  assign n3785 = ~n3782 & ~n3783;
  assign n3786 = ~n3781 & n3785;
  assign n3787 = ~n3784 & n3786;
  assign n3788 = pi23  & n3787;
  assign n3789 = ~pi23  & ~n3787;
  assign n3790 = ~n3788 & ~n3789;
  assign n3791 = ~n3780 & n3790;
  assign n3792 = n3780 & ~n3790;
  assign n3793 = ~n3791 & ~n3792;
  assign n3794 = ~n3725 & n3793;
  assign n3795 = n3725 & ~n3793;
  assign n3796 = ~n3794 & ~n3795;
  assign n3797 = pi77  & n1661;
  assign n3798 = pi78  & n1500;
  assign n3799 = pi79  & n1495;
  assign n3800 = n1048 & n1493;
  assign n3801 = ~n3798 & ~n3799;
  assign n3802 = ~n3797 & n3801;
  assign n3803 = ~n3800 & n3802;
  assign n3804 = pi20  & n3803;
  assign n3805 = ~pi20  & ~n3803;
  assign n3806 = ~n3804 & ~n3805;
  assign n3807 = n3796 & ~n3806;
  assign n3808 = ~n3796 & n3806;
  assign n3809 = ~n3807 & ~n3808;
  assign n3810 = ~n3724 & n3809;
  assign n3811 = n3724 & ~n3809;
  assign n3812 = ~n3810 & ~n3811;
  assign n3813 = ~n3723 & n3812;
  assign n3814 = n3723 & ~n3812;
  assign n3815 = ~n3813 & ~n3814;
  assign n3816 = n3713 & ~n3815;
  assign n3817 = ~n3713 & n3815;
  assign n3818 = ~n3816 & ~n3817;
  assign n3819 = pi83  & n1006;
  assign n3820 = pi84  & n897;
  assign n3821 = pi85  & n892;
  assign n3822 = n890 & n1831;
  assign n3823 = ~n3820 & ~n3821;
  assign n3824 = ~n3819 & n3823;
  assign n3825 = ~n3822 & n3824;
  assign n3826 = pi14  & n3825;
  assign n3827 = ~pi14  & ~n3825;
  assign n3828 = ~n3826 & ~n3827;
  assign n3829 = n3818 & ~n3828;
  assign n3830 = ~n3818 & n3828;
  assign n3831 = ~n3829 & ~n3830;
  assign n3832 = ~n3712 & n3831;
  assign n3833 = n3712 & ~n3831;
  assign n3834 = ~n3832 & ~n3833;
  assign n3835 = n3711 & ~n3834;
  assign n3836 = ~n3711 & n3834;
  assign n3837 = ~n3835 & ~n3836;
  assign n3838 = ~n3701 & n3837;
  assign n3839 = n3701 & ~n3837;
  assign n3840 = ~n3838 & ~n3839;
  assign n3841 = pi89  & n528;
  assign n3842 = pi90  & n490;
  assign n3843 = pi91  & n485;
  assign n3844 = n483 & n2746;
  assign n3845 = ~n3842 & ~n3843;
  assign n3846 = ~n3841 & n3845;
  assign n3847 = ~n3844 & n3846;
  assign n3848 = pi8  & n3847;
  assign n3849 = ~pi8  & ~n3847;
  assign n3850 = ~n3848 & ~n3849;
  assign n3851 = n3840 & ~n3850;
  assign n3852 = ~n3840 & n3850;
  assign n3853 = ~n3851 & ~n3852;
  assign n3854 = n3700 & ~n3853;
  assign n3855 = ~n3700 & n3853;
  assign n3856 = ~n3854 & ~n3855;
  assign n3857 = pi92  & n391;
  assign n3858 = pi93  & n353;
  assign n3859 = pi94  & n348;
  assign n3860 = n346 & n3280;
  assign n3861 = ~n3858 & ~n3859;
  assign n3862 = ~n3857 & n3861;
  assign n3863 = ~n3860 & n3862;
  assign n3864 = pi5  & n3863;
  assign n3865 = ~pi5  & ~n3863;
  assign n3866 = ~n3864 & ~n3865;
  assign n3867 = n3856 & ~n3866;
  assign n3868 = ~n3856 & n3866;
  assign n3869 = ~n3867 & ~n3868;
  assign n3870 = ~n3699 & n3869;
  assign n3871 = n3699 & ~n3869;
  assign n3872 = ~n3870 & ~n3871;
  assign n3873 = ~n3698 & n3872;
  assign n3874 = n3698 & ~n3872;
  assign n3875 = ~n3873 & ~n3874;
  assign n3876 = ~n3681 & n3875;
  assign n3877 = n3681 & ~n3875;
  assign po33  = ~n3876 & ~n3877;
  assign n3879 = ~n3873 & ~n3876;
  assign n3880 = pi98  & n269;
  assign n3881 = pi97  & n267;
  assign n3882 = pi96  & n282;
  assign n3883 = ~n3687 & ~n3689;
  assign n3884 = ~pi97  & ~pi98 ;
  assign n3885 = pi97  & pi98 ;
  assign n3886 = ~n3884 & ~n3885;
  assign n3887 = ~n3883 & n3886;
  assign n3888 = n3883 & ~n3886;
  assign n3889 = ~n3887 & ~n3888;
  assign n3890 = n262 & n3889;
  assign n3891 = ~n3880 & ~n3881;
  assign n3892 = ~n3882 & n3891;
  assign n3893 = ~n3890 & n3892;
  assign n3894 = pi2  & n3893;
  assign n3895 = ~pi2  & ~n3893;
  assign n3896 = ~n3894 & ~n3895;
  assign n3897 = ~n3867 & ~n3870;
  assign n3898 = ~n3851 & ~n3855;
  assign n3899 = ~n3836 & ~n3838;
  assign n3900 = ~n3829 & ~n3832;
  assign n3901 = ~n3813 & ~n3817;
  assign n3902 = ~n3807 & ~n3810;
  assign n3903 = ~n3792 & ~n3794;
  assign n3904 = ~n3775 & ~n3779;
  assign n3905 = ~n3769 & ~n3772;
  assign n3906 = pi69  & n3011;
  assign n3907 = pi70  & n2809;
  assign n3908 = pi71  & n2804;
  assign n3909 = n460 & n2802;
  assign n3910 = ~n3907 & ~n3908;
  assign n3911 = ~n3906 & n3910;
  assign n3912 = ~n3909 & n3911;
  assign n3913 = pi29  & n3912;
  assign n3914 = ~pi29  & ~n3912;
  assign n3915 = ~n3913 & ~n3914;
  assign n3916 = ~n3753 & ~n3756;
  assign n3917 = pi66  & n3553;
  assign n3918 = pi67  & n3334;
  assign n3919 = pi68  & n3329;
  assign n3920 = n334 & n3327;
  assign n3921 = ~n3918 & ~n3919;
  assign n3922 = ~n3917 & n3921;
  assign n3923 = ~n3920 & n3922;
  assign n3924 = pi32  & n3923;
  assign n3925 = ~pi32  & ~n3923;
  assign n3926 = ~n3924 & ~n3925;
  assign n3927 = pi35  & n3751;
  assign n3928 = ~pi34  & ~pi35 ;
  assign n3929 = pi34  & pi35 ;
  assign n3930 = ~n3928 & ~n3929;
  assign n3931 = n3750 & n3930;
  assign n3932 = n265 & n3931;
  assign n3933 = n3750 & ~n3930;
  assign n3934 = pi65  & n3933;
  assign n3935 = ~pi33  & ~pi34 ;
  assign n3936 = pi33  & pi34 ;
  assign n3937 = ~n3935 & ~n3936;
  assign n3938 = ~n3750 & n3937;
  assign n3939 = pi64  & n3938;
  assign n3940 = ~n3932 & ~n3934;
  assign n3941 = ~n3939 & n3940;
  assign n3942 = n3927 & ~n3941;
  assign n3943 = ~n3927 & n3941;
  assign n3944 = ~n3942 & ~n3943;
  assign n3945 = n3926 & ~n3944;
  assign n3946 = ~n3926 & n3944;
  assign n3947 = ~n3945 & ~n3946;
  assign n3948 = ~n3916 & n3947;
  assign n3949 = n3916 & ~n3947;
  assign n3950 = ~n3948 & ~n3949;
  assign n3951 = n3915 & ~n3950;
  assign n3952 = ~n3915 & n3950;
  assign n3953 = ~n3951 & ~n3952;
  assign n3954 = ~n3905 & n3953;
  assign n3955 = n3905 & ~n3953;
  assign n3956 = ~n3954 & ~n3955;
  assign n3957 = pi72  & n2510;
  assign n3958 = pi73  & n2342;
  assign n3959 = pi74  & n2337;
  assign n3960 = n689 & n2335;
  assign n3961 = ~n3958 & ~n3959;
  assign n3962 = ~n3957 & n3961;
  assign n3963 = ~n3960 & n3962;
  assign n3964 = pi26  & n3963;
  assign n3965 = ~pi26  & ~n3963;
  assign n3966 = ~n3964 & ~n3965;
  assign n3967 = n3956 & ~n3966;
  assign n3968 = ~n3956 & n3966;
  assign n3969 = ~n3967 & ~n3968;
  assign n3970 = n3904 & ~n3969;
  assign n3971 = ~n3904 & n3969;
  assign n3972 = ~n3970 & ~n3971;
  assign n3973 = pi75  & n2053;
  assign n3974 = pi76  & n1893;
  assign n3975 = pi77  & n1888;
  assign n3976 = n865 & n1886;
  assign n3977 = ~n3974 & ~n3975;
  assign n3978 = ~n3973 & n3977;
  assign n3979 = ~n3976 & n3978;
  assign n3980 = pi23  & n3979;
  assign n3981 = ~pi23  & ~n3979;
  assign n3982 = ~n3980 & ~n3981;
  assign n3983 = n3972 & ~n3982;
  assign n3984 = ~n3972 & n3982;
  assign n3985 = ~n3983 & ~n3984;
  assign n3986 = ~n3903 & n3985;
  assign n3987 = n3903 & ~n3985;
  assign n3988 = ~n3986 & ~n3987;
  assign n3989 = pi78  & n1661;
  assign n3990 = pi79  & n1500;
  assign n3991 = pi80  & n1495;
  assign n3992 = n1144 & n1493;
  assign n3993 = ~n3990 & ~n3991;
  assign n3994 = ~n3989 & n3993;
  assign n3995 = ~n3992 & n3994;
  assign n3996 = pi20  & n3995;
  assign n3997 = ~pi20  & ~n3995;
  assign n3998 = ~n3996 & ~n3997;
  assign n3999 = n3988 & ~n3998;
  assign n4000 = ~n3988 & n3998;
  assign n4001 = ~n3999 & ~n4000;
  assign n4002 = n3902 & ~n4001;
  assign n4003 = ~n3902 & n4001;
  assign n4004 = ~n4002 & ~n4003;
  assign n4005 = pi81  & n1296;
  assign n4006 = pi82  & n1207;
  assign n4007 = pi83  & n1202;
  assign n4008 = n1200 & n1577;
  assign n4009 = ~n4006 & ~n4007;
  assign n4010 = ~n4005 & n4009;
  assign n4011 = ~n4008 & n4010;
  assign n4012 = pi17  & n4011;
  assign n4013 = ~pi17  & ~n4011;
  assign n4014 = ~n4012 & ~n4013;
  assign n4015 = n4004 & ~n4014;
  assign n4016 = ~n4004 & n4014;
  assign n4017 = ~n4015 & ~n4016;
  assign n4018 = n3901 & ~n4017;
  assign n4019 = ~n3901 & n4017;
  assign n4020 = ~n4018 & ~n4019;
  assign n4021 = pi84  & n1006;
  assign n4022 = pi85  & n897;
  assign n4023 = pi86  & n892;
  assign n4024 = n890 & n1975;
  assign n4025 = ~n4022 & ~n4023;
  assign n4026 = ~n4021 & n4025;
  assign n4027 = ~n4024 & n4026;
  assign n4028 = pi14  & n4027;
  assign n4029 = ~pi14  & ~n4027;
  assign n4030 = ~n4028 & ~n4029;
  assign n4031 = n4020 & ~n4030;
  assign n4032 = ~n4020 & n4030;
  assign n4033 = ~n4031 & ~n4032;
  assign n4034 = n3900 & ~n4033;
  assign n4035 = ~n3900 & n4033;
  assign n4036 = ~n4034 & ~n4035;
  assign n4037 = pi87  & n750;
  assign n4038 = pi88  & n651;
  assign n4039 = pi89  & n646;
  assign n4040 = n644 & n2287;
  assign n4041 = ~n4038 & ~n4039;
  assign n4042 = ~n4037 & n4041;
  assign n4043 = ~n4040 & n4042;
  assign n4044 = pi11  & n4043;
  assign n4045 = ~pi11  & ~n4043;
  assign n4046 = ~n4044 & ~n4045;
  assign n4047 = n4036 & ~n4046;
  assign n4048 = ~n4036 & n4046;
  assign n4049 = ~n4047 & ~n4048;
  assign n4050 = ~n3899 & n4049;
  assign n4051 = n3899 & ~n4049;
  assign n4052 = ~n4050 & ~n4051;
  assign n4053 = pi90  & n528;
  assign n4054 = pi91  & n490;
  assign n4055 = pi92  & n485;
  assign n4056 = n483 & n2924;
  assign n4057 = ~n4054 & ~n4055;
  assign n4058 = ~n4053 & n4057;
  assign n4059 = ~n4056 & n4058;
  assign n4060 = pi8  & n4059;
  assign n4061 = ~pi8  & ~n4059;
  assign n4062 = ~n4060 & ~n4061;
  assign n4063 = n4052 & ~n4062;
  assign n4064 = ~n4052 & n4062;
  assign n4065 = ~n4063 & ~n4064;
  assign n4066 = n3898 & ~n4065;
  assign n4067 = ~n3898 & n4065;
  assign n4068 = ~n4066 & ~n4067;
  assign n4069 = pi93  & n391;
  assign n4070 = pi94  & n353;
  assign n4071 = pi95  & n348;
  assign n4072 = n346 & n3475;
  assign n4073 = ~n4070 & ~n4071;
  assign n4074 = ~n4069 & n4073;
  assign n4075 = ~n4072 & n4074;
  assign n4076 = pi5  & n4075;
  assign n4077 = ~pi5  & ~n4075;
  assign n4078 = ~n4076 & ~n4077;
  assign n4079 = n4068 & ~n4078;
  assign n4080 = ~n4068 & n4078;
  assign n4081 = ~n4079 & ~n4080;
  assign n4082 = ~n3897 & n4081;
  assign n4083 = n3897 & ~n4081;
  assign n4084 = ~n4082 & ~n4083;
  assign n4085 = ~n3896 & n4084;
  assign n4086 = n3896 & ~n4084;
  assign n4087 = ~n4085 & ~n4086;
  assign n4088 = ~n3879 & n4087;
  assign n4089 = n3879 & ~n4087;
  assign po34  = ~n4088 & ~n4089;
  assign n4091 = ~n4085 & ~n4088;
  assign n4092 = pi99  & n269;
  assign n4093 = pi98  & n267;
  assign n4094 = pi97  & n282;
  assign n4095 = ~n3885 & ~n3887;
  assign n4096 = ~pi98  & ~pi99 ;
  assign n4097 = pi98  & pi99 ;
  assign n4098 = ~n4096 & ~n4097;
  assign n4099 = ~n4095 & n4098;
  assign n4100 = n4095 & ~n4098;
  assign n4101 = ~n4099 & ~n4100;
  assign n4102 = n262 & n4101;
  assign n4103 = ~n4092 & ~n4093;
  assign n4104 = ~n4094 & n4103;
  assign n4105 = ~n4102 & n4104;
  assign n4106 = pi2  & n4105;
  assign n4107 = ~pi2  & ~n4105;
  assign n4108 = ~n4106 & ~n4107;
  assign n4109 = ~n4079 & ~n4082;
  assign n4110 = ~n4063 & ~n4067;
  assign n4111 = ~n4047 & ~n4050;
  assign n4112 = pi88  & n750;
  assign n4113 = pi89  & n651;
  assign n4114 = pi90  & n646;
  assign n4115 = n644 & n2448;
  assign n4116 = ~n4113 & ~n4114;
  assign n4117 = ~n4112 & n4116;
  assign n4118 = ~n4115 & n4117;
  assign n4119 = pi11  & n4118;
  assign n4120 = ~pi11  & ~n4118;
  assign n4121 = ~n4119 & ~n4120;
  assign n4122 = ~n4031 & ~n4035;
  assign n4123 = pi85  & n1006;
  assign n4124 = pi86  & n897;
  assign n4125 = pi87  & n892;
  assign n4126 = n890 & n2116;
  assign n4127 = ~n4124 & ~n4125;
  assign n4128 = ~n4123 & n4127;
  assign n4129 = ~n4126 & n4128;
  assign n4130 = pi14  & n4129;
  assign n4131 = ~pi14  & ~n4129;
  assign n4132 = ~n4130 & ~n4131;
  assign n4133 = ~n4015 & ~n4019;
  assign n4134 = ~n3999 & ~n4003;
  assign n4135 = ~n3983 & ~n3986;
  assign n4136 = pi76  & n2053;
  assign n4137 = pi77  & n1893;
  assign n4138 = pi78  & n1888;
  assign n4139 = n958 & n1886;
  assign n4140 = ~n4137 & ~n4138;
  assign n4141 = ~n4136 & n4140;
  assign n4142 = ~n4139 & n4141;
  assign n4143 = pi23  & n4142;
  assign n4144 = ~pi23  & ~n4142;
  assign n4145 = ~n4143 & ~n4144;
  assign n4146 = ~n3967 & ~n3971;
  assign n4147 = pi73  & n2510;
  assign n4148 = pi74  & n2342;
  assign n4149 = pi75  & n2337;
  assign n4150 = n713 & n2335;
  assign n4151 = ~n4148 & ~n4149;
  assign n4152 = ~n4147 & n4151;
  assign n4153 = ~n4150 & n4152;
  assign n4154 = pi26  & n4153;
  assign n4155 = ~pi26  & ~n4153;
  assign n4156 = ~n4154 & ~n4155;
  assign n4157 = ~n3952 & ~n3954;
  assign n4158 = ~n3946 & ~n3948;
  assign n4159 = pi67  & n3553;
  assign n4160 = pi68  & n3334;
  assign n4161 = pi69  & n3329;
  assign n4162 = n376 & n3327;
  assign n4163 = ~n4160 & ~n4161;
  assign n4164 = ~n4159 & n4163;
  assign n4165 = ~n4162 & n4164;
  assign n4166 = pi32  & n4165;
  assign n4167 = ~pi32  & ~n4165;
  assign n4168 = ~n4166 & ~n4167;
  assign n4169 = pi35  & ~n3751;
  assign n4170 = n3941 & n4169;
  assign n4171 = pi35  & ~n4170;
  assign n4172 = ~n287 & n3931;
  assign n4173 = pi65  & n3938;
  assign n4174 = pi66  & n3933;
  assign n4175 = ~n3750 & n3930;
  assign n4176 = ~n3937 & n4175;
  assign n4177 = pi64  & n4176;
  assign n4178 = ~n4172 & ~n4173;
  assign n4179 = ~n4174 & n4178;
  assign n4180 = ~n4177 & n4179;
  assign n4181 = ~n4171 & n4180;
  assign n4182 = n4171 & ~n4180;
  assign n4183 = ~n4181 & ~n4182;
  assign n4184 = ~n4168 & n4183;
  assign n4185 = n4168 & ~n4183;
  assign n4186 = ~n4184 & ~n4185;
  assign n4187 = ~n4158 & n4186;
  assign n4188 = n4158 & ~n4186;
  assign n4189 = ~n4187 & ~n4188;
  assign n4190 = pi70  & n3011;
  assign n4191 = pi71  & n2809;
  assign n4192 = pi72  & n2804;
  assign n4193 = n551 & n2802;
  assign n4194 = ~n4191 & ~n4192;
  assign n4195 = ~n4190 & n4194;
  assign n4196 = ~n4193 & n4195;
  assign n4197 = pi29  & n4196;
  assign n4198 = ~pi29  & ~n4196;
  assign n4199 = ~n4197 & ~n4198;
  assign n4200 = n4189 & ~n4199;
  assign n4201 = ~n4189 & n4199;
  assign n4202 = ~n4200 & ~n4201;
  assign n4203 = ~n4157 & n4202;
  assign n4204 = n4157 & ~n4202;
  assign n4205 = ~n4203 & ~n4204;
  assign n4206 = ~n4156 & n4205;
  assign n4207 = n4156 & ~n4205;
  assign n4208 = ~n4206 & ~n4207;
  assign n4209 = ~n4146 & n4208;
  assign n4210 = n4146 & ~n4208;
  assign n4211 = ~n4209 & ~n4210;
  assign n4212 = n4145 & ~n4211;
  assign n4213 = ~n4145 & n4211;
  assign n4214 = ~n4212 & ~n4213;
  assign n4215 = ~n4135 & n4214;
  assign n4216 = n4135 & ~n4214;
  assign n4217 = ~n4215 & ~n4216;
  assign n4218 = pi79  & n1661;
  assign n4219 = pi80  & n1500;
  assign n4220 = pi81  & n1495;
  assign n4221 = n1337 & n1493;
  assign n4222 = ~n4219 & ~n4220;
  assign n4223 = ~n4218 & n4222;
  assign n4224 = ~n4221 & n4223;
  assign n4225 = pi20  & n4224;
  assign n4226 = ~pi20  & ~n4224;
  assign n4227 = ~n4225 & ~n4226;
  assign n4228 = n4217 & ~n4227;
  assign n4229 = ~n4217 & n4227;
  assign n4230 = ~n4228 & ~n4229;
  assign n4231 = n4134 & ~n4230;
  assign n4232 = ~n4134 & n4230;
  assign n4233 = ~n4231 & ~n4232;
  assign n4234 = pi82  & n1296;
  assign n4235 = pi83  & n1207;
  assign n4236 = pi84  & n1202;
  assign n4237 = n1200 & n1601;
  assign n4238 = ~n4235 & ~n4236;
  assign n4239 = ~n4234 & n4238;
  assign n4240 = ~n4237 & n4239;
  assign n4241 = pi17  & n4240;
  assign n4242 = ~pi17  & ~n4240;
  assign n4243 = ~n4241 & ~n4242;
  assign n4244 = n4233 & ~n4243;
  assign n4245 = ~n4233 & n4243;
  assign n4246 = ~n4244 & ~n4245;
  assign n4247 = ~n4133 & n4246;
  assign n4248 = n4133 & ~n4246;
  assign n4249 = ~n4247 & ~n4248;
  assign n4250 = n4132 & ~n4249;
  assign n4251 = ~n4132 & n4249;
  assign n4252 = ~n4250 & ~n4251;
  assign n4253 = ~n4122 & n4252;
  assign n4254 = n4122 & ~n4252;
  assign n4255 = ~n4253 & ~n4254;
  assign n4256 = n4121 & ~n4255;
  assign n4257 = ~n4121 & n4255;
  assign n4258 = ~n4256 & ~n4257;
  assign n4259 = ~n4111 & n4258;
  assign n4260 = n4111 & ~n4258;
  assign n4261 = ~n4259 & ~n4260;
  assign n4262 = pi91  & n528;
  assign n4263 = pi92  & n490;
  assign n4264 = pi93  & n485;
  assign n4265 = n483 & n2948;
  assign n4266 = ~n4263 & ~n4264;
  assign n4267 = ~n4262 & n4266;
  assign n4268 = ~n4265 & n4267;
  assign n4269 = pi8  & n4268;
  assign n4270 = ~pi8  & ~n4268;
  assign n4271 = ~n4269 & ~n4270;
  assign n4272 = n4261 & ~n4271;
  assign n4273 = ~n4261 & n4271;
  assign n4274 = ~n4272 & ~n4273;
  assign n4275 = n4110 & ~n4274;
  assign n4276 = ~n4110 & n4274;
  assign n4277 = ~n4275 & ~n4276;
  assign n4278 = pi94  & n391;
  assign n4279 = pi95  & n353;
  assign n4280 = pi96  & n348;
  assign n4281 = n346 & n3499;
  assign n4282 = ~n4279 & ~n4280;
  assign n4283 = ~n4278 & n4282;
  assign n4284 = ~n4281 & n4283;
  assign n4285 = pi5  & n4284;
  assign n4286 = ~pi5  & ~n4284;
  assign n4287 = ~n4285 & ~n4286;
  assign n4288 = n4277 & ~n4287;
  assign n4289 = ~n4277 & n4287;
  assign n4290 = ~n4288 & ~n4289;
  assign n4291 = ~n4109 & n4290;
  assign n4292 = n4109 & ~n4290;
  assign n4293 = ~n4291 & ~n4292;
  assign n4294 = ~n4108 & n4293;
  assign n4295 = n4108 & ~n4293;
  assign n4296 = ~n4294 & ~n4295;
  assign n4297 = ~n4091 & n4296;
  assign n4298 = n4091 & ~n4296;
  assign po35  = ~n4297 & ~n4298;
  assign n4300 = ~n4294 & ~n4297;
  assign n4301 = ~n4288 & ~n4291;
  assign n4302 = pi95  & n391;
  assign n4303 = pi96  & n353;
  assign n4304 = pi97  & n348;
  assign n4305 = n346 & n3691;
  assign n4306 = ~n4303 & ~n4304;
  assign n4307 = ~n4302 & n4306;
  assign n4308 = ~n4305 & n4307;
  assign n4309 = pi5  & n4308;
  assign n4310 = ~pi5  & ~n4308;
  assign n4311 = ~n4309 & ~n4310;
  assign n4312 = ~n4272 & ~n4276;
  assign n4313 = pi92  & n528;
  assign n4314 = pi93  & n490;
  assign n4315 = pi94  & n485;
  assign n4316 = n483 & n3280;
  assign n4317 = ~n4314 & ~n4315;
  assign n4318 = ~n4313 & n4317;
  assign n4319 = ~n4316 & n4318;
  assign n4320 = pi8  & n4319;
  assign n4321 = ~pi8  & ~n4319;
  assign n4322 = ~n4320 & ~n4321;
  assign n4323 = ~n4257 & ~n4259;
  assign n4324 = ~n4251 & ~n4253;
  assign n4325 = pi86  & n1006;
  assign n4326 = pi87  & n897;
  assign n4327 = pi88  & n892;
  assign n4328 = n890 & n2140;
  assign n4329 = ~n4326 & ~n4327;
  assign n4330 = ~n4325 & n4329;
  assign n4331 = ~n4328 & n4330;
  assign n4332 = pi14  & n4331;
  assign n4333 = ~pi14  & ~n4331;
  assign n4334 = ~n4332 & ~n4333;
  assign n4335 = ~n4244 & ~n4247;
  assign n4336 = ~n4228 & ~n4232;
  assign n4337 = pi80  & n1661;
  assign n4338 = pi81  & n1500;
  assign n4339 = pi82  & n1495;
  assign n4340 = n1450 & n1493;
  assign n4341 = ~n4338 & ~n4339;
  assign n4342 = ~n4337 & n4341;
  assign n4343 = ~n4340 & n4342;
  assign n4344 = pi20  & n4343;
  assign n4345 = ~pi20  & ~n4343;
  assign n4346 = ~n4344 & ~n4345;
  assign n4347 = ~n4213 & ~n4215;
  assign n4348 = ~n4200 & ~n4203;
  assign n4349 = pi71  & n3011;
  assign n4350 = pi72  & n2809;
  assign n4351 = pi73  & n2804;
  assign n4352 = n613 & n2802;
  assign n4353 = ~n4350 & ~n4351;
  assign n4354 = ~n4349 & n4353;
  assign n4355 = ~n4352 & n4354;
  assign n4356 = pi29  & n4355;
  assign n4357 = ~pi29  & ~n4355;
  assign n4358 = ~n4356 & ~n4357;
  assign n4359 = ~n4184 & ~n4187;
  assign n4360 = pi65  & n4176;
  assign n4361 = pi66  & n3938;
  assign n4362 = pi67  & n3933;
  assign n4363 = n305 & n3931;
  assign n4364 = ~n4361 & ~n4362;
  assign n4365 = ~n4360 & n4364;
  assign n4366 = ~n4363 & n4365;
  assign n4367 = pi35  & n4366;
  assign n4368 = ~pi35  & ~n4366;
  assign n4369 = ~n4367 & ~n4368;
  assign n4370 = ~pi35  & ~pi36 ;
  assign n4371 = pi35  & pi36 ;
  assign n4372 = ~n4370 & ~n4371;
  assign n4373 = pi64  & n4372;
  assign n4374 = n4170 & n4180;
  assign n4375 = n4373 & n4374;
  assign n4376 = ~n4373 & ~n4374;
  assign n4377 = ~n4375 & ~n4376;
  assign n4378 = ~n4369 & n4377;
  assign n4379 = n4369 & ~n4377;
  assign n4380 = ~n4378 & ~n4379;
  assign n4381 = pi68  & n3553;
  assign n4382 = pi69  & n3334;
  assign n4383 = pi70  & n3329;
  assign n4384 = n415 & n3327;
  assign n4385 = ~n4382 & ~n4383;
  assign n4386 = ~n4381 & n4385;
  assign n4387 = ~n4384 & n4386;
  assign n4388 = pi32  & n4387;
  assign n4389 = ~pi32  & ~n4387;
  assign n4390 = ~n4388 & ~n4389;
  assign n4391 = n4380 & ~n4390;
  assign n4392 = ~n4380 & n4390;
  assign n4393 = ~n4391 & ~n4392;
  assign n4394 = ~n4359 & n4393;
  assign n4395 = n4359 & ~n4393;
  assign n4396 = ~n4394 & ~n4395;
  assign n4397 = ~n4358 & n4396;
  assign n4398 = n4358 & ~n4396;
  assign n4399 = ~n4397 & ~n4398;
  assign n4400 = n4348 & ~n4399;
  assign n4401 = ~n4348 & n4399;
  assign n4402 = ~n4400 & ~n4401;
  assign n4403 = pi74  & n2510;
  assign n4404 = pi75  & n2342;
  assign n4405 = pi76  & n2337;
  assign n4406 = n841 & n2335;
  assign n4407 = ~n4404 & ~n4405;
  assign n4408 = ~n4403 & n4407;
  assign n4409 = ~n4406 & n4408;
  assign n4410 = pi26  & n4409;
  assign n4411 = ~pi26  & ~n4409;
  assign n4412 = ~n4410 & ~n4411;
  assign n4413 = ~n4402 & n4412;
  assign n4414 = n4402 & ~n4412;
  assign n4415 = ~n4413 & ~n4414;
  assign n4416 = ~n4206 & ~n4209;
  assign n4417 = n4415 & ~n4416;
  assign n4418 = ~n4415 & n4416;
  assign n4419 = ~n4417 & ~n4418;
  assign n4420 = pi77  & n2053;
  assign n4421 = pi78  & n1893;
  assign n4422 = pi79  & n1888;
  assign n4423 = n1048 & n1886;
  assign n4424 = ~n4421 & ~n4422;
  assign n4425 = ~n4420 & n4424;
  assign n4426 = ~n4423 & n4425;
  assign n4427 = pi23  & n4426;
  assign n4428 = ~pi23  & ~n4426;
  assign n4429 = ~n4427 & ~n4428;
  assign n4430 = n4419 & ~n4429;
  assign n4431 = ~n4419 & n4429;
  assign n4432 = ~n4430 & ~n4431;
  assign n4433 = ~n4347 & n4432;
  assign n4434 = n4347 & ~n4432;
  assign n4435 = ~n4433 & ~n4434;
  assign n4436 = ~n4346 & n4435;
  assign n4437 = n4346 & ~n4435;
  assign n4438 = ~n4436 & ~n4437;
  assign n4439 = n4336 & ~n4438;
  assign n4440 = ~n4336 & n4438;
  assign n4441 = ~n4439 & ~n4440;
  assign n4442 = pi83  & n1296;
  assign n4443 = pi84  & n1207;
  assign n4444 = pi85  & n1202;
  assign n4445 = n1200 & n1831;
  assign n4446 = ~n4443 & ~n4444;
  assign n4447 = ~n4442 & n4446;
  assign n4448 = ~n4445 & n4447;
  assign n4449 = pi17  & n4448;
  assign n4450 = ~pi17  & ~n4448;
  assign n4451 = ~n4449 & ~n4450;
  assign n4452 = n4441 & ~n4451;
  assign n4453 = ~n4441 & n4451;
  assign n4454 = ~n4452 & ~n4453;
  assign n4455 = ~n4335 & n4454;
  assign n4456 = n4335 & ~n4454;
  assign n4457 = ~n4455 & ~n4456;
  assign n4458 = n4334 & ~n4457;
  assign n4459 = ~n4334 & n4457;
  assign n4460 = ~n4458 & ~n4459;
  assign n4461 = ~n4324 & n4460;
  assign n4462 = n4324 & ~n4460;
  assign n4463 = ~n4461 & ~n4462;
  assign n4464 = pi89  & n750;
  assign n4465 = pi90  & n651;
  assign n4466 = pi91  & n646;
  assign n4467 = n644 & n2746;
  assign n4468 = ~n4465 & ~n4466;
  assign n4469 = ~n4464 & n4468;
  assign n4470 = ~n4467 & n4469;
  assign n4471 = pi11  & n4470;
  assign n4472 = ~pi11  & ~n4470;
  assign n4473 = ~n4471 & ~n4472;
  assign n4474 = n4463 & ~n4473;
  assign n4475 = ~n4463 & n4473;
  assign n4476 = ~n4474 & ~n4475;
  assign n4477 = ~n4323 & n4476;
  assign n4478 = n4323 & ~n4476;
  assign n4479 = ~n4477 & ~n4478;
  assign n4480 = n4322 & ~n4479;
  assign n4481 = ~n4322 & n4479;
  assign n4482 = ~n4480 & ~n4481;
  assign n4483 = ~n4312 & n4482;
  assign n4484 = n4312 & ~n4482;
  assign n4485 = ~n4483 & ~n4484;
  assign n4486 = ~n4311 & n4485;
  assign n4487 = n4311 & ~n4485;
  assign n4488 = ~n4486 & ~n4487;
  assign n4489 = ~n4301 & n4488;
  assign n4490 = n4301 & ~n4488;
  assign n4491 = ~n4489 & ~n4490;
  assign n4492 = pi100  & n269;
  assign n4493 = pi99  & n267;
  assign n4494 = pi98  & n282;
  assign n4495 = ~n4097 & ~n4099;
  assign n4496 = ~pi99  & ~pi100 ;
  assign n4497 = pi99  & pi100 ;
  assign n4498 = ~n4496 & ~n4497;
  assign n4499 = ~n4495 & n4498;
  assign n4500 = n4495 & ~n4498;
  assign n4501 = ~n4499 & ~n4500;
  assign n4502 = n262 & n4501;
  assign n4503 = ~n4492 & ~n4493;
  assign n4504 = ~n4494 & n4503;
  assign n4505 = ~n4502 & n4504;
  assign n4506 = pi2  & n4505;
  assign n4507 = ~pi2  & ~n4505;
  assign n4508 = ~n4506 & ~n4507;
  assign n4509 = n4491 & ~n4508;
  assign n4510 = ~n4491 & n4508;
  assign n4511 = ~n4509 & ~n4510;
  assign n4512 = ~n4300 & n4511;
  assign n4513 = n4300 & ~n4511;
  assign po36  = ~n4512 & ~n4513;
  assign n4515 = ~n4509 & ~n4512;
  assign n4516 = ~n4486 & ~n4489;
  assign n4517 = ~n4481 & ~n4483;
  assign n4518 = pi93  & n528;
  assign n4519 = pi94  & n490;
  assign n4520 = pi95  & n485;
  assign n4521 = n483 & n3475;
  assign n4522 = ~n4519 & ~n4520;
  assign n4523 = ~n4518 & n4522;
  assign n4524 = ~n4521 & n4523;
  assign n4525 = pi8  & n4524;
  assign n4526 = ~pi8  & ~n4524;
  assign n4527 = ~n4525 & ~n4526;
  assign n4528 = ~n4474 & ~n4477;
  assign n4529 = pi90  & n750;
  assign n4530 = pi91  & n651;
  assign n4531 = pi92  & n646;
  assign n4532 = n644 & n2924;
  assign n4533 = ~n4530 & ~n4531;
  assign n4534 = ~n4529 & n4533;
  assign n4535 = ~n4532 & n4534;
  assign n4536 = pi11  & n4535;
  assign n4537 = ~pi11  & ~n4535;
  assign n4538 = ~n4536 & ~n4537;
  assign n4539 = ~n4459 & ~n4461;
  assign n4540 = ~n4452 & ~n4455;
  assign n4541 = ~n4436 & ~n4440;
  assign n4542 = ~n4430 & ~n4433;
  assign n4543 = ~n4414 & ~n4417;
  assign n4544 = pi75  & n2510;
  assign n4545 = pi76  & n2342;
  assign n4546 = pi77  & n2337;
  assign n4547 = n865 & n2335;
  assign n4548 = ~n4545 & ~n4546;
  assign n4549 = ~n4544 & n4548;
  assign n4550 = ~n4547 & n4549;
  assign n4551 = pi26  & n4550;
  assign n4552 = ~pi26  & ~n4550;
  assign n4553 = ~n4551 & ~n4552;
  assign n4554 = ~n4397 & ~n4401;
  assign n4555 = pi72  & n3011;
  assign n4556 = pi73  & n2809;
  assign n4557 = pi74  & n2804;
  assign n4558 = n689 & n2802;
  assign n4559 = ~n4556 & ~n4557;
  assign n4560 = ~n4555 & n4559;
  assign n4561 = ~n4558 & n4560;
  assign n4562 = pi29  & n4561;
  assign n4563 = ~pi29  & ~n4561;
  assign n4564 = ~n4562 & ~n4563;
  assign n4565 = ~n4391 & ~n4394;
  assign n4566 = pi69  & n3553;
  assign n4567 = pi70  & n3334;
  assign n4568 = pi71  & n3329;
  assign n4569 = n460 & n3327;
  assign n4570 = ~n4567 & ~n4568;
  assign n4571 = ~n4566 & n4570;
  assign n4572 = ~n4569 & n4571;
  assign n4573 = pi32  & n4572;
  assign n4574 = ~pi32  & ~n4572;
  assign n4575 = ~n4573 & ~n4574;
  assign n4576 = ~n4375 & ~n4378;
  assign n4577 = pi66  & n4176;
  assign n4578 = pi67  & n3938;
  assign n4579 = pi68  & n3933;
  assign n4580 = n334 & n3931;
  assign n4581 = ~n4578 & ~n4579;
  assign n4582 = ~n4577 & n4581;
  assign n4583 = ~n4580 & n4582;
  assign n4584 = pi35  & n4583;
  assign n4585 = ~pi35  & ~n4583;
  assign n4586 = ~n4584 & ~n4585;
  assign n4587 = pi38  & n4373;
  assign n4588 = ~pi37  & ~pi38 ;
  assign n4589 = pi37  & pi38 ;
  assign n4590 = ~n4588 & ~n4589;
  assign n4591 = n4372 & n4590;
  assign n4592 = n265 & n4591;
  assign n4593 = n4372 & ~n4590;
  assign n4594 = pi65  & n4593;
  assign n4595 = ~pi36  & ~pi37 ;
  assign n4596 = pi36  & pi37 ;
  assign n4597 = ~n4595 & ~n4596;
  assign n4598 = ~n4372 & n4597;
  assign n4599 = pi64  & n4598;
  assign n4600 = ~n4592 & ~n4594;
  assign n4601 = ~n4599 & n4600;
  assign n4602 = n4587 & ~n4601;
  assign n4603 = ~n4587 & n4601;
  assign n4604 = ~n4602 & ~n4603;
  assign n4605 = n4586 & ~n4604;
  assign n4606 = ~n4586 & n4604;
  assign n4607 = ~n4605 & ~n4606;
  assign n4608 = ~n4576 & n4607;
  assign n4609 = n4576 & ~n4607;
  assign n4610 = ~n4608 & ~n4609;
  assign n4611 = n4575 & ~n4610;
  assign n4612 = ~n4575 & n4610;
  assign n4613 = ~n4611 & ~n4612;
  assign n4614 = ~n4565 & n4613;
  assign n4615 = n4565 & ~n4613;
  assign n4616 = ~n4614 & ~n4615;
  assign n4617 = n4564 & ~n4616;
  assign n4618 = ~n4564 & n4616;
  assign n4619 = ~n4617 & ~n4618;
  assign n4620 = ~n4554 & n4619;
  assign n4621 = n4554 & ~n4619;
  assign n4622 = ~n4620 & ~n4621;
  assign n4623 = n4553 & ~n4622;
  assign n4624 = ~n4553 & n4622;
  assign n4625 = ~n4623 & ~n4624;
  assign n4626 = ~n4543 & n4625;
  assign n4627 = n4543 & ~n4625;
  assign n4628 = ~n4626 & ~n4627;
  assign n4629 = pi78  & n2053;
  assign n4630 = pi79  & n1893;
  assign n4631 = pi80  & n1888;
  assign n4632 = n1144 & n1886;
  assign n4633 = ~n4630 & ~n4631;
  assign n4634 = ~n4629 & n4633;
  assign n4635 = ~n4632 & n4634;
  assign n4636 = pi23  & n4635;
  assign n4637 = ~pi23  & ~n4635;
  assign n4638 = ~n4636 & ~n4637;
  assign n4639 = n4628 & ~n4638;
  assign n4640 = ~n4628 & n4638;
  assign n4641 = ~n4639 & ~n4640;
  assign n4642 = n4542 & ~n4641;
  assign n4643 = ~n4542 & n4641;
  assign n4644 = ~n4642 & ~n4643;
  assign n4645 = pi81  & n1661;
  assign n4646 = pi82  & n1500;
  assign n4647 = pi83  & n1495;
  assign n4648 = n1493 & n1577;
  assign n4649 = ~n4646 & ~n4647;
  assign n4650 = ~n4645 & n4649;
  assign n4651 = ~n4648 & n4650;
  assign n4652 = pi20  & n4651;
  assign n4653 = ~pi20  & ~n4651;
  assign n4654 = ~n4652 & ~n4653;
  assign n4655 = n4644 & ~n4654;
  assign n4656 = ~n4644 & n4654;
  assign n4657 = ~n4655 & ~n4656;
  assign n4658 = n4541 & ~n4657;
  assign n4659 = ~n4541 & n4657;
  assign n4660 = ~n4658 & ~n4659;
  assign n4661 = pi84  & n1296;
  assign n4662 = pi85  & n1207;
  assign n4663 = pi86  & n1202;
  assign n4664 = n1200 & n1975;
  assign n4665 = ~n4662 & ~n4663;
  assign n4666 = ~n4661 & n4665;
  assign n4667 = ~n4664 & n4666;
  assign n4668 = pi17  & n4667;
  assign n4669 = ~pi17  & ~n4667;
  assign n4670 = ~n4668 & ~n4669;
  assign n4671 = n4660 & ~n4670;
  assign n4672 = ~n4660 & n4670;
  assign n4673 = ~n4671 & ~n4672;
  assign n4674 = n4540 & ~n4673;
  assign n4675 = ~n4540 & n4673;
  assign n4676 = ~n4674 & ~n4675;
  assign n4677 = pi87  & n1006;
  assign n4678 = pi88  & n897;
  assign n4679 = pi89  & n892;
  assign n4680 = n890 & n2287;
  assign n4681 = ~n4678 & ~n4679;
  assign n4682 = ~n4677 & n4681;
  assign n4683 = ~n4680 & n4682;
  assign n4684 = pi14  & n4683;
  assign n4685 = ~pi14  & ~n4683;
  assign n4686 = ~n4684 & ~n4685;
  assign n4687 = n4676 & ~n4686;
  assign n4688 = ~n4676 & n4686;
  assign n4689 = ~n4687 & ~n4688;
  assign n4690 = ~n4539 & n4689;
  assign n4691 = n4539 & ~n4689;
  assign n4692 = ~n4690 & ~n4691;
  assign n4693 = n4538 & ~n4692;
  assign n4694 = ~n4538 & n4692;
  assign n4695 = ~n4693 & ~n4694;
  assign n4696 = ~n4528 & n4695;
  assign n4697 = n4528 & ~n4695;
  assign n4698 = ~n4696 & ~n4697;
  assign n4699 = n4527 & ~n4698;
  assign n4700 = ~n4527 & n4698;
  assign n4701 = ~n4699 & ~n4700;
  assign n4702 = ~n4517 & n4701;
  assign n4703 = n4517 & ~n4701;
  assign n4704 = ~n4702 & ~n4703;
  assign n4705 = pi96  & n391;
  assign n4706 = pi97  & n353;
  assign n4707 = pi98  & n348;
  assign n4708 = n346 & n3889;
  assign n4709 = ~n4706 & ~n4707;
  assign n4710 = ~n4705 & n4709;
  assign n4711 = ~n4708 & n4710;
  assign n4712 = pi5  & n4711;
  assign n4713 = ~pi5  & ~n4711;
  assign n4714 = ~n4712 & ~n4713;
  assign n4715 = n4704 & ~n4714;
  assign n4716 = ~n4704 & n4714;
  assign n4717 = ~n4715 & ~n4716;
  assign n4718 = n4516 & ~n4717;
  assign n4719 = ~n4516 & n4717;
  assign n4720 = ~n4718 & ~n4719;
  assign n4721 = pi101  & n269;
  assign n4722 = pi100  & n267;
  assign n4723 = pi99  & n282;
  assign n4724 = ~n4497 & ~n4499;
  assign n4725 = ~pi100  & ~pi101 ;
  assign n4726 = pi100  & pi101 ;
  assign n4727 = ~n4725 & ~n4726;
  assign n4728 = ~n4724 & n4727;
  assign n4729 = n4724 & ~n4727;
  assign n4730 = ~n4728 & ~n4729;
  assign n4731 = n262 & n4730;
  assign n4732 = ~n4721 & ~n4722;
  assign n4733 = ~n4723 & n4732;
  assign n4734 = ~n4731 & n4733;
  assign n4735 = pi2  & n4734;
  assign n4736 = ~pi2  & ~n4734;
  assign n4737 = ~n4735 & ~n4736;
  assign n4738 = ~n4720 & n4737;
  assign n4739 = n4720 & ~n4737;
  assign n4740 = ~n4738 & ~n4739;
  assign n4741 = ~n4515 & n4740;
  assign n4742 = n4515 & ~n4740;
  assign po37  = ~n4741 & ~n4742;
  assign n4744 = ~n4739 & ~n4741;
  assign n4745 = ~n4715 & ~n4719;
  assign n4746 = pi97  & n391;
  assign n4747 = pi98  & n353;
  assign n4748 = pi99  & n348;
  assign n4749 = n346 & n4101;
  assign n4750 = ~n4747 & ~n4748;
  assign n4751 = ~n4746 & n4750;
  assign n4752 = ~n4749 & n4751;
  assign n4753 = pi5  & n4752;
  assign n4754 = ~pi5  & ~n4752;
  assign n4755 = ~n4753 & ~n4754;
  assign n4756 = ~n4700 & ~n4702;
  assign n4757 = pi94  & n528;
  assign n4758 = pi95  & n490;
  assign n4759 = pi96  & n485;
  assign n4760 = n483 & n3499;
  assign n4761 = ~n4758 & ~n4759;
  assign n4762 = ~n4757 & n4761;
  assign n4763 = ~n4760 & n4762;
  assign n4764 = pi8  & n4763;
  assign n4765 = ~pi8  & ~n4763;
  assign n4766 = ~n4764 & ~n4765;
  assign n4767 = ~n4694 & ~n4696;
  assign n4768 = pi91  & n750;
  assign n4769 = pi92  & n651;
  assign n4770 = pi93  & n646;
  assign n4771 = n644 & n2948;
  assign n4772 = ~n4769 & ~n4770;
  assign n4773 = ~n4768 & n4772;
  assign n4774 = ~n4771 & n4773;
  assign n4775 = pi11  & n4774;
  assign n4776 = ~pi11  & ~n4774;
  assign n4777 = ~n4775 & ~n4776;
  assign n4778 = ~n4687 & ~n4690;
  assign n4779 = pi88  & n1006;
  assign n4780 = pi89  & n897;
  assign n4781 = pi90  & n892;
  assign n4782 = n890 & n2448;
  assign n4783 = ~n4780 & ~n4781;
  assign n4784 = ~n4779 & n4783;
  assign n4785 = ~n4782 & n4784;
  assign n4786 = pi14  & n4785;
  assign n4787 = ~pi14  & ~n4785;
  assign n4788 = ~n4786 & ~n4787;
  assign n4789 = ~n4671 & ~n4675;
  assign n4790 = ~n4655 & ~n4659;
  assign n4791 = ~n4639 & ~n4643;
  assign n4792 = ~n4624 & ~n4626;
  assign n4793 = pi76  & n2510;
  assign n4794 = pi77  & n2342;
  assign n4795 = pi78  & n2337;
  assign n4796 = n958 & n2335;
  assign n4797 = ~n4794 & ~n4795;
  assign n4798 = ~n4793 & n4797;
  assign n4799 = ~n4796 & n4798;
  assign n4800 = pi26  & n4799;
  assign n4801 = ~pi26  & ~n4799;
  assign n4802 = ~n4800 & ~n4801;
  assign n4803 = ~n4618 & ~n4620;
  assign n4804 = pi73  & n3011;
  assign n4805 = pi74  & n2809;
  assign n4806 = pi75  & n2804;
  assign n4807 = n713 & n2802;
  assign n4808 = ~n4805 & ~n4806;
  assign n4809 = ~n4804 & n4808;
  assign n4810 = ~n4807 & n4809;
  assign n4811 = pi29  & n4810;
  assign n4812 = ~pi29  & ~n4810;
  assign n4813 = ~n4811 & ~n4812;
  assign n4814 = ~n4612 & ~n4614;
  assign n4815 = pi70  & n3553;
  assign n4816 = pi71  & n3334;
  assign n4817 = pi72  & n3329;
  assign n4818 = n551 & n3327;
  assign n4819 = ~n4816 & ~n4817;
  assign n4820 = ~n4815 & n4819;
  assign n4821 = ~n4818 & n4820;
  assign n4822 = pi32  & n4821;
  assign n4823 = ~pi32  & ~n4821;
  assign n4824 = ~n4822 & ~n4823;
  assign n4825 = ~n4606 & ~n4608;
  assign n4826 = pi67  & n4176;
  assign n4827 = pi68  & n3938;
  assign n4828 = pi69  & n3933;
  assign n4829 = n376 & n3931;
  assign n4830 = ~n4827 & ~n4828;
  assign n4831 = ~n4826 & n4830;
  assign n4832 = ~n4829 & n4831;
  assign n4833 = pi35  & n4832;
  assign n4834 = ~pi35  & ~n4832;
  assign n4835 = ~n4833 & ~n4834;
  assign n4836 = pi38  & ~n4373;
  assign n4837 = n4601 & n4836;
  assign n4838 = pi38  & ~n4837;
  assign n4839 = ~n287 & n4591;
  assign n4840 = pi65  & n4598;
  assign n4841 = pi66  & n4593;
  assign n4842 = ~n4372 & n4590;
  assign n4843 = ~n4597 & n4842;
  assign n4844 = pi64  & n4843;
  assign n4845 = ~n4839 & ~n4840;
  assign n4846 = ~n4841 & n4845;
  assign n4847 = ~n4844 & n4846;
  assign n4848 = ~n4838 & n4847;
  assign n4849 = n4838 & ~n4847;
  assign n4850 = ~n4848 & ~n4849;
  assign n4851 = ~n4835 & n4850;
  assign n4852 = n4835 & ~n4850;
  assign n4853 = ~n4851 & ~n4852;
  assign n4854 = ~n4825 & n4853;
  assign n4855 = n4825 & ~n4853;
  assign n4856 = ~n4854 & ~n4855;
  assign n4857 = ~n4824 & n4856;
  assign n4858 = n4824 & ~n4856;
  assign n4859 = ~n4857 & ~n4858;
  assign n4860 = ~n4814 & n4859;
  assign n4861 = n4814 & ~n4859;
  assign n4862 = ~n4860 & ~n4861;
  assign n4863 = ~n4813 & n4862;
  assign n4864 = n4813 & ~n4862;
  assign n4865 = ~n4863 & ~n4864;
  assign n4866 = ~n4803 & n4865;
  assign n4867 = n4803 & ~n4865;
  assign n4868 = ~n4866 & ~n4867;
  assign n4869 = n4802 & ~n4868;
  assign n4870 = ~n4802 & n4868;
  assign n4871 = ~n4869 & ~n4870;
  assign n4872 = ~n4792 & n4871;
  assign n4873 = n4792 & ~n4871;
  assign n4874 = ~n4872 & ~n4873;
  assign n4875 = pi79  & n2053;
  assign n4876 = pi80  & n1893;
  assign n4877 = pi81  & n1888;
  assign n4878 = n1337 & n1886;
  assign n4879 = ~n4876 & ~n4877;
  assign n4880 = ~n4875 & n4879;
  assign n4881 = ~n4878 & n4880;
  assign n4882 = pi23  & n4881;
  assign n4883 = ~pi23  & ~n4881;
  assign n4884 = ~n4882 & ~n4883;
  assign n4885 = n4874 & ~n4884;
  assign n4886 = ~n4874 & n4884;
  assign n4887 = ~n4885 & ~n4886;
  assign n4888 = n4791 & ~n4887;
  assign n4889 = ~n4791 & n4887;
  assign n4890 = ~n4888 & ~n4889;
  assign n4891 = pi82  & n1661;
  assign n4892 = pi83  & n1500;
  assign n4893 = pi84  & n1495;
  assign n4894 = n1493 & n1601;
  assign n4895 = ~n4892 & ~n4893;
  assign n4896 = ~n4891 & n4895;
  assign n4897 = ~n4894 & n4896;
  assign n4898 = pi20  & n4897;
  assign n4899 = ~pi20  & ~n4897;
  assign n4900 = ~n4898 & ~n4899;
  assign n4901 = n4890 & ~n4900;
  assign n4902 = ~n4890 & n4900;
  assign n4903 = ~n4901 & ~n4902;
  assign n4904 = n4790 & ~n4903;
  assign n4905 = ~n4790 & n4903;
  assign n4906 = ~n4904 & ~n4905;
  assign n4907 = pi85  & n1296;
  assign n4908 = pi86  & n1207;
  assign n4909 = pi87  & n1202;
  assign n4910 = n1200 & n2116;
  assign n4911 = ~n4908 & ~n4909;
  assign n4912 = ~n4907 & n4911;
  assign n4913 = ~n4910 & n4912;
  assign n4914 = pi17  & n4913;
  assign n4915 = ~pi17  & ~n4913;
  assign n4916 = ~n4914 & ~n4915;
  assign n4917 = n4906 & ~n4916;
  assign n4918 = ~n4906 & n4916;
  assign n4919 = ~n4917 & ~n4918;
  assign n4920 = ~n4789 & n4919;
  assign n4921 = n4789 & ~n4919;
  assign n4922 = ~n4920 & ~n4921;
  assign n4923 = n4788 & ~n4922;
  assign n4924 = ~n4788 & n4922;
  assign n4925 = ~n4923 & ~n4924;
  assign n4926 = ~n4778 & n4925;
  assign n4927 = n4778 & ~n4925;
  assign n4928 = ~n4926 & ~n4927;
  assign n4929 = n4777 & ~n4928;
  assign n4930 = ~n4777 & n4928;
  assign n4931 = ~n4929 & ~n4930;
  assign n4932 = ~n4767 & n4931;
  assign n4933 = n4767 & ~n4931;
  assign n4934 = ~n4932 & ~n4933;
  assign n4935 = n4766 & ~n4934;
  assign n4936 = ~n4766 & n4934;
  assign n4937 = ~n4935 & ~n4936;
  assign n4938 = ~n4756 & n4937;
  assign n4939 = n4756 & ~n4937;
  assign n4940 = ~n4938 & ~n4939;
  assign n4941 = n4755 & ~n4940;
  assign n4942 = ~n4755 & n4940;
  assign n4943 = ~n4941 & ~n4942;
  assign n4944 = ~n4745 & n4943;
  assign n4945 = n4745 & ~n4943;
  assign n4946 = ~n4944 & ~n4945;
  assign n4947 = pi102  & n269;
  assign n4948 = pi101  & n267;
  assign n4949 = pi100  & n282;
  assign n4950 = ~n4726 & ~n4728;
  assign n4951 = ~pi101  & ~pi102 ;
  assign n4952 = pi101  & pi102 ;
  assign n4953 = ~n4951 & ~n4952;
  assign n4954 = ~n4950 & n4953;
  assign n4955 = n4950 & ~n4953;
  assign n4956 = ~n4954 & ~n4955;
  assign n4957 = n262 & n4956;
  assign n4958 = ~n4947 & ~n4948;
  assign n4959 = ~n4949 & n4958;
  assign n4960 = ~n4957 & n4959;
  assign n4961 = pi2  & n4960;
  assign n4962 = ~pi2  & ~n4960;
  assign n4963 = ~n4961 & ~n4962;
  assign n4964 = n4946 & ~n4963;
  assign n4965 = ~n4946 & n4963;
  assign n4966 = ~n4964 & ~n4965;
  assign n4967 = ~n4744 & n4966;
  assign n4968 = n4744 & ~n4966;
  assign po38  = ~n4967 & ~n4968;
  assign n4970 = ~n4964 & ~n4967;
  assign n4971 = ~n4942 & ~n4944;
  assign n4972 = pi98  & n391;
  assign n4973 = pi99  & n353;
  assign n4974 = pi100  & n348;
  assign n4975 = n346 & n4501;
  assign n4976 = ~n4973 & ~n4974;
  assign n4977 = ~n4972 & n4976;
  assign n4978 = ~n4975 & n4977;
  assign n4979 = pi5  & n4978;
  assign n4980 = ~pi5  & ~n4978;
  assign n4981 = ~n4979 & ~n4980;
  assign n4982 = ~n4936 & ~n4938;
  assign n4983 = ~n4930 & ~n4932;
  assign n4984 = pi92  & n750;
  assign n4985 = pi93  & n651;
  assign n4986 = pi94  & n646;
  assign n4987 = n644 & n3280;
  assign n4988 = ~n4985 & ~n4986;
  assign n4989 = ~n4984 & n4988;
  assign n4990 = ~n4987 & n4989;
  assign n4991 = pi11  & n4990;
  assign n4992 = ~pi11  & ~n4990;
  assign n4993 = ~n4991 & ~n4992;
  assign n4994 = ~n4924 & ~n4926;
  assign n4995 = ~n4917 & ~n4920;
  assign n4996 = ~n4901 & ~n4905;
  assign n4997 = ~n4885 & ~n4889;
  assign n4998 = pi80  & n2053;
  assign n4999 = pi81  & n1893;
  assign n5000 = pi82  & n1888;
  assign n5001 = n1450 & n1886;
  assign n5002 = ~n4999 & ~n5000;
  assign n5003 = ~n4998 & n5002;
  assign n5004 = ~n5001 & n5003;
  assign n5005 = pi23  & n5004;
  assign n5006 = ~pi23  & ~n5004;
  assign n5007 = ~n5005 & ~n5006;
  assign n5008 = ~n4870 & ~n4872;
  assign n5009 = ~n4857 & ~n4860;
  assign n5010 = ~n4851 & ~n4854;
  assign n5011 = pi65  & n4843;
  assign n5012 = pi66  & n4598;
  assign n5013 = pi67  & n4593;
  assign n5014 = n305 & n4591;
  assign n5015 = ~n5012 & ~n5013;
  assign n5016 = ~n5011 & n5015;
  assign n5017 = ~n5014 & n5016;
  assign n5018 = pi38  & n5017;
  assign n5019 = ~pi38  & ~n5017;
  assign n5020 = ~n5018 & ~n5019;
  assign n5021 = ~pi38  & ~pi39 ;
  assign n5022 = pi38  & pi39 ;
  assign n5023 = ~n5021 & ~n5022;
  assign n5024 = pi64  & n5023;
  assign n5025 = n4837 & n4847;
  assign n5026 = n5024 & n5025;
  assign n5027 = ~n5024 & ~n5025;
  assign n5028 = ~n5026 & ~n5027;
  assign n5029 = ~n5020 & n5028;
  assign n5030 = n5020 & ~n5028;
  assign n5031 = ~n5029 & ~n5030;
  assign n5032 = pi68  & n4176;
  assign n5033 = pi69  & n3938;
  assign n5034 = pi70  & n3933;
  assign n5035 = n415 & n3931;
  assign n5036 = ~n5033 & ~n5034;
  assign n5037 = ~n5032 & n5036;
  assign n5038 = ~n5035 & n5037;
  assign n5039 = pi35  & n5038;
  assign n5040 = ~pi35  & ~n5038;
  assign n5041 = ~n5039 & ~n5040;
  assign n5042 = n5031 & ~n5041;
  assign n5043 = ~n5031 & n5041;
  assign n5044 = ~n5042 & ~n5043;
  assign n5045 = n5010 & ~n5044;
  assign n5046 = ~n5010 & n5044;
  assign n5047 = ~n5045 & ~n5046;
  assign n5048 = pi71  & n3553;
  assign n5049 = pi72  & n3334;
  assign n5050 = pi73  & n3329;
  assign n5051 = n613 & n3327;
  assign n5052 = ~n5049 & ~n5050;
  assign n5053 = ~n5048 & n5052;
  assign n5054 = ~n5051 & n5053;
  assign n5055 = pi32  & n5054;
  assign n5056 = ~pi32  & ~n5054;
  assign n5057 = ~n5055 & ~n5056;
  assign n5058 = n5047 & ~n5057;
  assign n5059 = ~n5047 & n5057;
  assign n5060 = ~n5058 & ~n5059;
  assign n5061 = n5009 & ~n5060;
  assign n5062 = ~n5009 & n5060;
  assign n5063 = ~n5061 & ~n5062;
  assign n5064 = pi74  & n3011;
  assign n5065 = pi75  & n2809;
  assign n5066 = pi76  & n2804;
  assign n5067 = n841 & n2802;
  assign n5068 = ~n5065 & ~n5066;
  assign n5069 = ~n5064 & n5068;
  assign n5070 = ~n5067 & n5069;
  assign n5071 = pi29  & n5070;
  assign n5072 = ~pi29  & ~n5070;
  assign n5073 = ~n5071 & ~n5072;
  assign n5074 = ~n5063 & n5073;
  assign n5075 = n5063 & ~n5073;
  assign n5076 = ~n5074 & ~n5075;
  assign n5077 = ~n4863 & ~n4866;
  assign n5078 = n5076 & ~n5077;
  assign n5079 = ~n5076 & n5077;
  assign n5080 = ~n5078 & ~n5079;
  assign n5081 = pi77  & n2510;
  assign n5082 = pi78  & n2342;
  assign n5083 = pi79  & n2337;
  assign n5084 = n1048 & n2335;
  assign n5085 = ~n5082 & ~n5083;
  assign n5086 = ~n5081 & n5085;
  assign n5087 = ~n5084 & n5086;
  assign n5088 = pi26  & n5087;
  assign n5089 = ~pi26  & ~n5087;
  assign n5090 = ~n5088 & ~n5089;
  assign n5091 = n5080 & ~n5090;
  assign n5092 = ~n5080 & n5090;
  assign n5093 = ~n5091 & ~n5092;
  assign n5094 = ~n5008 & n5093;
  assign n5095 = n5008 & ~n5093;
  assign n5096 = ~n5094 & ~n5095;
  assign n5097 = ~n5007 & n5096;
  assign n5098 = n5007 & ~n5096;
  assign n5099 = ~n5097 & ~n5098;
  assign n5100 = n4997 & ~n5099;
  assign n5101 = ~n4997 & n5099;
  assign n5102 = ~n5100 & ~n5101;
  assign n5103 = pi83  & n1661;
  assign n5104 = pi84  & n1500;
  assign n5105 = pi85  & n1495;
  assign n5106 = n1493 & n1831;
  assign n5107 = ~n5104 & ~n5105;
  assign n5108 = ~n5103 & n5107;
  assign n5109 = ~n5106 & n5108;
  assign n5110 = pi20  & n5109;
  assign n5111 = ~pi20  & ~n5109;
  assign n5112 = ~n5110 & ~n5111;
  assign n5113 = n5102 & ~n5112;
  assign n5114 = ~n5102 & n5112;
  assign n5115 = ~n5113 & ~n5114;
  assign n5116 = n4996 & ~n5115;
  assign n5117 = ~n4996 & n5115;
  assign n5118 = ~n5116 & ~n5117;
  assign n5119 = pi86  & n1296;
  assign n5120 = pi87  & n1207;
  assign n5121 = pi88  & n1202;
  assign n5122 = n1200 & n2140;
  assign n5123 = ~n5120 & ~n5121;
  assign n5124 = ~n5119 & n5123;
  assign n5125 = ~n5122 & n5124;
  assign n5126 = pi17  & n5125;
  assign n5127 = ~pi17  & ~n5125;
  assign n5128 = ~n5126 & ~n5127;
  assign n5129 = ~n5118 & n5128;
  assign n5130 = n5118 & ~n5128;
  assign n5131 = ~n5129 & ~n5130;
  assign n5132 = ~n4995 & n5131;
  assign n5133 = n4995 & ~n5131;
  assign n5134 = ~n5132 & ~n5133;
  assign n5135 = pi89  & n1006;
  assign n5136 = pi90  & n897;
  assign n5137 = pi91  & n892;
  assign n5138 = n890 & n2746;
  assign n5139 = ~n5136 & ~n5137;
  assign n5140 = ~n5135 & n5139;
  assign n5141 = ~n5138 & n5140;
  assign n5142 = pi14  & n5141;
  assign n5143 = ~pi14  & ~n5141;
  assign n5144 = ~n5142 & ~n5143;
  assign n5145 = n5134 & ~n5144;
  assign n5146 = ~n5134 & n5144;
  assign n5147 = ~n5145 & ~n5146;
  assign n5148 = ~n4994 & n5147;
  assign n5149 = n4994 & ~n5147;
  assign n5150 = ~n5148 & ~n5149;
  assign n5151 = ~n4993 & n5150;
  assign n5152 = n4993 & ~n5150;
  assign n5153 = ~n5151 & ~n5152;
  assign n5154 = ~n4983 & n5153;
  assign n5155 = n4983 & ~n5153;
  assign n5156 = ~n5154 & ~n5155;
  assign n5157 = pi95  & n528;
  assign n5158 = pi96  & n490;
  assign n5159 = pi97  & n485;
  assign n5160 = n483 & n3691;
  assign n5161 = ~n5158 & ~n5159;
  assign n5162 = ~n5157 & n5161;
  assign n5163 = ~n5160 & n5162;
  assign n5164 = pi8  & n5163;
  assign n5165 = ~pi8  & ~n5163;
  assign n5166 = ~n5164 & ~n5165;
  assign n5167 = n5156 & ~n5166;
  assign n5168 = ~n5156 & n5166;
  assign n5169 = ~n5167 & ~n5168;
  assign n5170 = ~n4982 & n5169;
  assign n5171 = n4982 & ~n5169;
  assign n5172 = ~n5170 & ~n5171;
  assign n5173 = n4981 & ~n5172;
  assign n5174 = ~n4981 & n5172;
  assign n5175 = ~n5173 & ~n5174;
  assign n5176 = ~n4971 & n5175;
  assign n5177 = n4971 & ~n5175;
  assign n5178 = ~n5176 & ~n5177;
  assign n5179 = pi103  & n269;
  assign n5180 = pi102  & n267;
  assign n5181 = pi101  & n282;
  assign n5182 = ~n4952 & ~n4954;
  assign n5183 = ~pi102  & ~pi103 ;
  assign n5184 = pi102  & pi103 ;
  assign n5185 = ~n5183 & ~n5184;
  assign n5186 = ~n5182 & n5185;
  assign n5187 = n5182 & ~n5185;
  assign n5188 = ~n5186 & ~n5187;
  assign n5189 = n262 & n5188;
  assign n5190 = ~n5179 & ~n5180;
  assign n5191 = ~n5181 & n5190;
  assign n5192 = ~n5189 & n5191;
  assign n5193 = pi2  & n5192;
  assign n5194 = ~pi2  & ~n5192;
  assign n5195 = ~n5193 & ~n5194;
  assign n5196 = n5178 & ~n5195;
  assign n5197 = ~n5178 & n5195;
  assign n5198 = ~n5196 & ~n5197;
  assign n5199 = ~n4970 & n5198;
  assign n5200 = n4970 & ~n5198;
  assign po39  = ~n5199 & ~n5200;
  assign n5202 = ~n5196 & ~n5199;
  assign n5203 = pi104  & n269;
  assign n5204 = pi103  & n267;
  assign n5205 = pi102  & n282;
  assign n5206 = ~n5184 & ~n5186;
  assign n5207 = ~pi103  & ~pi104 ;
  assign n5208 = pi103  & pi104 ;
  assign n5209 = ~n5207 & ~n5208;
  assign n5210 = ~n5206 & n5209;
  assign n5211 = n5206 & ~n5209;
  assign n5212 = ~n5210 & ~n5211;
  assign n5213 = n262 & n5212;
  assign n5214 = ~n5203 & ~n5204;
  assign n5215 = ~n5205 & n5214;
  assign n5216 = ~n5213 & n5215;
  assign n5217 = pi2  & n5216;
  assign n5218 = ~pi2  & ~n5216;
  assign n5219 = ~n5217 & ~n5218;
  assign n5220 = ~n5174 & ~n5176;
  assign n5221 = ~n5167 & ~n5170;
  assign n5222 = pi96  & n528;
  assign n5223 = pi97  & n490;
  assign n5224 = pi98  & n485;
  assign n5225 = n483 & n3889;
  assign n5226 = ~n5223 & ~n5224;
  assign n5227 = ~n5222 & n5226;
  assign n5228 = ~n5225 & n5227;
  assign n5229 = pi8  & n5228;
  assign n5230 = ~pi8  & ~n5228;
  assign n5231 = ~n5229 & ~n5230;
  assign n5232 = ~n5151 & ~n5154;
  assign n5233 = pi93  & n750;
  assign n5234 = pi94  & n651;
  assign n5235 = pi95  & n646;
  assign n5236 = n644 & n3475;
  assign n5237 = ~n5234 & ~n5235;
  assign n5238 = ~n5233 & n5237;
  assign n5239 = ~n5236 & n5238;
  assign n5240 = pi11  & n5239;
  assign n5241 = ~pi11  & ~n5239;
  assign n5242 = ~n5240 & ~n5241;
  assign n5243 = ~n5145 & ~n5148;
  assign n5244 = pi90  & n1006;
  assign n5245 = pi91  & n897;
  assign n5246 = pi92  & n892;
  assign n5247 = n890 & n2924;
  assign n5248 = ~n5245 & ~n5246;
  assign n5249 = ~n5244 & n5248;
  assign n5250 = ~n5247 & n5249;
  assign n5251 = pi14  & n5250;
  assign n5252 = ~pi14  & ~n5250;
  assign n5253 = ~n5251 & ~n5252;
  assign n5254 = ~n5130 & ~n5132;
  assign n5255 = ~n5113 & ~n5117;
  assign n5256 = ~n5097 & ~n5101;
  assign n5257 = ~n5091 & ~n5094;
  assign n5258 = ~n5075 & ~n5078;
  assign n5259 = pi75  & n3011;
  assign n5260 = pi76  & n2809;
  assign n5261 = pi77  & n2804;
  assign n5262 = n865 & n2802;
  assign n5263 = ~n5260 & ~n5261;
  assign n5264 = ~n5259 & n5263;
  assign n5265 = ~n5262 & n5264;
  assign n5266 = pi29  & n5265;
  assign n5267 = ~pi29  & ~n5265;
  assign n5268 = ~n5266 & ~n5267;
  assign n5269 = ~n5058 & ~n5062;
  assign n5270 = ~n5042 & ~n5046;
  assign n5271 = ~n5026 & ~n5029;
  assign n5272 = pi66  & n4843;
  assign n5273 = pi67  & n4598;
  assign n5274 = pi68  & n4593;
  assign n5275 = n334 & n4591;
  assign n5276 = ~n5273 & ~n5274;
  assign n5277 = ~n5272 & n5276;
  assign n5278 = ~n5275 & n5277;
  assign n5279 = pi38  & n5278;
  assign n5280 = ~pi38  & ~n5278;
  assign n5281 = ~n5279 & ~n5280;
  assign n5282 = pi41  & n5024;
  assign n5283 = ~pi40  & ~pi41 ;
  assign n5284 = pi40  & pi41 ;
  assign n5285 = ~n5283 & ~n5284;
  assign n5286 = n5023 & n5285;
  assign n5287 = n265 & n5286;
  assign n5288 = n5023 & ~n5285;
  assign n5289 = pi65  & n5288;
  assign n5290 = ~pi39  & ~pi40 ;
  assign n5291 = pi39  & pi40 ;
  assign n5292 = ~n5290 & ~n5291;
  assign n5293 = ~n5023 & n5292;
  assign n5294 = pi64  & n5293;
  assign n5295 = ~n5287 & ~n5289;
  assign n5296 = ~n5294 & n5295;
  assign n5297 = n5282 & ~n5296;
  assign n5298 = ~n5282 & n5296;
  assign n5299 = ~n5297 & ~n5298;
  assign n5300 = n5281 & ~n5299;
  assign n5301 = ~n5281 & n5299;
  assign n5302 = ~n5300 & ~n5301;
  assign n5303 = ~n5271 & n5302;
  assign n5304 = n5271 & ~n5302;
  assign n5305 = ~n5303 & ~n5304;
  assign n5306 = pi69  & n4176;
  assign n5307 = pi70  & n3938;
  assign n5308 = pi71  & n3933;
  assign n5309 = n460 & n3931;
  assign n5310 = ~n5307 & ~n5308;
  assign n5311 = ~n5306 & n5310;
  assign n5312 = ~n5309 & n5311;
  assign n5313 = pi35  & n5312;
  assign n5314 = ~pi35  & ~n5312;
  assign n5315 = ~n5313 & ~n5314;
  assign n5316 = n5305 & ~n5315;
  assign n5317 = ~n5305 & n5315;
  assign n5318 = ~n5316 & ~n5317;
  assign n5319 = n5270 & ~n5318;
  assign n5320 = ~n5270 & n5318;
  assign n5321 = ~n5319 & ~n5320;
  assign n5322 = pi72  & n3553;
  assign n5323 = pi73  & n3334;
  assign n5324 = pi74  & n3329;
  assign n5325 = n689 & n3327;
  assign n5326 = ~n5323 & ~n5324;
  assign n5327 = ~n5322 & n5326;
  assign n5328 = ~n5325 & n5327;
  assign n5329 = pi32  & n5328;
  assign n5330 = ~pi32  & ~n5328;
  assign n5331 = ~n5329 & ~n5330;
  assign n5332 = n5321 & ~n5331;
  assign n5333 = ~n5321 & n5331;
  assign n5334 = ~n5332 & ~n5333;
  assign n5335 = ~n5269 & n5334;
  assign n5336 = n5269 & ~n5334;
  assign n5337 = ~n5335 & ~n5336;
  assign n5338 = n5268 & ~n5337;
  assign n5339 = ~n5268 & n5337;
  assign n5340 = ~n5338 & ~n5339;
  assign n5341 = ~n5258 & n5340;
  assign n5342 = n5258 & ~n5340;
  assign n5343 = ~n5341 & ~n5342;
  assign n5344 = pi78  & n2510;
  assign n5345 = pi79  & n2342;
  assign n5346 = pi80  & n2337;
  assign n5347 = n1144 & n2335;
  assign n5348 = ~n5345 & ~n5346;
  assign n5349 = ~n5344 & n5348;
  assign n5350 = ~n5347 & n5349;
  assign n5351 = pi26  & n5350;
  assign n5352 = ~pi26  & ~n5350;
  assign n5353 = ~n5351 & ~n5352;
  assign n5354 = n5343 & ~n5353;
  assign n5355 = ~n5343 & n5353;
  assign n5356 = ~n5354 & ~n5355;
  assign n5357 = n5257 & ~n5356;
  assign n5358 = ~n5257 & n5356;
  assign n5359 = ~n5357 & ~n5358;
  assign n5360 = pi81  & n2053;
  assign n5361 = pi82  & n1893;
  assign n5362 = pi83  & n1888;
  assign n5363 = n1577 & n1886;
  assign n5364 = ~n5361 & ~n5362;
  assign n5365 = ~n5360 & n5364;
  assign n5366 = ~n5363 & n5365;
  assign n5367 = pi23  & n5366;
  assign n5368 = ~pi23  & ~n5366;
  assign n5369 = ~n5367 & ~n5368;
  assign n5370 = n5359 & ~n5369;
  assign n5371 = ~n5359 & n5369;
  assign n5372 = ~n5370 & ~n5371;
  assign n5373 = n5256 & ~n5372;
  assign n5374 = ~n5256 & n5372;
  assign n5375 = ~n5373 & ~n5374;
  assign n5376 = pi84  & n1661;
  assign n5377 = pi85  & n1500;
  assign n5378 = pi86  & n1495;
  assign n5379 = n1493 & n1975;
  assign n5380 = ~n5377 & ~n5378;
  assign n5381 = ~n5376 & n5380;
  assign n5382 = ~n5379 & n5381;
  assign n5383 = pi20  & n5382;
  assign n5384 = ~pi20  & ~n5382;
  assign n5385 = ~n5383 & ~n5384;
  assign n5386 = n5375 & ~n5385;
  assign n5387 = ~n5375 & n5385;
  assign n5388 = ~n5386 & ~n5387;
  assign n5389 = n5255 & ~n5388;
  assign n5390 = ~n5255 & n5388;
  assign n5391 = ~n5389 & ~n5390;
  assign n5392 = pi87  & n1296;
  assign n5393 = pi88  & n1207;
  assign n5394 = pi89  & n1202;
  assign n5395 = n1200 & n2287;
  assign n5396 = ~n5393 & ~n5394;
  assign n5397 = ~n5392 & n5396;
  assign n5398 = ~n5395 & n5397;
  assign n5399 = pi17  & n5398;
  assign n5400 = ~pi17  & ~n5398;
  assign n5401 = ~n5399 & ~n5400;
  assign n5402 = n5391 & ~n5401;
  assign n5403 = ~n5391 & n5401;
  assign n5404 = ~n5402 & ~n5403;
  assign n5405 = ~n5254 & n5404;
  assign n5406 = n5254 & ~n5404;
  assign n5407 = ~n5405 & ~n5406;
  assign n5408 = ~n5253 & n5407;
  assign n5409 = n5253 & ~n5407;
  assign n5410 = ~n5408 & ~n5409;
  assign n5411 = ~n5243 & n5410;
  assign n5412 = n5243 & ~n5410;
  assign n5413 = ~n5411 & ~n5412;
  assign n5414 = n5242 & ~n5413;
  assign n5415 = ~n5242 & n5413;
  assign n5416 = ~n5414 & ~n5415;
  assign n5417 = ~n5232 & n5416;
  assign n5418 = n5232 & ~n5416;
  assign n5419 = ~n5417 & ~n5418;
  assign n5420 = n5231 & ~n5419;
  assign n5421 = ~n5231 & n5419;
  assign n5422 = ~n5420 & ~n5421;
  assign n5423 = ~n5221 & n5422;
  assign n5424 = n5221 & ~n5422;
  assign n5425 = ~n5423 & ~n5424;
  assign n5426 = pi99  & n391;
  assign n5427 = pi100  & n353;
  assign n5428 = pi101  & n348;
  assign n5429 = n346 & n4730;
  assign n5430 = ~n5427 & ~n5428;
  assign n5431 = ~n5426 & n5430;
  assign n5432 = ~n5429 & n5431;
  assign n5433 = pi5  & n5432;
  assign n5434 = ~pi5  & ~n5432;
  assign n5435 = ~n5433 & ~n5434;
  assign n5436 = n5425 & ~n5435;
  assign n5437 = ~n5425 & n5435;
  assign n5438 = ~n5436 & ~n5437;
  assign n5439 = ~n5220 & n5438;
  assign n5440 = n5220 & ~n5438;
  assign n5441 = ~n5439 & ~n5440;
  assign n5442 = ~n5219 & n5441;
  assign n5443 = n5219 & ~n5441;
  assign n5444 = ~n5442 & ~n5443;
  assign n5445 = ~n5202 & n5444;
  assign n5446 = n5202 & ~n5444;
  assign po40  = ~n5445 & ~n5446;
  assign n5448 = ~n5442 & ~n5445;
  assign n5449 = ~n5436 & ~n5439;
  assign n5450 = pi100  & n391;
  assign n5451 = pi101  & n353;
  assign n5452 = pi102  & n348;
  assign n5453 = n346 & n4956;
  assign n5454 = ~n5451 & ~n5452;
  assign n5455 = ~n5450 & n5454;
  assign n5456 = ~n5453 & n5455;
  assign n5457 = pi5  & n5456;
  assign n5458 = ~pi5  & ~n5456;
  assign n5459 = ~n5457 & ~n5458;
  assign n5460 = ~n5421 & ~n5423;
  assign n5461 = ~n5415 & ~n5417;
  assign n5462 = pi94  & n750;
  assign n5463 = pi95  & n651;
  assign n5464 = pi96  & n646;
  assign n5465 = n644 & n3499;
  assign n5466 = ~n5463 & ~n5464;
  assign n5467 = ~n5462 & n5466;
  assign n5468 = ~n5465 & n5467;
  assign n5469 = pi11  & n5468;
  assign n5470 = ~pi11  & ~n5468;
  assign n5471 = ~n5469 & ~n5470;
  assign n5472 = ~n5408 & ~n5411;
  assign n5473 = pi91  & n1006;
  assign n5474 = pi92  & n897;
  assign n5475 = pi93  & n892;
  assign n5476 = n890 & n2948;
  assign n5477 = ~n5474 & ~n5475;
  assign n5478 = ~n5473 & n5477;
  assign n5479 = ~n5476 & n5478;
  assign n5480 = pi14  & n5479;
  assign n5481 = ~pi14  & ~n5479;
  assign n5482 = ~n5480 & ~n5481;
  assign n5483 = ~n5402 & ~n5405;
  assign n5484 = pi88  & n1296;
  assign n5485 = pi89  & n1207;
  assign n5486 = pi90  & n1202;
  assign n5487 = n1200 & n2448;
  assign n5488 = ~n5485 & ~n5486;
  assign n5489 = ~n5484 & n5488;
  assign n5490 = ~n5487 & n5489;
  assign n5491 = pi17  & n5490;
  assign n5492 = ~pi17  & ~n5490;
  assign n5493 = ~n5491 & ~n5492;
  assign n5494 = ~n5386 & ~n5390;
  assign n5495 = ~n5370 & ~n5374;
  assign n5496 = ~n5354 & ~n5358;
  assign n5497 = pi79  & n2510;
  assign n5498 = pi80  & n2342;
  assign n5499 = pi81  & n2337;
  assign n5500 = n1337 & n2335;
  assign n5501 = ~n5498 & ~n5499;
  assign n5502 = ~n5497 & n5501;
  assign n5503 = ~n5500 & n5502;
  assign n5504 = pi26  & n5503;
  assign n5505 = ~pi26  & ~n5503;
  assign n5506 = ~n5504 & ~n5505;
  assign n5507 = ~n5339 & ~n5341;
  assign n5508 = pi76  & n3011;
  assign n5509 = pi77  & n2809;
  assign n5510 = pi78  & n2804;
  assign n5511 = n958 & n2802;
  assign n5512 = ~n5509 & ~n5510;
  assign n5513 = ~n5508 & n5512;
  assign n5514 = ~n5511 & n5513;
  assign n5515 = pi29  & n5514;
  assign n5516 = ~pi29  & ~n5514;
  assign n5517 = ~n5515 & ~n5516;
  assign n5518 = ~n5332 & ~n5335;
  assign n5519 = pi73  & n3553;
  assign n5520 = pi74  & n3334;
  assign n5521 = pi75  & n3329;
  assign n5522 = n713 & n3327;
  assign n5523 = ~n5520 & ~n5521;
  assign n5524 = ~n5519 & n5523;
  assign n5525 = ~n5522 & n5524;
  assign n5526 = pi32  & n5525;
  assign n5527 = ~pi32  & ~n5525;
  assign n5528 = ~n5526 & ~n5527;
  assign n5529 = ~n5316 & ~n5320;
  assign n5530 = pi70  & n4176;
  assign n5531 = pi71  & n3938;
  assign n5532 = pi72  & n3933;
  assign n5533 = n551 & n3931;
  assign n5534 = ~n5531 & ~n5532;
  assign n5535 = ~n5530 & n5534;
  assign n5536 = ~n5533 & n5535;
  assign n5537 = pi35  & n5536;
  assign n5538 = ~pi35  & ~n5536;
  assign n5539 = ~n5537 & ~n5538;
  assign n5540 = ~n5301 & ~n5303;
  assign n5541 = pi67  & n4843;
  assign n5542 = pi68  & n4598;
  assign n5543 = pi69  & n4593;
  assign n5544 = n376 & n4591;
  assign n5545 = ~n5542 & ~n5543;
  assign n5546 = ~n5541 & n5545;
  assign n5547 = ~n5544 & n5546;
  assign n5548 = pi38  & n5547;
  assign n5549 = ~pi38  & ~n5547;
  assign n5550 = ~n5548 & ~n5549;
  assign n5551 = pi41  & ~n5024;
  assign n5552 = n5296 & n5551;
  assign n5553 = pi41  & ~n5552;
  assign n5554 = ~n287 & n5286;
  assign n5555 = pi65  & n5293;
  assign n5556 = pi66  & n5288;
  assign n5557 = ~n5023 & n5285;
  assign n5558 = ~n5292 & n5557;
  assign n5559 = pi64  & n5558;
  assign n5560 = ~n5554 & ~n5555;
  assign n5561 = ~n5556 & n5560;
  assign n5562 = ~n5559 & n5561;
  assign n5563 = ~n5553 & n5562;
  assign n5564 = n5553 & ~n5562;
  assign n5565 = ~n5563 & ~n5564;
  assign n5566 = ~n5550 & n5565;
  assign n5567 = n5550 & ~n5565;
  assign n5568 = ~n5566 & ~n5567;
  assign n5569 = ~n5540 & n5568;
  assign n5570 = n5540 & ~n5568;
  assign n5571 = ~n5569 & ~n5570;
  assign n5572 = ~n5539 & n5571;
  assign n5573 = n5539 & ~n5571;
  assign n5574 = ~n5572 & ~n5573;
  assign n5575 = ~n5529 & n5574;
  assign n5576 = n5529 & ~n5574;
  assign n5577 = ~n5575 & ~n5576;
  assign n5578 = n5528 & ~n5577;
  assign n5579 = ~n5528 & n5577;
  assign n5580 = ~n5578 & ~n5579;
  assign n5581 = ~n5518 & n5580;
  assign n5582 = n5518 & ~n5580;
  assign n5583 = ~n5581 & ~n5582;
  assign n5584 = n5517 & ~n5583;
  assign n5585 = ~n5517 & n5583;
  assign n5586 = ~n5584 & ~n5585;
  assign n5587 = ~n5507 & n5586;
  assign n5588 = n5507 & ~n5586;
  assign n5589 = ~n5587 & ~n5588;
  assign n5590 = n5506 & ~n5589;
  assign n5591 = ~n5506 & n5589;
  assign n5592 = ~n5590 & ~n5591;
  assign n5593 = ~n5496 & n5592;
  assign n5594 = n5496 & ~n5592;
  assign n5595 = ~n5593 & ~n5594;
  assign n5596 = pi82  & n2053;
  assign n5597 = pi83  & n1893;
  assign n5598 = pi84  & n1888;
  assign n5599 = n1601 & n1886;
  assign n5600 = ~n5597 & ~n5598;
  assign n5601 = ~n5596 & n5600;
  assign n5602 = ~n5599 & n5601;
  assign n5603 = pi23  & n5602;
  assign n5604 = ~pi23  & ~n5602;
  assign n5605 = ~n5603 & ~n5604;
  assign n5606 = n5595 & ~n5605;
  assign n5607 = ~n5595 & n5605;
  assign n5608 = ~n5606 & ~n5607;
  assign n5609 = n5495 & ~n5608;
  assign n5610 = ~n5495 & n5608;
  assign n5611 = ~n5609 & ~n5610;
  assign n5612 = pi85  & n1661;
  assign n5613 = pi86  & n1500;
  assign n5614 = pi87  & n1495;
  assign n5615 = n1493 & n2116;
  assign n5616 = ~n5613 & ~n5614;
  assign n5617 = ~n5612 & n5616;
  assign n5618 = ~n5615 & n5617;
  assign n5619 = pi20  & n5618;
  assign n5620 = ~pi20  & ~n5618;
  assign n5621 = ~n5619 & ~n5620;
  assign n5622 = n5611 & ~n5621;
  assign n5623 = ~n5611 & n5621;
  assign n5624 = ~n5622 & ~n5623;
  assign n5625 = ~n5494 & n5624;
  assign n5626 = n5494 & ~n5624;
  assign n5627 = ~n5625 & ~n5626;
  assign n5628 = n5493 & ~n5627;
  assign n5629 = ~n5493 & n5627;
  assign n5630 = ~n5628 & ~n5629;
  assign n5631 = ~n5483 & n5630;
  assign n5632 = n5483 & ~n5630;
  assign n5633 = ~n5631 & ~n5632;
  assign n5634 = n5482 & ~n5633;
  assign n5635 = ~n5482 & n5633;
  assign n5636 = ~n5634 & ~n5635;
  assign n5637 = ~n5472 & n5636;
  assign n5638 = n5472 & ~n5636;
  assign n5639 = ~n5637 & ~n5638;
  assign n5640 = n5471 & ~n5639;
  assign n5641 = ~n5471 & n5639;
  assign n5642 = ~n5640 & ~n5641;
  assign n5643 = ~n5461 & n5642;
  assign n5644 = n5461 & ~n5642;
  assign n5645 = ~n5643 & ~n5644;
  assign n5646 = pi97  & n528;
  assign n5647 = pi98  & n490;
  assign n5648 = pi99  & n485;
  assign n5649 = n483 & n4101;
  assign n5650 = ~n5647 & ~n5648;
  assign n5651 = ~n5646 & n5650;
  assign n5652 = ~n5649 & n5651;
  assign n5653 = pi8  & n5652;
  assign n5654 = ~pi8  & ~n5652;
  assign n5655 = ~n5653 & ~n5654;
  assign n5656 = n5645 & ~n5655;
  assign n5657 = ~n5645 & n5655;
  assign n5658 = ~n5656 & ~n5657;
  assign n5659 = ~n5460 & n5658;
  assign n5660 = n5460 & ~n5658;
  assign n5661 = ~n5659 & ~n5660;
  assign n5662 = ~n5459 & n5661;
  assign n5663 = n5459 & ~n5661;
  assign n5664 = ~n5662 & ~n5663;
  assign n5665 = n5449 & ~n5664;
  assign n5666 = ~n5449 & n5664;
  assign n5667 = ~n5665 & ~n5666;
  assign n5668 = pi105  & n269;
  assign n5669 = pi104  & n267;
  assign n5670 = pi103  & n282;
  assign n5671 = ~n5208 & ~n5210;
  assign n5672 = ~pi104  & ~pi105 ;
  assign n5673 = pi104  & pi105 ;
  assign n5674 = ~n5672 & ~n5673;
  assign n5675 = ~n5671 & n5674;
  assign n5676 = n5671 & ~n5674;
  assign n5677 = ~n5675 & ~n5676;
  assign n5678 = n262 & n5677;
  assign n5679 = ~n5668 & ~n5669;
  assign n5680 = ~n5670 & n5679;
  assign n5681 = ~n5678 & n5680;
  assign n5682 = pi2  & n5681;
  assign n5683 = ~pi2  & ~n5681;
  assign n5684 = ~n5682 & ~n5683;
  assign n5685 = ~n5667 & n5684;
  assign n5686 = n5667 & ~n5684;
  assign n5687 = ~n5685 & ~n5686;
  assign n5688 = ~n5448 & n5687;
  assign n5689 = n5448 & ~n5687;
  assign po41  = ~n5688 & ~n5689;
  assign n5691 = ~n5686 & ~n5688;
  assign n5692 = pi106  & n269;
  assign n5693 = pi105  & n267;
  assign n5694 = pi104  & n282;
  assign n5695 = ~n5673 & ~n5675;
  assign n5696 = ~pi105  & ~pi106 ;
  assign n5697 = pi105  & pi106 ;
  assign n5698 = ~n5696 & ~n5697;
  assign n5699 = ~n5695 & n5698;
  assign n5700 = n5695 & ~n5698;
  assign n5701 = ~n5699 & ~n5700;
  assign n5702 = n262 & n5701;
  assign n5703 = ~n5692 & ~n5693;
  assign n5704 = ~n5694 & n5703;
  assign n5705 = ~n5702 & n5704;
  assign n5706 = pi2  & n5705;
  assign n5707 = ~pi2  & ~n5705;
  assign n5708 = ~n5706 & ~n5707;
  assign n5709 = ~n5662 & ~n5666;
  assign n5710 = pi101  & n391;
  assign n5711 = pi102  & n353;
  assign n5712 = pi103  & n348;
  assign n5713 = n346 & n5188;
  assign n5714 = ~n5711 & ~n5712;
  assign n5715 = ~n5710 & n5714;
  assign n5716 = ~n5713 & n5715;
  assign n5717 = pi5  & n5716;
  assign n5718 = ~pi5  & ~n5716;
  assign n5719 = ~n5717 & ~n5718;
  assign n5720 = ~n5656 & ~n5659;
  assign n5721 = pi98  & n528;
  assign n5722 = pi99  & n490;
  assign n5723 = pi100  & n485;
  assign n5724 = n483 & n4501;
  assign n5725 = ~n5722 & ~n5723;
  assign n5726 = ~n5721 & n5725;
  assign n5727 = ~n5724 & n5726;
  assign n5728 = pi8  & n5727;
  assign n5729 = ~pi8  & ~n5727;
  assign n5730 = ~n5728 & ~n5729;
  assign n5731 = ~n5641 & ~n5643;
  assign n5732 = ~n5635 & ~n5637;
  assign n5733 = pi92  & n1006;
  assign n5734 = pi93  & n897;
  assign n5735 = pi94  & n892;
  assign n5736 = n890 & n3280;
  assign n5737 = ~n5734 & ~n5735;
  assign n5738 = ~n5733 & n5737;
  assign n5739 = ~n5736 & n5738;
  assign n5740 = pi14  & n5739;
  assign n5741 = ~pi14  & ~n5739;
  assign n5742 = ~n5740 & ~n5741;
  assign n5743 = ~n5629 & ~n5631;
  assign n5744 = ~n5622 & ~n5625;
  assign n5745 = ~n5606 & ~n5610;
  assign n5746 = ~n5591 & ~n5593;
  assign n5747 = pi80  & n2510;
  assign n5748 = pi81  & n2342;
  assign n5749 = pi82  & n2337;
  assign n5750 = n1450 & n2335;
  assign n5751 = ~n5748 & ~n5749;
  assign n5752 = ~n5747 & n5751;
  assign n5753 = ~n5750 & n5752;
  assign n5754 = pi26  & n5753;
  assign n5755 = ~pi26  & ~n5753;
  assign n5756 = ~n5754 & ~n5755;
  assign n5757 = ~n5585 & ~n5587;
  assign n5758 = pi77  & n3011;
  assign n5759 = pi78  & n2809;
  assign n5760 = pi79  & n2804;
  assign n5761 = n1048 & n2802;
  assign n5762 = ~n5759 & ~n5760;
  assign n5763 = ~n5758 & n5762;
  assign n5764 = ~n5761 & n5763;
  assign n5765 = pi29  & n5764;
  assign n5766 = ~pi29  & ~n5764;
  assign n5767 = ~n5765 & ~n5766;
  assign n5768 = ~n5579 & ~n5581;
  assign n5769 = pi74  & n3553;
  assign n5770 = pi75  & n3334;
  assign n5771 = pi76  & n3329;
  assign n5772 = n841 & n3327;
  assign n5773 = ~n5770 & ~n5771;
  assign n5774 = ~n5769 & n5773;
  assign n5775 = ~n5772 & n5774;
  assign n5776 = pi32  & n5775;
  assign n5777 = ~pi32  & ~n5775;
  assign n5778 = ~n5776 & ~n5777;
  assign n5779 = ~n5572 & ~n5575;
  assign n5780 = ~n5566 & ~n5569;
  assign n5781 = pi65  & n5558;
  assign n5782 = pi66  & n5293;
  assign n5783 = pi67  & n5288;
  assign n5784 = n305 & n5286;
  assign n5785 = ~n5782 & ~n5783;
  assign n5786 = ~n5781 & n5785;
  assign n5787 = ~n5784 & n5786;
  assign n5788 = pi41  & n5787;
  assign n5789 = ~pi41  & ~n5787;
  assign n5790 = ~n5788 & ~n5789;
  assign n5791 = ~pi41  & ~pi42 ;
  assign n5792 = pi41  & pi42 ;
  assign n5793 = ~n5791 & ~n5792;
  assign n5794 = pi64  & n5793;
  assign n5795 = n5552 & n5562;
  assign n5796 = n5794 & n5795;
  assign n5797 = ~n5794 & ~n5795;
  assign n5798 = ~n5796 & ~n5797;
  assign n5799 = ~n5790 & n5798;
  assign n5800 = n5790 & ~n5798;
  assign n5801 = ~n5799 & ~n5800;
  assign n5802 = pi68  & n4843;
  assign n5803 = pi69  & n4598;
  assign n5804 = pi70  & n4593;
  assign n5805 = n415 & n4591;
  assign n5806 = ~n5803 & ~n5804;
  assign n5807 = ~n5802 & n5806;
  assign n5808 = ~n5805 & n5807;
  assign n5809 = pi38  & n5808;
  assign n5810 = ~pi38  & ~n5808;
  assign n5811 = ~n5809 & ~n5810;
  assign n5812 = n5801 & ~n5811;
  assign n5813 = ~n5801 & n5811;
  assign n5814 = ~n5812 & ~n5813;
  assign n5815 = n5780 & ~n5814;
  assign n5816 = ~n5780 & n5814;
  assign n5817 = ~n5815 & ~n5816;
  assign n5818 = pi71  & n4176;
  assign n5819 = pi72  & n3938;
  assign n5820 = pi73  & n3933;
  assign n5821 = n613 & n3931;
  assign n5822 = ~n5819 & ~n5820;
  assign n5823 = ~n5818 & n5822;
  assign n5824 = ~n5821 & n5823;
  assign n5825 = pi35  & n5824;
  assign n5826 = ~pi35  & ~n5824;
  assign n5827 = ~n5825 & ~n5826;
  assign n5828 = ~n5817 & n5827;
  assign n5829 = n5817 & ~n5827;
  assign n5830 = ~n5828 & ~n5829;
  assign n5831 = ~n5779 & n5830;
  assign n5832 = n5779 & ~n5830;
  assign n5833 = ~n5831 & ~n5832;
  assign n5834 = ~n5778 & n5833;
  assign n5835 = n5778 & ~n5833;
  assign n5836 = ~n5834 & ~n5835;
  assign n5837 = ~n5768 & n5836;
  assign n5838 = n5768 & ~n5836;
  assign n5839 = ~n5837 & ~n5838;
  assign n5840 = ~n5767 & n5839;
  assign n5841 = n5767 & ~n5839;
  assign n5842 = ~n5840 & ~n5841;
  assign n5843 = ~n5757 & n5842;
  assign n5844 = n5757 & ~n5842;
  assign n5845 = ~n5843 & ~n5844;
  assign n5846 = ~n5756 & n5845;
  assign n5847 = n5756 & ~n5845;
  assign n5848 = ~n5846 & ~n5847;
  assign n5849 = ~n5746 & n5848;
  assign n5850 = n5746 & ~n5848;
  assign n5851 = ~n5849 & ~n5850;
  assign n5852 = pi83  & n2053;
  assign n5853 = pi84  & n1893;
  assign n5854 = pi85  & n1888;
  assign n5855 = n1831 & n1886;
  assign n5856 = ~n5853 & ~n5854;
  assign n5857 = ~n5852 & n5856;
  assign n5858 = ~n5855 & n5857;
  assign n5859 = pi23  & n5858;
  assign n5860 = ~pi23  & ~n5858;
  assign n5861 = ~n5859 & ~n5860;
  assign n5862 = n5851 & ~n5861;
  assign n5863 = ~n5851 & n5861;
  assign n5864 = ~n5862 & ~n5863;
  assign n5865 = n5745 & ~n5864;
  assign n5866 = ~n5745 & n5864;
  assign n5867 = ~n5865 & ~n5866;
  assign n5868 = pi86  & n1661;
  assign n5869 = pi87  & n1500;
  assign n5870 = pi88  & n1495;
  assign n5871 = n1493 & n2140;
  assign n5872 = ~n5869 & ~n5870;
  assign n5873 = ~n5868 & n5872;
  assign n5874 = ~n5871 & n5873;
  assign n5875 = pi20  & n5874;
  assign n5876 = ~pi20  & ~n5874;
  assign n5877 = ~n5875 & ~n5876;
  assign n5878 = ~n5867 & n5877;
  assign n5879 = n5867 & ~n5877;
  assign n5880 = ~n5878 & ~n5879;
  assign n5881 = ~n5744 & n5880;
  assign n5882 = n5744 & ~n5880;
  assign n5883 = ~n5881 & ~n5882;
  assign n5884 = pi89  & n1296;
  assign n5885 = pi90  & n1207;
  assign n5886 = pi91  & n1202;
  assign n5887 = n1200 & n2746;
  assign n5888 = ~n5885 & ~n5886;
  assign n5889 = ~n5884 & n5888;
  assign n5890 = ~n5887 & n5889;
  assign n5891 = pi17  & n5890;
  assign n5892 = ~pi17  & ~n5890;
  assign n5893 = ~n5891 & ~n5892;
  assign n5894 = n5883 & ~n5893;
  assign n5895 = ~n5883 & n5893;
  assign n5896 = ~n5894 & ~n5895;
  assign n5897 = ~n5743 & n5896;
  assign n5898 = n5743 & ~n5896;
  assign n5899 = ~n5897 & ~n5898;
  assign n5900 = ~n5742 & n5899;
  assign n5901 = n5742 & ~n5899;
  assign n5902 = ~n5900 & ~n5901;
  assign n5903 = ~n5732 & n5902;
  assign n5904 = n5732 & ~n5902;
  assign n5905 = ~n5903 & ~n5904;
  assign n5906 = pi95  & n750;
  assign n5907 = pi96  & n651;
  assign n5908 = pi97  & n646;
  assign n5909 = n644 & n3691;
  assign n5910 = ~n5907 & ~n5908;
  assign n5911 = ~n5906 & n5910;
  assign n5912 = ~n5909 & n5911;
  assign n5913 = pi11  & n5912;
  assign n5914 = ~pi11  & ~n5912;
  assign n5915 = ~n5913 & ~n5914;
  assign n5916 = n5905 & ~n5915;
  assign n5917 = ~n5905 & n5915;
  assign n5918 = ~n5916 & ~n5917;
  assign n5919 = ~n5731 & n5918;
  assign n5920 = n5731 & ~n5918;
  assign n5921 = ~n5919 & ~n5920;
  assign n5922 = n5730 & ~n5921;
  assign n5923 = ~n5730 & n5921;
  assign n5924 = ~n5922 & ~n5923;
  assign n5925 = ~n5720 & n5924;
  assign n5926 = n5720 & ~n5924;
  assign n5927 = ~n5925 & ~n5926;
  assign n5928 = ~n5719 & n5927;
  assign n5929 = n5719 & ~n5927;
  assign n5930 = ~n5928 & ~n5929;
  assign n5931 = ~n5709 & n5930;
  assign n5932 = n5709 & ~n5930;
  assign n5933 = ~n5931 & ~n5932;
  assign n5934 = ~n5708 & n5933;
  assign n5935 = n5708 & ~n5933;
  assign n5936 = ~n5934 & ~n5935;
  assign n5937 = ~n5691 & n5936;
  assign n5938 = n5691 & ~n5936;
  assign po42  = ~n5937 & ~n5938;
  assign n5940 = ~n5934 & ~n5937;
  assign n5941 = ~n5928 & ~n5931;
  assign n5942 = pi102  & n391;
  assign n5943 = pi103  & n353;
  assign n5944 = pi104  & n348;
  assign n5945 = n346 & n5212;
  assign n5946 = ~n5943 & ~n5944;
  assign n5947 = ~n5942 & n5946;
  assign n5948 = ~n5945 & n5947;
  assign n5949 = pi5  & n5948;
  assign n5950 = ~pi5  & ~n5948;
  assign n5951 = ~n5949 & ~n5950;
  assign n5952 = ~n5923 & ~n5925;
  assign n5953 = ~n5916 & ~n5919;
  assign n5954 = ~n5900 & ~n5903;
  assign n5955 = pi93  & n1006;
  assign n5956 = pi94  & n897;
  assign n5957 = pi95  & n892;
  assign n5958 = n890 & n3475;
  assign n5959 = ~n5956 & ~n5957;
  assign n5960 = ~n5955 & n5959;
  assign n5961 = ~n5958 & n5960;
  assign n5962 = pi14  & n5961;
  assign n5963 = ~pi14  & ~n5961;
  assign n5964 = ~n5962 & ~n5963;
  assign n5965 = ~n5894 & ~n5897;
  assign n5966 = pi90  & n1296;
  assign n5967 = pi91  & n1207;
  assign n5968 = pi92  & n1202;
  assign n5969 = n1200 & n2924;
  assign n5970 = ~n5967 & ~n5968;
  assign n5971 = ~n5966 & n5970;
  assign n5972 = ~n5969 & n5971;
  assign n5973 = pi17  & n5972;
  assign n5974 = ~pi17  & ~n5972;
  assign n5975 = ~n5973 & ~n5974;
  assign n5976 = ~n5879 & ~n5881;
  assign n5977 = ~n5862 & ~n5866;
  assign n5978 = ~n5846 & ~n5849;
  assign n5979 = ~n5840 & ~n5843;
  assign n5980 = ~n5834 & ~n5837;
  assign n5981 = pi75  & n3553;
  assign n5982 = pi76  & n3334;
  assign n5983 = pi77  & n3329;
  assign n5984 = n865 & n3327;
  assign n5985 = ~n5982 & ~n5983;
  assign n5986 = ~n5981 & n5985;
  assign n5987 = ~n5984 & n5986;
  assign n5988 = pi32  & n5987;
  assign n5989 = ~pi32  & ~n5987;
  assign n5990 = ~n5988 & ~n5989;
  assign n5991 = ~n5829 & ~n5831;
  assign n5992 = ~n5812 & ~n5816;
  assign n5993 = ~n5796 & ~n5799;
  assign n5994 = pi66  & n5558;
  assign n5995 = pi67  & n5293;
  assign n5996 = pi68  & n5288;
  assign n5997 = n334 & n5286;
  assign n5998 = ~n5995 & ~n5996;
  assign n5999 = ~n5994 & n5998;
  assign n6000 = ~n5997 & n5999;
  assign n6001 = pi41  & n6000;
  assign n6002 = ~pi41  & ~n6000;
  assign n6003 = ~n6001 & ~n6002;
  assign n6004 = pi44  & n5794;
  assign n6005 = ~pi43  & ~pi44 ;
  assign n6006 = pi43  & pi44 ;
  assign n6007 = ~n6005 & ~n6006;
  assign n6008 = n5793 & n6007;
  assign n6009 = n265 & n6008;
  assign n6010 = n5793 & ~n6007;
  assign n6011 = pi65  & n6010;
  assign n6012 = ~pi42  & ~pi43 ;
  assign n6013 = pi42  & pi43 ;
  assign n6014 = ~n6012 & ~n6013;
  assign n6015 = ~n5793 & n6014;
  assign n6016 = pi64  & n6015;
  assign n6017 = ~n6009 & ~n6011;
  assign n6018 = ~n6016 & n6017;
  assign n6019 = n6004 & ~n6018;
  assign n6020 = ~n6004 & n6018;
  assign n6021 = ~n6019 & ~n6020;
  assign n6022 = n6003 & ~n6021;
  assign n6023 = ~n6003 & n6021;
  assign n6024 = ~n6022 & ~n6023;
  assign n6025 = ~n5993 & n6024;
  assign n6026 = n5993 & ~n6024;
  assign n6027 = ~n6025 & ~n6026;
  assign n6028 = pi69  & n4843;
  assign n6029 = pi70  & n4598;
  assign n6030 = pi71  & n4593;
  assign n6031 = n460 & n4591;
  assign n6032 = ~n6029 & ~n6030;
  assign n6033 = ~n6028 & n6032;
  assign n6034 = ~n6031 & n6033;
  assign n6035 = pi38  & n6034;
  assign n6036 = ~pi38  & ~n6034;
  assign n6037 = ~n6035 & ~n6036;
  assign n6038 = n6027 & ~n6037;
  assign n6039 = ~n6027 & n6037;
  assign n6040 = ~n6038 & ~n6039;
  assign n6041 = n5992 & ~n6040;
  assign n6042 = ~n5992 & n6040;
  assign n6043 = ~n6041 & ~n6042;
  assign n6044 = pi72  & n4176;
  assign n6045 = pi73  & n3938;
  assign n6046 = pi74  & n3933;
  assign n6047 = n689 & n3931;
  assign n6048 = ~n6045 & ~n6046;
  assign n6049 = ~n6044 & n6048;
  assign n6050 = ~n6047 & n6049;
  assign n6051 = pi35  & n6050;
  assign n6052 = ~pi35  & ~n6050;
  assign n6053 = ~n6051 & ~n6052;
  assign n6054 = n6043 & ~n6053;
  assign n6055 = ~n6043 & n6053;
  assign n6056 = ~n6054 & ~n6055;
  assign n6057 = ~n5991 & n6056;
  assign n6058 = n5991 & ~n6056;
  assign n6059 = ~n6057 & ~n6058;
  assign n6060 = n5990 & ~n6059;
  assign n6061 = ~n5990 & n6059;
  assign n6062 = ~n6060 & ~n6061;
  assign n6063 = ~n5980 & n6062;
  assign n6064 = n5980 & ~n6062;
  assign n6065 = ~n6063 & ~n6064;
  assign n6066 = pi78  & n3011;
  assign n6067 = pi79  & n2809;
  assign n6068 = pi80  & n2804;
  assign n6069 = n1144 & n2802;
  assign n6070 = ~n6067 & ~n6068;
  assign n6071 = ~n6066 & n6070;
  assign n6072 = ~n6069 & n6071;
  assign n6073 = pi29  & n6072;
  assign n6074 = ~pi29  & ~n6072;
  assign n6075 = ~n6073 & ~n6074;
  assign n6076 = n6065 & ~n6075;
  assign n6077 = ~n6065 & n6075;
  assign n6078 = ~n6076 & ~n6077;
  assign n6079 = n5979 & ~n6078;
  assign n6080 = ~n5979 & n6078;
  assign n6081 = ~n6079 & ~n6080;
  assign n6082 = pi81  & n2510;
  assign n6083 = pi82  & n2342;
  assign n6084 = pi83  & n2337;
  assign n6085 = n1577 & n2335;
  assign n6086 = ~n6083 & ~n6084;
  assign n6087 = ~n6082 & n6086;
  assign n6088 = ~n6085 & n6087;
  assign n6089 = pi26  & n6088;
  assign n6090 = ~pi26  & ~n6088;
  assign n6091 = ~n6089 & ~n6090;
  assign n6092 = n6081 & ~n6091;
  assign n6093 = ~n6081 & n6091;
  assign n6094 = ~n6092 & ~n6093;
  assign n6095 = n5978 & ~n6094;
  assign n6096 = ~n5978 & n6094;
  assign n6097 = ~n6095 & ~n6096;
  assign n6098 = pi84  & n2053;
  assign n6099 = pi85  & n1893;
  assign n6100 = pi86  & n1888;
  assign n6101 = n1886 & n1975;
  assign n6102 = ~n6099 & ~n6100;
  assign n6103 = ~n6098 & n6102;
  assign n6104 = ~n6101 & n6103;
  assign n6105 = pi23  & n6104;
  assign n6106 = ~pi23  & ~n6104;
  assign n6107 = ~n6105 & ~n6106;
  assign n6108 = n6097 & ~n6107;
  assign n6109 = ~n6097 & n6107;
  assign n6110 = ~n6108 & ~n6109;
  assign n6111 = n5977 & ~n6110;
  assign n6112 = ~n5977 & n6110;
  assign n6113 = ~n6111 & ~n6112;
  assign n6114 = pi87  & n1661;
  assign n6115 = pi88  & n1500;
  assign n6116 = pi89  & n1495;
  assign n6117 = n1493 & n2287;
  assign n6118 = ~n6115 & ~n6116;
  assign n6119 = ~n6114 & n6118;
  assign n6120 = ~n6117 & n6119;
  assign n6121 = pi20  & n6120;
  assign n6122 = ~pi20  & ~n6120;
  assign n6123 = ~n6121 & ~n6122;
  assign n6124 = n6113 & ~n6123;
  assign n6125 = ~n6113 & n6123;
  assign n6126 = ~n6124 & ~n6125;
  assign n6127 = ~n5976 & n6126;
  assign n6128 = n5976 & ~n6126;
  assign n6129 = ~n6127 & ~n6128;
  assign n6130 = ~n5975 & n6129;
  assign n6131 = n5975 & ~n6129;
  assign n6132 = ~n6130 & ~n6131;
  assign n6133 = ~n5965 & n6132;
  assign n6134 = n5965 & ~n6132;
  assign n6135 = ~n6133 & ~n6134;
  assign n6136 = n5964 & ~n6135;
  assign n6137 = ~n5964 & n6135;
  assign n6138 = ~n6136 & ~n6137;
  assign n6139 = ~n5954 & n6138;
  assign n6140 = n5954 & ~n6138;
  assign n6141 = ~n6139 & ~n6140;
  assign n6142 = pi96  & n750;
  assign n6143 = pi97  & n651;
  assign n6144 = pi98  & n646;
  assign n6145 = n644 & n3889;
  assign n6146 = ~n6143 & ~n6144;
  assign n6147 = ~n6142 & n6146;
  assign n6148 = ~n6145 & n6147;
  assign n6149 = pi11  & n6148;
  assign n6150 = ~pi11  & ~n6148;
  assign n6151 = ~n6149 & ~n6150;
  assign n6152 = n6141 & ~n6151;
  assign n6153 = ~n6141 & n6151;
  assign n6154 = ~n6152 & ~n6153;
  assign n6155 = n5953 & ~n6154;
  assign n6156 = ~n5953 & n6154;
  assign n6157 = ~n6155 & ~n6156;
  assign n6158 = pi99  & n528;
  assign n6159 = pi100  & n490;
  assign n6160 = pi101  & n485;
  assign n6161 = n483 & n4730;
  assign n6162 = ~n6159 & ~n6160;
  assign n6163 = ~n6158 & n6162;
  assign n6164 = ~n6161 & n6163;
  assign n6165 = pi8  & n6164;
  assign n6166 = ~pi8  & ~n6164;
  assign n6167 = ~n6165 & ~n6166;
  assign n6168 = n6157 & ~n6167;
  assign n6169 = ~n6157 & n6167;
  assign n6170 = ~n6168 & ~n6169;
  assign n6171 = ~n5952 & n6170;
  assign n6172 = n5952 & ~n6170;
  assign n6173 = ~n6171 & ~n6172;
  assign n6174 = n5951 & ~n6173;
  assign n6175 = ~n5951 & n6173;
  assign n6176 = ~n6174 & ~n6175;
  assign n6177 = ~n5941 & n6176;
  assign n6178 = n5941 & ~n6176;
  assign n6179 = ~n6177 & ~n6178;
  assign n6180 = pi107  & n269;
  assign n6181 = pi106  & n267;
  assign n6182 = pi105  & n282;
  assign n6183 = ~n5697 & ~n5699;
  assign n6184 = ~pi106  & ~pi107 ;
  assign n6185 = pi106  & pi107 ;
  assign n6186 = ~n6184 & ~n6185;
  assign n6187 = ~n6183 & n6186;
  assign n6188 = n6183 & ~n6186;
  assign n6189 = ~n6187 & ~n6188;
  assign n6190 = n262 & n6189;
  assign n6191 = ~n6180 & ~n6181;
  assign n6192 = ~n6182 & n6191;
  assign n6193 = ~n6190 & n6192;
  assign n6194 = pi2  & n6193;
  assign n6195 = ~pi2  & ~n6193;
  assign n6196 = ~n6194 & ~n6195;
  assign n6197 = n6179 & ~n6196;
  assign n6198 = ~n6179 & n6196;
  assign n6199 = ~n6197 & ~n6198;
  assign n6200 = ~n5940 & n6199;
  assign n6201 = n5940 & ~n6199;
  assign po43  = ~n6200 & ~n6201;
  assign n6203 = ~n6197 & ~n6200;
  assign n6204 = pi108  & n269;
  assign n6205 = pi107  & n267;
  assign n6206 = pi106  & n282;
  assign n6207 = ~n6185 & ~n6187;
  assign n6208 = ~pi107  & ~pi108 ;
  assign n6209 = pi107  & pi108 ;
  assign n6210 = ~n6208 & ~n6209;
  assign n6211 = ~n6207 & n6210;
  assign n6212 = n6207 & ~n6210;
  assign n6213 = ~n6211 & ~n6212;
  assign n6214 = n262 & n6213;
  assign n6215 = ~n6204 & ~n6205;
  assign n6216 = ~n6206 & n6215;
  assign n6217 = ~n6214 & n6216;
  assign n6218 = pi2  & n6217;
  assign n6219 = ~pi2  & ~n6217;
  assign n6220 = ~n6218 & ~n6219;
  assign n6221 = ~n6175 & ~n6177;
  assign n6222 = pi103  & n391;
  assign n6223 = pi104  & n353;
  assign n6224 = pi105  & n348;
  assign n6225 = n346 & n5677;
  assign n6226 = ~n6223 & ~n6224;
  assign n6227 = ~n6222 & n6226;
  assign n6228 = ~n6225 & n6227;
  assign n6229 = pi5  & n6228;
  assign n6230 = ~pi5  & ~n6228;
  assign n6231 = ~n6229 & ~n6230;
  assign n6232 = ~n6168 & ~n6171;
  assign n6233 = ~n6152 & ~n6156;
  assign n6234 = ~n6137 & ~n6139;
  assign n6235 = pi94  & n1006;
  assign n6236 = pi95  & n897;
  assign n6237 = pi96  & n892;
  assign n6238 = n890 & n3499;
  assign n6239 = ~n6236 & ~n6237;
  assign n6240 = ~n6235 & n6239;
  assign n6241 = ~n6238 & n6240;
  assign n6242 = pi14  & n6241;
  assign n6243 = ~pi14  & ~n6241;
  assign n6244 = ~n6242 & ~n6243;
  assign n6245 = ~n6130 & ~n6133;
  assign n6246 = pi91  & n1296;
  assign n6247 = pi92  & n1207;
  assign n6248 = pi93  & n1202;
  assign n6249 = n1200 & n2948;
  assign n6250 = ~n6247 & ~n6248;
  assign n6251 = ~n6246 & n6250;
  assign n6252 = ~n6249 & n6251;
  assign n6253 = pi17  & n6252;
  assign n6254 = ~pi17  & ~n6252;
  assign n6255 = ~n6253 & ~n6254;
  assign n6256 = ~n6124 & ~n6127;
  assign n6257 = pi88  & n1661;
  assign n6258 = pi89  & n1500;
  assign n6259 = pi90  & n1495;
  assign n6260 = n1493 & n2448;
  assign n6261 = ~n6258 & ~n6259;
  assign n6262 = ~n6257 & n6261;
  assign n6263 = ~n6260 & n6262;
  assign n6264 = pi20  & n6263;
  assign n6265 = ~pi20  & ~n6263;
  assign n6266 = ~n6264 & ~n6265;
  assign n6267 = ~n6108 & ~n6112;
  assign n6268 = ~n6092 & ~n6096;
  assign n6269 = ~n6076 & ~n6080;
  assign n6270 = pi79  & n3011;
  assign n6271 = pi80  & n2809;
  assign n6272 = pi81  & n2804;
  assign n6273 = n1337 & n2802;
  assign n6274 = ~n6271 & ~n6272;
  assign n6275 = ~n6270 & n6274;
  assign n6276 = ~n6273 & n6275;
  assign n6277 = pi29  & n6276;
  assign n6278 = ~pi29  & ~n6276;
  assign n6279 = ~n6277 & ~n6278;
  assign n6280 = ~n6061 & ~n6063;
  assign n6281 = pi76  & n3553;
  assign n6282 = pi77  & n3334;
  assign n6283 = pi78  & n3329;
  assign n6284 = n958 & n3327;
  assign n6285 = ~n6282 & ~n6283;
  assign n6286 = ~n6281 & n6285;
  assign n6287 = ~n6284 & n6286;
  assign n6288 = pi32  & n6287;
  assign n6289 = ~pi32  & ~n6287;
  assign n6290 = ~n6288 & ~n6289;
  assign n6291 = ~n6054 & ~n6057;
  assign n6292 = pi73  & n4176;
  assign n6293 = pi74  & n3938;
  assign n6294 = pi75  & n3933;
  assign n6295 = n713 & n3931;
  assign n6296 = ~n6293 & ~n6294;
  assign n6297 = ~n6292 & n6296;
  assign n6298 = ~n6295 & n6297;
  assign n6299 = pi35  & n6298;
  assign n6300 = ~pi35  & ~n6298;
  assign n6301 = ~n6299 & ~n6300;
  assign n6302 = ~n6038 & ~n6042;
  assign n6303 = pi70  & n4843;
  assign n6304 = pi71  & n4598;
  assign n6305 = pi72  & n4593;
  assign n6306 = n551 & n4591;
  assign n6307 = ~n6304 & ~n6305;
  assign n6308 = ~n6303 & n6307;
  assign n6309 = ~n6306 & n6308;
  assign n6310 = pi38  & n6309;
  assign n6311 = ~pi38  & ~n6309;
  assign n6312 = ~n6310 & ~n6311;
  assign n6313 = ~n6023 & ~n6025;
  assign n6314 = pi67  & n5558;
  assign n6315 = pi68  & n5293;
  assign n6316 = pi69  & n5288;
  assign n6317 = n376 & n5286;
  assign n6318 = ~n6315 & ~n6316;
  assign n6319 = ~n6314 & n6318;
  assign n6320 = ~n6317 & n6319;
  assign n6321 = pi41  & n6320;
  assign n6322 = ~pi41  & ~n6320;
  assign n6323 = ~n6321 & ~n6322;
  assign n6324 = pi44  & ~n5794;
  assign n6325 = n6018 & n6324;
  assign n6326 = pi44  & ~n6325;
  assign n6327 = ~n287 & n6008;
  assign n6328 = pi65  & n6015;
  assign n6329 = pi66  & n6010;
  assign n6330 = ~n5793 & n6007;
  assign n6331 = ~n6014 & n6330;
  assign n6332 = pi64  & n6331;
  assign n6333 = ~n6327 & ~n6328;
  assign n6334 = ~n6329 & n6333;
  assign n6335 = ~n6332 & n6334;
  assign n6336 = ~n6326 & n6335;
  assign n6337 = n6326 & ~n6335;
  assign n6338 = ~n6336 & ~n6337;
  assign n6339 = ~n6323 & n6338;
  assign n6340 = n6323 & ~n6338;
  assign n6341 = ~n6339 & ~n6340;
  assign n6342 = ~n6313 & n6341;
  assign n6343 = n6313 & ~n6341;
  assign n6344 = ~n6342 & ~n6343;
  assign n6345 = ~n6312 & n6344;
  assign n6346 = n6312 & ~n6344;
  assign n6347 = ~n6345 & ~n6346;
  assign n6348 = ~n6302 & n6347;
  assign n6349 = n6302 & ~n6347;
  assign n6350 = ~n6348 & ~n6349;
  assign n6351 = n6301 & ~n6350;
  assign n6352 = ~n6301 & n6350;
  assign n6353 = ~n6351 & ~n6352;
  assign n6354 = ~n6291 & n6353;
  assign n6355 = n6291 & ~n6353;
  assign n6356 = ~n6354 & ~n6355;
  assign n6357 = n6290 & ~n6356;
  assign n6358 = ~n6290 & n6356;
  assign n6359 = ~n6357 & ~n6358;
  assign n6360 = ~n6280 & n6359;
  assign n6361 = n6280 & ~n6359;
  assign n6362 = ~n6360 & ~n6361;
  assign n6363 = n6279 & ~n6362;
  assign n6364 = ~n6279 & n6362;
  assign n6365 = ~n6363 & ~n6364;
  assign n6366 = ~n6269 & n6365;
  assign n6367 = n6269 & ~n6365;
  assign n6368 = ~n6366 & ~n6367;
  assign n6369 = pi82  & n2510;
  assign n6370 = pi83  & n2342;
  assign n6371 = pi84  & n2337;
  assign n6372 = n1601 & n2335;
  assign n6373 = ~n6370 & ~n6371;
  assign n6374 = ~n6369 & n6373;
  assign n6375 = ~n6372 & n6374;
  assign n6376 = pi26  & n6375;
  assign n6377 = ~pi26  & ~n6375;
  assign n6378 = ~n6376 & ~n6377;
  assign n6379 = n6368 & ~n6378;
  assign n6380 = ~n6368 & n6378;
  assign n6381 = ~n6379 & ~n6380;
  assign n6382 = n6268 & ~n6381;
  assign n6383 = ~n6268 & n6381;
  assign n6384 = ~n6382 & ~n6383;
  assign n6385 = pi85  & n2053;
  assign n6386 = pi86  & n1893;
  assign n6387 = pi87  & n1888;
  assign n6388 = n1886 & n2116;
  assign n6389 = ~n6386 & ~n6387;
  assign n6390 = ~n6385 & n6389;
  assign n6391 = ~n6388 & n6390;
  assign n6392 = pi23  & n6391;
  assign n6393 = ~pi23  & ~n6391;
  assign n6394 = ~n6392 & ~n6393;
  assign n6395 = n6384 & ~n6394;
  assign n6396 = ~n6384 & n6394;
  assign n6397 = ~n6395 & ~n6396;
  assign n6398 = ~n6267 & n6397;
  assign n6399 = n6267 & ~n6397;
  assign n6400 = ~n6398 & ~n6399;
  assign n6401 = n6266 & ~n6400;
  assign n6402 = ~n6266 & n6400;
  assign n6403 = ~n6401 & ~n6402;
  assign n6404 = ~n6256 & n6403;
  assign n6405 = n6256 & ~n6403;
  assign n6406 = ~n6404 & ~n6405;
  assign n6407 = n6255 & ~n6406;
  assign n6408 = ~n6255 & n6406;
  assign n6409 = ~n6407 & ~n6408;
  assign n6410 = ~n6245 & n6409;
  assign n6411 = n6245 & ~n6409;
  assign n6412 = ~n6410 & ~n6411;
  assign n6413 = n6244 & ~n6412;
  assign n6414 = ~n6244 & n6412;
  assign n6415 = ~n6413 & ~n6414;
  assign n6416 = ~n6234 & n6415;
  assign n6417 = n6234 & ~n6415;
  assign n6418 = ~n6416 & ~n6417;
  assign n6419 = pi97  & n750;
  assign n6420 = pi98  & n651;
  assign n6421 = pi99  & n646;
  assign n6422 = n644 & n4101;
  assign n6423 = ~n6420 & ~n6421;
  assign n6424 = ~n6419 & n6423;
  assign n6425 = ~n6422 & n6424;
  assign n6426 = pi11  & n6425;
  assign n6427 = ~pi11  & ~n6425;
  assign n6428 = ~n6426 & ~n6427;
  assign n6429 = n6418 & ~n6428;
  assign n6430 = ~n6418 & n6428;
  assign n6431 = ~n6429 & ~n6430;
  assign n6432 = n6233 & ~n6431;
  assign n6433 = ~n6233 & n6431;
  assign n6434 = ~n6432 & ~n6433;
  assign n6435 = pi100  & n528;
  assign n6436 = pi101  & n490;
  assign n6437 = pi102  & n485;
  assign n6438 = n483 & n4956;
  assign n6439 = ~n6436 & ~n6437;
  assign n6440 = ~n6435 & n6439;
  assign n6441 = ~n6438 & n6440;
  assign n6442 = pi8  & n6441;
  assign n6443 = ~pi8  & ~n6441;
  assign n6444 = ~n6442 & ~n6443;
  assign n6445 = n6434 & ~n6444;
  assign n6446 = ~n6434 & n6444;
  assign n6447 = ~n6445 & ~n6446;
  assign n6448 = ~n6232 & n6447;
  assign n6449 = n6232 & ~n6447;
  assign n6450 = ~n6448 & ~n6449;
  assign n6451 = ~n6231 & n6450;
  assign n6452 = n6231 & ~n6450;
  assign n6453 = ~n6451 & ~n6452;
  assign n6454 = ~n6221 & n6453;
  assign n6455 = n6221 & ~n6453;
  assign n6456 = ~n6454 & ~n6455;
  assign n6457 = ~n6220 & n6456;
  assign n6458 = n6220 & ~n6456;
  assign n6459 = ~n6457 & ~n6458;
  assign n6460 = ~n6203 & n6459;
  assign n6461 = n6203 & ~n6459;
  assign po44  = ~n6460 & ~n6461;
  assign n6463 = ~n6457 & ~n6460;
  assign n6464 = ~n6451 & ~n6454;
  assign n6465 = ~n6445 & ~n6448;
  assign n6466 = ~n6429 & ~n6433;
  assign n6467 = pi98  & n750;
  assign n6468 = pi99  & n651;
  assign n6469 = pi100  & n646;
  assign n6470 = n644 & n4501;
  assign n6471 = ~n6468 & ~n6469;
  assign n6472 = ~n6467 & n6471;
  assign n6473 = ~n6470 & n6472;
  assign n6474 = pi11  & n6473;
  assign n6475 = ~pi11  & ~n6473;
  assign n6476 = ~n6474 & ~n6475;
  assign n6477 = ~n6414 & ~n6416;
  assign n6478 = ~n6408 & ~n6410;
  assign n6479 = pi92  & n1296;
  assign n6480 = pi93  & n1207;
  assign n6481 = pi94  & n1202;
  assign n6482 = n1200 & n3280;
  assign n6483 = ~n6480 & ~n6481;
  assign n6484 = ~n6479 & n6483;
  assign n6485 = ~n6482 & n6484;
  assign n6486 = pi17  & n6485;
  assign n6487 = ~pi17  & ~n6485;
  assign n6488 = ~n6486 & ~n6487;
  assign n6489 = ~n6402 & ~n6404;
  assign n6490 = ~n6395 & ~n6398;
  assign n6491 = ~n6379 & ~n6383;
  assign n6492 = ~n6364 & ~n6366;
  assign n6493 = pi80  & n3011;
  assign n6494 = pi81  & n2809;
  assign n6495 = pi82  & n2804;
  assign n6496 = n1450 & n2802;
  assign n6497 = ~n6494 & ~n6495;
  assign n6498 = ~n6493 & n6497;
  assign n6499 = ~n6496 & n6498;
  assign n6500 = pi29  & n6499;
  assign n6501 = ~pi29  & ~n6499;
  assign n6502 = ~n6500 & ~n6501;
  assign n6503 = ~n6358 & ~n6360;
  assign n6504 = pi77  & n3553;
  assign n6505 = pi78  & n3334;
  assign n6506 = pi79  & n3329;
  assign n6507 = n1048 & n3327;
  assign n6508 = ~n6505 & ~n6506;
  assign n6509 = ~n6504 & n6508;
  assign n6510 = ~n6507 & n6509;
  assign n6511 = pi32  & n6510;
  assign n6512 = ~pi32  & ~n6510;
  assign n6513 = ~n6511 & ~n6512;
  assign n6514 = ~n6352 & ~n6354;
  assign n6515 = pi74  & n4176;
  assign n6516 = pi75  & n3938;
  assign n6517 = pi76  & n3933;
  assign n6518 = n841 & n3931;
  assign n6519 = ~n6516 & ~n6517;
  assign n6520 = ~n6515 & n6519;
  assign n6521 = ~n6518 & n6520;
  assign n6522 = pi35  & n6521;
  assign n6523 = ~pi35  & ~n6521;
  assign n6524 = ~n6522 & ~n6523;
  assign n6525 = ~n6345 & ~n6348;
  assign n6526 = ~n6339 & ~n6342;
  assign n6527 = pi65  & n6331;
  assign n6528 = pi66  & n6015;
  assign n6529 = pi67  & n6010;
  assign n6530 = n305 & n6008;
  assign n6531 = ~n6528 & ~n6529;
  assign n6532 = ~n6527 & n6531;
  assign n6533 = ~n6530 & n6532;
  assign n6534 = pi44  & n6533;
  assign n6535 = ~pi44  & ~n6533;
  assign n6536 = ~n6534 & ~n6535;
  assign n6537 = ~pi44  & ~pi45 ;
  assign n6538 = pi44  & pi45 ;
  assign n6539 = ~n6537 & ~n6538;
  assign n6540 = pi64  & n6539;
  assign n6541 = n6325 & n6335;
  assign n6542 = n6540 & n6541;
  assign n6543 = ~n6540 & ~n6541;
  assign n6544 = ~n6542 & ~n6543;
  assign n6545 = ~n6536 & n6544;
  assign n6546 = n6536 & ~n6544;
  assign n6547 = ~n6545 & ~n6546;
  assign n6548 = pi68  & n5558;
  assign n6549 = pi69  & n5293;
  assign n6550 = pi70  & n5288;
  assign n6551 = n415 & n5286;
  assign n6552 = ~n6549 & ~n6550;
  assign n6553 = ~n6548 & n6552;
  assign n6554 = ~n6551 & n6553;
  assign n6555 = pi41  & n6554;
  assign n6556 = ~pi41  & ~n6554;
  assign n6557 = ~n6555 & ~n6556;
  assign n6558 = n6547 & ~n6557;
  assign n6559 = ~n6547 & n6557;
  assign n6560 = ~n6558 & ~n6559;
  assign n6561 = n6526 & ~n6560;
  assign n6562 = ~n6526 & n6560;
  assign n6563 = ~n6561 & ~n6562;
  assign n6564 = pi71  & n4843;
  assign n6565 = pi72  & n4598;
  assign n6566 = pi73  & n4593;
  assign n6567 = n613 & n4591;
  assign n6568 = ~n6565 & ~n6566;
  assign n6569 = ~n6564 & n6568;
  assign n6570 = ~n6567 & n6569;
  assign n6571 = pi38  & n6570;
  assign n6572 = ~pi38  & ~n6570;
  assign n6573 = ~n6571 & ~n6572;
  assign n6574 = ~n6563 & n6573;
  assign n6575 = n6563 & ~n6573;
  assign n6576 = ~n6574 & ~n6575;
  assign n6577 = ~n6525 & n6576;
  assign n6578 = n6525 & ~n6576;
  assign n6579 = ~n6577 & ~n6578;
  assign n6580 = ~n6524 & n6579;
  assign n6581 = n6524 & ~n6579;
  assign n6582 = ~n6580 & ~n6581;
  assign n6583 = ~n6514 & n6582;
  assign n6584 = n6514 & ~n6582;
  assign n6585 = ~n6583 & ~n6584;
  assign n6586 = ~n6513 & n6585;
  assign n6587 = n6513 & ~n6585;
  assign n6588 = ~n6586 & ~n6587;
  assign n6589 = ~n6503 & n6588;
  assign n6590 = n6503 & ~n6588;
  assign n6591 = ~n6589 & ~n6590;
  assign n6592 = ~n6502 & n6591;
  assign n6593 = n6502 & ~n6591;
  assign n6594 = ~n6592 & ~n6593;
  assign n6595 = ~n6492 & n6594;
  assign n6596 = n6492 & ~n6594;
  assign n6597 = ~n6595 & ~n6596;
  assign n6598 = pi83  & n2510;
  assign n6599 = pi84  & n2342;
  assign n6600 = pi85  & n2337;
  assign n6601 = n1831 & n2335;
  assign n6602 = ~n6599 & ~n6600;
  assign n6603 = ~n6598 & n6602;
  assign n6604 = ~n6601 & n6603;
  assign n6605 = pi26  & n6604;
  assign n6606 = ~pi26  & ~n6604;
  assign n6607 = ~n6605 & ~n6606;
  assign n6608 = n6597 & ~n6607;
  assign n6609 = ~n6597 & n6607;
  assign n6610 = ~n6608 & ~n6609;
  assign n6611 = n6491 & ~n6610;
  assign n6612 = ~n6491 & n6610;
  assign n6613 = ~n6611 & ~n6612;
  assign n6614 = pi86  & n2053;
  assign n6615 = pi87  & n1893;
  assign n6616 = pi88  & n1888;
  assign n6617 = n1886 & n2140;
  assign n6618 = ~n6615 & ~n6616;
  assign n6619 = ~n6614 & n6618;
  assign n6620 = ~n6617 & n6619;
  assign n6621 = pi23  & n6620;
  assign n6622 = ~pi23  & ~n6620;
  assign n6623 = ~n6621 & ~n6622;
  assign n6624 = ~n6613 & n6623;
  assign n6625 = n6613 & ~n6623;
  assign n6626 = ~n6624 & ~n6625;
  assign n6627 = ~n6490 & n6626;
  assign n6628 = n6490 & ~n6626;
  assign n6629 = ~n6627 & ~n6628;
  assign n6630 = pi89  & n1661;
  assign n6631 = pi90  & n1500;
  assign n6632 = pi91  & n1495;
  assign n6633 = n1493 & n2746;
  assign n6634 = ~n6631 & ~n6632;
  assign n6635 = ~n6630 & n6634;
  assign n6636 = ~n6633 & n6635;
  assign n6637 = pi20  & n6636;
  assign n6638 = ~pi20  & ~n6636;
  assign n6639 = ~n6637 & ~n6638;
  assign n6640 = n6629 & ~n6639;
  assign n6641 = ~n6629 & n6639;
  assign n6642 = ~n6640 & ~n6641;
  assign n6643 = ~n6489 & n6642;
  assign n6644 = n6489 & ~n6642;
  assign n6645 = ~n6643 & ~n6644;
  assign n6646 = ~n6488 & n6645;
  assign n6647 = n6488 & ~n6645;
  assign n6648 = ~n6646 & ~n6647;
  assign n6649 = ~n6478 & n6648;
  assign n6650 = n6478 & ~n6648;
  assign n6651 = ~n6649 & ~n6650;
  assign n6652 = pi95  & n1006;
  assign n6653 = pi96  & n897;
  assign n6654 = pi97  & n892;
  assign n6655 = n890 & n3691;
  assign n6656 = ~n6653 & ~n6654;
  assign n6657 = ~n6652 & n6656;
  assign n6658 = ~n6655 & n6657;
  assign n6659 = pi14  & n6658;
  assign n6660 = ~pi14  & ~n6658;
  assign n6661 = ~n6659 & ~n6660;
  assign n6662 = n6651 & ~n6661;
  assign n6663 = ~n6651 & n6661;
  assign n6664 = ~n6662 & ~n6663;
  assign n6665 = ~n6477 & n6664;
  assign n6666 = n6477 & ~n6664;
  assign n6667 = ~n6665 & ~n6666;
  assign n6668 = ~n6476 & n6667;
  assign n6669 = n6476 & ~n6667;
  assign n6670 = ~n6668 & ~n6669;
  assign n6671 = n6466 & ~n6670;
  assign n6672 = ~n6466 & n6670;
  assign n6673 = ~n6671 & ~n6672;
  assign n6674 = pi101  & n528;
  assign n6675 = pi102  & n490;
  assign n6676 = pi103  & n485;
  assign n6677 = n483 & n5188;
  assign n6678 = ~n6675 & ~n6676;
  assign n6679 = ~n6674 & n6678;
  assign n6680 = ~n6677 & n6679;
  assign n6681 = pi8  & n6680;
  assign n6682 = ~pi8  & ~n6680;
  assign n6683 = ~n6681 & ~n6682;
  assign n6684 = n6673 & ~n6683;
  assign n6685 = ~n6673 & n6683;
  assign n6686 = ~n6684 & ~n6685;
  assign n6687 = n6465 & ~n6686;
  assign n6688 = ~n6465 & n6686;
  assign n6689 = ~n6687 & ~n6688;
  assign n6690 = pi104  & n391;
  assign n6691 = pi105  & n353;
  assign n6692 = pi106  & n348;
  assign n6693 = n346 & n5701;
  assign n6694 = ~n6691 & ~n6692;
  assign n6695 = ~n6690 & n6694;
  assign n6696 = ~n6693 & n6695;
  assign n6697 = pi5  & n6696;
  assign n6698 = ~pi5  & ~n6696;
  assign n6699 = ~n6697 & ~n6698;
  assign n6700 = n6689 & ~n6699;
  assign n6701 = ~n6689 & n6699;
  assign n6702 = ~n6700 & ~n6701;
  assign n6703 = n6464 & ~n6702;
  assign n6704 = ~n6464 & n6702;
  assign n6705 = ~n6703 & ~n6704;
  assign n6706 = pi109  & n269;
  assign n6707 = pi108  & n267;
  assign n6708 = pi107  & n282;
  assign n6709 = ~n6209 & ~n6211;
  assign n6710 = ~pi108  & ~pi109 ;
  assign n6711 = pi108  & pi109 ;
  assign n6712 = ~n6710 & ~n6711;
  assign n6713 = ~n6709 & n6712;
  assign n6714 = n6709 & ~n6712;
  assign n6715 = ~n6713 & ~n6714;
  assign n6716 = n262 & n6715;
  assign n6717 = ~n6706 & ~n6707;
  assign n6718 = ~n6708 & n6717;
  assign n6719 = ~n6716 & n6718;
  assign n6720 = pi2  & n6719;
  assign n6721 = ~pi2  & ~n6719;
  assign n6722 = ~n6720 & ~n6721;
  assign n6723 = ~n6705 & n6722;
  assign n6724 = n6705 & ~n6722;
  assign n6725 = ~n6723 & ~n6724;
  assign n6726 = ~n6463 & n6725;
  assign n6727 = n6463 & ~n6725;
  assign po45  = ~n6726 & ~n6727;
  assign n6729 = ~n6724 & ~n6726;
  assign n6730 = ~n6700 & ~n6704;
  assign n6731 = ~n6684 & ~n6688;
  assign n6732 = ~n6668 & ~n6672;
  assign n6733 = ~n6662 & ~n6665;
  assign n6734 = ~n6646 & ~n6649;
  assign n6735 = pi93  & n1296;
  assign n6736 = pi94  & n1207;
  assign n6737 = pi95  & n1202;
  assign n6738 = n1200 & n3475;
  assign n6739 = ~n6736 & ~n6737;
  assign n6740 = ~n6735 & n6739;
  assign n6741 = ~n6738 & n6740;
  assign n6742 = pi17  & n6741;
  assign n6743 = ~pi17  & ~n6741;
  assign n6744 = ~n6742 & ~n6743;
  assign n6745 = ~n6640 & ~n6643;
  assign n6746 = pi90  & n1661;
  assign n6747 = pi91  & n1500;
  assign n6748 = pi92  & n1495;
  assign n6749 = n1493 & n2924;
  assign n6750 = ~n6747 & ~n6748;
  assign n6751 = ~n6746 & n6750;
  assign n6752 = ~n6749 & n6751;
  assign n6753 = pi20  & n6752;
  assign n6754 = ~pi20  & ~n6752;
  assign n6755 = ~n6753 & ~n6754;
  assign n6756 = ~n6625 & ~n6627;
  assign n6757 = ~n6608 & ~n6612;
  assign n6758 = ~n6592 & ~n6595;
  assign n6759 = ~n6586 & ~n6589;
  assign n6760 = ~n6580 & ~n6583;
  assign n6761 = pi75  & n4176;
  assign n6762 = pi76  & n3938;
  assign n6763 = pi77  & n3933;
  assign n6764 = n865 & n3931;
  assign n6765 = ~n6762 & ~n6763;
  assign n6766 = ~n6761 & n6765;
  assign n6767 = ~n6764 & n6766;
  assign n6768 = pi35  & n6767;
  assign n6769 = ~pi35  & ~n6767;
  assign n6770 = ~n6768 & ~n6769;
  assign n6771 = ~n6575 & ~n6577;
  assign n6772 = ~n6558 & ~n6562;
  assign n6773 = ~n6542 & ~n6545;
  assign n6774 = pi66  & n6331;
  assign n6775 = pi67  & n6015;
  assign n6776 = pi68  & n6010;
  assign n6777 = n334 & n6008;
  assign n6778 = ~n6775 & ~n6776;
  assign n6779 = ~n6774 & n6778;
  assign n6780 = ~n6777 & n6779;
  assign n6781 = pi44  & n6780;
  assign n6782 = ~pi44  & ~n6780;
  assign n6783 = ~n6781 & ~n6782;
  assign n6784 = pi47  & n6540;
  assign n6785 = ~pi46  & ~pi47 ;
  assign n6786 = pi46  & pi47 ;
  assign n6787 = ~n6785 & ~n6786;
  assign n6788 = n6539 & n6787;
  assign n6789 = n265 & n6788;
  assign n6790 = n6539 & ~n6787;
  assign n6791 = pi65  & n6790;
  assign n6792 = ~pi45  & ~pi46 ;
  assign n6793 = pi45  & pi46 ;
  assign n6794 = ~n6792 & ~n6793;
  assign n6795 = ~n6539 & n6794;
  assign n6796 = pi64  & n6795;
  assign n6797 = ~n6789 & ~n6791;
  assign n6798 = ~n6796 & n6797;
  assign n6799 = n6784 & ~n6798;
  assign n6800 = ~n6784 & n6798;
  assign n6801 = ~n6799 & ~n6800;
  assign n6802 = n6783 & ~n6801;
  assign n6803 = ~n6783 & n6801;
  assign n6804 = ~n6802 & ~n6803;
  assign n6805 = ~n6773 & n6804;
  assign n6806 = n6773 & ~n6804;
  assign n6807 = ~n6805 & ~n6806;
  assign n6808 = pi69  & n5558;
  assign n6809 = pi70  & n5293;
  assign n6810 = pi71  & n5288;
  assign n6811 = n460 & n5286;
  assign n6812 = ~n6809 & ~n6810;
  assign n6813 = ~n6808 & n6812;
  assign n6814 = ~n6811 & n6813;
  assign n6815 = pi41  & n6814;
  assign n6816 = ~pi41  & ~n6814;
  assign n6817 = ~n6815 & ~n6816;
  assign n6818 = n6807 & ~n6817;
  assign n6819 = ~n6807 & n6817;
  assign n6820 = ~n6818 & ~n6819;
  assign n6821 = n6772 & ~n6820;
  assign n6822 = ~n6772 & n6820;
  assign n6823 = ~n6821 & ~n6822;
  assign n6824 = pi72  & n4843;
  assign n6825 = pi73  & n4598;
  assign n6826 = pi74  & n4593;
  assign n6827 = n689 & n4591;
  assign n6828 = ~n6825 & ~n6826;
  assign n6829 = ~n6824 & n6828;
  assign n6830 = ~n6827 & n6829;
  assign n6831 = pi38  & n6830;
  assign n6832 = ~pi38  & ~n6830;
  assign n6833 = ~n6831 & ~n6832;
  assign n6834 = n6823 & ~n6833;
  assign n6835 = ~n6823 & n6833;
  assign n6836 = ~n6834 & ~n6835;
  assign n6837 = ~n6771 & n6836;
  assign n6838 = n6771 & ~n6836;
  assign n6839 = ~n6837 & ~n6838;
  assign n6840 = n6770 & ~n6839;
  assign n6841 = ~n6770 & n6839;
  assign n6842 = ~n6840 & ~n6841;
  assign n6843 = ~n6760 & n6842;
  assign n6844 = n6760 & ~n6842;
  assign n6845 = ~n6843 & ~n6844;
  assign n6846 = pi78  & n3553;
  assign n6847 = pi79  & n3334;
  assign n6848 = pi80  & n3329;
  assign n6849 = n1144 & n3327;
  assign n6850 = ~n6847 & ~n6848;
  assign n6851 = ~n6846 & n6850;
  assign n6852 = ~n6849 & n6851;
  assign n6853 = pi32  & n6852;
  assign n6854 = ~pi32  & ~n6852;
  assign n6855 = ~n6853 & ~n6854;
  assign n6856 = n6845 & ~n6855;
  assign n6857 = ~n6845 & n6855;
  assign n6858 = ~n6856 & ~n6857;
  assign n6859 = n6759 & ~n6858;
  assign n6860 = ~n6759 & n6858;
  assign n6861 = ~n6859 & ~n6860;
  assign n6862 = pi81  & n3011;
  assign n6863 = pi82  & n2809;
  assign n6864 = pi83  & n2804;
  assign n6865 = n1577 & n2802;
  assign n6866 = ~n6863 & ~n6864;
  assign n6867 = ~n6862 & n6866;
  assign n6868 = ~n6865 & n6867;
  assign n6869 = pi29  & n6868;
  assign n6870 = ~pi29  & ~n6868;
  assign n6871 = ~n6869 & ~n6870;
  assign n6872 = n6861 & ~n6871;
  assign n6873 = ~n6861 & n6871;
  assign n6874 = ~n6872 & ~n6873;
  assign n6875 = n6758 & ~n6874;
  assign n6876 = ~n6758 & n6874;
  assign n6877 = ~n6875 & ~n6876;
  assign n6878 = pi84  & n2510;
  assign n6879 = pi85  & n2342;
  assign n6880 = pi86  & n2337;
  assign n6881 = n1975 & n2335;
  assign n6882 = ~n6879 & ~n6880;
  assign n6883 = ~n6878 & n6882;
  assign n6884 = ~n6881 & n6883;
  assign n6885 = pi26  & n6884;
  assign n6886 = ~pi26  & ~n6884;
  assign n6887 = ~n6885 & ~n6886;
  assign n6888 = n6877 & ~n6887;
  assign n6889 = ~n6877 & n6887;
  assign n6890 = ~n6888 & ~n6889;
  assign n6891 = n6757 & ~n6890;
  assign n6892 = ~n6757 & n6890;
  assign n6893 = ~n6891 & ~n6892;
  assign n6894 = pi87  & n2053;
  assign n6895 = pi88  & n1893;
  assign n6896 = pi89  & n1888;
  assign n6897 = n1886 & n2287;
  assign n6898 = ~n6895 & ~n6896;
  assign n6899 = ~n6894 & n6898;
  assign n6900 = ~n6897 & n6899;
  assign n6901 = pi23  & n6900;
  assign n6902 = ~pi23  & ~n6900;
  assign n6903 = ~n6901 & ~n6902;
  assign n6904 = n6893 & ~n6903;
  assign n6905 = ~n6893 & n6903;
  assign n6906 = ~n6904 & ~n6905;
  assign n6907 = ~n6756 & n6906;
  assign n6908 = n6756 & ~n6906;
  assign n6909 = ~n6907 & ~n6908;
  assign n6910 = ~n6755 & n6909;
  assign n6911 = n6755 & ~n6909;
  assign n6912 = ~n6910 & ~n6911;
  assign n6913 = ~n6745 & n6912;
  assign n6914 = n6745 & ~n6912;
  assign n6915 = ~n6913 & ~n6914;
  assign n6916 = n6744 & ~n6915;
  assign n6917 = ~n6744 & n6915;
  assign n6918 = ~n6916 & ~n6917;
  assign n6919 = ~n6734 & n6918;
  assign n6920 = n6734 & ~n6918;
  assign n6921 = ~n6919 & ~n6920;
  assign n6922 = pi96  & n1006;
  assign n6923 = pi97  & n897;
  assign n6924 = pi98  & n892;
  assign n6925 = n890 & n3889;
  assign n6926 = ~n6923 & ~n6924;
  assign n6927 = ~n6922 & n6926;
  assign n6928 = ~n6925 & n6927;
  assign n6929 = pi14  & n6928;
  assign n6930 = ~pi14  & ~n6928;
  assign n6931 = ~n6929 & ~n6930;
  assign n6932 = n6921 & ~n6931;
  assign n6933 = ~n6921 & n6931;
  assign n6934 = ~n6932 & ~n6933;
  assign n6935 = n6733 & ~n6934;
  assign n6936 = ~n6733 & n6934;
  assign n6937 = ~n6935 & ~n6936;
  assign n6938 = pi99  & n750;
  assign n6939 = pi100  & n651;
  assign n6940 = pi101  & n646;
  assign n6941 = n644 & n4730;
  assign n6942 = ~n6939 & ~n6940;
  assign n6943 = ~n6938 & n6942;
  assign n6944 = ~n6941 & n6943;
  assign n6945 = pi11  & n6944;
  assign n6946 = ~pi11  & ~n6944;
  assign n6947 = ~n6945 & ~n6946;
  assign n6948 = n6937 & ~n6947;
  assign n6949 = ~n6937 & n6947;
  assign n6950 = ~n6948 & ~n6949;
  assign n6951 = n6732 & ~n6950;
  assign n6952 = ~n6732 & n6950;
  assign n6953 = ~n6951 & ~n6952;
  assign n6954 = pi102  & n528;
  assign n6955 = pi103  & n490;
  assign n6956 = pi104  & n485;
  assign n6957 = n483 & n5212;
  assign n6958 = ~n6955 & ~n6956;
  assign n6959 = ~n6954 & n6958;
  assign n6960 = ~n6957 & n6959;
  assign n6961 = pi8  & n6960;
  assign n6962 = ~pi8  & ~n6960;
  assign n6963 = ~n6961 & ~n6962;
  assign n6964 = n6953 & ~n6963;
  assign n6965 = ~n6953 & n6963;
  assign n6966 = ~n6964 & ~n6965;
  assign n6967 = ~n6731 & n6966;
  assign n6968 = n6731 & ~n6966;
  assign n6969 = ~n6967 & ~n6968;
  assign n6970 = pi105  & n391;
  assign n6971 = pi106  & n353;
  assign n6972 = pi107  & n348;
  assign n6973 = n346 & n6189;
  assign n6974 = ~n6971 & ~n6972;
  assign n6975 = ~n6970 & n6974;
  assign n6976 = ~n6973 & n6975;
  assign n6977 = pi5  & n6976;
  assign n6978 = ~pi5  & ~n6976;
  assign n6979 = ~n6977 & ~n6978;
  assign n6980 = n6969 & ~n6979;
  assign n6981 = ~n6969 & n6979;
  assign n6982 = ~n6980 & ~n6981;
  assign n6983 = n6730 & ~n6982;
  assign n6984 = ~n6730 & n6982;
  assign n6985 = ~n6983 & ~n6984;
  assign n6986 = pi110  & n269;
  assign n6987 = pi109  & n267;
  assign n6988 = pi108  & n282;
  assign n6989 = ~n6711 & ~n6713;
  assign n6990 = ~pi109  & ~pi110 ;
  assign n6991 = pi109  & pi110 ;
  assign n6992 = ~n6990 & ~n6991;
  assign n6993 = ~n6989 & n6992;
  assign n6994 = n6989 & ~n6992;
  assign n6995 = ~n6993 & ~n6994;
  assign n6996 = n262 & n6995;
  assign n6997 = ~n6986 & ~n6987;
  assign n6998 = ~n6988 & n6997;
  assign n6999 = ~n6996 & n6998;
  assign n7000 = pi2  & n6999;
  assign n7001 = ~pi2  & ~n6999;
  assign n7002 = ~n7000 & ~n7001;
  assign n7003 = n6985 & ~n7002;
  assign n7004 = ~n6985 & n7002;
  assign n7005 = ~n7003 & ~n7004;
  assign n7006 = ~n6729 & n7005;
  assign n7007 = n6729 & ~n7005;
  assign po46  = ~n7006 & ~n7007;
  assign n7009 = ~n7003 & ~n7006;
  assign n7010 = ~n6980 & ~n6984;
  assign n7011 = pi106  & n391;
  assign n7012 = pi107  & n353;
  assign n7013 = pi108  & n348;
  assign n7014 = n346 & n6213;
  assign n7015 = ~n7012 & ~n7013;
  assign n7016 = ~n7011 & n7015;
  assign n7017 = ~n7014 & n7016;
  assign n7018 = pi5  & n7017;
  assign n7019 = ~pi5  & ~n7017;
  assign n7020 = ~n7018 & ~n7019;
  assign n7021 = ~n6964 & ~n6967;
  assign n7022 = ~n6948 & ~n6952;
  assign n7023 = ~n6932 & ~n6936;
  assign n7024 = ~n6917 & ~n6919;
  assign n7025 = pi94  & n1296;
  assign n7026 = pi95  & n1207;
  assign n7027 = pi96  & n1202;
  assign n7028 = n1200 & n3499;
  assign n7029 = ~n7026 & ~n7027;
  assign n7030 = ~n7025 & n7029;
  assign n7031 = ~n7028 & n7030;
  assign n7032 = pi17  & n7031;
  assign n7033 = ~pi17  & ~n7031;
  assign n7034 = ~n7032 & ~n7033;
  assign n7035 = ~n6910 & ~n6913;
  assign n7036 = pi91  & n1661;
  assign n7037 = pi92  & n1500;
  assign n7038 = pi93  & n1495;
  assign n7039 = n1493 & n2948;
  assign n7040 = ~n7037 & ~n7038;
  assign n7041 = ~n7036 & n7040;
  assign n7042 = ~n7039 & n7041;
  assign n7043 = pi20  & n7042;
  assign n7044 = ~pi20  & ~n7042;
  assign n7045 = ~n7043 & ~n7044;
  assign n7046 = ~n6904 & ~n6907;
  assign n7047 = pi88  & n2053;
  assign n7048 = pi89  & n1893;
  assign n7049 = pi90  & n1888;
  assign n7050 = n1886 & n2448;
  assign n7051 = ~n7048 & ~n7049;
  assign n7052 = ~n7047 & n7051;
  assign n7053 = ~n7050 & n7052;
  assign n7054 = pi23  & n7053;
  assign n7055 = ~pi23  & ~n7053;
  assign n7056 = ~n7054 & ~n7055;
  assign n7057 = ~n6888 & ~n6892;
  assign n7058 = ~n6872 & ~n6876;
  assign n7059 = pi82  & n3011;
  assign n7060 = pi83  & n2809;
  assign n7061 = pi84  & n2804;
  assign n7062 = n1601 & n2802;
  assign n7063 = ~n7060 & ~n7061;
  assign n7064 = ~n7059 & n7063;
  assign n7065 = ~n7062 & n7064;
  assign n7066 = pi29  & n7065;
  assign n7067 = ~pi29  & ~n7065;
  assign n7068 = ~n7066 & ~n7067;
  assign n7069 = ~n6856 & ~n6860;
  assign n7070 = pi79  & n3553;
  assign n7071 = pi80  & n3334;
  assign n7072 = pi81  & n3329;
  assign n7073 = n1337 & n3327;
  assign n7074 = ~n7071 & ~n7072;
  assign n7075 = ~n7070 & n7074;
  assign n7076 = ~n7073 & n7075;
  assign n7077 = pi32  & n7076;
  assign n7078 = ~pi32  & ~n7076;
  assign n7079 = ~n7077 & ~n7078;
  assign n7080 = ~n6841 & ~n6843;
  assign n7081 = ~n6834 & ~n6837;
  assign n7082 = pi73  & n4843;
  assign n7083 = pi74  & n4598;
  assign n7084 = pi75  & n4593;
  assign n7085 = n713 & n4591;
  assign n7086 = ~n7083 & ~n7084;
  assign n7087 = ~n7082 & n7086;
  assign n7088 = ~n7085 & n7087;
  assign n7089 = pi38  & n7088;
  assign n7090 = ~pi38  & ~n7088;
  assign n7091 = ~n7089 & ~n7090;
  assign n7092 = ~n6818 & ~n6822;
  assign n7093 = pi70  & n5558;
  assign n7094 = pi71  & n5293;
  assign n7095 = pi72  & n5288;
  assign n7096 = n551 & n5286;
  assign n7097 = ~n7094 & ~n7095;
  assign n7098 = ~n7093 & n7097;
  assign n7099 = ~n7096 & n7098;
  assign n7100 = pi41  & n7099;
  assign n7101 = ~pi41  & ~n7099;
  assign n7102 = ~n7100 & ~n7101;
  assign n7103 = ~n6803 & ~n6805;
  assign n7104 = pi67  & n6331;
  assign n7105 = pi68  & n6015;
  assign n7106 = pi69  & n6010;
  assign n7107 = n376 & n6008;
  assign n7108 = ~n7105 & ~n7106;
  assign n7109 = ~n7104 & n7108;
  assign n7110 = ~n7107 & n7109;
  assign n7111 = pi44  & n7110;
  assign n7112 = ~pi44  & ~n7110;
  assign n7113 = ~n7111 & ~n7112;
  assign n7114 = pi47  & ~n6540;
  assign n7115 = n6798 & n7114;
  assign n7116 = pi47  & ~n7115;
  assign n7117 = ~n287 & n6788;
  assign n7118 = pi65  & n6795;
  assign n7119 = pi66  & n6790;
  assign n7120 = ~n6539 & n6787;
  assign n7121 = ~n6794 & n7120;
  assign n7122 = pi64  & n7121;
  assign n7123 = ~n7117 & ~n7118;
  assign n7124 = ~n7119 & n7123;
  assign n7125 = ~n7122 & n7124;
  assign n7126 = ~n7116 & n7125;
  assign n7127 = n7116 & ~n7125;
  assign n7128 = ~n7126 & ~n7127;
  assign n7129 = ~n7113 & n7128;
  assign n7130 = n7113 & ~n7128;
  assign n7131 = ~n7129 & ~n7130;
  assign n7132 = ~n7103 & n7131;
  assign n7133 = n7103 & ~n7131;
  assign n7134 = ~n7132 & ~n7133;
  assign n7135 = ~n7102 & n7134;
  assign n7136 = n7102 & ~n7134;
  assign n7137 = ~n7135 & ~n7136;
  assign n7138 = ~n7092 & n7137;
  assign n7139 = n7092 & ~n7137;
  assign n7140 = ~n7138 & ~n7139;
  assign n7141 = n7091 & ~n7140;
  assign n7142 = ~n7091 & n7140;
  assign n7143 = ~n7141 & ~n7142;
  assign n7144 = ~n7081 & n7143;
  assign n7145 = n7081 & ~n7143;
  assign n7146 = ~n7144 & ~n7145;
  assign n7147 = pi76  & n4176;
  assign n7148 = pi77  & n3938;
  assign n7149 = pi78  & n3933;
  assign n7150 = n958 & n3931;
  assign n7151 = ~n7148 & ~n7149;
  assign n7152 = ~n7147 & n7151;
  assign n7153 = ~n7150 & n7152;
  assign n7154 = pi35  & n7153;
  assign n7155 = ~pi35  & ~n7153;
  assign n7156 = ~n7154 & ~n7155;
  assign n7157 = n7146 & ~n7156;
  assign n7158 = ~n7146 & n7156;
  assign n7159 = ~n7157 & ~n7158;
  assign n7160 = ~n7080 & n7159;
  assign n7161 = n7080 & ~n7159;
  assign n7162 = ~n7160 & ~n7161;
  assign n7163 = ~n7079 & n7162;
  assign n7164 = n7079 & ~n7162;
  assign n7165 = ~n7163 & ~n7164;
  assign n7166 = ~n7069 & n7165;
  assign n7167 = n7069 & ~n7165;
  assign n7168 = ~n7166 & ~n7167;
  assign n7169 = ~n7068 & n7168;
  assign n7170 = n7068 & ~n7168;
  assign n7171 = ~n7169 & ~n7170;
  assign n7172 = n7058 & ~n7171;
  assign n7173 = ~n7058 & n7171;
  assign n7174 = ~n7172 & ~n7173;
  assign n7175 = pi85  & n2510;
  assign n7176 = pi86  & n2342;
  assign n7177 = pi87  & n2337;
  assign n7178 = n2116 & n2335;
  assign n7179 = ~n7176 & ~n7177;
  assign n7180 = ~n7175 & n7179;
  assign n7181 = ~n7178 & n7180;
  assign n7182 = pi26  & n7181;
  assign n7183 = ~pi26  & ~n7181;
  assign n7184 = ~n7182 & ~n7183;
  assign n7185 = n7174 & ~n7184;
  assign n7186 = ~n7174 & n7184;
  assign n7187 = ~n7185 & ~n7186;
  assign n7188 = ~n7057 & n7187;
  assign n7189 = n7057 & ~n7187;
  assign n7190 = ~n7188 & ~n7189;
  assign n7191 = n7056 & ~n7190;
  assign n7192 = ~n7056 & n7190;
  assign n7193 = ~n7191 & ~n7192;
  assign n7194 = ~n7046 & n7193;
  assign n7195 = n7046 & ~n7193;
  assign n7196 = ~n7194 & ~n7195;
  assign n7197 = n7045 & ~n7196;
  assign n7198 = ~n7045 & n7196;
  assign n7199 = ~n7197 & ~n7198;
  assign n7200 = ~n7035 & n7199;
  assign n7201 = n7035 & ~n7199;
  assign n7202 = ~n7200 & ~n7201;
  assign n7203 = n7034 & ~n7202;
  assign n7204 = ~n7034 & n7202;
  assign n7205 = ~n7203 & ~n7204;
  assign n7206 = ~n7024 & n7205;
  assign n7207 = n7024 & ~n7205;
  assign n7208 = ~n7206 & ~n7207;
  assign n7209 = pi97  & n1006;
  assign n7210 = pi98  & n897;
  assign n7211 = pi99  & n892;
  assign n7212 = n890 & n4101;
  assign n7213 = ~n7210 & ~n7211;
  assign n7214 = ~n7209 & n7213;
  assign n7215 = ~n7212 & n7214;
  assign n7216 = pi14  & n7215;
  assign n7217 = ~pi14  & ~n7215;
  assign n7218 = ~n7216 & ~n7217;
  assign n7219 = n7208 & ~n7218;
  assign n7220 = ~n7208 & n7218;
  assign n7221 = ~n7219 & ~n7220;
  assign n7222 = n7023 & ~n7221;
  assign n7223 = ~n7023 & n7221;
  assign n7224 = ~n7222 & ~n7223;
  assign n7225 = pi100  & n750;
  assign n7226 = pi101  & n651;
  assign n7227 = pi102  & n646;
  assign n7228 = n644 & n4956;
  assign n7229 = ~n7226 & ~n7227;
  assign n7230 = ~n7225 & n7229;
  assign n7231 = ~n7228 & n7230;
  assign n7232 = pi11  & n7231;
  assign n7233 = ~pi11  & ~n7231;
  assign n7234 = ~n7232 & ~n7233;
  assign n7235 = n7224 & ~n7234;
  assign n7236 = ~n7224 & n7234;
  assign n7237 = ~n7235 & ~n7236;
  assign n7238 = n7022 & ~n7237;
  assign n7239 = ~n7022 & n7237;
  assign n7240 = ~n7238 & ~n7239;
  assign n7241 = pi103  & n528;
  assign n7242 = pi104  & n490;
  assign n7243 = pi105  & n485;
  assign n7244 = n483 & n5677;
  assign n7245 = ~n7242 & ~n7243;
  assign n7246 = ~n7241 & n7245;
  assign n7247 = ~n7244 & n7246;
  assign n7248 = pi8  & n7247;
  assign n7249 = ~pi8  & ~n7247;
  assign n7250 = ~n7248 & ~n7249;
  assign n7251 = n7240 & ~n7250;
  assign n7252 = ~n7240 & n7250;
  assign n7253 = ~n7251 & ~n7252;
  assign n7254 = ~n7021 & n7253;
  assign n7255 = n7021 & ~n7253;
  assign n7256 = ~n7254 & ~n7255;
  assign n7257 = n7020 & ~n7256;
  assign n7258 = ~n7020 & n7256;
  assign n7259 = ~n7257 & ~n7258;
  assign n7260 = ~n7010 & n7259;
  assign n7261 = n7010 & ~n7259;
  assign n7262 = ~n7260 & ~n7261;
  assign n7263 = pi111  & n269;
  assign n7264 = pi110  & n267;
  assign n7265 = pi109  & n282;
  assign n7266 = ~n6991 & ~n6993;
  assign n7267 = ~pi110  & ~pi111 ;
  assign n7268 = pi110  & pi111 ;
  assign n7269 = ~n7267 & ~n7268;
  assign n7270 = ~n7266 & n7269;
  assign n7271 = n7266 & ~n7269;
  assign n7272 = ~n7270 & ~n7271;
  assign n7273 = n262 & n7272;
  assign n7274 = ~n7263 & ~n7264;
  assign n7275 = ~n7265 & n7274;
  assign n7276 = ~n7273 & n7275;
  assign n7277 = pi2  & n7276;
  assign n7278 = ~pi2  & ~n7276;
  assign n7279 = ~n7277 & ~n7278;
  assign n7280 = n7262 & ~n7279;
  assign n7281 = ~n7262 & n7279;
  assign n7282 = ~n7280 & ~n7281;
  assign n7283 = ~n7009 & n7282;
  assign n7284 = n7009 & ~n7282;
  assign po47  = ~n7283 & ~n7284;
  assign n7286 = ~n7280 & ~n7283;
  assign n7287 = pi112  & n269;
  assign n7288 = pi111  & n267;
  assign n7289 = pi110  & n282;
  assign n7290 = ~n7268 & ~n7270;
  assign n7291 = ~pi111  & ~pi112 ;
  assign n7292 = pi111  & pi112 ;
  assign n7293 = ~n7291 & ~n7292;
  assign n7294 = ~n7290 & n7293;
  assign n7295 = n7290 & ~n7293;
  assign n7296 = ~n7294 & ~n7295;
  assign n7297 = n262 & n7296;
  assign n7298 = ~n7287 & ~n7288;
  assign n7299 = ~n7289 & n7298;
  assign n7300 = ~n7297 & n7299;
  assign n7301 = pi2  & n7300;
  assign n7302 = ~pi2  & ~n7300;
  assign n7303 = ~n7301 & ~n7302;
  assign n7304 = ~n7258 & ~n7260;
  assign n7305 = pi107  & n391;
  assign n7306 = pi108  & n353;
  assign n7307 = pi109  & n348;
  assign n7308 = n346 & n6715;
  assign n7309 = ~n7306 & ~n7307;
  assign n7310 = ~n7305 & n7309;
  assign n7311 = ~n7308 & n7310;
  assign n7312 = pi5  & n7311;
  assign n7313 = ~pi5  & ~n7311;
  assign n7314 = ~n7312 & ~n7313;
  assign n7315 = ~n7251 & ~n7254;
  assign n7316 = ~n7235 & ~n7239;
  assign n7317 = ~n7219 & ~n7223;
  assign n7318 = pi98  & n1006;
  assign n7319 = pi99  & n897;
  assign n7320 = pi100  & n892;
  assign n7321 = n890 & n4501;
  assign n7322 = ~n7319 & ~n7320;
  assign n7323 = ~n7318 & n7322;
  assign n7324 = ~n7321 & n7323;
  assign n7325 = pi14  & n7324;
  assign n7326 = ~pi14  & ~n7324;
  assign n7327 = ~n7325 & ~n7326;
  assign n7328 = ~n7204 & ~n7206;
  assign n7329 = ~n7198 & ~n7200;
  assign n7330 = pi92  & n1661;
  assign n7331 = pi93  & n1500;
  assign n7332 = pi94  & n1495;
  assign n7333 = n1493 & n3280;
  assign n7334 = ~n7331 & ~n7332;
  assign n7335 = ~n7330 & n7334;
  assign n7336 = ~n7333 & n7335;
  assign n7337 = pi20  & n7336;
  assign n7338 = ~pi20  & ~n7336;
  assign n7339 = ~n7337 & ~n7338;
  assign n7340 = ~n7192 & ~n7194;
  assign n7341 = ~n7185 & ~n7188;
  assign n7342 = ~n7169 & ~n7173;
  assign n7343 = ~n7163 & ~n7166;
  assign n7344 = ~n7157 & ~n7160;
  assign n7345 = pi77  & n4176;
  assign n7346 = pi78  & n3938;
  assign n7347 = pi79  & n3933;
  assign n7348 = n1048 & n3931;
  assign n7349 = ~n7346 & ~n7347;
  assign n7350 = ~n7345 & n7349;
  assign n7351 = ~n7348 & n7350;
  assign n7352 = pi35  & n7351;
  assign n7353 = ~pi35  & ~n7351;
  assign n7354 = ~n7352 & ~n7353;
  assign n7355 = ~n7142 & ~n7144;
  assign n7356 = pi74  & n4843;
  assign n7357 = pi75  & n4598;
  assign n7358 = pi76  & n4593;
  assign n7359 = n841 & n4591;
  assign n7360 = ~n7357 & ~n7358;
  assign n7361 = ~n7356 & n7360;
  assign n7362 = ~n7359 & n7361;
  assign n7363 = pi38  & n7362;
  assign n7364 = ~pi38  & ~n7362;
  assign n7365 = ~n7363 & ~n7364;
  assign n7366 = ~n7135 & ~n7138;
  assign n7367 = ~n7129 & ~n7132;
  assign n7368 = pi65  & n7121;
  assign n7369 = pi66  & n6795;
  assign n7370 = pi67  & n6790;
  assign n7371 = n305 & n6788;
  assign n7372 = ~n7369 & ~n7370;
  assign n7373 = ~n7368 & n7372;
  assign n7374 = ~n7371 & n7373;
  assign n7375 = pi47  & n7374;
  assign n7376 = ~pi47  & ~n7374;
  assign n7377 = ~n7375 & ~n7376;
  assign n7378 = ~pi47  & ~pi48 ;
  assign n7379 = pi47  & pi48 ;
  assign n7380 = ~n7378 & ~n7379;
  assign n7381 = pi64  & n7380;
  assign n7382 = n7115 & n7125;
  assign n7383 = n7381 & n7382;
  assign n7384 = ~n7381 & ~n7382;
  assign n7385 = ~n7383 & ~n7384;
  assign n7386 = ~n7377 & n7385;
  assign n7387 = n7377 & ~n7385;
  assign n7388 = ~n7386 & ~n7387;
  assign n7389 = pi68  & n6331;
  assign n7390 = pi69  & n6015;
  assign n7391 = pi70  & n6010;
  assign n7392 = n415 & n6008;
  assign n7393 = ~n7390 & ~n7391;
  assign n7394 = ~n7389 & n7393;
  assign n7395 = ~n7392 & n7394;
  assign n7396 = pi44  & n7395;
  assign n7397 = ~pi44  & ~n7395;
  assign n7398 = ~n7396 & ~n7397;
  assign n7399 = n7388 & ~n7398;
  assign n7400 = ~n7388 & n7398;
  assign n7401 = ~n7399 & ~n7400;
  assign n7402 = n7367 & ~n7401;
  assign n7403 = ~n7367 & n7401;
  assign n7404 = ~n7402 & ~n7403;
  assign n7405 = pi71  & n5558;
  assign n7406 = pi72  & n5293;
  assign n7407 = pi73  & n5288;
  assign n7408 = n613 & n5286;
  assign n7409 = ~n7406 & ~n7407;
  assign n7410 = ~n7405 & n7409;
  assign n7411 = ~n7408 & n7410;
  assign n7412 = pi41  & n7411;
  assign n7413 = ~pi41  & ~n7411;
  assign n7414 = ~n7412 & ~n7413;
  assign n7415 = ~n7404 & n7414;
  assign n7416 = n7404 & ~n7414;
  assign n7417 = ~n7415 & ~n7416;
  assign n7418 = ~n7366 & n7417;
  assign n7419 = n7366 & ~n7417;
  assign n7420 = ~n7418 & ~n7419;
  assign n7421 = ~n7365 & n7420;
  assign n7422 = n7365 & ~n7420;
  assign n7423 = ~n7421 & ~n7422;
  assign n7424 = ~n7355 & n7423;
  assign n7425 = n7355 & ~n7423;
  assign n7426 = ~n7424 & ~n7425;
  assign n7427 = ~n7354 & n7426;
  assign n7428 = n7354 & ~n7426;
  assign n7429 = ~n7427 & ~n7428;
  assign n7430 = ~n7344 & n7429;
  assign n7431 = n7344 & ~n7429;
  assign n7432 = ~n7430 & ~n7431;
  assign n7433 = pi80  & n3553;
  assign n7434 = pi81  & n3334;
  assign n7435 = pi82  & n3329;
  assign n7436 = n1450 & n3327;
  assign n7437 = ~n7434 & ~n7435;
  assign n7438 = ~n7433 & n7437;
  assign n7439 = ~n7436 & n7438;
  assign n7440 = pi32  & n7439;
  assign n7441 = ~pi32  & ~n7439;
  assign n7442 = ~n7440 & ~n7441;
  assign n7443 = n7432 & ~n7442;
  assign n7444 = ~n7432 & n7442;
  assign n7445 = ~n7443 & ~n7444;
  assign n7446 = n7343 & ~n7445;
  assign n7447 = ~n7343 & n7445;
  assign n7448 = ~n7446 & ~n7447;
  assign n7449 = pi83  & n3011;
  assign n7450 = pi84  & n2809;
  assign n7451 = pi85  & n2804;
  assign n7452 = n1831 & n2802;
  assign n7453 = ~n7450 & ~n7451;
  assign n7454 = ~n7449 & n7453;
  assign n7455 = ~n7452 & n7454;
  assign n7456 = pi29  & n7455;
  assign n7457 = ~pi29  & ~n7455;
  assign n7458 = ~n7456 & ~n7457;
  assign n7459 = n7448 & ~n7458;
  assign n7460 = ~n7448 & n7458;
  assign n7461 = ~n7459 & ~n7460;
  assign n7462 = n7342 & ~n7461;
  assign n7463 = ~n7342 & n7461;
  assign n7464 = ~n7462 & ~n7463;
  assign n7465 = pi86  & n2510;
  assign n7466 = pi87  & n2342;
  assign n7467 = pi88  & n2337;
  assign n7468 = n2140 & n2335;
  assign n7469 = ~n7466 & ~n7467;
  assign n7470 = ~n7465 & n7469;
  assign n7471 = ~n7468 & n7470;
  assign n7472 = pi26  & n7471;
  assign n7473 = ~pi26  & ~n7471;
  assign n7474 = ~n7472 & ~n7473;
  assign n7475 = ~n7464 & n7474;
  assign n7476 = n7464 & ~n7474;
  assign n7477 = ~n7475 & ~n7476;
  assign n7478 = ~n7341 & n7477;
  assign n7479 = n7341 & ~n7477;
  assign n7480 = ~n7478 & ~n7479;
  assign n7481 = pi89  & n2053;
  assign n7482 = pi90  & n1893;
  assign n7483 = pi91  & n1888;
  assign n7484 = n1886 & n2746;
  assign n7485 = ~n7482 & ~n7483;
  assign n7486 = ~n7481 & n7485;
  assign n7487 = ~n7484 & n7486;
  assign n7488 = pi23  & n7487;
  assign n7489 = ~pi23  & ~n7487;
  assign n7490 = ~n7488 & ~n7489;
  assign n7491 = n7480 & ~n7490;
  assign n7492 = ~n7480 & n7490;
  assign n7493 = ~n7491 & ~n7492;
  assign n7494 = ~n7340 & n7493;
  assign n7495 = n7340 & ~n7493;
  assign n7496 = ~n7494 & ~n7495;
  assign n7497 = ~n7339 & n7496;
  assign n7498 = n7339 & ~n7496;
  assign n7499 = ~n7497 & ~n7498;
  assign n7500 = ~n7329 & n7499;
  assign n7501 = n7329 & ~n7499;
  assign n7502 = ~n7500 & ~n7501;
  assign n7503 = pi95  & n1296;
  assign n7504 = pi96  & n1207;
  assign n7505 = pi97  & n1202;
  assign n7506 = n1200 & n3691;
  assign n7507 = ~n7504 & ~n7505;
  assign n7508 = ~n7503 & n7507;
  assign n7509 = ~n7506 & n7508;
  assign n7510 = pi17  & n7509;
  assign n7511 = ~pi17  & ~n7509;
  assign n7512 = ~n7510 & ~n7511;
  assign n7513 = n7502 & ~n7512;
  assign n7514 = ~n7502 & n7512;
  assign n7515 = ~n7513 & ~n7514;
  assign n7516 = ~n7328 & n7515;
  assign n7517 = n7328 & ~n7515;
  assign n7518 = ~n7516 & ~n7517;
  assign n7519 = ~n7327 & n7518;
  assign n7520 = n7327 & ~n7518;
  assign n7521 = ~n7519 & ~n7520;
  assign n7522 = n7317 & ~n7521;
  assign n7523 = ~n7317 & n7521;
  assign n7524 = ~n7522 & ~n7523;
  assign n7525 = pi101  & n750;
  assign n7526 = pi102  & n651;
  assign n7527 = pi103  & n646;
  assign n7528 = n644 & n5188;
  assign n7529 = ~n7526 & ~n7527;
  assign n7530 = ~n7525 & n7529;
  assign n7531 = ~n7528 & n7530;
  assign n7532 = pi11  & n7531;
  assign n7533 = ~pi11  & ~n7531;
  assign n7534 = ~n7532 & ~n7533;
  assign n7535 = n7524 & ~n7534;
  assign n7536 = ~n7524 & n7534;
  assign n7537 = ~n7535 & ~n7536;
  assign n7538 = n7316 & ~n7537;
  assign n7539 = ~n7316 & n7537;
  assign n7540 = ~n7538 & ~n7539;
  assign n7541 = pi104  & n528;
  assign n7542 = pi105  & n490;
  assign n7543 = pi106  & n485;
  assign n7544 = n483 & n5701;
  assign n7545 = ~n7542 & ~n7543;
  assign n7546 = ~n7541 & n7545;
  assign n7547 = ~n7544 & n7546;
  assign n7548 = pi8  & n7547;
  assign n7549 = ~pi8  & ~n7547;
  assign n7550 = ~n7548 & ~n7549;
  assign n7551 = n7540 & ~n7550;
  assign n7552 = ~n7540 & n7550;
  assign n7553 = ~n7551 & ~n7552;
  assign n7554 = ~n7315 & n7553;
  assign n7555 = n7315 & ~n7553;
  assign n7556 = ~n7554 & ~n7555;
  assign n7557 = ~n7314 & n7556;
  assign n7558 = n7314 & ~n7556;
  assign n7559 = ~n7557 & ~n7558;
  assign n7560 = ~n7304 & n7559;
  assign n7561 = n7304 & ~n7559;
  assign n7562 = ~n7560 & ~n7561;
  assign n7563 = n7303 & ~n7562;
  assign n7564 = ~n7303 & n7562;
  assign n7565 = ~n7563 & ~n7564;
  assign n7566 = ~n7286 & n7565;
  assign n7567 = n7286 & ~n7565;
  assign po48  = ~n7566 & ~n7567;
  assign n7569 = ~n7564 & ~n7566;
  assign n7570 = ~n7557 & ~n7560;
  assign n7571 = ~n7551 & ~n7554;
  assign n7572 = ~n7535 & ~n7539;
  assign n7573 = ~n7519 & ~n7523;
  assign n7574 = ~n7513 & ~n7516;
  assign n7575 = ~n7497 & ~n7500;
  assign n7576 = pi93  & n1661;
  assign n7577 = pi94  & n1500;
  assign n7578 = pi95  & n1495;
  assign n7579 = n1493 & n3475;
  assign n7580 = ~n7577 & ~n7578;
  assign n7581 = ~n7576 & n7580;
  assign n7582 = ~n7579 & n7581;
  assign n7583 = pi20  & n7582;
  assign n7584 = ~pi20  & ~n7582;
  assign n7585 = ~n7583 & ~n7584;
  assign n7586 = ~n7491 & ~n7494;
  assign n7587 = pi90  & n2053;
  assign n7588 = pi91  & n1893;
  assign n7589 = pi92  & n1888;
  assign n7590 = n1886 & n2924;
  assign n7591 = ~n7588 & ~n7589;
  assign n7592 = ~n7587 & n7591;
  assign n7593 = ~n7590 & n7592;
  assign n7594 = pi23  & n7593;
  assign n7595 = ~pi23  & ~n7593;
  assign n7596 = ~n7594 & ~n7595;
  assign n7597 = ~n7476 & ~n7478;
  assign n7598 = ~n7459 & ~n7463;
  assign n7599 = ~n7443 & ~n7447;
  assign n7600 = ~n7427 & ~n7430;
  assign n7601 = ~n7421 & ~n7424;
  assign n7602 = pi75  & n4843;
  assign n7603 = pi76  & n4598;
  assign n7604 = pi77  & n4593;
  assign n7605 = n865 & n4591;
  assign n7606 = ~n7603 & ~n7604;
  assign n7607 = ~n7602 & n7606;
  assign n7608 = ~n7605 & n7607;
  assign n7609 = pi38  & n7608;
  assign n7610 = ~pi38  & ~n7608;
  assign n7611 = ~n7609 & ~n7610;
  assign n7612 = ~n7416 & ~n7418;
  assign n7613 = ~n7399 & ~n7403;
  assign n7614 = ~n7383 & ~n7386;
  assign n7615 = pi66  & n7121;
  assign n7616 = pi67  & n6795;
  assign n7617 = pi68  & n6790;
  assign n7618 = n334 & n6788;
  assign n7619 = ~n7616 & ~n7617;
  assign n7620 = ~n7615 & n7619;
  assign n7621 = ~n7618 & n7620;
  assign n7622 = pi47  & n7621;
  assign n7623 = ~pi47  & ~n7621;
  assign n7624 = ~n7622 & ~n7623;
  assign n7625 = pi50  & n7381;
  assign n7626 = ~pi49  & ~pi50 ;
  assign n7627 = pi49  & pi50 ;
  assign n7628 = ~n7626 & ~n7627;
  assign n7629 = n7380 & n7628;
  assign n7630 = n265 & n7629;
  assign n7631 = n7380 & ~n7628;
  assign n7632 = pi65  & n7631;
  assign n7633 = ~pi48  & ~pi49 ;
  assign n7634 = pi48  & pi49 ;
  assign n7635 = ~n7633 & ~n7634;
  assign n7636 = ~n7380 & n7635;
  assign n7637 = pi64  & n7636;
  assign n7638 = ~n7630 & ~n7632;
  assign n7639 = ~n7637 & n7638;
  assign n7640 = n7625 & ~n7639;
  assign n7641 = ~n7625 & n7639;
  assign n7642 = ~n7640 & ~n7641;
  assign n7643 = n7624 & ~n7642;
  assign n7644 = ~n7624 & n7642;
  assign n7645 = ~n7643 & ~n7644;
  assign n7646 = ~n7614 & n7645;
  assign n7647 = n7614 & ~n7645;
  assign n7648 = ~n7646 & ~n7647;
  assign n7649 = pi69  & n6331;
  assign n7650 = pi70  & n6015;
  assign n7651 = pi71  & n6010;
  assign n7652 = n460 & n6008;
  assign n7653 = ~n7650 & ~n7651;
  assign n7654 = ~n7649 & n7653;
  assign n7655 = ~n7652 & n7654;
  assign n7656 = pi44  & n7655;
  assign n7657 = ~pi44  & ~n7655;
  assign n7658 = ~n7656 & ~n7657;
  assign n7659 = n7648 & ~n7658;
  assign n7660 = ~n7648 & n7658;
  assign n7661 = ~n7659 & ~n7660;
  assign n7662 = n7613 & ~n7661;
  assign n7663 = ~n7613 & n7661;
  assign n7664 = ~n7662 & ~n7663;
  assign n7665 = pi72  & n5558;
  assign n7666 = pi73  & n5293;
  assign n7667 = pi74  & n5288;
  assign n7668 = n689 & n5286;
  assign n7669 = ~n7666 & ~n7667;
  assign n7670 = ~n7665 & n7669;
  assign n7671 = ~n7668 & n7670;
  assign n7672 = pi41  & n7671;
  assign n7673 = ~pi41  & ~n7671;
  assign n7674 = ~n7672 & ~n7673;
  assign n7675 = n7664 & ~n7674;
  assign n7676 = ~n7664 & n7674;
  assign n7677 = ~n7675 & ~n7676;
  assign n7678 = ~n7612 & n7677;
  assign n7679 = n7612 & ~n7677;
  assign n7680 = ~n7678 & ~n7679;
  assign n7681 = n7611 & ~n7680;
  assign n7682 = ~n7611 & n7680;
  assign n7683 = ~n7681 & ~n7682;
  assign n7684 = ~n7601 & n7683;
  assign n7685 = n7601 & ~n7683;
  assign n7686 = ~n7684 & ~n7685;
  assign n7687 = pi78  & n4176;
  assign n7688 = pi79  & n3938;
  assign n7689 = pi80  & n3933;
  assign n7690 = n1144 & n3931;
  assign n7691 = ~n7688 & ~n7689;
  assign n7692 = ~n7687 & n7691;
  assign n7693 = ~n7690 & n7692;
  assign n7694 = pi35  & n7693;
  assign n7695 = ~pi35  & ~n7693;
  assign n7696 = ~n7694 & ~n7695;
  assign n7697 = n7686 & ~n7696;
  assign n7698 = ~n7686 & n7696;
  assign n7699 = ~n7697 & ~n7698;
  assign n7700 = n7600 & ~n7699;
  assign n7701 = ~n7600 & n7699;
  assign n7702 = ~n7700 & ~n7701;
  assign n7703 = pi81  & n3553;
  assign n7704 = pi82  & n3334;
  assign n7705 = pi83  & n3329;
  assign n7706 = n1577 & n3327;
  assign n7707 = ~n7704 & ~n7705;
  assign n7708 = ~n7703 & n7707;
  assign n7709 = ~n7706 & n7708;
  assign n7710 = pi32  & n7709;
  assign n7711 = ~pi32  & ~n7709;
  assign n7712 = ~n7710 & ~n7711;
  assign n7713 = n7702 & ~n7712;
  assign n7714 = ~n7702 & n7712;
  assign n7715 = ~n7713 & ~n7714;
  assign n7716 = n7599 & ~n7715;
  assign n7717 = ~n7599 & n7715;
  assign n7718 = ~n7716 & ~n7717;
  assign n7719 = pi84  & n3011;
  assign n7720 = pi85  & n2809;
  assign n7721 = pi86  & n2804;
  assign n7722 = n1975 & n2802;
  assign n7723 = ~n7720 & ~n7721;
  assign n7724 = ~n7719 & n7723;
  assign n7725 = ~n7722 & n7724;
  assign n7726 = pi29  & n7725;
  assign n7727 = ~pi29  & ~n7725;
  assign n7728 = ~n7726 & ~n7727;
  assign n7729 = n7718 & ~n7728;
  assign n7730 = ~n7718 & n7728;
  assign n7731 = ~n7729 & ~n7730;
  assign n7732 = n7598 & ~n7731;
  assign n7733 = ~n7598 & n7731;
  assign n7734 = ~n7732 & ~n7733;
  assign n7735 = pi87  & n2510;
  assign n7736 = pi88  & n2342;
  assign n7737 = pi89  & n2337;
  assign n7738 = n2287 & n2335;
  assign n7739 = ~n7736 & ~n7737;
  assign n7740 = ~n7735 & n7739;
  assign n7741 = ~n7738 & n7740;
  assign n7742 = pi26  & n7741;
  assign n7743 = ~pi26  & ~n7741;
  assign n7744 = ~n7742 & ~n7743;
  assign n7745 = n7734 & ~n7744;
  assign n7746 = ~n7734 & n7744;
  assign n7747 = ~n7745 & ~n7746;
  assign n7748 = ~n7597 & n7747;
  assign n7749 = n7597 & ~n7747;
  assign n7750 = ~n7748 & ~n7749;
  assign n7751 = ~n7596 & n7750;
  assign n7752 = n7596 & ~n7750;
  assign n7753 = ~n7751 & ~n7752;
  assign n7754 = ~n7586 & n7753;
  assign n7755 = n7586 & ~n7753;
  assign n7756 = ~n7754 & ~n7755;
  assign n7757 = ~n7585 & n7756;
  assign n7758 = n7585 & ~n7756;
  assign n7759 = ~n7757 & ~n7758;
  assign n7760 = n7575 & ~n7759;
  assign n7761 = ~n7575 & n7759;
  assign n7762 = ~n7760 & ~n7761;
  assign n7763 = pi96  & n1296;
  assign n7764 = pi97  & n1207;
  assign n7765 = pi98  & n1202;
  assign n7766 = n1200 & n3889;
  assign n7767 = ~n7764 & ~n7765;
  assign n7768 = ~n7763 & n7767;
  assign n7769 = ~n7766 & n7768;
  assign n7770 = pi17  & n7769;
  assign n7771 = ~pi17  & ~n7769;
  assign n7772 = ~n7770 & ~n7771;
  assign n7773 = n7762 & ~n7772;
  assign n7774 = ~n7762 & n7772;
  assign n7775 = ~n7773 & ~n7774;
  assign n7776 = n7574 & ~n7775;
  assign n7777 = ~n7574 & n7775;
  assign n7778 = ~n7776 & ~n7777;
  assign n7779 = pi99  & n1006;
  assign n7780 = pi100  & n897;
  assign n7781 = pi101  & n892;
  assign n7782 = n890 & n4730;
  assign n7783 = ~n7780 & ~n7781;
  assign n7784 = ~n7779 & n7783;
  assign n7785 = ~n7782 & n7784;
  assign n7786 = pi14  & n7785;
  assign n7787 = ~pi14  & ~n7785;
  assign n7788 = ~n7786 & ~n7787;
  assign n7789 = n7778 & ~n7788;
  assign n7790 = ~n7778 & n7788;
  assign n7791 = ~n7789 & ~n7790;
  assign n7792 = n7573 & ~n7791;
  assign n7793 = ~n7573 & n7791;
  assign n7794 = ~n7792 & ~n7793;
  assign n7795 = pi102  & n750;
  assign n7796 = pi103  & n651;
  assign n7797 = pi104  & n646;
  assign n7798 = n644 & n5212;
  assign n7799 = ~n7796 & ~n7797;
  assign n7800 = ~n7795 & n7799;
  assign n7801 = ~n7798 & n7800;
  assign n7802 = pi11  & n7801;
  assign n7803 = ~pi11  & ~n7801;
  assign n7804 = ~n7802 & ~n7803;
  assign n7805 = n7794 & ~n7804;
  assign n7806 = ~n7794 & n7804;
  assign n7807 = ~n7805 & ~n7806;
  assign n7808 = n7572 & ~n7807;
  assign n7809 = ~n7572 & n7807;
  assign n7810 = ~n7808 & ~n7809;
  assign n7811 = pi105  & n528;
  assign n7812 = pi106  & n490;
  assign n7813 = pi107  & n485;
  assign n7814 = n483 & n6189;
  assign n7815 = ~n7812 & ~n7813;
  assign n7816 = ~n7811 & n7815;
  assign n7817 = ~n7814 & n7816;
  assign n7818 = pi8  & n7817;
  assign n7819 = ~pi8  & ~n7817;
  assign n7820 = ~n7818 & ~n7819;
  assign n7821 = n7810 & ~n7820;
  assign n7822 = ~n7810 & n7820;
  assign n7823 = ~n7821 & ~n7822;
  assign n7824 = n7571 & ~n7823;
  assign n7825 = ~n7571 & n7823;
  assign n7826 = ~n7824 & ~n7825;
  assign n7827 = pi108  & n391;
  assign n7828 = pi109  & n353;
  assign n7829 = pi110  & n348;
  assign n7830 = n346 & n6995;
  assign n7831 = ~n7828 & ~n7829;
  assign n7832 = ~n7827 & n7831;
  assign n7833 = ~n7830 & n7832;
  assign n7834 = pi5  & n7833;
  assign n7835 = ~pi5  & ~n7833;
  assign n7836 = ~n7834 & ~n7835;
  assign n7837 = n7826 & ~n7836;
  assign n7838 = ~n7826 & n7836;
  assign n7839 = ~n7837 & ~n7838;
  assign n7840 = n7570 & ~n7839;
  assign n7841 = ~n7570 & n7839;
  assign n7842 = ~n7840 & ~n7841;
  assign n7843 = pi113  & n269;
  assign n7844 = pi112  & n267;
  assign n7845 = pi111  & n282;
  assign n7846 = ~n7292 & ~n7294;
  assign n7847 = ~pi112  & ~pi113 ;
  assign n7848 = pi112  & pi113 ;
  assign n7849 = ~n7847 & ~n7848;
  assign n7850 = ~n7846 & n7849;
  assign n7851 = n7846 & ~n7849;
  assign n7852 = ~n7850 & ~n7851;
  assign n7853 = n262 & n7852;
  assign n7854 = ~n7843 & ~n7844;
  assign n7855 = ~n7845 & n7854;
  assign n7856 = ~n7853 & n7855;
  assign n7857 = pi2  & n7856;
  assign n7858 = ~pi2  & ~n7856;
  assign n7859 = ~n7857 & ~n7858;
  assign n7860 = ~n7842 & n7859;
  assign n7861 = n7842 & ~n7859;
  assign n7862 = ~n7860 & ~n7861;
  assign n7863 = ~n7569 & n7862;
  assign n7864 = n7569 & ~n7862;
  assign po49  = ~n7863 & ~n7864;
  assign n7866 = ~n7861 & ~n7863;
  assign n7867 = ~n7837 & ~n7841;
  assign n7868 = ~n7821 & ~n7825;
  assign n7869 = ~n7805 & ~n7809;
  assign n7870 = ~n7789 & ~n7793;
  assign n7871 = ~n7773 & ~n7777;
  assign n7872 = ~n7757 & ~n7761;
  assign n7873 = pi94  & n1661;
  assign n7874 = pi95  & n1500;
  assign n7875 = pi96  & n1495;
  assign n7876 = n1493 & n3499;
  assign n7877 = ~n7874 & ~n7875;
  assign n7878 = ~n7873 & n7877;
  assign n7879 = ~n7876 & n7878;
  assign n7880 = pi20  & n7879;
  assign n7881 = ~pi20  & ~n7879;
  assign n7882 = ~n7880 & ~n7881;
  assign n7883 = ~n7751 & ~n7754;
  assign n7884 = pi91  & n2053;
  assign n7885 = pi92  & n1893;
  assign n7886 = pi93  & n1888;
  assign n7887 = n1886 & n2948;
  assign n7888 = ~n7885 & ~n7886;
  assign n7889 = ~n7884 & n7888;
  assign n7890 = ~n7887 & n7889;
  assign n7891 = pi23  & n7890;
  assign n7892 = ~pi23  & ~n7890;
  assign n7893 = ~n7891 & ~n7892;
  assign n7894 = ~n7745 & ~n7748;
  assign n7895 = pi88  & n2510;
  assign n7896 = pi89  & n2342;
  assign n7897 = pi90  & n2337;
  assign n7898 = n2335 & n2448;
  assign n7899 = ~n7896 & ~n7897;
  assign n7900 = ~n7895 & n7899;
  assign n7901 = ~n7898 & n7900;
  assign n7902 = pi26  & n7901;
  assign n7903 = ~pi26  & ~n7901;
  assign n7904 = ~n7902 & ~n7903;
  assign n7905 = ~n7729 & ~n7733;
  assign n7906 = ~n7713 & ~n7717;
  assign n7907 = pi82  & n3553;
  assign n7908 = pi83  & n3334;
  assign n7909 = pi84  & n3329;
  assign n7910 = n1601 & n3327;
  assign n7911 = ~n7908 & ~n7909;
  assign n7912 = ~n7907 & n7911;
  assign n7913 = ~n7910 & n7912;
  assign n7914 = pi32  & n7913;
  assign n7915 = ~pi32  & ~n7913;
  assign n7916 = ~n7914 & ~n7915;
  assign n7917 = ~n7697 & ~n7701;
  assign n7918 = pi79  & n4176;
  assign n7919 = pi80  & n3938;
  assign n7920 = pi81  & n3933;
  assign n7921 = n1337 & n3931;
  assign n7922 = ~n7919 & ~n7920;
  assign n7923 = ~n7918 & n7922;
  assign n7924 = ~n7921 & n7923;
  assign n7925 = pi35  & n7924;
  assign n7926 = ~pi35  & ~n7924;
  assign n7927 = ~n7925 & ~n7926;
  assign n7928 = ~n7682 & ~n7684;
  assign n7929 = ~n7675 & ~n7678;
  assign n7930 = pi73  & n5558;
  assign n7931 = pi74  & n5293;
  assign n7932 = pi75  & n5288;
  assign n7933 = n713 & n5286;
  assign n7934 = ~n7931 & ~n7932;
  assign n7935 = ~n7930 & n7934;
  assign n7936 = ~n7933 & n7935;
  assign n7937 = pi41  & n7936;
  assign n7938 = ~pi41  & ~n7936;
  assign n7939 = ~n7937 & ~n7938;
  assign n7940 = ~n7659 & ~n7663;
  assign n7941 = pi70  & n6331;
  assign n7942 = pi71  & n6015;
  assign n7943 = pi72  & n6010;
  assign n7944 = n551 & n6008;
  assign n7945 = ~n7942 & ~n7943;
  assign n7946 = ~n7941 & n7945;
  assign n7947 = ~n7944 & n7946;
  assign n7948 = pi44  & n7947;
  assign n7949 = ~pi44  & ~n7947;
  assign n7950 = ~n7948 & ~n7949;
  assign n7951 = ~n7644 & ~n7646;
  assign n7952 = pi67  & n7121;
  assign n7953 = pi68  & n6795;
  assign n7954 = pi69  & n6790;
  assign n7955 = n376 & n6788;
  assign n7956 = ~n7953 & ~n7954;
  assign n7957 = ~n7952 & n7956;
  assign n7958 = ~n7955 & n7957;
  assign n7959 = pi47  & n7958;
  assign n7960 = ~pi47  & ~n7958;
  assign n7961 = ~n7959 & ~n7960;
  assign n7962 = pi50  & ~n7381;
  assign n7963 = n7639 & n7962;
  assign n7964 = pi50  & ~n7963;
  assign n7965 = ~n287 & n7629;
  assign n7966 = pi65  & n7636;
  assign n7967 = pi66  & n7631;
  assign n7968 = ~n7380 & n7628;
  assign n7969 = ~n7635 & n7968;
  assign n7970 = pi64  & n7969;
  assign n7971 = ~n7965 & ~n7966;
  assign n7972 = ~n7967 & n7971;
  assign n7973 = ~n7970 & n7972;
  assign n7974 = ~n7964 & n7973;
  assign n7975 = n7964 & ~n7973;
  assign n7976 = ~n7974 & ~n7975;
  assign n7977 = ~n7961 & n7976;
  assign n7978 = n7961 & ~n7976;
  assign n7979 = ~n7977 & ~n7978;
  assign n7980 = ~n7951 & n7979;
  assign n7981 = n7951 & ~n7979;
  assign n7982 = ~n7980 & ~n7981;
  assign n7983 = ~n7950 & n7982;
  assign n7984 = n7950 & ~n7982;
  assign n7985 = ~n7983 & ~n7984;
  assign n7986 = ~n7940 & n7985;
  assign n7987 = n7940 & ~n7985;
  assign n7988 = ~n7986 & ~n7987;
  assign n7989 = n7939 & ~n7988;
  assign n7990 = ~n7939 & n7988;
  assign n7991 = ~n7989 & ~n7990;
  assign n7992 = ~n7929 & n7991;
  assign n7993 = n7929 & ~n7991;
  assign n7994 = ~n7992 & ~n7993;
  assign n7995 = pi76  & n4843;
  assign n7996 = pi77  & n4598;
  assign n7997 = pi78  & n4593;
  assign n7998 = n958 & n4591;
  assign n7999 = ~n7996 & ~n7997;
  assign n8000 = ~n7995 & n7999;
  assign n8001 = ~n7998 & n8000;
  assign n8002 = pi38  & n8001;
  assign n8003 = ~pi38  & ~n8001;
  assign n8004 = ~n8002 & ~n8003;
  assign n8005 = n7994 & ~n8004;
  assign n8006 = ~n7994 & n8004;
  assign n8007 = ~n8005 & ~n8006;
  assign n8008 = ~n7928 & n8007;
  assign n8009 = n7928 & ~n8007;
  assign n8010 = ~n8008 & ~n8009;
  assign n8011 = ~n7927 & n8010;
  assign n8012 = n7927 & ~n8010;
  assign n8013 = ~n8011 & ~n8012;
  assign n8014 = ~n7917 & n8013;
  assign n8015 = n7917 & ~n8013;
  assign n8016 = ~n8014 & ~n8015;
  assign n8017 = ~n7916 & n8016;
  assign n8018 = n7916 & ~n8016;
  assign n8019 = ~n8017 & ~n8018;
  assign n8020 = n7906 & ~n8019;
  assign n8021 = ~n7906 & n8019;
  assign n8022 = ~n8020 & ~n8021;
  assign n8023 = pi85  & n3011;
  assign n8024 = pi86  & n2809;
  assign n8025 = pi87  & n2804;
  assign n8026 = n2116 & n2802;
  assign n8027 = ~n8024 & ~n8025;
  assign n8028 = ~n8023 & n8027;
  assign n8029 = ~n8026 & n8028;
  assign n8030 = pi29  & n8029;
  assign n8031 = ~pi29  & ~n8029;
  assign n8032 = ~n8030 & ~n8031;
  assign n8033 = n8022 & ~n8032;
  assign n8034 = ~n8022 & n8032;
  assign n8035 = ~n8033 & ~n8034;
  assign n8036 = ~n7905 & n8035;
  assign n8037 = n7905 & ~n8035;
  assign n8038 = ~n8036 & ~n8037;
  assign n8039 = n7904 & ~n8038;
  assign n8040 = ~n7904 & n8038;
  assign n8041 = ~n8039 & ~n8040;
  assign n8042 = ~n7894 & n8041;
  assign n8043 = n7894 & ~n8041;
  assign n8044 = ~n8042 & ~n8043;
  assign n8045 = n7893 & ~n8044;
  assign n8046 = ~n7893 & n8044;
  assign n8047 = ~n8045 & ~n8046;
  assign n8048 = ~n7883 & n8047;
  assign n8049 = n7883 & ~n8047;
  assign n8050 = ~n8048 & ~n8049;
  assign n8051 = n7882 & ~n8050;
  assign n8052 = ~n7882 & n8050;
  assign n8053 = ~n8051 & ~n8052;
  assign n8054 = ~n7872 & n8053;
  assign n8055 = n7872 & ~n8053;
  assign n8056 = ~n8054 & ~n8055;
  assign n8057 = pi97  & n1296;
  assign n8058 = pi98  & n1207;
  assign n8059 = pi99  & n1202;
  assign n8060 = n1200 & n4101;
  assign n8061 = ~n8058 & ~n8059;
  assign n8062 = ~n8057 & n8061;
  assign n8063 = ~n8060 & n8062;
  assign n8064 = pi17  & n8063;
  assign n8065 = ~pi17  & ~n8063;
  assign n8066 = ~n8064 & ~n8065;
  assign n8067 = n8056 & ~n8066;
  assign n8068 = ~n8056 & n8066;
  assign n8069 = ~n8067 & ~n8068;
  assign n8070 = n7871 & ~n8069;
  assign n8071 = ~n7871 & n8069;
  assign n8072 = ~n8070 & ~n8071;
  assign n8073 = pi100  & n1006;
  assign n8074 = pi101  & n897;
  assign n8075 = pi102  & n892;
  assign n8076 = n890 & n4956;
  assign n8077 = ~n8074 & ~n8075;
  assign n8078 = ~n8073 & n8077;
  assign n8079 = ~n8076 & n8078;
  assign n8080 = pi14  & n8079;
  assign n8081 = ~pi14  & ~n8079;
  assign n8082 = ~n8080 & ~n8081;
  assign n8083 = n8072 & ~n8082;
  assign n8084 = ~n8072 & n8082;
  assign n8085 = ~n8083 & ~n8084;
  assign n8086 = n7870 & ~n8085;
  assign n8087 = ~n7870 & n8085;
  assign n8088 = ~n8086 & ~n8087;
  assign n8089 = pi103  & n750;
  assign n8090 = pi104  & n651;
  assign n8091 = pi105  & n646;
  assign n8092 = n644 & n5677;
  assign n8093 = ~n8090 & ~n8091;
  assign n8094 = ~n8089 & n8093;
  assign n8095 = ~n8092 & n8094;
  assign n8096 = pi11  & n8095;
  assign n8097 = ~pi11  & ~n8095;
  assign n8098 = ~n8096 & ~n8097;
  assign n8099 = n8088 & ~n8098;
  assign n8100 = ~n8088 & n8098;
  assign n8101 = ~n8099 & ~n8100;
  assign n8102 = n7869 & ~n8101;
  assign n8103 = ~n7869 & n8101;
  assign n8104 = ~n8102 & ~n8103;
  assign n8105 = pi106  & n528;
  assign n8106 = pi107  & n490;
  assign n8107 = pi108  & n485;
  assign n8108 = n483 & n6213;
  assign n8109 = ~n8106 & ~n8107;
  assign n8110 = ~n8105 & n8109;
  assign n8111 = ~n8108 & n8110;
  assign n8112 = pi8  & n8111;
  assign n8113 = ~pi8  & ~n8111;
  assign n8114 = ~n8112 & ~n8113;
  assign n8115 = n8104 & ~n8114;
  assign n8116 = ~n8104 & n8114;
  assign n8117 = ~n8115 & ~n8116;
  assign n8118 = ~n7868 & n8117;
  assign n8119 = n7868 & ~n8117;
  assign n8120 = ~n8118 & ~n8119;
  assign n8121 = pi109  & n391;
  assign n8122 = pi110  & n353;
  assign n8123 = pi111  & n348;
  assign n8124 = n346 & n7272;
  assign n8125 = ~n8122 & ~n8123;
  assign n8126 = ~n8121 & n8125;
  assign n8127 = ~n8124 & n8126;
  assign n8128 = pi5  & n8127;
  assign n8129 = ~pi5  & ~n8127;
  assign n8130 = ~n8128 & ~n8129;
  assign n8131 = n8120 & ~n8130;
  assign n8132 = ~n8120 & n8130;
  assign n8133 = ~n8131 & ~n8132;
  assign n8134 = n7867 & ~n8133;
  assign n8135 = ~n7867 & n8133;
  assign n8136 = ~n8134 & ~n8135;
  assign n8137 = pi114  & n269;
  assign n8138 = pi113  & n267;
  assign n8139 = pi112  & n282;
  assign n8140 = ~n7848 & ~n7850;
  assign n8141 = ~pi113  & ~pi114 ;
  assign n8142 = pi113  & pi114 ;
  assign n8143 = ~n8141 & ~n8142;
  assign n8144 = ~n8140 & n8143;
  assign n8145 = n8140 & ~n8143;
  assign n8146 = ~n8144 & ~n8145;
  assign n8147 = n262 & n8146;
  assign n8148 = ~n8137 & ~n8138;
  assign n8149 = ~n8139 & n8148;
  assign n8150 = ~n8147 & n8149;
  assign n8151 = pi2  & n8150;
  assign n8152 = ~pi2  & ~n8150;
  assign n8153 = ~n8151 & ~n8152;
  assign n8154 = n8136 & ~n8153;
  assign n8155 = ~n8136 & n8153;
  assign n8156 = ~n8154 & ~n8155;
  assign n8157 = ~n7866 & n8156;
  assign n8158 = n7866 & ~n8156;
  assign po50  = ~n8157 & ~n8158;
  assign n8160 = ~n8154 & ~n8157;
  assign n8161 = pi115  & n269;
  assign n8162 = pi114  & n267;
  assign n8163 = pi113  & n282;
  assign n8164 = ~n8142 & ~n8144;
  assign n8165 = ~pi114  & ~pi115 ;
  assign n8166 = pi114  & pi115 ;
  assign n8167 = ~n8165 & ~n8166;
  assign n8168 = ~n8164 & n8167;
  assign n8169 = n8164 & ~n8167;
  assign n8170 = ~n8168 & ~n8169;
  assign n8171 = n262 & n8170;
  assign n8172 = ~n8161 & ~n8162;
  assign n8173 = ~n8163 & n8172;
  assign n8174 = ~n8171 & n8173;
  assign n8175 = pi2  & n8174;
  assign n8176 = ~pi2  & ~n8174;
  assign n8177 = ~n8175 & ~n8176;
  assign n8178 = ~n8131 & ~n8135;
  assign n8179 = pi110  & n391;
  assign n8180 = pi111  & n353;
  assign n8181 = pi112  & n348;
  assign n8182 = n346 & n7296;
  assign n8183 = ~n8180 & ~n8181;
  assign n8184 = ~n8179 & n8183;
  assign n8185 = ~n8182 & n8184;
  assign n8186 = pi5  & n8185;
  assign n8187 = ~pi5  & ~n8185;
  assign n8188 = ~n8186 & ~n8187;
  assign n8189 = ~n8115 & ~n8118;
  assign n8190 = ~n8083 & ~n8087;
  assign n8191 = ~n8067 & ~n8071;
  assign n8192 = pi98  & n1296;
  assign n8193 = pi99  & n1207;
  assign n8194 = pi100  & n1202;
  assign n8195 = n1200 & n4501;
  assign n8196 = ~n8193 & ~n8194;
  assign n8197 = ~n8192 & n8196;
  assign n8198 = ~n8195 & n8197;
  assign n8199 = pi17  & n8198;
  assign n8200 = ~pi17  & ~n8198;
  assign n8201 = ~n8199 & ~n8200;
  assign n8202 = ~n8052 & ~n8054;
  assign n8203 = ~n8046 & ~n8048;
  assign n8204 = pi92  & n2053;
  assign n8205 = pi93  & n1893;
  assign n8206 = pi94  & n1888;
  assign n8207 = n1886 & n3280;
  assign n8208 = ~n8205 & ~n8206;
  assign n8209 = ~n8204 & n8208;
  assign n8210 = ~n8207 & n8209;
  assign n8211 = pi23  & n8210;
  assign n8212 = ~pi23  & ~n8210;
  assign n8213 = ~n8211 & ~n8212;
  assign n8214 = ~n8040 & ~n8042;
  assign n8215 = ~n8033 & ~n8036;
  assign n8216 = ~n8017 & ~n8021;
  assign n8217 = ~n8011 & ~n8014;
  assign n8218 = pi80  & n4176;
  assign n8219 = pi81  & n3938;
  assign n8220 = pi82  & n3933;
  assign n8221 = n1450 & n3931;
  assign n8222 = ~n8219 & ~n8220;
  assign n8223 = ~n8218 & n8222;
  assign n8224 = ~n8221 & n8223;
  assign n8225 = pi35  & n8224;
  assign n8226 = ~pi35  & ~n8224;
  assign n8227 = ~n8225 & ~n8226;
  assign n8228 = ~n8005 & ~n8008;
  assign n8229 = pi77  & n4843;
  assign n8230 = pi78  & n4598;
  assign n8231 = pi79  & n4593;
  assign n8232 = n1048 & n4591;
  assign n8233 = ~n8230 & ~n8231;
  assign n8234 = ~n8229 & n8233;
  assign n8235 = ~n8232 & n8234;
  assign n8236 = pi38  & n8235;
  assign n8237 = ~pi38  & ~n8235;
  assign n8238 = ~n8236 & ~n8237;
  assign n8239 = ~n7990 & ~n7992;
  assign n8240 = pi74  & n5558;
  assign n8241 = pi75  & n5293;
  assign n8242 = pi76  & n5288;
  assign n8243 = n841 & n5286;
  assign n8244 = ~n8241 & ~n8242;
  assign n8245 = ~n8240 & n8244;
  assign n8246 = ~n8243 & n8245;
  assign n8247 = pi41  & n8246;
  assign n8248 = ~pi41  & ~n8246;
  assign n8249 = ~n8247 & ~n8248;
  assign n8250 = ~n7983 & ~n7986;
  assign n8251 = ~n7977 & ~n7980;
  assign n8252 = pi65  & n7969;
  assign n8253 = pi66  & n7636;
  assign n8254 = pi67  & n7631;
  assign n8255 = n305 & n7629;
  assign n8256 = ~n8253 & ~n8254;
  assign n8257 = ~n8252 & n8256;
  assign n8258 = ~n8255 & n8257;
  assign n8259 = pi50  & n8258;
  assign n8260 = ~pi50  & ~n8258;
  assign n8261 = ~n8259 & ~n8260;
  assign n8262 = ~pi50  & ~pi51 ;
  assign n8263 = pi50  & pi51 ;
  assign n8264 = ~n8262 & ~n8263;
  assign n8265 = pi64  & n8264;
  assign n8266 = n7963 & n7973;
  assign n8267 = n8265 & n8266;
  assign n8268 = ~n8265 & ~n8266;
  assign n8269 = ~n8267 & ~n8268;
  assign n8270 = ~n8261 & n8269;
  assign n8271 = n8261 & ~n8269;
  assign n8272 = ~n8270 & ~n8271;
  assign n8273 = pi68  & n7121;
  assign n8274 = pi69  & n6795;
  assign n8275 = pi70  & n6790;
  assign n8276 = n415 & n6788;
  assign n8277 = ~n8274 & ~n8275;
  assign n8278 = ~n8273 & n8277;
  assign n8279 = ~n8276 & n8278;
  assign n8280 = pi47  & n8279;
  assign n8281 = ~pi47  & ~n8279;
  assign n8282 = ~n8280 & ~n8281;
  assign n8283 = n8272 & ~n8282;
  assign n8284 = ~n8272 & n8282;
  assign n8285 = ~n8283 & ~n8284;
  assign n8286 = n8251 & ~n8285;
  assign n8287 = ~n8251 & n8285;
  assign n8288 = ~n8286 & ~n8287;
  assign n8289 = pi71  & n6331;
  assign n8290 = pi72  & n6015;
  assign n8291 = pi73  & n6010;
  assign n8292 = n613 & n6008;
  assign n8293 = ~n8290 & ~n8291;
  assign n8294 = ~n8289 & n8293;
  assign n8295 = ~n8292 & n8294;
  assign n8296 = pi44  & n8295;
  assign n8297 = ~pi44  & ~n8295;
  assign n8298 = ~n8296 & ~n8297;
  assign n8299 = ~n8288 & n8298;
  assign n8300 = n8288 & ~n8298;
  assign n8301 = ~n8299 & ~n8300;
  assign n8302 = ~n8250 & n8301;
  assign n8303 = n8250 & ~n8301;
  assign n8304 = ~n8302 & ~n8303;
  assign n8305 = ~n8249 & n8304;
  assign n8306 = n8249 & ~n8304;
  assign n8307 = ~n8305 & ~n8306;
  assign n8308 = ~n8239 & n8307;
  assign n8309 = n8239 & ~n8307;
  assign n8310 = ~n8308 & ~n8309;
  assign n8311 = ~n8238 & n8310;
  assign n8312 = n8238 & ~n8310;
  assign n8313 = ~n8311 & ~n8312;
  assign n8314 = ~n8228 & n8313;
  assign n8315 = n8228 & ~n8313;
  assign n8316 = ~n8314 & ~n8315;
  assign n8317 = ~n8227 & n8316;
  assign n8318 = n8227 & ~n8316;
  assign n8319 = ~n8317 & ~n8318;
  assign n8320 = ~n8217 & n8319;
  assign n8321 = n8217 & ~n8319;
  assign n8322 = ~n8320 & ~n8321;
  assign n8323 = pi83  & n3553;
  assign n8324 = pi84  & n3334;
  assign n8325 = pi85  & n3329;
  assign n8326 = n1831 & n3327;
  assign n8327 = ~n8324 & ~n8325;
  assign n8328 = ~n8323 & n8327;
  assign n8329 = ~n8326 & n8328;
  assign n8330 = pi32  & n8329;
  assign n8331 = ~pi32  & ~n8329;
  assign n8332 = ~n8330 & ~n8331;
  assign n8333 = n8322 & ~n8332;
  assign n8334 = ~n8322 & n8332;
  assign n8335 = ~n8333 & ~n8334;
  assign n8336 = n8216 & ~n8335;
  assign n8337 = ~n8216 & n8335;
  assign n8338 = ~n8336 & ~n8337;
  assign n8339 = pi86  & n3011;
  assign n8340 = pi87  & n2809;
  assign n8341 = pi88  & n2804;
  assign n8342 = n2140 & n2802;
  assign n8343 = ~n8340 & ~n8341;
  assign n8344 = ~n8339 & n8343;
  assign n8345 = ~n8342 & n8344;
  assign n8346 = pi29  & n8345;
  assign n8347 = ~pi29  & ~n8345;
  assign n8348 = ~n8346 & ~n8347;
  assign n8349 = ~n8338 & n8348;
  assign n8350 = n8338 & ~n8348;
  assign n8351 = ~n8349 & ~n8350;
  assign n8352 = ~n8215 & n8351;
  assign n8353 = n8215 & ~n8351;
  assign n8354 = ~n8352 & ~n8353;
  assign n8355 = pi89  & n2510;
  assign n8356 = pi90  & n2342;
  assign n8357 = pi91  & n2337;
  assign n8358 = n2335 & n2746;
  assign n8359 = ~n8356 & ~n8357;
  assign n8360 = ~n8355 & n8359;
  assign n8361 = ~n8358 & n8360;
  assign n8362 = pi26  & n8361;
  assign n8363 = ~pi26  & ~n8361;
  assign n8364 = ~n8362 & ~n8363;
  assign n8365 = n8354 & ~n8364;
  assign n8366 = ~n8354 & n8364;
  assign n8367 = ~n8365 & ~n8366;
  assign n8368 = ~n8214 & n8367;
  assign n8369 = n8214 & ~n8367;
  assign n8370 = ~n8368 & ~n8369;
  assign n8371 = ~n8213 & n8370;
  assign n8372 = n8213 & ~n8370;
  assign n8373 = ~n8371 & ~n8372;
  assign n8374 = ~n8203 & n8373;
  assign n8375 = n8203 & ~n8373;
  assign n8376 = ~n8374 & ~n8375;
  assign n8377 = pi95  & n1661;
  assign n8378 = pi96  & n1500;
  assign n8379 = pi97  & n1495;
  assign n8380 = n1493 & n3691;
  assign n8381 = ~n8378 & ~n8379;
  assign n8382 = ~n8377 & n8381;
  assign n8383 = ~n8380 & n8382;
  assign n8384 = pi20  & n8383;
  assign n8385 = ~pi20  & ~n8383;
  assign n8386 = ~n8384 & ~n8385;
  assign n8387 = n8376 & ~n8386;
  assign n8388 = ~n8376 & n8386;
  assign n8389 = ~n8387 & ~n8388;
  assign n8390 = ~n8202 & n8389;
  assign n8391 = n8202 & ~n8389;
  assign n8392 = ~n8390 & ~n8391;
  assign n8393 = ~n8201 & n8392;
  assign n8394 = n8201 & ~n8392;
  assign n8395 = ~n8393 & ~n8394;
  assign n8396 = n8191 & ~n8395;
  assign n8397 = ~n8191 & n8395;
  assign n8398 = ~n8396 & ~n8397;
  assign n8399 = pi101  & n1006;
  assign n8400 = pi102  & n897;
  assign n8401 = pi103  & n892;
  assign n8402 = n890 & n5188;
  assign n8403 = ~n8400 & ~n8401;
  assign n8404 = ~n8399 & n8403;
  assign n8405 = ~n8402 & n8404;
  assign n8406 = pi14  & n8405;
  assign n8407 = ~pi14  & ~n8405;
  assign n8408 = ~n8406 & ~n8407;
  assign n8409 = n8398 & ~n8408;
  assign n8410 = ~n8398 & n8408;
  assign n8411 = ~n8409 & ~n8410;
  assign n8412 = n8190 & ~n8411;
  assign n8413 = ~n8190 & n8411;
  assign n8414 = ~n8412 & ~n8413;
  assign n8415 = pi104  & n750;
  assign n8416 = pi105  & n651;
  assign n8417 = pi106  & n646;
  assign n8418 = n644 & n5701;
  assign n8419 = ~n8416 & ~n8417;
  assign n8420 = ~n8415 & n8419;
  assign n8421 = ~n8418 & n8420;
  assign n8422 = pi11  & n8421;
  assign n8423 = ~pi11  & ~n8421;
  assign n8424 = ~n8422 & ~n8423;
  assign n8425 = ~n8414 & n8424;
  assign n8426 = n8414 & ~n8424;
  assign n8427 = ~n8425 & ~n8426;
  assign n8428 = ~n8099 & ~n8103;
  assign n8429 = n8427 & ~n8428;
  assign n8430 = ~n8427 & n8428;
  assign n8431 = ~n8429 & ~n8430;
  assign n8432 = pi107  & n528;
  assign n8433 = pi108  & n490;
  assign n8434 = pi109  & n485;
  assign n8435 = n483 & n6715;
  assign n8436 = ~n8433 & ~n8434;
  assign n8437 = ~n8432 & n8436;
  assign n8438 = ~n8435 & n8437;
  assign n8439 = pi8  & n8438;
  assign n8440 = ~pi8  & ~n8438;
  assign n8441 = ~n8439 & ~n8440;
  assign n8442 = n8431 & ~n8441;
  assign n8443 = ~n8431 & n8441;
  assign n8444 = ~n8442 & ~n8443;
  assign n8445 = ~n8189 & n8444;
  assign n8446 = n8189 & ~n8444;
  assign n8447 = ~n8445 & ~n8446;
  assign n8448 = n8188 & ~n8447;
  assign n8449 = ~n8188 & n8447;
  assign n8450 = ~n8448 & ~n8449;
  assign n8451 = ~n8178 & n8450;
  assign n8452 = n8178 & ~n8450;
  assign n8453 = ~n8451 & ~n8452;
  assign n8454 = ~n8177 & n8453;
  assign n8455 = n8177 & ~n8453;
  assign n8456 = ~n8454 & ~n8455;
  assign n8457 = ~n8160 & n8456;
  assign n8458 = n8160 & ~n8456;
  assign po51  = ~n8457 & ~n8458;
  assign n8460 = ~n8454 & ~n8457;
  assign n8461 = pi116  & n269;
  assign n8462 = pi115  & n267;
  assign n8463 = pi114  & n282;
  assign n8464 = ~n8166 & ~n8168;
  assign n8465 = ~pi115  & ~pi116 ;
  assign n8466 = pi115  & pi116 ;
  assign n8467 = ~n8465 & ~n8466;
  assign n8468 = ~n8464 & n8467;
  assign n8469 = n8464 & ~n8467;
  assign n8470 = ~n8468 & ~n8469;
  assign n8471 = n262 & n8470;
  assign n8472 = ~n8461 & ~n8462;
  assign n8473 = ~n8463 & n8472;
  assign n8474 = ~n8471 & n8473;
  assign n8475 = pi2  & n8474;
  assign n8476 = ~pi2  & ~n8474;
  assign n8477 = ~n8475 & ~n8476;
  assign n8478 = ~n8449 & ~n8451;
  assign n8479 = ~n8442 & ~n8445;
  assign n8480 = ~n8426 & ~n8429;
  assign n8481 = ~n8409 & ~n8413;
  assign n8482 = ~n8393 & ~n8397;
  assign n8483 = ~n8387 & ~n8390;
  assign n8484 = ~n8371 & ~n8374;
  assign n8485 = ~n8365 & ~n8368;
  assign n8486 = pi90  & n2510;
  assign n8487 = pi91  & n2342;
  assign n8488 = pi92  & n2337;
  assign n8489 = n2335 & n2924;
  assign n8490 = ~n8487 & ~n8488;
  assign n8491 = ~n8486 & n8490;
  assign n8492 = ~n8489 & n8491;
  assign n8493 = pi26  & n8492;
  assign n8494 = ~pi26  & ~n8492;
  assign n8495 = ~n8493 & ~n8494;
  assign n8496 = ~n8350 & ~n8352;
  assign n8497 = ~n8333 & ~n8337;
  assign n8498 = ~n8317 & ~n8320;
  assign n8499 = ~n8311 & ~n8314;
  assign n8500 = ~n8305 & ~n8308;
  assign n8501 = pi75  & n5558;
  assign n8502 = pi76  & n5293;
  assign n8503 = pi77  & n5288;
  assign n8504 = n865 & n5286;
  assign n8505 = ~n8502 & ~n8503;
  assign n8506 = ~n8501 & n8505;
  assign n8507 = ~n8504 & n8506;
  assign n8508 = pi41  & n8507;
  assign n8509 = ~pi41  & ~n8507;
  assign n8510 = ~n8508 & ~n8509;
  assign n8511 = ~n8300 & ~n8302;
  assign n8512 = ~n8283 & ~n8287;
  assign n8513 = ~n8267 & ~n8270;
  assign n8514 = pi66  & n7969;
  assign n8515 = pi67  & n7636;
  assign n8516 = pi68  & n7631;
  assign n8517 = n334 & n7629;
  assign n8518 = ~n8515 & ~n8516;
  assign n8519 = ~n8514 & n8518;
  assign n8520 = ~n8517 & n8519;
  assign n8521 = pi50  & n8520;
  assign n8522 = ~pi50  & ~n8520;
  assign n8523 = ~n8521 & ~n8522;
  assign n8524 = pi53  & n8265;
  assign n8525 = ~pi52  & ~pi53 ;
  assign n8526 = pi52  & pi53 ;
  assign n8527 = ~n8525 & ~n8526;
  assign n8528 = n8264 & n8527;
  assign n8529 = n265 & n8528;
  assign n8530 = n8264 & ~n8527;
  assign n8531 = pi65  & n8530;
  assign n8532 = ~pi51  & ~pi52 ;
  assign n8533 = pi51  & pi52 ;
  assign n8534 = ~n8532 & ~n8533;
  assign n8535 = ~n8264 & n8534;
  assign n8536 = pi64  & n8535;
  assign n8537 = ~n8529 & ~n8531;
  assign n8538 = ~n8536 & n8537;
  assign n8539 = n8524 & ~n8538;
  assign n8540 = ~n8524 & n8538;
  assign n8541 = ~n8539 & ~n8540;
  assign n8542 = n8523 & ~n8541;
  assign n8543 = ~n8523 & n8541;
  assign n8544 = ~n8542 & ~n8543;
  assign n8545 = ~n8513 & n8544;
  assign n8546 = n8513 & ~n8544;
  assign n8547 = ~n8545 & ~n8546;
  assign n8548 = pi69  & n7121;
  assign n8549 = pi70  & n6795;
  assign n8550 = pi71  & n6790;
  assign n8551 = n460 & n6788;
  assign n8552 = ~n8549 & ~n8550;
  assign n8553 = ~n8548 & n8552;
  assign n8554 = ~n8551 & n8553;
  assign n8555 = pi47  & n8554;
  assign n8556 = ~pi47  & ~n8554;
  assign n8557 = ~n8555 & ~n8556;
  assign n8558 = n8547 & ~n8557;
  assign n8559 = ~n8547 & n8557;
  assign n8560 = ~n8558 & ~n8559;
  assign n8561 = n8512 & ~n8560;
  assign n8562 = ~n8512 & n8560;
  assign n8563 = ~n8561 & ~n8562;
  assign n8564 = pi72  & n6331;
  assign n8565 = pi73  & n6015;
  assign n8566 = pi74  & n6010;
  assign n8567 = n689 & n6008;
  assign n8568 = ~n8565 & ~n8566;
  assign n8569 = ~n8564 & n8568;
  assign n8570 = ~n8567 & n8569;
  assign n8571 = pi44  & n8570;
  assign n8572 = ~pi44  & ~n8570;
  assign n8573 = ~n8571 & ~n8572;
  assign n8574 = n8563 & ~n8573;
  assign n8575 = ~n8563 & n8573;
  assign n8576 = ~n8574 & ~n8575;
  assign n8577 = ~n8511 & n8576;
  assign n8578 = n8511 & ~n8576;
  assign n8579 = ~n8577 & ~n8578;
  assign n8580 = n8510 & ~n8579;
  assign n8581 = ~n8510 & n8579;
  assign n8582 = ~n8580 & ~n8581;
  assign n8583 = ~n8500 & n8582;
  assign n8584 = n8500 & ~n8582;
  assign n8585 = ~n8583 & ~n8584;
  assign n8586 = pi78  & n4843;
  assign n8587 = pi79  & n4598;
  assign n8588 = pi80  & n4593;
  assign n8589 = n1144 & n4591;
  assign n8590 = ~n8587 & ~n8588;
  assign n8591 = ~n8586 & n8590;
  assign n8592 = ~n8589 & n8591;
  assign n8593 = pi38  & n8592;
  assign n8594 = ~pi38  & ~n8592;
  assign n8595 = ~n8593 & ~n8594;
  assign n8596 = n8585 & ~n8595;
  assign n8597 = ~n8585 & n8595;
  assign n8598 = ~n8596 & ~n8597;
  assign n8599 = n8499 & ~n8598;
  assign n8600 = ~n8499 & n8598;
  assign n8601 = ~n8599 & ~n8600;
  assign n8602 = pi81  & n4176;
  assign n8603 = pi82  & n3938;
  assign n8604 = pi83  & n3933;
  assign n8605 = n1577 & n3931;
  assign n8606 = ~n8603 & ~n8604;
  assign n8607 = ~n8602 & n8606;
  assign n8608 = ~n8605 & n8607;
  assign n8609 = pi35  & n8608;
  assign n8610 = ~pi35  & ~n8608;
  assign n8611 = ~n8609 & ~n8610;
  assign n8612 = n8601 & ~n8611;
  assign n8613 = ~n8601 & n8611;
  assign n8614 = ~n8612 & ~n8613;
  assign n8615 = ~n8498 & n8614;
  assign n8616 = n8498 & ~n8614;
  assign n8617 = ~n8615 & ~n8616;
  assign n8618 = pi84  & n3553;
  assign n8619 = pi85  & n3334;
  assign n8620 = pi86  & n3329;
  assign n8621 = n1975 & n3327;
  assign n8622 = ~n8619 & ~n8620;
  assign n8623 = ~n8618 & n8622;
  assign n8624 = ~n8621 & n8623;
  assign n8625 = pi32  & n8624;
  assign n8626 = ~pi32  & ~n8624;
  assign n8627 = ~n8625 & ~n8626;
  assign n8628 = n8617 & ~n8627;
  assign n8629 = ~n8617 & n8627;
  assign n8630 = ~n8628 & ~n8629;
  assign n8631 = n8497 & ~n8630;
  assign n8632 = ~n8497 & n8630;
  assign n8633 = ~n8631 & ~n8632;
  assign n8634 = pi87  & n3011;
  assign n8635 = pi88  & n2809;
  assign n8636 = pi89  & n2804;
  assign n8637 = n2287 & n2802;
  assign n8638 = ~n8635 & ~n8636;
  assign n8639 = ~n8634 & n8638;
  assign n8640 = ~n8637 & n8639;
  assign n8641 = pi29  & n8640;
  assign n8642 = ~pi29  & ~n8640;
  assign n8643 = ~n8641 & ~n8642;
  assign n8644 = n8633 & ~n8643;
  assign n8645 = ~n8633 & n8643;
  assign n8646 = ~n8644 & ~n8645;
  assign n8647 = ~n8496 & n8646;
  assign n8648 = n8496 & ~n8646;
  assign n8649 = ~n8647 & ~n8648;
  assign n8650 = ~n8495 & n8649;
  assign n8651 = n8495 & ~n8649;
  assign n8652 = ~n8650 & ~n8651;
  assign n8653 = n8485 & ~n8652;
  assign n8654 = ~n8485 & n8652;
  assign n8655 = ~n8653 & ~n8654;
  assign n8656 = pi93  & n2053;
  assign n8657 = pi94  & n1893;
  assign n8658 = pi95  & n1888;
  assign n8659 = n1886 & n3475;
  assign n8660 = ~n8657 & ~n8658;
  assign n8661 = ~n8656 & n8660;
  assign n8662 = ~n8659 & n8661;
  assign n8663 = pi23  & n8662;
  assign n8664 = ~pi23  & ~n8662;
  assign n8665 = ~n8663 & ~n8664;
  assign n8666 = n8655 & ~n8665;
  assign n8667 = ~n8655 & n8665;
  assign n8668 = ~n8666 & ~n8667;
  assign n8669 = n8484 & ~n8668;
  assign n8670 = ~n8484 & n8668;
  assign n8671 = ~n8669 & ~n8670;
  assign n8672 = pi96  & n1661;
  assign n8673 = pi97  & n1500;
  assign n8674 = pi98  & n1495;
  assign n8675 = n1493 & n3889;
  assign n8676 = ~n8673 & ~n8674;
  assign n8677 = ~n8672 & n8676;
  assign n8678 = ~n8675 & n8677;
  assign n8679 = pi20  & n8678;
  assign n8680 = ~pi20  & ~n8678;
  assign n8681 = ~n8679 & ~n8680;
  assign n8682 = n8671 & ~n8681;
  assign n8683 = ~n8671 & n8681;
  assign n8684 = ~n8682 & ~n8683;
  assign n8685 = n8483 & ~n8684;
  assign n8686 = ~n8483 & n8684;
  assign n8687 = ~n8685 & ~n8686;
  assign n8688 = pi99  & n1296;
  assign n8689 = pi100  & n1207;
  assign n8690 = pi101  & n1202;
  assign n8691 = n1200 & n4730;
  assign n8692 = ~n8689 & ~n8690;
  assign n8693 = ~n8688 & n8692;
  assign n8694 = ~n8691 & n8693;
  assign n8695 = pi17  & n8694;
  assign n8696 = ~pi17  & ~n8694;
  assign n8697 = ~n8695 & ~n8696;
  assign n8698 = n8687 & ~n8697;
  assign n8699 = ~n8687 & n8697;
  assign n8700 = ~n8698 & ~n8699;
  assign n8701 = n8482 & ~n8700;
  assign n8702 = ~n8482 & n8700;
  assign n8703 = ~n8701 & ~n8702;
  assign n8704 = pi102  & n1006;
  assign n8705 = pi103  & n897;
  assign n8706 = pi104  & n892;
  assign n8707 = n890 & n5212;
  assign n8708 = ~n8705 & ~n8706;
  assign n8709 = ~n8704 & n8708;
  assign n8710 = ~n8707 & n8709;
  assign n8711 = pi14  & n8710;
  assign n8712 = ~pi14  & ~n8710;
  assign n8713 = ~n8711 & ~n8712;
  assign n8714 = n8703 & ~n8713;
  assign n8715 = ~n8703 & n8713;
  assign n8716 = ~n8714 & ~n8715;
  assign n8717 = n8481 & ~n8716;
  assign n8718 = ~n8481 & n8716;
  assign n8719 = ~n8717 & ~n8718;
  assign n8720 = pi105  & n750;
  assign n8721 = pi106  & n651;
  assign n8722 = pi107  & n646;
  assign n8723 = n644 & n6189;
  assign n8724 = ~n8721 & ~n8722;
  assign n8725 = ~n8720 & n8724;
  assign n8726 = ~n8723 & n8725;
  assign n8727 = pi11  & n8726;
  assign n8728 = ~pi11  & ~n8726;
  assign n8729 = ~n8727 & ~n8728;
  assign n8730 = n8719 & ~n8729;
  assign n8731 = ~n8719 & n8729;
  assign n8732 = ~n8730 & ~n8731;
  assign n8733 = ~n8480 & n8732;
  assign n8734 = n8480 & ~n8732;
  assign n8735 = ~n8733 & ~n8734;
  assign n8736 = pi108  & n528;
  assign n8737 = pi109  & n490;
  assign n8738 = pi110  & n485;
  assign n8739 = n483 & n6995;
  assign n8740 = ~n8737 & ~n8738;
  assign n8741 = ~n8736 & n8740;
  assign n8742 = ~n8739 & n8741;
  assign n8743 = pi8  & n8742;
  assign n8744 = ~pi8  & ~n8742;
  assign n8745 = ~n8743 & ~n8744;
  assign n8746 = n8735 & ~n8745;
  assign n8747 = ~n8735 & n8745;
  assign n8748 = ~n8746 & ~n8747;
  assign n8749 = n8479 & ~n8748;
  assign n8750 = ~n8479 & n8748;
  assign n8751 = ~n8749 & ~n8750;
  assign n8752 = pi111  & n391;
  assign n8753 = pi112  & n353;
  assign n8754 = pi113  & n348;
  assign n8755 = n346 & n7852;
  assign n8756 = ~n8753 & ~n8754;
  assign n8757 = ~n8752 & n8756;
  assign n8758 = ~n8755 & n8757;
  assign n8759 = pi5  & n8758;
  assign n8760 = ~pi5  & ~n8758;
  assign n8761 = ~n8759 & ~n8760;
  assign n8762 = n8751 & ~n8761;
  assign n8763 = ~n8751 & n8761;
  assign n8764 = ~n8762 & ~n8763;
  assign n8765 = ~n8478 & n8764;
  assign n8766 = n8478 & ~n8764;
  assign n8767 = ~n8765 & ~n8766;
  assign n8768 = ~n8477 & n8767;
  assign n8769 = n8477 & ~n8767;
  assign n8770 = ~n8768 & ~n8769;
  assign n8771 = ~n8460 & n8770;
  assign n8772 = n8460 & ~n8770;
  assign po52  = ~n8771 & ~n8772;
  assign n8774 = ~n8768 & ~n8771;
  assign n8775 = pi117  & n269;
  assign n8776 = pi116  & n267;
  assign n8777 = pi115  & n282;
  assign n8778 = ~n8466 & ~n8468;
  assign n8779 = ~pi116  & ~pi117 ;
  assign n8780 = pi116  & pi117 ;
  assign n8781 = ~n8779 & ~n8780;
  assign n8782 = ~n8778 & n8781;
  assign n8783 = n8778 & ~n8781;
  assign n8784 = ~n8782 & ~n8783;
  assign n8785 = n262 & n8784;
  assign n8786 = ~n8775 & ~n8776;
  assign n8787 = ~n8777 & n8786;
  assign n8788 = ~n8785 & n8787;
  assign n8789 = pi2  & n8788;
  assign n8790 = ~pi2  & ~n8788;
  assign n8791 = ~n8789 & ~n8790;
  assign n8792 = ~n8762 & ~n8765;
  assign n8793 = ~n8746 & ~n8750;
  assign n8794 = ~n8730 & ~n8733;
  assign n8795 = ~n8714 & ~n8718;
  assign n8796 = ~n8698 & ~n8702;
  assign n8797 = ~n8682 & ~n8686;
  assign n8798 = ~n8666 & ~n8670;
  assign n8799 = pi94  & n2053;
  assign n8800 = pi95  & n1893;
  assign n8801 = pi96  & n1888;
  assign n8802 = n1886 & n3499;
  assign n8803 = ~n8800 & ~n8801;
  assign n8804 = ~n8799 & n8803;
  assign n8805 = ~n8802 & n8804;
  assign n8806 = pi23  & n8805;
  assign n8807 = ~pi23  & ~n8805;
  assign n8808 = ~n8806 & ~n8807;
  assign n8809 = ~n8650 & ~n8654;
  assign n8810 = pi91  & n2510;
  assign n8811 = pi92  & n2342;
  assign n8812 = pi93  & n2337;
  assign n8813 = n2335 & n2948;
  assign n8814 = ~n8811 & ~n8812;
  assign n8815 = ~n8810 & n8814;
  assign n8816 = ~n8813 & n8815;
  assign n8817 = pi26  & n8816;
  assign n8818 = ~pi26  & ~n8816;
  assign n8819 = ~n8817 & ~n8818;
  assign n8820 = ~n8644 & ~n8647;
  assign n8821 = pi88  & n3011;
  assign n8822 = pi89  & n2809;
  assign n8823 = pi90  & n2804;
  assign n8824 = n2448 & n2802;
  assign n8825 = ~n8822 & ~n8823;
  assign n8826 = ~n8821 & n8825;
  assign n8827 = ~n8824 & n8826;
  assign n8828 = pi29  & n8827;
  assign n8829 = ~pi29  & ~n8827;
  assign n8830 = ~n8828 & ~n8829;
  assign n8831 = ~n8628 & ~n8632;
  assign n8832 = pi85  & n3553;
  assign n8833 = pi86  & n3334;
  assign n8834 = pi87  & n3329;
  assign n8835 = n2116 & n3327;
  assign n8836 = ~n8833 & ~n8834;
  assign n8837 = ~n8832 & n8836;
  assign n8838 = ~n8835 & n8837;
  assign n8839 = pi32  & n8838;
  assign n8840 = ~pi32  & ~n8838;
  assign n8841 = ~n8839 & ~n8840;
  assign n8842 = ~n8612 & ~n8615;
  assign n8843 = pi82  & n4176;
  assign n8844 = pi83  & n3938;
  assign n8845 = pi84  & n3933;
  assign n8846 = n1601 & n3931;
  assign n8847 = ~n8844 & ~n8845;
  assign n8848 = ~n8843 & n8847;
  assign n8849 = ~n8846 & n8848;
  assign n8850 = pi35  & n8849;
  assign n8851 = ~pi35  & ~n8849;
  assign n8852 = ~n8850 & ~n8851;
  assign n8853 = ~n8596 & ~n8600;
  assign n8854 = pi79  & n4843;
  assign n8855 = pi80  & n4598;
  assign n8856 = pi81  & n4593;
  assign n8857 = n1337 & n4591;
  assign n8858 = ~n8855 & ~n8856;
  assign n8859 = ~n8854 & n8858;
  assign n8860 = ~n8857 & n8859;
  assign n8861 = pi38  & n8860;
  assign n8862 = ~pi38  & ~n8860;
  assign n8863 = ~n8861 & ~n8862;
  assign n8864 = ~n8581 & ~n8583;
  assign n8865 = ~n8574 & ~n8577;
  assign n8866 = pi73  & n6331;
  assign n8867 = pi74  & n6015;
  assign n8868 = pi75  & n6010;
  assign n8869 = n713 & n6008;
  assign n8870 = ~n8867 & ~n8868;
  assign n8871 = ~n8866 & n8870;
  assign n8872 = ~n8869 & n8871;
  assign n8873 = pi44  & n8872;
  assign n8874 = ~pi44  & ~n8872;
  assign n8875 = ~n8873 & ~n8874;
  assign n8876 = ~n8558 & ~n8562;
  assign n8877 = pi70  & n7121;
  assign n8878 = pi71  & n6795;
  assign n8879 = pi72  & n6790;
  assign n8880 = n551 & n6788;
  assign n8881 = ~n8878 & ~n8879;
  assign n8882 = ~n8877 & n8881;
  assign n8883 = ~n8880 & n8882;
  assign n8884 = pi47  & n8883;
  assign n8885 = ~pi47  & ~n8883;
  assign n8886 = ~n8884 & ~n8885;
  assign n8887 = ~n8543 & ~n8545;
  assign n8888 = pi67  & n7969;
  assign n8889 = pi68  & n7636;
  assign n8890 = pi69  & n7631;
  assign n8891 = n376 & n7629;
  assign n8892 = ~n8889 & ~n8890;
  assign n8893 = ~n8888 & n8892;
  assign n8894 = ~n8891 & n8893;
  assign n8895 = pi50  & n8894;
  assign n8896 = ~pi50  & ~n8894;
  assign n8897 = ~n8895 & ~n8896;
  assign n8898 = pi53  & ~n8265;
  assign n8899 = n8538 & n8898;
  assign n8900 = pi53  & ~n8899;
  assign n8901 = ~n287 & n8528;
  assign n8902 = pi65  & n8535;
  assign n8903 = pi66  & n8530;
  assign n8904 = ~n8264 & n8527;
  assign n8905 = ~n8534 & n8904;
  assign n8906 = pi64  & n8905;
  assign n8907 = ~n8901 & ~n8902;
  assign n8908 = ~n8903 & n8907;
  assign n8909 = ~n8906 & n8908;
  assign n8910 = ~n8900 & n8909;
  assign n8911 = n8900 & ~n8909;
  assign n8912 = ~n8910 & ~n8911;
  assign n8913 = ~n8897 & n8912;
  assign n8914 = n8897 & ~n8912;
  assign n8915 = ~n8913 & ~n8914;
  assign n8916 = ~n8887 & n8915;
  assign n8917 = n8887 & ~n8915;
  assign n8918 = ~n8916 & ~n8917;
  assign n8919 = n8886 & ~n8918;
  assign n8920 = ~n8886 & n8918;
  assign n8921 = ~n8919 & ~n8920;
  assign n8922 = ~n8876 & n8921;
  assign n8923 = n8876 & ~n8921;
  assign n8924 = ~n8922 & ~n8923;
  assign n8925 = n8875 & ~n8924;
  assign n8926 = ~n8875 & n8924;
  assign n8927 = ~n8925 & ~n8926;
  assign n8928 = ~n8865 & n8927;
  assign n8929 = n8865 & ~n8927;
  assign n8930 = ~n8928 & ~n8929;
  assign n8931 = pi76  & n5558;
  assign n8932 = pi77  & n5293;
  assign n8933 = pi78  & n5288;
  assign n8934 = n958 & n5286;
  assign n8935 = ~n8932 & ~n8933;
  assign n8936 = ~n8931 & n8935;
  assign n8937 = ~n8934 & n8936;
  assign n8938 = pi41  & n8937;
  assign n8939 = ~pi41  & ~n8937;
  assign n8940 = ~n8938 & ~n8939;
  assign n8941 = n8930 & ~n8940;
  assign n8942 = ~n8930 & n8940;
  assign n8943 = ~n8941 & ~n8942;
  assign n8944 = ~n8864 & n8943;
  assign n8945 = n8864 & ~n8943;
  assign n8946 = ~n8944 & ~n8945;
  assign n8947 = ~n8863 & n8946;
  assign n8948 = n8863 & ~n8946;
  assign n8949 = ~n8947 & ~n8948;
  assign n8950 = ~n8853 & n8949;
  assign n8951 = n8853 & ~n8949;
  assign n8952 = ~n8950 & ~n8951;
  assign n8953 = ~n8852 & n8952;
  assign n8954 = n8852 & ~n8952;
  assign n8955 = ~n8953 & ~n8954;
  assign n8956 = ~n8842 & n8955;
  assign n8957 = n8842 & ~n8955;
  assign n8958 = ~n8956 & ~n8957;
  assign n8959 = ~n8841 & n8958;
  assign n8960 = n8841 & ~n8958;
  assign n8961 = ~n8959 & ~n8960;
  assign n8962 = ~n8831 & n8961;
  assign n8963 = n8831 & ~n8961;
  assign n8964 = ~n8962 & ~n8963;
  assign n8965 = n8830 & ~n8964;
  assign n8966 = ~n8830 & n8964;
  assign n8967 = ~n8965 & ~n8966;
  assign n8968 = ~n8820 & n8967;
  assign n8969 = n8820 & ~n8967;
  assign n8970 = ~n8968 & ~n8969;
  assign n8971 = n8819 & ~n8970;
  assign n8972 = ~n8819 & n8970;
  assign n8973 = ~n8971 & ~n8972;
  assign n8974 = ~n8809 & n8973;
  assign n8975 = n8809 & ~n8973;
  assign n8976 = ~n8974 & ~n8975;
  assign n8977 = n8808 & ~n8976;
  assign n8978 = ~n8808 & n8976;
  assign n8979 = ~n8977 & ~n8978;
  assign n8980 = ~n8798 & n8979;
  assign n8981 = n8798 & ~n8979;
  assign n8982 = ~n8980 & ~n8981;
  assign n8983 = pi97  & n1661;
  assign n8984 = pi98  & n1500;
  assign n8985 = pi99  & n1495;
  assign n8986 = n1493 & n4101;
  assign n8987 = ~n8984 & ~n8985;
  assign n8988 = ~n8983 & n8987;
  assign n8989 = ~n8986 & n8988;
  assign n8990 = pi20  & n8989;
  assign n8991 = ~pi20  & ~n8989;
  assign n8992 = ~n8990 & ~n8991;
  assign n8993 = n8982 & ~n8992;
  assign n8994 = ~n8982 & n8992;
  assign n8995 = ~n8993 & ~n8994;
  assign n8996 = n8797 & ~n8995;
  assign n8997 = ~n8797 & n8995;
  assign n8998 = ~n8996 & ~n8997;
  assign n8999 = pi100  & n1296;
  assign n9000 = pi101  & n1207;
  assign n9001 = pi102  & n1202;
  assign n9002 = n1200 & n4956;
  assign n9003 = ~n9000 & ~n9001;
  assign n9004 = ~n8999 & n9003;
  assign n9005 = ~n9002 & n9004;
  assign n9006 = pi17  & n9005;
  assign n9007 = ~pi17  & ~n9005;
  assign n9008 = ~n9006 & ~n9007;
  assign n9009 = n8998 & ~n9008;
  assign n9010 = ~n8998 & n9008;
  assign n9011 = ~n9009 & ~n9010;
  assign n9012 = n8796 & ~n9011;
  assign n9013 = ~n8796 & n9011;
  assign n9014 = ~n9012 & ~n9013;
  assign n9015 = pi103  & n1006;
  assign n9016 = pi104  & n897;
  assign n9017 = pi105  & n892;
  assign n9018 = n890 & n5677;
  assign n9019 = ~n9016 & ~n9017;
  assign n9020 = ~n9015 & n9019;
  assign n9021 = ~n9018 & n9020;
  assign n9022 = pi14  & n9021;
  assign n9023 = ~pi14  & ~n9021;
  assign n9024 = ~n9022 & ~n9023;
  assign n9025 = n9014 & ~n9024;
  assign n9026 = ~n9014 & n9024;
  assign n9027 = ~n9025 & ~n9026;
  assign n9028 = n8795 & ~n9027;
  assign n9029 = ~n8795 & n9027;
  assign n9030 = ~n9028 & ~n9029;
  assign n9031 = pi106  & n750;
  assign n9032 = pi107  & n651;
  assign n9033 = pi108  & n646;
  assign n9034 = n644 & n6213;
  assign n9035 = ~n9032 & ~n9033;
  assign n9036 = ~n9031 & n9035;
  assign n9037 = ~n9034 & n9036;
  assign n9038 = pi11  & n9037;
  assign n9039 = ~pi11  & ~n9037;
  assign n9040 = ~n9038 & ~n9039;
  assign n9041 = n9030 & ~n9040;
  assign n9042 = ~n9030 & n9040;
  assign n9043 = ~n9041 & ~n9042;
  assign n9044 = ~n8794 & n9043;
  assign n9045 = n8794 & ~n9043;
  assign n9046 = ~n9044 & ~n9045;
  assign n9047 = pi109  & n528;
  assign n9048 = pi110  & n490;
  assign n9049 = pi111  & n485;
  assign n9050 = n483 & n7272;
  assign n9051 = ~n9048 & ~n9049;
  assign n9052 = ~n9047 & n9051;
  assign n9053 = ~n9050 & n9052;
  assign n9054 = pi8  & n9053;
  assign n9055 = ~pi8  & ~n9053;
  assign n9056 = ~n9054 & ~n9055;
  assign n9057 = n9046 & ~n9056;
  assign n9058 = ~n9046 & n9056;
  assign n9059 = ~n9057 & ~n9058;
  assign n9060 = n8793 & ~n9059;
  assign n9061 = ~n8793 & n9059;
  assign n9062 = ~n9060 & ~n9061;
  assign n9063 = pi112  & n391;
  assign n9064 = pi113  & n353;
  assign n9065 = pi114  & n348;
  assign n9066 = n346 & n8146;
  assign n9067 = ~n9064 & ~n9065;
  assign n9068 = ~n9063 & n9067;
  assign n9069 = ~n9066 & n9068;
  assign n9070 = pi5  & n9069;
  assign n9071 = ~pi5  & ~n9069;
  assign n9072 = ~n9070 & ~n9071;
  assign n9073 = n9062 & ~n9072;
  assign n9074 = ~n9062 & n9072;
  assign n9075 = ~n9073 & ~n9074;
  assign n9076 = ~n8792 & n9075;
  assign n9077 = n8792 & ~n9075;
  assign n9078 = ~n9076 & ~n9077;
  assign n9079 = ~n8791 & n9078;
  assign n9080 = n8791 & ~n9078;
  assign n9081 = ~n9079 & ~n9080;
  assign n9082 = ~n8774 & n9081;
  assign n9083 = n8774 & ~n9081;
  assign po53  = ~n9082 & ~n9083;
  assign n9085 = ~n9079 & ~n9082;
  assign n9086 = pi118  & n269;
  assign n9087 = pi117  & n267;
  assign n9088 = pi116  & n282;
  assign n9089 = ~n8780 & ~n8782;
  assign n9090 = ~pi117  & ~pi118 ;
  assign n9091 = pi117  & pi118 ;
  assign n9092 = ~n9090 & ~n9091;
  assign n9093 = ~n9089 & n9092;
  assign n9094 = n9089 & ~n9092;
  assign n9095 = ~n9093 & ~n9094;
  assign n9096 = n262 & n9095;
  assign n9097 = ~n9086 & ~n9087;
  assign n9098 = ~n9088 & n9097;
  assign n9099 = ~n9096 & n9098;
  assign n9100 = pi2  & n9099;
  assign n9101 = ~pi2  & ~n9099;
  assign n9102 = ~n9100 & ~n9101;
  assign n9103 = ~n9073 & ~n9076;
  assign n9104 = ~n9057 & ~n9061;
  assign n9105 = pi110  & n528;
  assign n9106 = pi111  & n490;
  assign n9107 = pi112  & n485;
  assign n9108 = n483 & n7296;
  assign n9109 = ~n9106 & ~n9107;
  assign n9110 = ~n9105 & n9109;
  assign n9111 = ~n9108 & n9110;
  assign n9112 = pi8  & n9111;
  assign n9113 = ~pi8  & ~n9111;
  assign n9114 = ~n9112 & ~n9113;
  assign n9115 = ~n9041 & ~n9044;
  assign n9116 = pi107  & n750;
  assign n9117 = pi108  & n651;
  assign n9118 = pi109  & n646;
  assign n9119 = n644 & n6715;
  assign n9120 = ~n9117 & ~n9118;
  assign n9121 = ~n9116 & n9120;
  assign n9122 = ~n9119 & n9121;
  assign n9123 = pi11  & n9122;
  assign n9124 = ~pi11  & ~n9122;
  assign n9125 = ~n9123 & ~n9124;
  assign n9126 = ~n9025 & ~n9029;
  assign n9127 = ~n9009 & ~n9013;
  assign n9128 = ~n8993 & ~n8997;
  assign n9129 = pi98  & n1661;
  assign n9130 = pi99  & n1500;
  assign n9131 = pi100  & n1495;
  assign n9132 = n1493 & n4501;
  assign n9133 = ~n9130 & ~n9131;
  assign n9134 = ~n9129 & n9133;
  assign n9135 = ~n9132 & n9134;
  assign n9136 = pi20  & n9135;
  assign n9137 = ~pi20  & ~n9135;
  assign n9138 = ~n9136 & ~n9137;
  assign n9139 = ~n8978 & ~n8980;
  assign n9140 = ~n8972 & ~n8974;
  assign n9141 = pi92  & n2510;
  assign n9142 = pi93  & n2342;
  assign n9143 = pi94  & n2337;
  assign n9144 = n2335 & n3280;
  assign n9145 = ~n9142 & ~n9143;
  assign n9146 = ~n9141 & n9145;
  assign n9147 = ~n9144 & n9146;
  assign n9148 = pi26  & n9147;
  assign n9149 = ~pi26  & ~n9147;
  assign n9150 = ~n9148 & ~n9149;
  assign n9151 = ~n8966 & ~n8968;
  assign n9152 = pi89  & n3011;
  assign n9153 = pi90  & n2809;
  assign n9154 = pi91  & n2804;
  assign n9155 = n2746 & n2802;
  assign n9156 = ~n9153 & ~n9154;
  assign n9157 = ~n9152 & n9156;
  assign n9158 = ~n9155 & n9157;
  assign n9159 = pi29  & n9158;
  assign n9160 = ~pi29  & ~n9158;
  assign n9161 = ~n9159 & ~n9160;
  assign n9162 = ~n8959 & ~n8962;
  assign n9163 = pi86  & n3553;
  assign n9164 = pi87  & n3334;
  assign n9165 = pi88  & n3329;
  assign n9166 = n2140 & n3327;
  assign n9167 = ~n9164 & ~n9165;
  assign n9168 = ~n9163 & n9167;
  assign n9169 = ~n9166 & n9168;
  assign n9170 = pi32  & n9169;
  assign n9171 = ~pi32  & ~n9169;
  assign n9172 = ~n9170 & ~n9171;
  assign n9173 = ~n8953 & ~n8956;
  assign n9174 = pi83  & n4176;
  assign n9175 = pi84  & n3938;
  assign n9176 = pi85  & n3933;
  assign n9177 = n1831 & n3931;
  assign n9178 = ~n9175 & ~n9176;
  assign n9179 = ~n9174 & n9178;
  assign n9180 = ~n9177 & n9179;
  assign n9181 = pi35  & n9180;
  assign n9182 = ~pi35  & ~n9180;
  assign n9183 = ~n9181 & ~n9182;
  assign n9184 = ~n8947 & ~n8950;
  assign n9185 = pi80  & n4843;
  assign n9186 = pi81  & n4598;
  assign n9187 = pi82  & n4593;
  assign n9188 = n1450 & n4591;
  assign n9189 = ~n9186 & ~n9187;
  assign n9190 = ~n9185 & n9189;
  assign n9191 = ~n9188 & n9190;
  assign n9192 = pi38  & n9191;
  assign n9193 = ~pi38  & ~n9191;
  assign n9194 = ~n9192 & ~n9193;
  assign n9195 = ~n8941 & ~n8944;
  assign n9196 = pi77  & n5558;
  assign n9197 = pi78  & n5293;
  assign n9198 = pi79  & n5288;
  assign n9199 = n1048 & n5286;
  assign n9200 = ~n9197 & ~n9198;
  assign n9201 = ~n9196 & n9200;
  assign n9202 = ~n9199 & n9201;
  assign n9203 = pi41  & n9202;
  assign n9204 = ~pi41  & ~n9202;
  assign n9205 = ~n9203 & ~n9204;
  assign n9206 = ~n8926 & ~n8928;
  assign n9207 = pi74  & n6331;
  assign n9208 = pi75  & n6015;
  assign n9209 = pi76  & n6010;
  assign n9210 = n841 & n6008;
  assign n9211 = ~n9208 & ~n9209;
  assign n9212 = ~n9207 & n9211;
  assign n9213 = ~n9210 & n9212;
  assign n9214 = pi44  & n9213;
  assign n9215 = ~pi44  & ~n9213;
  assign n9216 = ~n9214 & ~n9215;
  assign n9217 = ~n8920 & ~n8922;
  assign n9218 = pi71  & n7121;
  assign n9219 = pi72  & n6795;
  assign n9220 = pi73  & n6790;
  assign n9221 = n613 & n6788;
  assign n9222 = ~n9219 & ~n9220;
  assign n9223 = ~n9218 & n9222;
  assign n9224 = ~n9221 & n9223;
  assign n9225 = pi47  & n9224;
  assign n9226 = ~pi47  & ~n9224;
  assign n9227 = ~n9225 & ~n9226;
  assign n9228 = ~n8913 & ~n8916;
  assign n9229 = pi65  & n8905;
  assign n9230 = pi66  & n8535;
  assign n9231 = pi67  & n8530;
  assign n9232 = n305 & n8528;
  assign n9233 = ~n9230 & ~n9231;
  assign n9234 = ~n9229 & n9233;
  assign n9235 = ~n9232 & n9234;
  assign n9236 = pi53  & n9235;
  assign n9237 = ~pi53  & ~n9235;
  assign n9238 = ~n9236 & ~n9237;
  assign n9239 = ~pi53  & ~pi54 ;
  assign n9240 = pi53  & pi54 ;
  assign n9241 = ~n9239 & ~n9240;
  assign n9242 = pi64  & n9241;
  assign n9243 = n8899 & n8909;
  assign n9244 = n9242 & n9243;
  assign n9245 = ~n9242 & ~n9243;
  assign n9246 = ~n9244 & ~n9245;
  assign n9247 = ~n9238 & n9246;
  assign n9248 = n9238 & ~n9246;
  assign n9249 = ~n9247 & ~n9248;
  assign n9250 = pi68  & n7969;
  assign n9251 = pi69  & n7636;
  assign n9252 = pi70  & n7631;
  assign n9253 = n415 & n7629;
  assign n9254 = ~n9251 & ~n9252;
  assign n9255 = ~n9250 & n9254;
  assign n9256 = ~n9253 & n9255;
  assign n9257 = pi50  & n9256;
  assign n9258 = ~pi50  & ~n9256;
  assign n9259 = ~n9257 & ~n9258;
  assign n9260 = n9249 & ~n9259;
  assign n9261 = ~n9249 & n9259;
  assign n9262 = ~n9260 & ~n9261;
  assign n9263 = ~n9228 & n9262;
  assign n9264 = n9228 & ~n9262;
  assign n9265 = ~n9263 & ~n9264;
  assign n9266 = ~n9227 & n9265;
  assign n9267 = n9227 & ~n9265;
  assign n9268 = ~n9266 & ~n9267;
  assign n9269 = ~n9217 & n9268;
  assign n9270 = n9217 & ~n9268;
  assign n9271 = ~n9269 & ~n9270;
  assign n9272 = ~n9216 & n9271;
  assign n9273 = n9216 & ~n9271;
  assign n9274 = ~n9272 & ~n9273;
  assign n9275 = ~n9206 & n9274;
  assign n9276 = n9206 & ~n9274;
  assign n9277 = ~n9275 & ~n9276;
  assign n9278 = ~n9205 & n9277;
  assign n9279 = n9205 & ~n9277;
  assign n9280 = ~n9278 & ~n9279;
  assign n9281 = ~n9195 & n9280;
  assign n9282 = n9195 & ~n9280;
  assign n9283 = ~n9281 & ~n9282;
  assign n9284 = ~n9194 & n9283;
  assign n9285 = n9194 & ~n9283;
  assign n9286 = ~n9284 & ~n9285;
  assign n9287 = ~n9184 & n9286;
  assign n9288 = n9184 & ~n9286;
  assign n9289 = ~n9287 & ~n9288;
  assign n9290 = ~n9183 & n9289;
  assign n9291 = n9183 & ~n9289;
  assign n9292 = ~n9290 & ~n9291;
  assign n9293 = ~n9173 & n9292;
  assign n9294 = n9173 & ~n9292;
  assign n9295 = ~n9293 & ~n9294;
  assign n9296 = ~n9172 & n9295;
  assign n9297 = n9172 & ~n9295;
  assign n9298 = ~n9296 & ~n9297;
  assign n9299 = ~n9162 & n9298;
  assign n9300 = n9162 & ~n9298;
  assign n9301 = ~n9299 & ~n9300;
  assign n9302 = ~n9161 & n9301;
  assign n9303 = n9161 & ~n9301;
  assign n9304 = ~n9302 & ~n9303;
  assign n9305 = ~n9151 & n9304;
  assign n9306 = n9151 & ~n9304;
  assign n9307 = ~n9305 & ~n9306;
  assign n9308 = ~n9150 & n9307;
  assign n9309 = n9150 & ~n9307;
  assign n9310 = ~n9308 & ~n9309;
  assign n9311 = ~n9140 & n9310;
  assign n9312 = n9140 & ~n9310;
  assign n9313 = ~n9311 & ~n9312;
  assign n9314 = pi95  & n2053;
  assign n9315 = pi96  & n1893;
  assign n9316 = pi97  & n1888;
  assign n9317 = n1886 & n3691;
  assign n9318 = ~n9315 & ~n9316;
  assign n9319 = ~n9314 & n9318;
  assign n9320 = ~n9317 & n9319;
  assign n9321 = pi23  & n9320;
  assign n9322 = ~pi23  & ~n9320;
  assign n9323 = ~n9321 & ~n9322;
  assign n9324 = n9313 & ~n9323;
  assign n9325 = ~n9313 & n9323;
  assign n9326 = ~n9324 & ~n9325;
  assign n9327 = ~n9139 & n9326;
  assign n9328 = n9139 & ~n9326;
  assign n9329 = ~n9327 & ~n9328;
  assign n9330 = ~n9138 & n9329;
  assign n9331 = n9138 & ~n9329;
  assign n9332 = ~n9330 & ~n9331;
  assign n9333 = n9128 & ~n9332;
  assign n9334 = ~n9128 & n9332;
  assign n9335 = ~n9333 & ~n9334;
  assign n9336 = pi101  & n1296;
  assign n9337 = pi102  & n1207;
  assign n9338 = pi103  & n1202;
  assign n9339 = n1200 & n5188;
  assign n9340 = ~n9337 & ~n9338;
  assign n9341 = ~n9336 & n9340;
  assign n9342 = ~n9339 & n9341;
  assign n9343 = pi17  & n9342;
  assign n9344 = ~pi17  & ~n9342;
  assign n9345 = ~n9343 & ~n9344;
  assign n9346 = n9335 & ~n9345;
  assign n9347 = ~n9335 & n9345;
  assign n9348 = ~n9346 & ~n9347;
  assign n9349 = n9127 & ~n9348;
  assign n9350 = ~n9127 & n9348;
  assign n9351 = ~n9349 & ~n9350;
  assign n9352 = pi104  & n1006;
  assign n9353 = pi105  & n897;
  assign n9354 = pi106  & n892;
  assign n9355 = n890 & n5701;
  assign n9356 = ~n9353 & ~n9354;
  assign n9357 = ~n9352 & n9356;
  assign n9358 = ~n9355 & n9357;
  assign n9359 = pi14  & n9358;
  assign n9360 = ~pi14  & ~n9358;
  assign n9361 = ~n9359 & ~n9360;
  assign n9362 = ~n9351 & n9361;
  assign n9363 = n9351 & ~n9361;
  assign n9364 = ~n9362 & ~n9363;
  assign n9365 = ~n9126 & n9364;
  assign n9366 = n9126 & ~n9364;
  assign n9367 = ~n9365 & ~n9366;
  assign n9368 = ~n9125 & n9367;
  assign n9369 = n9125 & ~n9367;
  assign n9370 = ~n9368 & ~n9369;
  assign n9371 = ~n9115 & n9370;
  assign n9372 = n9115 & ~n9370;
  assign n9373 = ~n9371 & ~n9372;
  assign n9374 = ~n9114 & n9373;
  assign n9375 = n9114 & ~n9373;
  assign n9376 = ~n9374 & ~n9375;
  assign n9377 = n9104 & ~n9376;
  assign n9378 = ~n9104 & n9376;
  assign n9379 = ~n9377 & ~n9378;
  assign n9380 = pi113  & n391;
  assign n9381 = pi114  & n353;
  assign n9382 = pi115  & n348;
  assign n9383 = n346 & n8170;
  assign n9384 = ~n9381 & ~n9382;
  assign n9385 = ~n9380 & n9384;
  assign n9386 = ~n9383 & n9385;
  assign n9387 = pi5  & n9386;
  assign n9388 = ~pi5  & ~n9386;
  assign n9389 = ~n9387 & ~n9388;
  assign n9390 = ~n9379 & n9389;
  assign n9391 = n9379 & ~n9389;
  assign n9392 = ~n9390 & ~n9391;
  assign n9393 = ~n9103 & n9392;
  assign n9394 = n9103 & ~n9392;
  assign n9395 = ~n9393 & ~n9394;
  assign n9396 = ~n9102 & n9395;
  assign n9397 = n9102 & ~n9395;
  assign n9398 = ~n9396 & ~n9397;
  assign n9399 = ~n9085 & n9398;
  assign n9400 = n9085 & ~n9398;
  assign po54  = ~n9399 & ~n9400;
  assign n9402 = ~n9396 & ~n9399;
  assign n9403 = pi119  & n269;
  assign n9404 = pi118  & n267;
  assign n9405 = pi117  & n282;
  assign n9406 = ~n9091 & ~n9093;
  assign n9407 = ~pi118  & ~pi119 ;
  assign n9408 = pi118  & pi119 ;
  assign n9409 = ~n9407 & ~n9408;
  assign n9410 = ~n9406 & n9409;
  assign n9411 = n9406 & ~n9409;
  assign n9412 = ~n9410 & ~n9411;
  assign n9413 = n262 & n9412;
  assign n9414 = ~n9403 & ~n9404;
  assign n9415 = ~n9405 & n9414;
  assign n9416 = ~n9413 & n9415;
  assign n9417 = pi2  & n9416;
  assign n9418 = ~pi2  & ~n9416;
  assign n9419 = ~n9417 & ~n9418;
  assign n9420 = ~n9391 & ~n9393;
  assign n9421 = ~n9374 & ~n9378;
  assign n9422 = pi111  & n528;
  assign n9423 = pi112  & n490;
  assign n9424 = pi113  & n485;
  assign n9425 = n483 & n7852;
  assign n9426 = ~n9423 & ~n9424;
  assign n9427 = ~n9422 & n9426;
  assign n9428 = ~n9425 & n9427;
  assign n9429 = pi8  & n9428;
  assign n9430 = ~pi8  & ~n9428;
  assign n9431 = ~n9429 & ~n9430;
  assign n9432 = ~n9368 & ~n9371;
  assign n9433 = pi108  & n750;
  assign n9434 = pi109  & n651;
  assign n9435 = pi110  & n646;
  assign n9436 = n644 & n6995;
  assign n9437 = ~n9434 & ~n9435;
  assign n9438 = ~n9433 & n9437;
  assign n9439 = ~n9436 & n9438;
  assign n9440 = pi11  & n9439;
  assign n9441 = ~pi11  & ~n9439;
  assign n9442 = ~n9440 & ~n9441;
  assign n9443 = ~n9363 & ~n9365;
  assign n9444 = ~n9346 & ~n9350;
  assign n9445 = ~n9330 & ~n9334;
  assign n9446 = ~n9324 & ~n9327;
  assign n9447 = ~n9308 & ~n9311;
  assign n9448 = ~n9302 & ~n9305;
  assign n9449 = ~n9296 & ~n9299;
  assign n9450 = ~n9290 & ~n9293;
  assign n9451 = ~n9284 & ~n9287;
  assign n9452 = ~n9278 & ~n9281;
  assign n9453 = ~n9272 & ~n9275;
  assign n9454 = pi75  & n6331;
  assign n9455 = pi76  & n6015;
  assign n9456 = pi77  & n6010;
  assign n9457 = n865 & n6008;
  assign n9458 = ~n9455 & ~n9456;
  assign n9459 = ~n9454 & n9458;
  assign n9460 = ~n9457 & n9459;
  assign n9461 = pi44  & n9460;
  assign n9462 = ~pi44  & ~n9460;
  assign n9463 = ~n9461 & ~n9462;
  assign n9464 = ~n9266 & ~n9269;
  assign n9465 = pi72  & n7121;
  assign n9466 = pi73  & n6795;
  assign n9467 = pi74  & n6790;
  assign n9468 = n689 & n6788;
  assign n9469 = ~n9466 & ~n9467;
  assign n9470 = ~n9465 & n9469;
  assign n9471 = ~n9468 & n9470;
  assign n9472 = pi47  & n9471;
  assign n9473 = ~pi47  & ~n9471;
  assign n9474 = ~n9472 & ~n9473;
  assign n9475 = ~n9260 & ~n9263;
  assign n9476 = pi69  & n7969;
  assign n9477 = pi70  & n7636;
  assign n9478 = pi71  & n7631;
  assign n9479 = n460 & n7629;
  assign n9480 = ~n9477 & ~n9478;
  assign n9481 = ~n9476 & n9480;
  assign n9482 = ~n9479 & n9481;
  assign n9483 = pi50  & n9482;
  assign n9484 = ~pi50  & ~n9482;
  assign n9485 = ~n9483 & ~n9484;
  assign n9486 = ~n9244 & ~n9247;
  assign n9487 = pi66  & n8905;
  assign n9488 = pi67  & n8535;
  assign n9489 = pi68  & n8530;
  assign n9490 = n334 & n8528;
  assign n9491 = ~n9488 & ~n9489;
  assign n9492 = ~n9487 & n9491;
  assign n9493 = ~n9490 & n9492;
  assign n9494 = pi53  & n9493;
  assign n9495 = ~pi53  & ~n9493;
  assign n9496 = ~n9494 & ~n9495;
  assign n9497 = pi56  & n9242;
  assign n9498 = ~pi55  & ~pi56 ;
  assign n9499 = pi55  & pi56 ;
  assign n9500 = ~n9498 & ~n9499;
  assign n9501 = n9241 & n9500;
  assign n9502 = n265 & n9501;
  assign n9503 = n9241 & ~n9500;
  assign n9504 = pi65  & n9503;
  assign n9505 = ~pi54  & ~pi55 ;
  assign n9506 = pi54  & pi55 ;
  assign n9507 = ~n9505 & ~n9506;
  assign n9508 = ~n9241 & n9507;
  assign n9509 = pi64  & n9508;
  assign n9510 = ~n9502 & ~n9504;
  assign n9511 = ~n9509 & n9510;
  assign n9512 = n9497 & ~n9511;
  assign n9513 = ~n9497 & n9511;
  assign n9514 = ~n9512 & ~n9513;
  assign n9515 = n9496 & ~n9514;
  assign n9516 = ~n9496 & n9514;
  assign n9517 = ~n9515 & ~n9516;
  assign n9518 = ~n9486 & n9517;
  assign n9519 = n9486 & ~n9517;
  assign n9520 = ~n9518 & ~n9519;
  assign n9521 = n9485 & ~n9520;
  assign n9522 = ~n9485 & n9520;
  assign n9523 = ~n9521 & ~n9522;
  assign n9524 = ~n9475 & n9523;
  assign n9525 = n9475 & ~n9523;
  assign n9526 = ~n9524 & ~n9525;
  assign n9527 = n9474 & ~n9526;
  assign n9528 = ~n9474 & n9526;
  assign n9529 = ~n9527 & ~n9528;
  assign n9530 = ~n9464 & n9529;
  assign n9531 = n9464 & ~n9529;
  assign n9532 = ~n9530 & ~n9531;
  assign n9533 = n9463 & ~n9532;
  assign n9534 = ~n9463 & n9532;
  assign n9535 = ~n9533 & ~n9534;
  assign n9536 = ~n9453 & n9535;
  assign n9537 = n9453 & ~n9535;
  assign n9538 = ~n9536 & ~n9537;
  assign n9539 = pi78  & n5558;
  assign n9540 = pi79  & n5293;
  assign n9541 = pi80  & n5288;
  assign n9542 = n1144 & n5286;
  assign n9543 = ~n9540 & ~n9541;
  assign n9544 = ~n9539 & n9543;
  assign n9545 = ~n9542 & n9544;
  assign n9546 = pi41  & n9545;
  assign n9547 = ~pi41  & ~n9545;
  assign n9548 = ~n9546 & ~n9547;
  assign n9549 = n9538 & ~n9548;
  assign n9550 = ~n9538 & n9548;
  assign n9551 = ~n9549 & ~n9550;
  assign n9552 = n9452 & ~n9551;
  assign n9553 = ~n9452 & n9551;
  assign n9554 = ~n9552 & ~n9553;
  assign n9555 = pi81  & n4843;
  assign n9556 = pi82  & n4598;
  assign n9557 = pi83  & n4593;
  assign n9558 = n1577 & n4591;
  assign n9559 = ~n9556 & ~n9557;
  assign n9560 = ~n9555 & n9559;
  assign n9561 = ~n9558 & n9560;
  assign n9562 = pi38  & n9561;
  assign n9563 = ~pi38  & ~n9561;
  assign n9564 = ~n9562 & ~n9563;
  assign n9565 = n9554 & ~n9564;
  assign n9566 = ~n9554 & n9564;
  assign n9567 = ~n9565 & ~n9566;
  assign n9568 = ~n9451 & n9567;
  assign n9569 = n9451 & ~n9567;
  assign n9570 = ~n9568 & ~n9569;
  assign n9571 = pi84  & n4176;
  assign n9572 = pi85  & n3938;
  assign n9573 = pi86  & n3933;
  assign n9574 = n1975 & n3931;
  assign n9575 = ~n9572 & ~n9573;
  assign n9576 = ~n9571 & n9575;
  assign n9577 = ~n9574 & n9576;
  assign n9578 = pi35  & n9577;
  assign n9579 = ~pi35  & ~n9577;
  assign n9580 = ~n9578 & ~n9579;
  assign n9581 = n9570 & ~n9580;
  assign n9582 = ~n9570 & n9580;
  assign n9583 = ~n9581 & ~n9582;
  assign n9584 = n9450 & ~n9583;
  assign n9585 = ~n9450 & n9583;
  assign n9586 = ~n9584 & ~n9585;
  assign n9587 = pi87  & n3553;
  assign n9588 = pi88  & n3334;
  assign n9589 = pi89  & n3329;
  assign n9590 = n2287 & n3327;
  assign n9591 = ~n9588 & ~n9589;
  assign n9592 = ~n9587 & n9591;
  assign n9593 = ~n9590 & n9592;
  assign n9594 = pi32  & n9593;
  assign n9595 = ~pi32  & ~n9593;
  assign n9596 = ~n9594 & ~n9595;
  assign n9597 = n9586 & ~n9596;
  assign n9598 = ~n9586 & n9596;
  assign n9599 = ~n9597 & ~n9598;
  assign n9600 = n9449 & ~n9599;
  assign n9601 = ~n9449 & n9599;
  assign n9602 = ~n9600 & ~n9601;
  assign n9603 = pi90  & n3011;
  assign n9604 = pi91  & n2809;
  assign n9605 = pi92  & n2804;
  assign n9606 = n2802 & n2924;
  assign n9607 = ~n9604 & ~n9605;
  assign n9608 = ~n9603 & n9607;
  assign n9609 = ~n9606 & n9608;
  assign n9610 = pi29  & n9609;
  assign n9611 = ~pi29  & ~n9609;
  assign n9612 = ~n9610 & ~n9611;
  assign n9613 = n9602 & ~n9612;
  assign n9614 = ~n9602 & n9612;
  assign n9615 = ~n9613 & ~n9614;
  assign n9616 = n9448 & ~n9615;
  assign n9617 = ~n9448 & n9615;
  assign n9618 = ~n9616 & ~n9617;
  assign n9619 = pi93  & n2510;
  assign n9620 = pi94  & n2342;
  assign n9621 = pi95  & n2337;
  assign n9622 = n2335 & n3475;
  assign n9623 = ~n9620 & ~n9621;
  assign n9624 = ~n9619 & n9623;
  assign n9625 = ~n9622 & n9624;
  assign n9626 = pi26  & n9625;
  assign n9627 = ~pi26  & ~n9625;
  assign n9628 = ~n9626 & ~n9627;
  assign n9629 = n9618 & ~n9628;
  assign n9630 = ~n9618 & n9628;
  assign n9631 = ~n9629 & ~n9630;
  assign n9632 = n9447 & ~n9631;
  assign n9633 = ~n9447 & n9631;
  assign n9634 = ~n9632 & ~n9633;
  assign n9635 = pi96  & n2053;
  assign n9636 = pi97  & n1893;
  assign n9637 = pi98  & n1888;
  assign n9638 = n1886 & n3889;
  assign n9639 = ~n9636 & ~n9637;
  assign n9640 = ~n9635 & n9639;
  assign n9641 = ~n9638 & n9640;
  assign n9642 = pi23  & n9641;
  assign n9643 = ~pi23  & ~n9641;
  assign n9644 = ~n9642 & ~n9643;
  assign n9645 = n9634 & ~n9644;
  assign n9646 = ~n9634 & n9644;
  assign n9647 = ~n9645 & ~n9646;
  assign n9648 = n9446 & ~n9647;
  assign n9649 = ~n9446 & n9647;
  assign n9650 = ~n9648 & ~n9649;
  assign n9651 = pi99  & n1661;
  assign n9652 = pi100  & n1500;
  assign n9653 = pi101  & n1495;
  assign n9654 = n1493 & n4730;
  assign n9655 = ~n9652 & ~n9653;
  assign n9656 = ~n9651 & n9655;
  assign n9657 = ~n9654 & n9656;
  assign n9658 = pi20  & n9657;
  assign n9659 = ~pi20  & ~n9657;
  assign n9660 = ~n9658 & ~n9659;
  assign n9661 = n9650 & ~n9660;
  assign n9662 = ~n9650 & n9660;
  assign n9663 = ~n9661 & ~n9662;
  assign n9664 = n9445 & ~n9663;
  assign n9665 = ~n9445 & n9663;
  assign n9666 = ~n9664 & ~n9665;
  assign n9667 = pi102  & n1296;
  assign n9668 = pi103  & n1207;
  assign n9669 = pi104  & n1202;
  assign n9670 = n1200 & n5212;
  assign n9671 = ~n9668 & ~n9669;
  assign n9672 = ~n9667 & n9671;
  assign n9673 = ~n9670 & n9672;
  assign n9674 = pi17  & n9673;
  assign n9675 = ~pi17  & ~n9673;
  assign n9676 = ~n9674 & ~n9675;
  assign n9677 = n9666 & ~n9676;
  assign n9678 = ~n9666 & n9676;
  assign n9679 = ~n9677 & ~n9678;
  assign n9680 = n9444 & ~n9679;
  assign n9681 = ~n9444 & n9679;
  assign n9682 = ~n9680 & ~n9681;
  assign n9683 = pi105  & n1006;
  assign n9684 = pi106  & n897;
  assign n9685 = pi107  & n892;
  assign n9686 = n890 & n6189;
  assign n9687 = ~n9684 & ~n9685;
  assign n9688 = ~n9683 & n9687;
  assign n9689 = ~n9686 & n9688;
  assign n9690 = pi14  & n9689;
  assign n9691 = ~pi14  & ~n9689;
  assign n9692 = ~n9690 & ~n9691;
  assign n9693 = n9682 & ~n9692;
  assign n9694 = ~n9682 & n9692;
  assign n9695 = ~n9693 & ~n9694;
  assign n9696 = ~n9443 & n9695;
  assign n9697 = n9443 & ~n9695;
  assign n9698 = ~n9696 & ~n9697;
  assign n9699 = n9442 & ~n9698;
  assign n9700 = ~n9442 & n9698;
  assign n9701 = ~n9699 & ~n9700;
  assign n9702 = ~n9432 & n9701;
  assign n9703 = n9432 & ~n9701;
  assign n9704 = ~n9702 & ~n9703;
  assign n9705 = n9431 & ~n9704;
  assign n9706 = ~n9431 & n9704;
  assign n9707 = ~n9705 & ~n9706;
  assign n9708 = ~n9421 & n9707;
  assign n9709 = n9421 & ~n9707;
  assign n9710 = ~n9708 & ~n9709;
  assign n9711 = pi114  & n391;
  assign n9712 = pi115  & n353;
  assign n9713 = pi116  & n348;
  assign n9714 = n346 & n8470;
  assign n9715 = ~n9712 & ~n9713;
  assign n9716 = ~n9711 & n9715;
  assign n9717 = ~n9714 & n9716;
  assign n9718 = pi5  & n9717;
  assign n9719 = ~pi5  & ~n9717;
  assign n9720 = ~n9718 & ~n9719;
  assign n9721 = n9710 & ~n9720;
  assign n9722 = ~n9710 & n9720;
  assign n9723 = ~n9721 & ~n9722;
  assign n9724 = ~n9420 & n9723;
  assign n9725 = n9420 & ~n9723;
  assign n9726 = ~n9724 & ~n9725;
  assign n9727 = ~n9419 & n9726;
  assign n9728 = n9419 & ~n9726;
  assign n9729 = ~n9727 & ~n9728;
  assign n9730 = ~n9402 & n9729;
  assign n9731 = n9402 & ~n9729;
  assign po55  = ~n9730 & ~n9731;
  assign n9733 = ~n9727 & ~n9730;
  assign n9734 = ~n9721 & ~n9724;
  assign n9735 = pi115  & n391;
  assign n9736 = pi116  & n353;
  assign n9737 = pi117  & n348;
  assign n9738 = n346 & n8784;
  assign n9739 = ~n9736 & ~n9737;
  assign n9740 = ~n9735 & n9739;
  assign n9741 = ~n9738 & n9740;
  assign n9742 = pi5  & n9741;
  assign n9743 = ~pi5  & ~n9741;
  assign n9744 = ~n9742 & ~n9743;
  assign n9745 = ~n9706 & ~n9708;
  assign n9746 = pi112  & n528;
  assign n9747 = pi113  & n490;
  assign n9748 = pi114  & n485;
  assign n9749 = n483 & n8146;
  assign n9750 = ~n9747 & ~n9748;
  assign n9751 = ~n9746 & n9750;
  assign n9752 = ~n9749 & n9751;
  assign n9753 = pi8  & n9752;
  assign n9754 = ~pi8  & ~n9752;
  assign n9755 = ~n9753 & ~n9754;
  assign n9756 = ~n9700 & ~n9702;
  assign n9757 = ~n9693 & ~n9696;
  assign n9758 = ~n9677 & ~n9681;
  assign n9759 = ~n9661 & ~n9665;
  assign n9760 = ~n9645 & ~n9649;
  assign n9761 = ~n9629 & ~n9633;
  assign n9762 = pi94  & n2510;
  assign n9763 = pi95  & n2342;
  assign n9764 = pi96  & n2337;
  assign n9765 = n2335 & n3499;
  assign n9766 = ~n9763 & ~n9764;
  assign n9767 = ~n9762 & n9766;
  assign n9768 = ~n9765 & n9767;
  assign n9769 = pi26  & n9768;
  assign n9770 = ~pi26  & ~n9768;
  assign n9771 = ~n9769 & ~n9770;
  assign n9772 = ~n9613 & ~n9617;
  assign n9773 = pi91  & n3011;
  assign n9774 = pi92  & n2809;
  assign n9775 = pi93  & n2804;
  assign n9776 = n2802 & n2948;
  assign n9777 = ~n9774 & ~n9775;
  assign n9778 = ~n9773 & n9777;
  assign n9779 = ~n9776 & n9778;
  assign n9780 = pi29  & n9779;
  assign n9781 = ~pi29  & ~n9779;
  assign n9782 = ~n9780 & ~n9781;
  assign n9783 = ~n9597 & ~n9601;
  assign n9784 = ~n9581 & ~n9585;
  assign n9785 = pi85  & n4176;
  assign n9786 = pi86  & n3938;
  assign n9787 = pi87  & n3933;
  assign n9788 = n2116 & n3931;
  assign n9789 = ~n9786 & ~n9787;
  assign n9790 = ~n9785 & n9789;
  assign n9791 = ~n9788 & n9790;
  assign n9792 = pi35  & n9791;
  assign n9793 = ~pi35  & ~n9791;
  assign n9794 = ~n9792 & ~n9793;
  assign n9795 = ~n9565 & ~n9568;
  assign n9796 = pi82  & n4843;
  assign n9797 = pi83  & n4598;
  assign n9798 = pi84  & n4593;
  assign n9799 = n1601 & n4591;
  assign n9800 = ~n9797 & ~n9798;
  assign n9801 = ~n9796 & n9800;
  assign n9802 = ~n9799 & n9801;
  assign n9803 = pi38  & n9802;
  assign n9804 = ~pi38  & ~n9802;
  assign n9805 = ~n9803 & ~n9804;
  assign n9806 = ~n9549 & ~n9553;
  assign n9807 = pi79  & n5558;
  assign n9808 = pi80  & n5293;
  assign n9809 = pi81  & n5288;
  assign n9810 = n1337 & n5286;
  assign n9811 = ~n9808 & ~n9809;
  assign n9812 = ~n9807 & n9811;
  assign n9813 = ~n9810 & n9812;
  assign n9814 = pi41  & n9813;
  assign n9815 = ~pi41  & ~n9813;
  assign n9816 = ~n9814 & ~n9815;
  assign n9817 = ~n9534 & ~n9536;
  assign n9818 = ~n9528 & ~n9530;
  assign n9819 = pi73  & n7121;
  assign n9820 = pi74  & n6795;
  assign n9821 = pi75  & n6790;
  assign n9822 = n713 & n6788;
  assign n9823 = ~n9820 & ~n9821;
  assign n9824 = ~n9819 & n9823;
  assign n9825 = ~n9822 & n9824;
  assign n9826 = pi47  & n9825;
  assign n9827 = ~pi47  & ~n9825;
  assign n9828 = ~n9826 & ~n9827;
  assign n9829 = ~n9522 & ~n9524;
  assign n9830 = pi70  & n7969;
  assign n9831 = pi71  & n7636;
  assign n9832 = pi72  & n7631;
  assign n9833 = n551 & n7629;
  assign n9834 = ~n9831 & ~n9832;
  assign n9835 = ~n9830 & n9834;
  assign n9836 = ~n9833 & n9835;
  assign n9837 = pi50  & n9836;
  assign n9838 = ~pi50  & ~n9836;
  assign n9839 = ~n9837 & ~n9838;
  assign n9840 = ~n9516 & ~n9518;
  assign n9841 = pi67  & n8905;
  assign n9842 = pi68  & n8535;
  assign n9843 = pi69  & n8530;
  assign n9844 = n376 & n8528;
  assign n9845 = ~n9842 & ~n9843;
  assign n9846 = ~n9841 & n9845;
  assign n9847 = ~n9844 & n9846;
  assign n9848 = pi53  & n9847;
  assign n9849 = ~pi53  & ~n9847;
  assign n9850 = ~n9848 & ~n9849;
  assign n9851 = pi56  & ~n9242;
  assign n9852 = n9511 & n9851;
  assign n9853 = pi56  & ~n9852;
  assign n9854 = ~n287 & n9501;
  assign n9855 = pi65  & n9508;
  assign n9856 = pi66  & n9503;
  assign n9857 = ~n9241 & n9500;
  assign n9858 = ~n9507 & n9857;
  assign n9859 = pi64  & n9858;
  assign n9860 = ~n9854 & ~n9855;
  assign n9861 = ~n9856 & n9860;
  assign n9862 = ~n9859 & n9861;
  assign n9863 = ~n9853 & n9862;
  assign n9864 = n9853 & ~n9862;
  assign n9865 = ~n9863 & ~n9864;
  assign n9866 = ~n9850 & n9865;
  assign n9867 = n9850 & ~n9865;
  assign n9868 = ~n9866 & ~n9867;
  assign n9869 = ~n9840 & n9868;
  assign n9870 = n9840 & ~n9868;
  assign n9871 = ~n9869 & ~n9870;
  assign n9872 = n9839 & ~n9871;
  assign n9873 = ~n9839 & n9871;
  assign n9874 = ~n9872 & ~n9873;
  assign n9875 = ~n9829 & n9874;
  assign n9876 = n9829 & ~n9874;
  assign n9877 = ~n9875 & ~n9876;
  assign n9878 = n9828 & ~n9877;
  assign n9879 = ~n9828 & n9877;
  assign n9880 = ~n9878 & ~n9879;
  assign n9881 = ~n9818 & n9880;
  assign n9882 = n9818 & ~n9880;
  assign n9883 = ~n9881 & ~n9882;
  assign n9884 = pi76  & n6331;
  assign n9885 = pi77  & n6015;
  assign n9886 = pi78  & n6010;
  assign n9887 = n958 & n6008;
  assign n9888 = ~n9885 & ~n9886;
  assign n9889 = ~n9884 & n9888;
  assign n9890 = ~n9887 & n9889;
  assign n9891 = pi44  & n9890;
  assign n9892 = ~pi44  & ~n9890;
  assign n9893 = ~n9891 & ~n9892;
  assign n9894 = n9883 & ~n9893;
  assign n9895 = ~n9883 & n9893;
  assign n9896 = ~n9894 & ~n9895;
  assign n9897 = ~n9817 & n9896;
  assign n9898 = n9817 & ~n9896;
  assign n9899 = ~n9897 & ~n9898;
  assign n9900 = ~n9816 & n9899;
  assign n9901 = n9816 & ~n9899;
  assign n9902 = ~n9900 & ~n9901;
  assign n9903 = ~n9806 & n9902;
  assign n9904 = n9806 & ~n9902;
  assign n9905 = ~n9903 & ~n9904;
  assign n9906 = ~n9805 & n9905;
  assign n9907 = n9805 & ~n9905;
  assign n9908 = ~n9906 & ~n9907;
  assign n9909 = ~n9795 & n9908;
  assign n9910 = n9795 & ~n9908;
  assign n9911 = ~n9909 & ~n9910;
  assign n9912 = ~n9794 & n9911;
  assign n9913 = n9794 & ~n9911;
  assign n9914 = ~n9912 & ~n9913;
  assign n9915 = n9784 & ~n9914;
  assign n9916 = ~n9784 & n9914;
  assign n9917 = ~n9915 & ~n9916;
  assign n9918 = pi88  & n3553;
  assign n9919 = pi89  & n3334;
  assign n9920 = pi90  & n3329;
  assign n9921 = n2448 & n3327;
  assign n9922 = ~n9919 & ~n9920;
  assign n9923 = ~n9918 & n9922;
  assign n9924 = ~n9921 & n9923;
  assign n9925 = pi32  & n9924;
  assign n9926 = ~pi32  & ~n9924;
  assign n9927 = ~n9925 & ~n9926;
  assign n9928 = n9917 & ~n9927;
  assign n9929 = ~n9917 & n9927;
  assign n9930 = ~n9928 & ~n9929;
  assign n9931 = ~n9783 & n9930;
  assign n9932 = n9783 & ~n9930;
  assign n9933 = ~n9931 & ~n9932;
  assign n9934 = n9782 & ~n9933;
  assign n9935 = ~n9782 & n9933;
  assign n9936 = ~n9934 & ~n9935;
  assign n9937 = ~n9772 & n9936;
  assign n9938 = n9772 & ~n9936;
  assign n9939 = ~n9937 & ~n9938;
  assign n9940 = n9771 & ~n9939;
  assign n9941 = ~n9771 & n9939;
  assign n9942 = ~n9940 & ~n9941;
  assign n9943 = ~n9761 & n9942;
  assign n9944 = n9761 & ~n9942;
  assign n9945 = ~n9943 & ~n9944;
  assign n9946 = pi97  & n2053;
  assign n9947 = pi98  & n1893;
  assign n9948 = pi99  & n1888;
  assign n9949 = n1886 & n4101;
  assign n9950 = ~n9947 & ~n9948;
  assign n9951 = ~n9946 & n9950;
  assign n9952 = ~n9949 & n9951;
  assign n9953 = pi23  & n9952;
  assign n9954 = ~pi23  & ~n9952;
  assign n9955 = ~n9953 & ~n9954;
  assign n9956 = n9945 & ~n9955;
  assign n9957 = ~n9945 & n9955;
  assign n9958 = ~n9956 & ~n9957;
  assign n9959 = n9760 & ~n9958;
  assign n9960 = ~n9760 & n9958;
  assign n9961 = ~n9959 & ~n9960;
  assign n9962 = pi100  & n1661;
  assign n9963 = pi101  & n1500;
  assign n9964 = pi102  & n1495;
  assign n9965 = n1493 & n4956;
  assign n9966 = ~n9963 & ~n9964;
  assign n9967 = ~n9962 & n9966;
  assign n9968 = ~n9965 & n9967;
  assign n9969 = pi20  & n9968;
  assign n9970 = ~pi20  & ~n9968;
  assign n9971 = ~n9969 & ~n9970;
  assign n9972 = n9961 & ~n9971;
  assign n9973 = ~n9961 & n9971;
  assign n9974 = ~n9972 & ~n9973;
  assign n9975 = n9759 & ~n9974;
  assign n9976 = ~n9759 & n9974;
  assign n9977 = ~n9975 & ~n9976;
  assign n9978 = pi103  & n1296;
  assign n9979 = pi104  & n1207;
  assign n9980 = pi105  & n1202;
  assign n9981 = n1200 & n5677;
  assign n9982 = ~n9979 & ~n9980;
  assign n9983 = ~n9978 & n9982;
  assign n9984 = ~n9981 & n9983;
  assign n9985 = pi17  & n9984;
  assign n9986 = ~pi17  & ~n9984;
  assign n9987 = ~n9985 & ~n9986;
  assign n9988 = n9977 & ~n9987;
  assign n9989 = ~n9977 & n9987;
  assign n9990 = ~n9988 & ~n9989;
  assign n9991 = n9758 & ~n9990;
  assign n9992 = ~n9758 & n9990;
  assign n9993 = ~n9991 & ~n9992;
  assign n9994 = pi106  & n1006;
  assign n9995 = pi107  & n897;
  assign n9996 = pi108  & n892;
  assign n9997 = n890 & n6213;
  assign n9998 = ~n9995 & ~n9996;
  assign n9999 = ~n9994 & n9998;
  assign n10000 = ~n9997 & n9999;
  assign n10001 = pi14  & n10000;
  assign n10002 = ~pi14  & ~n10000;
  assign n10003 = ~n10001 & ~n10002;
  assign n10004 = n9993 & ~n10003;
  assign n10005 = ~n9993 & n10003;
  assign n10006 = ~n10004 & ~n10005;
  assign n10007 = ~n9757 & n10006;
  assign n10008 = n9757 & ~n10006;
  assign n10009 = ~n10007 & ~n10008;
  assign n10010 = pi109  & n750;
  assign n10011 = pi110  & n651;
  assign n10012 = pi111  & n646;
  assign n10013 = n644 & n7272;
  assign n10014 = ~n10011 & ~n10012;
  assign n10015 = ~n10010 & n10014;
  assign n10016 = ~n10013 & n10015;
  assign n10017 = pi11  & n10016;
  assign n10018 = ~pi11  & ~n10016;
  assign n10019 = ~n10017 & ~n10018;
  assign n10020 = n10009 & ~n10019;
  assign n10021 = ~n10009 & n10019;
  assign n10022 = ~n10020 & ~n10021;
  assign n10023 = ~n9756 & n10022;
  assign n10024 = n9756 & ~n10022;
  assign n10025 = ~n10023 & ~n10024;
  assign n10026 = ~n9755 & n10025;
  assign n10027 = n9755 & ~n10025;
  assign n10028 = ~n10026 & ~n10027;
  assign n10029 = ~n9745 & n10028;
  assign n10030 = n9745 & ~n10028;
  assign n10031 = ~n10029 & ~n10030;
  assign n10032 = n9744 & ~n10031;
  assign n10033 = ~n9744 & n10031;
  assign n10034 = ~n10032 & ~n10033;
  assign n10035 = ~n9734 & n10034;
  assign n10036 = n9734 & ~n10034;
  assign n10037 = ~n10035 & ~n10036;
  assign n10038 = pi120  & n269;
  assign n10039 = pi119  & n267;
  assign n10040 = pi118  & n282;
  assign n10041 = ~n9408 & ~n9410;
  assign n10042 = ~pi119  & ~pi120 ;
  assign n10043 = pi119  & pi120 ;
  assign n10044 = ~n10042 & ~n10043;
  assign n10045 = ~n10041 & n10044;
  assign n10046 = n10041 & ~n10044;
  assign n10047 = ~n10045 & ~n10046;
  assign n10048 = n262 & n10047;
  assign n10049 = ~n10038 & ~n10039;
  assign n10050 = ~n10040 & n10049;
  assign n10051 = ~n10048 & n10050;
  assign n10052 = pi2  & n10051;
  assign n10053 = ~pi2  & ~n10051;
  assign n10054 = ~n10052 & ~n10053;
  assign n10055 = n10037 & ~n10054;
  assign n10056 = ~n10037 & n10054;
  assign n10057 = ~n10055 & ~n10056;
  assign n10058 = ~n9733 & n10057;
  assign n10059 = n9733 & ~n10057;
  assign po56  = ~n10058 & ~n10059;
  assign n10061 = ~n10055 & ~n10058;
  assign n10062 = pi121  & n269;
  assign n10063 = pi120  & n267;
  assign n10064 = pi119  & n282;
  assign n10065 = ~n10043 & ~n10045;
  assign n10066 = ~pi120  & ~pi121 ;
  assign n10067 = pi120  & pi121 ;
  assign n10068 = ~n10066 & ~n10067;
  assign n10069 = ~n10065 & n10068;
  assign n10070 = n10065 & ~n10068;
  assign n10071 = ~n10069 & ~n10070;
  assign n10072 = n262 & n10071;
  assign n10073 = ~n10062 & ~n10063;
  assign n10074 = ~n10064 & n10073;
  assign n10075 = ~n10072 & n10074;
  assign n10076 = pi2  & n10075;
  assign n10077 = ~pi2  & ~n10075;
  assign n10078 = ~n10076 & ~n10077;
  assign n10079 = ~n10033 & ~n10035;
  assign n10080 = pi116  & n391;
  assign n10081 = pi117  & n353;
  assign n10082 = pi118  & n348;
  assign n10083 = n346 & n9095;
  assign n10084 = ~n10081 & ~n10082;
  assign n10085 = ~n10080 & n10084;
  assign n10086 = ~n10083 & n10085;
  assign n10087 = pi5  & n10086;
  assign n10088 = ~pi5  & ~n10086;
  assign n10089 = ~n10087 & ~n10088;
  assign n10090 = ~n10026 & ~n10029;
  assign n10091 = pi113  & n528;
  assign n10092 = pi114  & n490;
  assign n10093 = pi115  & n485;
  assign n10094 = n483 & n8170;
  assign n10095 = ~n10092 & ~n10093;
  assign n10096 = ~n10091 & n10095;
  assign n10097 = ~n10094 & n10096;
  assign n10098 = pi8  & n10097;
  assign n10099 = ~pi8  & ~n10097;
  assign n10100 = ~n10098 & ~n10099;
  assign n10101 = ~n10020 & ~n10023;
  assign n10102 = pi110  & n750;
  assign n10103 = pi111  & n651;
  assign n10104 = pi112  & n646;
  assign n10105 = n644 & n7296;
  assign n10106 = ~n10103 & ~n10104;
  assign n10107 = ~n10102 & n10106;
  assign n10108 = ~n10105 & n10107;
  assign n10109 = pi11  & n10108;
  assign n10110 = ~pi11  & ~n10108;
  assign n10111 = ~n10109 & ~n10110;
  assign n10112 = ~n10004 & ~n10007;
  assign n10113 = pi107  & n1006;
  assign n10114 = pi108  & n897;
  assign n10115 = pi109  & n892;
  assign n10116 = n890 & n6715;
  assign n10117 = ~n10114 & ~n10115;
  assign n10118 = ~n10113 & n10117;
  assign n10119 = ~n10116 & n10118;
  assign n10120 = pi14  & n10119;
  assign n10121 = ~pi14  & ~n10119;
  assign n10122 = ~n10120 & ~n10121;
  assign n10123 = ~n9988 & ~n9992;
  assign n10124 = ~n9972 & ~n9976;
  assign n10125 = ~n9956 & ~n9960;
  assign n10126 = pi98  & n2053;
  assign n10127 = pi99  & n1893;
  assign n10128 = pi100  & n1888;
  assign n10129 = n1886 & n4501;
  assign n10130 = ~n10127 & ~n10128;
  assign n10131 = ~n10126 & n10130;
  assign n10132 = ~n10129 & n10131;
  assign n10133 = pi23  & n10132;
  assign n10134 = ~pi23  & ~n10132;
  assign n10135 = ~n10133 & ~n10134;
  assign n10136 = ~n9941 & ~n9943;
  assign n10137 = ~n9935 & ~n9937;
  assign n10138 = pi92  & n3011;
  assign n10139 = pi93  & n2809;
  assign n10140 = pi94  & n2804;
  assign n10141 = n2802 & n3280;
  assign n10142 = ~n10139 & ~n10140;
  assign n10143 = ~n10138 & n10142;
  assign n10144 = ~n10141 & n10143;
  assign n10145 = pi29  & n10144;
  assign n10146 = ~pi29  & ~n10144;
  assign n10147 = ~n10145 & ~n10146;
  assign n10148 = ~n9928 & ~n9931;
  assign n10149 = ~n9912 & ~n9916;
  assign n10150 = ~n9906 & ~n9909;
  assign n10151 = pi83  & n4843;
  assign n10152 = pi84  & n4598;
  assign n10153 = pi85  & n4593;
  assign n10154 = n1831 & n4591;
  assign n10155 = ~n10152 & ~n10153;
  assign n10156 = ~n10151 & n10155;
  assign n10157 = ~n10154 & n10156;
  assign n10158 = pi38  & n10157;
  assign n10159 = ~pi38  & ~n10157;
  assign n10160 = ~n10158 & ~n10159;
  assign n10161 = ~n9900 & ~n9903;
  assign n10162 = pi80  & n5558;
  assign n10163 = pi81  & n5293;
  assign n10164 = pi82  & n5288;
  assign n10165 = n1450 & n5286;
  assign n10166 = ~n10163 & ~n10164;
  assign n10167 = ~n10162 & n10166;
  assign n10168 = ~n10165 & n10167;
  assign n10169 = pi41  & n10168;
  assign n10170 = ~pi41  & ~n10168;
  assign n10171 = ~n10169 & ~n10170;
  assign n10172 = ~n9894 & ~n9897;
  assign n10173 = pi77  & n6331;
  assign n10174 = pi78  & n6015;
  assign n10175 = pi79  & n6010;
  assign n10176 = n1048 & n6008;
  assign n10177 = ~n10174 & ~n10175;
  assign n10178 = ~n10173 & n10177;
  assign n10179 = ~n10176 & n10178;
  assign n10180 = pi44  & n10179;
  assign n10181 = ~pi44  & ~n10179;
  assign n10182 = ~n10180 & ~n10181;
  assign n10183 = ~n9879 & ~n9881;
  assign n10184 = pi74  & n7121;
  assign n10185 = pi75  & n6795;
  assign n10186 = pi76  & n6790;
  assign n10187 = n841 & n6788;
  assign n10188 = ~n10185 & ~n10186;
  assign n10189 = ~n10184 & n10188;
  assign n10190 = ~n10187 & n10189;
  assign n10191 = pi47  & n10190;
  assign n10192 = ~pi47  & ~n10190;
  assign n10193 = ~n10191 & ~n10192;
  assign n10194 = ~n9873 & ~n9875;
  assign n10195 = pi71  & n7969;
  assign n10196 = pi72  & n7636;
  assign n10197 = pi73  & n7631;
  assign n10198 = n613 & n7629;
  assign n10199 = ~n10196 & ~n10197;
  assign n10200 = ~n10195 & n10199;
  assign n10201 = ~n10198 & n10200;
  assign n10202 = pi50  & n10201;
  assign n10203 = ~pi50  & ~n10201;
  assign n10204 = ~n10202 & ~n10203;
  assign n10205 = ~n9866 & ~n9869;
  assign n10206 = pi65  & n9858;
  assign n10207 = pi66  & n9508;
  assign n10208 = pi67  & n9503;
  assign n10209 = n305 & n9501;
  assign n10210 = ~n10207 & ~n10208;
  assign n10211 = ~n10206 & n10210;
  assign n10212 = ~n10209 & n10211;
  assign n10213 = pi56  & n10212;
  assign n10214 = ~pi56  & ~n10212;
  assign n10215 = ~n10213 & ~n10214;
  assign n10216 = ~pi56  & ~pi57 ;
  assign n10217 = pi56  & pi57 ;
  assign n10218 = ~n10216 & ~n10217;
  assign n10219 = pi64  & n10218;
  assign n10220 = n9852 & n9862;
  assign n10221 = n10219 & n10220;
  assign n10222 = ~n10219 & ~n10220;
  assign n10223 = ~n10221 & ~n10222;
  assign n10224 = ~n10215 & n10223;
  assign n10225 = n10215 & ~n10223;
  assign n10226 = ~n10224 & ~n10225;
  assign n10227 = pi68  & n8905;
  assign n10228 = pi69  & n8535;
  assign n10229 = pi70  & n8530;
  assign n10230 = n415 & n8528;
  assign n10231 = ~n10228 & ~n10229;
  assign n10232 = ~n10227 & n10231;
  assign n10233 = ~n10230 & n10232;
  assign n10234 = pi53  & n10233;
  assign n10235 = ~pi53  & ~n10233;
  assign n10236 = ~n10234 & ~n10235;
  assign n10237 = n10226 & ~n10236;
  assign n10238 = ~n10226 & n10236;
  assign n10239 = ~n10237 & ~n10238;
  assign n10240 = ~n10205 & n10239;
  assign n10241 = n10205 & ~n10239;
  assign n10242 = ~n10240 & ~n10241;
  assign n10243 = ~n10204 & n10242;
  assign n10244 = n10204 & ~n10242;
  assign n10245 = ~n10243 & ~n10244;
  assign n10246 = ~n10194 & n10245;
  assign n10247 = n10194 & ~n10245;
  assign n10248 = ~n10246 & ~n10247;
  assign n10249 = n10193 & ~n10248;
  assign n10250 = ~n10193 & n10248;
  assign n10251 = ~n10249 & ~n10250;
  assign n10252 = ~n10183 & n10251;
  assign n10253 = n10183 & ~n10251;
  assign n10254 = ~n10252 & ~n10253;
  assign n10255 = ~n10182 & n10254;
  assign n10256 = n10182 & ~n10254;
  assign n10257 = ~n10255 & ~n10256;
  assign n10258 = ~n10172 & n10257;
  assign n10259 = n10172 & ~n10257;
  assign n10260 = ~n10258 & ~n10259;
  assign n10261 = ~n10171 & n10260;
  assign n10262 = n10171 & ~n10260;
  assign n10263 = ~n10261 & ~n10262;
  assign n10264 = ~n10161 & n10263;
  assign n10265 = n10161 & ~n10263;
  assign n10266 = ~n10264 & ~n10265;
  assign n10267 = ~n10160 & n10266;
  assign n10268 = n10160 & ~n10266;
  assign n10269 = ~n10267 & ~n10268;
  assign n10270 = ~n10150 & n10269;
  assign n10271 = n10150 & ~n10269;
  assign n10272 = ~n10270 & ~n10271;
  assign n10273 = pi86  & n4176;
  assign n10274 = pi87  & n3938;
  assign n10275 = pi88  & n3933;
  assign n10276 = n2140 & n3931;
  assign n10277 = ~n10274 & ~n10275;
  assign n10278 = ~n10273 & n10277;
  assign n10279 = ~n10276 & n10278;
  assign n10280 = pi35  & n10279;
  assign n10281 = ~pi35  & ~n10279;
  assign n10282 = ~n10280 & ~n10281;
  assign n10283 = n10272 & ~n10282;
  assign n10284 = ~n10272 & n10282;
  assign n10285 = ~n10283 & ~n10284;
  assign n10286 = n10149 & ~n10285;
  assign n10287 = ~n10149 & n10285;
  assign n10288 = ~n10286 & ~n10287;
  assign n10289 = pi89  & n3553;
  assign n10290 = pi90  & n3334;
  assign n10291 = pi91  & n3329;
  assign n10292 = n2746 & n3327;
  assign n10293 = ~n10290 & ~n10291;
  assign n10294 = ~n10289 & n10293;
  assign n10295 = ~n10292 & n10294;
  assign n10296 = pi32  & n10295;
  assign n10297 = ~pi32  & ~n10295;
  assign n10298 = ~n10296 & ~n10297;
  assign n10299 = ~n10288 & n10298;
  assign n10300 = n10288 & ~n10298;
  assign n10301 = ~n10299 & ~n10300;
  assign n10302 = ~n10148 & n10301;
  assign n10303 = n10148 & ~n10301;
  assign n10304 = ~n10302 & ~n10303;
  assign n10305 = ~n10147 & n10304;
  assign n10306 = n10147 & ~n10304;
  assign n10307 = ~n10305 & ~n10306;
  assign n10308 = ~n10137 & n10307;
  assign n10309 = n10137 & ~n10307;
  assign n10310 = ~n10308 & ~n10309;
  assign n10311 = pi95  & n2510;
  assign n10312 = pi96  & n2342;
  assign n10313 = pi97  & n2337;
  assign n10314 = n2335 & n3691;
  assign n10315 = ~n10312 & ~n10313;
  assign n10316 = ~n10311 & n10315;
  assign n10317 = ~n10314 & n10316;
  assign n10318 = pi26  & n10317;
  assign n10319 = ~pi26  & ~n10317;
  assign n10320 = ~n10318 & ~n10319;
  assign n10321 = n10310 & ~n10320;
  assign n10322 = ~n10310 & n10320;
  assign n10323 = ~n10321 & ~n10322;
  assign n10324 = ~n10136 & n10323;
  assign n10325 = n10136 & ~n10323;
  assign n10326 = ~n10324 & ~n10325;
  assign n10327 = ~n10135 & n10326;
  assign n10328 = n10135 & ~n10326;
  assign n10329 = ~n10327 & ~n10328;
  assign n10330 = n10125 & ~n10329;
  assign n10331 = ~n10125 & n10329;
  assign n10332 = ~n10330 & ~n10331;
  assign n10333 = pi101  & n1661;
  assign n10334 = pi102  & n1500;
  assign n10335 = pi103  & n1495;
  assign n10336 = n1493 & n5188;
  assign n10337 = ~n10334 & ~n10335;
  assign n10338 = ~n10333 & n10337;
  assign n10339 = ~n10336 & n10338;
  assign n10340 = pi20  & n10339;
  assign n10341 = ~pi20  & ~n10339;
  assign n10342 = ~n10340 & ~n10341;
  assign n10343 = n10332 & ~n10342;
  assign n10344 = ~n10332 & n10342;
  assign n10345 = ~n10343 & ~n10344;
  assign n10346 = n10124 & ~n10345;
  assign n10347 = ~n10124 & n10345;
  assign n10348 = ~n10346 & ~n10347;
  assign n10349 = pi104  & n1296;
  assign n10350 = pi105  & n1207;
  assign n10351 = pi106  & n1202;
  assign n10352 = n1200 & n5701;
  assign n10353 = ~n10350 & ~n10351;
  assign n10354 = ~n10349 & n10353;
  assign n10355 = ~n10352 & n10354;
  assign n10356 = pi17  & n10355;
  assign n10357 = ~pi17  & ~n10355;
  assign n10358 = ~n10356 & ~n10357;
  assign n10359 = ~n10348 & n10358;
  assign n10360 = n10348 & ~n10358;
  assign n10361 = ~n10359 & ~n10360;
  assign n10362 = ~n10123 & n10361;
  assign n10363 = n10123 & ~n10361;
  assign n10364 = ~n10362 & ~n10363;
  assign n10365 = ~n10122 & n10364;
  assign n10366 = n10122 & ~n10364;
  assign n10367 = ~n10365 & ~n10366;
  assign n10368 = ~n10112 & n10367;
  assign n10369 = n10112 & ~n10367;
  assign n10370 = ~n10368 & ~n10369;
  assign n10371 = ~n10111 & n10370;
  assign n10372 = n10111 & ~n10370;
  assign n10373 = ~n10371 & ~n10372;
  assign n10374 = ~n10101 & n10373;
  assign n10375 = n10101 & ~n10373;
  assign n10376 = ~n10374 & ~n10375;
  assign n10377 = ~n10100 & n10376;
  assign n10378 = n10100 & ~n10376;
  assign n10379 = ~n10377 & ~n10378;
  assign n10380 = ~n10090 & n10379;
  assign n10381 = n10090 & ~n10379;
  assign n10382 = ~n10380 & ~n10381;
  assign n10383 = ~n10089 & n10382;
  assign n10384 = n10089 & ~n10382;
  assign n10385 = ~n10383 & ~n10384;
  assign n10386 = ~n10079 & n10385;
  assign n10387 = n10079 & ~n10385;
  assign n10388 = ~n10386 & ~n10387;
  assign n10389 = ~n10078 & n10388;
  assign n10390 = n10078 & ~n10388;
  assign n10391 = ~n10389 & ~n10390;
  assign n10392 = ~n10061 & n10391;
  assign n10393 = n10061 & ~n10391;
  assign po57  = ~n10392 & ~n10393;
  assign n10395 = ~n10389 & ~n10392;
  assign n10396 = ~n10383 & ~n10386;
  assign n10397 = pi117  & n391;
  assign n10398 = pi118  & n353;
  assign n10399 = pi119  & n348;
  assign n10400 = n346 & n9412;
  assign n10401 = ~n10398 & ~n10399;
  assign n10402 = ~n10397 & n10401;
  assign n10403 = ~n10400 & n10402;
  assign n10404 = pi5  & n10403;
  assign n10405 = ~pi5  & ~n10403;
  assign n10406 = ~n10404 & ~n10405;
  assign n10407 = ~n10377 & ~n10380;
  assign n10408 = pi114  & n528;
  assign n10409 = pi115  & n490;
  assign n10410 = pi116  & n485;
  assign n10411 = n483 & n8470;
  assign n10412 = ~n10409 & ~n10410;
  assign n10413 = ~n10408 & n10412;
  assign n10414 = ~n10411 & n10413;
  assign n10415 = pi8  & n10414;
  assign n10416 = ~pi8  & ~n10414;
  assign n10417 = ~n10415 & ~n10416;
  assign n10418 = ~n10371 & ~n10374;
  assign n10419 = pi111  & n750;
  assign n10420 = pi112  & n651;
  assign n10421 = pi113  & n646;
  assign n10422 = n644 & n7852;
  assign n10423 = ~n10420 & ~n10421;
  assign n10424 = ~n10419 & n10423;
  assign n10425 = ~n10422 & n10424;
  assign n10426 = pi11  & n10425;
  assign n10427 = ~pi11  & ~n10425;
  assign n10428 = ~n10426 & ~n10427;
  assign n10429 = ~n10365 & ~n10368;
  assign n10430 = pi108  & n1006;
  assign n10431 = pi109  & n897;
  assign n10432 = pi110  & n892;
  assign n10433 = n890 & n6995;
  assign n10434 = ~n10431 & ~n10432;
  assign n10435 = ~n10430 & n10434;
  assign n10436 = ~n10433 & n10435;
  assign n10437 = pi14  & n10436;
  assign n10438 = ~pi14  & ~n10436;
  assign n10439 = ~n10437 & ~n10438;
  assign n10440 = ~n10360 & ~n10362;
  assign n10441 = ~n10343 & ~n10347;
  assign n10442 = ~n10327 & ~n10331;
  assign n10443 = ~n10321 & ~n10324;
  assign n10444 = ~n10305 & ~n10308;
  assign n10445 = pi93  & n3011;
  assign n10446 = pi94  & n2809;
  assign n10447 = pi95  & n2804;
  assign n10448 = n2802 & n3475;
  assign n10449 = ~n10446 & ~n10447;
  assign n10450 = ~n10445 & n10449;
  assign n10451 = ~n10448 & n10450;
  assign n10452 = pi29  & n10451;
  assign n10453 = ~pi29  & ~n10451;
  assign n10454 = ~n10452 & ~n10453;
  assign n10455 = ~n10300 & ~n10302;
  assign n10456 = ~n10283 & ~n10287;
  assign n10457 = ~n10267 & ~n10270;
  assign n10458 = ~n10261 & ~n10264;
  assign n10459 = ~n10255 & ~n10258;
  assign n10460 = ~n10250 & ~n10252;
  assign n10461 = ~n10243 & ~n10246;
  assign n10462 = ~n10237 & ~n10240;
  assign n10463 = pi69  & n8905;
  assign n10464 = pi70  & n8535;
  assign n10465 = pi71  & n8530;
  assign n10466 = n460 & n8528;
  assign n10467 = ~n10464 & ~n10465;
  assign n10468 = ~n10463 & n10467;
  assign n10469 = ~n10466 & n10468;
  assign n10470 = pi53  & n10469;
  assign n10471 = ~pi53  & ~n10469;
  assign n10472 = ~n10470 & ~n10471;
  assign n10473 = ~n10221 & ~n10224;
  assign n10474 = pi66  & n9858;
  assign n10475 = pi67  & n9508;
  assign n10476 = pi68  & n9503;
  assign n10477 = n334 & n9501;
  assign n10478 = ~n10475 & ~n10476;
  assign n10479 = ~n10474 & n10478;
  assign n10480 = ~n10477 & n10479;
  assign n10481 = pi56  & n10480;
  assign n10482 = ~pi56  & ~n10480;
  assign n10483 = ~n10481 & ~n10482;
  assign n10484 = pi59  & n10219;
  assign n10485 = ~pi58  & ~pi59 ;
  assign n10486 = pi58  & pi59 ;
  assign n10487 = ~n10485 & ~n10486;
  assign n10488 = n10218 & n10487;
  assign n10489 = n265 & n10488;
  assign n10490 = n10218 & ~n10487;
  assign n10491 = pi65  & n10490;
  assign n10492 = ~pi57  & ~pi58 ;
  assign n10493 = pi57  & pi58 ;
  assign n10494 = ~n10492 & ~n10493;
  assign n10495 = ~n10218 & n10494;
  assign n10496 = pi64  & n10495;
  assign n10497 = ~n10489 & ~n10491;
  assign n10498 = ~n10496 & n10497;
  assign n10499 = n10484 & ~n10498;
  assign n10500 = ~n10484 & n10498;
  assign n10501 = ~n10499 & ~n10500;
  assign n10502 = n10483 & ~n10501;
  assign n10503 = ~n10483 & n10501;
  assign n10504 = ~n10502 & ~n10503;
  assign n10505 = ~n10473 & n10504;
  assign n10506 = n10473 & ~n10504;
  assign n10507 = ~n10505 & ~n10506;
  assign n10508 = n10472 & ~n10507;
  assign n10509 = ~n10472 & n10507;
  assign n10510 = ~n10508 & ~n10509;
  assign n10511 = ~n10462 & n10510;
  assign n10512 = n10462 & ~n10510;
  assign n10513 = ~n10511 & ~n10512;
  assign n10514 = pi72  & n7969;
  assign n10515 = pi73  & n7636;
  assign n10516 = pi74  & n7631;
  assign n10517 = n689 & n7629;
  assign n10518 = ~n10515 & ~n10516;
  assign n10519 = ~n10514 & n10518;
  assign n10520 = ~n10517 & n10519;
  assign n10521 = pi50  & n10520;
  assign n10522 = ~pi50  & ~n10520;
  assign n10523 = ~n10521 & ~n10522;
  assign n10524 = n10513 & ~n10523;
  assign n10525 = ~n10513 & n10523;
  assign n10526 = ~n10524 & ~n10525;
  assign n10527 = n10461 & ~n10526;
  assign n10528 = ~n10461 & n10526;
  assign n10529 = ~n10527 & ~n10528;
  assign n10530 = pi75  & n7121;
  assign n10531 = pi76  & n6795;
  assign n10532 = pi77  & n6790;
  assign n10533 = n865 & n6788;
  assign n10534 = ~n10531 & ~n10532;
  assign n10535 = ~n10530 & n10534;
  assign n10536 = ~n10533 & n10535;
  assign n10537 = pi47  & n10536;
  assign n10538 = ~pi47  & ~n10536;
  assign n10539 = ~n10537 & ~n10538;
  assign n10540 = n10529 & ~n10539;
  assign n10541 = ~n10529 & n10539;
  assign n10542 = ~n10540 & ~n10541;
  assign n10543 = ~n10460 & n10542;
  assign n10544 = n10460 & ~n10542;
  assign n10545 = ~n10543 & ~n10544;
  assign n10546 = pi78  & n6331;
  assign n10547 = pi79  & n6015;
  assign n10548 = pi80  & n6010;
  assign n10549 = n1144 & n6008;
  assign n10550 = ~n10547 & ~n10548;
  assign n10551 = ~n10546 & n10550;
  assign n10552 = ~n10549 & n10551;
  assign n10553 = pi44  & n10552;
  assign n10554 = ~pi44  & ~n10552;
  assign n10555 = ~n10553 & ~n10554;
  assign n10556 = n10545 & ~n10555;
  assign n10557 = ~n10545 & n10555;
  assign n10558 = ~n10556 & ~n10557;
  assign n10559 = n10459 & ~n10558;
  assign n10560 = ~n10459 & n10558;
  assign n10561 = ~n10559 & ~n10560;
  assign n10562 = pi81  & n5558;
  assign n10563 = pi82  & n5293;
  assign n10564 = pi83  & n5288;
  assign n10565 = n1577 & n5286;
  assign n10566 = ~n10563 & ~n10564;
  assign n10567 = ~n10562 & n10566;
  assign n10568 = ~n10565 & n10567;
  assign n10569 = pi41  & n10568;
  assign n10570 = ~pi41  & ~n10568;
  assign n10571 = ~n10569 & ~n10570;
  assign n10572 = n10561 & ~n10571;
  assign n10573 = ~n10561 & n10571;
  assign n10574 = ~n10572 & ~n10573;
  assign n10575 = ~n10458 & n10574;
  assign n10576 = n10458 & ~n10574;
  assign n10577 = ~n10575 & ~n10576;
  assign n10578 = pi84  & n4843;
  assign n10579 = pi85  & n4598;
  assign n10580 = pi86  & n4593;
  assign n10581 = n1975 & n4591;
  assign n10582 = ~n10579 & ~n10580;
  assign n10583 = ~n10578 & n10582;
  assign n10584 = ~n10581 & n10583;
  assign n10585 = pi38  & n10584;
  assign n10586 = ~pi38  & ~n10584;
  assign n10587 = ~n10585 & ~n10586;
  assign n10588 = n10577 & ~n10587;
  assign n10589 = ~n10577 & n10587;
  assign n10590 = ~n10588 & ~n10589;
  assign n10591 = n10457 & ~n10590;
  assign n10592 = ~n10457 & n10590;
  assign n10593 = ~n10591 & ~n10592;
  assign n10594 = pi87  & n4176;
  assign n10595 = pi88  & n3938;
  assign n10596 = pi89  & n3933;
  assign n10597 = n2287 & n3931;
  assign n10598 = ~n10595 & ~n10596;
  assign n10599 = ~n10594 & n10598;
  assign n10600 = ~n10597 & n10599;
  assign n10601 = pi35  & n10600;
  assign n10602 = ~pi35  & ~n10600;
  assign n10603 = ~n10601 & ~n10602;
  assign n10604 = n10593 & ~n10603;
  assign n10605 = ~n10593 & n10603;
  assign n10606 = ~n10604 & ~n10605;
  assign n10607 = n10456 & ~n10606;
  assign n10608 = ~n10456 & n10606;
  assign n10609 = ~n10607 & ~n10608;
  assign n10610 = pi90  & n3553;
  assign n10611 = pi91  & n3334;
  assign n10612 = pi92  & n3329;
  assign n10613 = n2924 & n3327;
  assign n10614 = ~n10611 & ~n10612;
  assign n10615 = ~n10610 & n10614;
  assign n10616 = ~n10613 & n10615;
  assign n10617 = pi32  & n10616;
  assign n10618 = ~pi32  & ~n10616;
  assign n10619 = ~n10617 & ~n10618;
  assign n10620 = n10609 & ~n10619;
  assign n10621 = ~n10609 & n10619;
  assign n10622 = ~n10620 & ~n10621;
  assign n10623 = ~n10455 & n10622;
  assign n10624 = n10455 & ~n10622;
  assign n10625 = ~n10623 & ~n10624;
  assign n10626 = ~n10454 & n10625;
  assign n10627 = n10454 & ~n10625;
  assign n10628 = ~n10626 & ~n10627;
  assign n10629 = n10444 & ~n10628;
  assign n10630 = ~n10444 & n10628;
  assign n10631 = ~n10629 & ~n10630;
  assign n10632 = pi96  & n2510;
  assign n10633 = pi97  & n2342;
  assign n10634 = pi98  & n2337;
  assign n10635 = n2335 & n3889;
  assign n10636 = ~n10633 & ~n10634;
  assign n10637 = ~n10632 & n10636;
  assign n10638 = ~n10635 & n10637;
  assign n10639 = pi26  & n10638;
  assign n10640 = ~pi26  & ~n10638;
  assign n10641 = ~n10639 & ~n10640;
  assign n10642 = n10631 & ~n10641;
  assign n10643 = ~n10631 & n10641;
  assign n10644 = ~n10642 & ~n10643;
  assign n10645 = n10443 & ~n10644;
  assign n10646 = ~n10443 & n10644;
  assign n10647 = ~n10645 & ~n10646;
  assign n10648 = pi99  & n2053;
  assign n10649 = pi100  & n1893;
  assign n10650 = pi101  & n1888;
  assign n10651 = n1886 & n4730;
  assign n10652 = ~n10649 & ~n10650;
  assign n10653 = ~n10648 & n10652;
  assign n10654 = ~n10651 & n10653;
  assign n10655 = pi23  & n10654;
  assign n10656 = ~pi23  & ~n10654;
  assign n10657 = ~n10655 & ~n10656;
  assign n10658 = n10647 & ~n10657;
  assign n10659 = ~n10647 & n10657;
  assign n10660 = ~n10658 & ~n10659;
  assign n10661 = n10442 & ~n10660;
  assign n10662 = ~n10442 & n10660;
  assign n10663 = ~n10661 & ~n10662;
  assign n10664 = pi102  & n1661;
  assign n10665 = pi103  & n1500;
  assign n10666 = pi104  & n1495;
  assign n10667 = n1493 & n5212;
  assign n10668 = ~n10665 & ~n10666;
  assign n10669 = ~n10664 & n10668;
  assign n10670 = ~n10667 & n10669;
  assign n10671 = pi20  & n10670;
  assign n10672 = ~pi20  & ~n10670;
  assign n10673 = ~n10671 & ~n10672;
  assign n10674 = n10663 & ~n10673;
  assign n10675 = ~n10663 & n10673;
  assign n10676 = ~n10674 & ~n10675;
  assign n10677 = n10441 & ~n10676;
  assign n10678 = ~n10441 & n10676;
  assign n10679 = ~n10677 & ~n10678;
  assign n10680 = pi105  & n1296;
  assign n10681 = pi106  & n1207;
  assign n10682 = pi107  & n1202;
  assign n10683 = n1200 & n6189;
  assign n10684 = ~n10681 & ~n10682;
  assign n10685 = ~n10680 & n10684;
  assign n10686 = ~n10683 & n10685;
  assign n10687 = pi17  & n10686;
  assign n10688 = ~pi17  & ~n10686;
  assign n10689 = ~n10687 & ~n10688;
  assign n10690 = n10679 & ~n10689;
  assign n10691 = ~n10679 & n10689;
  assign n10692 = ~n10690 & ~n10691;
  assign n10693 = ~n10440 & n10692;
  assign n10694 = n10440 & ~n10692;
  assign n10695 = ~n10693 & ~n10694;
  assign n10696 = n10439 & ~n10695;
  assign n10697 = ~n10439 & n10695;
  assign n10698 = ~n10696 & ~n10697;
  assign n10699 = ~n10429 & n10698;
  assign n10700 = n10429 & ~n10698;
  assign n10701 = ~n10699 & ~n10700;
  assign n10702 = n10428 & ~n10701;
  assign n10703 = ~n10428 & n10701;
  assign n10704 = ~n10702 & ~n10703;
  assign n10705 = ~n10418 & n10704;
  assign n10706 = n10418 & ~n10704;
  assign n10707 = ~n10705 & ~n10706;
  assign n10708 = n10417 & ~n10707;
  assign n10709 = ~n10417 & n10707;
  assign n10710 = ~n10708 & ~n10709;
  assign n10711 = ~n10407 & n10710;
  assign n10712 = n10407 & ~n10710;
  assign n10713 = ~n10711 & ~n10712;
  assign n10714 = n10406 & ~n10713;
  assign n10715 = ~n10406 & n10713;
  assign n10716 = ~n10714 & ~n10715;
  assign n10717 = ~n10396 & n10716;
  assign n10718 = n10396 & ~n10716;
  assign n10719 = ~n10717 & ~n10718;
  assign n10720 = pi122  & n269;
  assign n10721 = pi121  & n267;
  assign n10722 = pi120  & n282;
  assign n10723 = ~n10067 & ~n10069;
  assign n10724 = ~pi121  & ~pi122 ;
  assign n10725 = pi121  & pi122 ;
  assign n10726 = ~n10724 & ~n10725;
  assign n10727 = ~n10723 & n10726;
  assign n10728 = n10723 & ~n10726;
  assign n10729 = ~n10727 & ~n10728;
  assign n10730 = n262 & n10729;
  assign n10731 = ~n10720 & ~n10721;
  assign n10732 = ~n10722 & n10731;
  assign n10733 = ~n10730 & n10732;
  assign n10734 = pi2  & n10733;
  assign n10735 = ~pi2  & ~n10733;
  assign n10736 = ~n10734 & ~n10735;
  assign n10737 = n10719 & ~n10736;
  assign n10738 = ~n10719 & n10736;
  assign n10739 = ~n10737 & ~n10738;
  assign n10740 = ~n10395 & n10739;
  assign n10741 = n10395 & ~n10739;
  assign po58  = ~n10740 & ~n10741;
  assign n10743 = ~n10737 & ~n10740;
  assign n10744 = ~n10715 & ~n10717;
  assign n10745 = pi123  & n269;
  assign n10746 = pi122  & n267;
  assign n10747 = pi121  & n282;
  assign n10748 = ~n10725 & ~n10727;
  assign n10749 = ~pi122  & ~pi123 ;
  assign n10750 = pi122  & pi123 ;
  assign n10751 = ~n10749 & ~n10750;
  assign n10752 = ~n10748 & n10751;
  assign n10753 = n10748 & ~n10751;
  assign n10754 = ~n10752 & ~n10753;
  assign n10755 = n262 & n10754;
  assign n10756 = ~n10745 & ~n10746;
  assign n10757 = ~n10747 & n10756;
  assign n10758 = ~n10755 & n10757;
  assign n10759 = pi2  & n10758;
  assign n10760 = ~pi2  & ~n10758;
  assign n10761 = ~n10759 & ~n10760;
  assign n10762 = pi118  & n391;
  assign n10763 = pi119  & n353;
  assign n10764 = pi120  & n348;
  assign n10765 = n346 & n10047;
  assign n10766 = ~n10763 & ~n10764;
  assign n10767 = ~n10762 & n10766;
  assign n10768 = ~n10765 & n10767;
  assign n10769 = pi5  & n10768;
  assign n10770 = ~pi5  & ~n10768;
  assign n10771 = ~n10769 & ~n10770;
  assign n10772 = ~n10709 & ~n10711;
  assign n10773 = pi115  & n528;
  assign n10774 = pi116  & n490;
  assign n10775 = pi117  & n485;
  assign n10776 = n483 & n8784;
  assign n10777 = ~n10774 & ~n10775;
  assign n10778 = ~n10773 & n10777;
  assign n10779 = ~n10776 & n10778;
  assign n10780 = pi8  & n10779;
  assign n10781 = ~pi8  & ~n10779;
  assign n10782 = ~n10780 & ~n10781;
  assign n10783 = ~n10703 & ~n10705;
  assign n10784 = ~n10697 & ~n10699;
  assign n10785 = pi109  & n1006;
  assign n10786 = pi110  & n897;
  assign n10787 = pi111  & n892;
  assign n10788 = n890 & n7272;
  assign n10789 = ~n10786 & ~n10787;
  assign n10790 = ~n10785 & n10789;
  assign n10791 = ~n10788 & n10790;
  assign n10792 = pi14  & n10791;
  assign n10793 = ~pi14  & ~n10791;
  assign n10794 = ~n10792 & ~n10793;
  assign n10795 = ~n10690 & ~n10693;
  assign n10796 = ~n10674 & ~n10678;
  assign n10797 = ~n10658 & ~n10662;
  assign n10798 = ~n10642 & ~n10646;
  assign n10799 = ~n10626 & ~n10630;
  assign n10800 = pi94  & n3011;
  assign n10801 = pi95  & n2809;
  assign n10802 = pi96  & n2804;
  assign n10803 = n2802 & n3499;
  assign n10804 = ~n10801 & ~n10802;
  assign n10805 = ~n10800 & n10804;
  assign n10806 = ~n10803 & n10805;
  assign n10807 = pi29  & n10806;
  assign n10808 = ~pi29  & ~n10806;
  assign n10809 = ~n10807 & ~n10808;
  assign n10810 = ~n10620 & ~n10623;
  assign n10811 = ~n10604 & ~n10608;
  assign n10812 = ~n10588 & ~n10592;
  assign n10813 = pi85  & n4843;
  assign n10814 = pi86  & n4598;
  assign n10815 = pi87  & n4593;
  assign n10816 = n2116 & n4591;
  assign n10817 = ~n10814 & ~n10815;
  assign n10818 = ~n10813 & n10817;
  assign n10819 = ~n10816 & n10818;
  assign n10820 = pi38  & n10819;
  assign n10821 = ~pi38  & ~n10819;
  assign n10822 = ~n10820 & ~n10821;
  assign n10823 = ~n10572 & ~n10575;
  assign n10824 = pi82  & n5558;
  assign n10825 = pi83  & n5293;
  assign n10826 = pi84  & n5288;
  assign n10827 = n1601 & n5286;
  assign n10828 = ~n10825 & ~n10826;
  assign n10829 = ~n10824 & n10828;
  assign n10830 = ~n10827 & n10829;
  assign n10831 = pi41  & n10830;
  assign n10832 = ~pi41  & ~n10830;
  assign n10833 = ~n10831 & ~n10832;
  assign n10834 = ~n10556 & ~n10560;
  assign n10835 = pi79  & n6331;
  assign n10836 = pi80  & n6015;
  assign n10837 = pi81  & n6010;
  assign n10838 = n1337 & n6008;
  assign n10839 = ~n10836 & ~n10837;
  assign n10840 = ~n10835 & n10839;
  assign n10841 = ~n10838 & n10840;
  assign n10842 = pi44  & n10841;
  assign n10843 = ~pi44  & ~n10841;
  assign n10844 = ~n10842 & ~n10843;
  assign n10845 = ~n10540 & ~n10543;
  assign n10846 = ~n10524 & ~n10528;
  assign n10847 = pi73  & n7969;
  assign n10848 = pi74  & n7636;
  assign n10849 = pi75  & n7631;
  assign n10850 = n713 & n7629;
  assign n10851 = ~n10848 & ~n10849;
  assign n10852 = ~n10847 & n10851;
  assign n10853 = ~n10850 & n10852;
  assign n10854 = pi50  & n10853;
  assign n10855 = ~pi50  & ~n10853;
  assign n10856 = ~n10854 & ~n10855;
  assign n10857 = ~n10509 & ~n10511;
  assign n10858 = pi70  & n8905;
  assign n10859 = pi71  & n8535;
  assign n10860 = pi72  & n8530;
  assign n10861 = n551 & n8528;
  assign n10862 = ~n10859 & ~n10860;
  assign n10863 = ~n10858 & n10862;
  assign n10864 = ~n10861 & n10863;
  assign n10865 = pi53  & n10864;
  assign n10866 = ~pi53  & ~n10864;
  assign n10867 = ~n10865 & ~n10866;
  assign n10868 = ~n10503 & ~n10505;
  assign n10869 = pi67  & n9858;
  assign n10870 = pi68  & n9508;
  assign n10871 = pi69  & n9503;
  assign n10872 = n376 & n9501;
  assign n10873 = ~n10870 & ~n10871;
  assign n10874 = ~n10869 & n10873;
  assign n10875 = ~n10872 & n10874;
  assign n10876 = pi56  & n10875;
  assign n10877 = ~pi56  & ~n10875;
  assign n10878 = ~n10876 & ~n10877;
  assign n10879 = pi59  & ~n10219;
  assign n10880 = n10498 & n10879;
  assign n10881 = pi59  & ~n10880;
  assign n10882 = ~n287 & n10488;
  assign n10883 = pi65  & n10495;
  assign n10884 = pi66  & n10490;
  assign n10885 = ~n10218 & n10487;
  assign n10886 = ~n10494 & n10885;
  assign n10887 = pi64  & n10886;
  assign n10888 = ~n10882 & ~n10883;
  assign n10889 = ~n10884 & n10888;
  assign n10890 = ~n10887 & n10889;
  assign n10891 = ~n10881 & n10890;
  assign n10892 = n10881 & ~n10890;
  assign n10893 = ~n10891 & ~n10892;
  assign n10894 = ~n10878 & n10893;
  assign n10895 = n10878 & ~n10893;
  assign n10896 = ~n10894 & ~n10895;
  assign n10897 = ~n10868 & n10896;
  assign n10898 = n10868 & ~n10896;
  assign n10899 = ~n10897 & ~n10898;
  assign n10900 = n10867 & ~n10899;
  assign n10901 = ~n10867 & n10899;
  assign n10902 = ~n10900 & ~n10901;
  assign n10903 = ~n10857 & n10902;
  assign n10904 = n10857 & ~n10902;
  assign n10905 = ~n10903 & ~n10904;
  assign n10906 = n10856 & ~n10905;
  assign n10907 = ~n10856 & n10905;
  assign n10908 = ~n10906 & ~n10907;
  assign n10909 = ~n10846 & n10908;
  assign n10910 = n10846 & ~n10908;
  assign n10911 = ~n10909 & ~n10910;
  assign n10912 = pi76  & n7121;
  assign n10913 = pi77  & n6795;
  assign n10914 = pi78  & n6790;
  assign n10915 = n958 & n6788;
  assign n10916 = ~n10913 & ~n10914;
  assign n10917 = ~n10912 & n10916;
  assign n10918 = ~n10915 & n10917;
  assign n10919 = pi47  & n10918;
  assign n10920 = ~pi47  & ~n10918;
  assign n10921 = ~n10919 & ~n10920;
  assign n10922 = n10911 & ~n10921;
  assign n10923 = ~n10911 & n10921;
  assign n10924 = ~n10922 & ~n10923;
  assign n10925 = ~n10845 & n10924;
  assign n10926 = n10845 & ~n10924;
  assign n10927 = ~n10925 & ~n10926;
  assign n10928 = ~n10844 & n10927;
  assign n10929 = n10844 & ~n10927;
  assign n10930 = ~n10928 & ~n10929;
  assign n10931 = ~n10834 & n10930;
  assign n10932 = n10834 & ~n10930;
  assign n10933 = ~n10931 & ~n10932;
  assign n10934 = ~n10833 & n10933;
  assign n10935 = n10833 & ~n10933;
  assign n10936 = ~n10934 & ~n10935;
  assign n10937 = ~n10823 & n10936;
  assign n10938 = n10823 & ~n10936;
  assign n10939 = ~n10937 & ~n10938;
  assign n10940 = ~n10822 & n10939;
  assign n10941 = n10822 & ~n10939;
  assign n10942 = ~n10940 & ~n10941;
  assign n10943 = n10812 & ~n10942;
  assign n10944 = ~n10812 & n10942;
  assign n10945 = ~n10943 & ~n10944;
  assign n10946 = pi88  & n4176;
  assign n10947 = pi89  & n3938;
  assign n10948 = pi90  & n3933;
  assign n10949 = n2448 & n3931;
  assign n10950 = ~n10947 & ~n10948;
  assign n10951 = ~n10946 & n10950;
  assign n10952 = ~n10949 & n10951;
  assign n10953 = pi35  & n10952;
  assign n10954 = ~pi35  & ~n10952;
  assign n10955 = ~n10953 & ~n10954;
  assign n10956 = n10945 & ~n10955;
  assign n10957 = ~n10945 & n10955;
  assign n10958 = ~n10956 & ~n10957;
  assign n10959 = n10811 & ~n10958;
  assign n10960 = ~n10811 & n10958;
  assign n10961 = ~n10959 & ~n10960;
  assign n10962 = pi91  & n3553;
  assign n10963 = pi92  & n3334;
  assign n10964 = pi93  & n3329;
  assign n10965 = n2948 & n3327;
  assign n10966 = ~n10963 & ~n10964;
  assign n10967 = ~n10962 & n10966;
  assign n10968 = ~n10965 & n10967;
  assign n10969 = pi32  & n10968;
  assign n10970 = ~pi32  & ~n10968;
  assign n10971 = ~n10969 & ~n10970;
  assign n10972 = n10961 & ~n10971;
  assign n10973 = ~n10961 & n10971;
  assign n10974 = ~n10972 & ~n10973;
  assign n10975 = ~n10810 & n10974;
  assign n10976 = n10810 & ~n10974;
  assign n10977 = ~n10975 & ~n10976;
  assign n10978 = n10809 & ~n10977;
  assign n10979 = ~n10809 & n10977;
  assign n10980 = ~n10978 & ~n10979;
  assign n10981 = ~n10799 & n10980;
  assign n10982 = n10799 & ~n10980;
  assign n10983 = ~n10981 & ~n10982;
  assign n10984 = pi97  & n2510;
  assign n10985 = pi98  & n2342;
  assign n10986 = pi99  & n2337;
  assign n10987 = n2335 & n4101;
  assign n10988 = ~n10985 & ~n10986;
  assign n10989 = ~n10984 & n10988;
  assign n10990 = ~n10987 & n10989;
  assign n10991 = pi26  & n10990;
  assign n10992 = ~pi26  & ~n10990;
  assign n10993 = ~n10991 & ~n10992;
  assign n10994 = n10983 & ~n10993;
  assign n10995 = ~n10983 & n10993;
  assign n10996 = ~n10994 & ~n10995;
  assign n10997 = n10798 & ~n10996;
  assign n10998 = ~n10798 & n10996;
  assign n10999 = ~n10997 & ~n10998;
  assign n11000 = pi100  & n2053;
  assign n11001 = pi101  & n1893;
  assign n11002 = pi102  & n1888;
  assign n11003 = n1886 & n4956;
  assign n11004 = ~n11001 & ~n11002;
  assign n11005 = ~n11000 & n11004;
  assign n11006 = ~n11003 & n11005;
  assign n11007 = pi23  & n11006;
  assign n11008 = ~pi23  & ~n11006;
  assign n11009 = ~n11007 & ~n11008;
  assign n11010 = n10999 & ~n11009;
  assign n11011 = ~n10999 & n11009;
  assign n11012 = ~n11010 & ~n11011;
  assign n11013 = n10797 & ~n11012;
  assign n11014 = ~n10797 & n11012;
  assign n11015 = ~n11013 & ~n11014;
  assign n11016 = pi103  & n1661;
  assign n11017 = pi104  & n1500;
  assign n11018 = pi105  & n1495;
  assign n11019 = n1493 & n5677;
  assign n11020 = ~n11017 & ~n11018;
  assign n11021 = ~n11016 & n11020;
  assign n11022 = ~n11019 & n11021;
  assign n11023 = pi20  & n11022;
  assign n11024 = ~pi20  & ~n11022;
  assign n11025 = ~n11023 & ~n11024;
  assign n11026 = n11015 & ~n11025;
  assign n11027 = ~n11015 & n11025;
  assign n11028 = ~n11026 & ~n11027;
  assign n11029 = ~n10796 & n11028;
  assign n11030 = n10796 & ~n11028;
  assign n11031 = ~n11029 & ~n11030;
  assign n11032 = pi106  & n1296;
  assign n11033 = pi107  & n1207;
  assign n11034 = pi108  & n1202;
  assign n11035 = n1200 & n6213;
  assign n11036 = ~n11033 & ~n11034;
  assign n11037 = ~n11032 & n11036;
  assign n11038 = ~n11035 & n11037;
  assign n11039 = pi17  & n11038;
  assign n11040 = ~pi17  & ~n11038;
  assign n11041 = ~n11039 & ~n11040;
  assign n11042 = n11031 & ~n11041;
  assign n11043 = ~n11031 & n11041;
  assign n11044 = ~n11042 & ~n11043;
  assign n11045 = ~n10795 & n11044;
  assign n11046 = n10795 & ~n11044;
  assign n11047 = ~n11045 & ~n11046;
  assign n11048 = ~n10794 & n11047;
  assign n11049 = n10794 & ~n11047;
  assign n11050 = ~n11048 & ~n11049;
  assign n11051 = ~n10784 & n11050;
  assign n11052 = n10784 & ~n11050;
  assign n11053 = ~n11051 & ~n11052;
  assign n11054 = pi112  & n750;
  assign n11055 = pi113  & n651;
  assign n11056 = pi114  & n646;
  assign n11057 = n644 & n8146;
  assign n11058 = ~n11055 & ~n11056;
  assign n11059 = ~n11054 & n11058;
  assign n11060 = ~n11057 & n11059;
  assign n11061 = pi11  & n11060;
  assign n11062 = ~pi11  & ~n11060;
  assign n11063 = ~n11061 & ~n11062;
  assign n11064 = n11053 & ~n11063;
  assign n11065 = ~n11053 & n11063;
  assign n11066 = ~n11064 & ~n11065;
  assign n11067 = ~n10783 & n11066;
  assign n11068 = n10783 & ~n11066;
  assign n11069 = ~n11067 & ~n11068;
  assign n11070 = ~n10782 & n11069;
  assign n11071 = n10782 & ~n11069;
  assign n11072 = ~n11070 & ~n11071;
  assign n11073 = ~n10772 & n11072;
  assign n11074 = n10772 & ~n11072;
  assign n11075 = ~n11073 & ~n11074;
  assign n11076 = ~n10771 & n11075;
  assign n11077 = n10771 & ~n11075;
  assign n11078 = ~n11076 & ~n11077;
  assign n11079 = ~n10761 & n11078;
  assign n11080 = n10761 & ~n11078;
  assign n11081 = ~n11079 & ~n11080;
  assign n11082 = ~n10744 & n11081;
  assign n11083 = n10744 & ~n11081;
  assign n11084 = ~n11082 & ~n11083;
  assign n11085 = ~n10743 & n11084;
  assign n11086 = n10743 & ~n11084;
  assign po59  = ~n11085 & ~n11086;
  assign n11088 = ~n11082 & ~n11085;
  assign n11089 = ~n11076 & ~n11079;
  assign n11090 = pi124  & n269;
  assign n11091 = pi123  & n267;
  assign n11092 = pi122  & n282;
  assign n11093 = ~n10750 & ~n10752;
  assign n11094 = ~pi123  & ~pi124 ;
  assign n11095 = pi123  & pi124 ;
  assign n11096 = ~n11094 & ~n11095;
  assign n11097 = ~n11093 & n11096;
  assign n11098 = n11093 & ~n11096;
  assign n11099 = ~n11097 & ~n11098;
  assign n11100 = n262 & n11099;
  assign n11101 = ~n11090 & ~n11091;
  assign n11102 = ~n11092 & n11101;
  assign n11103 = ~n11100 & n11102;
  assign n11104 = pi2  & n11103;
  assign n11105 = ~pi2  & ~n11103;
  assign n11106 = ~n11104 & ~n11105;
  assign n11107 = pi119  & n391;
  assign n11108 = pi120  & n353;
  assign n11109 = pi121  & n348;
  assign n11110 = n346 & n10071;
  assign n11111 = ~n11108 & ~n11109;
  assign n11112 = ~n11107 & n11111;
  assign n11113 = ~n11110 & n11112;
  assign n11114 = pi5  & n11113;
  assign n11115 = ~pi5  & ~n11113;
  assign n11116 = ~n11114 & ~n11115;
  assign n11117 = ~n11070 & ~n11073;
  assign n11118 = pi116  & n528;
  assign n11119 = pi117  & n490;
  assign n11120 = pi118  & n485;
  assign n11121 = n483 & n9095;
  assign n11122 = ~n11119 & ~n11120;
  assign n11123 = ~n11118 & n11122;
  assign n11124 = ~n11121 & n11123;
  assign n11125 = pi8  & n11124;
  assign n11126 = ~pi8  & ~n11124;
  assign n11127 = ~n11125 & ~n11126;
  assign n11128 = ~n11064 & ~n11067;
  assign n11129 = pi113  & n750;
  assign n11130 = pi114  & n651;
  assign n11131 = pi115  & n646;
  assign n11132 = n644 & n8170;
  assign n11133 = ~n11130 & ~n11131;
  assign n11134 = ~n11129 & n11133;
  assign n11135 = ~n11132 & n11134;
  assign n11136 = pi11  & n11135;
  assign n11137 = ~pi11  & ~n11135;
  assign n11138 = ~n11136 & ~n11137;
  assign n11139 = ~n11048 & ~n11051;
  assign n11140 = pi110  & n1006;
  assign n11141 = pi111  & n897;
  assign n11142 = pi112  & n892;
  assign n11143 = n890 & n7296;
  assign n11144 = ~n11141 & ~n11142;
  assign n11145 = ~n11140 & n11144;
  assign n11146 = ~n11143 & n11145;
  assign n11147 = pi14  & n11146;
  assign n11148 = ~pi14  & ~n11146;
  assign n11149 = ~n11147 & ~n11148;
  assign n11150 = ~n11042 & ~n11045;
  assign n11151 = pi107  & n1296;
  assign n11152 = pi108  & n1207;
  assign n11153 = pi109  & n1202;
  assign n11154 = n1200 & n6715;
  assign n11155 = ~n11152 & ~n11153;
  assign n11156 = ~n11151 & n11155;
  assign n11157 = ~n11154 & n11156;
  assign n11158 = pi17  & n11157;
  assign n11159 = ~pi17  & ~n11157;
  assign n11160 = ~n11158 & ~n11159;
  assign n11161 = ~n11026 & ~n11029;
  assign n11162 = ~n11010 & ~n11014;
  assign n11163 = ~n10994 & ~n10998;
  assign n11164 = pi98  & n2510;
  assign n11165 = pi99  & n2342;
  assign n11166 = pi100  & n2337;
  assign n11167 = n2335 & n4501;
  assign n11168 = ~n11165 & ~n11166;
  assign n11169 = ~n11164 & n11168;
  assign n11170 = ~n11167 & n11169;
  assign n11171 = pi26  & n11170;
  assign n11172 = ~pi26  & ~n11170;
  assign n11173 = ~n11171 & ~n11172;
  assign n11174 = ~n10979 & ~n10981;
  assign n11175 = ~n10972 & ~n10975;
  assign n11176 = ~n10956 & ~n10960;
  assign n11177 = ~n10940 & ~n10944;
  assign n11178 = ~n10934 & ~n10937;
  assign n11179 = pi83  & n5558;
  assign n11180 = pi84  & n5293;
  assign n11181 = pi85  & n5288;
  assign n11182 = n1831 & n5286;
  assign n11183 = ~n11180 & ~n11181;
  assign n11184 = ~n11179 & n11183;
  assign n11185 = ~n11182 & n11184;
  assign n11186 = pi41  & n11185;
  assign n11187 = ~pi41  & ~n11185;
  assign n11188 = ~n11186 & ~n11187;
  assign n11189 = ~n10928 & ~n10931;
  assign n11190 = pi80  & n6331;
  assign n11191 = pi81  & n6015;
  assign n11192 = pi82  & n6010;
  assign n11193 = n1450 & n6008;
  assign n11194 = ~n11191 & ~n11192;
  assign n11195 = ~n11190 & n11194;
  assign n11196 = ~n11193 & n11195;
  assign n11197 = pi44  & n11196;
  assign n11198 = ~pi44  & ~n11196;
  assign n11199 = ~n11197 & ~n11198;
  assign n11200 = ~n10922 & ~n10925;
  assign n11201 = pi77  & n7121;
  assign n11202 = pi78  & n6795;
  assign n11203 = pi79  & n6790;
  assign n11204 = n1048 & n6788;
  assign n11205 = ~n11202 & ~n11203;
  assign n11206 = ~n11201 & n11205;
  assign n11207 = ~n11204 & n11206;
  assign n11208 = pi47  & n11207;
  assign n11209 = ~pi47  & ~n11207;
  assign n11210 = ~n11208 & ~n11209;
  assign n11211 = ~n10907 & ~n10909;
  assign n11212 = pi74  & n7969;
  assign n11213 = pi75  & n7636;
  assign n11214 = pi76  & n7631;
  assign n11215 = n841 & n7629;
  assign n11216 = ~n11213 & ~n11214;
  assign n11217 = ~n11212 & n11216;
  assign n11218 = ~n11215 & n11217;
  assign n11219 = pi50  & n11218;
  assign n11220 = ~pi50  & ~n11218;
  assign n11221 = ~n11219 & ~n11220;
  assign n11222 = ~n10901 & ~n10903;
  assign n11223 = pi71  & n8905;
  assign n11224 = pi72  & n8535;
  assign n11225 = pi73  & n8530;
  assign n11226 = n613 & n8528;
  assign n11227 = ~n11224 & ~n11225;
  assign n11228 = ~n11223 & n11227;
  assign n11229 = ~n11226 & n11228;
  assign n11230 = pi53  & n11229;
  assign n11231 = ~pi53  & ~n11229;
  assign n11232 = ~n11230 & ~n11231;
  assign n11233 = ~n10894 & ~n10897;
  assign n11234 = pi65  & n10886;
  assign n11235 = pi66  & n10495;
  assign n11236 = pi67  & n10490;
  assign n11237 = n305 & n10488;
  assign n11238 = ~n11235 & ~n11236;
  assign n11239 = ~n11234 & n11238;
  assign n11240 = ~n11237 & n11239;
  assign n11241 = pi59  & n11240;
  assign n11242 = ~pi59  & ~n11240;
  assign n11243 = ~n11241 & ~n11242;
  assign n11244 = ~pi59  & ~pi60 ;
  assign n11245 = pi59  & pi60 ;
  assign n11246 = ~n11244 & ~n11245;
  assign n11247 = pi64  & n11246;
  assign n11248 = n10880 & n10890;
  assign n11249 = n11247 & n11248;
  assign n11250 = ~n11247 & ~n11248;
  assign n11251 = ~n11249 & ~n11250;
  assign n11252 = ~n11243 & n11251;
  assign n11253 = n11243 & ~n11251;
  assign n11254 = ~n11252 & ~n11253;
  assign n11255 = pi68  & n9858;
  assign n11256 = pi69  & n9508;
  assign n11257 = pi70  & n9503;
  assign n11258 = n415 & n9501;
  assign n11259 = ~n11256 & ~n11257;
  assign n11260 = ~n11255 & n11259;
  assign n11261 = ~n11258 & n11260;
  assign n11262 = pi56  & n11261;
  assign n11263 = ~pi56  & ~n11261;
  assign n11264 = ~n11262 & ~n11263;
  assign n11265 = n11254 & ~n11264;
  assign n11266 = ~n11254 & n11264;
  assign n11267 = ~n11265 & ~n11266;
  assign n11268 = ~n11233 & n11267;
  assign n11269 = n11233 & ~n11267;
  assign n11270 = ~n11268 & ~n11269;
  assign n11271 = ~n11232 & n11270;
  assign n11272 = n11232 & ~n11270;
  assign n11273 = ~n11271 & ~n11272;
  assign n11274 = ~n11222 & n11273;
  assign n11275 = n11222 & ~n11273;
  assign n11276 = ~n11274 & ~n11275;
  assign n11277 = n11221 & ~n11276;
  assign n11278 = ~n11221 & n11276;
  assign n11279 = ~n11277 & ~n11278;
  assign n11280 = ~n11211 & n11279;
  assign n11281 = n11211 & ~n11279;
  assign n11282 = ~n11280 & ~n11281;
  assign n11283 = ~n11210 & n11282;
  assign n11284 = n11210 & ~n11282;
  assign n11285 = ~n11283 & ~n11284;
  assign n11286 = ~n11200 & n11285;
  assign n11287 = n11200 & ~n11285;
  assign n11288 = ~n11286 & ~n11287;
  assign n11289 = ~n11199 & n11288;
  assign n11290 = n11199 & ~n11288;
  assign n11291 = ~n11289 & ~n11290;
  assign n11292 = ~n11189 & n11291;
  assign n11293 = n11189 & ~n11291;
  assign n11294 = ~n11292 & ~n11293;
  assign n11295 = ~n11188 & n11294;
  assign n11296 = n11188 & ~n11294;
  assign n11297 = ~n11295 & ~n11296;
  assign n11298 = ~n11178 & n11297;
  assign n11299 = n11178 & ~n11297;
  assign n11300 = ~n11298 & ~n11299;
  assign n11301 = pi86  & n4843;
  assign n11302 = pi87  & n4598;
  assign n11303 = pi88  & n4593;
  assign n11304 = n2140 & n4591;
  assign n11305 = ~n11302 & ~n11303;
  assign n11306 = ~n11301 & n11305;
  assign n11307 = ~n11304 & n11306;
  assign n11308 = pi38  & n11307;
  assign n11309 = ~pi38  & ~n11307;
  assign n11310 = ~n11308 & ~n11309;
  assign n11311 = n11300 & ~n11310;
  assign n11312 = ~n11300 & n11310;
  assign n11313 = ~n11311 & ~n11312;
  assign n11314 = n11177 & ~n11313;
  assign n11315 = ~n11177 & n11313;
  assign n11316 = ~n11314 & ~n11315;
  assign n11317 = pi89  & n4176;
  assign n11318 = pi90  & n3938;
  assign n11319 = pi91  & n3933;
  assign n11320 = n2746 & n3931;
  assign n11321 = ~n11318 & ~n11319;
  assign n11322 = ~n11317 & n11321;
  assign n11323 = ~n11320 & n11322;
  assign n11324 = pi35  & n11323;
  assign n11325 = ~pi35  & ~n11323;
  assign n11326 = ~n11324 & ~n11325;
  assign n11327 = n11316 & ~n11326;
  assign n11328 = ~n11316 & n11326;
  assign n11329 = ~n11327 & ~n11328;
  assign n11330 = n11176 & ~n11329;
  assign n11331 = ~n11176 & n11329;
  assign n11332 = ~n11330 & ~n11331;
  assign n11333 = pi92  & n3553;
  assign n11334 = pi93  & n3334;
  assign n11335 = pi94  & n3329;
  assign n11336 = n3280 & n3327;
  assign n11337 = ~n11334 & ~n11335;
  assign n11338 = ~n11333 & n11337;
  assign n11339 = ~n11336 & n11338;
  assign n11340 = pi32  & n11339;
  assign n11341 = ~pi32  & ~n11339;
  assign n11342 = ~n11340 & ~n11341;
  assign n11343 = ~n11332 & n11342;
  assign n11344 = n11332 & ~n11342;
  assign n11345 = ~n11343 & ~n11344;
  assign n11346 = ~n11175 & n11345;
  assign n11347 = n11175 & ~n11345;
  assign n11348 = ~n11346 & ~n11347;
  assign n11349 = pi95  & n3011;
  assign n11350 = pi96  & n2809;
  assign n11351 = pi97  & n2804;
  assign n11352 = n2802 & n3691;
  assign n11353 = ~n11350 & ~n11351;
  assign n11354 = ~n11349 & n11353;
  assign n11355 = ~n11352 & n11354;
  assign n11356 = pi29  & n11355;
  assign n11357 = ~pi29  & ~n11355;
  assign n11358 = ~n11356 & ~n11357;
  assign n11359 = n11348 & ~n11358;
  assign n11360 = ~n11348 & n11358;
  assign n11361 = ~n11359 & ~n11360;
  assign n11362 = ~n11174 & n11361;
  assign n11363 = n11174 & ~n11361;
  assign n11364 = ~n11362 & ~n11363;
  assign n11365 = ~n11173 & n11364;
  assign n11366 = n11173 & ~n11364;
  assign n11367 = ~n11365 & ~n11366;
  assign n11368 = n11163 & ~n11367;
  assign n11369 = ~n11163 & n11367;
  assign n11370 = ~n11368 & ~n11369;
  assign n11371 = pi101  & n2053;
  assign n11372 = pi102  & n1893;
  assign n11373 = pi103  & n1888;
  assign n11374 = n1886 & n5188;
  assign n11375 = ~n11372 & ~n11373;
  assign n11376 = ~n11371 & n11375;
  assign n11377 = ~n11374 & n11376;
  assign n11378 = pi23  & n11377;
  assign n11379 = ~pi23  & ~n11377;
  assign n11380 = ~n11378 & ~n11379;
  assign n11381 = n11370 & ~n11380;
  assign n11382 = ~n11370 & n11380;
  assign n11383 = ~n11381 & ~n11382;
  assign n11384 = n11162 & ~n11383;
  assign n11385 = ~n11162 & n11383;
  assign n11386 = ~n11384 & ~n11385;
  assign n11387 = pi104  & n1661;
  assign n11388 = pi105  & n1500;
  assign n11389 = pi106  & n1495;
  assign n11390 = n1493 & n5701;
  assign n11391 = ~n11388 & ~n11389;
  assign n11392 = ~n11387 & n11391;
  assign n11393 = ~n11390 & n11392;
  assign n11394 = pi20  & n11393;
  assign n11395 = ~pi20  & ~n11393;
  assign n11396 = ~n11394 & ~n11395;
  assign n11397 = ~n11386 & n11396;
  assign n11398 = n11386 & ~n11396;
  assign n11399 = ~n11397 & ~n11398;
  assign n11400 = ~n11161 & n11399;
  assign n11401 = n11161 & ~n11399;
  assign n11402 = ~n11400 & ~n11401;
  assign n11403 = ~n11160 & n11402;
  assign n11404 = n11160 & ~n11402;
  assign n11405 = ~n11403 & ~n11404;
  assign n11406 = ~n11150 & n11405;
  assign n11407 = n11150 & ~n11405;
  assign n11408 = ~n11406 & ~n11407;
  assign n11409 = ~n11149 & n11408;
  assign n11410 = n11149 & ~n11408;
  assign n11411 = ~n11409 & ~n11410;
  assign n11412 = ~n11139 & n11411;
  assign n11413 = n11139 & ~n11411;
  assign n11414 = ~n11412 & ~n11413;
  assign n11415 = ~n11138 & n11414;
  assign n11416 = n11138 & ~n11414;
  assign n11417 = ~n11415 & ~n11416;
  assign n11418 = ~n11128 & n11417;
  assign n11419 = n11128 & ~n11417;
  assign n11420 = ~n11418 & ~n11419;
  assign n11421 = ~n11127 & n11420;
  assign n11422 = n11127 & ~n11420;
  assign n11423 = ~n11421 & ~n11422;
  assign n11424 = ~n11117 & n11423;
  assign n11425 = n11117 & ~n11423;
  assign n11426 = ~n11424 & ~n11425;
  assign n11427 = ~n11116 & n11426;
  assign n11428 = n11116 & ~n11426;
  assign n11429 = ~n11427 & ~n11428;
  assign n11430 = ~n11106 & n11429;
  assign n11431 = n11106 & ~n11429;
  assign n11432 = ~n11430 & ~n11431;
  assign n11433 = ~n11089 & n11432;
  assign n11434 = n11089 & ~n11432;
  assign n11435 = ~n11433 & ~n11434;
  assign n11436 = ~n11088 & n11435;
  assign n11437 = n11088 & ~n11435;
  assign po60  = ~n11436 & ~n11437;
  assign n11439 = ~n11427 & ~n11430;
  assign n11440 = ~n11421 & ~n11424;
  assign n11441 = ~n11415 & ~n11418;
  assign n11442 = pi114  & n750;
  assign n11443 = pi115  & n651;
  assign n11444 = pi116  & n646;
  assign n11445 = n644 & n8470;
  assign n11446 = ~n11443 & ~n11444;
  assign n11447 = ~n11442 & n11446;
  assign n11448 = ~n11445 & n11447;
  assign n11449 = pi11  & n11448;
  assign n11450 = ~pi11  & ~n11448;
  assign n11451 = ~n11449 & ~n11450;
  assign n11452 = ~n11409 & ~n11412;
  assign n11453 = pi111  & n1006;
  assign n11454 = pi112  & n897;
  assign n11455 = pi113  & n892;
  assign n11456 = n890 & n7852;
  assign n11457 = ~n11454 & ~n11455;
  assign n11458 = ~n11453 & n11457;
  assign n11459 = ~n11456 & n11458;
  assign n11460 = pi14  & n11459;
  assign n11461 = ~pi14  & ~n11459;
  assign n11462 = ~n11460 & ~n11461;
  assign n11463 = ~n11403 & ~n11406;
  assign n11464 = pi108  & n1296;
  assign n11465 = pi109  & n1207;
  assign n11466 = pi110  & n1202;
  assign n11467 = n1200 & n6995;
  assign n11468 = ~n11465 & ~n11466;
  assign n11469 = ~n11464 & n11468;
  assign n11470 = ~n11467 & n11469;
  assign n11471 = pi17  & n11470;
  assign n11472 = ~pi17  & ~n11470;
  assign n11473 = ~n11471 & ~n11472;
  assign n11474 = ~n11398 & ~n11400;
  assign n11475 = ~n11381 & ~n11385;
  assign n11476 = ~n11365 & ~n11369;
  assign n11477 = ~n11359 & ~n11362;
  assign n11478 = pi96  & n3011;
  assign n11479 = pi97  & n2809;
  assign n11480 = pi98  & n2804;
  assign n11481 = n2802 & n3889;
  assign n11482 = ~n11479 & ~n11480;
  assign n11483 = ~n11478 & n11482;
  assign n11484 = ~n11481 & n11483;
  assign n11485 = pi29  & n11484;
  assign n11486 = ~pi29  & ~n11484;
  assign n11487 = ~n11485 & ~n11486;
  assign n11488 = ~n11344 & ~n11346;
  assign n11489 = ~n11327 & ~n11331;
  assign n11490 = ~n11311 & ~n11315;
  assign n11491 = ~n11295 & ~n11298;
  assign n11492 = ~n11289 & ~n11292;
  assign n11493 = ~n11283 & ~n11286;
  assign n11494 = ~n11278 & ~n11280;
  assign n11495 = ~n11271 & ~n11274;
  assign n11496 = ~n11265 & ~n11268;
  assign n11497 = pi69  & n9858;
  assign n11498 = pi70  & n9508;
  assign n11499 = pi71  & n9503;
  assign n11500 = n460 & n9501;
  assign n11501 = ~n11498 & ~n11499;
  assign n11502 = ~n11497 & n11501;
  assign n11503 = ~n11500 & n11502;
  assign n11504 = pi56  & n11503;
  assign n11505 = ~pi56  & ~n11503;
  assign n11506 = ~n11504 & ~n11505;
  assign n11507 = ~n11249 & ~n11252;
  assign n11508 = pi66  & n10886;
  assign n11509 = pi67  & n10495;
  assign n11510 = pi68  & n10490;
  assign n11511 = n334 & n10488;
  assign n11512 = ~n11509 & ~n11510;
  assign n11513 = ~n11508 & n11512;
  assign n11514 = ~n11511 & n11513;
  assign n11515 = pi59  & n11514;
  assign n11516 = ~pi59  & ~n11514;
  assign n11517 = ~n11515 & ~n11516;
  assign n11518 = pi62  & n11247;
  assign n11519 = ~pi61  & ~pi62 ;
  assign n11520 = pi61  & pi62 ;
  assign n11521 = ~n11519 & ~n11520;
  assign n11522 = n11246 & n11521;
  assign n11523 = n265 & n11522;
  assign n11524 = n11246 & ~n11521;
  assign n11525 = pi65  & n11524;
  assign n11526 = ~pi60  & ~pi61 ;
  assign n11527 = pi60  & pi61 ;
  assign n11528 = ~n11526 & ~n11527;
  assign n11529 = ~n11246 & n11528;
  assign n11530 = pi64  & n11529;
  assign n11531 = ~n11523 & ~n11525;
  assign n11532 = ~n11530 & n11531;
  assign n11533 = n11518 & ~n11532;
  assign n11534 = ~n11518 & n11532;
  assign n11535 = ~n11533 & ~n11534;
  assign n11536 = n11517 & ~n11535;
  assign n11537 = ~n11517 & n11535;
  assign n11538 = ~n11536 & ~n11537;
  assign n11539 = ~n11507 & n11538;
  assign n11540 = n11507 & ~n11538;
  assign n11541 = ~n11539 & ~n11540;
  assign n11542 = n11506 & ~n11541;
  assign n11543 = ~n11506 & n11541;
  assign n11544 = ~n11542 & ~n11543;
  assign n11545 = ~n11496 & n11544;
  assign n11546 = n11496 & ~n11544;
  assign n11547 = ~n11545 & ~n11546;
  assign n11548 = pi72  & n8905;
  assign n11549 = pi73  & n8535;
  assign n11550 = pi74  & n8530;
  assign n11551 = n689 & n8528;
  assign n11552 = ~n11549 & ~n11550;
  assign n11553 = ~n11548 & n11552;
  assign n11554 = ~n11551 & n11553;
  assign n11555 = pi53  & n11554;
  assign n11556 = ~pi53  & ~n11554;
  assign n11557 = ~n11555 & ~n11556;
  assign n11558 = n11547 & ~n11557;
  assign n11559 = ~n11547 & n11557;
  assign n11560 = ~n11558 & ~n11559;
  assign n11561 = n11495 & ~n11560;
  assign n11562 = ~n11495 & n11560;
  assign n11563 = ~n11561 & ~n11562;
  assign n11564 = pi75  & n7969;
  assign n11565 = pi76  & n7636;
  assign n11566 = pi77  & n7631;
  assign n11567 = n865 & n7629;
  assign n11568 = ~n11565 & ~n11566;
  assign n11569 = ~n11564 & n11568;
  assign n11570 = ~n11567 & n11569;
  assign n11571 = pi50  & n11570;
  assign n11572 = ~pi50  & ~n11570;
  assign n11573 = ~n11571 & ~n11572;
  assign n11574 = n11563 & ~n11573;
  assign n11575 = ~n11563 & n11573;
  assign n11576 = ~n11574 & ~n11575;
  assign n11577 = ~n11494 & n11576;
  assign n11578 = n11494 & ~n11576;
  assign n11579 = ~n11577 & ~n11578;
  assign n11580 = pi78  & n7121;
  assign n11581 = pi79  & n6795;
  assign n11582 = pi80  & n6790;
  assign n11583 = n1144 & n6788;
  assign n11584 = ~n11581 & ~n11582;
  assign n11585 = ~n11580 & n11584;
  assign n11586 = ~n11583 & n11585;
  assign n11587 = pi47  & n11586;
  assign n11588 = ~pi47  & ~n11586;
  assign n11589 = ~n11587 & ~n11588;
  assign n11590 = n11579 & ~n11589;
  assign n11591 = ~n11579 & n11589;
  assign n11592 = ~n11590 & ~n11591;
  assign n11593 = n11493 & ~n11592;
  assign n11594 = ~n11493 & n11592;
  assign n11595 = ~n11593 & ~n11594;
  assign n11596 = pi81  & n6331;
  assign n11597 = pi82  & n6015;
  assign n11598 = pi83  & n6010;
  assign n11599 = n1577 & n6008;
  assign n11600 = ~n11597 & ~n11598;
  assign n11601 = ~n11596 & n11600;
  assign n11602 = ~n11599 & n11601;
  assign n11603 = pi44  & n11602;
  assign n11604 = ~pi44  & ~n11602;
  assign n11605 = ~n11603 & ~n11604;
  assign n11606 = n11595 & ~n11605;
  assign n11607 = ~n11595 & n11605;
  assign n11608 = ~n11606 & ~n11607;
  assign n11609 = ~n11492 & n11608;
  assign n11610 = n11492 & ~n11608;
  assign n11611 = ~n11609 & ~n11610;
  assign n11612 = pi84  & n5558;
  assign n11613 = pi85  & n5293;
  assign n11614 = pi86  & n5288;
  assign n11615 = n1975 & n5286;
  assign n11616 = ~n11613 & ~n11614;
  assign n11617 = ~n11612 & n11616;
  assign n11618 = ~n11615 & n11617;
  assign n11619 = pi41  & n11618;
  assign n11620 = ~pi41  & ~n11618;
  assign n11621 = ~n11619 & ~n11620;
  assign n11622 = n11611 & ~n11621;
  assign n11623 = ~n11611 & n11621;
  assign n11624 = ~n11622 & ~n11623;
  assign n11625 = n11491 & ~n11624;
  assign n11626 = ~n11491 & n11624;
  assign n11627 = ~n11625 & ~n11626;
  assign n11628 = pi87  & n4843;
  assign n11629 = pi88  & n4598;
  assign n11630 = pi89  & n4593;
  assign n11631 = n2287 & n4591;
  assign n11632 = ~n11629 & ~n11630;
  assign n11633 = ~n11628 & n11632;
  assign n11634 = ~n11631 & n11633;
  assign n11635 = pi38  & n11634;
  assign n11636 = ~pi38  & ~n11634;
  assign n11637 = ~n11635 & ~n11636;
  assign n11638 = n11627 & ~n11637;
  assign n11639 = ~n11627 & n11637;
  assign n11640 = ~n11638 & ~n11639;
  assign n11641 = n11490 & ~n11640;
  assign n11642 = ~n11490 & n11640;
  assign n11643 = ~n11641 & ~n11642;
  assign n11644 = pi90  & n4176;
  assign n11645 = pi91  & n3938;
  assign n11646 = pi92  & n3933;
  assign n11647 = n2924 & n3931;
  assign n11648 = ~n11645 & ~n11646;
  assign n11649 = ~n11644 & n11648;
  assign n11650 = ~n11647 & n11649;
  assign n11651 = pi35  & n11650;
  assign n11652 = ~pi35  & ~n11650;
  assign n11653 = ~n11651 & ~n11652;
  assign n11654 = n11643 & ~n11653;
  assign n11655 = ~n11643 & n11653;
  assign n11656 = ~n11654 & ~n11655;
  assign n11657 = n11489 & ~n11656;
  assign n11658 = ~n11489 & n11656;
  assign n11659 = ~n11657 & ~n11658;
  assign n11660 = pi93  & n3553;
  assign n11661 = pi94  & n3334;
  assign n11662 = pi95  & n3329;
  assign n11663 = n3327 & n3475;
  assign n11664 = ~n11661 & ~n11662;
  assign n11665 = ~n11660 & n11664;
  assign n11666 = ~n11663 & n11665;
  assign n11667 = pi32  & n11666;
  assign n11668 = ~pi32  & ~n11666;
  assign n11669 = ~n11667 & ~n11668;
  assign n11670 = n11659 & ~n11669;
  assign n11671 = ~n11659 & n11669;
  assign n11672 = ~n11670 & ~n11671;
  assign n11673 = ~n11488 & n11672;
  assign n11674 = n11488 & ~n11672;
  assign n11675 = ~n11673 & ~n11674;
  assign n11676 = ~n11487 & n11675;
  assign n11677 = n11487 & ~n11675;
  assign n11678 = ~n11676 & ~n11677;
  assign n11679 = n11477 & ~n11678;
  assign n11680 = ~n11477 & n11678;
  assign n11681 = ~n11679 & ~n11680;
  assign n11682 = pi99  & n2510;
  assign n11683 = pi100  & n2342;
  assign n11684 = pi101  & n2337;
  assign n11685 = n2335 & n4730;
  assign n11686 = ~n11683 & ~n11684;
  assign n11687 = ~n11682 & n11686;
  assign n11688 = ~n11685 & n11687;
  assign n11689 = pi26  & n11688;
  assign n11690 = ~pi26  & ~n11688;
  assign n11691 = ~n11689 & ~n11690;
  assign n11692 = n11681 & ~n11691;
  assign n11693 = ~n11681 & n11691;
  assign n11694 = ~n11692 & ~n11693;
  assign n11695 = n11476 & ~n11694;
  assign n11696 = ~n11476 & n11694;
  assign n11697 = ~n11695 & ~n11696;
  assign n11698 = pi102  & n2053;
  assign n11699 = pi103  & n1893;
  assign n11700 = pi104  & n1888;
  assign n11701 = n1886 & n5212;
  assign n11702 = ~n11699 & ~n11700;
  assign n11703 = ~n11698 & n11702;
  assign n11704 = ~n11701 & n11703;
  assign n11705 = pi23  & n11704;
  assign n11706 = ~pi23  & ~n11704;
  assign n11707 = ~n11705 & ~n11706;
  assign n11708 = n11697 & ~n11707;
  assign n11709 = ~n11697 & n11707;
  assign n11710 = ~n11708 & ~n11709;
  assign n11711 = n11475 & ~n11710;
  assign n11712 = ~n11475 & n11710;
  assign n11713 = ~n11711 & ~n11712;
  assign n11714 = pi105  & n1661;
  assign n11715 = pi106  & n1500;
  assign n11716 = pi107  & n1495;
  assign n11717 = n1493 & n6189;
  assign n11718 = ~n11715 & ~n11716;
  assign n11719 = ~n11714 & n11718;
  assign n11720 = ~n11717 & n11719;
  assign n11721 = pi20  & n11720;
  assign n11722 = ~pi20  & ~n11720;
  assign n11723 = ~n11721 & ~n11722;
  assign n11724 = n11713 & ~n11723;
  assign n11725 = ~n11713 & n11723;
  assign n11726 = ~n11724 & ~n11725;
  assign n11727 = ~n11474 & n11726;
  assign n11728 = n11474 & ~n11726;
  assign n11729 = ~n11727 & ~n11728;
  assign n11730 = n11473 & ~n11729;
  assign n11731 = ~n11473 & n11729;
  assign n11732 = ~n11730 & ~n11731;
  assign n11733 = ~n11463 & n11732;
  assign n11734 = n11463 & ~n11732;
  assign n11735 = ~n11733 & ~n11734;
  assign n11736 = n11462 & ~n11735;
  assign n11737 = ~n11462 & n11735;
  assign n11738 = ~n11736 & ~n11737;
  assign n11739 = ~n11452 & n11738;
  assign n11740 = n11452 & ~n11738;
  assign n11741 = ~n11739 & ~n11740;
  assign n11742 = n11451 & ~n11741;
  assign n11743 = ~n11451 & n11741;
  assign n11744 = ~n11742 & ~n11743;
  assign n11745 = ~n11441 & n11744;
  assign n11746 = n11441 & ~n11744;
  assign n11747 = ~n11745 & ~n11746;
  assign n11748 = pi117  & n528;
  assign n11749 = pi118  & n490;
  assign n11750 = pi119  & n485;
  assign n11751 = n483 & n9412;
  assign n11752 = ~n11749 & ~n11750;
  assign n11753 = ~n11748 & n11752;
  assign n11754 = ~n11751 & n11753;
  assign n11755 = pi8  & n11754;
  assign n11756 = ~pi8  & ~n11754;
  assign n11757 = ~n11755 & ~n11756;
  assign n11758 = n11747 & ~n11757;
  assign n11759 = ~n11747 & n11757;
  assign n11760 = ~n11758 & ~n11759;
  assign n11761 = n11440 & ~n11760;
  assign n11762 = ~n11440 & n11760;
  assign n11763 = ~n11761 & ~n11762;
  assign n11764 = pi120  & n391;
  assign n11765 = pi121  & n353;
  assign n11766 = pi122  & n348;
  assign n11767 = n346 & n10729;
  assign n11768 = ~n11765 & ~n11766;
  assign n11769 = ~n11764 & n11768;
  assign n11770 = ~n11767 & n11769;
  assign n11771 = pi5  & n11770;
  assign n11772 = ~pi5  & ~n11770;
  assign n11773 = ~n11771 & ~n11772;
  assign n11774 = ~n11763 & n11773;
  assign n11775 = n11763 & ~n11773;
  assign n11776 = ~n11774 & ~n11775;
  assign n11777 = pi125  & n269;
  assign n11778 = pi124  & n267;
  assign n11779 = pi123  & n282;
  assign n11780 = ~n11095 & ~n11097;
  assign n11781 = ~pi124  & ~pi125 ;
  assign n11782 = pi124  & pi125 ;
  assign n11783 = ~n11781 & ~n11782;
  assign n11784 = ~n11780 & n11783;
  assign n11785 = n11780 & ~n11783;
  assign n11786 = ~n11784 & ~n11785;
  assign n11787 = n262 & n11786;
  assign n11788 = ~n11777 & ~n11778;
  assign n11789 = ~n11779 & n11788;
  assign n11790 = ~n11787 & n11789;
  assign n11791 = pi2  & n11790;
  assign n11792 = ~pi2  & ~n11790;
  assign n11793 = ~n11791 & ~n11792;
  assign n11794 = n11776 & ~n11793;
  assign n11795 = ~n11776 & n11793;
  assign n11796 = ~n11794 & ~n11795;
  assign n11797 = n11439 & ~n11796;
  assign n11798 = ~n11439 & n11796;
  assign n11799 = ~n11797 & ~n11798;
  assign n11800 = ~n11433 & ~n11436;
  assign n11801 = n11799 & ~n11800;
  assign n11802 = ~n11799 & n11800;
  assign po61  = ~n11801 & ~n11802;
  assign n11804 = ~n11798 & ~n11801;
  assign n11805 = ~n11758 & ~n11762;
  assign n11806 = ~n11743 & ~n11745;
  assign n11807 = pi115  & n750;
  assign n11808 = pi116  & n651;
  assign n11809 = pi117  & n646;
  assign n11810 = n644 & n8784;
  assign n11811 = ~n11808 & ~n11809;
  assign n11812 = ~n11807 & n11811;
  assign n11813 = ~n11810 & n11812;
  assign n11814 = pi11  & n11813;
  assign n11815 = ~pi11  & ~n11813;
  assign n11816 = ~n11814 & ~n11815;
  assign n11817 = ~n11737 & ~n11739;
  assign n11818 = ~n11731 & ~n11733;
  assign n11819 = pi109  & n1296;
  assign n11820 = pi110  & n1207;
  assign n11821 = pi111  & n1202;
  assign n11822 = n1200 & n7272;
  assign n11823 = ~n11820 & ~n11821;
  assign n11824 = ~n11819 & n11823;
  assign n11825 = ~n11822 & n11824;
  assign n11826 = pi17  & n11825;
  assign n11827 = ~pi17  & ~n11825;
  assign n11828 = ~n11826 & ~n11827;
  assign n11829 = ~n11724 & ~n11727;
  assign n11830 = ~n11708 & ~n11712;
  assign n11831 = ~n11692 & ~n11696;
  assign n11832 = ~n11676 & ~n11680;
  assign n11833 = ~n11670 & ~n11673;
  assign n11834 = ~n11654 & ~n11658;
  assign n11835 = ~n11638 & ~n11642;
  assign n11836 = ~n11622 & ~n11626;
  assign n11837 = pi85  & n5558;
  assign n11838 = pi86  & n5293;
  assign n11839 = pi87  & n5288;
  assign n11840 = n2116 & n5286;
  assign n11841 = ~n11838 & ~n11839;
  assign n11842 = ~n11837 & n11841;
  assign n11843 = ~n11840 & n11842;
  assign n11844 = pi41  & n11843;
  assign n11845 = ~pi41  & ~n11843;
  assign n11846 = ~n11844 & ~n11845;
  assign n11847 = ~n11606 & ~n11609;
  assign n11848 = pi82  & n6331;
  assign n11849 = pi83  & n6015;
  assign n11850 = pi84  & n6010;
  assign n11851 = n1601 & n6008;
  assign n11852 = ~n11849 & ~n11850;
  assign n11853 = ~n11848 & n11852;
  assign n11854 = ~n11851 & n11853;
  assign n11855 = pi44  & n11854;
  assign n11856 = ~pi44  & ~n11854;
  assign n11857 = ~n11855 & ~n11856;
  assign n11858 = ~n11590 & ~n11594;
  assign n11859 = pi79  & n7121;
  assign n11860 = pi80  & n6795;
  assign n11861 = pi81  & n6790;
  assign n11862 = n1337 & n6788;
  assign n11863 = ~n11860 & ~n11861;
  assign n11864 = ~n11859 & n11863;
  assign n11865 = ~n11862 & n11864;
  assign n11866 = pi47  & n11865;
  assign n11867 = ~pi47  & ~n11865;
  assign n11868 = ~n11866 & ~n11867;
  assign n11869 = ~n11574 & ~n11577;
  assign n11870 = ~n11558 & ~n11562;
  assign n11871 = pi73  & n8905;
  assign n11872 = pi74  & n8535;
  assign n11873 = pi75  & n8530;
  assign n11874 = n713 & n8528;
  assign n11875 = ~n11872 & ~n11873;
  assign n11876 = ~n11871 & n11875;
  assign n11877 = ~n11874 & n11876;
  assign n11878 = pi53  & n11877;
  assign n11879 = ~pi53  & ~n11877;
  assign n11880 = ~n11878 & ~n11879;
  assign n11881 = ~n11543 & ~n11545;
  assign n11882 = pi70  & n9858;
  assign n11883 = pi71  & n9508;
  assign n11884 = pi72  & n9503;
  assign n11885 = n551 & n9501;
  assign n11886 = ~n11883 & ~n11884;
  assign n11887 = ~n11882 & n11886;
  assign n11888 = ~n11885 & n11887;
  assign n11889 = pi56  & n11888;
  assign n11890 = ~pi56  & ~n11888;
  assign n11891 = ~n11889 & ~n11890;
  assign n11892 = ~n11537 & ~n11539;
  assign n11893 = pi67  & n10886;
  assign n11894 = pi68  & n10495;
  assign n11895 = pi69  & n10490;
  assign n11896 = n376 & n10488;
  assign n11897 = ~n11894 & ~n11895;
  assign n11898 = ~n11893 & n11897;
  assign n11899 = ~n11896 & n11898;
  assign n11900 = pi59  & n11899;
  assign n11901 = ~pi59  & ~n11899;
  assign n11902 = ~n11900 & ~n11901;
  assign n11903 = pi62  & ~n11247;
  assign n11904 = n11532 & n11903;
  assign n11905 = pi62  & ~n11904;
  assign n11906 = ~n287 & n11522;
  assign n11907 = pi65  & n11529;
  assign n11908 = pi66  & n11524;
  assign n11909 = ~n11246 & n11521;
  assign n11910 = ~n11528 & n11909;
  assign n11911 = pi64  & n11910;
  assign n11912 = ~n11906 & ~n11907;
  assign n11913 = ~n11908 & n11912;
  assign n11914 = ~n11911 & n11913;
  assign n11915 = ~n11905 & n11914;
  assign n11916 = n11905 & ~n11914;
  assign n11917 = ~n11915 & ~n11916;
  assign n11918 = ~n11902 & n11917;
  assign n11919 = n11902 & ~n11917;
  assign n11920 = ~n11918 & ~n11919;
  assign n11921 = ~n11892 & n11920;
  assign n11922 = n11892 & ~n11920;
  assign n11923 = ~n11921 & ~n11922;
  assign n11924 = n11891 & ~n11923;
  assign n11925 = ~n11891 & n11923;
  assign n11926 = ~n11924 & ~n11925;
  assign n11927 = ~n11881 & n11926;
  assign n11928 = n11881 & ~n11926;
  assign n11929 = ~n11927 & ~n11928;
  assign n11930 = n11880 & ~n11929;
  assign n11931 = ~n11880 & n11929;
  assign n11932 = ~n11930 & ~n11931;
  assign n11933 = ~n11870 & n11932;
  assign n11934 = n11870 & ~n11932;
  assign n11935 = ~n11933 & ~n11934;
  assign n11936 = pi76  & n7969;
  assign n11937 = pi77  & n7636;
  assign n11938 = pi78  & n7631;
  assign n11939 = n958 & n7629;
  assign n11940 = ~n11937 & ~n11938;
  assign n11941 = ~n11936 & n11940;
  assign n11942 = ~n11939 & n11941;
  assign n11943 = pi50  & n11942;
  assign n11944 = ~pi50  & ~n11942;
  assign n11945 = ~n11943 & ~n11944;
  assign n11946 = n11935 & ~n11945;
  assign n11947 = ~n11935 & n11945;
  assign n11948 = ~n11946 & ~n11947;
  assign n11949 = ~n11869 & n11948;
  assign n11950 = n11869 & ~n11948;
  assign n11951 = ~n11949 & ~n11950;
  assign n11952 = ~n11868 & n11951;
  assign n11953 = n11868 & ~n11951;
  assign n11954 = ~n11952 & ~n11953;
  assign n11955 = ~n11858 & n11954;
  assign n11956 = n11858 & ~n11954;
  assign n11957 = ~n11955 & ~n11956;
  assign n11958 = ~n11857 & n11957;
  assign n11959 = n11857 & ~n11957;
  assign n11960 = ~n11958 & ~n11959;
  assign n11961 = ~n11847 & n11960;
  assign n11962 = n11847 & ~n11960;
  assign n11963 = ~n11961 & ~n11962;
  assign n11964 = ~n11846 & n11963;
  assign n11965 = n11846 & ~n11963;
  assign n11966 = ~n11964 & ~n11965;
  assign n11967 = n11836 & ~n11966;
  assign n11968 = ~n11836 & n11966;
  assign n11969 = ~n11967 & ~n11968;
  assign n11970 = pi88  & n4843;
  assign n11971 = pi89  & n4598;
  assign n11972 = pi90  & n4593;
  assign n11973 = n2448 & n4591;
  assign n11974 = ~n11971 & ~n11972;
  assign n11975 = ~n11970 & n11974;
  assign n11976 = ~n11973 & n11975;
  assign n11977 = pi38  & n11976;
  assign n11978 = ~pi38  & ~n11976;
  assign n11979 = ~n11977 & ~n11978;
  assign n11980 = n11969 & ~n11979;
  assign n11981 = ~n11969 & n11979;
  assign n11982 = ~n11980 & ~n11981;
  assign n11983 = n11835 & ~n11982;
  assign n11984 = ~n11835 & n11982;
  assign n11985 = ~n11983 & ~n11984;
  assign n11986 = pi91  & n4176;
  assign n11987 = pi92  & n3938;
  assign n11988 = pi93  & n3933;
  assign n11989 = n2948 & n3931;
  assign n11990 = ~n11987 & ~n11988;
  assign n11991 = ~n11986 & n11990;
  assign n11992 = ~n11989 & n11991;
  assign n11993 = pi35  & n11992;
  assign n11994 = ~pi35  & ~n11992;
  assign n11995 = ~n11993 & ~n11994;
  assign n11996 = n11985 & ~n11995;
  assign n11997 = ~n11985 & n11995;
  assign n11998 = ~n11996 & ~n11997;
  assign n11999 = n11834 & ~n11998;
  assign n12000 = ~n11834 & n11998;
  assign n12001 = ~n11999 & ~n12000;
  assign n12002 = pi94  & n3553;
  assign n12003 = pi95  & n3334;
  assign n12004 = pi96  & n3329;
  assign n12005 = n3327 & n3499;
  assign n12006 = ~n12003 & ~n12004;
  assign n12007 = ~n12002 & n12006;
  assign n12008 = ~n12005 & n12007;
  assign n12009 = pi32  & n12008;
  assign n12010 = ~pi32  & ~n12008;
  assign n12011 = ~n12009 & ~n12010;
  assign n12012 = n12001 & ~n12011;
  assign n12013 = ~n12001 & n12011;
  assign n12014 = ~n12012 & ~n12013;
  assign n12015 = ~n11833 & n12014;
  assign n12016 = n11833 & ~n12014;
  assign n12017 = ~n12015 & ~n12016;
  assign n12018 = pi97  & n3011;
  assign n12019 = pi98  & n2809;
  assign n12020 = pi99  & n2804;
  assign n12021 = n2802 & n4101;
  assign n12022 = ~n12019 & ~n12020;
  assign n12023 = ~n12018 & n12022;
  assign n12024 = ~n12021 & n12023;
  assign n12025 = pi29  & n12024;
  assign n12026 = ~pi29  & ~n12024;
  assign n12027 = ~n12025 & ~n12026;
  assign n12028 = n12017 & ~n12027;
  assign n12029 = ~n12017 & n12027;
  assign n12030 = ~n12028 & ~n12029;
  assign n12031 = n11832 & ~n12030;
  assign n12032 = ~n11832 & n12030;
  assign n12033 = ~n12031 & ~n12032;
  assign n12034 = pi100  & n2510;
  assign n12035 = pi101  & n2342;
  assign n12036 = pi102  & n2337;
  assign n12037 = n2335 & n4956;
  assign n12038 = ~n12035 & ~n12036;
  assign n12039 = ~n12034 & n12038;
  assign n12040 = ~n12037 & n12039;
  assign n12041 = pi26  & n12040;
  assign n12042 = ~pi26  & ~n12040;
  assign n12043 = ~n12041 & ~n12042;
  assign n12044 = n12033 & ~n12043;
  assign n12045 = ~n12033 & n12043;
  assign n12046 = ~n12044 & ~n12045;
  assign n12047 = n11831 & ~n12046;
  assign n12048 = ~n11831 & n12046;
  assign n12049 = ~n12047 & ~n12048;
  assign n12050 = pi103  & n2053;
  assign n12051 = pi104  & n1893;
  assign n12052 = pi105  & n1888;
  assign n12053 = n1886 & n5677;
  assign n12054 = ~n12051 & ~n12052;
  assign n12055 = ~n12050 & n12054;
  assign n12056 = ~n12053 & n12055;
  assign n12057 = pi23  & n12056;
  assign n12058 = ~pi23  & ~n12056;
  assign n12059 = ~n12057 & ~n12058;
  assign n12060 = n12049 & ~n12059;
  assign n12061 = ~n12049 & n12059;
  assign n12062 = ~n12060 & ~n12061;
  assign n12063 = ~n11830 & n12062;
  assign n12064 = n11830 & ~n12062;
  assign n12065 = ~n12063 & ~n12064;
  assign n12066 = pi106  & n1661;
  assign n12067 = pi107  & n1500;
  assign n12068 = pi108  & n1495;
  assign n12069 = n1493 & n6213;
  assign n12070 = ~n12067 & ~n12068;
  assign n12071 = ~n12066 & n12070;
  assign n12072 = ~n12069 & n12071;
  assign n12073 = pi20  & n12072;
  assign n12074 = ~pi20  & ~n12072;
  assign n12075 = ~n12073 & ~n12074;
  assign n12076 = n12065 & ~n12075;
  assign n12077 = ~n12065 & n12075;
  assign n12078 = ~n12076 & ~n12077;
  assign n12079 = ~n11829 & n12078;
  assign n12080 = n11829 & ~n12078;
  assign n12081 = ~n12079 & ~n12080;
  assign n12082 = ~n11828 & n12081;
  assign n12083 = n11828 & ~n12081;
  assign n12084 = ~n12082 & ~n12083;
  assign n12085 = ~n11818 & n12084;
  assign n12086 = n11818 & ~n12084;
  assign n12087 = ~n12085 & ~n12086;
  assign n12088 = pi112  & n1006;
  assign n12089 = pi113  & n897;
  assign n12090 = pi114  & n892;
  assign n12091 = n890 & n8146;
  assign n12092 = ~n12089 & ~n12090;
  assign n12093 = ~n12088 & n12092;
  assign n12094 = ~n12091 & n12093;
  assign n12095 = pi14  & n12094;
  assign n12096 = ~pi14  & ~n12094;
  assign n12097 = ~n12095 & ~n12096;
  assign n12098 = n12087 & ~n12097;
  assign n12099 = ~n12087 & n12097;
  assign n12100 = ~n12098 & ~n12099;
  assign n12101 = ~n11817 & n12100;
  assign n12102 = n11817 & ~n12100;
  assign n12103 = ~n12101 & ~n12102;
  assign n12104 = ~n11816 & n12103;
  assign n12105 = n11816 & ~n12103;
  assign n12106 = ~n12104 & ~n12105;
  assign n12107 = ~n11806 & n12106;
  assign n12108 = n11806 & ~n12106;
  assign n12109 = ~n12107 & ~n12108;
  assign n12110 = pi118  & n528;
  assign n12111 = pi119  & n490;
  assign n12112 = pi120  & n485;
  assign n12113 = n483 & n10047;
  assign n12114 = ~n12111 & ~n12112;
  assign n12115 = ~n12110 & n12114;
  assign n12116 = ~n12113 & n12115;
  assign n12117 = pi8  & n12116;
  assign n12118 = ~pi8  & ~n12116;
  assign n12119 = ~n12117 & ~n12118;
  assign n12120 = ~n12109 & n12119;
  assign n12121 = n12109 & ~n12119;
  assign n12122 = ~n12120 & ~n12121;
  assign n12123 = pi121  & n391;
  assign n12124 = pi122  & n353;
  assign n12125 = pi123  & n348;
  assign n12126 = n346 & n10754;
  assign n12127 = ~n12124 & ~n12125;
  assign n12128 = ~n12123 & n12127;
  assign n12129 = ~n12126 & n12128;
  assign n12130 = pi5  & n12129;
  assign n12131 = ~pi5  & ~n12129;
  assign n12132 = ~n12130 & ~n12131;
  assign n12133 = n12122 & ~n12132;
  assign n12134 = ~n12122 & n12132;
  assign n12135 = ~n12133 & ~n12134;
  assign n12136 = n11805 & ~n12135;
  assign n12137 = ~n11805 & n12135;
  assign n12138 = ~n12136 & ~n12137;
  assign n12139 = pi126  & n269;
  assign n12140 = pi125  & n267;
  assign n12141 = pi124  & n282;
  assign n12142 = ~n11782 & ~n11784;
  assign n12143 = ~pi125  & ~pi126 ;
  assign n12144 = pi125  & pi126 ;
  assign n12145 = ~n12143 & ~n12144;
  assign n12146 = ~n12142 & n12145;
  assign n12147 = n12142 & ~n12145;
  assign n12148 = ~n12146 & ~n12147;
  assign n12149 = n262 & n12148;
  assign n12150 = ~n12139 & ~n12140;
  assign n12151 = ~n12141 & n12150;
  assign n12152 = ~n12149 & n12151;
  assign n12153 = pi2  & n12152;
  assign n12154 = ~pi2  & ~n12152;
  assign n12155 = ~n12153 & ~n12154;
  assign n12156 = ~n12138 & n12155;
  assign n12157 = n12138 & ~n12155;
  assign n12158 = ~n12156 & ~n12157;
  assign n12159 = ~n11774 & ~n11793;
  assign n12160 = ~n11775 & ~n12159;
  assign n12161 = n12158 & ~n12160;
  assign n12162 = ~n12158 & n12160;
  assign n12163 = ~n12161 & ~n12162;
  assign n12164 = ~n11804 & n12163;
  assign n12165 = n11804 & ~n12163;
  assign po62  = ~n12164 & ~n12165;
  assign n12167 = ~n12161 & ~n12164;
  assign n12168 = ~n12137 & ~n12157;
  assign n12169 = pi122  & n391;
  assign n12170 = pi123  & n353;
  assign n12171 = pi124  & n348;
  assign n12172 = n346 & n11099;
  assign n12173 = ~n12170 & ~n12171;
  assign n12174 = ~n12169 & n12173;
  assign n12175 = ~n12172 & n12174;
  assign n12176 = pi5  & n12175;
  assign n12177 = ~pi5  & ~n12175;
  assign n12178 = ~n12176 & ~n12177;
  assign n12179 = ~n12104 & ~n12107;
  assign n12180 = ~n12098 & ~n12101;
  assign n12181 = pi113  & n1006;
  assign n12182 = pi114  & n897;
  assign n12183 = pi115  & n892;
  assign n12184 = n890 & n8170;
  assign n12185 = ~n12182 & ~n12183;
  assign n12186 = ~n12181 & n12185;
  assign n12187 = ~n12184 & n12186;
  assign n12188 = pi14  & n12187;
  assign n12189 = ~pi14  & ~n12187;
  assign n12190 = ~n12188 & ~n12189;
  assign n12191 = ~n12082 & ~n12085;
  assign n12192 = pi110  & n1296;
  assign n12193 = pi111  & n1207;
  assign n12194 = pi112  & n1202;
  assign n12195 = n1200 & n7296;
  assign n12196 = ~n12193 & ~n12194;
  assign n12197 = ~n12192 & n12196;
  assign n12198 = ~n12195 & n12197;
  assign n12199 = pi17  & n12198;
  assign n12200 = ~pi17  & ~n12198;
  assign n12201 = ~n12199 & ~n12200;
  assign n12202 = ~n12076 & ~n12079;
  assign n12203 = pi107  & n1661;
  assign n12204 = pi108  & n1500;
  assign n12205 = pi109  & n1495;
  assign n12206 = n1493 & n6715;
  assign n12207 = ~n12204 & ~n12205;
  assign n12208 = ~n12203 & n12207;
  assign n12209 = ~n12206 & n12208;
  assign n12210 = pi20  & n12209;
  assign n12211 = ~pi20  & ~n12209;
  assign n12212 = ~n12210 & ~n12211;
  assign n12213 = ~n12060 & ~n12063;
  assign n12214 = pi104  & n2053;
  assign n12215 = pi105  & n1893;
  assign n12216 = pi106  & n1888;
  assign n12217 = n1886 & n5701;
  assign n12218 = ~n12215 & ~n12216;
  assign n12219 = ~n12214 & n12218;
  assign n12220 = ~n12217 & n12219;
  assign n12221 = pi23  & n12220;
  assign n12222 = ~pi23  & ~n12220;
  assign n12223 = ~n12221 & ~n12222;
  assign n12224 = ~n12044 & ~n12048;
  assign n12225 = ~n12028 & ~n12032;
  assign n12226 = pi98  & n3011;
  assign n12227 = pi99  & n2809;
  assign n12228 = pi100  & n2804;
  assign n12229 = n2802 & n4501;
  assign n12230 = ~n12227 & ~n12228;
  assign n12231 = ~n12226 & n12230;
  assign n12232 = ~n12229 & n12231;
  assign n12233 = pi29  & n12232;
  assign n12234 = ~pi29  & ~n12232;
  assign n12235 = ~n12233 & ~n12234;
  assign n12236 = ~n12012 & ~n12015;
  assign n12237 = ~n11980 & ~n11984;
  assign n12238 = ~n11964 & ~n11968;
  assign n12239 = ~n11958 & ~n11961;
  assign n12240 = pi83  & n6331;
  assign n12241 = pi84  & n6015;
  assign n12242 = pi85  & n6010;
  assign n12243 = n1831 & n6008;
  assign n12244 = ~n12241 & ~n12242;
  assign n12245 = ~n12240 & n12244;
  assign n12246 = ~n12243 & n12245;
  assign n12247 = pi44  & n12246;
  assign n12248 = ~pi44  & ~n12246;
  assign n12249 = ~n12247 & ~n12248;
  assign n12250 = ~n11952 & ~n11955;
  assign n12251 = ~n11946 & ~n11949;
  assign n12252 = ~n11931 & ~n11933;
  assign n12253 = pi74  & n8905;
  assign n12254 = pi75  & n8535;
  assign n12255 = pi76  & n8530;
  assign n12256 = n841 & n8528;
  assign n12257 = ~n12254 & ~n12255;
  assign n12258 = ~n12253 & n12257;
  assign n12259 = ~n12256 & n12258;
  assign n12260 = pi53  & n12259;
  assign n12261 = ~pi53  & ~n12259;
  assign n12262 = ~n12260 & ~n12261;
  assign n12263 = ~n11925 & ~n11927;
  assign n12264 = ~n11918 & ~n11921;
  assign n12265 = pi68  & n10886;
  assign n12266 = pi69  & n10495;
  assign n12267 = pi70  & n10490;
  assign n12268 = n415 & n10488;
  assign n12269 = ~n12266 & ~n12267;
  assign n12270 = ~n12265 & n12269;
  assign n12271 = ~n12268 & n12270;
  assign n12272 = pi59  & n12271;
  assign n12273 = ~pi59  & ~n12271;
  assign n12274 = ~n12272 & ~n12273;
  assign n12275 = ~pi62  & ~pi63 ;
  assign n12276 = pi62  & pi63 ;
  assign n12277 = ~n12275 & ~n12276;
  assign n12278 = pi64  & n12277;
  assign n12279 = n11904 & n11914;
  assign n12280 = n12278 & n12279;
  assign n12281 = ~n12278 & ~n12279;
  assign n12282 = ~n12280 & ~n12281;
  assign n12283 = pi65  & n11910;
  assign n12284 = pi66  & n11529;
  assign n12285 = pi67  & n11524;
  assign n12286 = n305 & n11522;
  assign n12287 = ~n12284 & ~n12285;
  assign n12288 = ~n12283 & n12287;
  assign n12289 = ~n12286 & n12288;
  assign n12290 = pi62  & n12289;
  assign n12291 = ~pi62  & ~n12289;
  assign n12292 = ~n12290 & ~n12291;
  assign n12293 = n12282 & ~n12292;
  assign n12294 = ~n12282 & n12292;
  assign n12295 = ~n12293 & ~n12294;
  assign n12296 = n12274 & ~n12295;
  assign n12297 = ~n12274 & n12295;
  assign n12298 = ~n12296 & ~n12297;
  assign n12299 = ~n12264 & n12298;
  assign n12300 = n12264 & ~n12298;
  assign n12301 = ~n12299 & ~n12300;
  assign n12302 = pi71  & n9858;
  assign n12303 = pi72  & n9508;
  assign n12304 = pi73  & n9503;
  assign n12305 = n613 & n9501;
  assign n12306 = ~n12303 & ~n12304;
  assign n12307 = ~n12302 & n12306;
  assign n12308 = ~n12305 & n12307;
  assign n12309 = pi56  & n12308;
  assign n12310 = ~pi56  & ~n12308;
  assign n12311 = ~n12309 & ~n12310;
  assign n12312 = n12301 & ~n12311;
  assign n12313 = ~n12301 & n12311;
  assign n12314 = ~n12312 & ~n12313;
  assign n12315 = ~n12263 & n12314;
  assign n12316 = n12263 & ~n12314;
  assign n12317 = ~n12315 & ~n12316;
  assign n12318 = n12262 & ~n12317;
  assign n12319 = ~n12262 & n12317;
  assign n12320 = ~n12318 & ~n12319;
  assign n12321 = ~n12252 & n12320;
  assign n12322 = n12252 & ~n12320;
  assign n12323 = ~n12321 & ~n12322;
  assign n12324 = pi77  & n7969;
  assign n12325 = pi78  & n7636;
  assign n12326 = pi79  & n7631;
  assign n12327 = n1048 & n7629;
  assign n12328 = ~n12325 & ~n12326;
  assign n12329 = ~n12324 & n12328;
  assign n12330 = ~n12327 & n12329;
  assign n12331 = pi50  & n12330;
  assign n12332 = ~pi50  & ~n12330;
  assign n12333 = ~n12331 & ~n12332;
  assign n12334 = n12323 & ~n12333;
  assign n12335 = ~n12323 & n12333;
  assign n12336 = ~n12334 & ~n12335;
  assign n12337 = n12251 & ~n12336;
  assign n12338 = ~n12251 & n12336;
  assign n12339 = ~n12337 & ~n12338;
  assign n12340 = pi80  & n7121;
  assign n12341 = pi81  & n6795;
  assign n12342 = pi82  & n6790;
  assign n12343 = n1450 & n6788;
  assign n12344 = ~n12341 & ~n12342;
  assign n12345 = ~n12340 & n12344;
  assign n12346 = ~n12343 & n12345;
  assign n12347 = pi47  & n12346;
  assign n12348 = ~pi47  & ~n12346;
  assign n12349 = ~n12347 & ~n12348;
  assign n12350 = ~n12339 & n12349;
  assign n12351 = n12339 & ~n12349;
  assign n12352 = ~n12350 & ~n12351;
  assign n12353 = ~n12250 & n12352;
  assign n12354 = n12250 & ~n12352;
  assign n12355 = ~n12353 & ~n12354;
  assign n12356 = ~n12249 & n12355;
  assign n12357 = n12249 & ~n12355;
  assign n12358 = ~n12356 & ~n12357;
  assign n12359 = ~n12239 & n12358;
  assign n12360 = n12239 & ~n12358;
  assign n12361 = ~n12359 & ~n12360;
  assign n12362 = pi86  & n5558;
  assign n12363 = pi87  & n5293;
  assign n12364 = pi88  & n5288;
  assign n12365 = n2140 & n5286;
  assign n12366 = ~n12363 & ~n12364;
  assign n12367 = ~n12362 & n12366;
  assign n12368 = ~n12365 & n12367;
  assign n12369 = pi41  & n12368;
  assign n12370 = ~pi41  & ~n12368;
  assign n12371 = ~n12369 & ~n12370;
  assign n12372 = n12361 & ~n12371;
  assign n12373 = ~n12361 & n12371;
  assign n12374 = ~n12372 & ~n12373;
  assign n12375 = n12238 & ~n12374;
  assign n12376 = ~n12238 & n12374;
  assign n12377 = ~n12375 & ~n12376;
  assign n12378 = pi89  & n4843;
  assign n12379 = pi90  & n4598;
  assign n12380 = pi91  & n4593;
  assign n12381 = n2746 & n4591;
  assign n12382 = ~n12379 & ~n12380;
  assign n12383 = ~n12378 & n12382;
  assign n12384 = ~n12381 & n12383;
  assign n12385 = pi38  & n12384;
  assign n12386 = ~pi38  & ~n12384;
  assign n12387 = ~n12385 & ~n12386;
  assign n12388 = n12377 & ~n12387;
  assign n12389 = ~n12377 & n12387;
  assign n12390 = ~n12388 & ~n12389;
  assign n12391 = n12237 & ~n12390;
  assign n12392 = ~n12237 & n12390;
  assign n12393 = ~n12391 & ~n12392;
  assign n12394 = pi92  & n4176;
  assign n12395 = pi93  & n3938;
  assign n12396 = pi94  & n3933;
  assign n12397 = n3280 & n3931;
  assign n12398 = ~n12395 & ~n12396;
  assign n12399 = ~n12394 & n12398;
  assign n12400 = ~n12397 & n12399;
  assign n12401 = pi35  & n12400;
  assign n12402 = ~pi35  & ~n12400;
  assign n12403 = ~n12401 & ~n12402;
  assign n12404 = ~n12393 & n12403;
  assign n12405 = n12393 & ~n12403;
  assign n12406 = ~n12404 & ~n12405;
  assign n12407 = ~n11996 & ~n12000;
  assign n12408 = n12406 & ~n12407;
  assign n12409 = ~n12406 & n12407;
  assign n12410 = ~n12408 & ~n12409;
  assign n12411 = pi95  & n3553;
  assign n12412 = pi96  & n3334;
  assign n12413 = pi97  & n3329;
  assign n12414 = n3327 & n3691;
  assign n12415 = ~n12412 & ~n12413;
  assign n12416 = ~n12411 & n12415;
  assign n12417 = ~n12414 & n12416;
  assign n12418 = pi32  & n12417;
  assign n12419 = ~pi32  & ~n12417;
  assign n12420 = ~n12418 & ~n12419;
  assign n12421 = n12410 & ~n12420;
  assign n12422 = ~n12410 & n12420;
  assign n12423 = ~n12421 & ~n12422;
  assign n12424 = ~n12236 & n12423;
  assign n12425 = n12236 & ~n12423;
  assign n12426 = ~n12424 & ~n12425;
  assign n12427 = ~n12235 & n12426;
  assign n12428 = n12235 & ~n12426;
  assign n12429 = ~n12427 & ~n12428;
  assign n12430 = n12225 & ~n12429;
  assign n12431 = ~n12225 & n12429;
  assign n12432 = ~n12430 & ~n12431;
  assign n12433 = pi101  & n2510;
  assign n12434 = pi102  & n2342;
  assign n12435 = pi103  & n2337;
  assign n12436 = n2335 & n5188;
  assign n12437 = ~n12434 & ~n12435;
  assign n12438 = ~n12433 & n12437;
  assign n12439 = ~n12436 & n12438;
  assign n12440 = pi26  & n12439;
  assign n12441 = ~pi26  & ~n12439;
  assign n12442 = ~n12440 & ~n12441;
  assign n12443 = ~n12432 & n12442;
  assign n12444 = n12432 & ~n12442;
  assign n12445 = ~n12443 & ~n12444;
  assign n12446 = ~n12224 & n12445;
  assign n12447 = n12224 & ~n12445;
  assign n12448 = ~n12446 & ~n12447;
  assign n12449 = ~n12223 & n12448;
  assign n12450 = n12223 & ~n12448;
  assign n12451 = ~n12449 & ~n12450;
  assign n12452 = ~n12213 & n12451;
  assign n12453 = n12213 & ~n12451;
  assign n12454 = ~n12452 & ~n12453;
  assign n12455 = ~n12212 & n12454;
  assign n12456 = n12212 & ~n12454;
  assign n12457 = ~n12455 & ~n12456;
  assign n12458 = ~n12202 & n12457;
  assign n12459 = n12202 & ~n12457;
  assign n12460 = ~n12458 & ~n12459;
  assign n12461 = ~n12201 & n12460;
  assign n12462 = n12201 & ~n12460;
  assign n12463 = ~n12461 & ~n12462;
  assign n12464 = ~n12191 & n12463;
  assign n12465 = n12191 & ~n12463;
  assign n12466 = ~n12464 & ~n12465;
  assign n12467 = ~n12190 & n12466;
  assign n12468 = n12190 & ~n12466;
  assign n12469 = ~n12467 & ~n12468;
  assign n12470 = ~n12180 & n12469;
  assign n12471 = n12180 & ~n12469;
  assign n12472 = ~n12470 & ~n12471;
  assign n12473 = pi116  & n750;
  assign n12474 = pi117  & n651;
  assign n12475 = pi118  & n646;
  assign n12476 = n644 & n9095;
  assign n12477 = ~n12474 & ~n12475;
  assign n12478 = ~n12473 & n12477;
  assign n12479 = ~n12476 & n12478;
  assign n12480 = pi11  & n12479;
  assign n12481 = ~pi11  & ~n12479;
  assign n12482 = ~n12480 & ~n12481;
  assign n12483 = n12472 & ~n12482;
  assign n12484 = ~n12472 & n12482;
  assign n12485 = ~n12483 & ~n12484;
  assign n12486 = n12179 & ~n12485;
  assign n12487 = ~n12179 & n12485;
  assign n12488 = ~n12486 & ~n12487;
  assign n12489 = pi119  & n528;
  assign n12490 = pi120  & n490;
  assign n12491 = pi121  & n485;
  assign n12492 = n483 & n10071;
  assign n12493 = ~n12490 & ~n12491;
  assign n12494 = ~n12489 & n12493;
  assign n12495 = ~n12492 & n12494;
  assign n12496 = pi8  & n12495;
  assign n12497 = ~pi8  & ~n12495;
  assign n12498 = ~n12496 & ~n12497;
  assign n12499 = n12488 & ~n12498;
  assign n12500 = ~n12488 & n12498;
  assign n12501 = ~n12499 & ~n12500;
  assign n12502 = ~n12178 & n12501;
  assign n12503 = n12178 & ~n12501;
  assign n12504 = ~n12502 & ~n12503;
  assign n12505 = ~n12120 & ~n12132;
  assign n12506 = ~n12121 & ~n12505;
  assign n12507 = ~n12504 & n12506;
  assign n12508 = n12504 & ~n12506;
  assign n12509 = ~n12507 & ~n12508;
  assign n12510 = pi127  & n269;
  assign n12511 = pi126  & n267;
  assign n12512 = pi125  & n282;
  assign n12513 = ~n12144 & ~n12146;
  assign n12514 = ~pi126  & ~pi127 ;
  assign n12515 = pi126  & pi127 ;
  assign n12516 = ~n12514 & ~n12515;
  assign n12517 = n12513 & ~n12516;
  assign n12518 = ~n12513 & n12516;
  assign n12519 = ~n12517 & ~n12518;
  assign n12520 = n262 & n12519;
  assign n12521 = ~n12510 & ~n12511;
  assign n12522 = ~n12512 & n12521;
  assign n12523 = ~n12520 & n12522;
  assign n12524 = pi2  & n12523;
  assign n12525 = ~pi2  & ~n12523;
  assign n12526 = ~n12524 & ~n12525;
  assign n12527 = n12509 & ~n12526;
  assign n12528 = ~n12509 & n12526;
  assign n12529 = ~n12527 & ~n12528;
  assign n12530 = ~n12168 & n12529;
  assign n12531 = n12168 & ~n12529;
  assign n12532 = ~n12530 & ~n12531;
  assign n12533 = ~n12167 & n12532;
  assign n12534 = n12167 & ~n12532;
  assign po63  = ~n12533 & ~n12534;
  assign n12536 = ~n12530 & ~n12533;
  assign n12537 = pi126  & n282;
  assign n12538 = pi127  & n267;
  assign n12539 = ~pi126  & n12513;
  assign n12540 = pi126  & ~n12513;
  assign n12541 = ~n12539 & ~n12540;
  assign n12542 = n12516 & ~n12541;
  assign n12543 = n262 & n12542;
  assign n12544 = ~n12537 & ~n12538;
  assign n12545 = ~n12543 & n12544;
  assign n12546 = pi2  & n12545;
  assign n12547 = ~pi2  & ~n12545;
  assign n12548 = ~n12546 & ~n12547;
  assign n12549 = ~n12499 & ~n12502;
  assign n12550 = pi123  & n391;
  assign n12551 = pi124  & n353;
  assign n12552 = pi125  & n348;
  assign n12553 = n346 & n11786;
  assign n12554 = ~n12551 & ~n12552;
  assign n12555 = ~n12550 & n12554;
  assign n12556 = ~n12553 & n12555;
  assign n12557 = pi5  & n12556;
  assign n12558 = ~pi5  & ~n12556;
  assign n12559 = ~n12557 & ~n12558;
  assign n12560 = ~n12483 & ~n12487;
  assign n12561 = pi117  & n750;
  assign n12562 = pi118  & n651;
  assign n12563 = pi119  & n646;
  assign n12564 = n644 & n9412;
  assign n12565 = ~n12562 & ~n12563;
  assign n12566 = ~n12561 & n12565;
  assign n12567 = ~n12564 & n12566;
  assign n12568 = pi11  & n12567;
  assign n12569 = ~pi11  & ~n12567;
  assign n12570 = ~n12568 & ~n12569;
  assign n12571 = ~n12467 & ~n12470;
  assign n12572 = pi114  & n1006;
  assign n12573 = pi115  & n897;
  assign n12574 = pi116  & n892;
  assign n12575 = n890 & n8470;
  assign n12576 = ~n12573 & ~n12574;
  assign n12577 = ~n12572 & n12576;
  assign n12578 = ~n12575 & n12577;
  assign n12579 = pi14  & n12578;
  assign n12580 = ~pi14  & ~n12578;
  assign n12581 = ~n12579 & ~n12580;
  assign n12582 = ~n12461 & ~n12464;
  assign n12583 = pi111  & n1296;
  assign n12584 = pi112  & n1207;
  assign n12585 = pi113  & n1202;
  assign n12586 = n1200 & n7852;
  assign n12587 = ~n12584 & ~n12585;
  assign n12588 = ~n12583 & n12587;
  assign n12589 = ~n12586 & n12588;
  assign n12590 = pi17  & n12589;
  assign n12591 = ~pi17  & ~n12589;
  assign n12592 = ~n12590 & ~n12591;
  assign n12593 = ~n12455 & ~n12458;
  assign n12594 = pi108  & n1661;
  assign n12595 = pi109  & n1500;
  assign n12596 = pi110  & n1495;
  assign n12597 = n1493 & n6995;
  assign n12598 = ~n12595 & ~n12596;
  assign n12599 = ~n12594 & n12598;
  assign n12600 = ~n12597 & n12599;
  assign n12601 = pi20  & n12600;
  assign n12602 = ~pi20  & ~n12600;
  assign n12603 = ~n12601 & ~n12602;
  assign n12604 = ~n12449 & ~n12452;
  assign n12605 = pi105  & n2053;
  assign n12606 = pi106  & n1893;
  assign n12607 = pi107  & n1888;
  assign n12608 = n1886 & n6189;
  assign n12609 = ~n12606 & ~n12607;
  assign n12610 = ~n12605 & n12609;
  assign n12611 = ~n12608 & n12610;
  assign n12612 = pi23  & n12611;
  assign n12613 = ~pi23  & ~n12611;
  assign n12614 = ~n12612 & ~n12613;
  assign n12615 = ~n12444 & ~n12446;
  assign n12616 = ~n12427 & ~n12431;
  assign n12617 = ~n12421 & ~n12424;
  assign n12618 = ~n12388 & ~n12392;
  assign n12619 = ~n12372 & ~n12376;
  assign n12620 = ~n12356 & ~n12359;
  assign n12621 = ~n12334 & ~n12338;
  assign n12622 = ~n12312 & ~n12315;
  assign n12623 = ~n12297 & ~n12299;
  assign n12624 = pi66  & n11910;
  assign n12625 = pi67  & n11529;
  assign n12626 = pi68  & n11524;
  assign n12627 = n334 & n11522;
  assign n12628 = ~n12625 & ~n12626;
  assign n12629 = ~n12624 & n12628;
  assign n12630 = ~n12627 & n12629;
  assign n12631 = pi62  & n12630;
  assign n12632 = ~pi62  & ~n12630;
  assign n12633 = ~n12631 & ~n12632;
  assign n12634 = pi65  & n12277;
  assign n12635 = pi64  & n12276;
  assign n12636 = ~n12634 & ~n12635;
  assign n12637 = ~n12633 & ~n12636;
  assign n12638 = n12633 & n12636;
  assign n12639 = ~n12637 & ~n12638;
  assign n12640 = ~n12280 & n12292;
  assign n12641 = ~n12281 & ~n12640;
  assign n12642 = ~n12639 & ~n12641;
  assign n12643 = n12639 & n12641;
  assign n12644 = ~n12642 & ~n12643;
  assign n12645 = pi69  & n10886;
  assign n12646 = pi70  & n10495;
  assign n12647 = pi71  & n10490;
  assign n12648 = n460 & n10488;
  assign n12649 = ~n12646 & ~n12647;
  assign n12650 = ~n12645 & n12649;
  assign n12651 = ~n12648 & n12650;
  assign n12652 = pi59  & n12651;
  assign n12653 = ~pi59  & ~n12651;
  assign n12654 = ~n12652 & ~n12653;
  assign n12655 = ~n12644 & n12654;
  assign n12656 = n12644 & ~n12654;
  assign n12657 = ~n12655 & ~n12656;
  assign n12658 = ~n12623 & n12657;
  assign n12659 = n12623 & ~n12657;
  assign n12660 = ~n12658 & ~n12659;
  assign n12661 = pi72  & n9858;
  assign n12662 = pi73  & n9508;
  assign n12663 = pi74  & n9503;
  assign n12664 = n689 & n9501;
  assign n12665 = ~n12662 & ~n12663;
  assign n12666 = ~n12661 & n12665;
  assign n12667 = ~n12664 & n12666;
  assign n12668 = pi56  & n12667;
  assign n12669 = ~pi56  & ~n12667;
  assign n12670 = ~n12668 & ~n12669;
  assign n12671 = n12660 & ~n12670;
  assign n12672 = ~n12660 & n12670;
  assign n12673 = ~n12671 & ~n12672;
  assign n12674 = n12622 & ~n12673;
  assign n12675 = ~n12622 & n12673;
  assign n12676 = ~n12674 & ~n12675;
  assign n12677 = pi75  & n8905;
  assign n12678 = pi76  & n8535;
  assign n12679 = pi77  & n8530;
  assign n12680 = n865 & n8528;
  assign n12681 = ~n12678 & ~n12679;
  assign n12682 = ~n12677 & n12681;
  assign n12683 = ~n12680 & n12682;
  assign n12684 = pi53  & n12683;
  assign n12685 = ~pi53  & ~n12683;
  assign n12686 = ~n12684 & ~n12685;
  assign n12687 = ~n12676 & n12686;
  assign n12688 = n12676 & ~n12686;
  assign n12689 = ~n12687 & ~n12688;
  assign n12690 = ~n12319 & ~n12321;
  assign n12691 = n12689 & ~n12690;
  assign n12692 = ~n12689 & n12690;
  assign n12693 = ~n12691 & ~n12692;
  assign n12694 = pi78  & n7969;
  assign n12695 = pi79  & n7636;
  assign n12696 = pi80  & n7631;
  assign n12697 = n1144 & n7629;
  assign n12698 = ~n12695 & ~n12696;
  assign n12699 = ~n12694 & n12698;
  assign n12700 = ~n12697 & n12699;
  assign n12701 = pi50  & n12700;
  assign n12702 = ~pi50  & ~n12700;
  assign n12703 = ~n12701 & ~n12702;
  assign n12704 = n12693 & ~n12703;
  assign n12705 = ~n12693 & n12703;
  assign n12706 = ~n12704 & ~n12705;
  assign n12707 = n12621 & ~n12706;
  assign n12708 = ~n12621 & n12706;
  assign n12709 = ~n12707 & ~n12708;
  assign n12710 = pi81  & n7121;
  assign n12711 = pi82  & n6795;
  assign n12712 = pi83  & n6790;
  assign n12713 = n1577 & n6788;
  assign n12714 = ~n12711 & ~n12712;
  assign n12715 = ~n12710 & n12714;
  assign n12716 = ~n12713 & n12715;
  assign n12717 = pi47  & n12716;
  assign n12718 = ~pi47  & ~n12716;
  assign n12719 = ~n12717 & ~n12718;
  assign n12720 = ~n12709 & n12719;
  assign n12721 = n12709 & ~n12719;
  assign n12722 = ~n12720 & ~n12721;
  assign n12723 = ~n12351 & ~n12353;
  assign n12724 = n12722 & ~n12723;
  assign n12725 = ~n12722 & n12723;
  assign n12726 = ~n12724 & ~n12725;
  assign n12727 = pi84  & n6331;
  assign n12728 = pi85  & n6015;
  assign n12729 = pi86  & n6010;
  assign n12730 = n1975 & n6008;
  assign n12731 = ~n12728 & ~n12729;
  assign n12732 = ~n12727 & n12731;
  assign n12733 = ~n12730 & n12732;
  assign n12734 = pi44  & n12733;
  assign n12735 = ~pi44  & ~n12733;
  assign n12736 = ~n12734 & ~n12735;
  assign n12737 = n12726 & ~n12736;
  assign n12738 = ~n12726 & n12736;
  assign n12739 = ~n12737 & ~n12738;
  assign n12740 = n12620 & ~n12739;
  assign n12741 = ~n12620 & n12739;
  assign n12742 = ~n12740 & ~n12741;
  assign n12743 = pi87  & n5558;
  assign n12744 = pi88  & n5293;
  assign n12745 = pi89  & n5288;
  assign n12746 = n2287 & n5286;
  assign n12747 = ~n12744 & ~n12745;
  assign n12748 = ~n12743 & n12747;
  assign n12749 = ~n12746 & n12748;
  assign n12750 = pi41  & n12749;
  assign n12751 = ~pi41  & ~n12749;
  assign n12752 = ~n12750 & ~n12751;
  assign n12753 = n12742 & ~n12752;
  assign n12754 = ~n12742 & n12752;
  assign n12755 = ~n12753 & ~n12754;
  assign n12756 = n12619 & ~n12755;
  assign n12757 = ~n12619 & n12755;
  assign n12758 = ~n12756 & ~n12757;
  assign n12759 = pi90  & n4843;
  assign n12760 = pi91  & n4598;
  assign n12761 = pi92  & n4593;
  assign n12762 = n2924 & n4591;
  assign n12763 = ~n12760 & ~n12761;
  assign n12764 = ~n12759 & n12763;
  assign n12765 = ~n12762 & n12764;
  assign n12766 = pi38  & n12765;
  assign n12767 = ~pi38  & ~n12765;
  assign n12768 = ~n12766 & ~n12767;
  assign n12769 = n12758 & ~n12768;
  assign n12770 = ~n12758 & n12768;
  assign n12771 = ~n12769 & ~n12770;
  assign n12772 = n12618 & ~n12771;
  assign n12773 = ~n12618 & n12771;
  assign n12774 = ~n12772 & ~n12773;
  assign n12775 = pi93  & n4176;
  assign n12776 = pi94  & n3938;
  assign n12777 = pi95  & n3933;
  assign n12778 = n3475 & n3931;
  assign n12779 = ~n12776 & ~n12777;
  assign n12780 = ~n12775 & n12779;
  assign n12781 = ~n12778 & n12780;
  assign n12782 = pi35  & n12781;
  assign n12783 = ~pi35  & ~n12781;
  assign n12784 = ~n12782 & ~n12783;
  assign n12785 = ~n12774 & n12784;
  assign n12786 = n12774 & ~n12784;
  assign n12787 = ~n12785 & ~n12786;
  assign n12788 = ~n12405 & ~n12408;
  assign n12789 = n12787 & ~n12788;
  assign n12790 = ~n12787 & n12788;
  assign n12791 = ~n12789 & ~n12790;
  assign n12792 = pi96  & n3553;
  assign n12793 = pi97  & n3334;
  assign n12794 = pi98  & n3329;
  assign n12795 = n3327 & n3889;
  assign n12796 = ~n12793 & ~n12794;
  assign n12797 = ~n12792 & n12796;
  assign n12798 = ~n12795 & n12797;
  assign n12799 = pi32  & n12798;
  assign n12800 = ~pi32  & ~n12798;
  assign n12801 = ~n12799 & ~n12800;
  assign n12802 = n12791 & ~n12801;
  assign n12803 = ~n12791 & n12801;
  assign n12804 = ~n12802 & ~n12803;
  assign n12805 = n12617 & ~n12804;
  assign n12806 = ~n12617 & n12804;
  assign n12807 = ~n12805 & ~n12806;
  assign n12808 = pi99  & n3011;
  assign n12809 = pi100  & n2809;
  assign n12810 = pi101  & n2804;
  assign n12811 = n2802 & n4730;
  assign n12812 = ~n12809 & ~n12810;
  assign n12813 = ~n12808 & n12812;
  assign n12814 = ~n12811 & n12813;
  assign n12815 = pi29  & n12814;
  assign n12816 = ~pi29  & ~n12814;
  assign n12817 = ~n12815 & ~n12816;
  assign n12818 = n12807 & ~n12817;
  assign n12819 = ~n12807 & n12817;
  assign n12820 = ~n12818 & ~n12819;
  assign n12821 = n12616 & ~n12820;
  assign n12822 = ~n12616 & n12820;
  assign n12823 = ~n12821 & ~n12822;
  assign n12824 = pi102  & n2510;
  assign n12825 = pi103  & n2342;
  assign n12826 = pi104  & n2337;
  assign n12827 = n2335 & n5212;
  assign n12828 = ~n12825 & ~n12826;
  assign n12829 = ~n12824 & n12828;
  assign n12830 = ~n12827 & n12829;
  assign n12831 = pi26  & n12830;
  assign n12832 = ~pi26  & ~n12830;
  assign n12833 = ~n12831 & ~n12832;
  assign n12834 = n12823 & ~n12833;
  assign n12835 = ~n12823 & n12833;
  assign n12836 = ~n12834 & ~n12835;
  assign n12837 = ~n12615 & n12836;
  assign n12838 = n12615 & ~n12836;
  assign n12839 = ~n12837 & ~n12838;
  assign n12840 = ~n12614 & n12839;
  assign n12841 = n12614 & ~n12839;
  assign n12842 = ~n12840 & ~n12841;
  assign n12843 = ~n12604 & n12842;
  assign n12844 = n12604 & ~n12842;
  assign n12845 = ~n12843 & ~n12844;
  assign n12846 = ~n12603 & n12845;
  assign n12847 = n12603 & ~n12845;
  assign n12848 = ~n12846 & ~n12847;
  assign n12849 = ~n12593 & n12848;
  assign n12850 = n12593 & ~n12848;
  assign n12851 = ~n12849 & ~n12850;
  assign n12852 = ~n12592 & n12851;
  assign n12853 = n12592 & ~n12851;
  assign n12854 = ~n12852 & ~n12853;
  assign n12855 = ~n12582 & n12854;
  assign n12856 = n12582 & ~n12854;
  assign n12857 = ~n12855 & ~n12856;
  assign n12858 = ~n12581 & n12857;
  assign n12859 = n12581 & ~n12857;
  assign n12860 = ~n12858 & ~n12859;
  assign n12861 = ~n12571 & n12860;
  assign n12862 = n12571 & ~n12860;
  assign n12863 = ~n12861 & ~n12862;
  assign n12864 = ~n12570 & n12863;
  assign n12865 = n12570 & ~n12863;
  assign n12866 = ~n12864 & ~n12865;
  assign n12867 = ~n12560 & n12866;
  assign n12868 = n12560 & ~n12866;
  assign n12869 = ~n12867 & ~n12868;
  assign n12870 = pi120  & n528;
  assign n12871 = pi121  & n490;
  assign n12872 = pi122  & n485;
  assign n12873 = n483 & n10729;
  assign n12874 = ~n12871 & ~n12872;
  assign n12875 = ~n12870 & n12874;
  assign n12876 = ~n12873 & n12875;
  assign n12877 = pi8  & n12876;
  assign n12878 = ~pi8  & ~n12876;
  assign n12879 = ~n12877 & ~n12878;
  assign n12880 = n12869 & ~n12879;
  assign n12881 = ~n12869 & n12879;
  assign n12882 = ~n12880 & ~n12881;
  assign n12883 = ~n12559 & n12882;
  assign n12884 = n12559 & ~n12882;
  assign n12885 = ~n12883 & ~n12884;
  assign n12886 = ~n12549 & n12885;
  assign n12887 = n12549 & ~n12885;
  assign n12888 = ~n12886 & ~n12887;
  assign n12889 = ~n12548 & n12888;
  assign n12890 = n12548 & ~n12888;
  assign n12891 = ~n12889 & ~n12890;
  assign n12892 = ~n12507 & ~n12526;
  assign n12893 = ~n12508 & ~n12892;
  assign n12894 = n12891 & ~n12893;
  assign n12895 = ~n12891 & n12893;
  assign n12896 = ~n12894 & ~n12895;
  assign n12897 = ~n12536 & n12896;
  assign n12898 = n12536 & ~n12896;
  assign po64  = ~n12897 & ~n12898;
  assign n12900 = ~n12886 & ~n12889;
  assign n12901 = ~n12880 & ~n12883;
  assign n12902 = pi127  & n282;
  assign n12903 = pi127  & n262;
  assign n12904 = ~n12539 & n12903;
  assign n12905 = pi2  & ~n12902;
  assign n12906 = ~n12904 & n12905;
  assign n12907 = ~pi2  & n12904;
  assign n12908 = ~n12906 & ~n12907;
  assign n12909 = ~n12901 & ~n12908;
  assign n12910 = n12901 & n12908;
  assign n12911 = ~n12909 & ~n12910;
  assign n12912 = ~n12864 & ~n12867;
  assign n12913 = ~n12858 & ~n12861;
  assign n12914 = ~n12852 & ~n12855;
  assign n12915 = pi112  & n1296;
  assign n12916 = pi113  & n1207;
  assign n12917 = pi114  & n1202;
  assign n12918 = n1200 & n8146;
  assign n12919 = ~n12916 & ~n12917;
  assign n12920 = ~n12915 & n12919;
  assign n12921 = ~n12918 & n12920;
  assign n12922 = pi17  & n12921;
  assign n12923 = ~pi17  & ~n12921;
  assign n12924 = ~n12922 & ~n12923;
  assign n12925 = ~n12846 & ~n12849;
  assign n12926 = pi109  & n1661;
  assign n12927 = pi110  & n1500;
  assign n12928 = pi111  & n1495;
  assign n12929 = n1493 & n7272;
  assign n12930 = ~n12927 & ~n12928;
  assign n12931 = ~n12926 & n12930;
  assign n12932 = ~n12929 & n12931;
  assign n12933 = pi20  & n12932;
  assign n12934 = ~pi20  & ~n12932;
  assign n12935 = ~n12933 & ~n12934;
  assign n12936 = ~n12840 & ~n12843;
  assign n12937 = ~n12834 & ~n12837;
  assign n12938 = ~n12818 & ~n12822;
  assign n12939 = ~n12802 & ~n12806;
  assign n12940 = ~n12786 & ~n12789;
  assign n12941 = ~n12769 & ~n12773;
  assign n12942 = ~n12753 & ~n12757;
  assign n12943 = ~n12737 & ~n12741;
  assign n12944 = pi85  & n6331;
  assign n12945 = pi86  & n6015;
  assign n12946 = pi87  & n6010;
  assign n12947 = n2116 & n6008;
  assign n12948 = ~n12945 & ~n12946;
  assign n12949 = ~n12944 & n12948;
  assign n12950 = ~n12947 & n12949;
  assign n12951 = pi44  & n12950;
  assign n12952 = ~pi44  & ~n12950;
  assign n12953 = ~n12951 & ~n12952;
  assign n12954 = ~n12721 & ~n12724;
  assign n12955 = ~n12704 & ~n12708;
  assign n12956 = pi79  & n7969;
  assign n12957 = pi80  & n7636;
  assign n12958 = pi81  & n7631;
  assign n12959 = n1337 & n7629;
  assign n12960 = ~n12957 & ~n12958;
  assign n12961 = ~n12956 & n12960;
  assign n12962 = ~n12959 & n12961;
  assign n12963 = pi50  & n12962;
  assign n12964 = ~pi50  & ~n12962;
  assign n12965 = ~n12963 & ~n12964;
  assign n12966 = ~n12688 & ~n12691;
  assign n12967 = ~n12671 & ~n12675;
  assign n12968 = pi73  & n9858;
  assign n12969 = pi74  & n9508;
  assign n12970 = pi75  & n9503;
  assign n12971 = n713 & n9501;
  assign n12972 = ~n12969 & ~n12970;
  assign n12973 = ~n12968 & n12972;
  assign n12974 = ~n12971 & n12973;
  assign n12975 = pi56  & n12974;
  assign n12976 = ~pi56  & ~n12974;
  assign n12977 = ~n12975 & ~n12976;
  assign n12978 = ~n12656 & ~n12658;
  assign n12979 = ~n12637 & ~n12643;
  assign n12980 = pi67  & n11910;
  assign n12981 = pi68  & n11529;
  assign n12982 = pi69  & n11524;
  assign n12983 = n376 & n11522;
  assign n12984 = ~n12981 & ~n12982;
  assign n12985 = ~n12980 & n12984;
  assign n12986 = ~n12983 & n12985;
  assign n12987 = pi62  & n12986;
  assign n12988 = ~pi62  & ~n12986;
  assign n12989 = ~n12987 & ~n12988;
  assign n12990 = pi66  & n12277;
  assign n12991 = pi65  & n12276;
  assign n12992 = ~n12990 & ~n12991;
  assign n12993 = ~n12989 & ~n12992;
  assign n12994 = n12989 & n12992;
  assign n12995 = ~n12993 & ~n12994;
  assign n12996 = n12979 & ~n12995;
  assign n12997 = ~n12979 & n12995;
  assign n12998 = ~n12996 & ~n12997;
  assign n12999 = pi70  & n10886;
  assign n13000 = pi71  & n10495;
  assign n13001 = pi72  & n10490;
  assign n13002 = n551 & n10488;
  assign n13003 = ~n13000 & ~n13001;
  assign n13004 = ~n12999 & n13003;
  assign n13005 = ~n13002 & n13004;
  assign n13006 = pi59  & n13005;
  assign n13007 = ~pi59  & ~n13005;
  assign n13008 = ~n13006 & ~n13007;
  assign n13009 = n12998 & ~n13008;
  assign n13010 = ~n12998 & n13008;
  assign n13011 = ~n13009 & ~n13010;
  assign n13012 = ~n12978 & n13011;
  assign n13013 = n12978 & ~n13011;
  assign n13014 = ~n13012 & ~n13013;
  assign n13015 = n12977 & ~n13014;
  assign n13016 = ~n12977 & n13014;
  assign n13017 = ~n13015 & ~n13016;
  assign n13018 = ~n12967 & n13017;
  assign n13019 = n12967 & ~n13017;
  assign n13020 = ~n13018 & ~n13019;
  assign n13021 = pi76  & n8905;
  assign n13022 = pi77  & n8535;
  assign n13023 = pi78  & n8530;
  assign n13024 = n958 & n8528;
  assign n13025 = ~n13022 & ~n13023;
  assign n13026 = ~n13021 & n13025;
  assign n13027 = ~n13024 & n13026;
  assign n13028 = pi53  & n13027;
  assign n13029 = ~pi53  & ~n13027;
  assign n13030 = ~n13028 & ~n13029;
  assign n13031 = n13020 & ~n13030;
  assign n13032 = ~n13020 & n13030;
  assign n13033 = ~n13031 & ~n13032;
  assign n13034 = ~n12966 & n13033;
  assign n13035 = n12966 & ~n13033;
  assign n13036 = ~n13034 & ~n13035;
  assign n13037 = ~n12965 & n13036;
  assign n13038 = n12965 & ~n13036;
  assign n13039 = ~n13037 & ~n13038;
  assign n13040 = n12955 & ~n13039;
  assign n13041 = ~n12955 & n13039;
  assign n13042 = ~n13040 & ~n13041;
  assign n13043 = pi82  & n7121;
  assign n13044 = pi83  & n6795;
  assign n13045 = pi84  & n6790;
  assign n13046 = n1601 & n6788;
  assign n13047 = ~n13044 & ~n13045;
  assign n13048 = ~n13043 & n13047;
  assign n13049 = ~n13046 & n13048;
  assign n13050 = pi47  & n13049;
  assign n13051 = ~pi47  & ~n13049;
  assign n13052 = ~n13050 & ~n13051;
  assign n13053 = n13042 & ~n13052;
  assign n13054 = ~n13042 & n13052;
  assign n13055 = ~n13053 & ~n13054;
  assign n13056 = ~n12954 & n13055;
  assign n13057 = n12954 & ~n13055;
  assign n13058 = ~n13056 & ~n13057;
  assign n13059 = ~n12953 & n13058;
  assign n13060 = n12953 & ~n13058;
  assign n13061 = ~n13059 & ~n13060;
  assign n13062 = n12943 & ~n13061;
  assign n13063 = ~n12943 & n13061;
  assign n13064 = ~n13062 & ~n13063;
  assign n13065 = pi88  & n5558;
  assign n13066 = pi89  & n5293;
  assign n13067 = pi90  & n5288;
  assign n13068 = n2448 & n5286;
  assign n13069 = ~n13066 & ~n13067;
  assign n13070 = ~n13065 & n13069;
  assign n13071 = ~n13068 & n13070;
  assign n13072 = pi41  & n13071;
  assign n13073 = ~pi41  & ~n13071;
  assign n13074 = ~n13072 & ~n13073;
  assign n13075 = n13064 & ~n13074;
  assign n13076 = ~n13064 & n13074;
  assign n13077 = ~n13075 & ~n13076;
  assign n13078 = n12942 & ~n13077;
  assign n13079 = ~n12942 & n13077;
  assign n13080 = ~n13078 & ~n13079;
  assign n13081 = pi91  & n4843;
  assign n13082 = pi92  & n4598;
  assign n13083 = pi93  & n4593;
  assign n13084 = n2948 & n4591;
  assign n13085 = ~n13082 & ~n13083;
  assign n13086 = ~n13081 & n13085;
  assign n13087 = ~n13084 & n13086;
  assign n13088 = pi38  & n13087;
  assign n13089 = ~pi38  & ~n13087;
  assign n13090 = ~n13088 & ~n13089;
  assign n13091 = n13080 & ~n13090;
  assign n13092 = ~n13080 & n13090;
  assign n13093 = ~n13091 & ~n13092;
  assign n13094 = n12941 & ~n13093;
  assign n13095 = ~n12941 & n13093;
  assign n13096 = ~n13094 & ~n13095;
  assign n13097 = pi94  & n4176;
  assign n13098 = pi95  & n3938;
  assign n13099 = pi96  & n3933;
  assign n13100 = n3499 & n3931;
  assign n13101 = ~n13098 & ~n13099;
  assign n13102 = ~n13097 & n13101;
  assign n13103 = ~n13100 & n13102;
  assign n13104 = pi35  & n13103;
  assign n13105 = ~pi35  & ~n13103;
  assign n13106 = ~n13104 & ~n13105;
  assign n13107 = n13096 & ~n13106;
  assign n13108 = ~n13096 & n13106;
  assign n13109 = ~n13107 & ~n13108;
  assign n13110 = ~n12940 & n13109;
  assign n13111 = n12940 & ~n13109;
  assign n13112 = ~n13110 & ~n13111;
  assign n13113 = pi97  & n3553;
  assign n13114 = pi98  & n3334;
  assign n13115 = pi99  & n3329;
  assign n13116 = n3327 & n4101;
  assign n13117 = ~n13114 & ~n13115;
  assign n13118 = ~n13113 & n13117;
  assign n13119 = ~n13116 & n13118;
  assign n13120 = pi32  & n13119;
  assign n13121 = ~pi32  & ~n13119;
  assign n13122 = ~n13120 & ~n13121;
  assign n13123 = n13112 & ~n13122;
  assign n13124 = ~n13112 & n13122;
  assign n13125 = ~n13123 & ~n13124;
  assign n13126 = n12939 & ~n13125;
  assign n13127 = ~n12939 & n13125;
  assign n13128 = ~n13126 & ~n13127;
  assign n13129 = pi100  & n3011;
  assign n13130 = pi101  & n2809;
  assign n13131 = pi102  & n2804;
  assign n13132 = n2802 & n4956;
  assign n13133 = ~n13130 & ~n13131;
  assign n13134 = ~n13129 & n13133;
  assign n13135 = ~n13132 & n13134;
  assign n13136 = pi29  & n13135;
  assign n13137 = ~pi29  & ~n13135;
  assign n13138 = ~n13136 & ~n13137;
  assign n13139 = n13128 & ~n13138;
  assign n13140 = ~n13128 & n13138;
  assign n13141 = ~n13139 & ~n13140;
  assign n13142 = n12938 & ~n13141;
  assign n13143 = ~n12938 & n13141;
  assign n13144 = ~n13142 & ~n13143;
  assign n13145 = pi103  & n2510;
  assign n13146 = pi104  & n2342;
  assign n13147 = pi105  & n2337;
  assign n13148 = n2335 & n5677;
  assign n13149 = ~n13146 & ~n13147;
  assign n13150 = ~n13145 & n13149;
  assign n13151 = ~n13148 & n13150;
  assign n13152 = pi26  & n13151;
  assign n13153 = ~pi26  & ~n13151;
  assign n13154 = ~n13152 & ~n13153;
  assign n13155 = n13144 & ~n13154;
  assign n13156 = ~n13144 & n13154;
  assign n13157 = ~n13155 & ~n13156;
  assign n13158 = ~n12937 & n13157;
  assign n13159 = n12937 & ~n13157;
  assign n13160 = ~n13158 & ~n13159;
  assign n13161 = pi106  & n2053;
  assign n13162 = pi107  & n1893;
  assign n13163 = pi108  & n1888;
  assign n13164 = n1886 & n6213;
  assign n13165 = ~n13162 & ~n13163;
  assign n13166 = ~n13161 & n13165;
  assign n13167 = ~n13164 & n13166;
  assign n13168 = pi23  & n13167;
  assign n13169 = ~pi23  & ~n13167;
  assign n13170 = ~n13168 & ~n13169;
  assign n13171 = n13160 & ~n13170;
  assign n13172 = ~n13160 & n13170;
  assign n13173 = ~n13171 & ~n13172;
  assign n13174 = ~n12936 & n13173;
  assign n13175 = n12936 & ~n13173;
  assign n13176 = ~n13174 & ~n13175;
  assign n13177 = ~n12935 & n13176;
  assign n13178 = n12935 & ~n13176;
  assign n13179 = ~n13177 & ~n13178;
  assign n13180 = ~n12925 & n13179;
  assign n13181 = n12925 & ~n13179;
  assign n13182 = ~n13180 & ~n13181;
  assign n13183 = n12924 & ~n13182;
  assign n13184 = ~n12924 & n13182;
  assign n13185 = ~n13183 & ~n13184;
  assign n13186 = ~n12914 & n13185;
  assign n13187 = n12914 & ~n13185;
  assign n13188 = ~n13186 & ~n13187;
  assign n13189 = pi115  & n1006;
  assign n13190 = pi116  & n897;
  assign n13191 = pi117  & n892;
  assign n13192 = n890 & n8784;
  assign n13193 = ~n13190 & ~n13191;
  assign n13194 = ~n13189 & n13193;
  assign n13195 = ~n13192 & n13194;
  assign n13196 = pi14  & n13195;
  assign n13197 = ~pi14  & ~n13195;
  assign n13198 = ~n13196 & ~n13197;
  assign n13199 = n13188 & ~n13198;
  assign n13200 = ~n13188 & n13198;
  assign n13201 = ~n13199 & ~n13200;
  assign n13202 = n12913 & ~n13201;
  assign n13203 = ~n12913 & n13201;
  assign n13204 = ~n13202 & ~n13203;
  assign n13205 = pi118  & n750;
  assign n13206 = pi119  & n651;
  assign n13207 = pi120  & n646;
  assign n13208 = n644 & n10047;
  assign n13209 = ~n13206 & ~n13207;
  assign n13210 = ~n13205 & n13209;
  assign n13211 = ~n13208 & n13210;
  assign n13212 = pi11  & n13211;
  assign n13213 = ~pi11  & ~n13211;
  assign n13214 = ~n13212 & ~n13213;
  assign n13215 = ~n13204 & n13214;
  assign n13216 = n13204 & ~n13214;
  assign n13217 = ~n13215 & ~n13216;
  assign n13218 = pi121  & n528;
  assign n13219 = pi122  & n490;
  assign n13220 = pi123  & n485;
  assign n13221 = n483 & n10754;
  assign n13222 = ~n13219 & ~n13220;
  assign n13223 = ~n13218 & n13222;
  assign n13224 = ~n13221 & n13223;
  assign n13225 = pi8  & n13224;
  assign n13226 = ~pi8  & ~n13224;
  assign n13227 = ~n13225 & ~n13226;
  assign n13228 = n13217 & ~n13227;
  assign n13229 = ~n13217 & n13227;
  assign n13230 = ~n13228 & ~n13229;
  assign n13231 = n12912 & ~n13230;
  assign n13232 = ~n12912 & n13230;
  assign n13233 = ~n13231 & ~n13232;
  assign n13234 = pi124  & n391;
  assign n13235 = pi125  & n353;
  assign n13236 = pi126  & n348;
  assign n13237 = n346 & n12148;
  assign n13238 = ~n13235 & ~n13236;
  assign n13239 = ~n13234 & n13238;
  assign n13240 = ~n13237 & n13239;
  assign n13241 = pi5  & n13240;
  assign n13242 = ~pi5  & ~n13240;
  assign n13243 = ~n13241 & ~n13242;
  assign n13244 = n13233 & ~n13243;
  assign n13245 = ~n13233 & n13243;
  assign n13246 = ~n13244 & ~n13245;
  assign n13247 = n12911 & n13246;
  assign n13248 = ~n12911 & ~n13246;
  assign n13249 = ~n13247 & ~n13248;
  assign n13250 = n12900 & ~n13249;
  assign n13251 = ~n12900 & n13249;
  assign n13252 = ~n13250 & ~n13251;
  assign n13253 = ~n12894 & ~n12897;
  assign n13254 = n13252 & ~n13253;
  assign n13255 = ~n13252 & n13253;
  assign po65  = ~n13254 & ~n13255;
  assign n13257 = pi119  & n750;
  assign n13258 = pi120  & n651;
  assign n13259 = pi121  & n646;
  assign n13260 = n644 & n10071;
  assign n13261 = ~n13258 & ~n13259;
  assign n13262 = ~n13257 & n13261;
  assign n13263 = ~n13260 & n13262;
  assign n13264 = pi11  & n13263;
  assign n13265 = ~pi11  & ~n13263;
  assign n13266 = ~n13264 & ~n13265;
  assign n13267 = ~n13199 & ~n13203;
  assign n13268 = n13266 & n13267;
  assign n13269 = ~n13266 & ~n13267;
  assign n13270 = ~n13268 & ~n13269;
  assign n13271 = pi113  & n1296;
  assign n13272 = pi114  & n1207;
  assign n13273 = pi115  & n1202;
  assign n13274 = n1200 & n8170;
  assign n13275 = ~n13272 & ~n13273;
  assign n13276 = ~n13271 & n13275;
  assign n13277 = ~n13274 & n13276;
  assign n13278 = pi17  & n13277;
  assign n13279 = ~pi17  & ~n13277;
  assign n13280 = ~n13278 & ~n13279;
  assign n13281 = ~n13177 & ~n13180;
  assign n13282 = n13280 & n13281;
  assign n13283 = ~n13280 & ~n13281;
  assign n13284 = ~n13282 & ~n13283;
  assign n13285 = pi110  & n1661;
  assign n13286 = pi111  & n1500;
  assign n13287 = pi112  & n1495;
  assign n13288 = n1493 & n7296;
  assign n13289 = ~n13286 & ~n13287;
  assign n13290 = ~n13285 & n13289;
  assign n13291 = ~n13288 & n13290;
  assign n13292 = pi20  & n13291;
  assign n13293 = ~pi20  & ~n13291;
  assign n13294 = ~n13292 & ~n13293;
  assign n13295 = ~n13171 & ~n13174;
  assign n13296 = n13294 & n13295;
  assign n13297 = ~n13294 & ~n13295;
  assign n13298 = ~n13296 & ~n13297;
  assign n13299 = pi104  & n2510;
  assign n13300 = pi105  & n2342;
  assign n13301 = pi106  & n2337;
  assign n13302 = n2335 & n5701;
  assign n13303 = ~n13300 & ~n13301;
  assign n13304 = ~n13299 & n13303;
  assign n13305 = ~n13302 & n13304;
  assign n13306 = pi26  & n13305;
  assign n13307 = ~pi26  & ~n13305;
  assign n13308 = ~n13306 & ~n13307;
  assign n13309 = ~n13139 & ~n13143;
  assign n13310 = n13308 & n13309;
  assign n13311 = ~n13308 & ~n13309;
  assign n13312 = ~n13310 & ~n13311;
  assign n13313 = ~n13123 & ~n13127;
  assign n13314 = pi101  & n3011;
  assign n13315 = pi102  & n2809;
  assign n13316 = pi103  & n2804;
  assign n13317 = n2802 & n5188;
  assign n13318 = ~n13315 & ~n13316;
  assign n13319 = ~n13314 & n13318;
  assign n13320 = ~n13317 & n13319;
  assign n13321 = pi29  & n13320;
  assign n13322 = ~pi29  & ~n13320;
  assign n13323 = ~n13321 & ~n13322;
  assign n13324 = ~n13313 & ~n13323;
  assign n13325 = n13313 & n13323;
  assign n13326 = ~n13324 & ~n13325;
  assign n13327 = ~n13107 & ~n13110;
  assign n13328 = pi98  & n3553;
  assign n13329 = pi99  & n3334;
  assign n13330 = pi100  & n3329;
  assign n13331 = n3327 & n4501;
  assign n13332 = ~n13329 & ~n13330;
  assign n13333 = ~n13328 & n13332;
  assign n13334 = ~n13331 & n13333;
  assign n13335 = pi32  & n13334;
  assign n13336 = ~pi32  & ~n13334;
  assign n13337 = ~n13335 & ~n13336;
  assign n13338 = ~n13327 & ~n13337;
  assign n13339 = n13327 & n13337;
  assign n13340 = ~n13338 & ~n13339;
  assign n13341 = ~n13075 & ~n13079;
  assign n13342 = ~n13059 & ~n13063;
  assign n13343 = ~n13037 & ~n13041;
  assign n13344 = ~n13031 & ~n13034;
  assign n13345 = ~n13016 & ~n13018;
  assign n13346 = pi74  & n9858;
  assign n13347 = pi75  & n9508;
  assign n13348 = pi76  & n9503;
  assign n13349 = n841 & n9501;
  assign n13350 = ~n13347 & ~n13348;
  assign n13351 = ~n13346 & n13350;
  assign n13352 = ~n13349 & n13351;
  assign n13353 = pi56  & n13352;
  assign n13354 = ~pi56  & ~n13352;
  assign n13355 = ~n13353 & ~n13354;
  assign n13356 = ~n13009 & ~n13012;
  assign n13357 = ~n12993 & ~n12997;
  assign n13358 = pi67  & n12277;
  assign n13359 = pi66  & n12276;
  assign n13360 = ~n13358 & ~n13359;
  assign n13361 = pi2  & ~n13360;
  assign n13362 = ~pi2  & n13360;
  assign n13363 = ~n13361 & ~n13362;
  assign n13364 = pi68  & n11910;
  assign n13365 = pi69  & n11529;
  assign n13366 = pi70  & n11524;
  assign n13367 = n415 & n11522;
  assign n13368 = ~n13365 & ~n13366;
  assign n13369 = ~n13364 & n13368;
  assign n13370 = ~n13367 & n13369;
  assign n13371 = pi62  & n13370;
  assign n13372 = ~pi62  & ~n13370;
  assign n13373 = ~n13371 & ~n13372;
  assign n13374 = n13363 & ~n13373;
  assign n13375 = ~n13363 & n13373;
  assign n13376 = ~n13374 & ~n13375;
  assign n13377 = ~n13357 & n13376;
  assign n13378 = n13357 & ~n13376;
  assign n13379 = ~n13377 & ~n13378;
  assign n13380 = pi71  & n10886;
  assign n13381 = pi72  & n10495;
  assign n13382 = pi73  & n10490;
  assign n13383 = n613 & n10488;
  assign n13384 = ~n13381 & ~n13382;
  assign n13385 = ~n13380 & n13384;
  assign n13386 = ~n13383 & n13385;
  assign n13387 = pi59  & n13386;
  assign n13388 = ~pi59  & ~n13386;
  assign n13389 = ~n13387 & ~n13388;
  assign n13390 = n13379 & ~n13389;
  assign n13391 = ~n13379 & n13389;
  assign n13392 = ~n13390 & ~n13391;
  assign n13393 = ~n13356 & n13392;
  assign n13394 = n13356 & ~n13392;
  assign n13395 = ~n13393 & ~n13394;
  assign n13396 = n13355 & ~n13395;
  assign n13397 = ~n13355 & n13395;
  assign n13398 = ~n13396 & ~n13397;
  assign n13399 = ~n13345 & n13398;
  assign n13400 = n13345 & ~n13398;
  assign n13401 = ~n13399 & ~n13400;
  assign n13402 = pi77  & n8905;
  assign n13403 = pi78  & n8535;
  assign n13404 = pi79  & n8530;
  assign n13405 = n1048 & n8528;
  assign n13406 = ~n13403 & ~n13404;
  assign n13407 = ~n13402 & n13406;
  assign n13408 = ~n13405 & n13407;
  assign n13409 = pi53  & n13408;
  assign n13410 = ~pi53  & ~n13408;
  assign n13411 = ~n13409 & ~n13410;
  assign n13412 = n13401 & ~n13411;
  assign n13413 = ~n13401 & n13411;
  assign n13414 = ~n13412 & ~n13413;
  assign n13415 = n13344 & ~n13414;
  assign n13416 = ~n13344 & n13414;
  assign n13417 = ~n13415 & ~n13416;
  assign n13418 = pi80  & n7969;
  assign n13419 = pi81  & n7636;
  assign n13420 = pi82  & n7631;
  assign n13421 = n1450 & n7629;
  assign n13422 = ~n13419 & ~n13420;
  assign n13423 = ~n13418 & n13422;
  assign n13424 = ~n13421 & n13423;
  assign n13425 = pi50  & n13424;
  assign n13426 = ~pi50  & ~n13424;
  assign n13427 = ~n13425 & ~n13426;
  assign n13428 = n13417 & ~n13427;
  assign n13429 = ~n13417 & n13427;
  assign n13430 = ~n13428 & ~n13429;
  assign n13431 = n13343 & ~n13430;
  assign n13432 = ~n13343 & n13430;
  assign n13433 = ~n13431 & ~n13432;
  assign n13434 = pi83  & n7121;
  assign n13435 = pi84  & n6795;
  assign n13436 = pi85  & n6790;
  assign n13437 = n1831 & n6788;
  assign n13438 = ~n13435 & ~n13436;
  assign n13439 = ~n13434 & n13438;
  assign n13440 = ~n13437 & n13439;
  assign n13441 = pi47  & n13440;
  assign n13442 = ~pi47  & ~n13440;
  assign n13443 = ~n13441 & ~n13442;
  assign n13444 = ~n13433 & n13443;
  assign n13445 = n13433 & ~n13443;
  assign n13446 = ~n13444 & ~n13445;
  assign n13447 = ~n13053 & ~n13056;
  assign n13448 = n13446 & ~n13447;
  assign n13449 = ~n13446 & n13447;
  assign n13450 = ~n13448 & ~n13449;
  assign n13451 = pi86  & n6331;
  assign n13452 = pi87  & n6015;
  assign n13453 = pi88  & n6010;
  assign n13454 = n2140 & n6008;
  assign n13455 = ~n13452 & ~n13453;
  assign n13456 = ~n13451 & n13455;
  assign n13457 = ~n13454 & n13456;
  assign n13458 = pi44  & n13457;
  assign n13459 = ~pi44  & ~n13457;
  assign n13460 = ~n13458 & ~n13459;
  assign n13461 = n13450 & ~n13460;
  assign n13462 = ~n13450 & n13460;
  assign n13463 = ~n13461 & ~n13462;
  assign n13464 = n13342 & ~n13463;
  assign n13465 = ~n13342 & n13463;
  assign n13466 = ~n13464 & ~n13465;
  assign n13467 = pi89  & n5558;
  assign n13468 = pi90  & n5293;
  assign n13469 = pi91  & n5288;
  assign n13470 = n2746 & n5286;
  assign n13471 = ~n13468 & ~n13469;
  assign n13472 = ~n13467 & n13471;
  assign n13473 = ~n13470 & n13472;
  assign n13474 = pi41  & n13473;
  assign n13475 = ~pi41  & ~n13473;
  assign n13476 = ~n13474 & ~n13475;
  assign n13477 = n13466 & ~n13476;
  assign n13478 = ~n13466 & n13476;
  assign n13479 = ~n13477 & ~n13478;
  assign n13480 = n13341 & ~n13479;
  assign n13481 = ~n13341 & n13479;
  assign n13482 = ~n13480 & ~n13481;
  assign n13483 = pi92  & n4843;
  assign n13484 = pi93  & n4598;
  assign n13485 = pi94  & n4593;
  assign n13486 = n3280 & n4591;
  assign n13487 = ~n13484 & ~n13485;
  assign n13488 = ~n13483 & n13487;
  assign n13489 = ~n13486 & n13488;
  assign n13490 = pi38  & n13489;
  assign n13491 = ~pi38  & ~n13489;
  assign n13492 = ~n13490 & ~n13491;
  assign n13493 = ~n13482 & n13492;
  assign n13494 = n13482 & ~n13492;
  assign n13495 = ~n13493 & ~n13494;
  assign n13496 = ~n13091 & ~n13095;
  assign n13497 = n13495 & ~n13496;
  assign n13498 = ~n13495 & n13496;
  assign n13499 = ~n13497 & ~n13498;
  assign n13500 = pi95  & n4176;
  assign n13501 = pi96  & n3938;
  assign n13502 = pi97  & n3933;
  assign n13503 = n3691 & n3931;
  assign n13504 = ~n13501 & ~n13502;
  assign n13505 = ~n13500 & n13504;
  assign n13506 = ~n13503 & n13505;
  assign n13507 = pi35  & n13506;
  assign n13508 = ~pi35  & ~n13506;
  assign n13509 = ~n13507 & ~n13508;
  assign n13510 = n13499 & ~n13509;
  assign n13511 = ~n13499 & n13509;
  assign n13512 = ~n13510 & ~n13511;
  assign n13513 = n13340 & n13512;
  assign n13514 = ~n13340 & ~n13512;
  assign n13515 = ~n13513 & ~n13514;
  assign n13516 = n13326 & n13515;
  assign n13517 = ~n13326 & ~n13515;
  assign n13518 = ~n13516 & ~n13517;
  assign n13519 = n13312 & n13518;
  assign n13520 = ~n13312 & ~n13518;
  assign n13521 = ~n13519 & ~n13520;
  assign n13522 = ~n13155 & ~n13158;
  assign n13523 = pi107  & n2053;
  assign n13524 = pi108  & n1893;
  assign n13525 = pi109  & n1888;
  assign n13526 = n1886 & n6715;
  assign n13527 = ~n13524 & ~n13525;
  assign n13528 = ~n13523 & n13527;
  assign n13529 = ~n13526 & n13528;
  assign n13530 = pi23  & n13529;
  assign n13531 = ~pi23  & ~n13529;
  assign n13532 = ~n13530 & ~n13531;
  assign n13533 = ~n13522 & ~n13532;
  assign n13534 = n13522 & n13532;
  assign n13535 = ~n13533 & ~n13534;
  assign n13536 = n13521 & n13535;
  assign n13537 = ~n13521 & ~n13535;
  assign n13538 = ~n13536 & ~n13537;
  assign n13539 = n13298 & n13538;
  assign n13540 = ~n13298 & ~n13538;
  assign n13541 = ~n13539 & ~n13540;
  assign n13542 = n13284 & n13541;
  assign n13543 = ~n13284 & ~n13541;
  assign n13544 = ~n13542 & ~n13543;
  assign n13545 = ~n13184 & ~n13186;
  assign n13546 = pi116  & n1006;
  assign n13547 = pi117  & n897;
  assign n13548 = pi118  & n892;
  assign n13549 = n890 & n9095;
  assign n13550 = ~n13547 & ~n13548;
  assign n13551 = ~n13546 & n13550;
  assign n13552 = ~n13549 & n13551;
  assign n13553 = pi14  & n13552;
  assign n13554 = ~pi14  & ~n13552;
  assign n13555 = ~n13553 & ~n13554;
  assign n13556 = ~n13545 & ~n13555;
  assign n13557 = n13545 & n13555;
  assign n13558 = ~n13556 & ~n13557;
  assign n13559 = n13544 & n13558;
  assign n13560 = ~n13544 & ~n13558;
  assign n13561 = ~n13559 & ~n13560;
  assign n13562 = n13270 & ~n13561;
  assign n13563 = ~n13270 & n13561;
  assign n13564 = ~n13562 & ~n13563;
  assign n13565 = pi122  & n528;
  assign n13566 = pi123  & n490;
  assign n13567 = pi124  & n485;
  assign n13568 = n483 & n11099;
  assign n13569 = ~n13566 & ~n13567;
  assign n13570 = ~n13565 & n13569;
  assign n13571 = ~n13568 & n13570;
  assign n13572 = pi8  & n13571;
  assign n13573 = ~pi8  & ~n13571;
  assign n13574 = ~n13572 & ~n13573;
  assign n13575 = ~n13215 & ~n13227;
  assign n13576 = ~n13216 & ~n13575;
  assign n13577 = ~n13574 & ~n13576;
  assign n13578 = n13574 & n13576;
  assign n13579 = ~n13577 & ~n13578;
  assign n13580 = ~n13564 & n13579;
  assign n13581 = n13564 & ~n13579;
  assign n13582 = ~n13580 & ~n13581;
  assign n13583 = pi125  & n391;
  assign n13584 = pi126  & n353;
  assign n13585 = pi127  & n348;
  assign n13586 = n346 & n12519;
  assign n13587 = ~n13584 & ~n13585;
  assign n13588 = ~n13583 & n13587;
  assign n13589 = ~n13586 & n13588;
  assign n13590 = pi5  & n13589;
  assign n13591 = ~pi5  & ~n13589;
  assign n13592 = ~n13590 & ~n13591;
  assign n13593 = ~n13232 & n13243;
  assign n13594 = ~n13231 & ~n13593;
  assign n13595 = ~n13592 & n13594;
  assign n13596 = n13592 & ~n13594;
  assign n13597 = ~n13595 & ~n13596;
  assign n13598 = n13582 & n13597;
  assign n13599 = ~n13582 & ~n13597;
  assign n13600 = ~n13598 & ~n13599;
  assign n13601 = ~n12909 & ~n13246;
  assign n13602 = ~n12910 & ~n13601;
  assign n13603 = ~n13600 & ~n13602;
  assign n13604 = n13600 & n13602;
  assign n13605 = ~n13603 & ~n13604;
  assign n13606 = ~n13251 & ~n13254;
  assign n13607 = n13605 & ~n13606;
  assign n13608 = ~n13605 & n13606;
  assign po66  = ~n13607 & ~n13608;
  assign n13610 = ~n13604 & ~n13607;
  assign n13611 = ~n13595 & ~n13598;
  assign n13612 = pi117  & n1006;
  assign n13613 = pi118  & n897;
  assign n13614 = pi119  & n892;
  assign n13615 = n890 & n9412;
  assign n13616 = ~n13613 & ~n13614;
  assign n13617 = ~n13612 & n13616;
  assign n13618 = ~n13615 & n13617;
  assign n13619 = pi14  & n13618;
  assign n13620 = ~pi14  & ~n13618;
  assign n13621 = ~n13619 & ~n13620;
  assign n13622 = ~n13283 & ~n13542;
  assign n13623 = n13621 & n13622;
  assign n13624 = ~n13621 & ~n13622;
  assign n13625 = ~n13623 & ~n13624;
  assign n13626 = pi111  & n1661;
  assign n13627 = pi112  & n1500;
  assign n13628 = pi113  & n1495;
  assign n13629 = n1493 & n7852;
  assign n13630 = ~n13627 & ~n13628;
  assign n13631 = ~n13626 & n13630;
  assign n13632 = ~n13629 & n13631;
  assign n13633 = pi20  & n13632;
  assign n13634 = ~pi20  & ~n13632;
  assign n13635 = ~n13633 & ~n13634;
  assign n13636 = ~n13533 & ~n13536;
  assign n13637 = n13635 & n13636;
  assign n13638 = ~n13635 & ~n13636;
  assign n13639 = ~n13637 & ~n13638;
  assign n13640 = pi105  & n2510;
  assign n13641 = pi106  & n2342;
  assign n13642 = pi107  & n2337;
  assign n13643 = n2335 & n6189;
  assign n13644 = ~n13641 & ~n13642;
  assign n13645 = ~n13640 & n13644;
  assign n13646 = ~n13643 & n13645;
  assign n13647 = pi26  & n13646;
  assign n13648 = ~pi26  & ~n13646;
  assign n13649 = ~n13647 & ~n13648;
  assign n13650 = ~n13324 & ~n13516;
  assign n13651 = n13649 & n13650;
  assign n13652 = ~n13649 & ~n13650;
  assign n13653 = ~n13651 & ~n13652;
  assign n13654 = pi99  & n3553;
  assign n13655 = pi100  & n3334;
  assign n13656 = pi101  & n3329;
  assign n13657 = n3327 & n4730;
  assign n13658 = ~n13655 & ~n13656;
  assign n13659 = ~n13654 & n13658;
  assign n13660 = ~n13657 & n13659;
  assign n13661 = pi32  & n13660;
  assign n13662 = ~pi32  & ~n13660;
  assign n13663 = ~n13661 & ~n13662;
  assign n13664 = ~n13498 & ~n13509;
  assign n13665 = ~n13497 & ~n13664;
  assign n13666 = ~n13663 & ~n13665;
  assign n13667 = n13663 & n13665;
  assign n13668 = ~n13666 & ~n13667;
  assign n13669 = pi96  & n4176;
  assign n13670 = pi97  & n3938;
  assign n13671 = pi98  & n3933;
  assign n13672 = n3889 & n3931;
  assign n13673 = ~n13670 & ~n13671;
  assign n13674 = ~n13669 & n13673;
  assign n13675 = ~n13672 & n13674;
  assign n13676 = pi35  & n13675;
  assign n13677 = ~pi35  & ~n13675;
  assign n13678 = ~n13676 & ~n13677;
  assign n13679 = ~n13481 & ~n13494;
  assign n13680 = pi87  & n6331;
  assign n13681 = pi88  & n6015;
  assign n13682 = pi89  & n6010;
  assign n13683 = n2287 & n6008;
  assign n13684 = ~n13681 & ~n13682;
  assign n13685 = ~n13680 & n13684;
  assign n13686 = ~n13683 & n13685;
  assign n13687 = pi44  & n13686;
  assign n13688 = ~pi44  & ~n13686;
  assign n13689 = ~n13687 & ~n13688;
  assign n13690 = ~n13432 & ~n13445;
  assign n13691 = ~n13361 & ~n13374;
  assign n13692 = pi69  & n11910;
  assign n13693 = pi70  & n11529;
  assign n13694 = pi71  & n11524;
  assign n13695 = n460 & n11522;
  assign n13696 = ~n13693 & ~n13694;
  assign n13697 = ~n13692 & n13696;
  assign n13698 = ~n13695 & n13697;
  assign n13699 = pi62  & n13698;
  assign n13700 = ~pi62  & ~n13698;
  assign n13701 = ~n13699 & ~n13700;
  assign n13702 = pi68  & n12277;
  assign n13703 = pi67  & n12276;
  assign n13704 = ~n13702 & ~n13703;
  assign n13705 = pi2  & ~n13704;
  assign n13706 = ~pi2  & n13704;
  assign n13707 = ~n13705 & ~n13706;
  assign n13708 = ~n13701 & n13707;
  assign n13709 = n13701 & ~n13707;
  assign n13710 = ~n13708 & ~n13709;
  assign n13711 = n13691 & ~n13710;
  assign n13712 = ~n13691 & n13710;
  assign n13713 = ~n13711 & ~n13712;
  assign n13714 = pi72  & n10886;
  assign n13715 = pi73  & n10495;
  assign n13716 = pi74  & n10490;
  assign n13717 = n689 & n10488;
  assign n13718 = ~n13715 & ~n13716;
  assign n13719 = ~n13714 & n13718;
  assign n13720 = ~n13717 & n13719;
  assign n13721 = pi59  & n13720;
  assign n13722 = ~pi59  & ~n13720;
  assign n13723 = ~n13721 & ~n13722;
  assign n13724 = n13713 & ~n13723;
  assign n13725 = ~n13713 & n13723;
  assign n13726 = ~n13724 & ~n13725;
  assign n13727 = ~n13377 & n13389;
  assign n13728 = ~n13378 & ~n13727;
  assign n13729 = ~n13726 & ~n13728;
  assign n13730 = n13726 & n13728;
  assign n13731 = ~n13729 & ~n13730;
  assign n13732 = pi75  & n9858;
  assign n13733 = pi76  & n9508;
  assign n13734 = pi77  & n9503;
  assign n13735 = n865 & n9501;
  assign n13736 = ~n13733 & ~n13734;
  assign n13737 = ~n13732 & n13736;
  assign n13738 = ~n13735 & n13737;
  assign n13739 = pi56  & n13738;
  assign n13740 = ~pi56  & ~n13738;
  assign n13741 = ~n13739 & ~n13740;
  assign n13742 = ~n13731 & n13741;
  assign n13743 = n13731 & ~n13741;
  assign n13744 = ~n13742 & ~n13743;
  assign n13745 = ~n13393 & ~n13397;
  assign n13746 = n13744 & ~n13745;
  assign n13747 = ~n13744 & n13745;
  assign n13748 = ~n13746 & ~n13747;
  assign n13749 = pi78  & n8905;
  assign n13750 = pi79  & n8535;
  assign n13751 = pi80  & n8530;
  assign n13752 = n1144 & n8528;
  assign n13753 = ~n13750 & ~n13751;
  assign n13754 = ~n13749 & n13753;
  assign n13755 = ~n13752 & n13754;
  assign n13756 = pi53  & n13755;
  assign n13757 = ~pi53  & ~n13755;
  assign n13758 = ~n13756 & ~n13757;
  assign n13759 = n13748 & ~n13758;
  assign n13760 = ~n13748 & n13758;
  assign n13761 = ~n13759 & ~n13760;
  assign n13762 = ~n13399 & n13411;
  assign n13763 = ~n13400 & ~n13762;
  assign n13764 = ~n13761 & ~n13763;
  assign n13765 = n13761 & n13763;
  assign n13766 = ~n13764 & ~n13765;
  assign n13767 = pi81  & n7969;
  assign n13768 = pi82  & n7636;
  assign n13769 = pi83  & n7631;
  assign n13770 = n1577 & n7629;
  assign n13771 = ~n13768 & ~n13769;
  assign n13772 = ~n13767 & n13771;
  assign n13773 = ~n13770 & n13772;
  assign n13774 = pi50  & n13773;
  assign n13775 = ~pi50  & ~n13773;
  assign n13776 = ~n13774 & ~n13775;
  assign n13777 = n13766 & ~n13776;
  assign n13778 = ~n13766 & n13776;
  assign n13779 = ~n13777 & ~n13778;
  assign n13780 = ~n13416 & n13427;
  assign n13781 = ~n13415 & ~n13780;
  assign n13782 = ~n13779 & ~n13781;
  assign n13783 = n13779 & n13781;
  assign n13784 = ~n13782 & ~n13783;
  assign n13785 = pi84  & n7121;
  assign n13786 = pi85  & n6795;
  assign n13787 = pi86  & n6790;
  assign n13788 = n1975 & n6788;
  assign n13789 = ~n13786 & ~n13787;
  assign n13790 = ~n13785 & n13789;
  assign n13791 = ~n13788 & n13790;
  assign n13792 = pi47  & n13791;
  assign n13793 = ~pi47  & ~n13791;
  assign n13794 = ~n13792 & ~n13793;
  assign n13795 = n13784 & ~n13794;
  assign n13796 = ~n13784 & n13794;
  assign n13797 = ~n13795 & ~n13796;
  assign n13798 = ~n13690 & n13797;
  assign n13799 = n13690 & ~n13797;
  assign n13800 = ~n13798 & ~n13799;
  assign n13801 = ~n13689 & n13800;
  assign n13802 = n13689 & ~n13800;
  assign n13803 = ~n13801 & ~n13802;
  assign n13804 = ~n13449 & ~n13460;
  assign n13805 = ~n13448 & ~n13804;
  assign n13806 = ~n13803 & n13805;
  assign n13807 = n13803 & ~n13805;
  assign n13808 = ~n13806 & ~n13807;
  assign n13809 = pi90  & n5558;
  assign n13810 = pi91  & n5293;
  assign n13811 = pi92  & n5288;
  assign n13812 = n2924 & n5286;
  assign n13813 = ~n13810 & ~n13811;
  assign n13814 = ~n13809 & n13813;
  assign n13815 = ~n13812 & n13814;
  assign n13816 = pi41  & n13815;
  assign n13817 = ~pi41  & ~n13815;
  assign n13818 = ~n13816 & ~n13817;
  assign n13819 = n13808 & ~n13818;
  assign n13820 = ~n13808 & n13818;
  assign n13821 = ~n13819 & ~n13820;
  assign n13822 = ~n13465 & n13476;
  assign n13823 = ~n13464 & ~n13822;
  assign n13824 = ~n13821 & ~n13823;
  assign n13825 = n13821 & n13823;
  assign n13826 = ~n13824 & ~n13825;
  assign n13827 = pi93  & n4843;
  assign n13828 = pi94  & n4598;
  assign n13829 = pi95  & n4593;
  assign n13830 = n3475 & n4591;
  assign n13831 = ~n13828 & ~n13829;
  assign n13832 = ~n13827 & n13831;
  assign n13833 = ~n13830 & n13832;
  assign n13834 = pi38  & n13833;
  assign n13835 = ~pi38  & ~n13833;
  assign n13836 = ~n13834 & ~n13835;
  assign n13837 = ~n13826 & n13836;
  assign n13838 = n13826 & ~n13836;
  assign n13839 = ~n13837 & ~n13838;
  assign n13840 = ~n13679 & n13839;
  assign n13841 = n13679 & ~n13839;
  assign n13842 = ~n13840 & ~n13841;
  assign n13843 = n13678 & ~n13842;
  assign n13844 = ~n13678 & n13842;
  assign n13845 = ~n13843 & ~n13844;
  assign n13846 = ~n13668 & ~n13845;
  assign n13847 = n13668 & n13845;
  assign n13848 = ~n13846 & ~n13847;
  assign n13849 = ~n13338 & ~n13513;
  assign n13850 = pi102  & n3011;
  assign n13851 = pi103  & n2809;
  assign n13852 = pi104  & n2804;
  assign n13853 = n2802 & n5212;
  assign n13854 = ~n13851 & ~n13852;
  assign n13855 = ~n13850 & n13854;
  assign n13856 = ~n13853 & n13855;
  assign n13857 = pi29  & n13856;
  assign n13858 = ~pi29  & ~n13856;
  assign n13859 = ~n13857 & ~n13858;
  assign n13860 = ~n13849 & ~n13859;
  assign n13861 = n13849 & n13859;
  assign n13862 = ~n13860 & ~n13861;
  assign n13863 = n13848 & n13862;
  assign n13864 = ~n13848 & ~n13862;
  assign n13865 = ~n13863 & ~n13864;
  assign n13866 = n13653 & n13865;
  assign n13867 = ~n13653 & ~n13865;
  assign n13868 = ~n13866 & ~n13867;
  assign n13869 = pi108  & n2053;
  assign n13870 = pi109  & n1893;
  assign n13871 = pi110  & n1888;
  assign n13872 = n1886 & n6995;
  assign n13873 = ~n13870 & ~n13871;
  assign n13874 = ~n13869 & n13873;
  assign n13875 = ~n13872 & n13874;
  assign n13876 = pi23  & n13875;
  assign n13877 = ~pi23  & ~n13875;
  assign n13878 = ~n13876 & ~n13877;
  assign n13879 = ~n13311 & ~n13519;
  assign n13880 = ~n13878 & ~n13879;
  assign n13881 = n13878 & n13879;
  assign n13882 = ~n13880 & ~n13881;
  assign n13883 = n13868 & n13882;
  assign n13884 = ~n13868 & ~n13882;
  assign n13885 = ~n13883 & ~n13884;
  assign n13886 = n13639 & n13885;
  assign n13887 = ~n13639 & ~n13885;
  assign n13888 = ~n13886 & ~n13887;
  assign n13889 = pi114  & n1296;
  assign n13890 = pi115  & n1207;
  assign n13891 = pi116  & n1202;
  assign n13892 = n1200 & n8470;
  assign n13893 = ~n13890 & ~n13891;
  assign n13894 = ~n13889 & n13893;
  assign n13895 = ~n13892 & n13894;
  assign n13896 = pi17  & n13895;
  assign n13897 = ~pi17  & ~n13895;
  assign n13898 = ~n13896 & ~n13897;
  assign n13899 = ~n13297 & ~n13539;
  assign n13900 = ~n13898 & ~n13899;
  assign n13901 = n13898 & n13899;
  assign n13902 = ~n13900 & ~n13901;
  assign n13903 = n13888 & n13902;
  assign n13904 = ~n13888 & ~n13902;
  assign n13905 = ~n13903 & ~n13904;
  assign n13906 = n13625 & n13905;
  assign n13907 = ~n13625 & ~n13905;
  assign n13908 = ~n13906 & ~n13907;
  assign n13909 = ~n13556 & ~n13559;
  assign n13910 = pi120  & n750;
  assign n13911 = pi121  & n651;
  assign n13912 = pi122  & n646;
  assign n13913 = n644 & n10729;
  assign n13914 = ~n13911 & ~n13912;
  assign n13915 = ~n13910 & n13914;
  assign n13916 = ~n13913 & n13915;
  assign n13917 = pi11  & n13916;
  assign n13918 = ~pi11  & ~n13916;
  assign n13919 = ~n13917 & ~n13918;
  assign n13920 = ~n13909 & ~n13919;
  assign n13921 = n13909 & n13919;
  assign n13922 = ~n13920 & ~n13921;
  assign n13923 = n13908 & n13922;
  assign n13924 = ~n13908 & ~n13922;
  assign n13925 = ~n13923 & ~n13924;
  assign n13926 = pi123  & n528;
  assign n13927 = pi124  & n490;
  assign n13928 = pi125  & n485;
  assign n13929 = n483 & n11786;
  assign n13930 = ~n13927 & ~n13928;
  assign n13931 = ~n13926 & n13930;
  assign n13932 = ~n13929 & n13931;
  assign n13933 = pi8  & n13932;
  assign n13934 = ~pi8  & ~n13932;
  assign n13935 = ~n13933 & ~n13934;
  assign n13936 = ~n13269 & ~n13561;
  assign n13937 = ~n13268 & ~n13936;
  assign n13938 = ~n13935 & n13937;
  assign n13939 = n13935 & ~n13937;
  assign n13940 = ~n13938 & ~n13939;
  assign n13941 = n13925 & n13940;
  assign n13942 = ~n13925 & ~n13940;
  assign n13943 = ~n13941 & ~n13942;
  assign n13944 = ~n13577 & ~n13580;
  assign n13945 = pi126  & n391;
  assign n13946 = pi127  & n353;
  assign n13947 = n346 & n12542;
  assign n13948 = ~n13945 & ~n13946;
  assign n13949 = ~n13947 & n13948;
  assign n13950 = pi5  & n13949;
  assign n13951 = ~pi5  & ~n13949;
  assign n13952 = ~n13950 & ~n13951;
  assign n13953 = ~n13944 & ~n13952;
  assign n13954 = n13944 & n13952;
  assign n13955 = ~n13953 & ~n13954;
  assign n13956 = n13943 & n13955;
  assign n13957 = ~n13943 & ~n13955;
  assign n13958 = ~n13956 & ~n13957;
  assign n13959 = ~n13611 & n13958;
  assign n13960 = n13611 & ~n13958;
  assign n13961 = ~n13959 & ~n13960;
  assign n13962 = ~n13610 & n13961;
  assign n13963 = n13610 & ~n13961;
  assign po67  = ~n13962 & ~n13963;
  assign n13965 = ~n13959 & ~n13962;
  assign n13966 = ~n13953 & ~n13956;
  assign n13967 = pi121  & n750;
  assign n13968 = pi122  & n651;
  assign n13969 = pi123  & n646;
  assign n13970 = n644 & n10754;
  assign n13971 = ~n13968 & ~n13969;
  assign n13972 = ~n13967 & n13971;
  assign n13973 = ~n13970 & n13972;
  assign n13974 = pi11  & n13973;
  assign n13975 = ~pi11  & ~n13973;
  assign n13976 = ~n13974 & ~n13975;
  assign n13977 = ~n13624 & ~n13906;
  assign n13978 = n13976 & n13977;
  assign n13979 = ~n13976 & ~n13977;
  assign n13980 = ~n13978 & ~n13979;
  assign n13981 = ~n13638 & ~n13886;
  assign n13982 = pi115  & n1296;
  assign n13983 = pi116  & n1207;
  assign n13984 = pi117  & n1202;
  assign n13985 = n1200 & n8784;
  assign n13986 = ~n13983 & ~n13984;
  assign n13987 = ~n13982 & n13986;
  assign n13988 = ~n13985 & n13987;
  assign n13989 = pi17  & n13988;
  assign n13990 = ~pi17  & ~n13988;
  assign n13991 = ~n13989 & ~n13990;
  assign n13992 = ~n13981 & ~n13991;
  assign n13993 = n13981 & n13991;
  assign n13994 = ~n13992 & ~n13993;
  assign n13995 = pi109  & n2053;
  assign n13996 = pi110  & n1893;
  assign n13997 = pi111  & n1888;
  assign n13998 = n1886 & n7272;
  assign n13999 = ~n13996 & ~n13997;
  assign n14000 = ~n13995 & n13999;
  assign n14001 = ~n13998 & n14000;
  assign n14002 = pi23  & n14001;
  assign n14003 = ~pi23  & ~n14001;
  assign n14004 = ~n14002 & ~n14003;
  assign n14005 = ~n13652 & ~n13866;
  assign n14006 = n14004 & n14005;
  assign n14007 = ~n14004 & ~n14005;
  assign n14008 = ~n14006 & ~n14007;
  assign n14009 = ~n13860 & ~n13863;
  assign n14010 = pi106  & n2510;
  assign n14011 = pi107  & n2342;
  assign n14012 = pi108  & n2337;
  assign n14013 = n2335 & n6213;
  assign n14014 = ~n14011 & ~n14012;
  assign n14015 = ~n14010 & n14014;
  assign n14016 = ~n14013 & n14015;
  assign n14017 = pi26  & n14016;
  assign n14018 = ~pi26  & ~n14016;
  assign n14019 = ~n14017 & ~n14018;
  assign n14020 = ~n14009 & ~n14019;
  assign n14021 = n14009 & n14019;
  assign n14022 = ~n14020 & ~n14021;
  assign n14023 = pi103  & n3011;
  assign n14024 = pi104  & n2809;
  assign n14025 = pi105  & n2804;
  assign n14026 = n2802 & n5677;
  assign n14027 = ~n14024 & ~n14025;
  assign n14028 = ~n14023 & n14027;
  assign n14029 = ~n14026 & n14028;
  assign n14030 = pi29  & n14029;
  assign n14031 = ~pi29  & ~n14029;
  assign n14032 = ~n14030 & ~n14031;
  assign n14033 = ~n13666 & ~n13847;
  assign n14034 = n14032 & n14033;
  assign n14035 = ~n14032 & ~n14033;
  assign n14036 = ~n14034 & ~n14035;
  assign n14037 = pi100  & n3553;
  assign n14038 = pi101  & n3334;
  assign n14039 = pi102  & n3329;
  assign n14040 = n3327 & n4956;
  assign n14041 = ~n14038 & ~n14039;
  assign n14042 = ~n14037 & n14041;
  assign n14043 = ~n14040 & n14042;
  assign n14044 = pi32  & n14043;
  assign n14045 = ~pi32  & ~n14043;
  assign n14046 = ~n14044 & ~n14045;
  assign n14047 = n13678 & ~n13840;
  assign n14048 = ~n13841 & ~n14047;
  assign n14049 = ~n14046 & n14048;
  assign n14050 = n14046 & ~n14048;
  assign n14051 = ~n14049 & ~n14050;
  assign n14052 = ~n13806 & ~n13818;
  assign n14053 = ~n13807 & ~n14052;
  assign n14054 = ~n13798 & ~n13801;
  assign n14055 = ~n13747 & ~n13758;
  assign n14056 = ~n13746 & ~n14055;
  assign n14057 = pi79  & n8905;
  assign n14058 = pi80  & n8535;
  assign n14059 = pi81  & n8530;
  assign n14060 = n1337 & n8528;
  assign n14061 = ~n14058 & ~n14059;
  assign n14062 = ~n14057 & n14061;
  assign n14063 = ~n14060 & n14062;
  assign n14064 = pi53  & n14063;
  assign n14065 = ~pi53  & ~n14063;
  assign n14066 = ~n14064 & ~n14065;
  assign n14067 = ~n13730 & ~n13743;
  assign n14068 = ~n13705 & ~n13708;
  assign n14069 = pi70  & n11910;
  assign n14070 = pi71  & n11529;
  assign n14071 = pi72  & n11524;
  assign n14072 = n551 & n11522;
  assign n14073 = ~n14070 & ~n14071;
  assign n14074 = ~n14069 & n14073;
  assign n14075 = ~n14072 & n14074;
  assign n14076 = pi62  & n14075;
  assign n14077 = ~pi62  & ~n14075;
  assign n14078 = ~n14076 & ~n14077;
  assign n14079 = pi69  & n12277;
  assign n14080 = pi68  & n12276;
  assign n14081 = ~n14079 & ~n14080;
  assign n14082 = pi2  & ~n14081;
  assign n14083 = ~pi2  & n14081;
  assign n14084 = ~n14082 & ~n14083;
  assign n14085 = ~n14078 & n14084;
  assign n14086 = n14078 & ~n14084;
  assign n14087 = ~n14085 & ~n14086;
  assign n14088 = n14068 & ~n14087;
  assign n14089 = ~n14068 & n14087;
  assign n14090 = ~n14088 & ~n14089;
  assign n14091 = pi73  & n10886;
  assign n14092 = pi74  & n10495;
  assign n14093 = pi75  & n10490;
  assign n14094 = n713 & n10488;
  assign n14095 = ~n14092 & ~n14093;
  assign n14096 = ~n14091 & n14095;
  assign n14097 = ~n14094 & n14096;
  assign n14098 = pi59  & n14097;
  assign n14099 = ~pi59  & ~n14097;
  assign n14100 = ~n14098 & ~n14099;
  assign n14101 = ~n14090 & n14100;
  assign n14102 = n14090 & ~n14100;
  assign n14103 = ~n14101 & ~n14102;
  assign n14104 = ~n13712 & n13723;
  assign n14105 = ~n13711 & ~n14104;
  assign n14106 = n14103 & n14105;
  assign n14107 = ~n14103 & ~n14105;
  assign n14108 = ~n14106 & ~n14107;
  assign n14109 = pi76  & n9858;
  assign n14110 = pi77  & n9508;
  assign n14111 = pi78  & n9503;
  assign n14112 = n958 & n9501;
  assign n14113 = ~n14110 & ~n14111;
  assign n14114 = ~n14109 & n14113;
  assign n14115 = ~n14112 & n14114;
  assign n14116 = pi56  & n14115;
  assign n14117 = ~pi56  & ~n14115;
  assign n14118 = ~n14116 & ~n14117;
  assign n14119 = n14108 & ~n14118;
  assign n14120 = ~n14108 & n14118;
  assign n14121 = ~n14119 & ~n14120;
  assign n14122 = ~n14067 & n14121;
  assign n14123 = n14067 & ~n14121;
  assign n14124 = ~n14122 & ~n14123;
  assign n14125 = n14066 & ~n14124;
  assign n14126 = ~n14066 & n14124;
  assign n14127 = ~n14125 & ~n14126;
  assign n14128 = n14056 & ~n14127;
  assign n14129 = ~n14056 & n14127;
  assign n14130 = ~n14128 & ~n14129;
  assign n14131 = pi82  & n7969;
  assign n14132 = pi83  & n7636;
  assign n14133 = pi84  & n7631;
  assign n14134 = n1601 & n7629;
  assign n14135 = ~n14132 & ~n14133;
  assign n14136 = ~n14131 & n14135;
  assign n14137 = ~n14134 & n14136;
  assign n14138 = pi50  & n14137;
  assign n14139 = ~pi50  & ~n14137;
  assign n14140 = ~n14138 & ~n14139;
  assign n14141 = ~n14130 & n14140;
  assign n14142 = n14130 & ~n14140;
  assign n14143 = ~n14141 & ~n14142;
  assign n14144 = ~n13765 & n13776;
  assign n14145 = ~n13764 & ~n14144;
  assign n14146 = n14143 & n14145;
  assign n14147 = ~n14143 & ~n14145;
  assign n14148 = ~n14146 & ~n14147;
  assign n14149 = pi85  & n7121;
  assign n14150 = pi86  & n6795;
  assign n14151 = pi87  & n6790;
  assign n14152 = n2116 & n6788;
  assign n14153 = ~n14150 & ~n14151;
  assign n14154 = ~n14149 & n14153;
  assign n14155 = ~n14152 & n14154;
  assign n14156 = pi47  & n14155;
  assign n14157 = ~pi47  & ~n14155;
  assign n14158 = ~n14156 & ~n14157;
  assign n14159 = n14148 & ~n14158;
  assign n14160 = ~n14148 & n14158;
  assign n14161 = ~n14159 & ~n14160;
  assign n14162 = ~n13783 & n13794;
  assign n14163 = ~n13782 & ~n14162;
  assign n14164 = ~n14161 & ~n14163;
  assign n14165 = n14161 & n14163;
  assign n14166 = ~n14164 & ~n14165;
  assign n14167 = pi88  & n6331;
  assign n14168 = pi89  & n6015;
  assign n14169 = pi90  & n6010;
  assign n14170 = n2448 & n6008;
  assign n14171 = ~n14168 & ~n14169;
  assign n14172 = ~n14167 & n14171;
  assign n14173 = ~n14170 & n14172;
  assign n14174 = pi44  & n14173;
  assign n14175 = ~pi44  & ~n14173;
  assign n14176 = ~n14174 & ~n14175;
  assign n14177 = n14166 & ~n14176;
  assign n14178 = ~n14166 & n14176;
  assign n14179 = ~n14177 & ~n14178;
  assign n14180 = n14054 & ~n14179;
  assign n14181 = ~n14054 & n14179;
  assign n14182 = ~n14180 & ~n14181;
  assign n14183 = pi91  & n5558;
  assign n14184 = pi92  & n5293;
  assign n14185 = pi93  & n5288;
  assign n14186 = n2948 & n5286;
  assign n14187 = ~n14184 & ~n14185;
  assign n14188 = ~n14183 & n14187;
  assign n14189 = ~n14186 & n14188;
  assign n14190 = pi41  & n14189;
  assign n14191 = ~pi41  & ~n14189;
  assign n14192 = ~n14190 & ~n14191;
  assign n14193 = n14182 & ~n14192;
  assign n14194 = ~n14182 & n14192;
  assign n14195 = ~n14193 & ~n14194;
  assign n14196 = n14053 & ~n14195;
  assign n14197 = ~n14053 & n14195;
  assign n14198 = ~n14196 & ~n14197;
  assign n14199 = pi94  & n4843;
  assign n14200 = pi95  & n4598;
  assign n14201 = pi96  & n4593;
  assign n14202 = n3499 & n4591;
  assign n14203 = ~n14200 & ~n14201;
  assign n14204 = ~n14199 & n14203;
  assign n14205 = ~n14202 & n14204;
  assign n14206 = pi38  & n14205;
  assign n14207 = ~pi38  & ~n14205;
  assign n14208 = ~n14206 & ~n14207;
  assign n14209 = ~n14198 & n14208;
  assign n14210 = n14198 & ~n14208;
  assign n14211 = ~n14209 & ~n14210;
  assign n14212 = ~n13825 & ~n13838;
  assign n14213 = n14211 & ~n14212;
  assign n14214 = ~n14211 & n14212;
  assign n14215 = ~n14213 & ~n14214;
  assign n14216 = pi97  & n4176;
  assign n14217 = pi98  & n3938;
  assign n14218 = pi99  & n3933;
  assign n14219 = n3931 & n4101;
  assign n14220 = ~n14217 & ~n14218;
  assign n14221 = ~n14216 & n14220;
  assign n14222 = ~n14219 & n14221;
  assign n14223 = pi35  & n14222;
  assign n14224 = ~pi35  & ~n14222;
  assign n14225 = ~n14223 & ~n14224;
  assign n14226 = n14215 & ~n14225;
  assign n14227 = ~n14215 & n14225;
  assign n14228 = ~n14226 & ~n14227;
  assign n14229 = n14051 & n14228;
  assign n14230 = ~n14051 & ~n14228;
  assign n14231 = ~n14229 & ~n14230;
  assign n14232 = n14036 & n14231;
  assign n14233 = ~n14036 & ~n14231;
  assign n14234 = ~n14232 & ~n14233;
  assign n14235 = n14022 & n14234;
  assign n14236 = ~n14022 & ~n14234;
  assign n14237 = ~n14235 & ~n14236;
  assign n14238 = n14008 & n14237;
  assign n14239 = ~n14008 & ~n14237;
  assign n14240 = ~n14238 & ~n14239;
  assign n14241 = pi112  & n1661;
  assign n14242 = pi113  & n1500;
  assign n14243 = pi114  & n1495;
  assign n14244 = n1493 & n8146;
  assign n14245 = ~n14242 & ~n14243;
  assign n14246 = ~n14241 & n14245;
  assign n14247 = ~n14244 & n14246;
  assign n14248 = pi20  & n14247;
  assign n14249 = ~pi20  & ~n14247;
  assign n14250 = ~n14248 & ~n14249;
  assign n14251 = ~n13880 & ~n13883;
  assign n14252 = ~n14250 & ~n14251;
  assign n14253 = n14250 & n14251;
  assign n14254 = ~n14252 & ~n14253;
  assign n14255 = n14240 & n14254;
  assign n14256 = ~n14240 & ~n14254;
  assign n14257 = ~n14255 & ~n14256;
  assign n14258 = n13994 & n14257;
  assign n14259 = ~n13994 & ~n14257;
  assign n14260 = ~n14258 & ~n14259;
  assign n14261 = pi118  & n1006;
  assign n14262 = pi119  & n897;
  assign n14263 = pi120  & n892;
  assign n14264 = n890 & n10047;
  assign n14265 = ~n14262 & ~n14263;
  assign n14266 = ~n14261 & n14265;
  assign n14267 = ~n14264 & n14266;
  assign n14268 = pi14  & n14267;
  assign n14269 = ~pi14  & ~n14267;
  assign n14270 = ~n14268 & ~n14269;
  assign n14271 = ~n13900 & ~n13903;
  assign n14272 = ~n14270 & ~n14271;
  assign n14273 = n14270 & n14271;
  assign n14274 = ~n14272 & ~n14273;
  assign n14275 = n14260 & n14274;
  assign n14276 = ~n14260 & ~n14274;
  assign n14277 = ~n14275 & ~n14276;
  assign n14278 = n13980 & n14277;
  assign n14279 = ~n13980 & ~n14277;
  assign n14280 = ~n14278 & ~n14279;
  assign n14281 = ~n13920 & ~n13923;
  assign n14282 = pi124  & n528;
  assign n14283 = pi125  & n490;
  assign n14284 = pi126  & n485;
  assign n14285 = n483 & n12148;
  assign n14286 = ~n14283 & ~n14284;
  assign n14287 = ~n14282 & n14286;
  assign n14288 = ~n14285 & n14287;
  assign n14289 = pi8  & n14288;
  assign n14290 = ~pi8  & ~n14288;
  assign n14291 = ~n14289 & ~n14290;
  assign n14292 = ~n14281 & ~n14291;
  assign n14293 = n14281 & n14291;
  assign n14294 = ~n14292 & ~n14293;
  assign n14295 = n14280 & n14294;
  assign n14296 = ~n14280 & ~n14294;
  assign n14297 = ~n14295 & ~n14296;
  assign n14298 = ~n13938 & ~n13941;
  assign n14299 = n346 & ~n12539;
  assign n14300 = ~n391 & ~n14299;
  assign n14301 = pi127  & ~n14300;
  assign n14302 = pi5  & ~n14301;
  assign n14303 = ~pi5  & n14301;
  assign n14304 = ~n14302 & ~n14303;
  assign n14305 = ~n14298 & ~n14304;
  assign n14306 = n14298 & n14304;
  assign n14307 = ~n14305 & ~n14306;
  assign n14308 = n14297 & n14307;
  assign n14309 = ~n14297 & ~n14307;
  assign n14310 = ~n14308 & ~n14309;
  assign n14311 = ~n13966 & n14310;
  assign n14312 = n13966 & ~n14310;
  assign n14313 = ~n14311 & ~n14312;
  assign n14314 = ~n13965 & n14313;
  assign n14315 = n13965 & ~n14313;
  assign po68  = ~n14314 & ~n14315;
  assign n14317 = ~n14311 & ~n14314;
  assign n14318 = ~n14305 & ~n14308;
  assign n14319 = ~n14292 & ~n14295;
  assign n14320 = pi125  & n528;
  assign n14321 = pi126  & n490;
  assign n14322 = pi127  & n485;
  assign n14323 = n483 & n12519;
  assign n14324 = ~n14321 & ~n14322;
  assign n14325 = ~n14320 & n14324;
  assign n14326 = ~n14323 & n14325;
  assign n14327 = pi8  & n14326;
  assign n14328 = ~pi8  & ~n14326;
  assign n14329 = ~n14327 & ~n14328;
  assign n14330 = ~n14319 & ~n14329;
  assign n14331 = n14319 & n14329;
  assign n14332 = ~n14330 & ~n14331;
  assign n14333 = pi122  & n750;
  assign n14334 = pi123  & n651;
  assign n14335 = pi124  & n646;
  assign n14336 = n644 & n11099;
  assign n14337 = ~n14334 & ~n14335;
  assign n14338 = ~n14333 & n14337;
  assign n14339 = ~n14336 & n14338;
  assign n14340 = pi11  & n14339;
  assign n14341 = ~pi11  & ~n14339;
  assign n14342 = ~n14340 & ~n14341;
  assign n14343 = ~n13979 & ~n14278;
  assign n14344 = n14342 & n14343;
  assign n14345 = ~n14342 & ~n14343;
  assign n14346 = ~n14344 & ~n14345;
  assign n14347 = pi119  & n1006;
  assign n14348 = pi120  & n897;
  assign n14349 = pi121  & n892;
  assign n14350 = n890 & n10071;
  assign n14351 = ~n14348 & ~n14349;
  assign n14352 = ~n14347 & n14351;
  assign n14353 = ~n14350 & n14352;
  assign n14354 = pi14  & n14353;
  assign n14355 = ~pi14  & ~n14353;
  assign n14356 = ~n14354 & ~n14355;
  assign n14357 = ~n14272 & ~n14275;
  assign n14358 = ~n14356 & ~n14357;
  assign n14359 = n14356 & n14357;
  assign n14360 = ~n14358 & ~n14359;
  assign n14361 = pi113  & n1661;
  assign n14362 = pi114  & n1500;
  assign n14363 = pi115  & n1495;
  assign n14364 = n1493 & n8170;
  assign n14365 = ~n14362 & ~n14363;
  assign n14366 = ~n14361 & n14365;
  assign n14367 = ~n14364 & n14366;
  assign n14368 = pi20  & n14367;
  assign n14369 = ~pi20  & ~n14367;
  assign n14370 = ~n14368 & ~n14369;
  assign n14371 = ~n14252 & ~n14255;
  assign n14372 = ~n14370 & ~n14371;
  assign n14373 = n14370 & n14371;
  assign n14374 = ~n14372 & ~n14373;
  assign n14375 = pi110  & n2053;
  assign n14376 = pi111  & n1893;
  assign n14377 = pi112  & n1888;
  assign n14378 = n1886 & n7296;
  assign n14379 = ~n14376 & ~n14377;
  assign n14380 = ~n14375 & n14379;
  assign n14381 = ~n14378 & n14380;
  assign n14382 = pi23  & n14381;
  assign n14383 = ~pi23  & ~n14381;
  assign n14384 = ~n14382 & ~n14383;
  assign n14385 = ~n14007 & ~n14238;
  assign n14386 = n14384 & n14385;
  assign n14387 = ~n14384 & ~n14385;
  assign n14388 = ~n14386 & ~n14387;
  assign n14389 = pi104  & n3011;
  assign n14390 = pi105  & n2809;
  assign n14391 = pi106  & n2804;
  assign n14392 = n2802 & n5701;
  assign n14393 = ~n14390 & ~n14391;
  assign n14394 = ~n14389 & n14393;
  assign n14395 = ~n14392 & n14394;
  assign n14396 = pi29  & n14395;
  assign n14397 = ~pi29  & ~n14395;
  assign n14398 = ~n14396 & ~n14397;
  assign n14399 = ~n14035 & ~n14231;
  assign n14400 = ~n14034 & ~n14399;
  assign n14401 = n14398 & ~n14400;
  assign n14402 = ~n14398 & n14400;
  assign n14403 = ~n14401 & ~n14402;
  assign n14404 = pi98  & n4176;
  assign n14405 = pi99  & n3938;
  assign n14406 = pi100  & n3933;
  assign n14407 = n3931 & n4501;
  assign n14408 = ~n14405 & ~n14406;
  assign n14409 = ~n14404 & n14408;
  assign n14410 = ~n14407 & n14409;
  assign n14411 = pi35  & n14410;
  assign n14412 = ~pi35  & ~n14410;
  assign n14413 = ~n14411 & ~n14412;
  assign n14414 = ~n14197 & ~n14210;
  assign n14415 = pi95  & n4843;
  assign n14416 = pi96  & n4598;
  assign n14417 = pi97  & n4593;
  assign n14418 = n3691 & n4591;
  assign n14419 = ~n14416 & ~n14417;
  assign n14420 = ~n14415 & n14419;
  assign n14421 = ~n14418 & n14420;
  assign n14422 = pi38  & n14421;
  assign n14423 = ~pi38  & ~n14421;
  assign n14424 = ~n14422 & ~n14423;
  assign n14425 = pi86  & n7121;
  assign n14426 = pi87  & n6795;
  assign n14427 = pi88  & n6790;
  assign n14428 = n2140 & n6788;
  assign n14429 = ~n14426 & ~n14427;
  assign n14430 = ~n14425 & n14429;
  assign n14431 = ~n14428 & n14430;
  assign n14432 = pi47  & n14431;
  assign n14433 = ~pi47  & ~n14431;
  assign n14434 = ~n14432 & ~n14433;
  assign n14435 = ~n14129 & ~n14142;
  assign n14436 = pi77  & n9858;
  assign n14437 = pi78  & n9508;
  assign n14438 = pi79  & n9503;
  assign n14439 = n1048 & n9501;
  assign n14440 = ~n14437 & ~n14438;
  assign n14441 = ~n14436 & n14440;
  assign n14442 = ~n14439 & n14441;
  assign n14443 = pi56  & n14442;
  assign n14444 = ~pi56  & ~n14442;
  assign n14445 = ~n14443 & ~n14444;
  assign n14446 = ~n14089 & ~n14102;
  assign n14447 = pi74  & n10886;
  assign n14448 = pi75  & n10495;
  assign n14449 = pi76  & n10490;
  assign n14450 = n841 & n10488;
  assign n14451 = ~n14448 & ~n14449;
  assign n14452 = ~n14447 & n14451;
  assign n14453 = ~n14450 & n14452;
  assign n14454 = pi59  & n14453;
  assign n14455 = ~pi59  & ~n14453;
  assign n14456 = ~n14454 & ~n14455;
  assign n14457 = ~n14082 & ~n14085;
  assign n14458 = ~pi2  & ~pi5 ;
  assign n14459 = pi2  & pi5 ;
  assign n14460 = ~n14458 & ~n14459;
  assign n14461 = pi70  & n12277;
  assign n14462 = pi69  & n12276;
  assign n14463 = ~n14461 & ~n14462;
  assign n14464 = n14460 & ~n14463;
  assign n14465 = ~n14460 & n14463;
  assign n14466 = ~n14464 & ~n14465;
  assign n14467 = n14457 & ~n14466;
  assign n14468 = ~n14457 & n14466;
  assign n14469 = ~n14467 & ~n14468;
  assign n14470 = pi71  & n11910;
  assign n14471 = pi72  & n11529;
  assign n14472 = pi73  & n11524;
  assign n14473 = n613 & n11522;
  assign n14474 = ~n14471 & ~n14472;
  assign n14475 = ~n14470 & n14474;
  assign n14476 = ~n14473 & n14475;
  assign n14477 = pi62  & n14476;
  assign n14478 = ~pi62  & ~n14476;
  assign n14479 = ~n14477 & ~n14478;
  assign n14480 = ~n14469 & n14479;
  assign n14481 = n14469 & ~n14479;
  assign n14482 = ~n14480 & ~n14481;
  assign n14483 = ~n14456 & n14482;
  assign n14484 = n14456 & ~n14482;
  assign n14485 = ~n14483 & ~n14484;
  assign n14486 = ~n14446 & n14485;
  assign n14487 = n14446 & ~n14485;
  assign n14488 = ~n14486 & ~n14487;
  assign n14489 = ~n14445 & n14488;
  assign n14490 = n14445 & ~n14488;
  assign n14491 = ~n14489 & ~n14490;
  assign n14492 = ~n14106 & n14118;
  assign n14493 = ~n14107 & ~n14492;
  assign n14494 = ~n14491 & ~n14493;
  assign n14495 = n14491 & n14493;
  assign n14496 = ~n14494 & ~n14495;
  assign n14497 = pi80  & n8905;
  assign n14498 = pi81  & n8535;
  assign n14499 = pi82  & n8530;
  assign n14500 = n1450 & n8528;
  assign n14501 = ~n14498 & ~n14499;
  assign n14502 = ~n14497 & n14501;
  assign n14503 = ~n14500 & n14502;
  assign n14504 = pi53  & n14503;
  assign n14505 = ~pi53  & ~n14503;
  assign n14506 = ~n14504 & ~n14505;
  assign n14507 = n14496 & ~n14506;
  assign n14508 = ~n14496 & n14506;
  assign n14509 = ~n14507 & ~n14508;
  assign n14510 = n14066 & ~n14122;
  assign n14511 = ~n14123 & ~n14510;
  assign n14512 = ~n14509 & ~n14511;
  assign n14513 = n14509 & n14511;
  assign n14514 = ~n14512 & ~n14513;
  assign n14515 = pi83  & n7969;
  assign n14516 = pi84  & n7636;
  assign n14517 = pi85  & n7631;
  assign n14518 = n1831 & n7629;
  assign n14519 = ~n14516 & ~n14517;
  assign n14520 = ~n14515 & n14519;
  assign n14521 = ~n14518 & n14520;
  assign n14522 = pi50  & n14521;
  assign n14523 = ~pi50  & ~n14521;
  assign n14524 = ~n14522 & ~n14523;
  assign n14525 = n14514 & ~n14524;
  assign n14526 = ~n14514 & n14524;
  assign n14527 = ~n14525 & ~n14526;
  assign n14528 = ~n14435 & n14527;
  assign n14529 = n14435 & ~n14527;
  assign n14530 = ~n14528 & ~n14529;
  assign n14531 = ~n14434 & n14530;
  assign n14532 = n14434 & ~n14530;
  assign n14533 = ~n14531 & ~n14532;
  assign n14534 = ~n14146 & n14158;
  assign n14535 = ~n14147 & ~n14534;
  assign n14536 = ~n14533 & ~n14535;
  assign n14537 = n14533 & n14535;
  assign n14538 = ~n14536 & ~n14537;
  assign n14539 = pi89  & n6331;
  assign n14540 = pi90  & n6015;
  assign n14541 = pi91  & n6010;
  assign n14542 = n2746 & n6008;
  assign n14543 = ~n14540 & ~n14541;
  assign n14544 = ~n14539 & n14543;
  assign n14545 = ~n14542 & n14544;
  assign n14546 = pi44  & n14545;
  assign n14547 = ~pi44  & ~n14545;
  assign n14548 = ~n14546 & ~n14547;
  assign n14549 = n14538 & ~n14548;
  assign n14550 = ~n14538 & n14548;
  assign n14551 = ~n14549 & ~n14550;
  assign n14552 = ~n14165 & n14176;
  assign n14553 = ~n14164 & ~n14552;
  assign n14554 = ~n14551 & ~n14553;
  assign n14555 = n14551 & n14553;
  assign n14556 = ~n14554 & ~n14555;
  assign n14557 = pi92  & n5558;
  assign n14558 = pi93  & n5293;
  assign n14559 = pi94  & n5288;
  assign n14560 = n3280 & n5286;
  assign n14561 = ~n14558 & ~n14559;
  assign n14562 = ~n14557 & n14561;
  assign n14563 = ~n14560 & n14562;
  assign n14564 = pi41  & n14563;
  assign n14565 = ~pi41  & ~n14563;
  assign n14566 = ~n14564 & ~n14565;
  assign n14567 = n14556 & ~n14566;
  assign n14568 = ~n14556 & n14566;
  assign n14569 = ~n14567 & ~n14568;
  assign n14570 = ~n14181 & n14192;
  assign n14571 = ~n14180 & ~n14570;
  assign n14572 = n14569 & ~n14571;
  assign n14573 = ~n14569 & n14571;
  assign n14574 = ~n14572 & ~n14573;
  assign n14575 = ~n14424 & ~n14574;
  assign n14576 = n14424 & n14574;
  assign n14577 = ~n14575 & ~n14576;
  assign n14578 = ~n14414 & n14577;
  assign n14579 = n14414 & ~n14577;
  assign n14580 = ~n14578 & ~n14579;
  assign n14581 = ~n14413 & n14580;
  assign n14582 = n14413 & ~n14580;
  assign n14583 = ~n14581 & ~n14582;
  assign n14584 = ~n14214 & ~n14225;
  assign n14585 = ~n14213 & ~n14584;
  assign n14586 = ~n14583 & n14585;
  assign n14587 = n14583 & ~n14585;
  assign n14588 = ~n14586 & ~n14587;
  assign n14589 = pi101  & n3553;
  assign n14590 = pi102  & n3334;
  assign n14591 = pi103  & n3329;
  assign n14592 = n3327 & n5188;
  assign n14593 = ~n14590 & ~n14591;
  assign n14594 = ~n14589 & n14593;
  assign n14595 = ~n14592 & n14594;
  assign n14596 = pi32  & n14595;
  assign n14597 = ~pi32  & ~n14595;
  assign n14598 = ~n14596 & ~n14597;
  assign n14599 = ~n14049 & ~n14228;
  assign n14600 = ~n14050 & ~n14599;
  assign n14601 = n14598 & ~n14600;
  assign n14602 = ~n14598 & n14600;
  assign n14603 = ~n14601 & ~n14602;
  assign n14604 = n14588 & n14603;
  assign n14605 = ~n14588 & ~n14603;
  assign n14606 = ~n14604 & ~n14605;
  assign n14607 = n14403 & n14606;
  assign n14608 = ~n14403 & ~n14606;
  assign n14609 = ~n14607 & ~n14608;
  assign n14610 = ~n14020 & ~n14235;
  assign n14611 = pi107  & n2510;
  assign n14612 = pi108  & n2342;
  assign n14613 = pi109  & n2337;
  assign n14614 = n2335 & n6715;
  assign n14615 = ~n14612 & ~n14613;
  assign n14616 = ~n14611 & n14615;
  assign n14617 = ~n14614 & n14616;
  assign n14618 = pi26  & n14617;
  assign n14619 = ~pi26  & ~n14617;
  assign n14620 = ~n14618 & ~n14619;
  assign n14621 = ~n14610 & ~n14620;
  assign n14622 = n14610 & n14620;
  assign n14623 = ~n14621 & ~n14622;
  assign n14624 = n14609 & n14623;
  assign n14625 = ~n14609 & ~n14623;
  assign n14626 = ~n14624 & ~n14625;
  assign n14627 = n14388 & n14626;
  assign n14628 = ~n14388 & ~n14626;
  assign n14629 = ~n14627 & ~n14628;
  assign n14630 = n14374 & n14629;
  assign n14631 = ~n14374 & ~n14629;
  assign n14632 = ~n14630 & ~n14631;
  assign n14633 = ~n13992 & ~n14258;
  assign n14634 = pi116  & n1296;
  assign n14635 = pi117  & n1207;
  assign n14636 = pi118  & n1202;
  assign n14637 = n1200 & n9095;
  assign n14638 = ~n14635 & ~n14636;
  assign n14639 = ~n14634 & n14638;
  assign n14640 = ~n14637 & n14639;
  assign n14641 = pi17  & n14640;
  assign n14642 = ~pi17  & ~n14640;
  assign n14643 = ~n14641 & ~n14642;
  assign n14644 = ~n14633 & ~n14643;
  assign n14645 = n14633 & n14643;
  assign n14646 = ~n14644 & ~n14645;
  assign n14647 = n14632 & n14646;
  assign n14648 = ~n14632 & ~n14646;
  assign n14649 = ~n14647 & ~n14648;
  assign n14650 = ~n14360 & n14649;
  assign n14651 = n14360 & ~n14649;
  assign n14652 = ~n14650 & ~n14651;
  assign n14653 = n14346 & ~n14652;
  assign n14654 = ~n14346 & n14652;
  assign n14655 = ~n14653 & ~n14654;
  assign n14656 = n14332 & n14655;
  assign n14657 = ~n14332 & ~n14655;
  assign n14658 = ~n14656 & ~n14657;
  assign n14659 = ~n14318 & n14658;
  assign n14660 = n14318 & ~n14658;
  assign n14661 = ~n14659 & ~n14660;
  assign n14662 = ~n14317 & n14661;
  assign n14663 = n14317 & ~n14661;
  assign po69  = ~n14662 & ~n14663;
  assign n14665 = ~n14659 & ~n14662;
  assign n14666 = ~n14330 & ~n14656;
  assign n14667 = pi126  & n528;
  assign n14668 = pi127  & n490;
  assign n14669 = n483 & n12542;
  assign n14670 = ~n14667 & ~n14668;
  assign n14671 = ~n14669 & n14670;
  assign n14672 = pi8  & n14671;
  assign n14673 = ~pi8  & ~n14671;
  assign n14674 = ~n14672 & ~n14673;
  assign n14675 = ~n14345 & n14652;
  assign n14676 = ~n14344 & ~n14675;
  assign n14677 = ~n14674 & n14676;
  assign n14678 = n14674 & ~n14676;
  assign n14679 = ~n14677 & ~n14678;
  assign n14680 = pi123  & n750;
  assign n14681 = pi124  & n651;
  assign n14682 = pi125  & n646;
  assign n14683 = n644 & n11786;
  assign n14684 = ~n14681 & ~n14682;
  assign n14685 = ~n14680 & n14684;
  assign n14686 = ~n14683 & n14685;
  assign n14687 = pi11  & n14686;
  assign n14688 = ~pi11  & ~n14686;
  assign n14689 = ~n14687 & ~n14688;
  assign n14690 = ~n14358 & ~n14649;
  assign n14691 = ~n14359 & ~n14690;
  assign n14692 = n14689 & ~n14691;
  assign n14693 = ~n14689 & n14691;
  assign n14694 = ~n14692 & ~n14693;
  assign n14695 = ~n14644 & ~n14647;
  assign n14696 = pi120  & n1006;
  assign n14697 = pi121  & n897;
  assign n14698 = pi122  & n892;
  assign n14699 = n890 & n10729;
  assign n14700 = ~n14697 & ~n14698;
  assign n14701 = ~n14696 & n14700;
  assign n14702 = ~n14699 & n14701;
  assign n14703 = pi14  & n14702;
  assign n14704 = ~pi14  & ~n14702;
  assign n14705 = ~n14703 & ~n14704;
  assign n14706 = ~n14695 & ~n14705;
  assign n14707 = n14695 & n14705;
  assign n14708 = ~n14706 & ~n14707;
  assign n14709 = pi117  & n1296;
  assign n14710 = pi118  & n1207;
  assign n14711 = pi119  & n1202;
  assign n14712 = n1200 & n9412;
  assign n14713 = ~n14710 & ~n14711;
  assign n14714 = ~n14709 & n14713;
  assign n14715 = ~n14712 & n14714;
  assign n14716 = pi17  & n14715;
  assign n14717 = ~pi17  & ~n14715;
  assign n14718 = ~n14716 & ~n14717;
  assign n14719 = ~n14372 & ~n14630;
  assign n14720 = n14718 & n14719;
  assign n14721 = ~n14718 & ~n14719;
  assign n14722 = ~n14720 & ~n14721;
  assign n14723 = pi114  & n1661;
  assign n14724 = pi115  & n1500;
  assign n14725 = pi116  & n1495;
  assign n14726 = n1493 & n8470;
  assign n14727 = ~n14724 & ~n14725;
  assign n14728 = ~n14723 & n14727;
  assign n14729 = ~n14726 & n14728;
  assign n14730 = pi20  & n14729;
  assign n14731 = ~pi20  & ~n14729;
  assign n14732 = ~n14730 & ~n14731;
  assign n14733 = ~n14387 & ~n14627;
  assign n14734 = n14732 & n14733;
  assign n14735 = ~n14732 & ~n14733;
  assign n14736 = ~n14734 & ~n14735;
  assign n14737 = ~n14402 & ~n14607;
  assign n14738 = pi108  & n2510;
  assign n14739 = pi109  & n2342;
  assign n14740 = pi110  & n2337;
  assign n14741 = n2335 & n6995;
  assign n14742 = ~n14739 & ~n14740;
  assign n14743 = ~n14738 & n14742;
  assign n14744 = ~n14741 & n14743;
  assign n14745 = pi26  & n14744;
  assign n14746 = ~pi26  & ~n14744;
  assign n14747 = ~n14745 & ~n14746;
  assign n14748 = ~n14737 & ~n14747;
  assign n14749 = n14737 & n14747;
  assign n14750 = ~n14748 & ~n14749;
  assign n14751 = pi105  & n3011;
  assign n14752 = pi106  & n2809;
  assign n14753 = pi107  & n2804;
  assign n14754 = n2802 & n6189;
  assign n14755 = ~n14752 & ~n14753;
  assign n14756 = ~n14751 & n14755;
  assign n14757 = ~n14754 & n14756;
  assign n14758 = pi29  & n14757;
  assign n14759 = ~pi29  & ~n14757;
  assign n14760 = ~n14758 & ~n14759;
  assign n14761 = ~n14602 & ~n14604;
  assign n14762 = ~n14760 & ~n14761;
  assign n14763 = n14760 & n14761;
  assign n14764 = ~n14762 & ~n14763;
  assign n14765 = pi102  & n3553;
  assign n14766 = pi103  & n3334;
  assign n14767 = pi104  & n3329;
  assign n14768 = n3327 & n5212;
  assign n14769 = ~n14766 & ~n14767;
  assign n14770 = ~n14765 & n14769;
  assign n14771 = ~n14768 & n14770;
  assign n14772 = pi32  & n14771;
  assign n14773 = ~pi32  & ~n14771;
  assign n14774 = ~n14772 & ~n14773;
  assign n14775 = ~n14581 & ~n14587;
  assign n14776 = n14774 & n14775;
  assign n14777 = ~n14774 & ~n14775;
  assign n14778 = ~n14776 & ~n14777;
  assign n14779 = pi99  & n4176;
  assign n14780 = pi100  & n3938;
  assign n14781 = pi101  & n3933;
  assign n14782 = n3931 & n4730;
  assign n14783 = ~n14780 & ~n14781;
  assign n14784 = ~n14779 & n14783;
  assign n14785 = ~n14782 & n14784;
  assign n14786 = pi35  & n14785;
  assign n14787 = ~pi35  & ~n14785;
  assign n14788 = ~n14786 & ~n14787;
  assign n14789 = ~n14575 & ~n14578;
  assign n14790 = pi96  & n4843;
  assign n14791 = pi97  & n4598;
  assign n14792 = pi98  & n4593;
  assign n14793 = n3889 & n4591;
  assign n14794 = ~n14791 & ~n14792;
  assign n14795 = ~n14790 & n14794;
  assign n14796 = ~n14793 & n14795;
  assign n14797 = pi38  & n14796;
  assign n14798 = ~pi38  & ~n14796;
  assign n14799 = ~n14797 & ~n14798;
  assign n14800 = ~n14549 & ~n14555;
  assign n14801 = ~n14531 & ~n14537;
  assign n14802 = ~n14525 & ~n14528;
  assign n14803 = ~n14507 & ~n14513;
  assign n14804 = ~n14489 & ~n14495;
  assign n14805 = ~n14483 & ~n14486;
  assign n14806 = ~n14468 & ~n14481;
  assign n14807 = ~n14458 & ~n14464;
  assign n14808 = pi71  & n12277;
  assign n14809 = pi70  & n12276;
  assign n14810 = ~n14808 & ~n14809;
  assign n14811 = ~n14807 & n14810;
  assign n14812 = n14807 & ~n14810;
  assign n14813 = ~n14811 & ~n14812;
  assign n14814 = pi72  & n11910;
  assign n14815 = pi73  & n11529;
  assign n14816 = pi74  & n11524;
  assign n14817 = n689 & n11522;
  assign n14818 = ~n14815 & ~n14816;
  assign n14819 = ~n14814 & n14818;
  assign n14820 = ~n14817 & n14819;
  assign n14821 = pi62  & n14820;
  assign n14822 = ~pi62  & ~n14820;
  assign n14823 = ~n14821 & ~n14822;
  assign n14824 = n14813 & ~n14823;
  assign n14825 = ~n14813 & n14823;
  assign n14826 = ~n14824 & ~n14825;
  assign n14827 = ~n14806 & n14826;
  assign n14828 = n14806 & ~n14826;
  assign n14829 = ~n14827 & ~n14828;
  assign n14830 = pi75  & n10886;
  assign n14831 = pi76  & n10495;
  assign n14832 = pi77  & n10490;
  assign n14833 = n865 & n10488;
  assign n14834 = ~n14831 & ~n14832;
  assign n14835 = ~n14830 & n14834;
  assign n14836 = ~n14833 & n14835;
  assign n14837 = pi59  & n14836;
  assign n14838 = ~pi59  & ~n14836;
  assign n14839 = ~n14837 & ~n14838;
  assign n14840 = n14829 & ~n14839;
  assign n14841 = ~n14829 & n14839;
  assign n14842 = ~n14840 & ~n14841;
  assign n14843 = n14805 & ~n14842;
  assign n14844 = ~n14805 & n14842;
  assign n14845 = ~n14843 & ~n14844;
  assign n14846 = pi78  & n9858;
  assign n14847 = pi79  & n9508;
  assign n14848 = pi80  & n9503;
  assign n14849 = n1144 & n9501;
  assign n14850 = ~n14847 & ~n14848;
  assign n14851 = ~n14846 & n14850;
  assign n14852 = ~n14849 & n14851;
  assign n14853 = pi56  & n14852;
  assign n14854 = ~pi56  & ~n14852;
  assign n14855 = ~n14853 & ~n14854;
  assign n14856 = n14845 & ~n14855;
  assign n14857 = ~n14845 & n14855;
  assign n14858 = ~n14856 & ~n14857;
  assign n14859 = n14804 & ~n14858;
  assign n14860 = ~n14804 & n14858;
  assign n14861 = ~n14859 & ~n14860;
  assign n14862 = pi81  & n8905;
  assign n14863 = pi82  & n8535;
  assign n14864 = pi83  & n8530;
  assign n14865 = n1577 & n8528;
  assign n14866 = ~n14863 & ~n14864;
  assign n14867 = ~n14862 & n14866;
  assign n14868 = ~n14865 & n14867;
  assign n14869 = pi53  & n14868;
  assign n14870 = ~pi53  & ~n14868;
  assign n14871 = ~n14869 & ~n14870;
  assign n14872 = n14861 & ~n14871;
  assign n14873 = ~n14861 & n14871;
  assign n14874 = ~n14872 & ~n14873;
  assign n14875 = n14803 & ~n14874;
  assign n14876 = ~n14803 & n14874;
  assign n14877 = ~n14875 & ~n14876;
  assign n14878 = pi84  & n7969;
  assign n14879 = pi85  & n7636;
  assign n14880 = pi86  & n7631;
  assign n14881 = n1975 & n7629;
  assign n14882 = ~n14879 & ~n14880;
  assign n14883 = ~n14878 & n14882;
  assign n14884 = ~n14881 & n14883;
  assign n14885 = pi50  & n14884;
  assign n14886 = ~pi50  & ~n14884;
  assign n14887 = ~n14885 & ~n14886;
  assign n14888 = n14877 & ~n14887;
  assign n14889 = ~n14877 & n14887;
  assign n14890 = ~n14888 & ~n14889;
  assign n14891 = n14802 & ~n14890;
  assign n14892 = ~n14802 & n14890;
  assign n14893 = ~n14891 & ~n14892;
  assign n14894 = pi87  & n7121;
  assign n14895 = pi88  & n6795;
  assign n14896 = pi89  & n6790;
  assign n14897 = n2287 & n6788;
  assign n14898 = ~n14895 & ~n14896;
  assign n14899 = ~n14894 & n14898;
  assign n14900 = ~n14897 & n14899;
  assign n14901 = pi47  & n14900;
  assign n14902 = ~pi47  & ~n14900;
  assign n14903 = ~n14901 & ~n14902;
  assign n14904 = n14893 & ~n14903;
  assign n14905 = ~n14893 & n14903;
  assign n14906 = ~n14904 & ~n14905;
  assign n14907 = n14801 & ~n14906;
  assign n14908 = ~n14801 & n14906;
  assign n14909 = ~n14907 & ~n14908;
  assign n14910 = pi90  & n6331;
  assign n14911 = pi91  & n6015;
  assign n14912 = pi92  & n6010;
  assign n14913 = n2924 & n6008;
  assign n14914 = ~n14911 & ~n14912;
  assign n14915 = ~n14910 & n14914;
  assign n14916 = ~n14913 & n14915;
  assign n14917 = pi44  & n14916;
  assign n14918 = ~pi44  & ~n14916;
  assign n14919 = ~n14917 & ~n14918;
  assign n14920 = n14909 & ~n14919;
  assign n14921 = ~n14909 & n14919;
  assign n14922 = ~n14920 & ~n14921;
  assign n14923 = n14800 & ~n14922;
  assign n14924 = ~n14800 & n14922;
  assign n14925 = ~n14923 & ~n14924;
  assign n14926 = pi93  & n5558;
  assign n14927 = pi94  & n5293;
  assign n14928 = pi95  & n5288;
  assign n14929 = n3475 & n5286;
  assign n14930 = ~n14927 & ~n14928;
  assign n14931 = ~n14926 & n14930;
  assign n14932 = ~n14929 & n14931;
  assign n14933 = pi41  & n14932;
  assign n14934 = ~pi41  & ~n14932;
  assign n14935 = ~n14933 & ~n14934;
  assign n14936 = ~n14925 & n14935;
  assign n14937 = n14925 & ~n14935;
  assign n14938 = ~n14936 & ~n14937;
  assign n14939 = ~n14567 & ~n14571;
  assign n14940 = ~n14568 & ~n14939;
  assign n14941 = n14938 & n14940;
  assign n14942 = ~n14938 & ~n14940;
  assign n14943 = ~n14941 & ~n14942;
  assign n14944 = ~n14799 & n14943;
  assign n14945 = n14799 & ~n14943;
  assign n14946 = ~n14944 & ~n14945;
  assign n14947 = ~n14789 & n14946;
  assign n14948 = n14789 & ~n14946;
  assign n14949 = ~n14947 & ~n14948;
  assign n14950 = n14788 & ~n14949;
  assign n14951 = ~n14788 & n14949;
  assign n14952 = ~n14950 & ~n14951;
  assign n14953 = n14778 & n14952;
  assign n14954 = ~n14778 & ~n14952;
  assign n14955 = ~n14953 & ~n14954;
  assign n14956 = n14764 & n14955;
  assign n14957 = ~n14764 & ~n14955;
  assign n14958 = ~n14956 & ~n14957;
  assign n14959 = n14750 & n14958;
  assign n14960 = ~n14750 & ~n14958;
  assign n14961 = ~n14959 & ~n14960;
  assign n14962 = pi111  & n2053;
  assign n14963 = pi112  & n1893;
  assign n14964 = pi113  & n1888;
  assign n14965 = n1886 & n7852;
  assign n14966 = ~n14963 & ~n14964;
  assign n14967 = ~n14962 & n14966;
  assign n14968 = ~n14965 & n14967;
  assign n14969 = pi23  & n14968;
  assign n14970 = ~pi23  & ~n14968;
  assign n14971 = ~n14969 & ~n14970;
  assign n14972 = ~n14621 & ~n14624;
  assign n14973 = ~n14971 & ~n14972;
  assign n14974 = n14971 & n14972;
  assign n14975 = ~n14973 & ~n14974;
  assign n14976 = n14961 & n14975;
  assign n14977 = ~n14961 & ~n14975;
  assign n14978 = ~n14976 & ~n14977;
  assign n14979 = n14736 & n14978;
  assign n14980 = ~n14736 & ~n14978;
  assign n14981 = ~n14979 & ~n14980;
  assign n14982 = n14722 & n14981;
  assign n14983 = ~n14722 & ~n14981;
  assign n14984 = ~n14982 & ~n14983;
  assign n14985 = n14708 & n14984;
  assign n14986 = ~n14708 & ~n14984;
  assign n14987 = ~n14985 & ~n14986;
  assign n14988 = n14694 & n14987;
  assign n14989 = ~n14694 & ~n14987;
  assign n14990 = ~n14988 & ~n14989;
  assign n14991 = n14679 & n14990;
  assign n14992 = ~n14679 & ~n14990;
  assign n14993 = ~n14991 & ~n14992;
  assign n14994 = ~n14666 & n14993;
  assign n14995 = n14666 & ~n14993;
  assign n14996 = ~n14994 & ~n14995;
  assign n14997 = ~n14665 & n14996;
  assign n14998 = n14665 & ~n14996;
  assign po70  = ~n14997 & ~n14998;
  assign n15000 = ~n14994 & ~n14997;
  assign n15001 = pi118  & n1296;
  assign n15002 = pi119  & n1207;
  assign n15003 = pi120  & n1202;
  assign n15004 = n1200 & n10047;
  assign n15005 = ~n15002 & ~n15003;
  assign n15006 = ~n15001 & n15005;
  assign n15007 = ~n15004 & n15006;
  assign n15008 = pi17  & n15007;
  assign n15009 = ~pi17  & ~n15007;
  assign n15010 = ~n15008 & ~n15009;
  assign n15011 = ~n14735 & ~n14979;
  assign n15012 = n15010 & n15011;
  assign n15013 = ~n15010 & ~n15011;
  assign n15014 = ~n15012 & ~n15013;
  assign n15015 = pi112  & n2053;
  assign n15016 = pi113  & n1893;
  assign n15017 = pi114  & n1888;
  assign n15018 = n1886 & n8146;
  assign n15019 = ~n15016 & ~n15017;
  assign n15020 = ~n15015 & n15019;
  assign n15021 = ~n15018 & n15020;
  assign n15022 = pi23  & n15021;
  assign n15023 = ~pi23  & ~n15021;
  assign n15024 = ~n15022 & ~n15023;
  assign n15025 = ~n14748 & ~n14959;
  assign n15026 = n15024 & n15025;
  assign n15027 = ~n15024 & ~n15025;
  assign n15028 = ~n15026 & ~n15027;
  assign n15029 = pi109  & n2510;
  assign n15030 = pi110  & n2342;
  assign n15031 = pi111  & n2337;
  assign n15032 = n2335 & n7272;
  assign n15033 = ~n15030 & ~n15031;
  assign n15034 = ~n15029 & n15033;
  assign n15035 = ~n15032 & n15034;
  assign n15036 = pi26  & n15035;
  assign n15037 = ~pi26  & ~n15035;
  assign n15038 = ~n15036 & ~n15037;
  assign n15039 = ~n14762 & ~n14956;
  assign n15040 = ~n15038 & ~n15039;
  assign n15041 = n15038 & n15039;
  assign n15042 = ~n15040 & ~n15041;
  assign n15043 = pi103  & n3553;
  assign n15044 = pi104  & n3334;
  assign n15045 = pi105  & n3329;
  assign n15046 = n3327 & n5677;
  assign n15047 = ~n15044 & ~n15045;
  assign n15048 = ~n15043 & n15047;
  assign n15049 = ~n15046 & n15048;
  assign n15050 = pi32  & n15049;
  assign n15051 = ~pi32  & ~n15049;
  assign n15052 = ~n15050 & ~n15051;
  assign n15053 = n14788 & ~n14947;
  assign n15054 = ~n14948 & ~n15053;
  assign n15055 = n15052 & ~n15054;
  assign n15056 = ~n15052 & n15054;
  assign n15057 = ~n15055 & ~n15056;
  assign n15058 = ~n14941 & ~n14944;
  assign n15059 = pi85  & n7969;
  assign n15060 = pi86  & n7636;
  assign n15061 = pi87  & n7631;
  assign n15062 = n2116 & n7629;
  assign n15063 = ~n15060 & ~n15061;
  assign n15064 = ~n15059 & n15063;
  assign n15065 = ~n15062 & n15064;
  assign n15066 = pi50  & n15065;
  assign n15067 = ~pi50  & ~n15065;
  assign n15068 = ~n15066 & ~n15067;
  assign n15069 = pi76  & n10886;
  assign n15070 = pi77  & n10495;
  assign n15071 = pi78  & n10490;
  assign n15072 = n958 & n10488;
  assign n15073 = ~n15070 & ~n15071;
  assign n15074 = ~n15069 & n15073;
  assign n15075 = ~n15072 & n15074;
  assign n15076 = pi59  & n15075;
  assign n15077 = ~pi59  & ~n15075;
  assign n15078 = ~n15076 & ~n15077;
  assign n15079 = pi73  & n11910;
  assign n15080 = pi74  & n11529;
  assign n15081 = pi75  & n11524;
  assign n15082 = n713 & n11522;
  assign n15083 = ~n15080 & ~n15081;
  assign n15084 = ~n15079 & n15083;
  assign n15085 = ~n15082 & n15084;
  assign n15086 = pi62  & n15085;
  assign n15087 = ~pi62  & ~n15085;
  assign n15088 = ~n15086 & ~n15087;
  assign n15089 = ~n14811 & ~n14824;
  assign n15090 = pi72  & n12277;
  assign n15091 = pi71  & n12276;
  assign n15092 = ~n15090 & ~n15091;
  assign n15093 = n14810 & ~n15092;
  assign n15094 = ~n14810 & n15092;
  assign n15095 = ~n15093 & ~n15094;
  assign n15096 = ~n15089 & n15095;
  assign n15097 = n15089 & ~n15095;
  assign n15098 = ~n15096 & ~n15097;
  assign n15099 = ~n15088 & n15098;
  assign n15100 = n15088 & ~n15098;
  assign n15101 = ~n15099 & ~n15100;
  assign n15102 = ~n15078 & n15101;
  assign n15103 = n15078 & ~n15101;
  assign n15104 = ~n15102 & ~n15103;
  assign n15105 = ~n14827 & n14839;
  assign n15106 = ~n14828 & ~n15105;
  assign n15107 = ~n15104 & ~n15106;
  assign n15108 = n15104 & n15106;
  assign n15109 = ~n15107 & ~n15108;
  assign n15110 = pi79  & n9858;
  assign n15111 = pi80  & n9508;
  assign n15112 = pi81  & n9503;
  assign n15113 = n1337 & n9501;
  assign n15114 = ~n15111 & ~n15112;
  assign n15115 = ~n15110 & n15114;
  assign n15116 = ~n15113 & n15115;
  assign n15117 = pi56  & n15116;
  assign n15118 = ~pi56  & ~n15116;
  assign n15119 = ~n15117 & ~n15118;
  assign n15120 = n15109 & ~n15119;
  assign n15121 = ~n15109 & n15119;
  assign n15122 = ~n15120 & ~n15121;
  assign n15123 = ~n14844 & n14855;
  assign n15124 = ~n14843 & ~n15123;
  assign n15125 = ~n15122 & ~n15124;
  assign n15126 = n15122 & n15124;
  assign n15127 = ~n15125 & ~n15126;
  assign n15128 = pi82  & n8905;
  assign n15129 = pi83  & n8535;
  assign n15130 = pi84  & n8530;
  assign n15131 = n1601 & n8528;
  assign n15132 = ~n15129 & ~n15130;
  assign n15133 = ~n15128 & n15132;
  assign n15134 = ~n15131 & n15133;
  assign n15135 = pi53  & n15134;
  assign n15136 = ~pi53  & ~n15134;
  assign n15137 = ~n15135 & ~n15136;
  assign n15138 = ~n15127 & n15137;
  assign n15139 = n15127 & ~n15137;
  assign n15140 = ~n15138 & ~n15139;
  assign n15141 = ~n14860 & n14871;
  assign n15142 = ~n14859 & ~n15141;
  assign n15143 = n15140 & n15142;
  assign n15144 = ~n15140 & ~n15142;
  assign n15145 = ~n15143 & ~n15144;
  assign n15146 = ~n15068 & n15145;
  assign n15147 = n15068 & ~n15145;
  assign n15148 = ~n15146 & ~n15147;
  assign n15149 = ~n14876 & n14887;
  assign n15150 = ~n14875 & ~n15149;
  assign n15151 = n15148 & n15150;
  assign n15152 = ~n15148 & ~n15150;
  assign n15153 = ~n15151 & ~n15152;
  assign n15154 = pi88  & n7121;
  assign n15155 = pi89  & n6795;
  assign n15156 = pi90  & n6790;
  assign n15157 = n2448 & n6788;
  assign n15158 = ~n15155 & ~n15156;
  assign n15159 = ~n15154 & n15158;
  assign n15160 = ~n15157 & n15159;
  assign n15161 = pi47  & n15160;
  assign n15162 = ~pi47  & ~n15160;
  assign n15163 = ~n15161 & ~n15162;
  assign n15164 = n15153 & ~n15163;
  assign n15165 = ~n15153 & n15163;
  assign n15166 = ~n15164 & ~n15165;
  assign n15167 = ~n14892 & n14903;
  assign n15168 = ~n14891 & ~n15167;
  assign n15169 = ~n15166 & ~n15168;
  assign n15170 = n15166 & n15168;
  assign n15171 = ~n15169 & ~n15170;
  assign n15172 = pi91  & n6331;
  assign n15173 = pi92  & n6015;
  assign n15174 = pi93  & n6010;
  assign n15175 = n2948 & n6008;
  assign n15176 = ~n15173 & ~n15174;
  assign n15177 = ~n15172 & n15176;
  assign n15178 = ~n15175 & n15177;
  assign n15179 = pi44  & n15178;
  assign n15180 = ~pi44  & ~n15178;
  assign n15181 = ~n15179 & ~n15180;
  assign n15182 = n15171 & ~n15181;
  assign n15183 = ~n15171 & n15181;
  assign n15184 = ~n15182 & ~n15183;
  assign n15185 = ~n14908 & n14919;
  assign n15186 = ~n14907 & ~n15185;
  assign n15187 = ~n15184 & ~n15186;
  assign n15188 = n15184 & n15186;
  assign n15189 = ~n15187 & ~n15188;
  assign n15190 = pi94  & n5558;
  assign n15191 = pi95  & n5293;
  assign n15192 = pi96  & n5288;
  assign n15193 = n3499 & n5286;
  assign n15194 = ~n15191 & ~n15192;
  assign n15195 = ~n15190 & n15194;
  assign n15196 = ~n15193 & n15195;
  assign n15197 = pi41  & n15196;
  assign n15198 = ~pi41  & ~n15196;
  assign n15199 = ~n15197 & ~n15198;
  assign n15200 = ~n15189 & n15199;
  assign n15201 = n15189 & ~n15199;
  assign n15202 = ~n15200 & ~n15201;
  assign n15203 = ~n14924 & ~n14937;
  assign n15204 = n15202 & ~n15203;
  assign n15205 = ~n15202 & n15203;
  assign n15206 = ~n15204 & ~n15205;
  assign n15207 = pi97  & n4843;
  assign n15208 = pi98  & n4598;
  assign n15209 = pi99  & n4593;
  assign n15210 = n4101 & n4591;
  assign n15211 = ~n15208 & ~n15209;
  assign n15212 = ~n15207 & n15211;
  assign n15213 = ~n15210 & n15212;
  assign n15214 = pi38  & n15213;
  assign n15215 = ~pi38  & ~n15213;
  assign n15216 = ~n15214 & ~n15215;
  assign n15217 = n15206 & ~n15216;
  assign n15218 = ~n15206 & n15216;
  assign n15219 = ~n15217 & ~n15218;
  assign n15220 = n15058 & ~n15219;
  assign n15221 = ~n15058 & n15219;
  assign n15222 = ~n15220 & ~n15221;
  assign n15223 = pi100  & n4176;
  assign n15224 = pi101  & n3938;
  assign n15225 = pi102  & n3933;
  assign n15226 = n3931 & n4956;
  assign n15227 = ~n15224 & ~n15225;
  assign n15228 = ~n15223 & n15227;
  assign n15229 = ~n15226 & n15228;
  assign n15230 = pi35  & n15229;
  assign n15231 = ~pi35  & ~n15229;
  assign n15232 = ~n15230 & ~n15231;
  assign n15233 = n15222 & ~n15232;
  assign n15234 = ~n15222 & n15232;
  assign n15235 = ~n15233 & ~n15234;
  assign n15236 = n15057 & n15235;
  assign n15237 = ~n15057 & ~n15235;
  assign n15238 = ~n15236 & ~n15237;
  assign n15239 = pi106  & n3011;
  assign n15240 = pi107  & n2809;
  assign n15241 = pi108  & n2804;
  assign n15242 = n2802 & n6213;
  assign n15243 = ~n15240 & ~n15241;
  assign n15244 = ~n15239 & n15243;
  assign n15245 = ~n15242 & n15244;
  assign n15246 = pi29  & n15245;
  assign n15247 = ~pi29  & ~n15245;
  assign n15248 = ~n15246 & ~n15247;
  assign n15249 = ~n14777 & ~n14952;
  assign n15250 = ~n14776 & ~n15249;
  assign n15251 = ~n15248 & n15250;
  assign n15252 = n15248 & ~n15250;
  assign n15253 = ~n15251 & ~n15252;
  assign n15254 = n15238 & n15253;
  assign n15255 = ~n15238 & ~n15253;
  assign n15256 = ~n15254 & ~n15255;
  assign n15257 = n15042 & n15256;
  assign n15258 = ~n15042 & ~n15256;
  assign n15259 = ~n15257 & ~n15258;
  assign n15260 = ~n15028 & ~n15259;
  assign n15261 = n15028 & n15259;
  assign n15262 = ~n15260 & ~n15261;
  assign n15263 = ~n14973 & ~n14976;
  assign n15264 = pi115  & n1661;
  assign n15265 = pi116  & n1500;
  assign n15266 = pi117  & n1495;
  assign n15267 = n1493 & n8784;
  assign n15268 = ~n15265 & ~n15266;
  assign n15269 = ~n15264 & n15268;
  assign n15270 = ~n15267 & n15269;
  assign n15271 = pi20  & n15270;
  assign n15272 = ~pi20  & ~n15270;
  assign n15273 = ~n15271 & ~n15272;
  assign n15274 = ~n15263 & ~n15273;
  assign n15275 = n15263 & n15273;
  assign n15276 = ~n15274 & ~n15275;
  assign n15277 = n15262 & n15276;
  assign n15278 = ~n15262 & ~n15276;
  assign n15279 = ~n15277 & ~n15278;
  assign n15280 = n15014 & ~n15279;
  assign n15281 = ~n15014 & n15279;
  assign n15282 = ~n15280 & ~n15281;
  assign n15283 = pi121  & n1006;
  assign n15284 = pi122  & n897;
  assign n15285 = pi123  & n892;
  assign n15286 = n890 & n10754;
  assign n15287 = ~n15284 & ~n15285;
  assign n15288 = ~n15283 & n15287;
  assign n15289 = ~n15286 & n15288;
  assign n15290 = pi14  & n15289;
  assign n15291 = ~pi14  & ~n15289;
  assign n15292 = ~n15290 & ~n15291;
  assign n15293 = ~n14721 & ~n14982;
  assign n15294 = ~n15292 & ~n15293;
  assign n15295 = n15292 & n15293;
  assign n15296 = ~n15294 & ~n15295;
  assign n15297 = ~n15282 & n15296;
  assign n15298 = n15282 & ~n15296;
  assign n15299 = ~n15297 & ~n15298;
  assign n15300 = ~n14706 & ~n14985;
  assign n15301 = pi124  & n750;
  assign n15302 = pi125  & n651;
  assign n15303 = pi126  & n646;
  assign n15304 = n644 & n12148;
  assign n15305 = ~n15302 & ~n15303;
  assign n15306 = ~n15301 & n15305;
  assign n15307 = ~n15304 & n15306;
  assign n15308 = pi11  & n15307;
  assign n15309 = ~pi11  & ~n15307;
  assign n15310 = ~n15308 & ~n15309;
  assign n15311 = ~n15300 & ~n15310;
  assign n15312 = n15300 & n15310;
  assign n15313 = ~n15311 & ~n15312;
  assign n15314 = n15299 & n15313;
  assign n15315 = ~n15299 & ~n15313;
  assign n15316 = ~n15314 & ~n15315;
  assign n15317 = ~n14693 & ~n14988;
  assign n15318 = n483 & ~n12539;
  assign n15319 = ~n528 & ~n15318;
  assign n15320 = pi127  & ~n15319;
  assign n15321 = pi8  & ~n15320;
  assign n15322 = ~pi8  & n15320;
  assign n15323 = ~n15321 & ~n15322;
  assign n15324 = ~n15317 & ~n15323;
  assign n15325 = n15317 & n15323;
  assign n15326 = ~n15324 & ~n15325;
  assign n15327 = n15316 & n15326;
  assign n15328 = ~n15316 & ~n15326;
  assign n15329 = ~n15327 & ~n15328;
  assign n15330 = ~n14677 & ~n14990;
  assign n15331 = ~n14678 & ~n15330;
  assign n15332 = n15329 & n15331;
  assign n15333 = ~n15329 & ~n15331;
  assign n15334 = ~n15332 & ~n15333;
  assign n15335 = ~n15000 & n15334;
  assign n15336 = n15000 & ~n15334;
  assign po71  = ~n15335 & ~n15336;
  assign n15338 = ~n15332 & ~n15335;
  assign n15339 = ~n15324 & ~n15327;
  assign n15340 = pi119  & n1296;
  assign n15341 = pi120  & n1207;
  assign n15342 = pi121  & n1202;
  assign n15343 = n1200 & n10071;
  assign n15344 = ~n15341 & ~n15342;
  assign n15345 = ~n15340 & n15344;
  assign n15346 = ~n15343 & n15345;
  assign n15347 = pi17  & n15346;
  assign n15348 = ~pi17  & ~n15346;
  assign n15349 = ~n15347 & ~n15348;
  assign n15350 = ~n15013 & ~n15279;
  assign n15351 = ~n15012 & ~n15350;
  assign n15352 = n15349 & ~n15351;
  assign n15353 = ~n15349 & n15351;
  assign n15354 = ~n15352 & ~n15353;
  assign n15355 = pi113  & n2053;
  assign n15356 = pi114  & n1893;
  assign n15357 = pi115  & n1888;
  assign n15358 = n1886 & n8170;
  assign n15359 = ~n15356 & ~n15357;
  assign n15360 = ~n15355 & n15359;
  assign n15361 = ~n15358 & n15360;
  assign n15362 = pi23  & n15361;
  assign n15363 = ~pi23  & ~n15361;
  assign n15364 = ~n15362 & ~n15363;
  assign n15365 = ~n15027 & ~n15261;
  assign n15366 = ~n15364 & ~n15365;
  assign n15367 = n15364 & n15365;
  assign n15368 = ~n15366 & ~n15367;
  assign n15369 = pi110  & n2510;
  assign n15370 = pi111  & n2342;
  assign n15371 = pi112  & n2337;
  assign n15372 = n2335 & n7296;
  assign n15373 = ~n15370 & ~n15371;
  assign n15374 = ~n15369 & n15373;
  assign n15375 = ~n15372 & n15374;
  assign n15376 = pi26  & n15375;
  assign n15377 = ~pi26  & ~n15375;
  assign n15378 = ~n15376 & ~n15377;
  assign n15379 = ~n15040 & ~n15257;
  assign n15380 = n15378 & n15379;
  assign n15381 = ~n15378 & ~n15379;
  assign n15382 = ~n15380 & ~n15381;
  assign n15383 = ~n15251 & ~n15254;
  assign n15384 = pi107  & n3011;
  assign n15385 = pi108  & n2809;
  assign n15386 = pi109  & n2804;
  assign n15387 = n2802 & n6715;
  assign n15388 = ~n15385 & ~n15386;
  assign n15389 = ~n15384 & n15388;
  assign n15390 = ~n15387 & n15389;
  assign n15391 = pi29  & n15390;
  assign n15392 = ~pi29  & ~n15390;
  assign n15393 = ~n15391 & ~n15392;
  assign n15394 = ~n15383 & ~n15393;
  assign n15395 = n15383 & n15393;
  assign n15396 = ~n15394 & ~n15395;
  assign n15397 = ~n15221 & ~n15233;
  assign n15398 = pi98  & n4843;
  assign n15399 = pi99  & n4598;
  assign n15400 = pi100  & n4593;
  assign n15401 = n4501 & n4591;
  assign n15402 = ~n15399 & ~n15400;
  assign n15403 = ~n15398 & n15402;
  assign n15404 = ~n15401 & n15403;
  assign n15405 = pi38  & n15404;
  assign n15406 = ~pi38  & ~n15404;
  assign n15407 = ~n15405 & ~n15406;
  assign n15408 = ~n15188 & ~n15201;
  assign n15409 = pi95  & n5558;
  assign n15410 = pi96  & n5293;
  assign n15411 = pi97  & n5288;
  assign n15412 = n3691 & n5286;
  assign n15413 = ~n15410 & ~n15411;
  assign n15414 = ~n15409 & n15413;
  assign n15415 = ~n15412 & n15414;
  assign n15416 = pi41  & n15415;
  assign n15417 = ~pi41  & ~n15415;
  assign n15418 = ~n15416 & ~n15417;
  assign n15419 = pi89  & n7121;
  assign n15420 = pi90  & n6795;
  assign n15421 = pi91  & n6790;
  assign n15422 = n2746 & n6788;
  assign n15423 = ~n15420 & ~n15421;
  assign n15424 = ~n15419 & n15423;
  assign n15425 = ~n15422 & n15424;
  assign n15426 = pi47  & n15425;
  assign n15427 = ~pi47  & ~n15425;
  assign n15428 = ~n15426 & ~n15427;
  assign n15429 = ~n15143 & ~n15146;
  assign n15430 = pi86  & n7969;
  assign n15431 = pi87  & n7636;
  assign n15432 = pi88  & n7631;
  assign n15433 = n2140 & n7629;
  assign n15434 = ~n15431 & ~n15432;
  assign n15435 = ~n15430 & n15434;
  assign n15436 = ~n15433 & n15435;
  assign n15437 = pi50  & n15436;
  assign n15438 = ~pi50  & ~n15436;
  assign n15439 = ~n15437 & ~n15438;
  assign n15440 = ~n15126 & ~n15139;
  assign n15441 = ~n15099 & ~n15102;
  assign n15442 = pi77  & n10886;
  assign n15443 = pi78  & n10495;
  assign n15444 = pi79  & n10490;
  assign n15445 = n1048 & n10488;
  assign n15446 = ~n15443 & ~n15444;
  assign n15447 = ~n15442 & n15446;
  assign n15448 = ~n15445 & n15447;
  assign n15449 = pi59  & n15448;
  assign n15450 = ~pi59  & ~n15448;
  assign n15451 = ~n15449 & ~n15450;
  assign n15452 = pi74  & n11910;
  assign n15453 = pi75  & n11529;
  assign n15454 = pi76  & n11524;
  assign n15455 = n841 & n11522;
  assign n15456 = ~n15453 & ~n15454;
  assign n15457 = ~n15452 & n15456;
  assign n15458 = ~n15455 & n15457;
  assign n15459 = pi62  & n15458;
  assign n15460 = ~pi62  & ~n15458;
  assign n15461 = ~n15459 & ~n15460;
  assign n15462 = ~n15094 & ~n15096;
  assign n15463 = ~pi8  & ~n15092;
  assign n15464 = pi8  & n15092;
  assign n15465 = ~n15463 & ~n15464;
  assign n15466 = pi73  & n12277;
  assign n15467 = pi72  & n12276;
  assign n15468 = ~n15466 & ~n15467;
  assign n15469 = n15465 & ~n15468;
  assign n15470 = ~n15465 & n15468;
  assign n15471 = ~n15469 & ~n15470;
  assign n15472 = ~n15462 & n15471;
  assign n15473 = n15462 & ~n15471;
  assign n15474 = ~n15472 & ~n15473;
  assign n15475 = ~n15461 & n15474;
  assign n15476 = n15461 & ~n15474;
  assign n15477 = ~n15475 & ~n15476;
  assign n15478 = ~n15451 & n15477;
  assign n15479 = n15451 & ~n15477;
  assign n15480 = ~n15478 & ~n15479;
  assign n15481 = ~n15441 & n15480;
  assign n15482 = n15441 & ~n15480;
  assign n15483 = ~n15481 & ~n15482;
  assign n15484 = pi80  & n9858;
  assign n15485 = pi81  & n9508;
  assign n15486 = pi82  & n9503;
  assign n15487 = n1450 & n9501;
  assign n15488 = ~n15485 & ~n15486;
  assign n15489 = ~n15484 & n15488;
  assign n15490 = ~n15487 & n15489;
  assign n15491 = pi56  & n15490;
  assign n15492 = ~pi56  & ~n15490;
  assign n15493 = ~n15491 & ~n15492;
  assign n15494 = n15483 & ~n15493;
  assign n15495 = ~n15483 & n15493;
  assign n15496 = ~n15494 & ~n15495;
  assign n15497 = ~n15108 & n15119;
  assign n15498 = ~n15107 & ~n15497;
  assign n15499 = ~n15496 & ~n15498;
  assign n15500 = n15496 & n15498;
  assign n15501 = ~n15499 & ~n15500;
  assign n15502 = pi83  & n8905;
  assign n15503 = pi84  & n8535;
  assign n15504 = pi85  & n8530;
  assign n15505 = n1831 & n8528;
  assign n15506 = ~n15503 & ~n15504;
  assign n15507 = ~n15502 & n15506;
  assign n15508 = ~n15505 & n15507;
  assign n15509 = pi53  & n15508;
  assign n15510 = ~pi53  & ~n15508;
  assign n15511 = ~n15509 & ~n15510;
  assign n15512 = n15501 & ~n15511;
  assign n15513 = ~n15501 & n15511;
  assign n15514 = ~n15512 & ~n15513;
  assign n15515 = ~n15440 & n15514;
  assign n15516 = n15440 & ~n15514;
  assign n15517 = ~n15515 & ~n15516;
  assign n15518 = ~n15439 & n15517;
  assign n15519 = n15439 & ~n15517;
  assign n15520 = ~n15518 & ~n15519;
  assign n15521 = ~n15429 & n15520;
  assign n15522 = n15429 & ~n15520;
  assign n15523 = ~n15521 & ~n15522;
  assign n15524 = ~n15428 & n15523;
  assign n15525 = n15428 & ~n15523;
  assign n15526 = ~n15524 & ~n15525;
  assign n15527 = ~n15151 & n15163;
  assign n15528 = ~n15152 & ~n15527;
  assign n15529 = ~n15526 & ~n15528;
  assign n15530 = n15526 & n15528;
  assign n15531 = ~n15529 & ~n15530;
  assign n15532 = pi92  & n6331;
  assign n15533 = pi93  & n6015;
  assign n15534 = pi94  & n6010;
  assign n15535 = n3280 & n6008;
  assign n15536 = ~n15533 & ~n15534;
  assign n15537 = ~n15532 & n15536;
  assign n15538 = ~n15535 & n15537;
  assign n15539 = pi44  & n15538;
  assign n15540 = ~pi44  & ~n15538;
  assign n15541 = ~n15539 & ~n15540;
  assign n15542 = n15531 & ~n15541;
  assign n15543 = ~n15531 & n15541;
  assign n15544 = ~n15542 & ~n15543;
  assign n15545 = ~n15170 & n15181;
  assign n15546 = ~n15169 & ~n15545;
  assign n15547 = n15544 & ~n15546;
  assign n15548 = ~n15544 & n15546;
  assign n15549 = ~n15547 & ~n15548;
  assign n15550 = ~n15418 & ~n15549;
  assign n15551 = n15418 & n15549;
  assign n15552 = ~n15550 & ~n15551;
  assign n15553 = ~n15408 & n15552;
  assign n15554 = n15408 & ~n15552;
  assign n15555 = ~n15553 & ~n15554;
  assign n15556 = ~n15407 & n15555;
  assign n15557 = n15407 & ~n15555;
  assign n15558 = ~n15556 & ~n15557;
  assign n15559 = ~n15205 & ~n15216;
  assign n15560 = ~n15204 & ~n15559;
  assign n15561 = ~n15558 & n15560;
  assign n15562 = n15558 & ~n15560;
  assign n15563 = ~n15561 & ~n15562;
  assign n15564 = pi101  & n4176;
  assign n15565 = pi102  & n3938;
  assign n15566 = pi103  & n3933;
  assign n15567 = n3931 & n5188;
  assign n15568 = ~n15565 & ~n15566;
  assign n15569 = ~n15564 & n15568;
  assign n15570 = ~n15567 & n15569;
  assign n15571 = pi35  & n15570;
  assign n15572 = ~pi35  & ~n15570;
  assign n15573 = ~n15571 & ~n15572;
  assign n15574 = n15563 & ~n15573;
  assign n15575 = ~n15563 & n15573;
  assign n15576 = ~n15574 & ~n15575;
  assign n15577 = ~n15397 & n15576;
  assign n15578 = n15397 & ~n15576;
  assign n15579 = ~n15577 & ~n15578;
  assign n15580 = ~n15056 & ~n15236;
  assign n15581 = pi104  & n3553;
  assign n15582 = pi105  & n3334;
  assign n15583 = pi106  & n3329;
  assign n15584 = n3327 & n5701;
  assign n15585 = ~n15582 & ~n15583;
  assign n15586 = ~n15581 & n15585;
  assign n15587 = ~n15584 & n15586;
  assign n15588 = pi32  & n15587;
  assign n15589 = ~pi32  & ~n15587;
  assign n15590 = ~n15588 & ~n15589;
  assign n15591 = ~n15580 & ~n15590;
  assign n15592 = n15580 & n15590;
  assign n15593 = ~n15591 & ~n15592;
  assign n15594 = n15579 & n15593;
  assign n15595 = ~n15579 & ~n15593;
  assign n15596 = ~n15594 & ~n15595;
  assign n15597 = n15396 & n15596;
  assign n15598 = ~n15396 & ~n15596;
  assign n15599 = ~n15597 & ~n15598;
  assign n15600 = n15382 & n15599;
  assign n15601 = ~n15382 & ~n15599;
  assign n15602 = ~n15600 & ~n15601;
  assign n15603 = ~n15368 & n15602;
  assign n15604 = n15368 & ~n15602;
  assign n15605 = ~n15603 & ~n15604;
  assign n15606 = ~n15274 & ~n15277;
  assign n15607 = pi116  & n1661;
  assign n15608 = pi117  & n1500;
  assign n15609 = pi118  & n1495;
  assign n15610 = n1493 & n9095;
  assign n15611 = ~n15608 & ~n15609;
  assign n15612 = ~n15607 & n15611;
  assign n15613 = ~n15610 & n15612;
  assign n15614 = pi20  & n15613;
  assign n15615 = ~pi20  & ~n15613;
  assign n15616 = ~n15614 & ~n15615;
  assign n15617 = ~n15606 & ~n15616;
  assign n15618 = n15606 & n15616;
  assign n15619 = ~n15617 & ~n15618;
  assign n15620 = ~n15605 & n15619;
  assign n15621 = n15605 & ~n15619;
  assign n15622 = ~n15620 & ~n15621;
  assign n15623 = n15354 & n15622;
  assign n15624 = ~n15354 & ~n15622;
  assign n15625 = ~n15623 & ~n15624;
  assign n15626 = ~n15294 & ~n15297;
  assign n15627 = pi122  & n1006;
  assign n15628 = pi123  & n897;
  assign n15629 = pi124  & n892;
  assign n15630 = n890 & n11099;
  assign n15631 = ~n15628 & ~n15629;
  assign n15632 = ~n15627 & n15631;
  assign n15633 = ~n15630 & n15632;
  assign n15634 = pi14  & n15633;
  assign n15635 = ~pi14  & ~n15633;
  assign n15636 = ~n15634 & ~n15635;
  assign n15637 = ~n15626 & ~n15636;
  assign n15638 = n15626 & n15636;
  assign n15639 = ~n15637 & ~n15638;
  assign n15640 = n15625 & n15639;
  assign n15641 = ~n15625 & ~n15639;
  assign n15642 = ~n15640 & ~n15641;
  assign n15643 = ~n15311 & ~n15314;
  assign n15644 = pi125  & n750;
  assign n15645 = pi126  & n651;
  assign n15646 = pi127  & n646;
  assign n15647 = n644 & n12519;
  assign n15648 = ~n15645 & ~n15646;
  assign n15649 = ~n15644 & n15648;
  assign n15650 = ~n15647 & n15649;
  assign n15651 = pi11  & n15650;
  assign n15652 = ~pi11  & ~n15650;
  assign n15653 = ~n15651 & ~n15652;
  assign n15654 = ~n15643 & ~n15653;
  assign n15655 = n15643 & n15653;
  assign n15656 = ~n15654 & ~n15655;
  assign n15657 = n15642 & n15656;
  assign n15658 = ~n15642 & ~n15656;
  assign n15659 = ~n15657 & ~n15658;
  assign n15660 = ~n15339 & n15659;
  assign n15661 = n15339 & ~n15659;
  assign n15662 = ~n15660 & ~n15661;
  assign n15663 = ~n15338 & n15662;
  assign n15664 = n15338 & ~n15662;
  assign po72  = ~n15663 & ~n15664;
  assign n15666 = ~n15660 & ~n15663;
  assign n15667 = ~n15654 & ~n15657;
  assign n15668 = pi123  & n1006;
  assign n15669 = pi124  & n897;
  assign n15670 = pi125  & n892;
  assign n15671 = n890 & n11786;
  assign n15672 = ~n15669 & ~n15670;
  assign n15673 = ~n15668 & n15672;
  assign n15674 = ~n15671 & n15673;
  assign n15675 = pi14  & n15674;
  assign n15676 = ~pi14  & ~n15674;
  assign n15677 = ~n15675 & ~n15676;
  assign n15678 = ~n15353 & ~n15623;
  assign n15679 = ~n15677 & ~n15678;
  assign n15680 = n15677 & n15678;
  assign n15681 = ~n15679 & ~n15680;
  assign n15682 = pi117  & n1661;
  assign n15683 = pi118  & n1500;
  assign n15684 = pi119  & n1495;
  assign n15685 = n1493 & n9412;
  assign n15686 = ~n15683 & ~n15684;
  assign n15687 = ~n15682 & n15686;
  assign n15688 = ~n15685 & n15687;
  assign n15689 = pi20  & n15688;
  assign n15690 = ~pi20  & ~n15688;
  assign n15691 = ~n15689 & ~n15690;
  assign n15692 = ~n15366 & ~n15602;
  assign n15693 = ~n15367 & ~n15692;
  assign n15694 = n15691 & ~n15693;
  assign n15695 = ~n15691 & n15693;
  assign n15696 = ~n15694 & ~n15695;
  assign n15697 = pi114  & n2053;
  assign n15698 = pi115  & n1893;
  assign n15699 = pi116  & n1888;
  assign n15700 = n1886 & n8470;
  assign n15701 = ~n15698 & ~n15699;
  assign n15702 = ~n15697 & n15701;
  assign n15703 = ~n15700 & n15702;
  assign n15704 = pi23  & n15703;
  assign n15705 = ~pi23  & ~n15703;
  assign n15706 = ~n15704 & ~n15705;
  assign n15707 = ~n15381 & ~n15600;
  assign n15708 = n15706 & n15707;
  assign n15709 = ~n15706 & ~n15707;
  assign n15710 = ~n15708 & ~n15709;
  assign n15711 = ~n15591 & ~n15594;
  assign n15712 = pi108  & n3011;
  assign n15713 = pi109  & n2809;
  assign n15714 = pi110  & n2804;
  assign n15715 = n2802 & n6995;
  assign n15716 = ~n15713 & ~n15714;
  assign n15717 = ~n15712 & n15716;
  assign n15718 = ~n15715 & n15717;
  assign n15719 = pi29  & n15718;
  assign n15720 = ~pi29  & ~n15718;
  assign n15721 = ~n15719 & ~n15720;
  assign n15722 = ~n15711 & ~n15721;
  assign n15723 = n15711 & n15721;
  assign n15724 = ~n15722 & ~n15723;
  assign n15725 = pi105  & n3553;
  assign n15726 = pi106  & n3334;
  assign n15727 = pi107  & n3329;
  assign n15728 = n3327 & n6189;
  assign n15729 = ~n15726 & ~n15727;
  assign n15730 = ~n15725 & n15729;
  assign n15731 = ~n15728 & n15730;
  assign n15732 = pi32  & n15731;
  assign n15733 = ~pi32  & ~n15731;
  assign n15734 = ~n15732 & ~n15733;
  assign n15735 = ~n15574 & ~n15577;
  assign n15736 = n15734 & n15735;
  assign n15737 = ~n15734 & ~n15735;
  assign n15738 = ~n15736 & ~n15737;
  assign n15739 = pi102  & n4176;
  assign n15740 = pi103  & n3938;
  assign n15741 = pi104  & n3933;
  assign n15742 = n3931 & n5212;
  assign n15743 = ~n15740 & ~n15741;
  assign n15744 = ~n15739 & n15743;
  assign n15745 = ~n15742 & n15744;
  assign n15746 = pi35  & n15745;
  assign n15747 = ~pi35  & ~n15745;
  assign n15748 = ~n15746 & ~n15747;
  assign n15749 = ~n15556 & ~n15562;
  assign n15750 = pi99  & n4843;
  assign n15751 = pi100  & n4598;
  assign n15752 = pi101  & n4593;
  assign n15753 = n4591 & n4730;
  assign n15754 = ~n15751 & ~n15752;
  assign n15755 = ~n15750 & n15754;
  assign n15756 = ~n15753 & n15755;
  assign n15757 = pi38  & n15756;
  assign n15758 = ~pi38  & ~n15756;
  assign n15759 = ~n15757 & ~n15758;
  assign n15760 = ~n15550 & ~n15553;
  assign n15761 = pi96  & n5558;
  assign n15762 = pi97  & n5293;
  assign n15763 = pi98  & n5288;
  assign n15764 = n3889 & n5286;
  assign n15765 = ~n15762 & ~n15763;
  assign n15766 = ~n15761 & n15765;
  assign n15767 = ~n15764 & n15766;
  assign n15768 = pi41  & n15767;
  assign n15769 = ~pi41  & ~n15767;
  assign n15770 = ~n15768 & ~n15769;
  assign n15771 = ~n15524 & ~n15530;
  assign n15772 = ~n15518 & ~n15521;
  assign n15773 = ~n15512 & ~n15515;
  assign n15774 = ~n15494 & ~n15500;
  assign n15775 = ~n15478 & ~n15481;
  assign n15776 = pi78  & n10886;
  assign n15777 = pi79  & n10495;
  assign n15778 = pi80  & n10490;
  assign n15779 = n1144 & n10488;
  assign n15780 = ~n15777 & ~n15778;
  assign n15781 = ~n15776 & n15780;
  assign n15782 = ~n15779 & n15781;
  assign n15783 = pi59  & n15782;
  assign n15784 = ~pi59  & ~n15782;
  assign n15785 = ~n15783 & ~n15784;
  assign n15786 = ~n15472 & ~n15475;
  assign n15787 = pi75  & n11910;
  assign n15788 = pi76  & n11529;
  assign n15789 = pi77  & n11524;
  assign n15790 = n865 & n11522;
  assign n15791 = ~n15788 & ~n15789;
  assign n15792 = ~n15787 & n15791;
  assign n15793 = ~n15790 & n15792;
  assign n15794 = pi62  & n15793;
  assign n15795 = ~pi62  & ~n15793;
  assign n15796 = ~n15794 & ~n15795;
  assign n15797 = ~n15463 & ~n15469;
  assign n15798 = pi74  & n12277;
  assign n15799 = pi73  & n12276;
  assign n15800 = ~n15798 & ~n15799;
  assign n15801 = ~n15797 & n15800;
  assign n15802 = n15797 & ~n15800;
  assign n15803 = ~n15801 & ~n15802;
  assign n15804 = n15796 & ~n15803;
  assign n15805 = ~n15796 & n15803;
  assign n15806 = ~n15804 & ~n15805;
  assign n15807 = ~n15786 & n15806;
  assign n15808 = n15786 & ~n15806;
  assign n15809 = ~n15807 & ~n15808;
  assign n15810 = n15785 & ~n15809;
  assign n15811 = ~n15785 & n15809;
  assign n15812 = ~n15810 & ~n15811;
  assign n15813 = n15775 & ~n15812;
  assign n15814 = ~n15775 & n15812;
  assign n15815 = ~n15813 & ~n15814;
  assign n15816 = pi81  & n9858;
  assign n15817 = pi82  & n9508;
  assign n15818 = pi83  & n9503;
  assign n15819 = n1577 & n9501;
  assign n15820 = ~n15817 & ~n15818;
  assign n15821 = ~n15816 & n15820;
  assign n15822 = ~n15819 & n15821;
  assign n15823 = pi56  & n15822;
  assign n15824 = ~pi56  & ~n15822;
  assign n15825 = ~n15823 & ~n15824;
  assign n15826 = n15815 & ~n15825;
  assign n15827 = ~n15815 & n15825;
  assign n15828 = ~n15826 & ~n15827;
  assign n15829 = n15774 & ~n15828;
  assign n15830 = ~n15774 & n15828;
  assign n15831 = ~n15829 & ~n15830;
  assign n15832 = pi84  & n8905;
  assign n15833 = pi85  & n8535;
  assign n15834 = pi86  & n8530;
  assign n15835 = n1975 & n8528;
  assign n15836 = ~n15833 & ~n15834;
  assign n15837 = ~n15832 & n15836;
  assign n15838 = ~n15835 & n15837;
  assign n15839 = pi53  & n15838;
  assign n15840 = ~pi53  & ~n15838;
  assign n15841 = ~n15839 & ~n15840;
  assign n15842 = n15831 & ~n15841;
  assign n15843 = ~n15831 & n15841;
  assign n15844 = ~n15842 & ~n15843;
  assign n15845 = n15773 & ~n15844;
  assign n15846 = ~n15773 & n15844;
  assign n15847 = ~n15845 & ~n15846;
  assign n15848 = pi87  & n7969;
  assign n15849 = pi88  & n7636;
  assign n15850 = pi89  & n7631;
  assign n15851 = n2287 & n7629;
  assign n15852 = ~n15849 & ~n15850;
  assign n15853 = ~n15848 & n15852;
  assign n15854 = ~n15851 & n15853;
  assign n15855 = pi50  & n15854;
  assign n15856 = ~pi50  & ~n15854;
  assign n15857 = ~n15855 & ~n15856;
  assign n15858 = n15847 & ~n15857;
  assign n15859 = ~n15847 & n15857;
  assign n15860 = ~n15858 & ~n15859;
  assign n15861 = n15772 & ~n15860;
  assign n15862 = ~n15772 & n15860;
  assign n15863 = ~n15861 & ~n15862;
  assign n15864 = pi90  & n7121;
  assign n15865 = pi91  & n6795;
  assign n15866 = pi92  & n6790;
  assign n15867 = n2924 & n6788;
  assign n15868 = ~n15865 & ~n15866;
  assign n15869 = ~n15864 & n15868;
  assign n15870 = ~n15867 & n15869;
  assign n15871 = pi47  & n15870;
  assign n15872 = ~pi47  & ~n15870;
  assign n15873 = ~n15871 & ~n15872;
  assign n15874 = n15863 & ~n15873;
  assign n15875 = ~n15863 & n15873;
  assign n15876 = ~n15874 & ~n15875;
  assign n15877 = n15771 & ~n15876;
  assign n15878 = ~n15771 & n15876;
  assign n15879 = ~n15877 & ~n15878;
  assign n15880 = pi93  & n6331;
  assign n15881 = pi94  & n6015;
  assign n15882 = pi95  & n6010;
  assign n15883 = n3475 & n6008;
  assign n15884 = ~n15881 & ~n15882;
  assign n15885 = ~n15880 & n15884;
  assign n15886 = ~n15883 & n15885;
  assign n15887 = pi44  & n15886;
  assign n15888 = ~pi44  & ~n15886;
  assign n15889 = ~n15887 & ~n15888;
  assign n15890 = ~n15879 & n15889;
  assign n15891 = n15879 & ~n15889;
  assign n15892 = ~n15890 & ~n15891;
  assign n15893 = ~n15542 & ~n15546;
  assign n15894 = ~n15543 & ~n15893;
  assign n15895 = n15892 & n15894;
  assign n15896 = ~n15892 & ~n15894;
  assign n15897 = ~n15895 & ~n15896;
  assign n15898 = ~n15770 & n15897;
  assign n15899 = n15770 & ~n15897;
  assign n15900 = ~n15898 & ~n15899;
  assign n15901 = ~n15760 & n15900;
  assign n15902 = n15760 & ~n15900;
  assign n15903 = ~n15901 & ~n15902;
  assign n15904 = ~n15759 & n15903;
  assign n15905 = n15759 & ~n15903;
  assign n15906 = ~n15904 & ~n15905;
  assign n15907 = ~n15749 & n15906;
  assign n15908 = n15749 & ~n15906;
  assign n15909 = ~n15907 & ~n15908;
  assign n15910 = n15748 & ~n15909;
  assign n15911 = ~n15748 & n15909;
  assign n15912 = ~n15910 & ~n15911;
  assign n15913 = n15738 & n15912;
  assign n15914 = ~n15738 & ~n15912;
  assign n15915 = ~n15913 & ~n15914;
  assign n15916 = n15724 & n15915;
  assign n15917 = ~n15724 & ~n15915;
  assign n15918 = ~n15916 & ~n15917;
  assign n15919 = pi111  & n2510;
  assign n15920 = pi112  & n2342;
  assign n15921 = pi113  & n2337;
  assign n15922 = n2335 & n7852;
  assign n15923 = ~n15920 & ~n15921;
  assign n15924 = ~n15919 & n15923;
  assign n15925 = ~n15922 & n15924;
  assign n15926 = pi26  & n15925;
  assign n15927 = ~pi26  & ~n15925;
  assign n15928 = ~n15926 & ~n15927;
  assign n15929 = ~n15394 & ~n15597;
  assign n15930 = ~n15928 & ~n15929;
  assign n15931 = n15928 & n15929;
  assign n15932 = ~n15930 & ~n15931;
  assign n15933 = n15918 & n15932;
  assign n15934 = ~n15918 & ~n15932;
  assign n15935 = ~n15933 & ~n15934;
  assign n15936 = n15710 & n15935;
  assign n15937 = ~n15710 & ~n15935;
  assign n15938 = ~n15936 & ~n15937;
  assign n15939 = n15696 & n15938;
  assign n15940 = ~n15696 & ~n15938;
  assign n15941 = ~n15939 & ~n15940;
  assign n15942 = ~n15617 & ~n15620;
  assign n15943 = pi120  & n1296;
  assign n15944 = pi121  & n1207;
  assign n15945 = pi122  & n1202;
  assign n15946 = n1200 & n10729;
  assign n15947 = ~n15944 & ~n15945;
  assign n15948 = ~n15943 & n15947;
  assign n15949 = ~n15946 & n15948;
  assign n15950 = pi17  & n15949;
  assign n15951 = ~pi17  & ~n15949;
  assign n15952 = ~n15950 & ~n15951;
  assign n15953 = ~n15942 & ~n15952;
  assign n15954 = n15942 & n15952;
  assign n15955 = ~n15953 & ~n15954;
  assign n15956 = n15941 & n15955;
  assign n15957 = ~n15941 & ~n15955;
  assign n15958 = ~n15956 & ~n15957;
  assign n15959 = n15681 & n15958;
  assign n15960 = ~n15681 & ~n15958;
  assign n15961 = ~n15959 & ~n15960;
  assign n15962 = ~n15637 & ~n15640;
  assign n15963 = pi126  & n750;
  assign n15964 = pi127  & n651;
  assign n15965 = n644 & n12542;
  assign n15966 = ~n15963 & ~n15964;
  assign n15967 = ~n15965 & n15966;
  assign n15968 = pi11  & n15967;
  assign n15969 = ~pi11  & ~n15967;
  assign n15970 = ~n15968 & ~n15969;
  assign n15971 = ~n15962 & ~n15970;
  assign n15972 = n15962 & n15970;
  assign n15973 = ~n15971 & ~n15972;
  assign n15974 = n15961 & n15973;
  assign n15975 = ~n15961 & ~n15973;
  assign n15976 = ~n15974 & ~n15975;
  assign n15977 = ~n15667 & n15976;
  assign n15978 = n15667 & ~n15976;
  assign n15979 = ~n15977 & ~n15978;
  assign n15980 = ~n15666 & n15979;
  assign n15981 = n15666 & ~n15979;
  assign po73  = ~n15980 & ~n15981;
  assign n15983 = ~n15977 & ~n15980;
  assign n15984 = ~n15971 & ~n15974;
  assign n15985 = ~n15953 & ~n15956;
  assign n15986 = pi124  & n1006;
  assign n15987 = pi125  & n897;
  assign n15988 = pi126  & n892;
  assign n15989 = n890 & n12148;
  assign n15990 = ~n15987 & ~n15988;
  assign n15991 = ~n15986 & n15990;
  assign n15992 = ~n15989 & n15991;
  assign n15993 = pi14  & n15992;
  assign n15994 = ~pi14  & ~n15992;
  assign n15995 = ~n15993 & ~n15994;
  assign n15996 = ~n15985 & ~n15995;
  assign n15997 = n15985 & n15995;
  assign n15998 = ~n15996 & ~n15997;
  assign n15999 = pi121  & n1296;
  assign n16000 = pi122  & n1207;
  assign n16001 = pi123  & n1202;
  assign n16002 = n1200 & n10754;
  assign n16003 = ~n16000 & ~n16001;
  assign n16004 = ~n15999 & n16003;
  assign n16005 = ~n16002 & n16004;
  assign n16006 = pi17  & n16005;
  assign n16007 = ~pi17  & ~n16005;
  assign n16008 = ~n16006 & ~n16007;
  assign n16009 = ~n15695 & ~n15939;
  assign n16010 = n16008 & n16009;
  assign n16011 = ~n16008 & ~n16009;
  assign n16012 = ~n16010 & ~n16011;
  assign n16013 = pi118  & n1661;
  assign n16014 = pi119  & n1500;
  assign n16015 = pi120  & n1495;
  assign n16016 = n1493 & n10047;
  assign n16017 = ~n16014 & ~n16015;
  assign n16018 = ~n16013 & n16017;
  assign n16019 = ~n16016 & n16018;
  assign n16020 = pi20  & n16019;
  assign n16021 = ~pi20  & ~n16019;
  assign n16022 = ~n16020 & ~n16021;
  assign n16023 = ~n15709 & ~n15936;
  assign n16024 = ~n16022 & ~n16023;
  assign n16025 = n16022 & n16023;
  assign n16026 = ~n16024 & ~n16025;
  assign n16027 = ~n15722 & ~n15916;
  assign n16028 = pi112  & n2510;
  assign n16029 = pi113  & n2342;
  assign n16030 = pi114  & n2337;
  assign n16031 = n2335 & n8146;
  assign n16032 = ~n16029 & ~n16030;
  assign n16033 = ~n16028 & n16032;
  assign n16034 = ~n16031 & n16033;
  assign n16035 = pi26  & n16034;
  assign n16036 = ~pi26  & ~n16034;
  assign n16037 = ~n16035 & ~n16036;
  assign n16038 = ~n16027 & ~n16037;
  assign n16039 = n16027 & n16037;
  assign n16040 = ~n16038 & ~n16039;
  assign n16041 = pi109  & n3011;
  assign n16042 = pi110  & n2809;
  assign n16043 = pi111  & n2804;
  assign n16044 = n2802 & n7272;
  assign n16045 = ~n16042 & ~n16043;
  assign n16046 = ~n16041 & n16045;
  assign n16047 = ~n16044 & n16046;
  assign n16048 = pi29  & n16047;
  assign n16049 = ~pi29  & ~n16047;
  assign n16050 = ~n16048 & ~n16049;
  assign n16051 = ~n15737 & ~n15912;
  assign n16052 = ~n15736 & ~n16051;
  assign n16053 = n16050 & ~n16052;
  assign n16054 = ~n16050 & n16052;
  assign n16055 = ~n16053 & ~n16054;
  assign n16056 = pi106  & n3553;
  assign n16057 = pi107  & n3334;
  assign n16058 = pi108  & n3329;
  assign n16059 = n3327 & n6213;
  assign n16060 = ~n16057 & ~n16058;
  assign n16061 = ~n16056 & n16060;
  assign n16062 = ~n16059 & n16061;
  assign n16063 = pi32  & n16062;
  assign n16064 = ~pi32  & ~n16062;
  assign n16065 = ~n16063 & ~n16064;
  assign n16066 = n15748 & ~n15907;
  assign n16067 = ~n15908 & ~n16066;
  assign n16068 = ~n16065 & n16067;
  assign n16069 = n16065 & ~n16067;
  assign n16070 = ~n16068 & ~n16069;
  assign n16071 = pi103  & n4176;
  assign n16072 = pi104  & n3938;
  assign n16073 = pi105  & n3933;
  assign n16074 = n3931 & n5677;
  assign n16075 = ~n16072 & ~n16073;
  assign n16076 = ~n16071 & n16075;
  assign n16077 = ~n16074 & n16076;
  assign n16078 = pi35  & n16077;
  assign n16079 = ~pi35  & ~n16077;
  assign n16080 = ~n16078 & ~n16079;
  assign n16081 = ~n15901 & ~n15904;
  assign n16082 = ~n15895 & ~n15898;
  assign n16083 = pi88  & n7969;
  assign n16084 = pi89  & n7636;
  assign n16085 = pi90  & n7631;
  assign n16086 = n2448 & n7629;
  assign n16087 = ~n16084 & ~n16085;
  assign n16088 = ~n16083 & n16087;
  assign n16089 = ~n16086 & n16088;
  assign n16090 = pi50  & n16089;
  assign n16091 = ~pi50  & ~n16089;
  assign n16092 = ~n16090 & ~n16091;
  assign n16093 = pi85  & n8905;
  assign n16094 = pi86  & n8535;
  assign n16095 = pi87  & n8530;
  assign n16096 = n2116 & n8528;
  assign n16097 = ~n16094 & ~n16095;
  assign n16098 = ~n16093 & n16097;
  assign n16099 = ~n16096 & n16098;
  assign n16100 = pi53  & n16099;
  assign n16101 = ~pi53  & ~n16099;
  assign n16102 = ~n16100 & ~n16101;
  assign n16103 = pi79  & n10886;
  assign n16104 = pi80  & n10495;
  assign n16105 = pi81  & n10490;
  assign n16106 = n1337 & n10488;
  assign n16107 = ~n16104 & ~n16105;
  assign n16108 = ~n16103 & n16107;
  assign n16109 = ~n16106 & n16108;
  assign n16110 = pi59  & n16109;
  assign n16111 = ~pi59  & ~n16109;
  assign n16112 = ~n16110 & ~n16111;
  assign n16113 = pi76  & n11910;
  assign n16114 = pi77  & n11529;
  assign n16115 = pi78  & n11524;
  assign n16116 = n958 & n11522;
  assign n16117 = ~n16114 & ~n16115;
  assign n16118 = ~n16113 & n16117;
  assign n16119 = ~n16116 & n16118;
  assign n16120 = pi62  & n16119;
  assign n16121 = ~pi62  & ~n16119;
  assign n16122 = ~n16120 & ~n16121;
  assign n16123 = pi75  & n12277;
  assign n16124 = pi74  & n12276;
  assign n16125 = ~n16123 & ~n16124;
  assign n16126 = n15800 & ~n16125;
  assign n16127 = ~n15800 & n16125;
  assign n16128 = ~n16126 & ~n16127;
  assign n16129 = n15796 & ~n15801;
  assign n16130 = ~n15802 & ~n16129;
  assign n16131 = n16128 & n16130;
  assign n16132 = ~n16128 & ~n16130;
  assign n16133 = ~n16131 & ~n16132;
  assign n16134 = ~n16122 & n16133;
  assign n16135 = n16122 & ~n16133;
  assign n16136 = ~n16134 & ~n16135;
  assign n16137 = n16112 & ~n16136;
  assign n16138 = ~n16112 & n16136;
  assign n16139 = ~n16137 & ~n16138;
  assign n16140 = n15785 & ~n15807;
  assign n16141 = ~n15808 & ~n16140;
  assign n16142 = ~n16139 & ~n16141;
  assign n16143 = n16139 & n16141;
  assign n16144 = ~n16142 & ~n16143;
  assign n16145 = pi82  & n9858;
  assign n16146 = pi83  & n9508;
  assign n16147 = pi84  & n9503;
  assign n16148 = n1601 & n9501;
  assign n16149 = ~n16146 & ~n16147;
  assign n16150 = ~n16145 & n16149;
  assign n16151 = ~n16148 & n16150;
  assign n16152 = pi56  & n16151;
  assign n16153 = ~pi56  & ~n16151;
  assign n16154 = ~n16152 & ~n16153;
  assign n16155 = ~n16144 & n16154;
  assign n16156 = n16144 & ~n16154;
  assign n16157 = ~n16155 & ~n16156;
  assign n16158 = ~n15814 & n15825;
  assign n16159 = ~n15813 & ~n16158;
  assign n16160 = n16157 & n16159;
  assign n16161 = ~n16157 & ~n16159;
  assign n16162 = ~n16160 & ~n16161;
  assign n16163 = ~n16102 & n16162;
  assign n16164 = n16102 & ~n16162;
  assign n16165 = ~n16163 & ~n16164;
  assign n16166 = ~n15830 & n15841;
  assign n16167 = ~n15829 & ~n16166;
  assign n16168 = n16165 & n16167;
  assign n16169 = ~n16165 & ~n16167;
  assign n16170 = ~n16168 & ~n16169;
  assign n16171 = ~n16092 & n16170;
  assign n16172 = n16092 & ~n16170;
  assign n16173 = ~n16171 & ~n16172;
  assign n16174 = ~n15846 & n15857;
  assign n16175 = ~n15845 & ~n16174;
  assign n16176 = n16173 & n16175;
  assign n16177 = ~n16173 & ~n16175;
  assign n16178 = ~n16176 & ~n16177;
  assign n16179 = pi91  & n7121;
  assign n16180 = pi92  & n6795;
  assign n16181 = pi93  & n6790;
  assign n16182 = n2948 & n6788;
  assign n16183 = ~n16180 & ~n16181;
  assign n16184 = ~n16179 & n16183;
  assign n16185 = ~n16182 & n16184;
  assign n16186 = pi47  & n16185;
  assign n16187 = ~pi47  & ~n16185;
  assign n16188 = ~n16186 & ~n16187;
  assign n16189 = n16178 & ~n16188;
  assign n16190 = ~n16178 & n16188;
  assign n16191 = ~n16189 & ~n16190;
  assign n16192 = ~n15862 & n15873;
  assign n16193 = ~n15861 & ~n16192;
  assign n16194 = ~n16191 & ~n16193;
  assign n16195 = n16191 & n16193;
  assign n16196 = ~n16194 & ~n16195;
  assign n16197 = pi94  & n6331;
  assign n16198 = pi95  & n6015;
  assign n16199 = pi96  & n6010;
  assign n16200 = n3499 & n6008;
  assign n16201 = ~n16198 & ~n16199;
  assign n16202 = ~n16197 & n16201;
  assign n16203 = ~n16200 & n16202;
  assign n16204 = pi44  & n16203;
  assign n16205 = ~pi44  & ~n16203;
  assign n16206 = ~n16204 & ~n16205;
  assign n16207 = ~n16196 & n16206;
  assign n16208 = n16196 & ~n16206;
  assign n16209 = ~n16207 & ~n16208;
  assign n16210 = ~n15878 & ~n15891;
  assign n16211 = n16209 & ~n16210;
  assign n16212 = ~n16209 & n16210;
  assign n16213 = ~n16211 & ~n16212;
  assign n16214 = pi97  & n5558;
  assign n16215 = pi98  & n5293;
  assign n16216 = pi99  & n5288;
  assign n16217 = n4101 & n5286;
  assign n16218 = ~n16215 & ~n16216;
  assign n16219 = ~n16214 & n16218;
  assign n16220 = ~n16217 & n16219;
  assign n16221 = pi41  & n16220;
  assign n16222 = ~pi41  & ~n16220;
  assign n16223 = ~n16221 & ~n16222;
  assign n16224 = n16213 & ~n16223;
  assign n16225 = ~n16213 & n16223;
  assign n16226 = ~n16224 & ~n16225;
  assign n16227 = n16082 & ~n16226;
  assign n16228 = ~n16082 & n16226;
  assign n16229 = ~n16227 & ~n16228;
  assign n16230 = pi100  & n4843;
  assign n16231 = pi101  & n4598;
  assign n16232 = pi102  & n4593;
  assign n16233 = n4591 & n4956;
  assign n16234 = ~n16231 & ~n16232;
  assign n16235 = ~n16230 & n16234;
  assign n16236 = ~n16233 & n16235;
  assign n16237 = pi38  & n16236;
  assign n16238 = ~pi38  & ~n16236;
  assign n16239 = ~n16237 & ~n16238;
  assign n16240 = ~n16229 & n16239;
  assign n16241 = n16229 & ~n16239;
  assign n16242 = ~n16240 & ~n16241;
  assign n16243 = ~n16081 & n16242;
  assign n16244 = n16081 & ~n16242;
  assign n16245 = ~n16243 & ~n16244;
  assign n16246 = n16080 & ~n16245;
  assign n16247 = ~n16080 & n16245;
  assign n16248 = ~n16246 & ~n16247;
  assign n16249 = n16070 & n16248;
  assign n16250 = ~n16070 & ~n16248;
  assign n16251 = ~n16249 & ~n16250;
  assign n16252 = n16055 & n16251;
  assign n16253 = ~n16055 & ~n16251;
  assign n16254 = ~n16252 & ~n16253;
  assign n16255 = n16040 & n16254;
  assign n16256 = ~n16040 & ~n16254;
  assign n16257 = ~n16255 & ~n16256;
  assign n16258 = ~n15930 & ~n15933;
  assign n16259 = pi115  & n2053;
  assign n16260 = pi116  & n1893;
  assign n16261 = pi117  & n1888;
  assign n16262 = n1886 & n8784;
  assign n16263 = ~n16260 & ~n16261;
  assign n16264 = ~n16259 & n16263;
  assign n16265 = ~n16262 & n16264;
  assign n16266 = pi23  & n16265;
  assign n16267 = ~pi23  & ~n16265;
  assign n16268 = ~n16266 & ~n16267;
  assign n16269 = ~n16258 & ~n16268;
  assign n16270 = n16258 & n16268;
  assign n16271 = ~n16269 & ~n16270;
  assign n16272 = n16257 & n16271;
  assign n16273 = ~n16257 & ~n16271;
  assign n16274 = ~n16272 & ~n16273;
  assign n16275 = n16026 & n16274;
  assign n16276 = ~n16026 & ~n16274;
  assign n16277 = ~n16275 & ~n16276;
  assign n16278 = n16012 & n16277;
  assign n16279 = ~n16012 & ~n16277;
  assign n16280 = ~n16278 & ~n16279;
  assign n16281 = n15998 & n16280;
  assign n16282 = ~n15998 & ~n16280;
  assign n16283 = ~n16281 & ~n16282;
  assign n16284 = ~n15679 & ~n15959;
  assign n16285 = n644 & ~n12539;
  assign n16286 = ~n750 & ~n16285;
  assign n16287 = pi127  & ~n16286;
  assign n16288 = pi11  & ~n16287;
  assign n16289 = ~pi11  & n16287;
  assign n16290 = ~n16288 & ~n16289;
  assign n16291 = ~n16284 & ~n16290;
  assign n16292 = n16284 & n16290;
  assign n16293 = ~n16291 & ~n16292;
  assign n16294 = n16283 & n16293;
  assign n16295 = ~n16283 & ~n16293;
  assign n16296 = ~n16294 & ~n16295;
  assign n16297 = ~n15984 & n16296;
  assign n16298 = n15984 & ~n16296;
  assign n16299 = ~n16297 & ~n16298;
  assign n16300 = ~n15983 & n16299;
  assign n16301 = n15983 & ~n16299;
  assign po74  = ~n16300 & ~n16301;
  assign n16303 = ~n16297 & ~n16300;
  assign n16304 = ~n16291 & ~n16294;
  assign n16305 = pi119  & n1661;
  assign n16306 = pi120  & n1500;
  assign n16307 = pi121  & n1495;
  assign n16308 = n1493 & n10071;
  assign n16309 = ~n16306 & ~n16307;
  assign n16310 = ~n16305 & n16309;
  assign n16311 = ~n16308 & n16310;
  assign n16312 = pi20  & n16311;
  assign n16313 = ~pi20  & ~n16311;
  assign n16314 = ~n16312 & ~n16313;
  assign n16315 = ~n16024 & ~n16275;
  assign n16316 = n16314 & n16315;
  assign n16317 = ~n16314 & ~n16315;
  assign n16318 = ~n16316 & ~n16317;
  assign n16319 = pi113  & n2510;
  assign n16320 = pi114  & n2342;
  assign n16321 = pi115  & n2337;
  assign n16322 = n2335 & n8170;
  assign n16323 = ~n16320 & ~n16321;
  assign n16324 = ~n16319 & n16323;
  assign n16325 = ~n16322 & n16324;
  assign n16326 = pi26  & n16325;
  assign n16327 = ~pi26  & ~n16325;
  assign n16328 = ~n16326 & ~n16327;
  assign n16329 = ~n16038 & ~n16255;
  assign n16330 = n16328 & n16329;
  assign n16331 = ~n16328 & ~n16329;
  assign n16332 = ~n16330 & ~n16331;
  assign n16333 = pi104  & n4176;
  assign n16334 = pi105  & n3938;
  assign n16335 = pi106  & n3933;
  assign n16336 = n3931 & n5701;
  assign n16337 = ~n16334 & ~n16335;
  assign n16338 = ~n16333 & n16337;
  assign n16339 = ~n16336 & n16338;
  assign n16340 = pi35  & n16339;
  assign n16341 = ~pi35  & ~n16339;
  assign n16342 = ~n16340 & ~n16341;
  assign n16343 = ~n16228 & ~n16241;
  assign n16344 = pi98  & n5558;
  assign n16345 = pi99  & n5293;
  assign n16346 = pi100  & n5288;
  assign n16347 = n4501 & n5286;
  assign n16348 = ~n16345 & ~n16346;
  assign n16349 = ~n16344 & n16348;
  assign n16350 = ~n16347 & n16349;
  assign n16351 = pi41  & n16350;
  assign n16352 = ~pi41  & ~n16350;
  assign n16353 = ~n16351 & ~n16352;
  assign n16354 = ~n16195 & ~n16208;
  assign n16355 = pi95  & n6331;
  assign n16356 = pi96  & n6015;
  assign n16357 = pi97  & n6010;
  assign n16358 = n3691 & n6008;
  assign n16359 = ~n16356 & ~n16357;
  assign n16360 = ~n16355 & n16359;
  assign n16361 = ~n16358 & n16360;
  assign n16362 = pi44  & n16361;
  assign n16363 = ~pi44  & ~n16361;
  assign n16364 = ~n16362 & ~n16363;
  assign n16365 = ~n16168 & ~n16171;
  assign n16366 = pi89  & n7969;
  assign n16367 = pi90  & n7636;
  assign n16368 = pi91  & n7631;
  assign n16369 = n2746 & n7629;
  assign n16370 = ~n16367 & ~n16368;
  assign n16371 = ~n16366 & n16370;
  assign n16372 = ~n16369 & n16371;
  assign n16373 = pi50  & n16372;
  assign n16374 = ~pi50  & ~n16372;
  assign n16375 = ~n16373 & ~n16374;
  assign n16376 = ~n16160 & ~n16163;
  assign n16377 = pi86  & n8905;
  assign n16378 = pi87  & n8535;
  assign n16379 = pi88  & n8530;
  assign n16380 = n2140 & n8528;
  assign n16381 = ~n16378 & ~n16379;
  assign n16382 = ~n16377 & n16381;
  assign n16383 = ~n16380 & n16382;
  assign n16384 = pi53  & n16383;
  assign n16385 = ~pi53  & ~n16383;
  assign n16386 = ~n16384 & ~n16385;
  assign n16387 = ~n16143 & ~n16156;
  assign n16388 = pi80  & n10886;
  assign n16389 = pi81  & n10495;
  assign n16390 = pi82  & n10490;
  assign n16391 = n1450 & n10488;
  assign n16392 = ~n16389 & ~n16390;
  assign n16393 = ~n16388 & n16392;
  assign n16394 = ~n16391 & n16393;
  assign n16395 = pi59  & n16394;
  assign n16396 = ~pi59  & ~n16394;
  assign n16397 = ~n16395 & ~n16396;
  assign n16398 = ~n16126 & ~n16131;
  assign n16399 = pi77  & n11910;
  assign n16400 = pi78  & n11529;
  assign n16401 = pi79  & n11524;
  assign n16402 = n1048 & n11522;
  assign n16403 = ~n16400 & ~n16401;
  assign n16404 = ~n16399 & n16403;
  assign n16405 = ~n16402 & n16404;
  assign n16406 = pi62  & n16405;
  assign n16407 = ~pi62  & ~n16405;
  assign n16408 = ~n16406 & ~n16407;
  assign n16409 = ~pi11  & ~n15800;
  assign n16410 = pi11  & n15800;
  assign n16411 = ~n16409 & ~n16410;
  assign n16412 = pi76  & n12277;
  assign n16413 = pi75  & n12276;
  assign n16414 = ~n16412 & ~n16413;
  assign n16415 = n16411 & ~n16414;
  assign n16416 = ~n16411 & n16414;
  assign n16417 = ~n16415 & ~n16416;
  assign n16418 = ~n16408 & n16417;
  assign n16419 = n16408 & ~n16417;
  assign n16420 = ~n16418 & ~n16419;
  assign n16421 = ~n16398 & n16420;
  assign n16422 = n16398 & ~n16420;
  assign n16423 = ~n16421 & ~n16422;
  assign n16424 = ~n16397 & n16423;
  assign n16425 = n16397 & ~n16423;
  assign n16426 = ~n16424 & ~n16425;
  assign n16427 = n16112 & ~n16134;
  assign n16428 = ~n16135 & ~n16427;
  assign n16429 = ~n16426 & ~n16428;
  assign n16430 = n16426 & n16428;
  assign n16431 = ~n16429 & ~n16430;
  assign n16432 = pi83  & n9858;
  assign n16433 = pi84  & n9508;
  assign n16434 = pi85  & n9503;
  assign n16435 = n1831 & n9501;
  assign n16436 = ~n16433 & ~n16434;
  assign n16437 = ~n16432 & n16436;
  assign n16438 = ~n16435 & n16437;
  assign n16439 = pi56  & n16438;
  assign n16440 = ~pi56  & ~n16438;
  assign n16441 = ~n16439 & ~n16440;
  assign n16442 = n16431 & ~n16441;
  assign n16443 = ~n16431 & n16441;
  assign n16444 = ~n16442 & ~n16443;
  assign n16445 = ~n16387 & n16444;
  assign n16446 = n16387 & ~n16444;
  assign n16447 = ~n16445 & ~n16446;
  assign n16448 = ~n16386 & n16447;
  assign n16449 = n16386 & ~n16447;
  assign n16450 = ~n16448 & ~n16449;
  assign n16451 = ~n16376 & n16450;
  assign n16452 = n16376 & ~n16450;
  assign n16453 = ~n16451 & ~n16452;
  assign n16454 = ~n16375 & n16453;
  assign n16455 = n16375 & ~n16453;
  assign n16456 = ~n16454 & ~n16455;
  assign n16457 = n16365 & ~n16456;
  assign n16458 = ~n16365 & n16456;
  assign n16459 = ~n16457 & ~n16458;
  assign n16460 = pi92  & n7121;
  assign n16461 = pi93  & n6795;
  assign n16462 = pi94  & n6790;
  assign n16463 = n3280 & n6788;
  assign n16464 = ~n16461 & ~n16462;
  assign n16465 = ~n16460 & n16464;
  assign n16466 = ~n16463 & n16465;
  assign n16467 = pi47  & n16466;
  assign n16468 = ~pi47  & ~n16466;
  assign n16469 = ~n16467 & ~n16468;
  assign n16470 = n16459 & ~n16469;
  assign n16471 = ~n16459 & n16469;
  assign n16472 = ~n16470 & ~n16471;
  assign n16473 = ~n16176 & n16188;
  assign n16474 = ~n16177 & ~n16473;
  assign n16475 = n16472 & ~n16474;
  assign n16476 = ~n16472 & n16474;
  assign n16477 = ~n16475 & ~n16476;
  assign n16478 = ~n16364 & ~n16477;
  assign n16479 = n16364 & n16477;
  assign n16480 = ~n16478 & ~n16479;
  assign n16481 = ~n16354 & n16480;
  assign n16482 = n16354 & ~n16480;
  assign n16483 = ~n16481 & ~n16482;
  assign n16484 = ~n16353 & n16483;
  assign n16485 = n16353 & ~n16483;
  assign n16486 = ~n16484 & ~n16485;
  assign n16487 = ~n16212 & ~n16223;
  assign n16488 = ~n16211 & ~n16487;
  assign n16489 = ~n16486 & n16488;
  assign n16490 = n16486 & ~n16488;
  assign n16491 = ~n16489 & ~n16490;
  assign n16492 = pi101  & n4843;
  assign n16493 = pi102  & n4598;
  assign n16494 = pi103  & n4593;
  assign n16495 = n4591 & n5188;
  assign n16496 = ~n16493 & ~n16494;
  assign n16497 = ~n16492 & n16496;
  assign n16498 = ~n16495 & n16497;
  assign n16499 = pi38  & n16498;
  assign n16500 = ~pi38  & ~n16498;
  assign n16501 = ~n16499 & ~n16500;
  assign n16502 = n16491 & ~n16501;
  assign n16503 = ~n16491 & n16501;
  assign n16504 = ~n16502 & ~n16503;
  assign n16505 = ~n16343 & n16504;
  assign n16506 = n16343 & ~n16504;
  assign n16507 = ~n16505 & ~n16506;
  assign n16508 = ~n16342 & n16507;
  assign n16509 = n16342 & ~n16507;
  assign n16510 = ~n16508 & ~n16509;
  assign n16511 = n16080 & ~n16243;
  assign n16512 = ~n16244 & ~n16511;
  assign n16513 = ~n16510 & ~n16512;
  assign n16514 = n16510 & n16512;
  assign n16515 = ~n16513 & ~n16514;
  assign n16516 = pi107  & n3553;
  assign n16517 = pi108  & n3334;
  assign n16518 = pi109  & n3329;
  assign n16519 = n3327 & n6715;
  assign n16520 = ~n16517 & ~n16518;
  assign n16521 = ~n16516 & n16520;
  assign n16522 = ~n16519 & n16521;
  assign n16523 = pi32  & n16522;
  assign n16524 = ~pi32  & ~n16522;
  assign n16525 = ~n16523 & ~n16524;
  assign n16526 = ~n16068 & ~n16248;
  assign n16527 = ~n16069 & ~n16526;
  assign n16528 = ~n16525 & n16527;
  assign n16529 = n16525 & ~n16527;
  assign n16530 = ~n16528 & ~n16529;
  assign n16531 = n16515 & n16530;
  assign n16532 = ~n16515 & ~n16530;
  assign n16533 = ~n16531 & ~n16532;
  assign n16534 = ~n16054 & ~n16252;
  assign n16535 = pi110  & n3011;
  assign n16536 = pi111  & n2809;
  assign n16537 = pi112  & n2804;
  assign n16538 = n2802 & n7296;
  assign n16539 = ~n16536 & ~n16537;
  assign n16540 = ~n16535 & n16539;
  assign n16541 = ~n16538 & n16540;
  assign n16542 = pi29  & n16541;
  assign n16543 = ~pi29  & ~n16541;
  assign n16544 = ~n16542 & ~n16543;
  assign n16545 = ~n16534 & ~n16544;
  assign n16546 = n16534 & n16544;
  assign n16547 = ~n16545 & ~n16546;
  assign n16548 = n16533 & n16547;
  assign n16549 = ~n16533 & ~n16547;
  assign n16550 = ~n16548 & ~n16549;
  assign n16551 = n16332 & n16550;
  assign n16552 = ~n16332 & ~n16550;
  assign n16553 = ~n16551 & ~n16552;
  assign n16554 = ~n16269 & ~n16272;
  assign n16555 = pi116  & n2053;
  assign n16556 = pi117  & n1893;
  assign n16557 = pi118  & n1888;
  assign n16558 = n1886 & n9095;
  assign n16559 = ~n16556 & ~n16557;
  assign n16560 = ~n16555 & n16559;
  assign n16561 = ~n16558 & n16560;
  assign n16562 = pi23  & n16561;
  assign n16563 = ~pi23  & ~n16561;
  assign n16564 = ~n16562 & ~n16563;
  assign n16565 = ~n16554 & ~n16564;
  assign n16566 = n16554 & n16564;
  assign n16567 = ~n16565 & ~n16566;
  assign n16568 = n16553 & n16567;
  assign n16569 = ~n16553 & ~n16567;
  assign n16570 = ~n16568 & ~n16569;
  assign n16571 = n16318 & n16570;
  assign n16572 = ~n16318 & ~n16570;
  assign n16573 = ~n16571 & ~n16572;
  assign n16574 = ~n16011 & ~n16278;
  assign n16575 = pi122  & n1296;
  assign n16576 = pi123  & n1207;
  assign n16577 = pi124  & n1202;
  assign n16578 = n1200 & n11099;
  assign n16579 = ~n16576 & ~n16577;
  assign n16580 = ~n16575 & n16579;
  assign n16581 = ~n16578 & n16580;
  assign n16582 = pi17  & n16581;
  assign n16583 = ~pi17  & ~n16581;
  assign n16584 = ~n16582 & ~n16583;
  assign n16585 = ~n16574 & ~n16584;
  assign n16586 = n16574 & n16584;
  assign n16587 = ~n16585 & ~n16586;
  assign n16588 = n16573 & n16587;
  assign n16589 = ~n16573 & ~n16587;
  assign n16590 = ~n16588 & ~n16589;
  assign n16591 = ~n15996 & ~n16281;
  assign n16592 = pi125  & n1006;
  assign n16593 = pi126  & n897;
  assign n16594 = pi127  & n892;
  assign n16595 = n890 & n12519;
  assign n16596 = ~n16593 & ~n16594;
  assign n16597 = ~n16592 & n16596;
  assign n16598 = ~n16595 & n16597;
  assign n16599 = pi14  & n16598;
  assign n16600 = ~pi14  & ~n16598;
  assign n16601 = ~n16599 & ~n16600;
  assign n16602 = ~n16591 & ~n16601;
  assign n16603 = n16591 & n16601;
  assign n16604 = ~n16602 & ~n16603;
  assign n16605 = n16590 & n16604;
  assign n16606 = ~n16590 & ~n16604;
  assign n16607 = ~n16605 & ~n16606;
  assign n16608 = ~n16304 & n16607;
  assign n16609 = n16304 & ~n16607;
  assign n16610 = ~n16608 & ~n16609;
  assign n16611 = ~n16303 & n16610;
  assign n16612 = n16303 & ~n16610;
  assign po75  = ~n16611 & ~n16612;
  assign n16614 = ~n16608 & ~n16611;
  assign n16615 = ~n16602 & ~n16605;
  assign n16616 = pi123  & n1296;
  assign n16617 = pi124  & n1207;
  assign n16618 = pi125  & n1202;
  assign n16619 = n1200 & n11786;
  assign n16620 = ~n16617 & ~n16618;
  assign n16621 = ~n16616 & n16620;
  assign n16622 = ~n16619 & n16621;
  assign n16623 = pi17  & n16622;
  assign n16624 = ~pi17  & ~n16622;
  assign n16625 = ~n16623 & ~n16624;
  assign n16626 = ~n16317 & ~n16571;
  assign n16627 = ~n16625 & ~n16626;
  assign n16628 = n16625 & n16626;
  assign n16629 = ~n16627 & ~n16628;
  assign n16630 = ~n16545 & ~n16548;
  assign n16631 = pi114  & n2510;
  assign n16632 = pi115  & n2342;
  assign n16633 = pi116  & n2337;
  assign n16634 = n2335 & n8470;
  assign n16635 = ~n16632 & ~n16633;
  assign n16636 = ~n16631 & n16635;
  assign n16637 = ~n16634 & n16636;
  assign n16638 = pi26  & n16637;
  assign n16639 = ~pi26  & ~n16637;
  assign n16640 = ~n16638 & ~n16639;
  assign n16641 = ~n16630 & ~n16640;
  assign n16642 = n16630 & n16640;
  assign n16643 = ~n16641 & ~n16642;
  assign n16644 = ~n16508 & ~n16514;
  assign n16645 = pi108  & n3553;
  assign n16646 = pi109  & n3334;
  assign n16647 = pi110  & n3329;
  assign n16648 = n3327 & n6995;
  assign n16649 = ~n16646 & ~n16647;
  assign n16650 = ~n16645 & n16649;
  assign n16651 = ~n16648 & n16650;
  assign n16652 = pi32  & n16651;
  assign n16653 = ~pi32  & ~n16651;
  assign n16654 = ~n16652 & ~n16653;
  assign n16655 = ~n16644 & ~n16654;
  assign n16656 = n16644 & n16654;
  assign n16657 = ~n16655 & ~n16656;
  assign n16658 = ~n16502 & ~n16505;
  assign n16659 = pi102  & n4843;
  assign n16660 = pi103  & n4598;
  assign n16661 = pi104  & n4593;
  assign n16662 = n4591 & n5212;
  assign n16663 = ~n16660 & ~n16661;
  assign n16664 = ~n16659 & n16663;
  assign n16665 = ~n16662 & n16664;
  assign n16666 = pi38  & n16665;
  assign n16667 = ~pi38  & ~n16665;
  assign n16668 = ~n16666 & ~n16667;
  assign n16669 = ~n16484 & ~n16490;
  assign n16670 = pi99  & n5558;
  assign n16671 = pi100  & n5293;
  assign n16672 = pi101  & n5288;
  assign n16673 = n4730 & n5286;
  assign n16674 = ~n16671 & ~n16672;
  assign n16675 = ~n16670 & n16674;
  assign n16676 = ~n16673 & n16675;
  assign n16677 = pi41  & n16676;
  assign n16678 = ~pi41  & ~n16676;
  assign n16679 = ~n16677 & ~n16678;
  assign n16680 = ~n16478 & ~n16481;
  assign n16681 = pi96  & n6331;
  assign n16682 = pi97  & n6015;
  assign n16683 = pi98  & n6010;
  assign n16684 = n3889 & n6008;
  assign n16685 = ~n16682 & ~n16683;
  assign n16686 = ~n16681 & n16685;
  assign n16687 = ~n16684 & n16686;
  assign n16688 = pi44  & n16687;
  assign n16689 = ~pi44  & ~n16687;
  assign n16690 = ~n16688 & ~n16689;
  assign n16691 = pi93  & n7121;
  assign n16692 = pi94  & n6795;
  assign n16693 = pi95  & n6790;
  assign n16694 = n3475 & n6788;
  assign n16695 = ~n16692 & ~n16693;
  assign n16696 = ~n16691 & n16695;
  assign n16697 = ~n16694 & n16696;
  assign n16698 = pi47  & n16697;
  assign n16699 = ~pi47  & ~n16697;
  assign n16700 = ~n16698 & ~n16699;
  assign n16701 = ~n16454 & ~n16458;
  assign n16702 = ~n16448 & ~n16451;
  assign n16703 = ~n16442 & ~n16445;
  assign n16704 = ~n16424 & ~n16430;
  assign n16705 = ~n16418 & ~n16421;
  assign n16706 = pi78  & n11910;
  assign n16707 = pi79  & n11529;
  assign n16708 = pi80  & n11524;
  assign n16709 = n1144 & n11522;
  assign n16710 = ~n16707 & ~n16708;
  assign n16711 = ~n16706 & n16710;
  assign n16712 = ~n16709 & n16711;
  assign n16713 = pi62  & n16712;
  assign n16714 = ~pi62  & ~n16712;
  assign n16715 = ~n16713 & ~n16714;
  assign n16716 = ~n16409 & ~n16415;
  assign n16717 = pi77  & n12277;
  assign n16718 = pi76  & n12276;
  assign n16719 = ~n16717 & ~n16718;
  assign n16720 = ~n16716 & n16719;
  assign n16721 = n16716 & ~n16719;
  assign n16722 = ~n16720 & ~n16721;
  assign n16723 = ~n16715 & n16722;
  assign n16724 = n16715 & ~n16722;
  assign n16725 = ~n16723 & ~n16724;
  assign n16726 = n16705 & ~n16725;
  assign n16727 = ~n16705 & n16725;
  assign n16728 = ~n16726 & ~n16727;
  assign n16729 = pi81  & n10886;
  assign n16730 = pi82  & n10495;
  assign n16731 = pi83  & n10490;
  assign n16732 = n1577 & n10488;
  assign n16733 = ~n16730 & ~n16731;
  assign n16734 = ~n16729 & n16733;
  assign n16735 = ~n16732 & n16734;
  assign n16736 = pi59  & n16735;
  assign n16737 = ~pi59  & ~n16735;
  assign n16738 = ~n16736 & ~n16737;
  assign n16739 = n16728 & ~n16738;
  assign n16740 = ~n16728 & n16738;
  assign n16741 = ~n16739 & ~n16740;
  assign n16742 = n16704 & ~n16741;
  assign n16743 = ~n16704 & n16741;
  assign n16744 = ~n16742 & ~n16743;
  assign n16745 = pi84  & n9858;
  assign n16746 = pi85  & n9508;
  assign n16747 = pi86  & n9503;
  assign n16748 = n1975 & n9501;
  assign n16749 = ~n16746 & ~n16747;
  assign n16750 = ~n16745 & n16749;
  assign n16751 = ~n16748 & n16750;
  assign n16752 = pi56  & n16751;
  assign n16753 = ~pi56  & ~n16751;
  assign n16754 = ~n16752 & ~n16753;
  assign n16755 = n16744 & ~n16754;
  assign n16756 = ~n16744 & n16754;
  assign n16757 = ~n16755 & ~n16756;
  assign n16758 = n16703 & ~n16757;
  assign n16759 = ~n16703 & n16757;
  assign n16760 = ~n16758 & ~n16759;
  assign n16761 = pi87  & n8905;
  assign n16762 = pi88  & n8535;
  assign n16763 = pi89  & n8530;
  assign n16764 = n2287 & n8528;
  assign n16765 = ~n16762 & ~n16763;
  assign n16766 = ~n16761 & n16765;
  assign n16767 = ~n16764 & n16766;
  assign n16768 = pi53  & n16767;
  assign n16769 = ~pi53  & ~n16767;
  assign n16770 = ~n16768 & ~n16769;
  assign n16771 = n16760 & ~n16770;
  assign n16772 = ~n16760 & n16770;
  assign n16773 = ~n16771 & ~n16772;
  assign n16774 = n16702 & ~n16773;
  assign n16775 = ~n16702 & n16773;
  assign n16776 = ~n16774 & ~n16775;
  assign n16777 = pi90  & n7969;
  assign n16778 = pi91  & n7636;
  assign n16779 = pi92  & n7631;
  assign n16780 = n2924 & n7629;
  assign n16781 = ~n16778 & ~n16779;
  assign n16782 = ~n16777 & n16781;
  assign n16783 = ~n16780 & n16782;
  assign n16784 = pi50  & n16783;
  assign n16785 = ~pi50  & ~n16783;
  assign n16786 = ~n16784 & ~n16785;
  assign n16787 = ~n16776 & n16786;
  assign n16788 = n16776 & ~n16786;
  assign n16789 = ~n16787 & ~n16788;
  assign n16790 = ~n16701 & n16789;
  assign n16791 = n16701 & ~n16789;
  assign n16792 = ~n16790 & ~n16791;
  assign n16793 = ~n16700 & n16792;
  assign n16794 = n16700 & ~n16792;
  assign n16795 = ~n16793 & ~n16794;
  assign n16796 = ~n16470 & ~n16474;
  assign n16797 = ~n16471 & ~n16796;
  assign n16798 = n16795 & n16797;
  assign n16799 = ~n16795 & ~n16797;
  assign n16800 = ~n16798 & ~n16799;
  assign n16801 = ~n16690 & n16800;
  assign n16802 = n16690 & ~n16800;
  assign n16803 = ~n16801 & ~n16802;
  assign n16804 = ~n16680 & n16803;
  assign n16805 = n16680 & ~n16803;
  assign n16806 = ~n16804 & ~n16805;
  assign n16807 = ~n16679 & n16806;
  assign n16808 = n16679 & ~n16806;
  assign n16809 = ~n16807 & ~n16808;
  assign n16810 = ~n16669 & n16809;
  assign n16811 = n16669 & ~n16809;
  assign n16812 = ~n16810 & ~n16811;
  assign n16813 = ~n16668 & n16812;
  assign n16814 = n16668 & ~n16812;
  assign n16815 = ~n16813 & ~n16814;
  assign n16816 = ~n16658 & n16815;
  assign n16817 = n16658 & ~n16815;
  assign n16818 = ~n16816 & ~n16817;
  assign n16819 = pi105  & n4176;
  assign n16820 = pi106  & n3938;
  assign n16821 = pi107  & n3933;
  assign n16822 = n3931 & n6189;
  assign n16823 = ~n16820 & ~n16821;
  assign n16824 = ~n16819 & n16823;
  assign n16825 = ~n16822 & n16824;
  assign n16826 = pi35  & n16825;
  assign n16827 = ~pi35  & ~n16825;
  assign n16828 = ~n16826 & ~n16827;
  assign n16829 = n16818 & ~n16828;
  assign n16830 = ~n16818 & n16828;
  assign n16831 = ~n16829 & ~n16830;
  assign n16832 = n16657 & n16831;
  assign n16833 = ~n16657 & ~n16831;
  assign n16834 = ~n16832 & ~n16833;
  assign n16835 = pi111  & n3011;
  assign n16836 = pi112  & n2809;
  assign n16837 = pi113  & n2804;
  assign n16838 = n2802 & n7852;
  assign n16839 = ~n16836 & ~n16837;
  assign n16840 = ~n16835 & n16839;
  assign n16841 = ~n16838 & n16840;
  assign n16842 = pi29  & n16841;
  assign n16843 = ~pi29  & ~n16841;
  assign n16844 = ~n16842 & ~n16843;
  assign n16845 = ~n16528 & ~n16531;
  assign n16846 = ~n16844 & ~n16845;
  assign n16847 = n16844 & n16845;
  assign n16848 = ~n16846 & ~n16847;
  assign n16849 = n16834 & n16848;
  assign n16850 = ~n16834 & ~n16848;
  assign n16851 = ~n16849 & ~n16850;
  assign n16852 = ~n16643 & n16851;
  assign n16853 = n16643 & ~n16851;
  assign n16854 = ~n16852 & ~n16853;
  assign n16855 = pi117  & n2053;
  assign n16856 = pi118  & n1893;
  assign n16857 = pi119  & n1888;
  assign n16858 = n1886 & n9412;
  assign n16859 = ~n16856 & ~n16857;
  assign n16860 = ~n16855 & n16859;
  assign n16861 = ~n16858 & n16860;
  assign n16862 = pi23  & n16861;
  assign n16863 = ~pi23  & ~n16861;
  assign n16864 = ~n16862 & ~n16863;
  assign n16865 = ~n16331 & ~n16551;
  assign n16866 = ~n16864 & ~n16865;
  assign n16867 = n16864 & n16865;
  assign n16868 = ~n16866 & ~n16867;
  assign n16869 = ~n16854 & n16868;
  assign n16870 = n16854 & ~n16868;
  assign n16871 = ~n16869 & ~n16870;
  assign n16872 = ~n16565 & ~n16568;
  assign n16873 = pi120  & n1661;
  assign n16874 = pi121  & n1500;
  assign n16875 = pi122  & n1495;
  assign n16876 = n1493 & n10729;
  assign n16877 = ~n16874 & ~n16875;
  assign n16878 = ~n16873 & n16877;
  assign n16879 = ~n16876 & n16878;
  assign n16880 = pi20  & n16879;
  assign n16881 = ~pi20  & ~n16879;
  assign n16882 = ~n16880 & ~n16881;
  assign n16883 = ~n16872 & ~n16882;
  assign n16884 = n16872 & n16882;
  assign n16885 = ~n16883 & ~n16884;
  assign n16886 = n16871 & n16885;
  assign n16887 = ~n16871 & ~n16885;
  assign n16888 = ~n16886 & ~n16887;
  assign n16889 = n16629 & n16888;
  assign n16890 = ~n16629 & ~n16888;
  assign n16891 = ~n16889 & ~n16890;
  assign n16892 = ~n16585 & ~n16588;
  assign n16893 = pi126  & n1006;
  assign n16894 = pi127  & n897;
  assign n16895 = n890 & n12542;
  assign n16896 = ~n16893 & ~n16894;
  assign n16897 = ~n16895 & n16896;
  assign n16898 = pi14  & n16897;
  assign n16899 = ~pi14  & ~n16897;
  assign n16900 = ~n16898 & ~n16899;
  assign n16901 = ~n16892 & ~n16900;
  assign n16902 = n16892 & n16900;
  assign n16903 = ~n16901 & ~n16902;
  assign n16904 = n16891 & n16903;
  assign n16905 = ~n16891 & ~n16903;
  assign n16906 = ~n16904 & ~n16905;
  assign n16907 = ~n16615 & n16906;
  assign n16908 = n16615 & ~n16906;
  assign n16909 = ~n16907 & ~n16908;
  assign n16910 = ~n16614 & n16909;
  assign n16911 = n16614 & ~n16909;
  assign po76  = ~n16910 & ~n16911;
  assign n16913 = ~n16907 & ~n16910;
  assign n16914 = ~n16901 & ~n16904;
  assign n16915 = pi121  & n1661;
  assign n16916 = pi122  & n1500;
  assign n16917 = pi123  & n1495;
  assign n16918 = n1493 & n10754;
  assign n16919 = ~n16916 & ~n16917;
  assign n16920 = ~n16915 & n16919;
  assign n16921 = ~n16918 & n16920;
  assign n16922 = pi20  & n16921;
  assign n16923 = ~pi20  & ~n16921;
  assign n16924 = ~n16922 & ~n16923;
  assign n16925 = ~n16866 & ~n16869;
  assign n16926 = n16924 & n16925;
  assign n16927 = ~n16924 & ~n16925;
  assign n16928 = ~n16926 & ~n16927;
  assign n16929 = pi118  & n2053;
  assign n16930 = pi119  & n1893;
  assign n16931 = pi120  & n1888;
  assign n16932 = n1886 & n10047;
  assign n16933 = ~n16930 & ~n16931;
  assign n16934 = ~n16929 & n16933;
  assign n16935 = ~n16932 & n16934;
  assign n16936 = pi23  & n16935;
  assign n16937 = ~pi23  & ~n16935;
  assign n16938 = ~n16936 & ~n16937;
  assign n16939 = ~n16641 & ~n16851;
  assign n16940 = ~n16642 & ~n16939;
  assign n16941 = n16938 & ~n16940;
  assign n16942 = ~n16938 & n16940;
  assign n16943 = ~n16941 & ~n16942;
  assign n16944 = pi115  & n2510;
  assign n16945 = pi116  & n2342;
  assign n16946 = pi117  & n2337;
  assign n16947 = n2335 & n8784;
  assign n16948 = ~n16945 & ~n16946;
  assign n16949 = ~n16944 & n16948;
  assign n16950 = ~n16947 & n16949;
  assign n16951 = pi26  & n16950;
  assign n16952 = ~pi26  & ~n16950;
  assign n16953 = ~n16951 & ~n16952;
  assign n16954 = ~n16846 & ~n16849;
  assign n16955 = n16953 & n16954;
  assign n16956 = ~n16953 & ~n16954;
  assign n16957 = ~n16955 & ~n16956;
  assign n16958 = ~n16655 & ~n16832;
  assign n16959 = pi112  & n3011;
  assign n16960 = pi113  & n2809;
  assign n16961 = pi114  & n2804;
  assign n16962 = n2802 & n8146;
  assign n16963 = ~n16960 & ~n16961;
  assign n16964 = ~n16959 & n16963;
  assign n16965 = ~n16962 & n16964;
  assign n16966 = pi29  & n16965;
  assign n16967 = ~pi29  & ~n16965;
  assign n16968 = ~n16966 & ~n16967;
  assign n16969 = ~n16958 & ~n16968;
  assign n16970 = n16958 & n16968;
  assign n16971 = ~n16969 & ~n16970;
  assign n16972 = pi109  & n3553;
  assign n16973 = pi110  & n3334;
  assign n16974 = pi111  & n3329;
  assign n16975 = n3327 & n7272;
  assign n16976 = ~n16973 & ~n16974;
  assign n16977 = ~n16972 & n16976;
  assign n16978 = ~n16975 & n16977;
  assign n16979 = pi32  & n16978;
  assign n16980 = ~pi32  & ~n16978;
  assign n16981 = ~n16979 & ~n16980;
  assign n16982 = ~n16816 & n16828;
  assign n16983 = ~n16817 & ~n16982;
  assign n16984 = ~n16981 & n16983;
  assign n16985 = n16981 & ~n16983;
  assign n16986 = ~n16984 & ~n16985;
  assign n16987 = pi106  & n4176;
  assign n16988 = pi107  & n3938;
  assign n16989 = pi108  & n3933;
  assign n16990 = n3931 & n6213;
  assign n16991 = ~n16988 & ~n16989;
  assign n16992 = ~n16987 & n16991;
  assign n16993 = ~n16990 & n16992;
  assign n16994 = pi35  & n16993;
  assign n16995 = ~pi35  & ~n16993;
  assign n16996 = ~n16994 & ~n16995;
  assign n16997 = ~n16810 & ~n16813;
  assign n16998 = pi103  & n4843;
  assign n16999 = pi104  & n4598;
  assign n17000 = pi105  & n4593;
  assign n17001 = n4591 & n5677;
  assign n17002 = ~n16999 & ~n17000;
  assign n17003 = ~n16998 & n17002;
  assign n17004 = ~n17001 & n17003;
  assign n17005 = pi38  & n17004;
  assign n17006 = ~pi38  & ~n17004;
  assign n17007 = ~n17005 & ~n17006;
  assign n17008 = ~n16804 & ~n16807;
  assign n17009 = ~n16798 & ~n16801;
  assign n17010 = ~n16790 & ~n16793;
  assign n17011 = pi94  & n7121;
  assign n17012 = pi95  & n6795;
  assign n17013 = pi96  & n6790;
  assign n17014 = n3499 & n6788;
  assign n17015 = ~n17012 & ~n17013;
  assign n17016 = ~n17011 & n17015;
  assign n17017 = ~n17014 & n17016;
  assign n17018 = pi47  & n17017;
  assign n17019 = ~pi47  & ~n17017;
  assign n17020 = ~n17018 & ~n17019;
  assign n17021 = ~n16775 & ~n16788;
  assign n17022 = pi88  & n8905;
  assign n17023 = pi89  & n8535;
  assign n17024 = pi90  & n8530;
  assign n17025 = n2448 & n8528;
  assign n17026 = ~n17023 & ~n17024;
  assign n17027 = ~n17022 & n17026;
  assign n17028 = ~n17025 & n17027;
  assign n17029 = pi53  & n17028;
  assign n17030 = ~pi53  & ~n17028;
  assign n17031 = ~n17029 & ~n17030;
  assign n17032 = ~n16720 & ~n16723;
  assign n17033 = pi78  & n12277;
  assign n17034 = pi77  & n12276;
  assign n17035 = ~n17033 & ~n17034;
  assign n17036 = n16719 & ~n17035;
  assign n17037 = ~n16719 & n17035;
  assign n17038 = ~n17036 & ~n17037;
  assign n17039 = pi79  & n11910;
  assign n17040 = pi80  & n11529;
  assign n17041 = pi81  & n11524;
  assign n17042 = n1337 & n11522;
  assign n17043 = ~n17040 & ~n17041;
  assign n17044 = ~n17039 & n17043;
  assign n17045 = ~n17042 & n17044;
  assign n17046 = pi62  & n17045;
  assign n17047 = ~pi62  & ~n17045;
  assign n17048 = ~n17046 & ~n17047;
  assign n17049 = n17038 & ~n17048;
  assign n17050 = ~n17038 & n17048;
  assign n17051 = ~n17049 & ~n17050;
  assign n17052 = ~n17032 & n17051;
  assign n17053 = n17032 & ~n17051;
  assign n17054 = ~n17052 & ~n17053;
  assign n17055 = pi82  & n10886;
  assign n17056 = pi83  & n10495;
  assign n17057 = pi84  & n10490;
  assign n17058 = n1601 & n10488;
  assign n17059 = ~n17056 & ~n17057;
  assign n17060 = ~n17055 & n17059;
  assign n17061 = ~n17058 & n17060;
  assign n17062 = pi59  & n17061;
  assign n17063 = ~pi59  & ~n17061;
  assign n17064 = ~n17062 & ~n17063;
  assign n17065 = n17054 & ~n17064;
  assign n17066 = ~n17054 & n17064;
  assign n17067 = ~n17065 & ~n17066;
  assign n17068 = ~n16727 & n16738;
  assign n17069 = ~n16726 & ~n17068;
  assign n17070 = ~n17067 & ~n17069;
  assign n17071 = n17067 & n17069;
  assign n17072 = ~n17070 & ~n17071;
  assign n17073 = pi85  & n9858;
  assign n17074 = pi86  & n9508;
  assign n17075 = pi87  & n9503;
  assign n17076 = n2116 & n9501;
  assign n17077 = ~n17074 & ~n17075;
  assign n17078 = ~n17073 & n17077;
  assign n17079 = ~n17076 & n17078;
  assign n17080 = pi56  & n17079;
  assign n17081 = ~pi56  & ~n17079;
  assign n17082 = ~n17080 & ~n17081;
  assign n17083 = ~n17072 & n17082;
  assign n17084 = n17072 & ~n17082;
  assign n17085 = ~n17083 & ~n17084;
  assign n17086 = ~n16743 & n16754;
  assign n17087 = ~n16742 & ~n17086;
  assign n17088 = n17085 & n17087;
  assign n17089 = ~n17085 & ~n17087;
  assign n17090 = ~n17088 & ~n17089;
  assign n17091 = ~n17031 & n17090;
  assign n17092 = n17031 & ~n17090;
  assign n17093 = ~n17091 & ~n17092;
  assign n17094 = ~n16759 & n16770;
  assign n17095 = ~n16758 & ~n17094;
  assign n17096 = n17093 & n17095;
  assign n17097 = ~n17093 & ~n17095;
  assign n17098 = ~n17096 & ~n17097;
  assign n17099 = pi91  & n7969;
  assign n17100 = pi92  & n7636;
  assign n17101 = pi93  & n7631;
  assign n17102 = n2948 & n7629;
  assign n17103 = ~n17100 & ~n17101;
  assign n17104 = ~n17099 & n17103;
  assign n17105 = ~n17102 & n17104;
  assign n17106 = pi50  & n17105;
  assign n17107 = ~pi50  & ~n17105;
  assign n17108 = ~n17106 & ~n17107;
  assign n17109 = n17098 & ~n17108;
  assign n17110 = ~n17098 & n17108;
  assign n17111 = ~n17109 & ~n17110;
  assign n17112 = ~n17021 & n17111;
  assign n17113 = n17021 & ~n17111;
  assign n17114 = ~n17112 & ~n17113;
  assign n17115 = ~n17020 & n17114;
  assign n17116 = n17020 & ~n17114;
  assign n17117 = ~n17115 & ~n17116;
  assign n17118 = n17010 & ~n17117;
  assign n17119 = ~n17010 & n17117;
  assign n17120 = ~n17118 & ~n17119;
  assign n17121 = pi97  & n6331;
  assign n17122 = pi98  & n6015;
  assign n17123 = pi99  & n6010;
  assign n17124 = n4101 & n6008;
  assign n17125 = ~n17122 & ~n17123;
  assign n17126 = ~n17121 & n17125;
  assign n17127 = ~n17124 & n17126;
  assign n17128 = pi44  & n17127;
  assign n17129 = ~pi44  & ~n17127;
  assign n17130 = ~n17128 & ~n17129;
  assign n17131 = n17120 & ~n17130;
  assign n17132 = ~n17120 & n17130;
  assign n17133 = ~n17131 & ~n17132;
  assign n17134 = n17009 & ~n17133;
  assign n17135 = ~n17009 & n17133;
  assign n17136 = ~n17134 & ~n17135;
  assign n17137 = pi100  & n5558;
  assign n17138 = pi101  & n5293;
  assign n17139 = pi102  & n5288;
  assign n17140 = n4956 & n5286;
  assign n17141 = ~n17138 & ~n17139;
  assign n17142 = ~n17137 & n17141;
  assign n17143 = ~n17140 & n17142;
  assign n17144 = pi41  & n17143;
  assign n17145 = ~pi41  & ~n17143;
  assign n17146 = ~n17144 & ~n17145;
  assign n17147 = ~n17136 & n17146;
  assign n17148 = n17136 & ~n17146;
  assign n17149 = ~n17147 & ~n17148;
  assign n17150 = ~n17008 & n17149;
  assign n17151 = n17008 & ~n17149;
  assign n17152 = ~n17150 & ~n17151;
  assign n17153 = ~n17007 & n17152;
  assign n17154 = n17007 & ~n17152;
  assign n17155 = ~n17153 & ~n17154;
  assign n17156 = ~n16997 & n17155;
  assign n17157 = n16997 & ~n17155;
  assign n17158 = ~n17156 & ~n17157;
  assign n17159 = n16996 & ~n17158;
  assign n17160 = ~n16996 & n17158;
  assign n17161 = ~n17159 & ~n17160;
  assign n17162 = n16986 & n17161;
  assign n17163 = ~n16986 & ~n17161;
  assign n17164 = ~n17162 & ~n17163;
  assign n17165 = n16971 & n17164;
  assign n17166 = ~n16971 & ~n17164;
  assign n17167 = ~n17165 & ~n17166;
  assign n17168 = n16957 & ~n17167;
  assign n17169 = ~n16957 & n17167;
  assign n17170 = ~n17168 & ~n17169;
  assign n17171 = n16943 & ~n17170;
  assign n17172 = ~n16943 & n17170;
  assign n17173 = ~n17171 & ~n17172;
  assign n17174 = n16928 & n17173;
  assign n17175 = ~n16928 & ~n17173;
  assign n17176 = ~n17174 & ~n17175;
  assign n17177 = ~n16883 & ~n16886;
  assign n17178 = pi124  & n1296;
  assign n17179 = pi125  & n1207;
  assign n17180 = pi126  & n1202;
  assign n17181 = n1200 & n12148;
  assign n17182 = ~n17179 & ~n17180;
  assign n17183 = ~n17178 & n17182;
  assign n17184 = ~n17181 & n17183;
  assign n17185 = pi17  & n17184;
  assign n17186 = ~pi17  & ~n17184;
  assign n17187 = ~n17185 & ~n17186;
  assign n17188 = ~n17177 & ~n17187;
  assign n17189 = n17177 & n17187;
  assign n17190 = ~n17188 & ~n17189;
  assign n17191 = n17176 & n17190;
  assign n17192 = ~n17176 & ~n17190;
  assign n17193 = ~n17191 & ~n17192;
  assign n17194 = ~n16627 & ~n16889;
  assign n17195 = n890 & ~n12539;
  assign n17196 = ~n1006 & ~n17195;
  assign n17197 = pi127  & ~n17196;
  assign n17198 = pi14  & ~n17197;
  assign n17199 = ~pi14  & n17197;
  assign n17200 = ~n17198 & ~n17199;
  assign n17201 = ~n17194 & ~n17200;
  assign n17202 = n17194 & n17200;
  assign n17203 = ~n17201 & ~n17202;
  assign n17204 = n17193 & n17203;
  assign n17205 = ~n17193 & ~n17203;
  assign n17206 = ~n17204 & ~n17205;
  assign n17207 = ~n16914 & n17206;
  assign n17208 = n16914 & ~n17206;
  assign n17209 = ~n17207 & ~n17208;
  assign n17210 = ~n16913 & n17209;
  assign n17211 = n16913 & ~n17209;
  assign po77  = ~n17210 & ~n17211;
  assign n17213 = ~n17201 & ~n17204;
  assign n17214 = pi122  & n1661;
  assign n17215 = pi123  & n1500;
  assign n17216 = pi124  & n1495;
  assign n17217 = n1493 & n11099;
  assign n17218 = ~n17215 & ~n17216;
  assign n17219 = ~n17214 & n17218;
  assign n17220 = ~n17217 & n17219;
  assign n17221 = pi20  & n17220;
  assign n17222 = ~pi20  & ~n17220;
  assign n17223 = ~n17221 & ~n17222;
  assign n17224 = ~n16927 & ~n17174;
  assign n17225 = n17223 & n17224;
  assign n17226 = ~n17223 & ~n17224;
  assign n17227 = ~n17225 & ~n17226;
  assign n17228 = ~n16942 & ~n17171;
  assign n17229 = pi119  & n2053;
  assign n17230 = pi120  & n1893;
  assign n17231 = pi121  & n1888;
  assign n17232 = n1886 & n10071;
  assign n17233 = ~n17230 & ~n17231;
  assign n17234 = ~n17229 & n17233;
  assign n17235 = ~n17232 & n17234;
  assign n17236 = pi23  & n17235;
  assign n17237 = ~pi23  & ~n17235;
  assign n17238 = ~n17236 & ~n17237;
  assign n17239 = ~n17228 & ~n17238;
  assign n17240 = n17228 & n17238;
  assign n17241 = ~n17239 & ~n17240;
  assign n17242 = pi116  & n2510;
  assign n17243 = pi117  & n2342;
  assign n17244 = pi118  & n2337;
  assign n17245 = n2335 & n9095;
  assign n17246 = ~n17243 & ~n17244;
  assign n17247 = ~n17242 & n17246;
  assign n17248 = ~n17245 & n17247;
  assign n17249 = pi26  & n17248;
  assign n17250 = ~pi26  & ~n17248;
  assign n17251 = ~n17249 & ~n17250;
  assign n17252 = ~n16956 & ~n17167;
  assign n17253 = ~n16955 & ~n17252;
  assign n17254 = n17251 & ~n17253;
  assign n17255 = ~n17251 & n17253;
  assign n17256 = ~n17254 & ~n17255;
  assign n17257 = pi113  & n3011;
  assign n17258 = pi114  & n2809;
  assign n17259 = pi115  & n2804;
  assign n17260 = n2802 & n8170;
  assign n17261 = ~n17258 & ~n17259;
  assign n17262 = ~n17257 & n17261;
  assign n17263 = ~n17260 & n17262;
  assign n17264 = pi29  & n17263;
  assign n17265 = ~pi29  & ~n17263;
  assign n17266 = ~n17264 & ~n17265;
  assign n17267 = ~n16969 & ~n17164;
  assign n17268 = ~n16970 & ~n17267;
  assign n17269 = n17266 & ~n17268;
  assign n17270 = ~n17266 & n17268;
  assign n17271 = ~n17269 & ~n17270;
  assign n17272 = ~n17150 & ~n17153;
  assign n17273 = pi104  & n4843;
  assign n17274 = pi105  & n4598;
  assign n17275 = pi106  & n4593;
  assign n17276 = n4591 & n5701;
  assign n17277 = ~n17274 & ~n17275;
  assign n17278 = ~n17273 & n17277;
  assign n17279 = ~n17276 & n17278;
  assign n17280 = pi38  & n17279;
  assign n17281 = ~pi38  & ~n17279;
  assign n17282 = ~n17280 & ~n17281;
  assign n17283 = ~n17135 & ~n17148;
  assign n17284 = pi98  & n6331;
  assign n17285 = pi99  & n6015;
  assign n17286 = pi100  & n6010;
  assign n17287 = n4501 & n6008;
  assign n17288 = ~n17285 & ~n17286;
  assign n17289 = ~n17284 & n17288;
  assign n17290 = ~n17287 & n17289;
  assign n17291 = pi44  & n17290;
  assign n17292 = ~pi44  & ~n17290;
  assign n17293 = ~n17291 & ~n17292;
  assign n17294 = ~n17112 & ~n17115;
  assign n17295 = ~n17088 & ~n17091;
  assign n17296 = pi89  & n8905;
  assign n17297 = pi90  & n8535;
  assign n17298 = pi91  & n8530;
  assign n17299 = n2746 & n8528;
  assign n17300 = ~n17297 & ~n17298;
  assign n17301 = ~n17296 & n17300;
  assign n17302 = ~n17299 & n17301;
  assign n17303 = pi53  & n17302;
  assign n17304 = ~pi53  & ~n17302;
  assign n17305 = ~n17303 & ~n17304;
  assign n17306 = ~n17071 & ~n17084;
  assign n17307 = ~n17036 & ~n17049;
  assign n17308 = pi80  & n11910;
  assign n17309 = pi81  & n11529;
  assign n17310 = pi82  & n11524;
  assign n17311 = n1450 & n11522;
  assign n17312 = ~n17309 & ~n17310;
  assign n17313 = ~n17308 & n17312;
  assign n17314 = ~n17311 & n17313;
  assign n17315 = pi62  & n17314;
  assign n17316 = ~pi62  & ~n17314;
  assign n17317 = ~n17315 & ~n17316;
  assign n17318 = pi79  & n12277;
  assign n17319 = pi78  & n12276;
  assign n17320 = ~n17318 & ~n17319;
  assign n17321 = ~pi14  & ~n17320;
  assign n17322 = pi14  & n17320;
  assign n17323 = ~n17321 & ~n17322;
  assign n17324 = ~n16719 & n17323;
  assign n17325 = n16719 & ~n17323;
  assign n17326 = ~n17324 & ~n17325;
  assign n17327 = ~n17317 & n17326;
  assign n17328 = n17317 & ~n17326;
  assign n17329 = ~n17327 & ~n17328;
  assign n17330 = n17307 & ~n17329;
  assign n17331 = ~n17307 & n17329;
  assign n17332 = ~n17330 & ~n17331;
  assign n17333 = pi83  & n10886;
  assign n17334 = pi84  & n10495;
  assign n17335 = pi85  & n10490;
  assign n17336 = n1831 & n10488;
  assign n17337 = ~n17334 & ~n17335;
  assign n17338 = ~n17333 & n17337;
  assign n17339 = ~n17336 & n17338;
  assign n17340 = pi59  & n17339;
  assign n17341 = ~pi59  & ~n17339;
  assign n17342 = ~n17340 & ~n17341;
  assign n17343 = n17332 & ~n17342;
  assign n17344 = ~n17332 & n17342;
  assign n17345 = ~n17343 & ~n17344;
  assign n17346 = ~n17052 & n17064;
  assign n17347 = ~n17053 & ~n17346;
  assign n17348 = ~n17345 & ~n17347;
  assign n17349 = n17345 & n17347;
  assign n17350 = ~n17348 & ~n17349;
  assign n17351 = pi86  & n9858;
  assign n17352 = pi87  & n9508;
  assign n17353 = pi88  & n9503;
  assign n17354 = n2140 & n9501;
  assign n17355 = ~n17352 & ~n17353;
  assign n17356 = ~n17351 & n17355;
  assign n17357 = ~n17354 & n17356;
  assign n17358 = pi56  & n17357;
  assign n17359 = ~pi56  & ~n17357;
  assign n17360 = ~n17358 & ~n17359;
  assign n17361 = n17350 & ~n17360;
  assign n17362 = ~n17350 & n17360;
  assign n17363 = ~n17361 & ~n17362;
  assign n17364 = n17306 & n17363;
  assign n17365 = ~n17306 & ~n17363;
  assign n17366 = ~n17364 & ~n17365;
  assign n17367 = ~n17305 & ~n17366;
  assign n17368 = n17305 & n17366;
  assign n17369 = ~n17367 & ~n17368;
  assign n17370 = n17295 & ~n17369;
  assign n17371 = ~n17295 & n17369;
  assign n17372 = ~n17370 & ~n17371;
  assign n17373 = pi92  & n7969;
  assign n17374 = pi93  & n7636;
  assign n17375 = pi94  & n7631;
  assign n17376 = n3280 & n7629;
  assign n17377 = ~n17374 & ~n17375;
  assign n17378 = ~n17373 & n17377;
  assign n17379 = ~n17376 & n17378;
  assign n17380 = pi50  & n17379;
  assign n17381 = ~pi50  & ~n17379;
  assign n17382 = ~n17380 & ~n17381;
  assign n17383 = n17372 & ~n17382;
  assign n17384 = ~n17372 & n17382;
  assign n17385 = ~n17383 & ~n17384;
  assign n17386 = ~n17096 & n17108;
  assign n17387 = ~n17097 & ~n17386;
  assign n17388 = ~n17385 & ~n17387;
  assign n17389 = n17385 & n17387;
  assign n17390 = ~n17388 & ~n17389;
  assign n17391 = pi95  & n7121;
  assign n17392 = pi96  & n6795;
  assign n17393 = pi97  & n6790;
  assign n17394 = n3691 & n6788;
  assign n17395 = ~n17392 & ~n17393;
  assign n17396 = ~n17391 & n17395;
  assign n17397 = ~n17394 & n17396;
  assign n17398 = pi47  & n17397;
  assign n17399 = ~pi47  & ~n17397;
  assign n17400 = ~n17398 & ~n17399;
  assign n17401 = n17390 & ~n17400;
  assign n17402 = ~n17390 & n17400;
  assign n17403 = ~n17401 & ~n17402;
  assign n17404 = ~n17294 & n17403;
  assign n17405 = n17294 & ~n17403;
  assign n17406 = ~n17404 & ~n17405;
  assign n17407 = ~n17293 & n17406;
  assign n17408 = n17293 & ~n17406;
  assign n17409 = ~n17407 & ~n17408;
  assign n17410 = ~n17119 & n17130;
  assign n17411 = ~n17118 & ~n17410;
  assign n17412 = ~n17409 & ~n17411;
  assign n17413 = n17409 & n17411;
  assign n17414 = ~n17412 & ~n17413;
  assign n17415 = pi101  & n5558;
  assign n17416 = pi102  & n5293;
  assign n17417 = pi103  & n5288;
  assign n17418 = n5188 & n5286;
  assign n17419 = ~n17416 & ~n17417;
  assign n17420 = ~n17415 & n17419;
  assign n17421 = ~n17418 & n17420;
  assign n17422 = pi41  & n17421;
  assign n17423 = ~pi41  & ~n17421;
  assign n17424 = ~n17422 & ~n17423;
  assign n17425 = n17414 & ~n17424;
  assign n17426 = ~n17414 & n17424;
  assign n17427 = ~n17425 & ~n17426;
  assign n17428 = ~n17283 & n17427;
  assign n17429 = n17283 & ~n17427;
  assign n17430 = ~n17428 & ~n17429;
  assign n17431 = ~n17282 & n17430;
  assign n17432 = n17282 & ~n17430;
  assign n17433 = ~n17431 & ~n17432;
  assign n17434 = n17272 & ~n17433;
  assign n17435 = ~n17272 & n17433;
  assign n17436 = ~n17434 & ~n17435;
  assign n17437 = pi107  & n4176;
  assign n17438 = pi108  & n3938;
  assign n17439 = pi109  & n3933;
  assign n17440 = n3931 & n6715;
  assign n17441 = ~n17438 & ~n17439;
  assign n17442 = ~n17437 & n17441;
  assign n17443 = ~n17440 & n17442;
  assign n17444 = pi35  & n17443;
  assign n17445 = ~pi35  & ~n17443;
  assign n17446 = ~n17444 & ~n17445;
  assign n17447 = n17436 & ~n17446;
  assign n17448 = ~n17436 & n17446;
  assign n17449 = ~n17447 & ~n17448;
  assign n17450 = n16996 & ~n17156;
  assign n17451 = ~n17157 & ~n17450;
  assign n17452 = ~n17449 & ~n17451;
  assign n17453 = n17449 & n17451;
  assign n17454 = ~n17452 & ~n17453;
  assign n17455 = pi110  & n3553;
  assign n17456 = pi111  & n3334;
  assign n17457 = pi112  & n3329;
  assign n17458 = n3327 & n7296;
  assign n17459 = ~n17456 & ~n17457;
  assign n17460 = ~n17455 & n17459;
  assign n17461 = ~n17458 & n17460;
  assign n17462 = pi32  & n17461;
  assign n17463 = ~pi32  & ~n17461;
  assign n17464 = ~n17462 & ~n17463;
  assign n17465 = ~n16984 & ~n17161;
  assign n17466 = ~n16985 & ~n17465;
  assign n17467 = ~n17464 & n17466;
  assign n17468 = n17464 & ~n17466;
  assign n17469 = ~n17467 & ~n17468;
  assign n17470 = n17454 & n17469;
  assign n17471 = ~n17454 & ~n17469;
  assign n17472 = ~n17470 & ~n17471;
  assign n17473 = n17271 & n17472;
  assign n17474 = ~n17271 & ~n17472;
  assign n17475 = ~n17473 & ~n17474;
  assign n17476 = n17256 & n17475;
  assign n17477 = ~n17256 & ~n17475;
  assign n17478 = ~n17476 & ~n17477;
  assign n17479 = n17241 & n17478;
  assign n17480 = ~n17241 & ~n17478;
  assign n17481 = ~n17479 & ~n17480;
  assign n17482 = n17227 & n17481;
  assign n17483 = ~n17227 & ~n17481;
  assign n17484 = ~n17482 & ~n17483;
  assign n17485 = ~n17188 & ~n17191;
  assign n17486 = pi125  & n1296;
  assign n17487 = pi126  & n1207;
  assign n17488 = pi127  & n1202;
  assign n17489 = n1200 & n12519;
  assign n17490 = ~n17487 & ~n17488;
  assign n17491 = ~n17486 & n17490;
  assign n17492 = ~n17489 & n17491;
  assign n17493 = pi17  & n17492;
  assign n17494 = ~pi17  & ~n17492;
  assign n17495 = ~n17493 & ~n17494;
  assign n17496 = ~n17485 & ~n17495;
  assign n17497 = n17485 & n17495;
  assign n17498 = ~n17496 & ~n17497;
  assign n17499 = n17484 & n17498;
  assign n17500 = ~n17484 & ~n17498;
  assign n17501 = ~n17499 & ~n17500;
  assign n17502 = n17213 & ~n17501;
  assign n17503 = ~n17213 & n17501;
  assign n17504 = ~n17502 & ~n17503;
  assign n17505 = ~n17207 & ~n17210;
  assign n17506 = n17504 & ~n17505;
  assign n17507 = ~n17504 & n17505;
  assign po78  = ~n17506 & ~n17507;
  assign n17509 = ~n17496 & ~n17499;
  assign n17510 = ~n17226 & ~n17482;
  assign n17511 = pi126  & n1296;
  assign n17512 = pi127  & n1207;
  assign n17513 = n1200 & n12542;
  assign n17514 = ~n17511 & ~n17512;
  assign n17515 = ~n17513 & n17514;
  assign n17516 = pi17  & n17515;
  assign n17517 = ~pi17  & ~n17515;
  assign n17518 = ~n17516 & ~n17517;
  assign n17519 = ~n17510 & ~n17518;
  assign n17520 = n17510 & n17518;
  assign n17521 = ~n17519 & ~n17520;
  assign n17522 = pi123  & n1661;
  assign n17523 = pi124  & n1500;
  assign n17524 = pi125  & n1495;
  assign n17525 = n1493 & n11786;
  assign n17526 = ~n17523 & ~n17524;
  assign n17527 = ~n17522 & n17526;
  assign n17528 = ~n17525 & n17527;
  assign n17529 = pi20  & n17528;
  assign n17530 = ~pi20  & ~n17528;
  assign n17531 = ~n17529 & ~n17530;
  assign n17532 = ~n17239 & ~n17478;
  assign n17533 = ~n17240 & ~n17532;
  assign n17534 = n17531 & ~n17533;
  assign n17535 = ~n17531 & n17533;
  assign n17536 = ~n17534 & ~n17535;
  assign n17537 = ~n17255 & ~n17476;
  assign n17538 = pi120  & n2053;
  assign n17539 = pi121  & n1893;
  assign n17540 = pi122  & n1888;
  assign n17541 = n1886 & n10729;
  assign n17542 = ~n17539 & ~n17540;
  assign n17543 = ~n17538 & n17542;
  assign n17544 = ~n17541 & n17543;
  assign n17545 = pi23  & n17544;
  assign n17546 = ~pi23  & ~n17544;
  assign n17547 = ~n17545 & ~n17546;
  assign n17548 = ~n17537 & ~n17547;
  assign n17549 = n17537 & n17547;
  assign n17550 = ~n17548 & ~n17549;
  assign n17551 = pi117  & n2510;
  assign n17552 = pi118  & n2342;
  assign n17553 = pi119  & n2337;
  assign n17554 = n2335 & n9412;
  assign n17555 = ~n17552 & ~n17553;
  assign n17556 = ~n17551 & n17555;
  assign n17557 = ~n17554 & n17556;
  assign n17558 = pi26  & n17557;
  assign n17559 = ~pi26  & ~n17557;
  assign n17560 = ~n17558 & ~n17559;
  assign n17561 = ~n17270 & ~n17473;
  assign n17562 = n17560 & n17561;
  assign n17563 = ~n17560 & ~n17561;
  assign n17564 = ~n17562 & ~n17563;
  assign n17565 = pi111  & n3553;
  assign n17566 = pi112  & n3334;
  assign n17567 = pi113  & n3329;
  assign n17568 = n3327 & n7852;
  assign n17569 = ~n17566 & ~n17567;
  assign n17570 = ~n17565 & n17569;
  assign n17571 = ~n17568 & n17570;
  assign n17572 = pi32  & n17571;
  assign n17573 = ~pi32  & ~n17571;
  assign n17574 = ~n17572 & ~n17573;
  assign n17575 = ~n17447 & ~n17453;
  assign n17576 = n17574 & n17575;
  assign n17577 = ~n17574 & ~n17575;
  assign n17578 = ~n17576 & ~n17577;
  assign n17579 = ~n17431 & ~n17435;
  assign n17580 = ~n17425 & ~n17428;
  assign n17581 = pi102  & n5558;
  assign n17582 = pi103  & n5293;
  assign n17583 = pi104  & n5288;
  assign n17584 = n5212 & n5286;
  assign n17585 = ~n17582 & ~n17583;
  assign n17586 = ~n17581 & n17585;
  assign n17587 = ~n17584 & n17586;
  assign n17588 = pi41  & n17587;
  assign n17589 = ~pi41  & ~n17587;
  assign n17590 = ~n17588 & ~n17589;
  assign n17591 = ~n17407 & ~n17413;
  assign n17592 = pi99  & n6331;
  assign n17593 = pi100  & n6015;
  assign n17594 = pi101  & n6010;
  assign n17595 = n4730 & n6008;
  assign n17596 = ~n17593 & ~n17594;
  assign n17597 = ~n17592 & n17596;
  assign n17598 = ~n17595 & n17597;
  assign n17599 = pi44  & n17598;
  assign n17600 = ~pi44  & ~n17598;
  assign n17601 = ~n17599 & ~n17600;
  assign n17602 = ~n17401 & ~n17404;
  assign n17603 = ~n17383 & ~n17389;
  assign n17604 = pi90  & n8905;
  assign n17605 = pi91  & n8535;
  assign n17606 = pi92  & n8530;
  assign n17607 = n2924 & n8528;
  assign n17608 = ~n17605 & ~n17606;
  assign n17609 = ~n17604 & n17608;
  assign n17610 = ~n17607 & n17609;
  assign n17611 = pi53  & n17610;
  assign n17612 = ~pi53  & ~n17610;
  assign n17613 = ~n17611 & ~n17612;
  assign n17614 = ~n17343 & ~n17349;
  assign n17615 = ~n17327 & ~n17331;
  assign n17616 = ~n17321 & ~n17324;
  assign n17617 = pi80  & n12277;
  assign n17618 = pi79  & n12276;
  assign n17619 = ~n17617 & ~n17618;
  assign n17620 = n17616 & ~n17619;
  assign n17621 = ~n17616 & n17619;
  assign n17622 = ~n17620 & ~n17621;
  assign n17623 = pi81  & n11910;
  assign n17624 = pi82  & n11529;
  assign n17625 = pi83  & n11524;
  assign n17626 = n1577 & n11522;
  assign n17627 = ~n17624 & ~n17625;
  assign n17628 = ~n17623 & n17627;
  assign n17629 = ~n17626 & n17628;
  assign n17630 = pi62  & n17629;
  assign n17631 = ~pi62  & ~n17629;
  assign n17632 = ~n17630 & ~n17631;
  assign n17633 = n17622 & ~n17632;
  assign n17634 = ~n17622 & n17632;
  assign n17635 = ~n17633 & ~n17634;
  assign n17636 = ~n17615 & n17635;
  assign n17637 = n17615 & ~n17635;
  assign n17638 = ~n17636 & ~n17637;
  assign n17639 = pi84  & n10886;
  assign n17640 = pi85  & n10495;
  assign n17641 = pi86  & n10490;
  assign n17642 = n1975 & n10488;
  assign n17643 = ~n17640 & ~n17641;
  assign n17644 = ~n17639 & n17643;
  assign n17645 = ~n17642 & n17644;
  assign n17646 = pi59  & n17645;
  assign n17647 = ~pi59  & ~n17645;
  assign n17648 = ~n17646 & ~n17647;
  assign n17649 = n17638 & ~n17648;
  assign n17650 = ~n17638 & n17648;
  assign n17651 = ~n17649 & ~n17650;
  assign n17652 = n17614 & ~n17651;
  assign n17653 = ~n17614 & n17651;
  assign n17654 = ~n17652 & ~n17653;
  assign n17655 = pi87  & n9858;
  assign n17656 = pi88  & n9508;
  assign n17657 = pi89  & n9503;
  assign n17658 = n2287 & n9501;
  assign n17659 = ~n17656 & ~n17657;
  assign n17660 = ~n17655 & n17659;
  assign n17661 = ~n17658 & n17660;
  assign n17662 = pi56  & n17661;
  assign n17663 = ~pi56  & ~n17661;
  assign n17664 = ~n17662 & ~n17663;
  assign n17665 = n17654 & ~n17664;
  assign n17666 = ~n17654 & n17664;
  assign n17667 = ~n17665 & ~n17666;
  assign n17668 = n17306 & ~n17361;
  assign n17669 = ~n17362 & ~n17668;
  assign n17670 = n17667 & n17669;
  assign n17671 = ~n17667 & ~n17669;
  assign n17672 = ~n17670 & ~n17671;
  assign n17673 = n17613 & ~n17672;
  assign n17674 = ~n17613 & n17672;
  assign n17675 = ~n17673 & ~n17674;
  assign n17676 = ~n17367 & ~n17371;
  assign n17677 = n17675 & ~n17676;
  assign n17678 = ~n17675 & n17676;
  assign n17679 = ~n17677 & ~n17678;
  assign n17680 = pi93  & n7969;
  assign n17681 = pi94  & n7636;
  assign n17682 = pi95  & n7631;
  assign n17683 = n3475 & n7629;
  assign n17684 = ~n17681 & ~n17682;
  assign n17685 = ~n17680 & n17684;
  assign n17686 = ~n17683 & n17685;
  assign n17687 = pi50  & n17686;
  assign n17688 = ~pi50  & ~n17686;
  assign n17689 = ~n17687 & ~n17688;
  assign n17690 = n17679 & ~n17689;
  assign n17691 = ~n17679 & n17689;
  assign n17692 = ~n17690 & ~n17691;
  assign n17693 = n17603 & ~n17692;
  assign n17694 = ~n17603 & n17692;
  assign n17695 = ~n17693 & ~n17694;
  assign n17696 = pi96  & n7121;
  assign n17697 = pi97  & n6795;
  assign n17698 = pi98  & n6790;
  assign n17699 = n3889 & n6788;
  assign n17700 = ~n17697 & ~n17698;
  assign n17701 = ~n17696 & n17700;
  assign n17702 = ~n17699 & n17701;
  assign n17703 = pi47  & n17702;
  assign n17704 = ~pi47  & ~n17702;
  assign n17705 = ~n17703 & ~n17704;
  assign n17706 = ~n17695 & n17705;
  assign n17707 = n17695 & ~n17705;
  assign n17708 = ~n17706 & ~n17707;
  assign n17709 = ~n17602 & n17708;
  assign n17710 = n17602 & ~n17708;
  assign n17711 = ~n17709 & ~n17710;
  assign n17712 = ~n17601 & n17711;
  assign n17713 = n17601 & ~n17711;
  assign n17714 = ~n17712 & ~n17713;
  assign n17715 = ~n17591 & n17714;
  assign n17716 = n17591 & ~n17714;
  assign n17717 = ~n17715 & ~n17716;
  assign n17718 = ~n17590 & n17717;
  assign n17719 = n17590 & ~n17717;
  assign n17720 = ~n17718 & ~n17719;
  assign n17721 = ~n17580 & n17720;
  assign n17722 = n17580 & ~n17720;
  assign n17723 = ~n17721 & ~n17722;
  assign n17724 = pi105  & n4843;
  assign n17725 = pi106  & n4598;
  assign n17726 = pi107  & n4593;
  assign n17727 = n4591 & n6189;
  assign n17728 = ~n17725 & ~n17726;
  assign n17729 = ~n17724 & n17728;
  assign n17730 = ~n17727 & n17729;
  assign n17731 = pi38  & n17730;
  assign n17732 = ~pi38  & ~n17730;
  assign n17733 = ~n17731 & ~n17732;
  assign n17734 = n17723 & ~n17733;
  assign n17735 = ~n17723 & n17733;
  assign n17736 = ~n17734 & ~n17735;
  assign n17737 = n17579 & ~n17736;
  assign n17738 = ~n17579 & n17736;
  assign n17739 = ~n17737 & ~n17738;
  assign n17740 = pi108  & n4176;
  assign n17741 = pi109  & n3938;
  assign n17742 = pi110  & n3933;
  assign n17743 = n3931 & n6995;
  assign n17744 = ~n17741 & ~n17742;
  assign n17745 = ~n17740 & n17744;
  assign n17746 = ~n17743 & n17745;
  assign n17747 = pi35  & n17746;
  assign n17748 = ~pi35  & ~n17746;
  assign n17749 = ~n17747 & ~n17748;
  assign n17750 = n17739 & ~n17749;
  assign n17751 = ~n17739 & n17749;
  assign n17752 = ~n17750 & ~n17751;
  assign n17753 = n17578 & n17752;
  assign n17754 = ~n17578 & ~n17752;
  assign n17755 = ~n17753 & ~n17754;
  assign n17756 = pi114  & n3011;
  assign n17757 = pi115  & n2809;
  assign n17758 = pi116  & n2804;
  assign n17759 = n2802 & n8470;
  assign n17760 = ~n17757 & ~n17758;
  assign n17761 = ~n17756 & n17760;
  assign n17762 = ~n17759 & n17761;
  assign n17763 = pi29  & n17762;
  assign n17764 = ~pi29  & ~n17762;
  assign n17765 = ~n17763 & ~n17764;
  assign n17766 = ~n17467 & ~n17470;
  assign n17767 = ~n17765 & ~n17766;
  assign n17768 = n17765 & n17766;
  assign n17769 = ~n17767 & ~n17768;
  assign n17770 = n17755 & n17769;
  assign n17771 = ~n17755 & ~n17769;
  assign n17772 = ~n17770 & ~n17771;
  assign n17773 = n17564 & n17772;
  assign n17774 = ~n17564 & ~n17772;
  assign n17775 = ~n17773 & ~n17774;
  assign n17776 = n17550 & n17775;
  assign n17777 = ~n17550 & ~n17775;
  assign n17778 = ~n17776 & ~n17777;
  assign n17779 = n17536 & n17778;
  assign n17780 = ~n17536 & ~n17778;
  assign n17781 = ~n17779 & ~n17780;
  assign n17782 = n17521 & n17781;
  assign n17783 = ~n17521 & ~n17781;
  assign n17784 = ~n17782 & ~n17783;
  assign n17785 = n17509 & ~n17784;
  assign n17786 = ~n17509 & n17784;
  assign n17787 = ~n17785 & ~n17786;
  assign n17788 = ~n17503 & ~n17506;
  assign n17789 = n17787 & ~n17788;
  assign n17790 = ~n17787 & n17788;
  assign po79  = ~n17789 & ~n17790;
  assign n17792 = ~n17786 & ~n17789;
  assign n17793 = pi124  & n1661;
  assign n17794 = pi125  & n1500;
  assign n17795 = pi126  & n1495;
  assign n17796 = n1493 & n12148;
  assign n17797 = ~n17794 & ~n17795;
  assign n17798 = ~n17793 & n17797;
  assign n17799 = ~n17796 & n17798;
  assign n17800 = pi20  & n17799;
  assign n17801 = ~pi20  & ~n17799;
  assign n17802 = ~n17800 & ~n17801;
  assign n17803 = ~n17548 & ~n17776;
  assign n17804 = n17802 & n17803;
  assign n17805 = ~n17802 & ~n17803;
  assign n17806 = ~n17804 & ~n17805;
  assign n17807 = pi118  & n2510;
  assign n17808 = pi119  & n2342;
  assign n17809 = pi120  & n2337;
  assign n17810 = n2335 & n10047;
  assign n17811 = ~n17808 & ~n17809;
  assign n17812 = ~n17807 & n17811;
  assign n17813 = ~n17810 & n17812;
  assign n17814 = pi26  & n17813;
  assign n17815 = ~pi26  & ~n17813;
  assign n17816 = ~n17814 & ~n17815;
  assign n17817 = ~n17767 & ~n17770;
  assign n17818 = n17816 & n17817;
  assign n17819 = ~n17816 & ~n17817;
  assign n17820 = ~n17818 & ~n17819;
  assign n17821 = pi112  & n3553;
  assign n17822 = pi113  & n3334;
  assign n17823 = pi114  & n3329;
  assign n17824 = n3327 & n8146;
  assign n17825 = ~n17822 & ~n17823;
  assign n17826 = ~n17821 & n17825;
  assign n17827 = ~n17824 & n17826;
  assign n17828 = pi32  & n17827;
  assign n17829 = ~pi32  & ~n17827;
  assign n17830 = ~n17828 & ~n17829;
  assign n17831 = ~n17738 & n17749;
  assign n17832 = ~n17737 & ~n17831;
  assign n17833 = n17830 & ~n17832;
  assign n17834 = ~n17830 & n17832;
  assign n17835 = ~n17833 & ~n17834;
  assign n17836 = pi106  & n4843;
  assign n17837 = pi107  & n4598;
  assign n17838 = pi108  & n4593;
  assign n17839 = n4591 & n6213;
  assign n17840 = ~n17837 & ~n17838;
  assign n17841 = ~n17836 & n17840;
  assign n17842 = ~n17839 & n17841;
  assign n17843 = pi38  & n17842;
  assign n17844 = ~pi38  & ~n17842;
  assign n17845 = ~n17843 & ~n17844;
  assign n17846 = ~n17715 & ~n17718;
  assign n17847 = pi103  & n5558;
  assign n17848 = pi104  & n5293;
  assign n17849 = pi105  & n5288;
  assign n17850 = n5286 & n5677;
  assign n17851 = ~n17848 & ~n17849;
  assign n17852 = ~n17847 & n17851;
  assign n17853 = ~n17850 & n17852;
  assign n17854 = pi41  & n17853;
  assign n17855 = ~pi41  & ~n17853;
  assign n17856 = ~n17854 & ~n17855;
  assign n17857 = ~n17709 & ~n17712;
  assign n17858 = pi100  & n6331;
  assign n17859 = pi101  & n6015;
  assign n17860 = pi102  & n6010;
  assign n17861 = n4956 & n6008;
  assign n17862 = ~n17859 & ~n17860;
  assign n17863 = ~n17858 & n17862;
  assign n17864 = ~n17861 & n17863;
  assign n17865 = pi44  & n17864;
  assign n17866 = ~pi44  & ~n17864;
  assign n17867 = ~n17865 & ~n17866;
  assign n17868 = ~n17694 & ~n17707;
  assign n17869 = pi94  & n7969;
  assign n17870 = pi95  & n7636;
  assign n17871 = pi96  & n7631;
  assign n17872 = n3499 & n7629;
  assign n17873 = ~n17870 & ~n17871;
  assign n17874 = ~n17869 & n17873;
  assign n17875 = ~n17872 & n17874;
  assign n17876 = pi50  & n17875;
  assign n17877 = ~pi50  & ~n17875;
  assign n17878 = ~n17876 & ~n17877;
  assign n17879 = ~n17670 & ~n17674;
  assign n17880 = pi88  & n9858;
  assign n17881 = pi89  & n9508;
  assign n17882 = pi90  & n9503;
  assign n17883 = n2448 & n9501;
  assign n17884 = ~n17881 & ~n17882;
  assign n17885 = ~n17880 & n17884;
  assign n17886 = ~n17883 & n17885;
  assign n17887 = pi56  & n17886;
  assign n17888 = ~pi56  & ~n17886;
  assign n17889 = ~n17887 & ~n17888;
  assign n17890 = ~n17621 & ~n17633;
  assign n17891 = pi82  & n11910;
  assign n17892 = pi83  & n11529;
  assign n17893 = pi84  & n11524;
  assign n17894 = n1601 & n11522;
  assign n17895 = ~n17892 & ~n17893;
  assign n17896 = ~n17891 & n17895;
  assign n17897 = ~n17894 & n17896;
  assign n17898 = pi62  & n17897;
  assign n17899 = ~pi62  & ~n17897;
  assign n17900 = ~n17898 & ~n17899;
  assign n17901 = pi81  & n12277;
  assign n17902 = pi80  & n12276;
  assign n17903 = ~n17901 & ~n17902;
  assign n17904 = n17619 & ~n17903;
  assign n17905 = ~n17619 & n17903;
  assign n17906 = ~n17904 & ~n17905;
  assign n17907 = ~n17900 & n17906;
  assign n17908 = n17900 & ~n17906;
  assign n17909 = ~n17907 & ~n17908;
  assign n17910 = n17890 & ~n17909;
  assign n17911 = ~n17890 & n17909;
  assign n17912 = ~n17910 & ~n17911;
  assign n17913 = pi85  & n10886;
  assign n17914 = pi86  & n10495;
  assign n17915 = pi87  & n10490;
  assign n17916 = n2116 & n10488;
  assign n17917 = ~n17914 & ~n17915;
  assign n17918 = ~n17913 & n17917;
  assign n17919 = ~n17916 & n17918;
  assign n17920 = pi59  & n17919;
  assign n17921 = ~pi59  & ~n17919;
  assign n17922 = ~n17920 & ~n17921;
  assign n17923 = ~n17912 & n17922;
  assign n17924 = n17912 & ~n17922;
  assign n17925 = ~n17923 & ~n17924;
  assign n17926 = ~n17636 & n17648;
  assign n17927 = ~n17637 & ~n17926;
  assign n17928 = n17925 & n17927;
  assign n17929 = ~n17925 & ~n17927;
  assign n17930 = ~n17928 & ~n17929;
  assign n17931 = ~n17889 & n17930;
  assign n17932 = n17889 & ~n17930;
  assign n17933 = ~n17931 & ~n17932;
  assign n17934 = ~n17653 & n17664;
  assign n17935 = ~n17652 & ~n17934;
  assign n17936 = n17933 & n17935;
  assign n17937 = ~n17933 & ~n17935;
  assign n17938 = ~n17936 & ~n17937;
  assign n17939 = pi91  & n8905;
  assign n17940 = pi92  & n8535;
  assign n17941 = pi93  & n8530;
  assign n17942 = n2948 & n8528;
  assign n17943 = ~n17940 & ~n17941;
  assign n17944 = ~n17939 & n17943;
  assign n17945 = ~n17942 & n17944;
  assign n17946 = pi53  & n17945;
  assign n17947 = ~pi53  & ~n17945;
  assign n17948 = ~n17946 & ~n17947;
  assign n17949 = n17938 & ~n17948;
  assign n17950 = ~n17938 & n17948;
  assign n17951 = ~n17949 & ~n17950;
  assign n17952 = ~n17879 & n17951;
  assign n17953 = n17879 & ~n17951;
  assign n17954 = ~n17952 & ~n17953;
  assign n17955 = ~n17878 & n17954;
  assign n17956 = n17878 & ~n17954;
  assign n17957 = ~n17955 & ~n17956;
  assign n17958 = ~n17678 & ~n17689;
  assign n17959 = ~n17677 & ~n17958;
  assign n17960 = ~n17957 & n17959;
  assign n17961 = n17957 & ~n17959;
  assign n17962 = ~n17960 & ~n17961;
  assign n17963 = pi97  & n7121;
  assign n17964 = pi98  & n6795;
  assign n17965 = pi99  & n6790;
  assign n17966 = n4101 & n6788;
  assign n17967 = ~n17964 & ~n17965;
  assign n17968 = ~n17963 & n17967;
  assign n17969 = ~n17966 & n17968;
  assign n17970 = pi47  & n17969;
  assign n17971 = ~pi47  & ~n17969;
  assign n17972 = ~n17970 & ~n17971;
  assign n17973 = n17962 & ~n17972;
  assign n17974 = ~n17962 & n17972;
  assign n17975 = ~n17973 & ~n17974;
  assign n17976 = ~n17868 & n17975;
  assign n17977 = n17868 & ~n17975;
  assign n17978 = ~n17976 & ~n17977;
  assign n17979 = ~n17867 & n17978;
  assign n17980 = n17867 & ~n17978;
  assign n17981 = ~n17979 & ~n17980;
  assign n17982 = ~n17857 & n17981;
  assign n17983 = n17857 & ~n17981;
  assign n17984 = ~n17982 & ~n17983;
  assign n17985 = ~n17856 & n17984;
  assign n17986 = n17856 & ~n17984;
  assign n17987 = ~n17985 & ~n17986;
  assign n17988 = ~n17846 & n17987;
  assign n17989 = n17846 & ~n17987;
  assign n17990 = ~n17988 & ~n17989;
  assign n17991 = ~n17845 & n17990;
  assign n17992 = n17845 & ~n17990;
  assign n17993 = ~n17991 & ~n17992;
  assign n17994 = ~n17721 & n17733;
  assign n17995 = ~n17722 & ~n17994;
  assign n17996 = n17993 & n17995;
  assign n17997 = ~n17993 & ~n17995;
  assign n17998 = ~n17996 & ~n17997;
  assign n17999 = pi109  & n4176;
  assign n18000 = pi110  & n3938;
  assign n18001 = pi111  & n3933;
  assign n18002 = n3931 & n7272;
  assign n18003 = ~n18000 & ~n18001;
  assign n18004 = ~n17999 & n18003;
  assign n18005 = ~n18002 & n18004;
  assign n18006 = pi35  & n18005;
  assign n18007 = ~pi35  & ~n18005;
  assign n18008 = ~n18006 & ~n18007;
  assign n18009 = n17998 & ~n18008;
  assign n18010 = ~n17998 & n18008;
  assign n18011 = ~n18009 & ~n18010;
  assign n18012 = n17835 & n18011;
  assign n18013 = ~n17835 & ~n18011;
  assign n18014 = ~n18012 & ~n18013;
  assign n18015 = pi115  & n3011;
  assign n18016 = pi116  & n2809;
  assign n18017 = pi117  & n2804;
  assign n18018 = n2802 & n8784;
  assign n18019 = ~n18016 & ~n18017;
  assign n18020 = ~n18015 & n18019;
  assign n18021 = ~n18018 & n18020;
  assign n18022 = pi29  & n18021;
  assign n18023 = ~pi29  & ~n18021;
  assign n18024 = ~n18022 & ~n18023;
  assign n18025 = ~n17577 & ~n17753;
  assign n18026 = ~n18024 & ~n18025;
  assign n18027 = n18024 & n18025;
  assign n18028 = ~n18026 & ~n18027;
  assign n18029 = n18014 & n18028;
  assign n18030 = ~n18014 & ~n18028;
  assign n18031 = ~n18029 & ~n18030;
  assign n18032 = n17820 & n18031;
  assign n18033 = ~n17820 & ~n18031;
  assign n18034 = ~n18032 & ~n18033;
  assign n18035 = pi121  & n2053;
  assign n18036 = pi122  & n1893;
  assign n18037 = pi123  & n1888;
  assign n18038 = n1886 & n10754;
  assign n18039 = ~n18036 & ~n18037;
  assign n18040 = ~n18035 & n18039;
  assign n18041 = ~n18038 & n18040;
  assign n18042 = pi23  & n18041;
  assign n18043 = ~pi23  & ~n18041;
  assign n18044 = ~n18042 & ~n18043;
  assign n18045 = ~n17563 & ~n17773;
  assign n18046 = ~n18044 & ~n18045;
  assign n18047 = n18044 & n18045;
  assign n18048 = ~n18046 & ~n18047;
  assign n18049 = n18034 & n18048;
  assign n18050 = ~n18034 & ~n18048;
  assign n18051 = ~n18049 & ~n18050;
  assign n18052 = ~n17806 & ~n18051;
  assign n18053 = n17806 & n18051;
  assign n18054 = ~n18052 & ~n18053;
  assign n18055 = ~n17535 & ~n17779;
  assign n18056 = n1200 & ~n12539;
  assign n18057 = ~n1296 & ~n18056;
  assign n18058 = pi127  & ~n18057;
  assign n18059 = pi17  & ~n18058;
  assign n18060 = ~pi17  & n18058;
  assign n18061 = ~n18059 & ~n18060;
  assign n18062 = ~n18055 & ~n18061;
  assign n18063 = n18055 & n18061;
  assign n18064 = ~n18062 & ~n18063;
  assign n18065 = n18054 & n18064;
  assign n18066 = ~n18054 & ~n18064;
  assign n18067 = ~n18065 & ~n18066;
  assign n18068 = ~n17519 & ~n17781;
  assign n18069 = ~n17520 & ~n18068;
  assign n18070 = n18067 & n18069;
  assign n18071 = ~n18067 & ~n18069;
  assign n18072 = ~n18070 & ~n18071;
  assign n18073 = ~n17792 & n18072;
  assign n18074 = n17792 & ~n18072;
  assign po80  = ~n18073 & ~n18074;
  assign n18076 = ~n18070 & ~n18073;
  assign n18077 = ~n18062 & ~n18065;
  assign n18078 = ~n17805 & ~n18053;
  assign n18079 = pi125  & n1661;
  assign n18080 = pi126  & n1500;
  assign n18081 = pi127  & n1495;
  assign n18082 = n1493 & n12519;
  assign n18083 = ~n18080 & ~n18081;
  assign n18084 = ~n18079 & n18083;
  assign n18085 = ~n18082 & n18084;
  assign n18086 = pi20  & n18085;
  assign n18087 = ~pi20  & ~n18085;
  assign n18088 = ~n18086 & ~n18087;
  assign n18089 = ~n18078 & ~n18088;
  assign n18090 = n18078 & n18088;
  assign n18091 = ~n18089 & ~n18090;
  assign n18092 = pi122  & n2053;
  assign n18093 = pi123  & n1893;
  assign n18094 = pi124  & n1888;
  assign n18095 = n1886 & n11099;
  assign n18096 = ~n18093 & ~n18094;
  assign n18097 = ~n18092 & n18096;
  assign n18098 = ~n18095 & n18097;
  assign n18099 = pi23  & n18098;
  assign n18100 = ~pi23  & ~n18098;
  assign n18101 = ~n18099 & ~n18100;
  assign n18102 = ~n18046 & ~n18049;
  assign n18103 = n18101 & n18102;
  assign n18104 = ~n18101 & ~n18102;
  assign n18105 = ~n18103 & ~n18104;
  assign n18106 = pi116  & n3011;
  assign n18107 = pi117  & n2809;
  assign n18108 = pi118  & n2804;
  assign n18109 = n2802 & n9095;
  assign n18110 = ~n18107 & ~n18108;
  assign n18111 = ~n18106 & n18110;
  assign n18112 = ~n18109 & n18111;
  assign n18113 = pi29  & n18112;
  assign n18114 = ~pi29  & ~n18112;
  assign n18115 = ~n18113 & ~n18114;
  assign n18116 = ~n18026 & ~n18029;
  assign n18117 = n18115 & n18116;
  assign n18118 = ~n18115 & ~n18116;
  assign n18119 = ~n18117 & ~n18118;
  assign n18120 = ~n17988 & ~n17991;
  assign n18121 = ~n17982 & ~n17985;
  assign n18122 = pi104  & n5558;
  assign n18123 = pi105  & n5293;
  assign n18124 = pi106  & n5288;
  assign n18125 = n5286 & n5701;
  assign n18126 = ~n18123 & ~n18124;
  assign n18127 = ~n18122 & n18126;
  assign n18128 = ~n18125 & n18127;
  assign n18129 = pi41  & n18128;
  assign n18130 = ~pi41  & ~n18128;
  assign n18131 = ~n18129 & ~n18130;
  assign n18132 = ~n17976 & ~n17979;
  assign n18133 = pi98  & n7121;
  assign n18134 = pi99  & n6795;
  assign n18135 = pi100  & n6790;
  assign n18136 = n4501 & n6788;
  assign n18137 = ~n18134 & ~n18135;
  assign n18138 = ~n18133 & n18137;
  assign n18139 = ~n18136 & n18138;
  assign n18140 = pi47  & n18139;
  assign n18141 = ~pi47  & ~n18139;
  assign n18142 = ~n18140 & ~n18141;
  assign n18143 = ~n17928 & ~n17931;
  assign n18144 = ~n17911 & ~n17924;
  assign n18145 = pi86  & n10886;
  assign n18146 = pi87  & n10495;
  assign n18147 = pi88  & n10490;
  assign n18148 = n2140 & n10488;
  assign n18149 = ~n18146 & ~n18147;
  assign n18150 = ~n18145 & n18149;
  assign n18151 = ~n18148 & n18150;
  assign n18152 = pi59  & n18151;
  assign n18153 = ~pi59  & ~n18151;
  assign n18154 = ~n18152 & ~n18153;
  assign n18155 = ~n17905 & ~n17907;
  assign n18156 = pi83  & n11910;
  assign n18157 = pi84  & n11529;
  assign n18158 = pi85  & n11524;
  assign n18159 = n1831 & n11522;
  assign n18160 = ~n18157 & ~n18158;
  assign n18161 = ~n18156 & n18160;
  assign n18162 = ~n18159 & n18161;
  assign n18163 = pi62  & n18162;
  assign n18164 = ~pi62  & ~n18162;
  assign n18165 = ~n18163 & ~n18164;
  assign n18166 = pi82  & n12277;
  assign n18167 = pi81  & n12276;
  assign n18168 = ~n18166 & ~n18167;
  assign n18169 = ~pi17  & ~n18168;
  assign n18170 = pi17  & n18168;
  assign n18171 = ~n18169 & ~n18170;
  assign n18172 = ~n17903 & n18171;
  assign n18173 = n17903 & ~n18171;
  assign n18174 = ~n18172 & ~n18173;
  assign n18175 = ~n18165 & n18174;
  assign n18176 = n18165 & ~n18174;
  assign n18177 = ~n18175 & ~n18176;
  assign n18178 = ~n18155 & n18177;
  assign n18179 = n18155 & ~n18177;
  assign n18180 = ~n18178 & ~n18179;
  assign n18181 = n18154 & ~n18180;
  assign n18182 = ~n18154 & n18180;
  assign n18183 = ~n18181 & ~n18182;
  assign n18184 = ~n18144 & n18183;
  assign n18185 = n18144 & ~n18183;
  assign n18186 = ~n18184 & ~n18185;
  assign n18187 = pi89  & n9858;
  assign n18188 = pi90  & n9508;
  assign n18189 = pi91  & n9503;
  assign n18190 = n2746 & n9501;
  assign n18191 = ~n18188 & ~n18189;
  assign n18192 = ~n18187 & n18191;
  assign n18193 = ~n18190 & n18192;
  assign n18194 = pi56  & n18193;
  assign n18195 = ~pi56  & ~n18193;
  assign n18196 = ~n18194 & ~n18195;
  assign n18197 = n18186 & ~n18196;
  assign n18198 = ~n18186 & n18196;
  assign n18199 = ~n18197 & ~n18198;
  assign n18200 = n18143 & ~n18199;
  assign n18201 = ~n18143 & n18199;
  assign n18202 = ~n18200 & ~n18201;
  assign n18203 = pi92  & n8905;
  assign n18204 = pi93  & n8535;
  assign n18205 = pi94  & n8530;
  assign n18206 = n3280 & n8528;
  assign n18207 = ~n18204 & ~n18205;
  assign n18208 = ~n18203 & n18207;
  assign n18209 = ~n18206 & n18208;
  assign n18210 = pi53  & n18209;
  assign n18211 = ~pi53  & ~n18209;
  assign n18212 = ~n18210 & ~n18211;
  assign n18213 = n18202 & ~n18212;
  assign n18214 = ~n18202 & n18212;
  assign n18215 = ~n18213 & ~n18214;
  assign n18216 = ~n17936 & n17948;
  assign n18217 = ~n17937 & ~n18216;
  assign n18218 = ~n18215 & ~n18217;
  assign n18219 = n18215 & n18217;
  assign n18220 = ~n18218 & ~n18219;
  assign n18221 = pi95  & n7969;
  assign n18222 = pi96  & n7636;
  assign n18223 = pi97  & n7631;
  assign n18224 = n3691 & n7629;
  assign n18225 = ~n18222 & ~n18223;
  assign n18226 = ~n18221 & n18225;
  assign n18227 = ~n18224 & n18226;
  assign n18228 = pi50  & n18227;
  assign n18229 = ~pi50  & ~n18227;
  assign n18230 = ~n18228 & ~n18229;
  assign n18231 = ~n17952 & ~n17955;
  assign n18232 = ~n18230 & ~n18231;
  assign n18233 = n18230 & n18231;
  assign n18234 = ~n18232 & ~n18233;
  assign n18235 = n18220 & n18234;
  assign n18236 = ~n18220 & ~n18234;
  assign n18237 = ~n18235 & ~n18236;
  assign n18238 = ~n18142 & n18237;
  assign n18239 = n18142 & ~n18237;
  assign n18240 = ~n18238 & ~n18239;
  assign n18241 = ~n17960 & ~n17972;
  assign n18242 = ~n17961 & ~n18241;
  assign n18243 = ~n18240 & n18242;
  assign n18244 = n18240 & ~n18242;
  assign n18245 = ~n18243 & ~n18244;
  assign n18246 = pi101  & n6331;
  assign n18247 = pi102  & n6015;
  assign n18248 = pi103  & n6010;
  assign n18249 = n5188 & n6008;
  assign n18250 = ~n18247 & ~n18248;
  assign n18251 = ~n18246 & n18250;
  assign n18252 = ~n18249 & n18251;
  assign n18253 = pi44  & n18252;
  assign n18254 = ~pi44  & ~n18252;
  assign n18255 = ~n18253 & ~n18254;
  assign n18256 = n18245 & ~n18255;
  assign n18257 = ~n18245 & n18255;
  assign n18258 = ~n18256 & ~n18257;
  assign n18259 = ~n18132 & n18258;
  assign n18260 = n18132 & ~n18258;
  assign n18261 = ~n18259 & ~n18260;
  assign n18262 = ~n18131 & n18261;
  assign n18263 = n18131 & ~n18261;
  assign n18264 = ~n18262 & ~n18263;
  assign n18265 = n18121 & ~n18264;
  assign n18266 = ~n18121 & n18264;
  assign n18267 = ~n18265 & ~n18266;
  assign n18268 = pi107  & n4843;
  assign n18269 = pi108  & n4598;
  assign n18270 = pi109  & n4593;
  assign n18271 = n4591 & n6715;
  assign n18272 = ~n18269 & ~n18270;
  assign n18273 = ~n18268 & n18272;
  assign n18274 = ~n18271 & n18273;
  assign n18275 = pi38  & n18274;
  assign n18276 = ~pi38  & ~n18274;
  assign n18277 = ~n18275 & ~n18276;
  assign n18278 = n18267 & ~n18277;
  assign n18279 = ~n18267 & n18277;
  assign n18280 = ~n18278 & ~n18279;
  assign n18281 = n18120 & ~n18280;
  assign n18282 = ~n18120 & n18280;
  assign n18283 = ~n18281 & ~n18282;
  assign n18284 = pi110  & n4176;
  assign n18285 = pi111  & n3938;
  assign n18286 = pi112  & n3933;
  assign n18287 = n3931 & n7296;
  assign n18288 = ~n18285 & ~n18286;
  assign n18289 = ~n18284 & n18288;
  assign n18290 = ~n18287 & n18289;
  assign n18291 = pi35  & n18290;
  assign n18292 = ~pi35  & ~n18290;
  assign n18293 = ~n18291 & ~n18292;
  assign n18294 = n18283 & ~n18293;
  assign n18295 = ~n18283 & n18293;
  assign n18296 = ~n18294 & ~n18295;
  assign n18297 = ~n17996 & n18008;
  assign n18298 = ~n17997 & ~n18297;
  assign n18299 = ~n18296 & ~n18298;
  assign n18300 = n18296 & n18298;
  assign n18301 = ~n18299 & ~n18300;
  assign n18302 = pi113  & n3553;
  assign n18303 = pi114  & n3334;
  assign n18304 = pi115  & n3329;
  assign n18305 = n3327 & n8170;
  assign n18306 = ~n18303 & ~n18304;
  assign n18307 = ~n18302 & n18306;
  assign n18308 = ~n18305 & n18307;
  assign n18309 = pi32  & n18308;
  assign n18310 = ~pi32  & ~n18308;
  assign n18311 = ~n18309 & ~n18310;
  assign n18312 = ~n17834 & ~n18012;
  assign n18313 = ~n18311 & ~n18312;
  assign n18314 = n18311 & n18312;
  assign n18315 = ~n18313 & ~n18314;
  assign n18316 = n18301 & n18315;
  assign n18317 = ~n18301 & ~n18315;
  assign n18318 = ~n18316 & ~n18317;
  assign n18319 = n18119 & ~n18318;
  assign n18320 = ~n18119 & n18318;
  assign n18321 = ~n18319 & ~n18320;
  assign n18322 = pi119  & n2510;
  assign n18323 = pi120  & n2342;
  assign n18324 = pi121  & n2337;
  assign n18325 = n2335 & n10071;
  assign n18326 = ~n18323 & ~n18324;
  assign n18327 = ~n18322 & n18326;
  assign n18328 = ~n18325 & n18327;
  assign n18329 = pi26  & n18328;
  assign n18330 = ~pi26  & ~n18328;
  assign n18331 = ~n18329 & ~n18330;
  assign n18332 = ~n17819 & ~n18032;
  assign n18333 = ~n18331 & ~n18332;
  assign n18334 = n18331 & n18332;
  assign n18335 = ~n18333 & ~n18334;
  assign n18336 = n18321 & ~n18335;
  assign n18337 = ~n18321 & n18335;
  assign n18338 = ~n18336 & ~n18337;
  assign n18339 = n18105 & n18338;
  assign n18340 = ~n18105 & ~n18338;
  assign n18341 = ~n18339 & ~n18340;
  assign n18342 = n18091 & n18341;
  assign n18343 = ~n18091 & ~n18341;
  assign n18344 = ~n18342 & ~n18343;
  assign n18345 = ~n18077 & n18344;
  assign n18346 = n18077 & ~n18344;
  assign n18347 = ~n18345 & ~n18346;
  assign n18348 = ~n18076 & n18347;
  assign n18349 = n18076 & ~n18347;
  assign po81  = ~n18348 & ~n18349;
  assign n18351 = ~n18345 & ~n18348;
  assign n18352 = ~n18089 & ~n18342;
  assign n18353 = pi126  & n1661;
  assign n18354 = pi127  & n1500;
  assign n18355 = n1493 & n12542;
  assign n18356 = ~n18353 & ~n18354;
  assign n18357 = ~n18355 & n18356;
  assign n18358 = pi20  & n18357;
  assign n18359 = ~pi20  & ~n18357;
  assign n18360 = ~n18358 & ~n18359;
  assign n18361 = ~n18104 & ~n18338;
  assign n18362 = ~n18103 & ~n18361;
  assign n18363 = ~n18360 & n18362;
  assign n18364 = n18360 & ~n18362;
  assign n18365 = ~n18363 & ~n18364;
  assign n18366 = pi123  & n2053;
  assign n18367 = pi124  & n1893;
  assign n18368 = pi125  & n1888;
  assign n18369 = n1886 & n11786;
  assign n18370 = ~n18367 & ~n18368;
  assign n18371 = ~n18366 & n18370;
  assign n18372 = ~n18369 & n18371;
  assign n18373 = pi23  & n18372;
  assign n18374 = ~pi23  & ~n18372;
  assign n18375 = ~n18373 & ~n18374;
  assign n18376 = n18321 & ~n18333;
  assign n18377 = ~n18334 & ~n18376;
  assign n18378 = n18375 & ~n18377;
  assign n18379 = ~n18375 & n18377;
  assign n18380 = ~n18378 & ~n18379;
  assign n18381 = pi120  & n2510;
  assign n18382 = pi121  & n2342;
  assign n18383 = pi122  & n2337;
  assign n18384 = n2335 & n10729;
  assign n18385 = ~n18382 & ~n18383;
  assign n18386 = ~n18381 & n18385;
  assign n18387 = ~n18384 & n18386;
  assign n18388 = pi26  & n18387;
  assign n18389 = ~pi26  & ~n18387;
  assign n18390 = ~n18388 & ~n18389;
  assign n18391 = ~n18118 & ~n18318;
  assign n18392 = ~n18117 & ~n18391;
  assign n18393 = n18390 & ~n18392;
  assign n18394 = ~n18390 & n18392;
  assign n18395 = ~n18393 & ~n18394;
  assign n18396 = pi117  & n3011;
  assign n18397 = pi118  & n2809;
  assign n18398 = pi119  & n2804;
  assign n18399 = n2802 & n9412;
  assign n18400 = ~n18397 & ~n18398;
  assign n18401 = ~n18396 & n18400;
  assign n18402 = ~n18399 & n18401;
  assign n18403 = pi29  & n18402;
  assign n18404 = ~pi29  & ~n18402;
  assign n18405 = ~n18403 & ~n18404;
  assign n18406 = n18301 & ~n18314;
  assign n18407 = ~n18313 & ~n18406;
  assign n18408 = n18405 & n18407;
  assign n18409 = ~n18405 & ~n18407;
  assign n18410 = ~n18408 & ~n18409;
  assign n18411 = pi114  & n3553;
  assign n18412 = pi115  & n3334;
  assign n18413 = pi116  & n3329;
  assign n18414 = n3327 & n8470;
  assign n18415 = ~n18412 & ~n18413;
  assign n18416 = ~n18411 & n18415;
  assign n18417 = ~n18414 & n18416;
  assign n18418 = pi32  & n18417;
  assign n18419 = ~pi32  & ~n18417;
  assign n18420 = ~n18418 & ~n18419;
  assign n18421 = ~n18294 & ~n18300;
  assign n18422 = n18420 & n18421;
  assign n18423 = ~n18420 & ~n18421;
  assign n18424 = ~n18422 & ~n18423;
  assign n18425 = ~n18278 & ~n18282;
  assign n18426 = ~n18262 & ~n18266;
  assign n18427 = ~n18256 & ~n18259;
  assign n18428 = pi102  & n6331;
  assign n18429 = pi103  & n6015;
  assign n18430 = pi104  & n6010;
  assign n18431 = n5212 & n6008;
  assign n18432 = ~n18429 & ~n18430;
  assign n18433 = ~n18428 & n18432;
  assign n18434 = ~n18431 & n18433;
  assign n18435 = pi44  & n18434;
  assign n18436 = ~pi44  & ~n18434;
  assign n18437 = ~n18435 & ~n18436;
  assign n18438 = ~n18238 & ~n18244;
  assign n18439 = ~n18232 & ~n18235;
  assign n18440 = ~n18213 & ~n18219;
  assign n18441 = pi90  & n9858;
  assign n18442 = pi91  & n9508;
  assign n18443 = pi92  & n9503;
  assign n18444 = n2924 & n9501;
  assign n18445 = ~n18442 & ~n18443;
  assign n18446 = ~n18441 & n18445;
  assign n18447 = ~n18444 & n18446;
  assign n18448 = pi56  & n18447;
  assign n18449 = ~pi56  & ~n18447;
  assign n18450 = ~n18448 & ~n18449;
  assign n18451 = ~n18182 & ~n18184;
  assign n18452 = ~n18169 & ~n18172;
  assign n18453 = pi83  & n12277;
  assign n18454 = pi82  & n12276;
  assign n18455 = ~n18453 & ~n18454;
  assign n18456 = n18452 & ~n18455;
  assign n18457 = ~n18452 & n18455;
  assign n18458 = ~n18456 & ~n18457;
  assign n18459 = pi84  & n11910;
  assign n18460 = pi85  & n11529;
  assign n18461 = pi86  & n11524;
  assign n18462 = n1975 & n11522;
  assign n18463 = ~n18460 & ~n18461;
  assign n18464 = ~n18459 & n18463;
  assign n18465 = ~n18462 & n18464;
  assign n18466 = pi62  & n18465;
  assign n18467 = ~pi62  & ~n18465;
  assign n18468 = ~n18466 & ~n18467;
  assign n18469 = ~n18458 & n18468;
  assign n18470 = n18458 & ~n18468;
  assign n18471 = ~n18469 & ~n18470;
  assign n18472 = ~n18175 & ~n18178;
  assign n18473 = n18471 & ~n18472;
  assign n18474 = ~n18471 & n18472;
  assign n18475 = ~n18473 & ~n18474;
  assign n18476 = pi87  & n10886;
  assign n18477 = pi88  & n10495;
  assign n18478 = pi89  & n10490;
  assign n18479 = n2287 & n10488;
  assign n18480 = ~n18477 & ~n18478;
  assign n18481 = ~n18476 & n18480;
  assign n18482 = ~n18479 & n18481;
  assign n18483 = pi59  & n18482;
  assign n18484 = ~pi59  & ~n18482;
  assign n18485 = ~n18483 & ~n18484;
  assign n18486 = n18475 & ~n18485;
  assign n18487 = ~n18475 & n18485;
  assign n18488 = ~n18486 & ~n18487;
  assign n18489 = ~n18451 & n18488;
  assign n18490 = n18451 & ~n18488;
  assign n18491 = ~n18489 & ~n18490;
  assign n18492 = n18450 & ~n18491;
  assign n18493 = ~n18450 & n18491;
  assign n18494 = ~n18492 & ~n18493;
  assign n18495 = ~n18197 & ~n18201;
  assign n18496 = n18494 & ~n18495;
  assign n18497 = ~n18494 & n18495;
  assign n18498 = ~n18496 & ~n18497;
  assign n18499 = pi93  & n8905;
  assign n18500 = pi94  & n8535;
  assign n18501 = pi95  & n8530;
  assign n18502 = n3475 & n8528;
  assign n18503 = ~n18500 & ~n18501;
  assign n18504 = ~n18499 & n18503;
  assign n18505 = ~n18502 & n18504;
  assign n18506 = pi53  & n18505;
  assign n18507 = ~pi53  & ~n18505;
  assign n18508 = ~n18506 & ~n18507;
  assign n18509 = n18498 & ~n18508;
  assign n18510 = ~n18498 & n18508;
  assign n18511 = ~n18509 & ~n18510;
  assign n18512 = n18440 & ~n18511;
  assign n18513 = ~n18440 & n18511;
  assign n18514 = ~n18512 & ~n18513;
  assign n18515 = pi96  & n7969;
  assign n18516 = pi97  & n7636;
  assign n18517 = pi98  & n7631;
  assign n18518 = n3889 & n7629;
  assign n18519 = ~n18516 & ~n18517;
  assign n18520 = ~n18515 & n18519;
  assign n18521 = ~n18518 & n18520;
  assign n18522 = pi50  & n18521;
  assign n18523 = ~pi50  & ~n18521;
  assign n18524 = ~n18522 & ~n18523;
  assign n18525 = n18514 & ~n18524;
  assign n18526 = ~n18514 & n18524;
  assign n18527 = ~n18525 & ~n18526;
  assign n18528 = n18439 & ~n18527;
  assign n18529 = ~n18439 & n18527;
  assign n18530 = ~n18528 & ~n18529;
  assign n18531 = pi99  & n7121;
  assign n18532 = pi100  & n6795;
  assign n18533 = pi101  & n6790;
  assign n18534 = n4730 & n6788;
  assign n18535 = ~n18532 & ~n18533;
  assign n18536 = ~n18531 & n18535;
  assign n18537 = ~n18534 & n18536;
  assign n18538 = pi47  & n18537;
  assign n18539 = ~pi47  & ~n18537;
  assign n18540 = ~n18538 & ~n18539;
  assign n18541 = ~n18530 & n18540;
  assign n18542 = n18530 & ~n18540;
  assign n18543 = ~n18541 & ~n18542;
  assign n18544 = ~n18438 & n18543;
  assign n18545 = n18438 & ~n18543;
  assign n18546 = ~n18544 & ~n18545;
  assign n18547 = ~n18437 & n18546;
  assign n18548 = n18437 & ~n18546;
  assign n18549 = ~n18547 & ~n18548;
  assign n18550 = ~n18427 & n18549;
  assign n18551 = n18427 & ~n18549;
  assign n18552 = ~n18550 & ~n18551;
  assign n18553 = pi105  & n5558;
  assign n18554 = pi106  & n5293;
  assign n18555 = pi107  & n5288;
  assign n18556 = n5286 & n6189;
  assign n18557 = ~n18554 & ~n18555;
  assign n18558 = ~n18553 & n18557;
  assign n18559 = ~n18556 & n18558;
  assign n18560 = pi41  & n18559;
  assign n18561 = ~pi41  & ~n18559;
  assign n18562 = ~n18560 & ~n18561;
  assign n18563 = n18552 & ~n18562;
  assign n18564 = ~n18552 & n18562;
  assign n18565 = ~n18563 & ~n18564;
  assign n18566 = n18426 & ~n18565;
  assign n18567 = ~n18426 & n18565;
  assign n18568 = ~n18566 & ~n18567;
  assign n18569 = pi108  & n4843;
  assign n18570 = pi109  & n4598;
  assign n18571 = pi110  & n4593;
  assign n18572 = n4591 & n6995;
  assign n18573 = ~n18570 & ~n18571;
  assign n18574 = ~n18569 & n18573;
  assign n18575 = ~n18572 & n18574;
  assign n18576 = pi38  & n18575;
  assign n18577 = ~pi38  & ~n18575;
  assign n18578 = ~n18576 & ~n18577;
  assign n18579 = n18568 & ~n18578;
  assign n18580 = ~n18568 & n18578;
  assign n18581 = ~n18579 & ~n18580;
  assign n18582 = n18425 & ~n18581;
  assign n18583 = ~n18425 & n18581;
  assign n18584 = ~n18582 & ~n18583;
  assign n18585 = pi111  & n4176;
  assign n18586 = pi112  & n3938;
  assign n18587 = pi113  & n3933;
  assign n18588 = n3931 & n7852;
  assign n18589 = ~n18586 & ~n18587;
  assign n18590 = ~n18585 & n18589;
  assign n18591 = ~n18588 & n18590;
  assign n18592 = pi35  & n18591;
  assign n18593 = ~pi35  & ~n18591;
  assign n18594 = ~n18592 & ~n18593;
  assign n18595 = n18584 & ~n18594;
  assign n18596 = ~n18584 & n18594;
  assign n18597 = ~n18595 & ~n18596;
  assign n18598 = n18424 & n18597;
  assign n18599 = ~n18424 & ~n18597;
  assign n18600 = ~n18598 & ~n18599;
  assign n18601 = n18410 & n18600;
  assign n18602 = ~n18410 & ~n18600;
  assign n18603 = ~n18601 & ~n18602;
  assign n18604 = n18395 & n18603;
  assign n18605 = ~n18395 & ~n18603;
  assign n18606 = ~n18604 & ~n18605;
  assign n18607 = n18380 & n18606;
  assign n18608 = ~n18380 & ~n18606;
  assign n18609 = ~n18607 & ~n18608;
  assign n18610 = n18365 & n18609;
  assign n18611 = ~n18365 & ~n18609;
  assign n18612 = ~n18610 & ~n18611;
  assign n18613 = ~n18352 & n18612;
  assign n18614 = n18352 & ~n18612;
  assign n18615 = ~n18613 & ~n18614;
  assign n18616 = ~n18351 & n18615;
  assign n18617 = n18351 & ~n18615;
  assign po82  = ~n18616 & ~n18617;
  assign n18619 = ~n18613 & ~n18616;
  assign n18620 = ~n18363 & ~n18610;
  assign n18621 = pi121  & n2510;
  assign n18622 = pi122  & n2342;
  assign n18623 = pi123  & n2337;
  assign n18624 = n2335 & n10754;
  assign n18625 = ~n18622 & ~n18623;
  assign n18626 = ~n18621 & n18625;
  assign n18627 = ~n18624 & n18626;
  assign n18628 = pi26  & n18627;
  assign n18629 = ~pi26  & ~n18627;
  assign n18630 = ~n18628 & ~n18629;
  assign n18631 = ~n18409 & ~n18601;
  assign n18632 = n18630 & n18631;
  assign n18633 = ~n18630 & ~n18631;
  assign n18634 = ~n18632 & ~n18633;
  assign n18635 = pi115  & n3553;
  assign n18636 = pi116  & n3334;
  assign n18637 = pi117  & n3329;
  assign n18638 = n3327 & n8784;
  assign n18639 = ~n18636 & ~n18637;
  assign n18640 = ~n18635 & n18639;
  assign n18641 = ~n18638 & n18640;
  assign n18642 = pi32  & n18641;
  assign n18643 = ~pi32  & ~n18641;
  assign n18644 = ~n18642 & ~n18643;
  assign n18645 = ~n18583 & n18594;
  assign n18646 = ~n18582 & ~n18645;
  assign n18647 = n18644 & ~n18646;
  assign n18648 = ~n18644 & n18646;
  assign n18649 = ~n18647 & ~n18648;
  assign n18650 = pi106  & n5558;
  assign n18651 = pi107  & n5293;
  assign n18652 = pi108  & n5288;
  assign n18653 = n5286 & n6213;
  assign n18654 = ~n18651 & ~n18652;
  assign n18655 = ~n18650 & n18654;
  assign n18656 = ~n18653 & n18655;
  assign n18657 = pi41  & n18656;
  assign n18658 = ~pi41  & ~n18656;
  assign n18659 = ~n18657 & ~n18658;
  assign n18660 = ~n18544 & ~n18547;
  assign n18661 = pi103  & n6331;
  assign n18662 = pi104  & n6015;
  assign n18663 = pi105  & n6010;
  assign n18664 = n5677 & n6008;
  assign n18665 = ~n18662 & ~n18663;
  assign n18666 = ~n18661 & n18665;
  assign n18667 = ~n18664 & n18666;
  assign n18668 = pi44  & n18667;
  assign n18669 = ~pi44  & ~n18667;
  assign n18670 = ~n18668 & ~n18669;
  assign n18671 = ~n18529 & ~n18542;
  assign n18672 = pi100  & n7121;
  assign n18673 = pi101  & n6795;
  assign n18674 = pi102  & n6790;
  assign n18675 = n4956 & n6788;
  assign n18676 = ~n18673 & ~n18674;
  assign n18677 = ~n18672 & n18676;
  assign n18678 = ~n18675 & n18677;
  assign n18679 = pi47  & n18678;
  assign n18680 = ~pi47  & ~n18678;
  assign n18681 = ~n18679 & ~n18680;
  assign n18682 = pi97  & n7969;
  assign n18683 = pi98  & n7636;
  assign n18684 = pi99  & n7631;
  assign n18685 = n4101 & n7629;
  assign n18686 = ~n18683 & ~n18684;
  assign n18687 = ~n18682 & n18686;
  assign n18688 = ~n18685 & n18687;
  assign n18689 = pi50  & n18688;
  assign n18690 = ~pi50  & ~n18688;
  assign n18691 = ~n18689 & ~n18690;
  assign n18692 = pi94  & n8905;
  assign n18693 = pi95  & n8535;
  assign n18694 = pi96  & n8530;
  assign n18695 = n3499 & n8528;
  assign n18696 = ~n18693 & ~n18694;
  assign n18697 = ~n18692 & n18696;
  assign n18698 = ~n18695 & n18697;
  assign n18699 = pi53  & n18698;
  assign n18700 = ~pi53  & ~n18698;
  assign n18701 = ~n18699 & ~n18700;
  assign n18702 = ~n18489 & ~n18493;
  assign n18703 = pi88  & n10886;
  assign n18704 = pi89  & n10495;
  assign n18705 = pi90  & n10490;
  assign n18706 = n2448 & n10488;
  assign n18707 = ~n18704 & ~n18705;
  assign n18708 = ~n18703 & n18707;
  assign n18709 = ~n18706 & n18708;
  assign n18710 = pi59  & n18709;
  assign n18711 = ~pi59  & ~n18709;
  assign n18712 = ~n18710 & ~n18711;
  assign n18713 = ~n18457 & ~n18470;
  assign n18714 = pi84  & n12277;
  assign n18715 = pi83  & n12276;
  assign n18716 = ~n18714 & ~n18715;
  assign n18717 = ~n18455 & n18716;
  assign n18718 = n18455 & ~n18716;
  assign n18719 = ~n18717 & ~n18718;
  assign n18720 = pi85  & n11910;
  assign n18721 = pi86  & n11529;
  assign n18722 = pi87  & n11524;
  assign n18723 = n2116 & n11522;
  assign n18724 = ~n18721 & ~n18722;
  assign n18725 = ~n18720 & n18724;
  assign n18726 = ~n18723 & n18725;
  assign n18727 = pi62  & n18726;
  assign n18728 = ~pi62  & ~n18726;
  assign n18729 = ~n18727 & ~n18728;
  assign n18730 = n18719 & ~n18729;
  assign n18731 = ~n18719 & n18729;
  assign n18732 = ~n18730 & ~n18731;
  assign n18733 = ~n18713 & n18732;
  assign n18734 = n18713 & ~n18732;
  assign n18735 = ~n18733 & ~n18734;
  assign n18736 = ~n18712 & n18735;
  assign n18737 = n18712 & ~n18735;
  assign n18738 = ~n18736 & ~n18737;
  assign n18739 = ~n18474 & ~n18485;
  assign n18740 = ~n18473 & ~n18739;
  assign n18741 = n18738 & ~n18740;
  assign n18742 = ~n18738 & n18740;
  assign n18743 = ~n18741 & ~n18742;
  assign n18744 = pi91  & n9858;
  assign n18745 = pi92  & n9508;
  assign n18746 = pi93  & n9503;
  assign n18747 = n2948 & n9501;
  assign n18748 = ~n18745 & ~n18746;
  assign n18749 = ~n18744 & n18748;
  assign n18750 = ~n18747 & n18749;
  assign n18751 = pi56  & n18750;
  assign n18752 = ~pi56  & ~n18750;
  assign n18753 = ~n18751 & ~n18752;
  assign n18754 = n18743 & ~n18753;
  assign n18755 = ~n18743 & n18753;
  assign n18756 = ~n18754 & ~n18755;
  assign n18757 = ~n18702 & n18756;
  assign n18758 = n18702 & ~n18756;
  assign n18759 = ~n18757 & ~n18758;
  assign n18760 = ~n18701 & n18759;
  assign n18761 = n18701 & ~n18759;
  assign n18762 = ~n18760 & ~n18761;
  assign n18763 = ~n18497 & ~n18508;
  assign n18764 = ~n18496 & ~n18763;
  assign n18765 = n18762 & ~n18764;
  assign n18766 = ~n18762 & n18764;
  assign n18767 = ~n18765 & ~n18766;
  assign n18768 = ~n18691 & n18767;
  assign n18769 = n18691 & ~n18767;
  assign n18770 = ~n18768 & ~n18769;
  assign n18771 = ~n18513 & n18524;
  assign n18772 = ~n18512 & ~n18771;
  assign n18773 = n18770 & n18772;
  assign n18774 = ~n18770 & ~n18772;
  assign n18775 = ~n18773 & ~n18774;
  assign n18776 = ~n18681 & n18775;
  assign n18777 = n18681 & ~n18775;
  assign n18778 = ~n18776 & ~n18777;
  assign n18779 = ~n18671 & n18778;
  assign n18780 = n18671 & ~n18778;
  assign n18781 = ~n18779 & ~n18780;
  assign n18782 = ~n18670 & n18781;
  assign n18783 = n18670 & ~n18781;
  assign n18784 = ~n18782 & ~n18783;
  assign n18785 = ~n18660 & n18784;
  assign n18786 = n18660 & ~n18784;
  assign n18787 = ~n18785 & ~n18786;
  assign n18788 = ~n18659 & n18787;
  assign n18789 = n18659 & ~n18787;
  assign n18790 = ~n18788 & ~n18789;
  assign n18791 = ~n18550 & n18562;
  assign n18792 = ~n18551 & ~n18791;
  assign n18793 = n18790 & n18792;
  assign n18794 = ~n18790 & ~n18792;
  assign n18795 = ~n18793 & ~n18794;
  assign n18796 = pi109  & n4843;
  assign n18797 = pi110  & n4598;
  assign n18798 = pi111  & n4593;
  assign n18799 = n4591 & n7272;
  assign n18800 = ~n18797 & ~n18798;
  assign n18801 = ~n18796 & n18800;
  assign n18802 = ~n18799 & n18801;
  assign n18803 = pi38  & n18802;
  assign n18804 = ~pi38  & ~n18802;
  assign n18805 = ~n18803 & ~n18804;
  assign n18806 = n18795 & ~n18805;
  assign n18807 = ~n18795 & n18805;
  assign n18808 = ~n18806 & ~n18807;
  assign n18809 = ~n18567 & n18578;
  assign n18810 = ~n18566 & ~n18809;
  assign n18811 = ~n18808 & ~n18810;
  assign n18812 = n18808 & n18810;
  assign n18813 = ~n18811 & ~n18812;
  assign n18814 = pi112  & n4176;
  assign n18815 = pi113  & n3938;
  assign n18816 = pi114  & n3933;
  assign n18817 = n3931 & n8146;
  assign n18818 = ~n18815 & ~n18816;
  assign n18819 = ~n18814 & n18818;
  assign n18820 = ~n18817 & n18819;
  assign n18821 = pi35  & n18820;
  assign n18822 = ~pi35  & ~n18820;
  assign n18823 = ~n18821 & ~n18822;
  assign n18824 = n18813 & ~n18823;
  assign n18825 = ~n18813 & n18823;
  assign n18826 = ~n18824 & ~n18825;
  assign n18827 = n18649 & n18826;
  assign n18828 = ~n18649 & ~n18826;
  assign n18829 = ~n18827 & ~n18828;
  assign n18830 = pi118  & n3011;
  assign n18831 = pi119  & n2809;
  assign n18832 = pi120  & n2804;
  assign n18833 = n2802 & n10047;
  assign n18834 = ~n18831 & ~n18832;
  assign n18835 = ~n18830 & n18834;
  assign n18836 = ~n18833 & n18835;
  assign n18837 = pi29  & n18836;
  assign n18838 = ~pi29  & ~n18836;
  assign n18839 = ~n18837 & ~n18838;
  assign n18840 = ~n18423 & ~n18598;
  assign n18841 = ~n18839 & ~n18840;
  assign n18842 = n18839 & n18840;
  assign n18843 = ~n18841 & ~n18842;
  assign n18844 = n18829 & n18843;
  assign n18845 = ~n18829 & ~n18843;
  assign n18846 = ~n18844 & ~n18845;
  assign n18847 = n18634 & n18846;
  assign n18848 = ~n18634 & ~n18846;
  assign n18849 = ~n18847 & ~n18848;
  assign n18850 = pi124  & n2053;
  assign n18851 = pi125  & n1893;
  assign n18852 = pi126  & n1888;
  assign n18853 = n1886 & n12148;
  assign n18854 = ~n18851 & ~n18852;
  assign n18855 = ~n18850 & n18854;
  assign n18856 = ~n18853 & n18855;
  assign n18857 = pi23  & n18856;
  assign n18858 = ~pi23  & ~n18856;
  assign n18859 = ~n18857 & ~n18858;
  assign n18860 = ~n18394 & ~n18604;
  assign n18861 = ~n18859 & ~n18860;
  assign n18862 = n18859 & n18860;
  assign n18863 = ~n18861 & ~n18862;
  assign n18864 = n18849 & n18863;
  assign n18865 = ~n18849 & ~n18863;
  assign n18866 = ~n18864 & ~n18865;
  assign n18867 = n1493 & ~n12539;
  assign n18868 = ~n1661 & ~n18867;
  assign n18869 = pi127  & ~n18868;
  assign n18870 = pi20  & ~n18869;
  assign n18871 = ~pi20  & n18869;
  assign n18872 = ~n18870 & ~n18871;
  assign n18873 = ~n18379 & ~n18606;
  assign n18874 = ~n18378 & ~n18873;
  assign n18875 = ~n18872 & n18874;
  assign n18876 = n18872 & ~n18874;
  assign n18877 = ~n18875 & ~n18876;
  assign n18878 = n18866 & n18877;
  assign n18879 = ~n18866 & ~n18877;
  assign n18880 = ~n18878 & ~n18879;
  assign n18881 = ~n18620 & n18880;
  assign n18882 = n18620 & ~n18880;
  assign n18883 = ~n18881 & ~n18882;
  assign n18884 = ~n18619 & n18883;
  assign n18885 = n18619 & ~n18883;
  assign po83  = ~n18884 & ~n18885;
  assign n18887 = ~n18875 & ~n18878;
  assign n18888 = pi122  & n2510;
  assign n18889 = pi123  & n2342;
  assign n18890 = pi124  & n2337;
  assign n18891 = n2335 & n11099;
  assign n18892 = ~n18889 & ~n18890;
  assign n18893 = ~n18888 & n18892;
  assign n18894 = ~n18891 & n18893;
  assign n18895 = pi26  & n18894;
  assign n18896 = ~pi26  & ~n18894;
  assign n18897 = ~n18895 & ~n18896;
  assign n18898 = ~n18633 & ~n18847;
  assign n18899 = n18897 & n18898;
  assign n18900 = ~n18897 & ~n18898;
  assign n18901 = ~n18899 & ~n18900;
  assign n18902 = pi116  & n3553;
  assign n18903 = pi117  & n3334;
  assign n18904 = pi118  & n3329;
  assign n18905 = n3327 & n9095;
  assign n18906 = ~n18903 & ~n18904;
  assign n18907 = ~n18902 & n18906;
  assign n18908 = ~n18905 & n18907;
  assign n18909 = pi32  & n18908;
  assign n18910 = ~pi32  & ~n18908;
  assign n18911 = ~n18909 & ~n18910;
  assign n18912 = ~n18648 & ~n18827;
  assign n18913 = n18911 & n18912;
  assign n18914 = ~n18911 & ~n18912;
  assign n18915 = ~n18913 & ~n18914;
  assign n18916 = ~n18812 & ~n18824;
  assign n18917 = ~n18785 & ~n18788;
  assign n18918 = ~n18779 & ~n18782;
  assign n18919 = ~n18773 & ~n18776;
  assign n18920 = ~n18765 & ~n18768;
  assign n18921 = pi98  & n7969;
  assign n18922 = pi99  & n7636;
  assign n18923 = pi100  & n7631;
  assign n18924 = n4501 & n7629;
  assign n18925 = ~n18922 & ~n18923;
  assign n18926 = ~n18921 & n18925;
  assign n18927 = ~n18924 & n18926;
  assign n18928 = pi50  & n18927;
  assign n18929 = ~pi50  & ~n18927;
  assign n18930 = ~n18928 & ~n18929;
  assign n18931 = ~n18742 & ~n18753;
  assign n18932 = ~n18741 & ~n18931;
  assign n18933 = ~n18733 & ~n18736;
  assign n18934 = pi89  & n10886;
  assign n18935 = pi90  & n10495;
  assign n18936 = pi91  & n10490;
  assign n18937 = n2746 & n10488;
  assign n18938 = ~n18935 & ~n18936;
  assign n18939 = ~n18934 & n18938;
  assign n18940 = ~n18937 & n18939;
  assign n18941 = pi59  & n18940;
  assign n18942 = ~pi59  & ~n18940;
  assign n18943 = ~n18941 & ~n18942;
  assign n18944 = ~n18717 & ~n18730;
  assign n18945 = pi85  & n12277;
  assign n18946 = pi84  & n12276;
  assign n18947 = ~n18945 & ~n18946;
  assign n18948 = ~pi20  & ~n18947;
  assign n18949 = pi20  & n18947;
  assign n18950 = ~n18948 & ~n18949;
  assign n18951 = ~n18716 & n18950;
  assign n18952 = n18716 & ~n18950;
  assign n18953 = ~n18951 & ~n18952;
  assign n18954 = pi86  & n11910;
  assign n18955 = pi87  & n11529;
  assign n18956 = pi88  & n11524;
  assign n18957 = n2140 & n11522;
  assign n18958 = ~n18955 & ~n18956;
  assign n18959 = ~n18954 & n18958;
  assign n18960 = ~n18957 & n18959;
  assign n18961 = pi62  & n18960;
  assign n18962 = ~pi62  & ~n18960;
  assign n18963 = ~n18961 & ~n18962;
  assign n18964 = n18953 & ~n18963;
  assign n18965 = ~n18953 & n18963;
  assign n18966 = ~n18964 & ~n18965;
  assign n18967 = ~n18944 & n18966;
  assign n18968 = n18944 & ~n18966;
  assign n18969 = ~n18967 & ~n18968;
  assign n18970 = ~n18943 & n18969;
  assign n18971 = n18943 & ~n18969;
  assign n18972 = ~n18970 & ~n18971;
  assign n18973 = n18933 & ~n18972;
  assign n18974 = ~n18933 & n18972;
  assign n18975 = ~n18973 & ~n18974;
  assign n18976 = pi92  & n9858;
  assign n18977 = pi93  & n9508;
  assign n18978 = pi94  & n9503;
  assign n18979 = n3280 & n9501;
  assign n18980 = ~n18977 & ~n18978;
  assign n18981 = ~n18976 & n18980;
  assign n18982 = ~n18979 & n18981;
  assign n18983 = pi56  & n18982;
  assign n18984 = ~pi56  & ~n18982;
  assign n18985 = ~n18983 & ~n18984;
  assign n18986 = n18975 & ~n18985;
  assign n18987 = ~n18975 & n18985;
  assign n18988 = ~n18986 & ~n18987;
  assign n18989 = n18932 & ~n18988;
  assign n18990 = ~n18932 & n18988;
  assign n18991 = ~n18989 & ~n18990;
  assign n18992 = pi95  & n8905;
  assign n18993 = pi96  & n8535;
  assign n18994 = pi97  & n8530;
  assign n18995 = n3691 & n8528;
  assign n18996 = ~n18993 & ~n18994;
  assign n18997 = ~n18992 & n18996;
  assign n18998 = ~n18995 & n18997;
  assign n18999 = pi53  & n18998;
  assign n19000 = ~pi53  & ~n18998;
  assign n19001 = ~n18999 & ~n19000;
  assign n19002 = ~n18757 & ~n18760;
  assign n19003 = ~n19001 & ~n19002;
  assign n19004 = n19001 & n19002;
  assign n19005 = ~n19003 & ~n19004;
  assign n19006 = n18991 & n19005;
  assign n19007 = ~n18991 & ~n19005;
  assign n19008 = ~n19006 & ~n19007;
  assign n19009 = ~n18930 & n19008;
  assign n19010 = n18930 & ~n19008;
  assign n19011 = ~n19009 & ~n19010;
  assign n19012 = n18920 & ~n19011;
  assign n19013 = ~n18920 & n19011;
  assign n19014 = ~n19012 & ~n19013;
  assign n19015 = pi101  & n7121;
  assign n19016 = pi102  & n6795;
  assign n19017 = pi103  & n6790;
  assign n19018 = n5188 & n6788;
  assign n19019 = ~n19016 & ~n19017;
  assign n19020 = ~n19015 & n19019;
  assign n19021 = ~n19018 & n19020;
  assign n19022 = pi47  & n19021;
  assign n19023 = ~pi47  & ~n19021;
  assign n19024 = ~n19022 & ~n19023;
  assign n19025 = n19014 & ~n19024;
  assign n19026 = ~n19014 & n19024;
  assign n19027 = ~n19025 & ~n19026;
  assign n19028 = n18919 & ~n19027;
  assign n19029 = ~n18919 & n19027;
  assign n19030 = ~n19028 & ~n19029;
  assign n19031 = pi104  & n6331;
  assign n19032 = pi105  & n6015;
  assign n19033 = pi106  & n6010;
  assign n19034 = n5701 & n6008;
  assign n19035 = ~n19032 & ~n19033;
  assign n19036 = ~n19031 & n19035;
  assign n19037 = ~n19034 & n19036;
  assign n19038 = pi44  & n19037;
  assign n19039 = ~pi44  & ~n19037;
  assign n19040 = ~n19038 & ~n19039;
  assign n19041 = n19030 & ~n19040;
  assign n19042 = ~n19030 & n19040;
  assign n19043 = ~n19041 & ~n19042;
  assign n19044 = n18918 & ~n19043;
  assign n19045 = ~n18918 & n19043;
  assign n19046 = ~n19044 & ~n19045;
  assign n19047 = pi107  & n5558;
  assign n19048 = pi108  & n5293;
  assign n19049 = pi109  & n5288;
  assign n19050 = n5286 & n6715;
  assign n19051 = ~n19048 & ~n19049;
  assign n19052 = ~n19047 & n19051;
  assign n19053 = ~n19050 & n19052;
  assign n19054 = pi41  & n19053;
  assign n19055 = ~pi41  & ~n19053;
  assign n19056 = ~n19054 & ~n19055;
  assign n19057 = n19046 & ~n19056;
  assign n19058 = ~n19046 & n19056;
  assign n19059 = ~n19057 & ~n19058;
  assign n19060 = n18917 & ~n19059;
  assign n19061 = ~n18917 & n19059;
  assign n19062 = ~n19060 & ~n19061;
  assign n19063 = pi110  & n4843;
  assign n19064 = pi111  & n4598;
  assign n19065 = pi112  & n4593;
  assign n19066 = n4591 & n7296;
  assign n19067 = ~n19064 & ~n19065;
  assign n19068 = ~n19063 & n19067;
  assign n19069 = ~n19066 & n19068;
  assign n19070 = pi38  & n19069;
  assign n19071 = ~pi38  & ~n19069;
  assign n19072 = ~n19070 & ~n19071;
  assign n19073 = n19062 & ~n19072;
  assign n19074 = ~n19062 & n19072;
  assign n19075 = ~n19073 & ~n19074;
  assign n19076 = ~n18793 & n18805;
  assign n19077 = ~n18794 & ~n19076;
  assign n19078 = ~n19075 & ~n19077;
  assign n19079 = n19075 & n19077;
  assign n19080 = ~n19078 & ~n19079;
  assign n19081 = pi113  & n4176;
  assign n19082 = pi114  & n3938;
  assign n19083 = pi115  & n3933;
  assign n19084 = n3931 & n8170;
  assign n19085 = ~n19082 & ~n19083;
  assign n19086 = ~n19081 & n19085;
  assign n19087 = ~n19084 & n19086;
  assign n19088 = pi35  & n19087;
  assign n19089 = ~pi35  & ~n19087;
  assign n19090 = ~n19088 & ~n19089;
  assign n19091 = n19080 & ~n19090;
  assign n19092 = ~n19080 & n19090;
  assign n19093 = ~n19091 & ~n19092;
  assign n19094 = n18916 & n19093;
  assign n19095 = ~n18916 & ~n19093;
  assign n19096 = ~n19094 & ~n19095;
  assign n19097 = n18915 & ~n19096;
  assign n19098 = ~n18915 & n19096;
  assign n19099 = ~n19097 & ~n19098;
  assign n19100 = ~n18841 & ~n18844;
  assign n19101 = pi119  & n3011;
  assign n19102 = pi120  & n2809;
  assign n19103 = pi121  & n2804;
  assign n19104 = n2802 & n10071;
  assign n19105 = ~n19102 & ~n19103;
  assign n19106 = ~n19101 & n19105;
  assign n19107 = ~n19104 & n19106;
  assign n19108 = pi29  & n19107;
  assign n19109 = ~pi29  & ~n19107;
  assign n19110 = ~n19108 & ~n19109;
  assign n19111 = ~n19100 & ~n19110;
  assign n19112 = n19100 & n19110;
  assign n19113 = ~n19111 & ~n19112;
  assign n19114 = n19099 & n19113;
  assign n19115 = ~n19099 & ~n19113;
  assign n19116 = ~n19114 & ~n19115;
  assign n19117 = n18901 & n19116;
  assign n19118 = ~n18901 & ~n19116;
  assign n19119 = ~n19117 & ~n19118;
  assign n19120 = ~n18861 & ~n18864;
  assign n19121 = pi125  & n2053;
  assign n19122 = pi126  & n1893;
  assign n19123 = pi127  & n1888;
  assign n19124 = n1886 & n12519;
  assign n19125 = ~n19122 & ~n19123;
  assign n19126 = ~n19121 & n19125;
  assign n19127 = ~n19124 & n19126;
  assign n19128 = pi23  & n19127;
  assign n19129 = ~pi23  & ~n19127;
  assign n19130 = ~n19128 & ~n19129;
  assign n19131 = ~n19120 & ~n19130;
  assign n19132 = n19120 & n19130;
  assign n19133 = ~n19131 & ~n19132;
  assign n19134 = n19119 & n19133;
  assign n19135 = ~n19119 & ~n19133;
  assign n19136 = ~n19134 & ~n19135;
  assign n19137 = n18887 & ~n19136;
  assign n19138 = ~n18887 & n19136;
  assign n19139 = ~n19137 & ~n19138;
  assign n19140 = ~n18881 & ~n18884;
  assign n19141 = n19139 & ~n19140;
  assign n19142 = ~n19139 & n19140;
  assign po84  = ~n19141 & ~n19142;
  assign n19144 = ~n18900 & ~n19117;
  assign n19145 = pi126  & n2053;
  assign n19146 = pi127  & n1893;
  assign n19147 = n1886 & n12542;
  assign n19148 = ~n19145 & ~n19146;
  assign n19149 = ~n19147 & n19148;
  assign n19150 = pi23  & n19149;
  assign n19151 = ~pi23  & ~n19149;
  assign n19152 = ~n19150 & ~n19151;
  assign n19153 = ~n19144 & ~n19152;
  assign n19154 = n19144 & n19152;
  assign n19155 = ~n19153 & ~n19154;
  assign n19156 = pi123  & n2510;
  assign n19157 = pi124  & n2342;
  assign n19158 = pi125  & n2337;
  assign n19159 = n2335 & n11786;
  assign n19160 = ~n19157 & ~n19158;
  assign n19161 = ~n19156 & n19160;
  assign n19162 = ~n19159 & n19161;
  assign n19163 = pi26  & n19162;
  assign n19164 = ~pi26  & ~n19162;
  assign n19165 = ~n19163 & ~n19164;
  assign n19166 = ~n19111 & ~n19114;
  assign n19167 = n19165 & n19166;
  assign n19168 = ~n19165 & ~n19166;
  assign n19169 = ~n19167 & ~n19168;
  assign n19170 = ~n18914 & ~n19097;
  assign n19171 = pi120  & n3011;
  assign n19172 = pi121  & n2809;
  assign n19173 = pi122  & n2804;
  assign n19174 = n2802 & n10729;
  assign n19175 = ~n19172 & ~n19173;
  assign n19176 = ~n19171 & n19175;
  assign n19177 = ~n19174 & n19176;
  assign n19178 = pi29  & n19177;
  assign n19179 = ~pi29  & ~n19177;
  assign n19180 = ~n19178 & ~n19179;
  assign n19181 = ~n19170 & ~n19180;
  assign n19182 = n19170 & n19180;
  assign n19183 = ~n19181 & ~n19182;
  assign n19184 = pi117  & n3553;
  assign n19185 = pi118  & n3334;
  assign n19186 = pi119  & n3329;
  assign n19187 = n3327 & n9412;
  assign n19188 = ~n19185 & ~n19186;
  assign n19189 = ~n19184 & n19188;
  assign n19190 = ~n19187 & n19189;
  assign n19191 = pi32  & n19190;
  assign n19192 = ~pi32  & ~n19190;
  assign n19193 = ~n19191 & ~n19192;
  assign n19194 = n18916 & ~n19091;
  assign n19195 = ~n19092 & ~n19194;
  assign n19196 = ~n19193 & n19195;
  assign n19197 = n19193 & ~n19195;
  assign n19198 = ~n19196 & ~n19197;
  assign n19199 = ~n19073 & ~n19079;
  assign n19200 = ~n19057 & ~n19061;
  assign n19201 = ~n19041 & ~n19045;
  assign n19202 = ~n19025 & ~n19029;
  assign n19203 = pi102  & n7121;
  assign n19204 = pi103  & n6795;
  assign n19205 = pi104  & n6790;
  assign n19206 = n5212 & n6788;
  assign n19207 = ~n19204 & ~n19205;
  assign n19208 = ~n19203 & n19207;
  assign n19209 = ~n19206 & n19208;
  assign n19210 = pi47  & n19209;
  assign n19211 = ~pi47  & ~n19209;
  assign n19212 = ~n19210 & ~n19211;
  assign n19213 = ~n19009 & ~n19013;
  assign n19214 = ~n19003 & ~n19006;
  assign n19215 = ~n18986 & ~n18990;
  assign n19216 = ~n18970 & ~n18974;
  assign n19217 = pi90  & n10886;
  assign n19218 = pi91  & n10495;
  assign n19219 = pi92  & n10490;
  assign n19220 = n2924 & n10488;
  assign n19221 = ~n19218 & ~n19219;
  assign n19222 = ~n19217 & n19221;
  assign n19223 = ~n19220 & n19222;
  assign n19224 = pi59  & n19223;
  assign n19225 = ~pi59  & ~n19223;
  assign n19226 = ~n19224 & ~n19225;
  assign n19227 = ~n18964 & ~n18967;
  assign n19228 = ~n18948 & ~n18951;
  assign n19229 = pi86  & n12277;
  assign n19230 = pi85  & n12276;
  assign n19231 = ~n19229 & ~n19230;
  assign n19232 = n19228 & ~n19231;
  assign n19233 = ~n19228 & n19231;
  assign n19234 = ~n19232 & ~n19233;
  assign n19235 = pi87  & n11910;
  assign n19236 = pi88  & n11529;
  assign n19237 = pi89  & n11524;
  assign n19238 = n2287 & n11522;
  assign n19239 = ~n19236 & ~n19237;
  assign n19240 = ~n19235 & n19239;
  assign n19241 = ~n19238 & n19240;
  assign n19242 = pi62  & n19241;
  assign n19243 = ~pi62  & ~n19241;
  assign n19244 = ~n19242 & ~n19243;
  assign n19245 = n19234 & ~n19244;
  assign n19246 = ~n19234 & n19244;
  assign n19247 = ~n19245 & ~n19246;
  assign n19248 = ~n19227 & n19247;
  assign n19249 = n19227 & ~n19247;
  assign n19250 = ~n19248 & ~n19249;
  assign n19251 = ~n19226 & n19250;
  assign n19252 = n19226 & ~n19250;
  assign n19253 = ~n19251 & ~n19252;
  assign n19254 = ~n19216 & n19253;
  assign n19255 = n19216 & ~n19253;
  assign n19256 = ~n19254 & ~n19255;
  assign n19257 = pi93  & n9858;
  assign n19258 = pi94  & n9508;
  assign n19259 = pi95  & n9503;
  assign n19260 = n3475 & n9501;
  assign n19261 = ~n19258 & ~n19259;
  assign n19262 = ~n19257 & n19261;
  assign n19263 = ~n19260 & n19262;
  assign n19264 = pi56  & n19263;
  assign n19265 = ~pi56  & ~n19263;
  assign n19266 = ~n19264 & ~n19265;
  assign n19267 = n19256 & ~n19266;
  assign n19268 = ~n19256 & n19266;
  assign n19269 = ~n19267 & ~n19268;
  assign n19270 = n19215 & ~n19269;
  assign n19271 = ~n19215 & n19269;
  assign n19272 = ~n19270 & ~n19271;
  assign n19273 = pi96  & n8905;
  assign n19274 = pi97  & n8535;
  assign n19275 = pi98  & n8530;
  assign n19276 = n3889 & n8528;
  assign n19277 = ~n19274 & ~n19275;
  assign n19278 = ~n19273 & n19277;
  assign n19279 = ~n19276 & n19278;
  assign n19280 = pi53  & n19279;
  assign n19281 = ~pi53  & ~n19279;
  assign n19282 = ~n19280 & ~n19281;
  assign n19283 = n19272 & ~n19282;
  assign n19284 = ~n19272 & n19282;
  assign n19285 = ~n19283 & ~n19284;
  assign n19286 = n19214 & ~n19285;
  assign n19287 = ~n19214 & n19285;
  assign n19288 = ~n19286 & ~n19287;
  assign n19289 = pi99  & n7969;
  assign n19290 = pi100  & n7636;
  assign n19291 = pi101  & n7631;
  assign n19292 = n4730 & n7629;
  assign n19293 = ~n19290 & ~n19291;
  assign n19294 = ~n19289 & n19293;
  assign n19295 = ~n19292 & n19294;
  assign n19296 = pi50  & n19295;
  assign n19297 = ~pi50  & ~n19295;
  assign n19298 = ~n19296 & ~n19297;
  assign n19299 = ~n19288 & n19298;
  assign n19300 = n19288 & ~n19298;
  assign n19301 = ~n19299 & ~n19300;
  assign n19302 = ~n19213 & n19301;
  assign n19303 = n19213 & ~n19301;
  assign n19304 = ~n19302 & ~n19303;
  assign n19305 = ~n19212 & n19304;
  assign n19306 = n19212 & ~n19304;
  assign n19307 = ~n19305 & ~n19306;
  assign n19308 = ~n19202 & n19307;
  assign n19309 = n19202 & ~n19307;
  assign n19310 = ~n19308 & ~n19309;
  assign n19311 = pi105  & n6331;
  assign n19312 = pi106  & n6015;
  assign n19313 = pi107  & n6010;
  assign n19314 = n6008 & n6189;
  assign n19315 = ~n19312 & ~n19313;
  assign n19316 = ~n19311 & n19315;
  assign n19317 = ~n19314 & n19316;
  assign n19318 = pi44  & n19317;
  assign n19319 = ~pi44  & ~n19317;
  assign n19320 = ~n19318 & ~n19319;
  assign n19321 = n19310 & ~n19320;
  assign n19322 = ~n19310 & n19320;
  assign n19323 = ~n19321 & ~n19322;
  assign n19324 = n19201 & ~n19323;
  assign n19325 = ~n19201 & n19323;
  assign n19326 = ~n19324 & ~n19325;
  assign n19327 = pi108  & n5558;
  assign n19328 = pi109  & n5293;
  assign n19329 = pi110  & n5288;
  assign n19330 = n5286 & n6995;
  assign n19331 = ~n19328 & ~n19329;
  assign n19332 = ~n19327 & n19331;
  assign n19333 = ~n19330 & n19332;
  assign n19334 = pi41  & n19333;
  assign n19335 = ~pi41  & ~n19333;
  assign n19336 = ~n19334 & ~n19335;
  assign n19337 = n19326 & ~n19336;
  assign n19338 = ~n19326 & n19336;
  assign n19339 = ~n19337 & ~n19338;
  assign n19340 = n19200 & ~n19339;
  assign n19341 = ~n19200 & n19339;
  assign n19342 = ~n19340 & ~n19341;
  assign n19343 = pi111  & n4843;
  assign n19344 = pi112  & n4598;
  assign n19345 = pi113  & n4593;
  assign n19346 = n4591 & n7852;
  assign n19347 = ~n19344 & ~n19345;
  assign n19348 = ~n19343 & n19347;
  assign n19349 = ~n19346 & n19348;
  assign n19350 = pi38  & n19349;
  assign n19351 = ~pi38  & ~n19349;
  assign n19352 = ~n19350 & ~n19351;
  assign n19353 = n19342 & ~n19352;
  assign n19354 = ~n19342 & n19352;
  assign n19355 = ~n19353 & ~n19354;
  assign n19356 = n19199 & ~n19355;
  assign n19357 = ~n19199 & n19355;
  assign n19358 = ~n19356 & ~n19357;
  assign n19359 = pi114  & n4176;
  assign n19360 = pi115  & n3938;
  assign n19361 = pi116  & n3933;
  assign n19362 = n3931 & n8470;
  assign n19363 = ~n19360 & ~n19361;
  assign n19364 = ~n19359 & n19363;
  assign n19365 = ~n19362 & n19364;
  assign n19366 = pi35  & n19365;
  assign n19367 = ~pi35  & ~n19365;
  assign n19368 = ~n19366 & ~n19367;
  assign n19369 = n19358 & ~n19368;
  assign n19370 = ~n19358 & n19368;
  assign n19371 = ~n19369 & ~n19370;
  assign n19372 = n19198 & n19371;
  assign n19373 = ~n19198 & ~n19371;
  assign n19374 = ~n19372 & ~n19373;
  assign n19375 = n19183 & n19374;
  assign n19376 = ~n19183 & ~n19374;
  assign n19377 = ~n19375 & ~n19376;
  assign n19378 = n19169 & n19377;
  assign n19379 = ~n19169 & ~n19377;
  assign n19380 = ~n19378 & ~n19379;
  assign n19381 = n19155 & ~n19380;
  assign n19382 = ~n19155 & n19380;
  assign n19383 = ~n19381 & ~n19382;
  assign n19384 = ~n19131 & ~n19134;
  assign n19385 = n19383 & n19384;
  assign n19386 = ~n19383 & ~n19384;
  assign n19387 = ~n19385 & ~n19386;
  assign n19388 = ~n19138 & ~n19141;
  assign n19389 = n19387 & ~n19388;
  assign n19390 = ~n19387 & n19388;
  assign po85  = ~n19389 & ~n19390;
  assign n19392 = ~n19386 & ~n19389;
  assign n19393 = ~n19168 & ~n19378;
  assign n19394 = n1886 & ~n12539;
  assign n19395 = ~n2053 & ~n19394;
  assign n19396 = pi127  & ~n19395;
  assign n19397 = pi23  & ~n19396;
  assign n19398 = ~pi23  & n19396;
  assign n19399 = ~n19397 & ~n19398;
  assign n19400 = ~n19393 & ~n19399;
  assign n19401 = n19393 & n19399;
  assign n19402 = ~n19400 & ~n19401;
  assign n19403 = pi124  & n2510;
  assign n19404 = pi125  & n2342;
  assign n19405 = pi126  & n2337;
  assign n19406 = n2335 & n12148;
  assign n19407 = ~n19404 & ~n19405;
  assign n19408 = ~n19403 & n19407;
  assign n19409 = ~n19406 & n19408;
  assign n19410 = pi26  & n19409;
  assign n19411 = ~pi26  & ~n19409;
  assign n19412 = ~n19410 & ~n19411;
  assign n19413 = ~n19181 & ~n19375;
  assign n19414 = n19412 & n19413;
  assign n19415 = ~n19412 & ~n19413;
  assign n19416 = ~n19414 & ~n19415;
  assign n19417 = pi121  & n3011;
  assign n19418 = pi122  & n2809;
  assign n19419 = pi123  & n2804;
  assign n19420 = n2802 & n10754;
  assign n19421 = ~n19418 & ~n19419;
  assign n19422 = ~n19417 & n19421;
  assign n19423 = ~n19420 & n19422;
  assign n19424 = pi29  & n19423;
  assign n19425 = ~pi29  & ~n19423;
  assign n19426 = ~n19424 & ~n19425;
  assign n19427 = ~n19196 & ~n19372;
  assign n19428 = ~n19426 & ~n19427;
  assign n19429 = n19426 & n19427;
  assign n19430 = ~n19428 & ~n19429;
  assign n19431 = pi118  & n3553;
  assign n19432 = pi119  & n3334;
  assign n19433 = pi120  & n3329;
  assign n19434 = n3327 & n10047;
  assign n19435 = ~n19432 & ~n19433;
  assign n19436 = ~n19431 & n19435;
  assign n19437 = ~n19434 & n19436;
  assign n19438 = pi32  & n19437;
  assign n19439 = ~pi32  & ~n19437;
  assign n19440 = ~n19438 & ~n19439;
  assign n19441 = ~n19357 & n19368;
  assign n19442 = ~n19356 & ~n19441;
  assign n19443 = n19440 & ~n19442;
  assign n19444 = ~n19440 & n19442;
  assign n19445 = ~n19443 & ~n19444;
  assign n19446 = pi115  & n4176;
  assign n19447 = pi116  & n3938;
  assign n19448 = pi117  & n3933;
  assign n19449 = n3931 & n8784;
  assign n19450 = ~n19447 & ~n19448;
  assign n19451 = ~n19446 & n19450;
  assign n19452 = ~n19449 & n19451;
  assign n19453 = pi35  & n19452;
  assign n19454 = ~pi35  & ~n19452;
  assign n19455 = ~n19453 & ~n19454;
  assign n19456 = pi106  & n6331;
  assign n19457 = pi107  & n6015;
  assign n19458 = pi108  & n6010;
  assign n19459 = n6008 & n6213;
  assign n19460 = ~n19457 & ~n19458;
  assign n19461 = ~n19456 & n19460;
  assign n19462 = ~n19459 & n19461;
  assign n19463 = pi44  & n19462;
  assign n19464 = ~pi44  & ~n19462;
  assign n19465 = ~n19463 & ~n19464;
  assign n19466 = ~n19302 & ~n19305;
  assign n19467 = pi103  & n7121;
  assign n19468 = pi104  & n6795;
  assign n19469 = pi105  & n6790;
  assign n19470 = n5677 & n6788;
  assign n19471 = ~n19468 & ~n19469;
  assign n19472 = ~n19467 & n19471;
  assign n19473 = ~n19470 & n19472;
  assign n19474 = pi47  & n19473;
  assign n19475 = ~pi47  & ~n19473;
  assign n19476 = ~n19474 & ~n19475;
  assign n19477 = ~n19287 & ~n19300;
  assign n19478 = pi97  & n8905;
  assign n19479 = pi98  & n8535;
  assign n19480 = pi99  & n8530;
  assign n19481 = n4101 & n8528;
  assign n19482 = ~n19479 & ~n19480;
  assign n19483 = ~n19478 & n19482;
  assign n19484 = ~n19481 & n19483;
  assign n19485 = pi53  & n19484;
  assign n19486 = ~pi53  & ~n19484;
  assign n19487 = ~n19485 & ~n19486;
  assign n19488 = ~n19248 & ~n19251;
  assign n19489 = ~n19233 & ~n19245;
  assign n19490 = pi87  & n12277;
  assign n19491 = pi86  & n12276;
  assign n19492 = ~n19490 & ~n19491;
  assign n19493 = ~n19231 & n19492;
  assign n19494 = n19231 & ~n19492;
  assign n19495 = ~n19493 & ~n19494;
  assign n19496 = pi88  & n11910;
  assign n19497 = pi89  & n11529;
  assign n19498 = pi90  & n11524;
  assign n19499 = n2448 & n11522;
  assign n19500 = ~n19497 & ~n19498;
  assign n19501 = ~n19496 & n19500;
  assign n19502 = ~n19499 & n19501;
  assign n19503 = pi62  & n19502;
  assign n19504 = ~pi62  & ~n19502;
  assign n19505 = ~n19503 & ~n19504;
  assign n19506 = n19495 & ~n19505;
  assign n19507 = ~n19495 & n19505;
  assign n19508 = ~n19506 & ~n19507;
  assign n19509 = ~n19489 & n19508;
  assign n19510 = n19489 & ~n19508;
  assign n19511 = ~n19509 & ~n19510;
  assign n19512 = pi91  & n10886;
  assign n19513 = pi92  & n10495;
  assign n19514 = pi93  & n10490;
  assign n19515 = n2948 & n10488;
  assign n19516 = ~n19513 & ~n19514;
  assign n19517 = ~n19512 & n19516;
  assign n19518 = ~n19515 & n19517;
  assign n19519 = pi59  & n19518;
  assign n19520 = ~pi59  & ~n19518;
  assign n19521 = ~n19519 & ~n19520;
  assign n19522 = n19511 & ~n19521;
  assign n19523 = ~n19511 & n19521;
  assign n19524 = ~n19522 & ~n19523;
  assign n19525 = n19488 & ~n19524;
  assign n19526 = ~n19488 & n19524;
  assign n19527 = ~n19525 & ~n19526;
  assign n19528 = pi94  & n9858;
  assign n19529 = pi95  & n9508;
  assign n19530 = pi96  & n9503;
  assign n19531 = n3499 & n9501;
  assign n19532 = ~n19529 & ~n19530;
  assign n19533 = ~n19528 & n19532;
  assign n19534 = ~n19531 & n19533;
  assign n19535 = pi56  & n19534;
  assign n19536 = ~pi56  & ~n19534;
  assign n19537 = ~n19535 & ~n19536;
  assign n19538 = ~n19527 & n19537;
  assign n19539 = n19527 & ~n19537;
  assign n19540 = ~n19538 & ~n19539;
  assign n19541 = ~n19254 & n19266;
  assign n19542 = ~n19255 & ~n19541;
  assign n19543 = n19540 & n19542;
  assign n19544 = ~n19540 & ~n19542;
  assign n19545 = ~n19543 & ~n19544;
  assign n19546 = ~n19487 & n19545;
  assign n19547 = n19487 & ~n19545;
  assign n19548 = ~n19546 & ~n19547;
  assign n19549 = ~n19271 & n19282;
  assign n19550 = ~n19270 & ~n19549;
  assign n19551 = n19548 & n19550;
  assign n19552 = ~n19548 & ~n19550;
  assign n19553 = ~n19551 & ~n19552;
  assign n19554 = pi100  & n7969;
  assign n19555 = pi101  & n7636;
  assign n19556 = pi102  & n7631;
  assign n19557 = n4956 & n7629;
  assign n19558 = ~n19555 & ~n19556;
  assign n19559 = ~n19554 & n19558;
  assign n19560 = ~n19557 & n19559;
  assign n19561 = pi50  & n19560;
  assign n19562 = ~pi50  & ~n19560;
  assign n19563 = ~n19561 & ~n19562;
  assign n19564 = n19553 & ~n19563;
  assign n19565 = ~n19553 & n19563;
  assign n19566 = ~n19564 & ~n19565;
  assign n19567 = ~n19477 & n19566;
  assign n19568 = n19477 & ~n19566;
  assign n19569 = ~n19567 & ~n19568;
  assign n19570 = ~n19476 & n19569;
  assign n19571 = n19476 & ~n19569;
  assign n19572 = ~n19570 & ~n19571;
  assign n19573 = ~n19466 & n19572;
  assign n19574 = n19466 & ~n19572;
  assign n19575 = ~n19573 & ~n19574;
  assign n19576 = ~n19465 & n19575;
  assign n19577 = n19465 & ~n19575;
  assign n19578 = ~n19576 & ~n19577;
  assign n19579 = ~n19308 & n19320;
  assign n19580 = ~n19309 & ~n19579;
  assign n19581 = n19578 & n19580;
  assign n19582 = ~n19578 & ~n19580;
  assign n19583 = ~n19581 & ~n19582;
  assign n19584 = pi109  & n5558;
  assign n19585 = pi110  & n5293;
  assign n19586 = pi111  & n5288;
  assign n19587 = n5286 & n7272;
  assign n19588 = ~n19585 & ~n19586;
  assign n19589 = ~n19584 & n19588;
  assign n19590 = ~n19587 & n19589;
  assign n19591 = pi41  & n19590;
  assign n19592 = ~pi41  & ~n19590;
  assign n19593 = ~n19591 & ~n19592;
  assign n19594 = n19583 & ~n19593;
  assign n19595 = ~n19583 & n19593;
  assign n19596 = ~n19594 & ~n19595;
  assign n19597 = ~n19325 & n19336;
  assign n19598 = ~n19324 & ~n19597;
  assign n19599 = ~n19596 & ~n19598;
  assign n19600 = n19596 & n19598;
  assign n19601 = ~n19599 & ~n19600;
  assign n19602 = pi112  & n4843;
  assign n19603 = pi113  & n4598;
  assign n19604 = pi114  & n4593;
  assign n19605 = n4591 & n8146;
  assign n19606 = ~n19603 & ~n19604;
  assign n19607 = ~n19602 & n19606;
  assign n19608 = ~n19605 & n19607;
  assign n19609 = pi38  & n19608;
  assign n19610 = ~pi38  & ~n19608;
  assign n19611 = ~n19609 & ~n19610;
  assign n19612 = ~n19601 & n19611;
  assign n19613 = n19601 & ~n19611;
  assign n19614 = ~n19612 & ~n19613;
  assign n19615 = ~n19341 & n19352;
  assign n19616 = ~n19340 & ~n19615;
  assign n19617 = n19614 & n19616;
  assign n19618 = ~n19614 & ~n19616;
  assign n19619 = ~n19617 & ~n19618;
  assign n19620 = n19455 & ~n19619;
  assign n19621 = ~n19455 & n19619;
  assign n19622 = ~n19620 & ~n19621;
  assign n19623 = n19445 & n19622;
  assign n19624 = ~n19445 & ~n19622;
  assign n19625 = ~n19623 & ~n19624;
  assign n19626 = n19430 & n19625;
  assign n19627 = ~n19430 & ~n19625;
  assign n19628 = ~n19626 & ~n19627;
  assign n19629 = n19416 & n19628;
  assign n19630 = ~n19416 & ~n19628;
  assign n19631 = ~n19629 & ~n19630;
  assign n19632 = n19402 & n19631;
  assign n19633 = ~n19402 & ~n19631;
  assign n19634 = ~n19632 & ~n19633;
  assign n19635 = ~n19153 & ~n19380;
  assign n19636 = ~n19154 & ~n19635;
  assign n19637 = n19634 & n19636;
  assign n19638 = ~n19634 & ~n19636;
  assign n19639 = ~n19637 & ~n19638;
  assign n19640 = ~n19392 & n19639;
  assign n19641 = n19392 & ~n19639;
  assign po86  = ~n19640 & ~n19641;
  assign n19643 = ~n19637 & ~n19640;
  assign n19644 = ~n19400 & ~n19632;
  assign n19645 = ~n19428 & ~n19626;
  assign n19646 = pi122  & n3011;
  assign n19647 = pi123  & n2809;
  assign n19648 = pi124  & n2804;
  assign n19649 = n2802 & n11099;
  assign n19650 = ~n19647 & ~n19648;
  assign n19651 = ~n19646 & n19650;
  assign n19652 = ~n19649 & n19651;
  assign n19653 = pi29  & n19652;
  assign n19654 = ~pi29  & ~n19652;
  assign n19655 = ~n19653 & ~n19654;
  assign n19656 = ~n19645 & ~n19655;
  assign n19657 = n19645 & n19655;
  assign n19658 = ~n19656 & ~n19657;
  assign n19659 = pi119  & n3553;
  assign n19660 = pi120  & n3334;
  assign n19661 = pi121  & n3329;
  assign n19662 = n3327 & n10071;
  assign n19663 = ~n19660 & ~n19661;
  assign n19664 = ~n19659 & n19663;
  assign n19665 = ~n19662 & n19664;
  assign n19666 = pi32  & n19665;
  assign n19667 = ~pi32  & ~n19665;
  assign n19668 = ~n19666 & ~n19667;
  assign n19669 = ~n19444 & ~n19622;
  assign n19670 = ~n19443 & ~n19669;
  assign n19671 = n19668 & ~n19670;
  assign n19672 = ~n19668 & n19670;
  assign n19673 = ~n19671 & ~n19672;
  assign n19674 = pi116  & n4176;
  assign n19675 = pi117  & n3938;
  assign n19676 = pi118  & n3933;
  assign n19677 = n3931 & n9095;
  assign n19678 = ~n19675 & ~n19676;
  assign n19679 = ~n19674 & n19678;
  assign n19680 = ~n19677 & n19679;
  assign n19681 = pi35  & n19680;
  assign n19682 = ~pi35  & ~n19680;
  assign n19683 = ~n19681 & ~n19682;
  assign n19684 = ~n19600 & ~n19613;
  assign n19685 = ~n19573 & ~n19576;
  assign n19686 = pi107  & n6331;
  assign n19687 = pi108  & n6015;
  assign n19688 = pi109  & n6010;
  assign n19689 = n6008 & n6715;
  assign n19690 = ~n19687 & ~n19688;
  assign n19691 = ~n19686 & n19690;
  assign n19692 = ~n19689 & n19691;
  assign n19693 = pi44  & n19692;
  assign n19694 = ~pi44  & ~n19692;
  assign n19695 = ~n19693 & ~n19694;
  assign n19696 = ~n19567 & ~n19570;
  assign n19697 = ~n19543 & ~n19546;
  assign n19698 = pi92  & n10886;
  assign n19699 = pi93  & n10495;
  assign n19700 = pi94  & n10490;
  assign n19701 = n3280 & n10488;
  assign n19702 = ~n19699 & ~n19700;
  assign n19703 = ~n19698 & n19702;
  assign n19704 = ~n19701 & n19703;
  assign n19705 = pi59  & n19704;
  assign n19706 = ~pi59  & ~n19704;
  assign n19707 = ~n19705 & ~n19706;
  assign n19708 = ~n19493 & ~n19506;
  assign n19709 = pi88  & n12277;
  assign n19710 = pi87  & n12276;
  assign n19711 = ~n19709 & ~n19710;
  assign n19712 = ~pi23  & ~n19711;
  assign n19713 = pi23  & n19711;
  assign n19714 = ~n19712 & ~n19713;
  assign n19715 = ~n19492 & n19714;
  assign n19716 = n19492 & ~n19714;
  assign n19717 = ~n19715 & ~n19716;
  assign n19718 = pi89  & n11910;
  assign n19719 = pi90  & n11529;
  assign n19720 = pi91  & n11524;
  assign n19721 = n2746 & n11522;
  assign n19722 = ~n19719 & ~n19720;
  assign n19723 = ~n19718 & n19722;
  assign n19724 = ~n19721 & n19723;
  assign n19725 = pi62  & n19724;
  assign n19726 = ~pi62  & ~n19724;
  assign n19727 = ~n19725 & ~n19726;
  assign n19728 = n19717 & ~n19727;
  assign n19729 = ~n19717 & n19727;
  assign n19730 = ~n19728 & ~n19729;
  assign n19731 = ~n19708 & n19730;
  assign n19732 = n19708 & ~n19730;
  assign n19733 = ~n19731 & ~n19732;
  assign n19734 = ~n19707 & n19733;
  assign n19735 = n19707 & ~n19733;
  assign n19736 = ~n19734 & ~n19735;
  assign n19737 = ~n19509 & n19521;
  assign n19738 = ~n19510 & ~n19737;
  assign n19739 = ~n19736 & ~n19738;
  assign n19740 = n19736 & n19738;
  assign n19741 = ~n19739 & ~n19740;
  assign n19742 = pi95  & n9858;
  assign n19743 = pi96  & n9508;
  assign n19744 = pi97  & n9503;
  assign n19745 = n3691 & n9501;
  assign n19746 = ~n19743 & ~n19744;
  assign n19747 = ~n19742 & n19746;
  assign n19748 = ~n19745 & n19747;
  assign n19749 = pi56  & n19748;
  assign n19750 = ~pi56  & ~n19748;
  assign n19751 = ~n19749 & ~n19750;
  assign n19752 = ~n19526 & ~n19539;
  assign n19753 = ~n19751 & ~n19752;
  assign n19754 = n19751 & n19752;
  assign n19755 = ~n19753 & ~n19754;
  assign n19756 = n19741 & n19755;
  assign n19757 = ~n19741 & ~n19755;
  assign n19758 = ~n19756 & ~n19757;
  assign n19759 = pi98  & n8905;
  assign n19760 = pi99  & n8535;
  assign n19761 = pi100  & n8530;
  assign n19762 = n4501 & n8528;
  assign n19763 = ~n19760 & ~n19761;
  assign n19764 = ~n19759 & n19763;
  assign n19765 = ~n19762 & n19764;
  assign n19766 = pi53  & n19765;
  assign n19767 = ~pi53  & ~n19765;
  assign n19768 = ~n19766 & ~n19767;
  assign n19769 = n19758 & ~n19768;
  assign n19770 = ~n19758 & n19768;
  assign n19771 = ~n19769 & ~n19770;
  assign n19772 = n19697 & ~n19771;
  assign n19773 = ~n19697 & n19771;
  assign n19774 = ~n19772 & ~n19773;
  assign n19775 = pi101  & n7969;
  assign n19776 = pi102  & n7636;
  assign n19777 = pi103  & n7631;
  assign n19778 = n5188 & n7629;
  assign n19779 = ~n19776 & ~n19777;
  assign n19780 = ~n19775 & n19779;
  assign n19781 = ~n19778 & n19780;
  assign n19782 = pi50  & n19781;
  assign n19783 = ~pi50  & ~n19781;
  assign n19784 = ~n19782 & ~n19783;
  assign n19785 = n19774 & ~n19784;
  assign n19786 = ~n19774 & n19784;
  assign n19787 = ~n19785 & ~n19786;
  assign n19788 = ~n19551 & n19563;
  assign n19789 = ~n19552 & ~n19788;
  assign n19790 = ~n19787 & ~n19789;
  assign n19791 = n19787 & n19789;
  assign n19792 = ~n19790 & ~n19791;
  assign n19793 = pi104  & n7121;
  assign n19794 = pi105  & n6795;
  assign n19795 = pi106  & n6790;
  assign n19796 = n5701 & n6788;
  assign n19797 = ~n19794 & ~n19795;
  assign n19798 = ~n19793 & n19797;
  assign n19799 = ~n19796 & n19798;
  assign n19800 = pi47  & n19799;
  assign n19801 = ~pi47  & ~n19799;
  assign n19802 = ~n19800 & ~n19801;
  assign n19803 = n19792 & ~n19802;
  assign n19804 = ~n19792 & n19802;
  assign n19805 = ~n19803 & ~n19804;
  assign n19806 = ~n19696 & n19805;
  assign n19807 = n19696 & ~n19805;
  assign n19808 = ~n19806 & ~n19807;
  assign n19809 = ~n19695 & n19808;
  assign n19810 = n19695 & ~n19808;
  assign n19811 = ~n19809 & ~n19810;
  assign n19812 = n19685 & ~n19811;
  assign n19813 = ~n19685 & n19811;
  assign n19814 = ~n19812 & ~n19813;
  assign n19815 = pi110  & n5558;
  assign n19816 = pi111  & n5293;
  assign n19817 = pi112  & n5288;
  assign n19818 = n5286 & n7296;
  assign n19819 = ~n19816 & ~n19817;
  assign n19820 = ~n19815 & n19819;
  assign n19821 = ~n19818 & n19820;
  assign n19822 = pi41  & n19821;
  assign n19823 = ~pi41  & ~n19821;
  assign n19824 = ~n19822 & ~n19823;
  assign n19825 = n19814 & ~n19824;
  assign n19826 = ~n19814 & n19824;
  assign n19827 = ~n19825 & ~n19826;
  assign n19828 = ~n19581 & n19593;
  assign n19829 = ~n19582 & ~n19828;
  assign n19830 = ~n19827 & ~n19829;
  assign n19831 = n19827 & n19829;
  assign n19832 = ~n19830 & ~n19831;
  assign n19833 = pi113  & n4843;
  assign n19834 = pi114  & n4598;
  assign n19835 = pi115  & n4593;
  assign n19836 = n4591 & n8170;
  assign n19837 = ~n19834 & ~n19835;
  assign n19838 = ~n19833 & n19837;
  assign n19839 = ~n19836 & n19838;
  assign n19840 = pi38  & n19839;
  assign n19841 = ~pi38  & ~n19839;
  assign n19842 = ~n19840 & ~n19841;
  assign n19843 = n19832 & ~n19842;
  assign n19844 = ~n19832 & n19842;
  assign n19845 = ~n19843 & ~n19844;
  assign n19846 = n19684 & n19845;
  assign n19847 = ~n19684 & ~n19845;
  assign n19848 = ~n19846 & ~n19847;
  assign n19849 = n19683 & n19848;
  assign n19850 = ~n19683 & ~n19848;
  assign n19851 = ~n19849 & ~n19850;
  assign n19852 = n19455 & ~n19617;
  assign n19853 = ~n19618 & ~n19852;
  assign n19854 = n19851 & n19853;
  assign n19855 = ~n19851 & ~n19853;
  assign n19856 = ~n19854 & ~n19855;
  assign n19857 = n19673 & n19856;
  assign n19858 = ~n19673 & ~n19856;
  assign n19859 = ~n19857 & ~n19858;
  assign n19860 = n19658 & n19859;
  assign n19861 = ~n19658 & ~n19859;
  assign n19862 = ~n19860 & ~n19861;
  assign n19863 = ~n19415 & ~n19629;
  assign n19864 = pi125  & n2510;
  assign n19865 = pi126  & n2342;
  assign n19866 = pi127  & n2337;
  assign n19867 = n2335 & n12519;
  assign n19868 = ~n19865 & ~n19866;
  assign n19869 = ~n19864 & n19868;
  assign n19870 = ~n19867 & n19869;
  assign n19871 = pi26  & n19870;
  assign n19872 = ~pi26  & ~n19870;
  assign n19873 = ~n19871 & ~n19872;
  assign n19874 = ~n19863 & ~n19873;
  assign n19875 = n19863 & n19873;
  assign n19876 = ~n19874 & ~n19875;
  assign n19877 = n19862 & n19876;
  assign n19878 = ~n19862 & ~n19876;
  assign n19879 = ~n19877 & ~n19878;
  assign n19880 = ~n19644 & n19879;
  assign n19881 = n19644 & ~n19879;
  assign n19882 = ~n19880 & ~n19881;
  assign n19883 = ~n19643 & n19882;
  assign n19884 = n19643 & ~n19882;
  assign po87  = ~n19883 & ~n19884;
  assign n19886 = ~n19880 & ~n19883;
  assign n19887 = ~n19874 & ~n19877;
  assign n19888 = ~n19850 & ~n19854;
  assign n19889 = pi120  & n3553;
  assign n19890 = pi121  & n3334;
  assign n19891 = pi122  & n3329;
  assign n19892 = n3327 & n10729;
  assign n19893 = ~n19890 & ~n19891;
  assign n19894 = ~n19889 & n19893;
  assign n19895 = ~n19892 & n19894;
  assign n19896 = pi32  & n19895;
  assign n19897 = ~pi32  & ~n19895;
  assign n19898 = ~n19896 & ~n19897;
  assign n19899 = ~n19888 & ~n19898;
  assign n19900 = n19888 & n19898;
  assign n19901 = ~n19899 & ~n19900;
  assign n19902 = pi117  & n4176;
  assign n19903 = pi118  & n3938;
  assign n19904 = pi119  & n3933;
  assign n19905 = n3931 & n9412;
  assign n19906 = ~n19903 & ~n19904;
  assign n19907 = ~n19902 & n19906;
  assign n19908 = ~n19905 & n19907;
  assign n19909 = pi35  & n19908;
  assign n19910 = ~pi35  & ~n19908;
  assign n19911 = ~n19909 & ~n19910;
  assign n19912 = ~n19825 & ~n19831;
  assign n19913 = ~n19809 & ~n19813;
  assign n19914 = ~n19803 & ~n19806;
  assign n19915 = ~n19785 & ~n19791;
  assign n19916 = pi102  & n7969;
  assign n19917 = pi103  & n7636;
  assign n19918 = pi104  & n7631;
  assign n19919 = n5212 & n7629;
  assign n19920 = ~n19917 & ~n19918;
  assign n19921 = ~n19916 & n19920;
  assign n19922 = ~n19919 & n19921;
  assign n19923 = pi50  & n19922;
  assign n19924 = ~pi50  & ~n19922;
  assign n19925 = ~n19923 & ~n19924;
  assign n19926 = ~n19769 & ~n19773;
  assign n19927 = ~n19753 & ~n19756;
  assign n19928 = ~n19734 & ~n19740;
  assign n19929 = ~n19728 & ~n19731;
  assign n19930 = ~n19712 & ~n19715;
  assign n19931 = pi89  & n12277;
  assign n19932 = pi88  & n12276;
  assign n19933 = ~n19931 & ~n19932;
  assign n19934 = n19930 & ~n19933;
  assign n19935 = ~n19930 & n19933;
  assign n19936 = ~n19934 & ~n19935;
  assign n19937 = pi90  & n11910;
  assign n19938 = pi91  & n11529;
  assign n19939 = pi92  & n11524;
  assign n19940 = n2924 & n11522;
  assign n19941 = ~n19938 & ~n19939;
  assign n19942 = ~n19937 & n19941;
  assign n19943 = ~n19940 & n19942;
  assign n19944 = pi62  & n19943;
  assign n19945 = ~pi62  & ~n19943;
  assign n19946 = ~n19944 & ~n19945;
  assign n19947 = n19936 & ~n19946;
  assign n19948 = ~n19936 & n19946;
  assign n19949 = ~n19947 & ~n19948;
  assign n19950 = ~n19929 & n19949;
  assign n19951 = n19929 & ~n19949;
  assign n19952 = ~n19950 & ~n19951;
  assign n19953 = pi93  & n10886;
  assign n19954 = pi94  & n10495;
  assign n19955 = pi95  & n10490;
  assign n19956 = n3475 & n10488;
  assign n19957 = ~n19954 & ~n19955;
  assign n19958 = ~n19953 & n19957;
  assign n19959 = ~n19956 & n19958;
  assign n19960 = pi59  & n19959;
  assign n19961 = ~pi59  & ~n19959;
  assign n19962 = ~n19960 & ~n19961;
  assign n19963 = n19952 & ~n19962;
  assign n19964 = ~n19952 & n19962;
  assign n19965 = ~n19963 & ~n19964;
  assign n19966 = n19928 & ~n19965;
  assign n19967 = ~n19928 & n19965;
  assign n19968 = ~n19966 & ~n19967;
  assign n19969 = pi96  & n9858;
  assign n19970 = pi97  & n9508;
  assign n19971 = pi98  & n9503;
  assign n19972 = n3889 & n9501;
  assign n19973 = ~n19970 & ~n19971;
  assign n19974 = ~n19969 & n19973;
  assign n19975 = ~n19972 & n19974;
  assign n19976 = pi56  & n19975;
  assign n19977 = ~pi56  & ~n19975;
  assign n19978 = ~n19976 & ~n19977;
  assign n19979 = n19968 & ~n19978;
  assign n19980 = ~n19968 & n19978;
  assign n19981 = ~n19979 & ~n19980;
  assign n19982 = n19927 & ~n19981;
  assign n19983 = ~n19927 & n19981;
  assign n19984 = ~n19982 & ~n19983;
  assign n19985 = pi99  & n8905;
  assign n19986 = pi100  & n8535;
  assign n19987 = pi101  & n8530;
  assign n19988 = n4730 & n8528;
  assign n19989 = ~n19986 & ~n19987;
  assign n19990 = ~n19985 & n19989;
  assign n19991 = ~n19988 & n19990;
  assign n19992 = pi53  & n19991;
  assign n19993 = ~pi53  & ~n19991;
  assign n19994 = ~n19992 & ~n19993;
  assign n19995 = ~n19984 & n19994;
  assign n19996 = n19984 & ~n19994;
  assign n19997 = ~n19995 & ~n19996;
  assign n19998 = ~n19926 & n19997;
  assign n19999 = n19926 & ~n19997;
  assign n20000 = ~n19998 & ~n19999;
  assign n20001 = ~n19925 & n20000;
  assign n20002 = n19925 & ~n20000;
  assign n20003 = ~n20001 & ~n20002;
  assign n20004 = ~n19915 & n20003;
  assign n20005 = n19915 & ~n20003;
  assign n20006 = ~n20004 & ~n20005;
  assign n20007 = pi105  & n7121;
  assign n20008 = pi106  & n6795;
  assign n20009 = pi107  & n6790;
  assign n20010 = n6189 & n6788;
  assign n20011 = ~n20008 & ~n20009;
  assign n20012 = ~n20007 & n20011;
  assign n20013 = ~n20010 & n20012;
  assign n20014 = pi47  & n20013;
  assign n20015 = ~pi47  & ~n20013;
  assign n20016 = ~n20014 & ~n20015;
  assign n20017 = n20006 & ~n20016;
  assign n20018 = ~n20006 & n20016;
  assign n20019 = ~n20017 & ~n20018;
  assign n20020 = n19914 & ~n20019;
  assign n20021 = ~n19914 & n20019;
  assign n20022 = ~n20020 & ~n20021;
  assign n20023 = pi108  & n6331;
  assign n20024 = pi109  & n6015;
  assign n20025 = pi110  & n6010;
  assign n20026 = n6008 & n6995;
  assign n20027 = ~n20024 & ~n20025;
  assign n20028 = ~n20023 & n20027;
  assign n20029 = ~n20026 & n20028;
  assign n20030 = pi44  & n20029;
  assign n20031 = ~pi44  & ~n20029;
  assign n20032 = ~n20030 & ~n20031;
  assign n20033 = n20022 & ~n20032;
  assign n20034 = ~n20022 & n20032;
  assign n20035 = ~n20033 & ~n20034;
  assign n20036 = n19913 & ~n20035;
  assign n20037 = ~n19913 & n20035;
  assign n20038 = ~n20036 & ~n20037;
  assign n20039 = pi111  & n5558;
  assign n20040 = pi112  & n5293;
  assign n20041 = pi113  & n5288;
  assign n20042 = n5286 & n7852;
  assign n20043 = ~n20040 & ~n20041;
  assign n20044 = ~n20039 & n20043;
  assign n20045 = ~n20042 & n20044;
  assign n20046 = pi41  & n20045;
  assign n20047 = ~pi41  & ~n20045;
  assign n20048 = ~n20046 & ~n20047;
  assign n20049 = n20038 & ~n20048;
  assign n20050 = ~n20038 & n20048;
  assign n20051 = ~n20049 & ~n20050;
  assign n20052 = n19912 & ~n20051;
  assign n20053 = ~n19912 & n20051;
  assign n20054 = ~n20052 & ~n20053;
  assign n20055 = pi114  & n4843;
  assign n20056 = pi115  & n4598;
  assign n20057 = pi116  & n4593;
  assign n20058 = n4591 & n8470;
  assign n20059 = ~n20056 & ~n20057;
  assign n20060 = ~n20055 & n20059;
  assign n20061 = ~n20058 & n20060;
  assign n20062 = pi38  & n20061;
  assign n20063 = ~pi38  & ~n20061;
  assign n20064 = ~n20062 & ~n20063;
  assign n20065 = n20054 & ~n20064;
  assign n20066 = ~n20054 & n20064;
  assign n20067 = ~n20065 & ~n20066;
  assign n20068 = n19684 & ~n19843;
  assign n20069 = ~n19844 & ~n20068;
  assign n20070 = n20067 & n20069;
  assign n20071 = ~n20067 & ~n20069;
  assign n20072 = ~n20070 & ~n20071;
  assign n20073 = ~n19911 & n20072;
  assign n20074 = n19911 & ~n20072;
  assign n20075 = ~n20073 & ~n20074;
  assign n20076 = n19901 & n20075;
  assign n20077 = ~n19901 & ~n20075;
  assign n20078 = ~n20076 & ~n20077;
  assign n20079 = pi123  & n3011;
  assign n20080 = pi124  & n2809;
  assign n20081 = pi125  & n2804;
  assign n20082 = n2802 & n11786;
  assign n20083 = ~n20080 & ~n20081;
  assign n20084 = ~n20079 & n20083;
  assign n20085 = ~n20082 & n20084;
  assign n20086 = pi29  & n20085;
  assign n20087 = ~pi29  & ~n20085;
  assign n20088 = ~n20086 & ~n20087;
  assign n20089 = ~n19672 & ~n19857;
  assign n20090 = ~n20088 & ~n20089;
  assign n20091 = n20088 & n20089;
  assign n20092 = ~n20090 & ~n20091;
  assign n20093 = n20078 & n20092;
  assign n20094 = ~n20078 & ~n20092;
  assign n20095 = ~n20093 & ~n20094;
  assign n20096 = ~n19656 & ~n19860;
  assign n20097 = pi126  & n2510;
  assign n20098 = pi127  & n2342;
  assign n20099 = n2335 & n12542;
  assign n20100 = ~n20097 & ~n20098;
  assign n20101 = ~n20099 & n20100;
  assign n20102 = pi26  & n20101;
  assign n20103 = ~pi26  & ~n20101;
  assign n20104 = ~n20102 & ~n20103;
  assign n20105 = ~n20096 & ~n20104;
  assign n20106 = n20096 & n20104;
  assign n20107 = ~n20105 & ~n20106;
  assign n20108 = n20095 & n20107;
  assign n20109 = ~n20095 & ~n20107;
  assign n20110 = ~n20108 & ~n20109;
  assign n20111 = ~n19887 & n20110;
  assign n20112 = n19887 & ~n20110;
  assign n20113 = ~n20111 & ~n20112;
  assign n20114 = ~n19886 & n20113;
  assign n20115 = n19886 & ~n20113;
  assign po88  = ~n20114 & ~n20115;
  assign n20117 = ~n20111 & ~n20114;
  assign n20118 = ~n20105 & ~n20108;
  assign n20119 = pi124  & n3011;
  assign n20120 = pi125  & n2809;
  assign n20121 = pi126  & n2804;
  assign n20122 = n2802 & n12148;
  assign n20123 = ~n20120 & ~n20121;
  assign n20124 = ~n20119 & n20123;
  assign n20125 = ~n20122 & n20124;
  assign n20126 = pi29  & n20125;
  assign n20127 = ~pi29  & ~n20125;
  assign n20128 = ~n20126 & ~n20127;
  assign n20129 = ~n19899 & ~n20076;
  assign n20130 = n20128 & n20129;
  assign n20131 = ~n20128 & ~n20129;
  assign n20132 = ~n20130 & ~n20131;
  assign n20133 = pi121  & n3553;
  assign n20134 = pi122  & n3334;
  assign n20135 = pi123  & n3329;
  assign n20136 = n3327 & n10754;
  assign n20137 = ~n20134 & ~n20135;
  assign n20138 = ~n20133 & n20137;
  assign n20139 = ~n20136 & n20138;
  assign n20140 = pi32  & n20139;
  assign n20141 = ~pi32  & ~n20139;
  assign n20142 = ~n20140 & ~n20141;
  assign n20143 = ~n20070 & ~n20073;
  assign n20144 = n20142 & n20143;
  assign n20145 = ~n20142 & ~n20143;
  assign n20146 = ~n20144 & ~n20145;
  assign n20147 = pi118  & n4176;
  assign n20148 = pi119  & n3938;
  assign n20149 = pi120  & n3933;
  assign n20150 = n3931 & n10047;
  assign n20151 = ~n20148 & ~n20149;
  assign n20152 = ~n20147 & n20151;
  assign n20153 = ~n20150 & n20152;
  assign n20154 = pi35  & n20153;
  assign n20155 = ~pi35  & ~n20153;
  assign n20156 = ~n20154 & ~n20155;
  assign n20157 = pi115  & n4843;
  assign n20158 = pi116  & n4598;
  assign n20159 = pi117  & n4593;
  assign n20160 = n4591 & n8784;
  assign n20161 = ~n20158 & ~n20159;
  assign n20162 = ~n20157 & n20161;
  assign n20163 = ~n20160 & n20162;
  assign n20164 = pi38  & n20163;
  assign n20165 = ~pi38  & ~n20163;
  assign n20166 = ~n20164 & ~n20165;
  assign n20167 = pi106  & n7121;
  assign n20168 = pi107  & n6795;
  assign n20169 = pi108  & n6790;
  assign n20170 = n6213 & n6788;
  assign n20171 = ~n20168 & ~n20169;
  assign n20172 = ~n20167 & n20171;
  assign n20173 = ~n20170 & n20172;
  assign n20174 = pi47  & n20173;
  assign n20175 = ~pi47  & ~n20173;
  assign n20176 = ~n20174 & ~n20175;
  assign n20177 = ~n19998 & ~n20001;
  assign n20178 = pi103  & n7969;
  assign n20179 = pi104  & n7636;
  assign n20180 = pi105  & n7631;
  assign n20181 = n5677 & n7629;
  assign n20182 = ~n20179 & ~n20180;
  assign n20183 = ~n20178 & n20182;
  assign n20184 = ~n20181 & n20183;
  assign n20185 = pi50  & n20184;
  assign n20186 = ~pi50  & ~n20184;
  assign n20187 = ~n20185 & ~n20186;
  assign n20188 = ~n19983 & ~n19996;
  assign n20189 = pi97  & n9858;
  assign n20190 = pi98  & n9508;
  assign n20191 = pi99  & n9503;
  assign n20192 = n4101 & n9501;
  assign n20193 = ~n20190 & ~n20191;
  assign n20194 = ~n20189 & n20193;
  assign n20195 = ~n20192 & n20194;
  assign n20196 = pi56  & n20195;
  assign n20197 = ~pi56  & ~n20195;
  assign n20198 = ~n20196 & ~n20197;
  assign n20199 = pi94  & n10886;
  assign n20200 = pi95  & n10495;
  assign n20201 = pi96  & n10490;
  assign n20202 = n3499 & n10488;
  assign n20203 = ~n20200 & ~n20201;
  assign n20204 = ~n20199 & n20203;
  assign n20205 = ~n20202 & n20204;
  assign n20206 = pi59  & n20205;
  assign n20207 = ~pi59  & ~n20205;
  assign n20208 = ~n20206 & ~n20207;
  assign n20209 = ~n19935 & ~n19947;
  assign n20210 = pi90  & n12277;
  assign n20211 = pi89  & n12276;
  assign n20212 = ~n20210 & ~n20211;
  assign n20213 = ~n19933 & n20212;
  assign n20214 = n19933 & ~n20212;
  assign n20215 = ~n20213 & ~n20214;
  assign n20216 = pi91  & n11910;
  assign n20217 = pi92  & n11529;
  assign n20218 = pi93  & n11524;
  assign n20219 = n2948 & n11522;
  assign n20220 = ~n20217 & ~n20218;
  assign n20221 = ~n20216 & n20220;
  assign n20222 = ~n20219 & n20221;
  assign n20223 = pi62  & n20222;
  assign n20224 = ~pi62  & ~n20222;
  assign n20225 = ~n20223 & ~n20224;
  assign n20226 = n20215 & ~n20225;
  assign n20227 = ~n20215 & n20225;
  assign n20228 = ~n20226 & ~n20227;
  assign n20229 = ~n20209 & n20228;
  assign n20230 = n20209 & ~n20228;
  assign n20231 = ~n20229 & ~n20230;
  assign n20232 = ~n20208 & n20231;
  assign n20233 = n20208 & ~n20231;
  assign n20234 = ~n20232 & ~n20233;
  assign n20235 = ~n19950 & n19962;
  assign n20236 = ~n19951 & ~n20235;
  assign n20237 = n20234 & n20236;
  assign n20238 = ~n20234 & ~n20236;
  assign n20239 = ~n20237 & ~n20238;
  assign n20240 = ~n20198 & n20239;
  assign n20241 = n20198 & ~n20239;
  assign n20242 = ~n20240 & ~n20241;
  assign n20243 = ~n19967 & n19978;
  assign n20244 = ~n19966 & ~n20243;
  assign n20245 = n20242 & n20244;
  assign n20246 = ~n20242 & ~n20244;
  assign n20247 = ~n20245 & ~n20246;
  assign n20248 = pi100  & n8905;
  assign n20249 = pi101  & n8535;
  assign n20250 = pi102  & n8530;
  assign n20251 = n4956 & n8528;
  assign n20252 = ~n20249 & ~n20250;
  assign n20253 = ~n20248 & n20252;
  assign n20254 = ~n20251 & n20253;
  assign n20255 = pi53  & n20254;
  assign n20256 = ~pi53  & ~n20254;
  assign n20257 = ~n20255 & ~n20256;
  assign n20258 = n20247 & ~n20257;
  assign n20259 = ~n20247 & n20257;
  assign n20260 = ~n20258 & ~n20259;
  assign n20261 = ~n20188 & n20260;
  assign n20262 = n20188 & ~n20260;
  assign n20263 = ~n20261 & ~n20262;
  assign n20264 = ~n20187 & n20263;
  assign n20265 = n20187 & ~n20263;
  assign n20266 = ~n20264 & ~n20265;
  assign n20267 = ~n20177 & n20266;
  assign n20268 = n20177 & ~n20266;
  assign n20269 = ~n20267 & ~n20268;
  assign n20270 = ~n20176 & n20269;
  assign n20271 = n20176 & ~n20269;
  assign n20272 = ~n20270 & ~n20271;
  assign n20273 = ~n20004 & n20016;
  assign n20274 = ~n20005 & ~n20273;
  assign n20275 = n20272 & n20274;
  assign n20276 = ~n20272 & ~n20274;
  assign n20277 = ~n20275 & ~n20276;
  assign n20278 = pi109  & n6331;
  assign n20279 = pi110  & n6015;
  assign n20280 = pi111  & n6010;
  assign n20281 = n6008 & n7272;
  assign n20282 = ~n20279 & ~n20280;
  assign n20283 = ~n20278 & n20282;
  assign n20284 = ~n20281 & n20283;
  assign n20285 = pi44  & n20284;
  assign n20286 = ~pi44  & ~n20284;
  assign n20287 = ~n20285 & ~n20286;
  assign n20288 = n20277 & ~n20287;
  assign n20289 = ~n20277 & n20287;
  assign n20290 = ~n20288 & ~n20289;
  assign n20291 = ~n20021 & n20032;
  assign n20292 = ~n20020 & ~n20291;
  assign n20293 = ~n20290 & ~n20292;
  assign n20294 = n20290 & n20292;
  assign n20295 = ~n20293 & ~n20294;
  assign n20296 = pi112  & n5558;
  assign n20297 = pi113  & n5293;
  assign n20298 = pi114  & n5288;
  assign n20299 = n5286 & n8146;
  assign n20300 = ~n20297 & ~n20298;
  assign n20301 = ~n20296 & n20300;
  assign n20302 = ~n20299 & n20301;
  assign n20303 = pi41  & n20302;
  assign n20304 = ~pi41  & ~n20302;
  assign n20305 = ~n20303 & ~n20304;
  assign n20306 = ~n20295 & n20305;
  assign n20307 = n20295 & ~n20305;
  assign n20308 = ~n20306 & ~n20307;
  assign n20309 = ~n20037 & n20048;
  assign n20310 = ~n20036 & ~n20309;
  assign n20311 = n20308 & n20310;
  assign n20312 = ~n20308 & ~n20310;
  assign n20313 = ~n20311 & ~n20312;
  assign n20314 = ~n20166 & n20313;
  assign n20315 = n20166 & ~n20313;
  assign n20316 = ~n20314 & ~n20315;
  assign n20317 = ~n20053 & n20064;
  assign n20318 = ~n20052 & ~n20317;
  assign n20319 = n20316 & n20318;
  assign n20320 = ~n20316 & ~n20318;
  assign n20321 = ~n20319 & ~n20320;
  assign n20322 = n20156 & ~n20321;
  assign n20323 = ~n20156 & n20321;
  assign n20324 = ~n20322 & ~n20323;
  assign n20325 = n20146 & n20324;
  assign n20326 = ~n20146 & ~n20324;
  assign n20327 = ~n20325 & ~n20326;
  assign n20328 = ~n20132 & ~n20327;
  assign n20329 = n20132 & n20327;
  assign n20330 = ~n20328 & ~n20329;
  assign n20331 = ~n20090 & ~n20093;
  assign n20332 = n2335 & ~n12539;
  assign n20333 = ~n2510 & ~n20332;
  assign n20334 = pi127  & ~n20333;
  assign n20335 = pi26  & ~n20334;
  assign n20336 = ~pi26  & n20334;
  assign n20337 = ~n20335 & ~n20336;
  assign n20338 = ~n20331 & ~n20337;
  assign n20339 = n20331 & n20337;
  assign n20340 = ~n20338 & ~n20339;
  assign n20341 = n20330 & n20340;
  assign n20342 = ~n20330 & ~n20340;
  assign n20343 = ~n20341 & ~n20342;
  assign n20344 = ~n20118 & n20343;
  assign n20345 = n20118 & ~n20343;
  assign n20346 = ~n20344 & ~n20345;
  assign n20347 = ~n20117 & n20346;
  assign n20348 = n20117 & ~n20346;
  assign po89  = ~n20347 & ~n20348;
  assign n20350 = ~n20338 & ~n20341;
  assign n20351 = ~n20311 & ~n20314;
  assign n20352 = pi116  & n4843;
  assign n20353 = pi117  & n4598;
  assign n20354 = pi118  & n4593;
  assign n20355 = n4591 & n9095;
  assign n20356 = ~n20353 & ~n20354;
  assign n20357 = ~n20352 & n20356;
  assign n20358 = ~n20355 & n20357;
  assign n20359 = pi38  & n20358;
  assign n20360 = ~pi38  & ~n20358;
  assign n20361 = ~n20359 & ~n20360;
  assign n20362 = ~n20294 & ~n20307;
  assign n20363 = ~n20267 & ~n20270;
  assign n20364 = pi107  & n7121;
  assign n20365 = pi108  & n6795;
  assign n20366 = pi109  & n6790;
  assign n20367 = n6715 & n6788;
  assign n20368 = ~n20365 & ~n20366;
  assign n20369 = ~n20364 & n20368;
  assign n20370 = ~n20367 & n20369;
  assign n20371 = pi47  & n20370;
  assign n20372 = ~pi47  & ~n20370;
  assign n20373 = ~n20371 & ~n20372;
  assign n20374 = ~n20261 & ~n20264;
  assign n20375 = ~n20237 & ~n20240;
  assign n20376 = pi95  & n10886;
  assign n20377 = pi96  & n10495;
  assign n20378 = pi97  & n10490;
  assign n20379 = n3691 & n10488;
  assign n20380 = ~n20377 & ~n20378;
  assign n20381 = ~n20376 & n20380;
  assign n20382 = ~n20379 & n20381;
  assign n20383 = pi59  & n20382;
  assign n20384 = ~pi59  & ~n20382;
  assign n20385 = ~n20383 & ~n20384;
  assign n20386 = ~n20229 & ~n20232;
  assign n20387 = n20385 & n20386;
  assign n20388 = ~n20385 & ~n20386;
  assign n20389 = ~n20387 & ~n20388;
  assign n20390 = ~n20213 & ~n20226;
  assign n20391 = pi91  & n12277;
  assign n20392 = pi90  & n12276;
  assign n20393 = ~n20391 & ~n20392;
  assign n20394 = ~pi26  & ~n20393;
  assign n20395 = pi26  & n20393;
  assign n20396 = ~n20394 & ~n20395;
  assign n20397 = ~n20212 & n20396;
  assign n20398 = n20212 & ~n20396;
  assign n20399 = ~n20397 & ~n20398;
  assign n20400 = ~n20390 & n20399;
  assign n20401 = n20390 & ~n20399;
  assign n20402 = ~n20400 & ~n20401;
  assign n20403 = pi92  & n11910;
  assign n20404 = pi93  & n11529;
  assign n20405 = pi94  & n11524;
  assign n20406 = n3280 & n11522;
  assign n20407 = ~n20404 & ~n20405;
  assign n20408 = ~n20403 & n20407;
  assign n20409 = ~n20406 & n20408;
  assign n20410 = pi62  & n20409;
  assign n20411 = ~pi62  & ~n20409;
  assign n20412 = ~n20410 & ~n20411;
  assign n20413 = n20402 & ~n20412;
  assign n20414 = ~n20402 & n20412;
  assign n20415 = ~n20413 & ~n20414;
  assign n20416 = ~n20389 & ~n20415;
  assign n20417 = n20389 & n20415;
  assign n20418 = ~n20416 & ~n20417;
  assign n20419 = pi98  & n9858;
  assign n20420 = pi99  & n9508;
  assign n20421 = pi100  & n9503;
  assign n20422 = n4501 & n9501;
  assign n20423 = ~n20420 & ~n20421;
  assign n20424 = ~n20419 & n20423;
  assign n20425 = ~n20422 & n20424;
  assign n20426 = pi56  & n20425;
  assign n20427 = ~pi56  & ~n20425;
  assign n20428 = ~n20426 & ~n20427;
  assign n20429 = n20418 & ~n20428;
  assign n20430 = ~n20418 & n20428;
  assign n20431 = ~n20429 & ~n20430;
  assign n20432 = n20375 & ~n20431;
  assign n20433 = ~n20375 & n20431;
  assign n20434 = ~n20432 & ~n20433;
  assign n20435 = pi101  & n8905;
  assign n20436 = pi102  & n8535;
  assign n20437 = pi103  & n8530;
  assign n20438 = n5188 & n8528;
  assign n20439 = ~n20436 & ~n20437;
  assign n20440 = ~n20435 & n20439;
  assign n20441 = ~n20438 & n20440;
  assign n20442 = pi53  & n20441;
  assign n20443 = ~pi53  & ~n20441;
  assign n20444 = ~n20442 & ~n20443;
  assign n20445 = n20434 & ~n20444;
  assign n20446 = ~n20434 & n20444;
  assign n20447 = ~n20445 & ~n20446;
  assign n20448 = ~n20245 & n20257;
  assign n20449 = ~n20246 & ~n20448;
  assign n20450 = ~n20447 & ~n20449;
  assign n20451 = n20447 & n20449;
  assign n20452 = ~n20450 & ~n20451;
  assign n20453 = pi104  & n7969;
  assign n20454 = pi105  & n7636;
  assign n20455 = pi106  & n7631;
  assign n20456 = n5701 & n7629;
  assign n20457 = ~n20454 & ~n20455;
  assign n20458 = ~n20453 & n20457;
  assign n20459 = ~n20456 & n20458;
  assign n20460 = pi50  & n20459;
  assign n20461 = ~pi50  & ~n20459;
  assign n20462 = ~n20460 & ~n20461;
  assign n20463 = n20452 & ~n20462;
  assign n20464 = ~n20452 & n20462;
  assign n20465 = ~n20463 & ~n20464;
  assign n20466 = ~n20374 & n20465;
  assign n20467 = n20374 & ~n20465;
  assign n20468 = ~n20466 & ~n20467;
  assign n20469 = ~n20373 & n20468;
  assign n20470 = n20373 & ~n20468;
  assign n20471 = ~n20469 & ~n20470;
  assign n20472 = n20363 & ~n20471;
  assign n20473 = ~n20363 & n20471;
  assign n20474 = ~n20472 & ~n20473;
  assign n20475 = pi110  & n6331;
  assign n20476 = pi111  & n6015;
  assign n20477 = pi112  & n6010;
  assign n20478 = n6008 & n7296;
  assign n20479 = ~n20476 & ~n20477;
  assign n20480 = ~n20475 & n20479;
  assign n20481 = ~n20478 & n20480;
  assign n20482 = pi44  & n20481;
  assign n20483 = ~pi44  & ~n20481;
  assign n20484 = ~n20482 & ~n20483;
  assign n20485 = n20474 & ~n20484;
  assign n20486 = ~n20474 & n20484;
  assign n20487 = ~n20485 & ~n20486;
  assign n20488 = ~n20275 & n20287;
  assign n20489 = ~n20276 & ~n20488;
  assign n20490 = ~n20487 & ~n20489;
  assign n20491 = n20487 & n20489;
  assign n20492 = ~n20490 & ~n20491;
  assign n20493 = pi113  & n5558;
  assign n20494 = pi114  & n5293;
  assign n20495 = pi115  & n5288;
  assign n20496 = n5286 & n8170;
  assign n20497 = ~n20494 & ~n20495;
  assign n20498 = ~n20493 & n20497;
  assign n20499 = ~n20496 & n20498;
  assign n20500 = pi41  & n20499;
  assign n20501 = ~pi41  & ~n20499;
  assign n20502 = ~n20500 & ~n20501;
  assign n20503 = n20492 & ~n20502;
  assign n20504 = ~n20492 & n20502;
  assign n20505 = ~n20503 & ~n20504;
  assign n20506 = n20362 & n20505;
  assign n20507 = ~n20362 & ~n20505;
  assign n20508 = ~n20506 & ~n20507;
  assign n20509 = n20361 & n20508;
  assign n20510 = ~n20361 & ~n20508;
  assign n20511 = ~n20509 & ~n20510;
  assign n20512 = ~n20351 & n20511;
  assign n20513 = n20351 & ~n20511;
  assign n20514 = ~n20512 & ~n20513;
  assign n20515 = pi119  & n4176;
  assign n20516 = pi120  & n3938;
  assign n20517 = pi121  & n3933;
  assign n20518 = n3931 & n10071;
  assign n20519 = ~n20516 & ~n20517;
  assign n20520 = ~n20515 & n20519;
  assign n20521 = ~n20518 & n20520;
  assign n20522 = pi35  & n20521;
  assign n20523 = ~pi35  & ~n20521;
  assign n20524 = ~n20522 & ~n20523;
  assign n20525 = n20514 & ~n20524;
  assign n20526 = ~n20514 & n20524;
  assign n20527 = ~n20525 & ~n20526;
  assign n20528 = n20156 & ~n20319;
  assign n20529 = ~n20320 & ~n20528;
  assign n20530 = ~n20527 & ~n20529;
  assign n20531 = n20527 & n20529;
  assign n20532 = ~n20530 & ~n20531;
  assign n20533 = pi122  & n3553;
  assign n20534 = pi123  & n3334;
  assign n20535 = pi124  & n3329;
  assign n20536 = n3327 & n11099;
  assign n20537 = ~n20534 & ~n20535;
  assign n20538 = ~n20533 & n20537;
  assign n20539 = ~n20536 & n20538;
  assign n20540 = pi32  & n20539;
  assign n20541 = ~pi32  & ~n20539;
  assign n20542 = ~n20540 & ~n20541;
  assign n20543 = ~n20145 & ~n20324;
  assign n20544 = ~n20144 & ~n20543;
  assign n20545 = n20542 & ~n20544;
  assign n20546 = ~n20542 & n20544;
  assign n20547 = ~n20545 & ~n20546;
  assign n20548 = n20532 & n20547;
  assign n20549 = ~n20532 & ~n20547;
  assign n20550 = ~n20548 & ~n20549;
  assign n20551 = ~n20131 & ~n20329;
  assign n20552 = pi125  & n3011;
  assign n20553 = pi126  & n2809;
  assign n20554 = pi127  & n2804;
  assign n20555 = n2802 & n12519;
  assign n20556 = ~n20553 & ~n20554;
  assign n20557 = ~n20552 & n20556;
  assign n20558 = ~n20555 & n20557;
  assign n20559 = pi29  & n20558;
  assign n20560 = ~pi29  & ~n20558;
  assign n20561 = ~n20559 & ~n20560;
  assign n20562 = ~n20551 & ~n20561;
  assign n20563 = n20551 & n20561;
  assign n20564 = ~n20562 & ~n20563;
  assign n20565 = n20550 & n20564;
  assign n20566 = ~n20550 & ~n20564;
  assign n20567 = ~n20565 & ~n20566;
  assign n20568 = n20350 & ~n20567;
  assign n20569 = ~n20350 & n20567;
  assign n20570 = ~n20568 & ~n20569;
  assign n20571 = ~n20344 & ~n20347;
  assign n20572 = n20570 & ~n20571;
  assign n20573 = ~n20570 & n20571;
  assign po90  = ~n20572 & ~n20573;
  assign n20575 = ~n20562 & ~n20565;
  assign n20576 = ~n20546 & ~n20548;
  assign n20577 = pi126  & n3011;
  assign n20578 = pi127  & n2809;
  assign n20579 = n2802 & n12542;
  assign n20580 = ~n20577 & ~n20578;
  assign n20581 = ~n20579 & n20580;
  assign n20582 = pi29  & n20581;
  assign n20583 = ~pi29  & ~n20581;
  assign n20584 = ~n20582 & ~n20583;
  assign n20585 = ~n20576 & ~n20584;
  assign n20586 = n20576 & n20584;
  assign n20587 = ~n20585 & ~n20586;
  assign n20588 = pi123  & n3553;
  assign n20589 = pi124  & n3334;
  assign n20590 = pi125  & n3329;
  assign n20591 = n3327 & n11786;
  assign n20592 = ~n20589 & ~n20590;
  assign n20593 = ~n20588 & n20592;
  assign n20594 = ~n20591 & n20593;
  assign n20595 = pi32  & n20594;
  assign n20596 = ~pi32  & ~n20594;
  assign n20597 = ~n20595 & ~n20596;
  assign n20598 = ~n20525 & ~n20531;
  assign n20599 = n20597 & n20598;
  assign n20600 = ~n20597 & ~n20598;
  assign n20601 = ~n20599 & ~n20600;
  assign n20602 = ~n20510 & ~n20512;
  assign n20603 = pi117  & n4843;
  assign n20604 = pi118  & n4598;
  assign n20605 = pi119  & n4593;
  assign n20606 = n4591 & n9412;
  assign n20607 = ~n20604 & ~n20605;
  assign n20608 = ~n20603 & n20607;
  assign n20609 = ~n20606 & n20608;
  assign n20610 = pi38  & n20609;
  assign n20611 = ~pi38  & ~n20609;
  assign n20612 = ~n20610 & ~n20611;
  assign n20613 = ~n20485 & ~n20491;
  assign n20614 = ~n20469 & ~n20473;
  assign n20615 = ~n20463 & ~n20466;
  assign n20616 = ~n20445 & ~n20451;
  assign n20617 = pi102  & n8905;
  assign n20618 = pi103  & n8535;
  assign n20619 = pi104  & n8530;
  assign n20620 = n5212 & n8528;
  assign n20621 = ~n20618 & ~n20619;
  assign n20622 = ~n20617 & n20621;
  assign n20623 = ~n20620 & n20622;
  assign n20624 = pi53  & n20623;
  assign n20625 = ~pi53  & ~n20623;
  assign n20626 = ~n20624 & ~n20625;
  assign n20627 = ~n20429 & ~n20433;
  assign n20628 = pi99  & n9858;
  assign n20629 = pi100  & n9508;
  assign n20630 = pi101  & n9503;
  assign n20631 = n4730 & n9501;
  assign n20632 = ~n20629 & ~n20630;
  assign n20633 = ~n20628 & n20632;
  assign n20634 = ~n20631 & n20633;
  assign n20635 = pi56  & n20634;
  assign n20636 = ~pi56  & ~n20634;
  assign n20637 = ~n20635 & ~n20636;
  assign n20638 = ~n20388 & ~n20417;
  assign n20639 = ~n20394 & ~n20397;
  assign n20640 = pi92  & n12277;
  assign n20641 = pi91  & n12276;
  assign n20642 = ~n20640 & ~n20641;
  assign n20643 = n20639 & ~n20642;
  assign n20644 = ~n20639 & n20642;
  assign n20645 = ~n20643 & ~n20644;
  assign n20646 = pi93  & n11910;
  assign n20647 = pi94  & n11529;
  assign n20648 = pi95  & n11524;
  assign n20649 = n3475 & n11522;
  assign n20650 = ~n20647 & ~n20648;
  assign n20651 = ~n20646 & n20650;
  assign n20652 = ~n20649 & n20651;
  assign n20653 = pi62  & n20652;
  assign n20654 = ~pi62  & ~n20652;
  assign n20655 = ~n20653 & ~n20654;
  assign n20656 = ~n20645 & n20655;
  assign n20657 = n20645 & ~n20655;
  assign n20658 = ~n20656 & ~n20657;
  assign n20659 = ~n20400 & n20412;
  assign n20660 = ~n20401 & ~n20659;
  assign n20661 = n20658 & n20660;
  assign n20662 = ~n20658 & ~n20660;
  assign n20663 = ~n20661 & ~n20662;
  assign n20664 = pi96  & n10886;
  assign n20665 = pi97  & n10495;
  assign n20666 = pi98  & n10490;
  assign n20667 = n3889 & n10488;
  assign n20668 = ~n20665 & ~n20666;
  assign n20669 = ~n20664 & n20668;
  assign n20670 = ~n20667 & n20669;
  assign n20671 = pi59  & n20670;
  assign n20672 = ~pi59  & ~n20670;
  assign n20673 = ~n20671 & ~n20672;
  assign n20674 = n20663 & ~n20673;
  assign n20675 = ~n20663 & n20673;
  assign n20676 = ~n20674 & ~n20675;
  assign n20677 = ~n20638 & n20676;
  assign n20678 = n20638 & ~n20676;
  assign n20679 = ~n20677 & ~n20678;
  assign n20680 = ~n20637 & n20679;
  assign n20681 = n20637 & ~n20679;
  assign n20682 = ~n20680 & ~n20681;
  assign n20683 = ~n20627 & n20682;
  assign n20684 = n20627 & ~n20682;
  assign n20685 = ~n20683 & ~n20684;
  assign n20686 = ~n20626 & n20685;
  assign n20687 = n20626 & ~n20685;
  assign n20688 = ~n20686 & ~n20687;
  assign n20689 = ~n20616 & n20688;
  assign n20690 = n20616 & ~n20688;
  assign n20691 = ~n20689 & ~n20690;
  assign n20692 = pi105  & n7969;
  assign n20693 = pi106  & n7636;
  assign n20694 = pi107  & n7631;
  assign n20695 = n6189 & n7629;
  assign n20696 = ~n20693 & ~n20694;
  assign n20697 = ~n20692 & n20696;
  assign n20698 = ~n20695 & n20697;
  assign n20699 = pi50  & n20698;
  assign n20700 = ~pi50  & ~n20698;
  assign n20701 = ~n20699 & ~n20700;
  assign n20702 = n20691 & ~n20701;
  assign n20703 = ~n20691 & n20701;
  assign n20704 = ~n20702 & ~n20703;
  assign n20705 = n20615 & ~n20704;
  assign n20706 = ~n20615 & n20704;
  assign n20707 = ~n20705 & ~n20706;
  assign n20708 = pi108  & n7121;
  assign n20709 = pi109  & n6795;
  assign n20710 = pi110  & n6790;
  assign n20711 = n6788 & n6995;
  assign n20712 = ~n20709 & ~n20710;
  assign n20713 = ~n20708 & n20712;
  assign n20714 = ~n20711 & n20713;
  assign n20715 = pi47  & n20714;
  assign n20716 = ~pi47  & ~n20714;
  assign n20717 = ~n20715 & ~n20716;
  assign n20718 = n20707 & ~n20717;
  assign n20719 = ~n20707 & n20717;
  assign n20720 = ~n20718 & ~n20719;
  assign n20721 = n20614 & ~n20720;
  assign n20722 = ~n20614 & n20720;
  assign n20723 = ~n20721 & ~n20722;
  assign n20724 = pi111  & n6331;
  assign n20725 = pi112  & n6015;
  assign n20726 = pi113  & n6010;
  assign n20727 = n6008 & n7852;
  assign n20728 = ~n20725 & ~n20726;
  assign n20729 = ~n20724 & n20728;
  assign n20730 = ~n20727 & n20729;
  assign n20731 = pi44  & n20730;
  assign n20732 = ~pi44  & ~n20730;
  assign n20733 = ~n20731 & ~n20732;
  assign n20734 = n20723 & ~n20733;
  assign n20735 = ~n20723 & n20733;
  assign n20736 = ~n20734 & ~n20735;
  assign n20737 = n20613 & ~n20736;
  assign n20738 = ~n20613 & n20736;
  assign n20739 = ~n20737 & ~n20738;
  assign n20740 = pi114  & n5558;
  assign n20741 = pi115  & n5293;
  assign n20742 = pi116  & n5288;
  assign n20743 = n5286 & n8470;
  assign n20744 = ~n20741 & ~n20742;
  assign n20745 = ~n20740 & n20744;
  assign n20746 = ~n20743 & n20745;
  assign n20747 = pi41  & n20746;
  assign n20748 = ~pi41  & ~n20746;
  assign n20749 = ~n20747 & ~n20748;
  assign n20750 = n20739 & ~n20749;
  assign n20751 = ~n20739 & n20749;
  assign n20752 = ~n20750 & ~n20751;
  assign n20753 = n20362 & ~n20503;
  assign n20754 = ~n20504 & ~n20753;
  assign n20755 = n20752 & n20754;
  assign n20756 = ~n20752 & ~n20754;
  assign n20757 = ~n20755 & ~n20756;
  assign n20758 = ~n20612 & n20757;
  assign n20759 = n20612 & ~n20757;
  assign n20760 = ~n20758 & ~n20759;
  assign n20761 = ~n20602 & n20760;
  assign n20762 = n20602 & ~n20760;
  assign n20763 = ~n20761 & ~n20762;
  assign n20764 = pi120  & n4176;
  assign n20765 = pi121  & n3938;
  assign n20766 = pi122  & n3933;
  assign n20767 = n3931 & n10729;
  assign n20768 = ~n20765 & ~n20766;
  assign n20769 = ~n20764 & n20768;
  assign n20770 = ~n20767 & n20769;
  assign n20771 = pi35  & n20770;
  assign n20772 = ~pi35  & ~n20770;
  assign n20773 = ~n20771 & ~n20772;
  assign n20774 = n20763 & ~n20773;
  assign n20775 = ~n20763 & n20773;
  assign n20776 = ~n20774 & ~n20775;
  assign n20777 = n20601 & n20776;
  assign n20778 = ~n20601 & ~n20776;
  assign n20779 = ~n20777 & ~n20778;
  assign n20780 = n20587 & n20779;
  assign n20781 = ~n20587 & ~n20779;
  assign n20782 = ~n20780 & ~n20781;
  assign n20783 = n20575 & ~n20782;
  assign n20784 = ~n20575 & n20782;
  assign n20785 = ~n20783 & ~n20784;
  assign n20786 = ~n20569 & ~n20572;
  assign n20787 = n20785 & ~n20786;
  assign n20788 = ~n20785 & n20786;
  assign po91  = ~n20787 & ~n20788;
  assign n20790 = ~n20784 & ~n20787;
  assign n20791 = ~n20585 & ~n20780;
  assign n20792 = pi124  & n3553;
  assign n20793 = pi125  & n3334;
  assign n20794 = pi126  & n3329;
  assign n20795 = n3327 & n12148;
  assign n20796 = ~n20793 & ~n20794;
  assign n20797 = ~n20792 & n20796;
  assign n20798 = ~n20795 & n20797;
  assign n20799 = pi32  & n20798;
  assign n20800 = ~pi32  & ~n20798;
  assign n20801 = ~n20799 & ~n20800;
  assign n20802 = ~n20761 & n20773;
  assign n20803 = ~n20762 & ~n20802;
  assign n20804 = n20801 & ~n20803;
  assign n20805 = ~n20801 & n20803;
  assign n20806 = ~n20804 & ~n20805;
  assign n20807 = ~n20755 & ~n20758;
  assign n20808 = pi118  & n4843;
  assign n20809 = pi119  & n4598;
  assign n20810 = pi120  & n4593;
  assign n20811 = n4591 & n10047;
  assign n20812 = ~n20809 & ~n20810;
  assign n20813 = ~n20808 & n20812;
  assign n20814 = ~n20811 & n20813;
  assign n20815 = pi38  & n20814;
  assign n20816 = ~pi38  & ~n20814;
  assign n20817 = ~n20815 & ~n20816;
  assign n20818 = pi115  & n5558;
  assign n20819 = pi116  & n5293;
  assign n20820 = pi117  & n5288;
  assign n20821 = n5286 & n8784;
  assign n20822 = ~n20819 & ~n20820;
  assign n20823 = ~n20818 & n20822;
  assign n20824 = ~n20821 & n20823;
  assign n20825 = pi41  & n20824;
  assign n20826 = ~pi41  & ~n20824;
  assign n20827 = ~n20825 & ~n20826;
  assign n20828 = pi106  & n7969;
  assign n20829 = pi107  & n7636;
  assign n20830 = pi108  & n7631;
  assign n20831 = n6213 & n7629;
  assign n20832 = ~n20829 & ~n20830;
  assign n20833 = ~n20828 & n20832;
  assign n20834 = ~n20831 & n20833;
  assign n20835 = pi50  & n20834;
  assign n20836 = ~pi50  & ~n20834;
  assign n20837 = ~n20835 & ~n20836;
  assign n20838 = ~n20683 & ~n20686;
  assign n20839 = pi103  & n8905;
  assign n20840 = pi104  & n8535;
  assign n20841 = pi105  & n8530;
  assign n20842 = n5677 & n8528;
  assign n20843 = ~n20840 & ~n20841;
  assign n20844 = ~n20839 & n20843;
  assign n20845 = ~n20842 & n20844;
  assign n20846 = pi53  & n20845;
  assign n20847 = ~pi53  & ~n20845;
  assign n20848 = ~n20846 & ~n20847;
  assign n20849 = ~n20677 & ~n20680;
  assign n20850 = pi97  & n10886;
  assign n20851 = pi98  & n10495;
  assign n20852 = pi99  & n10490;
  assign n20853 = n4101 & n10488;
  assign n20854 = ~n20851 & ~n20852;
  assign n20855 = ~n20850 & n20854;
  assign n20856 = ~n20853 & n20855;
  assign n20857 = pi59  & n20856;
  assign n20858 = ~pi59  & ~n20856;
  assign n20859 = ~n20857 & ~n20858;
  assign n20860 = pi94  & n11910;
  assign n20861 = pi95  & n11529;
  assign n20862 = pi96  & n11524;
  assign n20863 = n3499 & n11522;
  assign n20864 = ~n20861 & ~n20862;
  assign n20865 = ~n20860 & n20864;
  assign n20866 = ~n20863 & n20865;
  assign n20867 = pi62  & n20866;
  assign n20868 = ~pi62  & ~n20866;
  assign n20869 = ~n20867 & ~n20868;
  assign n20870 = ~n20644 & ~n20657;
  assign n20871 = pi93  & n12277;
  assign n20872 = pi92  & n12276;
  assign n20873 = ~n20871 & ~n20872;
  assign n20874 = n20642 & ~n20873;
  assign n20875 = ~n20642 & n20873;
  assign n20876 = ~n20874 & ~n20875;
  assign n20877 = ~n20870 & n20876;
  assign n20878 = n20870 & ~n20876;
  assign n20879 = ~n20877 & ~n20878;
  assign n20880 = ~n20869 & n20879;
  assign n20881 = n20869 & ~n20879;
  assign n20882 = ~n20880 & ~n20881;
  assign n20883 = ~n20859 & n20882;
  assign n20884 = n20859 & ~n20882;
  assign n20885 = ~n20883 & ~n20884;
  assign n20886 = ~n20661 & n20673;
  assign n20887 = ~n20662 & ~n20886;
  assign n20888 = n20885 & n20887;
  assign n20889 = ~n20885 & ~n20887;
  assign n20890 = ~n20888 & ~n20889;
  assign n20891 = pi100  & n9858;
  assign n20892 = pi101  & n9508;
  assign n20893 = pi102  & n9503;
  assign n20894 = n4956 & n9501;
  assign n20895 = ~n20892 & ~n20893;
  assign n20896 = ~n20891 & n20895;
  assign n20897 = ~n20894 & n20896;
  assign n20898 = pi56  & n20897;
  assign n20899 = ~pi56  & ~n20897;
  assign n20900 = ~n20898 & ~n20899;
  assign n20901 = n20890 & ~n20900;
  assign n20902 = ~n20890 & n20900;
  assign n20903 = ~n20901 & ~n20902;
  assign n20904 = ~n20849 & n20903;
  assign n20905 = n20849 & ~n20903;
  assign n20906 = ~n20904 & ~n20905;
  assign n20907 = ~n20848 & n20906;
  assign n20908 = n20848 & ~n20906;
  assign n20909 = ~n20907 & ~n20908;
  assign n20910 = ~n20838 & n20909;
  assign n20911 = n20838 & ~n20909;
  assign n20912 = ~n20910 & ~n20911;
  assign n20913 = ~n20837 & n20912;
  assign n20914 = n20837 & ~n20912;
  assign n20915 = ~n20913 & ~n20914;
  assign n20916 = ~n20689 & n20701;
  assign n20917 = ~n20690 & ~n20916;
  assign n20918 = n20915 & n20917;
  assign n20919 = ~n20915 & ~n20917;
  assign n20920 = ~n20918 & ~n20919;
  assign n20921 = pi109  & n7121;
  assign n20922 = pi110  & n6795;
  assign n20923 = pi111  & n6790;
  assign n20924 = n6788 & n7272;
  assign n20925 = ~n20922 & ~n20923;
  assign n20926 = ~n20921 & n20925;
  assign n20927 = ~n20924 & n20926;
  assign n20928 = pi47  & n20927;
  assign n20929 = ~pi47  & ~n20927;
  assign n20930 = ~n20928 & ~n20929;
  assign n20931 = n20920 & ~n20930;
  assign n20932 = ~n20920 & n20930;
  assign n20933 = ~n20931 & ~n20932;
  assign n20934 = ~n20706 & n20717;
  assign n20935 = ~n20705 & ~n20934;
  assign n20936 = ~n20933 & ~n20935;
  assign n20937 = n20933 & n20935;
  assign n20938 = ~n20936 & ~n20937;
  assign n20939 = pi112  & n6331;
  assign n20940 = pi113  & n6015;
  assign n20941 = pi114  & n6010;
  assign n20942 = n6008 & n8146;
  assign n20943 = ~n20940 & ~n20941;
  assign n20944 = ~n20939 & n20943;
  assign n20945 = ~n20942 & n20944;
  assign n20946 = pi44  & n20945;
  assign n20947 = ~pi44  & ~n20945;
  assign n20948 = ~n20946 & ~n20947;
  assign n20949 = ~n20938 & n20948;
  assign n20950 = n20938 & ~n20948;
  assign n20951 = ~n20949 & ~n20950;
  assign n20952 = ~n20722 & n20733;
  assign n20953 = ~n20721 & ~n20952;
  assign n20954 = n20951 & n20953;
  assign n20955 = ~n20951 & ~n20953;
  assign n20956 = ~n20954 & ~n20955;
  assign n20957 = ~n20827 & n20956;
  assign n20958 = n20827 & ~n20956;
  assign n20959 = ~n20957 & ~n20958;
  assign n20960 = ~n20738 & n20749;
  assign n20961 = ~n20737 & ~n20960;
  assign n20962 = n20959 & n20961;
  assign n20963 = ~n20959 & ~n20961;
  assign n20964 = ~n20962 & ~n20963;
  assign n20965 = ~n20817 & n20964;
  assign n20966 = n20817 & ~n20964;
  assign n20967 = ~n20965 & ~n20966;
  assign n20968 = ~n20807 & n20967;
  assign n20969 = n20807 & ~n20967;
  assign n20970 = ~n20968 & ~n20969;
  assign n20971 = pi121  & n4176;
  assign n20972 = pi122  & n3938;
  assign n20973 = pi123  & n3933;
  assign n20974 = n3931 & n10754;
  assign n20975 = ~n20972 & ~n20973;
  assign n20976 = ~n20971 & n20975;
  assign n20977 = ~n20974 & n20976;
  assign n20978 = pi35  & n20977;
  assign n20979 = ~pi35  & ~n20977;
  assign n20980 = ~n20978 & ~n20979;
  assign n20981 = n20970 & ~n20980;
  assign n20982 = ~n20970 & n20980;
  assign n20983 = ~n20981 & ~n20982;
  assign n20984 = ~n20806 & ~n20983;
  assign n20985 = n20806 & n20983;
  assign n20986 = ~n20984 & ~n20985;
  assign n20987 = ~n20600 & ~n20777;
  assign n20988 = n2802 & ~n12539;
  assign n20989 = ~n3011 & ~n20988;
  assign n20990 = pi127  & ~n20989;
  assign n20991 = pi29  & ~n20990;
  assign n20992 = ~pi29  & n20990;
  assign n20993 = ~n20991 & ~n20992;
  assign n20994 = ~n20987 & ~n20993;
  assign n20995 = n20987 & n20993;
  assign n20996 = ~n20994 & ~n20995;
  assign n20997 = n20986 & n20996;
  assign n20998 = ~n20986 & ~n20996;
  assign n20999 = ~n20997 & ~n20998;
  assign n21000 = ~n20791 & n20999;
  assign n21001 = n20791 & ~n20999;
  assign n21002 = ~n21000 & ~n21001;
  assign n21003 = ~n20790 & n21002;
  assign n21004 = n20790 & ~n21002;
  assign po92  = ~n21003 & ~n21004;
  assign n21006 = ~n21000 & ~n21003;
  assign n21007 = ~n20994 & ~n20997;
  assign n21008 = ~n20962 & ~n20965;
  assign n21009 = ~n20954 & ~n20957;
  assign n21010 = pi116  & n5558;
  assign n21011 = pi117  & n5293;
  assign n21012 = pi118  & n5288;
  assign n21013 = n5286 & n9095;
  assign n21014 = ~n21011 & ~n21012;
  assign n21015 = ~n21010 & n21014;
  assign n21016 = ~n21013 & n21015;
  assign n21017 = pi41  & n21016;
  assign n21018 = ~pi41  & ~n21016;
  assign n21019 = ~n21017 & ~n21018;
  assign n21020 = ~n20937 & ~n20950;
  assign n21021 = ~n20910 & ~n20913;
  assign n21022 = pi107  & n7969;
  assign n21023 = pi108  & n7636;
  assign n21024 = pi109  & n7631;
  assign n21025 = n6715 & n7629;
  assign n21026 = ~n21023 & ~n21024;
  assign n21027 = ~n21022 & n21026;
  assign n21028 = ~n21025 & n21027;
  assign n21029 = pi50  & n21028;
  assign n21030 = ~pi50  & ~n21028;
  assign n21031 = ~n21029 & ~n21030;
  assign n21032 = ~n20904 & ~n20907;
  assign n21033 = ~n20880 & ~n20883;
  assign n21034 = pi98  & n10886;
  assign n21035 = pi99  & n10495;
  assign n21036 = pi100  & n10490;
  assign n21037 = n4501 & n10488;
  assign n21038 = ~n21035 & ~n21036;
  assign n21039 = ~n21034 & n21038;
  assign n21040 = ~n21037 & n21039;
  assign n21041 = pi59  & n21040;
  assign n21042 = ~pi59  & ~n21040;
  assign n21043 = ~n21041 & ~n21042;
  assign n21044 = pi95  & n11910;
  assign n21045 = pi96  & n11529;
  assign n21046 = pi97  & n11524;
  assign n21047 = n3691 & n11522;
  assign n21048 = ~n21045 & ~n21046;
  assign n21049 = ~n21044 & n21048;
  assign n21050 = ~n21047 & n21049;
  assign n21051 = pi62  & n21050;
  assign n21052 = ~pi62  & ~n21050;
  assign n21053 = ~n21051 & ~n21052;
  assign n21054 = ~n20875 & ~n20877;
  assign n21055 = pi94  & n12277;
  assign n21056 = pi93  & n12276;
  assign n21057 = ~n21055 & ~n21056;
  assign n21058 = ~pi29  & ~n21057;
  assign n21059 = pi29  & n21057;
  assign n21060 = ~n21058 & ~n21059;
  assign n21061 = ~n20873 & n21060;
  assign n21062 = n20873 & ~n21060;
  assign n21063 = ~n21061 & ~n21062;
  assign n21064 = ~n21054 & n21063;
  assign n21065 = n21054 & ~n21063;
  assign n21066 = ~n21064 & ~n21065;
  assign n21067 = ~n21053 & n21066;
  assign n21068 = n21053 & ~n21066;
  assign n21069 = ~n21067 & ~n21068;
  assign n21070 = ~n21043 & n21069;
  assign n21071 = n21043 & ~n21069;
  assign n21072 = ~n21070 & ~n21071;
  assign n21073 = ~n21033 & n21072;
  assign n21074 = n21033 & ~n21072;
  assign n21075 = ~n21073 & ~n21074;
  assign n21076 = pi101  & n9858;
  assign n21077 = pi102  & n9508;
  assign n21078 = pi103  & n9503;
  assign n21079 = n5188 & n9501;
  assign n21080 = ~n21077 & ~n21078;
  assign n21081 = ~n21076 & n21080;
  assign n21082 = ~n21079 & n21081;
  assign n21083 = pi56  & n21082;
  assign n21084 = ~pi56  & ~n21082;
  assign n21085 = ~n21083 & ~n21084;
  assign n21086 = n21075 & ~n21085;
  assign n21087 = ~n21075 & n21085;
  assign n21088 = ~n21086 & ~n21087;
  assign n21089 = ~n20888 & n20900;
  assign n21090 = ~n20889 & ~n21089;
  assign n21091 = ~n21088 & ~n21090;
  assign n21092 = n21088 & n21090;
  assign n21093 = ~n21091 & ~n21092;
  assign n21094 = pi104  & n8905;
  assign n21095 = pi105  & n8535;
  assign n21096 = pi106  & n8530;
  assign n21097 = n5701 & n8528;
  assign n21098 = ~n21095 & ~n21096;
  assign n21099 = ~n21094 & n21098;
  assign n21100 = ~n21097 & n21099;
  assign n21101 = pi53  & n21100;
  assign n21102 = ~pi53  & ~n21100;
  assign n21103 = ~n21101 & ~n21102;
  assign n21104 = n21093 & ~n21103;
  assign n21105 = ~n21093 & n21103;
  assign n21106 = ~n21104 & ~n21105;
  assign n21107 = ~n21032 & n21106;
  assign n21108 = n21032 & ~n21106;
  assign n21109 = ~n21107 & ~n21108;
  assign n21110 = ~n21031 & n21109;
  assign n21111 = n21031 & ~n21109;
  assign n21112 = ~n21110 & ~n21111;
  assign n21113 = n21021 & ~n21112;
  assign n21114 = ~n21021 & n21112;
  assign n21115 = ~n21113 & ~n21114;
  assign n21116 = pi110  & n7121;
  assign n21117 = pi111  & n6795;
  assign n21118 = pi112  & n6790;
  assign n21119 = n6788 & n7296;
  assign n21120 = ~n21117 & ~n21118;
  assign n21121 = ~n21116 & n21120;
  assign n21122 = ~n21119 & n21121;
  assign n21123 = pi47  & n21122;
  assign n21124 = ~pi47  & ~n21122;
  assign n21125 = ~n21123 & ~n21124;
  assign n21126 = n21115 & ~n21125;
  assign n21127 = ~n21115 & n21125;
  assign n21128 = ~n21126 & ~n21127;
  assign n21129 = ~n20918 & n20930;
  assign n21130 = ~n20919 & ~n21129;
  assign n21131 = ~n21128 & ~n21130;
  assign n21132 = n21128 & n21130;
  assign n21133 = ~n21131 & ~n21132;
  assign n21134 = pi113  & n6331;
  assign n21135 = pi114  & n6015;
  assign n21136 = pi115  & n6010;
  assign n21137 = n6008 & n8170;
  assign n21138 = ~n21135 & ~n21136;
  assign n21139 = ~n21134 & n21138;
  assign n21140 = ~n21137 & n21139;
  assign n21141 = pi44  & n21140;
  assign n21142 = ~pi44  & ~n21140;
  assign n21143 = ~n21141 & ~n21142;
  assign n21144 = n21133 & ~n21143;
  assign n21145 = ~n21133 & n21143;
  assign n21146 = ~n21144 & ~n21145;
  assign n21147 = n21020 & n21146;
  assign n21148 = ~n21020 & ~n21146;
  assign n21149 = ~n21147 & ~n21148;
  assign n21150 = n21019 & n21149;
  assign n21151 = ~n21019 & ~n21149;
  assign n21152 = ~n21150 & ~n21151;
  assign n21153 = ~n21009 & n21152;
  assign n21154 = n21009 & ~n21152;
  assign n21155 = ~n21153 & ~n21154;
  assign n21156 = pi119  & n4843;
  assign n21157 = pi120  & n4598;
  assign n21158 = pi121  & n4593;
  assign n21159 = n4591 & n10071;
  assign n21160 = ~n21157 & ~n21158;
  assign n21161 = ~n21156 & n21160;
  assign n21162 = ~n21159 & n21161;
  assign n21163 = pi38  & n21162;
  assign n21164 = ~pi38  & ~n21162;
  assign n21165 = ~n21163 & ~n21164;
  assign n21166 = n21155 & ~n21165;
  assign n21167 = ~n21155 & n21165;
  assign n21168 = ~n21166 & ~n21167;
  assign n21169 = n21008 & ~n21168;
  assign n21170 = ~n21008 & n21168;
  assign n21171 = ~n21169 & ~n21170;
  assign n21172 = pi122  & n4176;
  assign n21173 = pi123  & n3938;
  assign n21174 = pi124  & n3933;
  assign n21175 = n3931 & n11099;
  assign n21176 = ~n21173 & ~n21174;
  assign n21177 = ~n21172 & n21176;
  assign n21178 = ~n21175 & n21177;
  assign n21179 = pi35  & n21178;
  assign n21180 = ~pi35  & ~n21178;
  assign n21181 = ~n21179 & ~n21180;
  assign n21182 = n21171 & ~n21181;
  assign n21183 = ~n21171 & n21181;
  assign n21184 = ~n21182 & ~n21183;
  assign n21185 = ~n20968 & n20980;
  assign n21186 = ~n20969 & ~n21185;
  assign n21187 = ~n21184 & ~n21186;
  assign n21188 = n21184 & n21186;
  assign n21189 = ~n21187 & ~n21188;
  assign n21190 = ~n20805 & ~n20985;
  assign n21191 = pi125  & n3553;
  assign n21192 = pi126  & n3334;
  assign n21193 = pi127  & n3329;
  assign n21194 = n3327 & n12519;
  assign n21195 = ~n21192 & ~n21193;
  assign n21196 = ~n21191 & n21195;
  assign n21197 = ~n21194 & n21196;
  assign n21198 = pi32  & n21197;
  assign n21199 = ~pi32  & ~n21197;
  assign n21200 = ~n21198 & ~n21199;
  assign n21201 = ~n21190 & ~n21200;
  assign n21202 = n21190 & n21200;
  assign n21203 = ~n21201 & ~n21202;
  assign n21204 = ~n21189 & ~n21203;
  assign n21205 = n21189 & n21203;
  assign n21206 = ~n21204 & ~n21205;
  assign n21207 = ~n21007 & n21206;
  assign n21208 = n21007 & ~n21206;
  assign n21209 = ~n21207 & ~n21208;
  assign n21210 = ~n21006 & n21209;
  assign n21211 = n21006 & ~n21209;
  assign po93  = ~n21210 & ~n21211;
  assign n21213 = ~n21207 & ~n21210;
  assign n21214 = ~n21201 & ~n21205;
  assign n21215 = ~n21182 & ~n21188;
  assign n21216 = pi126  & n3553;
  assign n21217 = pi127  & n3334;
  assign n21218 = n3327 & n12542;
  assign n21219 = ~n21216 & ~n21217;
  assign n21220 = ~n21218 & n21219;
  assign n21221 = pi32  & n21220;
  assign n21222 = ~pi32  & ~n21220;
  assign n21223 = ~n21221 & ~n21222;
  assign n21224 = ~n21215 & ~n21223;
  assign n21225 = n21215 & n21223;
  assign n21226 = ~n21224 & ~n21225;
  assign n21227 = ~n21166 & ~n21170;
  assign n21228 = ~n21151 & ~n21153;
  assign n21229 = pi117  & n5558;
  assign n21230 = pi118  & n5293;
  assign n21231 = pi119  & n5288;
  assign n21232 = n5286 & n9412;
  assign n21233 = ~n21230 & ~n21231;
  assign n21234 = ~n21229 & n21233;
  assign n21235 = ~n21232 & n21234;
  assign n21236 = pi41  & n21235;
  assign n21237 = ~pi41  & ~n21235;
  assign n21238 = ~n21236 & ~n21237;
  assign n21239 = ~n21126 & ~n21132;
  assign n21240 = ~n21110 & ~n21114;
  assign n21241 = ~n21104 & ~n21107;
  assign n21242 = ~n21086 & ~n21092;
  assign n21243 = pi102  & n9858;
  assign n21244 = pi103  & n9508;
  assign n21245 = pi104  & n9503;
  assign n21246 = n5212 & n9501;
  assign n21247 = ~n21244 & ~n21245;
  assign n21248 = ~n21243 & n21247;
  assign n21249 = ~n21246 & n21248;
  assign n21250 = pi56  & n21249;
  assign n21251 = ~pi56  & ~n21249;
  assign n21252 = ~n21250 & ~n21251;
  assign n21253 = ~n21070 & ~n21073;
  assign n21254 = pi99  & n10886;
  assign n21255 = pi100  & n10495;
  assign n21256 = pi101  & n10490;
  assign n21257 = n4730 & n10488;
  assign n21258 = ~n21255 & ~n21256;
  assign n21259 = ~n21254 & n21258;
  assign n21260 = ~n21257 & n21259;
  assign n21261 = pi59  & n21260;
  assign n21262 = ~pi59  & ~n21260;
  assign n21263 = ~n21261 & ~n21262;
  assign n21264 = ~n21064 & ~n21067;
  assign n21265 = ~n20873 & ~n21059;
  assign n21266 = ~n21058 & ~n21265;
  assign n21267 = pi95  & n12277;
  assign n21268 = pi94  & n12276;
  assign n21269 = ~n21267 & ~n21268;
  assign n21270 = n21266 & ~n21269;
  assign n21271 = ~n21266 & n21269;
  assign n21272 = ~n21270 & ~n21271;
  assign n21273 = pi96  & n11910;
  assign n21274 = pi97  & n11529;
  assign n21275 = pi98  & n11524;
  assign n21276 = n3889 & n11522;
  assign n21277 = ~n21274 & ~n21275;
  assign n21278 = ~n21273 & n21277;
  assign n21279 = ~n21276 & n21278;
  assign n21280 = pi62  & n21279;
  assign n21281 = ~pi62  & ~n21279;
  assign n21282 = ~n21280 & ~n21281;
  assign n21283 = ~n21272 & n21282;
  assign n21284 = n21272 & ~n21282;
  assign n21285 = ~n21283 & ~n21284;
  assign n21286 = ~n21264 & n21285;
  assign n21287 = n21264 & ~n21285;
  assign n21288 = ~n21286 & ~n21287;
  assign n21289 = ~n21263 & n21288;
  assign n21290 = n21263 & ~n21288;
  assign n21291 = ~n21289 & ~n21290;
  assign n21292 = ~n21253 & n21291;
  assign n21293 = n21253 & ~n21291;
  assign n21294 = ~n21292 & ~n21293;
  assign n21295 = ~n21252 & n21294;
  assign n21296 = n21252 & ~n21294;
  assign n21297 = ~n21295 & ~n21296;
  assign n21298 = ~n21242 & n21297;
  assign n21299 = n21242 & ~n21297;
  assign n21300 = ~n21298 & ~n21299;
  assign n21301 = pi105  & n8905;
  assign n21302 = pi106  & n8535;
  assign n21303 = pi107  & n8530;
  assign n21304 = n6189 & n8528;
  assign n21305 = ~n21302 & ~n21303;
  assign n21306 = ~n21301 & n21305;
  assign n21307 = ~n21304 & n21306;
  assign n21308 = pi53  & n21307;
  assign n21309 = ~pi53  & ~n21307;
  assign n21310 = ~n21308 & ~n21309;
  assign n21311 = n21300 & ~n21310;
  assign n21312 = ~n21300 & n21310;
  assign n21313 = ~n21311 & ~n21312;
  assign n21314 = n21241 & ~n21313;
  assign n21315 = ~n21241 & n21313;
  assign n21316 = ~n21314 & ~n21315;
  assign n21317 = pi108  & n7969;
  assign n21318 = pi109  & n7636;
  assign n21319 = pi110  & n7631;
  assign n21320 = n6995 & n7629;
  assign n21321 = ~n21318 & ~n21319;
  assign n21322 = ~n21317 & n21321;
  assign n21323 = ~n21320 & n21322;
  assign n21324 = pi50  & n21323;
  assign n21325 = ~pi50  & ~n21323;
  assign n21326 = ~n21324 & ~n21325;
  assign n21327 = n21316 & ~n21326;
  assign n21328 = ~n21316 & n21326;
  assign n21329 = ~n21327 & ~n21328;
  assign n21330 = n21240 & ~n21329;
  assign n21331 = ~n21240 & n21329;
  assign n21332 = ~n21330 & ~n21331;
  assign n21333 = pi111  & n7121;
  assign n21334 = pi112  & n6795;
  assign n21335 = pi113  & n6790;
  assign n21336 = n6788 & n7852;
  assign n21337 = ~n21334 & ~n21335;
  assign n21338 = ~n21333 & n21337;
  assign n21339 = ~n21336 & n21338;
  assign n21340 = pi47  & n21339;
  assign n21341 = ~pi47  & ~n21339;
  assign n21342 = ~n21340 & ~n21341;
  assign n21343 = n21332 & ~n21342;
  assign n21344 = ~n21332 & n21342;
  assign n21345 = ~n21343 & ~n21344;
  assign n21346 = n21239 & ~n21345;
  assign n21347 = ~n21239 & n21345;
  assign n21348 = ~n21346 & ~n21347;
  assign n21349 = pi114  & n6331;
  assign n21350 = pi115  & n6015;
  assign n21351 = pi116  & n6010;
  assign n21352 = n6008 & n8470;
  assign n21353 = ~n21350 & ~n21351;
  assign n21354 = ~n21349 & n21353;
  assign n21355 = ~n21352 & n21354;
  assign n21356 = pi44  & n21355;
  assign n21357 = ~pi44  & ~n21355;
  assign n21358 = ~n21356 & ~n21357;
  assign n21359 = n21348 & ~n21358;
  assign n21360 = ~n21348 & n21358;
  assign n21361 = ~n21359 & ~n21360;
  assign n21362 = n21020 & ~n21144;
  assign n21363 = ~n21145 & ~n21362;
  assign n21364 = n21361 & n21363;
  assign n21365 = ~n21361 & ~n21363;
  assign n21366 = ~n21364 & ~n21365;
  assign n21367 = ~n21238 & n21366;
  assign n21368 = n21238 & ~n21366;
  assign n21369 = ~n21367 & ~n21368;
  assign n21370 = ~n21228 & n21369;
  assign n21371 = n21228 & ~n21369;
  assign n21372 = ~n21370 & ~n21371;
  assign n21373 = pi120  & n4843;
  assign n21374 = pi121  & n4598;
  assign n21375 = pi122  & n4593;
  assign n21376 = n4591 & n10729;
  assign n21377 = ~n21374 & ~n21375;
  assign n21378 = ~n21373 & n21377;
  assign n21379 = ~n21376 & n21378;
  assign n21380 = pi38  & n21379;
  assign n21381 = ~pi38  & ~n21379;
  assign n21382 = ~n21380 & ~n21381;
  assign n21383 = n21372 & ~n21382;
  assign n21384 = ~n21372 & n21382;
  assign n21385 = ~n21383 & ~n21384;
  assign n21386 = n21227 & ~n21385;
  assign n21387 = ~n21227 & n21385;
  assign n21388 = ~n21386 & ~n21387;
  assign n21389 = pi123  & n4176;
  assign n21390 = pi124  & n3938;
  assign n21391 = pi125  & n3933;
  assign n21392 = n3931 & n11786;
  assign n21393 = ~n21390 & ~n21391;
  assign n21394 = ~n21389 & n21393;
  assign n21395 = ~n21392 & n21394;
  assign n21396 = pi35  & n21395;
  assign n21397 = ~pi35  & ~n21395;
  assign n21398 = ~n21396 & ~n21397;
  assign n21399 = n21388 & ~n21398;
  assign n21400 = ~n21388 & n21398;
  assign n21401 = ~n21399 & ~n21400;
  assign n21402 = n21226 & n21401;
  assign n21403 = ~n21226 & ~n21401;
  assign n21404 = ~n21402 & ~n21403;
  assign n21405 = ~n21214 & n21404;
  assign n21406 = n21214 & ~n21404;
  assign n21407 = ~n21405 & ~n21406;
  assign n21408 = ~n21213 & n21407;
  assign n21409 = n21213 & ~n21407;
  assign po94  = ~n21408 & ~n21409;
  assign n21411 = ~n21405 & ~n21408;
  assign n21412 = ~n21224 & ~n21402;
  assign n21413 = ~n21387 & ~n21399;
  assign n21414 = n3327 & ~n12539;
  assign n21415 = ~n3553 & ~n21414;
  assign n21416 = pi127  & ~n21415;
  assign n21417 = pi32  & ~n21416;
  assign n21418 = ~pi32  & n21416;
  assign n21419 = ~n21417 & ~n21418;
  assign n21420 = ~n21413 & ~n21419;
  assign n21421 = n21413 & n21419;
  assign n21422 = ~n21420 & ~n21421;
  assign n21423 = ~n21364 & ~n21367;
  assign n21424 = pi118  & n5558;
  assign n21425 = pi119  & n5293;
  assign n21426 = pi120  & n5288;
  assign n21427 = n5286 & n10047;
  assign n21428 = ~n21425 & ~n21426;
  assign n21429 = ~n21424 & n21428;
  assign n21430 = ~n21427 & n21429;
  assign n21431 = pi41  & n21430;
  assign n21432 = ~pi41  & ~n21430;
  assign n21433 = ~n21431 & ~n21432;
  assign n21434 = pi115  & n6331;
  assign n21435 = pi116  & n6015;
  assign n21436 = pi117  & n6010;
  assign n21437 = n6008 & n8784;
  assign n21438 = ~n21435 & ~n21436;
  assign n21439 = ~n21434 & n21438;
  assign n21440 = ~n21437 & n21439;
  assign n21441 = pi44  & n21440;
  assign n21442 = ~pi44  & ~n21440;
  assign n21443 = ~n21441 & ~n21442;
  assign n21444 = pi106  & n8905;
  assign n21445 = pi107  & n8535;
  assign n21446 = pi108  & n8530;
  assign n21447 = n6213 & n8528;
  assign n21448 = ~n21445 & ~n21446;
  assign n21449 = ~n21444 & n21448;
  assign n21450 = ~n21447 & n21449;
  assign n21451 = pi53  & n21450;
  assign n21452 = ~pi53  & ~n21450;
  assign n21453 = ~n21451 & ~n21452;
  assign n21454 = ~n21292 & ~n21295;
  assign n21455 = pi103  & n9858;
  assign n21456 = pi104  & n9508;
  assign n21457 = pi105  & n9503;
  assign n21458 = n5677 & n9501;
  assign n21459 = ~n21456 & ~n21457;
  assign n21460 = ~n21455 & n21459;
  assign n21461 = ~n21458 & n21460;
  assign n21462 = pi56  & n21461;
  assign n21463 = ~pi56  & ~n21461;
  assign n21464 = ~n21462 & ~n21463;
  assign n21465 = ~n21286 & ~n21289;
  assign n21466 = pi100  & n10886;
  assign n21467 = pi101  & n10495;
  assign n21468 = pi102  & n10490;
  assign n21469 = n4956 & n10488;
  assign n21470 = ~n21467 & ~n21468;
  assign n21471 = ~n21466 & n21470;
  assign n21472 = ~n21469 & n21471;
  assign n21473 = pi59  & n21472;
  assign n21474 = ~pi59  & ~n21472;
  assign n21475 = ~n21473 & ~n21474;
  assign n21476 = ~n21271 & ~n21284;
  assign n21477 = pi96  & n12277;
  assign n21478 = pi95  & n12276;
  assign n21479 = ~n21477 & ~n21478;
  assign n21480 = ~n21269 & n21479;
  assign n21481 = n21269 & ~n21479;
  assign n21482 = ~n21480 & ~n21481;
  assign n21483 = ~n21476 & n21482;
  assign n21484 = n21476 & ~n21482;
  assign n21485 = ~n21483 & ~n21484;
  assign n21486 = pi97  & n11910;
  assign n21487 = pi98  & n11529;
  assign n21488 = pi99  & n11524;
  assign n21489 = n4101 & n11522;
  assign n21490 = ~n21487 & ~n21488;
  assign n21491 = ~n21486 & n21490;
  assign n21492 = ~n21489 & n21491;
  assign n21493 = pi62  & n21492;
  assign n21494 = ~pi62  & ~n21492;
  assign n21495 = ~n21493 & ~n21494;
  assign n21496 = n21485 & ~n21495;
  assign n21497 = ~n21485 & n21495;
  assign n21498 = ~n21496 & ~n21497;
  assign n21499 = ~n21475 & n21498;
  assign n21500 = n21475 & ~n21498;
  assign n21501 = ~n21499 & ~n21500;
  assign n21502 = ~n21465 & n21501;
  assign n21503 = n21465 & ~n21501;
  assign n21504 = ~n21502 & ~n21503;
  assign n21505 = ~n21464 & n21504;
  assign n21506 = n21464 & ~n21504;
  assign n21507 = ~n21505 & ~n21506;
  assign n21508 = ~n21454 & n21507;
  assign n21509 = n21454 & ~n21507;
  assign n21510 = ~n21508 & ~n21509;
  assign n21511 = ~n21453 & n21510;
  assign n21512 = n21453 & ~n21510;
  assign n21513 = ~n21511 & ~n21512;
  assign n21514 = ~n21298 & n21310;
  assign n21515 = ~n21299 & ~n21514;
  assign n21516 = n21513 & n21515;
  assign n21517 = ~n21513 & ~n21515;
  assign n21518 = ~n21516 & ~n21517;
  assign n21519 = pi109  & n7969;
  assign n21520 = pi110  & n7636;
  assign n21521 = pi111  & n7631;
  assign n21522 = n7272 & n7629;
  assign n21523 = ~n21520 & ~n21521;
  assign n21524 = ~n21519 & n21523;
  assign n21525 = ~n21522 & n21524;
  assign n21526 = pi50  & n21525;
  assign n21527 = ~pi50  & ~n21525;
  assign n21528 = ~n21526 & ~n21527;
  assign n21529 = n21518 & ~n21528;
  assign n21530 = ~n21518 & n21528;
  assign n21531 = ~n21529 & ~n21530;
  assign n21532 = ~n21315 & n21326;
  assign n21533 = ~n21314 & ~n21532;
  assign n21534 = ~n21531 & ~n21533;
  assign n21535 = n21531 & n21533;
  assign n21536 = ~n21534 & ~n21535;
  assign n21537 = pi112  & n7121;
  assign n21538 = pi113  & n6795;
  assign n21539 = pi114  & n6790;
  assign n21540 = n6788 & n8146;
  assign n21541 = ~n21538 & ~n21539;
  assign n21542 = ~n21537 & n21541;
  assign n21543 = ~n21540 & n21542;
  assign n21544 = pi47  & n21543;
  assign n21545 = ~pi47  & ~n21543;
  assign n21546 = ~n21544 & ~n21545;
  assign n21547 = ~n21536 & n21546;
  assign n21548 = n21536 & ~n21546;
  assign n21549 = ~n21547 & ~n21548;
  assign n21550 = ~n21331 & n21342;
  assign n21551 = ~n21330 & ~n21550;
  assign n21552 = n21549 & n21551;
  assign n21553 = ~n21549 & ~n21551;
  assign n21554 = ~n21552 & ~n21553;
  assign n21555 = ~n21443 & n21554;
  assign n21556 = n21443 & ~n21554;
  assign n21557 = ~n21555 & ~n21556;
  assign n21558 = ~n21347 & n21358;
  assign n21559 = ~n21346 & ~n21558;
  assign n21560 = n21557 & n21559;
  assign n21561 = ~n21557 & ~n21559;
  assign n21562 = ~n21560 & ~n21561;
  assign n21563 = ~n21433 & n21562;
  assign n21564 = n21433 & ~n21562;
  assign n21565 = ~n21563 & ~n21564;
  assign n21566 = ~n21423 & n21565;
  assign n21567 = n21423 & ~n21565;
  assign n21568 = ~n21566 & ~n21567;
  assign n21569 = pi121  & n4843;
  assign n21570 = pi122  & n4598;
  assign n21571 = pi123  & n4593;
  assign n21572 = n4591 & n10754;
  assign n21573 = ~n21570 & ~n21571;
  assign n21574 = ~n21569 & n21573;
  assign n21575 = ~n21572 & n21574;
  assign n21576 = pi38  & n21575;
  assign n21577 = ~pi38  & ~n21575;
  assign n21578 = ~n21576 & ~n21577;
  assign n21579 = n21568 & ~n21578;
  assign n21580 = ~n21568 & n21578;
  assign n21581 = ~n21579 & ~n21580;
  assign n21582 = ~n21370 & n21382;
  assign n21583 = ~n21371 & ~n21582;
  assign n21584 = ~n21581 & ~n21583;
  assign n21585 = n21581 & n21583;
  assign n21586 = ~n21584 & ~n21585;
  assign n21587 = pi124  & n4176;
  assign n21588 = pi125  & n3938;
  assign n21589 = pi126  & n3933;
  assign n21590 = n3931 & n12148;
  assign n21591 = ~n21588 & ~n21589;
  assign n21592 = ~n21587 & n21591;
  assign n21593 = ~n21590 & n21592;
  assign n21594 = pi35  & n21593;
  assign n21595 = ~pi35  & ~n21593;
  assign n21596 = ~n21594 & ~n21595;
  assign n21597 = n21586 & ~n21596;
  assign n21598 = ~n21586 & n21596;
  assign n21599 = ~n21597 & ~n21598;
  assign n21600 = n21422 & n21599;
  assign n21601 = ~n21422 & ~n21599;
  assign n21602 = ~n21600 & ~n21601;
  assign n21603 = ~n21412 & n21602;
  assign n21604 = n21412 & ~n21602;
  assign n21605 = ~n21603 & ~n21604;
  assign n21606 = ~n21411 & n21605;
  assign n21607 = n21411 & ~n21605;
  assign po95  = ~n21606 & ~n21607;
  assign n21609 = ~n21603 & ~n21606;
  assign n21610 = ~n21420 & ~n21600;
  assign n21611 = ~n21560 & ~n21563;
  assign n21612 = ~n21552 & ~n21555;
  assign n21613 = pi116  & n6331;
  assign n21614 = pi117  & n6015;
  assign n21615 = pi118  & n6010;
  assign n21616 = n6008 & n9095;
  assign n21617 = ~n21614 & ~n21615;
  assign n21618 = ~n21613 & n21617;
  assign n21619 = ~n21616 & n21618;
  assign n21620 = pi44  & n21619;
  assign n21621 = ~pi44  & ~n21619;
  assign n21622 = ~n21620 & ~n21621;
  assign n21623 = ~n21535 & ~n21548;
  assign n21624 = ~n21508 & ~n21511;
  assign n21625 = ~n21502 & ~n21505;
  assign n21626 = ~n21496 & ~n21499;
  assign n21627 = pi101  & n10886;
  assign n21628 = pi102  & n10495;
  assign n21629 = pi103  & n10490;
  assign n21630 = n5188 & n10488;
  assign n21631 = ~n21628 & ~n21629;
  assign n21632 = ~n21627 & n21631;
  assign n21633 = ~n21630 & n21632;
  assign n21634 = pi59  & n21633;
  assign n21635 = ~pi59  & ~n21633;
  assign n21636 = ~n21634 & ~n21635;
  assign n21637 = pi98  & n11910;
  assign n21638 = pi99  & n11529;
  assign n21639 = pi100  & n11524;
  assign n21640 = n4501 & n11522;
  assign n21641 = ~n21638 & ~n21639;
  assign n21642 = ~n21637 & n21641;
  assign n21643 = ~n21640 & n21642;
  assign n21644 = pi62  & n21643;
  assign n21645 = ~pi62  & ~n21643;
  assign n21646 = ~n21644 & ~n21645;
  assign n21647 = ~n21480 & ~n21483;
  assign n21648 = pi97  & n12277;
  assign n21649 = pi96  & n12276;
  assign n21650 = ~n21648 & ~n21649;
  assign n21651 = ~pi32  & ~n21650;
  assign n21652 = pi32  & n21650;
  assign n21653 = ~n21651 & ~n21652;
  assign n21654 = ~n21479 & n21653;
  assign n21655 = n21479 & ~n21653;
  assign n21656 = ~n21654 & ~n21655;
  assign n21657 = ~n21647 & n21656;
  assign n21658 = n21647 & ~n21656;
  assign n21659 = ~n21657 & ~n21658;
  assign n21660 = ~n21646 & n21659;
  assign n21661 = n21646 & ~n21659;
  assign n21662 = ~n21660 & ~n21661;
  assign n21663 = ~n21636 & n21662;
  assign n21664 = n21636 & ~n21662;
  assign n21665 = ~n21663 & ~n21664;
  assign n21666 = ~n21626 & n21665;
  assign n21667 = n21626 & ~n21665;
  assign n21668 = ~n21666 & ~n21667;
  assign n21669 = pi104  & n9858;
  assign n21670 = pi105  & n9508;
  assign n21671 = pi106  & n9503;
  assign n21672 = n5701 & n9501;
  assign n21673 = ~n21670 & ~n21671;
  assign n21674 = ~n21669 & n21673;
  assign n21675 = ~n21672 & n21674;
  assign n21676 = pi56  & n21675;
  assign n21677 = ~pi56  & ~n21675;
  assign n21678 = ~n21676 & ~n21677;
  assign n21679 = n21668 & ~n21678;
  assign n21680 = ~n21668 & n21678;
  assign n21681 = ~n21679 & ~n21680;
  assign n21682 = n21625 & ~n21681;
  assign n21683 = ~n21625 & n21681;
  assign n21684 = ~n21682 & ~n21683;
  assign n21685 = pi107  & n8905;
  assign n21686 = pi108  & n8535;
  assign n21687 = pi109  & n8530;
  assign n21688 = n6715 & n8528;
  assign n21689 = ~n21686 & ~n21687;
  assign n21690 = ~n21685 & n21689;
  assign n21691 = ~n21688 & n21690;
  assign n21692 = pi53  & n21691;
  assign n21693 = ~pi53  & ~n21691;
  assign n21694 = ~n21692 & ~n21693;
  assign n21695 = n21684 & ~n21694;
  assign n21696 = ~n21684 & n21694;
  assign n21697 = ~n21695 & ~n21696;
  assign n21698 = n21624 & ~n21697;
  assign n21699 = ~n21624 & n21697;
  assign n21700 = ~n21698 & ~n21699;
  assign n21701 = pi110  & n7969;
  assign n21702 = pi111  & n7636;
  assign n21703 = pi112  & n7631;
  assign n21704 = n7296 & n7629;
  assign n21705 = ~n21702 & ~n21703;
  assign n21706 = ~n21701 & n21705;
  assign n21707 = ~n21704 & n21706;
  assign n21708 = pi50  & n21707;
  assign n21709 = ~pi50  & ~n21707;
  assign n21710 = ~n21708 & ~n21709;
  assign n21711 = n21700 & ~n21710;
  assign n21712 = ~n21700 & n21710;
  assign n21713 = ~n21711 & ~n21712;
  assign n21714 = ~n21516 & n21528;
  assign n21715 = ~n21517 & ~n21714;
  assign n21716 = ~n21713 & ~n21715;
  assign n21717 = n21713 & n21715;
  assign n21718 = ~n21716 & ~n21717;
  assign n21719 = pi113  & n7121;
  assign n21720 = pi114  & n6795;
  assign n21721 = pi115  & n6790;
  assign n21722 = n6788 & n8170;
  assign n21723 = ~n21720 & ~n21721;
  assign n21724 = ~n21719 & n21723;
  assign n21725 = ~n21722 & n21724;
  assign n21726 = pi47  & n21725;
  assign n21727 = ~pi47  & ~n21725;
  assign n21728 = ~n21726 & ~n21727;
  assign n21729 = n21718 & ~n21728;
  assign n21730 = ~n21718 & n21728;
  assign n21731 = ~n21729 & ~n21730;
  assign n21732 = n21623 & n21731;
  assign n21733 = ~n21623 & ~n21731;
  assign n21734 = ~n21732 & ~n21733;
  assign n21735 = n21622 & n21734;
  assign n21736 = ~n21622 & ~n21734;
  assign n21737 = ~n21735 & ~n21736;
  assign n21738 = ~n21612 & n21737;
  assign n21739 = n21612 & ~n21737;
  assign n21740 = ~n21738 & ~n21739;
  assign n21741 = pi119  & n5558;
  assign n21742 = pi120  & n5293;
  assign n21743 = pi121  & n5288;
  assign n21744 = n5286 & n10071;
  assign n21745 = ~n21742 & ~n21743;
  assign n21746 = ~n21741 & n21745;
  assign n21747 = ~n21744 & n21746;
  assign n21748 = pi41  & n21747;
  assign n21749 = ~pi41  & ~n21747;
  assign n21750 = ~n21748 & ~n21749;
  assign n21751 = n21740 & ~n21750;
  assign n21752 = ~n21740 & n21750;
  assign n21753 = ~n21751 & ~n21752;
  assign n21754 = n21611 & ~n21753;
  assign n21755 = ~n21611 & n21753;
  assign n21756 = ~n21754 & ~n21755;
  assign n21757 = pi122  & n4843;
  assign n21758 = pi123  & n4598;
  assign n21759 = pi124  & n4593;
  assign n21760 = n4591 & n11099;
  assign n21761 = ~n21758 & ~n21759;
  assign n21762 = ~n21757 & n21761;
  assign n21763 = ~n21760 & n21762;
  assign n21764 = pi38  & n21763;
  assign n21765 = ~pi38  & ~n21763;
  assign n21766 = ~n21764 & ~n21765;
  assign n21767 = n21756 & ~n21766;
  assign n21768 = ~n21756 & n21766;
  assign n21769 = ~n21767 & ~n21768;
  assign n21770 = ~n21566 & n21578;
  assign n21771 = ~n21567 & ~n21770;
  assign n21772 = ~n21769 & ~n21771;
  assign n21773 = n21769 & n21771;
  assign n21774 = ~n21772 & ~n21773;
  assign n21775 = pi125  & n4176;
  assign n21776 = pi126  & n3938;
  assign n21777 = pi127  & n3933;
  assign n21778 = n3931 & n12519;
  assign n21779 = ~n21776 & ~n21777;
  assign n21780 = ~n21775 & n21779;
  assign n21781 = ~n21778 & n21780;
  assign n21782 = pi35  & n21781;
  assign n21783 = ~pi35  & ~n21781;
  assign n21784 = ~n21782 & ~n21783;
  assign n21785 = ~n21585 & n21596;
  assign n21786 = ~n21584 & ~n21785;
  assign n21787 = ~n21784 & n21786;
  assign n21788 = n21784 & ~n21786;
  assign n21789 = ~n21787 & ~n21788;
  assign n21790 = ~n21774 & ~n21789;
  assign n21791 = n21774 & n21789;
  assign n21792 = ~n21790 & ~n21791;
  assign n21793 = ~n21610 & n21792;
  assign n21794 = n21610 & ~n21792;
  assign n21795 = ~n21793 & ~n21794;
  assign n21796 = ~n21609 & n21795;
  assign n21797 = n21609 & ~n21795;
  assign po96  = ~n21796 & ~n21797;
  assign n21799 = ~n21793 & ~n21796;
  assign n21800 = ~n21787 & ~n21791;
  assign n21801 = ~n21767 & ~n21773;
  assign n21802 = pi126  & n4176;
  assign n21803 = pi127  & n3938;
  assign n21804 = n3931 & n12542;
  assign n21805 = ~n21802 & ~n21803;
  assign n21806 = ~n21804 & n21805;
  assign n21807 = pi35  & n21806;
  assign n21808 = ~pi35  & ~n21806;
  assign n21809 = ~n21807 & ~n21808;
  assign n21810 = ~n21801 & ~n21809;
  assign n21811 = n21801 & n21809;
  assign n21812 = ~n21810 & ~n21811;
  assign n21813 = ~n21751 & ~n21755;
  assign n21814 = ~n21736 & ~n21738;
  assign n21815 = pi117  & n6331;
  assign n21816 = pi118  & n6015;
  assign n21817 = pi119  & n6010;
  assign n21818 = n6008 & n9412;
  assign n21819 = ~n21816 & ~n21817;
  assign n21820 = ~n21815 & n21819;
  assign n21821 = ~n21818 & n21820;
  assign n21822 = pi44  & n21821;
  assign n21823 = ~pi44  & ~n21821;
  assign n21824 = ~n21822 & ~n21823;
  assign n21825 = ~n21711 & ~n21717;
  assign n21826 = ~n21695 & ~n21699;
  assign n21827 = ~n21679 & ~n21683;
  assign n21828 = ~n21663 & ~n21666;
  assign n21829 = pi102  & n10886;
  assign n21830 = pi103  & n10495;
  assign n21831 = pi104  & n10490;
  assign n21832 = n5212 & n10488;
  assign n21833 = ~n21830 & ~n21831;
  assign n21834 = ~n21829 & n21833;
  assign n21835 = ~n21832 & n21834;
  assign n21836 = pi59  & n21835;
  assign n21837 = ~pi59  & ~n21835;
  assign n21838 = ~n21836 & ~n21837;
  assign n21839 = ~n21657 & ~n21660;
  assign n21840 = ~n21479 & ~n21652;
  assign n21841 = ~n21651 & ~n21840;
  assign n21842 = pi98  & n12277;
  assign n21843 = pi97  & n12276;
  assign n21844 = ~n21842 & ~n21843;
  assign n21845 = n21841 & ~n21844;
  assign n21846 = ~n21841 & n21844;
  assign n21847 = ~n21845 & ~n21846;
  assign n21848 = pi99  & n11910;
  assign n21849 = pi100  & n11529;
  assign n21850 = pi101  & n11524;
  assign n21851 = n4730 & n11522;
  assign n21852 = ~n21849 & ~n21850;
  assign n21853 = ~n21848 & n21852;
  assign n21854 = ~n21851 & n21853;
  assign n21855 = pi62  & n21854;
  assign n21856 = ~pi62  & ~n21854;
  assign n21857 = ~n21855 & ~n21856;
  assign n21858 = ~n21847 & n21857;
  assign n21859 = n21847 & ~n21857;
  assign n21860 = ~n21858 & ~n21859;
  assign n21861 = ~n21839 & n21860;
  assign n21862 = n21839 & ~n21860;
  assign n21863 = ~n21861 & ~n21862;
  assign n21864 = ~n21838 & n21863;
  assign n21865 = n21838 & ~n21863;
  assign n21866 = ~n21864 & ~n21865;
  assign n21867 = ~n21828 & n21866;
  assign n21868 = n21828 & ~n21866;
  assign n21869 = ~n21867 & ~n21868;
  assign n21870 = pi105  & n9858;
  assign n21871 = pi106  & n9508;
  assign n21872 = pi107  & n9503;
  assign n21873 = n6189 & n9501;
  assign n21874 = ~n21871 & ~n21872;
  assign n21875 = ~n21870 & n21874;
  assign n21876 = ~n21873 & n21875;
  assign n21877 = pi56  & n21876;
  assign n21878 = ~pi56  & ~n21876;
  assign n21879 = ~n21877 & ~n21878;
  assign n21880 = n21869 & ~n21879;
  assign n21881 = ~n21869 & n21879;
  assign n21882 = ~n21880 & ~n21881;
  assign n21883 = n21827 & ~n21882;
  assign n21884 = ~n21827 & n21882;
  assign n21885 = ~n21883 & ~n21884;
  assign n21886 = pi108  & n8905;
  assign n21887 = pi109  & n8535;
  assign n21888 = pi110  & n8530;
  assign n21889 = n6995 & n8528;
  assign n21890 = ~n21887 & ~n21888;
  assign n21891 = ~n21886 & n21890;
  assign n21892 = ~n21889 & n21891;
  assign n21893 = pi53  & n21892;
  assign n21894 = ~pi53  & ~n21892;
  assign n21895 = ~n21893 & ~n21894;
  assign n21896 = n21885 & ~n21895;
  assign n21897 = ~n21885 & n21895;
  assign n21898 = ~n21896 & ~n21897;
  assign n21899 = n21826 & ~n21898;
  assign n21900 = ~n21826 & n21898;
  assign n21901 = ~n21899 & ~n21900;
  assign n21902 = pi111  & n7969;
  assign n21903 = pi112  & n7636;
  assign n21904 = pi113  & n7631;
  assign n21905 = n7629 & n7852;
  assign n21906 = ~n21903 & ~n21904;
  assign n21907 = ~n21902 & n21906;
  assign n21908 = ~n21905 & n21907;
  assign n21909 = pi50  & n21908;
  assign n21910 = ~pi50  & ~n21908;
  assign n21911 = ~n21909 & ~n21910;
  assign n21912 = n21901 & ~n21911;
  assign n21913 = ~n21901 & n21911;
  assign n21914 = ~n21912 & ~n21913;
  assign n21915 = n21825 & ~n21914;
  assign n21916 = ~n21825 & n21914;
  assign n21917 = ~n21915 & ~n21916;
  assign n21918 = pi114  & n7121;
  assign n21919 = pi115  & n6795;
  assign n21920 = pi116  & n6790;
  assign n21921 = n6788 & n8470;
  assign n21922 = ~n21919 & ~n21920;
  assign n21923 = ~n21918 & n21922;
  assign n21924 = ~n21921 & n21923;
  assign n21925 = pi47  & n21924;
  assign n21926 = ~pi47  & ~n21924;
  assign n21927 = ~n21925 & ~n21926;
  assign n21928 = n21917 & ~n21927;
  assign n21929 = ~n21917 & n21927;
  assign n21930 = ~n21928 & ~n21929;
  assign n21931 = n21623 & ~n21729;
  assign n21932 = ~n21730 & ~n21931;
  assign n21933 = n21930 & n21932;
  assign n21934 = ~n21930 & ~n21932;
  assign n21935 = ~n21933 & ~n21934;
  assign n21936 = ~n21824 & n21935;
  assign n21937 = n21824 & ~n21935;
  assign n21938 = ~n21936 & ~n21937;
  assign n21939 = ~n21814 & n21938;
  assign n21940 = n21814 & ~n21938;
  assign n21941 = ~n21939 & ~n21940;
  assign n21942 = pi120  & n5558;
  assign n21943 = pi121  & n5293;
  assign n21944 = pi122  & n5288;
  assign n21945 = n5286 & n10729;
  assign n21946 = ~n21943 & ~n21944;
  assign n21947 = ~n21942 & n21946;
  assign n21948 = ~n21945 & n21947;
  assign n21949 = pi41  & n21948;
  assign n21950 = ~pi41  & ~n21948;
  assign n21951 = ~n21949 & ~n21950;
  assign n21952 = n21941 & ~n21951;
  assign n21953 = ~n21941 & n21951;
  assign n21954 = ~n21952 & ~n21953;
  assign n21955 = n21813 & ~n21954;
  assign n21956 = ~n21813 & n21954;
  assign n21957 = ~n21955 & ~n21956;
  assign n21958 = pi123  & n4843;
  assign n21959 = pi124  & n4598;
  assign n21960 = pi125  & n4593;
  assign n21961 = n4591 & n11786;
  assign n21962 = ~n21959 & ~n21960;
  assign n21963 = ~n21958 & n21962;
  assign n21964 = ~n21961 & n21963;
  assign n21965 = pi38  & n21964;
  assign n21966 = ~pi38  & ~n21964;
  assign n21967 = ~n21965 & ~n21966;
  assign n21968 = n21957 & ~n21967;
  assign n21969 = ~n21957 & n21967;
  assign n21970 = ~n21968 & ~n21969;
  assign n21971 = n21812 & n21970;
  assign n21972 = ~n21812 & ~n21970;
  assign n21973 = ~n21971 & ~n21972;
  assign n21974 = ~n21800 & n21973;
  assign n21975 = n21800 & ~n21973;
  assign n21976 = ~n21974 & ~n21975;
  assign n21977 = ~n21799 & n21976;
  assign n21978 = n21799 & ~n21976;
  assign po97  = ~n21977 & ~n21978;
  assign n21980 = ~n21974 & ~n21977;
  assign n21981 = ~n21810 & ~n21971;
  assign n21982 = ~n21956 & ~n21968;
  assign n21983 = n3931 & ~n12539;
  assign n21984 = ~n4176 & ~n21983;
  assign n21985 = pi127  & ~n21984;
  assign n21986 = pi35  & ~n21985;
  assign n21987 = ~pi35  & n21985;
  assign n21988 = ~n21986 & ~n21987;
  assign n21989 = ~n21982 & ~n21988;
  assign n21990 = n21982 & n21988;
  assign n21991 = ~n21989 & ~n21990;
  assign n21992 = ~n21933 & ~n21936;
  assign n21993 = pi118  & n6331;
  assign n21994 = pi119  & n6015;
  assign n21995 = pi120  & n6010;
  assign n21996 = n6008 & n10047;
  assign n21997 = ~n21994 & ~n21995;
  assign n21998 = ~n21993 & n21997;
  assign n21999 = ~n21996 & n21998;
  assign n22000 = pi44  & n21999;
  assign n22001 = ~pi44  & ~n21999;
  assign n22002 = ~n22000 & ~n22001;
  assign n22003 = pi115  & n7121;
  assign n22004 = pi116  & n6795;
  assign n22005 = pi117  & n6790;
  assign n22006 = n6788 & n8784;
  assign n22007 = ~n22004 & ~n22005;
  assign n22008 = ~n22003 & n22007;
  assign n22009 = ~n22006 & n22008;
  assign n22010 = pi47  & n22009;
  assign n22011 = ~pi47  & ~n22009;
  assign n22012 = ~n22010 & ~n22011;
  assign n22013 = pi106  & n9858;
  assign n22014 = pi107  & n9508;
  assign n22015 = pi108  & n9503;
  assign n22016 = n6213 & n9501;
  assign n22017 = ~n22014 & ~n22015;
  assign n22018 = ~n22013 & n22017;
  assign n22019 = ~n22016 & n22018;
  assign n22020 = pi56  & n22019;
  assign n22021 = ~pi56  & ~n22019;
  assign n22022 = ~n22020 & ~n22021;
  assign n22023 = ~n21861 & ~n21864;
  assign n22024 = pi103  & n10886;
  assign n22025 = pi104  & n10495;
  assign n22026 = pi105  & n10490;
  assign n22027 = n5677 & n10488;
  assign n22028 = ~n22025 & ~n22026;
  assign n22029 = ~n22024 & n22028;
  assign n22030 = ~n22027 & n22029;
  assign n22031 = pi59  & n22030;
  assign n22032 = ~pi59  & ~n22030;
  assign n22033 = ~n22031 & ~n22032;
  assign n22034 = ~n21846 & ~n21859;
  assign n22035 = pi99  & n12277;
  assign n22036 = pi98  & n12276;
  assign n22037 = ~n22035 & ~n22036;
  assign n22038 = ~n21844 & n22037;
  assign n22039 = n21844 & ~n22037;
  assign n22040 = ~n22038 & ~n22039;
  assign n22041 = ~n22034 & n22040;
  assign n22042 = n22034 & ~n22040;
  assign n22043 = ~n22041 & ~n22042;
  assign n22044 = pi100  & n11910;
  assign n22045 = pi101  & n11529;
  assign n22046 = pi102  & n11524;
  assign n22047 = n4956 & n11522;
  assign n22048 = ~n22045 & ~n22046;
  assign n22049 = ~n22044 & n22048;
  assign n22050 = ~n22047 & n22049;
  assign n22051 = pi62  & n22050;
  assign n22052 = ~pi62  & ~n22050;
  assign n22053 = ~n22051 & ~n22052;
  assign n22054 = n22043 & ~n22053;
  assign n22055 = ~n22043 & n22053;
  assign n22056 = ~n22054 & ~n22055;
  assign n22057 = ~n22033 & n22056;
  assign n22058 = n22033 & ~n22056;
  assign n22059 = ~n22057 & ~n22058;
  assign n22060 = ~n22023 & n22059;
  assign n22061 = n22023 & ~n22059;
  assign n22062 = ~n22060 & ~n22061;
  assign n22063 = ~n22022 & n22062;
  assign n22064 = n22022 & ~n22062;
  assign n22065 = ~n22063 & ~n22064;
  assign n22066 = ~n21867 & n21879;
  assign n22067 = ~n21868 & ~n22066;
  assign n22068 = n22065 & n22067;
  assign n22069 = ~n22065 & ~n22067;
  assign n22070 = ~n22068 & ~n22069;
  assign n22071 = pi109  & n8905;
  assign n22072 = pi110  & n8535;
  assign n22073 = pi111  & n8530;
  assign n22074 = n7272 & n8528;
  assign n22075 = ~n22072 & ~n22073;
  assign n22076 = ~n22071 & n22075;
  assign n22077 = ~n22074 & n22076;
  assign n22078 = pi53  & n22077;
  assign n22079 = ~pi53  & ~n22077;
  assign n22080 = ~n22078 & ~n22079;
  assign n22081 = n22070 & ~n22080;
  assign n22082 = ~n22070 & n22080;
  assign n22083 = ~n22081 & ~n22082;
  assign n22084 = ~n21884 & n21895;
  assign n22085 = ~n21883 & ~n22084;
  assign n22086 = ~n22083 & ~n22085;
  assign n22087 = n22083 & n22085;
  assign n22088 = ~n22086 & ~n22087;
  assign n22089 = pi112  & n7969;
  assign n22090 = pi113  & n7636;
  assign n22091 = pi114  & n7631;
  assign n22092 = n7629 & n8146;
  assign n22093 = ~n22090 & ~n22091;
  assign n22094 = ~n22089 & n22093;
  assign n22095 = ~n22092 & n22094;
  assign n22096 = pi50  & n22095;
  assign n22097 = ~pi50  & ~n22095;
  assign n22098 = ~n22096 & ~n22097;
  assign n22099 = ~n22088 & n22098;
  assign n22100 = n22088 & ~n22098;
  assign n22101 = ~n22099 & ~n22100;
  assign n22102 = ~n21900 & n21911;
  assign n22103 = ~n21899 & ~n22102;
  assign n22104 = n22101 & n22103;
  assign n22105 = ~n22101 & ~n22103;
  assign n22106 = ~n22104 & ~n22105;
  assign n22107 = ~n22012 & n22106;
  assign n22108 = n22012 & ~n22106;
  assign n22109 = ~n22107 & ~n22108;
  assign n22110 = ~n21916 & n21927;
  assign n22111 = ~n21915 & ~n22110;
  assign n22112 = n22109 & n22111;
  assign n22113 = ~n22109 & ~n22111;
  assign n22114 = ~n22112 & ~n22113;
  assign n22115 = ~n22002 & n22114;
  assign n22116 = n22002 & ~n22114;
  assign n22117 = ~n22115 & ~n22116;
  assign n22118 = ~n21992 & n22117;
  assign n22119 = n21992 & ~n22117;
  assign n22120 = ~n22118 & ~n22119;
  assign n22121 = pi121  & n5558;
  assign n22122 = pi122  & n5293;
  assign n22123 = pi123  & n5288;
  assign n22124 = n5286 & n10754;
  assign n22125 = ~n22122 & ~n22123;
  assign n22126 = ~n22121 & n22125;
  assign n22127 = ~n22124 & n22126;
  assign n22128 = pi41  & n22127;
  assign n22129 = ~pi41  & ~n22127;
  assign n22130 = ~n22128 & ~n22129;
  assign n22131 = n22120 & ~n22130;
  assign n22132 = ~n22120 & n22130;
  assign n22133 = ~n22131 & ~n22132;
  assign n22134 = ~n21939 & n21951;
  assign n22135 = ~n21940 & ~n22134;
  assign n22136 = ~n22133 & ~n22135;
  assign n22137 = n22133 & n22135;
  assign n22138 = ~n22136 & ~n22137;
  assign n22139 = pi124  & n4843;
  assign n22140 = pi125  & n4598;
  assign n22141 = pi126  & n4593;
  assign n22142 = n4591 & n12148;
  assign n22143 = ~n22140 & ~n22141;
  assign n22144 = ~n22139 & n22143;
  assign n22145 = ~n22142 & n22144;
  assign n22146 = pi38  & n22145;
  assign n22147 = ~pi38  & ~n22145;
  assign n22148 = ~n22146 & ~n22147;
  assign n22149 = n22138 & ~n22148;
  assign n22150 = ~n22138 & n22148;
  assign n22151 = ~n22149 & ~n22150;
  assign n22152 = n21991 & n22151;
  assign n22153 = ~n21991 & ~n22151;
  assign n22154 = ~n22152 & ~n22153;
  assign n22155 = ~n21981 & n22154;
  assign n22156 = n21981 & ~n22154;
  assign n22157 = ~n22155 & ~n22156;
  assign n22158 = ~n21980 & n22157;
  assign n22159 = n21980 & ~n22157;
  assign po98  = ~n22158 & ~n22159;
  assign n22161 = ~n22155 & ~n22158;
  assign n22162 = ~n22112 & ~n22115;
  assign n22163 = ~n22104 & ~n22107;
  assign n22164 = pi116  & n7121;
  assign n22165 = pi117  & n6795;
  assign n22166 = pi118  & n6790;
  assign n22167 = n6788 & n9095;
  assign n22168 = ~n22165 & ~n22166;
  assign n22169 = ~n22164 & n22168;
  assign n22170 = ~n22167 & n22169;
  assign n22171 = pi47  & n22170;
  assign n22172 = ~pi47  & ~n22170;
  assign n22173 = ~n22171 & ~n22172;
  assign n22174 = ~n22087 & ~n22100;
  assign n22175 = ~n22060 & ~n22063;
  assign n22176 = pi107  & n9858;
  assign n22177 = pi108  & n9508;
  assign n22178 = pi109  & n9503;
  assign n22179 = n6715 & n9501;
  assign n22180 = ~n22177 & ~n22178;
  assign n22181 = ~n22176 & n22180;
  assign n22182 = ~n22179 & n22181;
  assign n22183 = pi56  & n22182;
  assign n22184 = ~pi56  & ~n22182;
  assign n22185 = ~n22183 & ~n22184;
  assign n22186 = ~n22054 & ~n22057;
  assign n22187 = ~n22038 & ~n22041;
  assign n22188 = ~pi35  & ~n22037;
  assign n22189 = pi35  & n22037;
  assign n22190 = ~n22188 & ~n22189;
  assign n22191 = pi100  & n12277;
  assign n22192 = pi99  & n12276;
  assign n22193 = ~n22191 & ~n22192;
  assign n22194 = n22190 & ~n22193;
  assign n22195 = ~n22190 & n22193;
  assign n22196 = ~n22194 & ~n22195;
  assign n22197 = ~n22187 & n22196;
  assign n22198 = n22187 & ~n22196;
  assign n22199 = ~n22197 & ~n22198;
  assign n22200 = pi101  & n11910;
  assign n22201 = pi102  & n11529;
  assign n22202 = pi103  & n11524;
  assign n22203 = n5188 & n11522;
  assign n22204 = ~n22201 & ~n22202;
  assign n22205 = ~n22200 & n22204;
  assign n22206 = ~n22203 & n22205;
  assign n22207 = pi62  & n22206;
  assign n22208 = ~pi62  & ~n22206;
  assign n22209 = ~n22207 & ~n22208;
  assign n22210 = ~n22199 & n22209;
  assign n22211 = n22199 & ~n22209;
  assign n22212 = ~n22210 & ~n22211;
  assign n22213 = pi104  & n10886;
  assign n22214 = pi105  & n10495;
  assign n22215 = pi106  & n10490;
  assign n22216 = n5701 & n10488;
  assign n22217 = ~n22214 & ~n22215;
  assign n22218 = ~n22213 & n22217;
  assign n22219 = ~n22216 & n22218;
  assign n22220 = pi59  & n22219;
  assign n22221 = ~pi59  & ~n22219;
  assign n22222 = ~n22220 & ~n22221;
  assign n22223 = n22212 & ~n22222;
  assign n22224 = ~n22212 & n22222;
  assign n22225 = ~n22223 & ~n22224;
  assign n22226 = ~n22186 & n22225;
  assign n22227 = n22186 & ~n22225;
  assign n22228 = ~n22226 & ~n22227;
  assign n22229 = ~n22185 & n22228;
  assign n22230 = n22185 & ~n22228;
  assign n22231 = ~n22229 & ~n22230;
  assign n22232 = n22175 & ~n22231;
  assign n22233 = ~n22175 & n22231;
  assign n22234 = ~n22232 & ~n22233;
  assign n22235 = pi110  & n8905;
  assign n22236 = pi111  & n8535;
  assign n22237 = pi112  & n8530;
  assign n22238 = n7296 & n8528;
  assign n22239 = ~n22236 & ~n22237;
  assign n22240 = ~n22235 & n22239;
  assign n22241 = ~n22238 & n22240;
  assign n22242 = pi53  & n22241;
  assign n22243 = ~pi53  & ~n22241;
  assign n22244 = ~n22242 & ~n22243;
  assign n22245 = n22234 & ~n22244;
  assign n22246 = ~n22234 & n22244;
  assign n22247 = ~n22245 & ~n22246;
  assign n22248 = ~n22068 & n22080;
  assign n22249 = ~n22069 & ~n22248;
  assign n22250 = ~n22247 & ~n22249;
  assign n22251 = n22247 & n22249;
  assign n22252 = ~n22250 & ~n22251;
  assign n22253 = pi113  & n7969;
  assign n22254 = pi114  & n7636;
  assign n22255 = pi115  & n7631;
  assign n22256 = n7629 & n8170;
  assign n22257 = ~n22254 & ~n22255;
  assign n22258 = ~n22253 & n22257;
  assign n22259 = ~n22256 & n22258;
  assign n22260 = pi50  & n22259;
  assign n22261 = ~pi50  & ~n22259;
  assign n22262 = ~n22260 & ~n22261;
  assign n22263 = ~n22252 & n22262;
  assign n22264 = n22252 & ~n22262;
  assign n22265 = ~n22263 & ~n22264;
  assign n22266 = ~n22174 & n22265;
  assign n22267 = n22174 & ~n22265;
  assign n22268 = ~n22266 & ~n22267;
  assign n22269 = ~n22173 & n22268;
  assign n22270 = n22173 & ~n22268;
  assign n22271 = ~n22269 & ~n22270;
  assign n22272 = ~n22163 & n22271;
  assign n22273 = n22163 & ~n22271;
  assign n22274 = ~n22272 & ~n22273;
  assign n22275 = pi119  & n6331;
  assign n22276 = pi120  & n6015;
  assign n22277 = pi121  & n6010;
  assign n22278 = n6008 & n10071;
  assign n22279 = ~n22276 & ~n22277;
  assign n22280 = ~n22275 & n22279;
  assign n22281 = ~n22278 & n22280;
  assign n22282 = pi44  & n22281;
  assign n22283 = ~pi44  & ~n22281;
  assign n22284 = ~n22282 & ~n22283;
  assign n22285 = n22274 & ~n22284;
  assign n22286 = ~n22274 & n22284;
  assign n22287 = ~n22285 & ~n22286;
  assign n22288 = n22162 & ~n22287;
  assign n22289 = ~n22162 & n22287;
  assign n22290 = ~n22288 & ~n22289;
  assign n22291 = pi122  & n5558;
  assign n22292 = pi123  & n5293;
  assign n22293 = pi124  & n5288;
  assign n22294 = n5286 & n11099;
  assign n22295 = ~n22292 & ~n22293;
  assign n22296 = ~n22291 & n22295;
  assign n22297 = ~n22294 & n22296;
  assign n22298 = pi41  & n22297;
  assign n22299 = ~pi41  & ~n22297;
  assign n22300 = ~n22298 & ~n22299;
  assign n22301 = n22290 & ~n22300;
  assign n22302 = ~n22290 & n22300;
  assign n22303 = ~n22301 & ~n22302;
  assign n22304 = ~n22118 & n22130;
  assign n22305 = ~n22119 & ~n22304;
  assign n22306 = ~n22303 & ~n22305;
  assign n22307 = n22303 & n22305;
  assign n22308 = ~n22306 & ~n22307;
  assign n22309 = pi125  & n4843;
  assign n22310 = pi126  & n4598;
  assign n22311 = pi127  & n4593;
  assign n22312 = n4591 & n12519;
  assign n22313 = ~n22310 & ~n22311;
  assign n22314 = ~n22309 & n22313;
  assign n22315 = ~n22312 & n22314;
  assign n22316 = pi38  & n22315;
  assign n22317 = ~pi38  & ~n22315;
  assign n22318 = ~n22316 & ~n22317;
  assign n22319 = n22308 & ~n22318;
  assign n22320 = ~n22308 & n22318;
  assign n22321 = ~n22319 & ~n22320;
  assign n22322 = ~n22137 & n22148;
  assign n22323 = ~n22136 & ~n22322;
  assign n22324 = ~n22321 & ~n22323;
  assign n22325 = n22321 & n22323;
  assign n22326 = ~n22324 & ~n22325;
  assign n22327 = ~n21989 & ~n22152;
  assign n22328 = n22326 & ~n22327;
  assign n22329 = ~n22326 & n22327;
  assign n22330 = ~n22328 & ~n22329;
  assign n22331 = ~n22161 & n22330;
  assign n22332 = n22161 & ~n22330;
  assign po99  = ~n22331 & ~n22332;
  assign n22334 = ~n22319 & ~n22325;
  assign n22335 = ~n22301 & ~n22307;
  assign n22336 = pi126  & n4843;
  assign n22337 = pi127  & n4598;
  assign n22338 = n4591 & n12542;
  assign n22339 = ~n22336 & ~n22337;
  assign n22340 = ~n22338 & n22339;
  assign n22341 = pi38  & n22340;
  assign n22342 = ~pi38  & ~n22340;
  assign n22343 = ~n22341 & ~n22342;
  assign n22344 = ~n22335 & ~n22343;
  assign n22345 = n22335 & n22343;
  assign n22346 = ~n22344 & ~n22345;
  assign n22347 = ~n22285 & ~n22289;
  assign n22348 = ~n22269 & ~n22272;
  assign n22349 = pi117  & n7121;
  assign n22350 = pi118  & n6795;
  assign n22351 = pi119  & n6790;
  assign n22352 = n6788 & n9412;
  assign n22353 = ~n22350 & ~n22351;
  assign n22354 = ~n22349 & n22353;
  assign n22355 = ~n22352 & n22354;
  assign n22356 = pi47  & n22355;
  assign n22357 = ~pi47  & ~n22355;
  assign n22358 = ~n22356 & ~n22357;
  assign n22359 = ~n22264 & ~n22266;
  assign n22360 = ~n22245 & ~n22251;
  assign n22361 = ~n22229 & ~n22233;
  assign n22362 = ~n22223 & ~n22226;
  assign n22363 = ~n22197 & ~n22211;
  assign n22364 = pi102  & n11910;
  assign n22365 = pi103  & n11529;
  assign n22366 = pi104  & n11524;
  assign n22367 = n5212 & n11522;
  assign n22368 = ~n22365 & ~n22366;
  assign n22369 = ~n22364 & n22368;
  assign n22370 = ~n22367 & n22369;
  assign n22371 = pi62  & n22370;
  assign n22372 = ~pi62  & ~n22370;
  assign n22373 = ~n22371 & ~n22372;
  assign n22374 = ~n22188 & ~n22194;
  assign n22375 = pi101  & n12277;
  assign n22376 = pi100  & n12276;
  assign n22377 = ~n22375 & ~n22376;
  assign n22378 = ~n22374 & n22377;
  assign n22379 = n22374 & ~n22377;
  assign n22380 = ~n22378 & ~n22379;
  assign n22381 = n22373 & ~n22380;
  assign n22382 = ~n22373 & n22380;
  assign n22383 = ~n22381 & ~n22382;
  assign n22384 = n22363 & ~n22383;
  assign n22385 = ~n22363 & n22383;
  assign n22386 = ~n22384 & ~n22385;
  assign n22387 = pi105  & n10886;
  assign n22388 = pi106  & n10495;
  assign n22389 = pi107  & n10490;
  assign n22390 = n6189 & n10488;
  assign n22391 = ~n22388 & ~n22389;
  assign n22392 = ~n22387 & n22391;
  assign n22393 = ~n22390 & n22392;
  assign n22394 = pi59  & n22393;
  assign n22395 = ~pi59  & ~n22393;
  assign n22396 = ~n22394 & ~n22395;
  assign n22397 = n22386 & ~n22396;
  assign n22398 = ~n22386 & n22396;
  assign n22399 = ~n22397 & ~n22398;
  assign n22400 = n22362 & ~n22399;
  assign n22401 = ~n22362 & n22399;
  assign n22402 = ~n22400 & ~n22401;
  assign n22403 = pi108  & n9858;
  assign n22404 = pi109  & n9508;
  assign n22405 = pi110  & n9503;
  assign n22406 = n6995 & n9501;
  assign n22407 = ~n22404 & ~n22405;
  assign n22408 = ~n22403 & n22407;
  assign n22409 = ~n22406 & n22408;
  assign n22410 = pi56  & n22409;
  assign n22411 = ~pi56  & ~n22409;
  assign n22412 = ~n22410 & ~n22411;
  assign n22413 = n22402 & ~n22412;
  assign n22414 = ~n22402 & n22412;
  assign n22415 = ~n22413 & ~n22414;
  assign n22416 = n22361 & ~n22415;
  assign n22417 = ~n22361 & n22415;
  assign n22418 = ~n22416 & ~n22417;
  assign n22419 = pi111  & n8905;
  assign n22420 = pi112  & n8535;
  assign n22421 = pi113  & n8530;
  assign n22422 = n7852 & n8528;
  assign n22423 = ~n22420 & ~n22421;
  assign n22424 = ~n22419 & n22423;
  assign n22425 = ~n22422 & n22424;
  assign n22426 = pi53  & n22425;
  assign n22427 = ~pi53  & ~n22425;
  assign n22428 = ~n22426 & ~n22427;
  assign n22429 = n22418 & ~n22428;
  assign n22430 = ~n22418 & n22428;
  assign n22431 = ~n22429 & ~n22430;
  assign n22432 = n22360 & ~n22431;
  assign n22433 = ~n22360 & n22431;
  assign n22434 = ~n22432 & ~n22433;
  assign n22435 = pi114  & n7969;
  assign n22436 = pi115  & n7636;
  assign n22437 = pi116  & n7631;
  assign n22438 = n7629 & n8470;
  assign n22439 = ~n22436 & ~n22437;
  assign n22440 = ~n22435 & n22439;
  assign n22441 = ~n22438 & n22440;
  assign n22442 = pi50  & n22441;
  assign n22443 = ~pi50  & ~n22441;
  assign n22444 = ~n22442 & ~n22443;
  assign n22445 = n22434 & ~n22444;
  assign n22446 = ~n22434 & n22444;
  assign n22447 = ~n22445 & ~n22446;
  assign n22448 = ~n22359 & n22447;
  assign n22449 = n22359 & ~n22447;
  assign n22450 = ~n22448 & ~n22449;
  assign n22451 = ~n22358 & n22450;
  assign n22452 = n22358 & ~n22450;
  assign n22453 = ~n22451 & ~n22452;
  assign n22454 = n22348 & ~n22453;
  assign n22455 = ~n22348 & n22453;
  assign n22456 = ~n22454 & ~n22455;
  assign n22457 = pi120  & n6331;
  assign n22458 = pi121  & n6015;
  assign n22459 = pi122  & n6010;
  assign n22460 = n6008 & n10729;
  assign n22461 = ~n22458 & ~n22459;
  assign n22462 = ~n22457 & n22461;
  assign n22463 = ~n22460 & n22462;
  assign n22464 = pi44  & n22463;
  assign n22465 = ~pi44  & ~n22463;
  assign n22466 = ~n22464 & ~n22465;
  assign n22467 = n22456 & ~n22466;
  assign n22468 = ~n22456 & n22466;
  assign n22469 = ~n22467 & ~n22468;
  assign n22470 = n22347 & ~n22469;
  assign n22471 = ~n22347 & n22469;
  assign n22472 = ~n22470 & ~n22471;
  assign n22473 = pi123  & n5558;
  assign n22474 = pi124  & n5293;
  assign n22475 = pi125  & n5288;
  assign n22476 = n5286 & n11786;
  assign n22477 = ~n22474 & ~n22475;
  assign n22478 = ~n22473 & n22477;
  assign n22479 = ~n22476 & n22478;
  assign n22480 = pi41  & n22479;
  assign n22481 = ~pi41  & ~n22479;
  assign n22482 = ~n22480 & ~n22481;
  assign n22483 = n22472 & ~n22482;
  assign n22484 = ~n22472 & n22482;
  assign n22485 = ~n22483 & ~n22484;
  assign n22486 = n22346 & n22485;
  assign n22487 = ~n22346 & ~n22485;
  assign n22488 = ~n22486 & ~n22487;
  assign n22489 = n22334 & ~n22488;
  assign n22490 = ~n22334 & n22488;
  assign n22491 = ~n22489 & ~n22490;
  assign n22492 = ~n22328 & ~n22331;
  assign n22493 = n22491 & ~n22492;
  assign n22494 = ~n22491 & n22492;
  assign po100  = ~n22493 & ~n22494;
  assign n22496 = ~n22490 & ~n22493;
  assign n22497 = ~n22344 & ~n22486;
  assign n22498 = ~n22471 & ~n22483;
  assign n22499 = n4591 & ~n12539;
  assign n22500 = ~n4843 & ~n22499;
  assign n22501 = pi127  & ~n22500;
  assign n22502 = pi38  & ~n22501;
  assign n22503 = ~pi38  & n22501;
  assign n22504 = ~n22502 & ~n22503;
  assign n22505 = ~n22498 & ~n22504;
  assign n22506 = n22498 & n22504;
  assign n22507 = ~n22505 & ~n22506;
  assign n22508 = ~n22448 & ~n22451;
  assign n22509 = pi118  & n7121;
  assign n22510 = pi119  & n6795;
  assign n22511 = pi120  & n6790;
  assign n22512 = n6788 & n10047;
  assign n22513 = ~n22510 & ~n22511;
  assign n22514 = ~n22509 & n22513;
  assign n22515 = ~n22512 & n22514;
  assign n22516 = pi47  & n22515;
  assign n22517 = ~pi47  & ~n22515;
  assign n22518 = ~n22516 & ~n22517;
  assign n22519 = pi115  & n7969;
  assign n22520 = pi116  & n7636;
  assign n22521 = pi117  & n7631;
  assign n22522 = n7629 & n8784;
  assign n22523 = ~n22520 & ~n22521;
  assign n22524 = ~n22519 & n22523;
  assign n22525 = ~n22522 & n22524;
  assign n22526 = pi50  & n22525;
  assign n22527 = ~pi50  & ~n22525;
  assign n22528 = ~n22526 & ~n22527;
  assign n22529 = pi106  & n10886;
  assign n22530 = pi107  & n10495;
  assign n22531 = pi108  & n10490;
  assign n22532 = n6213 & n10488;
  assign n22533 = ~n22530 & ~n22531;
  assign n22534 = ~n22529 & n22533;
  assign n22535 = ~n22532 & n22534;
  assign n22536 = pi59  & n22535;
  assign n22537 = ~pi59  & ~n22535;
  assign n22538 = ~n22536 & ~n22537;
  assign n22539 = pi103  & n11910;
  assign n22540 = pi104  & n11529;
  assign n22541 = pi105  & n11524;
  assign n22542 = n5677 & n11522;
  assign n22543 = ~n22540 & ~n22541;
  assign n22544 = ~n22539 & n22543;
  assign n22545 = ~n22542 & n22544;
  assign n22546 = pi62  & n22545;
  assign n22547 = ~pi62  & ~n22545;
  assign n22548 = ~n22546 & ~n22547;
  assign n22549 = pi102  & n12277;
  assign n22550 = pi101  & n12276;
  assign n22551 = ~n22549 & ~n22550;
  assign n22552 = n22377 & ~n22551;
  assign n22553 = ~n22377 & n22551;
  assign n22554 = ~n22552 & ~n22553;
  assign n22555 = n22373 & ~n22378;
  assign n22556 = ~n22379 & ~n22555;
  assign n22557 = n22554 & n22556;
  assign n22558 = ~n22554 & ~n22556;
  assign n22559 = ~n22557 & ~n22558;
  assign n22560 = ~n22548 & n22559;
  assign n22561 = n22548 & ~n22559;
  assign n22562 = ~n22560 & ~n22561;
  assign n22563 = ~n22538 & n22562;
  assign n22564 = n22538 & ~n22562;
  assign n22565 = ~n22563 & ~n22564;
  assign n22566 = ~n22385 & n22396;
  assign n22567 = ~n22384 & ~n22566;
  assign n22568 = ~n22565 & ~n22567;
  assign n22569 = n22565 & n22567;
  assign n22570 = ~n22568 & ~n22569;
  assign n22571 = pi109  & n9858;
  assign n22572 = pi110  & n9508;
  assign n22573 = pi111  & n9503;
  assign n22574 = n7272 & n9501;
  assign n22575 = ~n22572 & ~n22573;
  assign n22576 = ~n22571 & n22575;
  assign n22577 = ~n22574 & n22576;
  assign n22578 = pi56  & n22577;
  assign n22579 = ~pi56  & ~n22577;
  assign n22580 = ~n22578 & ~n22579;
  assign n22581 = n22570 & ~n22580;
  assign n22582 = ~n22570 & n22580;
  assign n22583 = ~n22581 & ~n22582;
  assign n22584 = ~n22401 & n22412;
  assign n22585 = ~n22400 & ~n22584;
  assign n22586 = ~n22583 & ~n22585;
  assign n22587 = n22583 & n22585;
  assign n22588 = ~n22586 & ~n22587;
  assign n22589 = pi112  & n8905;
  assign n22590 = pi113  & n8535;
  assign n22591 = pi114  & n8530;
  assign n22592 = n8146 & n8528;
  assign n22593 = ~n22590 & ~n22591;
  assign n22594 = ~n22589 & n22593;
  assign n22595 = ~n22592 & n22594;
  assign n22596 = pi53  & n22595;
  assign n22597 = ~pi53  & ~n22595;
  assign n22598 = ~n22596 & ~n22597;
  assign n22599 = ~n22588 & n22598;
  assign n22600 = n22588 & ~n22598;
  assign n22601 = ~n22599 & ~n22600;
  assign n22602 = ~n22417 & n22428;
  assign n22603 = ~n22416 & ~n22602;
  assign n22604 = n22601 & n22603;
  assign n22605 = ~n22601 & ~n22603;
  assign n22606 = ~n22604 & ~n22605;
  assign n22607 = ~n22528 & n22606;
  assign n22608 = n22528 & ~n22606;
  assign n22609 = ~n22607 & ~n22608;
  assign n22610 = ~n22433 & n22444;
  assign n22611 = ~n22432 & ~n22610;
  assign n22612 = n22609 & n22611;
  assign n22613 = ~n22609 & ~n22611;
  assign n22614 = ~n22612 & ~n22613;
  assign n22615 = ~n22518 & n22614;
  assign n22616 = n22518 & ~n22614;
  assign n22617 = ~n22615 & ~n22616;
  assign n22618 = ~n22508 & n22617;
  assign n22619 = n22508 & ~n22617;
  assign n22620 = ~n22618 & ~n22619;
  assign n22621 = pi121  & n6331;
  assign n22622 = pi122  & n6015;
  assign n22623 = pi123  & n6010;
  assign n22624 = n6008 & n10754;
  assign n22625 = ~n22622 & ~n22623;
  assign n22626 = ~n22621 & n22625;
  assign n22627 = ~n22624 & n22626;
  assign n22628 = pi44  & n22627;
  assign n22629 = ~pi44  & ~n22627;
  assign n22630 = ~n22628 & ~n22629;
  assign n22631 = n22620 & ~n22630;
  assign n22632 = ~n22620 & n22630;
  assign n22633 = ~n22631 & ~n22632;
  assign n22634 = ~n22455 & n22466;
  assign n22635 = ~n22454 & ~n22634;
  assign n22636 = ~n22633 & ~n22635;
  assign n22637 = n22633 & n22635;
  assign n22638 = ~n22636 & ~n22637;
  assign n22639 = pi124  & n5558;
  assign n22640 = pi125  & n5293;
  assign n22641 = pi126  & n5288;
  assign n22642 = n5286 & n12148;
  assign n22643 = ~n22640 & ~n22641;
  assign n22644 = ~n22639 & n22643;
  assign n22645 = ~n22642 & n22644;
  assign n22646 = pi41  & n22645;
  assign n22647 = ~pi41  & ~n22645;
  assign n22648 = ~n22646 & ~n22647;
  assign n22649 = n22638 & ~n22648;
  assign n22650 = ~n22638 & n22648;
  assign n22651 = ~n22649 & ~n22650;
  assign n22652 = n22507 & n22651;
  assign n22653 = ~n22507 & ~n22651;
  assign n22654 = ~n22652 & ~n22653;
  assign n22655 = ~n22497 & n22654;
  assign n22656 = n22497 & ~n22654;
  assign n22657 = ~n22655 & ~n22656;
  assign n22658 = ~n22496 & n22657;
  assign n22659 = n22496 & ~n22657;
  assign po101  = ~n22658 & ~n22659;
  assign n22661 = ~n22655 & ~n22658;
  assign n22662 = ~n22612 & ~n22615;
  assign n22663 = ~n22604 & ~n22607;
  assign n22664 = pi116  & n7969;
  assign n22665 = pi117  & n7636;
  assign n22666 = pi118  & n7631;
  assign n22667 = n7629 & n9095;
  assign n22668 = ~n22665 & ~n22666;
  assign n22669 = ~n22664 & n22668;
  assign n22670 = ~n22667 & n22669;
  assign n22671 = pi50  & n22670;
  assign n22672 = ~pi50  & ~n22670;
  assign n22673 = ~n22671 & ~n22672;
  assign n22674 = ~n22587 & ~n22600;
  assign n22675 = pi110  & n9858;
  assign n22676 = pi111  & n9508;
  assign n22677 = pi112  & n9503;
  assign n22678 = n7296 & n9501;
  assign n22679 = ~n22676 & ~n22677;
  assign n22680 = ~n22675 & n22679;
  assign n22681 = ~n22678 & n22680;
  assign n22682 = pi56  & n22681;
  assign n22683 = ~pi56  & ~n22681;
  assign n22684 = ~n22682 & ~n22683;
  assign n22685 = ~n22560 & ~n22563;
  assign n22686 = pi107  & n10886;
  assign n22687 = pi108  & n10495;
  assign n22688 = pi109  & n10490;
  assign n22689 = n6715 & n10488;
  assign n22690 = ~n22687 & ~n22688;
  assign n22691 = ~n22686 & n22690;
  assign n22692 = ~n22689 & n22691;
  assign n22693 = pi59  & n22692;
  assign n22694 = ~pi59  & ~n22692;
  assign n22695 = ~n22693 & ~n22694;
  assign n22696 = ~n22552 & ~n22557;
  assign n22697 = ~pi38  & ~n22377;
  assign n22698 = pi38  & n22377;
  assign n22699 = ~n22697 & ~n22698;
  assign n22700 = pi103  & n12277;
  assign n22701 = pi102  & n12276;
  assign n22702 = ~n22700 & ~n22701;
  assign n22703 = n22699 & ~n22702;
  assign n22704 = ~n22699 & n22702;
  assign n22705 = ~n22703 & ~n22704;
  assign n22706 = ~n22696 & n22705;
  assign n22707 = n22696 & ~n22705;
  assign n22708 = ~n22706 & ~n22707;
  assign n22709 = pi104  & n11910;
  assign n22710 = pi105  & n11529;
  assign n22711 = pi106  & n11524;
  assign n22712 = n5701 & n11522;
  assign n22713 = ~n22710 & ~n22711;
  assign n22714 = ~n22709 & n22713;
  assign n22715 = ~n22712 & n22714;
  assign n22716 = pi62  & n22715;
  assign n22717 = ~pi62  & ~n22715;
  assign n22718 = ~n22716 & ~n22717;
  assign n22719 = n22708 & ~n22718;
  assign n22720 = ~n22708 & n22718;
  assign n22721 = ~n22719 & ~n22720;
  assign n22722 = ~n22695 & n22721;
  assign n22723 = n22695 & ~n22721;
  assign n22724 = ~n22722 & ~n22723;
  assign n22725 = ~n22685 & n22724;
  assign n22726 = n22685 & ~n22724;
  assign n22727 = ~n22725 & ~n22726;
  assign n22728 = ~n22684 & n22727;
  assign n22729 = n22684 & ~n22727;
  assign n22730 = ~n22728 & ~n22729;
  assign n22731 = ~n22569 & n22580;
  assign n22732 = ~n22568 & ~n22731;
  assign n22733 = ~n22730 & ~n22732;
  assign n22734 = n22730 & n22732;
  assign n22735 = ~n22733 & ~n22734;
  assign n22736 = pi113  & n8905;
  assign n22737 = pi114  & n8535;
  assign n22738 = pi115  & n8530;
  assign n22739 = n8170 & n8528;
  assign n22740 = ~n22737 & ~n22738;
  assign n22741 = ~n22736 & n22740;
  assign n22742 = ~n22739 & n22741;
  assign n22743 = pi53  & n22742;
  assign n22744 = ~pi53  & ~n22742;
  assign n22745 = ~n22743 & ~n22744;
  assign n22746 = ~n22735 & n22745;
  assign n22747 = n22735 & ~n22745;
  assign n22748 = ~n22746 & ~n22747;
  assign n22749 = ~n22674 & n22748;
  assign n22750 = n22674 & ~n22748;
  assign n22751 = ~n22749 & ~n22750;
  assign n22752 = ~n22673 & n22751;
  assign n22753 = n22673 & ~n22751;
  assign n22754 = ~n22752 & ~n22753;
  assign n22755 = ~n22663 & n22754;
  assign n22756 = n22663 & ~n22754;
  assign n22757 = ~n22755 & ~n22756;
  assign n22758 = pi119  & n7121;
  assign n22759 = pi120  & n6795;
  assign n22760 = pi121  & n6790;
  assign n22761 = n6788 & n10071;
  assign n22762 = ~n22759 & ~n22760;
  assign n22763 = ~n22758 & n22762;
  assign n22764 = ~n22761 & n22763;
  assign n22765 = pi47  & n22764;
  assign n22766 = ~pi47  & ~n22764;
  assign n22767 = ~n22765 & ~n22766;
  assign n22768 = n22757 & ~n22767;
  assign n22769 = ~n22757 & n22767;
  assign n22770 = ~n22768 & ~n22769;
  assign n22771 = n22662 & ~n22770;
  assign n22772 = ~n22662 & n22770;
  assign n22773 = ~n22771 & ~n22772;
  assign n22774 = pi122  & n6331;
  assign n22775 = pi123  & n6015;
  assign n22776 = pi124  & n6010;
  assign n22777 = n6008 & n11099;
  assign n22778 = ~n22775 & ~n22776;
  assign n22779 = ~n22774 & n22778;
  assign n22780 = ~n22777 & n22779;
  assign n22781 = pi44  & n22780;
  assign n22782 = ~pi44  & ~n22780;
  assign n22783 = ~n22781 & ~n22782;
  assign n22784 = n22773 & ~n22783;
  assign n22785 = ~n22773 & n22783;
  assign n22786 = ~n22784 & ~n22785;
  assign n22787 = ~n22618 & n22630;
  assign n22788 = ~n22619 & ~n22787;
  assign n22789 = ~n22786 & ~n22788;
  assign n22790 = n22786 & n22788;
  assign n22791 = ~n22789 & ~n22790;
  assign n22792 = pi125  & n5558;
  assign n22793 = pi126  & n5293;
  assign n22794 = pi127  & n5288;
  assign n22795 = n5286 & n12519;
  assign n22796 = ~n22793 & ~n22794;
  assign n22797 = ~n22792 & n22796;
  assign n22798 = ~n22795 & n22797;
  assign n22799 = pi41  & n22798;
  assign n22800 = ~pi41  & ~n22798;
  assign n22801 = ~n22799 & ~n22800;
  assign n22802 = n22791 & ~n22801;
  assign n22803 = ~n22791 & n22801;
  assign n22804 = ~n22802 & ~n22803;
  assign n22805 = ~n22637 & n22648;
  assign n22806 = ~n22636 & ~n22805;
  assign n22807 = ~n22804 & ~n22806;
  assign n22808 = n22804 & n22806;
  assign n22809 = ~n22807 & ~n22808;
  assign n22810 = ~n22505 & ~n22652;
  assign n22811 = n22809 & ~n22810;
  assign n22812 = ~n22809 & n22810;
  assign n22813 = ~n22811 & ~n22812;
  assign n22814 = ~n22661 & n22813;
  assign n22815 = n22661 & ~n22813;
  assign po102  = ~n22814 & ~n22815;
  assign n22817 = ~n22802 & ~n22808;
  assign n22818 = ~n22784 & ~n22790;
  assign n22819 = pi126  & n5558;
  assign n22820 = pi127  & n5293;
  assign n22821 = n5286 & n12542;
  assign n22822 = ~n22819 & ~n22820;
  assign n22823 = ~n22821 & n22822;
  assign n22824 = pi41  & n22823;
  assign n22825 = ~pi41  & ~n22823;
  assign n22826 = ~n22824 & ~n22825;
  assign n22827 = ~n22818 & ~n22826;
  assign n22828 = n22818 & n22826;
  assign n22829 = ~n22827 & ~n22828;
  assign n22830 = ~n22768 & ~n22772;
  assign n22831 = ~n22752 & ~n22755;
  assign n22832 = pi117  & n7969;
  assign n22833 = pi118  & n7636;
  assign n22834 = pi119  & n7631;
  assign n22835 = n7629 & n9412;
  assign n22836 = ~n22833 & ~n22834;
  assign n22837 = ~n22832 & n22836;
  assign n22838 = ~n22835 & n22837;
  assign n22839 = pi50  & n22838;
  assign n22840 = ~pi50  & ~n22838;
  assign n22841 = ~n22839 & ~n22840;
  assign n22842 = ~n22747 & ~n22749;
  assign n22843 = ~n22728 & ~n22734;
  assign n22844 = ~n22722 & ~n22725;
  assign n22845 = ~n22697 & ~n22703;
  assign n22846 = pi104  & n12277;
  assign n22847 = pi103  & n12276;
  assign n22848 = ~n22846 & ~n22847;
  assign n22849 = ~n22845 & n22848;
  assign n22850 = n22845 & ~n22848;
  assign n22851 = ~n22849 & ~n22850;
  assign n22852 = pi105  & n11910;
  assign n22853 = pi106  & n11529;
  assign n22854 = pi107  & n11524;
  assign n22855 = n6189 & n11522;
  assign n22856 = ~n22853 & ~n22854;
  assign n22857 = ~n22852 & n22856;
  assign n22858 = ~n22855 & n22857;
  assign n22859 = pi62  & n22858;
  assign n22860 = ~pi62  & ~n22858;
  assign n22861 = ~n22859 & ~n22860;
  assign n22862 = n22851 & ~n22861;
  assign n22863 = ~n22851 & n22861;
  assign n22864 = ~n22862 & ~n22863;
  assign n22865 = ~n22706 & n22718;
  assign n22866 = ~n22707 & ~n22865;
  assign n22867 = n22864 & n22866;
  assign n22868 = ~n22864 & ~n22866;
  assign n22869 = ~n22867 & ~n22868;
  assign n22870 = pi108  & n10886;
  assign n22871 = pi109  & n10495;
  assign n22872 = pi110  & n10490;
  assign n22873 = n6995 & n10488;
  assign n22874 = ~n22871 & ~n22872;
  assign n22875 = ~n22870 & n22874;
  assign n22876 = ~n22873 & n22875;
  assign n22877 = pi59  & n22876;
  assign n22878 = ~pi59  & ~n22876;
  assign n22879 = ~n22877 & ~n22878;
  assign n22880 = n22869 & ~n22879;
  assign n22881 = ~n22869 & n22879;
  assign n22882 = ~n22880 & ~n22881;
  assign n22883 = n22844 & ~n22882;
  assign n22884 = ~n22844 & n22882;
  assign n22885 = ~n22883 & ~n22884;
  assign n22886 = pi111  & n9858;
  assign n22887 = pi112  & n9508;
  assign n22888 = pi113  & n9503;
  assign n22889 = n7852 & n9501;
  assign n22890 = ~n22887 & ~n22888;
  assign n22891 = ~n22886 & n22890;
  assign n22892 = ~n22889 & n22891;
  assign n22893 = pi56  & n22892;
  assign n22894 = ~pi56  & ~n22892;
  assign n22895 = ~n22893 & ~n22894;
  assign n22896 = n22885 & ~n22895;
  assign n22897 = ~n22885 & n22895;
  assign n22898 = ~n22896 & ~n22897;
  assign n22899 = n22843 & ~n22898;
  assign n22900 = ~n22843 & n22898;
  assign n22901 = ~n22899 & ~n22900;
  assign n22902 = pi114  & n8905;
  assign n22903 = pi115  & n8535;
  assign n22904 = pi116  & n8530;
  assign n22905 = n8470 & n8528;
  assign n22906 = ~n22903 & ~n22904;
  assign n22907 = ~n22902 & n22906;
  assign n22908 = ~n22905 & n22907;
  assign n22909 = pi53  & n22908;
  assign n22910 = ~pi53  & ~n22908;
  assign n22911 = ~n22909 & ~n22910;
  assign n22912 = n22901 & ~n22911;
  assign n22913 = ~n22901 & n22911;
  assign n22914 = ~n22912 & ~n22913;
  assign n22915 = ~n22842 & n22914;
  assign n22916 = n22842 & ~n22914;
  assign n22917 = ~n22915 & ~n22916;
  assign n22918 = ~n22841 & n22917;
  assign n22919 = n22841 & ~n22917;
  assign n22920 = ~n22918 & ~n22919;
  assign n22921 = n22831 & ~n22920;
  assign n22922 = ~n22831 & n22920;
  assign n22923 = ~n22921 & ~n22922;
  assign n22924 = pi120  & n7121;
  assign n22925 = pi121  & n6795;
  assign n22926 = pi122  & n6790;
  assign n22927 = n6788 & n10729;
  assign n22928 = ~n22925 & ~n22926;
  assign n22929 = ~n22924 & n22928;
  assign n22930 = ~n22927 & n22929;
  assign n22931 = pi47  & n22930;
  assign n22932 = ~pi47  & ~n22930;
  assign n22933 = ~n22931 & ~n22932;
  assign n22934 = n22923 & ~n22933;
  assign n22935 = ~n22923 & n22933;
  assign n22936 = ~n22934 & ~n22935;
  assign n22937 = n22830 & ~n22936;
  assign n22938 = ~n22830 & n22936;
  assign n22939 = ~n22937 & ~n22938;
  assign n22940 = pi123  & n6331;
  assign n22941 = pi124  & n6015;
  assign n22942 = pi125  & n6010;
  assign n22943 = n6008 & n11786;
  assign n22944 = ~n22941 & ~n22942;
  assign n22945 = ~n22940 & n22944;
  assign n22946 = ~n22943 & n22945;
  assign n22947 = pi44  & n22946;
  assign n22948 = ~pi44  & ~n22946;
  assign n22949 = ~n22947 & ~n22948;
  assign n22950 = n22939 & ~n22949;
  assign n22951 = ~n22939 & n22949;
  assign n22952 = ~n22950 & ~n22951;
  assign n22953 = n22829 & n22952;
  assign n22954 = ~n22829 & ~n22952;
  assign n22955 = ~n22953 & ~n22954;
  assign n22956 = n22817 & ~n22955;
  assign n22957 = ~n22817 & n22955;
  assign n22958 = ~n22956 & ~n22957;
  assign n22959 = ~n22811 & ~n22814;
  assign n22960 = n22958 & ~n22959;
  assign n22961 = ~n22958 & n22959;
  assign po103  = ~n22960 & ~n22961;
  assign n22963 = ~n22957 & ~n22960;
  assign n22964 = ~n22827 & ~n22953;
  assign n22965 = ~n22938 & ~n22950;
  assign n22966 = n5286 & ~n12539;
  assign n22967 = ~n5558 & ~n22966;
  assign n22968 = pi127  & ~n22967;
  assign n22969 = pi41  & ~n22968;
  assign n22970 = ~pi41  & n22968;
  assign n22971 = ~n22969 & ~n22970;
  assign n22972 = ~n22965 & ~n22971;
  assign n22973 = n22965 & n22971;
  assign n22974 = ~n22972 & ~n22973;
  assign n22975 = ~n22915 & ~n22918;
  assign n22976 = pi118  & n7969;
  assign n22977 = pi119  & n7636;
  assign n22978 = pi120  & n7631;
  assign n22979 = n7629 & n10047;
  assign n22980 = ~n22977 & ~n22978;
  assign n22981 = ~n22976 & n22980;
  assign n22982 = ~n22979 & n22981;
  assign n22983 = pi50  & n22982;
  assign n22984 = ~pi50  & ~n22982;
  assign n22985 = ~n22983 & ~n22984;
  assign n22986 = pi115  & n8905;
  assign n22987 = pi116  & n8535;
  assign n22988 = pi117  & n8530;
  assign n22989 = n8528 & n8784;
  assign n22990 = ~n22987 & ~n22988;
  assign n22991 = ~n22986 & n22990;
  assign n22992 = ~n22989 & n22991;
  assign n22993 = pi53  & n22992;
  assign n22994 = ~pi53  & ~n22992;
  assign n22995 = ~n22993 & ~n22994;
  assign n22996 = pi109  & n10886;
  assign n22997 = pi110  & n10495;
  assign n22998 = pi111  & n10490;
  assign n22999 = n7272 & n10488;
  assign n23000 = ~n22997 & ~n22998;
  assign n23001 = ~n22996 & n23000;
  assign n23002 = ~n22999 & n23001;
  assign n23003 = pi59  & n23002;
  assign n23004 = ~pi59  & ~n23002;
  assign n23005 = ~n23003 & ~n23004;
  assign n23006 = pi106  & n11910;
  assign n23007 = pi107  & n11529;
  assign n23008 = pi108  & n11524;
  assign n23009 = n6213 & n11522;
  assign n23010 = ~n23007 & ~n23008;
  assign n23011 = ~n23006 & n23010;
  assign n23012 = ~n23009 & n23011;
  assign n23013 = pi62  & n23012;
  assign n23014 = ~pi62  & ~n23012;
  assign n23015 = ~n23013 & ~n23014;
  assign n23016 = ~n22849 & ~n22862;
  assign n23017 = pi105  & n12277;
  assign n23018 = pi104  & n12276;
  assign n23019 = ~n23017 & ~n23018;
  assign n23020 = n22848 & ~n23019;
  assign n23021 = ~n22848 & n23019;
  assign n23022 = ~n23020 & ~n23021;
  assign n23023 = ~n23016 & n23022;
  assign n23024 = n23016 & ~n23022;
  assign n23025 = ~n23023 & ~n23024;
  assign n23026 = ~n23015 & n23025;
  assign n23027 = n23015 & ~n23025;
  assign n23028 = ~n23026 & ~n23027;
  assign n23029 = ~n23005 & n23028;
  assign n23030 = n23005 & ~n23028;
  assign n23031 = ~n23029 & ~n23030;
  assign n23032 = ~n22867 & n22879;
  assign n23033 = ~n22868 & ~n23032;
  assign n23034 = ~n23031 & ~n23033;
  assign n23035 = n23031 & n23033;
  assign n23036 = ~n23034 & ~n23035;
  assign n23037 = pi112  & n9858;
  assign n23038 = pi113  & n9508;
  assign n23039 = pi114  & n9503;
  assign n23040 = n8146 & n9501;
  assign n23041 = ~n23038 & ~n23039;
  assign n23042 = ~n23037 & n23041;
  assign n23043 = ~n23040 & n23042;
  assign n23044 = pi56  & n23043;
  assign n23045 = ~pi56  & ~n23043;
  assign n23046 = ~n23044 & ~n23045;
  assign n23047 = ~n23036 & n23046;
  assign n23048 = n23036 & ~n23046;
  assign n23049 = ~n23047 & ~n23048;
  assign n23050 = ~n22884 & n22895;
  assign n23051 = ~n22883 & ~n23050;
  assign n23052 = n23049 & n23051;
  assign n23053 = ~n23049 & ~n23051;
  assign n23054 = ~n23052 & ~n23053;
  assign n23055 = ~n22995 & n23054;
  assign n23056 = n22995 & ~n23054;
  assign n23057 = ~n23055 & ~n23056;
  assign n23058 = ~n22900 & n22911;
  assign n23059 = ~n22899 & ~n23058;
  assign n23060 = n23057 & n23059;
  assign n23061 = ~n23057 & ~n23059;
  assign n23062 = ~n23060 & ~n23061;
  assign n23063 = ~n22985 & n23062;
  assign n23064 = n22985 & ~n23062;
  assign n23065 = ~n23063 & ~n23064;
  assign n23066 = ~n22975 & n23065;
  assign n23067 = n22975 & ~n23065;
  assign n23068 = ~n23066 & ~n23067;
  assign n23069 = pi121  & n7121;
  assign n23070 = pi122  & n6795;
  assign n23071 = pi123  & n6790;
  assign n23072 = n6788 & n10754;
  assign n23073 = ~n23070 & ~n23071;
  assign n23074 = ~n23069 & n23073;
  assign n23075 = ~n23072 & n23074;
  assign n23076 = pi47  & n23075;
  assign n23077 = ~pi47  & ~n23075;
  assign n23078 = ~n23076 & ~n23077;
  assign n23079 = n23068 & ~n23078;
  assign n23080 = ~n23068 & n23078;
  assign n23081 = ~n23079 & ~n23080;
  assign n23082 = ~n22922 & n22933;
  assign n23083 = ~n22921 & ~n23082;
  assign n23084 = ~n23081 & ~n23083;
  assign n23085 = n23081 & n23083;
  assign n23086 = ~n23084 & ~n23085;
  assign n23087 = pi124  & n6331;
  assign n23088 = pi125  & n6015;
  assign n23089 = pi126  & n6010;
  assign n23090 = n6008 & n12148;
  assign n23091 = ~n23088 & ~n23089;
  assign n23092 = ~n23087 & n23091;
  assign n23093 = ~n23090 & n23092;
  assign n23094 = pi44  & n23093;
  assign n23095 = ~pi44  & ~n23093;
  assign n23096 = ~n23094 & ~n23095;
  assign n23097 = n23086 & ~n23096;
  assign n23098 = ~n23086 & n23096;
  assign n23099 = ~n23097 & ~n23098;
  assign n23100 = n22974 & n23099;
  assign n23101 = ~n22974 & ~n23099;
  assign n23102 = ~n23100 & ~n23101;
  assign n23103 = ~n22964 & n23102;
  assign n23104 = n22964 & ~n23102;
  assign n23105 = ~n23103 & ~n23104;
  assign n23106 = ~n22963 & n23105;
  assign n23107 = n22963 & ~n23105;
  assign po104  = ~n23106 & ~n23107;
  assign n23109 = ~n23103 & ~n23106;
  assign n23110 = ~n23060 & ~n23063;
  assign n23111 = pi119  & n7969;
  assign n23112 = pi120  & n7636;
  assign n23113 = pi121  & n7631;
  assign n23114 = n7629 & n10071;
  assign n23115 = ~n23112 & ~n23113;
  assign n23116 = ~n23111 & n23115;
  assign n23117 = ~n23114 & n23116;
  assign n23118 = pi50  & n23117;
  assign n23119 = ~pi50  & ~n23117;
  assign n23120 = ~n23118 & ~n23119;
  assign n23121 = ~n23052 & ~n23055;
  assign n23122 = pi116  & n8905;
  assign n23123 = pi117  & n8535;
  assign n23124 = pi118  & n8530;
  assign n23125 = n8528 & n9095;
  assign n23126 = ~n23123 & ~n23124;
  assign n23127 = ~n23122 & n23126;
  assign n23128 = ~n23125 & n23127;
  assign n23129 = pi53  & n23128;
  assign n23130 = ~pi53  & ~n23128;
  assign n23131 = ~n23129 & ~n23130;
  assign n23132 = ~n23035 & ~n23048;
  assign n23133 = pi113  & n9858;
  assign n23134 = pi114  & n9508;
  assign n23135 = pi115  & n9503;
  assign n23136 = n8170 & n9501;
  assign n23137 = ~n23134 & ~n23135;
  assign n23138 = ~n23133 & n23137;
  assign n23139 = ~n23136 & n23138;
  assign n23140 = pi56  & n23139;
  assign n23141 = ~pi56  & ~n23139;
  assign n23142 = ~n23140 & ~n23141;
  assign n23143 = ~n23026 & ~n23029;
  assign n23144 = ~n23020 & ~n23023;
  assign n23145 = ~pi41  & ~n22848;
  assign n23146 = pi41  & n22848;
  assign n23147 = ~n23145 & ~n23146;
  assign n23148 = pi106  & n12277;
  assign n23149 = pi105  & n12276;
  assign n23150 = ~n23148 & ~n23149;
  assign n23151 = ~n23147 & n23150;
  assign n23152 = n23147 & ~n23150;
  assign n23153 = ~n23151 & ~n23152;
  assign n23154 = pi107  & n11910;
  assign n23155 = pi108  & n11529;
  assign n23156 = pi109  & n11524;
  assign n23157 = n6715 & n11522;
  assign n23158 = ~n23155 & ~n23156;
  assign n23159 = ~n23154 & n23158;
  assign n23160 = ~n23157 & n23159;
  assign n23161 = pi62  & n23160;
  assign n23162 = ~pi62  & ~n23160;
  assign n23163 = ~n23161 & ~n23162;
  assign n23164 = n23153 & ~n23163;
  assign n23165 = ~n23153 & n23163;
  assign n23166 = ~n23164 & ~n23165;
  assign n23167 = n23144 & ~n23166;
  assign n23168 = ~n23144 & n23166;
  assign n23169 = ~n23167 & ~n23168;
  assign n23170 = pi110  & n10886;
  assign n23171 = pi111  & n10495;
  assign n23172 = pi112  & n10490;
  assign n23173 = n7296 & n10488;
  assign n23174 = ~n23171 & ~n23172;
  assign n23175 = ~n23170 & n23174;
  assign n23176 = ~n23173 & n23175;
  assign n23177 = pi59  & n23176;
  assign n23178 = ~pi59  & ~n23176;
  assign n23179 = ~n23177 & ~n23178;
  assign n23180 = n23169 & ~n23179;
  assign n23181 = ~n23169 & n23179;
  assign n23182 = ~n23180 & ~n23181;
  assign n23183 = ~n23143 & n23182;
  assign n23184 = n23143 & ~n23182;
  assign n23185 = ~n23183 & ~n23184;
  assign n23186 = ~n23142 & n23185;
  assign n23187 = n23142 & ~n23185;
  assign n23188 = ~n23186 & ~n23187;
  assign n23189 = ~n23132 & n23188;
  assign n23190 = n23132 & ~n23188;
  assign n23191 = ~n23189 & ~n23190;
  assign n23192 = n23131 & ~n23191;
  assign n23193 = ~n23131 & n23191;
  assign n23194 = ~n23192 & ~n23193;
  assign n23195 = ~n23121 & n23194;
  assign n23196 = n23121 & ~n23194;
  assign n23197 = ~n23195 & ~n23196;
  assign n23198 = n23120 & ~n23197;
  assign n23199 = ~n23120 & n23197;
  assign n23200 = ~n23198 & ~n23199;
  assign n23201 = ~n23110 & n23200;
  assign n23202 = n23110 & ~n23200;
  assign n23203 = ~n23201 & ~n23202;
  assign n23204 = pi122  & n7121;
  assign n23205 = pi123  & n6795;
  assign n23206 = pi124  & n6790;
  assign n23207 = n6788 & n11099;
  assign n23208 = ~n23205 & ~n23206;
  assign n23209 = ~n23204 & n23208;
  assign n23210 = ~n23207 & n23209;
  assign n23211 = pi47  & n23210;
  assign n23212 = ~pi47  & ~n23210;
  assign n23213 = ~n23211 & ~n23212;
  assign n23214 = n23203 & ~n23213;
  assign n23215 = ~n23203 & n23213;
  assign n23216 = ~n23214 & ~n23215;
  assign n23217 = ~n23066 & n23078;
  assign n23218 = ~n23067 & ~n23217;
  assign n23219 = ~n23216 & ~n23218;
  assign n23220 = n23216 & n23218;
  assign n23221 = ~n23219 & ~n23220;
  assign n23222 = pi125  & n6331;
  assign n23223 = pi126  & n6015;
  assign n23224 = pi127  & n6010;
  assign n23225 = n6008 & n12519;
  assign n23226 = ~n23223 & ~n23224;
  assign n23227 = ~n23222 & n23226;
  assign n23228 = ~n23225 & n23227;
  assign n23229 = pi44  & n23228;
  assign n23230 = ~pi44  & ~n23228;
  assign n23231 = ~n23229 & ~n23230;
  assign n23232 = n23221 & ~n23231;
  assign n23233 = ~n23221 & n23231;
  assign n23234 = ~n23232 & ~n23233;
  assign n23235 = ~n23085 & n23096;
  assign n23236 = ~n23084 & ~n23235;
  assign n23237 = ~n23234 & ~n23236;
  assign n23238 = n23234 & n23236;
  assign n23239 = ~n23237 & ~n23238;
  assign n23240 = ~n22972 & ~n23100;
  assign n23241 = n23239 & ~n23240;
  assign n23242 = ~n23239 & n23240;
  assign n23243 = ~n23241 & ~n23242;
  assign n23244 = ~n23109 & n23243;
  assign n23245 = n23109 & ~n23243;
  assign po105  = ~n23244 & ~n23245;
  assign n23247 = ~n23232 & ~n23238;
  assign n23248 = ~n23214 & ~n23220;
  assign n23249 = pi126  & n6331;
  assign n23250 = pi127  & n6015;
  assign n23251 = n6008 & n12542;
  assign n23252 = ~n23249 & ~n23250;
  assign n23253 = ~n23251 & n23252;
  assign n23254 = pi44  & n23253;
  assign n23255 = ~pi44  & ~n23253;
  assign n23256 = ~n23254 & ~n23255;
  assign n23257 = ~n23248 & ~n23256;
  assign n23258 = n23248 & n23256;
  assign n23259 = ~n23257 & ~n23258;
  assign n23260 = pi123  & n7121;
  assign n23261 = pi124  & n6795;
  assign n23262 = pi125  & n6790;
  assign n23263 = n6788 & n11786;
  assign n23264 = ~n23261 & ~n23262;
  assign n23265 = ~n23260 & n23264;
  assign n23266 = ~n23263 & n23265;
  assign n23267 = pi47  & n23266;
  assign n23268 = ~pi47  & ~n23266;
  assign n23269 = ~n23267 & ~n23268;
  assign n23270 = ~n23199 & ~n23201;
  assign n23271 = pi120  & n7969;
  assign n23272 = pi121  & n7636;
  assign n23273 = pi122  & n7631;
  assign n23274 = n7629 & n10729;
  assign n23275 = ~n23272 & ~n23273;
  assign n23276 = ~n23271 & n23275;
  assign n23277 = ~n23274 & n23276;
  assign n23278 = pi50  & n23277;
  assign n23279 = ~pi50  & ~n23277;
  assign n23280 = ~n23278 & ~n23279;
  assign n23281 = ~n23193 & ~n23195;
  assign n23282 = ~n23186 & ~n23189;
  assign n23283 = ~n23180 & ~n23183;
  assign n23284 = ~n23164 & ~n23168;
  assign n23285 = pi108  & n11910;
  assign n23286 = pi109  & n11529;
  assign n23287 = pi110  & n11524;
  assign n23288 = n6995 & n11522;
  assign n23289 = ~n23286 & ~n23287;
  assign n23290 = ~n23285 & n23289;
  assign n23291 = ~n23288 & n23290;
  assign n23292 = pi62  & n23291;
  assign n23293 = ~pi62  & ~n23291;
  assign n23294 = ~n23292 & ~n23293;
  assign n23295 = ~n23145 & ~n23152;
  assign n23296 = pi107  & n12277;
  assign n23297 = pi106  & n12276;
  assign n23298 = ~n23296 & ~n23297;
  assign n23299 = ~n23295 & n23298;
  assign n23300 = n23295 & ~n23298;
  assign n23301 = ~n23299 & ~n23300;
  assign n23302 = ~n23294 & n23301;
  assign n23303 = n23294 & ~n23301;
  assign n23304 = ~n23302 & ~n23303;
  assign n23305 = ~n23284 & n23304;
  assign n23306 = n23284 & ~n23304;
  assign n23307 = ~n23305 & ~n23306;
  assign n23308 = pi111  & n10886;
  assign n23309 = pi112  & n10495;
  assign n23310 = pi113  & n10490;
  assign n23311 = n7852 & n10488;
  assign n23312 = ~n23309 & ~n23310;
  assign n23313 = ~n23308 & n23312;
  assign n23314 = ~n23311 & n23313;
  assign n23315 = pi59  & n23314;
  assign n23316 = ~pi59  & ~n23314;
  assign n23317 = ~n23315 & ~n23316;
  assign n23318 = n23307 & ~n23317;
  assign n23319 = ~n23307 & n23317;
  assign n23320 = ~n23318 & ~n23319;
  assign n23321 = n23283 & ~n23320;
  assign n23322 = ~n23283 & n23320;
  assign n23323 = ~n23321 & ~n23322;
  assign n23324 = pi114  & n9858;
  assign n23325 = pi115  & n9508;
  assign n23326 = pi116  & n9503;
  assign n23327 = n8470 & n9501;
  assign n23328 = ~n23325 & ~n23326;
  assign n23329 = ~n23324 & n23328;
  assign n23330 = ~n23327 & n23329;
  assign n23331 = pi56  & n23330;
  assign n23332 = ~pi56  & ~n23330;
  assign n23333 = ~n23331 & ~n23332;
  assign n23334 = n23323 & ~n23333;
  assign n23335 = ~n23323 & n23333;
  assign n23336 = ~n23334 & ~n23335;
  assign n23337 = n23282 & ~n23336;
  assign n23338 = ~n23282 & n23336;
  assign n23339 = ~n23337 & ~n23338;
  assign n23340 = pi117  & n8905;
  assign n23341 = pi118  & n8535;
  assign n23342 = pi119  & n8530;
  assign n23343 = n8528 & n9412;
  assign n23344 = ~n23341 & ~n23342;
  assign n23345 = ~n23340 & n23344;
  assign n23346 = ~n23343 & n23345;
  assign n23347 = pi53  & n23346;
  assign n23348 = ~pi53  & ~n23346;
  assign n23349 = ~n23347 & ~n23348;
  assign n23350 = n23339 & ~n23349;
  assign n23351 = ~n23339 & n23349;
  assign n23352 = ~n23350 & ~n23351;
  assign n23353 = ~n23281 & n23352;
  assign n23354 = n23281 & ~n23352;
  assign n23355 = ~n23353 & ~n23354;
  assign n23356 = n23280 & ~n23355;
  assign n23357 = ~n23280 & n23355;
  assign n23358 = ~n23356 & ~n23357;
  assign n23359 = ~n23270 & n23358;
  assign n23360 = n23270 & ~n23358;
  assign n23361 = ~n23359 & ~n23360;
  assign n23362 = n23269 & ~n23361;
  assign n23363 = ~n23269 & n23361;
  assign n23364 = ~n23362 & ~n23363;
  assign n23365 = n23259 & n23364;
  assign n23366 = ~n23259 & ~n23364;
  assign n23367 = ~n23365 & ~n23366;
  assign n23368 = n23247 & ~n23367;
  assign n23369 = ~n23247 & n23367;
  assign n23370 = ~n23368 & ~n23369;
  assign n23371 = ~n23241 & ~n23244;
  assign n23372 = n23370 & ~n23371;
  assign n23373 = ~n23370 & n23371;
  assign po106  = ~n23372 & ~n23373;
  assign n23375 = ~n23369 & ~n23372;
  assign n23376 = n6008 & ~n12539;
  assign n23377 = ~n6331 & ~n23376;
  assign n23378 = pi127  & ~n23377;
  assign n23379 = pi44  & ~n23378;
  assign n23380 = ~pi44  & n23378;
  assign n23381 = ~n23379 & ~n23380;
  assign n23382 = n23269 & ~n23359;
  assign n23383 = ~n23360 & ~n23382;
  assign n23384 = ~n23381 & n23383;
  assign n23385 = n23381 & ~n23383;
  assign n23386 = ~n23384 & ~n23385;
  assign n23387 = pi124  & n7121;
  assign n23388 = pi125  & n6795;
  assign n23389 = pi126  & n6790;
  assign n23390 = n6788 & n12148;
  assign n23391 = ~n23388 & ~n23389;
  assign n23392 = ~n23387 & n23391;
  assign n23393 = ~n23390 & n23392;
  assign n23394 = pi47  & n23393;
  assign n23395 = ~pi47  & ~n23393;
  assign n23396 = ~n23394 & ~n23395;
  assign n23397 = ~n23353 & ~n23357;
  assign n23398 = pi118  & n8905;
  assign n23399 = pi119  & n8535;
  assign n23400 = pi120  & n8530;
  assign n23401 = n8528 & n10047;
  assign n23402 = ~n23399 & ~n23400;
  assign n23403 = ~n23398 & n23402;
  assign n23404 = ~n23401 & n23403;
  assign n23405 = pi53  & n23404;
  assign n23406 = ~pi53  & ~n23404;
  assign n23407 = ~n23405 & ~n23406;
  assign n23408 = pi115  & n9858;
  assign n23409 = pi116  & n9508;
  assign n23410 = pi117  & n9503;
  assign n23411 = n8784 & n9501;
  assign n23412 = ~n23409 & ~n23410;
  assign n23413 = ~n23408 & n23412;
  assign n23414 = ~n23411 & n23413;
  assign n23415 = pi56  & n23414;
  assign n23416 = ~pi56  & ~n23414;
  assign n23417 = ~n23415 & ~n23416;
  assign n23418 = pi112  & n10886;
  assign n23419 = pi113  & n10495;
  assign n23420 = pi114  & n10490;
  assign n23421 = n8146 & n10488;
  assign n23422 = ~n23419 & ~n23420;
  assign n23423 = ~n23418 & n23422;
  assign n23424 = ~n23421 & n23423;
  assign n23425 = pi59  & n23424;
  assign n23426 = ~pi59  & ~n23424;
  assign n23427 = ~n23425 & ~n23426;
  assign n23428 = ~n23299 & ~n23302;
  assign n23429 = pi108  & n12277;
  assign n23430 = pi107  & n12276;
  assign n23431 = ~n23429 & ~n23430;
  assign n23432 = n23298 & ~n23431;
  assign n23433 = ~n23298 & n23431;
  assign n23434 = ~n23432 & ~n23433;
  assign n23435 = pi109  & n11910;
  assign n23436 = pi110  & n11529;
  assign n23437 = pi111  & n11524;
  assign n23438 = n7272 & n11522;
  assign n23439 = ~n23436 & ~n23437;
  assign n23440 = ~n23435 & n23439;
  assign n23441 = ~n23438 & n23440;
  assign n23442 = pi62  & n23441;
  assign n23443 = ~pi62  & ~n23441;
  assign n23444 = ~n23442 & ~n23443;
  assign n23445 = n23434 & ~n23444;
  assign n23446 = ~n23434 & n23444;
  assign n23447 = ~n23445 & ~n23446;
  assign n23448 = ~n23428 & n23447;
  assign n23449 = n23428 & ~n23447;
  assign n23450 = ~n23448 & ~n23449;
  assign n23451 = ~n23427 & n23450;
  assign n23452 = n23427 & ~n23450;
  assign n23453 = ~n23451 & ~n23452;
  assign n23454 = ~n23305 & n23317;
  assign n23455 = ~n23306 & ~n23454;
  assign n23456 = n23453 & n23455;
  assign n23457 = ~n23453 & ~n23455;
  assign n23458 = ~n23456 & ~n23457;
  assign n23459 = ~n23417 & n23458;
  assign n23460 = n23417 & ~n23458;
  assign n23461 = ~n23459 & ~n23460;
  assign n23462 = ~n23322 & n23333;
  assign n23463 = ~n23321 & ~n23462;
  assign n23464 = n23461 & n23463;
  assign n23465 = ~n23461 & ~n23463;
  assign n23466 = ~n23464 & ~n23465;
  assign n23467 = ~n23407 & n23466;
  assign n23468 = n23407 & ~n23466;
  assign n23469 = ~n23467 & ~n23468;
  assign n23470 = ~n23338 & n23349;
  assign n23471 = ~n23337 & ~n23470;
  assign n23472 = n23469 & n23471;
  assign n23473 = ~n23469 & ~n23471;
  assign n23474 = ~n23472 & ~n23473;
  assign n23475 = pi121  & n7969;
  assign n23476 = pi122  & n7636;
  assign n23477 = pi123  & n7631;
  assign n23478 = n7629 & n10754;
  assign n23479 = ~n23476 & ~n23477;
  assign n23480 = ~n23475 & n23479;
  assign n23481 = ~n23478 & n23480;
  assign n23482 = pi50  & n23481;
  assign n23483 = ~pi50  & ~n23481;
  assign n23484 = ~n23482 & ~n23483;
  assign n23485 = n23474 & ~n23484;
  assign n23486 = ~n23474 & n23484;
  assign n23487 = ~n23485 & ~n23486;
  assign n23488 = ~n23397 & n23487;
  assign n23489 = n23397 & ~n23487;
  assign n23490 = ~n23488 & ~n23489;
  assign n23491 = n23396 & ~n23490;
  assign n23492 = ~n23396 & n23490;
  assign n23493 = ~n23491 & ~n23492;
  assign n23494 = n23386 & n23493;
  assign n23495 = ~n23386 & ~n23493;
  assign n23496 = ~n23494 & ~n23495;
  assign n23497 = ~n23257 & ~n23364;
  assign n23498 = ~n23258 & ~n23497;
  assign n23499 = n23496 & n23498;
  assign n23500 = ~n23496 & ~n23498;
  assign n23501 = ~n23499 & ~n23500;
  assign n23502 = ~n23375 & n23501;
  assign n23503 = n23375 & ~n23501;
  assign po107  = ~n23502 & ~n23503;
  assign n23505 = ~n23499 & ~n23502;
  assign n23506 = pi122  & n7969;
  assign n23507 = pi123  & n7636;
  assign n23508 = pi124  & n7631;
  assign n23509 = n7629 & n11099;
  assign n23510 = ~n23507 & ~n23508;
  assign n23511 = ~n23506 & n23510;
  assign n23512 = ~n23509 & n23511;
  assign n23513 = pi50  & n23512;
  assign n23514 = ~pi50  & ~n23512;
  assign n23515 = ~n23513 & ~n23514;
  assign n23516 = ~n23464 & ~n23467;
  assign n23517 = pi119  & n8905;
  assign n23518 = pi120  & n8535;
  assign n23519 = pi121  & n8530;
  assign n23520 = n8528 & n10071;
  assign n23521 = ~n23518 & ~n23519;
  assign n23522 = ~n23517 & n23521;
  assign n23523 = ~n23520 & n23522;
  assign n23524 = pi53  & n23523;
  assign n23525 = ~pi53  & ~n23523;
  assign n23526 = ~n23524 & ~n23525;
  assign n23527 = ~n23456 & ~n23459;
  assign n23528 = pi116  & n9858;
  assign n23529 = pi117  & n9508;
  assign n23530 = pi118  & n9503;
  assign n23531 = n9095 & n9501;
  assign n23532 = ~n23529 & ~n23530;
  assign n23533 = ~n23528 & n23532;
  assign n23534 = ~n23531 & n23533;
  assign n23535 = pi56  & n23534;
  assign n23536 = ~pi56  & ~n23534;
  assign n23537 = ~n23535 & ~n23536;
  assign n23538 = ~n23448 & ~n23451;
  assign n23539 = pi113  & n10886;
  assign n23540 = pi114  & n10495;
  assign n23541 = pi115  & n10490;
  assign n23542 = n8170 & n10488;
  assign n23543 = ~n23540 & ~n23541;
  assign n23544 = ~n23539 & n23543;
  assign n23545 = ~n23542 & n23544;
  assign n23546 = pi59  & n23545;
  assign n23547 = ~pi59  & ~n23545;
  assign n23548 = ~n23546 & ~n23547;
  assign n23549 = pi110  & n11910;
  assign n23550 = pi111  & n11529;
  assign n23551 = pi112  & n11524;
  assign n23552 = n7296 & n11522;
  assign n23553 = ~n23550 & ~n23551;
  assign n23554 = ~n23549 & n23553;
  assign n23555 = ~n23552 & n23554;
  assign n23556 = pi62  & n23555;
  assign n23557 = ~pi62  & ~n23555;
  assign n23558 = ~n23556 & ~n23557;
  assign n23559 = ~n23432 & ~n23445;
  assign n23560 = pi109  & n12277;
  assign n23561 = pi108  & n12276;
  assign n23562 = ~n23560 & ~n23561;
  assign n23563 = ~pi44  & ~n23562;
  assign n23564 = pi44  & n23562;
  assign n23565 = ~n23563 & ~n23564;
  assign n23566 = ~n23298 & n23565;
  assign n23567 = n23298 & ~n23565;
  assign n23568 = ~n23566 & ~n23567;
  assign n23569 = ~n23559 & n23568;
  assign n23570 = n23559 & ~n23568;
  assign n23571 = ~n23569 & ~n23570;
  assign n23572 = ~n23558 & n23571;
  assign n23573 = n23558 & ~n23571;
  assign n23574 = ~n23572 & ~n23573;
  assign n23575 = n23548 & ~n23574;
  assign n23576 = ~n23548 & n23574;
  assign n23577 = ~n23575 & ~n23576;
  assign n23578 = ~n23538 & n23577;
  assign n23579 = n23538 & ~n23577;
  assign n23580 = ~n23578 & ~n23579;
  assign n23581 = n23537 & ~n23580;
  assign n23582 = ~n23537 & n23580;
  assign n23583 = ~n23581 & ~n23582;
  assign n23584 = ~n23527 & n23583;
  assign n23585 = n23527 & ~n23583;
  assign n23586 = ~n23584 & ~n23585;
  assign n23587 = n23526 & ~n23586;
  assign n23588 = ~n23526 & n23586;
  assign n23589 = ~n23587 & ~n23588;
  assign n23590 = ~n23516 & n23589;
  assign n23591 = n23516 & ~n23589;
  assign n23592 = ~n23590 & ~n23591;
  assign n23593 = n23515 & ~n23592;
  assign n23594 = ~n23515 & n23592;
  assign n23595 = ~n23593 & ~n23594;
  assign n23596 = ~n23472 & n23484;
  assign n23597 = ~n23473 & ~n23596;
  assign n23598 = n23595 & n23597;
  assign n23599 = ~n23595 & ~n23597;
  assign n23600 = ~n23598 & ~n23599;
  assign n23601 = pi125  & n7121;
  assign n23602 = pi126  & n6795;
  assign n23603 = pi127  & n6790;
  assign n23604 = n6788 & n12519;
  assign n23605 = ~n23602 & ~n23603;
  assign n23606 = ~n23601 & n23605;
  assign n23607 = ~n23604 & n23606;
  assign n23608 = pi47  & n23607;
  assign n23609 = ~pi47  & ~n23607;
  assign n23610 = ~n23608 & ~n23609;
  assign n23611 = n23600 & ~n23610;
  assign n23612 = ~n23600 & n23610;
  assign n23613 = ~n23611 & ~n23612;
  assign n23614 = n23396 & ~n23488;
  assign n23615 = ~n23489 & ~n23614;
  assign n23616 = ~n23613 & ~n23615;
  assign n23617 = n23613 & n23615;
  assign n23618 = ~n23616 & ~n23617;
  assign n23619 = ~n23384 & ~n23494;
  assign n23620 = n23618 & ~n23619;
  assign n23621 = ~n23618 & n23619;
  assign n23622 = ~n23620 & ~n23621;
  assign n23623 = ~n23505 & n23622;
  assign n23624 = n23505 & ~n23622;
  assign po108  = ~n23623 & ~n23624;
  assign n23626 = ~n23611 & ~n23617;
  assign n23627 = ~n23594 & ~n23598;
  assign n23628 = pi126  & n7121;
  assign n23629 = pi127  & n6795;
  assign n23630 = n6788 & n12542;
  assign n23631 = ~n23628 & ~n23629;
  assign n23632 = ~n23630 & n23631;
  assign n23633 = pi47  & n23632;
  assign n23634 = ~pi47  & ~n23632;
  assign n23635 = ~n23633 & ~n23634;
  assign n23636 = ~n23627 & ~n23635;
  assign n23637 = n23627 & n23635;
  assign n23638 = ~n23636 & ~n23637;
  assign n23639 = pi123  & n7969;
  assign n23640 = pi124  & n7636;
  assign n23641 = pi125  & n7631;
  assign n23642 = n7629 & n11786;
  assign n23643 = ~n23640 & ~n23641;
  assign n23644 = ~n23639 & n23643;
  assign n23645 = ~n23642 & n23644;
  assign n23646 = pi50  & n23645;
  assign n23647 = ~pi50  & ~n23645;
  assign n23648 = ~n23646 & ~n23647;
  assign n23649 = ~n23588 & ~n23590;
  assign n23650 = pi120  & n8905;
  assign n23651 = pi121  & n8535;
  assign n23652 = pi122  & n8530;
  assign n23653 = n8528 & n10729;
  assign n23654 = ~n23651 & ~n23652;
  assign n23655 = ~n23650 & n23654;
  assign n23656 = ~n23653 & n23655;
  assign n23657 = pi53  & n23656;
  assign n23658 = ~pi53  & ~n23656;
  assign n23659 = ~n23657 & ~n23658;
  assign n23660 = ~n23582 & ~n23584;
  assign n23661 = ~n23576 & ~n23578;
  assign n23662 = pi114  & n10886;
  assign n23663 = pi115  & n10495;
  assign n23664 = pi116  & n10490;
  assign n23665 = n8470 & n10488;
  assign n23666 = ~n23663 & ~n23664;
  assign n23667 = ~n23662 & n23666;
  assign n23668 = ~n23665 & n23667;
  assign n23669 = pi59  & n23668;
  assign n23670 = ~pi59  & ~n23668;
  assign n23671 = ~n23669 & ~n23670;
  assign n23672 = ~n23569 & ~n23572;
  assign n23673 = ~n23298 & ~n23564;
  assign n23674 = ~n23563 & ~n23673;
  assign n23675 = pi110  & n12277;
  assign n23676 = pi109  & n12276;
  assign n23677 = ~n23675 & ~n23676;
  assign n23678 = n23674 & ~n23677;
  assign n23679 = ~n23674 & n23677;
  assign n23680 = ~n23678 & ~n23679;
  assign n23681 = pi111  & n11910;
  assign n23682 = pi112  & n11529;
  assign n23683 = pi113  & n11524;
  assign n23684 = n7852 & n11522;
  assign n23685 = ~n23682 & ~n23683;
  assign n23686 = ~n23681 & n23685;
  assign n23687 = ~n23684 & n23686;
  assign n23688 = pi62  & n23687;
  assign n23689 = ~pi62  & ~n23687;
  assign n23690 = ~n23688 & ~n23689;
  assign n23691 = ~n23680 & n23690;
  assign n23692 = n23680 & ~n23690;
  assign n23693 = ~n23691 & ~n23692;
  assign n23694 = ~n23672 & n23693;
  assign n23695 = n23672 & ~n23693;
  assign n23696 = ~n23694 & ~n23695;
  assign n23697 = ~n23671 & n23696;
  assign n23698 = n23671 & ~n23696;
  assign n23699 = ~n23697 & ~n23698;
  assign n23700 = ~n23661 & n23699;
  assign n23701 = n23661 & ~n23699;
  assign n23702 = ~n23700 & ~n23701;
  assign n23703 = pi117  & n9858;
  assign n23704 = pi118  & n9508;
  assign n23705 = pi119  & n9503;
  assign n23706 = n9412 & n9501;
  assign n23707 = ~n23704 & ~n23705;
  assign n23708 = ~n23703 & n23707;
  assign n23709 = ~n23706 & n23708;
  assign n23710 = pi56  & n23709;
  assign n23711 = ~pi56  & ~n23709;
  assign n23712 = ~n23710 & ~n23711;
  assign n23713 = n23702 & ~n23712;
  assign n23714 = ~n23702 & n23712;
  assign n23715 = ~n23713 & ~n23714;
  assign n23716 = ~n23660 & n23715;
  assign n23717 = n23660 & ~n23715;
  assign n23718 = ~n23716 & ~n23717;
  assign n23719 = n23659 & ~n23718;
  assign n23720 = ~n23659 & n23718;
  assign n23721 = ~n23719 & ~n23720;
  assign n23722 = ~n23649 & n23721;
  assign n23723 = n23649 & ~n23721;
  assign n23724 = ~n23722 & ~n23723;
  assign n23725 = n23648 & ~n23724;
  assign n23726 = ~n23648 & n23724;
  assign n23727 = ~n23725 & ~n23726;
  assign n23728 = n23638 & n23727;
  assign n23729 = ~n23638 & ~n23727;
  assign n23730 = ~n23728 & ~n23729;
  assign n23731 = n23626 & ~n23730;
  assign n23732 = ~n23626 & n23730;
  assign n23733 = ~n23731 & ~n23732;
  assign n23734 = ~n23620 & ~n23623;
  assign n23735 = n23733 & ~n23734;
  assign n23736 = ~n23733 & n23734;
  assign po109  = ~n23735 & ~n23736;
  assign n23738 = n6788 & ~n12539;
  assign n23739 = ~n7121 & ~n23738;
  assign n23740 = pi127  & ~n23739;
  assign n23741 = pi47  & ~n23740;
  assign n23742 = ~pi47  & n23740;
  assign n23743 = ~n23741 & ~n23742;
  assign n23744 = n23648 & ~n23722;
  assign n23745 = ~n23723 & ~n23744;
  assign n23746 = ~n23743 & n23745;
  assign n23747 = n23743 & ~n23745;
  assign n23748 = ~n23746 & ~n23747;
  assign n23749 = pi124  & n7969;
  assign n23750 = pi125  & n7636;
  assign n23751 = pi126  & n7631;
  assign n23752 = n7629 & n12148;
  assign n23753 = ~n23750 & ~n23751;
  assign n23754 = ~n23749 & n23753;
  assign n23755 = ~n23752 & n23754;
  assign n23756 = pi50  & n23755;
  assign n23757 = ~pi50  & ~n23755;
  assign n23758 = ~n23756 & ~n23757;
  assign n23759 = ~n23716 & ~n23720;
  assign n23760 = pi118  & n9858;
  assign n23761 = pi119  & n9508;
  assign n23762 = pi120  & n9503;
  assign n23763 = n9501 & n10047;
  assign n23764 = ~n23761 & ~n23762;
  assign n23765 = ~n23760 & n23764;
  assign n23766 = ~n23763 & n23765;
  assign n23767 = pi56  & n23766;
  assign n23768 = ~pi56  & ~n23766;
  assign n23769 = ~n23767 & ~n23768;
  assign n23770 = ~n23694 & ~n23697;
  assign n23771 = pi115  & n10886;
  assign n23772 = pi116  & n10495;
  assign n23773 = pi117  & n10490;
  assign n23774 = n8784 & n10488;
  assign n23775 = ~n23772 & ~n23773;
  assign n23776 = ~n23771 & n23775;
  assign n23777 = ~n23774 & n23776;
  assign n23778 = pi59  & n23777;
  assign n23779 = ~pi59  & ~n23777;
  assign n23780 = ~n23778 & ~n23779;
  assign n23781 = pi112  & n11910;
  assign n23782 = pi113  & n11529;
  assign n23783 = pi114  & n11524;
  assign n23784 = n8146 & n11522;
  assign n23785 = ~n23782 & ~n23783;
  assign n23786 = ~n23781 & n23785;
  assign n23787 = ~n23784 & n23786;
  assign n23788 = pi62  & n23787;
  assign n23789 = ~pi62  & ~n23787;
  assign n23790 = ~n23788 & ~n23789;
  assign n23791 = ~n23679 & ~n23692;
  assign n23792 = pi111  & n12277;
  assign n23793 = pi110  & n12276;
  assign n23794 = ~n23792 & ~n23793;
  assign n23795 = n23677 & ~n23794;
  assign n23796 = ~n23677 & n23794;
  assign n23797 = ~n23795 & ~n23796;
  assign n23798 = ~n23791 & n23797;
  assign n23799 = n23791 & ~n23797;
  assign n23800 = ~n23798 & ~n23799;
  assign n23801 = ~n23790 & n23800;
  assign n23802 = n23790 & ~n23800;
  assign n23803 = ~n23801 & ~n23802;
  assign n23804 = ~n23780 & n23803;
  assign n23805 = n23780 & ~n23803;
  assign n23806 = ~n23804 & ~n23805;
  assign n23807 = ~n23770 & n23806;
  assign n23808 = n23770 & ~n23806;
  assign n23809 = ~n23807 & ~n23808;
  assign n23810 = ~n23769 & n23809;
  assign n23811 = n23769 & ~n23809;
  assign n23812 = ~n23810 & ~n23811;
  assign n23813 = ~n23700 & n23712;
  assign n23814 = ~n23701 & ~n23813;
  assign n23815 = n23812 & n23814;
  assign n23816 = ~n23812 & ~n23814;
  assign n23817 = ~n23815 & ~n23816;
  assign n23818 = pi121  & n8905;
  assign n23819 = pi122  & n8535;
  assign n23820 = pi123  & n8530;
  assign n23821 = n8528 & n10754;
  assign n23822 = ~n23819 & ~n23820;
  assign n23823 = ~n23818 & n23822;
  assign n23824 = ~n23821 & n23823;
  assign n23825 = pi53  & n23824;
  assign n23826 = ~pi53  & ~n23824;
  assign n23827 = ~n23825 & ~n23826;
  assign n23828 = n23817 & ~n23827;
  assign n23829 = ~n23817 & n23827;
  assign n23830 = ~n23828 & ~n23829;
  assign n23831 = ~n23759 & n23830;
  assign n23832 = n23759 & ~n23830;
  assign n23833 = ~n23831 & ~n23832;
  assign n23834 = n23758 & ~n23833;
  assign n23835 = ~n23758 & n23833;
  assign n23836 = ~n23834 & ~n23835;
  assign n23837 = n23748 & n23836;
  assign n23838 = ~n23748 & ~n23836;
  assign n23839 = ~n23837 & ~n23838;
  assign n23840 = ~n23636 & ~n23727;
  assign n23841 = ~n23637 & ~n23840;
  assign n23842 = ~n23839 & ~n23841;
  assign n23843 = n23839 & n23841;
  assign n23844 = ~n23842 & ~n23843;
  assign n23845 = ~n23732 & ~n23735;
  assign n23846 = n23844 & ~n23845;
  assign n23847 = ~n23844 & n23845;
  assign po110  = ~n23846 & ~n23847;
  assign n23849 = pi122  & n8905;
  assign n23850 = pi123  & n8535;
  assign n23851 = pi124  & n8530;
  assign n23852 = n8528 & n11099;
  assign n23853 = ~n23850 & ~n23851;
  assign n23854 = ~n23849 & n23853;
  assign n23855 = ~n23852 & n23854;
  assign n23856 = pi53  & n23855;
  assign n23857 = ~pi53  & ~n23855;
  assign n23858 = ~n23856 & ~n23857;
  assign n23859 = ~n23807 & ~n23810;
  assign n23860 = pi119  & n9858;
  assign n23861 = pi120  & n9508;
  assign n23862 = pi121  & n9503;
  assign n23863 = n9501 & n10071;
  assign n23864 = ~n23861 & ~n23862;
  assign n23865 = ~n23860 & n23864;
  assign n23866 = ~n23863 & n23865;
  assign n23867 = pi56  & n23866;
  assign n23868 = ~pi56  & ~n23866;
  assign n23869 = ~n23867 & ~n23868;
  assign n23870 = ~n23801 & ~n23804;
  assign n23871 = pi116  & n10886;
  assign n23872 = pi117  & n10495;
  assign n23873 = pi118  & n10490;
  assign n23874 = n9095 & n10488;
  assign n23875 = ~n23872 & ~n23873;
  assign n23876 = ~n23871 & n23875;
  assign n23877 = ~n23874 & n23876;
  assign n23878 = pi59  & n23877;
  assign n23879 = ~pi59  & ~n23877;
  assign n23880 = ~n23878 & ~n23879;
  assign n23881 = ~n23796 & ~n23798;
  assign n23882 = pi113  & n11910;
  assign n23883 = pi114  & n11529;
  assign n23884 = pi115  & n11524;
  assign n23885 = n8170 & n11522;
  assign n23886 = ~n23883 & ~n23884;
  assign n23887 = ~n23882 & n23886;
  assign n23888 = ~n23885 & n23887;
  assign n23889 = pi62  & n23888;
  assign n23890 = ~pi62  & ~n23888;
  assign n23891 = ~n23889 & ~n23890;
  assign n23892 = ~pi47  & ~n23794;
  assign n23893 = pi47  & n23794;
  assign n23894 = ~n23892 & ~n23893;
  assign n23895 = pi112  & n12277;
  assign n23896 = pi111  & n12276;
  assign n23897 = ~n23895 & ~n23896;
  assign n23898 = n23894 & ~n23897;
  assign n23899 = ~n23894 & n23897;
  assign n23900 = ~n23898 & ~n23899;
  assign n23901 = ~n23891 & n23900;
  assign n23902 = n23891 & ~n23900;
  assign n23903 = ~n23901 & ~n23902;
  assign n23904 = ~n23881 & n23903;
  assign n23905 = n23881 & ~n23903;
  assign n23906 = ~n23904 & ~n23905;
  assign n23907 = n23880 & ~n23906;
  assign n23908 = ~n23880 & n23906;
  assign n23909 = ~n23907 & ~n23908;
  assign n23910 = ~n23870 & n23909;
  assign n23911 = n23870 & ~n23909;
  assign n23912 = ~n23910 & ~n23911;
  assign n23913 = n23869 & ~n23912;
  assign n23914 = ~n23869 & n23912;
  assign n23915 = ~n23913 & ~n23914;
  assign n23916 = ~n23859 & n23915;
  assign n23917 = n23859 & ~n23915;
  assign n23918 = ~n23916 & ~n23917;
  assign n23919 = n23858 & ~n23918;
  assign n23920 = ~n23858 & n23918;
  assign n23921 = ~n23919 & ~n23920;
  assign n23922 = ~n23815 & n23827;
  assign n23923 = ~n23816 & ~n23922;
  assign n23924 = n23921 & n23923;
  assign n23925 = ~n23921 & ~n23923;
  assign n23926 = ~n23924 & ~n23925;
  assign n23927 = pi125  & n7969;
  assign n23928 = pi126  & n7636;
  assign n23929 = pi127  & n7631;
  assign n23930 = n7629 & n12519;
  assign n23931 = ~n23928 & ~n23929;
  assign n23932 = ~n23927 & n23931;
  assign n23933 = ~n23930 & n23932;
  assign n23934 = pi50  & n23933;
  assign n23935 = ~pi50  & ~n23933;
  assign n23936 = ~n23934 & ~n23935;
  assign n23937 = n23926 & ~n23936;
  assign n23938 = ~n23926 & n23936;
  assign n23939 = ~n23937 & ~n23938;
  assign n23940 = n23758 & ~n23831;
  assign n23941 = ~n23832 & ~n23940;
  assign n23942 = ~n23939 & ~n23941;
  assign n23943 = n23939 & n23941;
  assign n23944 = ~n23942 & ~n23943;
  assign n23945 = ~n23746 & ~n23836;
  assign n23946 = ~n23747 & ~n23945;
  assign n23947 = ~n23944 & ~n23946;
  assign n23948 = n23944 & n23946;
  assign n23949 = ~n23947 & ~n23948;
  assign n23950 = ~n23843 & ~n23846;
  assign n23951 = n23949 & ~n23950;
  assign n23952 = ~n23949 & n23950;
  assign po111  = ~n23951 & ~n23952;
  assign n23954 = ~n23937 & ~n23943;
  assign n23955 = ~n23920 & ~n23924;
  assign n23956 = pi123  & n8905;
  assign n23957 = pi124  & n8535;
  assign n23958 = pi125  & n8530;
  assign n23959 = n8528 & n11786;
  assign n23960 = ~n23957 & ~n23958;
  assign n23961 = ~n23956 & n23960;
  assign n23962 = ~n23959 & n23961;
  assign n23963 = pi53  & n23962;
  assign n23964 = ~pi53  & ~n23962;
  assign n23965 = ~n23963 & ~n23964;
  assign n23966 = ~n23914 & ~n23916;
  assign n23967 = pi120  & n9858;
  assign n23968 = pi121  & n9508;
  assign n23969 = pi122  & n9503;
  assign n23970 = n9501 & n10729;
  assign n23971 = ~n23968 & ~n23969;
  assign n23972 = ~n23967 & n23971;
  assign n23973 = ~n23970 & n23972;
  assign n23974 = pi56  & n23973;
  assign n23975 = ~pi56  & ~n23973;
  assign n23976 = ~n23974 & ~n23975;
  assign n23977 = ~n23908 & ~n23910;
  assign n23978 = pi117  & n10886;
  assign n23979 = pi118  & n10495;
  assign n23980 = pi119  & n10490;
  assign n23981 = n9412 & n10488;
  assign n23982 = ~n23979 & ~n23980;
  assign n23983 = ~n23978 & n23982;
  assign n23984 = ~n23981 & n23983;
  assign n23985 = pi59  & n23984;
  assign n23986 = ~pi59  & ~n23984;
  assign n23987 = ~n23985 & ~n23986;
  assign n23988 = ~n23901 & ~n23904;
  assign n23989 = ~n23892 & ~n23898;
  assign n23990 = pi113  & n12277;
  assign n23991 = pi112  & n12276;
  assign n23992 = ~n23990 & ~n23991;
  assign n23993 = ~n23989 & n23992;
  assign n23994 = n23989 & ~n23992;
  assign n23995 = ~n23993 & ~n23994;
  assign n23996 = pi114  & n11910;
  assign n23997 = pi115  & n11529;
  assign n23998 = pi116  & n11524;
  assign n23999 = n8470 & n11522;
  assign n24000 = ~n23997 & ~n23998;
  assign n24001 = ~n23996 & n24000;
  assign n24002 = ~n23999 & n24001;
  assign n24003 = pi62  & n24002;
  assign n24004 = ~pi62  & ~n24002;
  assign n24005 = ~n24003 & ~n24004;
  assign n24006 = n23995 & ~n24005;
  assign n24007 = ~n23995 & n24005;
  assign n24008 = ~n24006 & ~n24007;
  assign n24009 = ~n23988 & n24008;
  assign n24010 = n23988 & ~n24008;
  assign n24011 = ~n24009 & ~n24010;
  assign n24012 = ~n23987 & n24011;
  assign n24013 = n23987 & ~n24011;
  assign n24014 = ~n24012 & ~n24013;
  assign n24015 = ~n23977 & n24014;
  assign n24016 = n23977 & ~n24014;
  assign n24017 = ~n24015 & ~n24016;
  assign n24018 = ~n23976 & n24017;
  assign n24019 = n23976 & ~n24017;
  assign n24020 = ~n24018 & ~n24019;
  assign n24021 = ~n23966 & n24020;
  assign n24022 = n23966 & ~n24020;
  assign n24023 = ~n24021 & ~n24022;
  assign n24024 = ~n23965 & n24023;
  assign n24025 = n23965 & ~n24023;
  assign n24026 = ~n24024 & ~n24025;
  assign n24027 = ~n23955 & n24026;
  assign n24028 = n23955 & ~n24026;
  assign n24029 = ~n24027 & ~n24028;
  assign n24030 = pi126  & n7969;
  assign n24031 = pi127  & n7636;
  assign n24032 = n7629 & n12542;
  assign n24033 = ~n24030 & ~n24031;
  assign n24034 = ~n24032 & n24033;
  assign n24035 = pi50  & n24034;
  assign n24036 = ~pi50  & ~n24034;
  assign n24037 = ~n24035 & ~n24036;
  assign n24038 = n24029 & ~n24037;
  assign n24039 = ~n24029 & n24037;
  assign n24040 = ~n24038 & ~n24039;
  assign n24041 = n23954 & ~n24040;
  assign n24042 = ~n23954 & n24040;
  assign n24043 = ~n24041 & ~n24042;
  assign n24044 = ~n23948 & ~n23951;
  assign n24045 = n24043 & ~n24044;
  assign n24046 = ~n24043 & n24044;
  assign po112  = ~n24045 & ~n24046;
  assign n24048 = ~n24021 & ~n24024;
  assign n24049 = n7629 & ~n12539;
  assign n24050 = ~n7969 & ~n24049;
  assign n24051 = pi127  & ~n24050;
  assign n24052 = pi50  & ~n24051;
  assign n24053 = ~pi50  & n24051;
  assign n24054 = ~n24052 & ~n24053;
  assign n24055 = ~n24048 & ~n24054;
  assign n24056 = n24048 & n24054;
  assign n24057 = ~n24055 & ~n24056;
  assign n24058 = ~n24015 & ~n24018;
  assign n24059 = ~n24009 & ~n24012;
  assign n24060 = ~n23993 & ~n24006;
  assign n24061 = pi115  & n11910;
  assign n24062 = pi116  & n11529;
  assign n24063 = pi117  & n11524;
  assign n24064 = n8784 & n11522;
  assign n24065 = ~n24062 & ~n24063;
  assign n24066 = ~n24061 & n24065;
  assign n24067 = ~n24064 & n24066;
  assign n24068 = pi62  & n24067;
  assign n24069 = ~pi62  & ~n24067;
  assign n24070 = ~n24068 & ~n24069;
  assign n24071 = pi114  & n12277;
  assign n24072 = pi113  & n12276;
  assign n24073 = ~n24071 & ~n24072;
  assign n24074 = n23992 & ~n24073;
  assign n24075 = ~n23992 & n24073;
  assign n24076 = ~n24074 & ~n24075;
  assign n24077 = ~n24070 & n24076;
  assign n24078 = n24070 & ~n24076;
  assign n24079 = ~n24077 & ~n24078;
  assign n24080 = n24060 & ~n24079;
  assign n24081 = ~n24060 & n24079;
  assign n24082 = ~n24080 & ~n24081;
  assign n24083 = pi118  & n10886;
  assign n24084 = pi119  & n10495;
  assign n24085 = pi120  & n10490;
  assign n24086 = n10047 & n10488;
  assign n24087 = ~n24084 & ~n24085;
  assign n24088 = ~n24083 & n24087;
  assign n24089 = ~n24086 & n24088;
  assign n24090 = pi59  & n24089;
  assign n24091 = ~pi59  & ~n24089;
  assign n24092 = ~n24090 & ~n24091;
  assign n24093 = ~n24082 & n24092;
  assign n24094 = n24082 & ~n24092;
  assign n24095 = ~n24093 & ~n24094;
  assign n24096 = ~n24059 & n24095;
  assign n24097 = n24059 & ~n24095;
  assign n24098 = ~n24096 & ~n24097;
  assign n24099 = pi121  & n9858;
  assign n24100 = pi122  & n9508;
  assign n24101 = pi123  & n9503;
  assign n24102 = n9501 & n10754;
  assign n24103 = ~n24100 & ~n24101;
  assign n24104 = ~n24099 & n24103;
  assign n24105 = ~n24102 & n24104;
  assign n24106 = pi56  & n24105;
  assign n24107 = ~pi56  & ~n24105;
  assign n24108 = ~n24106 & ~n24107;
  assign n24109 = n24098 & ~n24108;
  assign n24110 = ~n24098 & n24108;
  assign n24111 = ~n24109 & ~n24110;
  assign n24112 = n24058 & ~n24111;
  assign n24113 = ~n24058 & n24111;
  assign n24114 = ~n24112 & ~n24113;
  assign n24115 = pi124  & n8905;
  assign n24116 = pi125  & n8535;
  assign n24117 = pi126  & n8530;
  assign n24118 = n8528 & n12148;
  assign n24119 = ~n24116 & ~n24117;
  assign n24120 = ~n24115 & n24119;
  assign n24121 = ~n24118 & n24120;
  assign n24122 = pi53  & n24121;
  assign n24123 = ~pi53  & ~n24121;
  assign n24124 = ~n24122 & ~n24123;
  assign n24125 = n24114 & ~n24124;
  assign n24126 = ~n24114 & n24124;
  assign n24127 = ~n24125 & ~n24126;
  assign n24128 = n24057 & n24127;
  assign n24129 = ~n24057 & ~n24127;
  assign n24130 = ~n24128 & ~n24129;
  assign n24131 = ~n24027 & n24037;
  assign n24132 = ~n24028 & ~n24131;
  assign n24133 = ~n24130 & ~n24132;
  assign n24134 = n24130 & n24132;
  assign n24135 = ~n24133 & ~n24134;
  assign n24136 = ~n24042 & ~n24045;
  assign n24137 = n24135 & ~n24136;
  assign n24138 = ~n24135 & n24136;
  assign po113  = ~n24137 & ~n24138;
  assign n24140 = pi122  & n9858;
  assign n24141 = pi123  & n9508;
  assign n24142 = pi124  & n9503;
  assign n24143 = n9501 & n11099;
  assign n24144 = ~n24141 & ~n24142;
  assign n24145 = ~n24140 & n24144;
  assign n24146 = ~n24143 & n24145;
  assign n24147 = pi56  & n24146;
  assign n24148 = ~pi56  & ~n24146;
  assign n24149 = ~n24147 & ~n24148;
  assign n24150 = ~n24081 & ~n24094;
  assign n24151 = pi119  & n10886;
  assign n24152 = pi120  & n10495;
  assign n24153 = pi121  & n10490;
  assign n24154 = n10071 & n10488;
  assign n24155 = ~n24152 & ~n24153;
  assign n24156 = ~n24151 & n24155;
  assign n24157 = ~n24154 & n24156;
  assign n24158 = pi59  & n24157;
  assign n24159 = ~pi59  & ~n24157;
  assign n24160 = ~n24158 & ~n24159;
  assign n24161 = pi116  & n11910;
  assign n24162 = pi117  & n11529;
  assign n24163 = pi118  & n11524;
  assign n24164 = n9095 & n11522;
  assign n24165 = ~n24162 & ~n24163;
  assign n24166 = ~n24161 & n24165;
  assign n24167 = ~n24164 & n24166;
  assign n24168 = pi62  & n24167;
  assign n24169 = ~pi62  & ~n24167;
  assign n24170 = ~n24168 & ~n24169;
  assign n24171 = ~n24074 & ~n24077;
  assign n24172 = pi115  & n12277;
  assign n24173 = pi114  & n12276;
  assign n24174 = ~n24172 & ~n24173;
  assign n24175 = ~pi50  & ~n24174;
  assign n24176 = pi50  & n24174;
  assign n24177 = ~n24175 & ~n24176;
  assign n24178 = ~n23992 & n24177;
  assign n24179 = n23992 & ~n24177;
  assign n24180 = ~n24178 & ~n24179;
  assign n24181 = ~n24171 & n24180;
  assign n24182 = n24171 & ~n24180;
  assign n24183 = ~n24181 & ~n24182;
  assign n24184 = ~n24170 & n24183;
  assign n24185 = n24170 & ~n24183;
  assign n24186 = ~n24184 & ~n24185;
  assign n24187 = ~n24160 & n24186;
  assign n24188 = n24160 & ~n24186;
  assign n24189 = ~n24187 & ~n24188;
  assign n24190 = ~n24150 & n24189;
  assign n24191 = n24150 & ~n24189;
  assign n24192 = ~n24190 & ~n24191;
  assign n24193 = ~n24149 & n24192;
  assign n24194 = n24149 & ~n24192;
  assign n24195 = ~n24193 & ~n24194;
  assign n24196 = ~n24096 & n24108;
  assign n24197 = ~n24097 & ~n24196;
  assign n24198 = n24195 & n24197;
  assign n24199 = ~n24195 & ~n24197;
  assign n24200 = ~n24198 & ~n24199;
  assign n24201 = pi125  & n8905;
  assign n24202 = pi126  & n8535;
  assign n24203 = pi127  & n8530;
  assign n24204 = n8528 & n12519;
  assign n24205 = ~n24202 & ~n24203;
  assign n24206 = ~n24201 & n24205;
  assign n24207 = ~n24204 & n24206;
  assign n24208 = pi53  & n24207;
  assign n24209 = ~pi53  & ~n24207;
  assign n24210 = ~n24208 & ~n24209;
  assign n24211 = n24200 & ~n24210;
  assign n24212 = ~n24200 & n24210;
  assign n24213 = ~n24211 & ~n24212;
  assign n24214 = ~n24113 & n24124;
  assign n24215 = ~n24112 & ~n24214;
  assign n24216 = ~n24213 & ~n24215;
  assign n24217 = n24213 & n24215;
  assign n24218 = ~n24216 & ~n24217;
  assign n24219 = ~n24055 & ~n24127;
  assign n24220 = ~n24056 & ~n24219;
  assign n24221 = ~n24218 & ~n24220;
  assign n24222 = n24218 & n24220;
  assign n24223 = ~n24221 & ~n24222;
  assign n24224 = ~n24134 & ~n24137;
  assign n24225 = n24223 & ~n24224;
  assign n24226 = ~n24223 & n24224;
  assign po114  = ~n24225 & ~n24226;
  assign n24228 = ~n24211 & ~n24217;
  assign n24229 = ~n24193 & ~n24198;
  assign n24230 = pi123  & n9858;
  assign n24231 = pi124  & n9508;
  assign n24232 = pi125  & n9503;
  assign n24233 = n9501 & n11786;
  assign n24234 = ~n24231 & ~n24232;
  assign n24235 = ~n24230 & n24234;
  assign n24236 = ~n24233 & n24235;
  assign n24237 = pi56  & n24236;
  assign n24238 = ~pi56  & ~n24236;
  assign n24239 = ~n24237 & ~n24238;
  assign n24240 = ~n24187 & ~n24190;
  assign n24241 = pi120  & n10886;
  assign n24242 = pi121  & n10495;
  assign n24243 = pi122  & n10490;
  assign n24244 = n10488 & n10729;
  assign n24245 = ~n24242 & ~n24243;
  assign n24246 = ~n24241 & n24245;
  assign n24247 = ~n24244 & n24246;
  assign n24248 = pi59  & n24247;
  assign n24249 = ~pi59  & ~n24247;
  assign n24250 = ~n24248 & ~n24249;
  assign n24251 = ~n24181 & ~n24184;
  assign n24252 = ~n24175 & ~n24178;
  assign n24253 = pi116  & n12277;
  assign n24254 = pi115  & n12276;
  assign n24255 = ~n24253 & ~n24254;
  assign n24256 = n24252 & ~n24255;
  assign n24257 = ~n24252 & n24255;
  assign n24258 = ~n24256 & ~n24257;
  assign n24259 = pi117  & n11910;
  assign n24260 = pi118  & n11529;
  assign n24261 = pi119  & n11524;
  assign n24262 = n9412 & n11522;
  assign n24263 = ~n24260 & ~n24261;
  assign n24264 = ~n24259 & n24263;
  assign n24265 = ~n24262 & n24264;
  assign n24266 = pi62  & n24265;
  assign n24267 = ~pi62  & ~n24265;
  assign n24268 = ~n24266 & ~n24267;
  assign n24269 = ~n24258 & n24268;
  assign n24270 = n24258 & ~n24268;
  assign n24271 = ~n24269 & ~n24270;
  assign n24272 = ~n24251 & n24271;
  assign n24273 = n24251 & ~n24271;
  assign n24274 = ~n24272 & ~n24273;
  assign n24275 = ~n24250 & n24274;
  assign n24276 = n24250 & ~n24274;
  assign n24277 = ~n24275 & ~n24276;
  assign n24278 = ~n24240 & n24277;
  assign n24279 = n24240 & ~n24277;
  assign n24280 = ~n24278 & ~n24279;
  assign n24281 = ~n24239 & n24280;
  assign n24282 = n24239 & ~n24280;
  assign n24283 = ~n24281 & ~n24282;
  assign n24284 = ~n24229 & n24283;
  assign n24285 = n24229 & ~n24283;
  assign n24286 = ~n24284 & ~n24285;
  assign n24287 = pi126  & n8905;
  assign n24288 = pi127  & n8535;
  assign n24289 = n8528 & n12542;
  assign n24290 = ~n24287 & ~n24288;
  assign n24291 = ~n24289 & n24290;
  assign n24292 = pi53  & n24291;
  assign n24293 = ~pi53  & ~n24291;
  assign n24294 = ~n24292 & ~n24293;
  assign n24295 = n24286 & ~n24294;
  assign n24296 = ~n24286 & n24294;
  assign n24297 = ~n24295 & ~n24296;
  assign n24298 = n24228 & ~n24297;
  assign n24299 = ~n24228 & n24297;
  assign n24300 = ~n24298 & ~n24299;
  assign n24301 = ~n24222 & ~n24225;
  assign n24302 = n24300 & ~n24301;
  assign n24303 = ~n24300 & n24301;
  assign po115  = ~n24302 & ~n24303;
  assign n24305 = ~n24278 & ~n24281;
  assign n24306 = n8528 & ~n12539;
  assign n24307 = ~n8905 & ~n24306;
  assign n24308 = pi127  & ~n24307;
  assign n24309 = pi53  & ~n24308;
  assign n24310 = ~pi53  & n24308;
  assign n24311 = ~n24309 & ~n24310;
  assign n24312 = ~n24305 & ~n24311;
  assign n24313 = n24305 & n24311;
  assign n24314 = ~n24312 & ~n24313;
  assign n24315 = ~n24272 & ~n24275;
  assign n24316 = pi121  & n10886;
  assign n24317 = pi122  & n10495;
  assign n24318 = pi123  & n10490;
  assign n24319 = n10488 & n10754;
  assign n24320 = ~n24317 & ~n24318;
  assign n24321 = ~n24316 & n24320;
  assign n24322 = ~n24319 & n24321;
  assign n24323 = pi59  & n24322;
  assign n24324 = ~pi59  & ~n24322;
  assign n24325 = ~n24323 & ~n24324;
  assign n24326 = pi118  & n11910;
  assign n24327 = pi119  & n11529;
  assign n24328 = pi120  & n11524;
  assign n24329 = n10047 & n11522;
  assign n24330 = ~n24327 & ~n24328;
  assign n24331 = ~n24326 & n24330;
  assign n24332 = ~n24329 & n24331;
  assign n24333 = pi62  & n24332;
  assign n24334 = ~pi62  & ~n24332;
  assign n24335 = ~n24333 & ~n24334;
  assign n24336 = ~n24257 & ~n24270;
  assign n24337 = pi117  & n12277;
  assign n24338 = pi116  & n12276;
  assign n24339 = ~n24337 & ~n24338;
  assign n24340 = n24255 & ~n24339;
  assign n24341 = ~n24255 & n24339;
  assign n24342 = ~n24340 & ~n24341;
  assign n24343 = ~n24336 & n24342;
  assign n24344 = n24336 & ~n24342;
  assign n24345 = ~n24343 & ~n24344;
  assign n24346 = ~n24335 & n24345;
  assign n24347 = n24335 & ~n24345;
  assign n24348 = ~n24346 & ~n24347;
  assign n24349 = ~n24325 & n24348;
  assign n24350 = n24325 & ~n24348;
  assign n24351 = ~n24349 & ~n24350;
  assign n24352 = n24315 & ~n24351;
  assign n24353 = ~n24315 & n24351;
  assign n24354 = ~n24352 & ~n24353;
  assign n24355 = pi124  & n9858;
  assign n24356 = pi125  & n9508;
  assign n24357 = pi126  & n9503;
  assign n24358 = n9501 & n12148;
  assign n24359 = ~n24356 & ~n24357;
  assign n24360 = ~n24355 & n24359;
  assign n24361 = ~n24358 & n24360;
  assign n24362 = pi56  & n24361;
  assign n24363 = ~pi56  & ~n24361;
  assign n24364 = ~n24362 & ~n24363;
  assign n24365 = n24354 & ~n24364;
  assign n24366 = ~n24354 & n24364;
  assign n24367 = ~n24365 & ~n24366;
  assign n24368 = n24314 & n24367;
  assign n24369 = ~n24314 & ~n24367;
  assign n24370 = ~n24368 & ~n24369;
  assign n24371 = ~n24284 & n24294;
  assign n24372 = ~n24285 & ~n24371;
  assign n24373 = ~n24370 & ~n24372;
  assign n24374 = n24370 & n24372;
  assign n24375 = ~n24373 & ~n24374;
  assign n24376 = ~n24299 & ~n24302;
  assign n24377 = n24375 & ~n24376;
  assign n24378 = ~n24375 & n24376;
  assign po116  = ~n24377 & ~n24378;
  assign n24380 = ~n24374 & ~n24377;
  assign n24381 = pi125  & n9858;
  assign n24382 = pi126  & n9508;
  assign n24383 = pi127  & n9503;
  assign n24384 = n9501 & n12519;
  assign n24385 = ~n24382 & ~n24383;
  assign n24386 = ~n24381 & n24385;
  assign n24387 = ~n24384 & n24386;
  assign n24388 = pi56  & n24387;
  assign n24389 = ~pi56  & ~n24387;
  assign n24390 = ~n24388 & ~n24389;
  assign n24391 = ~n24353 & n24364;
  assign n24392 = ~n24352 & ~n24391;
  assign n24393 = ~n24390 & n24392;
  assign n24394 = n24390 & ~n24392;
  assign n24395 = ~n24393 & ~n24394;
  assign n24396 = ~n24346 & ~n24349;
  assign n24397 = pi122  & n10886;
  assign n24398 = pi123  & n10495;
  assign n24399 = pi124  & n10490;
  assign n24400 = n10488 & n11099;
  assign n24401 = ~n24398 & ~n24399;
  assign n24402 = ~n24397 & n24401;
  assign n24403 = ~n24400 & n24402;
  assign n24404 = pi59  & n24403;
  assign n24405 = ~pi59  & ~n24403;
  assign n24406 = ~n24404 & ~n24405;
  assign n24407 = ~n24341 & ~n24343;
  assign n24408 = ~pi53  & ~n24339;
  assign n24409 = pi53  & n24339;
  assign n24410 = ~n24408 & ~n24409;
  assign n24411 = pi118  & n12277;
  assign n24412 = pi117  & n12276;
  assign n24413 = ~n24411 & ~n24412;
  assign n24414 = ~n24410 & n24413;
  assign n24415 = n24410 & ~n24413;
  assign n24416 = ~n24414 & ~n24415;
  assign n24417 = pi119  & n11910;
  assign n24418 = pi120  & n11529;
  assign n24419 = pi121  & n11524;
  assign n24420 = n10071 & n11522;
  assign n24421 = ~n24418 & ~n24419;
  assign n24422 = ~n24417 & n24421;
  assign n24423 = ~n24420 & n24422;
  assign n24424 = pi62  & n24423;
  assign n24425 = ~pi62  & ~n24423;
  assign n24426 = ~n24424 & ~n24425;
  assign n24427 = n24416 & ~n24426;
  assign n24428 = ~n24416 & n24426;
  assign n24429 = ~n24427 & ~n24428;
  assign n24430 = ~n24407 & n24429;
  assign n24431 = n24407 & ~n24429;
  assign n24432 = ~n24430 & ~n24431;
  assign n24433 = ~n24406 & n24432;
  assign n24434 = n24406 & ~n24432;
  assign n24435 = ~n24433 & ~n24434;
  assign n24436 = ~n24396 & n24435;
  assign n24437 = n24396 & ~n24435;
  assign n24438 = ~n24436 & ~n24437;
  assign n24439 = n24395 & n24438;
  assign n24440 = ~n24395 & ~n24438;
  assign n24441 = ~n24439 & ~n24440;
  assign n24442 = ~n24312 & ~n24367;
  assign n24443 = ~n24313 & ~n24442;
  assign n24444 = n24441 & n24443;
  assign n24445 = ~n24441 & ~n24443;
  assign n24446 = ~n24444 & ~n24445;
  assign n24447 = ~n24380 & n24446;
  assign n24448 = n24380 & ~n24446;
  assign po117  = ~n24447 & ~n24448;
  assign n24450 = ~n24444 & ~n24447;
  assign n24451 = ~n24393 & ~n24439;
  assign n24452 = ~n24433 & ~n24436;
  assign n24453 = pi123  & n10886;
  assign n24454 = pi124  & n10495;
  assign n24455 = pi125  & n10490;
  assign n24456 = n10488 & n11786;
  assign n24457 = ~n24454 & ~n24455;
  assign n24458 = ~n24453 & n24457;
  assign n24459 = ~n24456 & n24458;
  assign n24460 = pi59  & n24459;
  assign n24461 = ~pi59  & ~n24459;
  assign n24462 = ~n24460 & ~n24461;
  assign n24463 = ~n24427 & ~n24430;
  assign n24464 = ~n24408 & ~n24415;
  assign n24465 = pi119  & n12277;
  assign n24466 = pi118  & n12276;
  assign n24467 = ~n24465 & ~n24466;
  assign n24468 = ~n24464 & n24467;
  assign n24469 = n24464 & ~n24467;
  assign n24470 = ~n24468 & ~n24469;
  assign n24471 = pi120  & n11910;
  assign n24472 = pi121  & n11529;
  assign n24473 = pi122  & n11524;
  assign n24474 = n10729 & n11522;
  assign n24475 = ~n24472 & ~n24473;
  assign n24476 = ~n24471 & n24475;
  assign n24477 = ~n24474 & n24476;
  assign n24478 = pi62  & n24477;
  assign n24479 = ~pi62  & ~n24477;
  assign n24480 = ~n24478 & ~n24479;
  assign n24481 = n24470 & ~n24480;
  assign n24482 = ~n24470 & n24480;
  assign n24483 = ~n24481 & ~n24482;
  assign n24484 = ~n24463 & n24483;
  assign n24485 = n24463 & ~n24483;
  assign n24486 = ~n24484 & ~n24485;
  assign n24487 = ~n24462 & n24486;
  assign n24488 = n24462 & ~n24486;
  assign n24489 = ~n24487 & ~n24488;
  assign n24490 = ~n24452 & n24489;
  assign n24491 = n24452 & ~n24489;
  assign n24492 = ~n24490 & ~n24491;
  assign n24493 = pi126  & n9858;
  assign n24494 = pi127  & n9508;
  assign n24495 = n9501 & n12542;
  assign n24496 = ~n24493 & ~n24494;
  assign n24497 = ~n24495 & n24496;
  assign n24498 = pi56  & n24497;
  assign n24499 = ~pi56  & ~n24497;
  assign n24500 = ~n24498 & ~n24499;
  assign n24501 = n24492 & ~n24500;
  assign n24502 = ~n24492 & n24500;
  assign n24503 = ~n24501 & ~n24502;
  assign n24504 = ~n24451 & n24503;
  assign n24505 = n24451 & ~n24503;
  assign n24506 = ~n24504 & ~n24505;
  assign n24507 = ~n24450 & n24506;
  assign n24508 = n24450 & ~n24506;
  assign po118  = ~n24507 & ~n24508;
  assign n24510 = ~n24484 & ~n24487;
  assign n24511 = n9501 & ~n12539;
  assign n24512 = ~n9858 & ~n24511;
  assign n24513 = pi127  & ~n24512;
  assign n24514 = pi56  & ~n24513;
  assign n24515 = ~pi56  & n24513;
  assign n24516 = ~n24514 & ~n24515;
  assign n24517 = ~n24510 & ~n24516;
  assign n24518 = n24510 & n24516;
  assign n24519 = ~n24517 & ~n24518;
  assign n24520 = ~n24468 & ~n24481;
  assign n24521 = pi121  & n11910;
  assign n24522 = pi122  & n11529;
  assign n24523 = pi123  & n11524;
  assign n24524 = n10754 & n11522;
  assign n24525 = ~n24522 & ~n24523;
  assign n24526 = ~n24521 & n24525;
  assign n24527 = ~n24524 & n24526;
  assign n24528 = pi62  & n24527;
  assign n24529 = ~pi62  & ~n24527;
  assign n24530 = ~n24528 & ~n24529;
  assign n24531 = pi120  & n12277;
  assign n24532 = pi119  & n12276;
  assign n24533 = ~n24531 & ~n24532;
  assign n24534 = n24467 & ~n24533;
  assign n24535 = ~n24467 & n24533;
  assign n24536 = ~n24534 & ~n24535;
  assign n24537 = ~n24530 & n24536;
  assign n24538 = n24530 & ~n24536;
  assign n24539 = ~n24537 & ~n24538;
  assign n24540 = n24520 & ~n24539;
  assign n24541 = ~n24520 & n24539;
  assign n24542 = ~n24540 & ~n24541;
  assign n24543 = pi124  & n10886;
  assign n24544 = pi125  & n10495;
  assign n24545 = pi126  & n10490;
  assign n24546 = n10488 & n12148;
  assign n24547 = ~n24544 & ~n24545;
  assign n24548 = ~n24543 & n24547;
  assign n24549 = ~n24546 & n24548;
  assign n24550 = pi59  & n24549;
  assign n24551 = ~pi59  & ~n24549;
  assign n24552 = ~n24550 & ~n24551;
  assign n24553 = n24542 & ~n24552;
  assign n24554 = ~n24542 & n24552;
  assign n24555 = ~n24553 & ~n24554;
  assign n24556 = n24519 & n24555;
  assign n24557 = ~n24519 & ~n24555;
  assign n24558 = ~n24556 & ~n24557;
  assign n24559 = ~n24490 & n24500;
  assign n24560 = ~n24491 & ~n24559;
  assign n24561 = ~n24558 & ~n24560;
  assign n24562 = n24558 & n24560;
  assign n24563 = ~n24561 & ~n24562;
  assign n24564 = ~n24504 & ~n24507;
  assign n24565 = n24563 & ~n24564;
  assign n24566 = ~n24563 & n24564;
  assign po119  = ~n24565 & ~n24566;
  assign n24568 = ~n24534 & ~n24537;
  assign n24569 = pi121  & n12277;
  assign n24570 = pi120  & n12276;
  assign n24571 = ~n24569 & ~n24570;
  assign n24572 = ~pi56  & ~n24571;
  assign n24573 = pi56  & n24571;
  assign n24574 = ~n24572 & ~n24573;
  assign n24575 = ~n24467 & n24574;
  assign n24576 = n24467 & ~n24574;
  assign n24577 = ~n24575 & ~n24576;
  assign n24578 = n24568 & ~n24577;
  assign n24579 = ~n24568 & n24577;
  assign n24580 = ~n24578 & ~n24579;
  assign n24581 = pi122  & n11910;
  assign n24582 = pi123  & n11529;
  assign n24583 = pi124  & n11524;
  assign n24584 = n11099 & n11522;
  assign n24585 = ~n24582 & ~n24583;
  assign n24586 = ~n24581 & n24585;
  assign n24587 = ~n24584 & n24586;
  assign n24588 = pi62  & n24587;
  assign n24589 = ~pi62  & ~n24587;
  assign n24590 = ~n24588 & ~n24589;
  assign n24591 = n24580 & ~n24590;
  assign n24592 = ~n24580 & n24590;
  assign n24593 = ~n24591 & ~n24592;
  assign n24594 = pi125  & n10886;
  assign n24595 = pi126  & n10495;
  assign n24596 = pi127  & n10490;
  assign n24597 = n10488 & n12519;
  assign n24598 = ~n24595 & ~n24596;
  assign n24599 = ~n24594 & n24598;
  assign n24600 = ~n24597 & n24599;
  assign n24601 = pi59  & n24600;
  assign n24602 = ~pi59  & ~n24600;
  assign n24603 = ~n24601 & ~n24602;
  assign n24604 = ~n24541 & n24552;
  assign n24605 = ~n24540 & ~n24604;
  assign n24606 = ~n24603 & n24605;
  assign n24607 = n24603 & ~n24605;
  assign n24608 = ~n24606 & ~n24607;
  assign n24609 = n24593 & n24608;
  assign n24610 = ~n24593 & ~n24608;
  assign n24611 = ~n24609 & ~n24610;
  assign n24612 = ~n24517 & ~n24555;
  assign n24613 = ~n24518 & ~n24612;
  assign n24614 = ~n24611 & ~n24613;
  assign n24615 = n24611 & n24613;
  assign n24616 = ~n24614 & ~n24615;
  assign n24617 = ~n24562 & ~n24565;
  assign n24618 = n24616 & ~n24617;
  assign n24619 = ~n24616 & n24617;
  assign po120  = ~n24618 & ~n24619;
  assign n24621 = ~n24606 & ~n24609;
  assign n24622 = ~n24579 & ~n24591;
  assign n24623 = ~n24572 & ~n24575;
  assign n24624 = pi122  & n12277;
  assign n24625 = pi121  & n12276;
  assign n24626 = ~n24624 & ~n24625;
  assign n24627 = n24623 & ~n24626;
  assign n24628 = ~n24623 & n24626;
  assign n24629 = ~n24627 & ~n24628;
  assign n24630 = pi123  & n11910;
  assign n24631 = pi124  & n11529;
  assign n24632 = pi125  & n11524;
  assign n24633 = n11522 & n11786;
  assign n24634 = ~n24631 & ~n24632;
  assign n24635 = ~n24630 & n24634;
  assign n24636 = ~n24633 & n24635;
  assign n24637 = pi62  & n24636;
  assign n24638 = ~pi62  & ~n24636;
  assign n24639 = ~n24637 & ~n24638;
  assign n24640 = n24629 & ~n24639;
  assign n24641 = ~n24629 & n24639;
  assign n24642 = ~n24640 & ~n24641;
  assign n24643 = ~n24622 & n24642;
  assign n24644 = n24622 & ~n24642;
  assign n24645 = ~n24643 & ~n24644;
  assign n24646 = pi126  & n10886;
  assign n24647 = pi127  & n10495;
  assign n24648 = n10488 & n12542;
  assign n24649 = ~n24646 & ~n24647;
  assign n24650 = ~n24648 & n24649;
  assign n24651 = pi59  & n24650;
  assign n24652 = ~pi59  & ~n24650;
  assign n24653 = ~n24651 & ~n24652;
  assign n24654 = n24645 & ~n24653;
  assign n24655 = ~n24645 & n24653;
  assign n24656 = ~n24654 & ~n24655;
  assign n24657 = n24621 & ~n24656;
  assign n24658 = ~n24621 & n24656;
  assign n24659 = ~n24657 & ~n24658;
  assign n24660 = ~n24615 & ~n24618;
  assign n24661 = n24659 & ~n24660;
  assign n24662 = ~n24659 & n24660;
  assign po121  = ~n24661 & ~n24662;
  assign n24664 = ~n24658 & ~n24661;
  assign n24665 = ~n24628 & ~n24640;
  assign n24666 = pi123  & n12277;
  assign n24667 = pi122  & n12276;
  assign n24668 = ~n24666 & ~n24667;
  assign n24669 = n24626 & ~n24668;
  assign n24670 = ~n24626 & n24668;
  assign n24671 = ~n24669 & ~n24670;
  assign n24672 = ~n24665 & n24671;
  assign n24673 = n24665 & ~n24671;
  assign n24674 = ~n24672 & ~n24673;
  assign n24675 = pi124  & n11910;
  assign n24676 = pi125  & n11529;
  assign n24677 = pi126  & n11524;
  assign n24678 = n11522 & n12148;
  assign n24679 = ~n24676 & ~n24677;
  assign n24680 = ~n24675 & n24679;
  assign n24681 = ~n24678 & n24680;
  assign n24682 = pi62  & n24681;
  assign n24683 = ~pi62  & ~n24681;
  assign n24684 = ~n24682 & ~n24683;
  assign n24685 = n10488 & ~n12539;
  assign n24686 = ~n10886 & ~n24685;
  assign n24687 = pi127  & ~n24686;
  assign n24688 = pi59  & ~n24687;
  assign n24689 = ~pi59  & n24687;
  assign n24690 = ~n24688 & ~n24689;
  assign n24691 = ~n24684 & ~n24690;
  assign n24692 = n24684 & n24690;
  assign n24693 = ~n24691 & ~n24692;
  assign n24694 = n24674 & n24693;
  assign n24695 = ~n24674 & ~n24693;
  assign n24696 = ~n24694 & ~n24695;
  assign n24697 = ~n24643 & n24653;
  assign n24698 = ~n24644 & ~n24697;
  assign n24699 = n24696 & n24698;
  assign n24700 = ~n24696 & ~n24698;
  assign n24701 = ~n24699 & ~n24700;
  assign n24702 = ~n24664 & n24701;
  assign n24703 = n24664 & ~n24701;
  assign po122  = ~n24702 & ~n24703;
  assign n24705 = ~n24699 & ~n24702;
  assign n24706 = ~n24691 & ~n24694;
  assign n24707 = ~n24670 & ~n24672;
  assign n24708 = ~pi59  & ~n24668;
  assign n24709 = pi59  & n24668;
  assign n24710 = ~n24708 & ~n24709;
  assign n24711 = pi124  & n12277;
  assign n24712 = pi123  & n12276;
  assign n24713 = ~n24711 & ~n24712;
  assign n24714 = ~n24710 & n24713;
  assign n24715 = n24710 & ~n24713;
  assign n24716 = ~n24714 & ~n24715;
  assign n24717 = pi125  & n11910;
  assign n24718 = pi126  & n11529;
  assign n24719 = pi127  & n11524;
  assign n24720 = n11522 & n12519;
  assign n24721 = ~n24718 & ~n24719;
  assign n24722 = ~n24717 & n24721;
  assign n24723 = ~n24720 & n24722;
  assign n24724 = pi62  & n24723;
  assign n24725 = ~pi62  & ~n24723;
  assign n24726 = ~n24724 & ~n24725;
  assign n24727 = n24716 & ~n24726;
  assign n24728 = ~n24716 & n24726;
  assign n24729 = ~n24727 & ~n24728;
  assign n24730 = ~n24707 & n24729;
  assign n24731 = n24707 & ~n24729;
  assign n24732 = ~n24730 & ~n24731;
  assign n24733 = ~n24706 & n24732;
  assign n24734 = n24706 & ~n24732;
  assign n24735 = ~n24733 & ~n24734;
  assign n24736 = ~n24705 & n24735;
  assign n24737 = n24705 & ~n24735;
  assign po123  = ~n24736 & ~n24737;
  assign n24739 = ~n24733 & ~n24736;
  assign n24740 = ~n24727 & ~n24730;
  assign n24741 = ~n24708 & ~n24715;
  assign n24742 = pi125  & n12277;
  assign n24743 = pi124  & n12276;
  assign n24744 = ~n24742 & ~n24743;
  assign n24745 = ~n24741 & n24744;
  assign n24746 = n24741 & ~n24744;
  assign n24747 = ~n24745 & ~n24746;
  assign n24748 = pi126  & n11910;
  assign n24749 = pi127  & n11529;
  assign n24750 = n11522 & n12542;
  assign n24751 = ~n24748 & ~n24749;
  assign n24752 = ~n24750 & n24751;
  assign n24753 = pi62  & n24752;
  assign n24754 = ~pi62  & ~n24752;
  assign n24755 = ~n24753 & ~n24754;
  assign n24756 = n24747 & ~n24755;
  assign n24757 = ~n24747 & n24755;
  assign n24758 = ~n24756 & ~n24757;
  assign n24759 = ~n24740 & n24758;
  assign n24760 = n24740 & ~n24758;
  assign n24761 = ~n24759 & ~n24760;
  assign n24762 = ~n24739 & n24761;
  assign n24763 = n24739 & ~n24761;
  assign po124  = ~n24762 & ~n24763;
  assign n24765 = ~n24759 & ~n24762;
  assign n24766 = ~n24745 & ~n24756;
  assign n24767 = pi126  & n12277;
  assign n24768 = pi125  & n12276;
  assign n24769 = ~n24767 & ~n24768;
  assign n24770 = n24744 & ~n24769;
  assign n24771 = ~n24744 & n24769;
  assign n24772 = ~n24770 & ~n24771;
  assign n24773 = n11522 & ~n12539;
  assign n24774 = ~n11910 & ~n24773;
  assign n24775 = pi127  & ~n24774;
  assign n24776 = pi62  & ~n24775;
  assign n24777 = ~pi62  & n24775;
  assign n24778 = ~n24776 & ~n24777;
  assign n24779 = n24772 & ~n24778;
  assign n24780 = ~n24772 & n24778;
  assign n24781 = ~n24779 & ~n24780;
  assign n24782 = ~n24766 & n24781;
  assign n24783 = n24766 & ~n24781;
  assign n24784 = ~n24782 & ~n24783;
  assign n24785 = ~n24765 & n24784;
  assign n24786 = n24765 & ~n24784;
  assign po125  = ~n24785 & ~n24786;
  assign n24788 = ~n24782 & ~n24785;
  assign n24789 = ~n24770 & ~n24779;
  assign n24790 = pi63  & pi127 ;
  assign n24791 = pi62  & ~pi127 ;
  assign n24792 = ~n24790 & ~n24791;
  assign n24793 = pi62  & pi126 ;
  assign n24794 = n12276 & n24793;
  assign n24795 = ~n24792 & ~n24794;
  assign n24796 = ~n24744 & ~n24795;
  assign n24797 = n24744 & n24795;
  assign n24798 = ~n24796 & ~n24797;
  assign n24799 = ~n24789 & n24798;
  assign n24800 = n24789 & ~n24798;
  assign n24801 = ~n24799 & ~n24800;
  assign n24802 = ~n24788 & n24801;
  assign n24803 = n24788 & ~n24801;
  assign po126  = ~n24802 & ~n24803;
  assign n24805 = ~n24799 & ~n24802;
  assign n24806 = n24790 & ~n24796;
  assign n24807 = pi62  & n24790;
  assign n24808 = n24796 & ~n24807;
  assign n24809 = ~n24806 & ~n24808;
  assign n24810 = n24805 & ~n24809;
  assign n24811 = ~n24805 & n24809;
  assign po127  = ~n24810 & ~n24811;
endmodule
