module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 , pi32 ,
    pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 , pi40 ,
    pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 , pi56 ,
    pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 , pi64 ,
    pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 , pi73 ,
    pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 , pi81 ,
    pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 , pi89 ,
    pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 , pi97 ,
    pi98 , pi99 , pi100 , pi101 , pi102 , pi103 , pi104 , pi105 ,
    pi106 , pi107 , pi108 , pi109 , pi110 , pi111 , pi112 , pi113 ,
    pi114 , pi115 , pi116 , pi117 , pi118 , pi119 , pi120 , pi121 ,
    pi122 , pi123 , pi124 , pi125 , pi126 , pi127 ,
    po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7 , po8 ,
    po9 , po10 , po11 , po12 , po13 , po14 , po15 , po16 ,
    po17 , po18 , po19 , po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 , po30 , po31 , po32 ,
    po33 , po34 , po35 , po36 , po37 , po38 , po39 , po40 ,
    po41 , po42 , po43 , po44 , po45 , po46 , po47 , po48 ,
    po49 , po50 , po51 , po52 , po53 , po54 , po55 , po56 ,
    po57 , po58 , po59 , po60 , po61 , po62 , po63 , po64 ,
    po65 , po66 , po67 , po68 , po69 , po70 , po71 , po72 ,
    po73 , po74 , po75 , po76 , po77 , po78 , po79 , po80 ,
    po81 , po82 , po83 , po84 , po85 , po86 , po87 , po88 ,
    po89 , po90 , po91 , po92 , po93 , po94 , po95 , po96 ,
    po97 , po98 , po99 , po100 , po101 , po102 , po103 ,
    po104 , po105 , po106 , po107 , po108 , po109 , po110 ,
    po111 , po112 , po113 , po114 , po115 , po116 , po117 ,
    po118 , po119 , po120 , po121 , po122 , po123 , po124 ,
    po125 , po126 , po127   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    pi32 , pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 ,
    pi56 , pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 ,
    pi64 , pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 ,
    pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 ,
    pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 ,
    pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 ,
    pi97 , pi98 , pi99 , pi100 , pi101 , pi102 , pi103 , pi104 ,
    pi105 , pi106 , pi107 , pi108 , pi109 , pi110 , pi111 , pi112 ,
    pi113 , pi114 , pi115 , pi116 , pi117 , pi118 , pi119 , pi120 ,
    pi121 , pi122 , pi123 , pi124 , pi125 , pi126 , pi127 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7 ,
    po8 , po9 , po10 , po11 , po12 , po13 , po14 , po15 ,
    po16 , po17 , po18 , po19 , po20 , po21 , po22 , po23 ,
    po24 , po25 , po26 , po27 , po28 , po29 , po30 , po31 ,
    po32 , po33 , po34 , po35 , po36 , po37 , po38 , po39 ,
    po40 , po41 , po42 , po43 , po44 , po45 , po46 , po47 ,
    po48 , po49 , po50 , po51 , po52 , po53 , po54 , po55 ,
    po56 , po57 , po58 , po59 , po60 , po61 , po62 , po63 ,
    po64 , po65 , po66 , po67 , po68 , po69 , po70 , po71 ,
    po72 , po73 , po74 , po75 , po76 , po77 , po78 , po79 ,
    po80 , po81 , po82 , po83 , po84 , po85 , po86 , po87 ,
    po88 , po89 , po90 , po91 , po92 , po93 , po94 , po95 ,
    po96 , po97 , po98 , po99 , po100 , po101 , po102 ,
    po103 , po104 , po105 , po106 , po107 , po108 , po109 ,
    po110 , po111 , po112 , po113 , po114 , po115 , po116 ,
    po117 , po118 , po119 , po120 , po121 , po122 , po123 ,
    po124 , po125 , po126 , po127 ;
  wire n257, n258, n259, n260, n261, n262, n263,
    n264, n265, n266, n267, n268, n269, n270,
    n271, n272, n273, n274, n275, n276, n277,
    n278, n279, n280, n281, n282, n283, n284,
    n285, n286, n287, n288, n289, n290, n291,
    n292, n293, n294, n295, n296, n297, n298,
    n299, n300, n301, n302, n303, n304, n305,
    n306, n307, n308, n309, n310, n311, n312,
    n313, n314, n315, n316, n317, n318, n319,
    n320, n321, n322, n323, n324, n325, n326,
    n327, n328, n329, n330, n331, n332, n333,
    n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403,
    n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416, n417,
    n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438,
    n439, n440, n441, n442, n443, n444, n445,
    n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487,
    n488, n489, n490, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501,
    n502, n503, n504, n505, n506, n507, n508,
    n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n541, n542, n543,
    n544, n545, n546, n547, n548, n549, n550,
    n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564,
    n565, n566, n567, n568, n569, n570, n571,
    n572, n573, n574, n575, n576, n577, n578,
    n579, n580, n581, n582, n583, n584, n585,
    n586, n587, n588, n589, n590, n591, n592,
    n593, n594, n595, n596, n597, n598, n599,
    n600, n601, n602, n603, n604, n605, n606,
    n607, n608, n609, n610, n611, n612, n613,
    n614, n615, n616, n617, n618, n619, n620,
    n621, n622, n623, n624, n625, n626, n627,
    n628, n629, n630, n631, n632, n633, n634,
    n635, n636, n637, n638, n639, n640, n641,
    n642, n643, n644, n645, n646, n647, n648,
    n649, n650, n651, n652, n653, n654, n655,
    n656, n657, n658, n659, n660, n661, n662,
    n663, n664, n665, n666, n667, n668, n669,
    n670, n671, n672, n673, n674, n675, n676,
    n677, n678, n679, n680, n681, n682, n683,
    n684, n685, n686, n687, n688, n689, n690,
    n691, n692, n693, n694, n695, n696, n697,
    n698, n699, n700, n701, n702, n703, n704,
    n705, n706, n707, n708, n709, n710, n711,
    n712, n713, n714, n715, n716, n717, n718,
    n719, n720, n721, n722, n723, n724, n725,
    n726, n727, n728, n729, n730, n731, n732,
    n733, n734, n735, n736, n737, n738, n739,
    n740, n741, n742, n743, n744, n745, n746,
    n747, n748, n749, n750, n751, n752, n753,
    n754, n755, n756, n757, n758, n759, n760,
    n761, n762, n763, n764, n765, n766, n767,
    n768, n769, n770, n771, n772, n773, n774,
    n775, n776, n777, n778, n779, n780, n781,
    n782, n783, n784, n785, n786, n787, n788,
    n789, n790, n791, n792, n793, n794, n795,
    n796, n797, n798, n799, n800, n801, n802,
    n803, n804, n805, n806, n807, n808, n809,
    n810, n811, n812, n813, n814, n815, n816,
    n817, n818, n819, n820, n821, n822, n823,
    n824, n825, n826, n827, n828, n829, n830,
    n831, n832, n833, n834, n835, n836, n837,
    n838, n839, n840, n841, n842, n843, n844,
    n845, n846, n847, n848, n849, n850, n851,
    n852, n853, n854, n855, n856, n857, n858,
    n859, n860, n861, n862, n863, n864, n865,
    n866, n867, n868, n869, n870, n871, n872,
    n873, n874, n875, n876, n877, n878, n879,
    n880, n881, n882, n883, n884, n885, n886,
    n887, n888, n889, n890, n891, n892, n893,
    n894, n895, n896, n897, n898, n899, n900,
    n901, n902, n903, n904, n905, n906, n907,
    n908, n909, n910, n911, n912, n913, n914,
    n915, n916, n917, n918, n919, n920, n921,
    n922, n923, n924, n925, n926, n927, n928,
    n929, n930, n931, n932, n933, n934, n935,
    n936, n937, n938, n939, n940, n941, n942,
    n943, n944, n945, n946, n947, n948, n949,
    n950, n951, n952, n953, n954, n955, n956,
    n957, n958, n959, n960, n961, n962, n963,
    n964, n965, n966, n967, n968, n969, n970,
    n971, n972, n973, n974, n975, n976, n977,
    n978, n979, n980, n981, n982, n983, n984,
    n985, n986, n987, n988, n989, n990, n991,
    n992, n993, n994, n995, n996, n997, n998,
    n999, n1000, n1001, n1002, n1003, n1004,
    n1005, n1006, n1007, n1008, n1009, n1010,
    n1011, n1012, n1013, n1014, n1015, n1016,
    n1017, n1018, n1019, n1020, n1021, n1022,
    n1023, n1024, n1025, n1026, n1027, n1028,
    n1029, n1030, n1031, n1032, n1033, n1034,
    n1035, n1036, n1037, n1038, n1039, n1040,
    n1041, n1042, n1043, n1044, n1045, n1046,
    n1047, n1048, n1049, n1050, n1051, n1052,
    n1053, n1054, n1055, n1056, n1057, n1058,
    n1059, n1060, n1061, n1062, n1063, n1064,
    n1065, n1066, n1067, n1068, n1069, n1070,
    n1071, n1072, n1073, n1074, n1075, n1076,
    n1077, n1078, n1079, n1080, n1081, n1082,
    n1083, n1084, n1085, n1086, n1087, n1088,
    n1089, n1090, n1091, n1092, n1093, n1094,
    n1095, n1096, n1097, n1098, n1099, n1100,
    n1101, n1102, n1103, n1104, n1105, n1106,
    n1107, n1108, n1109, n1110, n1111, n1112,
    n1113, n1114, n1115, n1116, n1117, n1118,
    n1119, n1120, n1121, n1122, n1123, n1124,
    n1125, n1126, n1127, n1128, n1129, n1130,
    n1131, n1132, n1133, n1134, n1135, n1136,
    n1137, n1138, n1139, n1140, n1141, n1142,
    n1143, n1144, n1145, n1146, n1147, n1148,
    n1149, n1150, n1151, n1152, n1153, n1154,
    n1155, n1156, n1157, n1158, n1159, n1160,
    n1161, n1162, n1163, n1164, n1165, n1166,
    n1167, n1168, n1169, n1170, n1171, n1172,
    n1173, n1174, n1175, n1176, n1177, n1178,
    n1179, n1180, n1181, n1182, n1183, n1184,
    n1185, n1186, n1187, n1188, n1189, n1190,
    n1191, n1192, n1193, n1194, n1195, n1196,
    n1197, n1198, n1199, n1200, n1201, n1202,
    n1203, n1204, n1205, n1206, n1207, n1208,
    n1209, n1210, n1211, n1212, n1213, n1214,
    n1215, n1216, n1217, n1218, n1219, n1220,
    n1221, n1222, n1223, n1224, n1225, n1226,
    n1227, n1228, n1229, n1230, n1231, n1232,
    n1233, n1234, n1235, n1236, n1237, n1238,
    n1239, n1240, n1241, n1242, n1243, n1244,
    n1245, n1246, n1247, n1248, n1249, n1250,
    n1251, n1252, n1253, n1254, n1255, n1256,
    n1257, n1258, n1259, n1260, n1261, n1262,
    n1263, n1264, n1265, n1266, n1267, n1268,
    n1269, n1270, n1271, n1272, n1273, n1274,
    n1275, n1276, n1277, n1278, n1279, n1280,
    n1281, n1282, n1283, n1284, n1285, n1286,
    n1287, n1288, n1289, n1290, n1291, n1292,
    n1293, n1294, n1295, n1296, n1297, n1298,
    n1299, n1300, n1301, n1302, n1303, n1304,
    n1305, n1306, n1307, n1308, n1309, n1310,
    n1311, n1312, n1313, n1314, n1315, n1316,
    n1317, n1318, n1319, n1320, n1321, n1322,
    n1323, n1324, n1325, n1326, n1327, n1328,
    n1329, n1330, n1331, n1332, n1333, n1334,
    n1335, n1336, n1337, n1338, n1339, n1340,
    n1341, n1342, n1343, n1344, n1345, n1346,
    n1347, n1348, n1349, n1350, n1351, n1352,
    n1353, n1354, n1355, n1356, n1357, n1358,
    n1359, n1360, n1361, n1362, n1363, n1364,
    n1365, n1366, n1367, n1368, n1369, n1370,
    n1371, n1372, n1373, n1374, n1375, n1376,
    n1377, n1378, n1379, n1380, n1381, n1382,
    n1383, n1384, n1385, n1386, n1387, n1388,
    n1389, n1390, n1391, n1392, n1393, n1394,
    n1395, n1396, n1397, n1398, n1399, n1400,
    n1401, n1402, n1403, n1404, n1405, n1406,
    n1407, n1408, n1409, n1410, n1411, n1412,
    n1413, n1414, n1415, n1416, n1417, n1418,
    n1419, n1420, n1421, n1422, n1423, n1424,
    n1425, n1426, n1427, n1428, n1429, n1430,
    n1431, n1432, n1433, n1434, n1435, n1436,
    n1437, n1438, n1439, n1440, n1441, n1442,
    n1443, n1444, n1445, n1446, n1447, n1448,
    n1449, n1450, n1451, n1452, n1453, n1454,
    n1455, n1456, n1457, n1458, n1459, n1460,
    n1461, n1462, n1463, n1464, n1465, n1466,
    n1467, n1468, n1469, n1470, n1471, n1472,
    n1473, n1474, n1475, n1476, n1477, n1478,
    n1479, n1480, n1481, n1482, n1483, n1484,
    n1485, n1486, n1487, n1488, n1489, n1490,
    n1491, n1492, n1493, n1494, n1495, n1496,
    n1497, n1498, n1499, n1500, n1501, n1502,
    n1503, n1504, n1505, n1506, n1507, n1508,
    n1509, n1510, n1511, n1512, n1513, n1514,
    n1515, n1516, n1517, n1518, n1519, n1520,
    n1521, n1522, n1523, n1524, n1525, n1526,
    n1527, n1528, n1529, n1530, n1531, n1532,
    n1533, n1534, n1535, n1536, n1537, n1538,
    n1539, n1540, n1541, n1542, n1543, n1544,
    n1545, n1546, n1547, n1548, n1549, n1550,
    n1551, n1552, n1553, n1554, n1555, n1556,
    n1557, n1558, n1559, n1560, n1561, n1562,
    n1563, n1564, n1565, n1566, n1567, n1568,
    n1569, n1570, n1571, n1572, n1573, n1574,
    n1575, n1576, n1577, n1578, n1579, n1580,
    n1581, n1582, n1583, n1584, n1585, n1586,
    n1587, n1588, n1589, n1590, n1591, n1592,
    n1593, n1594, n1595, n1596, n1597, n1598,
    n1599, n1600, n1601, n1602, n1603, n1604,
    n1605, n1606, n1607, n1608, n1609, n1610,
    n1611, n1612, n1613, n1614, n1615, n1616,
    n1617, n1618, n1619, n1620, n1621, n1622,
    n1623, n1624, n1625, n1626, n1627, n1628,
    n1629, n1630, n1631, n1632, n1633, n1634,
    n1635, n1636, n1637, n1638, n1639, n1640,
    n1641, n1642, n1643, n1644, n1645, n1646,
    n1647, n1648, n1649, n1650, n1651, n1652,
    n1653, n1654, n1655, n1656, n1657, n1658,
    n1659, n1660, n1661, n1662, n1663, n1664,
    n1665, n1666, n1667, n1668, n1669, n1670,
    n1671, n1672, n1673, n1674, n1675, n1676,
    n1677, n1678, n1679, n1680, n1681, n1682,
    n1683, n1684, n1685, n1686, n1687, n1688,
    n1689, n1690, n1691, n1692, n1693, n1694,
    n1695, n1696, n1697, n1698, n1699, n1700,
    n1701, n1702, n1703, n1704, n1705, n1706,
    n1707, n1708, n1709, n1710, n1711, n1712,
    n1713, n1714, n1715, n1716, n1717, n1718,
    n1719, n1720, n1721, n1722, n1723, n1724,
    n1725, n1726, n1727, n1728, n1729, n1730,
    n1731, n1732, n1733, n1734, n1735, n1736,
    n1737, n1738, n1739, n1740, n1741, n1742,
    n1743, n1744, n1745, n1746, n1747, n1748,
    n1749, n1750, n1751, n1752, n1753, n1754,
    n1755, n1756, n1757, n1758, n1759, n1760,
    n1761, n1762, n1763, n1764, n1765, n1766,
    n1767, n1768, n1769, n1770, n1771, n1772,
    n1773, n1774, n1775, n1776, n1777, n1778,
    n1779, n1780, n1781, n1782, n1783, n1784,
    n1785, n1786, n1787, n1788, n1789, n1790,
    n1791, n1792, n1793, n1794, n1795, n1796,
    n1797, n1798, n1799, n1800, n1801, n1802,
    n1803, n1804, n1805, n1806, n1807, n1808,
    n1809, n1810, n1811, n1812, n1813, n1814,
    n1815, n1816, n1817, n1818, n1819, n1820,
    n1821, n1822, n1823, n1824, n1825, n1826,
    n1827, n1828, n1829, n1830, n1831, n1832,
    n1833, n1834, n1835, n1836, n1837, n1838,
    n1839, n1840, n1841, n1842, n1843, n1844,
    n1845, n1846, n1847, n1848, n1849, n1850,
    n1851, n1852, n1853, n1854, n1855, n1856,
    n1857, n1858, n1859, n1860, n1861, n1862,
    n1863, n1864, n1865, n1866, n1867, n1868,
    n1869, n1870, n1871, n1872, n1873, n1874,
    n1875, n1876, n1877, n1878, n1879, n1880,
    n1881, n1882, n1883, n1884, n1885, n1886,
    n1887, n1888, n1889, n1890, n1891, n1892,
    n1893, n1894, n1895, n1896, n1897, n1898,
    n1899, n1900, n1901, n1902, n1903, n1904,
    n1905, n1906, n1907, n1908, n1909, n1910,
    n1911, n1912, n1913, n1914, n1915, n1916,
    n1917, n1918, n1919, n1920, n1921, n1922,
    n1923, n1924, n1925, n1926, n1927, n1928,
    n1929, n1930, n1931, n1932, n1933, n1934,
    n1935, n1936, n1937, n1938, n1939, n1940,
    n1941, n1942, n1943, n1944, n1945, n1946,
    n1947, n1948, n1949, n1950, n1951, n1952,
    n1953, n1954, n1955, n1956, n1957, n1958,
    n1959, n1960, n1961, n1962, n1963, n1964,
    n1965, n1966, n1967, n1968, n1969, n1970,
    n1971, n1972, n1973, n1974, n1975, n1976,
    n1977, n1978, n1979, n1980, n1981, n1982,
    n1983, n1984, n1985, n1986, n1987, n1988,
    n1989, n1990, n1991, n1992, n1993, n1994,
    n1995, n1996, n1997, n1998, n1999, n2000,
    n2001, n2002, n2003, n2004, n2005, n2006,
    n2007, n2008, n2009, n2010, n2011, n2012,
    n2013, n2014, n2015, n2016, n2017, n2018,
    n2019, n2020, n2021, n2022, n2023, n2024,
    n2025, n2026, n2027, n2028, n2029, n2030,
    n2031, n2032, n2033, n2034, n2035, n2036,
    n2037, n2038, n2039, n2040, n2041, n2042,
    n2043, n2044, n2045, n2046, n2047, n2048,
    n2049, n2050, n2051, n2052, n2053, n2054,
    n2055, n2056, n2057, n2058, n2059, n2060,
    n2061, n2062, n2063, n2064, n2065, n2066,
    n2067, n2068, n2069, n2070, n2071, n2072,
    n2073, n2074, n2075, n2076, n2077, n2078,
    n2079, n2080, n2081, n2082, n2083, n2084,
    n2085, n2086, n2087, n2088, n2089, n2090,
    n2091, n2092, n2093, n2094, n2095, n2096,
    n2097, n2098, n2099, n2100, n2101, n2102,
    n2103, n2104, n2105, n2106, n2107, n2108,
    n2109, n2110, n2111, n2112, n2113, n2114,
    n2115, n2116, n2117, n2118, n2119, n2120,
    n2121, n2122, n2123, n2124, n2125, n2126,
    n2127, n2128, n2129, n2130, n2131, n2132,
    n2133, n2134, n2135, n2136, n2137, n2138,
    n2139, n2140, n2141, n2142, n2143, n2144,
    n2145, n2146, n2147, n2148, n2149, n2150,
    n2151, n2152, n2153, n2154, n2155, n2156,
    n2157, n2158, n2159, n2160, n2161, n2162,
    n2163, n2164, n2165, n2166, n2167, n2168,
    n2169, n2170, n2171, n2172, n2173, n2174,
    n2175, n2176, n2177, n2178, n2179, n2180,
    n2181, n2182, n2183, n2184, n2185, n2186,
    n2187, n2188, n2189, n2190, n2191, n2192,
    n2193, n2194, n2195, n2196, n2197, n2198,
    n2199, n2200, n2201, n2202, n2203, n2204,
    n2205, n2206, n2207, n2208, n2209, n2210,
    n2211, n2212, n2213, n2214, n2215, n2216,
    n2217, n2218, n2219, n2220, n2221, n2222,
    n2223, n2224, n2225, n2226, n2227, n2228,
    n2229, n2230, n2231, n2232, n2233, n2234,
    n2235, n2236, n2237, n2238, n2239, n2240,
    n2241, n2242, n2243, n2244, n2245, n2246,
    n2247, n2248, n2249, n2250, n2251, n2252,
    n2253, n2254, n2255, n2256, n2257, n2258,
    n2259, n2260, n2261, n2262, n2263, n2264,
    n2265, n2266, n2267, n2268, n2269, n2270,
    n2271, n2272, n2273, n2274, n2275, n2276,
    n2277, n2278, n2279, n2280, n2281, n2282,
    n2283, n2284, n2285, n2286, n2287, n2288,
    n2289, n2290, n2291, n2292, n2293, n2294,
    n2295, n2296, n2297, n2298, n2299, n2300,
    n2301, n2302, n2303, n2304, n2305, n2306,
    n2307, n2308, n2309, n2310, n2311, n2312,
    n2313, n2314, n2315, n2316, n2317, n2318,
    n2319, n2320, n2321, n2322, n2323, n2324,
    n2325, n2326, n2327, n2328, n2329, n2330,
    n2331, n2332, n2333, n2334, n2335, n2336,
    n2337, n2338, n2339, n2340, n2341, n2342,
    n2343, n2344, n2345, n2346, n2347, n2348,
    n2349, n2350, n2351, n2352, n2353, n2354,
    n2355, n2356, n2357, n2358, n2359, n2360,
    n2361, n2362, n2363, n2364, n2365, n2366,
    n2367, n2368, n2369, n2370, n2371, n2372,
    n2373, n2374, n2375, n2376, n2377, n2378,
    n2379, n2380, n2381, n2382, n2383, n2384,
    n2385, n2386, n2387, n2388, n2389, n2390,
    n2391, n2392, n2393, n2394, n2395, n2396,
    n2397, n2398, n2399, n2400, n2401, n2402,
    n2403, n2404, n2405, n2406, n2407, n2408,
    n2409, n2410, n2411, n2412, n2413, n2414,
    n2415, n2416, n2417, n2418, n2419, n2420,
    n2421, n2422, n2423, n2424, n2425, n2426,
    n2427, n2428, n2429, n2430, n2431, n2432,
    n2433, n2434, n2435, n2436, n2437, n2438,
    n2439, n2440, n2441, n2442, n2443, n2444,
    n2445, n2446, n2447, n2448, n2449, n2450,
    n2451, n2452, n2453, n2454, n2455, n2456,
    n2457, n2458, n2459, n2460, n2461, n2462,
    n2463, n2464, n2465, n2466, n2467, n2468,
    n2469, n2470, n2471, n2472, n2473, n2474,
    n2475, n2476, n2477, n2478, n2479, n2480,
    n2481, n2482, n2483, n2484, n2485, n2486,
    n2487, n2488, n2489, n2490, n2491, n2492,
    n2493, n2494, n2495, n2496, n2497, n2498,
    n2499, n2500, n2501, n2502, n2503, n2504,
    n2505, n2506, n2507, n2508, n2509, n2510,
    n2511, n2512, n2513, n2514, n2515, n2516,
    n2517, n2518, n2519, n2520, n2521, n2522,
    n2523, n2524, n2525, n2526, n2527, n2528,
    n2529, n2530, n2531, n2532, n2533, n2534,
    n2535, n2536, n2537, n2538, n2539, n2540,
    n2541, n2542, n2543, n2544, n2545, n2546,
    n2547, n2548, n2549, n2550, n2551, n2552,
    n2553, n2554, n2555, n2556, n2557, n2558,
    n2559, n2560, n2561, n2562, n2563, n2564,
    n2565, n2566, n2567, n2568, n2569, n2570,
    n2571, n2572, n2573, n2574, n2575, n2576,
    n2577, n2578, n2579, n2580, n2581, n2582,
    n2583, n2584, n2585, n2586, n2587, n2588,
    n2589, n2590, n2591, n2592, n2593, n2594,
    n2595, n2596, n2597, n2598, n2599, n2600,
    n2601, n2602, n2603, n2604, n2605, n2606,
    n2607, n2608, n2609, n2610, n2611, n2612,
    n2613, n2614, n2615, n2616, n2617, n2618,
    n2619, n2620, n2621, n2622, n2623, n2624,
    n2625, n2626, n2627, n2628, n2629, n2630,
    n2631, n2632, n2633, n2634, n2635, n2636,
    n2637, n2638, n2639, n2640, n2641, n2642,
    n2643, n2644, n2645, n2646, n2647, n2648,
    n2649, n2650, n2651, n2652, n2653, n2654,
    n2655, n2656, n2657, n2658, n2659, n2660,
    n2661, n2662, n2663, n2664, n2665, n2666,
    n2667, n2668, n2669, n2670, n2671, n2672,
    n2673, n2674, n2675, n2676, n2677, n2678,
    n2679, n2680, n2681, n2682, n2683, n2684,
    n2685, n2686, n2687, n2688, n2689, n2690,
    n2691, n2692, n2693, n2694, n2695, n2696,
    n2697, n2698, n2699, n2700, n2701, n2702,
    n2703, n2704, n2705, n2706, n2707, n2708,
    n2709, n2710, n2711, n2712, n2713, n2714,
    n2715, n2716, n2717, n2718, n2719, n2720,
    n2721, n2722, n2723, n2724, n2725, n2726,
    n2727, n2728, n2729, n2730, n2731, n2732,
    n2733, n2734, n2735, n2736, n2737, n2738,
    n2739, n2740, n2741, n2742, n2743, n2744,
    n2745, n2746, n2747, n2748, n2749, n2750,
    n2751, n2752, n2753, n2754, n2755, n2756,
    n2757, n2758, n2759, n2760, n2761, n2762,
    n2763, n2764, n2765, n2766, n2767, n2768,
    n2769, n2770, n2771, n2772, n2773, n2774,
    n2775, n2776, n2777, n2778, n2779, n2780,
    n2781, n2782, n2783, n2784, n2785, n2786,
    n2787, n2788, n2789, n2790, n2791, n2792,
    n2793, n2794, n2795, n2796, n2797, n2798,
    n2799, n2800, n2801, n2802, n2803, n2804,
    n2805, n2806, n2807, n2808, n2809, n2810,
    n2811, n2812, n2813, n2814, n2815, n2816,
    n2817, n2818, n2819, n2820, n2821, n2822,
    n2823, n2824, n2825, n2826, n2827, n2828,
    n2829, n2830, n2831, n2832, n2833, n2834,
    n2835, n2836, n2837, n2838, n2839, n2840,
    n2841, n2842, n2843, n2844, n2845, n2846,
    n2847, n2848, n2849, n2850, n2851, n2852,
    n2853, n2854, n2855, n2856, n2857, n2858,
    n2859, n2860, n2861, n2862, n2863, n2864,
    n2865, n2866, n2867, n2868, n2869, n2870,
    n2871, n2872, n2873, n2874, n2875, n2876,
    n2877, n2878, n2879, n2880, n2881, n2882,
    n2883, n2884, n2885, n2886, n2887, n2888,
    n2889, n2890, n2891, n2892, n2893, n2894,
    n2895, n2896, n2897, n2898, n2899, n2900,
    n2901, n2902, n2903, n2904, n2905, n2906,
    n2907, n2908, n2909, n2910, n2911, n2912,
    n2913, n2914, n2915, n2916, n2917, n2918,
    n2919, n2920, n2921, n2922, n2923, n2924,
    n2925, n2926, n2927, n2928, n2929, n2930,
    n2931, n2932, n2933, n2934, n2935, n2936,
    n2937, n2938, n2939, n2940, n2941, n2942,
    n2943, n2944, n2945, n2946, n2947, n2948,
    n2949, n2950, n2951, n2952, n2953, n2954,
    n2955, n2956, n2957, n2958, n2959, n2960,
    n2961, n2962, n2963, n2964, n2965, n2966,
    n2967, n2968, n2969, n2970, n2971, n2972,
    n2973, n2974, n2975, n2976, n2977, n2978,
    n2979, n2980, n2981, n2982, n2983, n2984,
    n2985, n2986, n2987, n2988, n2989, n2990,
    n2991, n2992, n2993, n2994, n2995, n2996,
    n2997, n2998, n2999, n3000, n3001, n3002,
    n3003, n3004, n3005, n3006, n3007, n3008,
    n3009, n3010, n3011, n3012, n3013, n3014,
    n3015, n3016, n3017, n3018, n3019, n3020,
    n3021, n3022, n3023, n3024, n3025, n3026,
    n3027, n3028, n3029, n3030, n3031, n3032,
    n3033, n3034, n3035, n3036, n3037, n3038,
    n3039, n3040, n3041, n3042, n3043, n3044,
    n3045, n3046, n3047, n3048, n3049, n3050,
    n3051, n3052, n3053, n3054, n3055, n3056,
    n3057, n3058, n3059, n3060, n3061, n3062,
    n3063, n3064, n3065, n3066, n3067, n3068,
    n3069, n3070, n3071, n3072, n3073, n3074,
    n3075, n3076, n3077, n3078, n3079, n3080,
    n3081, n3082, n3083, n3084, n3085, n3086,
    n3087, n3088, n3089, n3090, n3091, n3092,
    n3093, n3094, n3095, n3096, n3097, n3098,
    n3099, n3100, n3101, n3102, n3103, n3104,
    n3105, n3106, n3107, n3108, n3109, n3110,
    n3111, n3112, n3113, n3114, n3115, n3116,
    n3117, n3118, n3119, n3120, n3121, n3122,
    n3123, n3124, n3125, n3126, n3127, n3128,
    n3129, n3130, n3131, n3132, n3133, n3134,
    n3135, n3136, n3137, n3138, n3139, n3140,
    n3141, n3142, n3143, n3144, n3145, n3146,
    n3147, n3148, n3149, n3150, n3151, n3152,
    n3153, n3154, n3155, n3156, n3157, n3158,
    n3159, n3160, n3161, n3162, n3163, n3164,
    n3165, n3166, n3167, n3168, n3169, n3170,
    n3171, n3172, n3173, n3174, n3175, n3176,
    n3177, n3178, n3179, n3180, n3181, n3182,
    n3183, n3184, n3185, n3186, n3187, n3188,
    n3189, n3190, n3191, n3192, n3193, n3194,
    n3195, n3196, n3197, n3198, n3199, n3200,
    n3201, n3202, n3203, n3204, n3205, n3206,
    n3207, n3208, n3209, n3210, n3211, n3212,
    n3213, n3214, n3215, n3216, n3217, n3218,
    n3219, n3220, n3221, n3222, n3223, n3224,
    n3225, n3226, n3227, n3228, n3229, n3230,
    n3231, n3232, n3233, n3234, n3235, n3236,
    n3237, n3238, n3239, n3240, n3241, n3242,
    n3243, n3244, n3245, n3246, n3247, n3248,
    n3249, n3250, n3251, n3252, n3253, n3254,
    n3255, n3256, n3257, n3258, n3259, n3260,
    n3261, n3262, n3263, n3264, n3265, n3266,
    n3267, n3268, n3269, n3270, n3271, n3272,
    n3273, n3274, n3275, n3276, n3277, n3278,
    n3279, n3280, n3281, n3282, n3283, n3284,
    n3285, n3286, n3287, n3288, n3289, n3290,
    n3291, n3292, n3293, n3294, n3295, n3296,
    n3297, n3298, n3299, n3300, n3301, n3302,
    n3303, n3304, n3305, n3306, n3307, n3308,
    n3309, n3310, n3311, n3312, n3313, n3314,
    n3315, n3316, n3317, n3318, n3319, n3320,
    n3321, n3322, n3323, n3324, n3325, n3326,
    n3327, n3328, n3329, n3330, n3331, n3332,
    n3333, n3334, n3335, n3336, n3337, n3338,
    n3339, n3340, n3341, n3342, n3343, n3344,
    n3345, n3346, n3347, n3348, n3349, n3350,
    n3351, n3352, n3353, n3354, n3355, n3356,
    n3357, n3358, n3359, n3360, n3361, n3362,
    n3363, n3364, n3365, n3366, n3367, n3368,
    n3369, n3370, n3371, n3372, n3373, n3374,
    n3375, n3376, n3377, n3378, n3379, n3380,
    n3381, n3382, n3383, n3384, n3385, n3386,
    n3387, n3388, n3389, n3390, n3391, n3392,
    n3393, n3394, n3395, n3396, n3397, n3398,
    n3399, n3400, n3401, n3402, n3403, n3404,
    n3405, n3406, n3407, n3408, n3409, n3410,
    n3411, n3412, n3413, n3414, n3415, n3416,
    n3417, n3418, n3419, n3420, n3421, n3422,
    n3423, n3424, n3425, n3426, n3427, n3428,
    n3429, n3430, n3431, n3432, n3433, n3434,
    n3435, n3436, n3437, n3438, n3439, n3440,
    n3441, n3442, n3443, n3444, n3445, n3446,
    n3447, n3448, n3449, n3450, n3451, n3452,
    n3453, n3454, n3455, n3456, n3457, n3458,
    n3459, n3460, n3461, n3462, n3463, n3464,
    n3465, n3466, n3467, n3468, n3469, n3470,
    n3471, n3472, n3473, n3474, n3475, n3476,
    n3477, n3478, n3479, n3480, n3481, n3482,
    n3483, n3484, n3485, n3486, n3487, n3488,
    n3489, n3490, n3491, n3492, n3493, n3494,
    n3495, n3496, n3497, n3498, n3499, n3500,
    n3501, n3502, n3503, n3504, n3505, n3506,
    n3507, n3508, n3509, n3510, n3511, n3512,
    n3513, n3514, n3515, n3516, n3517, n3518,
    n3519, n3520, n3521, n3522, n3523, n3524,
    n3525, n3526, n3527, n3528, n3529, n3530,
    n3531, n3532, n3533, n3534, n3535, n3536,
    n3537, n3538, n3539, n3540, n3541, n3542,
    n3543, n3544, n3545, n3546, n3547, n3548,
    n3549, n3550, n3551, n3552, n3553, n3554,
    n3555, n3556, n3557, n3558, n3559, n3560,
    n3561, n3562, n3563, n3564, n3565, n3566,
    n3567, n3568, n3569, n3570, n3571, n3572,
    n3573, n3574, n3575, n3576, n3577, n3578,
    n3579, n3580, n3581, n3582, n3583, n3584,
    n3585, n3586, n3587, n3588, n3589, n3590,
    n3591, n3592, n3593, n3594, n3595, n3596,
    n3597, n3598, n3599, n3600, n3601, n3602,
    n3603, n3604, n3605, n3606, n3607, n3608,
    n3609, n3610, n3611, n3612, n3613, n3614,
    n3615, n3616, n3617, n3618, n3619, n3620,
    n3621, n3622, n3623, n3624, n3625, n3626,
    n3627, n3628, n3629, n3630, n3631, n3632,
    n3633, n3634, n3635, n3636, n3637, n3638,
    n3639, n3640, n3641, n3642, n3643, n3644,
    n3645, n3646, n3647, n3648, n3649, n3650,
    n3651, n3652, n3653, n3654, n3655, n3656,
    n3657, n3658, n3659, n3660, n3661, n3662,
    n3663, n3664, n3665, n3666, n3667, n3668,
    n3669, n3670, n3671, n3672, n3673, n3674,
    n3675, n3676, n3677, n3678, n3679, n3680,
    n3681, n3682, n3683, n3684, n3685, n3686,
    n3687, n3688, n3689, n3690, n3691, n3692,
    n3693, n3694, n3695, n3696, n3697, n3698,
    n3699, n3700, n3701, n3702, n3703, n3704,
    n3705, n3706, n3707, n3708, n3709, n3710,
    n3711, n3712, n3713, n3714, n3715, n3716,
    n3717, n3718, n3719, n3720, n3721, n3722,
    n3723, n3724, n3725, n3726, n3727, n3728,
    n3729, n3730, n3731, n3732, n3733, n3734,
    n3735, n3736, n3737, n3738, n3739, n3740,
    n3741, n3742, n3743, n3744, n3745, n3746,
    n3747, n3748, n3749, n3750, n3751, n3752,
    n3753, n3754, n3755, n3756, n3757, n3758,
    n3759, n3760, n3761, n3762, n3763, n3764,
    n3765, n3766, n3767, n3768, n3769, n3770,
    n3771, n3772, n3773, n3774, n3775, n3776,
    n3777, n3778, n3779, n3780, n3781, n3782,
    n3783, n3784, n3785, n3786, n3787, n3788,
    n3789, n3790, n3791, n3792, n3793, n3794,
    n3795, n3796, n3797, n3798, n3799, n3800,
    n3801, n3802, n3803, n3804, n3805, n3806,
    n3807, n3808, n3809, n3810, n3811, n3812,
    n3813, n3814, n3815, n3816, n3817, n3818,
    n3819, n3820, n3821, n3822, n3823, n3824,
    n3825, n3826, n3827, n3828, n3829, n3830,
    n3831, n3832, n3833, n3834, n3835, n3836,
    n3837, n3838, n3839, n3840, n3841, n3842,
    n3843, n3844, n3845, n3846, n3847, n3848,
    n3849, n3850, n3851, n3852, n3853, n3854,
    n3855, n3856, n3857, n3858, n3859, n3860,
    n3861, n3862, n3863, n3864, n3865, n3866,
    n3867, n3868, n3869, n3870, n3871, n3872,
    n3873, n3874, n3875, n3876, n3877, n3878,
    n3879, n3880, n3881, n3882, n3883, n3884,
    n3885, n3886, n3887, n3888, n3889, n3890,
    n3891, n3892, n3893, n3894, n3895, n3896,
    n3897, n3898, n3899, n3900, n3901, n3902,
    n3903, n3904, n3905, n3906, n3907, n3908,
    n3909, n3910, n3911, n3912, n3913, n3914,
    n3915, n3916, n3917, n3918, n3919, n3920,
    n3921, n3922, n3923, n3924, n3925, n3926,
    n3927, n3928, n3929, n3930, n3931, n3932,
    n3933, n3934, n3935, n3936, n3937, n3938,
    n3939, n3940, n3941, n3942, n3943, n3944,
    n3945, n3946, n3947, n3948, n3949, n3950,
    n3951, n3952, n3953, n3954, n3955, n3956,
    n3957, n3958, n3959, n3960, n3961, n3962,
    n3963, n3964, n3965, n3966, n3967, n3968,
    n3969, n3970, n3971, n3972, n3973, n3974,
    n3975, n3976, n3977, n3978, n3979, n3980,
    n3981, n3982, n3983, n3984, n3985, n3986,
    n3987, n3988, n3989, n3990, n3991, n3992,
    n3993, n3994, n3995, n3996, n3997, n3998,
    n3999, n4000, n4001, n4002, n4003, n4004,
    n4005, n4006, n4007, n4008, n4009, n4010,
    n4011, n4012, n4013, n4014, n4015, n4016,
    n4017, n4018, n4019, n4020, n4021, n4022,
    n4023, n4024, n4025, n4026, n4027, n4028,
    n4029, n4030, n4031, n4032, n4033, n4034,
    n4035, n4036, n4037, n4038, n4039, n4040,
    n4041, n4042, n4043, n4044, n4045, n4046,
    n4047, n4048, n4049, n4050, n4051, n4052,
    n4053, n4054, n4055, n4056, n4057, n4058,
    n4059, n4060, n4061, n4062, n4063, n4064,
    n4065, n4066, n4067, n4068, n4069, n4070,
    n4071, n4072, n4073, n4074, n4075, n4076,
    n4077, n4078, n4079, n4080, n4081, n4082,
    n4083, n4084, n4085, n4086, n4087, n4088,
    n4089, n4090, n4091, n4092, n4093, n4094,
    n4095, n4096, n4097, n4098, n4099, n4100,
    n4101, n4102, n4103, n4104, n4105, n4106,
    n4107, n4108, n4109, n4110, n4111, n4112,
    n4113, n4114, n4115, n4116, n4117, n4118,
    n4119, n4120, n4121, n4122, n4123, n4124,
    n4125, n4126, n4127, n4128, n4129, n4130,
    n4131, n4132, n4133, n4134, n4135, n4136,
    n4137, n4138, n4139, n4140, n4141, n4142,
    n4143, n4144, n4145, n4146, n4147, n4148,
    n4149, n4150, n4151, n4152, n4153, n4154,
    n4155, n4156, n4157, n4158, n4159, n4160,
    n4161, n4162, n4163, n4164, n4165, n4166,
    n4167, n4168, n4169, n4170, n4171, n4172,
    n4173, n4174, n4175, n4176, n4177, n4178,
    n4179, n4180, n4181, n4182, n4183, n4184,
    n4185, n4186, n4187, n4188, n4189, n4190,
    n4191, n4192, n4193, n4194, n4195, n4196,
    n4197, n4198, n4199, n4200, n4201, n4202,
    n4203, n4204, n4205, n4206, n4207, n4208,
    n4209, n4210, n4211, n4212, n4213, n4214,
    n4215, n4216, n4217, n4218, n4219, n4220,
    n4221, n4222, n4223, n4224, n4225, n4226,
    n4227, n4228, n4229, n4230, n4231, n4232,
    n4233, n4234, n4235, n4236, n4237, n4238,
    n4239, n4240, n4241, n4242, n4243, n4244,
    n4245, n4246, n4247, n4248, n4249, n4250,
    n4251, n4252, n4253, n4254, n4255, n4256,
    n4257, n4258, n4259, n4260, n4261, n4262,
    n4263, n4264, n4265, n4266, n4267, n4268,
    n4269, n4270, n4271, n4272, n4273, n4274,
    n4275, n4276, n4277, n4278, n4279, n4280,
    n4281, n4282, n4283, n4284, n4285, n4286,
    n4287, n4288, n4289, n4290, n4291, n4292,
    n4293, n4294, n4295, n4296, n4297, n4298,
    n4299, n4300, n4301, n4302, n4303, n4304,
    n4305, n4306, n4307, n4308, n4309, n4310,
    n4311, n4312, n4313, n4314, n4315, n4316,
    n4317, n4318, n4319, n4320, n4321, n4322,
    n4323, n4324, n4325, n4326, n4327, n4328,
    n4329, n4330, n4331, n4332, n4333, n4334,
    n4335, n4336, n4337, n4338, n4339, n4340,
    n4341, n4342, n4343, n4344, n4345, n4346,
    n4347, n4348, n4349, n4350, n4351, n4352,
    n4353, n4354, n4355, n4356, n4357, n4358,
    n4359, n4360, n4361, n4362, n4363, n4364,
    n4365, n4366, n4367, n4368, n4369, n4370,
    n4371, n4372, n4373, n4374, n4375, n4376,
    n4377, n4378, n4379, n4380, n4381, n4382,
    n4383, n4384, n4385, n4386, n4387, n4388,
    n4389, n4390, n4391, n4392, n4393, n4394,
    n4395, n4396, n4397, n4398, n4399, n4400,
    n4401, n4402, n4403, n4404, n4405, n4406,
    n4407, n4408, n4409, n4410, n4411, n4412,
    n4413, n4414, n4415, n4416, n4417, n4418,
    n4419, n4420, n4421, n4422, n4423, n4424,
    n4425, n4426, n4427, n4428, n4429, n4430,
    n4431, n4432, n4433, n4434, n4435, n4436,
    n4437, n4438, n4439, n4440, n4441, n4442,
    n4443, n4444, n4445, n4446, n4447, n4448,
    n4449, n4450, n4451, n4452, n4453, n4454,
    n4455, n4456, n4457, n4458, n4459, n4460,
    n4461, n4462, n4463, n4464, n4465, n4466,
    n4467, n4468, n4469, n4470, n4471, n4472,
    n4473, n4474, n4475, n4476, n4477, n4478,
    n4479, n4480, n4481, n4482, n4483, n4484,
    n4485, n4486, n4487, n4488, n4489, n4490,
    n4491, n4492, n4493, n4494, n4495, n4496,
    n4497, n4498, n4499, n4500, n4501, n4502,
    n4503, n4504, n4505, n4506, n4507, n4508,
    n4509, n4510, n4511, n4512, n4513, n4514,
    n4515, n4516, n4517, n4518, n4519, n4520,
    n4521, n4522, n4523, n4524, n4525, n4526,
    n4527, n4528, n4529, n4530, n4531, n4532,
    n4533, n4534, n4535, n4536, n4537, n4538,
    n4539, n4540, n4541, n4542, n4543, n4544,
    n4545, n4546, n4547, n4548, n4549, n4550,
    n4551, n4552, n4553, n4554, n4555, n4556,
    n4557, n4558, n4559, n4560, n4561, n4562,
    n4563, n4564, n4565, n4566, n4567, n4568,
    n4569, n4570, n4571, n4572, n4573, n4574,
    n4575, n4576, n4577, n4578, n4579, n4580,
    n4581, n4582, n4583, n4584, n4585, n4586,
    n4587, n4588, n4589, n4590, n4591, n4592,
    n4593, n4594, n4595, n4596, n4597, n4598,
    n4599, n4600, n4601, n4602, n4603, n4604,
    n4605, n4606, n4607, n4608, n4609, n4610,
    n4611, n4612, n4613, n4614, n4615, n4616,
    n4617, n4618, n4619, n4620, n4621, n4622,
    n4623, n4624, n4625, n4626, n4627, n4628,
    n4629, n4630, n4631, n4632, n4633, n4634,
    n4635, n4636, n4637, n4638, n4639, n4640,
    n4641, n4642, n4643, n4644, n4645, n4646,
    n4647, n4648, n4649, n4650, n4651, n4652,
    n4653, n4654, n4655, n4656, n4657, n4658,
    n4659, n4660, n4661, n4662, n4663, n4664,
    n4665, n4666, n4667, n4668, n4669, n4670,
    n4671, n4672, n4673, n4674, n4675, n4676,
    n4677, n4678, n4679, n4680, n4681, n4682,
    n4683, n4684, n4685, n4686, n4687, n4688,
    n4689, n4690, n4691, n4692, n4693, n4694,
    n4695, n4696, n4697, n4698, n4699, n4700,
    n4701, n4702, n4703, n4704, n4705, n4706,
    n4707, n4708, n4709, n4710, n4711, n4712,
    n4713, n4714, n4715, n4716, n4717, n4718,
    n4719, n4720, n4721, n4722, n4723, n4724,
    n4725, n4726, n4727, n4728, n4729, n4730,
    n4731, n4732, n4733, n4734, n4735, n4736,
    n4737, n4738, n4739, n4740, n4741, n4742,
    n4743, n4744, n4745, n4746, n4747, n4748,
    n4749, n4750, n4751, n4752, n4753, n4754,
    n4755, n4756, n4757, n4758, n4759, n4760,
    n4761, n4762, n4763, n4764, n4765, n4766,
    n4767, n4768, n4769, n4770, n4771, n4772,
    n4773, n4774, n4775, n4776, n4777, n4778,
    n4779, n4780, n4781, n4782, n4783, n4784,
    n4785, n4786, n4787, n4788, n4789, n4790,
    n4791, n4792, n4793, n4794, n4795, n4796,
    n4797, n4798, n4799, n4800, n4801, n4802,
    n4803, n4804, n4805, n4806, n4807, n4808,
    n4809, n4810, n4811, n4812, n4813, n4814,
    n4815, n4816, n4817, n4818, n4819, n4820,
    n4821, n4822, n4823, n4824, n4825, n4826,
    n4827, n4828, n4829, n4830, n4831, n4832,
    n4833, n4834, n4835, n4836, n4837, n4838,
    n4839, n4840, n4841, n4842, n4843, n4844,
    n4845, n4846, n4847, n4848, n4849, n4850,
    n4851, n4852, n4853, n4854, n4855, n4856,
    n4857, n4858, n4859, n4860, n4861, n4862,
    n4863, n4864, n4865, n4866, n4867, n4868,
    n4869, n4870, n4871, n4872, n4873, n4874,
    n4875, n4876, n4877, n4878, n4879, n4880,
    n4881, n4882, n4883, n4884, n4885, n4886,
    n4887, n4888, n4889, n4890, n4891, n4892,
    n4893, n4894, n4895, n4896, n4897, n4898,
    n4899, n4900, n4901, n4902, n4903, n4904,
    n4905, n4906, n4907, n4908, n4909, n4910,
    n4911, n4912, n4913, n4914, n4915, n4916,
    n4917, n4918, n4919, n4920, n4921, n4922,
    n4923, n4924, n4925, n4926, n4927, n4928,
    n4929, n4930, n4931, n4932, n4933, n4934,
    n4935, n4936, n4937, n4938, n4939, n4940,
    n4941, n4942, n4943, n4944, n4945, n4946,
    n4947, n4948, n4949, n4950, n4951, n4952,
    n4953, n4954, n4955, n4956, n4957, n4958,
    n4959, n4960, n4961, n4962, n4963, n4964,
    n4965, n4966, n4967, n4968, n4969, n4970,
    n4971, n4972, n4973, n4974, n4975, n4976,
    n4977, n4978, n4979, n4980, n4981, n4982,
    n4983, n4984, n4985, n4986, n4987, n4988,
    n4989, n4990, n4991, n4992, n4993, n4994,
    n4995, n4996, n4997, n4998, n4999, n5000,
    n5001, n5002, n5003, n5004, n5005, n5006,
    n5007, n5008, n5009, n5010, n5011, n5012,
    n5013, n5014, n5015, n5016, n5017, n5018,
    n5019, n5020, n5021, n5022, n5023, n5024,
    n5025, n5026, n5027, n5028, n5029, n5030,
    n5031, n5032, n5033, n5034, n5035, n5036,
    n5037, n5038, n5039, n5040, n5041, n5042,
    n5043, n5044, n5045, n5046, n5047, n5048,
    n5049, n5050, n5051, n5052, n5053, n5054,
    n5055, n5056, n5057, n5058, n5059, n5060,
    n5061, n5062, n5063, n5064, n5065, n5066,
    n5067, n5068, n5069, n5070, n5071, n5072,
    n5073, n5074, n5075, n5076, n5077, n5078,
    n5079, n5080, n5081, n5082, n5083, n5084,
    n5085, n5086, n5087, n5088, n5089, n5090,
    n5091, n5092, n5093, n5094, n5095, n5096,
    n5097, n5098, n5099, n5100, n5101, n5102,
    n5103, n5104, n5105, n5106, n5107, n5108,
    n5109, n5110, n5111, n5112, n5113, n5114,
    n5115, n5116, n5117, n5118, n5119, n5120,
    n5121, n5122, n5123, n5124, n5125, n5126,
    n5127, n5128, n5129, n5130, n5131, n5132,
    n5133, n5134, n5135, n5136, n5137, n5138,
    n5139, n5140, n5141, n5142, n5143, n5144,
    n5145, n5146, n5147, n5148, n5149, n5150,
    n5151, n5152, n5153, n5154, n5155, n5156,
    n5157, n5158, n5159, n5160, n5161, n5162,
    n5163, n5164, n5165, n5166, n5167, n5168,
    n5169, n5170, n5171, n5172, n5173, n5174,
    n5175, n5176, n5177, n5178, n5179, n5180,
    n5181, n5182, n5183, n5184, n5185, n5186,
    n5187, n5188, n5189, n5190, n5191, n5192,
    n5193, n5194, n5195, n5196, n5197, n5198,
    n5199, n5200, n5201, n5202, n5203, n5204,
    n5205, n5206, n5207, n5208, n5209, n5210,
    n5211, n5212, n5213, n5214, n5215, n5216,
    n5217, n5218, n5219, n5220, n5221, n5222,
    n5223, n5224, n5225, n5226, n5227, n5228,
    n5229, n5230, n5231, n5232, n5233, n5234,
    n5235, n5236, n5237, n5238, n5239, n5240,
    n5241, n5242, n5243, n5244, n5245, n5246,
    n5247, n5248, n5249, n5250, n5251, n5252,
    n5253, n5254, n5255, n5256, n5257, n5258,
    n5259, n5260, n5261, n5262, n5263, n5264,
    n5265, n5266, n5267, n5268, n5269, n5270,
    n5271, n5272, n5273, n5274, n5275, n5276,
    n5277, n5278, n5279, n5280, n5281, n5282,
    n5283, n5284, n5285, n5286, n5287, n5288,
    n5289, n5290, n5291, n5292, n5293, n5294,
    n5295, n5296, n5297, n5298, n5299, n5300,
    n5301, n5302, n5303, n5304, n5305, n5306,
    n5307, n5308, n5309, n5310, n5311, n5312,
    n5313, n5314, n5315, n5316, n5317, n5318,
    n5319, n5320, n5321, n5322, n5323, n5324,
    n5325, n5326, n5327, n5328, n5329, n5330,
    n5331, n5332, n5333, n5334, n5335, n5336,
    n5337, n5338, n5339, n5340, n5341, n5342,
    n5343, n5344, n5345, n5346, n5347, n5348,
    n5349, n5350, n5351, n5352, n5353, n5354,
    n5355, n5356, n5357, n5358, n5359, n5360,
    n5361, n5362, n5363, n5364, n5365, n5366,
    n5367, n5368, n5369, n5370, n5371, n5372,
    n5373, n5374, n5375, n5376, n5377, n5378,
    n5379, n5380, n5381, n5382, n5383, n5384,
    n5385, n5386, n5387, n5388, n5389, n5390,
    n5391, n5392, n5393, n5394, n5395, n5396,
    n5397, n5398, n5399, n5400, n5401, n5402,
    n5403, n5404, n5405, n5406, n5407, n5408,
    n5409, n5410, n5411, n5412, n5413, n5414,
    n5415, n5416, n5417, n5418, n5419, n5420,
    n5421, n5422, n5423, n5424, n5425, n5426,
    n5427, n5428, n5429, n5430, n5431, n5432,
    n5433, n5434, n5435, n5436, n5437, n5438,
    n5439, n5440, n5441, n5442, n5443, n5444,
    n5445, n5446, n5447, n5448, n5449, n5450,
    n5451, n5452, n5453, n5454, n5455, n5456,
    n5457, n5458, n5459, n5460, n5461, n5462,
    n5463, n5464, n5465, n5466, n5467, n5468,
    n5469, n5470, n5471, n5472, n5473, n5474,
    n5475, n5476, n5477, n5478, n5479, n5480,
    n5481, n5482, n5483, n5484, n5485, n5486,
    n5487, n5488, n5489, n5490, n5491, n5492,
    n5493, n5494, n5495, n5496, n5497, n5498,
    n5499, n5500, n5501, n5502, n5503, n5504,
    n5505, n5506, n5507, n5508, n5509, n5510,
    n5511, n5512, n5513, n5514, n5515, n5516,
    n5517, n5518, n5519, n5520, n5521, n5522,
    n5523, n5524, n5525, n5526, n5527, n5528,
    n5529, n5530, n5531, n5532, n5533, n5534,
    n5535, n5536, n5537, n5538, n5539, n5540,
    n5541, n5542, n5543, n5544, n5545, n5546,
    n5547, n5548, n5549, n5550, n5551, n5552,
    n5553, n5554, n5555, n5556, n5557, n5558,
    n5559, n5560, n5561, n5562, n5563, n5564,
    n5565, n5566, n5567, n5568, n5569, n5570,
    n5571, n5572, n5573, n5574, n5575, n5576,
    n5577, n5578, n5579, n5580, n5581, n5582,
    n5583, n5584, n5585, n5586, n5587, n5588,
    n5589, n5590, n5591, n5592, n5593, n5594,
    n5595, n5596, n5597, n5598, n5599, n5600,
    n5601, n5602, n5603, n5604, n5605, n5606,
    n5607, n5608, n5609, n5610, n5611, n5612,
    n5613, n5614, n5615, n5616, n5617, n5618,
    n5619, n5620, n5621, n5622, n5623, n5624,
    n5625, n5626, n5627, n5628, n5629, n5630,
    n5631, n5632, n5633, n5634, n5635, n5636,
    n5637, n5638, n5639, n5640, n5641, n5642,
    n5643, n5644, n5645, n5646, n5647, n5648,
    n5649, n5650, n5651, n5652, n5653, n5654,
    n5655, n5656, n5657, n5658, n5659, n5660,
    n5661, n5662, n5663, n5664, n5665, n5666,
    n5667, n5668, n5669, n5670, n5671, n5672,
    n5673, n5674, n5675, n5676, n5677, n5678,
    n5679, n5680, n5681, n5682, n5683, n5684,
    n5685, n5686, n5687, n5688, n5689, n5690,
    n5691, n5692, n5693, n5694, n5695, n5696,
    n5697, n5698, n5699, n5700, n5701, n5702,
    n5703, n5704, n5705, n5706, n5707, n5708,
    n5709, n5710, n5711, n5712, n5713, n5714,
    n5715, n5716, n5717, n5718, n5719, n5720,
    n5721, n5722, n5723, n5724, n5725, n5726,
    n5727, n5728, n5729, n5730, n5731, n5732,
    n5733, n5734, n5735, n5736, n5737, n5738,
    n5739, n5740, n5741, n5742, n5743, n5744,
    n5745, n5746, n5747, n5748, n5749, n5750,
    n5751, n5752, n5753, n5754, n5755, n5756,
    n5757, n5758, n5759, n5760, n5761, n5762,
    n5763, n5764, n5765, n5766, n5767, n5768,
    n5769, n5770, n5771, n5772, n5773, n5774,
    n5775, n5776, n5777, n5778, n5779, n5780,
    n5781, n5782, n5783, n5784, n5785, n5786,
    n5787, n5788, n5789, n5790, n5791, n5792,
    n5793, n5794, n5795, n5796, n5797, n5798,
    n5799, n5800, n5801, n5802, n5803, n5804,
    n5805, n5806, n5807, n5808, n5809, n5810,
    n5811, n5812, n5813, n5814, n5815, n5816,
    n5817, n5818, n5819, n5820, n5821, n5822,
    n5823, n5824, n5825, n5826, n5827, n5828,
    n5829, n5830, n5831, n5832, n5833, n5834,
    n5835, n5836, n5837, n5838, n5839, n5840,
    n5841, n5842, n5843, n5844, n5845, n5846,
    n5847, n5848, n5849, n5850, n5851, n5852,
    n5853, n5854, n5855, n5856, n5857, n5858,
    n5859, n5860, n5861, n5862, n5863, n5864,
    n5865, n5866, n5867, n5868, n5869, n5870,
    n5871, n5872, n5873, n5874, n5875, n5876,
    n5877, n5878, n5879, n5880, n5881, n5882,
    n5883, n5884, n5885, n5886, n5887, n5888,
    n5889, n5890, n5891, n5892, n5893, n5894,
    n5895, n5896, n5897, n5898, n5899, n5900,
    n5901, n5902, n5903, n5904, n5905, n5906,
    n5907, n5908, n5909, n5910, n5911, n5912,
    n5913, n5914, n5915, n5916, n5917, n5918,
    n5919, n5920, n5921, n5922, n5923, n5924,
    n5925, n5926, n5927, n5928, n5929, n5930,
    n5931, n5932, n5933, n5934, n5935, n5936,
    n5937, n5938, n5939, n5940, n5941, n5942,
    n5943, n5944, n5945, n5946, n5947, n5948,
    n5949, n5950, n5951, n5952, n5953, n5954,
    n5955, n5956, n5957, n5958, n5959, n5960,
    n5961, n5962, n5963, n5964, n5965, n5966,
    n5967, n5968, n5969, n5970, n5971, n5972,
    n5973, n5974, n5975, n5976, n5977, n5978,
    n5979, n5980, n5981, n5982, n5983, n5984,
    n5985, n5986, n5987, n5988, n5989, n5990,
    n5991, n5992, n5993, n5994, n5995, n5996,
    n5997, n5998, n5999, n6000, n6001, n6002,
    n6003, n6004, n6005, n6006, n6007, n6008,
    n6009, n6010, n6011, n6012, n6013, n6014,
    n6015, n6016, n6017, n6018, n6019, n6020,
    n6021, n6022, n6023, n6024, n6025, n6026,
    n6027, n6028, n6029, n6030, n6031, n6032,
    n6033, n6034, n6035, n6036, n6037, n6038,
    n6039, n6040, n6041, n6042, n6043, n6044,
    n6045, n6046, n6047, n6048, n6049, n6050,
    n6051, n6052, n6053, n6054, n6055, n6056,
    n6057, n6058, n6059, n6060, n6061, n6062,
    n6063, n6064, n6065, n6066, n6067, n6068,
    n6069, n6070, n6071, n6072, n6073, n6074,
    n6075, n6076, n6077, n6078, n6079, n6080,
    n6081, n6082, n6083, n6084, n6085, n6086,
    n6087, n6088, n6089, n6090, n6091, n6092,
    n6093, n6094, n6095, n6096, n6097, n6098,
    n6099, n6100, n6101, n6102, n6103, n6104,
    n6105, n6106, n6107, n6108, n6109, n6110,
    n6111, n6112, n6113, n6114, n6115, n6116,
    n6117, n6118, n6119, n6120, n6121, n6122,
    n6123, n6124, n6125, n6126, n6127, n6128,
    n6129, n6130, n6131, n6132, n6133, n6134,
    n6135, n6136, n6137, n6138, n6139, n6140,
    n6141, n6142, n6143, n6144, n6145, n6146,
    n6147, n6148, n6149, n6150, n6151, n6152,
    n6153, n6154, n6155, n6156, n6157, n6158,
    n6159, n6160, n6161, n6162, n6163, n6164,
    n6165, n6166, n6167, n6168, n6169, n6170,
    n6171, n6172, n6173, n6174, n6175, n6176,
    n6177, n6178, n6179, n6180, n6181, n6182,
    n6183, n6184, n6185, n6186, n6187, n6188,
    n6189, n6190, n6191, n6192, n6193, n6194,
    n6195, n6196, n6197, n6198, n6199, n6200,
    n6201, n6202, n6203, n6204, n6205, n6206,
    n6207, n6208, n6209, n6210, n6211, n6212,
    n6213, n6214, n6215, n6216, n6217, n6218,
    n6219, n6220, n6221, n6222, n6223, n6224,
    n6225, n6226, n6227, n6228, n6229, n6230,
    n6231, n6232, n6233, n6234, n6235, n6236,
    n6237, n6238, n6239, n6240, n6241, n6242,
    n6243, n6244, n6245, n6246, n6247, n6248,
    n6249, n6250, n6251, n6252, n6253, n6254,
    n6255, n6256, n6257, n6258, n6259, n6260,
    n6261, n6262, n6263, n6264, n6265, n6266,
    n6267, n6268, n6269, n6270, n6271, n6272,
    n6273, n6274, n6275, n6276, n6277, n6278,
    n6279, n6280, n6281, n6282, n6283, n6284,
    n6285, n6286, n6287, n6288, n6289, n6290,
    n6291, n6292, n6293, n6294, n6295, n6296,
    n6297, n6298, n6299, n6300, n6301, n6302,
    n6303, n6304, n6305, n6306, n6307, n6308,
    n6309, n6310, n6311, n6312, n6313, n6314,
    n6315, n6316, n6317, n6318, n6319, n6320,
    n6321, n6322, n6323, n6324, n6325, n6326,
    n6327, n6328, n6329, n6330, n6331, n6332,
    n6333, n6334, n6335, n6336, n6337, n6338,
    n6339, n6340, n6341, n6342, n6343, n6344,
    n6345, n6346, n6347, n6348, n6349, n6350,
    n6351, n6352, n6353, n6354, n6355, n6356,
    n6357, n6358, n6359, n6360, n6361, n6362,
    n6363, n6364, n6365, n6366, n6367, n6368,
    n6369, n6370, n6371, n6372, n6373, n6374,
    n6375, n6376, n6377, n6378, n6379, n6380,
    n6381, n6382, n6383, n6384, n6385, n6386,
    n6387, n6388, n6389, n6390, n6391, n6392,
    n6393, n6394, n6395, n6396, n6397, n6398,
    n6399, n6400, n6401, n6402, n6403, n6404,
    n6405, n6406, n6407, n6408, n6409, n6410,
    n6411, n6412, n6413, n6414, n6415, n6416,
    n6417, n6418, n6419, n6420, n6421, n6422,
    n6423, n6424, n6425, n6426, n6427, n6428,
    n6429, n6430, n6431, n6432, n6433, n6434,
    n6435, n6436, n6437, n6438, n6439, n6440,
    n6441, n6442, n6443, n6444, n6445, n6446,
    n6447, n6448, n6449, n6450, n6451, n6452,
    n6453, n6454, n6455, n6456, n6457, n6458,
    n6459, n6460, n6461, n6462, n6463, n6464,
    n6465, n6466, n6467, n6468, n6469, n6470,
    n6471, n6472, n6473, n6474, n6475, n6476,
    n6477, n6478, n6479, n6480, n6481, n6482,
    n6483, n6484, n6485, n6486, n6487, n6488,
    n6489, n6490, n6491, n6492, n6493, n6494,
    n6495, n6496, n6497, n6498, n6499, n6500,
    n6501, n6502, n6503, n6504, n6505, n6506,
    n6507, n6508, n6509, n6510, n6511, n6512,
    n6513, n6514, n6515, n6516, n6517, n6518,
    n6519, n6520, n6521, n6522, n6523, n6524,
    n6525, n6526, n6527, n6528, n6529, n6530,
    n6531, n6532, n6533, n6534, n6535, n6536,
    n6537, n6538, n6539, n6540, n6541, n6542,
    n6543, n6544, n6545, n6546, n6547, n6548,
    n6549, n6550, n6551, n6552, n6553, n6554,
    n6555, n6556, n6557, n6558, n6559, n6560,
    n6561, n6562, n6563, n6564, n6565, n6566,
    n6567, n6568, n6569, n6570, n6571, n6572,
    n6573, n6574, n6575, n6576, n6577, n6578,
    n6579, n6580, n6581, n6582, n6583, n6584,
    n6585, n6586, n6587, n6588, n6589, n6590,
    n6591, n6592, n6593, n6594, n6595, n6596,
    n6597, n6598, n6599, n6600, n6601, n6602,
    n6603, n6604, n6605, n6606, n6607, n6608,
    n6609, n6610, n6611, n6612, n6613, n6614,
    n6615, n6616, n6617, n6618, n6619, n6620,
    n6621, n6622, n6623, n6624, n6625, n6626,
    n6627, n6628, n6629, n6630, n6631, n6632,
    n6633, n6634, n6635, n6636, n6637, n6638,
    n6639, n6640, n6641, n6642, n6643, n6644,
    n6645, n6646, n6647, n6648, n6649, n6650,
    n6651, n6652, n6653, n6654, n6655, n6656,
    n6657, n6658, n6659, n6660, n6661, n6662,
    n6663, n6664, n6665, n6666, n6667, n6668,
    n6669, n6670, n6671, n6672, n6673, n6674,
    n6675, n6676, n6677, n6678, n6679, n6680,
    n6681, n6682, n6683, n6684, n6685, n6686,
    n6687, n6688, n6689, n6690, n6691, n6692,
    n6693, n6694, n6695, n6696, n6697, n6698,
    n6699, n6700, n6701, n6702, n6703, n6704,
    n6705, n6706, n6707, n6708, n6709, n6710,
    n6711, n6712, n6713, n6714, n6715, n6716,
    n6717, n6718, n6719, n6720, n6721, n6722,
    n6723, n6724, n6725, n6726, n6727, n6728,
    n6729, n6730, n6731, n6732, n6733, n6734,
    n6735, n6736, n6737, n6738, n6739, n6740,
    n6741, n6742, n6743, n6744, n6745, n6746,
    n6747, n6748, n6749, n6750, n6751, n6752,
    n6753, n6754, n6755, n6756, n6757, n6758,
    n6759, n6760, n6761, n6762, n6763, n6764,
    n6765, n6766, n6767, n6768, n6769, n6770,
    n6771, n6772, n6773, n6774, n6775, n6776,
    n6777, n6778, n6779, n6780, n6781, n6782,
    n6783, n6784, n6785, n6786, n6787, n6788,
    n6789, n6790, n6791, n6792, n6793, n6794,
    n6795, n6796, n6797, n6798, n6799, n6800,
    n6801, n6802, n6803, n6804, n6805, n6806,
    n6807, n6808, n6809, n6810, n6811, n6812,
    n6813, n6814, n6815, n6816, n6817, n6818,
    n6819, n6820, n6821, n6822, n6823, n6824,
    n6825, n6826, n6827, n6828, n6829, n6830,
    n6831, n6832, n6833, n6834, n6835, n6836,
    n6837, n6838, n6839, n6840, n6841, n6842,
    n6843, n6844, n6845, n6846, n6847, n6848,
    n6849, n6850, n6851, n6852, n6853, n6854,
    n6855, n6856, n6857, n6858, n6859, n6860,
    n6861, n6862, n6863, n6864, n6865, n6866,
    n6867, n6868, n6869, n6870, n6871, n6872,
    n6873, n6874, n6875, n6876, n6877, n6878,
    n6879, n6880, n6881, n6882, n6883, n6884,
    n6885, n6886, n6887, n6888, n6889, n6890,
    n6891, n6892, n6893, n6894, n6895, n6896,
    n6897, n6898, n6899, n6900, n6901, n6902,
    n6903, n6904, n6905, n6906, n6907, n6908,
    n6909, n6910, n6911, n6912, n6913, n6914,
    n6915, n6916, n6917, n6918, n6919, n6920,
    n6921, n6922, n6923, n6924, n6925, n6926,
    n6927, n6928, n6929, n6930, n6931, n6932,
    n6933, n6934, n6935, n6936, n6937, n6938,
    n6939, n6940, n6941, n6942, n6943, n6944,
    n6945, n6946, n6947, n6948, n6949, n6950,
    n6951, n6952, n6953, n6954, n6955, n6956,
    n6957, n6958, n6959, n6960, n6961, n6962,
    n6963, n6964, n6965, n6966, n6967, n6968,
    n6969, n6970, n6971, n6972, n6973, n6974,
    n6975, n6976, n6977, n6978, n6979, n6980,
    n6981, n6982, n6983, n6984, n6985, n6986,
    n6987, n6988, n6989, n6990, n6991, n6992,
    n6993, n6994, n6995, n6996, n6997, n6998,
    n6999, n7000, n7001, n7002, n7003, n7004,
    n7005, n7006, n7007, n7008, n7009, n7010,
    n7011, n7012, n7013, n7014, n7015, n7016,
    n7017, n7018, n7019, n7020, n7021, n7022,
    n7023, n7024, n7025, n7026, n7027, n7028,
    n7029, n7030, n7031, n7032, n7033, n7034,
    n7035, n7036, n7037, n7038, n7039, n7040,
    n7041, n7042, n7043, n7044, n7045, n7046,
    n7047, n7048, n7049, n7050, n7051, n7052,
    n7053, n7054, n7055, n7056, n7057, n7058,
    n7059, n7060, n7061, n7062, n7063, n7064,
    n7065, n7066, n7067, n7068, n7069, n7070,
    n7071, n7072, n7073, n7074, n7075, n7076,
    n7077, n7078, n7079, n7080, n7081, n7082,
    n7083, n7084, n7085, n7086, n7087, n7088,
    n7089, n7090, n7091, n7092, n7093, n7094,
    n7095, n7096, n7097, n7098, n7099, n7100,
    n7101, n7102, n7103, n7104, n7105, n7106,
    n7107, n7108, n7109, n7110, n7111, n7112,
    n7113, n7114, n7115, n7116, n7117, n7118,
    n7119, n7120, n7121, n7122, n7123, n7124,
    n7125, n7126, n7127, n7128, n7129, n7130,
    n7131, n7132, n7133, n7134, n7135, n7136,
    n7137, n7138, n7139, n7140, n7141, n7142,
    n7143, n7144, n7145, n7146, n7147, n7148,
    n7149, n7150, n7151, n7152, n7153, n7154,
    n7155, n7156, n7157, n7158, n7159, n7160,
    n7161, n7162, n7163, n7164, n7165, n7166,
    n7167, n7168, n7169, n7170, n7171, n7172,
    n7173, n7174, n7175, n7176, n7177, n7178,
    n7179, n7180, n7181, n7182, n7183, n7184,
    n7185, n7186, n7187, n7188, n7189, n7190,
    n7191, n7192, n7193, n7194, n7195, n7196,
    n7197, n7198, n7199, n7200, n7201, n7202,
    n7203, n7204, n7205, n7206, n7207, n7208,
    n7209, n7210, n7211, n7212, n7213, n7214,
    n7215, n7216, n7217, n7218, n7219, n7220,
    n7221, n7222, n7223, n7224, n7225, n7226,
    n7227, n7228, n7229, n7230, n7231, n7232,
    n7233, n7234, n7235, n7236, n7237, n7238,
    n7239, n7240, n7241, n7242, n7243, n7244,
    n7245, n7246, n7247, n7248, n7249, n7250,
    n7251, n7252, n7253, n7254, n7255, n7256,
    n7257, n7258, n7259, n7260, n7261, n7262,
    n7263, n7264, n7265, n7266, n7267, n7268,
    n7269, n7270, n7271, n7272, n7273, n7274,
    n7275, n7276, n7277, n7278, n7279, n7280,
    n7281, n7282, n7283, n7284, n7285, n7286,
    n7287, n7288, n7289, n7290, n7291, n7292,
    n7293, n7294, n7295, n7296, n7297, n7298,
    n7299, n7300, n7301, n7302, n7303, n7304,
    n7305, n7306, n7307, n7308, n7309, n7310,
    n7311, n7312, n7313, n7314, n7315, n7316,
    n7317, n7318, n7319, n7320, n7321, n7322,
    n7323, n7324, n7325, n7326, n7327, n7328,
    n7329, n7330, n7331, n7332, n7333, n7334,
    n7335, n7336, n7337, n7338, n7339, n7340,
    n7341, n7342, n7343, n7344, n7345, n7346,
    n7347, n7348, n7349, n7350, n7351, n7352,
    n7353, n7354, n7355, n7356, n7357, n7358,
    n7359, n7360, n7361, n7362, n7363, n7364,
    n7365, n7366, n7367, n7368, n7369, n7370,
    n7371, n7372, n7373, n7374, n7375, n7376,
    n7377, n7378, n7379, n7380, n7381, n7382,
    n7383, n7384, n7385, n7386, n7387, n7388,
    n7389, n7390, n7391, n7392, n7393, n7394,
    n7395, n7396, n7397, n7398, n7399, n7400,
    n7401, n7402, n7403, n7404, n7405, n7406,
    n7407, n7408, n7409, n7410, n7411, n7412,
    n7413, n7414, n7415, n7416, n7417, n7418,
    n7419, n7420, n7421, n7422, n7423, n7424,
    n7425, n7426, n7427, n7428, n7429, n7430,
    n7431, n7432, n7433, n7434, n7435, n7436,
    n7437, n7438, n7439, n7440, n7441, n7442,
    n7443, n7444, n7445, n7446, n7447, n7448,
    n7449, n7450, n7451, n7452, n7453, n7454,
    n7455, n7456, n7457, n7458, n7459, n7460,
    n7461, n7462, n7463, n7464, n7465, n7466,
    n7467, n7468, n7469, n7470, n7471, n7472,
    n7473, n7474, n7475, n7476, n7477, n7478,
    n7479, n7480, n7481, n7482, n7483, n7484,
    n7485, n7486, n7487, n7488, n7489, n7490,
    n7491, n7492, n7493, n7494, n7495, n7496,
    n7497, n7498, n7499, n7500, n7501, n7502,
    n7503, n7504, n7505, n7506, n7507, n7508,
    n7509, n7510, n7511, n7512, n7513, n7514,
    n7515, n7516, n7517, n7518, n7519, n7520,
    n7521, n7522, n7523, n7524, n7525, n7526,
    n7527, n7528, n7529, n7530, n7531, n7532,
    n7533, n7534, n7535, n7536, n7537, n7538,
    n7539, n7540, n7541, n7542, n7543, n7544,
    n7545, n7546, n7547, n7548, n7549, n7550,
    n7551, n7552, n7553, n7554, n7555, n7556,
    n7557, n7558, n7559, n7560, n7561, n7562,
    n7563, n7564, n7565, n7566, n7567, n7568,
    n7569, n7570, n7571, n7572, n7573, n7574,
    n7575, n7576, n7577, n7578, n7579, n7580,
    n7581, n7582, n7583, n7584, n7585, n7586,
    n7587, n7588, n7589, n7590, n7591, n7592,
    n7593, n7594, n7595, n7596, n7597, n7598,
    n7599, n7600, n7601, n7602, n7603, n7604,
    n7605, n7606, n7607, n7608, n7609, n7610,
    n7611, n7612, n7613, n7614, n7615, n7616,
    n7617, n7618, n7619, n7620, n7621, n7622,
    n7623, n7624, n7625, n7626, n7627, n7628,
    n7629, n7630, n7631, n7632, n7633, n7634,
    n7635, n7636, n7637, n7638, n7639, n7640,
    n7641, n7642, n7643, n7644, n7645, n7646,
    n7647, n7648, n7649, n7650, n7651, n7652,
    n7653, n7654, n7655, n7656, n7657, n7658,
    n7659, n7660, n7661, n7662, n7663, n7664,
    n7665, n7666, n7667, n7668, n7669, n7670,
    n7671, n7672, n7673, n7674, n7675, n7676,
    n7677, n7678, n7679, n7680, n7681, n7682,
    n7683, n7684, n7685, n7686, n7687, n7688,
    n7689, n7690, n7691, n7692, n7693, n7694,
    n7695, n7696, n7697, n7698, n7699, n7700,
    n7701, n7702, n7703, n7704, n7705, n7706,
    n7707, n7708, n7709, n7710, n7711, n7712,
    n7713, n7714, n7715, n7716, n7717, n7718,
    n7719, n7720, n7721, n7722, n7723, n7724,
    n7725, n7726, n7727, n7728, n7729, n7730,
    n7731, n7732, n7733, n7734, n7735, n7736,
    n7737, n7738, n7739, n7740, n7741, n7742,
    n7743, n7744, n7745, n7746, n7747, n7748,
    n7749, n7750, n7751, n7752, n7753, n7754,
    n7755, n7756, n7757, n7758, n7759, n7760,
    n7761, n7762, n7763, n7764, n7765, n7766,
    n7767, n7768, n7769, n7770, n7771, n7772,
    n7773, n7774, n7775, n7776, n7777, n7778,
    n7779, n7780, n7781, n7782, n7783, n7784,
    n7785, n7786, n7787, n7788, n7789, n7790,
    n7791, n7792, n7793, n7794, n7795, n7796,
    n7797, n7798, n7799, n7800, n7801, n7802,
    n7803, n7804, n7805, n7806, n7807, n7808,
    n7809, n7810, n7811, n7812, n7813, n7814,
    n7815, n7816, n7817, n7818, n7819, n7820,
    n7821, n7822, n7823, n7824, n7825, n7826,
    n7827, n7828, n7829, n7830, n7831, n7832,
    n7833, n7834, n7835, n7836, n7837, n7838,
    n7839, n7840, n7841, n7842, n7843, n7844,
    n7845, n7846, n7847, n7848, n7849, n7850,
    n7851, n7852, n7853, n7854, n7855, n7856,
    n7857, n7858, n7859, n7860, n7861, n7862,
    n7863, n7864, n7865, n7866, n7867, n7868,
    n7869, n7870, n7871, n7872, n7873, n7874,
    n7875, n7876, n7877, n7878, n7879, n7880,
    n7881, n7882, n7883, n7884, n7885, n7886,
    n7887, n7888, n7889, n7890, n7891, n7892,
    n7893, n7894, n7895, n7896, n7897, n7898,
    n7899, n7900, n7901, n7902, n7903, n7904,
    n7905, n7906, n7907, n7908, n7909, n7910,
    n7911, n7912, n7913, n7914, n7915, n7916,
    n7917, n7918, n7919, n7920, n7921, n7922,
    n7923, n7924, n7925, n7926, n7927, n7928,
    n7929, n7930, n7931, n7932, n7933, n7934,
    n7935, n7936, n7937, n7938, n7939, n7940,
    n7941, n7942, n7943, n7944, n7945, n7946,
    n7947, n7948, n7949, n7950, n7951, n7952,
    n7953, n7954, n7955, n7956, n7957, n7958,
    n7959, n7960, n7961, n7962, n7963, n7964,
    n7965, n7966, n7967, n7968, n7969, n7970,
    n7971, n7972, n7973, n7974, n7975, n7976,
    n7977, n7978, n7979, n7980, n7981, n7982,
    n7983, n7984, n7985, n7986, n7987, n7988,
    n7989, n7990, n7991, n7992, n7993, n7994,
    n7995, n7996, n7997, n7998, n7999, n8000,
    n8001, n8002, n8003, n8004, n8005, n8006,
    n8007, n8008, n8009, n8010, n8011, n8012,
    n8013, n8014, n8015, n8016, n8017, n8018,
    n8019, n8020, n8021, n8022, n8023, n8024,
    n8025, n8026, n8027, n8028, n8029, n8030,
    n8031, n8032, n8033, n8034, n8035, n8036,
    n8037, n8038, n8039, n8040, n8041, n8042,
    n8043, n8044, n8045, n8046, n8047, n8048,
    n8049, n8050, n8051, n8052, n8053, n8054,
    n8055, n8056, n8057, n8058, n8059, n8060,
    n8061, n8062, n8063, n8064, n8065, n8066,
    n8067, n8068, n8069, n8070, n8071, n8072,
    n8073, n8074, n8075, n8076, n8077, n8078,
    n8079, n8080, n8081, n8082, n8083, n8084,
    n8085, n8086, n8087, n8088, n8089, n8090,
    n8091, n8092, n8093, n8094, n8095, n8096,
    n8097, n8098, n8099, n8100, n8101, n8102,
    n8103, n8104, n8105, n8106, n8107, n8108,
    n8109, n8110, n8111, n8112, n8113, n8114,
    n8115, n8116, n8117, n8118, n8119, n8120,
    n8121, n8122, n8123, n8124, n8125, n8126,
    n8127, n8128, n8129, n8130, n8131, n8132,
    n8133, n8134, n8135, n8136, n8137, n8138,
    n8139, n8140, n8141, n8142, n8143, n8144,
    n8145, n8146, n8147, n8148, n8149, n8150,
    n8151, n8152, n8153, n8154, n8155, n8156,
    n8157, n8158, n8159, n8160, n8161, n8162,
    n8163, n8164, n8165, n8166, n8167, n8168,
    n8169, n8170, n8171, n8172, n8173, n8174,
    n8175, n8176, n8177, n8178, n8179, n8180,
    n8181, n8182, n8183, n8184, n8185, n8186,
    n8187, n8188, n8189, n8190, n8191, n8192,
    n8193, n8194, n8195, n8196, n8197, n8198,
    n8199, n8200, n8201, n8202, n8203, n8204,
    n8205, n8206, n8207, n8208, n8209, n8210,
    n8211, n8212, n8213, n8214, n8215, n8216,
    n8217, n8218, n8219, n8220, n8221, n8222,
    n8223, n8224, n8225, n8226, n8227, n8228,
    n8229, n8230, n8231, n8232, n8233, n8234,
    n8235, n8236, n8237, n8238, n8239, n8240,
    n8241, n8242, n8243, n8244, n8245, n8246,
    n8247, n8248, n8249, n8250, n8251, n8252,
    n8253, n8254, n8255, n8256, n8257, n8258,
    n8259, n8260, n8261, n8262, n8263, n8264,
    n8265, n8266, n8267, n8268, n8269, n8270,
    n8271, n8272, n8273, n8274, n8275, n8276,
    n8277, n8278, n8279, n8280, n8281, n8282,
    n8283, n8284, n8285, n8286, n8287, n8288,
    n8289, n8290, n8291, n8292, n8293, n8294,
    n8295, n8296, n8297, n8298, n8299, n8300,
    n8301, n8302, n8303, n8304, n8305, n8306,
    n8307, n8308, n8309, n8310, n8311, n8312,
    n8313, n8314, n8315, n8316, n8317, n8318,
    n8319, n8320, n8321, n8322, n8323, n8324,
    n8325, n8326, n8327, n8328, n8329, n8330,
    n8331, n8332, n8333, n8334, n8335, n8336,
    n8337, n8338, n8339, n8340, n8341, n8342,
    n8343, n8344, n8345, n8346, n8347, n8348,
    n8349, n8350, n8351, n8352, n8353, n8354,
    n8355, n8356, n8357, n8358, n8359, n8360,
    n8361, n8362, n8363, n8364, n8365, n8366,
    n8367, n8368, n8369, n8370, n8371, n8372,
    n8373, n8374, n8375, n8376, n8377, n8378,
    n8379, n8380, n8381, n8382, n8383, n8384,
    n8385, n8386, n8387, n8388, n8389, n8390,
    n8391, n8392, n8393, n8394, n8395, n8396,
    n8397, n8398, n8399, n8400, n8401, n8402,
    n8403, n8404, n8405, n8406, n8407, n8408,
    n8409, n8410, n8411, n8412, n8413, n8414,
    n8415, n8416, n8417, n8418, n8419, n8420,
    n8421, n8422, n8423, n8424, n8425, n8426,
    n8427, n8428, n8429, n8430, n8431, n8432,
    n8433, n8434, n8435, n8436, n8437, n8438,
    n8439, n8440, n8441, n8442, n8443, n8444,
    n8445, n8446, n8447, n8448, n8449, n8450,
    n8451, n8452, n8453, n8454, n8455, n8456,
    n8457, n8458, n8459, n8460, n8461, n8462,
    n8463, n8464, n8465, n8466, n8467, n8468,
    n8469, n8470, n8471, n8472, n8473, n8474,
    n8475, n8476, n8477, n8478, n8479, n8480,
    n8481, n8482, n8483, n8484, n8485, n8486,
    n8487, n8488, n8489, n8490, n8491, n8492,
    n8493, n8494, n8495, n8496, n8497, n8498,
    n8499, n8500, n8501, n8502, n8503, n8504,
    n8505, n8506, n8507, n8508, n8509, n8510,
    n8511, n8512, n8513, n8514, n8515, n8516,
    n8517, n8518, n8519, n8520, n8521, n8522,
    n8523, n8524, n8525, n8526, n8527, n8528,
    n8529, n8530, n8531, n8532, n8533, n8534,
    n8535, n8536, n8537, n8538, n8539, n8540,
    n8541, n8542, n8543, n8544, n8545, n8546,
    n8547, n8548, n8549, n8550, n8551, n8552,
    n8553, n8554, n8555, n8556, n8557, n8558,
    n8559, n8560, n8561, n8562, n8563, n8564,
    n8565, n8566, n8567, n8568, n8569, n8570,
    n8571, n8572, n8573, n8574, n8575, n8576,
    n8577, n8578, n8579, n8580, n8581, n8582,
    n8583, n8584, n8585, n8586, n8587, n8588,
    n8589, n8590, n8591, n8592, n8593, n8594,
    n8595, n8596, n8597, n8598, n8599, n8600,
    n8601, n8602, n8603, n8604, n8605, n8606,
    n8607, n8608, n8609, n8610, n8611, n8612,
    n8613, n8614, n8615, n8616, n8617, n8618,
    n8619, n8620, n8621, n8622, n8623, n8624,
    n8625, n8626, n8627, n8628, n8629, n8630,
    n8631, n8632, n8633, n8634, n8635, n8636,
    n8637, n8638, n8639, n8640, n8641, n8642,
    n8643, n8644, n8645, n8646, n8647, n8648,
    n8649, n8650, n8651, n8652, n8653, n8654,
    n8655, n8656, n8657, n8658, n8659, n8660,
    n8661, n8662, n8663, n8664, n8665, n8666,
    n8667, n8668, n8669, n8670, n8671, n8672,
    n8673, n8674, n8675, n8676, n8677, n8678,
    n8679, n8680, n8681, n8682, n8683, n8684,
    n8685, n8686, n8687, n8688, n8689, n8690,
    n8691, n8692, n8693, n8694, n8695, n8696,
    n8697, n8698, n8699, n8700, n8701, n8702,
    n8703, n8704, n8705, n8706, n8707, n8708,
    n8709, n8710, n8711, n8712, n8713, n8714,
    n8715, n8716, n8717, n8718, n8719, n8720,
    n8721, n8722, n8723, n8724, n8725, n8726,
    n8727, n8728, n8729, n8730, n8731, n8732,
    n8733, n8734, n8735, n8736, n8737, n8738,
    n8739, n8740, n8741, n8742, n8743, n8744,
    n8745, n8746, n8747, n8748, n8749, n8750,
    n8751, n8752, n8753, n8754, n8755, n8756,
    n8757, n8758, n8759, n8760, n8761, n8762,
    n8763, n8764, n8765, n8766, n8767, n8768,
    n8769, n8770, n8771, n8772, n8773, n8774,
    n8775, n8776, n8777, n8778, n8779, n8780,
    n8781, n8782, n8783, n8784, n8785, n8786,
    n8787, n8788, n8789, n8790, n8791, n8792,
    n8793, n8794, n8795, n8796, n8797, n8798,
    n8799, n8800, n8801, n8802, n8803, n8804,
    n8805, n8806, n8807, n8808, n8809, n8810,
    n8811, n8812, n8813, n8814, n8815, n8816,
    n8817, n8818, n8819, n8820, n8821, n8822,
    n8823, n8824, n8825, n8826, n8827, n8828,
    n8829, n8830, n8831, n8832, n8833, n8834,
    n8835, n8836, n8837, n8838, n8839, n8840,
    n8841, n8842, n8843, n8844, n8845, n8846,
    n8847, n8848, n8849, n8850, n8851, n8852,
    n8853, n8854, n8855, n8856, n8857, n8858,
    n8859, n8860, n8861, n8862, n8863, n8864,
    n8865, n8866, n8867, n8868, n8869, n8870,
    n8871, n8872, n8873, n8874, n8875, n8876,
    n8877, n8878, n8879, n8880, n8881, n8882,
    n8883, n8884, n8885, n8886, n8887, n8888,
    n8889, n8890, n8891, n8892, n8893, n8894,
    n8895, n8896, n8897, n8898, n8899, n8900,
    n8901, n8902, n8903, n8904, n8905, n8906,
    n8907, n8908, n8909, n8910, n8911, n8912,
    n8913, n8914, n8915, n8916, n8917, n8918,
    n8919, n8920, n8921, n8922, n8923, n8924,
    n8925, n8926, n8927, n8928, n8929, n8930,
    n8931, n8932, n8933, n8934, n8935, n8936,
    n8937, n8938, n8939, n8940, n8941, n8942,
    n8943, n8944, n8945, n8946, n8947, n8948,
    n8949, n8950, n8951, n8952, n8953, n8954,
    n8955, n8956, n8957, n8958, n8959, n8960,
    n8961, n8962, n8963, n8964, n8965, n8966,
    n8967, n8968, n8969, n8970, n8971, n8972,
    n8973, n8974, n8975, n8976, n8977, n8978,
    n8979, n8980, n8981, n8982, n8983, n8984,
    n8985, n8986, n8987, n8988, n8989, n8990,
    n8991, n8992, n8993, n8994, n8995, n8996,
    n8997, n8998, n8999, n9000, n9001, n9002,
    n9003, n9004, n9005, n9006, n9007, n9008,
    n9009, n9010, n9011, n9012, n9013, n9014,
    n9015, n9016, n9017, n9018, n9019, n9020,
    n9021, n9022, n9023, n9024, n9025, n9026,
    n9027, n9028, n9029, n9030, n9031, n9032,
    n9033, n9034, n9035, n9036, n9037, n9038,
    n9039, n9040, n9041, n9042, n9043, n9044,
    n9045, n9046, n9047, n9048, n9049, n9050,
    n9051, n9052, n9053, n9054, n9055, n9056,
    n9057, n9058, n9059, n9060, n9061, n9062,
    n9063, n9064, n9065, n9066, n9067, n9068,
    n9069, n9070, n9071, n9072, n9073, n9074,
    n9075, n9076, n9077, n9078, n9079, n9080,
    n9081, n9082, n9083, n9084, n9085, n9086,
    n9087, n9088, n9089, n9090, n9091, n9092,
    n9093, n9094, n9095, n9096, n9097, n9098,
    n9099, n9100, n9101, n9102, n9103, n9104,
    n9105, n9106, n9107, n9108, n9109, n9110,
    n9111, n9112, n9113, n9114, n9115, n9116,
    n9117, n9118, n9119, n9120, n9121, n9122,
    n9123, n9124, n9125, n9126, n9127, n9128,
    n9129, n9130, n9131, n9132, n9133, n9134,
    n9135, n9136, n9137, n9138, n9139, n9140,
    n9141, n9142, n9143, n9144, n9145, n9146,
    n9147, n9148, n9149, n9150, n9151, n9152,
    n9153, n9154, n9155, n9156, n9157, n9158,
    n9159, n9160, n9161, n9162, n9163, n9164,
    n9165, n9166, n9167, n9168, n9169, n9170,
    n9171, n9172, n9173, n9174, n9175, n9176,
    n9177, n9178, n9179, n9180, n9181, n9182,
    n9183, n9184, n9185, n9186, n9187, n9188,
    n9189, n9190, n9191, n9192, n9193, n9194,
    n9195, n9196, n9197, n9198, n9199, n9200,
    n9201, n9202, n9203, n9204, n9205, n9206,
    n9207, n9208, n9209, n9210, n9211, n9212,
    n9213, n9214, n9215, n9216, n9217, n9218,
    n9219, n9220, n9221, n9222, n9223, n9224,
    n9225, n9226, n9227, n9228, n9229, n9230,
    n9231, n9232, n9233, n9234, n9235, n9236,
    n9237, n9238, n9239, n9240, n9241, n9242,
    n9243, n9244, n9245, n9246, n9247, n9248,
    n9249, n9250, n9251, n9252, n9253, n9254,
    n9255, n9256, n9257, n9258, n9259, n9260,
    n9261, n9262, n9263, n9264, n9265, n9266,
    n9267, n9268, n9269, n9270, n9271, n9272,
    n9273, n9274, n9275, n9276, n9277, n9278,
    n9279, n9280, n9281, n9282, n9283, n9284,
    n9285, n9286, n9287, n9288, n9289, n9290,
    n9291, n9292, n9293, n9294, n9295, n9296,
    n9297, n9298, n9299, n9300, n9301, n9302,
    n9303, n9304, n9305, n9306, n9307, n9308,
    n9309, n9310, n9311, n9312, n9313, n9314,
    n9315, n9316, n9317, n9318, n9319, n9320,
    n9321, n9322, n9323, n9324, n9325, n9326,
    n9327, n9328, n9329, n9330, n9331, n9332,
    n9333, n9334, n9335, n9336, n9337, n9338,
    n9339, n9340, n9341, n9342, n9343, n9344,
    n9345, n9346, n9347, n9348, n9349, n9350,
    n9351, n9352, n9353, n9354, n9355, n9356,
    n9357, n9358, n9359, n9360, n9361, n9362,
    n9363, n9364, n9365, n9366, n9367, n9368,
    n9369, n9370, n9371, n9372, n9373, n9374,
    n9375, n9376, n9377, n9378, n9379, n9380,
    n9381, n9382, n9383, n9384, n9385, n9386,
    n9387, n9388, n9389, n9390, n9391, n9392,
    n9393, n9394, n9395, n9396, n9397, n9398,
    n9399, n9400, n9401, n9402, n9403, n9404,
    n9405, n9406, n9407, n9408, n9409, n9410,
    n9411, n9412, n9413, n9414, n9415, n9416,
    n9417, n9418, n9419, n9420, n9421, n9422,
    n9423, n9424, n9425, n9426, n9427, n9428,
    n9429, n9430, n9431, n9432, n9433, n9434,
    n9435, n9436, n9437, n9438, n9439, n9440,
    n9441, n9442, n9443, n9444, n9445, n9446,
    n9447, n9448, n9449, n9450, n9451, n9452,
    n9453, n9454, n9455, n9456, n9457, n9458,
    n9459, n9460, n9461, n9462, n9463, n9464,
    n9465, n9466, n9467, n9468, n9469, n9470,
    n9471, n9472, n9473, n9474, n9475, n9476,
    n9477, n9478, n9479, n9480, n9481, n9482,
    n9483, n9484, n9485, n9486, n9487, n9488,
    n9489, n9490, n9491, n9492, n9493, n9494,
    n9495, n9496, n9497, n9498, n9499, n9500,
    n9501, n9502, n9503, n9504, n9505, n9506,
    n9507, n9508, n9509, n9510, n9511, n9512,
    n9513, n9514, n9515, n9516, n9517, n9518,
    n9519, n9520, n9521, n9522, n9523, n9524,
    n9525, n9526, n9527, n9528, n9529, n9530,
    n9531, n9532, n9533, n9534, n9535, n9536,
    n9537, n9538, n9539, n9540, n9541, n9542,
    n9543, n9544, n9545, n9546, n9547, n9548,
    n9549, n9550, n9551, n9552, n9553, n9554,
    n9555, n9556, n9557, n9558, n9559, n9560,
    n9561, n9562, n9563, n9564, n9565, n9566,
    n9567, n9568, n9569, n9570, n9571, n9572,
    n9573, n9574, n9575, n9576, n9577, n9578,
    n9579, n9580, n9581, n9582, n9583, n9584,
    n9585, n9586, n9587, n9588, n9589, n9590,
    n9591, n9592, n9593, n9594, n9595, n9596,
    n9597, n9598, n9599, n9600, n9601, n9602,
    n9603, n9604, n9605, n9606, n9607, n9608,
    n9609, n9610, n9611, n9612, n9613, n9614,
    n9615, n9616, n9617, n9618, n9619, n9620,
    n9621, n9622, n9623, n9624, n9625, n9626,
    n9627, n9628, n9629, n9630, n9631, n9632,
    n9633, n9634, n9635, n9636, n9637, n9638,
    n9639, n9640, n9641, n9642, n9643, n9644,
    n9645, n9646, n9647, n9648, n9649, n9650,
    n9651, n9652, n9653, n9654, n9655, n9656,
    n9657, n9658, n9659, n9660, n9661, n9662,
    n9663, n9664, n9665, n9666, n9667, n9668,
    n9669, n9670, n9671, n9672, n9673, n9674,
    n9675, n9676, n9677, n9678, n9679, n9680,
    n9681, n9682, n9683, n9684, n9685, n9686,
    n9687, n9688, n9689, n9690, n9691, n9692,
    n9693, n9694, n9695, n9696, n9697, n9698,
    n9699, n9700, n9701, n9702, n9703, n9704,
    n9705, n9706, n9707, n9708, n9709, n9710,
    n9711, n9712, n9713, n9714, n9715, n9716,
    n9717, n9718, n9719, n9720, n9721, n9722,
    n9723, n9724, n9725, n9726, n9727, n9728,
    n9729, n9730, n9731, n9732, n9733, n9734,
    n9735, n9736, n9737, n9738, n9739, n9740,
    n9741, n9742, n9743, n9744, n9745, n9746,
    n9747, n9748, n9749, n9750, n9751, n9752,
    n9753, n9754, n9755, n9756, n9757, n9758,
    n9759, n9760, n9761, n9762, n9763, n9764,
    n9765, n9766, n9767, n9768, n9769, n9770,
    n9771, n9772, n9773, n9774, n9775, n9776,
    n9777, n9778, n9779, n9780, n9781, n9782,
    n9783, n9784, n9785, n9786, n9787, n9788,
    n9789, n9790, n9791, n9792, n9793, n9794,
    n9795, n9796, n9797, n9798, n9799, n9800,
    n9801, n9802, n9803, n9804, n9805, n9806,
    n9807, n9808, n9809, n9810, n9811, n9812,
    n9813, n9814, n9815, n9816, n9817, n9818,
    n9819, n9820, n9821, n9822, n9823, n9824,
    n9825, n9826, n9827, n9828, n9829, n9830,
    n9831, n9832, n9833, n9834, n9835, n9836,
    n9837, n9838, n9839, n9840, n9841, n9842,
    n9843, n9844, n9845, n9846, n9847, n9848,
    n9849, n9850, n9851, n9852, n9853, n9854,
    n9855, n9856, n9857, n9858, n9859, n9860,
    n9861, n9862, n9863, n9864, n9865, n9866,
    n9867, n9868, n9869, n9870, n9871, n9872,
    n9873, n9874, n9875, n9876, n9877, n9878,
    n9879, n9880, n9881, n9882, n9883, n9884,
    n9885, n9886, n9887, n9888, n9889, n9890,
    n9891, n9892, n9893, n9894, n9895, n9896,
    n9897, n9898, n9899, n9900, n9901, n9902,
    n9903, n9904, n9905, n9906, n9907, n9908,
    n9909, n9910, n9911, n9912, n9913, n9914,
    n9915, n9916, n9917, n9918, n9919, n9920,
    n9921, n9922, n9923, n9924, n9925, n9926,
    n9927, n9928, n9929, n9930, n9931, n9932,
    n9933, n9934, n9935, n9936, n9937, n9938,
    n9939, n9940, n9941, n9942, n9943, n9944,
    n9945, n9946, n9947, n9948, n9949, n9950,
    n9951, n9952, n9953, n9954, n9955, n9956,
    n9957, n9958, n9959, n9960, n9961, n9962,
    n9963, n9964, n9965, n9966, n9967, n9968,
    n9969, n9970, n9971, n9972, n9973, n9974,
    n9975, n9976, n9977, n9978, n9979, n9980,
    n9981, n9982, n9983, n9984, n9985, n9986,
    n9987, n9988, n9989, n9990, n9991, n9992,
    n9993, n9994, n9995, n9996, n9997, n9998,
    n9999, n10000, n10001, n10002, n10003, n10004,
    n10005, n10006, n10007, n10008, n10009, n10010,
    n10011, n10012, n10013, n10014, n10015, n10016,
    n10017, n10018, n10019, n10020, n10021, n10022,
    n10023, n10024, n10025, n10026, n10027, n10028,
    n10029, n10030, n10031, n10032, n10033, n10034,
    n10035, n10036, n10037, n10038, n10039, n10040,
    n10041, n10042, n10043, n10044, n10045, n10046,
    n10047, n10048, n10049, n10050, n10051, n10052,
    n10053, n10054, n10055, n10056, n10057, n10058,
    n10059, n10060, n10061, n10062, n10063, n10064,
    n10065, n10066, n10067, n10068, n10069, n10070,
    n10071, n10072, n10073, n10074, n10075, n10076,
    n10077, n10078, n10079, n10080, n10081, n10082,
    n10083, n10084, n10085, n10086, n10087, n10088,
    n10089, n10090, n10091, n10092, n10093, n10094,
    n10095, n10096, n10097, n10098, n10099, n10100,
    n10101, n10102, n10103, n10104, n10105, n10106,
    n10107, n10108, n10109, n10110, n10111, n10112,
    n10113, n10114, n10115, n10116, n10117, n10118,
    n10119, n10120, n10121, n10122, n10123, n10124,
    n10125, n10126, n10127, n10128, n10129, n10130,
    n10131, n10132, n10133, n10134, n10135, n10136,
    n10137, n10138, n10139, n10140, n10141, n10142,
    n10143, n10144, n10145, n10146, n10147, n10148,
    n10149, n10150, n10151, n10152, n10153, n10154,
    n10155, n10156, n10157, n10158, n10159, n10160,
    n10161, n10162, n10163, n10164, n10165, n10166,
    n10167, n10168, n10169, n10170, n10171, n10172,
    n10173, n10174, n10175, n10176, n10177, n10178,
    n10179, n10180, n10181, n10182, n10183, n10184,
    n10185, n10186, n10187, n10188, n10189, n10190,
    n10191, n10192, n10193, n10194, n10195, n10196,
    n10197, n10198, n10199, n10200, n10201, n10202,
    n10203, n10204, n10205, n10206, n10207, n10208,
    n10209, n10210, n10211, n10212, n10213, n10214,
    n10215, n10216, n10217, n10218, n10219, n10220,
    n10221, n10222, n10223, n10224, n10225, n10226,
    n10227, n10228, n10229, n10230, n10231, n10232,
    n10233, n10234, n10235, n10236, n10237, n10238,
    n10239, n10240, n10241, n10242, n10243, n10244,
    n10245, n10246, n10247, n10248, n10249, n10250,
    n10251, n10252, n10253, n10254, n10255, n10256,
    n10257, n10258, n10259, n10260, n10261, n10262,
    n10263, n10264, n10265, n10266, n10267, n10268,
    n10269, n10270, n10271, n10272, n10273, n10274,
    n10275, n10276, n10277, n10278, n10279, n10280,
    n10281, n10282, n10283, n10284, n10285, n10286,
    n10287, n10288, n10289, n10290, n10291, n10292,
    n10293, n10294, n10295, n10296, n10297, n10298,
    n10299, n10300, n10301, n10302, n10303, n10304,
    n10305, n10306, n10307, n10308, n10309, n10310,
    n10311, n10312, n10313, n10314, n10315, n10316,
    n10317, n10318, n10319, n10320, n10321, n10322,
    n10323, n10324, n10325, n10326, n10327, n10328,
    n10329, n10330, n10331, n10332, n10333, n10334,
    n10335, n10336, n10337, n10338, n10339, n10340,
    n10341, n10342, n10343, n10344, n10345, n10346,
    n10347, n10348, n10349, n10350, n10351, n10352,
    n10353, n10354, n10355, n10356, n10357, n10358,
    n10359, n10360, n10361, n10362, n10363, n10364,
    n10365, n10366, n10367, n10368, n10369, n10370,
    n10371, n10372, n10373, n10374, n10375, n10376,
    n10377, n10378, n10379, n10380, n10381, n10382,
    n10383, n10384, n10385, n10386, n10387, n10388,
    n10389, n10390, n10391, n10392, n10393, n10394,
    n10395, n10396, n10397, n10398, n10399, n10400,
    n10401, n10402, n10403, n10404, n10405, n10406,
    n10407, n10408, n10409, n10410, n10411, n10412,
    n10413, n10414, n10415, n10416, n10417, n10418,
    n10419, n10420, n10421, n10422, n10423, n10424,
    n10425, n10426, n10427, n10428, n10429, n10430,
    n10431, n10432, n10433, n10434, n10435, n10436,
    n10437, n10438, n10439, n10440, n10441, n10442,
    n10443, n10444, n10445, n10446, n10447, n10448,
    n10449, n10450, n10451, n10452, n10453, n10454,
    n10455, n10456, n10457, n10458, n10459, n10460,
    n10461, n10462, n10463, n10464, n10465, n10466,
    n10467, n10468, n10469, n10470, n10471, n10472,
    n10473, n10474, n10475, n10476, n10477, n10478,
    n10479, n10480, n10481, n10482, n10483, n10484,
    n10485, n10486, n10487, n10488, n10489, n10490,
    n10491, n10492, n10493, n10494, n10495, n10496,
    n10497, n10498, n10499, n10500, n10501, n10502,
    n10503, n10504, n10505, n10506, n10507, n10508,
    n10509, n10510, n10511, n10512, n10513, n10514,
    n10515, n10516, n10517, n10518, n10519, n10520,
    n10521, n10522, n10523, n10524, n10525, n10526,
    n10527, n10528, n10529, n10530, n10531, n10532,
    n10533, n10534, n10535, n10536, n10537, n10538,
    n10539, n10540, n10541, n10542, n10543, n10544,
    n10545, n10546, n10547, n10548, n10549, n10550,
    n10551, n10552, n10553, n10554, n10555, n10556,
    n10557, n10558, n10559, n10560, n10561, n10562,
    n10563, n10564, n10565, n10566, n10567, n10568,
    n10569, n10570, n10571, n10572, n10573, n10574,
    n10575, n10576, n10577, n10578, n10579, n10580,
    n10581, n10582, n10583, n10584, n10585, n10586,
    n10587, n10588, n10589, n10590, n10591, n10592,
    n10593, n10594, n10595, n10596, n10597, n10598,
    n10599, n10600, n10601, n10602, n10603, n10604,
    n10605, n10606, n10607, n10608, n10609, n10610,
    n10611, n10612, n10613, n10614, n10615, n10616,
    n10617, n10618, n10619, n10620, n10621, n10622,
    n10623, n10624, n10625, n10626, n10627, n10628,
    n10629, n10630, n10631, n10632, n10633, n10634,
    n10635, n10636, n10637, n10638, n10639, n10640,
    n10641, n10642, n10643, n10644, n10645, n10646,
    n10647, n10648, n10649, n10650, n10651, n10652,
    n10653, n10654, n10655, n10656, n10657, n10658,
    n10659, n10660, n10661, n10662, n10663, n10664,
    n10665, n10666, n10667, n10668, n10669, n10670,
    n10671, n10672, n10673, n10674, n10675, n10676,
    n10677, n10678, n10679, n10680, n10681, n10682,
    n10683, n10684, n10685, n10686, n10687, n10688,
    n10689, n10690, n10691, n10692, n10693, n10694,
    n10695, n10696, n10697, n10698, n10699, n10700,
    n10701, n10702, n10703, n10704, n10705, n10706,
    n10707, n10708, n10709, n10710, n10711, n10712,
    n10713, n10714, n10715, n10716, n10717, n10718,
    n10719, n10720, n10721, n10722, n10723, n10724,
    n10725, n10726, n10727, n10728, n10729, n10730,
    n10731, n10732, n10733, n10734, n10735, n10736,
    n10737, n10738, n10739, n10740, n10741, n10742,
    n10743, n10744, n10745, n10746, n10747, n10748,
    n10749, n10750, n10751, n10752, n10753, n10754,
    n10755, n10756, n10757, n10758, n10759, n10760,
    n10761, n10762, n10763, n10764, n10765, n10766,
    n10767, n10768, n10769, n10770, n10771, n10772,
    n10773, n10774, n10775, n10776, n10777, n10778,
    n10779, n10780, n10781, n10782, n10783, n10784,
    n10785, n10786, n10787, n10788, n10789, n10790,
    n10791, n10792, n10793, n10794, n10795, n10796,
    n10797, n10798, n10799, n10800, n10801, n10802,
    n10803, n10804, n10805, n10806, n10807, n10808,
    n10809, n10810, n10811, n10812, n10813, n10814,
    n10815, n10816, n10817, n10818, n10819, n10820,
    n10821, n10822, n10823, n10824, n10825, n10826,
    n10827, n10828, n10829, n10830, n10831, n10832,
    n10833, n10834, n10835, n10836, n10837, n10838,
    n10839, n10840, n10841, n10842, n10843, n10844,
    n10845, n10846, n10847, n10848, n10849, n10850,
    n10851, n10852, n10853, n10854, n10855, n10856,
    n10857, n10858, n10859, n10860, n10861, n10862,
    n10863, n10864, n10865, n10866, n10867, n10868,
    n10869, n10870, n10871, n10872, n10873, n10874,
    n10875, n10876, n10877, n10878, n10879, n10880,
    n10881, n10882, n10883, n10884, n10885, n10886,
    n10887, n10888, n10889, n10890, n10891, n10892,
    n10893, n10894, n10895, n10896, n10897, n10898,
    n10899, n10900, n10901, n10902, n10903, n10904,
    n10905, n10906, n10907, n10908, n10909, n10910,
    n10911, n10912, n10913, n10914, n10915, n10916,
    n10917, n10918, n10919, n10920, n10921, n10922,
    n10923, n10924, n10925, n10926, n10927, n10928,
    n10929, n10930, n10931, n10932, n10933, n10934,
    n10935, n10936, n10937, n10938, n10939, n10940,
    n10941, n10942, n10943, n10944, n10945, n10946,
    n10947, n10948, n10949, n10950, n10951, n10952,
    n10953, n10954, n10955, n10956, n10957, n10958,
    n10959, n10960, n10961, n10962, n10963, n10964,
    n10965, n10966, n10967, n10968, n10969, n10970,
    n10971, n10972, n10973, n10974, n10975, n10976,
    n10977, n10978, n10979, n10980, n10981, n10982,
    n10983, n10984, n10985, n10986, n10987, n10988,
    n10989, n10990, n10991, n10992, n10993, n10994,
    n10995, n10996, n10997, n10998, n10999, n11000,
    n11001, n11002, n11003, n11004, n11005, n11006,
    n11007, n11008, n11009, n11010, n11011, n11012,
    n11013, n11014, n11015, n11016, n11017, n11018,
    n11019, n11020, n11021, n11022, n11023, n11024,
    n11025, n11026, n11027, n11028, n11029, n11030,
    n11031, n11032, n11033, n11034, n11035, n11036,
    n11037, n11038, n11039, n11040, n11041, n11042,
    n11043, n11044, n11045, n11046, n11047, n11048,
    n11049, n11050, n11051, n11052, n11053, n11054,
    n11055, n11056, n11057, n11058, n11059, n11060,
    n11061, n11062, n11063, n11064, n11065, n11066,
    n11067, n11068, n11069, n11070, n11071, n11072,
    n11073, n11074, n11075, n11076, n11077, n11078,
    n11079, n11080, n11081, n11082, n11083, n11084,
    n11085, n11086, n11087, n11088, n11089, n11090,
    n11091, n11092, n11093, n11094, n11095, n11096,
    n11097, n11098, n11099, n11100, n11101, n11102,
    n11103, n11104, n11105, n11106, n11107, n11108,
    n11109, n11110, n11111, n11112, n11113, n11114,
    n11115, n11116, n11117, n11118, n11119, n11120,
    n11121, n11122, n11123, n11124, n11125, n11126,
    n11127, n11128, n11129, n11130, n11131, n11132,
    n11133, n11134, n11135, n11136, n11137, n11138,
    n11139, n11140, n11141, n11142, n11143, n11144,
    n11145, n11146, n11147, n11148, n11149, n11150,
    n11151, n11152, n11153, n11154, n11155, n11156,
    n11157, n11158, n11159, n11160, n11161, n11162,
    n11163, n11164, n11165, n11166, n11167, n11168,
    n11169, n11170, n11171, n11172, n11173, n11174,
    n11175, n11176, n11177, n11178, n11179, n11180,
    n11181, n11182, n11183, n11184, n11185, n11186,
    n11187, n11188, n11189, n11190, n11191, n11192,
    n11193, n11194, n11195, n11196, n11197, n11198,
    n11199, n11200, n11201, n11202, n11203, n11204,
    n11205, n11206, n11207, n11208, n11209, n11210,
    n11211, n11212, n11213, n11214, n11215, n11216,
    n11217, n11218, n11219, n11220, n11221, n11222,
    n11223, n11224, n11225, n11226, n11227, n11228,
    n11229, n11230, n11231, n11232, n11233, n11234,
    n11235, n11236, n11237, n11238, n11239, n11240,
    n11241, n11242, n11243, n11244, n11245, n11246,
    n11247, n11248, n11249, n11250, n11251, n11252,
    n11253, n11254, n11255, n11256, n11257, n11258,
    n11259, n11260, n11261, n11262, n11263, n11264,
    n11265, n11266, n11267, n11268, n11269, n11270,
    n11271, n11272, n11273, n11274, n11275, n11276,
    n11277, n11278, n11279, n11280, n11281, n11282,
    n11283, n11284, n11285, n11286, n11287, n11288,
    n11289, n11290, n11291, n11292, n11293, n11294,
    n11295, n11296, n11297, n11298, n11299, n11300,
    n11301, n11302, n11303, n11304, n11305, n11306,
    n11307, n11308, n11309, n11310, n11311, n11312,
    n11313, n11314, n11315, n11316, n11317, n11318,
    n11319, n11320, n11321, n11322, n11323, n11324,
    n11325, n11326, n11327, n11328, n11329, n11330,
    n11331, n11332, n11333, n11334, n11335, n11336,
    n11337, n11338, n11339, n11340, n11341, n11342,
    n11343, n11344, n11345, n11346, n11347, n11348,
    n11349, n11350, n11351, n11352, n11353, n11354,
    n11355, n11356, n11357, n11358, n11359, n11360,
    n11361, n11362, n11363, n11364, n11365, n11366,
    n11367, n11368, n11369, n11370, n11371, n11372,
    n11373, n11374, n11375, n11376, n11377, n11378,
    n11379, n11380, n11381, n11382, n11383, n11384,
    n11385, n11386, n11387, n11388, n11389, n11390,
    n11391, n11392, n11393, n11394, n11395, n11396,
    n11397, n11398, n11399, n11400, n11401, n11402,
    n11403, n11404, n11405, n11406, n11407, n11408,
    n11409, n11410, n11411, n11412, n11413, n11414,
    n11415, n11416, n11417, n11418, n11419, n11420,
    n11421, n11422, n11423, n11424, n11425, n11426,
    n11427, n11428, n11429, n11430, n11431, n11432,
    n11433, n11434, n11435, n11436, n11437, n11438,
    n11439, n11440, n11441, n11442, n11443, n11444,
    n11445, n11446, n11447, n11448, n11449, n11450,
    n11451, n11452, n11453, n11454, n11455, n11456,
    n11457, n11458, n11459, n11460, n11461, n11462,
    n11463, n11464, n11465, n11466, n11467, n11468,
    n11469, n11470, n11471, n11472, n11473, n11474,
    n11475, n11476, n11477, n11478, n11479, n11480,
    n11481, n11482, n11483, n11484, n11485, n11486,
    n11487, n11488, n11489, n11490, n11491, n11492,
    n11493, n11494, n11495, n11496, n11497, n11498,
    n11499, n11500, n11501, n11502, n11503, n11504,
    n11505, n11506, n11507, n11508, n11509, n11510,
    n11511, n11512, n11513, n11514, n11515, n11516,
    n11517, n11518, n11519, n11520, n11521, n11522,
    n11523, n11524, n11525, n11526, n11527, n11528,
    n11529, n11530, n11531, n11532, n11533, n11534,
    n11535, n11536, n11537, n11538, n11539, n11540,
    n11541, n11542, n11543, n11544, n11545, n11546,
    n11547, n11548, n11549, n11550, n11551, n11552,
    n11553, n11554, n11555, n11556, n11557, n11558,
    n11559, n11560, n11561, n11562, n11563, n11564,
    n11565, n11566, n11567, n11568, n11569, n11570,
    n11571, n11572, n11573, n11574, n11575, n11576,
    n11577, n11578, n11579, n11580, n11581, n11582,
    n11583, n11584, n11585, n11586, n11587, n11588,
    n11589, n11590, n11591, n11592, n11593, n11594,
    n11595, n11596, n11597, n11598, n11599, n11600,
    n11601, n11602, n11603, n11604, n11605, n11606,
    n11607, n11608, n11609, n11610, n11611, n11612,
    n11613, n11614, n11615, n11616, n11617, n11618,
    n11619, n11620, n11621, n11622, n11623, n11624,
    n11625, n11626, n11627, n11628, n11629, n11630,
    n11631, n11632, n11633, n11634, n11635, n11636,
    n11637, n11638, n11639, n11640, n11641, n11642,
    n11643, n11644, n11645, n11646, n11647, n11648,
    n11649, n11650, n11651, n11652, n11653, n11654,
    n11655, n11656, n11657, n11658, n11659, n11660,
    n11661, n11662, n11663, n11664, n11665, n11666,
    n11667, n11668, n11669, n11670, n11671, n11672,
    n11673, n11674, n11675, n11676, n11677, n11678,
    n11679, n11680, n11681, n11682, n11683, n11684,
    n11685, n11686, n11687, n11688, n11689, n11690,
    n11691, n11692, n11693, n11694, n11695, n11696,
    n11697, n11698, n11699, n11700, n11701, n11702,
    n11703, n11704, n11705, n11706, n11707, n11708,
    n11709, n11710, n11711, n11712, n11713, n11714,
    n11715, n11716, n11717, n11718, n11719, n11720,
    n11721, n11722, n11723, n11724, n11725, n11726,
    n11727, n11728, n11729, n11730, n11731, n11732,
    n11733, n11734, n11735, n11736, n11737, n11738,
    n11739, n11740, n11741, n11742, n11743, n11744,
    n11745, n11746, n11747, n11748, n11749, n11750,
    n11751, n11752, n11753, n11754, n11755, n11756,
    n11757, n11758, n11759, n11760, n11761, n11762,
    n11763, n11764, n11765, n11766, n11767, n11768,
    n11769, n11770, n11771, n11772, n11773, n11774,
    n11775, n11776, n11777, n11778, n11779, n11780,
    n11781, n11782, n11783, n11784, n11785, n11786,
    n11787, n11788, n11789, n11790, n11791, n11792,
    n11793, n11794, n11795, n11796, n11797, n11798,
    n11799, n11800, n11801, n11802, n11803, n11804,
    n11805, n11806, n11807, n11808, n11809, n11810,
    n11811, n11812, n11813, n11814, n11815, n11816,
    n11817, n11818, n11819, n11820, n11821, n11822,
    n11823, n11824, n11825, n11826, n11827, n11828,
    n11829, n11830, n11831, n11832, n11833, n11834,
    n11835, n11836, n11837, n11838, n11839, n11840,
    n11841, n11842, n11843, n11844, n11845, n11846,
    n11847, n11848, n11849, n11850, n11851, n11852,
    n11853, n11854, n11855, n11856, n11857, n11858,
    n11859, n11860, n11861, n11862, n11863, n11864,
    n11865, n11866, n11867, n11868, n11869, n11870,
    n11871, n11872, n11873, n11874, n11875, n11876,
    n11877, n11878, n11879, n11880, n11881, n11882,
    n11883, n11884, n11885, n11886, n11887, n11888,
    n11889, n11890, n11891, n11892, n11893, n11894,
    n11895, n11896, n11897, n11898, n11899, n11900,
    n11901, n11902, n11903, n11904, n11905, n11906,
    n11907, n11908, n11909, n11910, n11911, n11912,
    n11913, n11914, n11915, n11916, n11917, n11918,
    n11919, n11920, n11921, n11922, n11923, n11924,
    n11925, n11926, n11927, n11928, n11929, n11930,
    n11931, n11932, n11933, n11934, n11935, n11936,
    n11937, n11938, n11939, n11940, n11941, n11942,
    n11943, n11944, n11945, n11946, n11947, n11948,
    n11949, n11950, n11951, n11952, n11953, n11954,
    n11955, n11956, n11957, n11958, n11959, n11960,
    n11961, n11962, n11963, n11964, n11965, n11966,
    n11967, n11968, n11969, n11970, n11971, n11972,
    n11973, n11974, n11975, n11976, n11977, n11978,
    n11979, n11980, n11981, n11982, n11983, n11984,
    n11985, n11986, n11987, n11988, n11989, n11990,
    n11991, n11992, n11993, n11994, n11995, n11996,
    n11997, n11998, n11999, n12000, n12001, n12002,
    n12003, n12004, n12005, n12006, n12007, n12008,
    n12009, n12010, n12011, n12012, n12013, n12014,
    n12015, n12016, n12017, n12018, n12019, n12020,
    n12021, n12022, n12023, n12024, n12025, n12026,
    n12027, n12028, n12029, n12030, n12031, n12032,
    n12033, n12034, n12035, n12036, n12037, n12038,
    n12039, n12040, n12041, n12042, n12043, n12044,
    n12045, n12046, n12047, n12048, n12049, n12050,
    n12051, n12052, n12053, n12054, n12055, n12056,
    n12057, n12058, n12059, n12060, n12061, n12062,
    n12063, n12064, n12065, n12066, n12067, n12068,
    n12069, n12070, n12071, n12072, n12073, n12074,
    n12075, n12076, n12077, n12078, n12079, n12080,
    n12081, n12082, n12083, n12084, n12085, n12086,
    n12087, n12088, n12089, n12090, n12091, n12092,
    n12093, n12094, n12095, n12096, n12097, n12098,
    n12099, n12100, n12101, n12102, n12103, n12104,
    n12105, n12106, n12107, n12108, n12109, n12110,
    n12111, n12112, n12113, n12114, n12115, n12116,
    n12117, n12118, n12119, n12120, n12121, n12122,
    n12123, n12124, n12125, n12126, n12127, n12128,
    n12129, n12130, n12131, n12132, n12133, n12134,
    n12135, n12136, n12137, n12138, n12139, n12140,
    n12141, n12142, n12143, n12144, n12145, n12146,
    n12147, n12148, n12149, n12150, n12151, n12152,
    n12153, n12154, n12155, n12156, n12157, n12158,
    n12159, n12160, n12161, n12162, n12163, n12164,
    n12165, n12166, n12167, n12168, n12169, n12170,
    n12171, n12172, n12173, n12174, n12175, n12176,
    n12177, n12178, n12179, n12180, n12181, n12182,
    n12183, n12184, n12185, n12186, n12187, n12188,
    n12189, n12190, n12191, n12192, n12193, n12194,
    n12195, n12196, n12197, n12198, n12199, n12200,
    n12201, n12202, n12203, n12204, n12205, n12206,
    n12207, n12208, n12209, n12210, n12211, n12212,
    n12213, n12214, n12215, n12216, n12217, n12218,
    n12219, n12220, n12221, n12222, n12223, n12224,
    n12225, n12226, n12227, n12228, n12229, n12230,
    n12231, n12232, n12233, n12234, n12235, n12236,
    n12237, n12238, n12239, n12240, n12241, n12242,
    n12243, n12244, n12245, n12246, n12247, n12248,
    n12249, n12250, n12251, n12252, n12253, n12254,
    n12255, n12256, n12257, n12258, n12259, n12260,
    n12261, n12262, n12263, n12264, n12265, n12266,
    n12267, n12268, n12269, n12270, n12271, n12272,
    n12273, n12274, n12275, n12276, n12277, n12278,
    n12279, n12280, n12281, n12282, n12283, n12284,
    n12285, n12286, n12287, n12288, n12289, n12290,
    n12291, n12292, n12293, n12294, n12295, n12296,
    n12297, n12298, n12299, n12300, n12301, n12302,
    n12303, n12304, n12305, n12306, n12307, n12308,
    n12309, n12310, n12311, n12312, n12313, n12314,
    n12315, n12316, n12317, n12318, n12319, n12320,
    n12321, n12322, n12323, n12324, n12325, n12326,
    n12327, n12328, n12329, n12330, n12331, n12332,
    n12333, n12334, n12335, n12336, n12337, n12338,
    n12339, n12340, n12341, n12342, n12343, n12344,
    n12345, n12346, n12347, n12348, n12349, n12350,
    n12351, n12352, n12353, n12354, n12355, n12356,
    n12357, n12358, n12359, n12360, n12361, n12362,
    n12363, n12364, n12365, n12366, n12367, n12368,
    n12369, n12370, n12371, n12372, n12373, n12374,
    n12375, n12376, n12377, n12378, n12379, n12380,
    n12381, n12382, n12383, n12384, n12385, n12386,
    n12387, n12388, n12389, n12390, n12391, n12392,
    n12393, n12394, n12395, n12396, n12397, n12398,
    n12399, n12400, n12401, n12402, n12403, n12404,
    n12405, n12406, n12407, n12408, n12409, n12410,
    n12411, n12412, n12413, n12414, n12415, n12416,
    n12417, n12418, n12419, n12420, n12421, n12422,
    n12423, n12424, n12425, n12426, n12427, n12428,
    n12429, n12430, n12431, n12432, n12433, n12434,
    n12435, n12436, n12437, n12438, n12439, n12440,
    n12441, n12442, n12443, n12444, n12445, n12446,
    n12447, n12448, n12449, n12450, n12451, n12452,
    n12453, n12454, n12455, n12456, n12457, n12458,
    n12459, n12460, n12461, n12462, n12463, n12464,
    n12465, n12466, n12467, n12468, n12469, n12470,
    n12471, n12472, n12473, n12474, n12475, n12476,
    n12477, n12478, n12479, n12480, n12481, n12482,
    n12483, n12484, n12485, n12486, n12487, n12488,
    n12489, n12490, n12491, n12492, n12493, n12494,
    n12495, n12496, n12497, n12498, n12499, n12500,
    n12501, n12502, n12503, n12504, n12505, n12506,
    n12507, n12508, n12509, n12510, n12511, n12512,
    n12513, n12514, n12515, n12516, n12517, n12518,
    n12519, n12520, n12521, n12522, n12523, n12524,
    n12525, n12526, n12527, n12528, n12529, n12530,
    n12531, n12532, n12533, n12534, n12535, n12536,
    n12537, n12538, n12539, n12540, n12541, n12542,
    n12543, n12544, n12545, n12546, n12547, n12548,
    n12549, n12550, n12551, n12552, n12553, n12554,
    n12555, n12556, n12557, n12558, n12559, n12560,
    n12561, n12562, n12563, n12564, n12565, n12566,
    n12567, n12568, n12569, n12570, n12571, n12572,
    n12573, n12574, n12575, n12576, n12577, n12578,
    n12579, n12580, n12581, n12582, n12583, n12584,
    n12585, n12586, n12587, n12588, n12589, n12590,
    n12591, n12592, n12593, n12594, n12595, n12596,
    n12597, n12598, n12599, n12600, n12601, n12602,
    n12603, n12604, n12605, n12606, n12607, n12608,
    n12609, n12610, n12611, n12612, n12613, n12614,
    n12615, n12616, n12617, n12618, n12619, n12620,
    n12621, n12622, n12623, n12624, n12625, n12626,
    n12627, n12628, n12629, n12630, n12631, n12632,
    n12633, n12634, n12635, n12636, n12637, n12638,
    n12639, n12640, n12641, n12642, n12643, n12644,
    n12645, n12646, n12647, n12648, n12649, n12650,
    n12651, n12652, n12653, n12654, n12655, n12656,
    n12657, n12658, n12659, n12660, n12661, n12662,
    n12663, n12664, n12665, n12666, n12667, n12668,
    n12669, n12670, n12671, n12672, n12673, n12674,
    n12675, n12676, n12677, n12678, n12679, n12680,
    n12681, n12682, n12683, n12684, n12685, n12686,
    n12687, n12688, n12689, n12690, n12691, n12692,
    n12693, n12694, n12695, n12696, n12697, n12698,
    n12699, n12700, n12701, n12702, n12703, n12704,
    n12705, n12706, n12707, n12708, n12709, n12710,
    n12711, n12712, n12713, n12714, n12715, n12716,
    n12717, n12718, n12719, n12720, n12721, n12722,
    n12723, n12724, n12725, n12726, n12727, n12728,
    n12729, n12730, n12731, n12732, n12733, n12734,
    n12735, n12736, n12737, n12738, n12739, n12740,
    n12741, n12742, n12743, n12744, n12745, n12746,
    n12747, n12748, n12749, n12750, n12751, n12752,
    n12753, n12754, n12755, n12756, n12757, n12758,
    n12759, n12760, n12761, n12762, n12763, n12764,
    n12765, n12766, n12767, n12768, n12769, n12770,
    n12771, n12772, n12773, n12774, n12775, n12776,
    n12777, n12778, n12779, n12780, n12781, n12782,
    n12783, n12784, n12785, n12786, n12787, n12788,
    n12789, n12790, n12791, n12792, n12793, n12794,
    n12795, n12796, n12797, n12798, n12799, n12800,
    n12801, n12802, n12803, n12804, n12805, n12806,
    n12807, n12808, n12809, n12810, n12811, n12812,
    n12813, n12814, n12815, n12816, n12817, n12818,
    n12819, n12820, n12821, n12822, n12823, n12824,
    n12825, n12826, n12827, n12828, n12829, n12830,
    n12831, n12832, n12833, n12834, n12835, n12836,
    n12837, n12838, n12839, n12840, n12841, n12842,
    n12843, n12844, n12845, n12846, n12847, n12848,
    n12849, n12850, n12851, n12852, n12853, n12854,
    n12855, n12856, n12857, n12858, n12859, n12860,
    n12861, n12862, n12863, n12864, n12865, n12866,
    n12867, n12868, n12869, n12870, n12871, n12872,
    n12873, n12874, n12875, n12876, n12877, n12878,
    n12879, n12880, n12881, n12882, n12883, n12884,
    n12885, n12886, n12887, n12888, n12889, n12890,
    n12891, n12892, n12893, n12894, n12895, n12896,
    n12897, n12898, n12899, n12900, n12901, n12902,
    n12903, n12904, n12905, n12906, n12907, n12908,
    n12909, n12910, n12911, n12912, n12913, n12914,
    n12915, n12916, n12917, n12918, n12919, n12920,
    n12921, n12922, n12923, n12924, n12925, n12926,
    n12927, n12928, n12929, n12930, n12931, n12932,
    n12933, n12934, n12935, n12936, n12937, n12938,
    n12939, n12940, n12941, n12942, n12943, n12944,
    n12945, n12946, n12947, n12948, n12949, n12950,
    n12951, n12952, n12953, n12954, n12955, n12956,
    n12957, n12958, n12959, n12960, n12961, n12962,
    n12963, n12964, n12965, n12966, n12967, n12968,
    n12969, n12970, n12971, n12972, n12973, n12974,
    n12975, n12976, n12977, n12978, n12979, n12980,
    n12981, n12982, n12983, n12984, n12985, n12986,
    n12987, n12988, n12989, n12990, n12991, n12992,
    n12993, n12994, n12995, n12996, n12997, n12998,
    n12999, n13000, n13001, n13002, n13003, n13004,
    n13005, n13006, n13007, n13008, n13009, n13010,
    n13011, n13012, n13013, n13014, n13015, n13016,
    n13017, n13018, n13019, n13020, n13021, n13022,
    n13023, n13024, n13025, n13026, n13027, n13028,
    n13029, n13030, n13031, n13032, n13033, n13034,
    n13035, n13036, n13037, n13038, n13039, n13040,
    n13041, n13042, n13043, n13044, n13045, n13046,
    n13047, n13048, n13049, n13050, n13051, n13052,
    n13053, n13054, n13055, n13056, n13057, n13058,
    n13059, n13060, n13061, n13062, n13063, n13064,
    n13065, n13066, n13067, n13068, n13069, n13070,
    n13071, n13072, n13073, n13074, n13075, n13076,
    n13077, n13078, n13079, n13080, n13081, n13082,
    n13083, n13084, n13085, n13086, n13087, n13088,
    n13089, n13090, n13091, n13092, n13093, n13094,
    n13095, n13096, n13097, n13098, n13099, n13100,
    n13101, n13102, n13103, n13104, n13105, n13106,
    n13107, n13108, n13109, n13110, n13111, n13112,
    n13113, n13114, n13115, n13116, n13117, n13118,
    n13119, n13120, n13121, n13122, n13123, n13124,
    n13125, n13126, n13127, n13128, n13129, n13130,
    n13131, n13132, n13133, n13134, n13135, n13136,
    n13137, n13138, n13139, n13140, n13141, n13142,
    n13143, n13144, n13145, n13146, n13147, n13148,
    n13149, n13150, n13151, n13152, n13153, n13154,
    n13155, n13156, n13157, n13158, n13159, n13160,
    n13161, n13162, n13163, n13164, n13165, n13166,
    n13167, n13168, n13169, n13170, n13171, n13172,
    n13173, n13174, n13175, n13176, n13177, n13178,
    n13179, n13180, n13181, n13182, n13183, n13184,
    n13185, n13186, n13187, n13188, n13189, n13190,
    n13191, n13192, n13193, n13194, n13195, n13196,
    n13197, n13198, n13199, n13200, n13201, n13202,
    n13203, n13204, n13205, n13206, n13207, n13208,
    n13209, n13210, n13211, n13212, n13213, n13214,
    n13215, n13216, n13217, n13218, n13219, n13220,
    n13221, n13222, n13223, n13224, n13225, n13226,
    n13227, n13228, n13229, n13230, n13231, n13232,
    n13233, n13234, n13235, n13236, n13237, n13238,
    n13239, n13240, n13241, n13242, n13243, n13244,
    n13245, n13246, n13247, n13248, n13249, n13250,
    n13251, n13252, n13253, n13254, n13255, n13256,
    n13257, n13258, n13259, n13260, n13261, n13262,
    n13263, n13264, n13265, n13266, n13267, n13268,
    n13269, n13270, n13271, n13272, n13273, n13274,
    n13275, n13276, n13277, n13278, n13279, n13280,
    n13281, n13282, n13283, n13284, n13285, n13286,
    n13287, n13288, n13289, n13290, n13291, n13292,
    n13293, n13294, n13295, n13296, n13297, n13298,
    n13299, n13300, n13301, n13302, n13303, n13304,
    n13305, n13306, n13307, n13308, n13309, n13310,
    n13311, n13312, n13313, n13314, n13315, n13316,
    n13317, n13318, n13319, n13320, n13321, n13322,
    n13323, n13324, n13325, n13326, n13327, n13328,
    n13329, n13330, n13331, n13332, n13333, n13334,
    n13335, n13336, n13337, n13338, n13339, n13340,
    n13341, n13342, n13343, n13344, n13345, n13346,
    n13347, n13348, n13349, n13350, n13351, n13352,
    n13353, n13354, n13355, n13356, n13357, n13358,
    n13359, n13360, n13361, n13362, n13363, n13364,
    n13365, n13366, n13367, n13368, n13369, n13370,
    n13371, n13372, n13373, n13374, n13375, n13376,
    n13377, n13378, n13379, n13380, n13381, n13382,
    n13383, n13384, n13385, n13386, n13387, n13388,
    n13389, n13390, n13391, n13392, n13393, n13394,
    n13395, n13396, n13397, n13398, n13399, n13400,
    n13401, n13402, n13403, n13404, n13405, n13406,
    n13407, n13408, n13409, n13410, n13411, n13412,
    n13413, n13414, n13415, n13416, n13417, n13418,
    n13419, n13420, n13421, n13422, n13423, n13424,
    n13425, n13426, n13427, n13428, n13429, n13430,
    n13431, n13432, n13433, n13434, n13435, n13436,
    n13437, n13438, n13439, n13440, n13441, n13442,
    n13443, n13444, n13445, n13446, n13447, n13448,
    n13449, n13450, n13451, n13452, n13453, n13454,
    n13455, n13456, n13457, n13458, n13459, n13460,
    n13461, n13462, n13463, n13464, n13465, n13466,
    n13467, n13468, n13469, n13470, n13471, n13472,
    n13473, n13474, n13475, n13476, n13477, n13478,
    n13479, n13480, n13481, n13482, n13483, n13484,
    n13485, n13486, n13487, n13488, n13489, n13490,
    n13491, n13492, n13493, n13494, n13495, n13496,
    n13497, n13498, n13499, n13500, n13501, n13502,
    n13503, n13504, n13505, n13506, n13507, n13508,
    n13509, n13510, n13511, n13512, n13513, n13514,
    n13515, n13516, n13517, n13518, n13519, n13520,
    n13521, n13522, n13523, n13524, n13525, n13526,
    n13527, n13528, n13529, n13530, n13531, n13532,
    n13533, n13534, n13535, n13536, n13537, n13538,
    n13539, n13540, n13541, n13542, n13543, n13544,
    n13545, n13546, n13547, n13548, n13549, n13550,
    n13551, n13552, n13553, n13554, n13555, n13556,
    n13557, n13558, n13559, n13560, n13561, n13562,
    n13563, n13564, n13565, n13566, n13567, n13568,
    n13569, n13570, n13571, n13572, n13573, n13574,
    n13575, n13576, n13577, n13578, n13579, n13580,
    n13581, n13582, n13583, n13584, n13585, n13586,
    n13587, n13588, n13589, n13590, n13591, n13592,
    n13593, n13594, n13595, n13596, n13597, n13598,
    n13599, n13600, n13601, n13602, n13603, n13604,
    n13605, n13606, n13607, n13608, n13609, n13610,
    n13611, n13612, n13613, n13614, n13615, n13616,
    n13617, n13618, n13619, n13620, n13621, n13622,
    n13623, n13624, n13625, n13626, n13627, n13628,
    n13629, n13630, n13631, n13632, n13633, n13634,
    n13635, n13636, n13637, n13638, n13639, n13640,
    n13641, n13642, n13643, n13644, n13645, n13646,
    n13647, n13648, n13649, n13650, n13651, n13652,
    n13653, n13654, n13655, n13656, n13657, n13658,
    n13659, n13660, n13661, n13662, n13663, n13664,
    n13665, n13666, n13667, n13668, n13669, n13670,
    n13671, n13672, n13673, n13674, n13675, n13676,
    n13677, n13678, n13679, n13680, n13681, n13682,
    n13683, n13684, n13685, n13686, n13687, n13688,
    n13689, n13690, n13691, n13692, n13693, n13694,
    n13695, n13696, n13697, n13698, n13699, n13700,
    n13701, n13702, n13703, n13704, n13705, n13706,
    n13707, n13708, n13709, n13710, n13711, n13712,
    n13713, n13714, n13715, n13716, n13717, n13718,
    n13719, n13720, n13721, n13722, n13723, n13724,
    n13725, n13726, n13727, n13728, n13729, n13730,
    n13731, n13732, n13733, n13734, n13735, n13736,
    n13737, n13738, n13739, n13740, n13741, n13742,
    n13743, n13744, n13745, n13746, n13747, n13748,
    n13749, n13750, n13751, n13752, n13753, n13754,
    n13755, n13756, n13757, n13758, n13759, n13760,
    n13761, n13762, n13763, n13764, n13765, n13766,
    n13767, n13768, n13769, n13770, n13771, n13772,
    n13773, n13774, n13775, n13776, n13777, n13778,
    n13779, n13780, n13781, n13782, n13783, n13784,
    n13785, n13786, n13787, n13788, n13789, n13790,
    n13791, n13792, n13793, n13794, n13795, n13796,
    n13797, n13798, n13799, n13800, n13801, n13802,
    n13803, n13804, n13805, n13806, n13807, n13808,
    n13809, n13810, n13811, n13812, n13813, n13814,
    n13815, n13816, n13817, n13818, n13819, n13820,
    n13821, n13822, n13823, n13824, n13825, n13826,
    n13827, n13828, n13829, n13830, n13831, n13832,
    n13833, n13834, n13835, n13836, n13837, n13838,
    n13839, n13840, n13841, n13842, n13843, n13844,
    n13845, n13846, n13847, n13848, n13849, n13850,
    n13851, n13852, n13853, n13854, n13855, n13856,
    n13857, n13858, n13859, n13860, n13861, n13862,
    n13863, n13864, n13865, n13866, n13867, n13868,
    n13869, n13870, n13871, n13872, n13873, n13874,
    n13875, n13876, n13877, n13878, n13879, n13880,
    n13881, n13882, n13883, n13884, n13885, n13886,
    n13887, n13888, n13889, n13890, n13891, n13892,
    n13893, n13894, n13895, n13896, n13897, n13898,
    n13899, n13900, n13901, n13902, n13903, n13904,
    n13905, n13906, n13907, n13908, n13909, n13910,
    n13911, n13912, n13913, n13914, n13915, n13916,
    n13917, n13918, n13919, n13920, n13921, n13922,
    n13923, n13924, n13925, n13926, n13927, n13928,
    n13929, n13930, n13931, n13932, n13933, n13934,
    n13935, n13936, n13937, n13938, n13939, n13940,
    n13941, n13942, n13943, n13944, n13945, n13946,
    n13947, n13948, n13949, n13950, n13951, n13952,
    n13953, n13954, n13955, n13956, n13957, n13958,
    n13959, n13960, n13961, n13962, n13963, n13964,
    n13965, n13966, n13967, n13968, n13969, n13970,
    n13971, n13972, n13973, n13974, n13975, n13976,
    n13977, n13978, n13979, n13980, n13981, n13982,
    n13983, n13984, n13985, n13986, n13987, n13988,
    n13989, n13990, n13991, n13992, n13993, n13994,
    n13995, n13996, n13997, n13998, n13999, n14000,
    n14001, n14002, n14003, n14004, n14005, n14006,
    n14007, n14008, n14009, n14010, n14011, n14012,
    n14013, n14014, n14015, n14016, n14017, n14018,
    n14019, n14020, n14021, n14022, n14023, n14024,
    n14025, n14026, n14027, n14028, n14029, n14030,
    n14031, n14032, n14033, n14034, n14035, n14036,
    n14037, n14038, n14039, n14040, n14041, n14042,
    n14043, n14044, n14045, n14046, n14047, n14048,
    n14049, n14050, n14051, n14052, n14053, n14054,
    n14055, n14056, n14057, n14058, n14059, n14060,
    n14061, n14062, n14063, n14064, n14065, n14066,
    n14067, n14068, n14069, n14070, n14071, n14072,
    n14073, n14074, n14075, n14076, n14077, n14078,
    n14079, n14080, n14081, n14082, n14083, n14084,
    n14085, n14086, n14087, n14088, n14089, n14090,
    n14091, n14092, n14093, n14094, n14095, n14096,
    n14097, n14098, n14099, n14100, n14101, n14102,
    n14103, n14104, n14105, n14106, n14107, n14108,
    n14109, n14110, n14111, n14112, n14113, n14114,
    n14115, n14116, n14117, n14118, n14119, n14120,
    n14121, n14122, n14123, n14124, n14125, n14126,
    n14127, n14128, n14129, n14130, n14131, n14132,
    n14133, n14134, n14135, n14136, n14137, n14138,
    n14139, n14140, n14141, n14142, n14143, n14144,
    n14145, n14146, n14147, n14148, n14149, n14150,
    n14151, n14152, n14153, n14154, n14155, n14156,
    n14157, n14158, n14159, n14160, n14161, n14162,
    n14163, n14164, n14165, n14166, n14167, n14168,
    n14169, n14170, n14171, n14172, n14173, n14174,
    n14175, n14176, n14177, n14178, n14179, n14180,
    n14181, n14182, n14183, n14184, n14185, n14186,
    n14187, n14188, n14189, n14190, n14191, n14192,
    n14193, n14194, n14195, n14196, n14197, n14198,
    n14199, n14200, n14201, n14202, n14203, n14204,
    n14205, n14206, n14207, n14208, n14209, n14210,
    n14211, n14212, n14213, n14214, n14215, n14216,
    n14217, n14218, n14219, n14220, n14221, n14222,
    n14223, n14224, n14225, n14226, n14227, n14228,
    n14229, n14230, n14231, n14232, n14233, n14234,
    n14235, n14236, n14237, n14238, n14239, n14240,
    n14241, n14242, n14243, n14244, n14245, n14246,
    n14247, n14248, n14249, n14250, n14251, n14252,
    n14253, n14254, n14255, n14256, n14257, n14258,
    n14259, n14260, n14261, n14262, n14263, n14264,
    n14265, n14266, n14267, n14268, n14269, n14270,
    n14271, n14272, n14273, n14274, n14275, n14276,
    n14277, n14278, n14279, n14280, n14281, n14282,
    n14283, n14284, n14285, n14286, n14287, n14288,
    n14289, n14290, n14291, n14292, n14293, n14294,
    n14295, n14296, n14297, n14298, n14299, n14300,
    n14301, n14302, n14303, n14304, n14305, n14306,
    n14307, n14308, n14309, n14310, n14311, n14312,
    n14313, n14314, n14315, n14316, n14317, n14318,
    n14319, n14320, n14321, n14322, n14323, n14324,
    n14325, n14326, n14327, n14328, n14329, n14330,
    n14331, n14332, n14333, n14334, n14335, n14336,
    n14337, n14338, n14339, n14340, n14341, n14342,
    n14343, n14344, n14345, n14346, n14347, n14348,
    n14349, n14350, n14351, n14352, n14353, n14354,
    n14355, n14356, n14357, n14358, n14359, n14360,
    n14361, n14362, n14363, n14364, n14365, n14366,
    n14367, n14368, n14369, n14370, n14371, n14372,
    n14373, n14374, n14375, n14376, n14377, n14378,
    n14379, n14380, n14381, n14382, n14383, n14384,
    n14385, n14386, n14387, n14388, n14389, n14390,
    n14391, n14392, n14393, n14394, n14395, n14396,
    n14397, n14398, n14399, n14400, n14401, n14402,
    n14403, n14404, n14405, n14406, n14407, n14408,
    n14409, n14410, n14411, n14412, n14413, n14414,
    n14415, n14416, n14417, n14418, n14419, n14420,
    n14421, n14422, n14423, n14424, n14425, n14426,
    n14427, n14428, n14429, n14430, n14431, n14432,
    n14433, n14434, n14435, n14436, n14437, n14438,
    n14439, n14440, n14441, n14442, n14443, n14444,
    n14445, n14446, n14447, n14448, n14449, n14450,
    n14451, n14452, n14453, n14454, n14455, n14456,
    n14457, n14458, n14459, n14460, n14461, n14462,
    n14463, n14464, n14465, n14466, n14467, n14468,
    n14469, n14470, n14471, n14472, n14473, n14474,
    n14475, n14476, n14477, n14478, n14479, n14480,
    n14481, n14482, n14483, n14484, n14485, n14486,
    n14487, n14488, n14489, n14490, n14491, n14492,
    n14493, n14494, n14495, n14496, n14497, n14498,
    n14499, n14500, n14501, n14502, n14503, n14504,
    n14505, n14506, n14507, n14508, n14509, n14510,
    n14511, n14512, n14513, n14514, n14515, n14516,
    n14517, n14518, n14519, n14520, n14521, n14522,
    n14523, n14524, n14525, n14526, n14527, n14528,
    n14529, n14530, n14531, n14532, n14533, n14534,
    n14535, n14536, n14537, n14538, n14539, n14540,
    n14541, n14542, n14543, n14544, n14545, n14546,
    n14547, n14548, n14549, n14550, n14551, n14552,
    n14553, n14554, n14555, n14556, n14557, n14558,
    n14559, n14560, n14561, n14562, n14563, n14564,
    n14565, n14566, n14567, n14568, n14569, n14570,
    n14571, n14572, n14573, n14574, n14575, n14576,
    n14577, n14578, n14579, n14580, n14581, n14582,
    n14583, n14584, n14585, n14586, n14587, n14588,
    n14589, n14590, n14591, n14592, n14593, n14594,
    n14595, n14596, n14597, n14598, n14599, n14600,
    n14601, n14602, n14603, n14604, n14605, n14606,
    n14607, n14608, n14609, n14610, n14611, n14612,
    n14613, n14614, n14615, n14616, n14617, n14618,
    n14619, n14620, n14621, n14622, n14623, n14624,
    n14625, n14626, n14627, n14628, n14629, n14630,
    n14631, n14632, n14633, n14634, n14635, n14636,
    n14637, n14638, n14639, n14640, n14641, n14642,
    n14643, n14644, n14645, n14646, n14647, n14648,
    n14649, n14650, n14651, n14652, n14653, n14654,
    n14655, n14656, n14657, n14658, n14659, n14660,
    n14661, n14662, n14663, n14664, n14665, n14666,
    n14667, n14668, n14669, n14670, n14671, n14672,
    n14673, n14674, n14675, n14676, n14677, n14678,
    n14679, n14680, n14681, n14682, n14683, n14684,
    n14685, n14686, n14687, n14688, n14689, n14690,
    n14691, n14692, n14693, n14694, n14695, n14696,
    n14697, n14698, n14699, n14700, n14701, n14702,
    n14703, n14704, n14705, n14706, n14707, n14708,
    n14709, n14710, n14711, n14712, n14713, n14714,
    n14715, n14716, n14717, n14718, n14719, n14720,
    n14721, n14722, n14723, n14724, n14725, n14726,
    n14727, n14728, n14729, n14730, n14731, n14732,
    n14733, n14734, n14735, n14736, n14737, n14738,
    n14739, n14740, n14741, n14742, n14743, n14744,
    n14745, n14746, n14747, n14748, n14749, n14750,
    n14751, n14752, n14753, n14754, n14755, n14756,
    n14757, n14758, n14759, n14760, n14761, n14762,
    n14763, n14764, n14765, n14766, n14767, n14768,
    n14769, n14770, n14771, n14772, n14773, n14774,
    n14775, n14776, n14777, n14778, n14779, n14780,
    n14781, n14782, n14783, n14784, n14785, n14786,
    n14787, n14788, n14789, n14790, n14791, n14792,
    n14793, n14794, n14795, n14796, n14797, n14798,
    n14799, n14800, n14801, n14802, n14803, n14804,
    n14805, n14806, n14807, n14808, n14809, n14810,
    n14811, n14812, n14813, n14814, n14815, n14816,
    n14817, n14818, n14819, n14820, n14821, n14822,
    n14823, n14824, n14825, n14826, n14827, n14828,
    n14829, n14830, n14831, n14832, n14833, n14834,
    n14835, n14836, n14837, n14838, n14839, n14840,
    n14841, n14842, n14843, n14844, n14845, n14846,
    n14847, n14848, n14849, n14850, n14851, n14852,
    n14853, n14854, n14855, n14856, n14857, n14858,
    n14859, n14860, n14861, n14862, n14863, n14864,
    n14865, n14866, n14867, n14868, n14869, n14870,
    n14871, n14872, n14873, n14874, n14875, n14876,
    n14877, n14878, n14879, n14880, n14881, n14882,
    n14883, n14884, n14885, n14886, n14887, n14888,
    n14889, n14890, n14891, n14892, n14893, n14894,
    n14895, n14896, n14897, n14898, n14899, n14900,
    n14901, n14902, n14903, n14904, n14905, n14906,
    n14907, n14908, n14909, n14910, n14911, n14912,
    n14913, n14914, n14915, n14916, n14917, n14918,
    n14919, n14920, n14921, n14922, n14923, n14924,
    n14925, n14926, n14927, n14928, n14929, n14930,
    n14931, n14932, n14933, n14934, n14935, n14936,
    n14937, n14938, n14939, n14940, n14941, n14942,
    n14943, n14944, n14945, n14946, n14947, n14948,
    n14949, n14950, n14951, n14952, n14953, n14954,
    n14955, n14956, n14957, n14958, n14959, n14960,
    n14961, n14962, n14963, n14964, n14965, n14966,
    n14967, n14968, n14969, n14970, n14971, n14972,
    n14973, n14974, n14975, n14976, n14977, n14978,
    n14979, n14980, n14981, n14982, n14983, n14984,
    n14985, n14986, n14987, n14988, n14989, n14990,
    n14991, n14992, n14993, n14994, n14995, n14996,
    n14997, n14998, n14999, n15000, n15001, n15002,
    n15003, n15004, n15005, n15006, n15007, n15008,
    n15009, n15010, n15011, n15012, n15013, n15014,
    n15015, n15016, n15017, n15018, n15019, n15020,
    n15021, n15022, n15023, n15024, n15025, n15026,
    n15027, n15028, n15029, n15030, n15031, n15032,
    n15033, n15034, n15035, n15036, n15037, n15038,
    n15039, n15040, n15041, n15042, n15043, n15044,
    n15045, n15046, n15047, n15048, n15049, n15050,
    n15051, n15052, n15053, n15054, n15055, n15056,
    n15057, n15058, n15059, n15060, n15061, n15062,
    n15063, n15064, n15065, n15066, n15067, n15068,
    n15069, n15070, n15071, n15072, n15073, n15074,
    n15075, n15076, n15077, n15078, n15079, n15080,
    n15081, n15082, n15083, n15084, n15085, n15086,
    n15087, n15088, n15089, n15090, n15091, n15092,
    n15093, n15094, n15095, n15096, n15097, n15098,
    n15099, n15100, n15101, n15102, n15103, n15104,
    n15105, n15106, n15107, n15108, n15109, n15110,
    n15111, n15112, n15113, n15114, n15115, n15116,
    n15117, n15118, n15119, n15120, n15121, n15122,
    n15123, n15124, n15125, n15126, n15127, n15128,
    n15129, n15130, n15131, n15132, n15133, n15134,
    n15135, n15136, n15137, n15138, n15139, n15140,
    n15141, n15142, n15143, n15144, n15145, n15146,
    n15147, n15148, n15149, n15150, n15151, n15152,
    n15153, n15154, n15155, n15156, n15157, n15158,
    n15159, n15160, n15161, n15162, n15163, n15164,
    n15165, n15166, n15167, n15168, n15169, n15170,
    n15171, n15172, n15173, n15174, n15175, n15176,
    n15177, n15178, n15179, n15180, n15181, n15182,
    n15183, n15184, n15185, n15186, n15187, n15188,
    n15189, n15190, n15191, n15192, n15193, n15194,
    n15195, n15196, n15197, n15198, n15199, n15200,
    n15201, n15202, n15203, n15204, n15205, n15206,
    n15207, n15208, n15209, n15210, n15211, n15212,
    n15213, n15214, n15215, n15216, n15217, n15218,
    n15219, n15220, n15221, n15222, n15223, n15224,
    n15225, n15226, n15227, n15228, n15229, n15230,
    n15231, n15232, n15233, n15234, n15235, n15236,
    n15237, n15238, n15239, n15240, n15241, n15242,
    n15243, n15244, n15245, n15246, n15247, n15248,
    n15249, n15250, n15251, n15252, n15253, n15254,
    n15255, n15256, n15257, n15258, n15259, n15260,
    n15261, n15262, n15263, n15264, n15265, n15266,
    n15267, n15268, n15269, n15270, n15271, n15272,
    n15273, n15274, n15275, n15276, n15277, n15278,
    n15279, n15280, n15281, n15282, n15283, n15284,
    n15285, n15286, n15287, n15288, n15289, n15290,
    n15291, n15292, n15293, n15294, n15295, n15296,
    n15297, n15298, n15299, n15300, n15301, n15302,
    n15303, n15304, n15305, n15306, n15307, n15308,
    n15309, n15310, n15311, n15312, n15313, n15314,
    n15315, n15316, n15317, n15318, n15319, n15320,
    n15321, n15322, n15323, n15324, n15325, n15326,
    n15327, n15328, n15329, n15330, n15331, n15332,
    n15333, n15334, n15335, n15336, n15337, n15338,
    n15339, n15340, n15341, n15342, n15343, n15344,
    n15345, n15346, n15347, n15348, n15349, n15350,
    n15351, n15352, n15353, n15354, n15355, n15356,
    n15357, n15358, n15359, n15360, n15361, n15362,
    n15363, n15364, n15365, n15366, n15367, n15368,
    n15369, n15370, n15371, n15372, n15373, n15374,
    n15375, n15376, n15377, n15378, n15379, n15380,
    n15381, n15382, n15383, n15384, n15385, n15386,
    n15387, n15388, n15389, n15390, n15391, n15392,
    n15393, n15394, n15395, n15396, n15397, n15398,
    n15399, n15400, n15401, n15402, n15403, n15404,
    n15405, n15406, n15407, n15408, n15409, n15410,
    n15411, n15412, n15413, n15414, n15415, n15416,
    n15417, n15418, n15419, n15420, n15421, n15422,
    n15423, n15424, n15425, n15426, n15427, n15428,
    n15429, n15430, n15431, n15432, n15433, n15434,
    n15435, n15436, n15437, n15438, n15439, n15440,
    n15441, n15442, n15443, n15444, n15445, n15446,
    n15447, n15448, n15449, n15450, n15451, n15452,
    n15453, n15454, n15455, n15456, n15457, n15458,
    n15459, n15460, n15461, n15462, n15463, n15464,
    n15465, n15466, n15467, n15468, n15469, n15470,
    n15471, n15472, n15473, n15474, n15475, n15476,
    n15477, n15478, n15479, n15480, n15481, n15482,
    n15483, n15484, n15485, n15486, n15487, n15488,
    n15489, n15490, n15491, n15492, n15493, n15494,
    n15495, n15496, n15497, n15498, n15499, n15500,
    n15501, n15502, n15503, n15504, n15505, n15506,
    n15507, n15508, n15509, n15510, n15511, n15512,
    n15513, n15514, n15515, n15516, n15517, n15518,
    n15519, n15520, n15521, n15522, n15523, n15524,
    n15525, n15526, n15527, n15528, n15529, n15530,
    n15531, n15532, n15533, n15534, n15535, n15536,
    n15537, n15538, n15539, n15540, n15541, n15542,
    n15543, n15544, n15545, n15546, n15547, n15548,
    n15549, n15550, n15551, n15552, n15553, n15554,
    n15555, n15556, n15557, n15558, n15559, n15560,
    n15561, n15562, n15563, n15564, n15565, n15566,
    n15567, n15568, n15569, n15570, n15571, n15572,
    n15573, n15574, n15575, n15576, n15577, n15578,
    n15579, n15580, n15581, n15582, n15583, n15584,
    n15585, n15586, n15587, n15588, n15589, n15590,
    n15591, n15592, n15593, n15594, n15595, n15596,
    n15597, n15598, n15599, n15600, n15601, n15602,
    n15603, n15604, n15605, n15606, n15607, n15608,
    n15609, n15610, n15611, n15612, n15613, n15614,
    n15615, n15616, n15617, n15618, n15619, n15620,
    n15621, n15622, n15623, n15624, n15625, n15626,
    n15627, n15628, n15629, n15630, n15631, n15632,
    n15633, n15634, n15635, n15636, n15637, n15638,
    n15639, n15640, n15641, n15642, n15643, n15644,
    n15645, n15646, n15647, n15648, n15649, n15650,
    n15651, n15652, n15653, n15654, n15655, n15656,
    n15657, n15658, n15659, n15660, n15661, n15662,
    n15663, n15664, n15665, n15666, n15667, n15668,
    n15669, n15670, n15671, n15672, n15673, n15674,
    n15675, n15676, n15677, n15678, n15679, n15680,
    n15681, n15682, n15683, n15684, n15685, n15686,
    n15687, n15688, n15689, n15690, n15691, n15692,
    n15693, n15694, n15695, n15696, n15697, n15698,
    n15699, n15700, n15701, n15702, n15703, n15704,
    n15705, n15706, n15707, n15708, n15709, n15710,
    n15711, n15712, n15713, n15714, n15715, n15716,
    n15717, n15718, n15719, n15720, n15721, n15722,
    n15723, n15724, n15725, n15726, n15727, n15728,
    n15729, n15730, n15731, n15732, n15733, n15734,
    n15735, n15736, n15737, n15738, n15739, n15740,
    n15741, n15742, n15743, n15744, n15745, n15746,
    n15747, n15748, n15749, n15750, n15751, n15752,
    n15753, n15754, n15755, n15756, n15757, n15758,
    n15759, n15760, n15761, n15762, n15763, n15764,
    n15765, n15766, n15767, n15768, n15769, n15770,
    n15771, n15772, n15773, n15774, n15775, n15776,
    n15777, n15778, n15779, n15780, n15781, n15782,
    n15783, n15784, n15785, n15786, n15787, n15788,
    n15789, n15790, n15791, n15792, n15793, n15794,
    n15795, n15796, n15797, n15798, n15799, n15800,
    n15801, n15802, n15803, n15804, n15805, n15806,
    n15807, n15808, n15809, n15810, n15811, n15812,
    n15813, n15814, n15815, n15816, n15817, n15818,
    n15819, n15820, n15821, n15822, n15823, n15824,
    n15825, n15826, n15827, n15828, n15829, n15830,
    n15831, n15832, n15833, n15834, n15835, n15836,
    n15837, n15838, n15839, n15840, n15841, n15842,
    n15843, n15844, n15845, n15846, n15847, n15848,
    n15849, n15850, n15851, n15852, n15853, n15854,
    n15855, n15856, n15857, n15858, n15859, n15860,
    n15861, n15862, n15863, n15864, n15865, n15866,
    n15867, n15868, n15869, n15870, n15871, n15872,
    n15873, n15874, n15875, n15876, n15877, n15878,
    n15879, n15880, n15881, n15882, n15883, n15884,
    n15885, n15886, n15887, n15888, n15889, n15890,
    n15891, n15892, n15893, n15894, n15895, n15896,
    n15897, n15898, n15899, n15900, n15901, n15902,
    n15903, n15904, n15905, n15906, n15907, n15908,
    n15909, n15910, n15911, n15912, n15913, n15914,
    n15915, n15916, n15917, n15918, n15919, n15920,
    n15921, n15922, n15923, n15924, n15925, n15926,
    n15927, n15928, n15929, n15930, n15931, n15932,
    n15933, n15934, n15935, n15936, n15937, n15938,
    n15939, n15940, n15941, n15942, n15943, n15944,
    n15945, n15946, n15947, n15948, n15949, n15950,
    n15951, n15952, n15953, n15954, n15955, n15956,
    n15957, n15958, n15959, n15960, n15961, n15962,
    n15963, n15964, n15965, n15966, n15967, n15968,
    n15969, n15970, n15971, n15972, n15973, n15974,
    n15975, n15976, n15977, n15978, n15979, n15980,
    n15981, n15982, n15983, n15984, n15985, n15986,
    n15987, n15988, n15989, n15990, n15991, n15992,
    n15993, n15994, n15995, n15996, n15997, n15998,
    n15999, n16000, n16001, n16002, n16003, n16004,
    n16005, n16006, n16007, n16008, n16009, n16010,
    n16011, n16012, n16013, n16014, n16015, n16016,
    n16017, n16018, n16019, n16020, n16021, n16022,
    n16023, n16024, n16025, n16026, n16027, n16028,
    n16029, n16030, n16031, n16032, n16033, n16034,
    n16035, n16036, n16037, n16038, n16039, n16040,
    n16041, n16042, n16043, n16044, n16045, n16046,
    n16047, n16048, n16049, n16050, n16051, n16052,
    n16053, n16054, n16055, n16056, n16057, n16058,
    n16059, n16060, n16061, n16062, n16063, n16064,
    n16065, n16066, n16067, n16068, n16069, n16070,
    n16071, n16072, n16073, n16074, n16075, n16076,
    n16077, n16078, n16079, n16080, n16081, n16082,
    n16083, n16084, n16085, n16086, n16087, n16088,
    n16089, n16090, n16091, n16092, n16093, n16094,
    n16095, n16096, n16097, n16098, n16099, n16100,
    n16101, n16102, n16103, n16104, n16105, n16106,
    n16107, n16108, n16109, n16110, n16111, n16112,
    n16113, n16114, n16115, n16116, n16117, n16118,
    n16119, n16120, n16121, n16122, n16123, n16124,
    n16125, n16126, n16127, n16128, n16129, n16130,
    n16131, n16132, n16133, n16134, n16135, n16136,
    n16137, n16138, n16139, n16140, n16141, n16142,
    n16143, n16144, n16145, n16146, n16147, n16148,
    n16149, n16150, n16151, n16152, n16153, n16154,
    n16155, n16156, n16157, n16158, n16159, n16160,
    n16161, n16162, n16163, n16164, n16165, n16166,
    n16167, n16168, n16169, n16170, n16171, n16172,
    n16173, n16174, n16175, n16176, n16177, n16178,
    n16179, n16180, n16181, n16182, n16183, n16184,
    n16185, n16186, n16187, n16188, n16189, n16190,
    n16191, n16192, n16193, n16194, n16195, n16196,
    n16197, n16198, n16199, n16200, n16201, n16202,
    n16203, n16204, n16205, n16206, n16207, n16208,
    n16209, n16210, n16211, n16212, n16213, n16214,
    n16215, n16216, n16217, n16218, n16219, n16220,
    n16221, n16222, n16223, n16224, n16225, n16226,
    n16227, n16228, n16229, n16230, n16231, n16232,
    n16233, n16234, n16235, n16236, n16237, n16238,
    n16239, n16240, n16241, n16242, n16243, n16244,
    n16245, n16246, n16247, n16248, n16249, n16250,
    n16251, n16252, n16253, n16254, n16255, n16256,
    n16257, n16258, n16259, n16260, n16261, n16262,
    n16263, n16264, n16265, n16266, n16267, n16268,
    n16269, n16270, n16271, n16272, n16273, n16274,
    n16275, n16276, n16277, n16278, n16279, n16280,
    n16281, n16282, n16283, n16284, n16285, n16286,
    n16287, n16288, n16289, n16290, n16291, n16292,
    n16293, n16294, n16295, n16296, n16297, n16298,
    n16299, n16300, n16301, n16302, n16303, n16304,
    n16305, n16306, n16307, n16308, n16309, n16310,
    n16311, n16312, n16313, n16314, n16315, n16316,
    n16317, n16318, n16319, n16320, n16321, n16322,
    n16323, n16324, n16325, n16326, n16327, n16328,
    n16329, n16330, n16331, n16332, n16333, n16334,
    n16335, n16336, n16337, n16338, n16339, n16340,
    n16341, n16342, n16343, n16344, n16345, n16346,
    n16347, n16348, n16349, n16350, n16351, n16352,
    n16353, n16354, n16355, n16356, n16357, n16358,
    n16359, n16360, n16361, n16362, n16363, n16364,
    n16365, n16366, n16367, n16368, n16369, n16370,
    n16371, n16372, n16373, n16374, n16375, n16376,
    n16377, n16378, n16379, n16380, n16381, n16382,
    n16383, n16384, n16385, n16386, n16387, n16388,
    n16389, n16390, n16391, n16392, n16393, n16394,
    n16395, n16396, n16397, n16398, n16399, n16400,
    n16401, n16402, n16403, n16404, n16405, n16406,
    n16407, n16408, n16409, n16410, n16411, n16412,
    n16413, n16414, n16415, n16416, n16417, n16418,
    n16419, n16420, n16421, n16422, n16423, n16424,
    n16425, n16426, n16427, n16428, n16429, n16430,
    n16431, n16432, n16433, n16434, n16435, n16436,
    n16437, n16438, n16439, n16440, n16441, n16442,
    n16443, n16444, n16445, n16446, n16447, n16448,
    n16449, n16450, n16451, n16452, n16453, n16454,
    n16455, n16456, n16457, n16458, n16459, n16460,
    n16461, n16462, n16463, n16464, n16465, n16466,
    n16467, n16468, n16469, n16470, n16471, n16472,
    n16473, n16474, n16475, n16476, n16477, n16478,
    n16479, n16480, n16481, n16482, n16483, n16484,
    n16485, n16486, n16487, n16488, n16489, n16490,
    n16491, n16492, n16493, n16494, n16495, n16496,
    n16497, n16498, n16499, n16500, n16501, n16502,
    n16503, n16504, n16505, n16506, n16507, n16508,
    n16509, n16510, n16511, n16512, n16513, n16514,
    n16515, n16516, n16517, n16518, n16519, n16520,
    n16521, n16522, n16523, n16524, n16525, n16526,
    n16527, n16528, n16529, n16530, n16531, n16532,
    n16533, n16534, n16535, n16536, n16537, n16538,
    n16539, n16540, n16541, n16542, n16543, n16544,
    n16545, n16546, n16547, n16548, n16549, n16550,
    n16551, n16552, n16553, n16554, n16555, n16556,
    n16557, n16558, n16559, n16560, n16561, n16562,
    n16563, n16564, n16565, n16566, n16567, n16568,
    n16569, n16570, n16571, n16572, n16573, n16574,
    n16575, n16576, n16577, n16578, n16579, n16580,
    n16581, n16582, n16583, n16584, n16585, n16586,
    n16587, n16588, n16589, n16590, n16591, n16592,
    n16593, n16594, n16595, n16596, n16597, n16598,
    n16599, n16600, n16601, n16602, n16603, n16604,
    n16605, n16606, n16607, n16608, n16609, n16610,
    n16611, n16612, n16613, n16614, n16615, n16616,
    n16617, n16618, n16619, n16620, n16621, n16622,
    n16623, n16624, n16625, n16626, n16627, n16628,
    n16629, n16630, n16631, n16632, n16633, n16634,
    n16635, n16636, n16637, n16638, n16639, n16640,
    n16641, n16642, n16643, n16644, n16645, n16646,
    n16647, n16648, n16649, n16650, n16651, n16652,
    n16653, n16654, n16655, n16656, n16657, n16658,
    n16659, n16660, n16661, n16662, n16663, n16664,
    n16665, n16666, n16667, n16668, n16669, n16670,
    n16671, n16672, n16673, n16674, n16675, n16676,
    n16677, n16678, n16679, n16680, n16681, n16682,
    n16683, n16684, n16685, n16686, n16687, n16688,
    n16689, n16690, n16691, n16692, n16693, n16694,
    n16695, n16696, n16697, n16698, n16699, n16700,
    n16701, n16702, n16703, n16704, n16705, n16706,
    n16707, n16708, n16709, n16710, n16711, n16712,
    n16713, n16714, n16715, n16716, n16717, n16718,
    n16719, n16720, n16721, n16722, n16723, n16724,
    n16725, n16726, n16727, n16728, n16729, n16730,
    n16731, n16732, n16733, n16734, n16735, n16736,
    n16737, n16738, n16739, n16740, n16741, n16742,
    n16743, n16744, n16745, n16746, n16747, n16748,
    n16749, n16750, n16751, n16752, n16753, n16754,
    n16755, n16756, n16757, n16758, n16759, n16760,
    n16761, n16762, n16763, n16764, n16765, n16766,
    n16767, n16768, n16769, n16770, n16771, n16772,
    n16773, n16774, n16775, n16776, n16777, n16778,
    n16779, n16780, n16781, n16782, n16783, n16784,
    n16785, n16786, n16787, n16788, n16789, n16790,
    n16791, n16792, n16793, n16794, n16795, n16796,
    n16797, n16798, n16799, n16800, n16801, n16802,
    n16803, n16804, n16805, n16806, n16807, n16808,
    n16809, n16810, n16811, n16812, n16813, n16814,
    n16815, n16816, n16817, n16818, n16819, n16820,
    n16821, n16822, n16823, n16824, n16825, n16826,
    n16827, n16828, n16829, n16830, n16831, n16832,
    n16833, n16834, n16835, n16836, n16837, n16838,
    n16839, n16840, n16841, n16842, n16843, n16844,
    n16845, n16846, n16847, n16848, n16849, n16850,
    n16851, n16852, n16853, n16854, n16855, n16856,
    n16857, n16858, n16859, n16860, n16861, n16862,
    n16863, n16864, n16865, n16866, n16867, n16868,
    n16869, n16870, n16871, n16872, n16873, n16874,
    n16875, n16876, n16877, n16878, n16879, n16880,
    n16881, n16882, n16883, n16884, n16885, n16886,
    n16887, n16888, n16889, n16890, n16891, n16892,
    n16893, n16894, n16895, n16896, n16897, n16898,
    n16899, n16900, n16901, n16902, n16903, n16904,
    n16905, n16906, n16907, n16908, n16909, n16910,
    n16911, n16912, n16913, n16914, n16915, n16916,
    n16917, n16918, n16919, n16920, n16921, n16922,
    n16923, n16924, n16925, n16926, n16927, n16928,
    n16929, n16930, n16931, n16932, n16933, n16934,
    n16935, n16936, n16937, n16938, n16939, n16940,
    n16941, n16942, n16943, n16944, n16945, n16946,
    n16947, n16948, n16949, n16950, n16951, n16952,
    n16953, n16954, n16955, n16956, n16957, n16958,
    n16959, n16960, n16961, n16962, n16963, n16964,
    n16965, n16966, n16967, n16968, n16969, n16970,
    n16971, n16972, n16973, n16974, n16975, n16976,
    n16977, n16978, n16979, n16980, n16981, n16982,
    n16983, n16984, n16985, n16986, n16987, n16988,
    n16989, n16990, n16991, n16992, n16993, n16994,
    n16995, n16996, n16997, n16998, n16999, n17000,
    n17001, n17002, n17003, n17004, n17005, n17006,
    n17007, n17008, n17009, n17010, n17011, n17012,
    n17013, n17014, n17015, n17016, n17017, n17018,
    n17019, n17020, n17021, n17022, n17023, n17024,
    n17025, n17026, n17027, n17028, n17029, n17030,
    n17031, n17032, n17033, n17034, n17035, n17036,
    n17037, n17038, n17039, n17040, n17041, n17042,
    n17043, n17044, n17045, n17046, n17047, n17048,
    n17049, n17050, n17051, n17052, n17053, n17054,
    n17055, n17056, n17057, n17058, n17059, n17060,
    n17061, n17062, n17063, n17064, n17065, n17066,
    n17067, n17068, n17069, n17070, n17071, n17072,
    n17073, n17074, n17075, n17076, n17077, n17078,
    n17079, n17080, n17081, n17082, n17083, n17084,
    n17085, n17086, n17087, n17088, n17089, n17090,
    n17091, n17092, n17093, n17094, n17095, n17096,
    n17097, n17098, n17099, n17100, n17101, n17102,
    n17103, n17104, n17105, n17106, n17107, n17108,
    n17109, n17110, n17111, n17112, n17113, n17114,
    n17115, n17116, n17117, n17118, n17119, n17120,
    n17121, n17122, n17123, n17124, n17125, n17126,
    n17127, n17128, n17129, n17130, n17131, n17132,
    n17133, n17134, n17135, n17136, n17137, n17138,
    n17139, n17140, n17141, n17142, n17143, n17144,
    n17145, n17146, n17147, n17148, n17149, n17150,
    n17151, n17152, n17153, n17154, n17155, n17156,
    n17157, n17158, n17159, n17160, n17161, n17162,
    n17163, n17164, n17165, n17166, n17167, n17168,
    n17169, n17170, n17171, n17172, n17173, n17174,
    n17175, n17176, n17177, n17178, n17179, n17180,
    n17181, n17182, n17183, n17184, n17185, n17186,
    n17187, n17188, n17189, n17190, n17191, n17192,
    n17193, n17194, n17195, n17196, n17197, n17198,
    n17199, n17200, n17201, n17202, n17203, n17204,
    n17205, n17206, n17207, n17208, n17209, n17210,
    n17211, n17212, n17213, n17214, n17215, n17216,
    n17217, n17218, n17219, n17220, n17221, n17222,
    n17223, n17224, n17225, n17226, n17227, n17228,
    n17229, n17230, n17231, n17232, n17233, n17234,
    n17235, n17236, n17237, n17238, n17239, n17240,
    n17241, n17242, n17243, n17244, n17245, n17246,
    n17247, n17248, n17249, n17250, n17251, n17252,
    n17253, n17254, n17255, n17256, n17257, n17258,
    n17259, n17260, n17261, n17262, n17263, n17264,
    n17265, n17266, n17267, n17268, n17269, n17270,
    n17271, n17272, n17273, n17274, n17275, n17276,
    n17277, n17278, n17279, n17280, n17281, n17282,
    n17283, n17284, n17285, n17286, n17287, n17288,
    n17289, n17290, n17291, n17292, n17293, n17294,
    n17295, n17296, n17297, n17298, n17299, n17300,
    n17301, n17302, n17303, n17304, n17305, n17306,
    n17307, n17308, n17309, n17310, n17311, n17312,
    n17313, n17314, n17315, n17316, n17317, n17318,
    n17319, n17320, n17321, n17322, n17323, n17324,
    n17325, n17326, n17327, n17328, n17329, n17330,
    n17331, n17332, n17333, n17334, n17335, n17336,
    n17337, n17338, n17339, n17340, n17341, n17342,
    n17343, n17344, n17345, n17346, n17347, n17348,
    n17349, n17350, n17351, n17352, n17353, n17354,
    n17355, n17356, n17357, n17358, n17359, n17360,
    n17361, n17362, n17363, n17364, n17365, n17366,
    n17367, n17368, n17369, n17370, n17371, n17372,
    n17373, n17374, n17375, n17376, n17377, n17378,
    n17379, n17380, n17381, n17382, n17383, n17384,
    n17385, n17386, n17387, n17388, n17389, n17390,
    n17391, n17392, n17393, n17394, n17395, n17396,
    n17397, n17398, n17399, n17400, n17401, n17402,
    n17403, n17404, n17405, n17406, n17407, n17408,
    n17409, n17410, n17411, n17412, n17413, n17414,
    n17415, n17416, n17417, n17418, n17419, n17420,
    n17421, n17422, n17423, n17424, n17425, n17426,
    n17427, n17428, n17429, n17430, n17431, n17432,
    n17433, n17434, n17435, n17436, n17437, n17438,
    n17439, n17440, n17441, n17442, n17443, n17444,
    n17445, n17446, n17447, n17448, n17449, n17450,
    n17451, n17452, n17453, n17454, n17455, n17456,
    n17457, n17458, n17459, n17460, n17461, n17462,
    n17463, n17464, n17465, n17466, n17467, n17468,
    n17469, n17470, n17471, n17472, n17473, n17474,
    n17475, n17476, n17477, n17478, n17479, n17480,
    n17481, n17482, n17483, n17484, n17485, n17486,
    n17487, n17488, n17489, n17490, n17491, n17492,
    n17493, n17494, n17495, n17496, n17497, n17498,
    n17499, n17500, n17501, n17502, n17503, n17504,
    n17505, n17506, n17507, n17508, n17509, n17510,
    n17511, n17512, n17513, n17514, n17515, n17516,
    n17517, n17518, n17519, n17520, n17521, n17522,
    n17523, n17524, n17525, n17526, n17527, n17528,
    n17529, n17530, n17531, n17532, n17533, n17534,
    n17535, n17536, n17537, n17538, n17539, n17540,
    n17541, n17542, n17543, n17544, n17545, n17546,
    n17547, n17548, n17549, n17550, n17551, n17552,
    n17553, n17554, n17555, n17556, n17557, n17558,
    n17559, n17560, n17561, n17562, n17563, n17564,
    n17565, n17566, n17567, n17568, n17569, n17570,
    n17571, n17572, n17573, n17574, n17575, n17576,
    n17577, n17578, n17579, n17580, n17581, n17582,
    n17583, n17584, n17585, n17586, n17587, n17588,
    n17589, n17590, n17591, n17592, n17593, n17594,
    n17595, n17596, n17597, n17598, n17599, n17600,
    n17601, n17602, n17603, n17604, n17605, n17606,
    n17607, n17608, n17609, n17610, n17611, n17612,
    n17613, n17614, n17615, n17616, n17617, n17618,
    n17619, n17620, n17621, n17622, n17623, n17624,
    n17625, n17626, n17627, n17628, n17629, n17630,
    n17631, n17632, n17633, n17634, n17635, n17636,
    n17637, n17638, n17639, n17640, n17641, n17642,
    n17643, n17644, n17645, n17646, n17647, n17648,
    n17649, n17650, n17651, n17652, n17653, n17654,
    n17655, n17656, n17657, n17658, n17659, n17660,
    n17661, n17662, n17663, n17664, n17665, n17666,
    n17667, n17668, n17669, n17670, n17671, n17672,
    n17673, n17674, n17675, n17676, n17677, n17678,
    n17679, n17680, n17681, n17682, n17683, n17684,
    n17685, n17686, n17687, n17688, n17689, n17690,
    n17691, n17692, n17693, n17694, n17695, n17696,
    n17698, n17699, n17700, n17701, n17702, n17703,
    n17704, n17705, n17706, n17707, n17708, n17709,
    n17710, n17711, n17712, n17713, n17714, n17715,
    n17716, n17717, n17718, n17719, n17720, n17721,
    n17722, n17723, n17724, n17725, n17726, n17727,
    n17728, n17729, n17730, n17731, n17732, n17733,
    n17734, n17735, n17736, n17737, n17738, n17739,
    n17740, n17741, n17742, n17743, n17744, n17745,
    n17746, n17747, n17748, n17749, n17750, n17751,
    n17752, n17753, n17754, n17755, n17756, n17757,
    n17758, n17759, n17760, n17761, n17762, n17763,
    n17764, n17765, n17766, n17767, n17768, n17769,
    n17770, n17771, n17772, n17773, n17774, n17775,
    n17776, n17777, n17778, n17779, n17780, n17781,
    n17782, n17783, n17784, n17785, n17786, n17787,
    n17788, n17789, n17790, n17791, n17792, n17793,
    n17794, n17795, n17796, n17797, n17798, n17799,
    n17800, n17801, n17802, n17803, n17804, n17805,
    n17806, n17807, n17808, n17809, n17810, n17811,
    n17812, n17813, n17814, n17815, n17816, n17817,
    n17818, n17819, n17820, n17821, n17822, n17823,
    n17824, n17825, n17826, n17827, n17828, n17829,
    n17830, n17831, n17832, n17833, n17834, n17835,
    n17836, n17837, n17838, n17839, n17840, n17841,
    n17842, n17843, n17844, n17845, n17846, n17847,
    n17848, n17849, n17850, n17851, n17852, n17853,
    n17854, n17855, n17856, n17857, n17858, n17859,
    n17860, n17861, n17862, n17863, n17864, n17865,
    n17866, n17867, n17868, n17869, n17870, n17871,
    n17872, n17873, n17874, n17875, n17876, n17877,
    n17878, n17879, n17880, n17881, n17882, n17883,
    n17884, n17885, n17886, n17887, n17888, n17889,
    n17890, n17891, n17892, n17893, n17894, n17895,
    n17896, n17897, n17898, n17899, n17900, n17901,
    n17902, n17903, n17904, n17905, n17906, n17907,
    n17908, n17909, n17910, n17911, n17912, n17913,
    n17914, n17915, n17916, n17917, n17918, n17919,
    n17920, n17921, n17922, n17923, n17924, n17925,
    n17926, n17927, n17928, n17929, n17930, n17931,
    n17932, n17933, n17934, n17935, n17936, n17937,
    n17938, n17939, n17940, n17941, n17942, n17943,
    n17944, n17945, n17946, n17947, n17948, n17949,
    n17950, n17951, n17952, n17953, n17954, n17955,
    n17956, n17957, n17958, n17959, n17960, n17961,
    n17962, n17963, n17964, n17965, n17966, n17967,
    n17968, n17969, n17970, n17971, n17972, n17973,
    n17974, n17975, n17976, n17977, n17978, n17979,
    n17980, n17981, n17982, n17983, n17984, n17985,
    n17986, n17987, n17988, n17989, n17990, n17991,
    n17992, n17993, n17994, n17995, n17996, n17997,
    n17998, n17999, n18000, n18001, n18002, n18003,
    n18004, n18005, n18006, n18007, n18008, n18009,
    n18010, n18011, n18012, n18013, n18014, n18015,
    n18016, n18017, n18018, n18019, n18020, n18021,
    n18022, n18023, n18024, n18025, n18026, n18027,
    n18028, n18029, n18030, n18031, n18032, n18033,
    n18034, n18035, n18036, n18037, n18038, n18039,
    n18040, n18041, n18042, n18043, n18044, n18045,
    n18046, n18047, n18048, n18049, n18050, n18051,
    n18052, n18053, n18054, n18055, n18056, n18057,
    n18058, n18059, n18060, n18061, n18062, n18063,
    n18064, n18065, n18066, n18067, n18068, n18069,
    n18070, n18071, n18072, n18073, n18074, n18075,
    n18076, n18077, n18078, n18079, n18080, n18081,
    n18082, n18083, n18084, n18085, n18086, n18087,
    n18088, n18089, n18090, n18091, n18092, n18093,
    n18094, n18095, n18096, n18097, n18098, n18099,
    n18100, n18101, n18102, n18103, n18104, n18105,
    n18106, n18107, n18108, n18109, n18110, n18111,
    n18112, n18113, n18114, n18115, n18116, n18117,
    n18118, n18119, n18120, n18121, n18122, n18123,
    n18124, n18125, n18126, n18127, n18128, n18129,
    n18130, n18131, n18132, n18133, n18134, n18135,
    n18136, n18137, n18138, n18139, n18140, n18141,
    n18142, n18143, n18144, n18145, n18146, n18147,
    n18148, n18149, n18150, n18151, n18152, n18153,
    n18154, n18155, n18156, n18157, n18158, n18159,
    n18160, n18161, n18162, n18163, n18164, n18165,
    n18166, n18167, n18168, n18169, n18170, n18171,
    n18172, n18173, n18174, n18175, n18176, n18177,
    n18178, n18179, n18180, n18181, n18182, n18183,
    n18184, n18185, n18186, n18187, n18188, n18189,
    n18190, n18191, n18192, n18193, n18194, n18195,
    n18196, n18197, n18198, n18199, n18200, n18201,
    n18202, n18203, n18204, n18205, n18206, n18207,
    n18208, n18209, n18210, n18211, n18212, n18213,
    n18214, n18215, n18216, n18217, n18218, n18219,
    n18220, n18221, n18222, n18223, n18224, n18225,
    n18226, n18227, n18228, n18229, n18230, n18231,
    n18232, n18233, n18234, n18235, n18236, n18237,
    n18238, n18239, n18240, n18241, n18242, n18243,
    n18244, n18245, n18246, n18247, n18248, n18249,
    n18250, n18251, n18252, n18253, n18254, n18255,
    n18256, n18257, n18258, n18259, n18260, n18261,
    n18262, n18263, n18264, n18265, n18266, n18267,
    n18268, n18269, n18270, n18271, n18272, n18273,
    n18274, n18275, n18276, n18277, n18278, n18279,
    n18280, n18281, n18282, n18283, n18284, n18285,
    n18286, n18287, n18288, n18289, n18290, n18291,
    n18292, n18293, n18294, n18295, n18296, n18297,
    n18298, n18299, n18300, n18301, n18302, n18303,
    n18304, n18305, n18306, n18307, n18308, n18309,
    n18310, n18311, n18312, n18313, n18314, n18315,
    n18316, n18317, n18318, n18319, n18320, n18321,
    n18322, n18323, n18324, n18325, n18326, n18327,
    n18328, n18329, n18330, n18331, n18332, n18333,
    n18334, n18335, n18336, n18337, n18338, n18339,
    n18340, n18341, n18342, n18343, n18344, n18345,
    n18346, n18347, n18348, n18349, n18350, n18351,
    n18352, n18353, n18354, n18355, n18356, n18357,
    n18358, n18359, n18360, n18361, n18362, n18363,
    n18364, n18365, n18366, n18367, n18368, n18369,
    n18370, n18371, n18372, n18373, n18374, n18375,
    n18376, n18377, n18378, n18379, n18380, n18381,
    n18382, n18383, n18384, n18385, n18386, n18387,
    n18388, n18389, n18390, n18391, n18392, n18393,
    n18394, n18395, n18396, n18397, n18398, n18399,
    n18400, n18401, n18402, n18403, n18404, n18405,
    n18406, n18407, n18408, n18409, n18410, n18411,
    n18412, n18413, n18414, n18415, n18416, n18417,
    n18418, n18419, n18420, n18421, n18422, n18423,
    n18424, n18425, n18426, n18427, n18428, n18429,
    n18430, n18431, n18432, n18433, n18434, n18435,
    n18436, n18437, n18438, n18439, n18440, n18441,
    n18442, n18443, n18444, n18445, n18446, n18447,
    n18448, n18449, n18450, n18451, n18452, n18453,
    n18454, n18455, n18456, n18457, n18458, n18459,
    n18460, n18461, n18462, n18463, n18464, n18465,
    n18466, n18467, n18468, n18469, n18470, n18471,
    n18472, n18473, n18474, n18475, n18476, n18477,
    n18478, n18479, n18480, n18481, n18482, n18483,
    n18484, n18485, n18486, n18487, n18488, n18489,
    n18490, n18491, n18492, n18493, n18494, n18495,
    n18496, n18497, n18498, n18499, n18500, n18501,
    n18502, n18503, n18504, n18505, n18506, n18507,
    n18508, n18509, n18510, n18511, n18512, n18513,
    n18514, n18515, n18516, n18517, n18518, n18519,
    n18520, n18521, n18522, n18523, n18524, n18525,
    n18526, n18527, n18528, n18529, n18530, n18531,
    n18532, n18533, n18534, n18535, n18536, n18537,
    n18538, n18539, n18540, n18541, n18542, n18543,
    n18544, n18545, n18546, n18547, n18548, n18549,
    n18550, n18551, n18552, n18553, n18554, n18555,
    n18556, n18557, n18558, n18559, n18560, n18561,
    n18562, n18563, n18564, n18565, n18566, n18567,
    n18568, n18569, n18570, n18571, n18572, n18573,
    n18574, n18575, n18576, n18577, n18578, n18579,
    n18580, n18581, n18582, n18583, n18584, n18585,
    n18586, n18587, n18588, n18589, n18590, n18591,
    n18592, n18593, n18594, n18595, n18596, n18597,
    n18598, n18599, n18600, n18601, n18602, n18603,
    n18604, n18605, n18606, n18607, n18608, n18609,
    n18610, n18611, n18612, n18613, n18614, n18615,
    n18616, n18617, n18618, n18619, n18620, n18621,
    n18622, n18623, n18624, n18625, n18626, n18627,
    n18628, n18629, n18630, n18631, n18632, n18633,
    n18634, n18635, n18636, n18637, n18638, n18639,
    n18640, n18641, n18642, n18643, n18644, n18645,
    n18646, n18647, n18648, n18649, n18650, n18651,
    n18652, n18653, n18654, n18655, n18656, n18657,
    n18658, n18659, n18660, n18661, n18662, n18663,
    n18664, n18665, n18666, n18667, n18668, n18669,
    n18670, n18672, n18673, n18674, n18675, n18676,
    n18677, n18678, n18679, n18680, n18681, n18682,
    n18683, n18684, n18685, n18686, n18687, n18688,
    n18689, n18690, n18691, n18692, n18693, n18694,
    n18695, n18696, n18697, n18698, n18699, n18700,
    n18701, n18702, n18703, n18704, n18705, n18706,
    n18707, n18708, n18709, n18710, n18711, n18712,
    n18713, n18714, n18715, n18716, n18717, n18718,
    n18719, n18720, n18721, n18722, n18723, n18724,
    n18725, n18726, n18727, n18728, n18729, n18730,
    n18731, n18732, n18733, n18734, n18735, n18736,
    n18737, n18738, n18739, n18740, n18741, n18742,
    n18743, n18744, n18745, n18746, n18747, n18748,
    n18749, n18750, n18751, n18752, n18753, n18754,
    n18755, n18756, n18757, n18758, n18759, n18760,
    n18761, n18762, n18763, n18764, n18765, n18766,
    n18767, n18768, n18769, n18770, n18771, n18772,
    n18773, n18774, n18775, n18776, n18777, n18778,
    n18779, n18780, n18781, n18782, n18783, n18784,
    n18785, n18786, n18787, n18788, n18789, n18790,
    n18791, n18792, n18793, n18794, n18795, n18796,
    n18797, n18798, n18799, n18800, n18801, n18802,
    n18803, n18804, n18805, n18806, n18807, n18808,
    n18809, n18810, n18811, n18812, n18813, n18814,
    n18815, n18816, n18817, n18818, n18819, n18820,
    n18821, n18822, n18823, n18824, n18825, n18826,
    n18827, n18828, n18829, n18830, n18831, n18832,
    n18833, n18834, n18835, n18836, n18837, n18838,
    n18839, n18840, n18841, n18842, n18843, n18844,
    n18845, n18846, n18847, n18848, n18849, n18850,
    n18851, n18852, n18853, n18854, n18855, n18856,
    n18857, n18858, n18859, n18860, n18861, n18862,
    n18863, n18864, n18865, n18866, n18867, n18868,
    n18869, n18870, n18871, n18872, n18873, n18874,
    n18875, n18876, n18877, n18878, n18879, n18880,
    n18881, n18882, n18883, n18884, n18885, n18886,
    n18887, n18888, n18889, n18890, n18891, n18892,
    n18893, n18894, n18895, n18896, n18897, n18898,
    n18899, n18900, n18901, n18902, n18903, n18904,
    n18905, n18906, n18907, n18908, n18909, n18910,
    n18911, n18912, n18913, n18914, n18915, n18916,
    n18917, n18918, n18919, n18920, n18921, n18922,
    n18923, n18924, n18925, n18926, n18927, n18928,
    n18929, n18930, n18931, n18932, n18933, n18934,
    n18935, n18936, n18937, n18938, n18939, n18940,
    n18941, n18942, n18943, n18944, n18945, n18946,
    n18947, n18948, n18949, n18950, n18951, n18952,
    n18953, n18954, n18955, n18956, n18957, n18958,
    n18959, n18960, n18961, n18962, n18963, n18964,
    n18965, n18966, n18967, n18968, n18969, n18970,
    n18971, n18972, n18973, n18974, n18975, n18976,
    n18977, n18978, n18979, n18980, n18981, n18982,
    n18983, n18984, n18985, n18986, n18987, n18988,
    n18989, n18990, n18991, n18992, n18993, n18994,
    n18995, n18996, n18997, n18998, n18999, n19000,
    n19001, n19002, n19003, n19004, n19005, n19006,
    n19007, n19008, n19009, n19010, n19011, n19012,
    n19013, n19014, n19015, n19016, n19017, n19018,
    n19019, n19020, n19021, n19022, n19023, n19024,
    n19025, n19026, n19027, n19028, n19029, n19030,
    n19031, n19032, n19033, n19034, n19035, n19036,
    n19037, n19038, n19039, n19040, n19041, n19042,
    n19043, n19044, n19045, n19046, n19047, n19048,
    n19049, n19050, n19051, n19052, n19053, n19054,
    n19055, n19056, n19057, n19058, n19059, n19060,
    n19061, n19062, n19063, n19064, n19065, n19066,
    n19067, n19068, n19069, n19070, n19071, n19072,
    n19073, n19074, n19075, n19076, n19077, n19078,
    n19079, n19080, n19081, n19082, n19083, n19084,
    n19085, n19086, n19087, n19088, n19089, n19090,
    n19091, n19092, n19093, n19094, n19095, n19096,
    n19097, n19098, n19099, n19100, n19101, n19102,
    n19103, n19104, n19105, n19106, n19107, n19108,
    n19109, n19110, n19111, n19112, n19113, n19114,
    n19115, n19116, n19117, n19118, n19119, n19120,
    n19121, n19122, n19123, n19124, n19125, n19126,
    n19127, n19128, n19129, n19130, n19131, n19132,
    n19133, n19134, n19135, n19136, n19137, n19138,
    n19139, n19140, n19141, n19142, n19143, n19144,
    n19145, n19146, n19147, n19148, n19149, n19150,
    n19151, n19152, n19153, n19154, n19155, n19156,
    n19157, n19158, n19159, n19160, n19161, n19162,
    n19163, n19164, n19165, n19166, n19167, n19168,
    n19169, n19170, n19171, n19172, n19173, n19174,
    n19175, n19176, n19177, n19178, n19179, n19180,
    n19181, n19182, n19183, n19184, n19185, n19186,
    n19187, n19188, n19189, n19190, n19191, n19192,
    n19193, n19194, n19195, n19196, n19197, n19198,
    n19199, n19200, n19201, n19202, n19203, n19204,
    n19205, n19206, n19207, n19208, n19209, n19210,
    n19211, n19212, n19213, n19214, n19215, n19216,
    n19217, n19218, n19219, n19220, n19222, n19223,
    n19224, n19225, n19226, n19227, n19228, n19229,
    n19230, n19231, n19232, n19233, n19234, n19235,
    n19236, n19237, n19238, n19239, n19240, n19241,
    n19242, n19243, n19244, n19245, n19246, n19247,
    n19248, n19249, n19250, n19251, n19252, n19253,
    n19254, n19255, n19256, n19257, n19258, n19259,
    n19260, n19261, n19262, n19263, n19264, n19265,
    n19266, n19267, n19268, n19269, n19270, n19271,
    n19272, n19273, n19274, n19275, n19276, n19277,
    n19278, n19279, n19280, n19281, n19282, n19283,
    n19284, n19285, n19286, n19287, n19288, n19289,
    n19290, n19291, n19292, n19293, n19294, n19295,
    n19296, n19297, n19298, n19299, n19300, n19301,
    n19302, n19303, n19304, n19305, n19306, n19307,
    n19308, n19309, n19310, n19311, n19312, n19313,
    n19314, n19315, n19316, n19317, n19318, n19319,
    n19320, n19321, n19322, n19323, n19324, n19325,
    n19326, n19327, n19328, n19329, n19330, n19331,
    n19332, n19333, n19334, n19335, n19336, n19337,
    n19338, n19339, n19340, n19341, n19342, n19343,
    n19344, n19345, n19346, n19347, n19348, n19349,
    n19350, n19351, n19352, n19353, n19354, n19355,
    n19356, n19357, n19358, n19359, n19360, n19361,
    n19362, n19363, n19364, n19365, n19366, n19367,
    n19368, n19369, n19370, n19371, n19372, n19373,
    n19374, n19375, n19376, n19377, n19378, n19379,
    n19380, n19381, n19382, n19383, n19384, n19385,
    n19386, n19387, n19388, n19389, n19390, n19391,
    n19392, n19393, n19394, n19395, n19396, n19397,
    n19398, n19399, n19400, n19401, n19402, n19403,
    n19404, n19405, n19406, n19407, n19408, n19409,
    n19410, n19411, n19412, n19413, n19414, n19415,
    n19416, n19417, n19418, n19419, n19420, n19421,
    n19422, n19423, n19424, n19425, n19426, n19427,
    n19428, n19429, n19430, n19431, n19432, n19433,
    n19434, n19435, n19436, n19437, n19438, n19439,
    n19440, n19441, n19442, n19443, n19444, n19445,
    n19446, n19447, n19448, n19449, n19450, n19451,
    n19452, n19453, n19454, n19455, n19456, n19457,
    n19458, n19459, n19460, n19461, n19462, n19463,
    n19464, n19465, n19466, n19467, n19468, n19469,
    n19470, n19471, n19472, n19473, n19474, n19475,
    n19476, n19477, n19478, n19479, n19480, n19481,
    n19482, n19483, n19484, n19485, n19486, n19487,
    n19488, n19489, n19490, n19491, n19492, n19493,
    n19494, n19495, n19496, n19497, n19498, n19499,
    n19500, n19501, n19502, n19503, n19504, n19505,
    n19506, n19507, n19508, n19509, n19510, n19511,
    n19512, n19513, n19514, n19515, n19516, n19517,
    n19518, n19519, n19520, n19521, n19522, n19523,
    n19524, n19525, n19526, n19527, n19528, n19529,
    n19530, n19531, n19532, n19533, n19534, n19535,
    n19536, n19537, n19538, n19539, n19540, n19541,
    n19542, n19543, n19544, n19545, n19546, n19547,
    n19548, n19549, n19550, n19551, n19552, n19553,
    n19554, n19555, n19556, n19557, n19558, n19559,
    n19560, n19561, n19562, n19563, n19564, n19565,
    n19566, n19567, n19568, n19569, n19570, n19571,
    n19572, n19573, n19574, n19575, n19576, n19577,
    n19578, n19579, n19580, n19581, n19582, n19583,
    n19584, n19585, n19586, n19587, n19588, n19589,
    n19590, n19591, n19592, n19593, n19594, n19595,
    n19596, n19597, n19598, n19599, n19600, n19601,
    n19602, n19603, n19604, n19605, n19606, n19607,
    n19608, n19609, n19610, n19611, n19612, n19613,
    n19614, n19615, n19616, n19617, n19618, n19619,
    n19620, n19621, n19622, n19623, n19624, n19625,
    n19626, n19627, n19628, n19629, n19630, n19631,
    n19632, n19633, n19634, n19635, n19636, n19637,
    n19638, n19639, n19640, n19641, n19642, n19643,
    n19644, n19645, n19646, n19647, n19648, n19649,
    n19650, n19651, n19652, n19653, n19654, n19655,
    n19656, n19657, n19658, n19659, n19660, n19661,
    n19662, n19663, n19664, n19665, n19666, n19667,
    n19668, n19669, n19670, n19671, n19672, n19673,
    n19674, n19675, n19676, n19677, n19678, n19679,
    n19680, n19681, n19682, n19683, n19684, n19685,
    n19686, n19687, n19688, n19689, n19690, n19691,
    n19692, n19693, n19694, n19695, n19696, n19697,
    n19698, n19699, n19700, n19701, n19702, n19703,
    n19704, n19705, n19706, n19707, n19708, n19709,
    n19710, n19711, n19712, n19713, n19714, n19715,
    n19716, n19717, n19718, n19719, n19720, n19721,
    n19722, n19723, n19724, n19725, n19726, n19727,
    n19728, n19729, n19730, n19731, n19732, n19733,
    n19734, n19735, n19736, n19737, n19738, n19739,
    n19740, n19741, n19742, n19743, n19744, n19745,
    n19746, n19747, n19748, n19749, n19750, n19751,
    n19752, n19753, n19754, n19755, n19756, n19757,
    n19758, n19759, n19760, n19761, n19762, n19763,
    n19764, n19765, n19766, n19767, n19768, n19769,
    n19770, n19771, n19772, n19773, n19775, n19776,
    n19777, n19778, n19779, n19780, n19781, n19782,
    n19783, n19784, n19785, n19786, n19787, n19788,
    n19789, n19790, n19791, n19792, n19793, n19794,
    n19795, n19796, n19797, n19798, n19799, n19800,
    n19801, n19802, n19803, n19804, n19805, n19806,
    n19807, n19808, n19809, n19810, n19811, n19812,
    n19813, n19814, n19815, n19816, n19817, n19818,
    n19819, n19820, n19821, n19822, n19823, n19824,
    n19825, n19826, n19827, n19828, n19829, n19830,
    n19831, n19832, n19833, n19834, n19835, n19836,
    n19837, n19838, n19839, n19840, n19841, n19842,
    n19843, n19844, n19845, n19846, n19847, n19848,
    n19849, n19850, n19851, n19852, n19853, n19854,
    n19855, n19856, n19857, n19858, n19859, n19860,
    n19861, n19862, n19863, n19864, n19865, n19866,
    n19867, n19868, n19869, n19870, n19871, n19872,
    n19873, n19874, n19875, n19876, n19877, n19878,
    n19879, n19880, n19881, n19882, n19883, n19884,
    n19885, n19886, n19887, n19888, n19889, n19890,
    n19891, n19892, n19893, n19894, n19895, n19896,
    n19897, n19898, n19899, n19900, n19901, n19902,
    n19903, n19904, n19905, n19906, n19907, n19908,
    n19909, n19910, n19911, n19912, n19913, n19914,
    n19915, n19916, n19917, n19918, n19919, n19920,
    n19921, n19922, n19923, n19924, n19925, n19926,
    n19927, n19928, n19929, n19930, n19931, n19932,
    n19933, n19934, n19935, n19936, n19937, n19938,
    n19939, n19940, n19941, n19942, n19943, n19944,
    n19945, n19946, n19947, n19948, n19949, n19950,
    n19951, n19952, n19953, n19954, n19955, n19956,
    n19957, n19958, n19959, n19960, n19961, n19962,
    n19963, n19964, n19965, n19966, n19967, n19968,
    n19969, n19970, n19971, n19972, n19973, n19974,
    n19975, n19976, n19977, n19978, n19979, n19980,
    n19981, n19982, n19983, n19984, n19985, n19986,
    n19987, n19988, n19989, n19990, n19991, n19992,
    n19993, n19994, n19995, n19996, n19997, n19998,
    n19999, n20000, n20001, n20002, n20003, n20004,
    n20005, n20006, n20007, n20008, n20009, n20010,
    n20011, n20012, n20013, n20014, n20015, n20016,
    n20017, n20018, n20019, n20020, n20021, n20022,
    n20023, n20024, n20025, n20026, n20027, n20028,
    n20029, n20030, n20031, n20032, n20033, n20034,
    n20035, n20036, n20037, n20038, n20039, n20040,
    n20041, n20042, n20043, n20044, n20045, n20046,
    n20047, n20048, n20049, n20050, n20051, n20052,
    n20053, n20054, n20055, n20056, n20057, n20058,
    n20059, n20060, n20061, n20062, n20063, n20064,
    n20065, n20066, n20067, n20068, n20069, n20070,
    n20071, n20072, n20073, n20074, n20075, n20076,
    n20077, n20078, n20079, n20080, n20081, n20082,
    n20083, n20084, n20085, n20086, n20087, n20088,
    n20089, n20090, n20091, n20092, n20093, n20094,
    n20095, n20096, n20097, n20098, n20099, n20100,
    n20101, n20102, n20103, n20104, n20105, n20106,
    n20107, n20108, n20109, n20110, n20111, n20112,
    n20113, n20114, n20115, n20116, n20117, n20118,
    n20119, n20120, n20121, n20122, n20123, n20124,
    n20125, n20126, n20127, n20128, n20129, n20130,
    n20131, n20132, n20133, n20134, n20135, n20136,
    n20137, n20138, n20139, n20140, n20141, n20142,
    n20143, n20144, n20145, n20146, n20147, n20148,
    n20149, n20150, n20151, n20152, n20153, n20154,
    n20155, n20156, n20157, n20158, n20159, n20160,
    n20161, n20162, n20163, n20164, n20165, n20166,
    n20167, n20168, n20169, n20170, n20171, n20172,
    n20173, n20174, n20175, n20176, n20177, n20178,
    n20179, n20180, n20181, n20182, n20183, n20184,
    n20185, n20186, n20187, n20188, n20189, n20190,
    n20191, n20192, n20193, n20194, n20195, n20196,
    n20197, n20198, n20199, n20200, n20201, n20202,
    n20203, n20204, n20205, n20206, n20207, n20208,
    n20209, n20210, n20211, n20212, n20213, n20214,
    n20215, n20216, n20217, n20218, n20219, n20220,
    n20221, n20222, n20223, n20224, n20225, n20226,
    n20227, n20228, n20229, n20230, n20231, n20232,
    n20233, n20234, n20235, n20236, n20237, n20238,
    n20239, n20240, n20241, n20242, n20243, n20244,
    n20245, n20246, n20247, n20248, n20249, n20250,
    n20251, n20252, n20253, n20254, n20255, n20256,
    n20257, n20258, n20259, n20260, n20261, n20262,
    n20263, n20264, n20265, n20266, n20267, n20268,
    n20269, n20270, n20271, n20272, n20273, n20274,
    n20275, n20276, n20277, n20278, n20279, n20280,
    n20281, n20282, n20283, n20284, n20285, n20286,
    n20287, n20288, n20289, n20290, n20291, n20292,
    n20293, n20294, n20295, n20296, n20297, n20298,
    n20299, n20300, n20301, n20302, n20303, n20304,
    n20305, n20306, n20307, n20308, n20310, n20311,
    n20312, n20313, n20314, n20315, n20316, n20317,
    n20318, n20319, n20320, n20321, n20322, n20323,
    n20324, n20325, n20326, n20327, n20328, n20329,
    n20330, n20331, n20332, n20333, n20334, n20335,
    n20336, n20337, n20338, n20339, n20340, n20341,
    n20342, n20343, n20344, n20345, n20346, n20347,
    n20348, n20349, n20350, n20351, n20352, n20353,
    n20354, n20355, n20356, n20357, n20358, n20359,
    n20360, n20361, n20362, n20363, n20364, n20365,
    n20366, n20367, n20368, n20369, n20370, n20371,
    n20372, n20373, n20374, n20375, n20376, n20377,
    n20378, n20379, n20380, n20381, n20382, n20383,
    n20384, n20385, n20386, n20387, n20388, n20389,
    n20390, n20391, n20392, n20393, n20394, n20395,
    n20396, n20397, n20398, n20399, n20400, n20401,
    n20402, n20403, n20404, n20405, n20406, n20407,
    n20408, n20409, n20410, n20411, n20412, n20413,
    n20414, n20415, n20416, n20417, n20418, n20419,
    n20420, n20421, n20422, n20423, n20424, n20425,
    n20426, n20427, n20428, n20429, n20430, n20431,
    n20432, n20433, n20434, n20435, n20436, n20437,
    n20438, n20439, n20440, n20441, n20442, n20443,
    n20444, n20445, n20446, n20447, n20448, n20449,
    n20450, n20451, n20452, n20453, n20454, n20455,
    n20456, n20457, n20458, n20459, n20460, n20461,
    n20462, n20463, n20464, n20465, n20466, n20467,
    n20468, n20469, n20470, n20471, n20472, n20473,
    n20474, n20475, n20476, n20477, n20478, n20479,
    n20480, n20481, n20482, n20483, n20484, n20485,
    n20486, n20487, n20488, n20489, n20490, n20491,
    n20492, n20493, n20494, n20495, n20496, n20497,
    n20498, n20499, n20500, n20501, n20502, n20503,
    n20504, n20505, n20506, n20507, n20508, n20509,
    n20510, n20511, n20512, n20513, n20514, n20515,
    n20516, n20517, n20518, n20519, n20520, n20521,
    n20522, n20523, n20524, n20525, n20526, n20527,
    n20528, n20529, n20530, n20531, n20532, n20533,
    n20534, n20535, n20536, n20537, n20538, n20539,
    n20540, n20541, n20542, n20543, n20544, n20545,
    n20546, n20547, n20548, n20549, n20550, n20551,
    n20552, n20553, n20554, n20555, n20556, n20557,
    n20558, n20559, n20560, n20561, n20562, n20563,
    n20564, n20565, n20566, n20567, n20568, n20569,
    n20570, n20571, n20572, n20573, n20574, n20575,
    n20576, n20577, n20578, n20579, n20580, n20581,
    n20582, n20583, n20584, n20585, n20586, n20587,
    n20588, n20589, n20590, n20591, n20592, n20593,
    n20594, n20595, n20596, n20597, n20598, n20599,
    n20600, n20601, n20602, n20603, n20604, n20605,
    n20606, n20607, n20608, n20609, n20610, n20611,
    n20612, n20613, n20614, n20615, n20616, n20617,
    n20618, n20619, n20620, n20621, n20622, n20623,
    n20624, n20625, n20626, n20627, n20628, n20629,
    n20630, n20631, n20632, n20633, n20634, n20635,
    n20636, n20637, n20638, n20639, n20640, n20641,
    n20642, n20643, n20644, n20645, n20646, n20647,
    n20648, n20649, n20650, n20651, n20652, n20653,
    n20654, n20655, n20656, n20657, n20658, n20659,
    n20660, n20661, n20662, n20663, n20664, n20665,
    n20666, n20667, n20668, n20669, n20670, n20671,
    n20672, n20673, n20674, n20675, n20676, n20677,
    n20678, n20679, n20680, n20681, n20682, n20683,
    n20684, n20685, n20686, n20687, n20688, n20689,
    n20690, n20691, n20692, n20693, n20694, n20695,
    n20696, n20697, n20698, n20699, n20700, n20701,
    n20702, n20703, n20704, n20705, n20706, n20707,
    n20708, n20709, n20710, n20711, n20712, n20713,
    n20714, n20715, n20716, n20717, n20718, n20719,
    n20720, n20721, n20722, n20723, n20724, n20725,
    n20726, n20727, n20728, n20729, n20730, n20731,
    n20732, n20733, n20734, n20735, n20736, n20737,
    n20738, n20739, n20740, n20741, n20742, n20743,
    n20744, n20745, n20746, n20747, n20748, n20749,
    n20750, n20751, n20752, n20753, n20754, n20755,
    n20756, n20757, n20758, n20759, n20760, n20761,
    n20762, n20763, n20764, n20765, n20766, n20767,
    n20768, n20769, n20770, n20771, n20772, n20773,
    n20774, n20775, n20776, n20777, n20778, n20779,
    n20780, n20781, n20782, n20783, n20784, n20785,
    n20786, n20787, n20788, n20789, n20790, n20791,
    n20792, n20793, n20794, n20795, n20796, n20797,
    n20798, n20799, n20800, n20801, n20802, n20803,
    n20804, n20805, n20806, n20807, n20808, n20809,
    n20810, n20811, n20812, n20813, n20814, n20815,
    n20816, n20817, n20818, n20819, n20820, n20821,
    n20822, n20823, n20824, n20825, n20826, n20827,
    n20828, n20829, n20830, n20831, n20832, n20833,
    n20834, n20835, n20836, n20837, n20838, n20839,
    n20840, n20841, n20842, n20843, n20844, n20845,
    n20846, n20847, n20848, n20849, n20850, n20851,
    n20852, n20853, n20854, n20855, n20856, n20857,
    n20858, n20859, n20860, n20861, n20862, n20863,
    n20864, n20865, n20866, n20867, n20868, n20869,
    n20870, n20871, n20872, n20874, n20875, n20876,
    n20877, n20878, n20879, n20880, n20881, n20882,
    n20883, n20884, n20885, n20886, n20887, n20888,
    n20889, n20890, n20891, n20892, n20893, n20894,
    n20895, n20896, n20897, n20898, n20899, n20900,
    n20901, n20902, n20903, n20904, n20905, n20906,
    n20907, n20908, n20909, n20910, n20911, n20912,
    n20913, n20914, n20915, n20916, n20917, n20918,
    n20919, n20920, n20921, n20922, n20923, n20924,
    n20925, n20926, n20927, n20928, n20929, n20930,
    n20931, n20932, n20933, n20934, n20935, n20936,
    n20937, n20938, n20939, n20940, n20941, n20942,
    n20943, n20944, n20945, n20946, n20947, n20948,
    n20949, n20950, n20951, n20952, n20953, n20954,
    n20955, n20956, n20957, n20958, n20959, n20960,
    n20961, n20962, n20963, n20964, n20965, n20966,
    n20967, n20968, n20969, n20970, n20971, n20972,
    n20973, n20974, n20975, n20976, n20977, n20978,
    n20979, n20980, n20981, n20982, n20983, n20984,
    n20985, n20986, n20987, n20988, n20989, n20990,
    n20991, n20992, n20993, n20994, n20995, n20996,
    n20997, n20998, n20999, n21000, n21001, n21002,
    n21003, n21004, n21005, n21006, n21007, n21008,
    n21009, n21010, n21011, n21012, n21013, n21014,
    n21015, n21016, n21017, n21018, n21019, n21020,
    n21021, n21022, n21023, n21024, n21025, n21026,
    n21027, n21028, n21029, n21030, n21031, n21032,
    n21033, n21034, n21035, n21036, n21037, n21038,
    n21039, n21040, n21041, n21042, n21043, n21044,
    n21045, n21046, n21047, n21048, n21049, n21050,
    n21051, n21052, n21053, n21054, n21055, n21056,
    n21057, n21058, n21059, n21060, n21061, n21062,
    n21063, n21064, n21065, n21066, n21067, n21068,
    n21069, n21070, n21071, n21072, n21073, n21074,
    n21075, n21076, n21077, n21078, n21079, n21080,
    n21081, n21082, n21083, n21084, n21085, n21086,
    n21087, n21088, n21089, n21090, n21091, n21092,
    n21093, n21094, n21095, n21096, n21097, n21098,
    n21099, n21100, n21101, n21102, n21103, n21104,
    n21105, n21106, n21107, n21108, n21109, n21110,
    n21111, n21112, n21113, n21114, n21115, n21116,
    n21117, n21118, n21119, n21120, n21121, n21122,
    n21123, n21124, n21125, n21126, n21127, n21128,
    n21129, n21130, n21131, n21132, n21133, n21134,
    n21135, n21136, n21137, n21138, n21139, n21140,
    n21141, n21142, n21143, n21144, n21145, n21146,
    n21147, n21148, n21149, n21150, n21151, n21152,
    n21153, n21154, n21155, n21156, n21157, n21158,
    n21159, n21160, n21161, n21162, n21163, n21164,
    n21165, n21166, n21167, n21168, n21169, n21170,
    n21171, n21172, n21173, n21174, n21175, n21176,
    n21177, n21178, n21179, n21180, n21181, n21182,
    n21183, n21184, n21185, n21186, n21187, n21188,
    n21189, n21190, n21191, n21192, n21193, n21194,
    n21195, n21196, n21197, n21198, n21199, n21200,
    n21201, n21202, n21203, n21204, n21205, n21206,
    n21207, n21208, n21209, n21210, n21211, n21212,
    n21213, n21214, n21215, n21216, n21217, n21218,
    n21219, n21220, n21221, n21222, n21223, n21224,
    n21225, n21226, n21227, n21228, n21229, n21230,
    n21231, n21232, n21233, n21234, n21235, n21236,
    n21237, n21238, n21239, n21240, n21241, n21242,
    n21243, n21244, n21245, n21246, n21247, n21248,
    n21249, n21250, n21251, n21252, n21253, n21254,
    n21255, n21256, n21257, n21258, n21259, n21260,
    n21261, n21262, n21263, n21264, n21265, n21266,
    n21267, n21268, n21269, n21270, n21271, n21272,
    n21273, n21274, n21275, n21276, n21277, n21278,
    n21279, n21280, n21281, n21282, n21283, n21284,
    n21285, n21286, n21287, n21288, n21289, n21290,
    n21291, n21292, n21293, n21294, n21295, n21296,
    n21297, n21298, n21299, n21300, n21301, n21302,
    n21303, n21304, n21305, n21306, n21307, n21308,
    n21309, n21310, n21311, n21312, n21313, n21314,
    n21315, n21316, n21317, n21318, n21319, n21320,
    n21321, n21322, n21323, n21324, n21325, n21326,
    n21327, n21328, n21329, n21330, n21331, n21332,
    n21333, n21334, n21335, n21336, n21337, n21338,
    n21339, n21340, n21341, n21342, n21343, n21344,
    n21345, n21346, n21347, n21348, n21349, n21350,
    n21351, n21352, n21353, n21354, n21355, n21356,
    n21357, n21358, n21359, n21360, n21361, n21362,
    n21363, n21364, n21365, n21366, n21367, n21368,
    n21369, n21370, n21371, n21372, n21373, n21374,
    n21375, n21376, n21377, n21378, n21379, n21380,
    n21381, n21382, n21383, n21384, n21385, n21386,
    n21387, n21388, n21389, n21390, n21391, n21392,
    n21393, n21394, n21395, n21396, n21397, n21398,
    n21399, n21400, n21401, n21402, n21403, n21404,
    n21405, n21406, n21407, n21408, n21409, n21410,
    n21411, n21412, n21413, n21414, n21415, n21416,
    n21417, n21418, n21419, n21420, n21421, n21422,
    n21424, n21425, n21426, n21427, n21428, n21429,
    n21430, n21431, n21432, n21433, n21434, n21435,
    n21436, n21437, n21438, n21439, n21440, n21441,
    n21442, n21443, n21444, n21445, n21446, n21447,
    n21448, n21449, n21450, n21451, n21452, n21453,
    n21454, n21455, n21456, n21457, n21458, n21459,
    n21460, n21461, n21462, n21463, n21464, n21465,
    n21466, n21467, n21468, n21469, n21470, n21471,
    n21472, n21473, n21474, n21475, n21476, n21477,
    n21478, n21479, n21480, n21481, n21482, n21483,
    n21484, n21485, n21486, n21487, n21488, n21489,
    n21490, n21491, n21492, n21493, n21494, n21495,
    n21496, n21497, n21498, n21499, n21500, n21501,
    n21502, n21503, n21504, n21505, n21506, n21507,
    n21508, n21509, n21510, n21511, n21512, n21513,
    n21514, n21515, n21516, n21517, n21518, n21519,
    n21520, n21521, n21522, n21523, n21524, n21525,
    n21526, n21527, n21528, n21529, n21530, n21531,
    n21532, n21533, n21534, n21535, n21536, n21537,
    n21538, n21539, n21540, n21541, n21542, n21543,
    n21544, n21545, n21546, n21547, n21548, n21549,
    n21550, n21551, n21552, n21553, n21554, n21555,
    n21556, n21557, n21558, n21559, n21560, n21561,
    n21562, n21563, n21564, n21565, n21566, n21567,
    n21568, n21569, n21570, n21571, n21572, n21573,
    n21574, n21575, n21576, n21577, n21578, n21579,
    n21580, n21581, n21582, n21583, n21584, n21585,
    n21586, n21587, n21588, n21589, n21590, n21591,
    n21592, n21593, n21594, n21595, n21596, n21597,
    n21598, n21599, n21600, n21601, n21602, n21603,
    n21604, n21605, n21606, n21607, n21608, n21609,
    n21610, n21611, n21612, n21613, n21614, n21615,
    n21616, n21617, n21618, n21619, n21620, n21621,
    n21622, n21623, n21624, n21625, n21626, n21627,
    n21628, n21629, n21630, n21631, n21632, n21633,
    n21634, n21635, n21636, n21637, n21638, n21639,
    n21640, n21641, n21642, n21643, n21644, n21645,
    n21646, n21647, n21648, n21649, n21650, n21651,
    n21652, n21653, n21654, n21655, n21656, n21657,
    n21658, n21659, n21660, n21661, n21662, n21663,
    n21664, n21665, n21666, n21667, n21668, n21669,
    n21670, n21671, n21672, n21673, n21674, n21675,
    n21676, n21677, n21678, n21679, n21680, n21681,
    n21682, n21683, n21684, n21685, n21686, n21687,
    n21688, n21689, n21690, n21691, n21692, n21693,
    n21694, n21695, n21696, n21697, n21698, n21699,
    n21700, n21701, n21702, n21703, n21704, n21705,
    n21706, n21707, n21708, n21709, n21710, n21711,
    n21712, n21713, n21714, n21715, n21716, n21717,
    n21718, n21719, n21720, n21721, n21722, n21723,
    n21724, n21725, n21726, n21727, n21728, n21729,
    n21730, n21731, n21732, n21733, n21734, n21735,
    n21736, n21737, n21738, n21739, n21740, n21741,
    n21742, n21743, n21744, n21745, n21746, n21747,
    n21748, n21749, n21750, n21751, n21752, n21753,
    n21754, n21755, n21756, n21757, n21758, n21759,
    n21760, n21761, n21762, n21763, n21764, n21765,
    n21766, n21767, n21768, n21769, n21770, n21771,
    n21772, n21773, n21774, n21775, n21776, n21777,
    n21778, n21779, n21780, n21781, n21782, n21783,
    n21784, n21785, n21786, n21787, n21788, n21789,
    n21790, n21791, n21792, n21793, n21794, n21795,
    n21796, n21797, n21798, n21799, n21800, n21801,
    n21802, n21803, n21804, n21805, n21806, n21807,
    n21808, n21809, n21810, n21811, n21812, n21813,
    n21814, n21815, n21816, n21817, n21818, n21819,
    n21820, n21821, n21822, n21823, n21824, n21825,
    n21826, n21827, n21828, n21829, n21830, n21831,
    n21832, n21833, n21834, n21835, n21836, n21837,
    n21838, n21839, n21840, n21841, n21842, n21843,
    n21844, n21845, n21846, n21847, n21848, n21849,
    n21850, n21851, n21852, n21853, n21854, n21855,
    n21856, n21857, n21858, n21859, n21860, n21861,
    n21862, n21863, n21864, n21865, n21866, n21867,
    n21868, n21869, n21870, n21871, n21872, n21873,
    n21874, n21875, n21876, n21877, n21878, n21879,
    n21880, n21881, n21882, n21883, n21884, n21885,
    n21886, n21887, n21888, n21889, n21890, n21891,
    n21892, n21893, n21894, n21895, n21896, n21897,
    n21898, n21899, n21900, n21901, n21902, n21903,
    n21904, n21905, n21906, n21907, n21908, n21909,
    n21910, n21911, n21912, n21913, n21914, n21915,
    n21916, n21917, n21918, n21919, n21920, n21921,
    n21922, n21923, n21924, n21925, n21926, n21927,
    n21928, n21929, n21930, n21931, n21932, n21933,
    n21934, n21935, n21936, n21937, n21938, n21939,
    n21940, n21941, n21942, n21943, n21944, n21945,
    n21946, n21947, n21948, n21949, n21950, n21951,
    n21952, n21953, n21954, n21955, n21956, n21957,
    n21958, n21959, n21960, n21961, n21962, n21963,
    n21964, n21966, n21967, n21968, n21969, n21970,
    n21971, n21972, n21973, n21974, n21975, n21976,
    n21977, n21978, n21979, n21980, n21981, n21982,
    n21983, n21984, n21985, n21986, n21987, n21988,
    n21989, n21990, n21991, n21992, n21993, n21994,
    n21995, n21996, n21997, n21998, n21999, n22000,
    n22001, n22002, n22003, n22004, n22005, n22006,
    n22007, n22008, n22009, n22010, n22011, n22012,
    n22013, n22014, n22015, n22016, n22017, n22018,
    n22019, n22020, n22021, n22022, n22023, n22024,
    n22025, n22026, n22027, n22028, n22029, n22030,
    n22031, n22032, n22033, n22034, n22035, n22036,
    n22037, n22038, n22039, n22040, n22041, n22042,
    n22043, n22044, n22045, n22046, n22047, n22048,
    n22049, n22050, n22051, n22052, n22053, n22054,
    n22055, n22056, n22057, n22058, n22059, n22060,
    n22061, n22062, n22063, n22064, n22065, n22066,
    n22067, n22068, n22069, n22070, n22071, n22072,
    n22073, n22074, n22075, n22076, n22077, n22078,
    n22079, n22080, n22081, n22082, n22083, n22084,
    n22085, n22086, n22087, n22088, n22089, n22090,
    n22091, n22092, n22093, n22094, n22095, n22096,
    n22097, n22098, n22099, n22100, n22101, n22102,
    n22103, n22104, n22105, n22106, n22107, n22108,
    n22109, n22110, n22111, n22112, n22113, n22114,
    n22115, n22116, n22117, n22118, n22119, n22120,
    n22121, n22122, n22123, n22124, n22125, n22126,
    n22127, n22128, n22129, n22130, n22131, n22132,
    n22133, n22134, n22135, n22136, n22137, n22138,
    n22139, n22140, n22141, n22142, n22143, n22144,
    n22145, n22146, n22147, n22148, n22149, n22150,
    n22151, n22152, n22153, n22154, n22155, n22156,
    n22157, n22158, n22159, n22160, n22161, n22162,
    n22163, n22164, n22165, n22166, n22167, n22168,
    n22169, n22170, n22171, n22172, n22173, n22174,
    n22175, n22176, n22177, n22178, n22179, n22180,
    n22181, n22182, n22183, n22184, n22185, n22186,
    n22187, n22188, n22189, n22190, n22191, n22192,
    n22193, n22194, n22195, n22196, n22197, n22198,
    n22199, n22200, n22201, n22202, n22203, n22204,
    n22205, n22206, n22207, n22208, n22209, n22210,
    n22211, n22212, n22213, n22214, n22215, n22216,
    n22217, n22218, n22219, n22220, n22221, n22222,
    n22223, n22224, n22225, n22226, n22227, n22228,
    n22229, n22230, n22231, n22232, n22233, n22234,
    n22235, n22236, n22237, n22238, n22239, n22240,
    n22241, n22242, n22243, n22244, n22245, n22246,
    n22247, n22248, n22249, n22250, n22251, n22252,
    n22253, n22254, n22255, n22256, n22257, n22258,
    n22259, n22260, n22261, n22262, n22263, n22264,
    n22265, n22266, n22267, n22268, n22269, n22270,
    n22271, n22272, n22273, n22274, n22275, n22276,
    n22277, n22278, n22279, n22280, n22281, n22282,
    n22283, n22284, n22285, n22286, n22287, n22288,
    n22289, n22290, n22291, n22292, n22293, n22294,
    n22295, n22296, n22297, n22298, n22299, n22300,
    n22301, n22302, n22303, n22304, n22305, n22306,
    n22307, n22308, n22309, n22310, n22311, n22312,
    n22313, n22314, n22315, n22316, n22317, n22318,
    n22319, n22320, n22321, n22322, n22323, n22324,
    n22325, n22326, n22327, n22328, n22329, n22330,
    n22331, n22332, n22333, n22334, n22335, n22336,
    n22337, n22338, n22339, n22340, n22341, n22342,
    n22343, n22344, n22345, n22346, n22347, n22348,
    n22349, n22350, n22351, n22352, n22353, n22354,
    n22355, n22356, n22357, n22358, n22359, n22360,
    n22361, n22362, n22363, n22364, n22365, n22366,
    n22367, n22368, n22369, n22370, n22371, n22372,
    n22373, n22374, n22375, n22376, n22377, n22378,
    n22379, n22380, n22381, n22382, n22383, n22384,
    n22385, n22386, n22387, n22388, n22389, n22390,
    n22391, n22392, n22393, n22394, n22395, n22396,
    n22397, n22398, n22399, n22400, n22401, n22402,
    n22403, n22404, n22405, n22406, n22407, n22408,
    n22409, n22410, n22411, n22412, n22413, n22414,
    n22415, n22416, n22417, n22418, n22419, n22420,
    n22421, n22422, n22423, n22424, n22425, n22426,
    n22427, n22428, n22429, n22430, n22431, n22432,
    n22433, n22434, n22435, n22436, n22437, n22438,
    n22439, n22440, n22441, n22442, n22443, n22444,
    n22445, n22446, n22447, n22448, n22449, n22450,
    n22451, n22452, n22453, n22454, n22455, n22456,
    n22457, n22459, n22460, n22461, n22462, n22463,
    n22464, n22465, n22466, n22467, n22468, n22469,
    n22470, n22471, n22472, n22473, n22474, n22475,
    n22476, n22477, n22478, n22479, n22480, n22481,
    n22482, n22483, n22484, n22485, n22486, n22487,
    n22488, n22489, n22490, n22491, n22492, n22493,
    n22494, n22495, n22496, n22497, n22498, n22499,
    n22500, n22501, n22502, n22503, n22504, n22505,
    n22506, n22507, n22508, n22509, n22510, n22511,
    n22512, n22513, n22514, n22515, n22516, n22517,
    n22518, n22519, n22520, n22521, n22522, n22523,
    n22524, n22525, n22526, n22527, n22528, n22529,
    n22530, n22531, n22532, n22533, n22534, n22535,
    n22536, n22537, n22538, n22539, n22540, n22541,
    n22542, n22543, n22544, n22545, n22546, n22547,
    n22548, n22549, n22550, n22551, n22552, n22553,
    n22554, n22555, n22556, n22557, n22558, n22559,
    n22560, n22561, n22562, n22563, n22564, n22565,
    n22566, n22567, n22568, n22569, n22570, n22571,
    n22572, n22573, n22574, n22575, n22576, n22577,
    n22578, n22579, n22580, n22581, n22582, n22583,
    n22584, n22585, n22586, n22587, n22588, n22589,
    n22590, n22591, n22592, n22593, n22594, n22595,
    n22596, n22597, n22598, n22599, n22600, n22601,
    n22602, n22603, n22604, n22605, n22606, n22607,
    n22608, n22609, n22610, n22611, n22612, n22613,
    n22614, n22615, n22616, n22617, n22618, n22619,
    n22620, n22621, n22622, n22623, n22624, n22625,
    n22626, n22627, n22628, n22629, n22630, n22631,
    n22632, n22633, n22634, n22635, n22636, n22637,
    n22638, n22639, n22640, n22641, n22642, n22643,
    n22644, n22645, n22646, n22647, n22648, n22649,
    n22650, n22651, n22652, n22653, n22654, n22655,
    n22656, n22657, n22658, n22659, n22660, n22661,
    n22662, n22663, n22664, n22665, n22666, n22667,
    n22668, n22669, n22670, n22671, n22672, n22673,
    n22674, n22675, n22676, n22677, n22678, n22679,
    n22680, n22681, n22682, n22683, n22684, n22685,
    n22686, n22687, n22688, n22689, n22690, n22691,
    n22692, n22693, n22694, n22695, n22696, n22697,
    n22698, n22699, n22700, n22701, n22702, n22703,
    n22704, n22705, n22706, n22707, n22708, n22709,
    n22710, n22711, n22712, n22713, n22714, n22715,
    n22716, n22717, n22718, n22719, n22720, n22721,
    n22722, n22723, n22724, n22725, n22726, n22727,
    n22728, n22729, n22730, n22731, n22732, n22733,
    n22734, n22735, n22736, n22737, n22738, n22739,
    n22740, n22741, n22742, n22743, n22744, n22745,
    n22746, n22747, n22748, n22749, n22750, n22751,
    n22752, n22753, n22754, n22755, n22756, n22757,
    n22758, n22759, n22760, n22761, n22762, n22763,
    n22764, n22765, n22766, n22767, n22768, n22769,
    n22770, n22771, n22772, n22773, n22774, n22775,
    n22776, n22777, n22778, n22779, n22780, n22781,
    n22782, n22783, n22784, n22785, n22786, n22787,
    n22788, n22789, n22790, n22791, n22792, n22793,
    n22794, n22795, n22796, n22797, n22798, n22799,
    n22800, n22801, n22802, n22803, n22804, n22805,
    n22806, n22807, n22808, n22809, n22810, n22811,
    n22812, n22813, n22814, n22815, n22816, n22817,
    n22818, n22819, n22820, n22821, n22822, n22823,
    n22824, n22825, n22826, n22827, n22828, n22829,
    n22830, n22831, n22832, n22833, n22834, n22835,
    n22836, n22837, n22838, n22839, n22840, n22841,
    n22842, n22843, n22844, n22845, n22846, n22847,
    n22848, n22849, n22850, n22851, n22852, n22853,
    n22854, n22855, n22856, n22857, n22858, n22859,
    n22860, n22861, n22862, n22863, n22864, n22865,
    n22866, n22867, n22868, n22869, n22870, n22871,
    n22872, n22873, n22874, n22875, n22876, n22877,
    n22878, n22879, n22880, n22881, n22882, n22883,
    n22884, n22885, n22886, n22887, n22888, n22889,
    n22890, n22891, n22892, n22893, n22894, n22895,
    n22896, n22897, n22898, n22899, n22900, n22901,
    n22902, n22903, n22904, n22905, n22906, n22907,
    n22908, n22909, n22910, n22911, n22912, n22913,
    n22914, n22915, n22916, n22917, n22918, n22919,
    n22920, n22921, n22922, n22923, n22924, n22925,
    n22926, n22927, n22928, n22929, n22930, n22931,
    n22932, n22933, n22934, n22935, n22936, n22937,
    n22938, n22939, n22940, n22941, n22942, n22943,
    n22944, n22945, n22946, n22947, n22948, n22949,
    n22950, n22951, n22952, n22953, n22954, n22955,
    n22956, n22957, n22958, n22959, n22960, n22961,
    n22962, n22963, n22964, n22965, n22966, n22967,
    n22968, n22969, n22970, n22971, n22972, n22973,
    n22974, n22975, n22976, n22977, n22978, n22979,
    n22980, n22981, n22982, n22983, n22984, n22985,
    n22986, n22987, n22988, n22989, n22990, n22991,
    n22993, n22994, n22995, n22996, n22997, n22998,
    n22999, n23000, n23001, n23002, n23003, n23004,
    n23005, n23006, n23007, n23008, n23009, n23010,
    n23011, n23012, n23013, n23014, n23015, n23016,
    n23017, n23018, n23019, n23020, n23021, n23022,
    n23023, n23024, n23025, n23026, n23027, n23028,
    n23029, n23030, n23031, n23032, n23033, n23034,
    n23035, n23036, n23037, n23038, n23039, n23040,
    n23041, n23042, n23043, n23044, n23045, n23046,
    n23047, n23048, n23049, n23050, n23051, n23052,
    n23053, n23054, n23055, n23056, n23057, n23058,
    n23059, n23060, n23061, n23062, n23063, n23064,
    n23065, n23066, n23067, n23068, n23069, n23070,
    n23071, n23072, n23073, n23074, n23075, n23076,
    n23077, n23078, n23079, n23080, n23081, n23082,
    n23083, n23084, n23085, n23086, n23087, n23088,
    n23089, n23090, n23091, n23092, n23093, n23094,
    n23095, n23096, n23097, n23098, n23099, n23100,
    n23101, n23102, n23103, n23104, n23105, n23106,
    n23107, n23108, n23109, n23110, n23111, n23112,
    n23113, n23114, n23115, n23116, n23117, n23118,
    n23119, n23120, n23121, n23122, n23123, n23124,
    n23125, n23126, n23127, n23128, n23129, n23130,
    n23131, n23132, n23133, n23134, n23135, n23136,
    n23137, n23138, n23139, n23140, n23141, n23142,
    n23143, n23144, n23145, n23146, n23147, n23148,
    n23149, n23150, n23151, n23152, n23153, n23154,
    n23155, n23156, n23157, n23158, n23159, n23160,
    n23161, n23162, n23163, n23164, n23165, n23166,
    n23167, n23168, n23169, n23170, n23171, n23172,
    n23173, n23174, n23175, n23176, n23177, n23178,
    n23179, n23180, n23181, n23182, n23183, n23184,
    n23185, n23186, n23187, n23188, n23189, n23190,
    n23191, n23192, n23193, n23194, n23195, n23196,
    n23197, n23198, n23199, n23200, n23201, n23202,
    n23203, n23204, n23205, n23206, n23207, n23208,
    n23209, n23210, n23211, n23212, n23213, n23214,
    n23215, n23216, n23217, n23218, n23219, n23220,
    n23221, n23222, n23223, n23224, n23225, n23226,
    n23227, n23228, n23229, n23230, n23231, n23232,
    n23233, n23234, n23235, n23236, n23237, n23238,
    n23239, n23240, n23241, n23242, n23243, n23244,
    n23245, n23246, n23247, n23248, n23249, n23250,
    n23251, n23252, n23253, n23254, n23255, n23256,
    n23257, n23258, n23259, n23260, n23261, n23262,
    n23263, n23264, n23265, n23266, n23267, n23268,
    n23269, n23270, n23271, n23272, n23273, n23274,
    n23275, n23276, n23277, n23278, n23279, n23280,
    n23281, n23282, n23283, n23284, n23285, n23286,
    n23287, n23288, n23289, n23290, n23291, n23292,
    n23293, n23294, n23295, n23296, n23297, n23298,
    n23299, n23300, n23301, n23302, n23303, n23304,
    n23305, n23306, n23307, n23308, n23309, n23310,
    n23311, n23312, n23313, n23314, n23315, n23316,
    n23317, n23318, n23319, n23320, n23321, n23322,
    n23323, n23324, n23325, n23326, n23327, n23328,
    n23329, n23330, n23331, n23332, n23333, n23334,
    n23335, n23336, n23337, n23338, n23339, n23340,
    n23341, n23342, n23343, n23344, n23345, n23346,
    n23347, n23348, n23349, n23350, n23351, n23352,
    n23353, n23354, n23355, n23356, n23357, n23358,
    n23359, n23360, n23361, n23362, n23363, n23364,
    n23365, n23366, n23367, n23368, n23369, n23370,
    n23371, n23372, n23373, n23374, n23375, n23376,
    n23377, n23378, n23379, n23380, n23381, n23382,
    n23383, n23384, n23385, n23386, n23387, n23388,
    n23389, n23390, n23391, n23392, n23393, n23394,
    n23395, n23396, n23397, n23398, n23399, n23400,
    n23401, n23402, n23403, n23404, n23405, n23406,
    n23407, n23408, n23409, n23410, n23411, n23412,
    n23413, n23414, n23415, n23416, n23417, n23418,
    n23419, n23420, n23421, n23422, n23423, n23424,
    n23425, n23426, n23427, n23428, n23429, n23430,
    n23431, n23432, n23433, n23434, n23435, n23436,
    n23437, n23438, n23439, n23440, n23441, n23442,
    n23443, n23444, n23445, n23446, n23447, n23448,
    n23449, n23450, n23451, n23452, n23453, n23454,
    n23455, n23456, n23457, n23458, n23459, n23460,
    n23461, n23462, n23463, n23464, n23465, n23466,
    n23467, n23468, n23469, n23470, n23471, n23472,
    n23473, n23474, n23475, n23476, n23477, n23478,
    n23479, n23480, n23481, n23482, n23483, n23484,
    n23485, n23486, n23487, n23488, n23489, n23490,
    n23491, n23492, n23493, n23494, n23495, n23496,
    n23497, n23498, n23499, n23500, n23501, n23502,
    n23503, n23504, n23505, n23506, n23507, n23508,
    n23509, n23510, n23511, n23512, n23513, n23514,
    n23515, n23516, n23517, n23518, n23519, n23520,
    n23522, n23523, n23524, n23525, n23526, n23527,
    n23528, n23529, n23530, n23531, n23532, n23533,
    n23534, n23535, n23536, n23537, n23538, n23539,
    n23540, n23541, n23542, n23543, n23544, n23545,
    n23546, n23547, n23548, n23549, n23550, n23551,
    n23552, n23553, n23554, n23555, n23556, n23557,
    n23558, n23559, n23560, n23561, n23562, n23563,
    n23564, n23565, n23566, n23567, n23568, n23569,
    n23570, n23571, n23572, n23573, n23574, n23575,
    n23576, n23577, n23578, n23579, n23580, n23581,
    n23582, n23583, n23584, n23585, n23586, n23587,
    n23588, n23589, n23590, n23591, n23592, n23593,
    n23594, n23595, n23596, n23597, n23598, n23599,
    n23600, n23601, n23602, n23603, n23604, n23605,
    n23606, n23607, n23608, n23609, n23610, n23611,
    n23612, n23613, n23614, n23615, n23616, n23617,
    n23618, n23619, n23620, n23621, n23622, n23623,
    n23624, n23625, n23626, n23627, n23628, n23629,
    n23630, n23631, n23632, n23633, n23634, n23635,
    n23636, n23637, n23638, n23639, n23640, n23641,
    n23642, n23643, n23644, n23645, n23646, n23647,
    n23648, n23649, n23650, n23651, n23652, n23653,
    n23654, n23655, n23656, n23657, n23658, n23659,
    n23660, n23661, n23662, n23663, n23664, n23665,
    n23666, n23667, n23668, n23669, n23670, n23671,
    n23672, n23673, n23674, n23675, n23676, n23677,
    n23678, n23679, n23680, n23681, n23682, n23683,
    n23684, n23685, n23686, n23687, n23688, n23689,
    n23690, n23691, n23692, n23693, n23694, n23695,
    n23696, n23697, n23698, n23699, n23700, n23701,
    n23702, n23703, n23704, n23705, n23706, n23707,
    n23708, n23709, n23710, n23711, n23712, n23713,
    n23714, n23715, n23716, n23717, n23718, n23719,
    n23720, n23721, n23722, n23723, n23724, n23725,
    n23726, n23727, n23728, n23729, n23730, n23731,
    n23732, n23733, n23734, n23735, n23736, n23737,
    n23738, n23739, n23740, n23741, n23742, n23743,
    n23744, n23745, n23746, n23747, n23748, n23749,
    n23750, n23751, n23752, n23753, n23754, n23755,
    n23756, n23757, n23758, n23759, n23760, n23761,
    n23762, n23763, n23764, n23765, n23766, n23767,
    n23768, n23769, n23770, n23771, n23772, n23773,
    n23774, n23775, n23776, n23777, n23778, n23779,
    n23780, n23781, n23782, n23783, n23784, n23785,
    n23786, n23787, n23788, n23789, n23790, n23791,
    n23792, n23793, n23794, n23795, n23796, n23797,
    n23798, n23799, n23800, n23801, n23802, n23803,
    n23804, n23805, n23806, n23807, n23808, n23809,
    n23810, n23811, n23812, n23813, n23814, n23815,
    n23816, n23817, n23818, n23819, n23820, n23821,
    n23822, n23823, n23824, n23825, n23826, n23827,
    n23828, n23829, n23830, n23831, n23832, n23833,
    n23834, n23835, n23836, n23837, n23838, n23839,
    n23840, n23841, n23842, n23843, n23844, n23845,
    n23846, n23847, n23848, n23849, n23850, n23851,
    n23852, n23853, n23854, n23855, n23856, n23857,
    n23858, n23859, n23860, n23861, n23862, n23863,
    n23864, n23865, n23866, n23867, n23868, n23869,
    n23870, n23871, n23872, n23873, n23874, n23875,
    n23876, n23877, n23878, n23879, n23880, n23881,
    n23882, n23883, n23884, n23885, n23886, n23887,
    n23888, n23889, n23890, n23891, n23892, n23893,
    n23894, n23895, n23896, n23897, n23898, n23899,
    n23900, n23901, n23902, n23903, n23904, n23905,
    n23906, n23907, n23908, n23909, n23910, n23911,
    n23912, n23913, n23914, n23915, n23916, n23917,
    n23918, n23919, n23920, n23921, n23922, n23923,
    n23924, n23925, n23926, n23927, n23928, n23929,
    n23930, n23931, n23932, n23933, n23934, n23935,
    n23936, n23937, n23938, n23939, n23940, n23941,
    n23942, n23943, n23944, n23945, n23946, n23947,
    n23948, n23949, n23950, n23951, n23952, n23953,
    n23954, n23955, n23956, n23957, n23958, n23959,
    n23960, n23961, n23962, n23963, n23964, n23965,
    n23966, n23967, n23968, n23969, n23970, n23971,
    n23972, n23973, n23974, n23975, n23976, n23977,
    n23978, n23979, n23980, n23981, n23982, n23983,
    n23984, n23985, n23986, n23987, n23988, n23989,
    n23990, n23991, n23992, n23993, n23994, n23995,
    n23996, n23997, n23998, n23999, n24000, n24001,
    n24002, n24003, n24004, n24005, n24006, n24007,
    n24008, n24009, n24010, n24011, n24012, n24013,
    n24014, n24015, n24016, n24017, n24018, n24019,
    n24020, n24021, n24022, n24023, n24025, n24026,
    n24027, n24028, n24029, n24030, n24031, n24032,
    n24033, n24034, n24035, n24036, n24037, n24038,
    n24039, n24040, n24041, n24042, n24043, n24044,
    n24045, n24046, n24047, n24048, n24049, n24050,
    n24051, n24052, n24053, n24054, n24055, n24056,
    n24057, n24058, n24059, n24060, n24061, n24062,
    n24063, n24064, n24065, n24066, n24067, n24068,
    n24069, n24070, n24071, n24072, n24073, n24074,
    n24075, n24076, n24077, n24078, n24079, n24080,
    n24081, n24082, n24083, n24084, n24085, n24086,
    n24087, n24088, n24089, n24090, n24091, n24092,
    n24093, n24094, n24095, n24096, n24097, n24098,
    n24099, n24100, n24101, n24102, n24103, n24104,
    n24105, n24106, n24107, n24108, n24109, n24110,
    n24111, n24112, n24113, n24114, n24115, n24116,
    n24117, n24118, n24119, n24120, n24121, n24122,
    n24123, n24124, n24125, n24126, n24127, n24128,
    n24129, n24130, n24131, n24132, n24133, n24134,
    n24135, n24136, n24137, n24138, n24139, n24140,
    n24141, n24142, n24143, n24144, n24145, n24146,
    n24147, n24148, n24149, n24150, n24151, n24152,
    n24153, n24154, n24155, n24156, n24157, n24158,
    n24159, n24160, n24161, n24162, n24163, n24164,
    n24165, n24166, n24167, n24168, n24169, n24170,
    n24171, n24172, n24173, n24174, n24175, n24176,
    n24177, n24178, n24179, n24180, n24181, n24182,
    n24183, n24184, n24185, n24186, n24187, n24188,
    n24189, n24190, n24191, n24192, n24193, n24194,
    n24195, n24196, n24197, n24198, n24199, n24200,
    n24201, n24202, n24203, n24204, n24205, n24206,
    n24207, n24208, n24209, n24210, n24211, n24212,
    n24213, n24214, n24215, n24216, n24217, n24218,
    n24219, n24220, n24221, n24222, n24223, n24224,
    n24225, n24226, n24227, n24228, n24229, n24230,
    n24231, n24232, n24233, n24234, n24235, n24236,
    n24237, n24238, n24239, n24240, n24241, n24242,
    n24243, n24244, n24245, n24246, n24247, n24248,
    n24249, n24250, n24251, n24252, n24253, n24254,
    n24255, n24256, n24257, n24258, n24259, n24260,
    n24261, n24262, n24263, n24264, n24265, n24266,
    n24267, n24268, n24269, n24270, n24271, n24272,
    n24273, n24274, n24275, n24276, n24277, n24278,
    n24279, n24280, n24281, n24282, n24283, n24284,
    n24285, n24286, n24287, n24288, n24289, n24290,
    n24291, n24292, n24293, n24294, n24295, n24296,
    n24297, n24298, n24299, n24300, n24301, n24302,
    n24303, n24304, n24305, n24306, n24307, n24308,
    n24309, n24310, n24311, n24312, n24313, n24314,
    n24315, n24316, n24317, n24318, n24319, n24320,
    n24321, n24322, n24323, n24324, n24325, n24326,
    n24327, n24328, n24329, n24330, n24331, n24332,
    n24333, n24334, n24335, n24336, n24337, n24338,
    n24339, n24340, n24341, n24342, n24343, n24344,
    n24345, n24346, n24347, n24348, n24349, n24350,
    n24351, n24352, n24353, n24354, n24355, n24356,
    n24357, n24358, n24359, n24360, n24361, n24362,
    n24363, n24364, n24365, n24366, n24367, n24368,
    n24369, n24370, n24371, n24372, n24373, n24374,
    n24375, n24376, n24377, n24378, n24379, n24380,
    n24381, n24382, n24383, n24384, n24385, n24386,
    n24387, n24388, n24389, n24390, n24391, n24392,
    n24393, n24394, n24395, n24396, n24397, n24398,
    n24399, n24400, n24401, n24402, n24403, n24404,
    n24405, n24406, n24407, n24408, n24409, n24410,
    n24411, n24412, n24413, n24414, n24415, n24416,
    n24417, n24418, n24419, n24420, n24421, n24422,
    n24423, n24424, n24425, n24426, n24427, n24428,
    n24429, n24430, n24431, n24432, n24433, n24434,
    n24435, n24436, n24437, n24438, n24439, n24440,
    n24441, n24442, n24443, n24444, n24445, n24446,
    n24447, n24448, n24449, n24450, n24451, n24452,
    n24453, n24454, n24455, n24456, n24457, n24458,
    n24459, n24460, n24461, n24462, n24463, n24464,
    n24465, n24466, n24467, n24468, n24469, n24470,
    n24471, n24472, n24473, n24474, n24475, n24476,
    n24477, n24478, n24479, n24480, n24481, n24482,
    n24483, n24484, n24485, n24486, n24487, n24488,
    n24489, n24490, n24491, n24492, n24493, n24494,
    n24495, n24496, n24497, n24498, n24499, n24500,
    n24501, n24502, n24503, n24504, n24505, n24506,
    n24507, n24508, n24509, n24510, n24511, n24512,
    n24513, n24514, n24515, n24516, n24518, n24519,
    n24520, n24521, n24522, n24523, n24524, n24525,
    n24526, n24527, n24528, n24529, n24530, n24531,
    n24532, n24533, n24534, n24535, n24536, n24537,
    n24538, n24539, n24540, n24541, n24542, n24543,
    n24544, n24545, n24546, n24547, n24548, n24549,
    n24550, n24551, n24552, n24553, n24554, n24555,
    n24556, n24557, n24558, n24559, n24560, n24561,
    n24562, n24563, n24564, n24565, n24566, n24567,
    n24568, n24569, n24570, n24571, n24572, n24573,
    n24574, n24575, n24576, n24577, n24578, n24579,
    n24580, n24581, n24582, n24583, n24584, n24585,
    n24586, n24587, n24588, n24589, n24590, n24591,
    n24592, n24593, n24594, n24595, n24596, n24597,
    n24598, n24599, n24600, n24601, n24602, n24603,
    n24604, n24605, n24606, n24607, n24608, n24609,
    n24610, n24611, n24612, n24613, n24614, n24615,
    n24616, n24617, n24618, n24619, n24620, n24621,
    n24622, n24623, n24624, n24625, n24626, n24627,
    n24628, n24629, n24630, n24631, n24632, n24633,
    n24634, n24635, n24636, n24637, n24638, n24639,
    n24640, n24641, n24642, n24643, n24644, n24645,
    n24646, n24647, n24648, n24649, n24650, n24651,
    n24652, n24653, n24654, n24655, n24656, n24657,
    n24658, n24659, n24660, n24661, n24662, n24663,
    n24664, n24665, n24666, n24667, n24668, n24669,
    n24670, n24671, n24672, n24673, n24674, n24675,
    n24676, n24677, n24678, n24679, n24680, n24681,
    n24682, n24683, n24684, n24685, n24686, n24687,
    n24688, n24689, n24690, n24691, n24692, n24693,
    n24694, n24695, n24696, n24697, n24698, n24699,
    n24700, n24701, n24702, n24703, n24704, n24705,
    n24706, n24707, n24708, n24709, n24710, n24711,
    n24712, n24713, n24714, n24715, n24716, n24717,
    n24718, n24719, n24720, n24721, n24722, n24723,
    n24724, n24725, n24726, n24727, n24728, n24729,
    n24730, n24731, n24732, n24733, n24734, n24735,
    n24736, n24737, n24738, n24739, n24740, n24741,
    n24742, n24743, n24744, n24745, n24746, n24747,
    n24748, n24749, n24750, n24751, n24752, n24753,
    n24754, n24755, n24756, n24757, n24758, n24759,
    n24760, n24761, n24762, n24763, n24764, n24765,
    n24766, n24767, n24768, n24769, n24770, n24771,
    n24772, n24773, n24774, n24775, n24776, n24777,
    n24778, n24779, n24780, n24781, n24782, n24783,
    n24784, n24785, n24786, n24787, n24788, n24789,
    n24790, n24791, n24792, n24793, n24794, n24795,
    n24796, n24797, n24798, n24799, n24800, n24801,
    n24802, n24803, n24804, n24805, n24806, n24807,
    n24808, n24809, n24810, n24811, n24812, n24813,
    n24814, n24815, n24816, n24817, n24818, n24819,
    n24820, n24821, n24822, n24823, n24824, n24825,
    n24826, n24827, n24828, n24829, n24830, n24831,
    n24832, n24833, n24834, n24835, n24836, n24837,
    n24838, n24839, n24840, n24841, n24842, n24843,
    n24844, n24845, n24846, n24847, n24848, n24849,
    n24850, n24851, n24852, n24853, n24854, n24855,
    n24856, n24857, n24858, n24859, n24860, n24861,
    n24862, n24863, n24864, n24865, n24866, n24867,
    n24868, n24869, n24870, n24871, n24872, n24873,
    n24874, n24875, n24876, n24877, n24878, n24879,
    n24880, n24881, n24882, n24883, n24884, n24885,
    n24886, n24887, n24888, n24889, n24890, n24891,
    n24892, n24893, n24894, n24895, n24896, n24897,
    n24898, n24899, n24900, n24901, n24902, n24903,
    n24904, n24905, n24906, n24907, n24908, n24909,
    n24910, n24911, n24912, n24913, n24914, n24915,
    n24916, n24917, n24918, n24919, n24920, n24921,
    n24922, n24923, n24924, n24925, n24926, n24927,
    n24928, n24929, n24930, n24931, n24932, n24933,
    n24934, n24935, n24936, n24937, n24938, n24939,
    n24940, n24941, n24942, n24943, n24944, n24945,
    n24946, n24947, n24948, n24949, n24950, n24951,
    n24952, n24953, n24954, n24955, n24956, n24957,
    n24958, n24959, n24960, n24961, n24962, n24963,
    n24964, n24965, n24966, n24967, n24968, n24969,
    n24970, n24971, n24972, n24973, n24974, n24975,
    n24976, n24977, n24978, n24979, n24980, n24981,
    n24982, n24983, n24984, n24985, n24986, n24987,
    n24988, n24989, n24990, n24991, n24992, n24993,
    n24994, n24995, n24996, n24997, n24998, n24999,
    n25000, n25001, n25002, n25003, n25004, n25005,
    n25006, n25007, n25008, n25009, n25010, n25011,
    n25012, n25013, n25014, n25015, n25016, n25017,
    n25018, n25019, n25020, n25021, n25022, n25023,
    n25024, n25025, n25026, n25028, n25029, n25030,
    n25031, n25032, n25033, n25034, n25035, n25036,
    n25037, n25038, n25039, n25040, n25041, n25042,
    n25043, n25044, n25045, n25046, n25047, n25048,
    n25049, n25050, n25051, n25052, n25053, n25054,
    n25055, n25056, n25057, n25058, n25059, n25060,
    n25061, n25062, n25063, n25064, n25065, n25066,
    n25067, n25068, n25069, n25070, n25071, n25072,
    n25073, n25074, n25075, n25076, n25077, n25078,
    n25079, n25080, n25081, n25082, n25083, n25084,
    n25085, n25086, n25087, n25088, n25089, n25090,
    n25091, n25092, n25093, n25094, n25095, n25096,
    n25097, n25098, n25099, n25100, n25101, n25102,
    n25103, n25104, n25105, n25106, n25107, n25108,
    n25109, n25110, n25111, n25112, n25113, n25114,
    n25115, n25116, n25117, n25118, n25119, n25120,
    n25121, n25122, n25123, n25124, n25125, n25126,
    n25127, n25128, n25129, n25130, n25131, n25132,
    n25133, n25134, n25135, n25136, n25137, n25138,
    n25139, n25140, n25141, n25142, n25143, n25144,
    n25145, n25146, n25147, n25148, n25149, n25150,
    n25151, n25152, n25153, n25154, n25155, n25156,
    n25157, n25158, n25159, n25160, n25161, n25162,
    n25163, n25164, n25165, n25166, n25167, n25168,
    n25169, n25170, n25171, n25172, n25173, n25174,
    n25175, n25176, n25177, n25178, n25179, n25180,
    n25181, n25182, n25183, n25184, n25185, n25186,
    n25187, n25188, n25189, n25190, n25191, n25192,
    n25193, n25194, n25195, n25196, n25197, n25198,
    n25199, n25200, n25201, n25202, n25203, n25204,
    n25205, n25206, n25207, n25208, n25209, n25210,
    n25211, n25212, n25213, n25214, n25215, n25216,
    n25217, n25218, n25219, n25220, n25221, n25222,
    n25223, n25224, n25225, n25226, n25227, n25228,
    n25229, n25230, n25231, n25232, n25233, n25234,
    n25235, n25236, n25237, n25238, n25239, n25240,
    n25241, n25242, n25243, n25244, n25245, n25246,
    n25247, n25248, n25249, n25250, n25251, n25252,
    n25253, n25254, n25255, n25256, n25257, n25258,
    n25259, n25260, n25261, n25262, n25263, n25264,
    n25265, n25266, n25267, n25268, n25269, n25270,
    n25271, n25272, n25273, n25274, n25275, n25276,
    n25277, n25278, n25279, n25280, n25281, n25282,
    n25283, n25284, n25285, n25286, n25287, n25288,
    n25289, n25290, n25291, n25292, n25293, n25294,
    n25295, n25296, n25297, n25298, n25299, n25300,
    n25301, n25302, n25303, n25304, n25305, n25306,
    n25307, n25308, n25309, n25310, n25311, n25312,
    n25313, n25314, n25315, n25316, n25317, n25318,
    n25319, n25320, n25321, n25322, n25323, n25324,
    n25325, n25326, n25327, n25328, n25329, n25330,
    n25331, n25332, n25333, n25334, n25335, n25336,
    n25337, n25338, n25339, n25340, n25341, n25342,
    n25343, n25344, n25345, n25346, n25347, n25348,
    n25349, n25350, n25351, n25352, n25353, n25354,
    n25355, n25356, n25357, n25358, n25359, n25360,
    n25361, n25362, n25363, n25364, n25365, n25366,
    n25367, n25368, n25369, n25370, n25371, n25372,
    n25373, n25374, n25375, n25376, n25377, n25378,
    n25379, n25380, n25381, n25382, n25383, n25384,
    n25385, n25386, n25387, n25388, n25389, n25390,
    n25391, n25392, n25393, n25394, n25395, n25396,
    n25397, n25398, n25399, n25400, n25401, n25402,
    n25403, n25404, n25405, n25406, n25407, n25408,
    n25409, n25410, n25411, n25412, n25413, n25414,
    n25415, n25416, n25417, n25418, n25419, n25420,
    n25421, n25422, n25423, n25424, n25425, n25426,
    n25427, n25428, n25429, n25430, n25431, n25432,
    n25433, n25434, n25435, n25436, n25437, n25438,
    n25439, n25440, n25441, n25442, n25443, n25444,
    n25445, n25446, n25447, n25448, n25449, n25450,
    n25451, n25452, n25453, n25454, n25455, n25456,
    n25457, n25458, n25459, n25460, n25461, n25462,
    n25463, n25464, n25465, n25466, n25467, n25468,
    n25469, n25470, n25471, n25472, n25473, n25474,
    n25475, n25476, n25477, n25478, n25479, n25480,
    n25481, n25482, n25483, n25484, n25485, n25486,
    n25487, n25488, n25489, n25490, n25491, n25492,
    n25493, n25494, n25495, n25496, n25497, n25498,
    n25499, n25500, n25502, n25503, n25504, n25505,
    n25506, n25507, n25508, n25509, n25510, n25511,
    n25512, n25513, n25514, n25515, n25516, n25517,
    n25518, n25519, n25520, n25521, n25522, n25523,
    n25524, n25525, n25526, n25527, n25528, n25529,
    n25530, n25531, n25532, n25533, n25534, n25535,
    n25536, n25537, n25538, n25539, n25540, n25541,
    n25542, n25543, n25544, n25545, n25546, n25547,
    n25548, n25549, n25550, n25551, n25552, n25553,
    n25554, n25555, n25556, n25557, n25558, n25559,
    n25560, n25561, n25562, n25563, n25564, n25565,
    n25566, n25567, n25568, n25569, n25570, n25571,
    n25572, n25573, n25574, n25575, n25576, n25577,
    n25578, n25579, n25580, n25581, n25582, n25583,
    n25584, n25585, n25586, n25587, n25588, n25589,
    n25590, n25591, n25592, n25593, n25594, n25595,
    n25596, n25597, n25598, n25599, n25600, n25601,
    n25602, n25603, n25604, n25605, n25606, n25607,
    n25608, n25609, n25610, n25611, n25612, n25613,
    n25614, n25615, n25616, n25617, n25618, n25619,
    n25620, n25621, n25622, n25623, n25624, n25625,
    n25626, n25627, n25628, n25629, n25630, n25631,
    n25632, n25633, n25634, n25635, n25636, n25637,
    n25638, n25639, n25640, n25641, n25642, n25643,
    n25644, n25645, n25646, n25647, n25648, n25649,
    n25650, n25651, n25652, n25653, n25654, n25655,
    n25656, n25657, n25658, n25659, n25660, n25661,
    n25662, n25663, n25664, n25665, n25666, n25667,
    n25668, n25669, n25670, n25671, n25672, n25673,
    n25674, n25675, n25676, n25677, n25678, n25679,
    n25680, n25681, n25682, n25683, n25684, n25685,
    n25686, n25687, n25688, n25689, n25690, n25691,
    n25692, n25693, n25694, n25695, n25696, n25697,
    n25698, n25699, n25700, n25701, n25702, n25703,
    n25704, n25705, n25706, n25707, n25708, n25709,
    n25710, n25711, n25712, n25713, n25714, n25715,
    n25716, n25717, n25718, n25719, n25720, n25721,
    n25722, n25723, n25724, n25725, n25726, n25727,
    n25728, n25729, n25730, n25731, n25732, n25733,
    n25734, n25735, n25736, n25737, n25738, n25739,
    n25740, n25741, n25742, n25743, n25744, n25745,
    n25746, n25747, n25748, n25749, n25750, n25751,
    n25752, n25753, n25754, n25755, n25756, n25757,
    n25758, n25759, n25760, n25761, n25762, n25763,
    n25764, n25765, n25766, n25767, n25768, n25769,
    n25770, n25771, n25772, n25773, n25774, n25775,
    n25776, n25777, n25778, n25779, n25780, n25781,
    n25782, n25783, n25784, n25785, n25786, n25787,
    n25788, n25789, n25790, n25791, n25792, n25793,
    n25794, n25795, n25796, n25797, n25798, n25799,
    n25800, n25801, n25802, n25803, n25804, n25805,
    n25806, n25807, n25808, n25809, n25810, n25811,
    n25812, n25813, n25814, n25815, n25816, n25817,
    n25818, n25819, n25820, n25821, n25822, n25823,
    n25824, n25825, n25826, n25827, n25828, n25829,
    n25830, n25831, n25832, n25833, n25834, n25835,
    n25836, n25837, n25838, n25839, n25840, n25841,
    n25842, n25843, n25844, n25845, n25846, n25847,
    n25848, n25849, n25850, n25851, n25852, n25853,
    n25854, n25855, n25856, n25857, n25858, n25859,
    n25860, n25861, n25862, n25863, n25864, n25865,
    n25866, n25867, n25868, n25869, n25870, n25871,
    n25872, n25873, n25874, n25875, n25876, n25877,
    n25878, n25879, n25880, n25881, n25882, n25883,
    n25884, n25885, n25886, n25887, n25888, n25889,
    n25890, n25891, n25892, n25893, n25894, n25895,
    n25896, n25897, n25898, n25899, n25900, n25901,
    n25902, n25903, n25904, n25905, n25906, n25907,
    n25908, n25909, n25910, n25911, n25912, n25913,
    n25914, n25915, n25916, n25917, n25918, n25919,
    n25920, n25921, n25922, n25923, n25924, n25925,
    n25926, n25927, n25928, n25929, n25930, n25931,
    n25932, n25933, n25934, n25935, n25936, n25937,
    n25938, n25939, n25940, n25941, n25943, n25944,
    n25945, n25946, n25947, n25948, n25949, n25950,
    n25951, n25952, n25953, n25954, n25955, n25956,
    n25957, n25958, n25959, n25960, n25961, n25962,
    n25963, n25964, n25965, n25966, n25967, n25968,
    n25969, n25970, n25971, n25972, n25973, n25974,
    n25975, n25976, n25977, n25978, n25979, n25980,
    n25981, n25982, n25983, n25984, n25985, n25986,
    n25987, n25988, n25989, n25990, n25991, n25992,
    n25993, n25994, n25995, n25996, n25997, n25998,
    n25999, n26000, n26001, n26002, n26003, n26004,
    n26005, n26006, n26007, n26008, n26009, n26010,
    n26011, n26012, n26013, n26014, n26015, n26016,
    n26017, n26018, n26019, n26020, n26021, n26022,
    n26023, n26024, n26025, n26026, n26027, n26028,
    n26029, n26030, n26031, n26032, n26033, n26034,
    n26035, n26036, n26037, n26038, n26039, n26040,
    n26041, n26042, n26043, n26044, n26045, n26046,
    n26047, n26048, n26049, n26050, n26051, n26052,
    n26053, n26054, n26055, n26056, n26057, n26058,
    n26059, n26060, n26061, n26062, n26063, n26064,
    n26065, n26066, n26067, n26068, n26069, n26070,
    n26071, n26072, n26073, n26074, n26075, n26076,
    n26077, n26078, n26079, n26080, n26081, n26082,
    n26083, n26084, n26085, n26086, n26087, n26088,
    n26089, n26090, n26091, n26092, n26093, n26094,
    n26095, n26096, n26097, n26098, n26099, n26100,
    n26101, n26102, n26103, n26104, n26105, n26106,
    n26107, n26108, n26109, n26110, n26111, n26112,
    n26113, n26114, n26115, n26116, n26117, n26118,
    n26119, n26120, n26121, n26122, n26123, n26124,
    n26125, n26126, n26127, n26128, n26129, n26130,
    n26131, n26132, n26133, n26134, n26135, n26136,
    n26137, n26138, n26139, n26140, n26141, n26142,
    n26143, n26144, n26145, n26146, n26147, n26148,
    n26149, n26150, n26151, n26152, n26153, n26154,
    n26155, n26156, n26157, n26158, n26159, n26160,
    n26161, n26162, n26163, n26164, n26165, n26166,
    n26167, n26168, n26169, n26170, n26171, n26172,
    n26173, n26174, n26175, n26176, n26177, n26178,
    n26179, n26180, n26181, n26182, n26183, n26184,
    n26185, n26186, n26187, n26188, n26189, n26190,
    n26191, n26192, n26193, n26194, n26195, n26196,
    n26197, n26198, n26199, n26200, n26201, n26202,
    n26203, n26204, n26205, n26206, n26207, n26208,
    n26209, n26210, n26211, n26212, n26213, n26214,
    n26215, n26216, n26217, n26218, n26219, n26220,
    n26221, n26222, n26223, n26224, n26225, n26226,
    n26227, n26228, n26229, n26230, n26231, n26232,
    n26233, n26234, n26235, n26236, n26237, n26238,
    n26239, n26240, n26241, n26242, n26243, n26244,
    n26245, n26246, n26247, n26248, n26249, n26250,
    n26251, n26252, n26253, n26254, n26255, n26256,
    n26257, n26258, n26259, n26260, n26261, n26262,
    n26263, n26264, n26265, n26266, n26267, n26268,
    n26269, n26270, n26271, n26272, n26273, n26274,
    n26275, n26276, n26277, n26278, n26279, n26280,
    n26281, n26282, n26283, n26284, n26285, n26286,
    n26287, n26288, n26289, n26290, n26291, n26292,
    n26293, n26294, n26295, n26296, n26297, n26298,
    n26299, n26300, n26301, n26302, n26303, n26304,
    n26305, n26306, n26307, n26308, n26309, n26310,
    n26311, n26312, n26313, n26314, n26315, n26316,
    n26317, n26318, n26319, n26320, n26321, n26322,
    n26323, n26324, n26325, n26326, n26327, n26328,
    n26329, n26330, n26331, n26332, n26333, n26334,
    n26335, n26336, n26337, n26338, n26339, n26340,
    n26341, n26342, n26343, n26344, n26345, n26346,
    n26347, n26348, n26349, n26350, n26351, n26352,
    n26353, n26354, n26355, n26356, n26357, n26358,
    n26359, n26360, n26361, n26362, n26363, n26364,
    n26365, n26366, n26367, n26368, n26369, n26370,
    n26371, n26372, n26373, n26374, n26375, n26376,
    n26377, n26378, n26379, n26380, n26381, n26382,
    n26383, n26384, n26385, n26386, n26387, n26388,
    n26389, n26390, n26391, n26392, n26393, n26394,
    n26395, n26396, n26397, n26398, n26399, n26400,
    n26401, n26402, n26403, n26404, n26405, n26406,
    n26407, n26408, n26409, n26410, n26411, n26412,
    n26413, n26414, n26415, n26416, n26417, n26418,
    n26419, n26420, n26421, n26423, n26424, n26425,
    n26426, n26427, n26428, n26429, n26430, n26431,
    n26432, n26433, n26434, n26435, n26436, n26437,
    n26438, n26439, n26440, n26441, n26442, n26443,
    n26444, n26445, n26446, n26447, n26448, n26449,
    n26450, n26451, n26452, n26453, n26454, n26455,
    n26456, n26457, n26458, n26459, n26460, n26461,
    n26462, n26463, n26464, n26465, n26466, n26467,
    n26468, n26469, n26470, n26471, n26472, n26473,
    n26474, n26475, n26476, n26477, n26478, n26479,
    n26480, n26481, n26482, n26483, n26484, n26485,
    n26486, n26487, n26488, n26489, n26490, n26491,
    n26492, n26493, n26494, n26495, n26496, n26497,
    n26498, n26499, n26500, n26501, n26502, n26503,
    n26504, n26505, n26506, n26507, n26508, n26509,
    n26510, n26511, n26512, n26513, n26514, n26515,
    n26516, n26517, n26518, n26519, n26520, n26521,
    n26522, n26523, n26524, n26525, n26526, n26527,
    n26528, n26529, n26530, n26531, n26532, n26533,
    n26534, n26535, n26536, n26537, n26538, n26539,
    n26540, n26541, n26542, n26543, n26544, n26545,
    n26546, n26547, n26548, n26549, n26550, n26551,
    n26552, n26553, n26554, n26555, n26556, n26557,
    n26558, n26559, n26560, n26561, n26562, n26563,
    n26564, n26565, n26566, n26567, n26568, n26569,
    n26570, n26571, n26572, n26573, n26574, n26575,
    n26576, n26577, n26578, n26579, n26580, n26581,
    n26582, n26583, n26584, n26585, n26586, n26587,
    n26588, n26589, n26590, n26591, n26592, n26593,
    n26594, n26595, n26596, n26597, n26598, n26599,
    n26600, n26601, n26602, n26603, n26604, n26605,
    n26606, n26607, n26608, n26609, n26610, n26611,
    n26612, n26613, n26614, n26615, n26616, n26617,
    n26618, n26619, n26620, n26621, n26622, n26623,
    n26624, n26625, n26626, n26627, n26628, n26629,
    n26630, n26631, n26632, n26633, n26634, n26635,
    n26636, n26637, n26638, n26639, n26640, n26641,
    n26642, n26643, n26644, n26645, n26646, n26647,
    n26648, n26649, n26650, n26651, n26652, n26653,
    n26654, n26655, n26656, n26657, n26658, n26659,
    n26660, n26661, n26662, n26663, n26664, n26665,
    n26666, n26667, n26668, n26669, n26670, n26671,
    n26672, n26673, n26674, n26675, n26676, n26677,
    n26678, n26679, n26680, n26681, n26682, n26683,
    n26684, n26685, n26686, n26687, n26688, n26689,
    n26690, n26691, n26692, n26693, n26694, n26695,
    n26696, n26697, n26698, n26699, n26700, n26701,
    n26702, n26703, n26704, n26705, n26706, n26707,
    n26708, n26709, n26710, n26711, n26712, n26713,
    n26714, n26715, n26716, n26717, n26718, n26719,
    n26720, n26721, n26722, n26723, n26724, n26725,
    n26726, n26727, n26728, n26729, n26730, n26731,
    n26732, n26733, n26734, n26735, n26736, n26737,
    n26738, n26739, n26740, n26741, n26742, n26743,
    n26744, n26745, n26746, n26747, n26748, n26749,
    n26750, n26751, n26752, n26753, n26754, n26755,
    n26756, n26757, n26758, n26759, n26760, n26761,
    n26762, n26763, n26764, n26765, n26766, n26767,
    n26768, n26769, n26770, n26771, n26772, n26773,
    n26774, n26775, n26776, n26777, n26778, n26779,
    n26780, n26781, n26782, n26783, n26784, n26785,
    n26786, n26787, n26788, n26789, n26790, n26791,
    n26792, n26793, n26794, n26795, n26796, n26797,
    n26798, n26799, n26800, n26801, n26802, n26803,
    n26804, n26805, n26806, n26807, n26808, n26809,
    n26810, n26811, n26812, n26813, n26814, n26815,
    n26816, n26817, n26818, n26819, n26820, n26821,
    n26822, n26823, n26824, n26825, n26826, n26827,
    n26828, n26829, n26830, n26831, n26832, n26833,
    n26835, n26836, n26837, n26838, n26839, n26840,
    n26841, n26842, n26843, n26844, n26845, n26846,
    n26847, n26848, n26849, n26850, n26851, n26852,
    n26853, n26854, n26855, n26856, n26857, n26858,
    n26859, n26860, n26861, n26862, n26863, n26864,
    n26865, n26866, n26867, n26868, n26869, n26870,
    n26871, n26872, n26873, n26874, n26875, n26876,
    n26877, n26878, n26879, n26880, n26881, n26882,
    n26883, n26884, n26885, n26886, n26887, n26888,
    n26889, n26890, n26891, n26892, n26893, n26894,
    n26895, n26896, n26897, n26898, n26899, n26900,
    n26901, n26902, n26903, n26904, n26905, n26906,
    n26907, n26908, n26909, n26910, n26911, n26912,
    n26913, n26914, n26915, n26916, n26917, n26918,
    n26919, n26920, n26921, n26922, n26923, n26924,
    n26925, n26926, n26927, n26928, n26929, n26930,
    n26931, n26932, n26933, n26934, n26935, n26936,
    n26937, n26938, n26939, n26940, n26941, n26942,
    n26943, n26944, n26945, n26946, n26947, n26948,
    n26949, n26950, n26951, n26952, n26953, n26954,
    n26955, n26956, n26957, n26958, n26959, n26960,
    n26961, n26962, n26963, n26964, n26965, n26966,
    n26967, n26968, n26969, n26970, n26971, n26972,
    n26973, n26974, n26975, n26976, n26977, n26978,
    n26979, n26980, n26981, n26982, n26983, n26984,
    n26985, n26986, n26987, n26988, n26989, n26990,
    n26991, n26992, n26993, n26994, n26995, n26996,
    n26997, n26998, n26999, n27000, n27001, n27002,
    n27003, n27004, n27005, n27006, n27007, n27008,
    n27009, n27010, n27011, n27012, n27013, n27014,
    n27015, n27016, n27017, n27018, n27019, n27020,
    n27021, n27022, n27023, n27024, n27025, n27026,
    n27027, n27028, n27029, n27030, n27031, n27032,
    n27033, n27034, n27035, n27036, n27037, n27038,
    n27039, n27040, n27041, n27042, n27043, n27044,
    n27045, n27046, n27047, n27048, n27049, n27050,
    n27051, n27052, n27053, n27054, n27055, n27056,
    n27057, n27058, n27059, n27060, n27061, n27062,
    n27063, n27064, n27065, n27066, n27067, n27068,
    n27069, n27070, n27071, n27072, n27073, n27074,
    n27075, n27076, n27077, n27078, n27079, n27080,
    n27081, n27082, n27083, n27084, n27085, n27086,
    n27087, n27088, n27089, n27090, n27091, n27092,
    n27093, n27094, n27095, n27096, n27097, n27098,
    n27099, n27100, n27101, n27102, n27103, n27104,
    n27105, n27106, n27107, n27108, n27109, n27110,
    n27111, n27112, n27113, n27114, n27115, n27116,
    n27117, n27118, n27119, n27120, n27121, n27122,
    n27123, n27124, n27125, n27126, n27127, n27128,
    n27129, n27130, n27131, n27132, n27133, n27134,
    n27135, n27136, n27137, n27138, n27139, n27140,
    n27141, n27142, n27143, n27144, n27145, n27146,
    n27147, n27148, n27149, n27150, n27151, n27152,
    n27153, n27154, n27155, n27156, n27157, n27158,
    n27159, n27160, n27161, n27162, n27163, n27164,
    n27165, n27166, n27167, n27168, n27169, n27170,
    n27171, n27172, n27173, n27174, n27175, n27176,
    n27177, n27178, n27179, n27180, n27181, n27182,
    n27183, n27184, n27185, n27186, n27187, n27188,
    n27189, n27190, n27191, n27192, n27193, n27194,
    n27195, n27196, n27197, n27198, n27199, n27200,
    n27201, n27202, n27203, n27204, n27205, n27206,
    n27207, n27208, n27209, n27210, n27211, n27212,
    n27213, n27214, n27215, n27216, n27217, n27218,
    n27219, n27220, n27221, n27222, n27223, n27224,
    n27225, n27226, n27227, n27228, n27229, n27230,
    n27231, n27232, n27233, n27234, n27235, n27236,
    n27237, n27238, n27239, n27240, n27241, n27242,
    n27243, n27244, n27245, n27246, n27247, n27248,
    n27249, n27250, n27251, n27252, n27253, n27254,
    n27255, n27256, n27257, n27258, n27259, n27260,
    n27261, n27262, n27263, n27264, n27265, n27267,
    n27268, n27269, n27270, n27271, n27272, n27273,
    n27274, n27275, n27276, n27277, n27278, n27279,
    n27280, n27281, n27282, n27283, n27284, n27285,
    n27286, n27287, n27288, n27289, n27290, n27291,
    n27292, n27293, n27294, n27295, n27296, n27297,
    n27298, n27299, n27300, n27301, n27302, n27303,
    n27304, n27305, n27306, n27307, n27308, n27309,
    n27310, n27311, n27312, n27313, n27314, n27315,
    n27316, n27317, n27318, n27319, n27320, n27321,
    n27322, n27323, n27324, n27325, n27326, n27327,
    n27328, n27329, n27330, n27331, n27332, n27333,
    n27334, n27335, n27336, n27337, n27338, n27339,
    n27340, n27341, n27342, n27343, n27344, n27345,
    n27346, n27347, n27348, n27349, n27350, n27351,
    n27352, n27353, n27354, n27355, n27356, n27357,
    n27358, n27359, n27360, n27361, n27362, n27363,
    n27364, n27365, n27366, n27367, n27368, n27369,
    n27370, n27371, n27372, n27373, n27374, n27375,
    n27376, n27377, n27378, n27379, n27380, n27381,
    n27382, n27383, n27384, n27385, n27386, n27387,
    n27388, n27389, n27390, n27391, n27392, n27393,
    n27394, n27395, n27396, n27397, n27398, n27399,
    n27400, n27401, n27402, n27403, n27404, n27405,
    n27406, n27407, n27408, n27409, n27410, n27411,
    n27412, n27413, n27414, n27415, n27416, n27417,
    n27418, n27419, n27420, n27421, n27422, n27423,
    n27424, n27425, n27426, n27427, n27428, n27429,
    n27430, n27431, n27432, n27433, n27434, n27435,
    n27436, n27437, n27438, n27439, n27440, n27441,
    n27442, n27443, n27444, n27445, n27446, n27447,
    n27448, n27449, n27450, n27451, n27452, n27453,
    n27454, n27455, n27456, n27457, n27458, n27459,
    n27460, n27461, n27462, n27463, n27464, n27465,
    n27466, n27467, n27468, n27469, n27470, n27471,
    n27472, n27473, n27474, n27475, n27476, n27477,
    n27478, n27479, n27480, n27481, n27482, n27483,
    n27484, n27485, n27486, n27487, n27488, n27489,
    n27490, n27491, n27492, n27493, n27494, n27495,
    n27496, n27497, n27498, n27499, n27500, n27501,
    n27502, n27503, n27504, n27505, n27506, n27507,
    n27508, n27509, n27510, n27511, n27512, n27513,
    n27514, n27515, n27516, n27517, n27518, n27519,
    n27520, n27521, n27522, n27523, n27524, n27525,
    n27526, n27527, n27528, n27529, n27530, n27531,
    n27532, n27533, n27534, n27535, n27536, n27537,
    n27538, n27539, n27540, n27541, n27542, n27543,
    n27544, n27545, n27546, n27547, n27548, n27549,
    n27550, n27551, n27552, n27553, n27554, n27555,
    n27556, n27557, n27558, n27559, n27560, n27561,
    n27562, n27563, n27564, n27565, n27566, n27567,
    n27568, n27569, n27570, n27571, n27572, n27573,
    n27574, n27575, n27576, n27577, n27578, n27579,
    n27580, n27581, n27582, n27583, n27584, n27585,
    n27586, n27587, n27588, n27589, n27590, n27591,
    n27592, n27593, n27594, n27595, n27596, n27597,
    n27598, n27599, n27600, n27601, n27602, n27603,
    n27604, n27605, n27606, n27607, n27608, n27609,
    n27610, n27611, n27612, n27613, n27614, n27615,
    n27616, n27617, n27618, n27619, n27620, n27621,
    n27622, n27623, n27624, n27625, n27626, n27627,
    n27628, n27629, n27630, n27631, n27632, n27633,
    n27634, n27635, n27636, n27637, n27638, n27639,
    n27640, n27641, n27642, n27643, n27644, n27645,
    n27646, n27647, n27648, n27649, n27650, n27651,
    n27652, n27653, n27654, n27655, n27656, n27657,
    n27658, n27659, n27660, n27661, n27662, n27663,
    n27664, n27665, n27666, n27667, n27668, n27669,
    n27670, n27671, n27672, n27673, n27674, n27675,
    n27676, n27677, n27678, n27679, n27680, n27681,
    n27682, n27683, n27684, n27685, n27686, n27687,
    n27689, n27690, n27691, n27692, n27693, n27694,
    n27695, n27696, n27697, n27698, n27699, n27700,
    n27701, n27702, n27703, n27704, n27705, n27706,
    n27707, n27708, n27709, n27710, n27711, n27712,
    n27713, n27714, n27715, n27716, n27717, n27718,
    n27719, n27720, n27721, n27722, n27723, n27724,
    n27725, n27726, n27727, n27728, n27729, n27730,
    n27731, n27732, n27733, n27734, n27735, n27736,
    n27737, n27738, n27739, n27740, n27741, n27742,
    n27743, n27744, n27745, n27746, n27747, n27748,
    n27749, n27750, n27751, n27752, n27753, n27754,
    n27755, n27756, n27757, n27758, n27759, n27760,
    n27761, n27762, n27763, n27764, n27765, n27766,
    n27767, n27768, n27769, n27770, n27771, n27772,
    n27773, n27774, n27775, n27776, n27777, n27778,
    n27779, n27780, n27781, n27782, n27783, n27784,
    n27785, n27786, n27787, n27788, n27789, n27790,
    n27791, n27792, n27793, n27794, n27795, n27796,
    n27797, n27798, n27799, n27800, n27801, n27802,
    n27803, n27804, n27805, n27806, n27807, n27808,
    n27809, n27810, n27811, n27812, n27813, n27814,
    n27815, n27816, n27817, n27818, n27819, n27820,
    n27821, n27822, n27823, n27824, n27825, n27826,
    n27827, n27828, n27829, n27830, n27831, n27832,
    n27833, n27834, n27835, n27836, n27837, n27838,
    n27839, n27840, n27841, n27842, n27843, n27844,
    n27845, n27846, n27847, n27848, n27849, n27850,
    n27851, n27852, n27853, n27854, n27855, n27856,
    n27857, n27858, n27859, n27860, n27861, n27862,
    n27863, n27864, n27865, n27866, n27867, n27868,
    n27869, n27870, n27871, n27872, n27873, n27874,
    n27875, n27876, n27877, n27878, n27879, n27880,
    n27881, n27882, n27883, n27884, n27885, n27886,
    n27887, n27888, n27889, n27890, n27891, n27892,
    n27893, n27894, n27895, n27896, n27897, n27898,
    n27899, n27900, n27901, n27902, n27903, n27904,
    n27905, n27906, n27907, n27908, n27909, n27910,
    n27911, n27912, n27913, n27914, n27915, n27916,
    n27917, n27918, n27919, n27920, n27921, n27922,
    n27923, n27924, n27925, n27926, n27927, n27928,
    n27929, n27930, n27931, n27932, n27933, n27934,
    n27935, n27936, n27937, n27938, n27939, n27940,
    n27941, n27942, n27943, n27944, n27945, n27946,
    n27947, n27948, n27949, n27950, n27951, n27952,
    n27953, n27954, n27955, n27956, n27957, n27958,
    n27959, n27960, n27961, n27962, n27963, n27964,
    n27965, n27966, n27967, n27968, n27969, n27970,
    n27971, n27972, n27973, n27974, n27975, n27976,
    n27977, n27978, n27979, n27980, n27981, n27982,
    n27983, n27984, n27985, n27986, n27987, n27988,
    n27989, n27990, n27991, n27992, n27993, n27994,
    n27995, n27996, n27997, n27998, n27999, n28000,
    n28001, n28002, n28003, n28004, n28005, n28006,
    n28007, n28008, n28009, n28010, n28011, n28012,
    n28013, n28014, n28015, n28016, n28017, n28018,
    n28019, n28020, n28021, n28022, n28023, n28024,
    n28025, n28026, n28027, n28028, n28029, n28030,
    n28031, n28032, n28033, n28034, n28035, n28036,
    n28037, n28038, n28039, n28040, n28041, n28042,
    n28043, n28044, n28045, n28046, n28047, n28048,
    n28049, n28050, n28051, n28052, n28053, n28054,
    n28055, n28056, n28057, n28058, n28059, n28060,
    n28061, n28062, n28063, n28064, n28065, n28066,
    n28067, n28068, n28069, n28070, n28071, n28072,
    n28073, n28074, n28075, n28076, n28077, n28078,
    n28079, n28080, n28081, n28082, n28083, n28084,
    n28085, n28086, n28087, n28088, n28090, n28091,
    n28092, n28093, n28094, n28095, n28096, n28097,
    n28098, n28099, n28100, n28101, n28102, n28103,
    n28104, n28105, n28106, n28107, n28108, n28109,
    n28110, n28111, n28112, n28113, n28114, n28115,
    n28116, n28117, n28118, n28119, n28120, n28121,
    n28122, n28123, n28124, n28125, n28126, n28127,
    n28128, n28129, n28130, n28131, n28132, n28133,
    n28134, n28135, n28136, n28137, n28138, n28139,
    n28140, n28141, n28142, n28143, n28144, n28145,
    n28146, n28147, n28148, n28149, n28150, n28151,
    n28152, n28153, n28154, n28155, n28156, n28157,
    n28158, n28159, n28160, n28161, n28162, n28163,
    n28164, n28165, n28166, n28167, n28168, n28169,
    n28170, n28171, n28172, n28173, n28174, n28175,
    n28176, n28177, n28178, n28179, n28180, n28181,
    n28182, n28183, n28184, n28185, n28186, n28187,
    n28188, n28189, n28190, n28191, n28192, n28193,
    n28194, n28195, n28196, n28197, n28198, n28199,
    n28200, n28201, n28202, n28203, n28204, n28205,
    n28206, n28207, n28208, n28209, n28210, n28211,
    n28212, n28213, n28214, n28215, n28216, n28217,
    n28218, n28219, n28220, n28221, n28222, n28223,
    n28224, n28225, n28226, n28227, n28228, n28229,
    n28230, n28231, n28232, n28233, n28234, n28235,
    n28236, n28237, n28238, n28239, n28240, n28241,
    n28242, n28243, n28244, n28245, n28246, n28247,
    n28248, n28249, n28250, n28251, n28252, n28253,
    n28254, n28255, n28256, n28257, n28258, n28259,
    n28260, n28261, n28262, n28263, n28264, n28265,
    n28266, n28267, n28268, n28269, n28270, n28271,
    n28272, n28273, n28274, n28275, n28276, n28277,
    n28278, n28279, n28280, n28281, n28282, n28283,
    n28284, n28285, n28286, n28287, n28288, n28289,
    n28290, n28291, n28292, n28293, n28294, n28295,
    n28296, n28297, n28298, n28299, n28300, n28301,
    n28302, n28303, n28304, n28305, n28306, n28307,
    n28308, n28309, n28310, n28311, n28312, n28313,
    n28314, n28315, n28316, n28317, n28318, n28319,
    n28320, n28321, n28322, n28323, n28324, n28325,
    n28326, n28327, n28328, n28329, n28330, n28331,
    n28332, n28333, n28334, n28335, n28336, n28337,
    n28338, n28339, n28340, n28341, n28342, n28343,
    n28344, n28345, n28346, n28347, n28348, n28349,
    n28350, n28351, n28352, n28353, n28354, n28355,
    n28356, n28357, n28358, n28359, n28360, n28361,
    n28362, n28363, n28364, n28365, n28366, n28367,
    n28368, n28369, n28370, n28371, n28372, n28373,
    n28374, n28375, n28376, n28377, n28378, n28379,
    n28380, n28381, n28382, n28383, n28384, n28385,
    n28386, n28387, n28388, n28389, n28390, n28391,
    n28392, n28393, n28394, n28395, n28396, n28397,
    n28398, n28399, n28400, n28401, n28402, n28403,
    n28404, n28405, n28406, n28407, n28408, n28409,
    n28410, n28411, n28412, n28413, n28414, n28415,
    n28416, n28417, n28418, n28419, n28420, n28421,
    n28422, n28423, n28424, n28425, n28426, n28427,
    n28428, n28429, n28430, n28431, n28432, n28433,
    n28434, n28435, n28436, n28437, n28438, n28439,
    n28440, n28441, n28442, n28443, n28444, n28445,
    n28446, n28447, n28448, n28449, n28450, n28451,
    n28452, n28453, n28454, n28455, n28456, n28457,
    n28458, n28459, n28460, n28461, n28462, n28463,
    n28464, n28465, n28466, n28467, n28468, n28469,
    n28470, n28471, n28472, n28473, n28474, n28475,
    n28476, n28477, n28478, n28479, n28480, n28481,
    n28482, n28484, n28485, n28486, n28487, n28488,
    n28489, n28490, n28491, n28492, n28493, n28494,
    n28495, n28496, n28497, n28498, n28499, n28500,
    n28501, n28502, n28503, n28504, n28505, n28506,
    n28507, n28508, n28509, n28510, n28511, n28512,
    n28513, n28514, n28515, n28516, n28517, n28518,
    n28519, n28520, n28521, n28522, n28523, n28524,
    n28525, n28526, n28527, n28528, n28529, n28530,
    n28531, n28532, n28533, n28534, n28535, n28536,
    n28537, n28538, n28539, n28540, n28541, n28542,
    n28543, n28544, n28545, n28546, n28547, n28548,
    n28549, n28550, n28551, n28552, n28553, n28554,
    n28555, n28556, n28557, n28558, n28559, n28560,
    n28561, n28562, n28563, n28564, n28565, n28566,
    n28567, n28568, n28569, n28570, n28571, n28572,
    n28573, n28574, n28575, n28576, n28577, n28578,
    n28579, n28580, n28581, n28582, n28583, n28584,
    n28585, n28586, n28587, n28588, n28589, n28590,
    n28591, n28592, n28593, n28594, n28595, n28596,
    n28597, n28598, n28599, n28600, n28601, n28602,
    n28603, n28604, n28605, n28606, n28607, n28608,
    n28609, n28610, n28611, n28612, n28613, n28614,
    n28615, n28616, n28617, n28618, n28619, n28620,
    n28621, n28622, n28623, n28624, n28625, n28626,
    n28627, n28628, n28629, n28630, n28631, n28632,
    n28633, n28634, n28635, n28636, n28637, n28638,
    n28639, n28640, n28641, n28642, n28643, n28644,
    n28645, n28646, n28647, n28648, n28649, n28650,
    n28651, n28652, n28653, n28654, n28655, n28656,
    n28657, n28658, n28659, n28660, n28661, n28662,
    n28663, n28664, n28665, n28666, n28667, n28668,
    n28669, n28670, n28671, n28672, n28673, n28674,
    n28675, n28676, n28677, n28678, n28679, n28680,
    n28681, n28682, n28683, n28684, n28685, n28686,
    n28687, n28688, n28689, n28690, n28691, n28692,
    n28693, n28694, n28695, n28696, n28697, n28698,
    n28699, n28700, n28701, n28702, n28703, n28704,
    n28705, n28706, n28707, n28708, n28709, n28710,
    n28711, n28712, n28713, n28714, n28715, n28716,
    n28717, n28718, n28719, n28720, n28721, n28722,
    n28723, n28724, n28725, n28726, n28727, n28728,
    n28729, n28730, n28731, n28732, n28733, n28734,
    n28735, n28736, n28737, n28738, n28739, n28740,
    n28741, n28742, n28743, n28744, n28745, n28746,
    n28747, n28748, n28749, n28750, n28751, n28752,
    n28753, n28754, n28755, n28756, n28757, n28758,
    n28759, n28760, n28761, n28762, n28763, n28764,
    n28765, n28766, n28767, n28768, n28769, n28770,
    n28771, n28772, n28773, n28774, n28775, n28776,
    n28777, n28778, n28779, n28780, n28781, n28782,
    n28783, n28784, n28785, n28786, n28787, n28788,
    n28789, n28790, n28791, n28792, n28793, n28794,
    n28795, n28796, n28797, n28798, n28799, n28800,
    n28801, n28802, n28803, n28804, n28805, n28806,
    n28807, n28808, n28809, n28810, n28811, n28812,
    n28813, n28814, n28815, n28816, n28817, n28818,
    n28819, n28820, n28821, n28822, n28823, n28824,
    n28825, n28826, n28827, n28828, n28829, n28830,
    n28831, n28832, n28833, n28834, n28835, n28836,
    n28837, n28838, n28839, n28840, n28841, n28842,
    n28843, n28844, n28845, n28846, n28847, n28848,
    n28849, n28850, n28851, n28852, n28853, n28854,
    n28855, n28856, n28857, n28858, n28859, n28860,
    n28861, n28862, n28863, n28864, n28865, n28866,
    n28867, n28868, n28869, n28870, n28871, n28872,
    n28873, n28874, n28875, n28876, n28877, n28878,
    n28879, n28880, n28881, n28882, n28883, n28884,
    n28885, n28886, n28887, n28888, n28889, n28890,
    n28891, n28892, n28894, n28895, n28896, n28897,
    n28898, n28899, n28900, n28901, n28902, n28903,
    n28904, n28905, n28906, n28907, n28908, n28909,
    n28910, n28911, n28912, n28913, n28914, n28915,
    n28916, n28917, n28918, n28919, n28920, n28921,
    n28922, n28923, n28924, n28925, n28926, n28927,
    n28928, n28929, n28930, n28931, n28932, n28933,
    n28934, n28935, n28936, n28937, n28938, n28939,
    n28940, n28941, n28942, n28943, n28944, n28945,
    n28946, n28947, n28948, n28949, n28950, n28951,
    n28952, n28953, n28954, n28955, n28956, n28957,
    n28958, n28959, n28960, n28961, n28962, n28963,
    n28964, n28965, n28966, n28967, n28968, n28969,
    n28970, n28971, n28972, n28973, n28974, n28975,
    n28976, n28977, n28978, n28979, n28980, n28981,
    n28982, n28983, n28984, n28985, n28986, n28987,
    n28988, n28989, n28990, n28991, n28992, n28993,
    n28994, n28995, n28996, n28997, n28998, n28999,
    n29000, n29001, n29002, n29003, n29004, n29005,
    n29006, n29007, n29008, n29009, n29010, n29011,
    n29012, n29013, n29014, n29015, n29016, n29017,
    n29018, n29019, n29020, n29021, n29022, n29023,
    n29024, n29025, n29026, n29027, n29028, n29029,
    n29030, n29031, n29032, n29033, n29034, n29035,
    n29036, n29037, n29038, n29039, n29040, n29041,
    n29042, n29043, n29044, n29045, n29046, n29047,
    n29048, n29049, n29050, n29051, n29052, n29053,
    n29054, n29055, n29056, n29057, n29058, n29059,
    n29060, n29061, n29062, n29063, n29064, n29065,
    n29066, n29067, n29068, n29069, n29070, n29071,
    n29072, n29073, n29074, n29075, n29076, n29077,
    n29078, n29079, n29080, n29081, n29082, n29083,
    n29084, n29085, n29086, n29087, n29088, n29089,
    n29090, n29091, n29092, n29093, n29094, n29095,
    n29096, n29097, n29098, n29099, n29100, n29101,
    n29102, n29103, n29104, n29105, n29106, n29107,
    n29108, n29109, n29110, n29111, n29112, n29113,
    n29114, n29115, n29116, n29117, n29118, n29119,
    n29120, n29121, n29122, n29123, n29124, n29125,
    n29126, n29127, n29128, n29129, n29130, n29131,
    n29132, n29133, n29134, n29135, n29136, n29137,
    n29138, n29139, n29140, n29141, n29142, n29143,
    n29144, n29145, n29146, n29147, n29148, n29149,
    n29150, n29151, n29152, n29153, n29154, n29155,
    n29156, n29157, n29158, n29159, n29160, n29161,
    n29162, n29163, n29164, n29165, n29166, n29167,
    n29168, n29169, n29170, n29171, n29172, n29173,
    n29174, n29175, n29176, n29177, n29178, n29179,
    n29180, n29181, n29182, n29183, n29184, n29185,
    n29186, n29187, n29188, n29189, n29190, n29191,
    n29192, n29193, n29194, n29195, n29196, n29197,
    n29198, n29199, n29200, n29201, n29202, n29203,
    n29204, n29205, n29206, n29207, n29208, n29209,
    n29210, n29211, n29212, n29213, n29214, n29215,
    n29216, n29217, n29218, n29219, n29220, n29221,
    n29222, n29223, n29224, n29225, n29226, n29227,
    n29228, n29229, n29230, n29231, n29232, n29233,
    n29234, n29235, n29236, n29237, n29238, n29239,
    n29240, n29241, n29242, n29243, n29244, n29245,
    n29246, n29247, n29248, n29250, n29251, n29252,
    n29253, n29254, n29255, n29256, n29257, n29258,
    n29259, n29260, n29261, n29262, n29263, n29264,
    n29265, n29266, n29267, n29268, n29269, n29270,
    n29271, n29272, n29273, n29274, n29275, n29276,
    n29277, n29278, n29279, n29280, n29281, n29282,
    n29283, n29284, n29285, n29286, n29287, n29288,
    n29289, n29290, n29291, n29292, n29293, n29294,
    n29295, n29296, n29297, n29298, n29299, n29300,
    n29301, n29302, n29303, n29304, n29305, n29306,
    n29307, n29308, n29309, n29310, n29311, n29312,
    n29313, n29314, n29315, n29316, n29317, n29318,
    n29319, n29320, n29321, n29322, n29323, n29324,
    n29325, n29326, n29327, n29328, n29329, n29330,
    n29331, n29332, n29333, n29334, n29335, n29336,
    n29337, n29338, n29339, n29340, n29341, n29342,
    n29343, n29344, n29345, n29346, n29347, n29348,
    n29349, n29350, n29351, n29352, n29353, n29354,
    n29355, n29356, n29357, n29358, n29359, n29360,
    n29361, n29362, n29363, n29364, n29365, n29366,
    n29367, n29368, n29369, n29370, n29371, n29372,
    n29373, n29374, n29375, n29376, n29377, n29378,
    n29379, n29380, n29381, n29382, n29383, n29384,
    n29385, n29386, n29387, n29388, n29389, n29390,
    n29391, n29392, n29393, n29394, n29395, n29396,
    n29397, n29398, n29399, n29400, n29401, n29402,
    n29403, n29404, n29405, n29406, n29407, n29408,
    n29409, n29410, n29411, n29412, n29413, n29414,
    n29415, n29416, n29417, n29418, n29419, n29420,
    n29421, n29422, n29423, n29424, n29425, n29426,
    n29427, n29428, n29429, n29430, n29431, n29432,
    n29433, n29434, n29435, n29436, n29437, n29438,
    n29439, n29440, n29441, n29442, n29443, n29444,
    n29445, n29446, n29447, n29448, n29449, n29450,
    n29451, n29452, n29453, n29454, n29455, n29456,
    n29457, n29458, n29459, n29460, n29461, n29462,
    n29463, n29464, n29465, n29466, n29467, n29468,
    n29469, n29470, n29471, n29472, n29473, n29474,
    n29475, n29476, n29477, n29478, n29479, n29480,
    n29481, n29482, n29483, n29484, n29485, n29486,
    n29487, n29488, n29489, n29490, n29491, n29492,
    n29493, n29494, n29495, n29496, n29497, n29498,
    n29499, n29500, n29501, n29502, n29503, n29504,
    n29505, n29506, n29507, n29508, n29509, n29510,
    n29511, n29512, n29513, n29514, n29515, n29516,
    n29517, n29518, n29519, n29520, n29521, n29522,
    n29523, n29524, n29525, n29526, n29527, n29528,
    n29529, n29530, n29531, n29532, n29533, n29534,
    n29535, n29536, n29537, n29538, n29539, n29540,
    n29541, n29542, n29543, n29544, n29545, n29546,
    n29547, n29548, n29549, n29550, n29551, n29552,
    n29553, n29554, n29555, n29556, n29557, n29558,
    n29559, n29560, n29561, n29562, n29563, n29564,
    n29565, n29566, n29567, n29568, n29569, n29570,
    n29571, n29572, n29573, n29574, n29575, n29576,
    n29577, n29578, n29579, n29580, n29581, n29582,
    n29583, n29584, n29585, n29586, n29587, n29588,
    n29589, n29590, n29591, n29592, n29593, n29594,
    n29595, n29596, n29597, n29598, n29599, n29600,
    n29601, n29602, n29603, n29604, n29605, n29606,
    n29607, n29608, n29609, n29610, n29611, n29612,
    n29613, n29614, n29615, n29616, n29617, n29618,
    n29619, n29620, n29621, n29622, n29623, n29625,
    n29626, n29627, n29628, n29629, n29630, n29631,
    n29632, n29633, n29634, n29635, n29636, n29637,
    n29638, n29639, n29640, n29641, n29642, n29643,
    n29644, n29645, n29646, n29647, n29648, n29649,
    n29650, n29651, n29652, n29653, n29654, n29655,
    n29656, n29657, n29658, n29659, n29660, n29661,
    n29662, n29663, n29664, n29665, n29666, n29667,
    n29668, n29669, n29670, n29671, n29672, n29673,
    n29674, n29675, n29676, n29677, n29678, n29679,
    n29680, n29681, n29682, n29683, n29684, n29685,
    n29686, n29687, n29688, n29689, n29690, n29691,
    n29692, n29693, n29694, n29695, n29696, n29697,
    n29698, n29699, n29700, n29701, n29702, n29703,
    n29704, n29705, n29706, n29707, n29708, n29709,
    n29710, n29711, n29712, n29713, n29714, n29715,
    n29716, n29717, n29718, n29719, n29720, n29721,
    n29722, n29723, n29724, n29725, n29726, n29727,
    n29728, n29729, n29730, n29731, n29732, n29733,
    n29734, n29735, n29736, n29737, n29738, n29739,
    n29740, n29741, n29742, n29743, n29744, n29745,
    n29746, n29747, n29748, n29749, n29750, n29751,
    n29752, n29753, n29754, n29755, n29756, n29757,
    n29758, n29759, n29760, n29761, n29762, n29763,
    n29764, n29765, n29766, n29767, n29768, n29769,
    n29770, n29771, n29772, n29773, n29774, n29775,
    n29776, n29777, n29778, n29779, n29780, n29781,
    n29782, n29783, n29784, n29785, n29786, n29787,
    n29788, n29789, n29790, n29791, n29792, n29793,
    n29794, n29795, n29796, n29797, n29798, n29799,
    n29800, n29801, n29802, n29803, n29804, n29805,
    n29806, n29807, n29808, n29809, n29810, n29811,
    n29812, n29813, n29814, n29815, n29816, n29817,
    n29818, n29819, n29820, n29821, n29822, n29823,
    n29824, n29825, n29826, n29827, n29828, n29829,
    n29830, n29831, n29832, n29833, n29834, n29835,
    n29836, n29837, n29838, n29839, n29840, n29841,
    n29842, n29843, n29844, n29845, n29846, n29847,
    n29848, n29849, n29850, n29851, n29852, n29853,
    n29854, n29855, n29856, n29857, n29858, n29859,
    n29860, n29861, n29862, n29863, n29864, n29865,
    n29866, n29867, n29868, n29869, n29870, n29871,
    n29872, n29873, n29874, n29875, n29876, n29877,
    n29878, n29879, n29880, n29881, n29882, n29883,
    n29884, n29885, n29886, n29887, n29888, n29889,
    n29890, n29891, n29892, n29893, n29894, n29895,
    n29896, n29897, n29898, n29899, n29900, n29901,
    n29902, n29903, n29904, n29905, n29906, n29907,
    n29908, n29909, n29910, n29911, n29912, n29913,
    n29914, n29915, n29916, n29917, n29918, n29919,
    n29920, n29921, n29922, n29923, n29924, n29925,
    n29926, n29927, n29928, n29929, n29930, n29931,
    n29932, n29933, n29934, n29935, n29936, n29937,
    n29938, n29939, n29940, n29941, n29942, n29943,
    n29944, n29945, n29946, n29947, n29948, n29949,
    n29950, n29951, n29952, n29953, n29954, n29955,
    n29956, n29957, n29958, n29959, n29960, n29961,
    n29962, n29963, n29964, n29965, n29966, n29967,
    n29968, n29969, n29970, n29971, n29972, n29973,
    n29974, n29975, n29976, n29977, n29978, n29979,
    n29980, n29981, n29982, n29983, n29984, n29985,
    n29986, n29987, n29988, n29989, n29990, n29991,
    n29992, n29993, n29994, n29995, n29996, n29997,
    n29998, n29999, n30000, n30001, n30002, n30003,
    n30004, n30005, n30006, n30008, n30009, n30010,
    n30011, n30012, n30013, n30014, n30015, n30016,
    n30017, n30018, n30019, n30020, n30021, n30022,
    n30023, n30024, n30025, n30026, n30027, n30028,
    n30029, n30030, n30031, n30032, n30033, n30034,
    n30035, n30036, n30037, n30038, n30039, n30040,
    n30041, n30042, n30043, n30044, n30045, n30046,
    n30047, n30048, n30049, n30050, n30051, n30052,
    n30053, n30054, n30055, n30056, n30057, n30058,
    n30059, n30060, n30061, n30062, n30063, n30064,
    n30065, n30066, n30067, n30068, n30069, n30070,
    n30071, n30072, n30073, n30074, n30075, n30076,
    n30077, n30078, n30079, n30080, n30081, n30082,
    n30083, n30084, n30085, n30086, n30087, n30088,
    n30089, n30090, n30091, n30092, n30093, n30094,
    n30095, n30096, n30097, n30098, n30099, n30100,
    n30101, n30102, n30103, n30104, n30105, n30106,
    n30107, n30108, n30109, n30110, n30111, n30112,
    n30113, n30114, n30115, n30116, n30117, n30118,
    n30119, n30120, n30121, n30122, n30123, n30124,
    n30125, n30126, n30127, n30128, n30129, n30130,
    n30131, n30132, n30133, n30134, n30135, n30136,
    n30137, n30138, n30139, n30140, n30141, n30142,
    n30143, n30144, n30145, n30146, n30147, n30148,
    n30149, n30150, n30151, n30152, n30153, n30154,
    n30155, n30156, n30157, n30158, n30159, n30160,
    n30161, n30162, n30163, n30164, n30165, n30166,
    n30167, n30168, n30169, n30170, n30171, n30172,
    n30173, n30174, n30175, n30176, n30177, n30178,
    n30179, n30180, n30181, n30182, n30183, n30184,
    n30185, n30186, n30187, n30188, n30189, n30190,
    n30191, n30192, n30193, n30194, n30195, n30196,
    n30197, n30198, n30199, n30200, n30201, n30202,
    n30203, n30204, n30205, n30206, n30207, n30208,
    n30209, n30210, n30211, n30212, n30213, n30214,
    n30215, n30216, n30217, n30218, n30219, n30220,
    n30221, n30222, n30223, n30224, n30225, n30226,
    n30227, n30228, n30229, n30230, n30231, n30232,
    n30233, n30234, n30235, n30236, n30237, n30238,
    n30239, n30240, n30241, n30242, n30243, n30244,
    n30245, n30246, n30247, n30248, n30249, n30250,
    n30251, n30252, n30253, n30254, n30255, n30256,
    n30257, n30258, n30259, n30260, n30261, n30262,
    n30263, n30264, n30265, n30266, n30267, n30268,
    n30269, n30270, n30271, n30272, n30273, n30274,
    n30275, n30276, n30277, n30278, n30279, n30280,
    n30281, n30282, n30283, n30284, n30285, n30286,
    n30287, n30288, n30289, n30290, n30291, n30292,
    n30293, n30294, n30295, n30296, n30297, n30298,
    n30299, n30300, n30301, n30302, n30303, n30304,
    n30305, n30306, n30307, n30308, n30309, n30310,
    n30311, n30312, n30313, n30314, n30315, n30316,
    n30317, n30318, n30319, n30320, n30321, n30322,
    n30323, n30324, n30325, n30326, n30327, n30328,
    n30329, n30330, n30331, n30332, n30333, n30334,
    n30335, n30336, n30337, n30338, n30339, n30340,
    n30341, n30342, n30343, n30344, n30345, n30346,
    n30347, n30348, n30350, n30351, n30352, n30353,
    n30354, n30355, n30356, n30357, n30358, n30359,
    n30360, n30361, n30362, n30363, n30364, n30365,
    n30366, n30367, n30368, n30369, n30370, n30371,
    n30372, n30373, n30374, n30375, n30376, n30377,
    n30378, n30379, n30380, n30381, n30382, n30383,
    n30384, n30385, n30386, n30387, n30388, n30389,
    n30390, n30391, n30392, n30393, n30394, n30395,
    n30396, n30397, n30398, n30399, n30400, n30401,
    n30402, n30403, n30404, n30405, n30406, n30407,
    n30408, n30409, n30410, n30411, n30412, n30413,
    n30414, n30415, n30416, n30417, n30418, n30419,
    n30420, n30421, n30422, n30423, n30424, n30425,
    n30426, n30427, n30428, n30429, n30430, n30431,
    n30432, n30433, n30434, n30435, n30436, n30437,
    n30438, n30439, n30440, n30441, n30442, n30443,
    n30444, n30445, n30446, n30447, n30448, n30449,
    n30450, n30451, n30452, n30453, n30454, n30455,
    n30456, n30457, n30458, n30459, n30460, n30461,
    n30462, n30463, n30464, n30465, n30466, n30467,
    n30468, n30469, n30470, n30471, n30472, n30473,
    n30474, n30475, n30476, n30477, n30478, n30479,
    n30480, n30481, n30482, n30483, n30484, n30485,
    n30486, n30487, n30488, n30489, n30490, n30491,
    n30492, n30493, n30494, n30495, n30496, n30497,
    n30498, n30499, n30500, n30501, n30502, n30503,
    n30504, n30505, n30506, n30507, n30508, n30509,
    n30510, n30511, n30512, n30513, n30514, n30515,
    n30516, n30517, n30518, n30519, n30520, n30521,
    n30522, n30523, n30524, n30525, n30526, n30527,
    n30528, n30529, n30530, n30531, n30532, n30533,
    n30534, n30535, n30536, n30537, n30538, n30539,
    n30540, n30541, n30542, n30543, n30544, n30545,
    n30546, n30547, n30548, n30549, n30550, n30551,
    n30552, n30553, n30554, n30555, n30556, n30557,
    n30558, n30559, n30560, n30561, n30562, n30563,
    n30564, n30565, n30566, n30567, n30568, n30569,
    n30570, n30571, n30572, n30573, n30574, n30575,
    n30576, n30577, n30578, n30579, n30580, n30581,
    n30582, n30583, n30584, n30585, n30586, n30587,
    n30588, n30589, n30590, n30591, n30592, n30593,
    n30594, n30595, n30596, n30597, n30598, n30599,
    n30600, n30601, n30602, n30603, n30604, n30605,
    n30606, n30607, n30608, n30609, n30610, n30611,
    n30612, n30613, n30614, n30615, n30616, n30617,
    n30618, n30619, n30620, n30621, n30622, n30623,
    n30624, n30625, n30626, n30627, n30628, n30629,
    n30630, n30631, n30632, n30633, n30634, n30635,
    n30636, n30637, n30638, n30639, n30640, n30641,
    n30642, n30643, n30644, n30645, n30646, n30647,
    n30648, n30649, n30650, n30651, n30652, n30653,
    n30654, n30655, n30656, n30657, n30658, n30659,
    n30660, n30661, n30662, n30663, n30664, n30665,
    n30666, n30667, n30668, n30669, n30670, n30671,
    n30672, n30673, n30674, n30675, n30676, n30677,
    n30678, n30679, n30681, n30682, n30683, n30684,
    n30685, n30686, n30687, n30688, n30689, n30690,
    n30691, n30692, n30693, n30694, n30695, n30696,
    n30697, n30698, n30699, n30700, n30701, n30702,
    n30703, n30704, n30705, n30706, n30707, n30708,
    n30709, n30710, n30711, n30712, n30713, n30714,
    n30715, n30716, n30717, n30718, n30719, n30720,
    n30721, n30722, n30723, n30724, n30725, n30726,
    n30727, n30728, n30729, n30730, n30731, n30732,
    n30733, n30734, n30735, n30736, n30737, n30738,
    n30739, n30740, n30741, n30742, n30743, n30744,
    n30745, n30746, n30747, n30748, n30749, n30750,
    n30751, n30752, n30753, n30754, n30755, n30756,
    n30757, n30758, n30759, n30760, n30761, n30762,
    n30763, n30764, n30765, n30766, n30767, n30768,
    n30769, n30770, n30771, n30772, n30773, n30774,
    n30775, n30776, n30777, n30778, n30779, n30780,
    n30781, n30782, n30783, n30784, n30785, n30786,
    n30787, n30788, n30789, n30790, n30791, n30792,
    n30793, n30794, n30795, n30796, n30797, n30798,
    n30799, n30800, n30801, n30802, n30803, n30804,
    n30805, n30806, n30807, n30808, n30809, n30810,
    n30811, n30812, n30813, n30814, n30815, n30816,
    n30817, n30818, n30819, n30820, n30821, n30822,
    n30823, n30824, n30825, n30826, n30827, n30828,
    n30829, n30830, n30831, n30832, n30833, n30834,
    n30835, n30836, n30837, n30838, n30839, n30840,
    n30841, n30842, n30843, n30844, n30845, n30846,
    n30847, n30848, n30849, n30850, n30851, n30852,
    n30853, n30854, n30855, n30856, n30857, n30858,
    n30859, n30860, n30861, n30862, n30863, n30864,
    n30865, n30866, n30867, n30868, n30869, n30870,
    n30871, n30872, n30873, n30874, n30875, n30876,
    n30877, n30878, n30879, n30880, n30881, n30882,
    n30883, n30884, n30885, n30886, n30887, n30888,
    n30889, n30890, n30891, n30892, n30893, n30894,
    n30895, n30896, n30897, n30898, n30899, n30900,
    n30901, n30902, n30903, n30904, n30905, n30906,
    n30907, n30908, n30909, n30910, n30911, n30912,
    n30913, n30914, n30915, n30916, n30917, n30918,
    n30919, n30920, n30921, n30922, n30923, n30924,
    n30925, n30926, n30927, n30928, n30929, n30930,
    n30931, n30932, n30933, n30934, n30935, n30936,
    n30937, n30938, n30939, n30940, n30941, n30942,
    n30943, n30944, n30945, n30946, n30947, n30948,
    n30949, n30950, n30951, n30952, n30953, n30954,
    n30955, n30956, n30957, n30958, n30959, n30960,
    n30961, n30962, n30963, n30964, n30965, n30966,
    n30967, n30968, n30969, n30970, n30971, n30972,
    n30973, n30974, n30975, n30976, n30977, n30978,
    n30979, n30980, n30981, n30982, n30983, n30984,
    n30985, n30986, n30987, n30988, n30989, n30990,
    n30991, n30992, n30993, n30994, n30995, n30996,
    n30997, n30998, n30999, n31000, n31001, n31002,
    n31003, n31004, n31005, n31006, n31007, n31008,
    n31009, n31010, n31011, n31012, n31013, n31014,
    n31015, n31016, n31017, n31018, n31019, n31020,
    n31021, n31023, n31024, n31025, n31026, n31027,
    n31028, n31029, n31030, n31031, n31032, n31033,
    n31034, n31035, n31036, n31037, n31038, n31039,
    n31040, n31041, n31042, n31043, n31044, n31045,
    n31046, n31047, n31048, n31049, n31050, n31051,
    n31052, n31053, n31054, n31055, n31056, n31057,
    n31058, n31059, n31060, n31061, n31062, n31063,
    n31064, n31065, n31066, n31067, n31068, n31069,
    n31070, n31071, n31072, n31073, n31074, n31075,
    n31076, n31077, n31078, n31079, n31080, n31081,
    n31082, n31083, n31084, n31085, n31086, n31087,
    n31088, n31089, n31090, n31091, n31092, n31093,
    n31094, n31095, n31096, n31097, n31098, n31099,
    n31100, n31101, n31102, n31103, n31104, n31105,
    n31106, n31107, n31108, n31109, n31110, n31111,
    n31112, n31113, n31114, n31115, n31116, n31117,
    n31118, n31119, n31120, n31121, n31122, n31123,
    n31124, n31125, n31126, n31127, n31128, n31129,
    n31130, n31131, n31132, n31133, n31134, n31135,
    n31136, n31137, n31138, n31139, n31140, n31141,
    n31142, n31143, n31144, n31145, n31146, n31147,
    n31148, n31149, n31150, n31151, n31152, n31153,
    n31154, n31155, n31156, n31157, n31158, n31159,
    n31160, n31161, n31162, n31163, n31164, n31165,
    n31166, n31167, n31168, n31169, n31170, n31171,
    n31172, n31173, n31174, n31175, n31176, n31177,
    n31178, n31179, n31180, n31181, n31182, n31183,
    n31184, n31185, n31186, n31187, n31188, n31189,
    n31190, n31191, n31192, n31193, n31194, n31195,
    n31196, n31197, n31198, n31199, n31200, n31201,
    n31202, n31203, n31204, n31205, n31206, n31207,
    n31208, n31209, n31210, n31211, n31212, n31213,
    n31214, n31215, n31216, n31217, n31218, n31219,
    n31220, n31221, n31222, n31223, n31224, n31225,
    n31226, n31227, n31228, n31229, n31230, n31231,
    n31232, n31233, n31234, n31235, n31236, n31237,
    n31238, n31239, n31240, n31241, n31242, n31243,
    n31244, n31245, n31246, n31247, n31248, n31249,
    n31250, n31251, n31252, n31253, n31254, n31255,
    n31256, n31257, n31258, n31259, n31260, n31261,
    n31262, n31263, n31264, n31265, n31266, n31267,
    n31268, n31269, n31270, n31271, n31272, n31273,
    n31274, n31275, n31276, n31277, n31278, n31279,
    n31280, n31281, n31282, n31283, n31284, n31285,
    n31286, n31287, n31288, n31289, n31290, n31291,
    n31292, n31293, n31294, n31295, n31296, n31297,
    n31298, n31299, n31300, n31301, n31302, n31303,
    n31304, n31305, n31306, n31307, n31308, n31309,
    n31310, n31311, n31312, n31313, n31314, n31315,
    n31316, n31317, n31318, n31319, n31320, n31321,
    n31322, n31323, n31324, n31325, n31326, n31327,
    n31328, n31329, n31330, n31331, n31332, n31333,
    n31334, n31336, n31337, n31338, n31339, n31340,
    n31341, n31342, n31343, n31344, n31345, n31346,
    n31347, n31348, n31349, n31350, n31351, n31352,
    n31353, n31354, n31355, n31356, n31357, n31358,
    n31359, n31360, n31361, n31362, n31363, n31364,
    n31365, n31366, n31367, n31368, n31369, n31370,
    n31371, n31372, n31373, n31374, n31375, n31376,
    n31377, n31378, n31379, n31380, n31381, n31382,
    n31383, n31384, n31385, n31386, n31387, n31388,
    n31389, n31390, n31391, n31392, n31393, n31394,
    n31395, n31396, n31397, n31398, n31399, n31400,
    n31401, n31402, n31403, n31404, n31405, n31406,
    n31407, n31408, n31409, n31410, n31411, n31412,
    n31413, n31414, n31415, n31416, n31417, n31418,
    n31419, n31420, n31421, n31422, n31423, n31424,
    n31425, n31426, n31427, n31428, n31429, n31430,
    n31431, n31432, n31433, n31434, n31435, n31436,
    n31437, n31438, n31439, n31440, n31441, n31442,
    n31443, n31444, n31445, n31446, n31447, n31448,
    n31449, n31450, n31451, n31452, n31453, n31454,
    n31455, n31456, n31457, n31458, n31459, n31460,
    n31461, n31462, n31463, n31464, n31465, n31466,
    n31467, n31468, n31469, n31470, n31471, n31472,
    n31473, n31474, n31475, n31476, n31477, n31478,
    n31479, n31480, n31481, n31482, n31483, n31484,
    n31485, n31486, n31487, n31488, n31489, n31490,
    n31491, n31492, n31493, n31494, n31495, n31496,
    n31497, n31498, n31499, n31500, n31501, n31502,
    n31503, n31504, n31505, n31506, n31507, n31508,
    n31509, n31510, n31511, n31512, n31513, n31514,
    n31515, n31516, n31517, n31518, n31519, n31520,
    n31521, n31522, n31523, n31524, n31525, n31526,
    n31527, n31528, n31529, n31530, n31531, n31532,
    n31533, n31534, n31535, n31536, n31537, n31538,
    n31539, n31540, n31541, n31542, n31543, n31544,
    n31545, n31546, n31547, n31548, n31549, n31550,
    n31551, n31552, n31553, n31554, n31555, n31556,
    n31557, n31558, n31559, n31560, n31561, n31562,
    n31563, n31564, n31565, n31566, n31567, n31568,
    n31569, n31570, n31571, n31572, n31573, n31574,
    n31575, n31576, n31577, n31578, n31579, n31580,
    n31581, n31582, n31583, n31584, n31585, n31586,
    n31587, n31588, n31589, n31590, n31591, n31592,
    n31593, n31594, n31595, n31596, n31597, n31598,
    n31599, n31600, n31601, n31602, n31603, n31604,
    n31605, n31606, n31607, n31608, n31609, n31610,
    n31611, n31612, n31613, n31614, n31615, n31616,
    n31617, n31618, n31619, n31620, n31621, n31622,
    n31623, n31624, n31625, n31626, n31627, n31628,
    n31629, n31630, n31631, n31632, n31633, n31634,
    n31635, n31636, n31637, n31638, n31639, n31640,
    n31641, n31642, n31643, n31644, n31645, n31646,
    n31647, n31648, n31649, n31650, n31651, n31652,
    n31653, n31654, n31655, n31656, n31658, n31659,
    n31660, n31661, n31662, n31663, n31664, n31665,
    n31666, n31667, n31668, n31669, n31670, n31671,
    n31672, n31673, n31674, n31675, n31676, n31677,
    n31678, n31679, n31680, n31681, n31682, n31683,
    n31684, n31685, n31686, n31687, n31688, n31689,
    n31690, n31691, n31692, n31693, n31694, n31695,
    n31696, n31697, n31698, n31699, n31700, n31701,
    n31702, n31703, n31704, n31705, n31706, n31707,
    n31708, n31709, n31710, n31711, n31712, n31713,
    n31714, n31715, n31716, n31717, n31718, n31719,
    n31720, n31721, n31722, n31723, n31724, n31725,
    n31726, n31727, n31728, n31729, n31730, n31731,
    n31732, n31733, n31734, n31735, n31736, n31737,
    n31738, n31739, n31740, n31741, n31742, n31743,
    n31744, n31745, n31746, n31747, n31748, n31749,
    n31750, n31751, n31752, n31753, n31754, n31755,
    n31756, n31757, n31758, n31759, n31760, n31761,
    n31762, n31763, n31764, n31765, n31766, n31767,
    n31768, n31769, n31770, n31771, n31772, n31773,
    n31774, n31775, n31776, n31777, n31778, n31779,
    n31780, n31781, n31782, n31783, n31784, n31785,
    n31786, n31787, n31788, n31789, n31790, n31791,
    n31792, n31793, n31794, n31795, n31796, n31797,
    n31798, n31799, n31800, n31801, n31802, n31803,
    n31804, n31805, n31806, n31807, n31808, n31809,
    n31810, n31811, n31812, n31813, n31814, n31815,
    n31816, n31817, n31818, n31819, n31820, n31821,
    n31822, n31823, n31824, n31825, n31826, n31827,
    n31828, n31829, n31830, n31831, n31832, n31833,
    n31834, n31835, n31836, n31837, n31838, n31839,
    n31840, n31841, n31842, n31843, n31844, n31845,
    n31846, n31847, n31848, n31849, n31850, n31851,
    n31852, n31853, n31854, n31855, n31856, n31857,
    n31858, n31859, n31860, n31861, n31862, n31863,
    n31864, n31865, n31866, n31867, n31868, n31869,
    n31870, n31871, n31872, n31873, n31874, n31875,
    n31876, n31877, n31878, n31879, n31880, n31881,
    n31882, n31883, n31884, n31885, n31886, n31887,
    n31888, n31889, n31890, n31891, n31892, n31893,
    n31894, n31895, n31896, n31897, n31898, n31899,
    n31900, n31901, n31902, n31903, n31904, n31905,
    n31906, n31907, n31908, n31909, n31910, n31911,
    n31912, n31913, n31914, n31915, n31916, n31917,
    n31918, n31919, n31920, n31921, n31922, n31923,
    n31924, n31925, n31926, n31927, n31928, n31929,
    n31930, n31931, n31932, n31933, n31934, n31935,
    n31936, n31937, n31938, n31939, n31940, n31941,
    n31942, n31943, n31944, n31945, n31946, n31947,
    n31948, n31949, n31950, n31951, n31952, n31953,
    n31954, n31955, n31956, n31957, n31958, n31959,
    n31960, n31961, n31962, n31963, n31964, n31965,
    n31966, n31967, n31968, n31969, n31970, n31971,
    n31972, n31973, n31974, n31975, n31976, n31977,
    n31978, n31980, n31981, n31982, n31983, n31984,
    n31985, n31986, n31987, n31988, n31989, n31990,
    n31991, n31992, n31993, n31994, n31995, n31996,
    n31997, n31998, n31999, n32000, n32001, n32002,
    n32003, n32004, n32005, n32006, n32007, n32008,
    n32009, n32010, n32011, n32012, n32013, n32014,
    n32015, n32016, n32017, n32018, n32019, n32020,
    n32021, n32022, n32023, n32024, n32025, n32026,
    n32027, n32028, n32029, n32030, n32031, n32032,
    n32033, n32034, n32035, n32036, n32037, n32038,
    n32039, n32040, n32041, n32042, n32043, n32044,
    n32045, n32046, n32047, n32048, n32049, n32050,
    n32051, n32052, n32053, n32054, n32055, n32056,
    n32057, n32058, n32059, n32060, n32061, n32062,
    n32063, n32064, n32065, n32066, n32067, n32068,
    n32069, n32070, n32071, n32072, n32073, n32074,
    n32075, n32076, n32077, n32078, n32079, n32080,
    n32081, n32082, n32083, n32084, n32085, n32086,
    n32087, n32088, n32089, n32090, n32091, n32092,
    n32093, n32094, n32095, n32096, n32097, n32098,
    n32099, n32100, n32101, n32102, n32103, n32104,
    n32105, n32106, n32107, n32108, n32109, n32110,
    n32111, n32112, n32113, n32114, n32115, n32116,
    n32117, n32118, n32119, n32120, n32121, n32122,
    n32123, n32124, n32125, n32126, n32127, n32128,
    n32129, n32130, n32131, n32132, n32133, n32134,
    n32135, n32136, n32137, n32138, n32139, n32140,
    n32141, n32142, n32143, n32144, n32145, n32146,
    n32147, n32148, n32149, n32150, n32151, n32152,
    n32153, n32154, n32155, n32156, n32157, n32158,
    n32159, n32160, n32161, n32162, n32163, n32164,
    n32165, n32166, n32167, n32168, n32169, n32170,
    n32171, n32172, n32173, n32174, n32175, n32176,
    n32177, n32178, n32179, n32180, n32181, n32182,
    n32183, n32184, n32185, n32186, n32187, n32188,
    n32189, n32190, n32191, n32192, n32193, n32194,
    n32195, n32196, n32197, n32198, n32199, n32200,
    n32201, n32202, n32203, n32204, n32205, n32206,
    n32207, n32208, n32209, n32210, n32211, n32212,
    n32213, n32214, n32215, n32216, n32217, n32218,
    n32219, n32220, n32221, n32222, n32223, n32224,
    n32225, n32226, n32227, n32228, n32229, n32230,
    n32231, n32232, n32233, n32234, n32235, n32236,
    n32237, n32238, n32239, n32240, n32241, n32242,
    n32243, n32244, n32245, n32246, n32247, n32248,
    n32249, n32250, n32251, n32252, n32253, n32254,
    n32255, n32256, n32257, n32258, n32259, n32260,
    n32261, n32262, n32263, n32264, n32265, n32267,
    n32268, n32269, n32270, n32271, n32272, n32273,
    n32274, n32275, n32276, n32277, n32278, n32279,
    n32280, n32281, n32282, n32283, n32284, n32285,
    n32286, n32287, n32288, n32289, n32290, n32291,
    n32292, n32293, n32294, n32295, n32296, n32297,
    n32298, n32299, n32300, n32301, n32302, n32303,
    n32304, n32305, n32306, n32307, n32308, n32309,
    n32310, n32311, n32312, n32313, n32314, n32315,
    n32316, n32317, n32318, n32319, n32320, n32321,
    n32322, n32323, n32324, n32325, n32326, n32327,
    n32328, n32329, n32330, n32331, n32332, n32333,
    n32334, n32335, n32336, n32337, n32338, n32339,
    n32340, n32341, n32342, n32343, n32344, n32345,
    n32346, n32347, n32348, n32349, n32350, n32351,
    n32352, n32353, n32354, n32355, n32356, n32357,
    n32358, n32359, n32360, n32361, n32362, n32363,
    n32364, n32365, n32366, n32367, n32368, n32369,
    n32370, n32371, n32372, n32373, n32374, n32375,
    n32376, n32377, n32378, n32379, n32380, n32381,
    n32382, n32383, n32384, n32385, n32386, n32387,
    n32388, n32389, n32390, n32391, n32392, n32393,
    n32394, n32395, n32396, n32397, n32398, n32399,
    n32400, n32401, n32402, n32403, n32404, n32405,
    n32406, n32407, n32408, n32409, n32410, n32411,
    n32412, n32413, n32414, n32415, n32416, n32417,
    n32418, n32419, n32420, n32421, n32422, n32423,
    n32424, n32425, n32426, n32427, n32428, n32429,
    n32430, n32431, n32432, n32433, n32434, n32435,
    n32436, n32437, n32438, n32439, n32440, n32441,
    n32442, n32443, n32444, n32445, n32446, n32447,
    n32448, n32449, n32450, n32451, n32452, n32453,
    n32454, n32455, n32456, n32457, n32458, n32459,
    n32460, n32461, n32462, n32463, n32464, n32465,
    n32466, n32467, n32468, n32469, n32470, n32471,
    n32472, n32473, n32474, n32475, n32476, n32477,
    n32478, n32479, n32480, n32481, n32482, n32483,
    n32484, n32485, n32486, n32487, n32488, n32489,
    n32490, n32491, n32492, n32493, n32494, n32495,
    n32496, n32497, n32498, n32499, n32500, n32501,
    n32502, n32503, n32504, n32505, n32506, n32507,
    n32508, n32509, n32510, n32511, n32512, n32513,
    n32514, n32515, n32516, n32517, n32518, n32519,
    n32520, n32521, n32522, n32523, n32524, n32525,
    n32526, n32527, n32528, n32529, n32530, n32531,
    n32532, n32533, n32534, n32535, n32536, n32537,
    n32538, n32539, n32540, n32541, n32542, n32543,
    n32544, n32545, n32546, n32547, n32548, n32549,
    n32550, n32551, n32552, n32553, n32554, n32555,
    n32556, n32557, n32558, n32559, n32560, n32561,
    n32562, n32563, n32565, n32566, n32567, n32568,
    n32569, n32570, n32571, n32572, n32573, n32574,
    n32575, n32576, n32577, n32578, n32579, n32580,
    n32581, n32582, n32583, n32584, n32585, n32586,
    n32587, n32588, n32589, n32590, n32591, n32592,
    n32593, n32594, n32595, n32596, n32597, n32598,
    n32599, n32600, n32601, n32602, n32603, n32604,
    n32605, n32606, n32607, n32608, n32609, n32610,
    n32611, n32612, n32613, n32614, n32615, n32616,
    n32617, n32618, n32619, n32620, n32621, n32622,
    n32623, n32624, n32625, n32626, n32627, n32628,
    n32629, n32630, n32631, n32632, n32633, n32634,
    n32635, n32636, n32637, n32638, n32639, n32640,
    n32641, n32642, n32643, n32644, n32645, n32646,
    n32647, n32648, n32649, n32650, n32651, n32652,
    n32653, n32654, n32655, n32656, n32657, n32658,
    n32659, n32660, n32661, n32662, n32663, n32664,
    n32665, n32666, n32667, n32668, n32669, n32670,
    n32671, n32672, n32673, n32674, n32675, n32676,
    n32677, n32678, n32679, n32680, n32681, n32682,
    n32683, n32684, n32685, n32686, n32687, n32688,
    n32689, n32690, n32691, n32692, n32693, n32694,
    n32695, n32696, n32697, n32698, n32699, n32700,
    n32701, n32702, n32703, n32704, n32705, n32706,
    n32707, n32708, n32709, n32710, n32711, n32712,
    n32713, n32714, n32715, n32716, n32717, n32718,
    n32719, n32720, n32721, n32722, n32723, n32724,
    n32725, n32726, n32727, n32728, n32729, n32730,
    n32731, n32732, n32733, n32734, n32735, n32736,
    n32737, n32738, n32739, n32740, n32741, n32742,
    n32743, n32744, n32745, n32746, n32747, n32748,
    n32749, n32750, n32751, n32752, n32753, n32754,
    n32755, n32756, n32757, n32758, n32759, n32760,
    n32761, n32762, n32763, n32764, n32765, n32766,
    n32767, n32768, n32769, n32770, n32771, n32772,
    n32773, n32774, n32775, n32776, n32777, n32778,
    n32779, n32780, n32781, n32782, n32783, n32784,
    n32785, n32786, n32787, n32788, n32789, n32790,
    n32791, n32792, n32793, n32794, n32795, n32796,
    n32797, n32798, n32799, n32800, n32801, n32802,
    n32803, n32804, n32805, n32806, n32807, n32808,
    n32809, n32810, n32811, n32812, n32813, n32814,
    n32815, n32816, n32817, n32818, n32819, n32820,
    n32821, n32822, n32823, n32824, n32825, n32826,
    n32827, n32828, n32829, n32830, n32831, n32832,
    n32833, n32834, n32835, n32836, n32837, n32838,
    n32839, n32840, n32841, n32842, n32843, n32844,
    n32845, n32846, n32847, n32848, n32849, n32850,
    n32851, n32852, n32853, n32854, n32855, n32856,
    n32857, n32858, n32859, n32860, n32862, n32863,
    n32864, n32865, n32866, n32867, n32868, n32869,
    n32870, n32871, n32872, n32873, n32874, n32875,
    n32876, n32877, n32878, n32879, n32880, n32881,
    n32882, n32883, n32884, n32885, n32886, n32887,
    n32888, n32889, n32890, n32891, n32892, n32893,
    n32894, n32895, n32896, n32897, n32898, n32899,
    n32900, n32901, n32902, n32903, n32904, n32905,
    n32906, n32907, n32908, n32909, n32910, n32911,
    n32912, n32913, n32914, n32915, n32916, n32917,
    n32918, n32919, n32920, n32921, n32922, n32923,
    n32924, n32925, n32926, n32927, n32928, n32929,
    n32930, n32931, n32932, n32933, n32934, n32935,
    n32936, n32937, n32938, n32939, n32940, n32941,
    n32942, n32943, n32944, n32945, n32946, n32947,
    n32948, n32949, n32950, n32951, n32952, n32953,
    n32954, n32955, n32956, n32957, n32958, n32959,
    n32960, n32961, n32962, n32963, n32964, n32965,
    n32966, n32967, n32968, n32969, n32970, n32971,
    n32972, n32973, n32974, n32975, n32976, n32977,
    n32978, n32979, n32980, n32981, n32982, n32983,
    n32984, n32985, n32986, n32987, n32988, n32989,
    n32990, n32991, n32992, n32993, n32994, n32995,
    n32996, n32997, n32998, n32999, n33000, n33001,
    n33002, n33003, n33004, n33005, n33006, n33007,
    n33008, n33009, n33010, n33011, n33012, n33013,
    n33014, n33015, n33016, n33017, n33018, n33019,
    n33020, n33021, n33022, n33023, n33024, n33025,
    n33026, n33027, n33028, n33029, n33030, n33031,
    n33032, n33033, n33034, n33035, n33036, n33037,
    n33038, n33039, n33040, n33041, n33042, n33043,
    n33044, n33045, n33046, n33047, n33048, n33049,
    n33050, n33051, n33052, n33053, n33054, n33055,
    n33056, n33057, n33058, n33059, n33060, n33061,
    n33062, n33063, n33064, n33065, n33066, n33067,
    n33068, n33069, n33070, n33071, n33072, n33073,
    n33074, n33075, n33076, n33077, n33078, n33079,
    n33080, n33081, n33082, n33083, n33084, n33085,
    n33086, n33087, n33088, n33089, n33090, n33091,
    n33092, n33093, n33094, n33095, n33096, n33097,
    n33098, n33099, n33100, n33101, n33102, n33103,
    n33104, n33105, n33106, n33107, n33108, n33109,
    n33110, n33111, n33112, n33113, n33114, n33115,
    n33116, n33117, n33118, n33119, n33120, n33122,
    n33123, n33124, n33125, n33126, n33127, n33128,
    n33129, n33130, n33131, n33132, n33133, n33134,
    n33135, n33136, n33137, n33138, n33139, n33140,
    n33141, n33142, n33143, n33144, n33145, n33146,
    n33147, n33148, n33149, n33150, n33151, n33152,
    n33153, n33154, n33155, n33156, n33157, n33158,
    n33159, n33160, n33161, n33162, n33163, n33164,
    n33165, n33166, n33167, n33168, n33169, n33170,
    n33171, n33172, n33173, n33174, n33175, n33176,
    n33177, n33178, n33179, n33180, n33181, n33182,
    n33183, n33184, n33185, n33186, n33187, n33188,
    n33189, n33190, n33191, n33192, n33193, n33194,
    n33195, n33196, n33197, n33198, n33199, n33200,
    n33201, n33202, n33203, n33204, n33205, n33206,
    n33207, n33208, n33209, n33210, n33211, n33212,
    n33213, n33214, n33215, n33216, n33217, n33218,
    n33219, n33220, n33221, n33222, n33223, n33224,
    n33225, n33226, n33227, n33228, n33229, n33230,
    n33231, n33232, n33233, n33234, n33235, n33236,
    n33237, n33238, n33239, n33240, n33241, n33242,
    n33243, n33244, n33245, n33246, n33247, n33248,
    n33249, n33250, n33251, n33252, n33253, n33254,
    n33255, n33256, n33257, n33258, n33259, n33260,
    n33261, n33262, n33263, n33264, n33265, n33266,
    n33267, n33268, n33269, n33270, n33271, n33272,
    n33273, n33274, n33275, n33276, n33277, n33278,
    n33279, n33280, n33281, n33282, n33283, n33284,
    n33285, n33286, n33287, n33288, n33289, n33290,
    n33291, n33292, n33293, n33294, n33295, n33296,
    n33297, n33298, n33299, n33300, n33301, n33302,
    n33303, n33304, n33305, n33306, n33307, n33308,
    n33309, n33310, n33311, n33312, n33313, n33314,
    n33315, n33316, n33317, n33318, n33319, n33320,
    n33321, n33322, n33323, n33324, n33325, n33326,
    n33327, n33328, n33329, n33330, n33331, n33332,
    n33333, n33334, n33335, n33336, n33337, n33338,
    n33339, n33340, n33341, n33342, n33343, n33344,
    n33345, n33346, n33347, n33348, n33349, n33350,
    n33351, n33352, n33353, n33354, n33355, n33356,
    n33357, n33358, n33359, n33360, n33361, n33362,
    n33363, n33364, n33365, n33366, n33367, n33368,
    n33369, n33370, n33371, n33372, n33373, n33374,
    n33375, n33376, n33377, n33378, n33379, n33380,
    n33381, n33382, n33383, n33384, n33385, n33386,
    n33387, n33388, n33389, n33390, n33391, n33393,
    n33394, n33395, n33396, n33397, n33398, n33399,
    n33400, n33401, n33402, n33403, n33404, n33405,
    n33406, n33407, n33408, n33409, n33410, n33411,
    n33412, n33413, n33414, n33415, n33416, n33417,
    n33418, n33419, n33420, n33421, n33422, n33423,
    n33424, n33425, n33426, n33427, n33428, n33429,
    n33430, n33431, n33432, n33433, n33434, n33435,
    n33436, n33437, n33438, n33439, n33440, n33441,
    n33442, n33443, n33444, n33445, n33446, n33447,
    n33448, n33449, n33450, n33451, n33452, n33453,
    n33454, n33455, n33456, n33457, n33458, n33459,
    n33460, n33461, n33462, n33463, n33464, n33465,
    n33466, n33467, n33468, n33469, n33470, n33471,
    n33472, n33473, n33474, n33475, n33476, n33477,
    n33478, n33479, n33480, n33481, n33482, n33483,
    n33484, n33485, n33486, n33487, n33488, n33489,
    n33490, n33491, n33492, n33493, n33494, n33495,
    n33496, n33497, n33498, n33499, n33500, n33501,
    n33502, n33503, n33504, n33505, n33506, n33507,
    n33508, n33509, n33510, n33511, n33512, n33513,
    n33514, n33515, n33516, n33517, n33518, n33519,
    n33520, n33521, n33522, n33523, n33524, n33525,
    n33526, n33527, n33528, n33529, n33530, n33531,
    n33532, n33533, n33534, n33535, n33536, n33537,
    n33538, n33539, n33540, n33541, n33542, n33543,
    n33544, n33545, n33546, n33547, n33548, n33549,
    n33550, n33551, n33552, n33553, n33554, n33555,
    n33556, n33557, n33558, n33559, n33560, n33561,
    n33562, n33563, n33564, n33565, n33566, n33567,
    n33568, n33569, n33570, n33571, n33572, n33573,
    n33574, n33575, n33576, n33577, n33578, n33579,
    n33580, n33581, n33582, n33583, n33584, n33585,
    n33586, n33587, n33588, n33589, n33590, n33591,
    n33592, n33593, n33594, n33595, n33596, n33597,
    n33598, n33599, n33600, n33601, n33602, n33603,
    n33604, n33605, n33606, n33607, n33608, n33609,
    n33610, n33611, n33612, n33613, n33614, n33615,
    n33616, n33617, n33618, n33619, n33620, n33621,
    n33622, n33623, n33624, n33625, n33626, n33627,
    n33628, n33629, n33630, n33631, n33632, n33633,
    n33634, n33635, n33636, n33637, n33638, n33639,
    n33640, n33641, n33642, n33643, n33644, n33645,
    n33646, n33647, n33648, n33649, n33651, n33652,
    n33653, n33654, n33655, n33656, n33657, n33658,
    n33659, n33660, n33661, n33662, n33663, n33664,
    n33665, n33666, n33667, n33668, n33669, n33670,
    n33671, n33672, n33673, n33674, n33675, n33676,
    n33677, n33678, n33679, n33680, n33681, n33682,
    n33683, n33684, n33685, n33686, n33687, n33688,
    n33689, n33690, n33691, n33692, n33693, n33694,
    n33695, n33696, n33697, n33698, n33699, n33700,
    n33701, n33702, n33703, n33704, n33705, n33706,
    n33707, n33708, n33709, n33710, n33711, n33712,
    n33713, n33714, n33715, n33716, n33717, n33718,
    n33719, n33720, n33721, n33722, n33723, n33724,
    n33725, n33726, n33727, n33728, n33729, n33730,
    n33731, n33732, n33733, n33734, n33735, n33736,
    n33737, n33738, n33739, n33740, n33741, n33742,
    n33743, n33744, n33745, n33746, n33747, n33748,
    n33749, n33750, n33751, n33752, n33753, n33754,
    n33755, n33756, n33757, n33758, n33759, n33760,
    n33761, n33762, n33763, n33764, n33765, n33766,
    n33767, n33768, n33769, n33770, n33771, n33772,
    n33773, n33774, n33775, n33776, n33777, n33778,
    n33779, n33780, n33781, n33782, n33783, n33784,
    n33785, n33786, n33787, n33788, n33789, n33790,
    n33791, n33792, n33793, n33794, n33795, n33796,
    n33797, n33798, n33799, n33800, n33801, n33802,
    n33803, n33804, n33805, n33806, n33807, n33808,
    n33809, n33810, n33811, n33812, n33813, n33814,
    n33815, n33816, n33817, n33818, n33819, n33820,
    n33821, n33822, n33823, n33824, n33825, n33826,
    n33827, n33828, n33829, n33830, n33831, n33832,
    n33833, n33834, n33835, n33836, n33837, n33838,
    n33839, n33840, n33841, n33842, n33843, n33844,
    n33845, n33846, n33847, n33848, n33849, n33850,
    n33851, n33852, n33853, n33854, n33855, n33856,
    n33857, n33858, n33859, n33860, n33861, n33862,
    n33863, n33864, n33865, n33866, n33867, n33868,
    n33869, n33870, n33871, n33872, n33873, n33874,
    n33875, n33876, n33877, n33878, n33879, n33880,
    n33881, n33882, n33883, n33884, n33885, n33886,
    n33887, n33888, n33889, n33890, n33891, n33892,
    n33894, n33895, n33896, n33897, n33898, n33899,
    n33900, n33901, n33902, n33903, n33904, n33905,
    n33906, n33907, n33908, n33909, n33910, n33911,
    n33912, n33913, n33914, n33915, n33916, n33917,
    n33918, n33919, n33920, n33921, n33922, n33923,
    n33924, n33925, n33926, n33927, n33928, n33929,
    n33930, n33931, n33932, n33933, n33934, n33935,
    n33936, n33937, n33938, n33939, n33940, n33941,
    n33942, n33943, n33944, n33945, n33946, n33947,
    n33948, n33949, n33950, n33951, n33952, n33953,
    n33954, n33955, n33956, n33957, n33958, n33959,
    n33960, n33961, n33962, n33963, n33964, n33965,
    n33966, n33967, n33968, n33969, n33970, n33971,
    n33972, n33973, n33974, n33975, n33976, n33977,
    n33978, n33979, n33980, n33981, n33982, n33983,
    n33984, n33985, n33986, n33987, n33988, n33989,
    n33990, n33991, n33992, n33993, n33994, n33995,
    n33996, n33997, n33998, n33999, n34000, n34001,
    n34002, n34003, n34004, n34005, n34006, n34007,
    n34008, n34009, n34010, n34011, n34012, n34013,
    n34014, n34015, n34016, n34017, n34018, n34019,
    n34020, n34021, n34022, n34023, n34024, n34025,
    n34026, n34027, n34028, n34029, n34030, n34031,
    n34032, n34033, n34034, n34035, n34036, n34037,
    n34038, n34039, n34040, n34041, n34042, n34043,
    n34044, n34045, n34046, n34047, n34048, n34049,
    n34050, n34051, n34052, n34053, n34054, n34055,
    n34056, n34057, n34058, n34059, n34060, n34061,
    n34062, n34063, n34064, n34065, n34066, n34067,
    n34068, n34069, n34070, n34071, n34072, n34073,
    n34074, n34075, n34076, n34077, n34078, n34079,
    n34080, n34081, n34082, n34083, n34084, n34085,
    n34086, n34087, n34088, n34089, n34090, n34091,
    n34092, n34093, n34094, n34095, n34096, n34097,
    n34098, n34099, n34100, n34101, n34102, n34103,
    n34104, n34105, n34106, n34107, n34108, n34109,
    n34110, n34111, n34112, n34113, n34114, n34115,
    n34116, n34117, n34118, n34119, n34120, n34121,
    n34122, n34123, n34124, n34125, n34126, n34127,
    n34128, n34129, n34130, n34131, n34132, n34133,
    n34134, n34135, n34136, n34137, n34138, n34139,
    n34140, n34141, n34142, n34143, n34145, n34146,
    n34147, n34148, n34149, n34150, n34151, n34152,
    n34153, n34154, n34155, n34156, n34157, n34158,
    n34159, n34160, n34161, n34162, n34163, n34164,
    n34165, n34166, n34167, n34168, n34169, n34170,
    n34171, n34172, n34173, n34174, n34175, n34176,
    n34177, n34178, n34179, n34180, n34181, n34182,
    n34183, n34184, n34185, n34186, n34187, n34188,
    n34189, n34190, n34191, n34192, n34193, n34194,
    n34195, n34196, n34197, n34198, n34199, n34200,
    n34201, n34202, n34203, n34204, n34205, n34206,
    n34207, n34208, n34209, n34210, n34211, n34212,
    n34213, n34214, n34215, n34216, n34217, n34218,
    n34219, n34220, n34221, n34222, n34223, n34224,
    n34225, n34226, n34227, n34228, n34229, n34230,
    n34231, n34232, n34233, n34234, n34235, n34236,
    n34237, n34238, n34239, n34240, n34241, n34242,
    n34243, n34244, n34245, n34246, n34247, n34248,
    n34249, n34250, n34251, n34252, n34253, n34254,
    n34255, n34256, n34257, n34258, n34259, n34260,
    n34261, n34262, n34263, n34264, n34265, n34266,
    n34267, n34268, n34269, n34270, n34271, n34272,
    n34273, n34274, n34275, n34276, n34277, n34278,
    n34279, n34280, n34281, n34282, n34283, n34284,
    n34285, n34286, n34287, n34288, n34289, n34290,
    n34291, n34292, n34293, n34294, n34295, n34296,
    n34297, n34298, n34299, n34300, n34301, n34302,
    n34303, n34304, n34305, n34306, n34307, n34308,
    n34309, n34310, n34311, n34312, n34313, n34314,
    n34315, n34316, n34317, n34318, n34319, n34320,
    n34321, n34322, n34323, n34324, n34325, n34326,
    n34327, n34328, n34329, n34330, n34331, n34332,
    n34333, n34334, n34335, n34336, n34337, n34338,
    n34339, n34340, n34341, n34342, n34343, n34344,
    n34345, n34346, n34347, n34348, n34349, n34350,
    n34351, n34352, n34353, n34354, n34355, n34356,
    n34357, n34358, n34359, n34360, n34361, n34362,
    n34363, n34364, n34365, n34366, n34367, n34368,
    n34369, n34370, n34371, n34372, n34373, n34374,
    n34375, n34376, n34377, n34378, n34380, n34381,
    n34382, n34383, n34384, n34385, n34386, n34387,
    n34388, n34389, n34390, n34391, n34392, n34393,
    n34394, n34395, n34396, n34397, n34398, n34399,
    n34400, n34401, n34402, n34403, n34404, n34405,
    n34406, n34407, n34408, n34409, n34410, n34411,
    n34412, n34413, n34414, n34415, n34416, n34417,
    n34418, n34419, n34420, n34421, n34422, n34423,
    n34424, n34425, n34426, n34427, n34428, n34429,
    n34430, n34431, n34432, n34433, n34434, n34435,
    n34436, n34437, n34438, n34439, n34440, n34441,
    n34442, n34443, n34444, n34445, n34446, n34447,
    n34448, n34449, n34450, n34451, n34452, n34453,
    n34454, n34455, n34456, n34457, n34458, n34459,
    n34460, n34461, n34462, n34463, n34464, n34465,
    n34466, n34467, n34468, n34469, n34470, n34471,
    n34472, n34473, n34474, n34475, n34476, n34477,
    n34478, n34479, n34480, n34481, n34482, n34483,
    n34484, n34485, n34486, n34487, n34488, n34489,
    n34490, n34491, n34492, n34493, n34494, n34495,
    n34496, n34497, n34498, n34499, n34500, n34501,
    n34502, n34503, n34504, n34505, n34506, n34507,
    n34508, n34509, n34510, n34511, n34512, n34513,
    n34514, n34515, n34516, n34517, n34518, n34519,
    n34520, n34521, n34522, n34523, n34524, n34525,
    n34526, n34527, n34528, n34529, n34530, n34531,
    n34532, n34533, n34534, n34535, n34536, n34537,
    n34538, n34539, n34540, n34541, n34542, n34543,
    n34544, n34545, n34546, n34547, n34548, n34549,
    n34550, n34551, n34552, n34553, n34554, n34555,
    n34556, n34557, n34558, n34559, n34560, n34561,
    n34562, n34563, n34564, n34565, n34566, n34567,
    n34568, n34569, n34570, n34571, n34572, n34573,
    n34574, n34575, n34576, n34577, n34578, n34579,
    n34580, n34581, n34582, n34583, n34584, n34585,
    n34586, n34587, n34588, n34590, n34591, n34592,
    n34593, n34594, n34595, n34596, n34597, n34598,
    n34599, n34600, n34601, n34602, n34603, n34604,
    n34605, n34606, n34607, n34608, n34609, n34610,
    n34611, n34612, n34613, n34614, n34615, n34616,
    n34617, n34618, n34619, n34620, n34621, n34622,
    n34623, n34624, n34625, n34626, n34627, n34628,
    n34629, n34630, n34631, n34632, n34633, n34634,
    n34635, n34636, n34637, n34638, n34639, n34640,
    n34641, n34642, n34643, n34644, n34645, n34646,
    n34647, n34648, n34649, n34650, n34651, n34652,
    n34653, n34654, n34655, n34656, n34657, n34658,
    n34659, n34660, n34661, n34662, n34663, n34664,
    n34665, n34666, n34667, n34668, n34669, n34670,
    n34671, n34672, n34673, n34674, n34675, n34676,
    n34677, n34678, n34679, n34680, n34681, n34682,
    n34683, n34684, n34685, n34686, n34687, n34688,
    n34689, n34690, n34691, n34692, n34693, n34694,
    n34695, n34696, n34697, n34698, n34699, n34700,
    n34701, n34702, n34703, n34704, n34705, n34706,
    n34707, n34708, n34709, n34710, n34711, n34712,
    n34713, n34714, n34715, n34716, n34717, n34718,
    n34719, n34720, n34721, n34722, n34723, n34724,
    n34725, n34726, n34727, n34728, n34729, n34730,
    n34731, n34732, n34733, n34734, n34735, n34736,
    n34737, n34738, n34739, n34740, n34741, n34742,
    n34743, n34744, n34745, n34746, n34747, n34748,
    n34749, n34750, n34751, n34752, n34753, n34754,
    n34755, n34756, n34757, n34758, n34759, n34760,
    n34761, n34762, n34763, n34764, n34765, n34766,
    n34767, n34768, n34769, n34770, n34771, n34772,
    n34773, n34774, n34775, n34776, n34777, n34778,
    n34779, n34780, n34781, n34782, n34783, n34784,
    n34785, n34786, n34787, n34788, n34789, n34790,
    n34791, n34792, n34793, n34794, n34795, n34796,
    n34797, n34798, n34799, n34800, n34801, n34802,
    n34803, n34804, n34805, n34806, n34807, n34808,
    n34809, n34810, n34811, n34812, n34813, n34814,
    n34816, n34817, n34818, n34819, n34820, n34821,
    n34822, n34823, n34824, n34825, n34826, n34827,
    n34828, n34829, n34830, n34831, n34832, n34833,
    n34834, n34835, n34836, n34837, n34838, n34839,
    n34840, n34841, n34842, n34843, n34844, n34845,
    n34846, n34847, n34848, n34849, n34850, n34851,
    n34852, n34853, n34854, n34855, n34856, n34857,
    n34858, n34859, n34860, n34861, n34862, n34863,
    n34864, n34865, n34866, n34867, n34868, n34869,
    n34870, n34871, n34872, n34873, n34874, n34875,
    n34876, n34877, n34878, n34879, n34880, n34881,
    n34882, n34883, n34884, n34885, n34886, n34887,
    n34888, n34889, n34890, n34891, n34892, n34893,
    n34894, n34895, n34896, n34897, n34898, n34899,
    n34900, n34901, n34902, n34903, n34904, n34905,
    n34906, n34907, n34908, n34909, n34910, n34911,
    n34912, n34913, n34914, n34915, n34916, n34917,
    n34918, n34919, n34920, n34921, n34922, n34923,
    n34924, n34925, n34926, n34927, n34928, n34929,
    n34930, n34931, n34932, n34933, n34934, n34935,
    n34936, n34937, n34938, n34939, n34940, n34941,
    n34942, n34943, n34944, n34945, n34946, n34947,
    n34948, n34949, n34950, n34951, n34952, n34953,
    n34954, n34955, n34956, n34957, n34958, n34959,
    n34960, n34961, n34962, n34963, n34964, n34965,
    n34966, n34967, n34968, n34969, n34970, n34971,
    n34972, n34973, n34974, n34975, n34976, n34977,
    n34978, n34979, n34980, n34981, n34982, n34983,
    n34984, n34985, n34986, n34987, n34988, n34989,
    n34990, n34991, n34992, n34993, n34994, n34995,
    n34996, n34997, n34998, n34999, n35000, n35001,
    n35002, n35003, n35004, n35005, n35006, n35007,
    n35008, n35009, n35010, n35011, n35012, n35013,
    n35014, n35015, n35016, n35017, n35018, n35019,
    n35020, n35021, n35022, n35023, n35024, n35026,
    n35027, n35028, n35029, n35030, n35031, n35032,
    n35033, n35034, n35035, n35036, n35037, n35038,
    n35039, n35040, n35041, n35042, n35043, n35044,
    n35045, n35046, n35047, n35048, n35049, n35050,
    n35051, n35052, n35053, n35054, n35055, n35056,
    n35057, n35058, n35059, n35060, n35061, n35062,
    n35063, n35064, n35065, n35066, n35067, n35068,
    n35069, n35070, n35071, n35072, n35073, n35074,
    n35075, n35076, n35077, n35078, n35079, n35080,
    n35081, n35082, n35083, n35084, n35085, n35086,
    n35087, n35088, n35089, n35090, n35091, n35092,
    n35093, n35094, n35095, n35096, n35097, n35098,
    n35099, n35100, n35101, n35102, n35103, n35104,
    n35105, n35106, n35107, n35108, n35109, n35110,
    n35111, n35112, n35113, n35114, n35115, n35116,
    n35117, n35118, n35119, n35120, n35121, n35122,
    n35123, n35124, n35125, n35126, n35127, n35128,
    n35129, n35130, n35131, n35132, n35133, n35134,
    n35135, n35136, n35137, n35138, n35139, n35140,
    n35141, n35142, n35143, n35144, n35145, n35146,
    n35147, n35148, n35149, n35150, n35151, n35152,
    n35153, n35154, n35155, n35156, n35157, n35158,
    n35159, n35160, n35161, n35162, n35163, n35164,
    n35165, n35166, n35167, n35168, n35169, n35170,
    n35171, n35172, n35173, n35174, n35175, n35176,
    n35177, n35178, n35179, n35180, n35181, n35182,
    n35183, n35184, n35185, n35186, n35187, n35188,
    n35189, n35190, n35191, n35192, n35193, n35194,
    n35195, n35196, n35197, n35198, n35199, n35200,
    n35201, n35202, n35203, n35204, n35205, n35206,
    n35207, n35208, n35209, n35210, n35211, n35213,
    n35214, n35215, n35216, n35217, n35218, n35219,
    n35220, n35221, n35222, n35223, n35224, n35225,
    n35226, n35227, n35228, n35229, n35230, n35231,
    n35232, n35233, n35234, n35235, n35236, n35237,
    n35238, n35239, n35240, n35241, n35242, n35243,
    n35244, n35245, n35246, n35247, n35248, n35249,
    n35250, n35251, n35252, n35253, n35254, n35255,
    n35256, n35257, n35258, n35259, n35260, n35261,
    n35262, n35263, n35264, n35265, n35266, n35267,
    n35268, n35269, n35270, n35271, n35272, n35273,
    n35274, n35275, n35276, n35277, n35278, n35279,
    n35280, n35281, n35282, n35283, n35284, n35285,
    n35286, n35287, n35288, n35289, n35290, n35291,
    n35292, n35293, n35294, n35295, n35296, n35297,
    n35298, n35299, n35300, n35301, n35302, n35303,
    n35304, n35305, n35306, n35307, n35308, n35309,
    n35310, n35311, n35312, n35313, n35314, n35315,
    n35316, n35317, n35318, n35319, n35320, n35321,
    n35322, n35323, n35324, n35325, n35326, n35327,
    n35328, n35329, n35330, n35331, n35332, n35333,
    n35334, n35335, n35336, n35337, n35338, n35339,
    n35340, n35341, n35342, n35343, n35344, n35345,
    n35346, n35347, n35348, n35349, n35350, n35351,
    n35352, n35353, n35354, n35355, n35356, n35357,
    n35358, n35359, n35360, n35361, n35362, n35363,
    n35364, n35365, n35366, n35367, n35368, n35369,
    n35370, n35371, n35372, n35373, n35374, n35375,
    n35376, n35377, n35378, n35379, n35380, n35381,
    n35382, n35383, n35384, n35385, n35386, n35387,
    n35388, n35389, n35390, n35391, n35392, n35393,
    n35394, n35395, n35396, n35397, n35398, n35399,
    n35400, n35401, n35402, n35403, n35404, n35405,
    n35406, n35407, n35408, n35409, n35410, n35411,
    n35412, n35413, n35414, n35416, n35417, n35418,
    n35419, n35420, n35421, n35422, n35423, n35424,
    n35425, n35426, n35427, n35428, n35429, n35430,
    n35431, n35432, n35433, n35434, n35435, n35436,
    n35437, n35438, n35439, n35440, n35441, n35442,
    n35443, n35444, n35445, n35446, n35447, n35448,
    n35449, n35450, n35451, n35452, n35453, n35454,
    n35455, n35456, n35457, n35458, n35459, n35460,
    n35461, n35462, n35463, n35464, n35465, n35466,
    n35467, n35468, n35469, n35470, n35471, n35472,
    n35473, n35474, n35475, n35476, n35477, n35478,
    n35479, n35480, n35481, n35482, n35483, n35484,
    n35485, n35486, n35487, n35488, n35489, n35490,
    n35491, n35492, n35493, n35494, n35495, n35496,
    n35497, n35498, n35499, n35500, n35501, n35502,
    n35503, n35504, n35505, n35506, n35507, n35508,
    n35509, n35510, n35511, n35512, n35513, n35514,
    n35515, n35516, n35517, n35518, n35519, n35520,
    n35521, n35522, n35523, n35524, n35525, n35526,
    n35527, n35528, n35529, n35530, n35531, n35532,
    n35533, n35534, n35535, n35536, n35537, n35538,
    n35539, n35540, n35541, n35542, n35543, n35544,
    n35545, n35546, n35547, n35548, n35549, n35550,
    n35551, n35552, n35553, n35554, n35555, n35556,
    n35557, n35558, n35559, n35560, n35561, n35562,
    n35563, n35564, n35565, n35566, n35567, n35568,
    n35569, n35570, n35571, n35572, n35573, n35574,
    n35575, n35576, n35577, n35578, n35579, n35580,
    n35581, n35582, n35583, n35584, n35585, n35587,
    n35588, n35589, n35590, n35591, n35592, n35593,
    n35594, n35595, n35596, n35597, n35598, n35599,
    n35600, n35601, n35602, n35603, n35604, n35605,
    n35606, n35607, n35608, n35609, n35610, n35611,
    n35612, n35613, n35614, n35615, n35616, n35617,
    n35618, n35619, n35620, n35621, n35622, n35623,
    n35624, n35625, n35626, n35627, n35628, n35629,
    n35630, n35631, n35632, n35633, n35634, n35635,
    n35636, n35637, n35638, n35639, n35640, n35641,
    n35642, n35643, n35644, n35645, n35646, n35647,
    n35648, n35649, n35650, n35651, n35652, n35653,
    n35654, n35655, n35656, n35657, n35658, n35659,
    n35660, n35661, n35662, n35663, n35664, n35665,
    n35666, n35667, n35668, n35669, n35670, n35671,
    n35672, n35673, n35674, n35675, n35676, n35677,
    n35678, n35679, n35680, n35681, n35682, n35683,
    n35684, n35685, n35686, n35687, n35688, n35689,
    n35690, n35691, n35692, n35693, n35694, n35695,
    n35696, n35697, n35698, n35699, n35700, n35701,
    n35702, n35703, n35704, n35705, n35706, n35707,
    n35708, n35709, n35710, n35711, n35712, n35713,
    n35714, n35715, n35716, n35717, n35718, n35719,
    n35720, n35721, n35722, n35723, n35724, n35725,
    n35726, n35727, n35728, n35729, n35730, n35731,
    n35732, n35733, n35734, n35735, n35736, n35737,
    n35738, n35739, n35740, n35741, n35742, n35743,
    n35744, n35745, n35747, n35748, n35749, n35750,
    n35751, n35752, n35753, n35754, n35755, n35756,
    n35757, n35758, n35759, n35760, n35761, n35762,
    n35763, n35764, n35765, n35766, n35767, n35768,
    n35769, n35770, n35771, n35772, n35773, n35774,
    n35775, n35776, n35777, n35778, n35779, n35780,
    n35781, n35782, n35783, n35784, n35785, n35786,
    n35787, n35788, n35789, n35790, n35791, n35792,
    n35793, n35794, n35795, n35796, n35797, n35798,
    n35799, n35800, n35801, n35802, n35803, n35804,
    n35805, n35806, n35807, n35808, n35809, n35810,
    n35811, n35812, n35813, n35814, n35815, n35816,
    n35817, n35818, n35819, n35820, n35821, n35822,
    n35823, n35824, n35825, n35826, n35827, n35828,
    n35829, n35830, n35831, n35832, n35833, n35834,
    n35835, n35836, n35837, n35838, n35839, n35840,
    n35841, n35842, n35843, n35844, n35845, n35846,
    n35847, n35848, n35849, n35850, n35851, n35852,
    n35853, n35854, n35855, n35856, n35857, n35858,
    n35859, n35860, n35861, n35862, n35863, n35864,
    n35865, n35866, n35867, n35868, n35869, n35870,
    n35871, n35872, n35873, n35874, n35875, n35876,
    n35877, n35878, n35879, n35880, n35881, n35882,
    n35883, n35884, n35885, n35886, n35887, n35888,
    n35889, n35890, n35891, n35892, n35893, n35894,
    n35895, n35896, n35897, n35898, n35899, n35900,
    n35901, n35902, n35903, n35904, n35905, n35906,
    n35907, n35908, n35909, n35910, n35911, n35912,
    n35913, n35914, n35915, n35916, n35918, n35919,
    n35920, n35921, n35922, n35923, n35924, n35925,
    n35926, n35927, n35928, n35929, n35930, n35931,
    n35932, n35933, n35934, n35935, n35936, n35937,
    n35938, n35939, n35940, n35941, n35942, n35943,
    n35944, n35945, n35946, n35947, n35948, n35949,
    n35950, n35951, n35952, n35953, n35954, n35955,
    n35956, n35957, n35958, n35959, n35960, n35961,
    n35962, n35963, n35964, n35965, n35966, n35967,
    n35968, n35969, n35970, n35971, n35972, n35973,
    n35974, n35975, n35976, n35977, n35978, n35979,
    n35980, n35981, n35982, n35983, n35984, n35985,
    n35986, n35987, n35988, n35989, n35990, n35991,
    n35992, n35993, n35994, n35995, n35996, n35997,
    n35998, n35999, n36000, n36001, n36002, n36003,
    n36004, n36005, n36006, n36007, n36008, n36009,
    n36010, n36011, n36012, n36013, n36014, n36015,
    n36016, n36017, n36018, n36019, n36020, n36021,
    n36022, n36023, n36024, n36025, n36026, n36027,
    n36028, n36029, n36030, n36031, n36032, n36033,
    n36034, n36035, n36036, n36037, n36038, n36039,
    n36040, n36041, n36042, n36043, n36044, n36045,
    n36046, n36047, n36048, n36049, n36050, n36051,
    n36052, n36053, n36054, n36055, n36056, n36057,
    n36058, n36059, n36060, n36061, n36062, n36063,
    n36064, n36065, n36066, n36068, n36069, n36070,
    n36071, n36072, n36073, n36074, n36075, n36076,
    n36077, n36078, n36079, n36080, n36081, n36082,
    n36083, n36084, n36085, n36086, n36087, n36088,
    n36089, n36090, n36091, n36092, n36093, n36094,
    n36095, n36096, n36097, n36098, n36099, n36100,
    n36101, n36102, n36103, n36104, n36105, n36106,
    n36107, n36108, n36109, n36110, n36111, n36112,
    n36113, n36114, n36115, n36116, n36117, n36118,
    n36119, n36120, n36121, n36122, n36123, n36124,
    n36125, n36126, n36127, n36128, n36129, n36130,
    n36131, n36132, n36133, n36134, n36135, n36136,
    n36137, n36138, n36139, n36140, n36141, n36142,
    n36143, n36144, n36145, n36146, n36147, n36148,
    n36149, n36150, n36151, n36152, n36153, n36154,
    n36155, n36156, n36157, n36158, n36159, n36160,
    n36161, n36162, n36163, n36164, n36165, n36166,
    n36167, n36168, n36169, n36170, n36171, n36172,
    n36173, n36174, n36175, n36176, n36177, n36178,
    n36179, n36180, n36181, n36182, n36183, n36184,
    n36185, n36186, n36187, n36188, n36189, n36190,
    n36191, n36192, n36193, n36194, n36195, n36196,
    n36198, n36199, n36200, n36201, n36202, n36203,
    n36204, n36205, n36206, n36207, n36208, n36209,
    n36210, n36211, n36212, n36213, n36214, n36215,
    n36216, n36217, n36218, n36219, n36220, n36221,
    n36222, n36223, n36224, n36225, n36226, n36227,
    n36228, n36229, n36230, n36231, n36232, n36233,
    n36234, n36235, n36236, n36237, n36238, n36239,
    n36240, n36241, n36242, n36243, n36244, n36245,
    n36246, n36247, n36248, n36249, n36250, n36251,
    n36252, n36253, n36254, n36255, n36256, n36257,
    n36258, n36259, n36260, n36261, n36262, n36263,
    n36264, n36265, n36266, n36267, n36268, n36269,
    n36270, n36271, n36272, n36273, n36274, n36275,
    n36276, n36277, n36278, n36279, n36280, n36281,
    n36282, n36283, n36284, n36285, n36286, n36287,
    n36288, n36289, n36290, n36291, n36292, n36293,
    n36294, n36295, n36296, n36297, n36298, n36299,
    n36300, n36301, n36302, n36303, n36304, n36305,
    n36306, n36307, n36308, n36309, n36310, n36311,
    n36312, n36313, n36314, n36315, n36316, n36317,
    n36318, n36319, n36320, n36321, n36322, n36323,
    n36324, n36325, n36326, n36327, n36328, n36329,
    n36330, n36331, n36332, n36334, n36335, n36336,
    n36337, n36338, n36339, n36340, n36341, n36342,
    n36343, n36344, n36345, n36346, n36347, n36348,
    n36349, n36350, n36351, n36352, n36353, n36354,
    n36355, n36356, n36357, n36358, n36359, n36360,
    n36361, n36362, n36363, n36364, n36365, n36366,
    n36367, n36368, n36369, n36370, n36371, n36372,
    n36373, n36374, n36375, n36376, n36377, n36378,
    n36379, n36380, n36381, n36382, n36383, n36384,
    n36385, n36386, n36387, n36388, n36389, n36390,
    n36391, n36392, n36393, n36394, n36395, n36396,
    n36397, n36398, n36399, n36400, n36401, n36402,
    n36403, n36404, n36405, n36406, n36407, n36408,
    n36409, n36410, n36411, n36412, n36413, n36414,
    n36415, n36416, n36417, n36418, n36419, n36420,
    n36421, n36422, n36423, n36424, n36425, n36426,
    n36427, n36428, n36429, n36430, n36431, n36432,
    n36433, n36434, n36435, n36436, n36437, n36438,
    n36439, n36440, n36441, n36442, n36443, n36444,
    n36445, n36446, n36447, n36448, n36449, n36450,
    n36451, n36452, n36453, n36454, n36455, n36456,
    n36457, n36458, n36459, n36460, n36461, n36462,
    n36463, n36464, n36465, n36466, n36468, n36469,
    n36470, n36471, n36472, n36473, n36474, n36475,
    n36476, n36477, n36478, n36479, n36480, n36481,
    n36482, n36483, n36484, n36485, n36486, n36487,
    n36488, n36489, n36490, n36491, n36492, n36493,
    n36494, n36495, n36496, n36497, n36498, n36499,
    n36500, n36501, n36502, n36503, n36504, n36505,
    n36506, n36507, n36508, n36509, n36510, n36511,
    n36512, n36513, n36514, n36515, n36516, n36517,
    n36518, n36519, n36520, n36521, n36522, n36523,
    n36524, n36525, n36526, n36527, n36528, n36529,
    n36530, n36531, n36532, n36533, n36534, n36535,
    n36536, n36537, n36538, n36539, n36540, n36541,
    n36542, n36543, n36544, n36545, n36546, n36547,
    n36548, n36549, n36550, n36551, n36552, n36553,
    n36554, n36555, n36556, n36557, n36558, n36559,
    n36560, n36561, n36562, n36563, n36564, n36565,
    n36566, n36567, n36568, n36569, n36571, n36572,
    n36573, n36574, n36575, n36576, n36577, n36578,
    n36579, n36580, n36581, n36582, n36583, n36584,
    n36585, n36586, n36587, n36588, n36589, n36590,
    n36591, n36592, n36593, n36594, n36595, n36596,
    n36597, n36598, n36599, n36600, n36601, n36602,
    n36603, n36604, n36605, n36606, n36607, n36608,
    n36609, n36610, n36611, n36612, n36613, n36614,
    n36615, n36616, n36617, n36618, n36619, n36620,
    n36621, n36622, n36623, n36624, n36625, n36626,
    n36627, n36628, n36629, n36630, n36631, n36632,
    n36633, n36634, n36635, n36636, n36637, n36638,
    n36639, n36640, n36641, n36642, n36643, n36644,
    n36645, n36646, n36647, n36648, n36649, n36650,
    n36651, n36652, n36653, n36654, n36655, n36656,
    n36657, n36658, n36659, n36660, n36661, n36662,
    n36663, n36664, n36665, n36666, n36667, n36668,
    n36669, n36670, n36671, n36672, n36673, n36674,
    n36675, n36676, n36677, n36678, n36679, n36681,
    n36682, n36683, n36684, n36685, n36686, n36687,
    n36688, n36689, n36690, n36691, n36692, n36693,
    n36694, n36695, n36696, n36697, n36698, n36699,
    n36700, n36701, n36702, n36703, n36704, n36705,
    n36706, n36707, n36708, n36709, n36710, n36711,
    n36712, n36713, n36714, n36715, n36716, n36717,
    n36718, n36719, n36720, n36721, n36722, n36723,
    n36724, n36725, n36726, n36727, n36728, n36729,
    n36730, n36731, n36732, n36733, n36734, n36735,
    n36736, n36737, n36738, n36739, n36740, n36741,
    n36742, n36743, n36744, n36745, n36746, n36747,
    n36748, n36749, n36750, n36751, n36752, n36753,
    n36754, n36755, n36756, n36757, n36758, n36759,
    n36760, n36761, n36762, n36763, n36764, n36765,
    n36766, n36767, n36768, n36769, n36770, n36771,
    n36772, n36773, n36774, n36775, n36776, n36777,
    n36778, n36779, n36780, n36781, n36782, n36783,
    n36784, n36785, n36786, n36787, n36788, n36789,
    n36790, n36791, n36793, n36794, n36795, n36796,
    n36797, n36798, n36799, n36800, n36801, n36802,
    n36803, n36804, n36805, n36806, n36807, n36808,
    n36809, n36810, n36811, n36812, n36813, n36814,
    n36815, n36816, n36817, n36818, n36819, n36820,
    n36821, n36822, n36823, n36824, n36825, n36826,
    n36827, n36828, n36829, n36830, n36831, n36832,
    n36833, n36834, n36835, n36836, n36837, n36838,
    n36839, n36840, n36841, n36842, n36843, n36844,
    n36845, n36846, n36847, n36848, n36849, n36850,
    n36851, n36852, n36853, n36854, n36855, n36856,
    n36857, n36858, n36859, n36860, n36861, n36862,
    n36863, n36864, n36865, n36866, n36867, n36868,
    n36869, n36870, n36871, n36872, n36873, n36874,
    n36875, n36877, n36878, n36879, n36880, n36881,
    n36882, n36883, n36884, n36885, n36886, n36887,
    n36888, n36889, n36890, n36891, n36892, n36893,
    n36894, n36895, n36896, n36897, n36898, n36899,
    n36900, n36901, n36902, n36903, n36904, n36905,
    n36906, n36907, n36908, n36909, n36910, n36911,
    n36912, n36913, n36914, n36915, n36916, n36917,
    n36918, n36919, n36920, n36921, n36922, n36923,
    n36924, n36925, n36926, n36927, n36928, n36929,
    n36930, n36931, n36932, n36933, n36934, n36935,
    n36936, n36937, n36938, n36939, n36940, n36941,
    n36942, n36943, n36944, n36945, n36946, n36947,
    n36948, n36949, n36950, n36951, n36952, n36953,
    n36954, n36955, n36956, n36957, n36958, n36959,
    n36960, n36961, n36962, n36963, n36964, n36966,
    n36967, n36968, n36969, n36970, n36971, n36972,
    n36973, n36974, n36975, n36976, n36977, n36978,
    n36979, n36980, n36981, n36982, n36983, n36984,
    n36985, n36986, n36987, n36988, n36989, n36990,
    n36991, n36992, n36993, n36994, n36995, n36996,
    n36997, n36998, n36999, n37000, n37001, n37002,
    n37003, n37004, n37005, n37006, n37007, n37008,
    n37009, n37010, n37011, n37012, n37013, n37014,
    n37015, n37016, n37017, n37018, n37019, n37020,
    n37021, n37022, n37023, n37024, n37025, n37026,
    n37027, n37028, n37029, n37030, n37031, n37032,
    n37033, n37034, n37035, n37036, n37037, n37038,
    n37039, n37040, n37041, n37042, n37043, n37044,
    n37045, n37046, n37047, n37048, n37049, n37051,
    n37052, n37053, n37054, n37055, n37056, n37057,
    n37058, n37059, n37060, n37061, n37062, n37063,
    n37064, n37065, n37066, n37067, n37068, n37069,
    n37070, n37071, n37072, n37073, n37074, n37075,
    n37076, n37077, n37078, n37079, n37080, n37081,
    n37082, n37083, n37084, n37085, n37086, n37087,
    n37088, n37089, n37090, n37091, n37092, n37093,
    n37094, n37095, n37096, n37097, n37098, n37099,
    n37100, n37101, n37102, n37103, n37105, n37106,
    n37107, n37108, n37109, n37110, n37111, n37112,
    n37113, n37114, n37115, n37116, n37117, n37118,
    n37119, n37120, n37121, n37122, n37123, n37124,
    n37125, n37126, n37127, n37128, n37129, n37130,
    n37131, n37132, n37133, n37134, n37135, n37136,
    n37137, n37138, n37139, n37140, n37141, n37142,
    n37143, n37144, n37145, n37146, n37147, n37148,
    n37149, n37150, n37151, n37152, n37153, n37154,
    n37155, n37156, n37157, n37158, n37159, n37160,
    n37161, n37162, n37163, n37164, n37165, n37166,
    n37167, n37168, n37169, n37170, n37171, n37172,
    n37173, n37175, n37176, n37177, n37178, n37179,
    n37180, n37181, n37182, n37183, n37184, n37185,
    n37186, n37187, n37188, n37189, n37190, n37191,
    n37192, n37193, n37194, n37195, n37196, n37197,
    n37198, n37199, n37200, n37201, n37202, n37203,
    n37204, n37205, n37206, n37207, n37208, n37209,
    n37210, n37211, n37212, n37213, n37214, n37215,
    n37216, n37217, n37218, n37219, n37220, n37221,
    n37222, n37223, n37224, n37226, n37227, n37228,
    n37229, n37230, n37231, n37232, n37233, n37234,
    n37235, n37236, n37237, n37238, n37239, n37240,
    n37241, n37242, n37243, n37244, n37245, n37246,
    n37247, n37248, n37249, n37250, n37251, n37252,
    n37253, n37254, n37255, n37256, n37257, n37258,
    n37260, n37261, n37262, n37263, n37264, n37265,
    n37266, n37267, n37268, n37269, n37270, n37271,
    n37272, n37273, n37274, n37275, n37276, n37277,
    n37278, n37279, n37280, n37281, n37282, n37283,
    n37284, n37285, n37286, n37287, n37288, n37289,
    n37290, n37292, n37293, n37294, n37295, n37296,
    n37297, n37298, n37299, n37300, n37301, n37302,
    n37303, n37304, n37305, n37306, n37307, n37308,
    n37309, n37310, n37311, n37312, n37313, n37315,
    n37316, n37317, n37318, n37319, n37320, n37321,
    n37322, n37323, n37324, n37325, n37326, n37327,
    n37328, n37329, n37330, n37331, n37332, n37333,
    n37334, n37336, n37338, n37340, n37341, n37342,
    n37344, n37346, n37348, n37350, n37352, n37354,
    n37356, n37358, n37360, n37362, n37364, n37366,
    n37368, n37370, n37372, n37374, n37376, n37378,
    n37380, n37382, n37384, n37386, n37388, n37390,
    n37392, n37394, n37396, n37398, n37400, n37402,
    n37404, n37406, n37408, n37410, n37412, n37414,
    n37416, n37418, n37420, n37422, n37424, n37426,
    n37428, n37430, n37431, n37432, n37434, n37436,
    n37438, n37440, n37442, n37444, n37446, n37448,
    n37450, n37452, n37454, n37456, n37458, n37459,
    n37460, n37461, n37462, n37463, n37464, n37465,
    n37466, n37467, n37468, n37469, n37470, n37471,
    n37472, n37473, n37474, n37475, n37476, n37477,
    n37478, n37479, n37480, n37481, n37482, n37483,
    n37484, n37485, n37486, n37487, n37488, n37489,
    n37490, n37491, n37492, n37493, n37494, n37495,
    n37496, n37497, n37498, n37499, n37500, n37501,
    n37502, n37503, n37504, n37505, n37506, n37507,
    n37508, n37509, n37510, n37511, n37512, n37513,
    n37514, n37515, n37516, n37517, n37518, n37519,
    n37520, n37521, n37522, n37523, n37524, n37525,
    n37526, n37527, n37528, n37529, n37530, n37531,
    n37532, n37533, n37534, n37535, n37536, n37537,
    n37538, n37539, n37540, n37541, n37542, n37543,
    n37544, n37545, n37546, n37547, n37548, n37549,
    n37550, n37551, n37552, n37553, n37554, n37555,
    n37556, n37557, n37558, n37559, n37560, n37561,
    n37562, n37563, n37564, n37565, n37566, n37567,
    n37568, n37569, n37570, n37571, n37572, n37573,
    n37574, n37575, n37576, n37577, n37578, n37579,
    n37580, n37581, n37582, n37583, n37584, n37585,
    n37586, n37587, n37588, n37589, n37590, n37591,
    n37592, n37593, n37594, n37595, n37596, n37597,
    n37598, n37599, n37600, n37601, n37602, n37603,
    n37604, n37605, n37606, n37607, n37608, n37609,
    n37610, n37611, n37612, n37613, n37614, n37615,
    n37616, n37617, n37618, n37619, n37620, n37621,
    n37622, n37623, n37624, n37625, n37626, n37627,
    n37628, n37629, n37630, n37631, n37632, n37633,
    n37634, n37635, n37636, n37637, n37638, n37639,
    n37640, n37641, n37642, n37643, n37644, n37645,
    n37646, n37647, n37648, n37649, n37650, n37651,
    n37652, n37653, n37654, n37655, n37656, n37657,
    n37658, n37659, n37660, n37661, n37662, n37663,
    n37664, n37665, n37666, n37667, n37668, n37669,
    n37670, n37671, n37672, n37673, n37674, n37675,
    n37676, n37677, n37678, n37679, n37680, n37681,
    n37682, n37683, n37684, n37685, n37686, n37687,
    n37688, n37689, n37690, n37691, n37692, n37693,
    n37694, n37695, n37696, n37697, n37698, n37699,
    n37700, n37701, n37702, n37703, n37704, n37705,
    n37706, n37707, n37708, n37709, n37710, n37711,
    n37712, n37713, n37714, n37715, n37716, n37717,
    n37718, n37719, n37720, n37721, n37722, n37723,
    n37724, n37725, n37726, n37727, n37728, n37729,
    n37730, n37731, n37732, n37733, n37734, n37735,
    n37736, n37737, n37738, n37739, n37740, n37741,
    n37742, n37743, n37744, n37745, n37746, n37747,
    n37748, n37749, n37750, n37751, n37752, n37753,
    n37754, n37755, n37756, n37757, n37758, n37759,
    n37760, n37761, n37762, n37763, n37764, n37765,
    n37766, n37767, n37768, n37769, n37770, n37771,
    n37772, n37773, n37774, n37775, n37776, n37777,
    n37778, n37779, n37780, n37781, n37782, n37783,
    n37784, n37785, n37786, n37787, n37788, n37789,
    n37790, n37791, n37792, n37793, n37794, n37795,
    n37796, n37797, n37798, n37799, n37800, n37801,
    n37802, n37803, n37804, n37805, n37806, n37807,
    n37808, n37809, n37810, n37811, n37812, n37813,
    n37814, n37815, n37816, n37817, n37818, n37819,
    n37820, n37821, n37822, n37823, n37824, n37825,
    n37826, n37827, n37828, n37829, n37830, n37831,
    n37832, n37833, n37834, n37835, n37836, n37837,
    n37838, n37839, n37840, n37841, n37842, n37843,
    n37844, n37845, n37846, n37847, n37848, n37849,
    n37850, n37851, n37852, n37853, n37854, n37855,
    n37856, n37857, n37858, n37859, n37860, n37861,
    n37862, n37863, n37864, n37865, n37866, n37867,
    n37868, n37869, n37870, n37871, n37872, n37873,
    n37874, n37875, n37876, n37877, n37878, n37879,
    n37880, n37881, n37882, n37883, n37884, n37885,
    n37886, n37887, n37888, n37889, n37890, n37891,
    n37892, n37893, n37894, n37895, n37896, n37897,
    n37898, n37899, n37900, n37901, n37902, n37903,
    n37904, n37905, n37906, n37907, n37908, n37909,
    n37910, n37911, n37912, n37913, n37914, n37915,
    n37916, n37917, n37918, n37919, n37920, n37921,
    n37922, n37923, n37924, n37925, n37926, n37927,
    n37928, n37929, n37930, n37931, n37932, n37933,
    n37934, n37935, n37936, n37937, n37938, n37939,
    n37940, n37941, n37942, n37943, n37944, n37945,
    n37946, n37947, n37948, n37949, n37950, n37951,
    n37952, n37953, n37954, n37955, n37956, n37957,
    n37958, n37959, n37960, n37961, n37962, n37963,
    n37964, n37965, n37966, n37967, n37968, n37969,
    n37970, n37971, n37972, n37973, n37974, n37975,
    n37976, n37977, n37978, n37979, n37980, n37981,
    n37982, n37983, n37984, n37985, n37986, n37987,
    n37988, n37989, n37990, n37991, n37992, n37993,
    n37994, n37995, n37996, n37997, n37998, n37999,
    n38000, n38001, n38002, n38003, n38004, n38005,
    n38006, n38007, n38008, n38009, n38010, n38011,
    n38012, n38013, n38014, n38015, n38016, n38017,
    n38018, n38019, n38020, n38021, n38022, n38023,
    n38024, n38025, n38026, n38027, n38028, n38029,
    n38030, n38031, n38032, n38033, n38034, n38035,
    n38036, n38037, n38038, n38039, n38040, n38041,
    n38042, n38043, n38044, n38045, n38046, n38047,
    n38048, n38049, n38050, n38051, n38052, n38053,
    n38054, n38055, n38056, n38057, n38058, n38059,
    n38060, n38061, n38062, n38063, n38064, n38065,
    n38066, n38067, n38068, n38069, n38070, n38071,
    n38072, n38073, n38074, n38075, n38076, n38077,
    n38078, n38079, n38080, n38081, n38082, n38083,
    n38084, n38085, n38086, n38087, n38088, n38089,
    n38090, n38091, n38092, n38093, n38094, n38095,
    n38096, n38097, n38098, n38099, n38100, n38101,
    n38102, n38103, n38104, n38105, n38106, n38107,
    n38108, n38109, n38110, n38111, n38112, n38113,
    n38114, n38115, n38116, n38117, n38118, n38119,
    n38120, n38121, n38122, n38123, n38124, n38125,
    n38126, n38127, n38128, n38129, n38130, n38131,
    n38132, n38133, n38134, n38135, n38136, n38137,
    n38138, n38139, n38140, n38141, n38142, n38143,
    n38144, n38145, n38146, n38147, n38148, n38149,
    n38150, n38151, n38152, n38153, n38154, n38155,
    n38156, n38157, n38158, n38159, n38160, n38161,
    n38162, n38163, n38164, n38165, n38166, n38167,
    n38168, n38169, n38170, n38171, n38172, n38173,
    n38174, n38175, n38176, n38177, n38178, n38179,
    n38180, n38181, n38182, n38183, n38184, n38185,
    n38186, n38187, n38188, n38189, n38190, n38191,
    n38192, n38193, n38194, n38195, n38196, n38197,
    n38198, n38199, n38200, n38201, n38202, n38203,
    n38204, n38205, n38206, n38207, n38208, n38209,
    n38210, n38211, n38212, n38213, n38214, n38215,
    n38216, n38217, n38218, n38219, n38220, n38221,
    n38222, n38223, n38224, n38225, n38226, n38227,
    n38228, n38229, n38230, n38231, n38232, n38233,
    n38234, n38235, n38236, n38237, n38238, n38239,
    n38240, n38241, n38242, n38243, n38244, n38245,
    n38246, n38247, n38248, n38249, n38250, n38251,
    n38252, n38253, n38254, n38255, n38256, n38257,
    n38258, n38259, n38260, n38261, n38262, n38263,
    n38264, n38265, n38266, n38267, n38268, n38269,
    n38270, n38271, n38272, n38273, n38274, n38275,
    n38276, n38277, n38278, n38279, n38280, n38281,
    n38282, n38283, n38284, n38285, n38286, n38287,
    n38288, n38289, n38290, n38291, n38292, n38293,
    n38294, n38295, n38296, n38297, n38298, n38299,
    n38300, n38301, n38302, n38303, n38304, n38305,
    n38306, n38307, n38308, n38309, n38310, n38311,
    n38312, n38313, n38314, n38315, n38316, n38317,
    n38318, n38319, n38320, n38321, n38322, n38323,
    n38324, n38325, n38326, n38327, n38328, n38329,
    n38330, n38331, n38332, n38333, n38334, n38335,
    n38336, n38337, n38338, n38339, n38340, n38341,
    n38342, n38343, n38344, n38345, n38346, n38347,
    n38348, n38349, n38350, n38351, n38352, n38353,
    n38354, n38355, n38356, n38357, n38358, n38359,
    n38360, n38361, n38362, n38363, n38364, n38365,
    n38366, n38367, n38368, n38369, n38370, n38371,
    n38372, n38373, n38374, n38375, n38376, n38377,
    n38378, n38379, n38380, n38381, n38382, n38383,
    n38384, n38385, n38386, n38387, n38388, n38389,
    n38390, n38391, n38392, n38393, n38394, n38395,
    n38396, n38397, n38398, n38399, n38400, n38401,
    n38402, n38403, n38404, n38405, n38406, n38407,
    n38408, n38409, n38410, n38411, n38412, n38413,
    n38414, n38415, n38416, n38417, n38418, n38419,
    n38420, n38421, n38422, n38423, n38424, n38425,
    n38426, n38427, n38428, n38429, n38430, n38431,
    n38432, n38433, n38434, n38435, n38436, n38437,
    n38438, n38439, n38440, n38441, n38442, n38443,
    n38444, n38445, n38446, n38447, n38448, n38449,
    n38450, n38451, n38452, n38453, n38454, n38455,
    n38456, n38457, n38458, n38459, n38460, n38461,
    n38462, n38463, n38464, n38465, n38466, n38467,
    n38468, n38469, n38470, n38471, n38472, n38473,
    n38474, n38475, n38476, n38477, n38478, n38479,
    n38480, n38481, n38482, n38483, n38484, n38485,
    n38486, n38487, n38488, n38489, n38490, n38491,
    n38492, n38493, n38494, n38495, n38496, n38497,
    n38498, n38499, n38500, n38501, n38502, n38503,
    n38504, n38505, n38506, n38507, n38508, n38509,
    n38510, n38511, n38512, n38513, n38514, n38515,
    n38516, n38517, n38518, n38519, n38520, n38521,
    n38522, n38523, n38524, n38525, n38526, n38527,
    n38528, n38529, n38530, n38531, n38532, n38533,
    n38534, n38535, n38536, n38537, n38538, n38539,
    n38540, n38541, n38542, n38543, n38544, n38545,
    n38546, n38547, n38548, n38549, n38550, n38551,
    n38552, n38553, n38554, n38555, n38556, n38557,
    n38558, n38559, n38560, n38561, n38562, n38563,
    n38564, n38565, n38566, n38567, n38568, n38569,
    n38570, n38571, n38572, n38573, n38574, n38575,
    n38576, n38577, n38578, n38579, n38580, n38581,
    n38582, n38583, n38584, n38585, n38586, n38587,
    n38588, n38589, n38590, n38591, n38592, n38593,
    n38594, n38595, n38596, n38597, n38598, n38599,
    n38600, n38601, n38602, n38603, n38604, n38605,
    n38606, n38607, n38608, n38609, n38610, n38611,
    n38612, n38613, n38614, n38615, n38616, n38617,
    n38618, n38619, n38620, n38621, n38622, n38623,
    n38624, n38625, n38626, n38627, n38628, n38629,
    n38630, n38631, n38632, n38633, n38634, n38635,
    n38636, n38637, n38638, n38639, n38640, n38641,
    n38642, n38643, n38644, n38645, n38646, n38647,
    n38648, n38649, n38650, n38651, n38652, n38653,
    n38654, n38655, n38656, n38657, n38658, n38659,
    n38660, n38661, n38662, n38663, n38664, n38665,
    n38666, n38667, n38668, n38669, n38670, n38671,
    n38672, n38673, n38674, n38675, n38676, n38677,
    n38678, n38679, n38680, n38681, n38682, n38683,
    n38684, n38685, n38686, n38687, n38688, n38689,
    n38690, n38691, n38692, n38693, n38694, n38695,
    n38696, n38697, n38698, n38699, n38700, n38701,
    n38702, n38703, n38704, n38705, n38706, n38707,
    n38708, n38709, n38710, n38711, n38712, n38713,
    n38714, n38715, n38716, n38717, n38718, n38719,
    n38720, n38721, n38722, n38723, n38724, n38725,
    n38726, n38727, n38728, n38729, n38730, n38731,
    n38732, n38733, n38734, n38735, n38736, n38737,
    n38738, n38739, n38740, n38741, n38742, n38743,
    n38744, n38745, n38746, n38747, n38748, n38749,
    n38750, n38751, n38752, n38753, n38754, n38755,
    n38756, n38757, n38758, n38759, n38760, n38761,
    n38762, n38763, n38764, n38765, n38766, n38767,
    n38768, n38769, n38770, n38771, n38772, n38773,
    n38774, n38775, n38776, n38777, n38778, n38779,
    n38780, n38781, n38782, n38783, n38784, n38785,
    n38786, n38787, n38788, n38789, n38790, n38791,
    n38792, n38793, n38794, n38795, n38796, n38797,
    n38798, n38799, n38800, n38801, n38802, n38803,
    n38804, n38805, n38806, n38807, n38808, n38809,
    n38810, n38811, n38812, n38813, n38814, n38815,
    n38816, n38817, n38818, n38819, n38820, n38821,
    n38822, n38823, n38824, n38825, n38826, n38827,
    n38828, n38829, n38830, n38831, n38832, n38833,
    n38834, n38835, n38836, n38837, n38838, n38839,
    n38840, n38841, n38842, n38843, n38844, n38845,
    n38846, n38847, n38848, n38849, n38850, n38851,
    n38852, n38853, n38854, n38855, n38856, n38857,
    n38858, n38859, n38860, n38861, n38862, n38863,
    n38864, n38865, n38866, n38867, n38868, n38869,
    n38870, n38871, n38872, n38873, n38874, n38875,
    n38876, n38877, n38878, n38879, n38880, n38881,
    n38882, n38883, n38884, n38885, n38886, n38887,
    n38888, n38889, n38890, n38891, n38892, n38893,
    n38894, n38895, n38896, n38897, n38898, n38899,
    n38900, n38901, n38902, n38903, n38904, n38905,
    n38906, n38907, n38908, n38909, n38910, n38911,
    n38912, n38913, n38914, n38915, n38916, n38917,
    n38918, n38919, n38920, n38921, n38922, n38923,
    n38924, n38925, n38926, n38927, n38928, n38929,
    n38930, n38931, n38932, n38933, n38934, n38935,
    n38936, n38937, n38938, n38939, n38940, n38941,
    n38942, n38943, n38944, n38945, n38946, n38947,
    n38948, n38949, n38950, n38951, n38952, n38953,
    n38954, n38955, n38956, n38957, n38958, n38959,
    n38960, n38961, n38962, n38963, n38964, n38965,
    n38966, n38967, n38968, n38969, n38970, n38971,
    n38972, n38973, n38974, n38975, n38976, n38977,
    n38978, n38979, n38980, n38981, n38982, n38983,
    n38984, n38985, n38986, n38987, n38988, n38989,
    n38990, n38991, n38992, n38993, n38994, n38995,
    n38996, n38997, n38998, n38999, n39000, n39001,
    n39002, n39003, n39004, n39005, n39006, n39007,
    n39008, n39009, n39010, n39011, n39012, n39013,
    n39014, n39015, n39016, n39017, n39018, n39019,
    n39020, n39021, n39022, n39023, n39024, n39025,
    n39026, n39027, n39028, n39029, n39030, n39031,
    n39032, n39033, n39034, n39035, n39036, n39037,
    n39038, n39039, n39040, n39041, n39042, n39043,
    n39044, n39045, n39046, n39047, n39048, n39049,
    n39050, n39051, n39052, n39053, n39054, n39055,
    n39056, n39057, n39058, n39059, n39060, n39061,
    n39062, n39063, n39064, n39065, n39066, n39067,
    n39068, n39069, n39070, n39071, n39072, n39073,
    n39074, n39075, n39076, n39077, n39078, n39079,
    n39080, n39081, n39082, n39083, n39084, n39085,
    n39086, n39087, n39088, n39089, n39090, n39091,
    n39092, n39093, n39094, n39095, n39096, n39097,
    n39098, n39099, n39100, n39101, n39102, n39103,
    n39104, n39105, n39106, n39107, n39108, n39109,
    n39110, n39111, n39112, n39113, n39114, n39115,
    n39116, n39117, n39118, n39119, n39120, n39121,
    n39122, n39123, n39124, n39125, n39126, n39127,
    n39128, n39129, n39130, n39131, n39132, n39133,
    n39134, n39135, n39136, n39137, n39138, n39139,
    n39140, n39141, n39142, n39143, n39144, n39145,
    n39146, n39147, n39148, n39149, n39150, n39151,
    n39152, n39153, n39154, n39155, n39156, n39157,
    n39158, n39159, n39160, n39161, n39162, n39163,
    n39164, n39165, n39166, n39167, n39168, n39169,
    n39170, n39171, n39172, n39173, n39174, n39175,
    n39176, n39177, n39178, n39179, n39180, n39181,
    n39182, n39183, n39184, n39185, n39186, n39187,
    n39188, n39189, n39190, n39191, n39192, n39193,
    n39194, n39195, n39196, n39197, n39198, n39199,
    n39200, n39201, n39202, n39203, n39204, n39205,
    n39206, n39207, n39208, n39209, n39210, n39211,
    n39212, n39213, n39214, n39215, n39216, n39217,
    n39218, n39219, n39220, n39221, n39222, n39223,
    n39224, n39225, n39226, n39227, n39228, n39229,
    n39230, n39231, n39232, n39233, n39234, n39235,
    n39236, n39237, n39238, n39239, n39240, n39241,
    n39242, n39243, n39244, n39245, n39246, n39247,
    n39248, n39249, n39250, n39251, n39252, n39253,
    n39254, n39255, n39256, n39257, n39258, n39259,
    n39260, n39261, n39262, n39263, n39264, n39265,
    n39266, n39267, n39268, n39269, n39270, n39271,
    n39272, n39273, n39274, n39275, n39276, n39277,
    n39278, n39279, n39280, n39281, n39282, n39283,
    n39284, n39285, n39286, n39287, n39288, n39289,
    n39290, n39291, n39292, n39293, n39294, n39295,
    n39296, n39297, n39298, n39299, n39300, n39301,
    n39302, n39303, n39304, n39305, n39306, n39307,
    n39308, n39309, n39310, n39311, n39312, n39313,
    n39314, n39315, n39316, n39317, n39318, n39319,
    n39320, n39321, n39322, n39323, n39324, n39325,
    n39326, n39327, n39328, n39329, n39330, n39331,
    n39332, n39333, n39334, n39335, n39336, n39337,
    n39338, n39339, n39340, n39341, n39342, n39343,
    n39344, n39345, n39346, n39347, n39348, n39349,
    n39350, n39351, n39352, n39353, n39354, n39355,
    n39356, n39357, n39358, n39359, n39360, n39361,
    n39362, n39363, n39364, n39365, n39366, n39367,
    n39368, n39369, n39370, n39371, n39372, n39373,
    n39374, n39375, n39376, n39377, n39378, n39379,
    n39380, n39381, n39382, n39383, n39384, n39385,
    n39386, n39387, n39388, n39389, n39390, n39391,
    n39392, n39393, n39394, n39395, n39396, n39397,
    n39398, n39399, n39400, n39401, n39402, n39403,
    n39404, n39405, n39406, n39407, n39408, n39409,
    n39410, n39411, n39412, n39413, n39414, n39415,
    n39416, n39417, n39418, n39419, n39420, n39421,
    n39422, n39423, n39424, n39425, n39426, n39427,
    n39428, n39429, n39430, n39431, n39432, n39433,
    n39434, n39435, n39436, n39437, n39438, n39439,
    n39440, n39441, n39442, n39443, n39444, n39445,
    n39446, n39447, n39448, n39449, n39450, n39451,
    n39452, n39453, n39454, n39455, n39456, n39457,
    n39458, n39459, n39460, n39461, n39462, n39463,
    n39464, n39465, n39466, n39467, n39468, n39469,
    n39470, n39471, n39472, n39473, n39474, n39475,
    n39476, n39477, n39478, n39479, n39480, n39481,
    n39482, n39483, n39484, n39485, n39486, n39487,
    n39488, n39489, n39490, n39491, n39492, n39493,
    n39494, n39495, n39496, n39497, n39498, n39499,
    n39500, n39501, n39502, n39503, n39504, n39505,
    n39506, n39507, n39508, n39509, n39510, n39511,
    n39512, n39513, n39514, n39515, n39516, n39517,
    n39518, n39519, n39520, n39521, n39522, n39523,
    n39524, n39525, n39526, n39527, n39528, n39529,
    n39530, n39531, n39532, n39533, n39534, n39535,
    n39536, n39537, n39538, n39539, n39540, n39541,
    n39542, n39543, n39544, n39545, n39546, n39547,
    n39548, n39549, n39550, n39551, n39552, n39553,
    n39554, n39555, n39556, n39557, n39558, n39559,
    n39560, n39561, n39562, n39563, n39564, n39565,
    n39566, n39567, n39568, n39569, n39570, n39571,
    n39572, n39573, n39574, n39575, n39576, n39577,
    n39578, n39579, n39580, n39581, n39582, n39583,
    n39584, n39585, n39586, n39587, n39588, n39589,
    n39590, n39591, n39592, n39593, n39594, n39595,
    n39596, n39597, n39598, n39599, n39600, n39601,
    n39602, n39603, n39604, n39605, n39606, n39607,
    n39608, n39609, n39610, n39611, n39612, n39613,
    n39614, n39615, n39616, n39617, n39618, n39619,
    n39620, n39621, n39622, n39623, n39624, n39625,
    n39626, n39627, n39628, n39629, n39630, n39631,
    n39632, n39633, n39634, n39635, n39636, n39637,
    n39638, n39639, n39640, n39641, n39642, n39643,
    n39644, n39645, n39646, n39647, n39648, n39649,
    n39650, n39651, n39652, n39653, n39654, n39655,
    n39656, n39657, n39658, n39659, n39660, n39661,
    n39662, n39663, n39664, n39665, n39666, n39667,
    n39668, n39669, n39670, n39671, n39672, n39673,
    n39674, n39675, n39676, n39677, n39678, n39679,
    n39680, n39681, n39682, n39683, n39684, n39685,
    n39686, n39687, n39688, n39689, n39690, n39691,
    n39692, n39693, n39694, n39695, n39696, n39697,
    n39698, n39699, n39700, n39701, n39702, n39703,
    n39704, n39705, n39706, n39707, n39708, n39709,
    n39710, n39711, n39712, n39713, n39714, n39715,
    n39716, n39717, n39718, n39719, n39720, n39721,
    n39722, n39723, n39724, n39725, n39726, n39727,
    n39728, n39729, n39730, n39731, n39732, n39733,
    n39734, n39735, n39736, n39737, n39738, n39739,
    n39740, n39741, n39742, n39743, n39744, n39745,
    n39746, n39747, n39748, n39749, n39750, n39751,
    n39752, n39753, n39754, n39755, n39756, n39757,
    n39758, n39759, n39760, n39761, n39762, n39763,
    n39764, n39765, n39766, n39767, n39768, n39769,
    n39770, n39771, n39772, n39773, n39774, n39775,
    n39776, n39777, n39778, n39779, n39780, n39781,
    n39782, n39783, n39784, n39785, n39786, n39787,
    n39788, n39789, n39790, n39791, n39792, n39793,
    n39794, n39795, n39796, n39797, n39798, n39799,
    n39800, n39801, n39802, n39803, n39804, n39805,
    n39806, n39807, n39808, n39809, n39810, n39811,
    n39812, n39813, n39814, n39815, n39816, n39817,
    n39818, n39819, n39820, n39821, n39822, n39823,
    n39824, n39825, n39826, n39827, n39828, n39829,
    n39830, n39831, n39832, n39833, n39834, n39835,
    n39836, n39837, n39838, n39839, n39840, n39841,
    n39842, n39843, n39844, n39845, n39846, n39847,
    n39848, n39849, n39850, n39851, n39852, n39853,
    n39854, n39855, n39856, n39857, n39858, n39859,
    n39860, n39861, n39862, n39863, n39864, n39865,
    n39866, n39867, n39868, n39869, n39870, n39871,
    n39872, n39873, n39874, n39875, n39876, n39877,
    n39878, n39879, n39880, n39881, n39882, n39883,
    n39884, n39885, n39886, n39887, n39888, n39889,
    n39890, n39891, n39892, n39893, n39894, n39895,
    n39896, n39897, n39898, n39899, n39900, n39901,
    n39902, n39903, n39904, n39905, n39906, n39907,
    n39908, n39909, n39910, n39911, n39912, n39913,
    n39914, n39915, n39916, n39917, n39918, n39919,
    n39920, n39921, n39922, n39923, n39924, n39925,
    n39926, n39927, n39928, n39929, n39930, n39931,
    n39932, n39933, n39934, n39935, n39936, n39937,
    n39938, n39939, n39940, n39941, n39942, n39943,
    n39944, n39945, n39946, n39947, n39948, n39949,
    n39950, n39951, n39952, n39953, n39954, n39955,
    n39956, n39957, n39958, n39959, n39960, n39961,
    n39962, n39963, n39964, n39965, n39966, n39967,
    n39968, n39969, n39970, n39971, n39972, n39973,
    n39974, n39975, n39976, n39977, n39978, n39979,
    n39980, n39981, n39982, n39983, n39984, n39985,
    n39986, n39987, n39988, n39989, n39990, n39991,
    n39992, n39993, n39994, n39995, n39996, n39997,
    n39998, n39999, n40000, n40001, n40002, n40003,
    n40004, n40005, n40006, n40007, n40008, n40009,
    n40010, n40011, n40012, n40013, n40014, n40015,
    n40016, n40017, n40018, n40019, n40020, n40021,
    n40022, n40023, n40024, n40025, n40026, n40027,
    n40028, n40029, n40030, n40031, n40032, n40033,
    n40034, n40035, n40036, n40037, n40038, n40039,
    n40040, n40041, n40042, n40043, n40044, n40045,
    n40046, n40047, n40048, n40049, n40050, n40051,
    n40052, n40053, n40054, n40055, n40056, n40057,
    n40058, n40059, n40060, n40061, n40062, n40063,
    n40064, n40065, n40066, n40067, n40068, n40069,
    n40070, n40071, n40072, n40073, n40074, n40075,
    n40076, n40077, n40078, n40079, n40080, n40081,
    n40082, n40083, n40084, n40085, n40086, n40087,
    n40088, n40089, n40090, n40091, n40092, n40093,
    n40094, n40095, n40096, n40097, n40098, n40099,
    n40100, n40101, n40102, n40103, n40104, n40105,
    n40106, n40107, n40108, n40109, n40110, n40111,
    n40112, n40113, n40114, n40115, n40116, n40117,
    n40118, n40119, n40120, n40121, n40122, n40123,
    n40124, n40125, n40126, n40127, n40128, n40129,
    n40130, n40131, n40132, n40133, n40134, n40135,
    n40136, n40137, n40138, n40139, n40140, n40141,
    n40142, n40143, n40144, n40145, n40146, n40147,
    n40148, n40149, n40150, n40151, n40152, n40153,
    n40154, n40155, n40156, n40157, n40158, n40159,
    n40160, n40161, n40162, n40163, n40164, n40165,
    n40166, n40167, n40168, n40169, n40170, n40171,
    n40172, n40173, n40174, n40175, n40176, n40177,
    n40178, n40179, n40180, n40181, n40182, n40183,
    n40184, n40185, n40186, n40187, n40188, n40189,
    n40190, n40191, n40192, n40193, n40194, n40195,
    n40196, n40197, n40198, n40199, n40200, n40201,
    n40202, n40203, n40204, n40205, n40206, n40207,
    n40208, n40209, n40210, n40211, n40212, n40213,
    n40214, n40215, n40216, n40217, n40218, n40219,
    n40220, n40221, n40222, n40223, n40224, n40225,
    n40226, n40227, n40228, n40229, n40230, n40231,
    n40232, n40233, n40234, n40235, n40236, n40237,
    n40238, n40239, n40240, n40241, n40242, n40243,
    n40244, n40245, n40246, n40247, n40248, n40249,
    n40250, n40251, n40252, n40253, n40254, n40255,
    n40256, n40257, n40258, n40259, n40260, n40261,
    n40262, n40263, n40264, n40265, n40266, n40267,
    n40268, n40269, n40270, n40271, n40272, n40273,
    n40274, n40275, n40276, n40277, n40278, n40279,
    n40280, n40281, n40282, n40283, n40284, n40285,
    n40286, n40287, n40288, n40289, n40290, n40291,
    n40292, n40293, n40294, n40295, n40296, n40297,
    n40298, n40299, n40300, n40301, n40302, n40303,
    n40304, n40305, n40306, n40307, n40308, n40309,
    n40310, n40311, n40312, n40313, n40314, n40315,
    n40316, n40317, n40318, n40319, n40320, n40321,
    n40322, n40323, n40324, n40325, n40326, n40327,
    n40328, n40329, n40330, n40331, n40332, n40333,
    n40334, n40335, n40336, n40337, n40338, n40339,
    n40340, n40341, n40342, n40343, n40344, n40345,
    n40346, n40347, n40348, n40349, n40350, n40351,
    n40352, n40353, n40354, n40355, n40356, n40357,
    n40358, n40359, n40360, n40361, n40362, n40363,
    n40364, n40365, n40366, n40367, n40368, n40369,
    n40370, n40371, n40372, n40373, n40374, n40375,
    n40376, n40377, n40378, n40379, n40380, n40381,
    n40382, n40383, n40384, n40385, n40386, n40387,
    n40388, n40389, n40390, n40391, n40392, n40393,
    n40394, n40395, n40396, n40397, n40398, n40399,
    n40400, n40401, n40402, n40403, n40404, n40405,
    n40406, n40407, n40408, n40409, n40410, n40411,
    n40412, n40413, n40414, n40415, n40416, n40417,
    n40418, n40419, n40420, n40421, n40422, n40423,
    n40424, n40425, n40426, n40427, n40428, n40429,
    n40430, n40431, n40432, n40433, n40434, n40435,
    n40436, n40437, n40438, n40439, n40440, n40441,
    n40442, n40443, n40444, n40445, n40446, n40447,
    n40448, n40449, n40450, n40451, n40452, n40453,
    n40454, n40455, n40456, n40457, n40458, n40459,
    n40460, n40461, n40462, n40463, n40464, n40465,
    n40466, n40467, n40468, n40469, n40470, n40471,
    n40472, n40473, n40474, n40475, n40476, n40477,
    n40478, n40479, n40480, n40481, n40482, n40483,
    n40484, n40485, n40486, n40487, n40488, n40489,
    n40490, n40491, n40492, n40493, n40494, n40495,
    n40496, n40497, n40498, n40499, n40500, n40501,
    n40502, n40503, n40504, n40505, n40506, n40507,
    n40508, n40509, n40510, n40511, n40512, n40513,
    n40514, n40515, n40516, n40517, n40518, n40519,
    n40520, n40521, n40522, n40523, n40524, n40525,
    n40526, n40527, n40528, n40529, n40530, n40531,
    n40532, n40533, n40534, n40535, n40536, n40537,
    n40538, n40539, n40540, n40541, n40542, n40543,
    n40544, n40545, n40546, n40547, n40548, n40549,
    n40550, n40551, n40552, n40553, n40554, n40555,
    n40556, n40557, n40558, n40559, n40560, n40561,
    n40562, n40563, n40564, n40565, n40566, n40567,
    n40568, n40569, n40570, n40571, n40572, n40573,
    n40574, n40575, n40576, n40577, n40578, n40579,
    n40580, n40581, n40582, n40583, n40584, n40585,
    n40586, n40587, n40588, n40589, n40590, n40591,
    n40592, n40593, n40594, n40595, n40596, n40597,
    n40598, n40599, n40600, n40601, n40602, n40603,
    n40604, n40605, n40606, n40607, n40608, n40609,
    n40610, n40611, n40612, n40613, n40614, n40615,
    n40616, n40617, n40618, n40619, n40620, n40621,
    n40622, n40623, n40624, n40625, n40626, n40627,
    n40628, n40629, n40630, n40631, n40632, n40633,
    n40634, n40635, n40636, n40637, n40638, n40639,
    n40640, n40641, n40642, n40643, n40644, n40645,
    n40646, n40647, n40648, n40649, n40650, n40651,
    n40652, n40653, n40654, n40655, n40656, n40657,
    n40658, n40659, n40660, n40661, n40662, n40663,
    n40664, n40665, n40666, n40667, n40668, n40669,
    n40670, n40671, n40672, n40673, n40674, n40675,
    n40676, n40677, n40678, n40679, n40680, n40681,
    n40682, n40683, n40684, n40685, n40686, n40687,
    n40688, n40689, n40690, n40691, n40692, n40693,
    n40694, n40695, n40696, n40697, n40698, n40699,
    n40700, n40701, n40702, n40703, n40704, n40705,
    n40706, n40707, n40708, n40709, n40710, n40711,
    n40712, n40713, n40714, n40715, n40716, n40717,
    n40718, n40719, n40720, n40721, n40722, n40723,
    n40724, n40725, n40726, n40727, n40728, n40729,
    n40730, n40731, n40732, n40733, n40734, n40735,
    n40736, n40737, n40738, n40739, n40740, n40741,
    n40742, n40743, n40744, n40745, n40746, n40747,
    n40748, n40749, n40750, n40751, n40752, n40753,
    n40754, n40755, n40756, n40757, n40758, n40759,
    n40760, n40761, n40762, n40763, n40764, n40765,
    n40766, n40767, n40768, n40769, n40770, n40771,
    n40772, n40773, n40774, n40775, n40776, n40777,
    n40778, n40779, n40780, n40781, n40782, n40783,
    n40784, n40785, n40786, n40787, n40788, n40789,
    n40790, n40791, n40792, n40793, n40794, n40795,
    n40796, n40797, n40798, n40799, n40800, n40801,
    n40802, n40803, n40804, n40805, n40806, n40807,
    n40808, n40809, n40810, n40811, n40812, n40813,
    n40814, n40815, n40816, n40817, n40818, n40819,
    n40820, n40821, n40822, n40823, n40824, n40825,
    n40826, n40827, n40828, n40829, n40830, n40831,
    n40832, n40833, n40834, n40835, n40836, n40837,
    n40838, n40839, n40840, n40841, n40842, n40843,
    n40844, n40845, n40846, n40847, n40848, n40849,
    n40850, n40851, n40852, n40853, n40854, n40855,
    n40856, n40857, n40858, n40859, n40860, n40861,
    n40862, n40863, n40864, n40865, n40866, n40867,
    n40868, n40869, n40870, n40871, n40872, n40873,
    n40874, n40875, n40876, n40877, n40878, n40879,
    n40880, n40881, n40882, n40883, n40884, n40885,
    n40886, n40887, n40888, n40889, n40890, n40891,
    n40892, n40893, n40894, n40895, n40896, n40897,
    n40898, n40899, n40900, n40901, n40902, n40903,
    n40904, n40905, n40906, n40907, n40908, n40909,
    n40910, n40911, n40912, n40913, n40914, n40915,
    n40916, n40917, n40918, n40919, n40920, n40921,
    n40922, n40923, n40924, n40925, n40926, n40927,
    n40928, n40929, n40930, n40931, n40932, n40933,
    n40934, n40935, n40936, n40937, n40938, n40939,
    n40940, n40941, n40942, n40943, n40944, n40945,
    n40946, n40947, n40948, n40949, n40950, n40951,
    n40952, n40953, n40954, n40955, n40956, n40957,
    n40958, n40959, n40960, n40961, n40962, n40963,
    n40964, n40965, n40966, n40967, n40968, n40969,
    n40970, n40971, n40972, n40973, n40974, n40975,
    n40976, n40977, n40978, n40979, n40980, n40981,
    n40982, n40983, n40984, n40985, n40986, n40987,
    n40988, n40989, n40990, n40991, n40992, n40993,
    n40994, n40995, n40996, n40997, n40998, n40999,
    n41000, n41001, n41002, n41003, n41004, n41005,
    n41006, n41007, n41008, n41009, n41010, n41011,
    n41012, n41013, n41014, n41015, n41016, n41017,
    n41018, n41019, n41020, n41021, n41022, n41023,
    n41024, n41025, n41026, n41027, n41028, n41029,
    n41030, n41031, n41032, n41033, n41034, n41035,
    n41036, n41037, n41038, n41039, n41040, n41041,
    n41042, n41043, n41044, n41045, n41046, n41047,
    n41048, n41049, n41050, n41051, n41052, n41053,
    n41054, n41055, n41056, n41057, n41058, n41059,
    n41060, n41061, n41062, n41063, n41064, n41065,
    n41066, n41067, n41068, n41069, n41070, n41071,
    n41072, n41073, n41074, n41075, n41076, n41077,
    n41078, n41079, n41080, n41081, n41082, n41083,
    n41084, n41085, n41086, n41087, n41088, n41089,
    n41090, n41091, n41092, n41093, n41094, n41095,
    n41096, n41097, n41098, n41099, n41100, n41101,
    n41102, n41103, n41104, n41105, n41106, n41107,
    n41108, n41109, n41110, n41111, n41112, n41113,
    n41114, n41115, n41116, n41117, n41118, n41119,
    n41120, n41121, n41122, n41123, n41124, n41125,
    n41126, n41127, n41128, n41129, n41130, n41131,
    n41132, n41133, n41134, n41135, n41136, n41137,
    n41138, n41139, n41140, n41141, n41142, n41143,
    n41144, n41145, n41146, n41147, n41148, n41149,
    n41150, n41151, n41152, n41153, n41154, n41155,
    n41156, n41157, n41158, n41159, n41160, n41161,
    n41162, n41163, n41164, n41165, n41166, n41167,
    n41168, n41169, n41170, n41171, n41172, n41173,
    n41174, n41175, n41176, n41177, n41178, n41179,
    n41180, n41181, n41182, n41183, n41184, n41185,
    n41186, n41187, n41188, n41189, n41190, n41191,
    n41192, n41193, n41194, n41195, n41196, n41197,
    n41198, n41199, n41200, n41201, n41202, n41203,
    n41204, n41205, n41206, n41207, n41208, n41209,
    n41210, n41211, n41212, n41213, n41214, n41215,
    n41216, n41217, n41218, n41219, n41220, n41221,
    n41222, n41223, n41224, n41225, n41226, n41227,
    n41228, n41229, n41230, n41231, n41232, n41233,
    n41234, n41235, n41236, n41237, n41238, n41239,
    n41240, n41241, n41242, n41243, n41244, n41245,
    n41246, n41247, n41248, n41249, n41250, n41251,
    n41252, n41253, n41254, n41255, n41256, n41257,
    n41258, n41259, n41260, n41261, n41262, n41263,
    n41264, n41265, n41266, n41267, n41268, n41269,
    n41270, n41271, n41272, n41273, n41274, n41275,
    n41276, n41277, n41278, n41279, n41280, n41281,
    n41282, n41283, n41284, n41285, n41286, n41287,
    n41288, n41289, n41290, n41291, n41292, n41293,
    n41294, n41295, n41296, n41297, n41298, n41299,
    n41300, n41301, n41302, n41303, n41304, n41305,
    n41306, n41307, n41308, n41309, n41310, n41311,
    n41312, n41313, n41314, n41315, n41316, n41317,
    n41318, n41319, n41320, n41321, n41322, n41323,
    n41324, n41325, n41326, n41327, n41328, n41329,
    n41330, n41331, n41332, n41333, n41334, n41335,
    n41336, n41337, n41338, n41339, n41340, n41341,
    n41342, n41343, n41344, n41345, n41346, n41347,
    n41348, n41349, n41350, n41351, n41352, n41353,
    n41354, n41355, n41356, n41357, n41358, n41359,
    n41360, n41361, n41362, n41363, n41364, n41365,
    n41366, n41367, n41368, n41369, n41370, n41371,
    n41372, n41373, n41374, n41375, n41376, n41377,
    n41378, n41379, n41380, n41381, n41382, n41383,
    n41384, n41385, n41386, n41387, n41388, n41389,
    n41390, n41391, n41392, n41393, n41394, n41395,
    n41396, n41397, n41398, n41399, n41400, n41401,
    n41402, n41403, n41404, n41405, n41406, n41407,
    n41408, n41409, n41410, n41411, n41412, n41413,
    n41414, n41415, n41416, n41417, n41418, n41419,
    n41420, n41421, n41422, n41423, n41424, n41425,
    n41426, n41427, n41428, n41429, n41430, n41431,
    n41432, n41433, n41434, n41435, n41436, n41437,
    n41438, n41439, n41440, n41441, n41442, n41443,
    n41444, n41445, n41446, n41447, n41448, n41449,
    n41450, n41451, n41452, n41453, n41454, n41455,
    n41456, n41457, n41458, n41459, n41460, n41461,
    n41462, n41463, n41464, n41465, n41466, n41467,
    n41468, n41469, n41470, n41471, n41472, n41473,
    n41474, n41475, n41476, n41477, n41478, n41479,
    n41480, n41481, n41482, n41483, n41484, n41485,
    n41486, n41487, n41488, n41489, n41490, n41491,
    n41492, n41493, n41494, n41495, n41496, n41497,
    n41498, n41499, n41500, n41501, n41502, n41503,
    n41504, n41505, n41506, n41507, n41508, n41509,
    n41510, n41511, n41512, n41513, n41514, n41515,
    n41516, n41517, n41518, n41519, n41520, n41521,
    n41522, n41523, n41524, n41525, n41526, n41527,
    n41528, n41529, n41530, n41531, n41532, n41533,
    n41534, n41535, n41536, n41537, n41538, n41539,
    n41540, n41541, n41542, n41543, n41544, n41545,
    n41546, n41547, n41548, n41549, n41550, n41551,
    n41552, n41553, n41554, n41555, n41556, n41557,
    n41558, n41559, n41560, n41561, n41562, n41563,
    n41564, n41565, n41566, n41567, n41568, n41569,
    n41570, n41571, n41572, n41573, n41574, n41575,
    n41576, n41577, n41578, n41579, n41580, n41581,
    n41582, n41583, n41584, n41585, n41586, n41587,
    n41588, n41589, n41590, n41591, n41592, n41593,
    n41594, n41595, n41596, n41597, n41598, n41599,
    n41600, n41601, n41602, n41603, n41604, n41605,
    n41606, n41607, n41608, n41609, n41610, n41611,
    n41612, n41613, n41614, n41615, n41616, n41617,
    n41618, n41619, n41620, n41621, n41622, n41623,
    n41624, n41625, n41626, n41627, n41628, n41629,
    n41630, n41631, n41632, n41633, n41634, n41635,
    n41636, n41637, n41638, n41639, n41640, n41641,
    n41642, n41643, n41644, n41645, n41646, n41647,
    n41648, n41649, n41650, n41651, n41652, n41653,
    n41654, n41655, n41656, n41657, n41658, n41659,
    n41660, n41661, n41662, n41663, n41664, n41665,
    n41666, n41667, n41668, n41669, n41670, n41671,
    n41672, n41673, n41674, n41675, n41676, n41677,
    n41678, n41679, n41680, n41681, n41682, n41683,
    n41684, n41685, n41686, n41687, n41688, n41689,
    n41690, n41691, n41692, n41693, n41694, n41695,
    n41696, n41697, n41698, n41699, n41700, n41701,
    n41702, n41703, n41704, n41705, n41706, n41707,
    n41708, n41709, n41710, n41711, n41712, n41713,
    n41714, n41715, n41716, n41717, n41718, n41719,
    n41720, n41721, n41722, n41723, n41724, n41725,
    n41726, n41727, n41728, n41729, n41730, n41731,
    n41732, n41733, n41734, n41735, n41736, n41737,
    n41738, n41739, n41740, n41741, n41742, n41743,
    n41744, n41745, n41746, n41747, n41748, n41749,
    n41750, n41751, n41752, n41753, n41754, n41755,
    n41756, n41757, n41758, n41759, n41760, n41761,
    n41762, n41763, n41764, n41765, n41766, n41767,
    n41768, n41769, n41770, n41771, n41772, n41773,
    n41774, n41775, n41776, n41777, n41778, n41779,
    n41780, n41781, n41782, n41783, n41784, n41785,
    n41786, n41787, n41788, n41789, n41790, n41791,
    n41792, n41793, n41794, n41795, n41796, n41797,
    n41798, n41799, n41800, n41801, n41802, n41803,
    n41804, n41805, n41806, n41807, n41808, n41809,
    n41810, n41811, n41812, n41813, n41814, n41815,
    n41816, n41817, n41818, n41819, n41820, n41821,
    n41822, n41823, n41824, n41825, n41826, n41827,
    n41828, n41829, n41830, n41831, n41832, n41833,
    n41834, n41835, n41836, n41837, n41838, n41839,
    n41840, n41841, n41842, n41843, n41844, n41845,
    n41846, n41847, n41848, n41849, n41850, n41851,
    n41852, n41853, n41854, n41855, n41856, n41857,
    n41858, n41859, n41860, n41861, n41862, n41863,
    n41864, n41865, n41866, n41867, n41868, n41869,
    n41870, n41871, n41872, n41873, n41874, n41875,
    n41876, n41877, n41878, n41879, n41880, n41881,
    n41882, n41883, n41884, n41885, n41886, n41887,
    n41888, n41889, n41890, n41891, n41892, n41893,
    n41894, n41895, n41896, n41897, n41898, n41899,
    n41900, n41901, n41902, n41903, n41904, n41905,
    n41906, n41907, n41908, n41909, n41910, n41911,
    n41912, n41913, n41914, n41915, n41916, n41917,
    n41918, n41919, n41920, n41921, n41922, n41923,
    n41924, n41925, n41926, n41927, n41928, n41929,
    n41930, n41931, n41932, n41933, n41934, n41935,
    n41936, n41937, n41938, n41939, n41940, n41941,
    n41942, n41943, n41944, n41945, n41946, n41947,
    n41948, n41949, n41950, n41951, n41952, n41953,
    n41954, n41955, n41956, n41957, n41958, n41959,
    n41960, n41961, n41962, n41963, n41964, n41965,
    n41966, n41967, n41968, n41969, n41970, n41971,
    n41972, n41973, n41974, n41975, n41976, n41977,
    n41978, n41979, n41980, n41981, n41982, n41983,
    n41984, n41985, n41986, n41987, n41988, n41989,
    n41990, n41991, n41992, n41993, n41994, n41995,
    n41996, n41997, n41998, n41999, n42000, n42001,
    n42002, n42003, n42004, n42005, n42006, n42007,
    n42008, n42009, n42010, n42011, n42012, n42013,
    n42014, n42015, n42016, n42017, n42018, n42019,
    n42020, n42021, n42022, n42023, n42024, n42025,
    n42026, n42027, n42028, n42029, n42030, n42031,
    n42032, n42033, n42034, n42035, n42036, n42037,
    n42038, n42039, n42040, n42041, n42042, n42043,
    n42044, n42045, n42046, n42047, n42048, n42049,
    n42050, n42051, n42052, n42053, n42054, n42055,
    n42056, n42057, n42058, n42059, n42060, n42061,
    n42062, n42063, n42064, n42065, n42066, n42067,
    n42068, n42069, n42070, n42071, n42072, n42073,
    n42074, n42075, n42076, n42077, n42078, n42079,
    n42080, n42081, n42082, n42083, n42084, n42085,
    n42086, n42087, n42088, n42089, n42090, n42091,
    n42092, n42093, n42094, n42095, n42096, n42097,
    n42098, n42099, n42100, n42101, n42102, n42103,
    n42104, n42105, n42106, n42107, n42108, n42109,
    n42110, n42111, n42112, n42113, n42114, n42115,
    n42116, n42117, n42118, n42119, n42120, n42121,
    n42122, n42123, n42124, n42125, n42126, n42127,
    n42128, n42129, n42130, n42131, n42132, n42133,
    n42134, n42135, n42136, n42137, n42138, n42139,
    n42140, n42141, n42142, n42143, n42144, n42145,
    n42146, n42147, n42148, n42149, n42150, n42151,
    n42152, n42153, n42154, n42155, n42156, n42157,
    n42158, n42159, n42160, n42161, n42162, n42163,
    n42164, n42165, n42166, n42167, n42168, n42169,
    n42170, n42171, n42172, n42173, n42174, n42175,
    n42176, n42177, n42178, n42179, n42180, n42181,
    n42182, n42183, n42184, n42185, n42186, n42187,
    n42188, n42189, n42190, n42191, n42192, n42193,
    n42194, n42195, n42196, n42197, n42198, n42199,
    n42200, n42201, n42202, n42203, n42204, n42205,
    n42206, n42207, n42208, n42209, n42210, n42211,
    n42212, n42213, n42214, n42215, n42216, n42217,
    n42218, n42219, n42220, n42221, n42222, n42223,
    n42224, n42225, n42226, n42227, n42228, n42229,
    n42230, n42231, n42232, n42233, n42234, n42235,
    n42236, n42237, n42238, n42239, n42240, n42241,
    n42242, n42243, n42244, n42245, n42246, n42247,
    n42248, n42249, n42250, n42251, n42252, n42253,
    n42254, n42255, n42256, n42257, n42258, n42259,
    n42260, n42261, n42262, n42263, n42264, n42265,
    n42266, n42267, n42268, n42269, n42270, n42271,
    n42272, n42273, n42274, n42275, n42276, n42277,
    n42278, n42279, n42280, n42281, n42282, n42283,
    n42284, n42285, n42286, n42287, n42288, n42289,
    n42290, n42291, n42292, n42293, n42294, n42295,
    n42296, n42297, n42298, n42299, n42300, n42301,
    n42302, n42303, n42304, n42305, n42306, n42307,
    n42308, n42309, n42310, n42311, n42312, n42313,
    n42314, n42315, n42316, n42317, n42318, n42319,
    n42320, n42321, n42322, n42323, n42324, n42325,
    n42326, n42327, n42328, n42329, n42330, n42331,
    n42332, n42333, n42334, n42335, n42336, n42337,
    n42338, n42339, n42340, n42341, n42342, n42343,
    n42344, n42345, n42346, n42347, n42348, n42349,
    n42350, n42351, n42352, n42353, n42354, n42355,
    n42356, n42357, n42358, n42359, n42360, n42361,
    n42362, n42363, n42364, n42365, n42366, n42367,
    n42368, n42369, n42370, n42371, n42372, n42373,
    n42374, n42375, n42376, n42377, n42378, n42379,
    n42380, n42381, n42382, n42383, n42384, n42385,
    n42386, n42387, n42388, n42389, n42390, n42391,
    n42392, n42393, n42394, n42395, n42396, n42397,
    n42398, n42399, n42400, n42401, n42402, n42403,
    n42404, n42405, n42406, n42407, n42408, n42409,
    n42410, n42411, n42412, n42413, n42414, n42415,
    n42416, n42417, n42418, n42419, n42420, n42421,
    n42422, n42423, n42424, n42425, n42426, n42427,
    n42428, n42429, n42430, n42431, n42432, n42433,
    n42434, n42435, n42436, n42437, n42438, n42439,
    n42440, n42441, n42442, n42443, n42444, n42445,
    n42446, n42447, n42448, n42449, n42450, n42451,
    n42452, n42453, n42454, n42455, n42456, n42457,
    n42458, n42459, n42460, n42461, n42462, n42463,
    n42464, n42465, n42466, n42467, n42468, n42469,
    n42470, n42471, n42472, n42473, n42474, n42475,
    n42476, n42477, n42478, n42479, n42480, n42481,
    n42482, n42483, n42484, n42485, n42486, n42487,
    n42488, n42489, n42490, n42491, n42492, n42493,
    n42494, n42495, n42496, n42497, n42498, n42499,
    n42500, n42501, n42502, n42503, n42504, n42505,
    n42506, n42507, n42508, n42509, n42510, n42511,
    n42512, n42513, n42514, n42515, n42516, n42517,
    n42518, n42519, n42520, n42521, n42522, n42523,
    n42524, n42525, n42526, n42527, n42528, n42529,
    n42530, n42531, n42532, n42533, n42534, n42535,
    n42536, n42537, n42538, n42539, n42540, n42541,
    n42542, n42543, n42544, n42545, n42546, n42547,
    n42548, n42549, n42550, n42551, n42552, n42553,
    n42554, n42555, n42556, n42557, n42558, n42559,
    n42560, n42561, n42562, n42563, n42564, n42565,
    n42566, n42567, n42568, n42569, n42570, n42571,
    n42572, n42573, n42574, n42575, n42576, n42577,
    n42578, n42579, n42580, n42581, n42582, n42583,
    n42584, n42585, n42586, n42587, n42588, n42589,
    n42590, n42591, n42592, n42593, n42594, n42595,
    n42596, n42597, n42598, n42599, n42600, n42601,
    n42602, n42603, n42604, n42605, n42606, n42607,
    n42608, n42609, n42610, n42611, n42612, n42613,
    n42614, n42615, n42616, n42617, n42618, n42619,
    n42620, n42621, n42622, n42623, n42624, n42625,
    n42626, n42627, n42628, n42629, n42630, n42631,
    n42632, n42633, n42634, n42635, n42636, n42637,
    n42638, n42639, n42640, n42641, n42642, n42643,
    n42644, n42645, n42646, n42647, n42648, n42649,
    n42650, n42651, n42652, n42653, n42654, n42655,
    n42656, n42657, n42658, n42659, n42660, n42661,
    n42662, n42663, n42664, n42665, n42666, n42667,
    n42668, n42669, n42670, n42671, n42672, n42673,
    n42674, n42675, n42676, n42677, n42678, n42679,
    n42680, n42681, n42682, n42683, n42684, n42685,
    n42686, n42687, n42688, n42689, n42690, n42691,
    n42692, n42693, n42694, n42695, n42696, n42697,
    n42698, n42699, n42700, n42701, n42702, n42703,
    n42704, n42705, n42706, n42707, n42708, n42709,
    n42710, n42711, n42712, n42713, n42714, n42715,
    n42716, n42717, n42718, n42719, n42720, n42721,
    n42722, n42723, n42724, n42725, n42726, n42727,
    n42728, n42729, n42730, n42731, n42732, n42733,
    n42734, n42735, n42736, n42737, n42738, n42739,
    n42740, n42741, n42742, n42743, n42744, n42745,
    n42746, n42747, n42748, n42749, n42750, n42751,
    n42752, n42753, n42754, n42755, n42756, n42757,
    n42758, n42759, n42760, n42761, n42762, n42763,
    n42764, n42765, n42766, n42767, n42768, n42769,
    n42770, n42771, n42772, n42773, n42774, n42775,
    n42776, n42777, n42778, n42779, n42780, n42781,
    n42782, n42783, n42784, n42785, n42786, n42787,
    n42788, n42789, n42790, n42791, n42792, n42793,
    n42794, n42795, n42796, n42797, n42798, n42799,
    n42800, n42801, n42802, n42803, n42804, n42805,
    n42806, n42807, n42808, n42809, n42810, n42811,
    n42812, n42813, n42814, n42815, n42816, n42817,
    n42818, n42819, n42820, n42821, n42822, n42823,
    n42824, n42825, n42826, n42827, n42828, n42829,
    n42830, n42831, n42832, n42833, n42834, n42835,
    n42836, n42837, n42838, n42839, n42840, n42841,
    n42842, n42843, n42844, n42845, n42846, n42847,
    n42848, n42849, n42850, n42851, n42852, n42853,
    n42854, n42855, n42856, n42857, n42858, n42859,
    n42860, n42861, n42862, n42863, n42864, n42865,
    n42866, n42867, n42868, n42869, n42870, n42871,
    n42872, n42873, n42874, n42875, n42876, n42877,
    n42878, n42879, n42880, n42881, n42882, n42883,
    n42884, n42885, n42886, n42887, n42888, n42889,
    n42890, n42891, n42892, n42893, n42894, n42895,
    n42896, n42897, n42898, n42899, n42900, n42901,
    n42902, n42903, n42904, n42905, n42906, n42907,
    n42908, n42909, n42910, n42911, n42912, n42913,
    n42914, n42915, n42916, n42917, n42918, n42919,
    n42920, n42921, n42922, n42923, n42924, n42925,
    n42926, n42927, n42928, n42929, n42930, n42931,
    n42932, n42933, n42934, n42935, n42936, n42937,
    n42938, n42939, n42940, n42941, n42942, n42943,
    n42944, n42945, n42946, n42947, n42948, n42949,
    n42950, n42951, n42952, n42953, n42954, n42955,
    n42956, n42957, n42958, n42959, n42960, n42961,
    n42962, n42963, n42964, n42965, n42966, n42967,
    n42968, n42969, n42970, n42971, n42972, n42973,
    n42974, n42975, n42976, n42977, n42978, n42979,
    n42980, n42981, n42982, n42983, n42984, n42985,
    n42986, n42987, n42988, n42989, n42990, n42991,
    n42992, n42993, n42994, n42995, n42996, n42997,
    n42998, n42999, n43000, n43001, n43002, n43003,
    n43004, n43005, n43006, n43007, n43008, n43009,
    n43010, n43011, n43012, n43013, n43014, n43015,
    n43016, n43017, n43018, n43019, n43020, n43021,
    n43022, n43023, n43024, n43025, n43026, n43027,
    n43028, n43029, n43030, n43031, n43032, n43033,
    n43034, n43035, n43036, n43037, n43038, n43039,
    n43040, n43041, n43042, n43043, n43044, n43045,
    n43046, n43047, n43048, n43049, n43050, n43051,
    n43052, n43053, n43054, n43055, n43056, n43057,
    n43058, n43059, n43060, n43061, n43062, n43063,
    n43064, n43065, n43066, n43067, n43068, n43069,
    n43070, n43071, n43072, n43073, n43074, n43075,
    n43076, n43077, n43078, n43079, n43080, n43081,
    n43082, n43083, n43084, n43085, n43086, n43087,
    n43088, n43089, n43090, n43091, n43092, n43093,
    n43094, n43095, n43096, n43097, n43098, n43099,
    n43100, n43101, n43102, n43103, n43104, n43105,
    n43106, n43107, n43108, n43109, n43110, n43111,
    n43112, n43113, n43114, n43115, n43116, n43117,
    n43118, n43119, n43120, n43121, n43122, n43123,
    n43124, n43125, n43126, n43127, n43128, n43129,
    n43130, n43131, n43132, n43133, n43134, n43135,
    n43136, n43137, n43138, n43139, n43140, n43141,
    n43142, n43143, n43144, n43145, n43146, n43147,
    n43148, n43149, n43150, n43151, n43152, n43153,
    n43154, n43155, n43156, n43157, n43158, n43159,
    n43160, n43161, n43162, n43163, n43164, n43165,
    n43166, n43167, n43168, n43169, n43170, n43171,
    n43172, n43173, n43174, n43175, n43176, n43177,
    n43178, n43179, n43180, n43181, n43182, n43183,
    n43184, n43185, n43186, n43187, n43188, n43189,
    n43190, n43191, n43192, n43193, n43194, n43195,
    n43196, n43197, n43198, n43199, n43200, n43201,
    n43202, n43203, n43204, n43205, n43206, n43207,
    n43208, n43209, n43210, n43211, n43212, n43213,
    n43214, n43215, n43216, n43217, n43218, n43219,
    n43220, n43221, n43222, n43223, n43224, n43225,
    n43226, n43227, n43228, n43229, n43230, n43231,
    n43232, n43233, n43234, n43235, n43236, n43237,
    n43238, n43239, n43240, n43241, n43242, n43243,
    n43244, n43245, n43246, n43247, n43248, n43249,
    n43250, n43251, n43252, n43253, n43254, n43255,
    n43256, n43257, n43258, n43259, n43260, n43261,
    n43262, n43263, n43264, n43265, n43266, n43267,
    n43268, n43269, n43270, n43271, n43272, n43273,
    n43274, n43275, n43276, n43277, n43278, n43279,
    n43280, n43281, n43282, n43283, n43284, n43285,
    n43286, n43287, n43288, n43289, n43290, n43291,
    n43292, n43293, n43294, n43295, n43296, n43297,
    n43298, n43299, n43300, n43301, n43302, n43303,
    n43304, n43305, n43306, n43307, n43308, n43309,
    n43310, n43311, n43312, n43313, n43314, n43315,
    n43316, n43317, n43318, n43319, n43320, n43321,
    n43322, n43323, n43324, n43325, n43326, n43327,
    n43328, n43329, n43330, n43331, n43332, n43333,
    n43334, n43335, n43336, n43337, n43338, n43339,
    n43340, n43341, n43342, n43343, n43344, n43345,
    n43346, n43347, n43348, n43349, n43350, n43351,
    n43352, n43353, n43354, n43355, n43356, n43357,
    n43358, n43359, n43360, n43361, n43362, n43363,
    n43364, n43365, n43366, n43367, n43368, n43369,
    n43370, n43371, n43372, n43373, n43374, n43375,
    n43376, n43377, n43378, n43379, n43380, n43381,
    n43382, n43383, n43384, n43385, n43386, n43387,
    n43388, n43389, n43390, n43391, n43392, n43393,
    n43394, n43395, n43396, n43397, n43398, n43399,
    n43400, n43401, n43402, n43403, n43404, n43405,
    n43406, n43407, n43408, n43409, n43410, n43411,
    n43412, n43413, n43414, n43415, n43416, n43417,
    n43418, n43419, n43420, n43421, n43422, n43423,
    n43424, n43425, n43426, n43427, n43428, n43429,
    n43430, n43431, n43432, n43433, n43434, n43435,
    n43436, n43437, n43438, n43439, n43440, n43441,
    n43442, n43443, n43444, n43445, n43446, n43447,
    n43448, n43449, n43450, n43451, n43452, n43453,
    n43454, n43455, n43456, n43457, n43458, n43459,
    n43460, n43461, n43462, n43463, n43464, n43465,
    n43466, n43467, n43468, n43469, n43470, n43471,
    n43472, n43473, n43474, n43475, n43476, n43477,
    n43478, n43479, n43480, n43481, n43482, n43483,
    n43484, n43485, n43486, n43487, n43488, n43489,
    n43490, n43491, n43492, n43493, n43494, n43495,
    n43496, n43497, n43498, n43499, n43500, n43501,
    n43502, n43503, n43504, n43505, n43506, n43507,
    n43508, n43509, n43510, n43511, n43512, n43513,
    n43514, n43515, n43516, n43517, n43518, n43519,
    n43520, n43521, n43522, n43523, n43524, n43525,
    n43526, n43527, n43528, n43529, n43530, n43531,
    n43532, n43533, n43534, n43535, n43536, n43537,
    n43538, n43539, n43540, n43541, n43542, n43543,
    n43544, n43545, n43546, n43547, n43548, n43549,
    n43550, n43551, n43552, n43553, n43554, n43555,
    n43556, n43557, n43558, n43559, n43560, n43561,
    n43562, n43563, n43564, n43565, n43566, n43567,
    n43568, n43569, n43570, n43571, n43572, n43573,
    n43574, n43575, n43576, n43577, n43578, n43579,
    n43580, n43581, n43582, n43583, n43584, n43585,
    n43586, n43587, n43588, n43589, n43590, n43591,
    n43592, n43593, n43594, n43595, n43596, n43597,
    n43598, n43599, n43600, n43601, n43602, n43603,
    n43604, n43605, n43606, n43607, n43608, n43609,
    n43610, n43611, n43612, n43613, n43614, n43615,
    n43616, n43617, n43618, n43619, n43620, n43621,
    n43622, n43623, n43624, n43625, n43626, n43627,
    n43628, n43629, n43630, n43631, n43632, n43633,
    n43634, n43635, n43636, n43637, n43638, n43639,
    n43640, n43641, n43642, n43643, n43644, n43645,
    n43646, n43647, n43648, n43649, n43650, n43651,
    n43652, n43653, n43654, n43655, n43656, n43657,
    n43658, n43659, n43660, n43661, n43662, n43663,
    n43664, n43665, n43666, n43667, n43668, n43669,
    n43670, n43671, n43672, n43673, n43674, n43675,
    n43676, n43677, n43678, n43679, n43680, n43681,
    n43682, n43683, n43684, n43685, n43686, n43687,
    n43688, n43689, n43690, n43691, n43692, n43693,
    n43694, n43695, n43696, n43697, n43698, n43699,
    n43700, n43701, n43702, n43703, n43704, n43705,
    n43706, n43707, n43708, n43709, n43710, n43711,
    n43712, n43713, n43714, n43715, n43716, n43717,
    n43718, n43719, n43720, n43721, n43722, n43723,
    n43724, n43725, n43726, n43727, n43728, n43729,
    n43730, n43731, n43732, n43733, n43734, n43735,
    n43736, n43737, n43738, n43739, n43740, n43741,
    n43742, n43743, n43744, n43745, n43746, n43747,
    n43748, n43749, n43750, n43751, n43752, n43753,
    n43754, n43755, n43756, n43757, n43758, n43759,
    n43760, n43761, n43762, n43763, n43764, n43765,
    n43766, n43767, n43768, n43769, n43770, n43771,
    n43772, n43773, n43774, n43775, n43776, n43777,
    n43778, n43779, n43780, n43781, n43782, n43783,
    n43784, n43785, n43786, n43787, n43788, n43789,
    n43790, n43791, n43792, n43793, n43794, n43795,
    n43796, n43797, n43798, n43799, n43800, n43801,
    n43802, n43803, n43804, n43805, n43806, n43807,
    n43808, n43809, n43810, n43811, n43812, n43813,
    n43814, n43815, n43816, n43817, n43818, n43819,
    n43820, n43821, n43822, n43823, n43824, n43825,
    n43826, n43827, n43828, n43829, n43830, n43831,
    n43832, n43833, n43834, n43835, n43836, n43837,
    n43838, n43839, n43840, n43841, n43842, n43843,
    n43844, n43845, n43846, n43847, n43848, n43849,
    n43850, n43851, n43852, n43853, n43854, n43855,
    n43856, n43857, n43858, n43859, n43860, n43861,
    n43862, n43863, n43864, n43865, n43866, n43867,
    n43868, n43869, n43870, n43871, n43872, n43873,
    n43874, n43875, n43876, n43877, n43878, n43879,
    n43880, n43881, n43882, n43883, n43884, n43885,
    n43886, n43887, n43888, n43889, n43890, n43891,
    n43892, n43893, n43894, n43895, n43896, n43897,
    n43898, n43899, n43900, n43901, n43902, n43903,
    n43904, n43905, n43906, n43907, n43908, n43909,
    n43910, n43911, n43912, n43913, n43914, n43915,
    n43916, n43917, n43918, n43919, n43920, n43921,
    n43922, n43923, n43924, n43925, n43926, n43927,
    n43928, n43929, n43930, n43931, n43932, n43933,
    n43934, n43935, n43936, n43937, n43938, n43939,
    n43940, n43941, n43942, n43943, n43944, n43945,
    n43946, n43947, n43948, n43949, n43950, n43951,
    n43952, n43953, n43954, n43955, n43956, n43957,
    n43958, n43959, n43960, n43961, n43962, n43963,
    n43964, n43965, n43966, n43967, n43968, n43969,
    n43970, n43971, n43972, n43973, n43974, n43975,
    n43976, n43977, n43978, n43979, n43980, n43981,
    n43982, n43983, n43984, n43985, n43986, n43987,
    n43988, n43989, n43990, n43991, n43992, n43993,
    n43994, n43995, n43996, n43997, n43998, n43999,
    n44000, n44001, n44002, n44003, n44004, n44005,
    n44006, n44007, n44008, n44009, n44010, n44011,
    n44012, n44013, n44014, n44015, n44016, n44017,
    n44018, n44019, n44020, n44021, n44022, n44023,
    n44024, n44025, n44026, n44027, n44028, n44029,
    n44030, n44031, n44032, n44033, n44034, n44035,
    n44036, n44037, n44038, n44039, n44040, n44041,
    n44042, n44043, n44044, n44045, n44046, n44047,
    n44048, n44049, n44050, n44051, n44052, n44053,
    n44054, n44055, n44056, n44057, n44058, n44059,
    n44060, n44061, n44062, n44063, n44064, n44065,
    n44066, n44067, n44068, n44069, n44070, n44071,
    n44072, n44073, n44074, n44075, n44076, n44077,
    n44078, n44079, n44080, n44081, n44082, n44083,
    n44084, n44085, n44086, n44087, n44088, n44089,
    n44090, n44091, n44092, n44093, n44094, n44095,
    n44096, n44097, n44098, n44099, n44100, n44101,
    n44102, n44103, n44104, n44105, n44106, n44107,
    n44108, n44109, n44110, n44111, n44112, n44113,
    n44114, n44115, n44116, n44117, n44118, n44119,
    n44120, n44121, n44122, n44123, n44124, n44125,
    n44126, n44127, n44128, n44129, n44130, n44131,
    n44132, n44133, n44134, n44135, n44136, n44137,
    n44138, n44139, n44140, n44141, n44142, n44143,
    n44144, n44145, n44146, n44147, n44148, n44149,
    n44150, n44151, n44152, n44153, n44154, n44155,
    n44156, n44157, n44158, n44159, n44160, n44161,
    n44162, n44163, n44164, n44165, n44166, n44167,
    n44168, n44169, n44170, n44171, n44172, n44173,
    n44174, n44175, n44176, n44177, n44178, n44179,
    n44180, n44181, n44182, n44183, n44184, n44185,
    n44186, n44187, n44188, n44189, n44190, n44191,
    n44192, n44193, n44194, n44195, n44196, n44197,
    n44198, n44199, n44200, n44201, n44202, n44203,
    n44204, n44205, n44206, n44207, n44208, n44209,
    n44210, n44211, n44212, n44213, n44214, n44215,
    n44216, n44217, n44218, n44219, n44220, n44221,
    n44222, n44223, n44224, n44225, n44226, n44227,
    n44228, n44229, n44230, n44231, n44232, n44233,
    n44234, n44235, n44236, n44237, n44238, n44239,
    n44240, n44241, n44242, n44243, n44244, n44245,
    n44246, n44247, n44248, n44249, n44250, n44251,
    n44252, n44253, n44254, n44255, n44256, n44257,
    n44258, n44259, n44260, n44261, n44262, n44263,
    n44264, n44265, n44266, n44267, n44268, n44269,
    n44270, n44271, n44272, n44273, n44274, n44275,
    n44276, n44277, n44278, n44279, n44280, n44281,
    n44282, n44283, n44284, n44285, n44286, n44287,
    n44288, n44289, n44290, n44291, n44292, n44293,
    n44294, n44295, n44296, n44297, n44298, n44299,
    n44300, n44301, n44302, n44303, n44304, n44305,
    n44307, n44308;
  assign n257 = pi8  & ~pi9 ;
  assign n258 = ~pi8  & pi9 ;
  assign n259 = ~pi8  & ~pi9 ;
  assign n260 = pi8  & pi9 ;
  assign n261 = ~n259 & ~n260;
  assign n262 = ~n257 & ~n258;
  assign n263 = pi10  & ~pi11 ;
  assign n264 = ~pi10  & pi11 ;
  assign n265 = ~pi10  & ~pi11 ;
  assign n266 = pi10  & pi11 ;
  assign n267 = ~n265 & ~n266;
  assign n268 = ~n263 & ~n264;
  assign n269 = n37470 & n37471;
  assign n270 = pi113  & pi114 ;
  assign n271 = pi112  & pi113 ;
  assign n272 = pi111  & pi112 ;
  assign n273 = pi110  & pi111 ;
  assign n274 = pi109  & pi110 ;
  assign n275 = pi108  & pi109 ;
  assign n276 = pi107  & pi108 ;
  assign n277 = pi106  & pi107 ;
  assign n278 = pi105  & pi106 ;
  assign n279 = pi104  & pi105 ;
  assign n280 = pi103  & pi104 ;
  assign n281 = pi102  & pi103 ;
  assign n282 = pi101  & pi102 ;
  assign n283 = pi100  & pi101 ;
  assign n284 = pi99  & pi100 ;
  assign n285 = pi98  & pi99 ;
  assign n286 = pi97  & pi98 ;
  assign n287 = pi96  & pi97 ;
  assign n288 = pi95  & pi96 ;
  assign n289 = pi94  & pi95 ;
  assign n290 = pi93  & pi94 ;
  assign n291 = pi92  & pi93 ;
  assign n292 = pi91  & pi92 ;
  assign n293 = pi90  & pi91 ;
  assign n294 = pi89  & pi90 ;
  assign n295 = pi88  & pi89 ;
  assign n296 = pi87  & pi88 ;
  assign n297 = pi86  & pi87 ;
  assign n298 = pi85  & pi86 ;
  assign n299 = pi84  & pi85 ;
  assign n300 = pi83  & pi84 ;
  assign n301 = pi82  & pi83 ;
  assign n302 = pi81  & pi82 ;
  assign n303 = pi80  & pi81 ;
  assign n304 = pi79  & pi80 ;
  assign n305 = pi78  & pi79 ;
  assign n306 = pi77  & pi78 ;
  assign n307 = pi76  & pi77 ;
  assign n308 = pi75  & pi76 ;
  assign n309 = pi74  & pi75 ;
  assign n310 = pi73  & pi74 ;
  assign n311 = pi72  & pi73 ;
  assign n312 = pi71  & pi72 ;
  assign n313 = pi70  & pi71 ;
  assign n314 = pi69  & pi70 ;
  assign n315 = pi68  & pi69 ;
  assign n316 = pi67  & pi68 ;
  assign n317 = pi66  & pi67 ;
  assign n318 = ~pi66  & ~pi67 ;
  assign n319 = ~n317 & ~n318;
  assign n320 = ~pi64  & ~pi66 ;
  assign n321 = pi64  & pi65 ;
  assign n322 = pi64  & ~pi66 ;
  assign n323 = pi65  & n322;
  assign n324 = ~pi66  & n321;
  assign n325 = pi65  & pi66 ;
  assign n326 = ~n37472 & ~n325;
  assign n327 = pi65  & ~n320;
  assign n328 = n319 & ~n37473;
  assign n329 = ~n317 & ~n328;
  assign n330 = ~pi67  & ~pi68 ;
  assign n331 = ~n316 & ~n330;
  assign n332 = ~n329 & n331;
  assign n333 = ~n316 & ~n332;
  assign n334 = ~pi68  & ~pi69 ;
  assign n335 = ~n315 & ~n334;
  assign n336 = ~n333 & n335;
  assign n337 = ~n315 & ~n336;
  assign n338 = ~pi69  & ~pi70 ;
  assign n339 = ~n314 & ~n338;
  assign n340 = ~n337 & n339;
  assign n341 = ~n314 & ~n340;
  assign n342 = ~pi70  & ~pi71 ;
  assign n343 = ~n313 & ~n342;
  assign n344 = ~n341 & n343;
  assign n345 = ~n313 & ~n344;
  assign n346 = ~pi71  & ~pi72 ;
  assign n347 = ~n312 & ~n346;
  assign n348 = ~n345 & n347;
  assign n349 = ~n312 & ~n348;
  assign n350 = ~pi72  & ~pi73 ;
  assign n351 = ~n311 & ~n350;
  assign n352 = ~n349 & n351;
  assign n353 = ~n311 & ~n352;
  assign n354 = ~pi73  & ~pi74 ;
  assign n355 = ~n310 & ~n354;
  assign n356 = ~n353 & n355;
  assign n357 = ~n310 & ~n356;
  assign n358 = ~pi74  & ~pi75 ;
  assign n359 = ~n309 & ~n358;
  assign n360 = ~n357 & n359;
  assign n361 = ~n309 & ~n360;
  assign n362 = ~pi75  & ~pi76 ;
  assign n363 = ~n308 & ~n362;
  assign n364 = ~n361 & n363;
  assign n365 = ~n308 & ~n364;
  assign n366 = ~pi76  & ~pi77 ;
  assign n367 = ~n307 & ~n366;
  assign n368 = ~n365 & n367;
  assign n369 = ~n307 & ~n368;
  assign n370 = ~pi77  & ~pi78 ;
  assign n371 = ~n306 & ~n370;
  assign n372 = ~n369 & n371;
  assign n373 = ~n306 & ~n372;
  assign n374 = ~pi78  & ~pi79 ;
  assign n375 = ~n305 & ~n374;
  assign n376 = ~n373 & n375;
  assign n377 = ~n305 & ~n376;
  assign n378 = ~pi79  & ~pi80 ;
  assign n379 = ~n304 & ~n378;
  assign n380 = ~n377 & n379;
  assign n381 = ~n304 & ~n380;
  assign n382 = ~pi80  & ~pi81 ;
  assign n383 = ~n303 & ~n382;
  assign n384 = ~n381 & n383;
  assign n385 = ~n303 & ~n384;
  assign n386 = ~pi81  & ~pi82 ;
  assign n387 = ~n302 & ~n386;
  assign n388 = ~n385 & n387;
  assign n389 = ~n302 & ~n388;
  assign n390 = ~pi82  & ~pi83 ;
  assign n391 = ~n301 & ~n390;
  assign n392 = ~n389 & n391;
  assign n393 = ~n301 & ~n392;
  assign n394 = ~pi83  & ~pi84 ;
  assign n395 = ~n300 & ~n394;
  assign n396 = ~n393 & n395;
  assign n397 = ~n300 & ~n396;
  assign n398 = ~pi84  & ~pi85 ;
  assign n399 = ~n299 & ~n398;
  assign n400 = ~n397 & n399;
  assign n401 = ~n299 & ~n400;
  assign n402 = ~pi85  & ~pi86 ;
  assign n403 = ~n298 & ~n402;
  assign n404 = ~n401 & n403;
  assign n405 = ~n298 & ~n404;
  assign n406 = ~pi86  & ~pi87 ;
  assign n407 = ~n297 & ~n406;
  assign n408 = ~n405 & n407;
  assign n409 = ~n297 & ~n408;
  assign n410 = ~pi87  & ~pi88 ;
  assign n411 = ~n296 & ~n410;
  assign n412 = ~n409 & n411;
  assign n413 = ~n296 & ~n412;
  assign n414 = ~pi88  & ~pi89 ;
  assign n415 = ~n295 & ~n414;
  assign n416 = ~n413 & n415;
  assign n417 = ~n295 & ~n416;
  assign n418 = ~pi89  & ~pi90 ;
  assign n419 = ~n294 & ~n418;
  assign n420 = ~n417 & n419;
  assign n421 = ~n294 & ~n420;
  assign n422 = ~pi90  & ~pi91 ;
  assign n423 = ~n293 & ~n422;
  assign n424 = ~n421 & n423;
  assign n425 = ~n293 & ~n424;
  assign n426 = ~pi91  & ~pi92 ;
  assign n427 = ~n292 & ~n426;
  assign n428 = ~n425 & n427;
  assign n429 = ~n292 & ~n428;
  assign n430 = ~pi92  & ~pi93 ;
  assign n431 = ~n291 & ~n430;
  assign n432 = ~n429 & n431;
  assign n433 = ~n291 & ~n432;
  assign n434 = ~pi93  & ~pi94 ;
  assign n435 = ~n290 & ~n434;
  assign n436 = ~n433 & n435;
  assign n437 = ~n290 & ~n436;
  assign n438 = ~pi94  & ~pi95 ;
  assign n439 = ~n289 & ~n438;
  assign n440 = ~n437 & n439;
  assign n441 = ~n289 & ~n440;
  assign n442 = ~pi95  & ~pi96 ;
  assign n443 = ~n288 & ~n442;
  assign n444 = ~n441 & n443;
  assign n445 = ~n288 & ~n444;
  assign n446 = ~pi96  & ~pi97 ;
  assign n447 = ~n287 & ~n446;
  assign n448 = ~n445 & n447;
  assign n449 = ~n287 & ~n448;
  assign n450 = ~pi97  & ~pi98 ;
  assign n451 = ~n286 & ~n450;
  assign n452 = ~n449 & n451;
  assign n453 = ~n286 & ~n452;
  assign n454 = ~pi98  & ~pi99 ;
  assign n455 = ~n285 & ~n454;
  assign n456 = ~n453 & n455;
  assign n457 = ~n285 & ~n456;
  assign n458 = ~pi99  & ~pi100 ;
  assign n459 = ~n284 & ~n458;
  assign n460 = ~n457 & n459;
  assign n461 = ~n284 & ~n460;
  assign n462 = ~pi100  & ~pi101 ;
  assign n463 = ~n283 & ~n462;
  assign n464 = ~n461 & n463;
  assign n465 = ~n283 & ~n464;
  assign n466 = ~pi101  & ~pi102 ;
  assign n467 = ~n282 & ~n466;
  assign n468 = ~n465 & n467;
  assign n469 = ~n282 & ~n468;
  assign n470 = ~pi102  & ~pi103 ;
  assign n471 = ~n281 & ~n470;
  assign n472 = ~n469 & n471;
  assign n473 = ~n281 & ~n472;
  assign n474 = ~pi103  & ~pi104 ;
  assign n475 = ~n280 & ~n474;
  assign n476 = ~n473 & n475;
  assign n477 = ~n280 & ~n476;
  assign n478 = ~pi104  & ~pi105 ;
  assign n479 = ~n279 & ~n478;
  assign n480 = ~n477 & n479;
  assign n481 = ~n279 & ~n480;
  assign n482 = ~pi105  & ~pi106 ;
  assign n483 = ~n278 & ~n482;
  assign n484 = ~n481 & n483;
  assign n485 = ~n278 & ~n484;
  assign n486 = ~pi106  & ~pi107 ;
  assign n487 = ~n277 & ~n486;
  assign n488 = ~n485 & n487;
  assign n489 = ~n277 & ~n488;
  assign n490 = ~pi107  & ~pi108 ;
  assign n491 = ~n276 & ~n490;
  assign n492 = ~n489 & n491;
  assign n493 = ~n276 & ~n492;
  assign n494 = ~pi108  & ~pi109 ;
  assign n495 = ~n275 & ~n494;
  assign n496 = ~n493 & n495;
  assign n497 = ~n275 & ~n496;
  assign n498 = ~pi109  & ~pi110 ;
  assign n499 = ~n274 & ~n498;
  assign n500 = ~n497 & n499;
  assign n501 = ~n274 & ~n500;
  assign n502 = ~pi110  & ~pi111 ;
  assign n503 = ~n273 & ~n502;
  assign n504 = ~n501 & n503;
  assign n505 = ~n273 & ~n504;
  assign n506 = ~pi111  & ~pi112 ;
  assign n507 = ~n272 & ~n506;
  assign n508 = ~n505 & n507;
  assign n509 = ~n272 & ~n508;
  assign n510 = ~pi112  & ~pi113 ;
  assign n511 = ~n271 & ~n510;
  assign n512 = ~n509 & n511;
  assign n513 = ~n271 & ~n512;
  assign n514 = ~pi113  & ~pi114 ;
  assign n515 = ~n270 & ~n514;
  assign n516 = ~n513 & n515;
  assign n517 = ~n270 & ~n516;
  assign n518 = ~pi114  & ~pi115 ;
  assign n519 = pi114  & pi115 ;
  assign n520 = ~n518 & ~n519;
  assign n521 = ~n517 & n520;
  assign n522 = n517 & ~n520;
  assign n523 = ~n521 & ~n522;
  assign n524 = n269 & n523;
  assign n525 = pi9  & ~pi10 ;
  assign n526 = ~pi9  & pi10 ;
  assign n527 = ~pi9  & ~pi10 ;
  assign n528 = pi9  & pi10 ;
  assign n529 = ~n527 & ~n528;
  assign n530 = ~n525 & ~n526;
  assign n531 = ~n37470 & n37471;
  assign n532 = ~n37470 & ~n37474;
  assign n533 = n37471 & n532;
  assign n534 = ~n37474 & n531;
  assign n535 = pi113  & n37475;
  assign n536 = n37470 & ~n37471;
  assign n537 = pi115  & n536;
  assign n538 = ~n37470 & n37474;
  assign n539 = pi114  & n538;
  assign n540 = ~n537 & ~n539;
  assign n541 = ~n535 & ~n539;
  assign n542 = ~n537 & n541;
  assign n543 = ~n535 & n540;
  assign n544 = ~n524 & n37476;
  assign n545 = pi11  & ~n544;
  assign n546 = pi11  & ~n545;
  assign n547 = pi11  & n544;
  assign n548 = ~n544 & ~n545;
  assign n549 = ~pi11  & ~n544;
  assign n550 = ~n37477 & ~n37478;
  assign n551 = pi11  & ~pi12 ;
  assign n552 = ~pi11  & pi12 ;
  assign n553 = ~pi11  & ~pi12 ;
  assign n554 = pi11  & pi12 ;
  assign n555 = ~n553 & ~n554;
  assign n556 = ~n551 & ~n552;
  assign n557 = pi13  & ~pi14 ;
  assign n558 = ~pi13  & pi14 ;
  assign n559 = ~pi13  & ~pi14 ;
  assign n560 = pi13  & pi14 ;
  assign n561 = ~n559 & ~n560;
  assign n562 = ~n557 & ~n558;
  assign n563 = n37479 & n37480;
  assign n564 = n501 & ~n503;
  assign n565 = ~n504 & ~n564;
  assign n566 = n563 & n565;
  assign n567 = pi12  & ~pi13 ;
  assign n568 = ~pi12  & pi13 ;
  assign n569 = ~pi12  & ~pi13 ;
  assign n570 = pi12  & pi13 ;
  assign n571 = ~n569 & ~n570;
  assign n572 = ~n567 & ~n568;
  assign n573 = ~n37479 & n37480;
  assign n574 = ~n37479 & ~n37481;
  assign n575 = n37480 & n574;
  assign n576 = ~n37481 & n573;
  assign n577 = pi109  & n37482;
  assign n578 = n37479 & ~n37480;
  assign n579 = pi111  & n578;
  assign n580 = ~n37479 & n37481;
  assign n581 = pi110  & n580;
  assign n582 = ~n579 & ~n581;
  assign n583 = ~n577 & ~n581;
  assign n584 = ~n579 & n583;
  assign n585 = ~n577 & n582;
  assign n586 = ~n566 & n37483;
  assign n587 = pi14  & ~n586;
  assign n588 = pi14  & ~n587;
  assign n589 = pi14  & n586;
  assign n590 = ~n586 & ~n587;
  assign n591 = ~pi14  & ~n586;
  assign n592 = ~n37484 & ~n37485;
  assign n593 = n421 & ~n423;
  assign n594 = ~n424 & ~n593;
  assign n595 = pi26  & ~pi27 ;
  assign n596 = ~pi26  & pi27 ;
  assign n597 = ~pi26  & ~pi27 ;
  assign n598 = pi26  & pi27 ;
  assign n599 = ~n597 & ~n598;
  assign n600 = ~n595 & ~n596;
  assign n601 = pi28  & ~pi29 ;
  assign n602 = ~pi28  & pi29 ;
  assign n603 = ~pi28  & ~pi29 ;
  assign n604 = pi28  & pi29 ;
  assign n605 = ~n603 & ~n604;
  assign n606 = ~n601 & ~n602;
  assign n607 = n37486 & n37487;
  assign n608 = n594 & n607;
  assign n609 = pi27  & ~pi28 ;
  assign n610 = ~pi27  & pi28 ;
  assign n611 = ~pi27  & ~pi28 ;
  assign n612 = pi27  & pi28 ;
  assign n613 = ~n611 & ~n612;
  assign n614 = ~n609 & ~n610;
  assign n615 = ~n37486 & n37487;
  assign n616 = ~n37486 & ~n37488;
  assign n617 = n37487 & n616;
  assign n618 = ~n37488 & n615;
  assign n619 = pi89  & n37489;
  assign n620 = n37486 & ~n37487;
  assign n621 = pi91  & n620;
  assign n622 = ~n37486 & n37488;
  assign n623 = pi90  & n622;
  assign n624 = ~n621 & ~n623;
  assign n625 = ~n619 & ~n623;
  assign n626 = ~n621 & n625;
  assign n627 = ~n619 & n624;
  assign n628 = ~n608 & n37490;
  assign n629 = pi29  & ~n628;
  assign n630 = pi29  & ~n629;
  assign n631 = pi29  & n628;
  assign n632 = ~n628 & ~n629;
  assign n633 = ~pi29  & ~n628;
  assign n634 = ~n37491 & ~n37492;
  assign n635 = n405 & ~n407;
  assign n636 = ~n408 & ~n635;
  assign n637 = pi29  & ~pi30 ;
  assign n638 = ~pi29  & pi30 ;
  assign n639 = ~pi29  & ~pi30 ;
  assign n640 = pi29  & pi30 ;
  assign n641 = ~n639 & ~n640;
  assign n642 = ~n637 & ~n638;
  assign n643 = pi31  & ~pi32 ;
  assign n644 = ~pi31  & pi32 ;
  assign n645 = ~pi31  & ~pi32 ;
  assign n646 = pi31  & pi32 ;
  assign n647 = ~n645 & ~n646;
  assign n648 = ~n643 & ~n644;
  assign n649 = n37493 & n37494;
  assign n650 = n636 & n649;
  assign n651 = pi30  & ~pi31 ;
  assign n652 = ~pi30  & pi31 ;
  assign n653 = ~pi30  & ~pi31 ;
  assign n654 = pi30  & pi31 ;
  assign n655 = ~n653 & ~n654;
  assign n656 = ~n651 & ~n652;
  assign n657 = ~n37493 & n37494;
  assign n658 = ~n37493 & ~n37495;
  assign n659 = n37494 & n658;
  assign n660 = ~n37495 & n657;
  assign n661 = pi85  & n37496;
  assign n662 = n37493 & ~n37494;
  assign n663 = pi87  & n662;
  assign n664 = ~n37493 & n37495;
  assign n665 = pi86  & n664;
  assign n666 = ~n663 & ~n665;
  assign n667 = ~n661 & ~n665;
  assign n668 = ~n663 & n667;
  assign n669 = ~n661 & n666;
  assign n670 = ~n650 & n37497;
  assign n671 = pi32  & ~n670;
  assign n672 = pi32  & ~n671;
  assign n673 = pi32  & n670;
  assign n674 = ~n670 & ~n671;
  assign n675 = ~pi32  & ~n670;
  assign n676 = ~n37498 & ~n37499;
  assign n677 = n373 & ~n375;
  assign n678 = ~n376 & ~n677;
  assign n679 = pi35  & ~pi36 ;
  assign n680 = ~pi35  & pi36 ;
  assign n681 = ~pi35  & ~pi36 ;
  assign n682 = pi35  & pi36 ;
  assign n683 = ~n681 & ~n682;
  assign n684 = ~n679 & ~n680;
  assign n685 = pi37  & ~pi38 ;
  assign n686 = ~pi37  & pi38 ;
  assign n687 = ~pi37  & ~pi38 ;
  assign n688 = pi37  & pi38 ;
  assign n689 = ~n687 & ~n688;
  assign n690 = ~n685 & ~n686;
  assign n691 = n37500 & n37501;
  assign n692 = n678 & n691;
  assign n693 = pi36  & ~pi37 ;
  assign n694 = ~pi36  & pi37 ;
  assign n695 = ~pi36  & ~pi37 ;
  assign n696 = pi36  & pi37 ;
  assign n697 = ~n695 & ~n696;
  assign n698 = ~n693 & ~n694;
  assign n699 = ~n37500 & n37501;
  assign n700 = ~n37500 & ~n37502;
  assign n701 = n37501 & n700;
  assign n702 = ~n37502 & n699;
  assign n703 = pi77  & n37503;
  assign n704 = n37500 & ~n37501;
  assign n705 = pi79  & n704;
  assign n706 = ~n37500 & n37502;
  assign n707 = pi78  & n706;
  assign n708 = ~n705 & ~n707;
  assign n709 = ~n703 & ~n707;
  assign n710 = ~n705 & n709;
  assign n711 = ~n703 & n708;
  assign n712 = ~n692 & n37504;
  assign n713 = pi38  & ~n712;
  assign n714 = pi38  & ~n713;
  assign n715 = pi38  & n712;
  assign n716 = ~n712 & ~n713;
  assign n717 = ~pi38  & ~n712;
  assign n718 = ~n37505 & ~n37506;
  assign n719 = n357 & ~n359;
  assign n720 = ~n360 & ~n719;
  assign n721 = pi38  & ~pi39 ;
  assign n722 = ~pi38  & pi39 ;
  assign n723 = ~pi38  & ~pi39 ;
  assign n724 = pi38  & pi39 ;
  assign n725 = ~n723 & ~n724;
  assign n726 = ~n721 & ~n722;
  assign n727 = pi40  & ~pi41 ;
  assign n728 = ~pi40  & pi41 ;
  assign n729 = ~pi40  & ~pi41 ;
  assign n730 = pi40  & pi41 ;
  assign n731 = ~n729 & ~n730;
  assign n732 = ~n727 & ~n728;
  assign n733 = n37507 & n37508;
  assign n734 = n720 & n733;
  assign n735 = pi39  & ~pi40 ;
  assign n736 = ~pi39  & pi40 ;
  assign n737 = ~pi39  & ~pi40 ;
  assign n738 = pi39  & pi40 ;
  assign n739 = ~n737 & ~n738;
  assign n740 = ~n735 & ~n736;
  assign n741 = ~n37507 & n37508;
  assign n742 = ~n37507 & ~n37509;
  assign n743 = n37508 & n742;
  assign n744 = ~n37509 & n741;
  assign n745 = pi73  & n37510;
  assign n746 = n37507 & ~n37508;
  assign n747 = pi75  & n746;
  assign n748 = ~n37507 & n37509;
  assign n749 = pi74  & n748;
  assign n750 = ~n747 & ~n749;
  assign n751 = ~n745 & ~n749;
  assign n752 = ~n747 & n751;
  assign n753 = ~n745 & n750;
  assign n754 = ~n734 & n37511;
  assign n755 = pi41  & ~n754;
  assign n756 = pi41  & ~n755;
  assign n757 = pi41  & n754;
  assign n758 = ~n754 & ~n755;
  assign n759 = ~pi41  & ~n754;
  assign n760 = ~n37512 & ~n37513;
  assign n761 = pi47  & ~pi48 ;
  assign n762 = ~pi47  & pi48 ;
  assign n763 = ~pi47  & ~pi48 ;
  assign n764 = pi47  & pi48 ;
  assign n765 = ~n763 & ~n764;
  assign n766 = ~n761 & ~n762;
  assign n767 = pi64  & n37514;
  assign n768 = ~pi64  & pi65 ;
  assign n769 = pi64  & ~pi65 ;
  assign n770 = ~pi64  & ~pi65 ;
  assign n771 = ~n321 & ~n770;
  assign n772 = ~n768 & ~n769;
  assign n773 = pi44  & ~pi45 ;
  assign n774 = ~pi44  & pi45 ;
  assign n775 = ~pi44  & ~pi45 ;
  assign n776 = pi44  & pi45 ;
  assign n777 = ~n775 & ~n776;
  assign n778 = ~n773 & ~n774;
  assign n779 = pi46  & ~pi47 ;
  assign n780 = ~pi46  & pi47 ;
  assign n781 = ~pi46  & ~pi47 ;
  assign n782 = pi46  & pi47 ;
  assign n783 = ~n781 & ~n782;
  assign n784 = ~n779 & ~n780;
  assign n785 = n37516 & n37517;
  assign n786 = n37515 & n785;
  assign n787 = n37516 & ~n37517;
  assign n788 = pi65  & n787;
  assign n789 = pi45  & ~pi46 ;
  assign n790 = ~pi45  & pi46 ;
  assign n791 = ~pi45  & ~pi46 ;
  assign n792 = pi45  & pi46 ;
  assign n793 = ~n791 & ~n792;
  assign n794 = ~n789 & ~n790;
  assign n795 = ~n37516 & n37518;
  assign n796 = pi64  & n795;
  assign n797 = ~n788 & ~n796;
  assign n798 = ~n786 & n797;
  assign n799 = pi64  & n37516;
  assign n800 = pi47  & ~n799;
  assign n801 = pi47  & ~n798;
  assign n802 = pi47  & ~n801;
  assign n803 = ~n798 & ~n801;
  assign n804 = ~n802 & ~n803;
  assign n805 = n800 & ~n804;
  assign n806 = n798 & n800;
  assign n807 = ~n37516 & n37517;
  assign n808 = ~n37516 & ~n37518;
  assign n809 = n37517 & n808;
  assign n810 = ~n37518 & n807;
  assign n811 = pi64  & n37520;
  assign n812 = pi65  & n795;
  assign n813 = ~pi66  & ~n768;
  assign n814 = pi66  & n768;
  assign n815 = pi66  & ~n768;
  assign n816 = ~pi66  & n768;
  assign n817 = ~n815 & ~n816;
  assign n818 = ~pi65  & pi66 ;
  assign n819 = pi65  & ~pi66 ;
  assign n820 = ~n321 & ~n819;
  assign n821 = ~n818 & ~n819;
  assign n822 = ~n321 & n821;
  assign n823 = ~n818 & n820;
  assign n824 = ~n37472 & ~n37522;
  assign n825 = ~n813 & ~n814;
  assign n826 = n785 & ~n37521;
  assign n827 = pi66  & n787;
  assign n828 = ~n826 & ~n827;
  assign n829 = ~n812 & ~n826;
  assign n830 = ~n827 & n829;
  assign n831 = ~n812 & ~n827;
  assign n832 = ~n826 & n831;
  assign n833 = ~n812 & n828;
  assign n834 = ~n811 & ~n812;
  assign n835 = ~n827 & n834;
  assign n836 = ~n811 & n831;
  assign n837 = ~n826 & n37524;
  assign n838 = ~n811 & n37523;
  assign n839 = pi47  & ~n37525;
  assign n840 = pi47  & ~n839;
  assign n841 = ~n37525 & ~n839;
  assign n842 = ~n840 & ~n841;
  assign n843 = n37519 & ~n842;
  assign n844 = n37519 & n37525;
  assign n845 = n767 & n37526;
  assign n846 = ~n319 & n37473;
  assign n847 = ~n328 & ~n846;
  assign n848 = n785 & n847;
  assign n849 = pi65  & n37520;
  assign n850 = pi67  & n787;
  assign n851 = pi66  & n795;
  assign n852 = ~n850 & ~n851;
  assign n853 = ~n849 & ~n851;
  assign n854 = ~n850 & n853;
  assign n855 = ~n849 & n852;
  assign n856 = ~n848 & n37527;
  assign n857 = pi47  & ~n856;
  assign n858 = pi47  & ~n857;
  assign n859 = pi47  & n856;
  assign n860 = ~n856 & ~n857;
  assign n861 = ~pi47  & ~n856;
  assign n862 = ~n37528 & ~n37529;
  assign n863 = ~n767 & ~n37526;
  assign n864 = n767 & ~n37526;
  assign n865 = ~n767 & n37526;
  assign n866 = ~n864 & ~n865;
  assign n867 = ~n845 & ~n863;
  assign n868 = ~n862 & ~n37530;
  assign n869 = ~n845 & ~n868;
  assign n870 = n329 & ~n331;
  assign n871 = ~n332 & ~n870;
  assign n872 = n785 & n871;
  assign n873 = pi66  & n37520;
  assign n874 = pi68  & n787;
  assign n875 = pi67  & n795;
  assign n876 = ~n874 & ~n875;
  assign n877 = ~n873 & ~n875;
  assign n878 = ~n874 & n877;
  assign n879 = ~n873 & n876;
  assign n880 = ~n872 & n37531;
  assign n881 = pi47  & ~n880;
  assign n882 = pi47  & ~n881;
  assign n883 = pi47  & n880;
  assign n884 = ~n880 & ~n881;
  assign n885 = ~pi47  & ~n880;
  assign n886 = ~n37532 & ~n37533;
  assign n887 = pi50  & n767;
  assign n888 = pi49  & ~pi50 ;
  assign n889 = ~pi49  & pi50 ;
  assign n890 = ~pi49  & ~pi50 ;
  assign n891 = pi49  & pi50 ;
  assign n892 = ~n890 & ~n891;
  assign n893 = ~n888 & ~n889;
  assign n894 = n37514 & n37534;
  assign n895 = n37515 & n894;
  assign n896 = n37514 & ~n37534;
  assign n897 = pi65  & n896;
  assign n898 = pi48  & ~pi49 ;
  assign n899 = ~pi48  & pi49 ;
  assign n900 = ~pi48  & ~pi49 ;
  assign n901 = pi48  & pi49 ;
  assign n902 = ~n900 & ~n901;
  assign n903 = ~n898 & ~n899;
  assign n904 = ~n37514 & n37535;
  assign n905 = pi64  & n904;
  assign n906 = ~n897 & ~n905;
  assign n907 = ~n895 & n906;
  assign n908 = n887 & ~n907;
  assign n909 = ~n887 & n907;
  assign n910 = pi50  & ~n767;
  assign n911 = pi50  & ~n907;
  assign n912 = pi50  & ~n911;
  assign n913 = ~n907 & ~n911;
  assign n914 = ~n912 & ~n913;
  assign n915 = n910 & ~n914;
  assign n916 = n907 & n910;
  assign n917 = ~n910 & n914;
  assign n918 = ~n37536 & ~n917;
  assign n919 = ~n908 & ~n909;
  assign n920 = n886 & ~n37537;
  assign n921 = ~n886 & n37537;
  assign n922 = ~n920 & ~n921;
  assign n923 = ~n869 & n922;
  assign n924 = n869 & ~n922;
  assign n925 = ~n923 & ~n924;
  assign n926 = n341 & ~n343;
  assign n927 = ~n344 & ~n926;
  assign n928 = pi41  & ~pi42 ;
  assign n929 = ~pi41  & pi42 ;
  assign n930 = ~pi41  & ~pi42 ;
  assign n931 = pi41  & pi42 ;
  assign n932 = ~n930 & ~n931;
  assign n933 = ~n928 & ~n929;
  assign n934 = pi43  & ~pi44 ;
  assign n935 = ~pi43  & pi44 ;
  assign n936 = ~pi43  & ~pi44 ;
  assign n937 = pi43  & pi44 ;
  assign n938 = ~n936 & ~n937;
  assign n939 = ~n934 & ~n935;
  assign n940 = n37538 & n37539;
  assign n941 = n927 & n940;
  assign n942 = pi42  & ~pi43 ;
  assign n943 = ~pi42  & pi43 ;
  assign n944 = ~pi42  & ~pi43 ;
  assign n945 = pi42  & pi43 ;
  assign n946 = ~n944 & ~n945;
  assign n947 = ~n942 & ~n943;
  assign n948 = ~n37538 & n37539;
  assign n949 = ~n37538 & ~n37540;
  assign n950 = n37539 & n949;
  assign n951 = ~n37540 & n948;
  assign n952 = pi69  & n37541;
  assign n953 = n37538 & ~n37539;
  assign n954 = pi71  & n953;
  assign n955 = ~n37538 & n37540;
  assign n956 = pi70  & n955;
  assign n957 = ~n954 & ~n956;
  assign n958 = ~n952 & ~n956;
  assign n959 = ~n954 & n958;
  assign n960 = ~n952 & n957;
  assign n961 = ~n941 & n37542;
  assign n962 = pi44  & ~n961;
  assign n963 = pi44  & ~n962;
  assign n964 = pi44  & n961;
  assign n965 = ~n961 & ~n962;
  assign n966 = ~pi44  & ~n961;
  assign n967 = ~n37543 & ~n37544;
  assign n968 = n925 & ~n967;
  assign n969 = n862 & n37530;
  assign n970 = ~n868 & ~n969;
  assign n971 = n337 & ~n339;
  assign n972 = ~n340 & ~n971;
  assign n973 = n940 & n972;
  assign n974 = pi68  & n37541;
  assign n975 = pi70  & n953;
  assign n976 = pi69  & n955;
  assign n977 = ~n975 & ~n976;
  assign n978 = ~n974 & ~n976;
  assign n979 = ~n975 & n978;
  assign n980 = ~n974 & n977;
  assign n981 = ~n973 & n37545;
  assign n982 = pi44  & ~n981;
  assign n983 = pi44  & ~n982;
  assign n984 = pi44  & n981;
  assign n985 = ~n981 & ~n982;
  assign n986 = ~pi44  & ~n981;
  assign n987 = ~n37546 & ~n37547;
  assign n988 = n970 & ~n987;
  assign n989 = n333 & ~n335;
  assign n990 = ~n336 & ~n989;
  assign n991 = n940 & n990;
  assign n992 = pi67  & n37541;
  assign n993 = pi69  & n953;
  assign n994 = pi68  & n955;
  assign n995 = ~n993 & ~n994;
  assign n996 = ~n992 & ~n994;
  assign n997 = ~n993 & n996;
  assign n998 = ~n992 & n995;
  assign n999 = ~n991 & n37548;
  assign n1000 = pi44  & ~n999;
  assign n1001 = pi44  & ~n1000;
  assign n1002 = pi44  & n999;
  assign n1003 = ~n999 & ~n1000;
  assign n1004 = ~pi44  & ~n999;
  assign n1005 = ~n37549 & ~n37550;
  assign n1006 = pi47  & ~n37519;
  assign n1007 = n37525 & ~n1006;
  assign n1008 = ~n37525 & n1006;
  assign n1009 = ~n37519 & n842;
  assign n1010 = ~n37526 & ~n1009;
  assign n1011 = ~n1007 & ~n1008;
  assign n1012 = ~n1005 & n37551;
  assign n1013 = n871 & n940;
  assign n1014 = pi66  & n37541;
  assign n1015 = pi68  & n953;
  assign n1016 = pi67  & n955;
  assign n1017 = ~n1015 & ~n1016;
  assign n1018 = ~n1014 & ~n1016;
  assign n1019 = ~n1015 & n1018;
  assign n1020 = ~n1014 & n1017;
  assign n1021 = ~n1013 & n37552;
  assign n1022 = pi44  & ~n1021;
  assign n1023 = pi44  & ~n1022;
  assign n1024 = pi44  & n1021;
  assign n1025 = ~n1021 & ~n1022;
  assign n1026 = ~pi44  & ~n1021;
  assign n1027 = ~n37553 & ~n37554;
  assign n1028 = pi47  & n799;
  assign n1029 = ~n798 & n1028;
  assign n1030 = n798 & ~n1028;
  assign n1031 = ~n800 & n804;
  assign n1032 = ~n37519 & ~n1031;
  assign n1033 = ~n1029 & ~n1030;
  assign n1034 = ~n1027 & n37555;
  assign n1035 = n37515 & n940;
  assign n1036 = pi65  & n953;
  assign n1037 = pi64  & n955;
  assign n1038 = ~n1036 & ~n1037;
  assign n1039 = ~n1035 & n1038;
  assign n1040 = pi64  & n37538;
  assign n1041 = pi44  & ~n1040;
  assign n1042 = pi44  & ~n1039;
  assign n1043 = pi44  & ~n1042;
  assign n1044 = ~n1039 & ~n1042;
  assign n1045 = ~n1043 & ~n1044;
  assign n1046 = n1041 & ~n1045;
  assign n1047 = n1039 & n1041;
  assign n1048 = pi64  & n37541;
  assign n1049 = pi65  & n955;
  assign n1050 = ~n37521 & n940;
  assign n1051 = pi66  & n953;
  assign n1052 = ~n1050 & ~n1051;
  assign n1053 = ~n1049 & ~n1050;
  assign n1054 = ~n1051 & n1053;
  assign n1055 = ~n1049 & ~n1051;
  assign n1056 = ~n1050 & n1055;
  assign n1057 = ~n1049 & n1052;
  assign n1058 = ~n1048 & ~n1049;
  assign n1059 = ~n1051 & n1058;
  assign n1060 = ~n1048 & n1055;
  assign n1061 = ~n1050 & n37558;
  assign n1062 = ~n1048 & n37557;
  assign n1063 = pi44  & ~n37559;
  assign n1064 = pi44  & ~n1063;
  assign n1065 = ~n37559 & ~n1063;
  assign n1066 = ~n1064 & ~n1065;
  assign n1067 = n37556 & ~n1066;
  assign n1068 = n37556 & n37559;
  assign n1069 = n799 & n37560;
  assign n1070 = n847 & n940;
  assign n1071 = pi65  & n37541;
  assign n1072 = pi67  & n953;
  assign n1073 = pi66  & n955;
  assign n1074 = ~n1072 & ~n1073;
  assign n1075 = ~n1071 & ~n1073;
  assign n1076 = ~n1072 & n1075;
  assign n1077 = ~n1071 & n1074;
  assign n1078 = ~n1070 & n37561;
  assign n1079 = pi44  & ~n1078;
  assign n1080 = pi44  & ~n1079;
  assign n1081 = pi44  & n1078;
  assign n1082 = ~n1078 & ~n1079;
  assign n1083 = ~pi44  & ~n1078;
  assign n1084 = ~n37562 & ~n37563;
  assign n1085 = ~n799 & ~n37560;
  assign n1086 = n799 & ~n37560;
  assign n1087 = ~n799 & n37560;
  assign n1088 = ~n1086 & ~n1087;
  assign n1089 = ~n1069 & ~n1085;
  assign n1090 = ~n1084 & ~n37564;
  assign n1091 = ~n1069 & ~n1090;
  assign n1092 = n1027 & ~n37555;
  assign n1093 = ~n1034 & ~n1092;
  assign n1094 = ~n1091 & n1093;
  assign n1095 = ~n1034 & ~n1094;
  assign n1096 = n1005 & ~n37551;
  assign n1097 = n37551 & ~n1012;
  assign n1098 = n1005 & n37551;
  assign n1099 = ~n1005 & ~n1012;
  assign n1100 = ~n1005 & ~n37551;
  assign n1101 = ~n37565 & ~n37566;
  assign n1102 = ~n1012 & ~n1096;
  assign n1103 = ~n1095 & ~n37567;
  assign n1104 = ~n1012 & ~n1103;
  assign n1105 = ~n970 & n987;
  assign n1106 = n970 & ~n988;
  assign n1107 = n970 & n987;
  assign n1108 = ~n987 & ~n988;
  assign n1109 = ~n970 & ~n987;
  assign n1110 = ~n37568 & ~n37569;
  assign n1111 = ~n988 & ~n1105;
  assign n1112 = ~n1104 & ~n37570;
  assign n1113 = ~n988 & ~n1112;
  assign n1114 = ~n925 & n967;
  assign n1115 = n925 & ~n968;
  assign n1116 = n925 & n967;
  assign n1117 = ~n967 & ~n968;
  assign n1118 = ~n925 & ~n967;
  assign n1119 = ~n37571 & ~n37572;
  assign n1120 = ~n968 & ~n1114;
  assign n1121 = ~n1113 & ~n37573;
  assign n1122 = ~n968 & ~n1121;
  assign n1123 = n345 & ~n347;
  assign n1124 = ~n348 & ~n1123;
  assign n1125 = n940 & n1124;
  assign n1126 = pi70  & n37541;
  assign n1127 = pi72  & n953;
  assign n1128 = pi71  & n955;
  assign n1129 = ~n1127 & ~n1128;
  assign n1130 = ~n1126 & ~n1128;
  assign n1131 = ~n1127 & n1130;
  assign n1132 = ~n1126 & n1129;
  assign n1133 = ~n1125 & n37574;
  assign n1134 = pi44  & ~n1133;
  assign n1135 = pi44  & ~n1134;
  assign n1136 = pi44  & n1133;
  assign n1137 = ~n1133 & ~n1134;
  assign n1138 = ~pi44  & ~n1133;
  assign n1139 = ~n37575 & ~n37576;
  assign n1140 = ~n921 & ~n923;
  assign n1141 = n785 & n990;
  assign n1142 = pi67  & n37520;
  assign n1143 = pi69  & n787;
  assign n1144 = pi68  & n795;
  assign n1145 = ~n1143 & ~n1144;
  assign n1146 = ~n1142 & ~n1144;
  assign n1147 = ~n1143 & n1146;
  assign n1148 = ~n1142 & n1145;
  assign n1149 = ~n1141 & n37577;
  assign n1150 = pi47  & ~n1149;
  assign n1151 = pi47  & ~n1150;
  assign n1152 = pi47  & n1149;
  assign n1153 = ~n1149 & ~n1150;
  assign n1154 = ~pi47  & ~n1149;
  assign n1155 = ~n37578 & ~n37579;
  assign n1156 = pi50  & ~n37536;
  assign n1157 = ~n37514 & n37534;
  assign n1158 = ~n37514 & ~n37535;
  assign n1159 = n37534 & n1158;
  assign n1160 = ~n37535 & n1157;
  assign n1161 = pi64  & n37580;
  assign n1162 = pi65  & n904;
  assign n1163 = ~n37521 & n894;
  assign n1164 = pi66  & n896;
  assign n1165 = ~n1163 & ~n1164;
  assign n1166 = ~n1162 & ~n1163;
  assign n1167 = ~n1164 & n1166;
  assign n1168 = ~n1162 & ~n1164;
  assign n1169 = ~n1163 & n1168;
  assign n1170 = ~n1162 & n1165;
  assign n1171 = ~n1161 & ~n1162;
  assign n1172 = ~n1164 & n1171;
  assign n1173 = ~n1161 & n1168;
  assign n1174 = ~n1163 & n37582;
  assign n1175 = ~n1161 & n37581;
  assign n1176 = ~n1156 & n37583;
  assign n1177 = n1156 & ~n37583;
  assign n1178 = pi50  & ~n37583;
  assign n1179 = pi50  & ~n1178;
  assign n1180 = ~n37583 & ~n1178;
  assign n1181 = ~n1179 & ~n1180;
  assign n1182 = n37536 & ~n1181;
  assign n1183 = n37536 & n37583;
  assign n1184 = ~n37536 & n1181;
  assign n1185 = ~n37584 & ~n1184;
  assign n1186 = ~n1176 & ~n1177;
  assign n1187 = ~n1155 & n37585;
  assign n1188 = n1155 & ~n37585;
  assign n1189 = n37585 & ~n1187;
  assign n1190 = n1155 & n37585;
  assign n1191 = ~n1155 & ~n1187;
  assign n1192 = ~n1155 & ~n37585;
  assign n1193 = ~n37586 & ~n37587;
  assign n1194 = ~n1187 & ~n1188;
  assign n1195 = ~n1140 & ~n37588;
  assign n1196 = n1140 & n37588;
  assign n1197 = ~n1195 & ~n1196;
  assign n1198 = ~n1139 & n1197;
  assign n1199 = n1139 & ~n1197;
  assign n1200 = ~n1139 & ~n1198;
  assign n1201 = ~n1139 & ~n1197;
  assign n1202 = n1197 & ~n1198;
  assign n1203 = n1139 & n1197;
  assign n1204 = ~n37589 & ~n37590;
  assign n1205 = ~n1198 & ~n1199;
  assign n1206 = ~n1122 & ~n37591;
  assign n1207 = n1122 & n37591;
  assign n1208 = ~n1122 & ~n1206;
  assign n1209 = ~n1122 & n37591;
  assign n1210 = ~n37591 & ~n1206;
  assign n1211 = n1122 & ~n37591;
  assign n1212 = ~n37592 & ~n37593;
  assign n1213 = ~n1206 & ~n1207;
  assign n1214 = ~n760 & ~n37594;
  assign n1215 = n1113 & n37573;
  assign n1216 = ~n1121 & ~n1215;
  assign n1217 = n353 & ~n355;
  assign n1218 = ~n356 & ~n1217;
  assign n1219 = n733 & n1218;
  assign n1220 = pi72  & n37510;
  assign n1221 = pi74  & n746;
  assign n1222 = pi73  & n748;
  assign n1223 = ~n1221 & ~n1222;
  assign n1224 = ~n1220 & ~n1222;
  assign n1225 = ~n1221 & n1224;
  assign n1226 = ~n1220 & n1223;
  assign n1227 = ~n1219 & n37595;
  assign n1228 = pi41  & ~n1227;
  assign n1229 = pi41  & ~n1228;
  assign n1230 = pi41  & n1227;
  assign n1231 = ~n1227 & ~n1228;
  assign n1232 = ~pi41  & ~n1227;
  assign n1233 = ~n37596 & ~n37597;
  assign n1234 = n1216 & ~n1233;
  assign n1235 = n1104 & n37570;
  assign n1236 = ~n1112 & ~n1235;
  assign n1237 = n349 & ~n351;
  assign n1238 = ~n352 & ~n1237;
  assign n1239 = n733 & n1238;
  assign n1240 = pi71  & n37510;
  assign n1241 = pi73  & n746;
  assign n1242 = pi72  & n748;
  assign n1243 = ~n1241 & ~n1242;
  assign n1244 = ~n1240 & ~n1242;
  assign n1245 = ~n1241 & n1244;
  assign n1246 = ~n1240 & n1243;
  assign n1247 = ~n1239 & n37598;
  assign n1248 = pi41  & ~n1247;
  assign n1249 = pi41  & ~n1248;
  assign n1250 = pi41  & n1247;
  assign n1251 = ~n1247 & ~n1248;
  assign n1252 = ~pi41  & ~n1247;
  assign n1253 = ~n37599 & ~n37600;
  assign n1254 = n1236 & ~n1253;
  assign n1255 = n733 & n1124;
  assign n1256 = pi70  & n37510;
  assign n1257 = pi72  & n746;
  assign n1258 = pi71  & n748;
  assign n1259 = ~n1257 & ~n1258;
  assign n1260 = ~n1256 & ~n1258;
  assign n1261 = ~n1257 & n1260;
  assign n1262 = ~n1256 & n1259;
  assign n1263 = ~n1255 & n37601;
  assign n1264 = pi41  & ~n1263;
  assign n1265 = pi41  & ~n1264;
  assign n1266 = pi41  & n1263;
  assign n1267 = ~n1263 & ~n1264;
  assign n1268 = ~pi41  & ~n1263;
  assign n1269 = ~n37602 & ~n37603;
  assign n1270 = n1095 & n37567;
  assign n1271 = ~n1103 & ~n1270;
  assign n1272 = ~n1269 & n1271;
  assign n1273 = n1091 & ~n1093;
  assign n1274 = ~n1094 & ~n1273;
  assign n1275 = n733 & n927;
  assign n1276 = pi69  & n37510;
  assign n1277 = pi71  & n746;
  assign n1278 = pi70  & n748;
  assign n1279 = ~n1277 & ~n1278;
  assign n1280 = ~n1276 & ~n1278;
  assign n1281 = ~n1277 & n1280;
  assign n1282 = ~n1276 & n1279;
  assign n1283 = ~n1275 & n37604;
  assign n1284 = pi41  & ~n1283;
  assign n1285 = pi41  & ~n1284;
  assign n1286 = pi41  & n1283;
  assign n1287 = ~n1283 & ~n1284;
  assign n1288 = ~pi41  & ~n1283;
  assign n1289 = ~n37605 & ~n37606;
  assign n1290 = n1274 & ~n1289;
  assign n1291 = n1084 & n37564;
  assign n1292 = ~n1090 & ~n1291;
  assign n1293 = n733 & n972;
  assign n1294 = pi68  & n37510;
  assign n1295 = pi70  & n746;
  assign n1296 = pi69  & n748;
  assign n1297 = ~n1295 & ~n1296;
  assign n1298 = ~n1294 & ~n1296;
  assign n1299 = ~n1295 & n1298;
  assign n1300 = ~n1294 & n1297;
  assign n1301 = ~n1293 & n37607;
  assign n1302 = pi41  & ~n1301;
  assign n1303 = pi41  & ~n1302;
  assign n1304 = pi41  & n1301;
  assign n1305 = ~n1301 & ~n1302;
  assign n1306 = ~pi41  & ~n1301;
  assign n1307 = ~n37608 & ~n37609;
  assign n1308 = n1292 & ~n1307;
  assign n1309 = n733 & n990;
  assign n1310 = pi67  & n37510;
  assign n1311 = pi69  & n746;
  assign n1312 = pi68  & n748;
  assign n1313 = ~n1311 & ~n1312;
  assign n1314 = ~n1310 & ~n1312;
  assign n1315 = ~n1311 & n1314;
  assign n1316 = ~n1310 & n1313;
  assign n1317 = ~n1309 & n37610;
  assign n1318 = pi41  & ~n1317;
  assign n1319 = pi41  & ~n1318;
  assign n1320 = pi41  & n1317;
  assign n1321 = ~n1317 & ~n1318;
  assign n1322 = ~pi41  & ~n1317;
  assign n1323 = ~n37611 & ~n37612;
  assign n1324 = pi44  & ~n37556;
  assign n1325 = n37559 & ~n1324;
  assign n1326 = ~n37559 & n1324;
  assign n1327 = ~n37556 & n1066;
  assign n1328 = ~n37560 & ~n1327;
  assign n1329 = ~n1325 & ~n1326;
  assign n1330 = ~n1323 & n37613;
  assign n1331 = n733 & n871;
  assign n1332 = pi66  & n37510;
  assign n1333 = pi68  & n746;
  assign n1334 = pi67  & n748;
  assign n1335 = ~n1333 & ~n1334;
  assign n1336 = ~n1332 & ~n1334;
  assign n1337 = ~n1333 & n1336;
  assign n1338 = ~n1332 & n1335;
  assign n1339 = ~n1331 & n37614;
  assign n1340 = pi41  & ~n1339;
  assign n1341 = pi41  & ~n1340;
  assign n1342 = pi41  & n1339;
  assign n1343 = ~n1339 & ~n1340;
  assign n1344 = ~pi41  & ~n1339;
  assign n1345 = ~n37615 & ~n37616;
  assign n1346 = pi44  & n1040;
  assign n1347 = ~n1039 & n1346;
  assign n1348 = n1039 & ~n1346;
  assign n1349 = ~n1041 & n1045;
  assign n1350 = ~n37556 & ~n1349;
  assign n1351 = ~n1347 & ~n1348;
  assign n1352 = ~n1345 & n37617;
  assign n1353 = n733 & n37515;
  assign n1354 = pi65  & n746;
  assign n1355 = pi64  & n748;
  assign n1356 = ~n1354 & ~n1355;
  assign n1357 = ~n1353 & n1356;
  assign n1358 = pi64  & n37507;
  assign n1359 = pi41  & ~n1358;
  assign n1360 = pi41  & ~n1357;
  assign n1361 = pi41  & ~n1360;
  assign n1362 = ~n1357 & ~n1360;
  assign n1363 = ~n1361 & ~n1362;
  assign n1364 = n1359 & ~n1363;
  assign n1365 = n1357 & n1359;
  assign n1366 = pi64  & n37510;
  assign n1367 = pi65  & n748;
  assign n1368 = n733 & ~n37521;
  assign n1369 = pi66  & n746;
  assign n1370 = ~n1368 & ~n1369;
  assign n1371 = ~n1367 & ~n1368;
  assign n1372 = ~n1369 & n1371;
  assign n1373 = ~n1367 & ~n1369;
  assign n1374 = ~n1368 & n1373;
  assign n1375 = ~n1367 & n1370;
  assign n1376 = ~n1366 & ~n1367;
  assign n1377 = ~n1369 & n1376;
  assign n1378 = ~n1366 & n1373;
  assign n1379 = ~n1368 & n37620;
  assign n1380 = ~n1366 & n37619;
  assign n1381 = pi41  & ~n37621;
  assign n1382 = pi41  & ~n1381;
  assign n1383 = ~n37621 & ~n1381;
  assign n1384 = ~n1382 & ~n1383;
  assign n1385 = n37618 & ~n1384;
  assign n1386 = n37618 & n37621;
  assign n1387 = n1040 & n37622;
  assign n1388 = n733 & n847;
  assign n1389 = pi65  & n37510;
  assign n1390 = pi67  & n746;
  assign n1391 = pi66  & n748;
  assign n1392 = ~n1390 & ~n1391;
  assign n1393 = ~n1389 & ~n1391;
  assign n1394 = ~n1390 & n1393;
  assign n1395 = ~n1389 & n1392;
  assign n1396 = ~n1388 & n37623;
  assign n1397 = pi41  & ~n1396;
  assign n1398 = pi41  & ~n1397;
  assign n1399 = pi41  & n1396;
  assign n1400 = ~n1396 & ~n1397;
  assign n1401 = ~pi41  & ~n1396;
  assign n1402 = ~n37624 & ~n37625;
  assign n1403 = ~n1040 & ~n37622;
  assign n1404 = n1040 & ~n37622;
  assign n1405 = ~n1040 & n37622;
  assign n1406 = ~n1404 & ~n1405;
  assign n1407 = ~n1387 & ~n1403;
  assign n1408 = ~n1402 & ~n37626;
  assign n1409 = ~n1387 & ~n1408;
  assign n1410 = n1345 & ~n37617;
  assign n1411 = ~n1352 & ~n1410;
  assign n1412 = ~n1409 & n1411;
  assign n1413 = ~n1352 & ~n1412;
  assign n1414 = n1323 & ~n37613;
  assign n1415 = n37613 & ~n1330;
  assign n1416 = n1323 & n37613;
  assign n1417 = ~n1323 & ~n1330;
  assign n1418 = ~n1323 & ~n37613;
  assign n1419 = ~n37627 & ~n37628;
  assign n1420 = ~n1330 & ~n1414;
  assign n1421 = ~n1413 & ~n37629;
  assign n1422 = ~n1330 & ~n1421;
  assign n1423 = ~n1292 & n1307;
  assign n1424 = n1292 & ~n1308;
  assign n1425 = n1292 & n1307;
  assign n1426 = ~n1307 & ~n1308;
  assign n1427 = ~n1292 & ~n1307;
  assign n1428 = ~n37630 & ~n37631;
  assign n1429 = ~n1308 & ~n1423;
  assign n1430 = ~n1422 & ~n37632;
  assign n1431 = ~n1308 & ~n1430;
  assign n1432 = ~n1274 & n1289;
  assign n1433 = n1274 & ~n1290;
  assign n1434 = n1274 & n1289;
  assign n1435 = ~n1289 & ~n1290;
  assign n1436 = ~n1274 & ~n1289;
  assign n1437 = ~n37633 & ~n37634;
  assign n1438 = ~n1290 & ~n1432;
  assign n1439 = ~n1431 & ~n37635;
  assign n1440 = ~n1290 & ~n1439;
  assign n1441 = n1269 & ~n1271;
  assign n1442 = ~n1269 & ~n1272;
  assign n1443 = ~n1269 & ~n1271;
  assign n1444 = n1271 & ~n1272;
  assign n1445 = n1269 & n1271;
  assign n1446 = ~n37636 & ~n37637;
  assign n1447 = ~n1272 & ~n1441;
  assign n1448 = ~n1440 & ~n37638;
  assign n1449 = ~n1272 & ~n1448;
  assign n1450 = ~n1236 & n1253;
  assign n1451 = ~n1254 & ~n1450;
  assign n1452 = ~n1449 & n1451;
  assign n1453 = ~n1254 & ~n1452;
  assign n1454 = ~n1216 & n1233;
  assign n1455 = ~n1234 & ~n1454;
  assign n1456 = ~n1453 & ~n1454;
  assign n1457 = ~n1234 & n1456;
  assign n1458 = ~n1453 & n1455;
  assign n1459 = ~n1234 & ~n37639;
  assign n1460 = n760 & n37594;
  assign n1461 = ~n1214 & ~n1460;
  assign n1462 = ~n1459 & n1461;
  assign n1463 = ~n1214 & ~n1462;
  assign n1464 = n361 & ~n363;
  assign n1465 = ~n364 & ~n1464;
  assign n1466 = n733 & n1465;
  assign n1467 = pi74  & n37510;
  assign n1468 = pi76  & n746;
  assign n1469 = pi75  & n748;
  assign n1470 = ~n1468 & ~n1469;
  assign n1471 = ~n1467 & ~n1469;
  assign n1472 = ~n1468 & n1471;
  assign n1473 = ~n1467 & n1470;
  assign n1474 = ~n1466 & n37640;
  assign n1475 = pi41  & ~n1474;
  assign n1476 = pi41  & ~n1475;
  assign n1477 = pi41  & n1474;
  assign n1478 = ~n1474 & ~n1475;
  assign n1479 = ~pi41  & ~n1474;
  assign n1480 = ~n37641 & ~n37642;
  assign n1481 = ~n1198 & ~n1206;
  assign n1482 = ~n1187 & ~n1195;
  assign n1483 = n847 & n894;
  assign n1484 = pi65  & n37580;
  assign n1485 = pi67  & n896;
  assign n1486 = pi66  & n904;
  assign n1487 = ~n1485 & ~n1486;
  assign n1488 = ~n1484 & ~n1486;
  assign n1489 = ~n1485 & n1488;
  assign n1490 = ~n1484 & n1487;
  assign n1491 = ~n1483 & n37643;
  assign n1492 = pi50  & ~n1491;
  assign n1493 = pi50  & ~n1492;
  assign n1494 = pi50  & n1491;
  assign n1495 = ~n1491 & ~n1492;
  assign n1496 = ~pi50  & ~n1491;
  assign n1497 = ~n37644 & ~n37645;
  assign n1498 = pi50  & ~pi51 ;
  assign n1499 = ~pi50  & pi51 ;
  assign n1500 = ~pi50  & ~pi51 ;
  assign n1501 = pi50  & pi51 ;
  assign n1502 = ~n1500 & ~n1501;
  assign n1503 = ~n1498 & ~n1499;
  assign n1504 = pi64  & n37646;
  assign n1505 = n37584 & n1504;
  assign n1506 = ~n37584 & ~n1504;
  assign n1507 = ~n37584 & n1504;
  assign n1508 = n37584 & ~n1504;
  assign n1509 = ~n1507 & ~n1508;
  assign n1510 = ~n1505 & ~n1506;
  assign n1511 = ~n1497 & ~n37647;
  assign n1512 = n1497 & n37647;
  assign n1513 = ~n1511 & ~n1512;
  assign n1514 = n785 & n972;
  assign n1515 = pi68  & n37520;
  assign n1516 = pi70  & n787;
  assign n1517 = pi69  & n795;
  assign n1518 = ~n1516 & ~n1517;
  assign n1519 = ~n1515 & ~n1517;
  assign n1520 = ~n1516 & n1519;
  assign n1521 = ~n1515 & n1518;
  assign n1522 = ~n1514 & n37648;
  assign n1523 = pi47  & ~n1522;
  assign n1524 = pi47  & ~n1523;
  assign n1525 = pi47  & n1522;
  assign n1526 = ~n1522 & ~n1523;
  assign n1527 = ~pi47  & ~n1522;
  assign n1528 = ~n37649 & ~n37650;
  assign n1529 = n1513 & ~n1528;
  assign n1530 = ~n1513 & n1528;
  assign n1531 = n1513 & ~n1529;
  assign n1532 = n1513 & n1528;
  assign n1533 = ~n1528 & ~n1529;
  assign n1534 = ~n1513 & ~n1528;
  assign n1535 = ~n37651 & ~n37652;
  assign n1536 = ~n1529 & ~n1530;
  assign n1537 = n1482 & n37653;
  assign n1538 = ~n1482 & ~n37653;
  assign n1539 = ~n1537 & ~n1538;
  assign n1540 = n940 & n1238;
  assign n1541 = pi71  & n37541;
  assign n1542 = pi73  & n953;
  assign n1543 = pi72  & n955;
  assign n1544 = ~n1542 & ~n1543;
  assign n1545 = ~n1541 & ~n1543;
  assign n1546 = ~n1542 & n1545;
  assign n1547 = ~n1541 & n1544;
  assign n1548 = ~n1540 & n37654;
  assign n1549 = pi44  & ~n1548;
  assign n1550 = pi44  & ~n1549;
  assign n1551 = pi44  & n1548;
  assign n1552 = ~n1548 & ~n1549;
  assign n1553 = ~pi44  & ~n1548;
  assign n1554 = ~n37655 & ~n37656;
  assign n1555 = ~n1539 & n1554;
  assign n1556 = n1539 & ~n1554;
  assign n1557 = ~n1555 & ~n1556;
  assign n1558 = ~n1481 & n1557;
  assign n1559 = n1481 & ~n1557;
  assign n1560 = ~n1558 & ~n1559;
  assign n1561 = ~n1480 & n1560;
  assign n1562 = n1480 & ~n1560;
  assign n1563 = ~n1480 & ~n1561;
  assign n1564 = ~n1480 & ~n1560;
  assign n1565 = n1560 & ~n1561;
  assign n1566 = n1480 & n1560;
  assign n1567 = ~n37657 & ~n37658;
  assign n1568 = ~n1561 & ~n1562;
  assign n1569 = ~n1463 & ~n37659;
  assign n1570 = n1463 & ~n37658;
  assign n1571 = ~n37657 & n1570;
  assign n1572 = n1463 & n37659;
  assign n1573 = ~n1569 & ~n37660;
  assign n1574 = ~n718 & n1573;
  assign n1575 = n1459 & ~n1461;
  assign n1576 = ~n1462 & ~n1575;
  assign n1577 = n369 & ~n371;
  assign n1578 = ~n372 & ~n1577;
  assign n1579 = n691 & n1578;
  assign n1580 = pi76  & n37503;
  assign n1581 = pi78  & n704;
  assign n1582 = pi77  & n706;
  assign n1583 = ~n1581 & ~n1582;
  assign n1584 = ~n1580 & ~n1582;
  assign n1585 = ~n1581 & n1584;
  assign n1586 = ~n1580 & n1583;
  assign n1587 = ~n1579 & n37661;
  assign n1588 = pi38  & ~n1587;
  assign n1589 = pi38  & ~n1588;
  assign n1590 = pi38  & n1587;
  assign n1591 = ~n1587 & ~n1588;
  assign n1592 = ~pi38  & ~n1587;
  assign n1593 = ~n37662 & ~n37663;
  assign n1594 = n1576 & ~n1593;
  assign n1595 = n365 & ~n367;
  assign n1596 = ~n368 & ~n1595;
  assign n1597 = n691 & n1596;
  assign n1598 = pi75  & n37503;
  assign n1599 = pi77  & n704;
  assign n1600 = pi76  & n706;
  assign n1601 = ~n1599 & ~n1600;
  assign n1602 = ~n1598 & ~n1600;
  assign n1603 = ~n1599 & n1602;
  assign n1604 = ~n1598 & n1601;
  assign n1605 = ~n1597 & n37664;
  assign n1606 = pi38  & ~n1605;
  assign n1607 = pi38  & ~n1606;
  assign n1608 = pi38  & n1605;
  assign n1609 = ~n1605 & ~n1606;
  assign n1610 = ~pi38  & ~n1605;
  assign n1611 = ~n37665 & ~n37666;
  assign n1612 = n1453 & ~n1455;
  assign n1613 = ~n1453 & ~n37639;
  assign n1614 = ~n1454 & n1459;
  assign n1615 = ~n1613 & ~n1614;
  assign n1616 = ~n37639 & ~n1612;
  assign n1617 = ~n1611 & ~n37667;
  assign n1618 = n691 & n1465;
  assign n1619 = pi74  & n37503;
  assign n1620 = pi76  & n704;
  assign n1621 = pi75  & n706;
  assign n1622 = ~n1620 & ~n1621;
  assign n1623 = ~n1619 & ~n1621;
  assign n1624 = ~n1620 & n1623;
  assign n1625 = ~n1619 & n1622;
  assign n1626 = ~n1618 & n37668;
  assign n1627 = pi38  & ~n1626;
  assign n1628 = pi38  & ~n1627;
  assign n1629 = pi38  & n1626;
  assign n1630 = ~n1626 & ~n1627;
  assign n1631 = ~pi38  & ~n1626;
  assign n1632 = ~n37669 & ~n37670;
  assign n1633 = n1449 & ~n1451;
  assign n1634 = ~n1452 & ~n1633;
  assign n1635 = ~n1632 & n1634;
  assign n1636 = n691 & n720;
  assign n1637 = pi73  & n37503;
  assign n1638 = pi75  & n704;
  assign n1639 = pi74  & n706;
  assign n1640 = ~n1638 & ~n1639;
  assign n1641 = ~n1637 & ~n1639;
  assign n1642 = ~n1638 & n1641;
  assign n1643 = ~n1637 & n1640;
  assign n1644 = ~n1636 & n37671;
  assign n1645 = pi38  & ~n1644;
  assign n1646 = pi38  & ~n1645;
  assign n1647 = pi38  & n1644;
  assign n1648 = ~n1644 & ~n1645;
  assign n1649 = ~pi38  & ~n1644;
  assign n1650 = ~n37672 & ~n37673;
  assign n1651 = n1440 & n37638;
  assign n1652 = ~n1440 & ~n1448;
  assign n1653 = ~n1440 & n37638;
  assign n1654 = ~n37638 & ~n1448;
  assign n1655 = n1440 & ~n37638;
  assign n1656 = ~n37674 & ~n37675;
  assign n1657 = ~n1448 & ~n1651;
  assign n1658 = ~n1650 & ~n37676;
  assign n1659 = n1431 & n37635;
  assign n1660 = ~n1439 & ~n1659;
  assign n1661 = n691 & n1218;
  assign n1662 = pi72  & n37503;
  assign n1663 = pi74  & n704;
  assign n1664 = pi73  & n706;
  assign n1665 = ~n1663 & ~n1664;
  assign n1666 = ~n1662 & ~n1664;
  assign n1667 = ~n1663 & n1666;
  assign n1668 = ~n1662 & n1665;
  assign n1669 = ~n1661 & n37677;
  assign n1670 = pi38  & ~n1669;
  assign n1671 = pi38  & ~n1670;
  assign n1672 = pi38  & n1669;
  assign n1673 = ~n1669 & ~n1670;
  assign n1674 = ~pi38  & ~n1669;
  assign n1675 = ~n37678 & ~n37679;
  assign n1676 = n1660 & ~n1675;
  assign n1677 = n1422 & n37632;
  assign n1678 = ~n1430 & ~n1677;
  assign n1679 = n691 & n1238;
  assign n1680 = pi71  & n37503;
  assign n1681 = pi73  & n704;
  assign n1682 = pi72  & n706;
  assign n1683 = ~n1681 & ~n1682;
  assign n1684 = ~n1680 & ~n1682;
  assign n1685 = ~n1681 & n1684;
  assign n1686 = ~n1680 & n1683;
  assign n1687 = ~n1679 & n37680;
  assign n1688 = pi38  & ~n1687;
  assign n1689 = pi38  & ~n1688;
  assign n1690 = pi38  & n1687;
  assign n1691 = ~n1687 & ~n1688;
  assign n1692 = ~pi38  & ~n1687;
  assign n1693 = ~n37681 & ~n37682;
  assign n1694 = n1678 & ~n1693;
  assign n1695 = n691 & n1124;
  assign n1696 = pi70  & n37503;
  assign n1697 = pi72  & n704;
  assign n1698 = pi71  & n706;
  assign n1699 = ~n1697 & ~n1698;
  assign n1700 = ~n1696 & ~n1698;
  assign n1701 = ~n1697 & n1700;
  assign n1702 = ~n1696 & n1699;
  assign n1703 = ~n1695 & n37683;
  assign n1704 = pi38  & ~n1703;
  assign n1705 = pi38  & ~n1704;
  assign n1706 = pi38  & n1703;
  assign n1707 = ~n1703 & ~n1704;
  assign n1708 = ~pi38  & ~n1703;
  assign n1709 = ~n37684 & ~n37685;
  assign n1710 = n1413 & n37629;
  assign n1711 = ~n1421 & ~n1710;
  assign n1712 = ~n1709 & n1711;
  assign n1713 = n1409 & ~n1411;
  assign n1714 = ~n1412 & ~n1713;
  assign n1715 = n691 & n927;
  assign n1716 = pi69  & n37503;
  assign n1717 = pi71  & n704;
  assign n1718 = pi70  & n706;
  assign n1719 = ~n1717 & ~n1718;
  assign n1720 = ~n1716 & ~n1718;
  assign n1721 = ~n1717 & n1720;
  assign n1722 = ~n1716 & n1719;
  assign n1723 = ~n1715 & n37686;
  assign n1724 = pi38  & ~n1723;
  assign n1725 = pi38  & ~n1724;
  assign n1726 = pi38  & n1723;
  assign n1727 = ~n1723 & ~n1724;
  assign n1728 = ~pi38  & ~n1723;
  assign n1729 = ~n37687 & ~n37688;
  assign n1730 = n1714 & ~n1729;
  assign n1731 = n1402 & n37626;
  assign n1732 = ~n1408 & ~n1731;
  assign n1733 = n691 & n972;
  assign n1734 = pi68  & n37503;
  assign n1735 = pi70  & n704;
  assign n1736 = pi69  & n706;
  assign n1737 = ~n1735 & ~n1736;
  assign n1738 = ~n1734 & ~n1736;
  assign n1739 = ~n1735 & n1738;
  assign n1740 = ~n1734 & n1737;
  assign n1741 = ~n1733 & n37689;
  assign n1742 = pi38  & ~n1741;
  assign n1743 = pi38  & ~n1742;
  assign n1744 = pi38  & n1741;
  assign n1745 = ~n1741 & ~n1742;
  assign n1746 = ~pi38  & ~n1741;
  assign n1747 = ~n37690 & ~n37691;
  assign n1748 = n1732 & ~n1747;
  assign n1749 = n691 & n990;
  assign n1750 = pi67  & n37503;
  assign n1751 = pi69  & n704;
  assign n1752 = pi68  & n706;
  assign n1753 = ~n1751 & ~n1752;
  assign n1754 = ~n1750 & ~n1752;
  assign n1755 = ~n1751 & n1754;
  assign n1756 = ~n1750 & n1753;
  assign n1757 = ~n1749 & n37692;
  assign n1758 = pi38  & ~n1757;
  assign n1759 = pi38  & ~n1758;
  assign n1760 = pi38  & n1757;
  assign n1761 = ~n1757 & ~n1758;
  assign n1762 = ~pi38  & ~n1757;
  assign n1763 = ~n37693 & ~n37694;
  assign n1764 = pi41  & ~n37618;
  assign n1765 = n37621 & ~n1764;
  assign n1766 = ~n37621 & n1764;
  assign n1767 = ~n37618 & n1384;
  assign n1768 = ~n37622 & ~n1767;
  assign n1769 = ~n1765 & ~n1766;
  assign n1770 = ~n1763 & n37695;
  assign n1771 = n691 & n871;
  assign n1772 = pi66  & n37503;
  assign n1773 = pi68  & n704;
  assign n1774 = pi67  & n706;
  assign n1775 = ~n1773 & ~n1774;
  assign n1776 = ~n1772 & ~n1774;
  assign n1777 = ~n1773 & n1776;
  assign n1778 = ~n1772 & n1775;
  assign n1779 = ~n1771 & n37696;
  assign n1780 = pi38  & ~n1779;
  assign n1781 = pi38  & ~n1780;
  assign n1782 = pi38  & n1779;
  assign n1783 = ~n1779 & ~n1780;
  assign n1784 = ~pi38  & ~n1779;
  assign n1785 = ~n37697 & ~n37698;
  assign n1786 = pi41  & n1358;
  assign n1787 = ~n1357 & n1786;
  assign n1788 = n1357 & ~n1786;
  assign n1789 = ~n1359 & n1363;
  assign n1790 = ~n37618 & ~n1789;
  assign n1791 = ~n1787 & ~n1788;
  assign n1792 = ~n1785 & n37699;
  assign n1793 = n691 & n37515;
  assign n1794 = pi65  & n704;
  assign n1795 = pi64  & n706;
  assign n1796 = ~n1794 & ~n1795;
  assign n1797 = ~n1793 & n1796;
  assign n1798 = pi64  & n37500;
  assign n1799 = pi38  & ~n1798;
  assign n1800 = pi38  & ~n1797;
  assign n1801 = pi38  & ~n1800;
  assign n1802 = ~n1797 & ~n1800;
  assign n1803 = ~n1801 & ~n1802;
  assign n1804 = n1799 & ~n1803;
  assign n1805 = n1797 & n1799;
  assign n1806 = pi64  & n37503;
  assign n1807 = pi65  & n706;
  assign n1808 = n691 & ~n37521;
  assign n1809 = pi66  & n704;
  assign n1810 = ~n1808 & ~n1809;
  assign n1811 = ~n1807 & ~n1808;
  assign n1812 = ~n1809 & n1811;
  assign n1813 = ~n1807 & ~n1809;
  assign n1814 = ~n1808 & n1813;
  assign n1815 = ~n1807 & n1810;
  assign n1816 = ~n1806 & ~n1807;
  assign n1817 = ~n1809 & n1816;
  assign n1818 = ~n1806 & n1813;
  assign n1819 = ~n1808 & n37702;
  assign n1820 = ~n1806 & n37701;
  assign n1821 = pi38  & ~n37703;
  assign n1822 = pi38  & ~n1821;
  assign n1823 = ~n37703 & ~n1821;
  assign n1824 = ~n1822 & ~n1823;
  assign n1825 = n37700 & ~n1824;
  assign n1826 = n37700 & n37703;
  assign n1827 = n1358 & n37704;
  assign n1828 = n691 & n847;
  assign n1829 = pi65  & n37503;
  assign n1830 = pi67  & n704;
  assign n1831 = pi66  & n706;
  assign n1832 = ~n1830 & ~n1831;
  assign n1833 = ~n1829 & ~n1831;
  assign n1834 = ~n1830 & n1833;
  assign n1835 = ~n1829 & n1832;
  assign n1836 = ~n1828 & n37705;
  assign n1837 = pi38  & ~n1836;
  assign n1838 = pi38  & ~n1837;
  assign n1839 = pi38  & n1836;
  assign n1840 = ~n1836 & ~n1837;
  assign n1841 = ~pi38  & ~n1836;
  assign n1842 = ~n37706 & ~n37707;
  assign n1843 = ~n1358 & ~n37704;
  assign n1844 = n1358 & ~n37704;
  assign n1845 = ~n1358 & n37704;
  assign n1846 = ~n1844 & ~n1845;
  assign n1847 = ~n1827 & ~n1843;
  assign n1848 = ~n1842 & ~n37708;
  assign n1849 = ~n1827 & ~n1848;
  assign n1850 = n1785 & ~n37699;
  assign n1851 = ~n1792 & ~n1850;
  assign n1852 = ~n1849 & n1851;
  assign n1853 = ~n1792 & ~n1852;
  assign n1854 = n1763 & ~n37695;
  assign n1855 = n37695 & ~n1770;
  assign n1856 = n1763 & n37695;
  assign n1857 = ~n1763 & ~n1770;
  assign n1858 = ~n1763 & ~n37695;
  assign n1859 = ~n37709 & ~n37710;
  assign n1860 = ~n1770 & ~n1854;
  assign n1861 = ~n1853 & ~n37711;
  assign n1862 = ~n1770 & ~n1861;
  assign n1863 = ~n1732 & n1747;
  assign n1864 = n1732 & ~n1748;
  assign n1865 = n1732 & n1747;
  assign n1866 = ~n1747 & ~n1748;
  assign n1867 = ~n1732 & ~n1747;
  assign n1868 = ~n37712 & ~n37713;
  assign n1869 = ~n1748 & ~n1863;
  assign n1870 = ~n1862 & ~n37714;
  assign n1871 = ~n1748 & ~n1870;
  assign n1872 = ~n1714 & n1729;
  assign n1873 = n1714 & ~n1730;
  assign n1874 = n1714 & n1729;
  assign n1875 = ~n1729 & ~n1730;
  assign n1876 = ~n1714 & ~n1729;
  assign n1877 = ~n37715 & ~n37716;
  assign n1878 = ~n1730 & ~n1872;
  assign n1879 = ~n1871 & ~n37717;
  assign n1880 = ~n1730 & ~n1879;
  assign n1881 = n1709 & ~n1711;
  assign n1882 = ~n1709 & ~n1712;
  assign n1883 = ~n1709 & ~n1711;
  assign n1884 = n1711 & ~n1712;
  assign n1885 = n1709 & n1711;
  assign n1886 = ~n37718 & ~n37719;
  assign n1887 = ~n1712 & ~n1881;
  assign n1888 = ~n1880 & ~n37720;
  assign n1889 = ~n1712 & ~n1888;
  assign n1890 = ~n1678 & n1693;
  assign n1891 = ~n1694 & ~n1890;
  assign n1892 = ~n1889 & n1891;
  assign n1893 = ~n1694 & ~n1892;
  assign n1894 = ~n1660 & n1675;
  assign n1895 = ~n1676 & ~n1894;
  assign n1896 = ~n1893 & ~n1894;
  assign n1897 = ~n1676 & n1896;
  assign n1898 = ~n1893 & n1895;
  assign n1899 = ~n1676 & ~n37721;
  assign n1900 = n1650 & n37676;
  assign n1901 = ~n1658 & ~n1900;
  assign n1902 = ~n1899 & n1901;
  assign n1903 = ~n1658 & ~n1902;
  assign n1904 = n1632 & ~n1634;
  assign n1905 = ~n1632 & ~n1635;
  assign n1906 = ~n1632 & ~n1634;
  assign n1907 = n1634 & ~n1635;
  assign n1908 = n1632 & n1634;
  assign n1909 = ~n37722 & ~n37723;
  assign n1910 = ~n1635 & ~n1904;
  assign n1911 = ~n1903 & ~n37724;
  assign n1912 = ~n1635 & ~n1911;
  assign n1913 = n1611 & n37667;
  assign n1914 = ~n1617 & ~n1913;
  assign n1915 = ~n1912 & n1914;
  assign n1916 = ~n1617 & ~n1915;
  assign n1917 = ~n1576 & n1593;
  assign n1918 = n1576 & ~n1594;
  assign n1919 = n1576 & n1593;
  assign n1920 = ~n1593 & ~n1594;
  assign n1921 = ~n1576 & ~n1593;
  assign n1922 = ~n37725 & ~n37726;
  assign n1923 = ~n1594 & ~n1917;
  assign n1924 = ~n1916 & ~n37727;
  assign n1925 = ~n1594 & ~n1924;
  assign n1926 = n718 & ~n1573;
  assign n1927 = ~n1574 & ~n1926;
  assign n1928 = ~n1925 & n1927;
  assign n1929 = ~n1574 & ~n1928;
  assign n1930 = ~n1561 & ~n1569;
  assign n1931 = n733 & n1596;
  assign n1932 = pi75  & n37510;
  assign n1933 = pi77  & n746;
  assign n1934 = pi76  & n748;
  assign n1935 = ~n1933 & ~n1934;
  assign n1936 = ~n1932 & ~n1934;
  assign n1937 = ~n1933 & n1936;
  assign n1938 = ~n1932 & n1935;
  assign n1939 = ~n1931 & n37728;
  assign n1940 = pi41  & ~n1939;
  assign n1941 = pi41  & ~n1940;
  assign n1942 = pi41  & n1939;
  assign n1943 = ~n1939 & ~n1940;
  assign n1944 = ~pi41  & ~n1939;
  assign n1945 = ~n37729 & ~n37730;
  assign n1946 = ~n1556 & ~n1558;
  assign n1947 = ~n1529 & ~n1538;
  assign n1948 = ~n1505 & ~n1511;
  assign n1949 = n871 & n894;
  assign n1950 = pi66  & n37580;
  assign n1951 = pi68  & n896;
  assign n1952 = pi67  & n904;
  assign n1953 = ~n1951 & ~n1952;
  assign n1954 = ~n1950 & ~n1952;
  assign n1955 = ~n1951 & n1954;
  assign n1956 = ~n1950 & n1953;
  assign n1957 = ~n1949 & n37731;
  assign n1958 = pi50  & ~n1957;
  assign n1959 = pi50  & ~n1958;
  assign n1960 = pi50  & n1957;
  assign n1961 = ~n1957 & ~n1958;
  assign n1962 = ~pi50  & ~n1957;
  assign n1963 = ~n37732 & ~n37733;
  assign n1964 = pi53  & n1504;
  assign n1965 = pi52  & ~pi53 ;
  assign n1966 = ~pi52  & pi53 ;
  assign n1967 = ~pi52  & ~pi53 ;
  assign n1968 = pi52  & pi53 ;
  assign n1969 = ~n1967 & ~n1968;
  assign n1970 = ~n1965 & ~n1966;
  assign n1971 = n37646 & n37734;
  assign n1972 = n37515 & n1971;
  assign n1973 = n37646 & ~n37734;
  assign n1974 = pi65  & n1973;
  assign n1975 = pi51  & ~pi52 ;
  assign n1976 = ~pi51  & pi52 ;
  assign n1977 = ~pi51  & ~pi52 ;
  assign n1978 = pi51  & pi52 ;
  assign n1979 = ~n1977 & ~n1978;
  assign n1980 = ~n1975 & ~n1976;
  assign n1981 = ~n37646 & n37735;
  assign n1982 = pi64  & n1981;
  assign n1983 = ~n1974 & ~n1982;
  assign n1984 = ~n1972 & n1983;
  assign n1985 = n1964 & ~n1984;
  assign n1986 = ~n1964 & n1984;
  assign n1987 = pi53  & ~n1504;
  assign n1988 = pi53  & ~n1984;
  assign n1989 = pi53  & ~n1988;
  assign n1990 = ~n1984 & ~n1988;
  assign n1991 = ~n1989 & ~n1990;
  assign n1992 = n1987 & ~n1991;
  assign n1993 = n1984 & n1987;
  assign n1994 = ~n1987 & n1991;
  assign n1995 = ~n37736 & ~n1994;
  assign n1996 = ~n1985 & ~n1986;
  assign n1997 = n1963 & ~n37737;
  assign n1998 = ~n1963 & n37737;
  assign n1999 = ~n1997 & ~n1998;
  assign n2000 = ~n1948 & n1999;
  assign n2001 = n1948 & ~n1999;
  assign n2002 = ~n2000 & ~n2001;
  assign n2003 = n785 & n927;
  assign n2004 = pi69  & n37520;
  assign n2005 = pi71  & n787;
  assign n2006 = pi70  & n795;
  assign n2007 = ~n2005 & ~n2006;
  assign n2008 = ~n2004 & ~n2006;
  assign n2009 = ~n2005 & n2008;
  assign n2010 = ~n2004 & n2007;
  assign n2011 = ~n2003 & n37738;
  assign n2012 = pi47  & ~n2011;
  assign n2013 = pi47  & ~n2012;
  assign n2014 = pi47  & n2011;
  assign n2015 = ~n2011 & ~n2012;
  assign n2016 = ~pi47  & ~n2011;
  assign n2017 = ~n37739 & ~n37740;
  assign n2018 = n2002 & ~n2017;
  assign n2019 = ~n2002 & n2017;
  assign n2020 = n2002 & ~n2018;
  assign n2021 = n2002 & n2017;
  assign n2022 = ~n2017 & ~n2018;
  assign n2023 = ~n2002 & ~n2017;
  assign n2024 = ~n37741 & ~n37742;
  assign n2025 = ~n2018 & ~n2019;
  assign n2026 = n1947 & n37743;
  assign n2027 = ~n1947 & ~n37743;
  assign n2028 = ~n2026 & ~n2027;
  assign n2029 = n940 & n1218;
  assign n2030 = pi72  & n37541;
  assign n2031 = pi74  & n953;
  assign n2032 = pi73  & n955;
  assign n2033 = ~n2031 & ~n2032;
  assign n2034 = ~n2030 & ~n2032;
  assign n2035 = ~n2031 & n2034;
  assign n2036 = ~n2030 & n2033;
  assign n2037 = ~n2029 & n37744;
  assign n2038 = pi44  & ~n2037;
  assign n2039 = pi44  & ~n2038;
  assign n2040 = pi44  & n2037;
  assign n2041 = ~n2037 & ~n2038;
  assign n2042 = ~pi44  & ~n2037;
  assign n2043 = ~n37745 & ~n37746;
  assign n2044 = n2028 & ~n2043;
  assign n2045 = ~n2028 & n2043;
  assign n2046 = ~n2044 & ~n2045;
  assign n2047 = ~n1946 & ~n2045;
  assign n2048 = ~n2044 & n2047;
  assign n2049 = ~n1946 & n2046;
  assign n2050 = n1946 & ~n2046;
  assign n2051 = ~n1946 & ~n37747;
  assign n2052 = ~n2044 & ~n37747;
  assign n2053 = ~n2045 & n2052;
  assign n2054 = ~n2051 & ~n2053;
  assign n2055 = ~n37747 & ~n2050;
  assign n2056 = n1945 & n37748;
  assign n2057 = ~n1945 & ~n37748;
  assign n2058 = ~n2056 & ~n2057;
  assign n2059 = ~n1930 & n2058;
  assign n2060 = n1930 & ~n2058;
  assign n2061 = ~n2059 & ~n2060;
  assign n2062 = n377 & ~n379;
  assign n2063 = ~n380 & ~n2062;
  assign n2064 = n691 & n2063;
  assign n2065 = pi78  & n37503;
  assign n2066 = pi80  & n704;
  assign n2067 = pi79  & n706;
  assign n2068 = ~n2066 & ~n2067;
  assign n2069 = ~n2065 & ~n2067;
  assign n2070 = ~n2066 & n2069;
  assign n2071 = ~n2065 & n2068;
  assign n2072 = ~n2064 & n37749;
  assign n2073 = pi38  & ~n2072;
  assign n2074 = pi38  & ~n2073;
  assign n2075 = pi38  & n2072;
  assign n2076 = ~n2072 & ~n2073;
  assign n2077 = ~pi38  & ~n2072;
  assign n2078 = ~n37750 & ~n37751;
  assign n2079 = n2061 & ~n2078;
  assign n2080 = ~n2061 & n2078;
  assign n2081 = n2061 & ~n2079;
  assign n2082 = n2061 & n2078;
  assign n2083 = ~n2078 & ~n2079;
  assign n2084 = ~n2061 & ~n2078;
  assign n2085 = ~n37752 & ~n37753;
  assign n2086 = ~n2079 & ~n2080;
  assign n2087 = n1929 & n37754;
  assign n2088 = ~n1929 & ~n37754;
  assign n2089 = ~n2087 & ~n2088;
  assign n2090 = n389 & ~n391;
  assign n2091 = ~n392 & ~n2090;
  assign n2092 = pi32  & ~pi33 ;
  assign n2093 = ~pi32  & pi33 ;
  assign n2094 = ~pi32  & ~pi33 ;
  assign n2095 = pi32  & pi33 ;
  assign n2096 = ~n2094 & ~n2095;
  assign n2097 = ~n2092 & ~n2093;
  assign n2098 = pi34  & ~pi35 ;
  assign n2099 = ~pi34  & pi35 ;
  assign n2100 = ~pi34  & ~pi35 ;
  assign n2101 = pi34  & pi35 ;
  assign n2102 = ~n2100 & ~n2101;
  assign n2103 = ~n2098 & ~n2099;
  assign n2104 = n37755 & n37756;
  assign n2105 = n2091 & n2104;
  assign n2106 = pi33  & ~pi34 ;
  assign n2107 = ~pi33  & pi34 ;
  assign n2108 = ~pi33  & ~pi34 ;
  assign n2109 = pi33  & pi34 ;
  assign n2110 = ~n2108 & ~n2109;
  assign n2111 = ~n2106 & ~n2107;
  assign n2112 = ~n37755 & n37756;
  assign n2113 = ~n37755 & ~n37757;
  assign n2114 = n37756 & n2113;
  assign n2115 = ~n37757 & n2112;
  assign n2116 = pi81  & n37758;
  assign n2117 = n37755 & ~n37756;
  assign n2118 = pi83  & n2117;
  assign n2119 = ~n37755 & n37757;
  assign n2120 = pi82  & n2119;
  assign n2121 = ~n2118 & ~n2120;
  assign n2122 = ~n2116 & ~n2120;
  assign n2123 = ~n2118 & n2122;
  assign n2124 = ~n2116 & n2121;
  assign n2125 = ~n2105 & n37759;
  assign n2126 = pi35  & ~n2125;
  assign n2127 = pi35  & ~n2126;
  assign n2128 = pi35  & n2125;
  assign n2129 = ~n2125 & ~n2126;
  assign n2130 = ~pi35  & ~n2125;
  assign n2131 = ~n37760 & ~n37761;
  assign n2132 = n2089 & ~n2131;
  assign n2133 = n385 & ~n387;
  assign n2134 = ~n388 & ~n2133;
  assign n2135 = n2104 & n2134;
  assign n2136 = pi80  & n37758;
  assign n2137 = pi82  & n2117;
  assign n2138 = pi81  & n2119;
  assign n2139 = ~n2137 & ~n2138;
  assign n2140 = ~n2136 & ~n2138;
  assign n2141 = ~n2137 & n2140;
  assign n2142 = ~n2136 & n2139;
  assign n2143 = ~n2135 & n37762;
  assign n2144 = pi35  & ~n2143;
  assign n2145 = pi35  & ~n2144;
  assign n2146 = pi35  & n2143;
  assign n2147 = ~n2143 & ~n2144;
  assign n2148 = ~pi35  & ~n2143;
  assign n2149 = ~n37763 & ~n37764;
  assign n2150 = n1925 & ~n1927;
  assign n2151 = ~n1928 & ~n2150;
  assign n2152 = ~n2149 & n2151;
  assign n2153 = n381 & ~n383;
  assign n2154 = ~n384 & ~n2153;
  assign n2155 = n2104 & n2154;
  assign n2156 = pi79  & n37758;
  assign n2157 = pi81  & n2117;
  assign n2158 = pi80  & n2119;
  assign n2159 = ~n2157 & ~n2158;
  assign n2160 = ~n2156 & ~n2158;
  assign n2161 = ~n2157 & n2160;
  assign n2162 = ~n2156 & n2159;
  assign n2163 = ~n2155 & n37765;
  assign n2164 = pi35  & ~n2163;
  assign n2165 = pi35  & ~n2164;
  assign n2166 = pi35  & n2163;
  assign n2167 = ~n2163 & ~n2164;
  assign n2168 = ~pi35  & ~n2163;
  assign n2169 = ~n37766 & ~n37767;
  assign n2170 = n1916 & n37727;
  assign n2171 = ~n1924 & ~n2170;
  assign n2172 = ~n2169 & n2171;
  assign n2173 = n1912 & ~n1914;
  assign n2174 = ~n1915 & ~n2173;
  assign n2175 = n2063 & n2104;
  assign n2176 = pi78  & n37758;
  assign n2177 = pi80  & n2117;
  assign n2178 = pi79  & n2119;
  assign n2179 = ~n2177 & ~n2178;
  assign n2180 = ~n2176 & ~n2178;
  assign n2181 = ~n2177 & n2180;
  assign n2182 = ~n2176 & n2179;
  assign n2183 = ~n2175 & n37768;
  assign n2184 = pi35  & ~n2183;
  assign n2185 = pi35  & ~n2184;
  assign n2186 = pi35  & n2183;
  assign n2187 = ~n2183 & ~n2184;
  assign n2188 = ~pi35  & ~n2183;
  assign n2189 = ~n37769 & ~n37770;
  assign n2190 = n2174 & ~n2189;
  assign n2191 = n678 & n2104;
  assign n2192 = pi77  & n37758;
  assign n2193 = pi79  & n2117;
  assign n2194 = pi78  & n2119;
  assign n2195 = ~n2193 & ~n2194;
  assign n2196 = ~n2192 & ~n2194;
  assign n2197 = ~n2193 & n2196;
  assign n2198 = ~n2192 & n2195;
  assign n2199 = ~n2191 & n37771;
  assign n2200 = pi35  & ~n2199;
  assign n2201 = pi35  & ~n2200;
  assign n2202 = pi35  & n2199;
  assign n2203 = ~n2199 & ~n2200;
  assign n2204 = ~pi35  & ~n2199;
  assign n2205 = ~n37772 & ~n37773;
  assign n2206 = n1903 & ~n37723;
  assign n2207 = ~n37722 & n2206;
  assign n2208 = n1903 & n37724;
  assign n2209 = ~n1911 & ~n37774;
  assign n2210 = ~n2205 & n2209;
  assign n2211 = n1899 & ~n1901;
  assign n2212 = ~n1902 & ~n2211;
  assign n2213 = n1578 & n2104;
  assign n2214 = pi76  & n37758;
  assign n2215 = pi78  & n2117;
  assign n2216 = pi77  & n2119;
  assign n2217 = ~n2215 & ~n2216;
  assign n2218 = ~n2214 & ~n2216;
  assign n2219 = ~n2215 & n2218;
  assign n2220 = ~n2214 & n2217;
  assign n2221 = ~n2213 & n37775;
  assign n2222 = pi35  & ~n2221;
  assign n2223 = pi35  & ~n2222;
  assign n2224 = pi35  & n2221;
  assign n2225 = ~n2221 & ~n2222;
  assign n2226 = ~pi35  & ~n2221;
  assign n2227 = ~n37776 & ~n37777;
  assign n2228 = n2212 & ~n2227;
  assign n2229 = n1596 & n2104;
  assign n2230 = pi75  & n37758;
  assign n2231 = pi77  & n2117;
  assign n2232 = pi76  & n2119;
  assign n2233 = ~n2231 & ~n2232;
  assign n2234 = ~n2230 & ~n2232;
  assign n2235 = ~n2231 & n2234;
  assign n2236 = ~n2230 & n2233;
  assign n2237 = ~n2229 & n37778;
  assign n2238 = pi35  & ~n2237;
  assign n2239 = pi35  & ~n2238;
  assign n2240 = pi35  & n2237;
  assign n2241 = ~n2237 & ~n2238;
  assign n2242 = ~pi35  & ~n2237;
  assign n2243 = ~n37779 & ~n37780;
  assign n2244 = n1893 & ~n1895;
  assign n2245 = ~n1893 & ~n37721;
  assign n2246 = ~n1894 & n1899;
  assign n2247 = ~n2245 & ~n2246;
  assign n2248 = ~n37721 & ~n2244;
  assign n2249 = ~n2243 & ~n37781;
  assign n2250 = n1465 & n2104;
  assign n2251 = pi74  & n37758;
  assign n2252 = pi76  & n2117;
  assign n2253 = pi75  & n2119;
  assign n2254 = ~n2252 & ~n2253;
  assign n2255 = ~n2251 & ~n2253;
  assign n2256 = ~n2252 & n2255;
  assign n2257 = ~n2251 & n2254;
  assign n2258 = ~n2250 & n37782;
  assign n2259 = pi35  & ~n2258;
  assign n2260 = pi35  & ~n2259;
  assign n2261 = pi35  & n2258;
  assign n2262 = ~n2258 & ~n2259;
  assign n2263 = ~pi35  & ~n2258;
  assign n2264 = ~n37783 & ~n37784;
  assign n2265 = n1889 & ~n1891;
  assign n2266 = ~n1892 & ~n2265;
  assign n2267 = ~n2264 & n2266;
  assign n2268 = n720 & n2104;
  assign n2269 = pi73  & n37758;
  assign n2270 = pi75  & n2117;
  assign n2271 = pi74  & n2119;
  assign n2272 = ~n2270 & ~n2271;
  assign n2273 = ~n2269 & ~n2271;
  assign n2274 = ~n2270 & n2273;
  assign n2275 = ~n2269 & n2272;
  assign n2276 = ~n2268 & n37785;
  assign n2277 = pi35  & ~n2276;
  assign n2278 = pi35  & ~n2277;
  assign n2279 = pi35  & n2276;
  assign n2280 = ~n2276 & ~n2277;
  assign n2281 = ~pi35  & ~n2276;
  assign n2282 = ~n37786 & ~n37787;
  assign n2283 = n1880 & n37720;
  assign n2284 = ~n1880 & ~n1888;
  assign n2285 = ~n1880 & n37720;
  assign n2286 = ~n37720 & ~n1888;
  assign n2287 = n1880 & ~n37720;
  assign n2288 = ~n37788 & ~n37789;
  assign n2289 = ~n1888 & ~n2283;
  assign n2290 = ~n2282 & ~n37790;
  assign n2291 = n1871 & n37717;
  assign n2292 = ~n1879 & ~n2291;
  assign n2293 = n1218 & n2104;
  assign n2294 = pi72  & n37758;
  assign n2295 = pi74  & n2117;
  assign n2296 = pi73  & n2119;
  assign n2297 = ~n2295 & ~n2296;
  assign n2298 = ~n2294 & ~n2296;
  assign n2299 = ~n2295 & n2298;
  assign n2300 = ~n2294 & n2297;
  assign n2301 = ~n2293 & n37791;
  assign n2302 = pi35  & ~n2301;
  assign n2303 = pi35  & ~n2302;
  assign n2304 = pi35  & n2301;
  assign n2305 = ~n2301 & ~n2302;
  assign n2306 = ~pi35  & ~n2301;
  assign n2307 = ~n37792 & ~n37793;
  assign n2308 = n2292 & ~n2307;
  assign n2309 = n1862 & n37714;
  assign n2310 = ~n1870 & ~n2309;
  assign n2311 = n1238 & n2104;
  assign n2312 = pi71  & n37758;
  assign n2313 = pi73  & n2117;
  assign n2314 = pi72  & n2119;
  assign n2315 = ~n2313 & ~n2314;
  assign n2316 = ~n2312 & ~n2314;
  assign n2317 = ~n2313 & n2316;
  assign n2318 = ~n2312 & n2315;
  assign n2319 = ~n2311 & n37794;
  assign n2320 = pi35  & ~n2319;
  assign n2321 = pi35  & ~n2320;
  assign n2322 = pi35  & n2319;
  assign n2323 = ~n2319 & ~n2320;
  assign n2324 = ~pi35  & ~n2319;
  assign n2325 = ~n37795 & ~n37796;
  assign n2326 = n2310 & ~n2325;
  assign n2327 = n1124 & n2104;
  assign n2328 = pi70  & n37758;
  assign n2329 = pi72  & n2117;
  assign n2330 = pi71  & n2119;
  assign n2331 = ~n2329 & ~n2330;
  assign n2332 = ~n2328 & ~n2330;
  assign n2333 = ~n2329 & n2332;
  assign n2334 = ~n2328 & n2331;
  assign n2335 = ~n2327 & n37797;
  assign n2336 = pi35  & ~n2335;
  assign n2337 = pi35  & ~n2336;
  assign n2338 = pi35  & n2335;
  assign n2339 = ~n2335 & ~n2336;
  assign n2340 = ~pi35  & ~n2335;
  assign n2341 = ~n37798 & ~n37799;
  assign n2342 = n1853 & n37711;
  assign n2343 = ~n1861 & ~n2342;
  assign n2344 = ~n2341 & n2343;
  assign n2345 = n1849 & ~n1851;
  assign n2346 = ~n1852 & ~n2345;
  assign n2347 = n927 & n2104;
  assign n2348 = pi69  & n37758;
  assign n2349 = pi71  & n2117;
  assign n2350 = pi70  & n2119;
  assign n2351 = ~n2349 & ~n2350;
  assign n2352 = ~n2348 & ~n2350;
  assign n2353 = ~n2349 & n2352;
  assign n2354 = ~n2348 & n2351;
  assign n2355 = ~n2347 & n37800;
  assign n2356 = pi35  & ~n2355;
  assign n2357 = pi35  & ~n2356;
  assign n2358 = pi35  & n2355;
  assign n2359 = ~n2355 & ~n2356;
  assign n2360 = ~pi35  & ~n2355;
  assign n2361 = ~n37801 & ~n37802;
  assign n2362 = n2346 & ~n2361;
  assign n2363 = n1842 & n37708;
  assign n2364 = ~n1848 & ~n2363;
  assign n2365 = n972 & n2104;
  assign n2366 = pi68  & n37758;
  assign n2367 = pi70  & n2117;
  assign n2368 = pi69  & n2119;
  assign n2369 = ~n2367 & ~n2368;
  assign n2370 = ~n2366 & ~n2368;
  assign n2371 = ~n2367 & n2370;
  assign n2372 = ~n2366 & n2369;
  assign n2373 = ~n2365 & n37803;
  assign n2374 = pi35  & ~n2373;
  assign n2375 = pi35  & ~n2374;
  assign n2376 = pi35  & n2373;
  assign n2377 = ~n2373 & ~n2374;
  assign n2378 = ~pi35  & ~n2373;
  assign n2379 = ~n37804 & ~n37805;
  assign n2380 = n2364 & ~n2379;
  assign n2381 = n990 & n2104;
  assign n2382 = pi67  & n37758;
  assign n2383 = pi69  & n2117;
  assign n2384 = pi68  & n2119;
  assign n2385 = ~n2383 & ~n2384;
  assign n2386 = ~n2382 & ~n2384;
  assign n2387 = ~n2383 & n2386;
  assign n2388 = ~n2382 & n2385;
  assign n2389 = ~n2381 & n37806;
  assign n2390 = pi35  & ~n2389;
  assign n2391 = pi35  & ~n2390;
  assign n2392 = pi35  & n2389;
  assign n2393 = ~n2389 & ~n2390;
  assign n2394 = ~pi35  & ~n2389;
  assign n2395 = ~n37807 & ~n37808;
  assign n2396 = pi38  & ~n37700;
  assign n2397 = n37703 & ~n2396;
  assign n2398 = ~n37703 & n2396;
  assign n2399 = ~n37700 & n1824;
  assign n2400 = ~n37704 & ~n2399;
  assign n2401 = ~n2397 & ~n2398;
  assign n2402 = ~n2395 & n37809;
  assign n2403 = n871 & n2104;
  assign n2404 = pi66  & n37758;
  assign n2405 = pi68  & n2117;
  assign n2406 = pi67  & n2119;
  assign n2407 = ~n2405 & ~n2406;
  assign n2408 = ~n2404 & ~n2406;
  assign n2409 = ~n2405 & n2408;
  assign n2410 = ~n2404 & n2407;
  assign n2411 = ~n2403 & n37810;
  assign n2412 = pi35  & ~n2411;
  assign n2413 = pi35  & ~n2412;
  assign n2414 = pi35  & n2411;
  assign n2415 = ~n2411 & ~n2412;
  assign n2416 = ~pi35  & ~n2411;
  assign n2417 = ~n37811 & ~n37812;
  assign n2418 = pi38  & n1798;
  assign n2419 = ~n1797 & n2418;
  assign n2420 = n1797 & ~n2418;
  assign n2421 = ~n1799 & n1803;
  assign n2422 = ~n37700 & ~n2421;
  assign n2423 = ~n2419 & ~n2420;
  assign n2424 = ~n2417 & n37813;
  assign n2425 = n37515 & n2104;
  assign n2426 = pi65  & n2117;
  assign n2427 = pi64  & n2119;
  assign n2428 = ~n2426 & ~n2427;
  assign n2429 = ~n2425 & n2428;
  assign n2430 = pi64  & n37755;
  assign n2431 = pi35  & ~n2430;
  assign n2432 = pi35  & ~n2429;
  assign n2433 = pi35  & ~n2432;
  assign n2434 = ~n2429 & ~n2432;
  assign n2435 = ~n2433 & ~n2434;
  assign n2436 = n2431 & ~n2435;
  assign n2437 = n2429 & n2431;
  assign n2438 = pi64  & n37758;
  assign n2439 = pi65  & n2119;
  assign n2440 = ~n37521 & n2104;
  assign n2441 = pi66  & n2117;
  assign n2442 = ~n2440 & ~n2441;
  assign n2443 = ~n2439 & ~n2440;
  assign n2444 = ~n2441 & n2443;
  assign n2445 = ~n2439 & ~n2441;
  assign n2446 = ~n2440 & n2445;
  assign n2447 = ~n2439 & n2442;
  assign n2448 = ~n2438 & ~n2439;
  assign n2449 = ~n2441 & n2448;
  assign n2450 = ~n2438 & n2445;
  assign n2451 = ~n2440 & n37816;
  assign n2452 = ~n2438 & n37815;
  assign n2453 = pi35  & ~n37817;
  assign n2454 = pi35  & ~n2453;
  assign n2455 = ~n37817 & ~n2453;
  assign n2456 = ~n2454 & ~n2455;
  assign n2457 = n37814 & ~n2456;
  assign n2458 = n37814 & n37817;
  assign n2459 = n1798 & n37818;
  assign n2460 = n847 & n2104;
  assign n2461 = pi65  & n37758;
  assign n2462 = pi67  & n2117;
  assign n2463 = pi66  & n2119;
  assign n2464 = ~n2462 & ~n2463;
  assign n2465 = ~n2461 & ~n2463;
  assign n2466 = ~n2462 & n2465;
  assign n2467 = ~n2461 & n2464;
  assign n2468 = ~n2460 & n37819;
  assign n2469 = pi35  & ~n2468;
  assign n2470 = pi35  & ~n2469;
  assign n2471 = pi35  & n2468;
  assign n2472 = ~n2468 & ~n2469;
  assign n2473 = ~pi35  & ~n2468;
  assign n2474 = ~n37820 & ~n37821;
  assign n2475 = ~n1798 & ~n37818;
  assign n2476 = n1798 & ~n37818;
  assign n2477 = ~n1798 & n37818;
  assign n2478 = ~n2476 & ~n2477;
  assign n2479 = ~n2459 & ~n2475;
  assign n2480 = ~n2474 & ~n37822;
  assign n2481 = ~n2459 & ~n2480;
  assign n2482 = n2417 & ~n37813;
  assign n2483 = ~n2424 & ~n2482;
  assign n2484 = ~n2481 & n2483;
  assign n2485 = ~n2424 & ~n2484;
  assign n2486 = n2395 & ~n37809;
  assign n2487 = n37809 & ~n2402;
  assign n2488 = n2395 & n37809;
  assign n2489 = ~n2395 & ~n2402;
  assign n2490 = ~n2395 & ~n37809;
  assign n2491 = ~n37823 & ~n37824;
  assign n2492 = ~n2402 & ~n2486;
  assign n2493 = ~n2485 & ~n37825;
  assign n2494 = ~n2402 & ~n2493;
  assign n2495 = ~n2364 & n2379;
  assign n2496 = n2364 & ~n2380;
  assign n2497 = n2364 & n2379;
  assign n2498 = ~n2379 & ~n2380;
  assign n2499 = ~n2364 & ~n2379;
  assign n2500 = ~n37826 & ~n37827;
  assign n2501 = ~n2380 & ~n2495;
  assign n2502 = ~n2494 & ~n37828;
  assign n2503 = ~n2380 & ~n2502;
  assign n2504 = ~n2346 & n2361;
  assign n2505 = n2346 & ~n2362;
  assign n2506 = n2346 & n2361;
  assign n2507 = ~n2361 & ~n2362;
  assign n2508 = ~n2346 & ~n2361;
  assign n2509 = ~n37829 & ~n37830;
  assign n2510 = ~n2362 & ~n2504;
  assign n2511 = ~n2503 & ~n37831;
  assign n2512 = ~n2362 & ~n2511;
  assign n2513 = n2341 & ~n2343;
  assign n2514 = ~n2341 & ~n2344;
  assign n2515 = ~n2341 & ~n2343;
  assign n2516 = n2343 & ~n2344;
  assign n2517 = n2341 & n2343;
  assign n2518 = ~n37832 & ~n37833;
  assign n2519 = ~n2344 & ~n2513;
  assign n2520 = ~n2512 & ~n37834;
  assign n2521 = ~n2344 & ~n2520;
  assign n2522 = ~n2310 & n2325;
  assign n2523 = ~n2326 & ~n2522;
  assign n2524 = ~n2521 & n2523;
  assign n2525 = ~n2326 & ~n2524;
  assign n2526 = ~n2292 & n2307;
  assign n2527 = ~n2308 & ~n2526;
  assign n2528 = ~n2525 & ~n2526;
  assign n2529 = ~n2308 & n2528;
  assign n2530 = ~n2525 & n2527;
  assign n2531 = ~n2308 & ~n37835;
  assign n2532 = n2282 & n37790;
  assign n2533 = ~n2290 & ~n2532;
  assign n2534 = ~n2531 & n2533;
  assign n2535 = ~n2290 & ~n2534;
  assign n2536 = n2264 & ~n2266;
  assign n2537 = ~n2264 & ~n2267;
  assign n2538 = ~n2264 & ~n2266;
  assign n2539 = n2266 & ~n2267;
  assign n2540 = n2264 & n2266;
  assign n2541 = ~n37836 & ~n37837;
  assign n2542 = ~n2267 & ~n2536;
  assign n2543 = ~n2535 & ~n37838;
  assign n2544 = ~n2267 & ~n2543;
  assign n2545 = n2243 & n37781;
  assign n2546 = ~n2249 & ~n2545;
  assign n2547 = ~n2544 & n2546;
  assign n2548 = ~n2249 & ~n2547;
  assign n2549 = ~n2212 & n2227;
  assign n2550 = n2212 & ~n2228;
  assign n2551 = n2212 & n2227;
  assign n2552 = ~n2227 & ~n2228;
  assign n2553 = ~n2212 & ~n2227;
  assign n2554 = ~n37839 & ~n37840;
  assign n2555 = ~n2228 & ~n2549;
  assign n2556 = ~n2548 & ~n37841;
  assign n2557 = ~n2228 & ~n2556;
  assign n2558 = n2205 & ~n2209;
  assign n2559 = ~n2210 & ~n2558;
  assign n2560 = ~n2557 & n2559;
  assign n2561 = ~n2210 & ~n2560;
  assign n2562 = ~n2174 & n2189;
  assign n2563 = n2174 & ~n2190;
  assign n2564 = n2174 & n2189;
  assign n2565 = ~n2189 & ~n2190;
  assign n2566 = ~n2174 & ~n2189;
  assign n2567 = ~n37842 & ~n37843;
  assign n2568 = ~n2190 & ~n2562;
  assign n2569 = ~n2561 & ~n37844;
  assign n2570 = ~n2190 & ~n2569;
  assign n2571 = n2169 & ~n2171;
  assign n2572 = ~n2169 & ~n2172;
  assign n2573 = ~n2169 & ~n2171;
  assign n2574 = n2171 & ~n2172;
  assign n2575 = n2169 & n2171;
  assign n2576 = ~n37845 & ~n37846;
  assign n2577 = ~n2172 & ~n2571;
  assign n2578 = ~n2570 & ~n37847;
  assign n2579 = ~n2172 & ~n2578;
  assign n2580 = n2149 & ~n2151;
  assign n2581 = ~n2152 & ~n2580;
  assign n2582 = ~n2579 & n2581;
  assign n2583 = ~n2152 & ~n2582;
  assign n2584 = ~n2089 & n2131;
  assign n2585 = ~n2132 & ~n2584;
  assign n2586 = ~n2583 & ~n2584;
  assign n2587 = ~n2132 & n2586;
  assign n2588 = ~n2583 & n2585;
  assign n2589 = ~n2132 & ~n37848;
  assign n2590 = n393 & ~n395;
  assign n2591 = ~n396 & ~n2590;
  assign n2592 = n2104 & n2591;
  assign n2593 = pi82  & n37758;
  assign n2594 = pi84  & n2117;
  assign n2595 = pi83  & n2119;
  assign n2596 = ~n2594 & ~n2595;
  assign n2597 = ~n2593 & ~n2595;
  assign n2598 = ~n2594 & n2597;
  assign n2599 = ~n2593 & n2596;
  assign n2600 = ~n2592 & n37849;
  assign n2601 = pi35  & ~n2600;
  assign n2602 = pi35  & ~n2601;
  assign n2603 = pi35  & n2600;
  assign n2604 = ~n2600 & ~n2601;
  assign n2605 = ~pi35  & ~n2600;
  assign n2606 = ~n37850 & ~n37851;
  assign n2607 = ~n2079 & ~n2088;
  assign n2608 = n691 & n2154;
  assign n2609 = pi79  & n37503;
  assign n2610 = pi81  & n704;
  assign n2611 = pi80  & n706;
  assign n2612 = ~n2610 & ~n2611;
  assign n2613 = ~n2609 & ~n2611;
  assign n2614 = ~n2610 & n2613;
  assign n2615 = ~n2609 & n2612;
  assign n2616 = ~n2608 & n37852;
  assign n2617 = pi38  & ~n2616;
  assign n2618 = pi38  & ~n2617;
  assign n2619 = pi38  & n2616;
  assign n2620 = ~n2616 & ~n2617;
  assign n2621 = ~pi38  & ~n2616;
  assign n2622 = ~n37853 & ~n37854;
  assign n2623 = ~n2057 & ~n2059;
  assign n2624 = n720 & n940;
  assign n2625 = pi73  & n37541;
  assign n2626 = pi75  & n953;
  assign n2627 = pi74  & n955;
  assign n2628 = ~n2626 & ~n2627;
  assign n2629 = ~n2625 & ~n2627;
  assign n2630 = ~n2626 & n2629;
  assign n2631 = ~n2625 & n2628;
  assign n2632 = ~n2624 & n37855;
  assign n2633 = pi44  & ~n2632;
  assign n2634 = pi44  & ~n2633;
  assign n2635 = pi44  & n2632;
  assign n2636 = ~n2632 & ~n2633;
  assign n2637 = ~pi44  & ~n2632;
  assign n2638 = ~n37856 & ~n37857;
  assign n2639 = ~n2018 & ~n2027;
  assign n2640 = n785 & n1124;
  assign n2641 = pi70  & n37520;
  assign n2642 = pi72  & n787;
  assign n2643 = pi71  & n795;
  assign n2644 = ~n2642 & ~n2643;
  assign n2645 = ~n2641 & ~n2643;
  assign n2646 = ~n2642 & n2645;
  assign n2647 = ~n2641 & n2644;
  assign n2648 = ~n2640 & n37858;
  assign n2649 = pi47  & ~n2648;
  assign n2650 = pi47  & ~n2649;
  assign n2651 = pi47  & n2648;
  assign n2652 = ~n2648 & ~n2649;
  assign n2653 = ~pi47  & ~n2648;
  assign n2654 = ~n37859 & ~n37860;
  assign n2655 = ~n1998 & ~n2000;
  assign n2656 = n894 & n990;
  assign n2657 = pi67  & n37580;
  assign n2658 = pi69  & n896;
  assign n2659 = pi68  & n904;
  assign n2660 = ~n2658 & ~n2659;
  assign n2661 = ~n2657 & ~n2659;
  assign n2662 = ~n2658 & n2661;
  assign n2663 = ~n2657 & n2660;
  assign n2664 = ~n2656 & n37861;
  assign n2665 = pi50  & ~n2664;
  assign n2666 = pi50  & ~n2665;
  assign n2667 = pi50  & n2664;
  assign n2668 = ~n2664 & ~n2665;
  assign n2669 = ~pi50  & ~n2664;
  assign n2670 = ~n37862 & ~n37863;
  assign n2671 = pi53  & ~n37736;
  assign n2672 = ~n37646 & n37734;
  assign n2673 = ~n37646 & ~n37735;
  assign n2674 = n37734 & n2673;
  assign n2675 = ~n37735 & n2672;
  assign n2676 = pi64  & n37864;
  assign n2677 = pi65  & n1981;
  assign n2678 = ~n37521 & n1971;
  assign n2679 = pi66  & n1973;
  assign n2680 = ~n2678 & ~n2679;
  assign n2681 = ~n2677 & ~n2678;
  assign n2682 = ~n2679 & n2681;
  assign n2683 = ~n2677 & ~n2679;
  assign n2684 = ~n2678 & n2683;
  assign n2685 = ~n2677 & n2680;
  assign n2686 = ~n2676 & ~n2677;
  assign n2687 = ~n2679 & n2686;
  assign n2688 = ~n2676 & n2683;
  assign n2689 = ~n2678 & n37866;
  assign n2690 = ~n2676 & n37865;
  assign n2691 = ~n2671 & n37867;
  assign n2692 = n2671 & ~n37867;
  assign n2693 = pi53  & ~n37867;
  assign n2694 = pi53  & ~n2693;
  assign n2695 = ~n37867 & ~n2693;
  assign n2696 = ~n2694 & ~n2695;
  assign n2697 = n37736 & ~n2696;
  assign n2698 = n37736 & n37867;
  assign n2699 = ~n37736 & n2696;
  assign n2700 = ~n37868 & ~n2699;
  assign n2701 = ~n2691 & ~n2692;
  assign n2702 = ~n2670 & n37869;
  assign n2703 = n2670 & ~n37869;
  assign n2704 = ~n2702 & ~n2703;
  assign n2705 = ~n2655 & ~n2703;
  assign n2706 = ~n2702 & n2705;
  assign n2707 = ~n2655 & n2704;
  assign n2708 = n2655 & ~n2704;
  assign n2709 = ~n2655 & ~n37870;
  assign n2710 = ~n2702 & ~n37870;
  assign n2711 = ~n2703 & n2710;
  assign n2712 = ~n2709 & ~n2711;
  assign n2713 = ~n37870 & ~n2708;
  assign n2714 = n2654 & n37871;
  assign n2715 = ~n2654 & ~n37871;
  assign n2716 = ~n2714 & ~n2715;
  assign n2717 = ~n2639 & n2716;
  assign n2718 = n2639 & ~n2716;
  assign n2719 = ~n2717 & ~n2718;
  assign n2720 = n2638 & ~n2719;
  assign n2721 = ~n2638 & n2719;
  assign n2722 = ~n2720 & ~n2721;
  assign n2723 = ~n2052 & n2722;
  assign n2724 = n2052 & ~n2722;
  assign n2725 = ~n2723 & ~n2724;
  assign n2726 = n733 & n1578;
  assign n2727 = pi76  & n37510;
  assign n2728 = pi78  & n746;
  assign n2729 = pi77  & n748;
  assign n2730 = ~n2728 & ~n2729;
  assign n2731 = ~n2727 & ~n2729;
  assign n2732 = ~n2728 & n2731;
  assign n2733 = ~n2727 & n2730;
  assign n2734 = ~n2726 & n37872;
  assign n2735 = pi41  & ~n2734;
  assign n2736 = pi41  & ~n2735;
  assign n2737 = pi41  & n2734;
  assign n2738 = ~n2734 & ~n2735;
  assign n2739 = ~pi41  & ~n2734;
  assign n2740 = ~n37873 & ~n37874;
  assign n2741 = n2725 & ~n2740;
  assign n2742 = ~n2725 & n2740;
  assign n2743 = n2725 & ~n2741;
  assign n2744 = n2725 & n2740;
  assign n2745 = ~n2740 & ~n2741;
  assign n2746 = ~n2725 & ~n2740;
  assign n2747 = ~n37875 & ~n37876;
  assign n2748 = ~n2741 & ~n2742;
  assign n2749 = ~n2623 & ~n37877;
  assign n2750 = n2623 & n37877;
  assign n2751 = ~n2749 & ~n2750;
  assign n2752 = ~n2622 & n2751;
  assign n2753 = n2622 & ~n2751;
  assign n2754 = ~n2622 & ~n2752;
  assign n2755 = ~n2622 & ~n2751;
  assign n2756 = n2751 & ~n2752;
  assign n2757 = n2622 & n2751;
  assign n2758 = ~n37878 & ~n37879;
  assign n2759 = ~n2752 & ~n2753;
  assign n2760 = ~n2607 & ~n37880;
  assign n2761 = n2607 & n37880;
  assign n2762 = ~n2607 & ~n2760;
  assign n2763 = ~n2607 & n37880;
  assign n2764 = ~n37880 & ~n2760;
  assign n2765 = n2607 & ~n37880;
  assign n2766 = ~n37881 & ~n37882;
  assign n2767 = ~n2760 & ~n2761;
  assign n2768 = ~n2606 & ~n37883;
  assign n2769 = n2606 & n37883;
  assign n2770 = ~n37883 & ~n2768;
  assign n2771 = ~n2606 & ~n2768;
  assign n2772 = ~n2770 & ~n2771;
  assign n2773 = ~n2768 & ~n2769;
  assign n2774 = ~n2589 & ~n37884;
  assign n2775 = n2589 & n37884;
  assign n2776 = ~n2774 & ~n2775;
  assign n2777 = ~n676 & n2776;
  assign n2778 = n401 & ~n403;
  assign n2779 = ~n404 & ~n2778;
  assign n2780 = n649 & n2779;
  assign n2781 = pi84  & n37496;
  assign n2782 = pi86  & n662;
  assign n2783 = pi85  & n664;
  assign n2784 = ~n2782 & ~n2783;
  assign n2785 = ~n2781 & ~n2783;
  assign n2786 = ~n2782 & n2785;
  assign n2787 = ~n2781 & n2784;
  assign n2788 = ~n2780 & n37885;
  assign n2789 = pi32  & ~n2788;
  assign n2790 = pi32  & ~n2789;
  assign n2791 = pi32  & n2788;
  assign n2792 = ~n2788 & ~n2789;
  assign n2793 = ~pi32  & ~n2788;
  assign n2794 = ~n37886 & ~n37887;
  assign n2795 = n2583 & ~n2585;
  assign n2796 = ~n2583 & ~n37848;
  assign n2797 = ~n2584 & n2589;
  assign n2798 = ~n2796 & ~n2797;
  assign n2799 = ~n37848 & ~n2795;
  assign n2800 = ~n2794 & ~n37888;
  assign n2801 = n2579 & ~n2581;
  assign n2802 = ~n2582 & ~n2801;
  assign n2803 = n397 & ~n399;
  assign n2804 = ~n400 & ~n2803;
  assign n2805 = n649 & n2804;
  assign n2806 = pi83  & n37496;
  assign n2807 = pi85  & n662;
  assign n2808 = pi84  & n664;
  assign n2809 = ~n2807 & ~n2808;
  assign n2810 = ~n2806 & ~n2808;
  assign n2811 = ~n2807 & n2810;
  assign n2812 = ~n2806 & n2809;
  assign n2813 = ~n2805 & n37889;
  assign n2814 = pi32  & ~n2813;
  assign n2815 = pi32  & ~n2814;
  assign n2816 = pi32  & n2813;
  assign n2817 = ~n2813 & ~n2814;
  assign n2818 = ~pi32  & ~n2813;
  assign n2819 = ~n37890 & ~n37891;
  assign n2820 = n2802 & ~n2819;
  assign n2821 = n649 & n2591;
  assign n2822 = pi82  & n37496;
  assign n2823 = pi84  & n662;
  assign n2824 = pi83  & n664;
  assign n2825 = ~n2823 & ~n2824;
  assign n2826 = ~n2822 & ~n2824;
  assign n2827 = ~n2823 & n2826;
  assign n2828 = ~n2822 & n2825;
  assign n2829 = ~n2821 & n37892;
  assign n2830 = pi32  & ~n2829;
  assign n2831 = pi32  & ~n2830;
  assign n2832 = pi32  & n2829;
  assign n2833 = ~n2829 & ~n2830;
  assign n2834 = ~pi32  & ~n2829;
  assign n2835 = ~n37893 & ~n37894;
  assign n2836 = n2570 & n37847;
  assign n2837 = ~n2570 & ~n2578;
  assign n2838 = ~n2570 & n37847;
  assign n2839 = ~n37847 & ~n2578;
  assign n2840 = n2570 & ~n37847;
  assign n2841 = ~n37895 & ~n37896;
  assign n2842 = ~n2578 & ~n2836;
  assign n2843 = ~n2835 & ~n37897;
  assign n2844 = n2561 & n37844;
  assign n2845 = ~n2569 & ~n2844;
  assign n2846 = n649 & n2091;
  assign n2847 = pi81  & n37496;
  assign n2848 = pi83  & n662;
  assign n2849 = pi82  & n664;
  assign n2850 = ~n2848 & ~n2849;
  assign n2851 = ~n2847 & ~n2849;
  assign n2852 = ~n2848 & n2851;
  assign n2853 = ~n2847 & n2850;
  assign n2854 = ~n2846 & n37898;
  assign n2855 = pi32  & ~n2854;
  assign n2856 = pi32  & ~n2855;
  assign n2857 = pi32  & n2854;
  assign n2858 = ~n2854 & ~n2855;
  assign n2859 = ~pi32  & ~n2854;
  assign n2860 = ~n37899 & ~n37900;
  assign n2861 = n2845 & ~n2860;
  assign n2862 = n2557 & ~n2559;
  assign n2863 = ~n2560 & ~n2862;
  assign n2864 = n649 & n2134;
  assign n2865 = pi80  & n37496;
  assign n2866 = pi82  & n662;
  assign n2867 = pi81  & n664;
  assign n2868 = ~n2866 & ~n2867;
  assign n2869 = ~n2865 & ~n2867;
  assign n2870 = ~n2866 & n2869;
  assign n2871 = ~n2865 & n2868;
  assign n2872 = ~n2864 & n37901;
  assign n2873 = pi32  & ~n2872;
  assign n2874 = pi32  & ~n2873;
  assign n2875 = pi32  & n2872;
  assign n2876 = ~n2872 & ~n2873;
  assign n2877 = ~pi32  & ~n2872;
  assign n2878 = ~n37902 & ~n37903;
  assign n2879 = n2863 & ~n2878;
  assign n2880 = n649 & n2154;
  assign n2881 = pi79  & n37496;
  assign n2882 = pi81  & n662;
  assign n2883 = pi80  & n664;
  assign n2884 = ~n2882 & ~n2883;
  assign n2885 = ~n2881 & ~n2883;
  assign n2886 = ~n2882 & n2885;
  assign n2887 = ~n2881 & n2884;
  assign n2888 = ~n2880 & n37904;
  assign n2889 = pi32  & ~n2888;
  assign n2890 = pi32  & ~n2889;
  assign n2891 = pi32  & n2888;
  assign n2892 = ~n2888 & ~n2889;
  assign n2893 = ~pi32  & ~n2888;
  assign n2894 = ~n37905 & ~n37906;
  assign n2895 = n2548 & n37841;
  assign n2896 = ~n2556 & ~n2895;
  assign n2897 = ~n2894 & n2896;
  assign n2898 = n2544 & ~n2546;
  assign n2899 = ~n2547 & ~n2898;
  assign n2900 = n649 & n2063;
  assign n2901 = pi78  & n37496;
  assign n2902 = pi80  & n662;
  assign n2903 = pi79  & n664;
  assign n2904 = ~n2902 & ~n2903;
  assign n2905 = ~n2901 & ~n2903;
  assign n2906 = ~n2902 & n2905;
  assign n2907 = ~n2901 & n2904;
  assign n2908 = ~n2900 & n37907;
  assign n2909 = pi32  & ~n2908;
  assign n2910 = pi32  & ~n2909;
  assign n2911 = pi32  & n2908;
  assign n2912 = ~n2908 & ~n2909;
  assign n2913 = ~pi32  & ~n2908;
  assign n2914 = ~n37908 & ~n37909;
  assign n2915 = n2899 & ~n2914;
  assign n2916 = n649 & n678;
  assign n2917 = pi77  & n37496;
  assign n2918 = pi79  & n662;
  assign n2919 = pi78  & n664;
  assign n2920 = ~n2918 & ~n2919;
  assign n2921 = ~n2917 & ~n2919;
  assign n2922 = ~n2918 & n2921;
  assign n2923 = ~n2917 & n2920;
  assign n2924 = ~n2916 & n37910;
  assign n2925 = pi32  & ~n2924;
  assign n2926 = pi32  & ~n2925;
  assign n2927 = pi32  & n2924;
  assign n2928 = ~n2924 & ~n2925;
  assign n2929 = ~pi32  & ~n2924;
  assign n2930 = ~n37911 & ~n37912;
  assign n2931 = n2535 & n37838;
  assign n2932 = ~n2535 & ~n2543;
  assign n2933 = ~n37838 & ~n2543;
  assign n2934 = ~n2932 & ~n2933;
  assign n2935 = ~n2543 & ~n2931;
  assign n2936 = ~n2930 & ~n37913;
  assign n2937 = n649 & n1578;
  assign n2938 = pi76  & n37496;
  assign n2939 = pi78  & n662;
  assign n2940 = pi77  & n664;
  assign n2941 = ~n2939 & ~n2940;
  assign n2942 = ~n2938 & ~n2940;
  assign n2943 = ~n2939 & n2942;
  assign n2944 = ~n2938 & n2941;
  assign n2945 = ~n2937 & n37914;
  assign n2946 = pi32  & ~n2945;
  assign n2947 = pi32  & ~n2946;
  assign n2948 = pi32  & n2945;
  assign n2949 = ~n2945 & ~n2946;
  assign n2950 = ~pi32  & ~n2945;
  assign n2951 = ~n37915 & ~n37916;
  assign n2952 = n2531 & ~n2533;
  assign n2953 = ~n2534 & ~n2952;
  assign n2954 = ~n2951 & n2953;
  assign n2955 = n649 & n1596;
  assign n2956 = pi75  & n37496;
  assign n2957 = pi77  & n662;
  assign n2958 = pi76  & n664;
  assign n2959 = ~n2957 & ~n2958;
  assign n2960 = ~n2956 & ~n2958;
  assign n2961 = ~n2957 & n2960;
  assign n2962 = ~n2956 & n2959;
  assign n2963 = ~n2955 & n37917;
  assign n2964 = pi32  & ~n2963;
  assign n2965 = pi32  & ~n2964;
  assign n2966 = pi32  & n2963;
  assign n2967 = ~n2963 & ~n2964;
  assign n2968 = ~pi32  & ~n2963;
  assign n2969 = ~n37918 & ~n37919;
  assign n2970 = n2525 & ~n2527;
  assign n2971 = ~n2525 & ~n37835;
  assign n2972 = ~n2526 & n2531;
  assign n2973 = ~n2971 & ~n2972;
  assign n2974 = ~n37835 & ~n2970;
  assign n2975 = ~n2969 & ~n37920;
  assign n2976 = n649 & n1465;
  assign n2977 = pi74  & n37496;
  assign n2978 = pi76  & n662;
  assign n2979 = pi75  & n664;
  assign n2980 = ~n2978 & ~n2979;
  assign n2981 = ~n2977 & ~n2979;
  assign n2982 = ~n2978 & n2981;
  assign n2983 = ~n2977 & n2980;
  assign n2984 = ~n2976 & n37921;
  assign n2985 = pi32  & ~n2984;
  assign n2986 = pi32  & ~n2985;
  assign n2987 = pi32  & n2984;
  assign n2988 = ~n2984 & ~n2985;
  assign n2989 = ~pi32  & ~n2984;
  assign n2990 = ~n37922 & ~n37923;
  assign n2991 = n2521 & ~n2523;
  assign n2992 = ~n2524 & ~n2991;
  assign n2993 = ~n2990 & n2992;
  assign n2994 = n649 & n720;
  assign n2995 = pi73  & n37496;
  assign n2996 = pi75  & n662;
  assign n2997 = pi74  & n664;
  assign n2998 = ~n2996 & ~n2997;
  assign n2999 = ~n2995 & ~n2997;
  assign n3000 = ~n2996 & n2999;
  assign n3001 = ~n2995 & n2998;
  assign n3002 = ~n2994 & n37924;
  assign n3003 = pi32  & ~n3002;
  assign n3004 = pi32  & ~n3003;
  assign n3005 = pi32  & n3002;
  assign n3006 = ~n3002 & ~n3003;
  assign n3007 = ~pi32  & ~n3002;
  assign n3008 = ~n37925 & ~n37926;
  assign n3009 = n2512 & n37834;
  assign n3010 = ~n2512 & ~n2520;
  assign n3011 = ~n2512 & n37834;
  assign n3012 = ~n37834 & ~n2520;
  assign n3013 = n2512 & ~n37834;
  assign n3014 = ~n37927 & ~n37928;
  assign n3015 = ~n2520 & ~n3009;
  assign n3016 = ~n3008 & ~n37929;
  assign n3017 = n2503 & n37831;
  assign n3018 = ~n2511 & ~n3017;
  assign n3019 = n649 & n1218;
  assign n3020 = pi72  & n37496;
  assign n3021 = pi74  & n662;
  assign n3022 = pi73  & n664;
  assign n3023 = ~n3021 & ~n3022;
  assign n3024 = ~n3020 & ~n3022;
  assign n3025 = ~n3021 & n3024;
  assign n3026 = ~n3020 & n3023;
  assign n3027 = ~n3019 & n37930;
  assign n3028 = pi32  & ~n3027;
  assign n3029 = pi32  & ~n3028;
  assign n3030 = pi32  & n3027;
  assign n3031 = ~n3027 & ~n3028;
  assign n3032 = ~pi32  & ~n3027;
  assign n3033 = ~n37931 & ~n37932;
  assign n3034 = n3018 & ~n3033;
  assign n3035 = n2494 & n37828;
  assign n3036 = ~n2502 & ~n3035;
  assign n3037 = n649 & n1238;
  assign n3038 = pi71  & n37496;
  assign n3039 = pi73  & n662;
  assign n3040 = pi72  & n664;
  assign n3041 = ~n3039 & ~n3040;
  assign n3042 = ~n3038 & ~n3040;
  assign n3043 = ~n3039 & n3042;
  assign n3044 = ~n3038 & n3041;
  assign n3045 = ~n3037 & n37933;
  assign n3046 = pi32  & ~n3045;
  assign n3047 = pi32  & ~n3046;
  assign n3048 = pi32  & n3045;
  assign n3049 = ~n3045 & ~n3046;
  assign n3050 = ~pi32  & ~n3045;
  assign n3051 = ~n37934 & ~n37935;
  assign n3052 = n3036 & ~n3051;
  assign n3053 = n649 & n1124;
  assign n3054 = pi70  & n37496;
  assign n3055 = pi72  & n662;
  assign n3056 = pi71  & n664;
  assign n3057 = ~n3055 & ~n3056;
  assign n3058 = ~n3054 & ~n3056;
  assign n3059 = ~n3055 & n3058;
  assign n3060 = ~n3054 & n3057;
  assign n3061 = ~n3053 & n37936;
  assign n3062 = pi32  & ~n3061;
  assign n3063 = pi32  & ~n3062;
  assign n3064 = pi32  & n3061;
  assign n3065 = ~n3061 & ~n3062;
  assign n3066 = ~pi32  & ~n3061;
  assign n3067 = ~n37937 & ~n37938;
  assign n3068 = n2485 & n37825;
  assign n3069 = ~n2485 & n37825;
  assign n3070 = n2485 & ~n37825;
  assign n3071 = ~n3069 & ~n3070;
  assign n3072 = ~n2493 & ~n3068;
  assign n3073 = ~n3067 & ~n37939;
  assign n3074 = n649 & n927;
  assign n3075 = pi69  & n37496;
  assign n3076 = pi71  & n662;
  assign n3077 = pi70  & n664;
  assign n3078 = ~n3076 & ~n3077;
  assign n3079 = ~n3075 & ~n3077;
  assign n3080 = ~n3076 & n3079;
  assign n3081 = ~n3075 & n3078;
  assign n3082 = ~n3074 & n37940;
  assign n3083 = pi32  & ~n3082;
  assign n3084 = pi32  & ~n3083;
  assign n3085 = pi32  & n3082;
  assign n3086 = ~n3082 & ~n3083;
  assign n3087 = ~pi32  & ~n3082;
  assign n3088 = ~n37941 & ~n37942;
  assign n3089 = n2481 & ~n2483;
  assign n3090 = ~n2484 & ~n3089;
  assign n3091 = ~n3088 & n3090;
  assign n3092 = n2474 & n37822;
  assign n3093 = ~n2480 & ~n3092;
  assign n3094 = n649 & n972;
  assign n3095 = pi68  & n37496;
  assign n3096 = pi70  & n662;
  assign n3097 = pi69  & n664;
  assign n3098 = ~n3096 & ~n3097;
  assign n3099 = ~n3095 & ~n3097;
  assign n3100 = ~n3096 & n3099;
  assign n3101 = ~n3095 & n3098;
  assign n3102 = ~n3094 & n37943;
  assign n3103 = pi32  & ~n3102;
  assign n3104 = pi32  & ~n3103;
  assign n3105 = pi32  & n3102;
  assign n3106 = ~n3102 & ~n3103;
  assign n3107 = ~pi32  & ~n3102;
  assign n3108 = ~n37944 & ~n37945;
  assign n3109 = n3093 & ~n3108;
  assign n3110 = n649 & n990;
  assign n3111 = pi67  & n37496;
  assign n3112 = pi69  & n662;
  assign n3113 = pi68  & n664;
  assign n3114 = ~n3112 & ~n3113;
  assign n3115 = ~n3111 & ~n3113;
  assign n3116 = ~n3112 & n3115;
  assign n3117 = ~n3111 & n3114;
  assign n3118 = ~n3110 & n37946;
  assign n3119 = pi32  & ~n3118;
  assign n3120 = pi32  & ~n3119;
  assign n3121 = pi32  & n3118;
  assign n3122 = ~n3118 & ~n3119;
  assign n3123 = ~pi32  & ~n3118;
  assign n3124 = ~n37947 & ~n37948;
  assign n3125 = pi35  & ~n37814;
  assign n3126 = n37817 & ~n3125;
  assign n3127 = ~n37817 & n3125;
  assign n3128 = ~n37814 & n2456;
  assign n3129 = ~n37818 & ~n3128;
  assign n3130 = ~n3126 & ~n3127;
  assign n3131 = ~n3124 & n37949;
  assign n3132 = n649 & n871;
  assign n3133 = pi66  & n37496;
  assign n3134 = pi68  & n662;
  assign n3135 = pi67  & n664;
  assign n3136 = ~n3134 & ~n3135;
  assign n3137 = ~n3133 & ~n3135;
  assign n3138 = ~n3134 & n3137;
  assign n3139 = ~n3133 & n3136;
  assign n3140 = ~n3132 & n37950;
  assign n3141 = pi32  & ~n3140;
  assign n3142 = pi32  & ~n3141;
  assign n3143 = pi32  & n3140;
  assign n3144 = ~n3140 & ~n3141;
  assign n3145 = ~pi32  & ~n3140;
  assign n3146 = ~n37951 & ~n37952;
  assign n3147 = pi35  & n2430;
  assign n3148 = ~n2429 & n3147;
  assign n3149 = n2429 & ~n3147;
  assign n3150 = ~n2431 & n2435;
  assign n3151 = ~n37814 & ~n3150;
  assign n3152 = ~n3148 & ~n3149;
  assign n3153 = ~n3146 & n37953;
  assign n3154 = n649 & n37515;
  assign n3155 = pi65  & n662;
  assign n3156 = pi64  & n664;
  assign n3157 = ~n3155 & ~n3156;
  assign n3158 = ~n3154 & n3157;
  assign n3159 = pi64  & n37493;
  assign n3160 = pi32  & ~n3159;
  assign n3161 = pi32  & ~n3158;
  assign n3162 = pi32  & ~n3161;
  assign n3163 = ~n3158 & ~n3161;
  assign n3164 = ~n3162 & ~n3163;
  assign n3165 = n3160 & ~n3164;
  assign n3166 = n3158 & n3160;
  assign n3167 = pi64  & n37496;
  assign n3168 = pi65  & n664;
  assign n3169 = n649 & ~n37521;
  assign n3170 = pi66  & n662;
  assign n3171 = ~n3169 & ~n3170;
  assign n3172 = ~n3168 & ~n3169;
  assign n3173 = ~n3170 & n3172;
  assign n3174 = ~n3168 & ~n3170;
  assign n3175 = ~n3169 & n3174;
  assign n3176 = ~n3168 & n3171;
  assign n3177 = ~n3167 & ~n3168;
  assign n3178 = ~n3170 & n3177;
  assign n3179 = ~n3167 & n3174;
  assign n3180 = ~n3169 & n37956;
  assign n3181 = ~n3167 & n37955;
  assign n3182 = pi32  & ~n37957;
  assign n3183 = pi32  & ~n3182;
  assign n3184 = ~n37957 & ~n3182;
  assign n3185 = ~n3183 & ~n3184;
  assign n3186 = n37954 & ~n3185;
  assign n3187 = n37954 & n37957;
  assign n3188 = n2430 & n37958;
  assign n3189 = n649 & n847;
  assign n3190 = pi65  & n37496;
  assign n3191 = pi67  & n662;
  assign n3192 = pi66  & n664;
  assign n3193 = ~n3191 & ~n3192;
  assign n3194 = ~n3190 & ~n3192;
  assign n3195 = ~n3191 & n3194;
  assign n3196 = ~n3190 & n3193;
  assign n3197 = ~n3189 & n37959;
  assign n3198 = pi32  & ~n3197;
  assign n3199 = pi32  & ~n3198;
  assign n3200 = pi32  & n3197;
  assign n3201 = ~n3197 & ~n3198;
  assign n3202 = ~pi32  & ~n3197;
  assign n3203 = ~n37960 & ~n37961;
  assign n3204 = ~n2430 & ~n37958;
  assign n3205 = n2430 & ~n37958;
  assign n3206 = ~n2430 & n37958;
  assign n3207 = ~n3205 & ~n3206;
  assign n3208 = ~n3188 & ~n3204;
  assign n3209 = ~n3203 & ~n37962;
  assign n3210 = ~n3188 & ~n3209;
  assign n3211 = n3146 & ~n37953;
  assign n3212 = ~n3153 & ~n3211;
  assign n3213 = ~n3210 & n3212;
  assign n3214 = ~n3153 & ~n3213;
  assign n3215 = n3124 & ~n37949;
  assign n3216 = ~n3131 & ~n3215;
  assign n3217 = ~n3214 & ~n3215;
  assign n3218 = ~n3131 & n3217;
  assign n3219 = ~n3214 & n3216;
  assign n3220 = ~n3131 & ~n37963;
  assign n3221 = ~n3093 & n3108;
  assign n3222 = n3093 & ~n3109;
  assign n3223 = n3093 & n3108;
  assign n3224 = ~n3108 & ~n3109;
  assign n3225 = ~n3093 & ~n3108;
  assign n3226 = ~n37964 & ~n37965;
  assign n3227 = ~n3109 & ~n3221;
  assign n3228 = ~n3220 & ~n37966;
  assign n3229 = ~n3109 & ~n3228;
  assign n3230 = n3088 & ~n3090;
  assign n3231 = ~n3091 & ~n3230;
  assign n3232 = ~n3229 & n3231;
  assign n3233 = ~n3091 & ~n3232;
  assign n3234 = n3067 & n37939;
  assign n3235 = ~n3073 & ~n3234;
  assign n3236 = ~n3233 & n3235;
  assign n3237 = ~n3073 & ~n3236;
  assign n3238 = ~n3036 & n3051;
  assign n3239 = n3036 & ~n3052;
  assign n3240 = n3036 & n3051;
  assign n3241 = ~n3051 & ~n3052;
  assign n3242 = ~n3036 & ~n3051;
  assign n3243 = ~n37967 & ~n37968;
  assign n3244 = ~n3052 & ~n3238;
  assign n3245 = ~n3237 & ~n37969;
  assign n3246 = ~n3052 & ~n3245;
  assign n3247 = ~n3018 & n3033;
  assign n3248 = ~n3034 & ~n3247;
  assign n3249 = ~n3246 & ~n3247;
  assign n3250 = ~n3034 & n3249;
  assign n3251 = ~n3246 & n3248;
  assign n3252 = ~n3034 & ~n37970;
  assign n3253 = n3008 & n37929;
  assign n3254 = ~n3016 & ~n3253;
  assign n3255 = ~n3252 & n3254;
  assign n3256 = ~n3016 & ~n3255;
  assign n3257 = n2990 & ~n2992;
  assign n3258 = ~n2990 & ~n2993;
  assign n3259 = ~n2990 & ~n2992;
  assign n3260 = n2992 & ~n2993;
  assign n3261 = n2990 & n2992;
  assign n3262 = ~n37971 & ~n37972;
  assign n3263 = ~n2993 & ~n3257;
  assign n3264 = ~n3256 & ~n37973;
  assign n3265 = ~n2993 & ~n3264;
  assign n3266 = n2969 & n37920;
  assign n3267 = ~n2975 & ~n3266;
  assign n3268 = ~n3265 & n3267;
  assign n3269 = ~n2975 & ~n3268;
  assign n3270 = n2951 & ~n2953;
  assign n3271 = ~n2954 & ~n3270;
  assign n3272 = ~n3269 & n3271;
  assign n3273 = ~n2954 & ~n3272;
  assign n3274 = n2930 & n37913;
  assign n3275 = ~n37913 & ~n2936;
  assign n3276 = n2930 & ~n37913;
  assign n3277 = ~n2930 & ~n2936;
  assign n3278 = ~n2930 & n37913;
  assign n3279 = ~n37974 & ~n37975;
  assign n3280 = ~n2936 & ~n3274;
  assign n3281 = ~n3273 & ~n37976;
  assign n3282 = ~n2936 & ~n3281;
  assign n3283 = ~n2899 & n2914;
  assign n3284 = n2899 & ~n2915;
  assign n3285 = n2899 & n2914;
  assign n3286 = ~n2914 & ~n2915;
  assign n3287 = ~n2899 & ~n2914;
  assign n3288 = ~n37977 & ~n37978;
  assign n3289 = ~n2915 & ~n3283;
  assign n3290 = ~n3282 & ~n37979;
  assign n3291 = ~n2915 & ~n3290;
  assign n3292 = n2894 & ~n2896;
  assign n3293 = ~n2894 & ~n2897;
  assign n3294 = ~n2894 & ~n2896;
  assign n3295 = n2896 & ~n2897;
  assign n3296 = n2894 & n2896;
  assign n3297 = ~n37980 & ~n37981;
  assign n3298 = ~n2897 & ~n3292;
  assign n3299 = ~n3291 & ~n37982;
  assign n3300 = ~n2897 & ~n3299;
  assign n3301 = ~n2863 & n2878;
  assign n3302 = n2863 & ~n2879;
  assign n3303 = n2863 & n2878;
  assign n3304 = ~n2878 & ~n2879;
  assign n3305 = ~n2863 & ~n2878;
  assign n3306 = ~n37983 & ~n37984;
  assign n3307 = ~n2879 & ~n3301;
  assign n3308 = ~n3300 & ~n37985;
  assign n3309 = ~n2879 & ~n3308;
  assign n3310 = ~n2845 & n2860;
  assign n3311 = n2845 & ~n2861;
  assign n3312 = n2845 & n2860;
  assign n3313 = ~n2860 & ~n2861;
  assign n3314 = ~n2845 & ~n2860;
  assign n3315 = ~n37986 & ~n37987;
  assign n3316 = ~n2861 & ~n3310;
  assign n3317 = ~n3309 & ~n37988;
  assign n3318 = ~n2861 & ~n3317;
  assign n3319 = n2835 & n37897;
  assign n3320 = ~n37897 & ~n2843;
  assign n3321 = ~n2835 & ~n2843;
  assign n3322 = ~n3320 & ~n3321;
  assign n3323 = ~n2843 & ~n3319;
  assign n3324 = ~n3318 & ~n37989;
  assign n3325 = ~n2843 & ~n3324;
  assign n3326 = ~n2802 & n2819;
  assign n3327 = n2802 & ~n2820;
  assign n3328 = n2802 & n2819;
  assign n3329 = ~n2819 & ~n2820;
  assign n3330 = ~n2802 & ~n2819;
  assign n3331 = ~n37990 & ~n37991;
  assign n3332 = ~n2820 & ~n3326;
  assign n3333 = ~n3325 & ~n37992;
  assign n3334 = ~n2820 & ~n3333;
  assign n3335 = n2794 & n37888;
  assign n3336 = ~n37888 & ~n2800;
  assign n3337 = n2794 & ~n37888;
  assign n3338 = ~n2794 & ~n2800;
  assign n3339 = ~n2794 & n37888;
  assign n3340 = ~n37993 & ~n37994;
  assign n3341 = ~n2800 & ~n3335;
  assign n3342 = ~n3334 & ~n37995;
  assign n3343 = ~n2800 & ~n3342;
  assign n3344 = n676 & ~n2776;
  assign n3345 = ~n676 & ~n2777;
  assign n3346 = ~n676 & ~n2776;
  assign n3347 = n2776 & ~n2777;
  assign n3348 = n676 & n2776;
  assign n3349 = ~n37996 & ~n37997;
  assign n3350 = ~n2777 & ~n3344;
  assign n3351 = ~n3343 & ~n37998;
  assign n3352 = ~n2777 & ~n3351;
  assign n3353 = n409 & ~n411;
  assign n3354 = ~n412 & ~n3353;
  assign n3355 = n649 & n3354;
  assign n3356 = pi86  & n37496;
  assign n3357 = pi88  & n662;
  assign n3358 = pi87  & n664;
  assign n3359 = ~n3357 & ~n3358;
  assign n3360 = ~n3356 & ~n3358;
  assign n3361 = ~n3357 & n3360;
  assign n3362 = ~n3356 & n3359;
  assign n3363 = ~n3355 & n37999;
  assign n3364 = pi32  & ~n3363;
  assign n3365 = pi32  & ~n3364;
  assign n3366 = pi32  & n3363;
  assign n3367 = ~n3363 & ~n3364;
  assign n3368 = ~pi32  & ~n3363;
  assign n3369 = ~n38000 & ~n38001;
  assign n3370 = ~n2768 & ~n2774;
  assign n3371 = n2104 & n2804;
  assign n3372 = pi83  & n37758;
  assign n3373 = pi85  & n2117;
  assign n3374 = pi84  & n2119;
  assign n3375 = ~n3373 & ~n3374;
  assign n3376 = ~n3372 & ~n3374;
  assign n3377 = ~n3373 & n3376;
  assign n3378 = ~n3372 & n3375;
  assign n3379 = ~n3371 & n38002;
  assign n3380 = pi35  & ~n3379;
  assign n3381 = pi35  & ~n3380;
  assign n3382 = pi35  & n3379;
  assign n3383 = ~n3379 & ~n3380;
  assign n3384 = ~pi35  & ~n3379;
  assign n3385 = ~n38003 & ~n38004;
  assign n3386 = ~n2752 & ~n2760;
  assign n3387 = n691 & n2134;
  assign n3388 = pi80  & n37503;
  assign n3389 = pi82  & n704;
  assign n3390 = pi81  & n706;
  assign n3391 = ~n3389 & ~n3390;
  assign n3392 = ~n3388 & ~n3390;
  assign n3393 = ~n3389 & n3392;
  assign n3394 = ~n3388 & n3391;
  assign n3395 = ~n3387 & n38005;
  assign n3396 = pi38  & ~n3395;
  assign n3397 = pi38  & ~n3396;
  assign n3398 = pi38  & n3395;
  assign n3399 = ~n3395 & ~n3396;
  assign n3400 = ~pi38  & ~n3395;
  assign n3401 = ~n38006 & ~n38007;
  assign n3402 = ~n2741 & ~n2749;
  assign n3403 = n678 & n733;
  assign n3404 = pi77  & n37510;
  assign n3405 = pi79  & n746;
  assign n3406 = pi78  & n748;
  assign n3407 = ~n3405 & ~n3406;
  assign n3408 = ~n3404 & ~n3406;
  assign n3409 = ~n3405 & n3408;
  assign n3410 = ~n3404 & n3407;
  assign n3411 = ~n3403 & n38008;
  assign n3412 = pi41  & ~n3411;
  assign n3413 = pi41  & ~n3412;
  assign n3414 = pi41  & n3411;
  assign n3415 = ~n3411 & ~n3412;
  assign n3416 = ~pi41  & ~n3411;
  assign n3417 = ~n38009 & ~n38010;
  assign n3418 = ~n2721 & ~n2723;
  assign n3419 = n940 & n1465;
  assign n3420 = pi74  & n37541;
  assign n3421 = pi76  & n953;
  assign n3422 = pi75  & n955;
  assign n3423 = ~n3421 & ~n3422;
  assign n3424 = ~n3420 & ~n3422;
  assign n3425 = ~n3421 & n3424;
  assign n3426 = ~n3420 & n3423;
  assign n3427 = ~n3419 & n38011;
  assign n3428 = pi44  & ~n3427;
  assign n3429 = pi44  & ~n3428;
  assign n3430 = pi44  & n3427;
  assign n3431 = ~n3427 & ~n3428;
  assign n3432 = ~pi44  & ~n3427;
  assign n3433 = ~n38012 & ~n38013;
  assign n3434 = ~n2715 & ~n2717;
  assign n3435 = n785 & n1238;
  assign n3436 = pi71  & n37520;
  assign n3437 = pi73  & n787;
  assign n3438 = pi72  & n795;
  assign n3439 = ~n3437 & ~n3438;
  assign n3440 = ~n3436 & ~n3438;
  assign n3441 = ~n3437 & n3440;
  assign n3442 = ~n3436 & n3439;
  assign n3443 = ~n3435 & n38014;
  assign n3444 = pi47  & ~n3443;
  assign n3445 = pi47  & ~n3444;
  assign n3446 = pi47  & n3443;
  assign n3447 = ~n3443 & ~n3444;
  assign n3448 = ~pi47  & ~n3443;
  assign n3449 = ~n38015 & ~n38016;
  assign n3450 = n847 & n1971;
  assign n3451 = pi65  & n37864;
  assign n3452 = pi67  & n1973;
  assign n3453 = pi66  & n1981;
  assign n3454 = ~n3452 & ~n3453;
  assign n3455 = ~n3451 & ~n3453;
  assign n3456 = ~n3452 & n3455;
  assign n3457 = ~n3451 & n3454;
  assign n3458 = ~n3450 & n38017;
  assign n3459 = pi53  & ~n3458;
  assign n3460 = pi53  & ~n3459;
  assign n3461 = pi53  & n3458;
  assign n3462 = ~n3458 & ~n3459;
  assign n3463 = ~pi53  & ~n3458;
  assign n3464 = ~n38018 & ~n38019;
  assign n3465 = pi53  & ~pi54 ;
  assign n3466 = ~pi53  & pi54 ;
  assign n3467 = ~pi53  & ~pi54 ;
  assign n3468 = pi53  & pi54 ;
  assign n3469 = ~n3467 & ~n3468;
  assign n3470 = ~n3465 & ~n3466;
  assign n3471 = pi64  & n38020;
  assign n3472 = n37868 & n3471;
  assign n3473 = ~n37868 & ~n3471;
  assign n3474 = ~n37868 & n3471;
  assign n3475 = n37868 & ~n3471;
  assign n3476 = ~n3474 & ~n3475;
  assign n3477 = ~n3472 & ~n3473;
  assign n3478 = ~n3464 & ~n38021;
  assign n3479 = n3464 & n38021;
  assign n3480 = ~n3478 & ~n3479;
  assign n3481 = n894 & n972;
  assign n3482 = pi68  & n37580;
  assign n3483 = pi70  & n896;
  assign n3484 = pi69  & n904;
  assign n3485 = ~n3483 & ~n3484;
  assign n3486 = ~n3482 & ~n3484;
  assign n3487 = ~n3483 & n3486;
  assign n3488 = ~n3482 & n3485;
  assign n3489 = ~n3481 & n38022;
  assign n3490 = pi50  & ~n3489;
  assign n3491 = pi50  & ~n3490;
  assign n3492 = pi50  & n3489;
  assign n3493 = ~n3489 & ~n3490;
  assign n3494 = ~pi50  & ~n3489;
  assign n3495 = ~n38023 & ~n38024;
  assign n3496 = n3480 & ~n3495;
  assign n3497 = ~n3480 & n3495;
  assign n3498 = n3480 & ~n3496;
  assign n3499 = n3480 & n3495;
  assign n3500 = ~n3495 & ~n3496;
  assign n3501 = ~n3480 & ~n3495;
  assign n3502 = ~n38025 & ~n38026;
  assign n3503 = ~n3496 & ~n3497;
  assign n3504 = ~n2710 & ~n38027;
  assign n3505 = n2710 & n38027;
  assign n3506 = ~n3504 & ~n3505;
  assign n3507 = ~n3449 & n3506;
  assign n3508 = n3449 & ~n3506;
  assign n3509 = ~n3449 & ~n3507;
  assign n3510 = ~n3449 & ~n3506;
  assign n3511 = n3506 & ~n3507;
  assign n3512 = n3449 & n3506;
  assign n3513 = ~n38028 & ~n38029;
  assign n3514 = ~n3507 & ~n3508;
  assign n3515 = ~n3434 & ~n38030;
  assign n3516 = n3434 & ~n38029;
  assign n3517 = ~n38028 & n3516;
  assign n3518 = n3434 & n38030;
  assign n3519 = ~n3515 & ~n38031;
  assign n3520 = ~n3433 & n3519;
  assign n3521 = n3433 & ~n3519;
  assign n3522 = ~n3433 & ~n3520;
  assign n3523 = ~n3433 & ~n3519;
  assign n3524 = n3519 & ~n3520;
  assign n3525 = n3433 & n3519;
  assign n3526 = ~n38032 & ~n38033;
  assign n3527 = ~n3520 & ~n3521;
  assign n3528 = ~n3418 & ~n38034;
  assign n3529 = n3418 & ~n38033;
  assign n3530 = ~n38032 & n3529;
  assign n3531 = n3418 & n38034;
  assign n3532 = ~n3528 & ~n38035;
  assign n3533 = ~n3417 & n3532;
  assign n3534 = n3417 & ~n3532;
  assign n3535 = ~n3533 & ~n3534;
  assign n3536 = ~n3402 & n3535;
  assign n3537 = n3402 & ~n3535;
  assign n3538 = ~n3536 & ~n3537;
  assign n3539 = ~n3401 & n3538;
  assign n3540 = n3401 & ~n3538;
  assign n3541 = ~n3401 & ~n3539;
  assign n3542 = ~n3401 & ~n3538;
  assign n3543 = n3538 & ~n3539;
  assign n3544 = n3401 & n3538;
  assign n3545 = ~n38036 & ~n38037;
  assign n3546 = ~n3539 & ~n3540;
  assign n3547 = ~n3386 & ~n38038;
  assign n3548 = n3386 & ~n38037;
  assign n3549 = ~n38036 & n3548;
  assign n3550 = n3386 & n38038;
  assign n3551 = ~n3547 & ~n38039;
  assign n3552 = ~n3385 & n3551;
  assign n3553 = n3385 & ~n3551;
  assign n3554 = ~n3552 & ~n3553;
  assign n3555 = ~n3370 & n3554;
  assign n3556 = n3370 & ~n3554;
  assign n3557 = ~n3555 & ~n3556;
  assign n3558 = ~n3369 & n3557;
  assign n3559 = n3369 & ~n3557;
  assign n3560 = ~n3558 & ~n3559;
  assign n3561 = ~n3352 & n3560;
  assign n3562 = n3352 & ~n3560;
  assign n3563 = ~n3561 & ~n3562;
  assign n3564 = ~n634 & n3563;
  assign n3565 = n417 & ~n419;
  assign n3566 = ~n420 & ~n3565;
  assign n3567 = n607 & n3566;
  assign n3568 = pi88  & n37489;
  assign n3569 = pi90  & n620;
  assign n3570 = pi89  & n622;
  assign n3571 = ~n3569 & ~n3570;
  assign n3572 = ~n3568 & ~n3570;
  assign n3573 = ~n3569 & n3572;
  assign n3574 = ~n3568 & n3571;
  assign n3575 = ~n3567 & n38040;
  assign n3576 = pi29  & ~n3575;
  assign n3577 = pi29  & ~n3576;
  assign n3578 = pi29  & n3575;
  assign n3579 = ~n3575 & ~n3576;
  assign n3580 = ~pi29  & ~n3575;
  assign n3581 = ~n38041 & ~n38042;
  assign n3582 = n3343 & n37998;
  assign n3583 = ~n3343 & ~n3351;
  assign n3584 = ~n37998 & ~n3351;
  assign n3585 = ~n3583 & ~n3584;
  assign n3586 = ~n3351 & ~n3582;
  assign n3587 = ~n3581 & ~n38043;
  assign n3588 = n3334 & n37995;
  assign n3589 = ~n3342 & ~n3588;
  assign n3590 = n413 & ~n415;
  assign n3591 = ~n416 & ~n3590;
  assign n3592 = n607 & n3591;
  assign n3593 = pi87  & n37489;
  assign n3594 = pi89  & n620;
  assign n3595 = pi88  & n622;
  assign n3596 = ~n3594 & ~n3595;
  assign n3597 = ~n3593 & ~n3595;
  assign n3598 = ~n3594 & n3597;
  assign n3599 = ~n3593 & n3596;
  assign n3600 = ~n3592 & n38044;
  assign n3601 = pi29  & ~n3600;
  assign n3602 = pi29  & ~n3601;
  assign n3603 = pi29  & n3600;
  assign n3604 = ~n3600 & ~n3601;
  assign n3605 = ~pi29  & ~n3600;
  assign n3606 = ~n38045 & ~n38046;
  assign n3607 = n3589 & ~n3606;
  assign n3608 = n3325 & n37992;
  assign n3609 = ~n3333 & ~n3608;
  assign n3610 = n607 & n3354;
  assign n3611 = pi86  & n37489;
  assign n3612 = pi88  & n620;
  assign n3613 = pi87  & n622;
  assign n3614 = ~n3612 & ~n3613;
  assign n3615 = ~n3611 & ~n3613;
  assign n3616 = ~n3612 & n3615;
  assign n3617 = ~n3611 & n3614;
  assign n3618 = ~n3610 & n38047;
  assign n3619 = pi29  & ~n3618;
  assign n3620 = pi29  & ~n3619;
  assign n3621 = pi29  & n3618;
  assign n3622 = ~n3618 & ~n3619;
  assign n3623 = ~pi29  & ~n3618;
  assign n3624 = ~n38048 & ~n38049;
  assign n3625 = n3609 & ~n3624;
  assign n3626 = n3318 & n37989;
  assign n3627 = ~n3324 & ~n3626;
  assign n3628 = n607 & n636;
  assign n3629 = pi85  & n37489;
  assign n3630 = pi87  & n620;
  assign n3631 = pi86  & n622;
  assign n3632 = ~n3630 & ~n3631;
  assign n3633 = ~n3629 & ~n3631;
  assign n3634 = ~n3630 & n3633;
  assign n3635 = ~n3629 & n3632;
  assign n3636 = ~n3628 & n38050;
  assign n3637 = pi29  & ~n3636;
  assign n3638 = pi29  & ~n3637;
  assign n3639 = pi29  & n3636;
  assign n3640 = ~n3636 & ~n3637;
  assign n3641 = ~pi29  & ~n3636;
  assign n3642 = ~n38051 & ~n38052;
  assign n3643 = n3627 & ~n3642;
  assign n3644 = n3309 & n37988;
  assign n3645 = ~n3317 & ~n3644;
  assign n3646 = n607 & n2779;
  assign n3647 = pi84  & n37489;
  assign n3648 = pi86  & n620;
  assign n3649 = pi85  & n622;
  assign n3650 = ~n3648 & ~n3649;
  assign n3651 = ~n3647 & ~n3649;
  assign n3652 = ~n3648 & n3651;
  assign n3653 = ~n3647 & n3650;
  assign n3654 = ~n3646 & n38053;
  assign n3655 = pi29  & ~n3654;
  assign n3656 = pi29  & ~n3655;
  assign n3657 = pi29  & n3654;
  assign n3658 = ~n3654 & ~n3655;
  assign n3659 = ~pi29  & ~n3654;
  assign n3660 = ~n38054 & ~n38055;
  assign n3661 = n3645 & ~n3660;
  assign n3662 = n3300 & n37985;
  assign n3663 = ~n3308 & ~n3662;
  assign n3664 = n607 & n2804;
  assign n3665 = pi83  & n37489;
  assign n3666 = pi85  & n620;
  assign n3667 = pi84  & n622;
  assign n3668 = ~n3666 & ~n3667;
  assign n3669 = ~n3665 & ~n3667;
  assign n3670 = ~n3666 & n3669;
  assign n3671 = ~n3665 & n3668;
  assign n3672 = ~n3664 & n38056;
  assign n3673 = pi29  & ~n3672;
  assign n3674 = pi29  & ~n3673;
  assign n3675 = pi29  & n3672;
  assign n3676 = ~n3672 & ~n3673;
  assign n3677 = ~pi29  & ~n3672;
  assign n3678 = ~n38057 & ~n38058;
  assign n3679 = n3663 & ~n3678;
  assign n3680 = n607 & n2591;
  assign n3681 = pi82  & n37489;
  assign n3682 = pi84  & n620;
  assign n3683 = pi83  & n622;
  assign n3684 = ~n3682 & ~n3683;
  assign n3685 = ~n3681 & ~n3683;
  assign n3686 = ~n3682 & n3685;
  assign n3687 = ~n3681 & n3684;
  assign n3688 = ~n3680 & n38059;
  assign n3689 = pi29  & ~n3688;
  assign n3690 = pi29  & ~n3689;
  assign n3691 = pi29  & n3688;
  assign n3692 = ~n3688 & ~n3689;
  assign n3693 = ~pi29  & ~n3688;
  assign n3694 = ~n38060 & ~n38061;
  assign n3695 = n3291 & n37982;
  assign n3696 = ~n3291 & ~n3299;
  assign n3697 = ~n3291 & n37982;
  assign n3698 = ~n37982 & ~n3299;
  assign n3699 = n3291 & ~n37982;
  assign n3700 = ~n38062 & ~n38063;
  assign n3701 = ~n3299 & ~n3695;
  assign n3702 = ~n3694 & ~n38064;
  assign n3703 = n3282 & n37979;
  assign n3704 = ~n3290 & ~n3703;
  assign n3705 = n607 & n2091;
  assign n3706 = pi81  & n37489;
  assign n3707 = pi83  & n620;
  assign n3708 = pi82  & n622;
  assign n3709 = ~n3707 & ~n3708;
  assign n3710 = ~n3706 & ~n3708;
  assign n3711 = ~n3707 & n3710;
  assign n3712 = ~n3706 & n3709;
  assign n3713 = ~n3705 & n38065;
  assign n3714 = pi29  & ~n3713;
  assign n3715 = pi29  & ~n3714;
  assign n3716 = pi29  & n3713;
  assign n3717 = ~n3713 & ~n3714;
  assign n3718 = ~pi29  & ~n3713;
  assign n3719 = ~n38066 & ~n38067;
  assign n3720 = n3704 & ~n3719;
  assign n3721 = n607 & n2134;
  assign n3722 = pi80  & n37489;
  assign n3723 = pi82  & n620;
  assign n3724 = pi81  & n622;
  assign n3725 = ~n3723 & ~n3724;
  assign n3726 = ~n3722 & ~n3724;
  assign n3727 = ~n3723 & n3726;
  assign n3728 = ~n3722 & n3725;
  assign n3729 = ~n3721 & n38068;
  assign n3730 = pi29  & ~n3729;
  assign n3731 = pi29  & ~n3730;
  assign n3732 = pi29  & n3729;
  assign n3733 = ~n3729 & ~n3730;
  assign n3734 = ~pi29  & ~n3729;
  assign n3735 = ~n38069 & ~n38070;
  assign n3736 = n3273 & n37976;
  assign n3737 = ~n3273 & n37976;
  assign n3738 = n3273 & ~n37976;
  assign n3739 = ~n3737 & ~n3738;
  assign n3740 = ~n3281 & ~n3736;
  assign n3741 = ~n3735 & ~n38071;
  assign n3742 = n607 & n2154;
  assign n3743 = pi79  & n37489;
  assign n3744 = pi81  & n620;
  assign n3745 = pi80  & n622;
  assign n3746 = ~n3744 & ~n3745;
  assign n3747 = ~n3743 & ~n3745;
  assign n3748 = ~n3744 & n3747;
  assign n3749 = ~n3743 & n3746;
  assign n3750 = ~n3742 & n38072;
  assign n3751 = pi29  & ~n3750;
  assign n3752 = pi29  & ~n3751;
  assign n3753 = pi29  & n3750;
  assign n3754 = ~n3750 & ~n3751;
  assign n3755 = ~pi29  & ~n3750;
  assign n3756 = ~n38073 & ~n38074;
  assign n3757 = n3269 & ~n3271;
  assign n3758 = ~n3272 & ~n3757;
  assign n3759 = ~n3756 & n3758;
  assign n3760 = n3265 & ~n3267;
  assign n3761 = ~n3268 & ~n3760;
  assign n3762 = n607 & n2063;
  assign n3763 = pi78  & n37489;
  assign n3764 = pi80  & n620;
  assign n3765 = pi79  & n622;
  assign n3766 = ~n3764 & ~n3765;
  assign n3767 = ~n3763 & ~n3765;
  assign n3768 = ~n3764 & n3767;
  assign n3769 = ~n3763 & n3766;
  assign n3770 = ~n3762 & n38075;
  assign n3771 = pi29  & ~n3770;
  assign n3772 = pi29  & ~n3771;
  assign n3773 = pi29  & n3770;
  assign n3774 = ~n3770 & ~n3771;
  assign n3775 = ~pi29  & ~n3770;
  assign n3776 = ~n38076 & ~n38077;
  assign n3777 = n3761 & ~n3776;
  assign n3778 = n607 & n678;
  assign n3779 = pi77  & n37489;
  assign n3780 = pi79  & n620;
  assign n3781 = pi78  & n622;
  assign n3782 = ~n3780 & ~n3781;
  assign n3783 = ~n3779 & ~n3781;
  assign n3784 = ~n3780 & n3783;
  assign n3785 = ~n3779 & n3782;
  assign n3786 = ~n3778 & n38078;
  assign n3787 = pi29  & ~n3786;
  assign n3788 = pi29  & ~n3787;
  assign n3789 = pi29  & n3786;
  assign n3790 = ~n3786 & ~n3787;
  assign n3791 = ~pi29  & ~n3786;
  assign n3792 = ~n38079 & ~n38080;
  assign n3793 = n3256 & n37973;
  assign n3794 = ~n3256 & ~n3264;
  assign n3795 = ~n37973 & ~n3264;
  assign n3796 = ~n3794 & ~n3795;
  assign n3797 = ~n3264 & ~n3793;
  assign n3798 = ~n3792 & ~n38081;
  assign n3799 = n607 & n1578;
  assign n3800 = pi76  & n37489;
  assign n3801 = pi78  & n620;
  assign n3802 = pi77  & n622;
  assign n3803 = ~n3801 & ~n3802;
  assign n3804 = ~n3800 & ~n3802;
  assign n3805 = ~n3801 & n3804;
  assign n3806 = ~n3800 & n3803;
  assign n3807 = ~n3799 & n38082;
  assign n3808 = pi29  & ~n3807;
  assign n3809 = pi29  & ~n3808;
  assign n3810 = pi29  & n3807;
  assign n3811 = ~n3807 & ~n3808;
  assign n3812 = ~pi29  & ~n3807;
  assign n3813 = ~n38083 & ~n38084;
  assign n3814 = n3252 & ~n3254;
  assign n3815 = ~n3255 & ~n3814;
  assign n3816 = ~n3813 & n3815;
  assign n3817 = n607 & n1596;
  assign n3818 = pi75  & n37489;
  assign n3819 = pi77  & n620;
  assign n3820 = pi76  & n622;
  assign n3821 = ~n3819 & ~n3820;
  assign n3822 = ~n3818 & ~n3820;
  assign n3823 = ~n3819 & n3822;
  assign n3824 = ~n3818 & n3821;
  assign n3825 = ~n3817 & n38085;
  assign n3826 = pi29  & ~n3825;
  assign n3827 = pi29  & ~n3826;
  assign n3828 = pi29  & n3825;
  assign n3829 = ~n3825 & ~n3826;
  assign n3830 = ~pi29  & ~n3825;
  assign n3831 = ~n38086 & ~n38087;
  assign n3832 = n3246 & ~n3248;
  assign n3833 = ~n3246 & ~n37970;
  assign n3834 = ~n3247 & n3252;
  assign n3835 = ~n3833 & ~n3834;
  assign n3836 = ~n37970 & ~n3832;
  assign n3837 = ~n3831 & ~n38088;
  assign n3838 = n3237 & n37969;
  assign n3839 = ~n3245 & ~n3838;
  assign n3840 = n607 & n1465;
  assign n3841 = pi74  & n37489;
  assign n3842 = pi76  & n620;
  assign n3843 = pi75  & n622;
  assign n3844 = ~n3842 & ~n3843;
  assign n3845 = ~n3841 & ~n3843;
  assign n3846 = ~n3842 & n3845;
  assign n3847 = ~n3841 & n3844;
  assign n3848 = ~n3840 & n38089;
  assign n3849 = pi29  & ~n3848;
  assign n3850 = pi29  & ~n3849;
  assign n3851 = pi29  & n3848;
  assign n3852 = ~n3848 & ~n3849;
  assign n3853 = ~pi29  & ~n3848;
  assign n3854 = ~n38090 & ~n38091;
  assign n3855 = n3839 & ~n3854;
  assign n3856 = ~n3839 & n3854;
  assign n3857 = ~n3855 & ~n3856;
  assign n3858 = n607 & n720;
  assign n3859 = pi73  & n37489;
  assign n3860 = pi75  & n620;
  assign n3861 = pi74  & n622;
  assign n3862 = ~n3860 & ~n3861;
  assign n3863 = ~n3859 & ~n3861;
  assign n3864 = ~n3860 & n3863;
  assign n3865 = ~n3859 & n3862;
  assign n3866 = ~n3858 & n38092;
  assign n3867 = pi29  & ~n3866;
  assign n3868 = pi29  & ~n3867;
  assign n3869 = pi29  & n3866;
  assign n3870 = ~n3866 & ~n3867;
  assign n3871 = ~pi29  & ~n3866;
  assign n3872 = ~n38093 & ~n38094;
  assign n3873 = n3233 & ~n3235;
  assign n3874 = ~n3236 & ~n3873;
  assign n3875 = ~n3872 & n3874;
  assign n3876 = n607 & n1218;
  assign n3877 = pi72  & n37489;
  assign n3878 = pi74  & n620;
  assign n3879 = pi73  & n622;
  assign n3880 = ~n3878 & ~n3879;
  assign n3881 = ~n3877 & ~n3879;
  assign n3882 = ~n3878 & n3881;
  assign n3883 = ~n3877 & n3880;
  assign n3884 = ~n3876 & n38095;
  assign n3885 = pi29  & ~n3884;
  assign n3886 = pi29  & ~n3885;
  assign n3887 = pi29  & n3884;
  assign n3888 = ~n3884 & ~n3885;
  assign n3889 = ~pi29  & ~n3884;
  assign n3890 = ~n38096 & ~n38097;
  assign n3891 = n3229 & ~n3231;
  assign n3892 = ~n3232 & ~n3891;
  assign n3893 = ~n3890 & n3892;
  assign n3894 = n607 & n1238;
  assign n3895 = pi71  & n37489;
  assign n3896 = pi73  & n620;
  assign n3897 = pi72  & n622;
  assign n3898 = ~n3896 & ~n3897;
  assign n3899 = ~n3895 & ~n3897;
  assign n3900 = ~n3896 & n3899;
  assign n3901 = ~n3895 & n3898;
  assign n3902 = ~n3894 & n38098;
  assign n3903 = pi29  & ~n3902;
  assign n3904 = pi29  & ~n3903;
  assign n3905 = pi29  & n3902;
  assign n3906 = ~n3902 & ~n3903;
  assign n3907 = ~pi29  & ~n3902;
  assign n3908 = ~n38099 & ~n38100;
  assign n3909 = n3220 & n37966;
  assign n3910 = ~n3220 & n37966;
  assign n3911 = n3220 & ~n37966;
  assign n3912 = ~n3910 & ~n3911;
  assign n3913 = ~n3228 & ~n3909;
  assign n3914 = ~n3908 & ~n38101;
  assign n3915 = n607 & n1124;
  assign n3916 = pi70  & n37489;
  assign n3917 = pi72  & n620;
  assign n3918 = pi71  & n622;
  assign n3919 = ~n3917 & ~n3918;
  assign n3920 = ~n3916 & ~n3918;
  assign n3921 = ~n3917 & n3920;
  assign n3922 = ~n3916 & n3919;
  assign n3923 = ~n3915 & n38102;
  assign n3924 = pi29  & ~n3923;
  assign n3925 = pi29  & ~n3924;
  assign n3926 = pi29  & n3923;
  assign n3927 = ~n3923 & ~n3924;
  assign n3928 = ~pi29  & ~n3923;
  assign n3929 = ~n38103 & ~n38104;
  assign n3930 = n3214 & ~n3216;
  assign n3931 = ~n3214 & ~n37963;
  assign n3932 = ~n3215 & n3220;
  assign n3933 = ~n3931 & ~n3932;
  assign n3934 = ~n37963 & ~n3930;
  assign n3935 = ~n3929 & ~n38105;
  assign n3936 = n607 & n927;
  assign n3937 = pi69  & n37489;
  assign n3938 = pi71  & n620;
  assign n3939 = pi70  & n622;
  assign n3940 = ~n3938 & ~n3939;
  assign n3941 = ~n3937 & ~n3939;
  assign n3942 = ~n3938 & n3941;
  assign n3943 = ~n3937 & n3940;
  assign n3944 = ~n3936 & n38106;
  assign n3945 = pi29  & ~n3944;
  assign n3946 = pi29  & ~n3945;
  assign n3947 = pi29  & n3944;
  assign n3948 = ~n3944 & ~n3945;
  assign n3949 = ~pi29  & ~n3944;
  assign n3950 = ~n38107 & ~n38108;
  assign n3951 = n3210 & ~n3212;
  assign n3952 = ~n3213 & ~n3951;
  assign n3953 = ~n3950 & n3952;
  assign n3954 = n3203 & n37962;
  assign n3955 = ~n3209 & ~n3954;
  assign n3956 = n607 & n972;
  assign n3957 = pi68  & n37489;
  assign n3958 = pi70  & n620;
  assign n3959 = pi69  & n622;
  assign n3960 = ~n3958 & ~n3959;
  assign n3961 = ~n3957 & ~n3959;
  assign n3962 = ~n3958 & n3961;
  assign n3963 = ~n3957 & n3960;
  assign n3964 = ~n3956 & n38109;
  assign n3965 = pi29  & ~n3964;
  assign n3966 = pi29  & ~n3965;
  assign n3967 = pi29  & n3964;
  assign n3968 = ~n3964 & ~n3965;
  assign n3969 = ~pi29  & ~n3964;
  assign n3970 = ~n38110 & ~n38111;
  assign n3971 = n3955 & ~n3970;
  assign n3972 = n607 & n990;
  assign n3973 = pi67  & n37489;
  assign n3974 = pi69  & n620;
  assign n3975 = pi68  & n622;
  assign n3976 = ~n3974 & ~n3975;
  assign n3977 = ~n3973 & ~n3975;
  assign n3978 = ~n3974 & n3977;
  assign n3979 = ~n3973 & n3976;
  assign n3980 = ~n3972 & n38112;
  assign n3981 = pi29  & ~n3980;
  assign n3982 = pi29  & ~n3981;
  assign n3983 = pi29  & n3980;
  assign n3984 = ~n3980 & ~n3981;
  assign n3985 = ~pi29  & ~n3980;
  assign n3986 = ~n38113 & ~n38114;
  assign n3987 = pi32  & ~n37954;
  assign n3988 = n37957 & ~n3987;
  assign n3989 = ~n37957 & n3987;
  assign n3990 = ~n37954 & n3185;
  assign n3991 = ~n37958 & ~n3990;
  assign n3992 = ~n3988 & ~n3989;
  assign n3993 = ~n3986 & n38115;
  assign n3994 = n607 & n871;
  assign n3995 = pi66  & n37489;
  assign n3996 = pi68  & n620;
  assign n3997 = pi67  & n622;
  assign n3998 = ~n3996 & ~n3997;
  assign n3999 = ~n3995 & ~n3997;
  assign n4000 = ~n3996 & n3999;
  assign n4001 = ~n3995 & n3998;
  assign n4002 = ~n3994 & n38116;
  assign n4003 = pi29  & ~n4002;
  assign n4004 = pi29  & ~n4003;
  assign n4005 = pi29  & n4002;
  assign n4006 = ~n4002 & ~n4003;
  assign n4007 = ~pi29  & ~n4002;
  assign n4008 = ~n38117 & ~n38118;
  assign n4009 = pi32  & n3159;
  assign n4010 = ~n3158 & n4009;
  assign n4011 = n3158 & ~n4009;
  assign n4012 = ~n3160 & n3164;
  assign n4013 = ~n37954 & ~n4012;
  assign n4014 = ~n4010 & ~n4011;
  assign n4015 = ~n4008 & n38119;
  assign n4016 = n607 & n37515;
  assign n4017 = pi65  & n620;
  assign n4018 = pi64  & n622;
  assign n4019 = ~n4017 & ~n4018;
  assign n4020 = ~n4016 & n4019;
  assign n4021 = pi64  & n37486;
  assign n4022 = pi29  & ~n4021;
  assign n4023 = pi29  & ~n4020;
  assign n4024 = pi29  & ~n4023;
  assign n4025 = ~n4020 & ~n4023;
  assign n4026 = ~n4024 & ~n4025;
  assign n4027 = n4022 & ~n4026;
  assign n4028 = n4020 & n4022;
  assign n4029 = pi64  & n37489;
  assign n4030 = pi65  & n622;
  assign n4031 = n607 & ~n37521;
  assign n4032 = pi66  & n620;
  assign n4033 = ~n4031 & ~n4032;
  assign n4034 = ~n4030 & ~n4031;
  assign n4035 = ~n4032 & n4034;
  assign n4036 = ~n4030 & ~n4032;
  assign n4037 = ~n4031 & n4036;
  assign n4038 = ~n4030 & n4033;
  assign n4039 = ~n4029 & ~n4030;
  assign n4040 = ~n4032 & n4039;
  assign n4041 = ~n4029 & n4036;
  assign n4042 = ~n4031 & n38122;
  assign n4043 = ~n4029 & n38121;
  assign n4044 = pi29  & ~n38123;
  assign n4045 = pi29  & ~n4044;
  assign n4046 = ~n38123 & ~n4044;
  assign n4047 = ~n4045 & ~n4046;
  assign n4048 = n38120 & ~n4047;
  assign n4049 = n38120 & n38123;
  assign n4050 = n3159 & n38124;
  assign n4051 = n607 & n847;
  assign n4052 = pi65  & n37489;
  assign n4053 = pi67  & n620;
  assign n4054 = pi66  & n622;
  assign n4055 = ~n4053 & ~n4054;
  assign n4056 = ~n4052 & ~n4054;
  assign n4057 = ~n4053 & n4056;
  assign n4058 = ~n4052 & n4055;
  assign n4059 = ~n4051 & n38125;
  assign n4060 = pi29  & ~n4059;
  assign n4061 = pi29  & ~n4060;
  assign n4062 = pi29  & n4059;
  assign n4063 = ~n4059 & ~n4060;
  assign n4064 = ~pi29  & ~n4059;
  assign n4065 = ~n38126 & ~n38127;
  assign n4066 = ~n3159 & ~n38124;
  assign n4067 = n3159 & ~n38124;
  assign n4068 = ~n3159 & n38124;
  assign n4069 = ~n4067 & ~n4068;
  assign n4070 = ~n4050 & ~n4066;
  assign n4071 = ~n4065 & ~n38128;
  assign n4072 = ~n4050 & ~n4071;
  assign n4073 = n4008 & ~n38119;
  assign n4074 = n4008 & n38119;
  assign n4075 = ~n4008 & ~n38119;
  assign n4076 = ~n4074 & ~n4075;
  assign n4077 = ~n4015 & ~n4073;
  assign n4078 = ~n4072 & ~n38129;
  assign n4079 = ~n4015 & ~n4078;
  assign n4080 = n3986 & ~n38115;
  assign n4081 = ~n3993 & ~n4080;
  assign n4082 = ~n4079 & ~n4080;
  assign n4083 = ~n3993 & n4082;
  assign n4084 = ~n4079 & n4081;
  assign n4085 = ~n3993 & ~n38130;
  assign n4086 = ~n3955 & n3970;
  assign n4087 = n3955 & ~n3971;
  assign n4088 = n3955 & n3970;
  assign n4089 = ~n3970 & ~n3971;
  assign n4090 = ~n3955 & ~n3970;
  assign n4091 = ~n38131 & ~n38132;
  assign n4092 = ~n3971 & ~n4086;
  assign n4093 = ~n4085 & ~n38133;
  assign n4094 = ~n3971 & ~n4093;
  assign n4095 = n3950 & ~n3952;
  assign n4096 = ~n3953 & ~n4095;
  assign n4097 = ~n4094 & n4096;
  assign n4098 = ~n3953 & ~n4097;
  assign n4099 = n3929 & n38105;
  assign n4100 = ~n38105 & ~n3935;
  assign n4101 = n3929 & ~n38105;
  assign n4102 = ~n3929 & ~n3935;
  assign n4103 = ~n3929 & n38105;
  assign n4104 = ~n38134 & ~n38135;
  assign n4105 = ~n3935 & ~n4099;
  assign n4106 = ~n4098 & ~n38136;
  assign n4107 = ~n3935 & ~n4106;
  assign n4108 = n3908 & n38101;
  assign n4109 = ~n3914 & ~n4108;
  assign n4110 = ~n4107 & n4109;
  assign n4111 = ~n3914 & ~n4110;
  assign n4112 = n3890 & ~n3892;
  assign n4113 = ~n3893 & ~n4112;
  assign n4114 = ~n4111 & n4113;
  assign n4115 = ~n3893 & ~n4114;
  assign n4116 = n3872 & ~n3874;
  assign n4117 = ~n3872 & ~n3875;
  assign n4118 = ~n3872 & ~n3874;
  assign n4119 = n3874 & ~n3875;
  assign n4120 = n3872 & n3874;
  assign n4121 = ~n38137 & ~n38138;
  assign n4122 = ~n3875 & ~n4116;
  assign n4123 = ~n4115 & ~n38139;
  assign n4124 = ~n3875 & ~n4123;
  assign n4125 = n3857 & ~n4124;
  assign n4126 = ~n3855 & ~n4125;
  assign n4127 = n3831 & n38088;
  assign n4128 = ~n3837 & ~n4127;
  assign n4129 = ~n4126 & n4128;
  assign n4130 = ~n3837 & ~n4129;
  assign n4131 = n3813 & ~n3815;
  assign n4132 = ~n3816 & ~n4131;
  assign n4133 = ~n4130 & n4132;
  assign n4134 = ~n3816 & ~n4133;
  assign n4135 = n3792 & n38081;
  assign n4136 = ~n38081 & ~n3798;
  assign n4137 = n3792 & ~n38081;
  assign n4138 = ~n3792 & ~n3798;
  assign n4139 = ~n3792 & n38081;
  assign n4140 = ~n38140 & ~n38141;
  assign n4141 = ~n3798 & ~n4135;
  assign n4142 = ~n4134 & ~n38142;
  assign n4143 = ~n3798 & ~n4142;
  assign n4144 = ~n3761 & n3776;
  assign n4145 = n3761 & ~n3777;
  assign n4146 = n3761 & n3776;
  assign n4147 = ~n3776 & ~n3777;
  assign n4148 = ~n3761 & ~n3776;
  assign n4149 = ~n38143 & ~n38144;
  assign n4150 = ~n3777 & ~n4144;
  assign n4151 = ~n4143 & ~n38145;
  assign n4152 = ~n3777 & ~n4151;
  assign n4153 = n3756 & ~n3758;
  assign n4154 = ~n3759 & ~n4153;
  assign n4155 = ~n4152 & n4154;
  assign n4156 = ~n3759 & ~n4155;
  assign n4157 = n3735 & n38071;
  assign n4158 = ~n3741 & ~n4157;
  assign n4159 = ~n4156 & n4158;
  assign n4160 = ~n3741 & ~n4159;
  assign n4161 = ~n3704 & n3719;
  assign n4162 = n3704 & ~n3720;
  assign n4163 = n3704 & n3719;
  assign n4164 = ~n3719 & ~n3720;
  assign n4165 = ~n3704 & ~n3719;
  assign n4166 = ~n38146 & ~n38147;
  assign n4167 = ~n3720 & ~n4161;
  assign n4168 = ~n4160 & ~n38148;
  assign n4169 = ~n3720 & ~n4168;
  assign n4170 = n3694 & n38064;
  assign n4171 = ~n38064 & ~n3702;
  assign n4172 = ~n3694 & ~n3702;
  assign n4173 = ~n4171 & ~n4172;
  assign n4174 = ~n3702 & ~n4170;
  assign n4175 = ~n4169 & ~n38149;
  assign n4176 = ~n3702 & ~n4175;
  assign n4177 = ~n3663 & n3678;
  assign n4178 = n3663 & ~n3679;
  assign n4179 = n3663 & n3678;
  assign n4180 = ~n3678 & ~n3679;
  assign n4181 = ~n3663 & ~n3678;
  assign n4182 = ~n38150 & ~n38151;
  assign n4183 = ~n3679 & ~n4177;
  assign n4184 = ~n4176 & ~n38152;
  assign n4185 = ~n3679 & ~n4184;
  assign n4186 = ~n3645 & n3660;
  assign n4187 = n3645 & ~n3661;
  assign n4188 = n3645 & n3660;
  assign n4189 = ~n3660 & ~n3661;
  assign n4190 = ~n3645 & ~n3660;
  assign n4191 = ~n38153 & ~n38154;
  assign n4192 = ~n3661 & ~n4186;
  assign n4193 = ~n4185 & ~n38155;
  assign n4194 = ~n3661 & ~n4193;
  assign n4195 = ~n3627 & n3642;
  assign n4196 = ~n3643 & ~n4195;
  assign n4197 = ~n4194 & ~n4195;
  assign n4198 = ~n3643 & n4197;
  assign n4199 = ~n4194 & n4196;
  assign n4200 = ~n3643 & ~n38156;
  assign n4201 = ~n3609 & n3624;
  assign n4202 = ~n3625 & ~n4201;
  assign n4203 = ~n4200 & n4202;
  assign n4204 = ~n3625 & ~n4203;
  assign n4205 = ~n3589 & n3606;
  assign n4206 = n3589 & ~n3607;
  assign n4207 = n3589 & n3606;
  assign n4208 = ~n3606 & ~n3607;
  assign n4209 = ~n3589 & ~n3606;
  assign n4210 = ~n38157 & ~n38158;
  assign n4211 = ~n3607 & ~n4205;
  assign n4212 = ~n4204 & ~n38159;
  assign n4213 = ~n3607 & ~n4212;
  assign n4214 = n3581 & n38043;
  assign n4215 = ~n3587 & ~n4214;
  assign n4216 = ~n4213 & n4215;
  assign n4217 = ~n3587 & ~n4216;
  assign n4218 = n634 & ~n3563;
  assign n4219 = ~n3564 & ~n4218;
  assign n4220 = ~n4217 & n4219;
  assign n4221 = ~n3564 & ~n4220;
  assign n4222 = ~n3558 & ~n3561;
  assign n4223 = ~n3552 & ~n3555;
  assign n4224 = n2104 & n2779;
  assign n4225 = pi84  & n37758;
  assign n4226 = pi86  & n2117;
  assign n4227 = pi85  & n2119;
  assign n4228 = ~n4226 & ~n4227;
  assign n4229 = ~n4225 & ~n4227;
  assign n4230 = ~n4226 & n4229;
  assign n4231 = ~n4225 & n4228;
  assign n4232 = ~n4224 & n38160;
  assign n4233 = pi35  & ~n4232;
  assign n4234 = pi35  & ~n4233;
  assign n4235 = pi35  & n4232;
  assign n4236 = ~n4232 & ~n4233;
  assign n4237 = ~pi35  & ~n4232;
  assign n4238 = ~n38161 & ~n38162;
  assign n4239 = ~n3539 & ~n3547;
  assign n4240 = ~n3533 & ~n3536;
  assign n4241 = ~n3520 & ~n3528;
  assign n4242 = n940 & n1596;
  assign n4243 = pi75  & n37541;
  assign n4244 = pi77  & n953;
  assign n4245 = pi76  & n955;
  assign n4246 = ~n4244 & ~n4245;
  assign n4247 = ~n4243 & ~n4245;
  assign n4248 = ~n4244 & n4247;
  assign n4249 = ~n4243 & n4246;
  assign n4250 = ~n4242 & n38163;
  assign n4251 = pi44  & ~n4250;
  assign n4252 = pi44  & ~n4251;
  assign n4253 = pi44  & n4250;
  assign n4254 = ~n4250 & ~n4251;
  assign n4255 = ~pi44  & ~n4250;
  assign n4256 = ~n38164 & ~n38165;
  assign n4257 = ~n3507 & ~n3515;
  assign n4258 = n785 & n1218;
  assign n4259 = pi72  & n37520;
  assign n4260 = pi74  & n787;
  assign n4261 = pi73  & n795;
  assign n4262 = ~n4260 & ~n4261;
  assign n4263 = ~n4259 & ~n4261;
  assign n4264 = ~n4260 & n4263;
  assign n4265 = ~n4259 & n4262;
  assign n4266 = ~n4258 & n38166;
  assign n4267 = pi47  & ~n4266;
  assign n4268 = pi47  & ~n4267;
  assign n4269 = pi47  & n4266;
  assign n4270 = ~n4266 & ~n4267;
  assign n4271 = ~pi47  & ~n4266;
  assign n4272 = ~n38167 & ~n38168;
  assign n4273 = ~n3496 & ~n3504;
  assign n4274 = n894 & n927;
  assign n4275 = pi69  & n37580;
  assign n4276 = pi71  & n896;
  assign n4277 = pi70  & n904;
  assign n4278 = ~n4276 & ~n4277;
  assign n4279 = ~n4275 & ~n4277;
  assign n4280 = ~n4276 & n4279;
  assign n4281 = ~n4275 & n4278;
  assign n4282 = ~n4274 & n38169;
  assign n4283 = pi50  & ~n4282;
  assign n4284 = pi50  & ~n4283;
  assign n4285 = pi50  & n4282;
  assign n4286 = ~n4282 & ~n4283;
  assign n4287 = ~pi50  & ~n4282;
  assign n4288 = ~n38170 & ~n38171;
  assign n4289 = ~n3472 & ~n3478;
  assign n4290 = n871 & n1971;
  assign n4291 = pi66  & n37864;
  assign n4292 = pi68  & n1973;
  assign n4293 = pi67  & n1981;
  assign n4294 = ~n4292 & ~n4293;
  assign n4295 = ~n4291 & ~n4293;
  assign n4296 = ~n4292 & n4295;
  assign n4297 = ~n4291 & n4294;
  assign n4298 = ~n4290 & n38172;
  assign n4299 = pi53  & ~n4298;
  assign n4300 = pi53  & ~n4299;
  assign n4301 = pi53  & n4298;
  assign n4302 = ~n4298 & ~n4299;
  assign n4303 = ~pi53  & ~n4298;
  assign n4304 = ~n38173 & ~n38174;
  assign n4305 = pi56  & n3471;
  assign n4306 = pi55  & ~pi56 ;
  assign n4307 = ~pi55  & pi56 ;
  assign n4308 = ~pi55  & ~pi56 ;
  assign n4309 = pi55  & pi56 ;
  assign n4310 = ~n4308 & ~n4309;
  assign n4311 = ~n4306 & ~n4307;
  assign n4312 = n38020 & n38175;
  assign n4313 = n37515 & n4312;
  assign n4314 = n38020 & ~n38175;
  assign n4315 = pi65  & n4314;
  assign n4316 = pi54  & ~pi55 ;
  assign n4317 = ~pi54  & pi55 ;
  assign n4318 = ~pi54  & ~pi55 ;
  assign n4319 = pi54  & pi55 ;
  assign n4320 = ~n4318 & ~n4319;
  assign n4321 = ~n4316 & ~n4317;
  assign n4322 = ~n38020 & n38176;
  assign n4323 = pi64  & n4322;
  assign n4324 = ~n4315 & ~n4323;
  assign n4325 = ~n4313 & n4324;
  assign n4326 = n4305 & ~n4325;
  assign n4327 = ~n4305 & n4325;
  assign n4328 = pi56  & ~n3471;
  assign n4329 = pi56  & ~n4325;
  assign n4330 = pi56  & ~n4329;
  assign n4331 = ~n4325 & ~n4329;
  assign n4332 = ~n4330 & ~n4331;
  assign n4333 = n4328 & ~n4332;
  assign n4334 = n4325 & n4328;
  assign n4335 = ~n4328 & n4332;
  assign n4336 = ~n38177 & ~n4335;
  assign n4337 = ~n4326 & ~n4327;
  assign n4338 = n4304 & ~n38178;
  assign n4339 = ~n4304 & n38178;
  assign n4340 = ~n4338 & ~n4339;
  assign n4341 = ~n4289 & n4340;
  assign n4342 = n4289 & ~n4340;
  assign n4343 = ~n4341 & ~n4342;
  assign n4344 = n4288 & ~n4343;
  assign n4345 = ~n4288 & n4343;
  assign n4346 = ~n4344 & ~n4345;
  assign n4347 = ~n4273 & n4346;
  assign n4348 = n4273 & ~n4346;
  assign n4349 = ~n4347 & ~n4348;
  assign n4350 = n4272 & ~n4349;
  assign n4351 = ~n4272 & n4349;
  assign n4352 = ~n4350 & ~n4351;
  assign n4353 = ~n4257 & n4352;
  assign n4354 = n4257 & ~n4352;
  assign n4355 = ~n4353 & ~n4354;
  assign n4356 = n4256 & ~n4355;
  assign n4357 = ~n4256 & n4355;
  assign n4358 = ~n4356 & ~n4357;
  assign n4359 = ~n4241 & n4358;
  assign n4360 = n4241 & ~n4358;
  assign n4361 = ~n4359 & ~n4360;
  assign n4362 = n733 & n2063;
  assign n4363 = pi78  & n37510;
  assign n4364 = pi80  & n746;
  assign n4365 = pi79  & n748;
  assign n4366 = ~n4364 & ~n4365;
  assign n4367 = ~n4363 & ~n4365;
  assign n4368 = ~n4364 & n4367;
  assign n4369 = ~n4363 & n4366;
  assign n4370 = ~n4362 & n38179;
  assign n4371 = pi41  & ~n4370;
  assign n4372 = pi41  & ~n4371;
  assign n4373 = pi41  & n4370;
  assign n4374 = ~n4370 & ~n4371;
  assign n4375 = ~pi41  & ~n4370;
  assign n4376 = ~n38180 & ~n38181;
  assign n4377 = n4361 & ~n4376;
  assign n4378 = ~n4361 & n4376;
  assign n4379 = n4361 & ~n4377;
  assign n4380 = n4361 & n4376;
  assign n4381 = ~n4376 & ~n4377;
  assign n4382 = ~n4361 & ~n4376;
  assign n4383 = ~n38182 & ~n38183;
  assign n4384 = ~n4377 & ~n4378;
  assign n4385 = n4240 & n38184;
  assign n4386 = ~n4240 & ~n38184;
  assign n4387 = ~n4385 & ~n4386;
  assign n4388 = n691 & n2091;
  assign n4389 = pi81  & n37503;
  assign n4390 = pi83  & n704;
  assign n4391 = pi82  & n706;
  assign n4392 = ~n4390 & ~n4391;
  assign n4393 = ~n4389 & ~n4391;
  assign n4394 = ~n4390 & n4393;
  assign n4395 = ~n4389 & n4392;
  assign n4396 = ~n4388 & n38185;
  assign n4397 = pi38  & ~n4396;
  assign n4398 = pi38  & ~n4397;
  assign n4399 = pi38  & n4396;
  assign n4400 = ~n4396 & ~n4397;
  assign n4401 = ~pi38  & ~n4396;
  assign n4402 = ~n38186 & ~n38187;
  assign n4403 = n4387 & ~n4402;
  assign n4404 = ~n4387 & n4402;
  assign n4405 = ~n4403 & ~n4404;
  assign n4406 = ~n4239 & ~n4404;
  assign n4407 = ~n4403 & n4406;
  assign n4408 = ~n4239 & n4405;
  assign n4409 = n4239 & ~n4405;
  assign n4410 = ~n4239 & ~n38188;
  assign n4411 = ~n4403 & ~n38188;
  assign n4412 = ~n4404 & n4411;
  assign n4413 = ~n4410 & ~n4412;
  assign n4414 = ~n38188 & ~n4409;
  assign n4415 = ~n4238 & ~n38189;
  assign n4416 = n4238 & n38189;
  assign n4417 = ~n38189 & ~n4415;
  assign n4418 = n4238 & ~n38189;
  assign n4419 = ~n4238 & ~n4415;
  assign n4420 = ~n4238 & n38189;
  assign n4421 = ~n38190 & ~n38191;
  assign n4422 = ~n4415 & ~n4416;
  assign n4423 = n4223 & n38192;
  assign n4424 = ~n4223 & ~n38192;
  assign n4425 = ~n4423 & ~n4424;
  assign n4426 = n649 & n3591;
  assign n4427 = pi87  & n37496;
  assign n4428 = pi89  & n662;
  assign n4429 = pi88  & n664;
  assign n4430 = ~n4428 & ~n4429;
  assign n4431 = ~n4427 & ~n4429;
  assign n4432 = ~n4428 & n4431;
  assign n4433 = ~n4427 & n4430;
  assign n4434 = ~n4426 & n38193;
  assign n4435 = pi32  & ~n4434;
  assign n4436 = pi32  & ~n4435;
  assign n4437 = pi32  & n4434;
  assign n4438 = ~n4434 & ~n4435;
  assign n4439 = ~pi32  & ~n4434;
  assign n4440 = ~n38194 & ~n38195;
  assign n4441 = n4425 & ~n4440;
  assign n4442 = ~n4425 & n4440;
  assign n4443 = n4425 & ~n4441;
  assign n4444 = n4425 & n4440;
  assign n4445 = ~n4440 & ~n4441;
  assign n4446 = ~n4425 & ~n4440;
  assign n4447 = ~n38196 & ~n38197;
  assign n4448 = ~n4441 & ~n4442;
  assign n4449 = n4222 & n38198;
  assign n4450 = ~n4222 & ~n38198;
  assign n4451 = ~n4449 & ~n4450;
  assign n4452 = n425 & ~n427;
  assign n4453 = ~n428 & ~n4452;
  assign n4454 = n607 & n4453;
  assign n4455 = pi90  & n37489;
  assign n4456 = pi92  & n620;
  assign n4457 = pi91  & n622;
  assign n4458 = ~n4456 & ~n4457;
  assign n4459 = ~n4455 & ~n4457;
  assign n4460 = ~n4456 & n4459;
  assign n4461 = ~n4455 & n4458;
  assign n4462 = ~n4454 & n38199;
  assign n4463 = pi29  & ~n4462;
  assign n4464 = pi29  & ~n4463;
  assign n4465 = pi29  & n4462;
  assign n4466 = ~n4462 & ~n4463;
  assign n4467 = ~pi29  & ~n4462;
  assign n4468 = ~n38200 & ~n38201;
  assign n4469 = n4451 & ~n4468;
  assign n4470 = ~n4451 & n4468;
  assign n4471 = n4451 & ~n4469;
  assign n4472 = n4451 & n4468;
  assign n4473 = ~n4468 & ~n4469;
  assign n4474 = ~n4451 & ~n4468;
  assign n4475 = ~n38202 & ~n38203;
  assign n4476 = ~n4469 & ~n4470;
  assign n4477 = n4221 & n38204;
  assign n4478 = ~n4221 & ~n38204;
  assign n4479 = ~n4477 & ~n4478;
  assign n4480 = pi23  & ~pi24 ;
  assign n4481 = ~pi23  & pi24 ;
  assign n4482 = ~pi23  & ~pi24 ;
  assign n4483 = pi23  & pi24 ;
  assign n4484 = ~n4482 & ~n4483;
  assign n4485 = ~n4480 & ~n4481;
  assign n4486 = pi25  & ~pi26 ;
  assign n4487 = ~pi25  & pi26 ;
  assign n4488 = ~pi25  & ~pi26 ;
  assign n4489 = pi25  & pi26 ;
  assign n4490 = ~n4488 & ~n4489;
  assign n4491 = ~n4486 & ~n4487;
  assign n4492 = n38205 & n38206;
  assign n4493 = n437 & ~n439;
  assign n4494 = ~n440 & ~n4493;
  assign n4495 = n4492 & n4494;
  assign n4496 = pi24  & ~pi25 ;
  assign n4497 = ~pi24  & pi25 ;
  assign n4498 = ~pi24  & ~pi25 ;
  assign n4499 = pi24  & pi25 ;
  assign n4500 = ~n4498 & ~n4499;
  assign n4501 = ~n4496 & ~n4497;
  assign n4502 = ~n38205 & n38206;
  assign n4503 = ~n38205 & ~n38207;
  assign n4504 = n38206 & n4503;
  assign n4505 = ~n38207 & n4502;
  assign n4506 = pi93  & n38208;
  assign n4507 = n38205 & ~n38206;
  assign n4508 = pi95  & n4507;
  assign n4509 = ~n38205 & n38207;
  assign n4510 = pi94  & n4509;
  assign n4511 = ~n4508 & ~n4510;
  assign n4512 = ~n4506 & ~n4510;
  assign n4513 = ~n4508 & n4512;
  assign n4514 = ~n4506 & n4511;
  assign n4515 = ~n4495 & n38209;
  assign n4516 = pi26  & ~n4515;
  assign n4517 = pi26  & ~n4516;
  assign n4518 = pi26  & n4515;
  assign n4519 = ~n4515 & ~n4516;
  assign n4520 = ~pi26  & ~n4515;
  assign n4521 = ~n38210 & ~n38211;
  assign n4522 = n4479 & ~n4521;
  assign n4523 = n433 & ~n435;
  assign n4524 = ~n436 & ~n4523;
  assign n4525 = n4492 & n4524;
  assign n4526 = pi92  & n38208;
  assign n4527 = pi94  & n4507;
  assign n4528 = pi93  & n4509;
  assign n4529 = ~n4527 & ~n4528;
  assign n4530 = ~n4526 & ~n4528;
  assign n4531 = ~n4527 & n4530;
  assign n4532 = ~n4526 & n4529;
  assign n4533 = ~n4525 & n38212;
  assign n4534 = pi26  & ~n4533;
  assign n4535 = pi26  & ~n4534;
  assign n4536 = pi26  & n4533;
  assign n4537 = ~n4533 & ~n4534;
  assign n4538 = ~pi26  & ~n4533;
  assign n4539 = ~n38213 & ~n38214;
  assign n4540 = n4217 & ~n4219;
  assign n4541 = ~n4220 & ~n4540;
  assign n4542 = ~n4539 & n4541;
  assign n4543 = n429 & ~n431;
  assign n4544 = ~n432 & ~n4543;
  assign n4545 = n4492 & n4544;
  assign n4546 = pi91  & n38208;
  assign n4547 = pi93  & n4507;
  assign n4548 = pi92  & n4509;
  assign n4549 = ~n4547 & ~n4548;
  assign n4550 = ~n4546 & ~n4548;
  assign n4551 = ~n4547 & n4550;
  assign n4552 = ~n4546 & n4549;
  assign n4553 = ~n4545 & n38215;
  assign n4554 = pi26  & ~n4553;
  assign n4555 = pi26  & ~n4554;
  assign n4556 = pi26  & n4553;
  assign n4557 = ~n4553 & ~n4554;
  assign n4558 = ~pi26  & ~n4553;
  assign n4559 = ~n38216 & ~n38217;
  assign n4560 = n4213 & ~n4215;
  assign n4561 = ~n4216 & ~n4560;
  assign n4562 = ~n4559 & n4561;
  assign n4563 = n4453 & n4492;
  assign n4564 = pi90  & n38208;
  assign n4565 = pi92  & n4507;
  assign n4566 = pi91  & n4509;
  assign n4567 = ~n4565 & ~n4566;
  assign n4568 = ~n4564 & ~n4566;
  assign n4569 = ~n4565 & n4568;
  assign n4570 = ~n4564 & n4567;
  assign n4571 = ~n4563 & n38218;
  assign n4572 = pi26  & ~n4571;
  assign n4573 = pi26  & ~n4572;
  assign n4574 = pi26  & n4571;
  assign n4575 = ~n4571 & ~n4572;
  assign n4576 = ~pi26  & ~n4571;
  assign n4577 = ~n38219 & ~n38220;
  assign n4578 = n4204 & n38159;
  assign n4579 = ~n4204 & n38159;
  assign n4580 = n4204 & ~n38159;
  assign n4581 = ~n4579 & ~n4580;
  assign n4582 = ~n4212 & ~n4578;
  assign n4583 = ~n4577 & ~n38221;
  assign n4584 = n4200 & ~n4202;
  assign n4585 = ~n4203 & ~n4584;
  assign n4586 = n594 & n4492;
  assign n4587 = pi89  & n38208;
  assign n4588 = pi91  & n4507;
  assign n4589 = pi90  & n4509;
  assign n4590 = ~n4588 & ~n4589;
  assign n4591 = ~n4587 & ~n4589;
  assign n4592 = ~n4588 & n4591;
  assign n4593 = ~n4587 & n4590;
  assign n4594 = ~n4586 & n38222;
  assign n4595 = pi26  & ~n4594;
  assign n4596 = pi26  & ~n4595;
  assign n4597 = pi26  & n4594;
  assign n4598 = ~n4594 & ~n4595;
  assign n4599 = ~pi26  & ~n4594;
  assign n4600 = ~n38223 & ~n38224;
  assign n4601 = n4585 & ~n4600;
  assign n4602 = n3566 & n4492;
  assign n4603 = pi88  & n38208;
  assign n4604 = pi90  & n4507;
  assign n4605 = pi89  & n4509;
  assign n4606 = ~n4604 & ~n4605;
  assign n4607 = ~n4603 & ~n4605;
  assign n4608 = ~n4604 & n4607;
  assign n4609 = ~n4603 & n4606;
  assign n4610 = ~n4602 & n38225;
  assign n4611 = pi26  & ~n4610;
  assign n4612 = pi26  & ~n4611;
  assign n4613 = pi26  & n4610;
  assign n4614 = ~n4610 & ~n4611;
  assign n4615 = ~pi26  & ~n4610;
  assign n4616 = ~n38226 & ~n38227;
  assign n4617 = n4194 & ~n4196;
  assign n4618 = ~n4194 & ~n38156;
  assign n4619 = ~n4195 & n4200;
  assign n4620 = ~n4618 & ~n4619;
  assign n4621 = ~n38156 & ~n4617;
  assign n4622 = ~n4616 & ~n38228;
  assign n4623 = n4185 & n38155;
  assign n4624 = ~n4193 & ~n4623;
  assign n4625 = n3591 & n4492;
  assign n4626 = pi87  & n38208;
  assign n4627 = pi89  & n4507;
  assign n4628 = pi88  & n4509;
  assign n4629 = ~n4627 & ~n4628;
  assign n4630 = ~n4626 & ~n4628;
  assign n4631 = ~n4627 & n4630;
  assign n4632 = ~n4626 & n4629;
  assign n4633 = ~n4625 & n38229;
  assign n4634 = pi26  & ~n4633;
  assign n4635 = pi26  & ~n4634;
  assign n4636 = pi26  & n4633;
  assign n4637 = ~n4633 & ~n4634;
  assign n4638 = ~pi26  & ~n4633;
  assign n4639 = ~n38230 & ~n38231;
  assign n4640 = n4624 & ~n4639;
  assign n4641 = n4176 & n38152;
  assign n4642 = ~n4184 & ~n4641;
  assign n4643 = n3354 & n4492;
  assign n4644 = pi86  & n38208;
  assign n4645 = pi88  & n4507;
  assign n4646 = pi87  & n4509;
  assign n4647 = ~n4645 & ~n4646;
  assign n4648 = ~n4644 & ~n4646;
  assign n4649 = ~n4645 & n4648;
  assign n4650 = ~n4644 & n4647;
  assign n4651 = ~n4643 & n38232;
  assign n4652 = pi26  & ~n4651;
  assign n4653 = pi26  & ~n4652;
  assign n4654 = pi26  & n4651;
  assign n4655 = ~n4651 & ~n4652;
  assign n4656 = ~pi26  & ~n4651;
  assign n4657 = ~n38233 & ~n38234;
  assign n4658 = n4642 & ~n4657;
  assign n4659 = n4169 & n38149;
  assign n4660 = ~n4175 & ~n4659;
  assign n4661 = n636 & n4492;
  assign n4662 = pi85  & n38208;
  assign n4663 = pi87  & n4507;
  assign n4664 = pi86  & n4509;
  assign n4665 = ~n4663 & ~n4664;
  assign n4666 = ~n4662 & ~n4664;
  assign n4667 = ~n4663 & n4666;
  assign n4668 = ~n4662 & n4665;
  assign n4669 = ~n4661 & n38235;
  assign n4670 = pi26  & ~n4669;
  assign n4671 = pi26  & ~n4670;
  assign n4672 = pi26  & n4669;
  assign n4673 = ~n4669 & ~n4670;
  assign n4674 = ~pi26  & ~n4669;
  assign n4675 = ~n38236 & ~n38237;
  assign n4676 = n4660 & ~n4675;
  assign n4677 = n4160 & n38148;
  assign n4678 = ~n4168 & ~n4677;
  assign n4679 = n2779 & n4492;
  assign n4680 = pi84  & n38208;
  assign n4681 = pi86  & n4507;
  assign n4682 = pi85  & n4509;
  assign n4683 = ~n4681 & ~n4682;
  assign n4684 = ~n4680 & ~n4682;
  assign n4685 = ~n4681 & n4684;
  assign n4686 = ~n4680 & n4683;
  assign n4687 = ~n4679 & n38238;
  assign n4688 = pi26  & ~n4687;
  assign n4689 = pi26  & ~n4688;
  assign n4690 = pi26  & n4687;
  assign n4691 = ~n4687 & ~n4688;
  assign n4692 = ~pi26  & ~n4687;
  assign n4693 = ~n38239 & ~n38240;
  assign n4694 = n4678 & ~n4693;
  assign n4695 = n4156 & ~n4158;
  assign n4696 = ~n4159 & ~n4695;
  assign n4697 = n2804 & n4492;
  assign n4698 = pi83  & n38208;
  assign n4699 = pi85  & n4507;
  assign n4700 = pi84  & n4509;
  assign n4701 = ~n4699 & ~n4700;
  assign n4702 = ~n4698 & ~n4700;
  assign n4703 = ~n4699 & n4702;
  assign n4704 = ~n4698 & n4701;
  assign n4705 = ~n4697 & n38241;
  assign n4706 = pi26  & ~n4705;
  assign n4707 = pi26  & ~n4706;
  assign n4708 = pi26  & n4705;
  assign n4709 = ~n4705 & ~n4706;
  assign n4710 = ~pi26  & ~n4705;
  assign n4711 = ~n38242 & ~n38243;
  assign n4712 = n4696 & ~n4711;
  assign n4713 = n4152 & ~n4154;
  assign n4714 = ~n4155 & ~n4713;
  assign n4715 = n2591 & n4492;
  assign n4716 = pi82  & n38208;
  assign n4717 = pi84  & n4507;
  assign n4718 = pi83  & n4509;
  assign n4719 = ~n4717 & ~n4718;
  assign n4720 = ~n4716 & ~n4718;
  assign n4721 = ~n4717 & n4720;
  assign n4722 = ~n4716 & n4719;
  assign n4723 = ~n4715 & n38244;
  assign n4724 = pi26  & ~n4723;
  assign n4725 = pi26  & ~n4724;
  assign n4726 = pi26  & n4723;
  assign n4727 = ~n4723 & ~n4724;
  assign n4728 = ~pi26  & ~n4723;
  assign n4729 = ~n38245 & ~n38246;
  assign n4730 = n4714 & ~n4729;
  assign n4731 = n4143 & n38145;
  assign n4732 = ~n4151 & ~n4731;
  assign n4733 = n2091 & n4492;
  assign n4734 = pi81  & n38208;
  assign n4735 = pi83  & n4507;
  assign n4736 = pi82  & n4509;
  assign n4737 = ~n4735 & ~n4736;
  assign n4738 = ~n4734 & ~n4736;
  assign n4739 = ~n4735 & n4738;
  assign n4740 = ~n4734 & n4737;
  assign n4741 = ~n4733 & n38247;
  assign n4742 = pi26  & ~n4741;
  assign n4743 = pi26  & ~n4742;
  assign n4744 = pi26  & n4741;
  assign n4745 = ~n4741 & ~n4742;
  assign n4746 = ~pi26  & ~n4741;
  assign n4747 = ~n38248 & ~n38249;
  assign n4748 = n4732 & ~n4747;
  assign n4749 = n2134 & n4492;
  assign n4750 = pi80  & n38208;
  assign n4751 = pi82  & n4507;
  assign n4752 = pi81  & n4509;
  assign n4753 = ~n4751 & ~n4752;
  assign n4754 = ~n4750 & ~n4752;
  assign n4755 = ~n4751 & n4754;
  assign n4756 = ~n4750 & n4753;
  assign n4757 = ~n4749 & n38250;
  assign n4758 = pi26  & ~n4757;
  assign n4759 = pi26  & ~n4758;
  assign n4760 = pi26  & n4757;
  assign n4761 = ~n4757 & ~n4758;
  assign n4762 = ~pi26  & ~n4757;
  assign n4763 = ~n38251 & ~n38252;
  assign n4764 = n4134 & n38142;
  assign n4765 = ~n4134 & n38142;
  assign n4766 = n4134 & ~n38142;
  assign n4767 = ~n4765 & ~n4766;
  assign n4768 = ~n4142 & ~n4764;
  assign n4769 = ~n4763 & ~n38253;
  assign n4770 = n2154 & n4492;
  assign n4771 = pi79  & n38208;
  assign n4772 = pi81  & n4507;
  assign n4773 = pi80  & n4509;
  assign n4774 = ~n4772 & ~n4773;
  assign n4775 = ~n4771 & ~n4773;
  assign n4776 = ~n4772 & n4775;
  assign n4777 = ~n4771 & n4774;
  assign n4778 = ~n4770 & n38254;
  assign n4779 = pi26  & ~n4778;
  assign n4780 = pi26  & ~n4779;
  assign n4781 = pi26  & n4778;
  assign n4782 = ~n4778 & ~n4779;
  assign n4783 = ~pi26  & ~n4778;
  assign n4784 = ~n38255 & ~n38256;
  assign n4785 = n4130 & ~n4132;
  assign n4786 = ~n4133 & ~n4785;
  assign n4787 = ~n4784 & n4786;
  assign n4788 = n4126 & ~n4128;
  assign n4789 = ~n4129 & ~n4788;
  assign n4790 = n2063 & n4492;
  assign n4791 = pi78  & n38208;
  assign n4792 = pi80  & n4507;
  assign n4793 = pi79  & n4509;
  assign n4794 = ~n4792 & ~n4793;
  assign n4795 = ~n4791 & ~n4793;
  assign n4796 = ~n4792 & n4795;
  assign n4797 = ~n4791 & n4794;
  assign n4798 = ~n4790 & n38257;
  assign n4799 = pi26  & ~n4798;
  assign n4800 = pi26  & ~n4799;
  assign n4801 = pi26  & n4798;
  assign n4802 = ~n4798 & ~n4799;
  assign n4803 = ~pi26  & ~n4798;
  assign n4804 = ~n38258 & ~n38259;
  assign n4805 = n4789 & ~n4804;
  assign n4806 = ~n3857 & n4124;
  assign n4807 = ~n4125 & ~n4806;
  assign n4808 = n678 & n4492;
  assign n4809 = pi77  & n38208;
  assign n4810 = pi79  & n4507;
  assign n4811 = pi78  & n4509;
  assign n4812 = ~n4810 & ~n4811;
  assign n4813 = ~n4809 & ~n4811;
  assign n4814 = ~n4810 & n4813;
  assign n4815 = ~n4809 & n4812;
  assign n4816 = ~n4808 & n38260;
  assign n4817 = pi26  & ~n4816;
  assign n4818 = pi26  & ~n4817;
  assign n4819 = pi26  & n4816;
  assign n4820 = ~n4816 & ~n4817;
  assign n4821 = ~pi26  & ~n4816;
  assign n4822 = ~n38261 & ~n38262;
  assign n4823 = n4807 & ~n4822;
  assign n4824 = n1578 & n4492;
  assign n4825 = pi76  & n38208;
  assign n4826 = pi78  & n4507;
  assign n4827 = pi77  & n4509;
  assign n4828 = ~n4826 & ~n4827;
  assign n4829 = ~n4825 & ~n4827;
  assign n4830 = ~n4826 & n4829;
  assign n4831 = ~n4825 & n4828;
  assign n4832 = ~n4824 & n38263;
  assign n4833 = pi26  & ~n4832;
  assign n4834 = pi26  & ~n4833;
  assign n4835 = pi26  & n4832;
  assign n4836 = ~n4832 & ~n4833;
  assign n4837 = ~pi26  & ~n4832;
  assign n4838 = ~n38264 & ~n38265;
  assign n4839 = n4115 & n38139;
  assign n4840 = ~n4115 & ~n4123;
  assign n4841 = ~n38139 & ~n4123;
  assign n4842 = ~n4840 & ~n4841;
  assign n4843 = ~n4123 & ~n4839;
  assign n4844 = ~n4838 & ~n38266;
  assign n4845 = n1596 & n4492;
  assign n4846 = pi75  & n38208;
  assign n4847 = pi77  & n4507;
  assign n4848 = pi76  & n4509;
  assign n4849 = ~n4847 & ~n4848;
  assign n4850 = ~n4846 & ~n4848;
  assign n4851 = ~n4847 & n4850;
  assign n4852 = ~n4846 & n4849;
  assign n4853 = ~n4845 & n38267;
  assign n4854 = pi26  & ~n4853;
  assign n4855 = pi26  & ~n4854;
  assign n4856 = pi26  & n4853;
  assign n4857 = ~n4853 & ~n4854;
  assign n4858 = ~pi26  & ~n4853;
  assign n4859 = ~n38268 & ~n38269;
  assign n4860 = n4111 & ~n4113;
  assign n4861 = ~n4114 & ~n4860;
  assign n4862 = ~n4859 & n4861;
  assign n4863 = n4107 & ~n4109;
  assign n4864 = ~n4110 & ~n4863;
  assign n4865 = n1465 & n4492;
  assign n4866 = pi74  & n38208;
  assign n4867 = pi76  & n4507;
  assign n4868 = pi75  & n4509;
  assign n4869 = ~n4867 & ~n4868;
  assign n4870 = ~n4866 & ~n4868;
  assign n4871 = ~n4867 & n4870;
  assign n4872 = ~n4866 & n4869;
  assign n4873 = ~n4865 & n38270;
  assign n4874 = pi26  & ~n4873;
  assign n4875 = pi26  & ~n4874;
  assign n4876 = pi26  & n4873;
  assign n4877 = ~n4873 & ~n4874;
  assign n4878 = ~pi26  & ~n4873;
  assign n4879 = ~n38271 & ~n38272;
  assign n4880 = n4864 & ~n4879;
  assign n4881 = ~n4864 & n4879;
  assign n4882 = ~n4880 & ~n4881;
  assign n4883 = n720 & n4492;
  assign n4884 = pi73  & n38208;
  assign n4885 = pi75  & n4507;
  assign n4886 = pi74  & n4509;
  assign n4887 = ~n4885 & ~n4886;
  assign n4888 = ~n4884 & ~n4886;
  assign n4889 = ~n4885 & n4888;
  assign n4890 = ~n4884 & n4887;
  assign n4891 = ~n4883 & n38273;
  assign n4892 = pi26  & ~n4891;
  assign n4893 = pi26  & ~n4892;
  assign n4894 = pi26  & n4891;
  assign n4895 = ~n4891 & ~n4892;
  assign n4896 = ~pi26  & ~n4891;
  assign n4897 = ~n38274 & ~n38275;
  assign n4898 = n4098 & n38136;
  assign n4899 = ~n4106 & ~n4898;
  assign n4900 = ~n4897 & n4899;
  assign n4901 = n4094 & ~n4096;
  assign n4902 = ~n4097 & ~n4901;
  assign n4903 = n1218 & n4492;
  assign n4904 = pi72  & n38208;
  assign n4905 = pi74  & n4507;
  assign n4906 = pi73  & n4509;
  assign n4907 = ~n4905 & ~n4906;
  assign n4908 = ~n4904 & ~n4906;
  assign n4909 = ~n4905 & n4908;
  assign n4910 = ~n4904 & n4907;
  assign n4911 = ~n4903 & n38276;
  assign n4912 = pi26  & ~n4911;
  assign n4913 = pi26  & ~n4912;
  assign n4914 = pi26  & n4911;
  assign n4915 = ~n4911 & ~n4912;
  assign n4916 = ~pi26  & ~n4911;
  assign n4917 = ~n38277 & ~n38278;
  assign n4918 = n4902 & ~n4917;
  assign n4919 = n1238 & n4492;
  assign n4920 = pi71  & n38208;
  assign n4921 = pi73  & n4507;
  assign n4922 = pi72  & n4509;
  assign n4923 = ~n4921 & ~n4922;
  assign n4924 = ~n4920 & ~n4922;
  assign n4925 = ~n4921 & n4924;
  assign n4926 = ~n4920 & n4923;
  assign n4927 = ~n4919 & n38279;
  assign n4928 = pi26  & ~n4927;
  assign n4929 = pi26  & ~n4928;
  assign n4930 = pi26  & n4927;
  assign n4931 = ~n4927 & ~n4928;
  assign n4932 = ~pi26  & ~n4927;
  assign n4933 = ~n38280 & ~n38281;
  assign n4934 = n4085 & n38133;
  assign n4935 = ~n4085 & n38133;
  assign n4936 = n4085 & ~n38133;
  assign n4937 = ~n4935 & ~n4936;
  assign n4938 = ~n4093 & ~n4934;
  assign n4939 = ~n4933 & ~n38282;
  assign n4940 = n1124 & n4492;
  assign n4941 = pi70  & n38208;
  assign n4942 = pi72  & n4507;
  assign n4943 = pi71  & n4509;
  assign n4944 = ~n4942 & ~n4943;
  assign n4945 = ~n4941 & ~n4943;
  assign n4946 = ~n4942 & n4945;
  assign n4947 = ~n4941 & n4944;
  assign n4948 = ~n4940 & n38283;
  assign n4949 = pi26  & ~n4948;
  assign n4950 = pi26  & ~n4949;
  assign n4951 = pi26  & n4948;
  assign n4952 = ~n4948 & ~n4949;
  assign n4953 = ~pi26  & ~n4948;
  assign n4954 = ~n38284 & ~n38285;
  assign n4955 = n4079 & ~n4081;
  assign n4956 = ~n4079 & ~n38130;
  assign n4957 = ~n4080 & n4085;
  assign n4958 = ~n4956 & ~n4957;
  assign n4959 = ~n38130 & ~n4955;
  assign n4960 = ~n4954 & ~n38286;
  assign n4961 = n927 & n4492;
  assign n4962 = pi69  & n38208;
  assign n4963 = pi71  & n4507;
  assign n4964 = pi70  & n4509;
  assign n4965 = ~n4963 & ~n4964;
  assign n4966 = ~n4962 & ~n4964;
  assign n4967 = ~n4963 & n4966;
  assign n4968 = ~n4962 & n4965;
  assign n4969 = ~n4961 & n38287;
  assign n4970 = pi26  & ~n4969;
  assign n4971 = pi26  & ~n4970;
  assign n4972 = pi26  & n4969;
  assign n4973 = ~n4969 & ~n4970;
  assign n4974 = ~pi26  & ~n4969;
  assign n4975 = ~n38288 & ~n38289;
  assign n4976 = n4072 & n38129;
  assign n4977 = ~n4078 & ~n4976;
  assign n4978 = ~n4975 & n4977;
  assign n4979 = n4065 & n38128;
  assign n4980 = ~n4071 & ~n4979;
  assign n4981 = n972 & n4492;
  assign n4982 = pi68  & n38208;
  assign n4983 = pi70  & n4507;
  assign n4984 = pi69  & n4509;
  assign n4985 = ~n4983 & ~n4984;
  assign n4986 = ~n4982 & ~n4984;
  assign n4987 = ~n4983 & n4986;
  assign n4988 = ~n4982 & n4985;
  assign n4989 = ~n4981 & n38290;
  assign n4990 = pi26  & ~n4989;
  assign n4991 = pi26  & ~n4990;
  assign n4992 = pi26  & n4989;
  assign n4993 = ~n4989 & ~n4990;
  assign n4994 = ~pi26  & ~n4989;
  assign n4995 = ~n38291 & ~n38292;
  assign n4996 = n4980 & ~n4995;
  assign n4997 = n990 & n4492;
  assign n4998 = pi67  & n38208;
  assign n4999 = pi69  & n4507;
  assign n5000 = pi68  & n4509;
  assign n5001 = ~n4999 & ~n5000;
  assign n5002 = ~n4998 & ~n5000;
  assign n5003 = ~n4999 & n5002;
  assign n5004 = ~n4998 & n5001;
  assign n5005 = ~n4997 & n38293;
  assign n5006 = pi26  & ~n5005;
  assign n5007 = pi26  & ~n5006;
  assign n5008 = pi26  & n5005;
  assign n5009 = ~n5005 & ~n5006;
  assign n5010 = ~pi26  & ~n5005;
  assign n5011 = ~n38294 & ~n38295;
  assign n5012 = pi29  & ~n38120;
  assign n5013 = n38123 & ~n5012;
  assign n5014 = ~n38123 & n5012;
  assign n5015 = ~n38120 & n4047;
  assign n5016 = ~n38124 & ~n5015;
  assign n5017 = ~n5013 & ~n5014;
  assign n5018 = ~n5011 & n38296;
  assign n5019 = n871 & n4492;
  assign n5020 = pi66  & n38208;
  assign n5021 = pi68  & n4507;
  assign n5022 = pi67  & n4509;
  assign n5023 = ~n5021 & ~n5022;
  assign n5024 = ~n5020 & ~n5022;
  assign n5025 = ~n5021 & n5024;
  assign n5026 = ~n5020 & n5023;
  assign n5027 = ~n5019 & n38297;
  assign n5028 = pi26  & ~n5027;
  assign n5029 = pi26  & ~n5028;
  assign n5030 = pi26  & n5027;
  assign n5031 = ~n5027 & ~n5028;
  assign n5032 = ~pi26  & ~n5027;
  assign n5033 = ~n38298 & ~n38299;
  assign n5034 = pi29  & n4021;
  assign n5035 = ~n4020 & n5034;
  assign n5036 = n4020 & ~n5034;
  assign n5037 = ~n4022 & n4026;
  assign n5038 = ~n38120 & ~n5037;
  assign n5039 = ~n5035 & ~n5036;
  assign n5040 = ~n5033 & n38300;
  assign n5041 = n37515 & n4492;
  assign n5042 = pi65  & n4507;
  assign n5043 = pi64  & n4509;
  assign n5044 = ~n5042 & ~n5043;
  assign n5045 = ~n5041 & n5044;
  assign n5046 = pi64  & n38205;
  assign n5047 = pi26  & ~n5046;
  assign n5048 = pi26  & ~n5045;
  assign n5049 = pi26  & ~n5048;
  assign n5050 = ~n5045 & ~n5048;
  assign n5051 = ~n5049 & ~n5050;
  assign n5052 = n5047 & ~n5051;
  assign n5053 = n5045 & n5047;
  assign n5054 = pi64  & n38208;
  assign n5055 = pi65  & n4509;
  assign n5056 = ~n37521 & n4492;
  assign n5057 = pi66  & n4507;
  assign n5058 = ~n5056 & ~n5057;
  assign n5059 = ~n5055 & ~n5056;
  assign n5060 = ~n5057 & n5059;
  assign n5061 = ~n5055 & ~n5057;
  assign n5062 = ~n5056 & n5061;
  assign n5063 = ~n5055 & n5058;
  assign n5064 = ~n5054 & ~n5055;
  assign n5065 = ~n5057 & n5064;
  assign n5066 = ~n5054 & n5061;
  assign n5067 = ~n5056 & n38303;
  assign n5068 = ~n5054 & n38302;
  assign n5069 = pi26  & ~n38304;
  assign n5070 = pi26  & ~n5069;
  assign n5071 = ~n38304 & ~n5069;
  assign n5072 = ~n5070 & ~n5071;
  assign n5073 = n38301 & ~n5072;
  assign n5074 = n38301 & n38304;
  assign n5075 = n4021 & n38305;
  assign n5076 = n847 & n4492;
  assign n5077 = pi65  & n38208;
  assign n5078 = pi67  & n4507;
  assign n5079 = pi66  & n4509;
  assign n5080 = ~n5078 & ~n5079;
  assign n5081 = ~n5077 & ~n5079;
  assign n5082 = ~n5078 & n5081;
  assign n5083 = ~n5077 & n5080;
  assign n5084 = ~n5076 & n38306;
  assign n5085 = pi26  & ~n5084;
  assign n5086 = pi26  & ~n5085;
  assign n5087 = pi26  & n5084;
  assign n5088 = ~n5084 & ~n5085;
  assign n5089 = ~pi26  & ~n5084;
  assign n5090 = ~n38307 & ~n38308;
  assign n5091 = ~n4021 & ~n38305;
  assign n5092 = n4021 & ~n38305;
  assign n5093 = ~n4021 & n38305;
  assign n5094 = ~n5092 & ~n5093;
  assign n5095 = ~n5075 & ~n5091;
  assign n5096 = ~n5090 & ~n38309;
  assign n5097 = ~n5075 & ~n5096;
  assign n5098 = n5033 & ~n38300;
  assign n5099 = n5033 & n38300;
  assign n5100 = ~n5033 & ~n38300;
  assign n5101 = ~n5099 & ~n5100;
  assign n5102 = ~n5040 & ~n5098;
  assign n5103 = ~n5097 & ~n38310;
  assign n5104 = ~n5040 & ~n5103;
  assign n5105 = n5011 & ~n38296;
  assign n5106 = ~n5018 & ~n5105;
  assign n5107 = ~n5104 & ~n5105;
  assign n5108 = ~n5018 & n5107;
  assign n5109 = ~n5104 & n5106;
  assign n5110 = ~n5018 & ~n38311;
  assign n5111 = ~n4980 & n4995;
  assign n5112 = n4980 & ~n4996;
  assign n5113 = n4980 & n4995;
  assign n5114 = ~n4995 & ~n4996;
  assign n5115 = ~n4980 & ~n4995;
  assign n5116 = ~n38312 & ~n38313;
  assign n5117 = ~n4996 & ~n5111;
  assign n5118 = ~n5110 & ~n38314;
  assign n5119 = ~n4996 & ~n5118;
  assign n5120 = n4975 & ~n4977;
  assign n5121 = ~n4978 & ~n5120;
  assign n5122 = ~n5119 & n5121;
  assign n5123 = ~n4978 & ~n5122;
  assign n5124 = n4954 & n38286;
  assign n5125 = ~n38286 & ~n4960;
  assign n5126 = n4954 & ~n38286;
  assign n5127 = ~n4954 & ~n4960;
  assign n5128 = ~n4954 & n38286;
  assign n5129 = ~n38315 & ~n38316;
  assign n5130 = ~n4960 & ~n5124;
  assign n5131 = ~n5123 & ~n38317;
  assign n5132 = ~n4960 & ~n5131;
  assign n5133 = n4933 & n38282;
  assign n5134 = ~n4939 & ~n5133;
  assign n5135 = ~n5132 & n5134;
  assign n5136 = ~n4939 & ~n5135;
  assign n5137 = ~n4902 & n4917;
  assign n5138 = n4902 & ~n4918;
  assign n5139 = n4902 & n4917;
  assign n5140 = ~n4917 & ~n4918;
  assign n5141 = ~n4902 & ~n4917;
  assign n5142 = ~n38318 & ~n38319;
  assign n5143 = ~n4918 & ~n5137;
  assign n5144 = ~n5136 & ~n38320;
  assign n5145 = ~n4918 & ~n5144;
  assign n5146 = n4897 & ~n4899;
  assign n5147 = ~n4897 & ~n4900;
  assign n5148 = ~n4897 & ~n4899;
  assign n5149 = n4899 & ~n4900;
  assign n5150 = n4897 & n4899;
  assign n5151 = ~n38321 & ~n38322;
  assign n5152 = ~n4900 & ~n5146;
  assign n5153 = ~n5145 & ~n38323;
  assign n5154 = ~n4900 & ~n5153;
  assign n5155 = n4882 & ~n5154;
  assign n5156 = ~n4880 & ~n5155;
  assign n5157 = n4859 & ~n4861;
  assign n5158 = ~n4862 & ~n5157;
  assign n5159 = ~n5156 & n5158;
  assign n5160 = ~n4862 & ~n5159;
  assign n5161 = n4838 & n38266;
  assign n5162 = ~n4844 & ~n5161;
  assign n5163 = ~n5160 & n5162;
  assign n5164 = ~n4844 & ~n5163;
  assign n5165 = ~n4807 & n4822;
  assign n5166 = n4807 & ~n4823;
  assign n5167 = n4807 & n4822;
  assign n5168 = ~n4822 & ~n4823;
  assign n5169 = ~n4807 & ~n4822;
  assign n5170 = ~n38324 & ~n38325;
  assign n5171 = ~n4823 & ~n5165;
  assign n5172 = ~n5164 & ~n38326;
  assign n5173 = ~n4823 & ~n5172;
  assign n5174 = ~n4789 & n4804;
  assign n5175 = n4789 & ~n4805;
  assign n5176 = n4789 & n4804;
  assign n5177 = ~n4804 & ~n4805;
  assign n5178 = ~n4789 & ~n4804;
  assign n5179 = ~n38327 & ~n38328;
  assign n5180 = ~n4805 & ~n5174;
  assign n5181 = ~n5173 & ~n38329;
  assign n5182 = ~n4805 & ~n5181;
  assign n5183 = n4784 & ~n4786;
  assign n5184 = ~n4787 & ~n5183;
  assign n5185 = ~n5182 & n5184;
  assign n5186 = ~n4787 & ~n5185;
  assign n5187 = n4763 & n38253;
  assign n5188 = ~n4769 & ~n5187;
  assign n5189 = ~n5186 & n5188;
  assign n5190 = ~n4769 & ~n5189;
  assign n5191 = ~n4732 & n4747;
  assign n5192 = n4732 & ~n4748;
  assign n5193 = n4732 & n4747;
  assign n5194 = ~n4747 & ~n4748;
  assign n5195 = ~n4732 & ~n4747;
  assign n5196 = ~n38330 & ~n38331;
  assign n5197 = ~n4748 & ~n5191;
  assign n5198 = ~n5190 & ~n38332;
  assign n5199 = ~n4748 & ~n5198;
  assign n5200 = ~n4714 & n4729;
  assign n5201 = n4714 & ~n4730;
  assign n5202 = n4714 & n4729;
  assign n5203 = ~n4729 & ~n4730;
  assign n5204 = ~n4714 & ~n4729;
  assign n5205 = ~n38333 & ~n38334;
  assign n5206 = ~n4730 & ~n5200;
  assign n5207 = ~n5199 & ~n38335;
  assign n5208 = ~n4730 & ~n5207;
  assign n5209 = ~n4696 & n4711;
  assign n5210 = n4696 & ~n4712;
  assign n5211 = n4696 & n4711;
  assign n5212 = ~n4711 & ~n4712;
  assign n5213 = ~n4696 & ~n4711;
  assign n5214 = ~n38336 & ~n38337;
  assign n5215 = ~n4712 & ~n5209;
  assign n5216 = ~n5208 & ~n38338;
  assign n5217 = ~n4712 & ~n5216;
  assign n5218 = ~n4678 & n4693;
  assign n5219 = n4678 & ~n4694;
  assign n5220 = n4678 & n4693;
  assign n5221 = ~n4693 & ~n4694;
  assign n5222 = ~n4678 & ~n4693;
  assign n5223 = ~n38339 & ~n38340;
  assign n5224 = ~n4694 & ~n5218;
  assign n5225 = ~n5217 & ~n38341;
  assign n5226 = ~n4694 & ~n5225;
  assign n5227 = ~n4660 & n4675;
  assign n5228 = ~n4676 & ~n5227;
  assign n5229 = ~n5226 & ~n5227;
  assign n5230 = ~n4676 & n5229;
  assign n5231 = ~n5226 & n5228;
  assign n5232 = ~n4676 & ~n38342;
  assign n5233 = ~n4642 & n4657;
  assign n5234 = ~n4658 & ~n5233;
  assign n5235 = ~n5232 & n5234;
  assign n5236 = ~n4658 & ~n5235;
  assign n5237 = ~n4624 & n4639;
  assign n5238 = n4624 & ~n4640;
  assign n5239 = n4624 & n4639;
  assign n5240 = ~n4639 & ~n4640;
  assign n5241 = ~n4624 & ~n4639;
  assign n5242 = ~n38343 & ~n38344;
  assign n5243 = ~n4640 & ~n5237;
  assign n5244 = ~n5236 & ~n38345;
  assign n5245 = ~n4640 & ~n5244;
  assign n5246 = n4616 & n38228;
  assign n5247 = ~n4622 & ~n5246;
  assign n5248 = ~n5245 & n5247;
  assign n5249 = ~n4622 & ~n5248;
  assign n5250 = ~n4585 & n4600;
  assign n5251 = n4585 & ~n4601;
  assign n5252 = n4585 & n4600;
  assign n5253 = ~n4600 & ~n4601;
  assign n5254 = ~n4585 & ~n4600;
  assign n5255 = ~n38346 & ~n38347;
  assign n5256 = ~n4601 & ~n5250;
  assign n5257 = ~n5249 & ~n38348;
  assign n5258 = ~n4601 & ~n5257;
  assign n5259 = n4577 & n38221;
  assign n5260 = ~n4583 & ~n5259;
  assign n5261 = ~n5258 & n5260;
  assign n5262 = ~n4583 & ~n5261;
  assign n5263 = n4559 & ~n4561;
  assign n5264 = ~n4562 & ~n5263;
  assign n5265 = ~n5262 & n5264;
  assign n5266 = ~n4562 & ~n5265;
  assign n5267 = n4539 & ~n4541;
  assign n5268 = ~n4542 & ~n5267;
  assign n5269 = ~n5266 & n5268;
  assign n5270 = ~n4542 & ~n5269;
  assign n5271 = ~n4479 & n4521;
  assign n5272 = n4479 & ~n4522;
  assign n5273 = n4479 & n4521;
  assign n5274 = ~n4521 & ~n4522;
  assign n5275 = ~n4479 & ~n4521;
  assign n5276 = ~n38349 & ~n38350;
  assign n5277 = ~n4522 & ~n5271;
  assign n5278 = ~n5270 & ~n38351;
  assign n5279 = ~n4522 & ~n5278;
  assign n5280 = n441 & ~n443;
  assign n5281 = ~n444 & ~n5280;
  assign n5282 = n4492 & n5281;
  assign n5283 = pi94  & n38208;
  assign n5284 = pi96  & n4507;
  assign n5285 = pi95  & n4509;
  assign n5286 = ~n5284 & ~n5285;
  assign n5287 = ~n5283 & ~n5285;
  assign n5288 = ~n5284 & n5287;
  assign n5289 = ~n5283 & n5286;
  assign n5290 = ~n5282 & n38352;
  assign n5291 = pi26  & ~n5290;
  assign n5292 = pi26  & ~n5291;
  assign n5293 = pi26  & n5290;
  assign n5294 = ~n5290 & ~n5291;
  assign n5295 = ~pi26  & ~n5290;
  assign n5296 = ~n38353 & ~n38354;
  assign n5297 = ~n4469 & ~n4478;
  assign n5298 = n607 & n4544;
  assign n5299 = pi91  & n37489;
  assign n5300 = pi93  & n620;
  assign n5301 = pi92  & n622;
  assign n5302 = ~n5300 & ~n5301;
  assign n5303 = ~n5299 & ~n5301;
  assign n5304 = ~n5300 & n5303;
  assign n5305 = ~n5299 & n5302;
  assign n5306 = ~n5298 & n38355;
  assign n5307 = pi29  & ~n5306;
  assign n5308 = pi29  & ~n5307;
  assign n5309 = pi29  & n5306;
  assign n5310 = ~n5306 & ~n5307;
  assign n5311 = ~pi29  & ~n5306;
  assign n5312 = ~n38356 & ~n38357;
  assign n5313 = ~n4441 & ~n4450;
  assign n5314 = ~n4415 & ~n4424;
  assign n5315 = n636 & n2104;
  assign n5316 = pi85  & n37758;
  assign n5317 = pi87  & n2117;
  assign n5318 = pi86  & n2119;
  assign n5319 = ~n5317 & ~n5318;
  assign n5320 = ~n5316 & ~n5318;
  assign n5321 = ~n5317 & n5320;
  assign n5322 = ~n5316 & n5319;
  assign n5323 = ~n5315 & n38358;
  assign n5324 = pi35  & ~n5323;
  assign n5325 = pi35  & ~n5324;
  assign n5326 = pi35  & n5323;
  assign n5327 = ~n5323 & ~n5324;
  assign n5328 = ~pi35  & ~n5323;
  assign n5329 = ~n38359 & ~n38360;
  assign n5330 = n691 & n2591;
  assign n5331 = pi82  & n37503;
  assign n5332 = pi84  & n704;
  assign n5333 = pi83  & n706;
  assign n5334 = ~n5332 & ~n5333;
  assign n5335 = ~n5331 & ~n5333;
  assign n5336 = ~n5332 & n5335;
  assign n5337 = ~n5331 & n5334;
  assign n5338 = ~n5330 & n38361;
  assign n5339 = pi38  & ~n5338;
  assign n5340 = pi38  & ~n5339;
  assign n5341 = pi38  & n5338;
  assign n5342 = ~n5338 & ~n5339;
  assign n5343 = ~pi38  & ~n5338;
  assign n5344 = ~n38362 & ~n38363;
  assign n5345 = ~n4377 & ~n4386;
  assign n5346 = n733 & n2154;
  assign n5347 = pi79  & n37510;
  assign n5348 = pi81  & n746;
  assign n5349 = pi80  & n748;
  assign n5350 = ~n5348 & ~n5349;
  assign n5351 = ~n5347 & ~n5349;
  assign n5352 = ~n5348 & n5351;
  assign n5353 = ~n5347 & n5350;
  assign n5354 = ~n5346 & n38364;
  assign n5355 = pi41  & ~n5354;
  assign n5356 = pi41  & ~n5355;
  assign n5357 = pi41  & n5354;
  assign n5358 = ~n5354 & ~n5355;
  assign n5359 = ~pi41  & ~n5354;
  assign n5360 = ~n38365 & ~n38366;
  assign n5361 = ~n4357 & ~n4359;
  assign n5362 = ~n4351 & ~n4353;
  assign n5363 = n720 & n785;
  assign n5364 = pi73  & n37520;
  assign n5365 = pi75  & n787;
  assign n5366 = pi74  & n795;
  assign n5367 = ~n5365 & ~n5366;
  assign n5368 = ~n5364 & ~n5366;
  assign n5369 = ~n5365 & n5368;
  assign n5370 = ~n5364 & n5367;
  assign n5371 = ~n5363 & n38367;
  assign n5372 = pi47  & ~n5371;
  assign n5373 = pi47  & ~n5372;
  assign n5374 = pi47  & n5371;
  assign n5375 = ~n5371 & ~n5372;
  assign n5376 = ~pi47  & ~n5371;
  assign n5377 = ~n38368 & ~n38369;
  assign n5378 = ~n4345 & ~n4347;
  assign n5379 = n894 & n1124;
  assign n5380 = pi70  & n37580;
  assign n5381 = pi72  & n896;
  assign n5382 = pi71  & n904;
  assign n5383 = ~n5381 & ~n5382;
  assign n5384 = ~n5380 & ~n5382;
  assign n5385 = ~n5381 & n5384;
  assign n5386 = ~n5380 & n5383;
  assign n5387 = ~n5379 & n38370;
  assign n5388 = pi50  & ~n5387;
  assign n5389 = pi50  & ~n5388;
  assign n5390 = pi50  & n5387;
  assign n5391 = ~n5387 & ~n5388;
  assign n5392 = ~pi50  & ~n5387;
  assign n5393 = ~n38371 & ~n38372;
  assign n5394 = ~n4339 & ~n4341;
  assign n5395 = n990 & n1971;
  assign n5396 = pi67  & n37864;
  assign n5397 = pi69  & n1973;
  assign n5398 = pi68  & n1981;
  assign n5399 = ~n5397 & ~n5398;
  assign n5400 = ~n5396 & ~n5398;
  assign n5401 = ~n5397 & n5400;
  assign n5402 = ~n5396 & n5399;
  assign n5403 = ~n5395 & n38373;
  assign n5404 = pi53  & ~n5403;
  assign n5405 = pi53  & ~n5404;
  assign n5406 = pi53  & n5403;
  assign n5407 = ~n5403 & ~n5404;
  assign n5408 = ~pi53  & ~n5403;
  assign n5409 = ~n38374 & ~n38375;
  assign n5410 = pi56  & ~n38177;
  assign n5411 = ~n38020 & n38175;
  assign n5412 = ~n38020 & ~n38176;
  assign n5413 = n38175 & n5412;
  assign n5414 = ~n38176 & n5411;
  assign n5415 = pi64  & n38376;
  assign n5416 = pi65  & n4322;
  assign n5417 = ~n37521 & n4312;
  assign n5418 = pi66  & n4314;
  assign n5419 = ~n5417 & ~n5418;
  assign n5420 = ~n5416 & ~n5417;
  assign n5421 = ~n5418 & n5420;
  assign n5422 = ~n5416 & ~n5418;
  assign n5423 = ~n5417 & n5422;
  assign n5424 = ~n5416 & n5419;
  assign n5425 = ~n5415 & ~n5416;
  assign n5426 = ~n5418 & n5425;
  assign n5427 = ~n5415 & n5422;
  assign n5428 = ~n5417 & n38378;
  assign n5429 = ~n5415 & n38377;
  assign n5430 = ~n5410 & n38379;
  assign n5431 = n5410 & ~n38379;
  assign n5432 = pi56  & ~n38379;
  assign n5433 = pi56  & ~n5432;
  assign n5434 = ~n38379 & ~n5432;
  assign n5435 = ~n5433 & ~n5434;
  assign n5436 = n38177 & ~n5435;
  assign n5437 = n38177 & n38379;
  assign n5438 = ~n38177 & n5435;
  assign n5439 = ~n38380 & ~n5438;
  assign n5440 = ~n5430 & ~n5431;
  assign n5441 = ~n5409 & n38381;
  assign n5442 = n5409 & ~n38381;
  assign n5443 = ~n5441 & ~n5442;
  assign n5444 = ~n5394 & ~n5442;
  assign n5445 = ~n5441 & n5444;
  assign n5446 = ~n5394 & n5443;
  assign n5447 = n5394 & ~n5443;
  assign n5448 = ~n5394 & ~n38382;
  assign n5449 = ~n5441 & ~n38382;
  assign n5450 = ~n5442 & n5449;
  assign n5451 = ~n5448 & ~n5450;
  assign n5452 = ~n38382 & ~n5447;
  assign n5453 = n5393 & n38383;
  assign n5454 = ~n5393 & ~n38383;
  assign n5455 = ~n5453 & ~n5454;
  assign n5456 = ~n5378 & n5455;
  assign n5457 = n5378 & ~n5455;
  assign n5458 = ~n5456 & ~n5457;
  assign n5459 = n5377 & ~n5458;
  assign n5460 = ~n5377 & n5458;
  assign n5461 = ~n5459 & ~n5460;
  assign n5462 = ~n5362 & n5461;
  assign n5463 = n5362 & ~n5461;
  assign n5464 = ~n5462 & ~n5463;
  assign n5465 = n940 & n1578;
  assign n5466 = pi76  & n37541;
  assign n5467 = pi78  & n953;
  assign n5468 = pi77  & n955;
  assign n5469 = ~n5467 & ~n5468;
  assign n5470 = ~n5466 & ~n5468;
  assign n5471 = ~n5467 & n5470;
  assign n5472 = ~n5466 & n5469;
  assign n5473 = ~n5465 & n38384;
  assign n5474 = pi44  & ~n5473;
  assign n5475 = pi44  & ~n5474;
  assign n5476 = pi44  & n5473;
  assign n5477 = ~n5473 & ~n5474;
  assign n5478 = ~pi44  & ~n5473;
  assign n5479 = ~n38385 & ~n38386;
  assign n5480 = n5464 & ~n5479;
  assign n5481 = ~n5464 & n5479;
  assign n5482 = n5464 & ~n5480;
  assign n5483 = n5464 & n5479;
  assign n5484 = ~n5479 & ~n5480;
  assign n5485 = ~n5464 & ~n5479;
  assign n5486 = ~n38387 & ~n38388;
  assign n5487 = ~n5480 & ~n5481;
  assign n5488 = ~n5361 & ~n38389;
  assign n5489 = n5361 & n38389;
  assign n5490 = ~n5488 & ~n5489;
  assign n5491 = ~n5360 & n5490;
  assign n5492 = n5360 & ~n5490;
  assign n5493 = ~n5360 & ~n5491;
  assign n5494 = ~n5360 & ~n5490;
  assign n5495 = n5490 & ~n5491;
  assign n5496 = n5360 & n5490;
  assign n5497 = ~n38390 & ~n38391;
  assign n5498 = ~n5491 & ~n5492;
  assign n5499 = ~n5345 & ~n38392;
  assign n5500 = n5345 & n38392;
  assign n5501 = ~n5345 & ~n5499;
  assign n5502 = ~n5345 & n38392;
  assign n5503 = ~n38392 & ~n5499;
  assign n5504 = n5345 & ~n38392;
  assign n5505 = ~n38393 & ~n38394;
  assign n5506 = ~n5499 & ~n5500;
  assign n5507 = ~n5344 & ~n38395;
  assign n5508 = n5344 & n38395;
  assign n5509 = ~n38395 & ~n5507;
  assign n5510 = ~n5344 & ~n5507;
  assign n5511 = ~n5509 & ~n5510;
  assign n5512 = ~n5507 & ~n5508;
  assign n5513 = ~n4411 & ~n38396;
  assign n5514 = n4411 & n38396;
  assign n5515 = ~n4411 & n38396;
  assign n5516 = n4411 & ~n38396;
  assign n5517 = ~n5515 & ~n5516;
  assign n5518 = ~n5513 & ~n5514;
  assign n5519 = ~n5329 & ~n38397;
  assign n5520 = n5329 & n38397;
  assign n5521 = ~n5519 & ~n5520;
  assign n5522 = n5314 & ~n5521;
  assign n5523 = ~n5314 & n5521;
  assign n5524 = ~n5522 & ~n5523;
  assign n5525 = n649 & n3566;
  assign n5526 = pi88  & n37496;
  assign n5527 = pi90  & n662;
  assign n5528 = pi89  & n664;
  assign n5529 = ~n5527 & ~n5528;
  assign n5530 = ~n5526 & ~n5528;
  assign n5531 = ~n5527 & n5530;
  assign n5532 = ~n5526 & n5529;
  assign n5533 = ~n5525 & n38398;
  assign n5534 = pi32  & ~n5533;
  assign n5535 = pi32  & ~n5534;
  assign n5536 = pi32  & n5533;
  assign n5537 = ~n5533 & ~n5534;
  assign n5538 = ~pi32  & ~n5533;
  assign n5539 = ~n38399 & ~n38400;
  assign n5540 = n5524 & ~n5539;
  assign n5541 = ~n5524 & n5539;
  assign n5542 = ~n5540 & ~n5541;
  assign n5543 = ~n5313 & ~n5541;
  assign n5544 = ~n5540 & n5543;
  assign n5545 = ~n5313 & n5542;
  assign n5546 = n5313 & ~n5542;
  assign n5547 = ~n5313 & ~n38401;
  assign n5548 = ~n5540 & ~n38401;
  assign n5549 = ~n5541 & n5548;
  assign n5550 = ~n5547 & ~n5549;
  assign n5551 = ~n38401 & ~n5546;
  assign n5552 = n5312 & n38402;
  assign n5553 = ~n5312 & ~n38402;
  assign n5554 = ~n5552 & ~n5553;
  assign n5555 = ~n5297 & n5554;
  assign n5556 = n5297 & ~n5554;
  assign n5557 = ~n5555 & ~n5556;
  assign n5558 = n5296 & ~n5557;
  assign n5559 = ~n5296 & n5557;
  assign n5560 = ~n5558 & ~n5559;
  assign n5561 = ~n5279 & n5560;
  assign n5562 = n5279 & ~n5560;
  assign n5563 = ~n5561 & ~n5562;
  assign n5564 = pi20  & ~pi21 ;
  assign n5565 = ~pi20  & pi21 ;
  assign n5566 = ~pi20  & ~pi21 ;
  assign n5567 = pi20  & pi21 ;
  assign n5568 = ~n5566 & ~n5567;
  assign n5569 = ~n5564 & ~n5565;
  assign n5570 = pi22  & ~pi23 ;
  assign n5571 = ~pi22  & pi23 ;
  assign n5572 = ~pi22  & ~pi23 ;
  assign n5573 = pi22  & pi23 ;
  assign n5574 = ~n5572 & ~n5573;
  assign n5575 = ~n5570 & ~n5571;
  assign n5576 = n38403 & n38404;
  assign n5577 = n453 & ~n455;
  assign n5578 = ~n456 & ~n5577;
  assign n5579 = n5576 & n5578;
  assign n5580 = pi21  & ~pi22 ;
  assign n5581 = ~pi21  & pi22 ;
  assign n5582 = ~pi21  & ~pi22 ;
  assign n5583 = pi21  & pi22 ;
  assign n5584 = ~n5582 & ~n5583;
  assign n5585 = ~n5580 & ~n5581;
  assign n5586 = ~n38403 & n38404;
  assign n5587 = ~n38403 & ~n38405;
  assign n5588 = n38404 & n5587;
  assign n5589 = ~n38405 & n5586;
  assign n5590 = pi97  & n38406;
  assign n5591 = n38403 & ~n38404;
  assign n5592 = pi99  & n5591;
  assign n5593 = ~n38403 & n38405;
  assign n5594 = pi98  & n5593;
  assign n5595 = ~n5592 & ~n5594;
  assign n5596 = ~n5590 & ~n5594;
  assign n5597 = ~n5592 & n5596;
  assign n5598 = ~n5590 & n5595;
  assign n5599 = ~n5579 & n38407;
  assign n5600 = pi23  & ~n5599;
  assign n5601 = pi23  & ~n5600;
  assign n5602 = pi23  & n5599;
  assign n5603 = ~n5599 & ~n5600;
  assign n5604 = ~pi23  & ~n5599;
  assign n5605 = ~n38408 & ~n38409;
  assign n5606 = n5563 & ~n5605;
  assign n5607 = n5270 & n38351;
  assign n5608 = ~n5278 & ~n5607;
  assign n5609 = n449 & ~n451;
  assign n5610 = ~n452 & ~n5609;
  assign n5611 = n5576 & n5610;
  assign n5612 = pi96  & n38406;
  assign n5613 = pi98  & n5591;
  assign n5614 = pi97  & n5593;
  assign n5615 = ~n5613 & ~n5614;
  assign n5616 = ~n5612 & ~n5614;
  assign n5617 = ~n5613 & n5616;
  assign n5618 = ~n5612 & n5615;
  assign n5619 = ~n5611 & n38410;
  assign n5620 = pi23  & ~n5619;
  assign n5621 = pi23  & ~n5620;
  assign n5622 = pi23  & n5619;
  assign n5623 = ~n5619 & ~n5620;
  assign n5624 = ~pi23  & ~n5619;
  assign n5625 = ~n38411 & ~n38412;
  assign n5626 = n5608 & ~n5625;
  assign n5627 = n5266 & ~n5268;
  assign n5628 = ~n5269 & ~n5627;
  assign n5629 = n445 & ~n447;
  assign n5630 = ~n448 & ~n5629;
  assign n5631 = n5576 & n5630;
  assign n5632 = pi95  & n38406;
  assign n5633 = pi97  & n5591;
  assign n5634 = pi96  & n5593;
  assign n5635 = ~n5633 & ~n5634;
  assign n5636 = ~n5632 & ~n5634;
  assign n5637 = ~n5633 & n5636;
  assign n5638 = ~n5632 & n5635;
  assign n5639 = ~n5631 & n38413;
  assign n5640 = pi23  & ~n5639;
  assign n5641 = pi23  & ~n5640;
  assign n5642 = pi23  & n5639;
  assign n5643 = ~n5639 & ~n5640;
  assign n5644 = ~pi23  & ~n5639;
  assign n5645 = ~n38414 & ~n38415;
  assign n5646 = n5628 & ~n5645;
  assign n5647 = n5281 & n5576;
  assign n5648 = pi94  & n38406;
  assign n5649 = pi96  & n5591;
  assign n5650 = pi95  & n5593;
  assign n5651 = ~n5649 & ~n5650;
  assign n5652 = ~n5648 & ~n5650;
  assign n5653 = ~n5649 & n5652;
  assign n5654 = ~n5648 & n5651;
  assign n5655 = ~n5647 & n38416;
  assign n5656 = pi23  & ~n5655;
  assign n5657 = pi23  & ~n5656;
  assign n5658 = pi23  & n5655;
  assign n5659 = ~n5655 & ~n5656;
  assign n5660 = ~pi23  & ~n5655;
  assign n5661 = ~n38417 & ~n38418;
  assign n5662 = n5262 & ~n5264;
  assign n5663 = ~n5265 & ~n5662;
  assign n5664 = ~n5661 & n5663;
  assign n5665 = n5258 & ~n5260;
  assign n5666 = ~n5261 & ~n5665;
  assign n5667 = n4494 & n5576;
  assign n5668 = pi93  & n38406;
  assign n5669 = pi95  & n5591;
  assign n5670 = pi94  & n5593;
  assign n5671 = ~n5669 & ~n5670;
  assign n5672 = ~n5668 & ~n5670;
  assign n5673 = ~n5669 & n5672;
  assign n5674 = ~n5668 & n5671;
  assign n5675 = ~n5667 & n38419;
  assign n5676 = pi23  & ~n5675;
  assign n5677 = pi23  & ~n5676;
  assign n5678 = pi23  & n5675;
  assign n5679 = ~n5675 & ~n5676;
  assign n5680 = ~pi23  & ~n5675;
  assign n5681 = ~n38420 & ~n38421;
  assign n5682 = n5666 & ~n5681;
  assign n5683 = n4524 & n5576;
  assign n5684 = pi92  & n38406;
  assign n5685 = pi94  & n5591;
  assign n5686 = pi93  & n5593;
  assign n5687 = ~n5685 & ~n5686;
  assign n5688 = ~n5684 & ~n5686;
  assign n5689 = ~n5685 & n5688;
  assign n5690 = ~n5684 & n5687;
  assign n5691 = ~n5683 & n38422;
  assign n5692 = pi23  & ~n5691;
  assign n5693 = pi23  & ~n5692;
  assign n5694 = pi23  & n5691;
  assign n5695 = ~n5691 & ~n5692;
  assign n5696 = ~pi23  & ~n5691;
  assign n5697 = ~n38423 & ~n38424;
  assign n5698 = n5249 & n38348;
  assign n5699 = ~n5249 & n38348;
  assign n5700 = n5249 & ~n38348;
  assign n5701 = ~n5699 & ~n5700;
  assign n5702 = ~n5257 & ~n5698;
  assign n5703 = ~n5697 & ~n38425;
  assign n5704 = n4544 & n5576;
  assign n5705 = pi91  & n38406;
  assign n5706 = pi93  & n5591;
  assign n5707 = pi92  & n5593;
  assign n5708 = ~n5706 & ~n5707;
  assign n5709 = ~n5705 & ~n5707;
  assign n5710 = ~n5706 & n5709;
  assign n5711 = ~n5705 & n5708;
  assign n5712 = ~n5704 & n38426;
  assign n5713 = pi23  & ~n5712;
  assign n5714 = pi23  & ~n5713;
  assign n5715 = pi23  & n5712;
  assign n5716 = ~n5712 & ~n5713;
  assign n5717 = ~pi23  & ~n5712;
  assign n5718 = ~n38427 & ~n38428;
  assign n5719 = n5245 & ~n5247;
  assign n5720 = ~n5248 & ~n5719;
  assign n5721 = ~n5718 & n5720;
  assign n5722 = n4453 & n5576;
  assign n5723 = pi90  & n38406;
  assign n5724 = pi92  & n5591;
  assign n5725 = pi91  & n5593;
  assign n5726 = ~n5724 & ~n5725;
  assign n5727 = ~n5723 & ~n5725;
  assign n5728 = ~n5724 & n5727;
  assign n5729 = ~n5723 & n5726;
  assign n5730 = ~n5722 & n38429;
  assign n5731 = pi23  & ~n5730;
  assign n5732 = pi23  & ~n5731;
  assign n5733 = pi23  & n5730;
  assign n5734 = ~n5730 & ~n5731;
  assign n5735 = ~pi23  & ~n5730;
  assign n5736 = ~n38430 & ~n38431;
  assign n5737 = n5236 & n38345;
  assign n5738 = ~n5244 & ~n5737;
  assign n5739 = ~n5736 & n5738;
  assign n5740 = n5232 & ~n5234;
  assign n5741 = ~n5235 & ~n5740;
  assign n5742 = n594 & n5576;
  assign n5743 = pi89  & n38406;
  assign n5744 = pi91  & n5591;
  assign n5745 = pi90  & n5593;
  assign n5746 = ~n5744 & ~n5745;
  assign n5747 = ~n5743 & ~n5745;
  assign n5748 = ~n5744 & n5747;
  assign n5749 = ~n5743 & n5746;
  assign n5750 = ~n5742 & n38432;
  assign n5751 = pi23  & ~n5750;
  assign n5752 = pi23  & ~n5751;
  assign n5753 = pi23  & n5750;
  assign n5754 = ~n5750 & ~n5751;
  assign n5755 = ~pi23  & ~n5750;
  assign n5756 = ~n38433 & ~n38434;
  assign n5757 = n5741 & ~n5756;
  assign n5758 = n3566 & n5576;
  assign n5759 = pi88  & n38406;
  assign n5760 = pi90  & n5591;
  assign n5761 = pi89  & n5593;
  assign n5762 = ~n5760 & ~n5761;
  assign n5763 = ~n5759 & ~n5761;
  assign n5764 = ~n5760 & n5763;
  assign n5765 = ~n5759 & n5762;
  assign n5766 = ~n5758 & n38435;
  assign n5767 = pi23  & ~n5766;
  assign n5768 = pi23  & ~n5767;
  assign n5769 = pi23  & n5766;
  assign n5770 = ~n5766 & ~n5767;
  assign n5771 = ~pi23  & ~n5766;
  assign n5772 = ~n38436 & ~n38437;
  assign n5773 = n5226 & ~n5228;
  assign n5774 = ~n5226 & ~n38342;
  assign n5775 = ~n5227 & n5232;
  assign n5776 = ~n5774 & ~n5775;
  assign n5777 = ~n38342 & ~n5773;
  assign n5778 = ~n5772 & ~n38438;
  assign n5779 = n5217 & n38341;
  assign n5780 = ~n5225 & ~n5779;
  assign n5781 = n3591 & n5576;
  assign n5782 = pi87  & n38406;
  assign n5783 = pi89  & n5591;
  assign n5784 = pi88  & n5593;
  assign n5785 = ~n5783 & ~n5784;
  assign n5786 = ~n5782 & ~n5784;
  assign n5787 = ~n5783 & n5786;
  assign n5788 = ~n5782 & n5785;
  assign n5789 = ~n5781 & n38439;
  assign n5790 = pi23  & ~n5789;
  assign n5791 = pi23  & ~n5790;
  assign n5792 = pi23  & n5789;
  assign n5793 = ~n5789 & ~n5790;
  assign n5794 = ~pi23  & ~n5789;
  assign n5795 = ~n38440 & ~n38441;
  assign n5796 = n5780 & ~n5795;
  assign n5797 = n5208 & n38338;
  assign n5798 = ~n5216 & ~n5797;
  assign n5799 = n3354 & n5576;
  assign n5800 = pi86  & n38406;
  assign n5801 = pi88  & n5591;
  assign n5802 = pi87  & n5593;
  assign n5803 = ~n5801 & ~n5802;
  assign n5804 = ~n5800 & ~n5802;
  assign n5805 = ~n5801 & n5804;
  assign n5806 = ~n5800 & n5803;
  assign n5807 = ~n5799 & n38442;
  assign n5808 = pi23  & ~n5807;
  assign n5809 = pi23  & ~n5808;
  assign n5810 = pi23  & n5807;
  assign n5811 = ~n5807 & ~n5808;
  assign n5812 = ~pi23  & ~n5807;
  assign n5813 = ~n38443 & ~n38444;
  assign n5814 = n5798 & ~n5813;
  assign n5815 = n5199 & n38335;
  assign n5816 = ~n5207 & ~n5815;
  assign n5817 = n636 & n5576;
  assign n5818 = pi85  & n38406;
  assign n5819 = pi87  & n5591;
  assign n5820 = pi86  & n5593;
  assign n5821 = ~n5819 & ~n5820;
  assign n5822 = ~n5818 & ~n5820;
  assign n5823 = ~n5819 & n5822;
  assign n5824 = ~n5818 & n5821;
  assign n5825 = ~n5817 & n38445;
  assign n5826 = pi23  & ~n5825;
  assign n5827 = pi23  & ~n5826;
  assign n5828 = pi23  & n5825;
  assign n5829 = ~n5825 & ~n5826;
  assign n5830 = ~pi23  & ~n5825;
  assign n5831 = ~n38446 & ~n38447;
  assign n5832 = n5816 & ~n5831;
  assign n5833 = n5190 & n38332;
  assign n5834 = ~n5198 & ~n5833;
  assign n5835 = n2779 & n5576;
  assign n5836 = pi84  & n38406;
  assign n5837 = pi86  & n5591;
  assign n5838 = pi85  & n5593;
  assign n5839 = ~n5837 & ~n5838;
  assign n5840 = ~n5836 & ~n5838;
  assign n5841 = ~n5837 & n5840;
  assign n5842 = ~n5836 & n5839;
  assign n5843 = ~n5835 & n38448;
  assign n5844 = pi23  & ~n5843;
  assign n5845 = pi23  & ~n5844;
  assign n5846 = pi23  & n5843;
  assign n5847 = ~n5843 & ~n5844;
  assign n5848 = ~pi23  & ~n5843;
  assign n5849 = ~n38449 & ~n38450;
  assign n5850 = n5834 & ~n5849;
  assign n5851 = n5186 & ~n5188;
  assign n5852 = ~n5189 & ~n5851;
  assign n5853 = n2804 & n5576;
  assign n5854 = pi83  & n38406;
  assign n5855 = pi85  & n5591;
  assign n5856 = pi84  & n5593;
  assign n5857 = ~n5855 & ~n5856;
  assign n5858 = ~n5854 & ~n5856;
  assign n5859 = ~n5855 & n5858;
  assign n5860 = ~n5854 & n5857;
  assign n5861 = ~n5853 & n38451;
  assign n5862 = pi23  & ~n5861;
  assign n5863 = pi23  & ~n5862;
  assign n5864 = pi23  & n5861;
  assign n5865 = ~n5861 & ~n5862;
  assign n5866 = ~pi23  & ~n5861;
  assign n5867 = ~n38452 & ~n38453;
  assign n5868 = n5852 & ~n5867;
  assign n5869 = n5182 & ~n5184;
  assign n5870 = ~n5185 & ~n5869;
  assign n5871 = n2591 & n5576;
  assign n5872 = pi82  & n38406;
  assign n5873 = pi84  & n5591;
  assign n5874 = pi83  & n5593;
  assign n5875 = ~n5873 & ~n5874;
  assign n5876 = ~n5872 & ~n5874;
  assign n5877 = ~n5873 & n5876;
  assign n5878 = ~n5872 & n5875;
  assign n5879 = ~n5871 & n38454;
  assign n5880 = pi23  & ~n5879;
  assign n5881 = pi23  & ~n5880;
  assign n5882 = pi23  & n5879;
  assign n5883 = ~n5879 & ~n5880;
  assign n5884 = ~pi23  & ~n5879;
  assign n5885 = ~n38455 & ~n38456;
  assign n5886 = n5870 & ~n5885;
  assign n5887 = n5173 & n38329;
  assign n5888 = ~n5181 & ~n5887;
  assign n5889 = n2091 & n5576;
  assign n5890 = pi81  & n38406;
  assign n5891 = pi83  & n5591;
  assign n5892 = pi82  & n5593;
  assign n5893 = ~n5891 & ~n5892;
  assign n5894 = ~n5890 & ~n5892;
  assign n5895 = ~n5891 & n5894;
  assign n5896 = ~n5890 & n5893;
  assign n5897 = ~n5889 & n38457;
  assign n5898 = pi23  & ~n5897;
  assign n5899 = pi23  & ~n5898;
  assign n5900 = pi23  & n5897;
  assign n5901 = ~n5897 & ~n5898;
  assign n5902 = ~pi23  & ~n5897;
  assign n5903 = ~n38458 & ~n38459;
  assign n5904 = n5888 & ~n5903;
  assign n5905 = n2134 & n5576;
  assign n5906 = pi80  & n38406;
  assign n5907 = pi82  & n5591;
  assign n5908 = pi81  & n5593;
  assign n5909 = ~n5907 & ~n5908;
  assign n5910 = ~n5906 & ~n5908;
  assign n5911 = ~n5907 & n5910;
  assign n5912 = ~n5906 & n5909;
  assign n5913 = ~n5905 & n38460;
  assign n5914 = pi23  & ~n5913;
  assign n5915 = pi23  & ~n5914;
  assign n5916 = pi23  & n5913;
  assign n5917 = ~n5913 & ~n5914;
  assign n5918 = ~pi23  & ~n5913;
  assign n5919 = ~n38461 & ~n38462;
  assign n5920 = n5164 & n38326;
  assign n5921 = ~n5164 & n38326;
  assign n5922 = n5164 & ~n38326;
  assign n5923 = ~n5921 & ~n5922;
  assign n5924 = ~n5172 & ~n5920;
  assign n5925 = ~n5919 & ~n38463;
  assign n5926 = n5160 & ~n5162;
  assign n5927 = ~n5163 & ~n5926;
  assign n5928 = n2154 & n5576;
  assign n5929 = pi79  & n38406;
  assign n5930 = pi81  & n5591;
  assign n5931 = pi80  & n5593;
  assign n5932 = ~n5930 & ~n5931;
  assign n5933 = ~n5929 & ~n5931;
  assign n5934 = ~n5930 & n5933;
  assign n5935 = ~n5929 & n5932;
  assign n5936 = ~n5928 & n38464;
  assign n5937 = pi23  & ~n5936;
  assign n5938 = pi23  & ~n5937;
  assign n5939 = pi23  & n5936;
  assign n5940 = ~n5936 & ~n5937;
  assign n5941 = ~pi23  & ~n5936;
  assign n5942 = ~n38465 & ~n38466;
  assign n5943 = n5927 & ~n5942;
  assign n5944 = n5156 & ~n5158;
  assign n5945 = ~n5159 & ~n5944;
  assign n5946 = n2063 & n5576;
  assign n5947 = pi78  & n38406;
  assign n5948 = pi80  & n5591;
  assign n5949 = pi79  & n5593;
  assign n5950 = ~n5948 & ~n5949;
  assign n5951 = ~n5947 & ~n5949;
  assign n5952 = ~n5948 & n5951;
  assign n5953 = ~n5947 & n5950;
  assign n5954 = ~n5946 & n38467;
  assign n5955 = pi23  & ~n5954;
  assign n5956 = pi23  & ~n5955;
  assign n5957 = pi23  & n5954;
  assign n5958 = ~n5954 & ~n5955;
  assign n5959 = ~pi23  & ~n5954;
  assign n5960 = ~n38468 & ~n38469;
  assign n5961 = n5945 & ~n5960;
  assign n5962 = ~n4882 & n5154;
  assign n5963 = ~n5155 & ~n5962;
  assign n5964 = n678 & n5576;
  assign n5965 = pi77  & n38406;
  assign n5966 = pi79  & n5591;
  assign n5967 = pi78  & n5593;
  assign n5968 = ~n5966 & ~n5967;
  assign n5969 = ~n5965 & ~n5967;
  assign n5970 = ~n5966 & n5969;
  assign n5971 = ~n5965 & n5968;
  assign n5972 = ~n5964 & n38470;
  assign n5973 = pi23  & ~n5972;
  assign n5974 = pi23  & ~n5973;
  assign n5975 = pi23  & n5972;
  assign n5976 = ~n5972 & ~n5973;
  assign n5977 = ~pi23  & ~n5972;
  assign n5978 = ~n38471 & ~n38472;
  assign n5979 = n5963 & ~n5978;
  assign n5980 = n1578 & n5576;
  assign n5981 = pi76  & n38406;
  assign n5982 = pi78  & n5591;
  assign n5983 = pi77  & n5593;
  assign n5984 = ~n5982 & ~n5983;
  assign n5985 = ~n5981 & ~n5983;
  assign n5986 = ~n5982 & n5985;
  assign n5987 = ~n5981 & n5984;
  assign n5988 = ~n5980 & n38473;
  assign n5989 = pi23  & ~n5988;
  assign n5990 = pi23  & ~n5989;
  assign n5991 = pi23  & n5988;
  assign n5992 = ~n5988 & ~n5989;
  assign n5993 = ~pi23  & ~n5988;
  assign n5994 = ~n38474 & ~n38475;
  assign n5995 = n5145 & n38323;
  assign n5996 = ~n5145 & ~n5153;
  assign n5997 = ~n5145 & n38323;
  assign n5998 = ~n38323 & ~n5153;
  assign n5999 = n5145 & ~n38323;
  assign n6000 = ~n38476 & ~n38477;
  assign n6001 = ~n5153 & ~n5995;
  assign n6002 = ~n5994 & ~n38478;
  assign n6003 = n5136 & n38320;
  assign n6004 = ~n5144 & ~n6003;
  assign n6005 = n1596 & n5576;
  assign n6006 = pi75  & n38406;
  assign n6007 = pi77  & n5591;
  assign n6008 = pi76  & n5593;
  assign n6009 = ~n6007 & ~n6008;
  assign n6010 = ~n6006 & ~n6008;
  assign n6011 = ~n6007 & n6010;
  assign n6012 = ~n6006 & n6009;
  assign n6013 = ~n6005 & n38479;
  assign n6014 = pi23  & ~n6013;
  assign n6015 = pi23  & ~n6014;
  assign n6016 = pi23  & n6013;
  assign n6017 = ~n6013 & ~n6014;
  assign n6018 = ~pi23  & ~n6013;
  assign n6019 = ~n38480 & ~n38481;
  assign n6020 = n6004 & ~n6019;
  assign n6021 = n5132 & ~n5134;
  assign n6022 = ~n5135 & ~n6021;
  assign n6023 = n1465 & n5576;
  assign n6024 = pi74  & n38406;
  assign n6025 = pi76  & n5591;
  assign n6026 = pi75  & n5593;
  assign n6027 = ~n6025 & ~n6026;
  assign n6028 = ~n6024 & ~n6026;
  assign n6029 = ~n6025 & n6028;
  assign n6030 = ~n6024 & n6027;
  assign n6031 = ~n6023 & n38482;
  assign n6032 = pi23  & ~n6031;
  assign n6033 = pi23  & ~n6032;
  assign n6034 = pi23  & n6031;
  assign n6035 = ~n6031 & ~n6032;
  assign n6036 = ~pi23  & ~n6031;
  assign n6037 = ~n38483 & ~n38484;
  assign n6038 = n6022 & ~n6037;
  assign n6039 = n5123 & n38317;
  assign n6040 = ~n5131 & ~n6039;
  assign n6041 = n720 & n5576;
  assign n6042 = pi73  & n38406;
  assign n6043 = pi75  & n5591;
  assign n6044 = pi74  & n5593;
  assign n6045 = ~n6043 & ~n6044;
  assign n6046 = ~n6042 & ~n6044;
  assign n6047 = ~n6043 & n6046;
  assign n6048 = ~n6042 & n6045;
  assign n6049 = ~n6041 & n38485;
  assign n6050 = pi23  & ~n6049;
  assign n6051 = pi23  & ~n6050;
  assign n6052 = pi23  & n6049;
  assign n6053 = ~n6049 & ~n6050;
  assign n6054 = ~pi23  & ~n6049;
  assign n6055 = ~n38486 & ~n38487;
  assign n6056 = n6040 & ~n6055;
  assign n6057 = n5119 & ~n5121;
  assign n6058 = ~n5122 & ~n6057;
  assign n6059 = n1218 & n5576;
  assign n6060 = pi72  & n38406;
  assign n6061 = pi74  & n5591;
  assign n6062 = pi73  & n5593;
  assign n6063 = ~n6061 & ~n6062;
  assign n6064 = ~n6060 & ~n6062;
  assign n6065 = ~n6061 & n6064;
  assign n6066 = ~n6060 & n6063;
  assign n6067 = ~n6059 & n38488;
  assign n6068 = pi23  & ~n6067;
  assign n6069 = pi23  & ~n6068;
  assign n6070 = pi23  & n6067;
  assign n6071 = ~n6067 & ~n6068;
  assign n6072 = ~pi23  & ~n6067;
  assign n6073 = ~n38489 & ~n38490;
  assign n6074 = n6058 & ~n6073;
  assign n6075 = n1238 & n5576;
  assign n6076 = pi71  & n38406;
  assign n6077 = pi73  & n5591;
  assign n6078 = pi72  & n5593;
  assign n6079 = ~n6077 & ~n6078;
  assign n6080 = ~n6076 & ~n6078;
  assign n6081 = ~n6077 & n6080;
  assign n6082 = ~n6076 & n6079;
  assign n6083 = ~n6075 & n38491;
  assign n6084 = pi23  & ~n6083;
  assign n6085 = pi23  & ~n6084;
  assign n6086 = pi23  & n6083;
  assign n6087 = ~n6083 & ~n6084;
  assign n6088 = ~pi23  & ~n6083;
  assign n6089 = ~n38492 & ~n38493;
  assign n6090 = n5110 & n38314;
  assign n6091 = ~n5110 & n38314;
  assign n6092 = n5110 & ~n38314;
  assign n6093 = ~n6091 & ~n6092;
  assign n6094 = ~n5118 & ~n6090;
  assign n6095 = ~n6089 & ~n38494;
  assign n6096 = n1124 & n5576;
  assign n6097 = pi70  & n38406;
  assign n6098 = pi72  & n5591;
  assign n6099 = pi71  & n5593;
  assign n6100 = ~n6098 & ~n6099;
  assign n6101 = ~n6097 & ~n6099;
  assign n6102 = ~n6098 & n6101;
  assign n6103 = ~n6097 & n6100;
  assign n6104 = ~n6096 & n38495;
  assign n6105 = pi23  & ~n6104;
  assign n6106 = pi23  & ~n6105;
  assign n6107 = pi23  & n6104;
  assign n6108 = ~n6104 & ~n6105;
  assign n6109 = ~pi23  & ~n6104;
  assign n6110 = ~n38496 & ~n38497;
  assign n6111 = n5104 & ~n5106;
  assign n6112 = ~n5104 & ~n38311;
  assign n6113 = ~n5105 & n5110;
  assign n6114 = ~n6112 & ~n6113;
  assign n6115 = ~n38311 & ~n6111;
  assign n6116 = ~n6110 & ~n38498;
  assign n6117 = n927 & n5576;
  assign n6118 = pi69  & n38406;
  assign n6119 = pi71  & n5591;
  assign n6120 = pi70  & n5593;
  assign n6121 = ~n6119 & ~n6120;
  assign n6122 = ~n6118 & ~n6120;
  assign n6123 = ~n6119 & n6122;
  assign n6124 = ~n6118 & n6121;
  assign n6125 = ~n6117 & n38499;
  assign n6126 = pi23  & ~n6125;
  assign n6127 = pi23  & ~n6126;
  assign n6128 = pi23  & n6125;
  assign n6129 = ~n6125 & ~n6126;
  assign n6130 = ~pi23  & ~n6125;
  assign n6131 = ~n38500 & ~n38501;
  assign n6132 = n5097 & n38310;
  assign n6133 = ~n5103 & ~n6132;
  assign n6134 = ~n6131 & n6133;
  assign n6135 = n5090 & n38309;
  assign n6136 = ~n5096 & ~n6135;
  assign n6137 = n972 & n5576;
  assign n6138 = pi68  & n38406;
  assign n6139 = pi70  & n5591;
  assign n6140 = pi69  & n5593;
  assign n6141 = ~n6139 & ~n6140;
  assign n6142 = ~n6138 & ~n6140;
  assign n6143 = ~n6139 & n6142;
  assign n6144 = ~n6138 & n6141;
  assign n6145 = ~n6137 & n38502;
  assign n6146 = pi23  & ~n6145;
  assign n6147 = pi23  & ~n6146;
  assign n6148 = pi23  & n6145;
  assign n6149 = ~n6145 & ~n6146;
  assign n6150 = ~pi23  & ~n6145;
  assign n6151 = ~n38503 & ~n38504;
  assign n6152 = n6136 & ~n6151;
  assign n6153 = n990 & n5576;
  assign n6154 = pi67  & n38406;
  assign n6155 = pi69  & n5591;
  assign n6156 = pi68  & n5593;
  assign n6157 = ~n6155 & ~n6156;
  assign n6158 = ~n6154 & ~n6156;
  assign n6159 = ~n6155 & n6158;
  assign n6160 = ~n6154 & n6157;
  assign n6161 = ~n6153 & n38505;
  assign n6162 = pi23  & ~n6161;
  assign n6163 = pi23  & ~n6162;
  assign n6164 = pi23  & n6161;
  assign n6165 = ~n6161 & ~n6162;
  assign n6166 = ~pi23  & ~n6161;
  assign n6167 = ~n38506 & ~n38507;
  assign n6168 = pi26  & ~n38301;
  assign n6169 = n38304 & ~n6168;
  assign n6170 = ~n38304 & n6168;
  assign n6171 = ~n38301 & n5072;
  assign n6172 = ~n38305 & ~n6171;
  assign n6173 = ~n6169 & ~n6170;
  assign n6174 = ~n6167 & n38508;
  assign n6175 = n871 & n5576;
  assign n6176 = pi66  & n38406;
  assign n6177 = pi68  & n5591;
  assign n6178 = pi67  & n5593;
  assign n6179 = ~n6177 & ~n6178;
  assign n6180 = ~n6176 & ~n6178;
  assign n6181 = ~n6177 & n6180;
  assign n6182 = ~n6176 & n6179;
  assign n6183 = ~n6175 & n38509;
  assign n6184 = pi23  & ~n6183;
  assign n6185 = pi23  & ~n6184;
  assign n6186 = pi23  & n6183;
  assign n6187 = ~n6183 & ~n6184;
  assign n6188 = ~pi23  & ~n6183;
  assign n6189 = ~n38510 & ~n38511;
  assign n6190 = pi26  & n5046;
  assign n6191 = ~n5045 & n6190;
  assign n6192 = n5045 & ~n6190;
  assign n6193 = ~n5047 & n5051;
  assign n6194 = ~n38301 & ~n6193;
  assign n6195 = ~n6191 & ~n6192;
  assign n6196 = ~n6189 & n38512;
  assign n6197 = n37515 & n5576;
  assign n6198 = pi65  & n5591;
  assign n6199 = pi64  & n5593;
  assign n6200 = ~n6198 & ~n6199;
  assign n6201 = ~n6197 & n6200;
  assign n6202 = pi64  & n38403;
  assign n6203 = pi23  & ~n6202;
  assign n6204 = pi23  & ~n6201;
  assign n6205 = pi23  & ~n6204;
  assign n6206 = ~n6201 & ~n6204;
  assign n6207 = ~n6205 & ~n6206;
  assign n6208 = n6203 & ~n6207;
  assign n6209 = n6201 & n6203;
  assign n6210 = pi64  & n38406;
  assign n6211 = pi65  & n5593;
  assign n6212 = ~n37521 & n5576;
  assign n6213 = pi66  & n5591;
  assign n6214 = ~n6212 & ~n6213;
  assign n6215 = ~n6211 & ~n6212;
  assign n6216 = ~n6213 & n6215;
  assign n6217 = ~n6211 & ~n6213;
  assign n6218 = ~n6212 & n6217;
  assign n6219 = ~n6211 & n6214;
  assign n6220 = ~n6210 & ~n6211;
  assign n6221 = ~n6213 & n6220;
  assign n6222 = ~n6210 & n6217;
  assign n6223 = ~n6212 & n38515;
  assign n6224 = ~n6210 & n38514;
  assign n6225 = pi23  & ~n38516;
  assign n6226 = pi23  & ~n6225;
  assign n6227 = ~n38516 & ~n6225;
  assign n6228 = ~n6226 & ~n6227;
  assign n6229 = n38513 & ~n6228;
  assign n6230 = n38513 & n38516;
  assign n6231 = n5046 & n38517;
  assign n6232 = n847 & n5576;
  assign n6233 = pi65  & n38406;
  assign n6234 = pi67  & n5591;
  assign n6235 = pi66  & n5593;
  assign n6236 = ~n6234 & ~n6235;
  assign n6237 = ~n6233 & ~n6235;
  assign n6238 = ~n6234 & n6237;
  assign n6239 = ~n6233 & n6236;
  assign n6240 = ~n6232 & n38518;
  assign n6241 = pi23  & ~n6240;
  assign n6242 = pi23  & ~n6241;
  assign n6243 = pi23  & n6240;
  assign n6244 = ~n6240 & ~n6241;
  assign n6245 = ~pi23  & ~n6240;
  assign n6246 = ~n38519 & ~n38520;
  assign n6247 = ~n5046 & ~n38517;
  assign n6248 = n5046 & ~n38517;
  assign n6249 = ~n5046 & n38517;
  assign n6250 = ~n6248 & ~n6249;
  assign n6251 = ~n6231 & ~n6247;
  assign n6252 = ~n6246 & ~n38521;
  assign n6253 = ~n6231 & ~n6252;
  assign n6254 = n6189 & ~n38512;
  assign n6255 = n6189 & n38512;
  assign n6256 = ~n6189 & ~n38512;
  assign n6257 = ~n6255 & ~n6256;
  assign n6258 = ~n6196 & ~n6254;
  assign n6259 = ~n6253 & ~n38522;
  assign n6260 = ~n6196 & ~n6259;
  assign n6261 = n6167 & ~n38508;
  assign n6262 = ~n6174 & ~n6261;
  assign n6263 = ~n6260 & ~n6261;
  assign n6264 = ~n6174 & n6263;
  assign n6265 = ~n6260 & n6262;
  assign n6266 = ~n6174 & ~n38523;
  assign n6267 = ~n6136 & n6151;
  assign n6268 = n6136 & ~n6152;
  assign n6269 = n6136 & n6151;
  assign n6270 = ~n6151 & ~n6152;
  assign n6271 = ~n6136 & ~n6151;
  assign n6272 = ~n38524 & ~n38525;
  assign n6273 = ~n6152 & ~n6267;
  assign n6274 = ~n6266 & ~n38526;
  assign n6275 = ~n6152 & ~n6274;
  assign n6276 = n6131 & ~n6133;
  assign n6277 = ~n6134 & ~n6276;
  assign n6278 = ~n6275 & n6277;
  assign n6279 = ~n6134 & ~n6278;
  assign n6280 = n6110 & n38498;
  assign n6281 = ~n6116 & ~n6280;
  assign n6282 = ~n6279 & n6281;
  assign n6283 = ~n6116 & ~n6282;
  assign n6284 = n6089 & n38494;
  assign n6285 = ~n6095 & ~n6284;
  assign n6286 = ~n6283 & n6285;
  assign n6287 = ~n6095 & ~n6286;
  assign n6288 = ~n6058 & n6073;
  assign n6289 = n6058 & ~n6074;
  assign n6290 = n6058 & n6073;
  assign n6291 = ~n6073 & ~n6074;
  assign n6292 = ~n6058 & ~n6073;
  assign n6293 = ~n38527 & ~n38528;
  assign n6294 = ~n6074 & ~n6288;
  assign n6295 = ~n6287 & ~n38529;
  assign n6296 = ~n6074 & ~n6295;
  assign n6297 = ~n6040 & n6055;
  assign n6298 = ~n6056 & ~n6297;
  assign n6299 = ~n6296 & ~n6297;
  assign n6300 = ~n6056 & n6299;
  assign n6301 = ~n6296 & n6298;
  assign n6302 = ~n6056 & ~n38530;
  assign n6303 = ~n6022 & n6037;
  assign n6304 = ~n6038 & ~n6303;
  assign n6305 = ~n6302 & n6304;
  assign n6306 = ~n6038 & ~n6305;
  assign n6307 = ~n6004 & n6019;
  assign n6308 = ~n6020 & ~n6307;
  assign n6309 = ~n6306 & ~n6307;
  assign n6310 = ~n6020 & n6309;
  assign n6311 = ~n6306 & n6308;
  assign n6312 = ~n6020 & ~n38531;
  assign n6313 = n5994 & n38478;
  assign n6314 = ~n6002 & ~n6313;
  assign n6315 = ~n6312 & n6314;
  assign n6316 = ~n6002 & ~n6315;
  assign n6317 = ~n5963 & n5978;
  assign n6318 = n5963 & ~n5979;
  assign n6319 = n5963 & n5978;
  assign n6320 = ~n5978 & ~n5979;
  assign n6321 = ~n5963 & ~n5978;
  assign n6322 = ~n38532 & ~n38533;
  assign n6323 = ~n5979 & ~n6317;
  assign n6324 = ~n6316 & ~n38534;
  assign n6325 = ~n5979 & ~n6324;
  assign n6326 = ~n5945 & n5960;
  assign n6327 = n5945 & ~n5961;
  assign n6328 = n5945 & n5960;
  assign n6329 = ~n5960 & ~n5961;
  assign n6330 = ~n5945 & ~n5960;
  assign n6331 = ~n38535 & ~n38536;
  assign n6332 = ~n5961 & ~n6326;
  assign n6333 = ~n6325 & ~n38537;
  assign n6334 = ~n5961 & ~n6333;
  assign n6335 = ~n5927 & n5942;
  assign n6336 = n5927 & ~n5943;
  assign n6337 = n5927 & n5942;
  assign n6338 = ~n5942 & ~n5943;
  assign n6339 = ~n5927 & ~n5942;
  assign n6340 = ~n38538 & ~n38539;
  assign n6341 = ~n5943 & ~n6335;
  assign n6342 = ~n6334 & ~n38540;
  assign n6343 = ~n5943 & ~n6342;
  assign n6344 = n5919 & n38463;
  assign n6345 = ~n5925 & ~n6344;
  assign n6346 = ~n6343 & n6345;
  assign n6347 = ~n5925 & ~n6346;
  assign n6348 = ~n5888 & n5903;
  assign n6349 = n5888 & ~n5904;
  assign n6350 = n5888 & n5903;
  assign n6351 = ~n5903 & ~n5904;
  assign n6352 = ~n5888 & ~n5903;
  assign n6353 = ~n38541 & ~n38542;
  assign n6354 = ~n5904 & ~n6348;
  assign n6355 = ~n6347 & ~n38543;
  assign n6356 = ~n5904 & ~n6355;
  assign n6357 = ~n5870 & n5885;
  assign n6358 = n5870 & ~n5886;
  assign n6359 = n5870 & n5885;
  assign n6360 = ~n5885 & ~n5886;
  assign n6361 = ~n5870 & ~n5885;
  assign n6362 = ~n38544 & ~n38545;
  assign n6363 = ~n5886 & ~n6357;
  assign n6364 = ~n6356 & ~n38546;
  assign n6365 = ~n5886 & ~n6364;
  assign n6366 = ~n5852 & n5867;
  assign n6367 = n5852 & ~n5868;
  assign n6368 = n5852 & n5867;
  assign n6369 = ~n5867 & ~n5868;
  assign n6370 = ~n5852 & ~n5867;
  assign n6371 = ~n38547 & ~n38548;
  assign n6372 = ~n5868 & ~n6366;
  assign n6373 = ~n6365 & ~n38549;
  assign n6374 = ~n5868 & ~n6373;
  assign n6375 = ~n5834 & n5849;
  assign n6376 = n5834 & ~n5850;
  assign n6377 = n5834 & n5849;
  assign n6378 = ~n5849 & ~n5850;
  assign n6379 = ~n5834 & ~n5849;
  assign n6380 = ~n38550 & ~n38551;
  assign n6381 = ~n5850 & ~n6375;
  assign n6382 = ~n6374 & ~n38552;
  assign n6383 = ~n5850 & ~n6382;
  assign n6384 = ~n5816 & n5831;
  assign n6385 = ~n5832 & ~n6384;
  assign n6386 = ~n6383 & ~n6384;
  assign n6387 = ~n5832 & n6386;
  assign n6388 = ~n6383 & n6385;
  assign n6389 = ~n5832 & ~n38553;
  assign n6390 = ~n5798 & n5813;
  assign n6391 = ~n5814 & ~n6390;
  assign n6392 = ~n6389 & n6391;
  assign n6393 = ~n5814 & ~n6392;
  assign n6394 = ~n5780 & n5795;
  assign n6395 = n5780 & ~n5796;
  assign n6396 = n5780 & n5795;
  assign n6397 = ~n5795 & ~n5796;
  assign n6398 = ~n5780 & ~n5795;
  assign n6399 = ~n38554 & ~n38555;
  assign n6400 = ~n5796 & ~n6394;
  assign n6401 = ~n6393 & ~n38556;
  assign n6402 = ~n5796 & ~n6401;
  assign n6403 = n5772 & n38438;
  assign n6404 = ~n5778 & ~n6403;
  assign n6405 = ~n6402 & n6404;
  assign n6406 = ~n5778 & ~n6405;
  assign n6407 = ~n5741 & n5756;
  assign n6408 = n5741 & ~n5757;
  assign n6409 = n5741 & n5756;
  assign n6410 = ~n5756 & ~n5757;
  assign n6411 = ~n5741 & ~n5756;
  assign n6412 = ~n38557 & ~n38558;
  assign n6413 = ~n5757 & ~n6407;
  assign n6414 = ~n6406 & ~n38559;
  assign n6415 = ~n5757 & ~n6414;
  assign n6416 = n5736 & ~n5738;
  assign n6417 = ~n5736 & ~n5739;
  assign n6418 = ~n5736 & ~n5738;
  assign n6419 = n5738 & ~n5739;
  assign n6420 = n5736 & n5738;
  assign n6421 = ~n38560 & ~n38561;
  assign n6422 = ~n5739 & ~n6416;
  assign n6423 = ~n6415 & ~n38562;
  assign n6424 = ~n5739 & ~n6423;
  assign n6425 = n5718 & ~n5720;
  assign n6426 = ~n5721 & ~n6425;
  assign n6427 = ~n6424 & n6426;
  assign n6428 = ~n5721 & ~n6427;
  assign n6429 = n5697 & n38425;
  assign n6430 = ~n5703 & ~n6429;
  assign n6431 = ~n6428 & n6430;
  assign n6432 = ~n5703 & ~n6431;
  assign n6433 = ~n5666 & n5681;
  assign n6434 = n5666 & ~n5682;
  assign n6435 = n5666 & n5681;
  assign n6436 = ~n5681 & ~n5682;
  assign n6437 = ~n5666 & ~n5681;
  assign n6438 = ~n38563 & ~n38564;
  assign n6439 = ~n5682 & ~n6433;
  assign n6440 = ~n6432 & ~n38565;
  assign n6441 = ~n5682 & ~n6440;
  assign n6442 = n5661 & ~n5663;
  assign n6443 = ~n5664 & ~n6442;
  assign n6444 = ~n6441 & n6443;
  assign n6445 = ~n5664 & ~n6444;
  assign n6446 = ~n5628 & n5645;
  assign n6447 = n5628 & ~n5646;
  assign n6448 = n5628 & n5645;
  assign n6449 = ~n5645 & ~n5646;
  assign n6450 = ~n5628 & ~n5645;
  assign n6451 = ~n38566 & ~n38567;
  assign n6452 = ~n5646 & ~n6446;
  assign n6453 = ~n6445 & ~n38568;
  assign n6454 = ~n5646 & ~n6453;
  assign n6455 = ~n5608 & n5625;
  assign n6456 = n5608 & ~n5626;
  assign n6457 = n5608 & n5625;
  assign n6458 = ~n5625 & ~n5626;
  assign n6459 = ~n5608 & ~n5625;
  assign n6460 = ~n38569 & ~n38570;
  assign n6461 = ~n5626 & ~n6455;
  assign n6462 = ~n6454 & ~n38571;
  assign n6463 = ~n5626 & ~n6462;
  assign n6464 = ~n5563 & n5605;
  assign n6465 = n5563 & ~n5606;
  assign n6466 = n5563 & n5605;
  assign n6467 = ~n5605 & ~n5606;
  assign n6468 = ~n5563 & ~n5605;
  assign n6469 = ~n38572 & ~n38573;
  assign n6470 = ~n5606 & ~n6464;
  assign n6471 = ~n6463 & ~n38574;
  assign n6472 = ~n5606 & ~n6471;
  assign n6473 = n457 & ~n459;
  assign n6474 = ~n460 & ~n6473;
  assign n6475 = n5576 & n6474;
  assign n6476 = pi98  & n38406;
  assign n6477 = pi100  & n5591;
  assign n6478 = pi99  & n5593;
  assign n6479 = ~n6477 & ~n6478;
  assign n6480 = ~n6476 & ~n6478;
  assign n6481 = ~n6477 & n6480;
  assign n6482 = ~n6476 & n6479;
  assign n6483 = ~n6475 & n38575;
  assign n6484 = pi23  & ~n6483;
  assign n6485 = pi23  & ~n6484;
  assign n6486 = pi23  & n6483;
  assign n6487 = ~n6483 & ~n6484;
  assign n6488 = ~pi23  & ~n6483;
  assign n6489 = ~n38576 & ~n38577;
  assign n6490 = ~n5559 & ~n5561;
  assign n6491 = ~n5553 & ~n5555;
  assign n6492 = n607 & n4524;
  assign n6493 = pi92  & n37489;
  assign n6494 = pi94  & n620;
  assign n6495 = pi93  & n622;
  assign n6496 = ~n6494 & ~n6495;
  assign n6497 = ~n6493 & ~n6495;
  assign n6498 = ~n6494 & n6497;
  assign n6499 = ~n6493 & n6496;
  assign n6500 = ~n6492 & n38578;
  assign n6501 = pi29  & ~n6500;
  assign n6502 = pi29  & ~n6501;
  assign n6503 = pi29  & n6500;
  assign n6504 = ~n6500 & ~n6501;
  assign n6505 = ~pi29  & ~n6500;
  assign n6506 = ~n38579 & ~n38580;
  assign n6507 = ~n5519 & ~n5523;
  assign n6508 = ~n5507 & ~n5513;
  assign n6509 = n691 & n2804;
  assign n6510 = pi83  & n37503;
  assign n6511 = pi85  & n704;
  assign n6512 = pi84  & n706;
  assign n6513 = ~n6511 & ~n6512;
  assign n6514 = ~n6510 & ~n6512;
  assign n6515 = ~n6511 & n6514;
  assign n6516 = ~n6510 & n6513;
  assign n6517 = ~n6509 & n38581;
  assign n6518 = pi38  & ~n6517;
  assign n6519 = pi38  & ~n6518;
  assign n6520 = pi38  & n6517;
  assign n6521 = ~n6517 & ~n6518;
  assign n6522 = ~pi38  & ~n6517;
  assign n6523 = ~n38582 & ~n38583;
  assign n6524 = ~n5491 & ~n5499;
  assign n6525 = n733 & n2134;
  assign n6526 = pi80  & n37510;
  assign n6527 = pi82  & n746;
  assign n6528 = pi81  & n748;
  assign n6529 = ~n6527 & ~n6528;
  assign n6530 = ~n6526 & ~n6528;
  assign n6531 = ~n6527 & n6530;
  assign n6532 = ~n6526 & n6529;
  assign n6533 = ~n6525 & n38584;
  assign n6534 = pi41  & ~n6533;
  assign n6535 = pi41  & ~n6534;
  assign n6536 = pi41  & n6533;
  assign n6537 = ~n6533 & ~n6534;
  assign n6538 = ~pi41  & ~n6533;
  assign n6539 = ~n38585 & ~n38586;
  assign n6540 = ~n5480 & ~n5488;
  assign n6541 = n678 & n940;
  assign n6542 = pi77  & n37541;
  assign n6543 = pi79  & n953;
  assign n6544 = pi78  & n955;
  assign n6545 = ~n6543 & ~n6544;
  assign n6546 = ~n6542 & ~n6544;
  assign n6547 = ~n6543 & n6546;
  assign n6548 = ~n6542 & n6545;
  assign n6549 = ~n6541 & n38587;
  assign n6550 = pi44  & ~n6549;
  assign n6551 = pi44  & ~n6550;
  assign n6552 = pi44  & n6549;
  assign n6553 = ~n6549 & ~n6550;
  assign n6554 = ~pi44  & ~n6549;
  assign n6555 = ~n38588 & ~n38589;
  assign n6556 = ~n5460 & ~n5462;
  assign n6557 = n785 & n1465;
  assign n6558 = pi74  & n37520;
  assign n6559 = pi76  & n787;
  assign n6560 = pi75  & n795;
  assign n6561 = ~n6559 & ~n6560;
  assign n6562 = ~n6558 & ~n6560;
  assign n6563 = ~n6559 & n6562;
  assign n6564 = ~n6558 & n6561;
  assign n6565 = ~n6557 & n38590;
  assign n6566 = pi47  & ~n6565;
  assign n6567 = pi47  & ~n6566;
  assign n6568 = pi47  & n6565;
  assign n6569 = ~n6565 & ~n6566;
  assign n6570 = ~pi47  & ~n6565;
  assign n6571 = ~n38591 & ~n38592;
  assign n6572 = ~n5454 & ~n5456;
  assign n6573 = n894 & n1238;
  assign n6574 = pi71  & n37580;
  assign n6575 = pi73  & n896;
  assign n6576 = pi72  & n904;
  assign n6577 = ~n6575 & ~n6576;
  assign n6578 = ~n6574 & ~n6576;
  assign n6579 = ~n6575 & n6578;
  assign n6580 = ~n6574 & n6577;
  assign n6581 = ~n6573 & n38593;
  assign n6582 = pi50  & ~n6581;
  assign n6583 = pi50  & ~n6582;
  assign n6584 = pi50  & n6581;
  assign n6585 = ~n6581 & ~n6582;
  assign n6586 = ~pi50  & ~n6581;
  assign n6587 = ~n38594 & ~n38595;
  assign n6588 = n847 & n4312;
  assign n6589 = pi65  & n38376;
  assign n6590 = pi67  & n4314;
  assign n6591 = pi66  & n4322;
  assign n6592 = ~n6590 & ~n6591;
  assign n6593 = ~n6589 & ~n6591;
  assign n6594 = ~n6590 & n6593;
  assign n6595 = ~n6589 & n6592;
  assign n6596 = ~n6588 & n38596;
  assign n6597 = pi56  & ~n6596;
  assign n6598 = pi56  & ~n6597;
  assign n6599 = pi56  & n6596;
  assign n6600 = ~n6596 & ~n6597;
  assign n6601 = ~pi56  & ~n6596;
  assign n6602 = ~n38597 & ~n38598;
  assign n6603 = pi56  & ~pi57 ;
  assign n6604 = ~pi56  & pi57 ;
  assign n6605 = ~pi56  & ~pi57 ;
  assign n6606 = pi56  & pi57 ;
  assign n6607 = ~n6605 & ~n6606;
  assign n6608 = ~n6603 & ~n6604;
  assign n6609 = pi64  & n38599;
  assign n6610 = n38380 & n6609;
  assign n6611 = ~n38380 & ~n6609;
  assign n6612 = ~n38380 & n6609;
  assign n6613 = n38380 & ~n6609;
  assign n6614 = ~n6612 & ~n6613;
  assign n6615 = ~n6610 & ~n6611;
  assign n6616 = ~n6602 & ~n38600;
  assign n6617 = n6602 & n38600;
  assign n6618 = ~n6616 & ~n6617;
  assign n6619 = n972 & n1971;
  assign n6620 = pi68  & n37864;
  assign n6621 = pi70  & n1973;
  assign n6622 = pi69  & n1981;
  assign n6623 = ~n6621 & ~n6622;
  assign n6624 = ~n6620 & ~n6622;
  assign n6625 = ~n6621 & n6624;
  assign n6626 = ~n6620 & n6623;
  assign n6627 = ~n6619 & n38601;
  assign n6628 = pi53  & ~n6627;
  assign n6629 = pi53  & ~n6628;
  assign n6630 = pi53  & n6627;
  assign n6631 = ~n6627 & ~n6628;
  assign n6632 = ~pi53  & ~n6627;
  assign n6633 = ~n38602 & ~n38603;
  assign n6634 = n6618 & ~n6633;
  assign n6635 = ~n6618 & n6633;
  assign n6636 = n6618 & ~n6634;
  assign n6637 = n6618 & n6633;
  assign n6638 = ~n6633 & ~n6634;
  assign n6639 = ~n6618 & ~n6633;
  assign n6640 = ~n38604 & ~n38605;
  assign n6641 = ~n6634 & ~n6635;
  assign n6642 = ~n5449 & ~n38606;
  assign n6643 = n5449 & n38606;
  assign n6644 = ~n5449 & n38606;
  assign n6645 = n5449 & ~n38606;
  assign n6646 = ~n6644 & ~n6645;
  assign n6647 = ~n6642 & ~n6643;
  assign n6648 = ~n6587 & ~n38607;
  assign n6649 = n6587 & n38607;
  assign n6650 = ~n6648 & ~n6649;
  assign n6651 = ~n6572 & n6650;
  assign n6652 = n6572 & ~n6650;
  assign n6653 = ~n6651 & ~n6652;
  assign n6654 = n6571 & ~n6653;
  assign n6655 = ~n6571 & n6653;
  assign n6656 = ~n6654 & ~n6655;
  assign n6657 = ~n6556 & n6656;
  assign n6658 = n6556 & ~n6656;
  assign n6659 = ~n6657 & ~n6658;
  assign n6660 = ~n6555 & n6659;
  assign n6661 = n6555 & ~n6659;
  assign n6662 = ~n6660 & ~n6661;
  assign n6663 = ~n6540 & n6662;
  assign n6664 = n6540 & ~n6662;
  assign n6665 = ~n6663 & ~n6664;
  assign n6666 = ~n6539 & n6665;
  assign n6667 = n6539 & ~n6665;
  assign n6668 = ~n6539 & ~n6666;
  assign n6669 = ~n6539 & ~n6665;
  assign n6670 = n6665 & ~n6666;
  assign n6671 = n6539 & n6665;
  assign n6672 = ~n38608 & ~n38609;
  assign n6673 = ~n6666 & ~n6667;
  assign n6674 = ~n6524 & ~n38610;
  assign n6675 = n6524 & ~n38609;
  assign n6676 = ~n38608 & n6675;
  assign n6677 = n6524 & n38610;
  assign n6678 = ~n6674 & ~n38611;
  assign n6679 = ~n6523 & n6678;
  assign n6680 = n6523 & ~n6678;
  assign n6681 = ~n6679 & ~n6680;
  assign n6682 = ~n6508 & n6681;
  assign n6683 = n6508 & ~n6681;
  assign n6684 = ~n6682 & ~n6683;
  assign n6685 = n2104 & n3354;
  assign n6686 = pi86  & n37758;
  assign n6687 = pi88  & n2117;
  assign n6688 = pi87  & n2119;
  assign n6689 = ~n6687 & ~n6688;
  assign n6690 = ~n6686 & ~n6688;
  assign n6691 = ~n6687 & n6690;
  assign n6692 = ~n6686 & n6689;
  assign n6693 = ~n6685 & n38612;
  assign n6694 = pi35  & ~n6693;
  assign n6695 = pi35  & ~n6694;
  assign n6696 = pi35  & n6693;
  assign n6697 = ~n6693 & ~n6694;
  assign n6698 = ~pi35  & ~n6693;
  assign n6699 = ~n38613 & ~n38614;
  assign n6700 = n6684 & ~n6699;
  assign n6701 = ~n6684 & n6699;
  assign n6702 = n6684 & ~n6700;
  assign n6703 = n6684 & n6699;
  assign n6704 = ~n6699 & ~n6700;
  assign n6705 = ~n6684 & ~n6699;
  assign n6706 = ~n38615 & ~n38616;
  assign n6707 = ~n6700 & ~n6701;
  assign n6708 = n6507 & n38617;
  assign n6709 = ~n6507 & ~n38617;
  assign n6710 = ~n6708 & ~n6709;
  assign n6711 = n594 & n649;
  assign n6712 = pi89  & n37496;
  assign n6713 = pi91  & n662;
  assign n6714 = pi90  & n664;
  assign n6715 = ~n6713 & ~n6714;
  assign n6716 = ~n6712 & ~n6714;
  assign n6717 = ~n6713 & n6716;
  assign n6718 = ~n6712 & n6715;
  assign n6719 = ~n6711 & n38618;
  assign n6720 = pi32  & ~n6719;
  assign n6721 = pi32  & ~n6720;
  assign n6722 = pi32  & n6719;
  assign n6723 = ~n6719 & ~n6720;
  assign n6724 = ~pi32  & ~n6719;
  assign n6725 = ~n38619 & ~n38620;
  assign n6726 = ~n6710 & n6725;
  assign n6727 = n6710 & ~n6725;
  assign n6728 = ~n6726 & ~n6727;
  assign n6729 = ~n5548 & n6728;
  assign n6730 = n5548 & ~n6728;
  assign n6731 = ~n6729 & ~n6730;
  assign n6732 = ~n6506 & n6731;
  assign n6733 = n6506 & ~n6731;
  assign n6734 = ~n6732 & ~n6733;
  assign n6735 = ~n6491 & n6734;
  assign n6736 = n6491 & ~n6734;
  assign n6737 = ~n6735 & ~n6736;
  assign n6738 = n4492 & n5630;
  assign n6739 = pi95  & n38208;
  assign n6740 = pi97  & n4507;
  assign n6741 = pi96  & n4509;
  assign n6742 = ~n6740 & ~n6741;
  assign n6743 = ~n6739 & ~n6741;
  assign n6744 = ~n6740 & n6743;
  assign n6745 = ~n6739 & n6742;
  assign n6746 = ~n6738 & n38621;
  assign n6747 = pi26  & ~n6746;
  assign n6748 = pi26  & ~n6747;
  assign n6749 = pi26  & n6746;
  assign n6750 = ~n6746 & ~n6747;
  assign n6751 = ~pi26  & ~n6746;
  assign n6752 = ~n38622 & ~n38623;
  assign n6753 = n6737 & ~n6752;
  assign n6754 = ~n6737 & n6752;
  assign n6755 = n6737 & ~n6753;
  assign n6756 = n6737 & n6752;
  assign n6757 = ~n6752 & ~n6753;
  assign n6758 = ~n6737 & ~n6752;
  assign n6759 = ~n38624 & ~n38625;
  assign n6760 = ~n6753 & ~n6754;
  assign n6761 = ~n6490 & ~n38626;
  assign n6762 = n6490 & n38626;
  assign n6763 = ~n6490 & n38626;
  assign n6764 = n6490 & ~n38626;
  assign n6765 = ~n6763 & ~n6764;
  assign n6766 = ~n6761 & ~n6762;
  assign n6767 = ~n6489 & ~n38627;
  assign n6768 = n6489 & n38627;
  assign n6769 = ~n6767 & ~n6768;
  assign n6770 = n6472 & ~n6769;
  assign n6771 = ~n6472 & n6769;
  assign n6772 = ~n6770 & ~n6771;
  assign n6773 = pi17  & ~pi18 ;
  assign n6774 = ~pi17  & pi18 ;
  assign n6775 = ~pi17  & ~pi18 ;
  assign n6776 = pi17  & pi18 ;
  assign n6777 = ~n6775 & ~n6776;
  assign n6778 = ~n6773 & ~n6774;
  assign n6779 = pi19  & ~pi20 ;
  assign n6780 = ~pi19  & pi20 ;
  assign n6781 = ~pi19  & ~pi20 ;
  assign n6782 = pi19  & pi20 ;
  assign n6783 = ~n6781 & ~n6782;
  assign n6784 = ~n6779 & ~n6780;
  assign n6785 = n38628 & n38629;
  assign n6786 = n469 & ~n471;
  assign n6787 = ~n472 & ~n6786;
  assign n6788 = n6785 & n6787;
  assign n6789 = pi18  & ~pi19 ;
  assign n6790 = ~pi18  & pi19 ;
  assign n6791 = ~pi18  & ~pi19 ;
  assign n6792 = pi18  & pi19 ;
  assign n6793 = ~n6791 & ~n6792;
  assign n6794 = ~n6789 & ~n6790;
  assign n6795 = ~n38628 & n38629;
  assign n6796 = ~n38628 & ~n38630;
  assign n6797 = n38629 & n6796;
  assign n6798 = ~n38630 & n6795;
  assign n6799 = pi101  & n38631;
  assign n6800 = n38628 & ~n38629;
  assign n6801 = pi103  & n6800;
  assign n6802 = ~n38628 & n38630;
  assign n6803 = pi102  & n6802;
  assign n6804 = ~n6801 & ~n6803;
  assign n6805 = ~n6799 & ~n6803;
  assign n6806 = ~n6801 & n6805;
  assign n6807 = ~n6799 & n6804;
  assign n6808 = ~n6788 & n38632;
  assign n6809 = pi20  & ~n6808;
  assign n6810 = pi20  & ~n6809;
  assign n6811 = pi20  & n6808;
  assign n6812 = ~n6808 & ~n6809;
  assign n6813 = ~pi20  & ~n6808;
  assign n6814 = ~n38633 & ~n38634;
  assign n6815 = n6772 & ~n6814;
  assign n6816 = n6463 & n38574;
  assign n6817 = ~n6471 & ~n6816;
  assign n6818 = n465 & ~n467;
  assign n6819 = ~n468 & ~n6818;
  assign n6820 = n6785 & n6819;
  assign n6821 = pi100  & n38631;
  assign n6822 = pi102  & n6800;
  assign n6823 = pi101  & n6802;
  assign n6824 = ~n6822 & ~n6823;
  assign n6825 = ~n6821 & ~n6823;
  assign n6826 = ~n6822 & n6825;
  assign n6827 = ~n6821 & n6824;
  assign n6828 = ~n6820 & n38635;
  assign n6829 = pi20  & ~n6828;
  assign n6830 = pi20  & ~n6829;
  assign n6831 = pi20  & n6828;
  assign n6832 = ~n6828 & ~n6829;
  assign n6833 = ~pi20  & ~n6828;
  assign n6834 = ~n38636 & ~n38637;
  assign n6835 = n6817 & ~n6834;
  assign n6836 = n6454 & n38571;
  assign n6837 = ~n6462 & ~n6836;
  assign n6838 = n461 & ~n463;
  assign n6839 = ~n464 & ~n6838;
  assign n6840 = n6785 & n6839;
  assign n6841 = pi99  & n38631;
  assign n6842 = pi101  & n6800;
  assign n6843 = pi100  & n6802;
  assign n6844 = ~n6842 & ~n6843;
  assign n6845 = ~n6841 & ~n6843;
  assign n6846 = ~n6842 & n6845;
  assign n6847 = ~n6841 & n6844;
  assign n6848 = ~n6840 & n38638;
  assign n6849 = pi20  & ~n6848;
  assign n6850 = pi20  & ~n6849;
  assign n6851 = pi20  & n6848;
  assign n6852 = ~n6848 & ~n6849;
  assign n6853 = ~pi20  & ~n6848;
  assign n6854 = ~n38639 & ~n38640;
  assign n6855 = n6837 & ~n6854;
  assign n6856 = n6474 & n6785;
  assign n6857 = pi98  & n38631;
  assign n6858 = pi100  & n6800;
  assign n6859 = pi99  & n6802;
  assign n6860 = ~n6858 & ~n6859;
  assign n6861 = ~n6857 & ~n6859;
  assign n6862 = ~n6858 & n6861;
  assign n6863 = ~n6857 & n6860;
  assign n6864 = ~n6856 & n38641;
  assign n6865 = pi20  & ~n6864;
  assign n6866 = pi20  & ~n6865;
  assign n6867 = pi20  & n6864;
  assign n6868 = ~n6864 & ~n6865;
  assign n6869 = ~pi20  & ~n6864;
  assign n6870 = ~n38642 & ~n38643;
  assign n6871 = n6445 & n38568;
  assign n6872 = ~n6445 & n38568;
  assign n6873 = n6445 & ~n38568;
  assign n6874 = ~n6872 & ~n6873;
  assign n6875 = ~n6453 & ~n6871;
  assign n6876 = ~n6870 & ~n38644;
  assign n6877 = n6441 & ~n6443;
  assign n6878 = ~n6444 & ~n6877;
  assign n6879 = n5578 & n6785;
  assign n6880 = pi97  & n38631;
  assign n6881 = pi99  & n6800;
  assign n6882 = pi98  & n6802;
  assign n6883 = ~n6881 & ~n6882;
  assign n6884 = ~n6880 & ~n6882;
  assign n6885 = ~n6881 & n6884;
  assign n6886 = ~n6880 & n6883;
  assign n6887 = ~n6879 & n38645;
  assign n6888 = pi20  & ~n6887;
  assign n6889 = pi20  & ~n6888;
  assign n6890 = pi20  & n6887;
  assign n6891 = ~n6887 & ~n6888;
  assign n6892 = ~pi20  & ~n6887;
  assign n6893 = ~n38646 & ~n38647;
  assign n6894 = n6878 & ~n6893;
  assign n6895 = n6432 & n38565;
  assign n6896 = ~n6440 & ~n6895;
  assign n6897 = n5610 & n6785;
  assign n6898 = pi96  & n38631;
  assign n6899 = pi98  & n6800;
  assign n6900 = pi97  & n6802;
  assign n6901 = ~n6899 & ~n6900;
  assign n6902 = ~n6898 & ~n6900;
  assign n6903 = ~n6899 & n6902;
  assign n6904 = ~n6898 & n6901;
  assign n6905 = ~n6897 & n38648;
  assign n6906 = pi20  & ~n6905;
  assign n6907 = pi20  & ~n6906;
  assign n6908 = pi20  & n6905;
  assign n6909 = ~n6905 & ~n6906;
  assign n6910 = ~pi20  & ~n6905;
  assign n6911 = ~n38649 & ~n38650;
  assign n6912 = n6896 & ~n6911;
  assign n6913 = n6428 & ~n6430;
  assign n6914 = ~n6431 & ~n6913;
  assign n6915 = n5630 & n6785;
  assign n6916 = pi95  & n38631;
  assign n6917 = pi97  & n6800;
  assign n6918 = pi96  & n6802;
  assign n6919 = ~n6917 & ~n6918;
  assign n6920 = ~n6916 & ~n6918;
  assign n6921 = ~n6917 & n6920;
  assign n6922 = ~n6916 & n6919;
  assign n6923 = ~n6915 & n38651;
  assign n6924 = pi20  & ~n6923;
  assign n6925 = pi20  & ~n6924;
  assign n6926 = pi20  & n6923;
  assign n6927 = ~n6923 & ~n6924;
  assign n6928 = ~pi20  & ~n6923;
  assign n6929 = ~n38652 & ~n38653;
  assign n6930 = n6914 & ~n6929;
  assign n6931 = n5281 & n6785;
  assign n6932 = pi94  & n38631;
  assign n6933 = pi96  & n6800;
  assign n6934 = pi95  & n6802;
  assign n6935 = ~n6933 & ~n6934;
  assign n6936 = ~n6932 & ~n6934;
  assign n6937 = ~n6933 & n6936;
  assign n6938 = ~n6932 & n6935;
  assign n6939 = ~n6931 & n38654;
  assign n6940 = pi20  & ~n6939;
  assign n6941 = pi20  & ~n6940;
  assign n6942 = pi20  & n6939;
  assign n6943 = ~n6939 & ~n6940;
  assign n6944 = ~pi20  & ~n6939;
  assign n6945 = ~n38655 & ~n38656;
  assign n6946 = n6424 & ~n6426;
  assign n6947 = ~n6427 & ~n6946;
  assign n6948 = ~n6945 & n6947;
  assign n6949 = n4494 & n6785;
  assign n6950 = pi93  & n38631;
  assign n6951 = pi95  & n6800;
  assign n6952 = pi94  & n6802;
  assign n6953 = ~n6951 & ~n6952;
  assign n6954 = ~n6950 & ~n6952;
  assign n6955 = ~n6951 & n6954;
  assign n6956 = ~n6950 & n6953;
  assign n6957 = ~n6949 & n38657;
  assign n6958 = pi20  & ~n6957;
  assign n6959 = pi20  & ~n6958;
  assign n6960 = pi20  & n6957;
  assign n6961 = ~n6957 & ~n6958;
  assign n6962 = ~pi20  & ~n6957;
  assign n6963 = ~n38658 & ~n38659;
  assign n6964 = n6415 & n38562;
  assign n6965 = ~n6415 & ~n6423;
  assign n6966 = ~n6415 & n38562;
  assign n6967 = ~n38562 & ~n6423;
  assign n6968 = n6415 & ~n38562;
  assign n6969 = ~n38660 & ~n38661;
  assign n6970 = ~n6423 & ~n6964;
  assign n6971 = ~n6963 & ~n38662;
  assign n6972 = n4524 & n6785;
  assign n6973 = pi92  & n38631;
  assign n6974 = pi94  & n6800;
  assign n6975 = pi93  & n6802;
  assign n6976 = ~n6974 & ~n6975;
  assign n6977 = ~n6973 & ~n6975;
  assign n6978 = ~n6974 & n6977;
  assign n6979 = ~n6973 & n6976;
  assign n6980 = ~n6972 & n38663;
  assign n6981 = pi20  & ~n6980;
  assign n6982 = pi20  & ~n6981;
  assign n6983 = pi20  & n6980;
  assign n6984 = ~n6980 & ~n6981;
  assign n6985 = ~pi20  & ~n6980;
  assign n6986 = ~n38664 & ~n38665;
  assign n6987 = n6406 & n38559;
  assign n6988 = ~n6406 & n38559;
  assign n6989 = n6406 & ~n38559;
  assign n6990 = ~n6988 & ~n6989;
  assign n6991 = ~n6414 & ~n6987;
  assign n6992 = ~n6986 & ~n38666;
  assign n6993 = n4544 & n6785;
  assign n6994 = pi91  & n38631;
  assign n6995 = pi93  & n6800;
  assign n6996 = pi92  & n6802;
  assign n6997 = ~n6995 & ~n6996;
  assign n6998 = ~n6994 & ~n6996;
  assign n6999 = ~n6995 & n6998;
  assign n7000 = ~n6994 & n6997;
  assign n7001 = ~n6993 & n38667;
  assign n7002 = pi20  & ~n7001;
  assign n7003 = pi20  & ~n7002;
  assign n7004 = pi20  & n7001;
  assign n7005 = ~n7001 & ~n7002;
  assign n7006 = ~pi20  & ~n7001;
  assign n7007 = ~n38668 & ~n38669;
  assign n7008 = n6402 & ~n6404;
  assign n7009 = ~n6405 & ~n7008;
  assign n7010 = ~n7007 & n7009;
  assign n7011 = n4453 & n6785;
  assign n7012 = pi90  & n38631;
  assign n7013 = pi92  & n6800;
  assign n7014 = pi91  & n6802;
  assign n7015 = ~n7013 & ~n7014;
  assign n7016 = ~n7012 & ~n7014;
  assign n7017 = ~n7013 & n7016;
  assign n7018 = ~n7012 & n7015;
  assign n7019 = ~n7011 & n38670;
  assign n7020 = pi20  & ~n7019;
  assign n7021 = pi20  & ~n7020;
  assign n7022 = pi20  & n7019;
  assign n7023 = ~n7019 & ~n7020;
  assign n7024 = ~pi20  & ~n7019;
  assign n7025 = ~n38671 & ~n38672;
  assign n7026 = n6393 & n38556;
  assign n7027 = ~n6401 & ~n7026;
  assign n7028 = ~n7025 & n7027;
  assign n7029 = n6389 & ~n6391;
  assign n7030 = ~n6392 & ~n7029;
  assign n7031 = n594 & n6785;
  assign n7032 = pi89  & n38631;
  assign n7033 = pi91  & n6800;
  assign n7034 = pi90  & n6802;
  assign n7035 = ~n7033 & ~n7034;
  assign n7036 = ~n7032 & ~n7034;
  assign n7037 = ~n7033 & n7036;
  assign n7038 = ~n7032 & n7035;
  assign n7039 = ~n7031 & n38673;
  assign n7040 = pi20  & ~n7039;
  assign n7041 = pi20  & ~n7040;
  assign n7042 = pi20  & n7039;
  assign n7043 = ~n7039 & ~n7040;
  assign n7044 = ~pi20  & ~n7039;
  assign n7045 = ~n38674 & ~n38675;
  assign n7046 = n7030 & ~n7045;
  assign n7047 = n3566 & n6785;
  assign n7048 = pi88  & n38631;
  assign n7049 = pi90  & n6800;
  assign n7050 = pi89  & n6802;
  assign n7051 = ~n7049 & ~n7050;
  assign n7052 = ~n7048 & ~n7050;
  assign n7053 = ~n7049 & n7052;
  assign n7054 = ~n7048 & n7051;
  assign n7055 = ~n7047 & n38676;
  assign n7056 = pi20  & ~n7055;
  assign n7057 = pi20  & ~n7056;
  assign n7058 = pi20  & n7055;
  assign n7059 = ~n7055 & ~n7056;
  assign n7060 = ~pi20  & ~n7055;
  assign n7061 = ~n38677 & ~n38678;
  assign n7062 = n6383 & ~n6385;
  assign n7063 = ~n6383 & ~n38553;
  assign n7064 = ~n6384 & n6389;
  assign n7065 = ~n7063 & ~n7064;
  assign n7066 = ~n38553 & ~n7062;
  assign n7067 = ~n7061 & ~n38679;
  assign n7068 = n6374 & n38552;
  assign n7069 = ~n6382 & ~n7068;
  assign n7070 = n3591 & n6785;
  assign n7071 = pi87  & n38631;
  assign n7072 = pi89  & n6800;
  assign n7073 = pi88  & n6802;
  assign n7074 = ~n7072 & ~n7073;
  assign n7075 = ~n7071 & ~n7073;
  assign n7076 = ~n7072 & n7075;
  assign n7077 = ~n7071 & n7074;
  assign n7078 = ~n7070 & n38680;
  assign n7079 = pi20  & ~n7078;
  assign n7080 = pi20  & ~n7079;
  assign n7081 = pi20  & n7078;
  assign n7082 = ~n7078 & ~n7079;
  assign n7083 = ~pi20  & ~n7078;
  assign n7084 = ~n38681 & ~n38682;
  assign n7085 = n7069 & ~n7084;
  assign n7086 = n6365 & n38549;
  assign n7087 = ~n6373 & ~n7086;
  assign n7088 = n3354 & n6785;
  assign n7089 = pi86  & n38631;
  assign n7090 = pi88  & n6800;
  assign n7091 = pi87  & n6802;
  assign n7092 = ~n7090 & ~n7091;
  assign n7093 = ~n7089 & ~n7091;
  assign n7094 = ~n7090 & n7093;
  assign n7095 = ~n7089 & n7092;
  assign n7096 = ~n7088 & n38683;
  assign n7097 = pi20  & ~n7096;
  assign n7098 = pi20  & ~n7097;
  assign n7099 = pi20  & n7096;
  assign n7100 = ~n7096 & ~n7097;
  assign n7101 = ~pi20  & ~n7096;
  assign n7102 = ~n38684 & ~n38685;
  assign n7103 = n7087 & ~n7102;
  assign n7104 = n6356 & n38546;
  assign n7105 = ~n6364 & ~n7104;
  assign n7106 = n636 & n6785;
  assign n7107 = pi85  & n38631;
  assign n7108 = pi87  & n6800;
  assign n7109 = pi86  & n6802;
  assign n7110 = ~n7108 & ~n7109;
  assign n7111 = ~n7107 & ~n7109;
  assign n7112 = ~n7108 & n7111;
  assign n7113 = ~n7107 & n7110;
  assign n7114 = ~n7106 & n38686;
  assign n7115 = pi20  & ~n7114;
  assign n7116 = pi20  & ~n7115;
  assign n7117 = pi20  & n7114;
  assign n7118 = ~n7114 & ~n7115;
  assign n7119 = ~pi20  & ~n7114;
  assign n7120 = ~n38687 & ~n38688;
  assign n7121 = n7105 & ~n7120;
  assign n7122 = n6347 & n38543;
  assign n7123 = ~n6355 & ~n7122;
  assign n7124 = n2779 & n6785;
  assign n7125 = pi84  & n38631;
  assign n7126 = pi86  & n6800;
  assign n7127 = pi85  & n6802;
  assign n7128 = ~n7126 & ~n7127;
  assign n7129 = ~n7125 & ~n7127;
  assign n7130 = ~n7126 & n7129;
  assign n7131 = ~n7125 & n7128;
  assign n7132 = ~n7124 & n38689;
  assign n7133 = pi20  & ~n7132;
  assign n7134 = pi20  & ~n7133;
  assign n7135 = pi20  & n7132;
  assign n7136 = ~n7132 & ~n7133;
  assign n7137 = ~pi20  & ~n7132;
  assign n7138 = ~n38690 & ~n38691;
  assign n7139 = n7123 & ~n7138;
  assign n7140 = n6343 & ~n6345;
  assign n7141 = ~n6346 & ~n7140;
  assign n7142 = n2804 & n6785;
  assign n7143 = pi83  & n38631;
  assign n7144 = pi85  & n6800;
  assign n7145 = pi84  & n6802;
  assign n7146 = ~n7144 & ~n7145;
  assign n7147 = ~n7143 & ~n7145;
  assign n7148 = ~n7144 & n7147;
  assign n7149 = ~n7143 & n7146;
  assign n7150 = ~n7142 & n38692;
  assign n7151 = pi20  & ~n7150;
  assign n7152 = pi20  & ~n7151;
  assign n7153 = pi20  & n7150;
  assign n7154 = ~n7150 & ~n7151;
  assign n7155 = ~pi20  & ~n7150;
  assign n7156 = ~n38693 & ~n38694;
  assign n7157 = n7141 & ~n7156;
  assign n7158 = n6334 & n38540;
  assign n7159 = ~n6342 & ~n7158;
  assign n7160 = n2591 & n6785;
  assign n7161 = pi82  & n38631;
  assign n7162 = pi84  & n6800;
  assign n7163 = pi83  & n6802;
  assign n7164 = ~n7162 & ~n7163;
  assign n7165 = ~n7161 & ~n7163;
  assign n7166 = ~n7162 & n7165;
  assign n7167 = ~n7161 & n7164;
  assign n7168 = ~n7160 & n38695;
  assign n7169 = pi20  & ~n7168;
  assign n7170 = pi20  & ~n7169;
  assign n7171 = pi20  & n7168;
  assign n7172 = ~n7168 & ~n7169;
  assign n7173 = ~pi20  & ~n7168;
  assign n7174 = ~n38696 & ~n38697;
  assign n7175 = n7159 & ~n7174;
  assign n7176 = n6325 & n38537;
  assign n7177 = ~n6333 & ~n7176;
  assign n7178 = n2091 & n6785;
  assign n7179 = pi81  & n38631;
  assign n7180 = pi83  & n6800;
  assign n7181 = pi82  & n6802;
  assign n7182 = ~n7180 & ~n7181;
  assign n7183 = ~n7179 & ~n7181;
  assign n7184 = ~n7180 & n7183;
  assign n7185 = ~n7179 & n7182;
  assign n7186 = ~n7178 & n38698;
  assign n7187 = pi20  & ~n7186;
  assign n7188 = pi20  & ~n7187;
  assign n7189 = pi20  & n7186;
  assign n7190 = ~n7186 & ~n7187;
  assign n7191 = ~pi20  & ~n7186;
  assign n7192 = ~n38699 & ~n38700;
  assign n7193 = n7177 & ~n7192;
  assign n7194 = n2134 & n6785;
  assign n7195 = pi80  & n38631;
  assign n7196 = pi82  & n6800;
  assign n7197 = pi81  & n6802;
  assign n7198 = ~n7196 & ~n7197;
  assign n7199 = ~n7195 & ~n7197;
  assign n7200 = ~n7196 & n7199;
  assign n7201 = ~n7195 & n7198;
  assign n7202 = ~n7194 & n38701;
  assign n7203 = pi20  & ~n7202;
  assign n7204 = pi20  & ~n7203;
  assign n7205 = pi20  & n7202;
  assign n7206 = ~n7202 & ~n7203;
  assign n7207 = ~pi20  & ~n7202;
  assign n7208 = ~n38702 & ~n38703;
  assign n7209 = n6316 & n38534;
  assign n7210 = ~n6316 & n38534;
  assign n7211 = n6316 & ~n38534;
  assign n7212 = ~n7210 & ~n7211;
  assign n7213 = ~n6324 & ~n7209;
  assign n7214 = ~n7208 & ~n38704;
  assign n7215 = n6312 & ~n6314;
  assign n7216 = ~n6315 & ~n7215;
  assign n7217 = n2154 & n6785;
  assign n7218 = pi79  & n38631;
  assign n7219 = pi81  & n6800;
  assign n7220 = pi80  & n6802;
  assign n7221 = ~n7219 & ~n7220;
  assign n7222 = ~n7218 & ~n7220;
  assign n7223 = ~n7219 & n7222;
  assign n7224 = ~n7218 & n7221;
  assign n7225 = ~n7217 & n38705;
  assign n7226 = pi20  & ~n7225;
  assign n7227 = pi20  & ~n7226;
  assign n7228 = pi20  & n7225;
  assign n7229 = ~n7225 & ~n7226;
  assign n7230 = ~pi20  & ~n7225;
  assign n7231 = ~n38706 & ~n38707;
  assign n7232 = n7216 & ~n7231;
  assign n7233 = n2063 & n6785;
  assign n7234 = pi78  & n38631;
  assign n7235 = pi80  & n6800;
  assign n7236 = pi79  & n6802;
  assign n7237 = ~n7235 & ~n7236;
  assign n7238 = ~n7234 & ~n7236;
  assign n7239 = ~n7235 & n7238;
  assign n7240 = ~n7234 & n7237;
  assign n7241 = ~n7233 & n38708;
  assign n7242 = pi20  & ~n7241;
  assign n7243 = pi20  & ~n7242;
  assign n7244 = pi20  & n7241;
  assign n7245 = ~n7241 & ~n7242;
  assign n7246 = ~pi20  & ~n7241;
  assign n7247 = ~n38709 & ~n38710;
  assign n7248 = n6306 & ~n6308;
  assign n7249 = ~n6306 & ~n38531;
  assign n7250 = ~n6307 & n6312;
  assign n7251 = ~n7249 & ~n7250;
  assign n7252 = ~n38531 & ~n7248;
  assign n7253 = ~n7247 & ~n38711;
  assign n7254 = n6302 & ~n6304;
  assign n7255 = ~n6305 & ~n7254;
  assign n7256 = n678 & n6785;
  assign n7257 = pi77  & n38631;
  assign n7258 = pi79  & n6800;
  assign n7259 = pi78  & n6802;
  assign n7260 = ~n7258 & ~n7259;
  assign n7261 = ~n7257 & ~n7259;
  assign n7262 = ~n7258 & n7261;
  assign n7263 = ~n7257 & n7260;
  assign n7264 = ~n7256 & n38712;
  assign n7265 = pi20  & ~n7264;
  assign n7266 = pi20  & ~n7265;
  assign n7267 = pi20  & n7264;
  assign n7268 = ~n7264 & ~n7265;
  assign n7269 = ~pi20  & ~n7264;
  assign n7270 = ~n38713 & ~n38714;
  assign n7271 = n7255 & ~n7270;
  assign n7272 = n1578 & n6785;
  assign n7273 = pi76  & n38631;
  assign n7274 = pi78  & n6800;
  assign n7275 = pi77  & n6802;
  assign n7276 = ~n7274 & ~n7275;
  assign n7277 = ~n7273 & ~n7275;
  assign n7278 = ~n7274 & n7277;
  assign n7279 = ~n7273 & n7276;
  assign n7280 = ~n7272 & n38715;
  assign n7281 = pi20  & ~n7280;
  assign n7282 = pi20  & ~n7281;
  assign n7283 = pi20  & n7280;
  assign n7284 = ~n7280 & ~n7281;
  assign n7285 = ~pi20  & ~n7280;
  assign n7286 = ~n38716 & ~n38717;
  assign n7287 = n6296 & ~n6298;
  assign n7288 = ~n6296 & ~n38530;
  assign n7289 = ~n6297 & n6302;
  assign n7290 = ~n7288 & ~n7289;
  assign n7291 = ~n38530 & ~n7287;
  assign n7292 = ~n7286 & ~n38718;
  assign n7293 = n6287 & n38529;
  assign n7294 = ~n6295 & ~n7293;
  assign n7295 = n1596 & n6785;
  assign n7296 = pi75  & n38631;
  assign n7297 = pi77  & n6800;
  assign n7298 = pi76  & n6802;
  assign n7299 = ~n7297 & ~n7298;
  assign n7300 = ~n7296 & ~n7298;
  assign n7301 = ~n7297 & n7300;
  assign n7302 = ~n7296 & n7299;
  assign n7303 = ~n7295 & n38719;
  assign n7304 = pi20  & ~n7303;
  assign n7305 = pi20  & ~n7304;
  assign n7306 = pi20  & n7303;
  assign n7307 = ~n7303 & ~n7304;
  assign n7308 = ~pi20  & ~n7303;
  assign n7309 = ~n38720 & ~n38721;
  assign n7310 = n7294 & ~n7309;
  assign n7311 = ~n7294 & n7309;
  assign n7312 = ~n7310 & ~n7311;
  assign n7313 = n1465 & n6785;
  assign n7314 = pi74  & n38631;
  assign n7315 = pi76  & n6800;
  assign n7316 = pi75  & n6802;
  assign n7317 = ~n7315 & ~n7316;
  assign n7318 = ~n7314 & ~n7316;
  assign n7319 = ~n7315 & n7318;
  assign n7320 = ~n7314 & n7317;
  assign n7321 = ~n7313 & n38722;
  assign n7322 = pi20  & ~n7321;
  assign n7323 = pi20  & ~n7322;
  assign n7324 = pi20  & n7321;
  assign n7325 = ~n7321 & ~n7322;
  assign n7326 = ~pi20  & ~n7321;
  assign n7327 = ~n38723 & ~n38724;
  assign n7328 = n6283 & ~n6285;
  assign n7329 = ~n6286 & ~n7328;
  assign n7330 = ~n7327 & n7329;
  assign n7331 = n720 & n6785;
  assign n7332 = pi73  & n38631;
  assign n7333 = pi75  & n6800;
  assign n7334 = pi74  & n6802;
  assign n7335 = ~n7333 & ~n7334;
  assign n7336 = ~n7332 & ~n7334;
  assign n7337 = ~n7333 & n7336;
  assign n7338 = ~n7332 & n7335;
  assign n7339 = ~n7331 & n38725;
  assign n7340 = pi20  & ~n7339;
  assign n7341 = pi20  & ~n7340;
  assign n7342 = pi20  & n7339;
  assign n7343 = ~n7339 & ~n7340;
  assign n7344 = ~pi20  & ~n7339;
  assign n7345 = ~n38726 & ~n38727;
  assign n7346 = n6279 & ~n6281;
  assign n7347 = ~n6282 & ~n7346;
  assign n7348 = ~n7345 & n7347;
  assign n7349 = n6275 & ~n6277;
  assign n7350 = ~n6278 & ~n7349;
  assign n7351 = n1218 & n6785;
  assign n7352 = pi72  & n38631;
  assign n7353 = pi74  & n6800;
  assign n7354 = pi73  & n6802;
  assign n7355 = ~n7353 & ~n7354;
  assign n7356 = ~n7352 & ~n7354;
  assign n7357 = ~n7353 & n7356;
  assign n7358 = ~n7352 & n7355;
  assign n7359 = ~n7351 & n38728;
  assign n7360 = pi20  & ~n7359;
  assign n7361 = pi20  & ~n7360;
  assign n7362 = pi20  & n7359;
  assign n7363 = ~n7359 & ~n7360;
  assign n7364 = ~pi20  & ~n7359;
  assign n7365 = ~n38729 & ~n38730;
  assign n7366 = n7350 & ~n7365;
  assign n7367 = n1238 & n6785;
  assign n7368 = pi71  & n38631;
  assign n7369 = pi73  & n6800;
  assign n7370 = pi72  & n6802;
  assign n7371 = ~n7369 & ~n7370;
  assign n7372 = ~n7368 & ~n7370;
  assign n7373 = ~n7369 & n7372;
  assign n7374 = ~n7368 & n7371;
  assign n7375 = ~n7367 & n38731;
  assign n7376 = pi20  & ~n7375;
  assign n7377 = pi20  & ~n7376;
  assign n7378 = pi20  & n7375;
  assign n7379 = ~n7375 & ~n7376;
  assign n7380 = ~pi20  & ~n7375;
  assign n7381 = ~n38732 & ~n38733;
  assign n7382 = n6266 & n38526;
  assign n7383 = ~n6266 & n38526;
  assign n7384 = n6266 & ~n38526;
  assign n7385 = ~n7383 & ~n7384;
  assign n7386 = ~n6274 & ~n7382;
  assign n7387 = ~n7381 & ~n38734;
  assign n7388 = n1124 & n6785;
  assign n7389 = pi70  & n38631;
  assign n7390 = pi72  & n6800;
  assign n7391 = pi71  & n6802;
  assign n7392 = ~n7390 & ~n7391;
  assign n7393 = ~n7389 & ~n7391;
  assign n7394 = ~n7390 & n7393;
  assign n7395 = ~n7389 & n7392;
  assign n7396 = ~n7388 & n38735;
  assign n7397 = pi20  & ~n7396;
  assign n7398 = pi20  & ~n7397;
  assign n7399 = pi20  & n7396;
  assign n7400 = ~n7396 & ~n7397;
  assign n7401 = ~pi20  & ~n7396;
  assign n7402 = ~n38736 & ~n38737;
  assign n7403 = n6260 & ~n6262;
  assign n7404 = ~n6260 & ~n38523;
  assign n7405 = ~n6261 & n6266;
  assign n7406 = ~n7404 & ~n7405;
  assign n7407 = ~n38523 & ~n7403;
  assign n7408 = ~n7402 & ~n38738;
  assign n7409 = n927 & n6785;
  assign n7410 = pi69  & n38631;
  assign n7411 = pi71  & n6800;
  assign n7412 = pi70  & n6802;
  assign n7413 = ~n7411 & ~n7412;
  assign n7414 = ~n7410 & ~n7412;
  assign n7415 = ~n7411 & n7414;
  assign n7416 = ~n7410 & n7413;
  assign n7417 = ~n7409 & n38739;
  assign n7418 = pi20  & ~n7417;
  assign n7419 = pi20  & ~n7418;
  assign n7420 = pi20  & n7417;
  assign n7421 = ~n7417 & ~n7418;
  assign n7422 = ~pi20  & ~n7417;
  assign n7423 = ~n38740 & ~n38741;
  assign n7424 = n6253 & n38522;
  assign n7425 = ~n6259 & ~n7424;
  assign n7426 = ~n7423 & n7425;
  assign n7427 = n6246 & n38521;
  assign n7428 = ~n6252 & ~n7427;
  assign n7429 = n972 & n6785;
  assign n7430 = pi68  & n38631;
  assign n7431 = pi70  & n6800;
  assign n7432 = pi69  & n6802;
  assign n7433 = ~n7431 & ~n7432;
  assign n7434 = ~n7430 & ~n7432;
  assign n7435 = ~n7431 & n7434;
  assign n7436 = ~n7430 & n7433;
  assign n7437 = ~n7429 & n38742;
  assign n7438 = pi20  & ~n7437;
  assign n7439 = pi20  & ~n7438;
  assign n7440 = pi20  & n7437;
  assign n7441 = ~n7437 & ~n7438;
  assign n7442 = ~pi20  & ~n7437;
  assign n7443 = ~n38743 & ~n38744;
  assign n7444 = n7428 & ~n7443;
  assign n7445 = n990 & n6785;
  assign n7446 = pi67  & n38631;
  assign n7447 = pi69  & n6800;
  assign n7448 = pi68  & n6802;
  assign n7449 = ~n7447 & ~n7448;
  assign n7450 = ~n7446 & ~n7448;
  assign n7451 = ~n7447 & n7450;
  assign n7452 = ~n7446 & n7449;
  assign n7453 = ~n7445 & n38745;
  assign n7454 = pi20  & ~n7453;
  assign n7455 = pi20  & ~n7454;
  assign n7456 = pi20  & n7453;
  assign n7457 = ~n7453 & ~n7454;
  assign n7458 = ~pi20  & ~n7453;
  assign n7459 = ~n38746 & ~n38747;
  assign n7460 = pi23  & ~n38513;
  assign n7461 = n38516 & ~n7460;
  assign n7462 = ~n38516 & n7460;
  assign n7463 = ~n38513 & n6228;
  assign n7464 = ~n38517 & ~n7463;
  assign n7465 = ~n7461 & ~n7462;
  assign n7466 = ~n7459 & n38748;
  assign n7467 = n871 & n6785;
  assign n7468 = pi66  & n38631;
  assign n7469 = pi68  & n6800;
  assign n7470 = pi67  & n6802;
  assign n7471 = ~n7469 & ~n7470;
  assign n7472 = ~n7468 & ~n7470;
  assign n7473 = ~n7469 & n7472;
  assign n7474 = ~n7468 & n7471;
  assign n7475 = ~n7467 & n38749;
  assign n7476 = pi20  & ~n7475;
  assign n7477 = pi20  & ~n7476;
  assign n7478 = pi20  & n7475;
  assign n7479 = ~n7475 & ~n7476;
  assign n7480 = ~pi20  & ~n7475;
  assign n7481 = ~n38750 & ~n38751;
  assign n7482 = pi23  & n6202;
  assign n7483 = ~n6201 & n7482;
  assign n7484 = n6201 & ~n7482;
  assign n7485 = ~n6203 & n6207;
  assign n7486 = ~n38513 & ~n7485;
  assign n7487 = ~n7483 & ~n7484;
  assign n7488 = ~n7481 & n38752;
  assign n7489 = n37515 & n6785;
  assign n7490 = pi65  & n6800;
  assign n7491 = pi64  & n6802;
  assign n7492 = ~n7490 & ~n7491;
  assign n7493 = ~n7489 & n7492;
  assign n7494 = pi64  & n38628;
  assign n7495 = pi20  & ~n7494;
  assign n7496 = pi20  & ~n7493;
  assign n7497 = pi20  & ~n7496;
  assign n7498 = ~n7493 & ~n7496;
  assign n7499 = ~n7497 & ~n7498;
  assign n7500 = n7495 & ~n7499;
  assign n7501 = n7493 & n7495;
  assign n7502 = pi64  & n38631;
  assign n7503 = pi65  & n6802;
  assign n7504 = ~n37521 & n6785;
  assign n7505 = pi66  & n6800;
  assign n7506 = ~n7504 & ~n7505;
  assign n7507 = ~n7503 & ~n7504;
  assign n7508 = ~n7505 & n7507;
  assign n7509 = ~n7503 & ~n7505;
  assign n7510 = ~n7504 & n7509;
  assign n7511 = ~n7503 & n7506;
  assign n7512 = ~n7502 & ~n7503;
  assign n7513 = ~n7505 & n7512;
  assign n7514 = ~n7502 & n7509;
  assign n7515 = ~n7504 & n38755;
  assign n7516 = ~n7502 & n38754;
  assign n7517 = pi20  & ~n38756;
  assign n7518 = pi20  & ~n7517;
  assign n7519 = ~n38756 & ~n7517;
  assign n7520 = ~n7518 & ~n7519;
  assign n7521 = n38753 & ~n7520;
  assign n7522 = n38753 & n38756;
  assign n7523 = n6202 & n38757;
  assign n7524 = n847 & n6785;
  assign n7525 = pi65  & n38631;
  assign n7526 = pi67  & n6800;
  assign n7527 = pi66  & n6802;
  assign n7528 = ~n7526 & ~n7527;
  assign n7529 = ~n7525 & ~n7527;
  assign n7530 = ~n7526 & n7529;
  assign n7531 = ~n7525 & n7528;
  assign n7532 = ~n7524 & n38758;
  assign n7533 = pi20  & ~n7532;
  assign n7534 = pi20  & ~n7533;
  assign n7535 = pi20  & n7532;
  assign n7536 = ~n7532 & ~n7533;
  assign n7537 = ~pi20  & ~n7532;
  assign n7538 = ~n38759 & ~n38760;
  assign n7539 = ~n6202 & ~n38757;
  assign n7540 = n6202 & ~n38757;
  assign n7541 = ~n6202 & n38757;
  assign n7542 = ~n7540 & ~n7541;
  assign n7543 = ~n7523 & ~n7539;
  assign n7544 = ~n7538 & ~n38761;
  assign n7545 = ~n7523 & ~n7544;
  assign n7546 = n7481 & ~n38752;
  assign n7547 = n7481 & n38752;
  assign n7548 = ~n7481 & ~n38752;
  assign n7549 = ~n7547 & ~n7548;
  assign n7550 = ~n7488 & ~n7546;
  assign n7551 = ~n7545 & ~n38762;
  assign n7552 = ~n7488 & ~n7551;
  assign n7553 = n7459 & ~n38748;
  assign n7554 = ~n7466 & ~n7553;
  assign n7555 = ~n7552 & ~n7553;
  assign n7556 = ~n7466 & n7555;
  assign n7557 = ~n7552 & n7554;
  assign n7558 = ~n7466 & ~n38763;
  assign n7559 = ~n7428 & n7443;
  assign n7560 = n7428 & ~n7444;
  assign n7561 = n7428 & n7443;
  assign n7562 = ~n7443 & ~n7444;
  assign n7563 = ~n7428 & ~n7443;
  assign n7564 = ~n38764 & ~n38765;
  assign n7565 = ~n7444 & ~n7559;
  assign n7566 = ~n7558 & ~n38766;
  assign n7567 = ~n7444 & ~n7566;
  assign n7568 = n7423 & ~n7425;
  assign n7569 = ~n7426 & ~n7568;
  assign n7570 = ~n7567 & n7569;
  assign n7571 = ~n7426 & ~n7570;
  assign n7572 = n7402 & n38738;
  assign n7573 = ~n7408 & ~n7572;
  assign n7574 = ~n7571 & n7573;
  assign n7575 = ~n7408 & ~n7574;
  assign n7576 = n7381 & n38734;
  assign n7577 = ~n7387 & ~n7576;
  assign n7578 = ~n7575 & n7577;
  assign n7579 = ~n7387 & ~n7578;
  assign n7580 = ~n7350 & n7365;
  assign n7581 = n7350 & ~n7366;
  assign n7582 = n7350 & n7365;
  assign n7583 = ~n7365 & ~n7366;
  assign n7584 = ~n7350 & ~n7365;
  assign n7585 = ~n38767 & ~n38768;
  assign n7586 = ~n7366 & ~n7580;
  assign n7587 = ~n7579 & ~n38769;
  assign n7588 = ~n7366 & ~n7587;
  assign n7589 = n7345 & ~n7347;
  assign n7590 = ~n7348 & ~n7589;
  assign n7591 = ~n7588 & n7590;
  assign n7592 = ~n7348 & ~n7591;
  assign n7593 = n7327 & ~n7329;
  assign n7594 = ~n7330 & ~n7593;
  assign n7595 = ~n7592 & n7594;
  assign n7596 = ~n7330 & ~n7595;
  assign n7597 = n7312 & ~n7596;
  assign n7598 = ~n7310 & ~n7597;
  assign n7599 = n7286 & n38718;
  assign n7600 = ~n7292 & ~n7599;
  assign n7601 = ~n7598 & n7600;
  assign n7602 = ~n7292 & ~n7601;
  assign n7603 = ~n7255 & n7270;
  assign n7604 = n7255 & ~n7271;
  assign n7605 = n7255 & n7270;
  assign n7606 = ~n7270 & ~n7271;
  assign n7607 = ~n7255 & ~n7270;
  assign n7608 = ~n38770 & ~n38771;
  assign n7609 = ~n7271 & ~n7603;
  assign n7610 = ~n7602 & ~n38772;
  assign n7611 = ~n7271 & ~n7610;
  assign n7612 = n7247 & n38711;
  assign n7613 = ~n38711 & ~n7253;
  assign n7614 = n7247 & ~n38711;
  assign n7615 = ~n7247 & ~n7253;
  assign n7616 = ~n7247 & n38711;
  assign n7617 = ~n38773 & ~n38774;
  assign n7618 = ~n7253 & ~n7612;
  assign n7619 = ~n7611 & ~n38775;
  assign n7620 = ~n7253 & ~n7619;
  assign n7621 = ~n7216 & n7231;
  assign n7622 = n7216 & ~n7232;
  assign n7623 = n7216 & n7231;
  assign n7624 = ~n7231 & ~n7232;
  assign n7625 = ~n7216 & ~n7231;
  assign n7626 = ~n38776 & ~n38777;
  assign n7627 = ~n7232 & ~n7621;
  assign n7628 = ~n7620 & ~n38778;
  assign n7629 = ~n7232 & ~n7628;
  assign n7630 = n7208 & n38704;
  assign n7631 = ~n7214 & ~n7630;
  assign n7632 = ~n7629 & n7631;
  assign n7633 = ~n7214 & ~n7632;
  assign n7634 = ~n7177 & n7192;
  assign n7635 = n7177 & ~n7193;
  assign n7636 = n7177 & n7192;
  assign n7637 = ~n7192 & ~n7193;
  assign n7638 = ~n7177 & ~n7192;
  assign n7639 = ~n38779 & ~n38780;
  assign n7640 = ~n7193 & ~n7634;
  assign n7641 = ~n7633 & ~n38781;
  assign n7642 = ~n7193 & ~n7641;
  assign n7643 = ~n7159 & n7174;
  assign n7644 = n7159 & ~n7175;
  assign n7645 = n7159 & n7174;
  assign n7646 = ~n7174 & ~n7175;
  assign n7647 = ~n7159 & ~n7174;
  assign n7648 = ~n38782 & ~n38783;
  assign n7649 = ~n7175 & ~n7643;
  assign n7650 = ~n7642 & ~n38784;
  assign n7651 = ~n7175 & ~n7650;
  assign n7652 = ~n7141 & n7156;
  assign n7653 = n7141 & ~n7157;
  assign n7654 = n7141 & n7156;
  assign n7655 = ~n7156 & ~n7157;
  assign n7656 = ~n7141 & ~n7156;
  assign n7657 = ~n38785 & ~n38786;
  assign n7658 = ~n7157 & ~n7652;
  assign n7659 = ~n7651 & ~n38787;
  assign n7660 = ~n7157 & ~n7659;
  assign n7661 = ~n7123 & n7138;
  assign n7662 = n7123 & ~n7139;
  assign n7663 = n7123 & n7138;
  assign n7664 = ~n7138 & ~n7139;
  assign n7665 = ~n7123 & ~n7138;
  assign n7666 = ~n38788 & ~n38789;
  assign n7667 = ~n7139 & ~n7661;
  assign n7668 = ~n7660 & ~n38790;
  assign n7669 = ~n7139 & ~n7668;
  assign n7670 = ~n7105 & n7120;
  assign n7671 = ~n7121 & ~n7670;
  assign n7672 = ~n7669 & ~n7670;
  assign n7673 = ~n7121 & n7672;
  assign n7674 = ~n7669 & n7671;
  assign n7675 = ~n7121 & ~n38791;
  assign n7676 = ~n7087 & n7102;
  assign n7677 = ~n7103 & ~n7676;
  assign n7678 = ~n7675 & n7677;
  assign n7679 = ~n7103 & ~n7678;
  assign n7680 = ~n7069 & n7084;
  assign n7681 = n7069 & ~n7085;
  assign n7682 = n7069 & n7084;
  assign n7683 = ~n7084 & ~n7085;
  assign n7684 = ~n7069 & ~n7084;
  assign n7685 = ~n38792 & ~n38793;
  assign n7686 = ~n7085 & ~n7680;
  assign n7687 = ~n7679 & ~n38794;
  assign n7688 = ~n7085 & ~n7687;
  assign n7689 = n7061 & n38679;
  assign n7690 = ~n7067 & ~n7689;
  assign n7691 = ~n7688 & n7690;
  assign n7692 = ~n7067 & ~n7691;
  assign n7693 = ~n7030 & n7045;
  assign n7694 = n7030 & ~n7046;
  assign n7695 = n7030 & n7045;
  assign n7696 = ~n7045 & ~n7046;
  assign n7697 = ~n7030 & ~n7045;
  assign n7698 = ~n38795 & ~n38796;
  assign n7699 = ~n7046 & ~n7693;
  assign n7700 = ~n7692 & ~n38797;
  assign n7701 = ~n7046 & ~n7700;
  assign n7702 = n7025 & ~n7027;
  assign n7703 = ~n7025 & ~n7028;
  assign n7704 = ~n7025 & ~n7027;
  assign n7705 = n7027 & ~n7028;
  assign n7706 = n7025 & n7027;
  assign n7707 = ~n38798 & ~n38799;
  assign n7708 = ~n7028 & ~n7702;
  assign n7709 = ~n7701 & ~n38800;
  assign n7710 = ~n7028 & ~n7709;
  assign n7711 = n7007 & ~n7009;
  assign n7712 = ~n7010 & ~n7711;
  assign n7713 = ~n7710 & n7712;
  assign n7714 = ~n7010 & ~n7713;
  assign n7715 = n6986 & n38666;
  assign n7716 = ~n6992 & ~n7715;
  assign n7717 = ~n7714 & n7716;
  assign n7718 = ~n6992 & ~n7717;
  assign n7719 = n6963 & n38662;
  assign n7720 = ~n38662 & ~n6971;
  assign n7721 = ~n6963 & ~n6971;
  assign n7722 = ~n7720 & ~n7721;
  assign n7723 = ~n6971 & ~n7719;
  assign n7724 = ~n7718 & ~n38801;
  assign n7725 = ~n6971 & ~n7724;
  assign n7726 = n6945 & ~n6947;
  assign n7727 = ~n6948 & ~n7726;
  assign n7728 = ~n7725 & n7727;
  assign n7729 = ~n6948 & ~n7728;
  assign n7730 = ~n6914 & n6929;
  assign n7731 = n6914 & ~n6930;
  assign n7732 = n6914 & n6929;
  assign n7733 = ~n6929 & ~n6930;
  assign n7734 = ~n6914 & ~n6929;
  assign n7735 = ~n38802 & ~n38803;
  assign n7736 = ~n6930 & ~n7730;
  assign n7737 = ~n7729 & ~n38804;
  assign n7738 = ~n6930 & ~n7737;
  assign n7739 = ~n6896 & n6911;
  assign n7740 = n6896 & ~n6912;
  assign n7741 = n6896 & n6911;
  assign n7742 = ~n6911 & ~n6912;
  assign n7743 = ~n6896 & ~n6911;
  assign n7744 = ~n38805 & ~n38806;
  assign n7745 = ~n6912 & ~n7739;
  assign n7746 = ~n7738 & ~n38807;
  assign n7747 = ~n6912 & ~n7746;
  assign n7748 = ~n6878 & n6893;
  assign n7749 = n6878 & ~n6894;
  assign n7750 = n6878 & n6893;
  assign n7751 = ~n6893 & ~n6894;
  assign n7752 = ~n6878 & ~n6893;
  assign n7753 = ~n38808 & ~n38809;
  assign n7754 = ~n6894 & ~n7748;
  assign n7755 = ~n7747 & ~n38810;
  assign n7756 = ~n6894 & ~n7755;
  assign n7757 = n6870 & n38644;
  assign n7758 = ~n6876 & ~n7757;
  assign n7759 = ~n7756 & n7758;
  assign n7760 = ~n6876 & ~n7759;
  assign n7761 = ~n6837 & n6854;
  assign n7762 = n6837 & ~n6855;
  assign n7763 = n6837 & n6854;
  assign n7764 = ~n6854 & ~n6855;
  assign n7765 = ~n6837 & ~n6854;
  assign n7766 = ~n38811 & ~n38812;
  assign n7767 = ~n6855 & ~n7761;
  assign n7768 = ~n7760 & ~n38813;
  assign n7769 = ~n6855 & ~n7768;
  assign n7770 = ~n6817 & n6834;
  assign n7771 = n6817 & ~n6835;
  assign n7772 = n6817 & n6834;
  assign n7773 = ~n6834 & ~n6835;
  assign n7774 = ~n6817 & ~n6834;
  assign n7775 = ~n38814 & ~n38815;
  assign n7776 = ~n6835 & ~n7770;
  assign n7777 = ~n7769 & ~n38816;
  assign n7778 = ~n6835 & ~n7777;
  assign n7779 = ~n6772 & n6814;
  assign n7780 = n6772 & ~n6815;
  assign n7781 = n6772 & n6814;
  assign n7782 = ~n6814 & ~n6815;
  assign n7783 = ~n6772 & ~n6814;
  assign n7784 = ~n38817 & ~n38818;
  assign n7785 = ~n6815 & ~n7779;
  assign n7786 = ~n7778 & ~n38819;
  assign n7787 = ~n6815 & ~n7786;
  assign n7788 = ~n6767 & ~n6771;
  assign n7789 = ~n6753 & ~n6761;
  assign n7790 = ~n6732 & ~n6735;
  assign n7791 = n607 & n4494;
  assign n7792 = pi93  & n37489;
  assign n7793 = pi95  & n620;
  assign n7794 = pi94  & n622;
  assign n7795 = ~n7793 & ~n7794;
  assign n7796 = ~n7792 & ~n7794;
  assign n7797 = ~n7793 & n7796;
  assign n7798 = ~n7792 & n7795;
  assign n7799 = ~n7791 & n38820;
  assign n7800 = pi29  & ~n7799;
  assign n7801 = pi29  & ~n7800;
  assign n7802 = pi29  & n7799;
  assign n7803 = ~n7799 & ~n7800;
  assign n7804 = ~pi29  & ~n7799;
  assign n7805 = ~n38821 & ~n38822;
  assign n7806 = ~n6727 & ~n6729;
  assign n7807 = ~n6700 & ~n6709;
  assign n7808 = ~n6679 & ~n6682;
  assign n7809 = n691 & n2779;
  assign n7810 = pi84  & n37503;
  assign n7811 = pi86  & n704;
  assign n7812 = pi85  & n706;
  assign n7813 = ~n7811 & ~n7812;
  assign n7814 = ~n7810 & ~n7812;
  assign n7815 = ~n7811 & n7814;
  assign n7816 = ~n7810 & n7813;
  assign n7817 = ~n7809 & n38823;
  assign n7818 = pi38  & ~n7817;
  assign n7819 = pi38  & ~n7818;
  assign n7820 = pi38  & n7817;
  assign n7821 = ~n7817 & ~n7818;
  assign n7822 = ~pi38  & ~n7817;
  assign n7823 = ~n38824 & ~n38825;
  assign n7824 = ~n6666 & ~n6674;
  assign n7825 = ~n6660 & ~n6663;
  assign n7826 = n940 & n2063;
  assign n7827 = pi78  & n37541;
  assign n7828 = pi80  & n953;
  assign n7829 = pi79  & n955;
  assign n7830 = ~n7828 & ~n7829;
  assign n7831 = ~n7827 & ~n7829;
  assign n7832 = ~n7828 & n7831;
  assign n7833 = ~n7827 & n7830;
  assign n7834 = ~n7826 & n38826;
  assign n7835 = pi44  & ~n7834;
  assign n7836 = pi44  & ~n7835;
  assign n7837 = pi44  & n7834;
  assign n7838 = ~n7834 & ~n7835;
  assign n7839 = ~pi44  & ~n7834;
  assign n7840 = ~n38827 & ~n38828;
  assign n7841 = ~n6655 & ~n6657;
  assign n7842 = ~n6648 & ~n6651;
  assign n7843 = ~n6634 & ~n6642;
  assign n7844 = n927 & n1971;
  assign n7845 = pi69  & n37864;
  assign n7846 = pi71  & n1973;
  assign n7847 = pi70  & n1981;
  assign n7848 = ~n7846 & ~n7847;
  assign n7849 = ~n7845 & ~n7847;
  assign n7850 = ~n7846 & n7849;
  assign n7851 = ~n7845 & n7848;
  assign n7852 = ~n7844 & n38829;
  assign n7853 = pi53  & ~n7852;
  assign n7854 = pi53  & ~n7853;
  assign n7855 = pi53  & n7852;
  assign n7856 = ~n7852 & ~n7853;
  assign n7857 = ~pi53  & ~n7852;
  assign n7858 = ~n38830 & ~n38831;
  assign n7859 = ~n6610 & ~n6616;
  assign n7860 = n871 & n4312;
  assign n7861 = pi66  & n38376;
  assign n7862 = pi68  & n4314;
  assign n7863 = pi67  & n4322;
  assign n7864 = ~n7862 & ~n7863;
  assign n7865 = ~n7861 & ~n7863;
  assign n7866 = ~n7862 & n7865;
  assign n7867 = ~n7861 & n7864;
  assign n7868 = ~n7860 & n38832;
  assign n7869 = pi56  & ~n7868;
  assign n7870 = pi56  & ~n7869;
  assign n7871 = pi56  & n7868;
  assign n7872 = ~n7868 & ~n7869;
  assign n7873 = ~pi56  & ~n7868;
  assign n7874 = ~n38833 & ~n38834;
  assign n7875 = pi59  & n6609;
  assign n7876 = pi58  & ~pi59 ;
  assign n7877 = ~pi58  & pi59 ;
  assign n7878 = ~pi58  & ~pi59 ;
  assign n7879 = pi58  & pi59 ;
  assign n7880 = ~n7878 & ~n7879;
  assign n7881 = ~n7876 & ~n7877;
  assign n7882 = n38599 & n38835;
  assign n7883 = n37515 & n7882;
  assign n7884 = n38599 & ~n38835;
  assign n7885 = pi65  & n7884;
  assign n7886 = pi57  & ~pi58 ;
  assign n7887 = ~pi57  & pi58 ;
  assign n7888 = ~pi57  & ~pi58 ;
  assign n7889 = pi57  & pi58 ;
  assign n7890 = ~n7888 & ~n7889;
  assign n7891 = ~n7886 & ~n7887;
  assign n7892 = ~n38599 & n38836;
  assign n7893 = pi64  & n7892;
  assign n7894 = ~n7885 & ~n7893;
  assign n7895 = ~n7883 & n7894;
  assign n7896 = n7875 & ~n7895;
  assign n7897 = ~n7875 & n7895;
  assign n7898 = pi59  & ~n6609;
  assign n7899 = pi59  & ~n7895;
  assign n7900 = pi59  & ~n7899;
  assign n7901 = ~n7895 & ~n7899;
  assign n7902 = ~n7900 & ~n7901;
  assign n7903 = n7898 & ~n7902;
  assign n7904 = n7895 & n7898;
  assign n7905 = ~n7898 & n7902;
  assign n7906 = ~n38837 & ~n7905;
  assign n7907 = ~n7896 & ~n7897;
  assign n7908 = n7874 & ~n38838;
  assign n7909 = ~n7874 & n38838;
  assign n7910 = ~n7908 & ~n7909;
  assign n7911 = ~n7859 & n7910;
  assign n7912 = n7859 & ~n7910;
  assign n7913 = ~n7911 & ~n7912;
  assign n7914 = n7858 & ~n7913;
  assign n7915 = ~n7858 & n7913;
  assign n7916 = ~n7914 & ~n7915;
  assign n7917 = ~n7843 & n7916;
  assign n7918 = n7843 & ~n7916;
  assign n7919 = ~n7917 & ~n7918;
  assign n7920 = n894 & n1218;
  assign n7921 = pi72  & n37580;
  assign n7922 = pi74  & n896;
  assign n7923 = pi73  & n904;
  assign n7924 = ~n7922 & ~n7923;
  assign n7925 = ~n7921 & ~n7923;
  assign n7926 = ~n7922 & n7925;
  assign n7927 = ~n7921 & n7924;
  assign n7928 = ~n7920 & n38839;
  assign n7929 = pi50  & ~n7928;
  assign n7930 = pi50  & ~n7929;
  assign n7931 = pi50  & n7928;
  assign n7932 = ~n7928 & ~n7929;
  assign n7933 = ~pi50  & ~n7928;
  assign n7934 = ~n38840 & ~n38841;
  assign n7935 = n7919 & ~n7934;
  assign n7936 = ~n7919 & n7934;
  assign n7937 = n7919 & ~n7935;
  assign n7938 = n7919 & n7934;
  assign n7939 = ~n7934 & ~n7935;
  assign n7940 = ~n7919 & ~n7934;
  assign n7941 = ~n38842 & ~n38843;
  assign n7942 = ~n7935 & ~n7936;
  assign n7943 = n7842 & n38844;
  assign n7944 = ~n7842 & ~n38844;
  assign n7945 = ~n7943 & ~n7944;
  assign n7946 = n785 & n1596;
  assign n7947 = pi75  & n37520;
  assign n7948 = pi77  & n787;
  assign n7949 = pi76  & n795;
  assign n7950 = ~n7948 & ~n7949;
  assign n7951 = ~n7947 & ~n7949;
  assign n7952 = ~n7948 & n7951;
  assign n7953 = ~n7947 & n7950;
  assign n7954 = ~n7946 & n38845;
  assign n7955 = pi47  & ~n7954;
  assign n7956 = pi47  & ~n7955;
  assign n7957 = pi47  & n7954;
  assign n7958 = ~n7954 & ~n7955;
  assign n7959 = ~pi47  & ~n7954;
  assign n7960 = ~n38846 & ~n38847;
  assign n7961 = n7945 & ~n7960;
  assign n7962 = ~n7945 & n7960;
  assign n7963 = ~n7961 & ~n7962;
  assign n7964 = ~n7841 & ~n7962;
  assign n7965 = ~n7961 & n7964;
  assign n7966 = ~n7841 & n7963;
  assign n7967 = n7841 & ~n7963;
  assign n7968 = ~n7841 & ~n38848;
  assign n7969 = ~n7961 & ~n38848;
  assign n7970 = ~n7962 & n7969;
  assign n7971 = ~n7968 & ~n7970;
  assign n7972 = ~n38848 & ~n7967;
  assign n7973 = ~n7840 & ~n38849;
  assign n7974 = n7840 & n38849;
  assign n7975 = ~n38849 & ~n7973;
  assign n7976 = n7840 & ~n38849;
  assign n7977 = ~n7840 & ~n7973;
  assign n7978 = ~n7840 & n38849;
  assign n7979 = ~n38850 & ~n38851;
  assign n7980 = ~n7973 & ~n7974;
  assign n7981 = n7825 & n38852;
  assign n7982 = ~n7825 & ~n38852;
  assign n7983 = ~n7981 & ~n7982;
  assign n7984 = n733 & n2091;
  assign n7985 = pi81  & n37510;
  assign n7986 = pi83  & n746;
  assign n7987 = pi82  & n748;
  assign n7988 = ~n7986 & ~n7987;
  assign n7989 = ~n7985 & ~n7987;
  assign n7990 = ~n7986 & n7989;
  assign n7991 = ~n7985 & n7988;
  assign n7992 = ~n7984 & n38853;
  assign n7993 = pi41  & ~n7992;
  assign n7994 = pi41  & ~n7993;
  assign n7995 = pi41  & n7992;
  assign n7996 = ~n7992 & ~n7993;
  assign n7997 = ~pi41  & ~n7992;
  assign n7998 = ~n38854 & ~n38855;
  assign n7999 = n7983 & ~n7998;
  assign n8000 = ~n7983 & n7998;
  assign n8001 = ~n7999 & ~n8000;
  assign n8002 = ~n7824 & ~n8000;
  assign n8003 = ~n7999 & n8002;
  assign n8004 = ~n7824 & n8001;
  assign n8005 = n7824 & ~n8001;
  assign n8006 = ~n7824 & ~n38856;
  assign n8007 = ~n7999 & ~n38856;
  assign n8008 = ~n8000 & n8007;
  assign n8009 = ~n8006 & ~n8008;
  assign n8010 = ~n38856 & ~n8005;
  assign n8011 = ~n7823 & ~n38857;
  assign n8012 = n7823 & n38857;
  assign n8013 = ~n38857 & ~n8011;
  assign n8014 = n7823 & ~n38857;
  assign n8015 = ~n7823 & ~n8011;
  assign n8016 = ~n7823 & n38857;
  assign n8017 = ~n38858 & ~n38859;
  assign n8018 = ~n8011 & ~n8012;
  assign n8019 = n7808 & n38860;
  assign n8020 = ~n7808 & ~n38860;
  assign n8021 = ~n8019 & ~n8020;
  assign n8022 = n2104 & n3591;
  assign n8023 = pi87  & n37758;
  assign n8024 = pi89  & n2117;
  assign n8025 = pi88  & n2119;
  assign n8026 = ~n8024 & ~n8025;
  assign n8027 = ~n8023 & ~n8025;
  assign n8028 = ~n8024 & n8027;
  assign n8029 = ~n8023 & n8026;
  assign n8030 = ~n8022 & n38861;
  assign n8031 = pi35  & ~n8030;
  assign n8032 = pi35  & ~n8031;
  assign n8033 = pi35  & n8030;
  assign n8034 = ~n8030 & ~n8031;
  assign n8035 = ~pi35  & ~n8030;
  assign n8036 = ~n38862 & ~n38863;
  assign n8037 = n8021 & ~n8036;
  assign n8038 = ~n8021 & n8036;
  assign n8039 = n8021 & ~n8037;
  assign n8040 = n8021 & n8036;
  assign n8041 = ~n8036 & ~n8037;
  assign n8042 = ~n8021 & ~n8036;
  assign n8043 = ~n38864 & ~n38865;
  assign n8044 = ~n8037 & ~n8038;
  assign n8045 = n7807 & n38866;
  assign n8046 = ~n7807 & ~n38866;
  assign n8047 = ~n8045 & ~n8046;
  assign n8048 = n649 & n4453;
  assign n8049 = pi90  & n37496;
  assign n8050 = pi92  & n662;
  assign n8051 = pi91  & n664;
  assign n8052 = ~n8050 & ~n8051;
  assign n8053 = ~n8049 & ~n8051;
  assign n8054 = ~n8050 & n8053;
  assign n8055 = ~n8049 & n8052;
  assign n8056 = ~n8048 & n38867;
  assign n8057 = pi32  & ~n8056;
  assign n8058 = pi32  & ~n8057;
  assign n8059 = pi32  & n8056;
  assign n8060 = ~n8056 & ~n8057;
  assign n8061 = ~pi32  & ~n8056;
  assign n8062 = ~n38868 & ~n38869;
  assign n8063 = n8047 & ~n8062;
  assign n8064 = ~n8047 & n8062;
  assign n8065 = n8047 & ~n8063;
  assign n8066 = n8047 & n8062;
  assign n8067 = ~n8062 & ~n8063;
  assign n8068 = ~n8047 & ~n8062;
  assign n8069 = ~n38870 & ~n38871;
  assign n8070 = ~n8063 & ~n8064;
  assign n8071 = ~n7806 & ~n38872;
  assign n8072 = n7806 & n38872;
  assign n8073 = ~n7806 & n38872;
  assign n8074 = n7806 & ~n38872;
  assign n8075 = ~n8073 & ~n8074;
  assign n8076 = ~n8071 & ~n8072;
  assign n8077 = ~n7805 & ~n38873;
  assign n8078 = n7805 & n38873;
  assign n8079 = ~n8077 & ~n8078;
  assign n8080 = n7790 & ~n8079;
  assign n8081 = ~n7790 & n8079;
  assign n8082 = ~n8080 & ~n8081;
  assign n8083 = n4492 & n5610;
  assign n8084 = pi96  & n38208;
  assign n8085 = pi98  & n4507;
  assign n8086 = pi97  & n4509;
  assign n8087 = ~n8085 & ~n8086;
  assign n8088 = ~n8084 & ~n8086;
  assign n8089 = ~n8085 & n8088;
  assign n8090 = ~n8084 & n8087;
  assign n8091 = ~n8083 & n38874;
  assign n8092 = pi26  & ~n8091;
  assign n8093 = pi26  & ~n8092;
  assign n8094 = pi26  & n8091;
  assign n8095 = ~n8091 & ~n8092;
  assign n8096 = ~pi26  & ~n8091;
  assign n8097 = ~n38875 & ~n38876;
  assign n8098 = n8082 & ~n8097;
  assign n8099 = ~n8082 & n8097;
  assign n8100 = n8082 & ~n8098;
  assign n8101 = n8082 & n8097;
  assign n8102 = ~n8097 & ~n8098;
  assign n8103 = ~n8082 & ~n8097;
  assign n8104 = ~n38877 & ~n38878;
  assign n8105 = ~n8098 & ~n8099;
  assign n8106 = n7789 & n38879;
  assign n8107 = ~n7789 & ~n38879;
  assign n8108 = ~n8106 & ~n8107;
  assign n8109 = n5576 & n6839;
  assign n8110 = pi99  & n38406;
  assign n8111 = pi101  & n5591;
  assign n8112 = pi100  & n5593;
  assign n8113 = ~n8111 & ~n8112;
  assign n8114 = ~n8110 & ~n8112;
  assign n8115 = ~n8111 & n8114;
  assign n8116 = ~n8110 & n8113;
  assign n8117 = ~n8109 & n38880;
  assign n8118 = pi23  & ~n8117;
  assign n8119 = pi23  & ~n8118;
  assign n8120 = pi23  & n8117;
  assign n8121 = ~n8117 & ~n8118;
  assign n8122 = ~pi23  & ~n8117;
  assign n8123 = ~n38881 & ~n38882;
  assign n8124 = n8108 & ~n8123;
  assign n8125 = ~n8108 & n8123;
  assign n8126 = n8108 & ~n8124;
  assign n8127 = n8108 & n8123;
  assign n8128 = ~n8123 & ~n8124;
  assign n8129 = ~n8108 & ~n8123;
  assign n8130 = ~n38883 & ~n38884;
  assign n8131 = ~n8124 & ~n8125;
  assign n8132 = n7788 & n38885;
  assign n8133 = ~n7788 & ~n38885;
  assign n8134 = ~n8132 & ~n8133;
  assign n8135 = n473 & ~n475;
  assign n8136 = ~n476 & ~n8135;
  assign n8137 = n6785 & n8136;
  assign n8138 = pi102  & n38631;
  assign n8139 = pi104  & n6800;
  assign n8140 = pi103  & n6802;
  assign n8141 = ~n8139 & ~n8140;
  assign n8142 = ~n8138 & ~n8140;
  assign n8143 = ~n8139 & n8142;
  assign n8144 = ~n8138 & n8141;
  assign n8145 = ~n8137 & n38886;
  assign n8146 = pi20  & ~n8145;
  assign n8147 = pi20  & ~n8146;
  assign n8148 = pi20  & n8145;
  assign n8149 = ~n8145 & ~n8146;
  assign n8150 = ~pi20  & ~n8145;
  assign n8151 = ~n38887 & ~n38888;
  assign n8152 = n8134 & ~n8151;
  assign n8153 = ~n8134 & n8151;
  assign n8154 = n8134 & ~n8152;
  assign n8155 = n8134 & n8151;
  assign n8156 = ~n8151 & ~n8152;
  assign n8157 = ~n8134 & ~n8151;
  assign n8158 = ~n38889 & ~n38890;
  assign n8159 = ~n8152 & ~n8153;
  assign n8160 = n7787 & n38891;
  assign n8161 = ~n7787 & ~n38891;
  assign n8162 = ~n8160 & ~n8161;
  assign n8163 = pi14  & ~pi15 ;
  assign n8164 = ~pi14  & pi15 ;
  assign n8165 = ~pi14  & ~pi15 ;
  assign n8166 = pi14  & pi15 ;
  assign n8167 = ~n8165 & ~n8166;
  assign n8168 = ~n8163 & ~n8164;
  assign n8169 = pi16  & ~pi17 ;
  assign n8170 = ~pi16  & pi17 ;
  assign n8171 = ~pi16  & ~pi17 ;
  assign n8172 = pi16  & pi17 ;
  assign n8173 = ~n8171 & ~n8172;
  assign n8174 = ~n8169 & ~n8170;
  assign n8175 = n38892 & n38893;
  assign n8176 = n485 & ~n487;
  assign n8177 = ~n488 & ~n8176;
  assign n8178 = n8175 & n8177;
  assign n8179 = pi15  & ~pi16 ;
  assign n8180 = ~pi15  & pi16 ;
  assign n8181 = ~pi15  & ~pi16 ;
  assign n8182 = pi15  & pi16 ;
  assign n8183 = ~n8181 & ~n8182;
  assign n8184 = ~n8179 & ~n8180;
  assign n8185 = ~n38892 & n38893;
  assign n8186 = ~n38892 & ~n38894;
  assign n8187 = n38893 & n8186;
  assign n8188 = ~n38894 & n8185;
  assign n8189 = pi105  & n38895;
  assign n8190 = n38892 & ~n38893;
  assign n8191 = pi107  & n8190;
  assign n8192 = ~n38892 & n38894;
  assign n8193 = pi106  & n8192;
  assign n8194 = ~n8191 & ~n8193;
  assign n8195 = ~n8189 & ~n8193;
  assign n8196 = ~n8191 & n8195;
  assign n8197 = ~n8189 & n8194;
  assign n8198 = ~n8178 & n38896;
  assign n8199 = pi17  & ~n8198;
  assign n8200 = pi17  & ~n8199;
  assign n8201 = pi17  & n8198;
  assign n8202 = ~n8198 & ~n8199;
  assign n8203 = ~pi17  & ~n8198;
  assign n8204 = ~n38897 & ~n38898;
  assign n8205 = n8162 & ~n8204;
  assign n8206 = n7778 & n38819;
  assign n8207 = ~n7786 & ~n8206;
  assign n8208 = n481 & ~n483;
  assign n8209 = ~n484 & ~n8208;
  assign n8210 = n8175 & n8209;
  assign n8211 = pi104  & n38895;
  assign n8212 = pi106  & n8190;
  assign n8213 = pi105  & n8192;
  assign n8214 = ~n8212 & ~n8213;
  assign n8215 = ~n8211 & ~n8213;
  assign n8216 = ~n8212 & n8215;
  assign n8217 = ~n8211 & n8214;
  assign n8218 = ~n8210 & n38899;
  assign n8219 = pi17  & ~n8218;
  assign n8220 = pi17  & ~n8219;
  assign n8221 = pi17  & n8218;
  assign n8222 = ~n8218 & ~n8219;
  assign n8223 = ~pi17  & ~n8218;
  assign n8224 = ~n38900 & ~n38901;
  assign n8225 = n8207 & ~n8224;
  assign n8226 = n7769 & n38816;
  assign n8227 = ~n7777 & ~n8226;
  assign n8228 = n477 & ~n479;
  assign n8229 = ~n480 & ~n8228;
  assign n8230 = n8175 & n8229;
  assign n8231 = pi103  & n38895;
  assign n8232 = pi105  & n8190;
  assign n8233 = pi104  & n8192;
  assign n8234 = ~n8232 & ~n8233;
  assign n8235 = ~n8231 & ~n8233;
  assign n8236 = ~n8232 & n8235;
  assign n8237 = ~n8231 & n8234;
  assign n8238 = ~n8230 & n38902;
  assign n8239 = pi17  & ~n8238;
  assign n8240 = pi17  & ~n8239;
  assign n8241 = pi17  & n8238;
  assign n8242 = ~n8238 & ~n8239;
  assign n8243 = ~pi17  & ~n8238;
  assign n8244 = ~n38903 & ~n38904;
  assign n8245 = n8227 & ~n8244;
  assign n8246 = n7760 & n38813;
  assign n8247 = ~n7768 & ~n8246;
  assign n8248 = n8136 & n8175;
  assign n8249 = pi102  & n38895;
  assign n8250 = pi104  & n8190;
  assign n8251 = pi103  & n8192;
  assign n8252 = ~n8250 & ~n8251;
  assign n8253 = ~n8249 & ~n8251;
  assign n8254 = ~n8250 & n8253;
  assign n8255 = ~n8249 & n8252;
  assign n8256 = ~n8248 & n38905;
  assign n8257 = pi17  & ~n8256;
  assign n8258 = pi17  & ~n8257;
  assign n8259 = pi17  & n8256;
  assign n8260 = ~n8256 & ~n8257;
  assign n8261 = ~pi17  & ~n8256;
  assign n8262 = ~n38906 & ~n38907;
  assign n8263 = n8247 & ~n8262;
  assign n8264 = n7756 & ~n7758;
  assign n8265 = ~n7759 & ~n8264;
  assign n8266 = n6787 & n8175;
  assign n8267 = pi101  & n38895;
  assign n8268 = pi103  & n8190;
  assign n8269 = pi102  & n8192;
  assign n8270 = ~n8268 & ~n8269;
  assign n8271 = ~n8267 & ~n8269;
  assign n8272 = ~n8268 & n8271;
  assign n8273 = ~n8267 & n8270;
  assign n8274 = ~n8266 & n38908;
  assign n8275 = pi17  & ~n8274;
  assign n8276 = pi17  & ~n8275;
  assign n8277 = pi17  & n8274;
  assign n8278 = ~n8274 & ~n8275;
  assign n8279 = ~pi17  & ~n8274;
  assign n8280 = ~n38909 & ~n38910;
  assign n8281 = n8265 & ~n8280;
  assign n8282 = n7747 & n38810;
  assign n8283 = ~n7755 & ~n8282;
  assign n8284 = n6819 & n8175;
  assign n8285 = pi100  & n38895;
  assign n8286 = pi102  & n8190;
  assign n8287 = pi101  & n8192;
  assign n8288 = ~n8286 & ~n8287;
  assign n8289 = ~n8285 & ~n8287;
  assign n8290 = ~n8286 & n8289;
  assign n8291 = ~n8285 & n8288;
  assign n8292 = ~n8284 & n38911;
  assign n8293 = pi17  & ~n8292;
  assign n8294 = pi17  & ~n8293;
  assign n8295 = pi17  & n8292;
  assign n8296 = ~n8292 & ~n8293;
  assign n8297 = ~pi17  & ~n8292;
  assign n8298 = ~n38912 & ~n38913;
  assign n8299 = n8283 & ~n8298;
  assign n8300 = n7738 & n38807;
  assign n8301 = ~n7746 & ~n8300;
  assign n8302 = n6839 & n8175;
  assign n8303 = pi99  & n38895;
  assign n8304 = pi101  & n8190;
  assign n8305 = pi100  & n8192;
  assign n8306 = ~n8304 & ~n8305;
  assign n8307 = ~n8303 & ~n8305;
  assign n8308 = ~n8304 & n8307;
  assign n8309 = ~n8303 & n8306;
  assign n8310 = ~n8302 & n38914;
  assign n8311 = pi17  & ~n8310;
  assign n8312 = pi17  & ~n8311;
  assign n8313 = pi17  & n8310;
  assign n8314 = ~n8310 & ~n8311;
  assign n8315 = ~pi17  & ~n8310;
  assign n8316 = ~n38915 & ~n38916;
  assign n8317 = n8301 & ~n8316;
  assign n8318 = n6474 & n8175;
  assign n8319 = pi98  & n38895;
  assign n8320 = pi100  & n8190;
  assign n8321 = pi99  & n8192;
  assign n8322 = ~n8320 & ~n8321;
  assign n8323 = ~n8319 & ~n8321;
  assign n8324 = ~n8320 & n8323;
  assign n8325 = ~n8319 & n8322;
  assign n8326 = ~n8318 & n38917;
  assign n8327 = pi17  & ~n8326;
  assign n8328 = pi17  & ~n8327;
  assign n8329 = pi17  & n8326;
  assign n8330 = ~n8326 & ~n8327;
  assign n8331 = ~pi17  & ~n8326;
  assign n8332 = ~n38918 & ~n38919;
  assign n8333 = n7729 & n38804;
  assign n8334 = ~n7729 & n38804;
  assign n8335 = n7729 & ~n38804;
  assign n8336 = ~n8334 & ~n8335;
  assign n8337 = ~n7737 & ~n8333;
  assign n8338 = ~n8332 & ~n38920;
  assign n8339 = n7725 & ~n7727;
  assign n8340 = ~n7728 & ~n8339;
  assign n8341 = n5578 & n8175;
  assign n8342 = pi97  & n38895;
  assign n8343 = pi99  & n8190;
  assign n8344 = pi98  & n8192;
  assign n8345 = ~n8343 & ~n8344;
  assign n8346 = ~n8342 & ~n8344;
  assign n8347 = ~n8343 & n8346;
  assign n8348 = ~n8342 & n8345;
  assign n8349 = ~n8341 & n38921;
  assign n8350 = pi17  & ~n8349;
  assign n8351 = pi17  & ~n8350;
  assign n8352 = pi17  & n8349;
  assign n8353 = ~n8349 & ~n8350;
  assign n8354 = ~pi17  & ~n8349;
  assign n8355 = ~n38922 & ~n38923;
  assign n8356 = n8340 & ~n8355;
  assign n8357 = n7718 & n38801;
  assign n8358 = ~n7724 & ~n8357;
  assign n8359 = n5610 & n8175;
  assign n8360 = pi96  & n38895;
  assign n8361 = pi98  & n8190;
  assign n8362 = pi97  & n8192;
  assign n8363 = ~n8361 & ~n8362;
  assign n8364 = ~n8360 & ~n8362;
  assign n8365 = ~n8361 & n8364;
  assign n8366 = ~n8360 & n8363;
  assign n8367 = ~n8359 & n38924;
  assign n8368 = pi17  & ~n8367;
  assign n8369 = pi17  & ~n8368;
  assign n8370 = pi17  & n8367;
  assign n8371 = ~n8367 & ~n8368;
  assign n8372 = ~pi17  & ~n8367;
  assign n8373 = ~n38925 & ~n38926;
  assign n8374 = n8358 & ~n8373;
  assign n8375 = n7714 & ~n7716;
  assign n8376 = ~n7717 & ~n8375;
  assign n8377 = n5630 & n8175;
  assign n8378 = pi95  & n38895;
  assign n8379 = pi97  & n8190;
  assign n8380 = pi96  & n8192;
  assign n8381 = ~n8379 & ~n8380;
  assign n8382 = ~n8378 & ~n8380;
  assign n8383 = ~n8379 & n8382;
  assign n8384 = ~n8378 & n8381;
  assign n8385 = ~n8377 & n38927;
  assign n8386 = pi17  & ~n8385;
  assign n8387 = pi17  & ~n8386;
  assign n8388 = pi17  & n8385;
  assign n8389 = ~n8385 & ~n8386;
  assign n8390 = ~pi17  & ~n8385;
  assign n8391 = ~n38928 & ~n38929;
  assign n8392 = n8376 & ~n8391;
  assign n8393 = n5281 & n8175;
  assign n8394 = pi94  & n38895;
  assign n8395 = pi96  & n8190;
  assign n8396 = pi95  & n8192;
  assign n8397 = ~n8395 & ~n8396;
  assign n8398 = ~n8394 & ~n8396;
  assign n8399 = ~n8395 & n8398;
  assign n8400 = ~n8394 & n8397;
  assign n8401 = ~n8393 & n38930;
  assign n8402 = pi17  & ~n8401;
  assign n8403 = pi17  & ~n8402;
  assign n8404 = pi17  & n8401;
  assign n8405 = ~n8401 & ~n8402;
  assign n8406 = ~pi17  & ~n8401;
  assign n8407 = ~n38931 & ~n38932;
  assign n8408 = n7710 & ~n7712;
  assign n8409 = ~n7713 & ~n8408;
  assign n8410 = ~n8407 & n8409;
  assign n8411 = n4494 & n8175;
  assign n8412 = pi93  & n38895;
  assign n8413 = pi95  & n8190;
  assign n8414 = pi94  & n8192;
  assign n8415 = ~n8413 & ~n8414;
  assign n8416 = ~n8412 & ~n8414;
  assign n8417 = ~n8413 & n8416;
  assign n8418 = ~n8412 & n8415;
  assign n8419 = ~n8411 & n38933;
  assign n8420 = pi17  & ~n8419;
  assign n8421 = pi17  & ~n8420;
  assign n8422 = pi17  & n8419;
  assign n8423 = ~n8419 & ~n8420;
  assign n8424 = ~pi17  & ~n8419;
  assign n8425 = ~n38934 & ~n38935;
  assign n8426 = n7701 & n38800;
  assign n8427 = ~n7701 & ~n7709;
  assign n8428 = ~n7701 & n38800;
  assign n8429 = ~n38800 & ~n7709;
  assign n8430 = n7701 & ~n38800;
  assign n8431 = ~n38936 & ~n38937;
  assign n8432 = ~n7709 & ~n8426;
  assign n8433 = ~n8425 & ~n38938;
  assign n8434 = n4524 & n8175;
  assign n8435 = pi92  & n38895;
  assign n8436 = pi94  & n8190;
  assign n8437 = pi93  & n8192;
  assign n8438 = ~n8436 & ~n8437;
  assign n8439 = ~n8435 & ~n8437;
  assign n8440 = ~n8436 & n8439;
  assign n8441 = ~n8435 & n8438;
  assign n8442 = ~n8434 & n38939;
  assign n8443 = pi17  & ~n8442;
  assign n8444 = pi17  & ~n8443;
  assign n8445 = pi17  & n8442;
  assign n8446 = ~n8442 & ~n8443;
  assign n8447 = ~pi17  & ~n8442;
  assign n8448 = ~n38940 & ~n38941;
  assign n8449 = n7692 & n38797;
  assign n8450 = ~n7692 & n38797;
  assign n8451 = n7692 & ~n38797;
  assign n8452 = ~n8450 & ~n8451;
  assign n8453 = ~n7700 & ~n8449;
  assign n8454 = ~n8448 & ~n38942;
  assign n8455 = n4544 & n8175;
  assign n8456 = pi91  & n38895;
  assign n8457 = pi93  & n8190;
  assign n8458 = pi92  & n8192;
  assign n8459 = ~n8457 & ~n8458;
  assign n8460 = ~n8456 & ~n8458;
  assign n8461 = ~n8457 & n8460;
  assign n8462 = ~n8456 & n8459;
  assign n8463 = ~n8455 & n38943;
  assign n8464 = pi17  & ~n8463;
  assign n8465 = pi17  & ~n8464;
  assign n8466 = pi17  & n8463;
  assign n8467 = ~n8463 & ~n8464;
  assign n8468 = ~pi17  & ~n8463;
  assign n8469 = ~n38944 & ~n38945;
  assign n8470 = n7688 & ~n7690;
  assign n8471 = ~n7691 & ~n8470;
  assign n8472 = ~n8469 & n8471;
  assign n8473 = n4453 & n8175;
  assign n8474 = pi90  & n38895;
  assign n8475 = pi92  & n8190;
  assign n8476 = pi91  & n8192;
  assign n8477 = ~n8475 & ~n8476;
  assign n8478 = ~n8474 & ~n8476;
  assign n8479 = ~n8475 & n8478;
  assign n8480 = ~n8474 & n8477;
  assign n8481 = ~n8473 & n38946;
  assign n8482 = pi17  & ~n8481;
  assign n8483 = pi17  & ~n8482;
  assign n8484 = pi17  & n8481;
  assign n8485 = ~n8481 & ~n8482;
  assign n8486 = ~pi17  & ~n8481;
  assign n8487 = ~n38947 & ~n38948;
  assign n8488 = n7679 & n38794;
  assign n8489 = ~n7687 & ~n8488;
  assign n8490 = ~n8487 & n8489;
  assign n8491 = n7675 & ~n7677;
  assign n8492 = ~n7678 & ~n8491;
  assign n8493 = n594 & n8175;
  assign n8494 = pi89  & n38895;
  assign n8495 = pi91  & n8190;
  assign n8496 = pi90  & n8192;
  assign n8497 = ~n8495 & ~n8496;
  assign n8498 = ~n8494 & ~n8496;
  assign n8499 = ~n8495 & n8498;
  assign n8500 = ~n8494 & n8497;
  assign n8501 = ~n8493 & n38949;
  assign n8502 = pi17  & ~n8501;
  assign n8503 = pi17  & ~n8502;
  assign n8504 = pi17  & n8501;
  assign n8505 = ~n8501 & ~n8502;
  assign n8506 = ~pi17  & ~n8501;
  assign n8507 = ~n38950 & ~n38951;
  assign n8508 = n8492 & ~n8507;
  assign n8509 = n3566 & n8175;
  assign n8510 = pi88  & n38895;
  assign n8511 = pi90  & n8190;
  assign n8512 = pi89  & n8192;
  assign n8513 = ~n8511 & ~n8512;
  assign n8514 = ~n8510 & ~n8512;
  assign n8515 = ~n8511 & n8514;
  assign n8516 = ~n8510 & n8513;
  assign n8517 = ~n8509 & n38952;
  assign n8518 = pi17  & ~n8517;
  assign n8519 = pi17  & ~n8518;
  assign n8520 = pi17  & n8517;
  assign n8521 = ~n8517 & ~n8518;
  assign n8522 = ~pi17  & ~n8517;
  assign n8523 = ~n38953 & ~n38954;
  assign n8524 = n7669 & ~n7671;
  assign n8525 = ~n7669 & ~n38791;
  assign n8526 = ~n7670 & n7675;
  assign n8527 = ~n8525 & ~n8526;
  assign n8528 = ~n38791 & ~n8524;
  assign n8529 = ~n8523 & ~n38955;
  assign n8530 = n7660 & n38790;
  assign n8531 = ~n7668 & ~n8530;
  assign n8532 = n3591 & n8175;
  assign n8533 = pi87  & n38895;
  assign n8534 = pi89  & n8190;
  assign n8535 = pi88  & n8192;
  assign n8536 = ~n8534 & ~n8535;
  assign n8537 = ~n8533 & ~n8535;
  assign n8538 = ~n8534 & n8537;
  assign n8539 = ~n8533 & n8536;
  assign n8540 = ~n8532 & n38956;
  assign n8541 = pi17  & ~n8540;
  assign n8542 = pi17  & ~n8541;
  assign n8543 = pi17  & n8540;
  assign n8544 = ~n8540 & ~n8541;
  assign n8545 = ~pi17  & ~n8540;
  assign n8546 = ~n38957 & ~n38958;
  assign n8547 = n8531 & ~n8546;
  assign n8548 = n7651 & n38787;
  assign n8549 = ~n7659 & ~n8548;
  assign n8550 = n3354 & n8175;
  assign n8551 = pi86  & n38895;
  assign n8552 = pi88  & n8190;
  assign n8553 = pi87  & n8192;
  assign n8554 = ~n8552 & ~n8553;
  assign n8555 = ~n8551 & ~n8553;
  assign n8556 = ~n8552 & n8555;
  assign n8557 = ~n8551 & n8554;
  assign n8558 = ~n8550 & n38959;
  assign n8559 = pi17  & ~n8558;
  assign n8560 = pi17  & ~n8559;
  assign n8561 = pi17  & n8558;
  assign n8562 = ~n8558 & ~n8559;
  assign n8563 = ~pi17  & ~n8558;
  assign n8564 = ~n38960 & ~n38961;
  assign n8565 = n8549 & ~n8564;
  assign n8566 = n7642 & n38784;
  assign n8567 = ~n7650 & ~n8566;
  assign n8568 = n636 & n8175;
  assign n8569 = pi85  & n38895;
  assign n8570 = pi87  & n8190;
  assign n8571 = pi86  & n8192;
  assign n8572 = ~n8570 & ~n8571;
  assign n8573 = ~n8569 & ~n8571;
  assign n8574 = ~n8570 & n8573;
  assign n8575 = ~n8569 & n8572;
  assign n8576 = ~n8568 & n38962;
  assign n8577 = pi17  & ~n8576;
  assign n8578 = pi17  & ~n8577;
  assign n8579 = pi17  & n8576;
  assign n8580 = ~n8576 & ~n8577;
  assign n8581 = ~pi17  & ~n8576;
  assign n8582 = ~n38963 & ~n38964;
  assign n8583 = n8567 & ~n8582;
  assign n8584 = n7633 & n38781;
  assign n8585 = ~n7641 & ~n8584;
  assign n8586 = n2779 & n8175;
  assign n8587 = pi84  & n38895;
  assign n8588 = pi86  & n8190;
  assign n8589 = pi85  & n8192;
  assign n8590 = ~n8588 & ~n8589;
  assign n8591 = ~n8587 & ~n8589;
  assign n8592 = ~n8588 & n8591;
  assign n8593 = ~n8587 & n8590;
  assign n8594 = ~n8586 & n38965;
  assign n8595 = pi17  & ~n8594;
  assign n8596 = pi17  & ~n8595;
  assign n8597 = pi17  & n8594;
  assign n8598 = ~n8594 & ~n8595;
  assign n8599 = ~pi17  & ~n8594;
  assign n8600 = ~n38966 & ~n38967;
  assign n8601 = n8585 & ~n8600;
  assign n8602 = n7629 & ~n7631;
  assign n8603 = ~n7632 & ~n8602;
  assign n8604 = n2804 & n8175;
  assign n8605 = pi83  & n38895;
  assign n8606 = pi85  & n8190;
  assign n8607 = pi84  & n8192;
  assign n8608 = ~n8606 & ~n8607;
  assign n8609 = ~n8605 & ~n8607;
  assign n8610 = ~n8606 & n8609;
  assign n8611 = ~n8605 & n8608;
  assign n8612 = ~n8604 & n38968;
  assign n8613 = pi17  & ~n8612;
  assign n8614 = pi17  & ~n8613;
  assign n8615 = pi17  & n8612;
  assign n8616 = ~n8612 & ~n8613;
  assign n8617 = ~pi17  & ~n8612;
  assign n8618 = ~n38969 & ~n38970;
  assign n8619 = n8603 & ~n8618;
  assign n8620 = n7620 & n38778;
  assign n8621 = ~n7628 & ~n8620;
  assign n8622 = n2591 & n8175;
  assign n8623 = pi82  & n38895;
  assign n8624 = pi84  & n8190;
  assign n8625 = pi83  & n8192;
  assign n8626 = ~n8624 & ~n8625;
  assign n8627 = ~n8623 & ~n8625;
  assign n8628 = ~n8624 & n8627;
  assign n8629 = ~n8623 & n8626;
  assign n8630 = ~n8622 & n38971;
  assign n8631 = pi17  & ~n8630;
  assign n8632 = pi17  & ~n8631;
  assign n8633 = pi17  & n8630;
  assign n8634 = ~n8630 & ~n8631;
  assign n8635 = ~pi17  & ~n8630;
  assign n8636 = ~n38972 & ~n38973;
  assign n8637 = n8621 & ~n8636;
  assign n8638 = n7611 & n38775;
  assign n8639 = ~n7619 & ~n8638;
  assign n8640 = n2091 & n8175;
  assign n8641 = pi81  & n38895;
  assign n8642 = pi83  & n8190;
  assign n8643 = pi82  & n8192;
  assign n8644 = ~n8642 & ~n8643;
  assign n8645 = ~n8641 & ~n8643;
  assign n8646 = ~n8642 & n8645;
  assign n8647 = ~n8641 & n8644;
  assign n8648 = ~n8640 & n38974;
  assign n8649 = pi17  & ~n8648;
  assign n8650 = pi17  & ~n8649;
  assign n8651 = pi17  & n8648;
  assign n8652 = ~n8648 & ~n8649;
  assign n8653 = ~pi17  & ~n8648;
  assign n8654 = ~n38975 & ~n38976;
  assign n8655 = n8639 & ~n8654;
  assign n8656 = n2134 & n8175;
  assign n8657 = pi80  & n38895;
  assign n8658 = pi82  & n8190;
  assign n8659 = pi81  & n8192;
  assign n8660 = ~n8658 & ~n8659;
  assign n8661 = ~n8657 & ~n8659;
  assign n8662 = ~n8658 & n8661;
  assign n8663 = ~n8657 & n8660;
  assign n8664 = ~n8656 & n38977;
  assign n8665 = pi17  & ~n8664;
  assign n8666 = pi17  & ~n8665;
  assign n8667 = pi17  & n8664;
  assign n8668 = ~n8664 & ~n8665;
  assign n8669 = ~pi17  & ~n8664;
  assign n8670 = ~n38978 & ~n38979;
  assign n8671 = n7602 & n38772;
  assign n8672 = ~n7602 & n38772;
  assign n8673 = n7602 & ~n38772;
  assign n8674 = ~n8672 & ~n8673;
  assign n8675 = ~n7610 & ~n8671;
  assign n8676 = ~n8670 & ~n38980;
  assign n8677 = n7598 & ~n7600;
  assign n8678 = ~n7601 & ~n8677;
  assign n8679 = n2154 & n8175;
  assign n8680 = pi79  & n38895;
  assign n8681 = pi81  & n8190;
  assign n8682 = pi80  & n8192;
  assign n8683 = ~n8681 & ~n8682;
  assign n8684 = ~n8680 & ~n8682;
  assign n8685 = ~n8681 & n8684;
  assign n8686 = ~n8680 & n8683;
  assign n8687 = ~n8679 & n38981;
  assign n8688 = pi17  & ~n8687;
  assign n8689 = pi17  & ~n8688;
  assign n8690 = pi17  & n8687;
  assign n8691 = ~n8687 & ~n8688;
  assign n8692 = ~pi17  & ~n8687;
  assign n8693 = ~n38982 & ~n38983;
  assign n8694 = n8678 & ~n8693;
  assign n8695 = ~n7312 & n7596;
  assign n8696 = ~n7597 & ~n8695;
  assign n8697 = n2063 & n8175;
  assign n8698 = pi78  & n38895;
  assign n8699 = pi80  & n8190;
  assign n8700 = pi79  & n8192;
  assign n8701 = ~n8699 & ~n8700;
  assign n8702 = ~n8698 & ~n8700;
  assign n8703 = ~n8699 & n8702;
  assign n8704 = ~n8698 & n8701;
  assign n8705 = ~n8697 & n38984;
  assign n8706 = pi17  & ~n8705;
  assign n8707 = pi17  & ~n8706;
  assign n8708 = pi17  & n8705;
  assign n8709 = ~n8705 & ~n8706;
  assign n8710 = ~pi17  & ~n8705;
  assign n8711 = ~n38985 & ~n38986;
  assign n8712 = n8696 & ~n8711;
  assign n8713 = n7592 & ~n7594;
  assign n8714 = ~n7595 & ~n8713;
  assign n8715 = n678 & n8175;
  assign n8716 = pi77  & n38895;
  assign n8717 = pi79  & n8190;
  assign n8718 = pi78  & n8192;
  assign n8719 = ~n8717 & ~n8718;
  assign n8720 = ~n8716 & ~n8718;
  assign n8721 = ~n8717 & n8720;
  assign n8722 = ~n8716 & n8719;
  assign n8723 = ~n8715 & n38987;
  assign n8724 = pi17  & ~n8723;
  assign n8725 = pi17  & ~n8724;
  assign n8726 = pi17  & n8723;
  assign n8727 = ~n8723 & ~n8724;
  assign n8728 = ~pi17  & ~n8723;
  assign n8729 = ~n38988 & ~n38989;
  assign n8730 = n8714 & ~n8729;
  assign n8731 = n7588 & ~n7590;
  assign n8732 = ~n7591 & ~n8731;
  assign n8733 = n1578 & n8175;
  assign n8734 = pi76  & n38895;
  assign n8735 = pi78  & n8190;
  assign n8736 = pi77  & n8192;
  assign n8737 = ~n8735 & ~n8736;
  assign n8738 = ~n8734 & ~n8736;
  assign n8739 = ~n8735 & n8738;
  assign n8740 = ~n8734 & n8737;
  assign n8741 = ~n8733 & n38990;
  assign n8742 = pi17  & ~n8741;
  assign n8743 = pi17  & ~n8742;
  assign n8744 = pi17  & n8741;
  assign n8745 = ~n8741 & ~n8742;
  assign n8746 = ~pi17  & ~n8741;
  assign n8747 = ~n38991 & ~n38992;
  assign n8748 = n8732 & ~n8747;
  assign n8749 = n7579 & n38769;
  assign n8750 = ~n7587 & ~n8749;
  assign n8751 = n1596 & n8175;
  assign n8752 = pi75  & n38895;
  assign n8753 = pi77  & n8190;
  assign n8754 = pi76  & n8192;
  assign n8755 = ~n8753 & ~n8754;
  assign n8756 = ~n8752 & ~n8754;
  assign n8757 = ~n8753 & n8756;
  assign n8758 = ~n8752 & n8755;
  assign n8759 = ~n8751 & n38993;
  assign n8760 = pi17  & ~n8759;
  assign n8761 = pi17  & ~n8760;
  assign n8762 = pi17  & n8759;
  assign n8763 = ~n8759 & ~n8760;
  assign n8764 = ~pi17  & ~n8759;
  assign n8765 = ~n38994 & ~n38995;
  assign n8766 = n8750 & ~n8765;
  assign n8767 = n1465 & n8175;
  assign n8768 = pi74  & n38895;
  assign n8769 = pi76  & n8190;
  assign n8770 = pi75  & n8192;
  assign n8771 = ~n8769 & ~n8770;
  assign n8772 = ~n8768 & ~n8770;
  assign n8773 = ~n8769 & n8772;
  assign n8774 = ~n8768 & n8771;
  assign n8775 = ~n8767 & n38996;
  assign n8776 = pi17  & ~n8775;
  assign n8777 = pi17  & ~n8776;
  assign n8778 = pi17  & n8775;
  assign n8779 = ~n8775 & ~n8776;
  assign n8780 = ~pi17  & ~n8775;
  assign n8781 = ~n38997 & ~n38998;
  assign n8782 = n7575 & ~n7577;
  assign n8783 = ~n7578 & ~n8782;
  assign n8784 = ~n8781 & n8783;
  assign n8785 = n720 & n8175;
  assign n8786 = pi73  & n38895;
  assign n8787 = pi75  & n8190;
  assign n8788 = pi74  & n8192;
  assign n8789 = ~n8787 & ~n8788;
  assign n8790 = ~n8786 & ~n8788;
  assign n8791 = ~n8787 & n8790;
  assign n8792 = ~n8786 & n8789;
  assign n8793 = ~n8785 & n38999;
  assign n8794 = pi17  & ~n8793;
  assign n8795 = pi17  & ~n8794;
  assign n8796 = pi17  & n8793;
  assign n8797 = ~n8793 & ~n8794;
  assign n8798 = ~pi17  & ~n8793;
  assign n8799 = ~n39000 & ~n39001;
  assign n8800 = n7571 & ~n7573;
  assign n8801 = ~n7574 & ~n8800;
  assign n8802 = ~n8799 & n8801;
  assign n8803 = n7567 & ~n7569;
  assign n8804 = ~n7570 & ~n8803;
  assign n8805 = n1218 & n8175;
  assign n8806 = pi72  & n38895;
  assign n8807 = pi74  & n8190;
  assign n8808 = pi73  & n8192;
  assign n8809 = ~n8807 & ~n8808;
  assign n8810 = ~n8806 & ~n8808;
  assign n8811 = ~n8807 & n8810;
  assign n8812 = ~n8806 & n8809;
  assign n8813 = ~n8805 & n39002;
  assign n8814 = pi17  & ~n8813;
  assign n8815 = pi17  & ~n8814;
  assign n8816 = pi17  & n8813;
  assign n8817 = ~n8813 & ~n8814;
  assign n8818 = ~pi17  & ~n8813;
  assign n8819 = ~n39003 & ~n39004;
  assign n8820 = n8804 & ~n8819;
  assign n8821 = n1238 & n8175;
  assign n8822 = pi71  & n38895;
  assign n8823 = pi73  & n8190;
  assign n8824 = pi72  & n8192;
  assign n8825 = ~n8823 & ~n8824;
  assign n8826 = ~n8822 & ~n8824;
  assign n8827 = ~n8823 & n8826;
  assign n8828 = ~n8822 & n8825;
  assign n8829 = ~n8821 & n39005;
  assign n8830 = pi17  & ~n8829;
  assign n8831 = pi17  & ~n8830;
  assign n8832 = pi17  & n8829;
  assign n8833 = ~n8829 & ~n8830;
  assign n8834 = ~pi17  & ~n8829;
  assign n8835 = ~n39006 & ~n39007;
  assign n8836 = n7558 & n38766;
  assign n8837 = ~n7558 & n38766;
  assign n8838 = n7558 & ~n38766;
  assign n8839 = ~n8837 & ~n8838;
  assign n8840 = ~n7566 & ~n8836;
  assign n8841 = ~n8835 & ~n39008;
  assign n8842 = n1124 & n8175;
  assign n8843 = pi70  & n38895;
  assign n8844 = pi72  & n8190;
  assign n8845 = pi71  & n8192;
  assign n8846 = ~n8844 & ~n8845;
  assign n8847 = ~n8843 & ~n8845;
  assign n8848 = ~n8844 & n8847;
  assign n8849 = ~n8843 & n8846;
  assign n8850 = ~n8842 & n39009;
  assign n8851 = pi17  & ~n8850;
  assign n8852 = pi17  & ~n8851;
  assign n8853 = pi17  & n8850;
  assign n8854 = ~n8850 & ~n8851;
  assign n8855 = ~pi17  & ~n8850;
  assign n8856 = ~n39010 & ~n39011;
  assign n8857 = n7552 & ~n7554;
  assign n8858 = ~n7552 & ~n38763;
  assign n8859 = ~n7553 & n7558;
  assign n8860 = ~n8858 & ~n8859;
  assign n8861 = ~n38763 & ~n8857;
  assign n8862 = ~n8856 & ~n39012;
  assign n8863 = n927 & n8175;
  assign n8864 = pi69  & n38895;
  assign n8865 = pi71  & n8190;
  assign n8866 = pi70  & n8192;
  assign n8867 = ~n8865 & ~n8866;
  assign n8868 = ~n8864 & ~n8866;
  assign n8869 = ~n8865 & n8868;
  assign n8870 = ~n8864 & n8867;
  assign n8871 = ~n8863 & n39013;
  assign n8872 = pi17  & ~n8871;
  assign n8873 = pi17  & ~n8872;
  assign n8874 = pi17  & n8871;
  assign n8875 = ~n8871 & ~n8872;
  assign n8876 = ~pi17  & ~n8871;
  assign n8877 = ~n39014 & ~n39015;
  assign n8878 = n7545 & n38762;
  assign n8879 = ~n7551 & ~n8878;
  assign n8880 = ~n8877 & n8879;
  assign n8881 = n7538 & n38761;
  assign n8882 = ~n7544 & ~n8881;
  assign n8883 = n972 & n8175;
  assign n8884 = pi68  & n38895;
  assign n8885 = pi70  & n8190;
  assign n8886 = pi69  & n8192;
  assign n8887 = ~n8885 & ~n8886;
  assign n8888 = ~n8884 & ~n8886;
  assign n8889 = ~n8885 & n8888;
  assign n8890 = ~n8884 & n8887;
  assign n8891 = ~n8883 & n39016;
  assign n8892 = pi17  & ~n8891;
  assign n8893 = pi17  & ~n8892;
  assign n8894 = pi17  & n8891;
  assign n8895 = ~n8891 & ~n8892;
  assign n8896 = ~pi17  & ~n8891;
  assign n8897 = ~n39017 & ~n39018;
  assign n8898 = n8882 & ~n8897;
  assign n8899 = n990 & n8175;
  assign n8900 = pi67  & n38895;
  assign n8901 = pi69  & n8190;
  assign n8902 = pi68  & n8192;
  assign n8903 = ~n8901 & ~n8902;
  assign n8904 = ~n8900 & ~n8902;
  assign n8905 = ~n8901 & n8904;
  assign n8906 = ~n8900 & n8903;
  assign n8907 = ~n8899 & n39019;
  assign n8908 = pi17  & ~n8907;
  assign n8909 = pi17  & ~n8908;
  assign n8910 = pi17  & n8907;
  assign n8911 = ~n8907 & ~n8908;
  assign n8912 = ~pi17  & ~n8907;
  assign n8913 = ~n39020 & ~n39021;
  assign n8914 = pi20  & ~n38753;
  assign n8915 = n38756 & ~n8914;
  assign n8916 = ~n38756 & n8914;
  assign n8917 = ~n38753 & n7520;
  assign n8918 = ~n38757 & ~n8917;
  assign n8919 = ~n8915 & ~n8916;
  assign n8920 = ~n8913 & n39022;
  assign n8921 = n871 & n8175;
  assign n8922 = pi66  & n38895;
  assign n8923 = pi68  & n8190;
  assign n8924 = pi67  & n8192;
  assign n8925 = ~n8923 & ~n8924;
  assign n8926 = ~n8922 & ~n8924;
  assign n8927 = ~n8923 & n8926;
  assign n8928 = ~n8922 & n8925;
  assign n8929 = ~n8921 & n39023;
  assign n8930 = pi17  & ~n8929;
  assign n8931 = pi17  & ~n8930;
  assign n8932 = pi17  & n8929;
  assign n8933 = ~n8929 & ~n8930;
  assign n8934 = ~pi17  & ~n8929;
  assign n8935 = ~n39024 & ~n39025;
  assign n8936 = pi20  & n7494;
  assign n8937 = ~n7493 & n8936;
  assign n8938 = n7493 & ~n8936;
  assign n8939 = ~n7495 & n7499;
  assign n8940 = ~n38753 & ~n8939;
  assign n8941 = ~n8937 & ~n8938;
  assign n8942 = ~n8935 & n39026;
  assign n8943 = n37515 & n8175;
  assign n8944 = pi65  & n8190;
  assign n8945 = pi64  & n8192;
  assign n8946 = ~n8944 & ~n8945;
  assign n8947 = ~n8943 & n8946;
  assign n8948 = pi64  & n38892;
  assign n8949 = pi17  & ~n8948;
  assign n8950 = pi17  & ~n8947;
  assign n8951 = pi17  & ~n8950;
  assign n8952 = ~n8947 & ~n8950;
  assign n8953 = ~n8951 & ~n8952;
  assign n8954 = n8949 & ~n8953;
  assign n8955 = n8947 & n8949;
  assign n8956 = pi64  & n38895;
  assign n8957 = pi65  & n8192;
  assign n8958 = ~n37521 & n8175;
  assign n8959 = pi66  & n8190;
  assign n8960 = ~n8958 & ~n8959;
  assign n8961 = ~n8957 & ~n8958;
  assign n8962 = ~n8959 & n8961;
  assign n8963 = ~n8957 & ~n8959;
  assign n8964 = ~n8958 & n8963;
  assign n8965 = ~n8957 & n8960;
  assign n8966 = ~n8956 & ~n8957;
  assign n8967 = ~n8959 & n8966;
  assign n8968 = ~n8956 & n8963;
  assign n8969 = ~n8958 & n39029;
  assign n8970 = ~n8956 & n39028;
  assign n8971 = pi17  & ~n39030;
  assign n8972 = pi17  & ~n8971;
  assign n8973 = ~n39030 & ~n8971;
  assign n8974 = ~n8972 & ~n8973;
  assign n8975 = n39027 & ~n8974;
  assign n8976 = n39027 & n39030;
  assign n8977 = n7494 & n39031;
  assign n8978 = n847 & n8175;
  assign n8979 = pi65  & n38895;
  assign n8980 = pi67  & n8190;
  assign n8981 = pi66  & n8192;
  assign n8982 = ~n8980 & ~n8981;
  assign n8983 = ~n8979 & ~n8981;
  assign n8984 = ~n8980 & n8983;
  assign n8985 = ~n8979 & n8982;
  assign n8986 = ~n8978 & n39032;
  assign n8987 = pi17  & ~n8986;
  assign n8988 = pi17  & ~n8987;
  assign n8989 = pi17  & n8986;
  assign n8990 = ~n8986 & ~n8987;
  assign n8991 = ~pi17  & ~n8986;
  assign n8992 = ~n39033 & ~n39034;
  assign n8993 = ~n7494 & ~n39031;
  assign n8994 = n7494 & ~n39031;
  assign n8995 = ~n7494 & n39031;
  assign n8996 = ~n8994 & ~n8995;
  assign n8997 = ~n8977 & ~n8993;
  assign n8998 = ~n8992 & ~n39035;
  assign n8999 = ~n8977 & ~n8998;
  assign n9000 = n8935 & ~n39026;
  assign n9001 = n8935 & n39026;
  assign n9002 = ~n8935 & ~n39026;
  assign n9003 = ~n9001 & ~n9002;
  assign n9004 = ~n8942 & ~n9000;
  assign n9005 = ~n8999 & ~n39036;
  assign n9006 = ~n8942 & ~n9005;
  assign n9007 = n8913 & ~n39022;
  assign n9008 = ~n8920 & ~n9007;
  assign n9009 = ~n9006 & ~n9007;
  assign n9010 = ~n8920 & n9009;
  assign n9011 = ~n9006 & n9008;
  assign n9012 = ~n8920 & ~n39037;
  assign n9013 = ~n8882 & n8897;
  assign n9014 = n8882 & ~n8898;
  assign n9015 = n8882 & n8897;
  assign n9016 = ~n8897 & ~n8898;
  assign n9017 = ~n8882 & ~n8897;
  assign n9018 = ~n39038 & ~n39039;
  assign n9019 = ~n8898 & ~n9013;
  assign n9020 = ~n9012 & ~n39040;
  assign n9021 = ~n8898 & ~n9020;
  assign n9022 = n8877 & ~n8879;
  assign n9023 = ~n8880 & ~n9022;
  assign n9024 = ~n9021 & n9023;
  assign n9025 = ~n8880 & ~n9024;
  assign n9026 = n8856 & n39012;
  assign n9027 = ~n8862 & ~n9026;
  assign n9028 = ~n9025 & n9027;
  assign n9029 = ~n8862 & ~n9028;
  assign n9030 = n8835 & n39008;
  assign n9031 = ~n8841 & ~n9030;
  assign n9032 = ~n9029 & n9031;
  assign n9033 = ~n8841 & ~n9032;
  assign n9034 = ~n8804 & n8819;
  assign n9035 = n8804 & ~n8820;
  assign n9036 = n8804 & n8819;
  assign n9037 = ~n8819 & ~n8820;
  assign n9038 = ~n8804 & ~n8819;
  assign n9039 = ~n39041 & ~n39042;
  assign n9040 = ~n8820 & ~n9034;
  assign n9041 = ~n9033 & ~n39043;
  assign n9042 = ~n8820 & ~n9041;
  assign n9043 = n8799 & ~n8801;
  assign n9044 = ~n8802 & ~n9043;
  assign n9045 = ~n9042 & n9044;
  assign n9046 = ~n8802 & ~n9045;
  assign n9047 = n8781 & ~n8783;
  assign n9048 = ~n8784 & ~n9047;
  assign n9049 = ~n9046 & n9048;
  assign n9050 = ~n8784 & ~n9049;
  assign n9051 = ~n8750 & n8765;
  assign n9052 = n8750 & ~n8766;
  assign n9053 = n8750 & n8765;
  assign n9054 = ~n8765 & ~n8766;
  assign n9055 = ~n8750 & ~n8765;
  assign n9056 = ~n39044 & ~n39045;
  assign n9057 = ~n8766 & ~n9051;
  assign n9058 = ~n9050 & ~n39046;
  assign n9059 = ~n8766 & ~n9058;
  assign n9060 = ~n8732 & n8747;
  assign n9061 = n8732 & ~n8748;
  assign n9062 = n8732 & n8747;
  assign n9063 = ~n8747 & ~n8748;
  assign n9064 = ~n8732 & ~n8747;
  assign n9065 = ~n39047 & ~n39048;
  assign n9066 = ~n8748 & ~n9060;
  assign n9067 = ~n9059 & ~n39049;
  assign n9068 = ~n8748 & ~n9067;
  assign n9069 = ~n8714 & n8729;
  assign n9070 = n8714 & ~n8730;
  assign n9071 = n8714 & n8729;
  assign n9072 = ~n8729 & ~n8730;
  assign n9073 = ~n8714 & ~n8729;
  assign n9074 = ~n39050 & ~n39051;
  assign n9075 = ~n8730 & ~n9069;
  assign n9076 = ~n9068 & ~n39052;
  assign n9077 = ~n8730 & ~n9076;
  assign n9078 = ~n8696 & n8711;
  assign n9079 = n8696 & ~n8712;
  assign n9080 = n8696 & n8711;
  assign n9081 = ~n8711 & ~n8712;
  assign n9082 = ~n8696 & ~n8711;
  assign n9083 = ~n39053 & ~n39054;
  assign n9084 = ~n8712 & ~n9078;
  assign n9085 = ~n9077 & ~n39055;
  assign n9086 = ~n8712 & ~n9085;
  assign n9087 = ~n8678 & n8693;
  assign n9088 = n8678 & ~n8694;
  assign n9089 = n8678 & n8693;
  assign n9090 = ~n8693 & ~n8694;
  assign n9091 = ~n8678 & ~n8693;
  assign n9092 = ~n39056 & ~n39057;
  assign n9093 = ~n8694 & ~n9087;
  assign n9094 = ~n9086 & ~n39058;
  assign n9095 = ~n8694 & ~n9094;
  assign n9096 = n8670 & n38980;
  assign n9097 = ~n8676 & ~n9096;
  assign n9098 = ~n9095 & n9097;
  assign n9099 = ~n8676 & ~n9098;
  assign n9100 = ~n8639 & n8654;
  assign n9101 = n8639 & ~n8655;
  assign n9102 = n8639 & n8654;
  assign n9103 = ~n8654 & ~n8655;
  assign n9104 = ~n8639 & ~n8654;
  assign n9105 = ~n39059 & ~n39060;
  assign n9106 = ~n8655 & ~n9100;
  assign n9107 = ~n9099 & ~n39061;
  assign n9108 = ~n8655 & ~n9107;
  assign n9109 = ~n8621 & n8636;
  assign n9110 = ~n8637 & ~n9109;
  assign n9111 = ~n9108 & ~n9109;
  assign n9112 = ~n8637 & n9111;
  assign n9113 = ~n9108 & n9110;
  assign n9114 = ~n8637 & ~n39062;
  assign n9115 = ~n8603 & n8618;
  assign n9116 = n8603 & ~n8619;
  assign n9117 = n8603 & n8618;
  assign n9118 = ~n8618 & ~n8619;
  assign n9119 = ~n8603 & ~n8618;
  assign n9120 = ~n39063 & ~n39064;
  assign n9121 = ~n8619 & ~n9115;
  assign n9122 = ~n9114 & ~n39065;
  assign n9123 = ~n8619 & ~n9122;
  assign n9124 = ~n8585 & n8600;
  assign n9125 = n8585 & ~n8601;
  assign n9126 = n8585 & n8600;
  assign n9127 = ~n8600 & ~n8601;
  assign n9128 = ~n8585 & ~n8600;
  assign n9129 = ~n39066 & ~n39067;
  assign n9130 = ~n8601 & ~n9124;
  assign n9131 = ~n9123 & ~n39068;
  assign n9132 = ~n8601 & ~n9131;
  assign n9133 = ~n8567 & n8582;
  assign n9134 = ~n8583 & ~n9133;
  assign n9135 = ~n9132 & ~n9133;
  assign n9136 = ~n8583 & n9135;
  assign n9137 = ~n9132 & n9134;
  assign n9138 = ~n8583 & ~n39069;
  assign n9139 = ~n8549 & n8564;
  assign n9140 = ~n8565 & ~n9139;
  assign n9141 = ~n9138 & n9140;
  assign n9142 = ~n8565 & ~n9141;
  assign n9143 = ~n8531 & n8546;
  assign n9144 = n8531 & ~n8547;
  assign n9145 = n8531 & n8546;
  assign n9146 = ~n8546 & ~n8547;
  assign n9147 = ~n8531 & ~n8546;
  assign n9148 = ~n39070 & ~n39071;
  assign n9149 = ~n8547 & ~n9143;
  assign n9150 = ~n9142 & ~n39072;
  assign n9151 = ~n8547 & ~n9150;
  assign n9152 = n8523 & n38955;
  assign n9153 = ~n8529 & ~n9152;
  assign n9154 = ~n9151 & n9153;
  assign n9155 = ~n8529 & ~n9154;
  assign n9156 = ~n8492 & n8507;
  assign n9157 = n8492 & ~n8508;
  assign n9158 = n8492 & n8507;
  assign n9159 = ~n8507 & ~n8508;
  assign n9160 = ~n8492 & ~n8507;
  assign n9161 = ~n39073 & ~n39074;
  assign n9162 = ~n8508 & ~n9156;
  assign n9163 = ~n9155 & ~n39075;
  assign n9164 = ~n8508 & ~n9163;
  assign n9165 = n8487 & ~n8489;
  assign n9166 = ~n8487 & ~n8490;
  assign n9167 = ~n8487 & ~n8489;
  assign n9168 = n8489 & ~n8490;
  assign n9169 = n8487 & n8489;
  assign n9170 = ~n39076 & ~n39077;
  assign n9171 = ~n8490 & ~n9165;
  assign n9172 = ~n9164 & ~n39078;
  assign n9173 = ~n8490 & ~n9172;
  assign n9174 = n8469 & ~n8471;
  assign n9175 = ~n8472 & ~n9174;
  assign n9176 = ~n9173 & n9175;
  assign n9177 = ~n8472 & ~n9176;
  assign n9178 = n8448 & n38942;
  assign n9179 = ~n8454 & ~n9178;
  assign n9180 = ~n9177 & n9179;
  assign n9181 = ~n8454 & ~n9180;
  assign n9182 = n8425 & n38938;
  assign n9183 = ~n8433 & ~n9182;
  assign n9184 = ~n9181 & n9183;
  assign n9185 = ~n8433 & ~n9184;
  assign n9186 = n8407 & ~n8409;
  assign n9187 = ~n8410 & ~n9186;
  assign n9188 = ~n9185 & n9187;
  assign n9189 = ~n8410 & ~n9188;
  assign n9190 = ~n8376 & n8391;
  assign n9191 = n8376 & ~n8392;
  assign n9192 = n8376 & n8391;
  assign n9193 = ~n8391 & ~n8392;
  assign n9194 = ~n8376 & ~n8391;
  assign n9195 = ~n39079 & ~n39080;
  assign n9196 = ~n8392 & ~n9190;
  assign n9197 = ~n9189 & ~n39081;
  assign n9198 = ~n8392 & ~n9197;
  assign n9199 = ~n8358 & n8373;
  assign n9200 = n8358 & ~n8374;
  assign n9201 = n8358 & n8373;
  assign n9202 = ~n8373 & ~n8374;
  assign n9203 = ~n8358 & ~n8373;
  assign n9204 = ~n39082 & ~n39083;
  assign n9205 = ~n8374 & ~n9199;
  assign n9206 = ~n9198 & ~n39084;
  assign n9207 = ~n8374 & ~n9206;
  assign n9208 = ~n8340 & n8355;
  assign n9209 = n8340 & ~n8356;
  assign n9210 = n8340 & n8355;
  assign n9211 = ~n8355 & ~n8356;
  assign n9212 = ~n8340 & ~n8355;
  assign n9213 = ~n39085 & ~n39086;
  assign n9214 = ~n8356 & ~n9208;
  assign n9215 = ~n9207 & ~n39087;
  assign n9216 = ~n8356 & ~n9215;
  assign n9217 = n8332 & n38920;
  assign n9218 = ~n8338 & ~n9217;
  assign n9219 = ~n9216 & n9218;
  assign n9220 = ~n8338 & ~n9219;
  assign n9221 = ~n8301 & n8316;
  assign n9222 = n8301 & ~n8317;
  assign n9223 = n8301 & n8316;
  assign n9224 = ~n8316 & ~n8317;
  assign n9225 = ~n8301 & ~n8316;
  assign n9226 = ~n39088 & ~n39089;
  assign n9227 = ~n8317 & ~n9221;
  assign n9228 = ~n9220 & ~n39090;
  assign n9229 = ~n8317 & ~n9228;
  assign n9230 = ~n8283 & n8298;
  assign n9231 = n8283 & ~n8299;
  assign n9232 = n8283 & n8298;
  assign n9233 = ~n8298 & ~n8299;
  assign n9234 = ~n8283 & ~n8298;
  assign n9235 = ~n39091 & ~n39092;
  assign n9236 = ~n8299 & ~n9230;
  assign n9237 = ~n9229 & ~n39093;
  assign n9238 = ~n8299 & ~n9237;
  assign n9239 = ~n8265 & n8280;
  assign n9240 = n8265 & ~n8281;
  assign n9241 = n8265 & n8280;
  assign n9242 = ~n8280 & ~n8281;
  assign n9243 = ~n8265 & ~n8280;
  assign n9244 = ~n39094 & ~n39095;
  assign n9245 = ~n8281 & ~n9239;
  assign n9246 = ~n9238 & ~n39096;
  assign n9247 = ~n8281 & ~n9246;
  assign n9248 = ~n8247 & n8262;
  assign n9249 = n8247 & ~n8263;
  assign n9250 = n8247 & n8262;
  assign n9251 = ~n8262 & ~n8263;
  assign n9252 = ~n8247 & ~n8262;
  assign n9253 = ~n39097 & ~n39098;
  assign n9254 = ~n8263 & ~n9248;
  assign n9255 = ~n9247 & ~n39099;
  assign n9256 = ~n8263 & ~n9255;
  assign n9257 = ~n8227 & n8244;
  assign n9258 = n8227 & ~n8245;
  assign n9259 = n8227 & n8244;
  assign n9260 = ~n8244 & ~n8245;
  assign n9261 = ~n8227 & ~n8244;
  assign n9262 = ~n39100 & ~n39101;
  assign n9263 = ~n8245 & ~n9257;
  assign n9264 = ~n9256 & ~n39102;
  assign n9265 = ~n8245 & ~n9264;
  assign n9266 = ~n8207 & n8224;
  assign n9267 = ~n8225 & ~n9266;
  assign n9268 = ~n9265 & n9267;
  assign n9269 = ~n8225 & ~n9268;
  assign n9270 = ~n8162 & n8204;
  assign n9271 = ~n8205 & ~n9270;
  assign n9272 = ~n9269 & ~n9270;
  assign n9273 = ~n8205 & n9272;
  assign n9274 = ~n9269 & n9271;
  assign n9275 = ~n8205 & ~n39103;
  assign n9276 = n489 & ~n491;
  assign n9277 = ~n492 & ~n9276;
  assign n9278 = n8175 & n9277;
  assign n9279 = pi106  & n38895;
  assign n9280 = pi108  & n8190;
  assign n9281 = pi107  & n8192;
  assign n9282 = ~n9280 & ~n9281;
  assign n9283 = ~n9279 & ~n9281;
  assign n9284 = ~n9280 & n9283;
  assign n9285 = ~n9279 & n9282;
  assign n9286 = ~n9278 & n39104;
  assign n9287 = pi17  & ~n9286;
  assign n9288 = pi17  & ~n9287;
  assign n9289 = pi17  & n9286;
  assign n9290 = ~n9286 & ~n9287;
  assign n9291 = ~pi17  & ~n9286;
  assign n9292 = ~n39105 & ~n39106;
  assign n9293 = ~n8152 & ~n8161;
  assign n9294 = ~n8124 & ~n8133;
  assign n9295 = ~n8098 & ~n8107;
  assign n9296 = ~n8077 & ~n8081;
  assign n9297 = n607 & n5281;
  assign n9298 = pi94  & n37489;
  assign n9299 = pi96  & n620;
  assign n9300 = pi95  & n622;
  assign n9301 = ~n9299 & ~n9300;
  assign n9302 = ~n9298 & ~n9300;
  assign n9303 = ~n9299 & n9302;
  assign n9304 = ~n9298 & n9301;
  assign n9305 = ~n9297 & n39107;
  assign n9306 = pi29  & ~n9305;
  assign n9307 = pi29  & ~n9306;
  assign n9308 = pi29  & n9305;
  assign n9309 = ~n9305 & ~n9306;
  assign n9310 = ~pi29  & ~n9305;
  assign n9311 = ~n39108 & ~n39109;
  assign n9312 = ~n8063 & ~n8071;
  assign n9313 = ~n8037 & ~n8046;
  assign n9314 = ~n8011 & ~n8020;
  assign n9315 = n636 & n691;
  assign n9316 = pi85  & n37503;
  assign n9317 = pi87  & n704;
  assign n9318 = pi86  & n706;
  assign n9319 = ~n9317 & ~n9318;
  assign n9320 = ~n9316 & ~n9318;
  assign n9321 = ~n9317 & n9320;
  assign n9322 = ~n9316 & n9319;
  assign n9323 = ~n9315 & n39110;
  assign n9324 = pi38  & ~n9323;
  assign n9325 = pi38  & ~n9324;
  assign n9326 = pi38  & n9323;
  assign n9327 = ~n9323 & ~n9324;
  assign n9328 = ~pi38  & ~n9323;
  assign n9329 = ~n39111 & ~n39112;
  assign n9330 = n733 & n2591;
  assign n9331 = pi82  & n37510;
  assign n9332 = pi84  & n746;
  assign n9333 = pi83  & n748;
  assign n9334 = ~n9332 & ~n9333;
  assign n9335 = ~n9331 & ~n9333;
  assign n9336 = ~n9332 & n9335;
  assign n9337 = ~n9331 & n9334;
  assign n9338 = ~n9330 & n39113;
  assign n9339 = pi41  & ~n9338;
  assign n9340 = pi41  & ~n9339;
  assign n9341 = pi41  & n9338;
  assign n9342 = ~n9338 & ~n9339;
  assign n9343 = ~pi41  & ~n9338;
  assign n9344 = ~n39114 & ~n39115;
  assign n9345 = ~n7973 & ~n7982;
  assign n9346 = n940 & n2154;
  assign n9347 = pi79  & n37541;
  assign n9348 = pi81  & n953;
  assign n9349 = pi80  & n955;
  assign n9350 = ~n9348 & ~n9349;
  assign n9351 = ~n9347 & ~n9349;
  assign n9352 = ~n9348 & n9351;
  assign n9353 = ~n9347 & n9350;
  assign n9354 = ~n9346 & n39116;
  assign n9355 = pi44  & ~n9354;
  assign n9356 = pi44  & ~n9355;
  assign n9357 = pi44  & n9354;
  assign n9358 = ~n9354 & ~n9355;
  assign n9359 = ~pi44  & ~n9354;
  assign n9360 = ~n39117 & ~n39118;
  assign n9361 = ~n7935 & ~n7944;
  assign n9362 = n720 & n894;
  assign n9363 = pi73  & n37580;
  assign n9364 = pi75  & n896;
  assign n9365 = pi74  & n904;
  assign n9366 = ~n9364 & ~n9365;
  assign n9367 = ~n9363 & ~n9365;
  assign n9368 = ~n9364 & n9367;
  assign n9369 = ~n9363 & n9366;
  assign n9370 = ~n9362 & n39119;
  assign n9371 = pi50  & ~n9370;
  assign n9372 = pi50  & ~n9371;
  assign n9373 = pi50  & n9370;
  assign n9374 = ~n9370 & ~n9371;
  assign n9375 = ~pi50  & ~n9370;
  assign n9376 = ~n39120 & ~n39121;
  assign n9377 = ~n7915 & ~n7917;
  assign n9378 = n1124 & n1971;
  assign n9379 = pi70  & n37864;
  assign n9380 = pi72  & n1973;
  assign n9381 = pi71  & n1981;
  assign n9382 = ~n9380 & ~n9381;
  assign n9383 = ~n9379 & ~n9381;
  assign n9384 = ~n9380 & n9383;
  assign n9385 = ~n9379 & n9382;
  assign n9386 = ~n9378 & n39122;
  assign n9387 = pi53  & ~n9386;
  assign n9388 = pi53  & ~n9387;
  assign n9389 = pi53  & n9386;
  assign n9390 = ~n9386 & ~n9387;
  assign n9391 = ~pi53  & ~n9386;
  assign n9392 = ~n39123 & ~n39124;
  assign n9393 = ~n7909 & ~n7911;
  assign n9394 = n990 & n4312;
  assign n9395 = pi67  & n38376;
  assign n9396 = pi69  & n4314;
  assign n9397 = pi68  & n4322;
  assign n9398 = ~n9396 & ~n9397;
  assign n9399 = ~n9395 & ~n9397;
  assign n9400 = ~n9396 & n9399;
  assign n9401 = ~n9395 & n9398;
  assign n9402 = ~n9394 & n39125;
  assign n9403 = pi56  & ~n9402;
  assign n9404 = pi56  & ~n9403;
  assign n9405 = pi56  & n9402;
  assign n9406 = ~n9402 & ~n9403;
  assign n9407 = ~pi56  & ~n9402;
  assign n9408 = ~n39126 & ~n39127;
  assign n9409 = pi59  & ~n38837;
  assign n9410 = ~n38599 & n38835;
  assign n9411 = ~n38599 & ~n38836;
  assign n9412 = n38835 & n9411;
  assign n9413 = ~n38836 & n9410;
  assign n9414 = pi64  & n39128;
  assign n9415 = pi65  & n7892;
  assign n9416 = ~n37521 & n7882;
  assign n9417 = pi66  & n7884;
  assign n9418 = ~n9416 & ~n9417;
  assign n9419 = ~n9415 & ~n9416;
  assign n9420 = ~n9417 & n9419;
  assign n9421 = ~n9415 & ~n9417;
  assign n9422 = ~n9416 & n9421;
  assign n9423 = ~n9415 & n9418;
  assign n9424 = ~n9414 & ~n9415;
  assign n9425 = ~n9417 & n9424;
  assign n9426 = ~n9414 & n9421;
  assign n9427 = ~n9416 & n39130;
  assign n9428 = ~n9414 & n39129;
  assign n9429 = ~n9409 & n39131;
  assign n9430 = n9409 & ~n39131;
  assign n9431 = pi59  & ~n39131;
  assign n9432 = pi59  & ~n9431;
  assign n9433 = ~n39131 & ~n9431;
  assign n9434 = ~n9432 & ~n9433;
  assign n9435 = n38837 & ~n9434;
  assign n9436 = n38837 & n39131;
  assign n9437 = ~n38837 & n9434;
  assign n9438 = ~n39132 & ~n9437;
  assign n9439 = ~n9429 & ~n9430;
  assign n9440 = ~n9408 & n39133;
  assign n9441 = n9408 & ~n39133;
  assign n9442 = ~n9440 & ~n9441;
  assign n9443 = ~n9393 & ~n9441;
  assign n9444 = ~n9440 & n9443;
  assign n9445 = ~n9393 & n9442;
  assign n9446 = n9393 & ~n9442;
  assign n9447 = ~n9393 & ~n39134;
  assign n9448 = ~n9440 & ~n39134;
  assign n9449 = ~n9441 & n9448;
  assign n9450 = ~n9447 & ~n9449;
  assign n9451 = ~n39134 & ~n9446;
  assign n9452 = n9392 & n39135;
  assign n9453 = ~n9392 & ~n39135;
  assign n9454 = ~n9452 & ~n9453;
  assign n9455 = ~n9377 & n9454;
  assign n9456 = n9377 & ~n9454;
  assign n9457 = ~n9455 & ~n9456;
  assign n9458 = n9376 & ~n9457;
  assign n9459 = ~n9376 & n9457;
  assign n9460 = ~n9458 & ~n9459;
  assign n9461 = ~n9361 & n9460;
  assign n9462 = n9361 & ~n9460;
  assign n9463 = ~n9461 & ~n9462;
  assign n9464 = n785 & n1578;
  assign n9465 = pi76  & n37520;
  assign n9466 = pi78  & n787;
  assign n9467 = pi77  & n795;
  assign n9468 = ~n9466 & ~n9467;
  assign n9469 = ~n9465 & ~n9467;
  assign n9470 = ~n9466 & n9469;
  assign n9471 = ~n9465 & n9468;
  assign n9472 = ~n9464 & n39136;
  assign n9473 = pi47  & ~n9472;
  assign n9474 = pi47  & ~n9473;
  assign n9475 = pi47  & n9472;
  assign n9476 = ~n9472 & ~n9473;
  assign n9477 = ~pi47  & ~n9472;
  assign n9478 = ~n39137 & ~n39138;
  assign n9479 = n9463 & ~n9478;
  assign n9480 = ~n9463 & n9478;
  assign n9481 = n9463 & ~n9479;
  assign n9482 = n9463 & n9478;
  assign n9483 = ~n9478 & ~n9479;
  assign n9484 = ~n9463 & ~n9478;
  assign n9485 = ~n39139 & ~n39140;
  assign n9486 = ~n9479 & ~n9480;
  assign n9487 = ~n7969 & ~n39141;
  assign n9488 = n7969 & n39141;
  assign n9489 = ~n9487 & ~n9488;
  assign n9490 = ~n9360 & n9489;
  assign n9491 = n9360 & ~n9489;
  assign n9492 = ~n9360 & ~n9490;
  assign n9493 = ~n9360 & ~n9489;
  assign n9494 = n9489 & ~n9490;
  assign n9495 = n9360 & n9489;
  assign n9496 = ~n39142 & ~n39143;
  assign n9497 = ~n9490 & ~n9491;
  assign n9498 = ~n9345 & ~n39144;
  assign n9499 = n9345 & n39144;
  assign n9500 = ~n9345 & ~n9498;
  assign n9501 = ~n9345 & n39144;
  assign n9502 = ~n39144 & ~n9498;
  assign n9503 = n9345 & ~n39144;
  assign n9504 = ~n39145 & ~n39146;
  assign n9505 = ~n9498 & ~n9499;
  assign n9506 = ~n9344 & ~n39147;
  assign n9507 = n9344 & n39147;
  assign n9508 = ~n39147 & ~n9506;
  assign n9509 = ~n9344 & ~n9506;
  assign n9510 = ~n9508 & ~n9509;
  assign n9511 = ~n9506 & ~n9507;
  assign n9512 = ~n8007 & ~n39148;
  assign n9513 = n8007 & n39148;
  assign n9514 = ~n8007 & n39148;
  assign n9515 = n8007 & ~n39148;
  assign n9516 = ~n9514 & ~n9515;
  assign n9517 = ~n9512 & ~n9513;
  assign n9518 = ~n9329 & ~n39149;
  assign n9519 = n9329 & n39149;
  assign n9520 = ~n9518 & ~n9519;
  assign n9521 = n9314 & ~n9520;
  assign n9522 = ~n9314 & n9520;
  assign n9523 = ~n9521 & ~n9522;
  assign n9524 = n2104 & n3566;
  assign n9525 = pi88  & n37758;
  assign n9526 = pi90  & n2117;
  assign n9527 = pi89  & n2119;
  assign n9528 = ~n9526 & ~n9527;
  assign n9529 = ~n9525 & ~n9527;
  assign n9530 = ~n9526 & n9529;
  assign n9531 = ~n9525 & n9528;
  assign n9532 = ~n9524 & n39150;
  assign n9533 = pi35  & ~n9532;
  assign n9534 = pi35  & ~n9533;
  assign n9535 = pi35  & n9532;
  assign n9536 = ~n9532 & ~n9533;
  assign n9537 = ~pi35  & ~n9532;
  assign n9538 = ~n39151 & ~n39152;
  assign n9539 = n9523 & ~n9538;
  assign n9540 = ~n9523 & n9538;
  assign n9541 = n9523 & ~n9539;
  assign n9542 = n9523 & n9538;
  assign n9543 = ~n9538 & ~n9539;
  assign n9544 = ~n9523 & ~n9538;
  assign n9545 = ~n39153 & ~n39154;
  assign n9546 = ~n9539 & ~n9540;
  assign n9547 = n9313 & n39155;
  assign n9548 = ~n9313 & ~n39155;
  assign n9549 = ~n9547 & ~n9548;
  assign n9550 = n649 & n4544;
  assign n9551 = pi91  & n37496;
  assign n9552 = pi93  & n662;
  assign n9553 = pi92  & n664;
  assign n9554 = ~n9552 & ~n9553;
  assign n9555 = ~n9551 & ~n9553;
  assign n9556 = ~n9552 & n9555;
  assign n9557 = ~n9551 & n9554;
  assign n9558 = ~n9550 & n39156;
  assign n9559 = pi32  & ~n9558;
  assign n9560 = pi32  & ~n9559;
  assign n9561 = pi32  & n9558;
  assign n9562 = ~n9558 & ~n9559;
  assign n9563 = ~pi32  & ~n9558;
  assign n9564 = ~n39157 & ~n39158;
  assign n9565 = n9549 & ~n9564;
  assign n9566 = ~n9549 & n9564;
  assign n9567 = ~n9565 & ~n9566;
  assign n9568 = ~n9312 & ~n9566;
  assign n9569 = ~n9565 & n9568;
  assign n9570 = ~n9312 & n9567;
  assign n9571 = n9312 & ~n9567;
  assign n9572 = ~n9312 & ~n39159;
  assign n9573 = ~n9565 & ~n39159;
  assign n9574 = ~n9566 & n9573;
  assign n9575 = ~n9572 & ~n9574;
  assign n9576 = ~n39159 & ~n9571;
  assign n9577 = n9311 & n39160;
  assign n9578 = ~n9311 & ~n39160;
  assign n9579 = ~n9577 & ~n9578;
  assign n9580 = ~n9296 & n9579;
  assign n9581 = n9296 & ~n9579;
  assign n9582 = ~n9580 & ~n9581;
  assign n9583 = n4492 & n5578;
  assign n9584 = pi97  & n38208;
  assign n9585 = pi99  & n4507;
  assign n9586 = pi98  & n4509;
  assign n9587 = ~n9585 & ~n9586;
  assign n9588 = ~n9584 & ~n9586;
  assign n9589 = ~n9585 & n9588;
  assign n9590 = ~n9584 & n9587;
  assign n9591 = ~n9583 & n39161;
  assign n9592 = pi26  & ~n9591;
  assign n9593 = pi26  & ~n9592;
  assign n9594 = pi26  & n9591;
  assign n9595 = ~n9591 & ~n9592;
  assign n9596 = ~pi26  & ~n9591;
  assign n9597 = ~n39162 & ~n39163;
  assign n9598 = n9582 & ~n9597;
  assign n9599 = ~n9582 & n9597;
  assign n9600 = n9582 & ~n9598;
  assign n9601 = n9582 & n9597;
  assign n9602 = ~n9597 & ~n9598;
  assign n9603 = ~n9582 & ~n9597;
  assign n9604 = ~n39164 & ~n39165;
  assign n9605 = ~n9598 & ~n9599;
  assign n9606 = n9295 & n39166;
  assign n9607 = ~n9295 & ~n39166;
  assign n9608 = ~n9606 & ~n9607;
  assign n9609 = n5576 & n6819;
  assign n9610 = pi100  & n38406;
  assign n9611 = pi102  & n5591;
  assign n9612 = pi101  & n5593;
  assign n9613 = ~n9611 & ~n9612;
  assign n9614 = ~n9610 & ~n9612;
  assign n9615 = ~n9611 & n9614;
  assign n9616 = ~n9610 & n9613;
  assign n9617 = ~n9609 & n39167;
  assign n9618 = pi23  & ~n9617;
  assign n9619 = pi23  & ~n9618;
  assign n9620 = pi23  & n9617;
  assign n9621 = ~n9617 & ~n9618;
  assign n9622 = ~pi23  & ~n9617;
  assign n9623 = ~n39168 & ~n39169;
  assign n9624 = n9608 & ~n9623;
  assign n9625 = ~n9608 & n9623;
  assign n9626 = n9608 & ~n9624;
  assign n9627 = n9608 & n9623;
  assign n9628 = ~n9623 & ~n9624;
  assign n9629 = ~n9608 & ~n9623;
  assign n9630 = ~n39170 & ~n39171;
  assign n9631 = ~n9624 & ~n9625;
  assign n9632 = n9294 & n39172;
  assign n9633 = ~n9294 & ~n39172;
  assign n9634 = ~n9632 & ~n9633;
  assign n9635 = n6785 & n8229;
  assign n9636 = pi103  & n38631;
  assign n9637 = pi105  & n6800;
  assign n9638 = pi104  & n6802;
  assign n9639 = ~n9637 & ~n9638;
  assign n9640 = ~n9636 & ~n9638;
  assign n9641 = ~n9637 & n9640;
  assign n9642 = ~n9636 & n9639;
  assign n9643 = ~n9635 & n39173;
  assign n9644 = pi20  & ~n9643;
  assign n9645 = pi20  & ~n9644;
  assign n9646 = pi20  & n9643;
  assign n9647 = ~n9643 & ~n9644;
  assign n9648 = ~pi20  & ~n9643;
  assign n9649 = ~n39174 & ~n39175;
  assign n9650 = n9634 & ~n9649;
  assign n9651 = ~n9634 & n9649;
  assign n9652 = ~n9650 & ~n9651;
  assign n9653 = ~n9293 & ~n9651;
  assign n9654 = ~n9650 & n9653;
  assign n9655 = ~n9293 & n9652;
  assign n9656 = n9293 & ~n9652;
  assign n9657 = ~n9293 & ~n39176;
  assign n9658 = ~n9650 & ~n39176;
  assign n9659 = ~n9651 & n9658;
  assign n9660 = ~n9657 & ~n9659;
  assign n9661 = ~n39176 & ~n9656;
  assign n9662 = ~n9292 & ~n39177;
  assign n9663 = n9292 & n39177;
  assign n9664 = ~n39177 & ~n9662;
  assign n9665 = n9292 & ~n39177;
  assign n9666 = ~n9292 & ~n9662;
  assign n9667 = ~n9292 & n39177;
  assign n9668 = ~n39178 & ~n39179;
  assign n9669 = ~n9662 & ~n9663;
  assign n9670 = ~n9275 & ~n39180;
  assign n9671 = n9275 & n39180;
  assign n9672 = ~n9275 & n39180;
  assign n9673 = n9275 & ~n39180;
  assign n9674 = ~n9672 & ~n9673;
  assign n9675 = ~n9670 & ~n9671;
  assign n9676 = ~n592 & ~n39181;
  assign n9677 = n497 & ~n499;
  assign n9678 = ~n500 & ~n9677;
  assign n9679 = n563 & n9678;
  assign n9680 = pi108  & n37482;
  assign n9681 = pi110  & n578;
  assign n9682 = pi109  & n580;
  assign n9683 = ~n9681 & ~n9682;
  assign n9684 = ~n9680 & ~n9682;
  assign n9685 = ~n9681 & n9684;
  assign n9686 = ~n9680 & n9683;
  assign n9687 = ~n9679 & n39182;
  assign n9688 = pi14  & ~n9687;
  assign n9689 = pi14  & ~n9688;
  assign n9690 = pi14  & n9687;
  assign n9691 = ~n9687 & ~n9688;
  assign n9692 = ~pi14  & ~n9687;
  assign n9693 = ~n39183 & ~n39184;
  assign n9694 = n9269 & ~n9271;
  assign n9695 = ~n9269 & ~n39103;
  assign n9696 = ~n9270 & n9275;
  assign n9697 = ~n9695 & ~n9696;
  assign n9698 = ~n39103 & ~n9694;
  assign n9699 = ~n9693 & ~n39185;
  assign n9700 = n493 & ~n495;
  assign n9701 = ~n496 & ~n9700;
  assign n9702 = n563 & n9701;
  assign n9703 = pi107  & n37482;
  assign n9704 = pi109  & n578;
  assign n9705 = pi108  & n580;
  assign n9706 = ~n9704 & ~n9705;
  assign n9707 = ~n9703 & ~n9705;
  assign n9708 = ~n9704 & n9707;
  assign n9709 = ~n9703 & n9706;
  assign n9710 = ~n9702 & n39186;
  assign n9711 = pi14  & ~n9710;
  assign n9712 = pi14  & ~n9711;
  assign n9713 = pi14  & n9710;
  assign n9714 = ~n9710 & ~n9711;
  assign n9715 = ~pi14  & ~n9710;
  assign n9716 = ~n39187 & ~n39188;
  assign n9717 = n9265 & ~n9267;
  assign n9718 = ~n9268 & ~n9717;
  assign n9719 = ~n9716 & n9718;
  assign n9720 = n9256 & n39102;
  assign n9721 = ~n9264 & ~n9720;
  assign n9722 = n563 & n9277;
  assign n9723 = pi106  & n37482;
  assign n9724 = pi108  & n578;
  assign n9725 = pi107  & n580;
  assign n9726 = ~n9724 & ~n9725;
  assign n9727 = ~n9723 & ~n9725;
  assign n9728 = ~n9724 & n9727;
  assign n9729 = ~n9723 & n9726;
  assign n9730 = ~n9722 & n39189;
  assign n9731 = pi14  & ~n9730;
  assign n9732 = pi14  & ~n9731;
  assign n9733 = pi14  & n9730;
  assign n9734 = ~n9730 & ~n9731;
  assign n9735 = ~pi14  & ~n9730;
  assign n9736 = ~n39190 & ~n39191;
  assign n9737 = n9721 & ~n9736;
  assign n9738 = n9247 & n39099;
  assign n9739 = ~n9255 & ~n9738;
  assign n9740 = n563 & n8177;
  assign n9741 = pi105  & n37482;
  assign n9742 = pi107  & n578;
  assign n9743 = pi106  & n580;
  assign n9744 = ~n9742 & ~n9743;
  assign n9745 = ~n9741 & ~n9743;
  assign n9746 = ~n9742 & n9745;
  assign n9747 = ~n9741 & n9744;
  assign n9748 = ~n9740 & n39192;
  assign n9749 = pi14  & ~n9748;
  assign n9750 = pi14  & ~n9749;
  assign n9751 = pi14  & n9748;
  assign n9752 = ~n9748 & ~n9749;
  assign n9753 = ~pi14  & ~n9748;
  assign n9754 = ~n39193 & ~n39194;
  assign n9755 = n9739 & ~n9754;
  assign n9756 = n9238 & n39096;
  assign n9757 = ~n9246 & ~n9756;
  assign n9758 = n563 & n8209;
  assign n9759 = pi104  & n37482;
  assign n9760 = pi106  & n578;
  assign n9761 = pi105  & n580;
  assign n9762 = ~n9760 & ~n9761;
  assign n9763 = ~n9759 & ~n9761;
  assign n9764 = ~n9760 & n9763;
  assign n9765 = ~n9759 & n9762;
  assign n9766 = ~n9758 & n39195;
  assign n9767 = pi14  & ~n9766;
  assign n9768 = pi14  & ~n9767;
  assign n9769 = pi14  & n9766;
  assign n9770 = ~n9766 & ~n9767;
  assign n9771 = ~pi14  & ~n9766;
  assign n9772 = ~n39196 & ~n39197;
  assign n9773 = n9757 & ~n9772;
  assign n9774 = n9229 & n39093;
  assign n9775 = ~n9237 & ~n9774;
  assign n9776 = n563 & n8229;
  assign n9777 = pi103  & n37482;
  assign n9778 = pi105  & n578;
  assign n9779 = pi104  & n580;
  assign n9780 = ~n9778 & ~n9779;
  assign n9781 = ~n9777 & ~n9779;
  assign n9782 = ~n9778 & n9781;
  assign n9783 = ~n9777 & n9780;
  assign n9784 = ~n9776 & n39198;
  assign n9785 = pi14  & ~n9784;
  assign n9786 = pi14  & ~n9785;
  assign n9787 = pi14  & n9784;
  assign n9788 = ~n9784 & ~n9785;
  assign n9789 = ~pi14  & ~n9784;
  assign n9790 = ~n39199 & ~n39200;
  assign n9791 = n9775 & ~n9790;
  assign n9792 = n9220 & n39090;
  assign n9793 = ~n9228 & ~n9792;
  assign n9794 = n563 & n8136;
  assign n9795 = pi102  & n37482;
  assign n9796 = pi104  & n578;
  assign n9797 = pi103  & n580;
  assign n9798 = ~n9796 & ~n9797;
  assign n9799 = ~n9795 & ~n9797;
  assign n9800 = ~n9796 & n9799;
  assign n9801 = ~n9795 & n9798;
  assign n9802 = ~n9794 & n39201;
  assign n9803 = pi14  & ~n9802;
  assign n9804 = pi14  & ~n9803;
  assign n9805 = pi14  & n9802;
  assign n9806 = ~n9802 & ~n9803;
  assign n9807 = ~pi14  & ~n9802;
  assign n9808 = ~n39202 & ~n39203;
  assign n9809 = n9793 & ~n9808;
  assign n9810 = n9216 & ~n9218;
  assign n9811 = ~n9219 & ~n9810;
  assign n9812 = n563 & n6787;
  assign n9813 = pi101  & n37482;
  assign n9814 = pi103  & n578;
  assign n9815 = pi102  & n580;
  assign n9816 = ~n9814 & ~n9815;
  assign n9817 = ~n9813 & ~n9815;
  assign n9818 = ~n9814 & n9817;
  assign n9819 = ~n9813 & n9816;
  assign n9820 = ~n9812 & n39204;
  assign n9821 = pi14  & ~n9820;
  assign n9822 = pi14  & ~n9821;
  assign n9823 = pi14  & n9820;
  assign n9824 = ~n9820 & ~n9821;
  assign n9825 = ~pi14  & ~n9820;
  assign n9826 = ~n39205 & ~n39206;
  assign n9827 = n9811 & ~n9826;
  assign n9828 = n9207 & n39087;
  assign n9829 = ~n9215 & ~n9828;
  assign n9830 = n563 & n6819;
  assign n9831 = pi100  & n37482;
  assign n9832 = pi102  & n578;
  assign n9833 = pi101  & n580;
  assign n9834 = ~n9832 & ~n9833;
  assign n9835 = ~n9831 & ~n9833;
  assign n9836 = ~n9832 & n9835;
  assign n9837 = ~n9831 & n9834;
  assign n9838 = ~n9830 & n39207;
  assign n9839 = pi14  & ~n9838;
  assign n9840 = pi14  & ~n9839;
  assign n9841 = pi14  & n9838;
  assign n9842 = ~n9838 & ~n9839;
  assign n9843 = ~pi14  & ~n9838;
  assign n9844 = ~n39208 & ~n39209;
  assign n9845 = n9829 & ~n9844;
  assign n9846 = n9198 & n39084;
  assign n9847 = ~n9206 & ~n9846;
  assign n9848 = n563 & n6839;
  assign n9849 = pi99  & n37482;
  assign n9850 = pi101  & n578;
  assign n9851 = pi100  & n580;
  assign n9852 = ~n9850 & ~n9851;
  assign n9853 = ~n9849 & ~n9851;
  assign n9854 = ~n9850 & n9853;
  assign n9855 = ~n9849 & n9852;
  assign n9856 = ~n9848 & n39210;
  assign n9857 = pi14  & ~n9856;
  assign n9858 = pi14  & ~n9857;
  assign n9859 = pi14  & n9856;
  assign n9860 = ~n9856 & ~n9857;
  assign n9861 = ~pi14  & ~n9856;
  assign n9862 = ~n39211 & ~n39212;
  assign n9863 = n9847 & ~n9862;
  assign n9864 = n563 & n6474;
  assign n9865 = pi98  & n37482;
  assign n9866 = pi100  & n578;
  assign n9867 = pi99  & n580;
  assign n9868 = ~n9866 & ~n9867;
  assign n9869 = ~n9865 & ~n9867;
  assign n9870 = ~n9866 & n9869;
  assign n9871 = ~n9865 & n9868;
  assign n9872 = ~n9864 & n39213;
  assign n9873 = pi14  & ~n9872;
  assign n9874 = pi14  & ~n9873;
  assign n9875 = pi14  & n9872;
  assign n9876 = ~n9872 & ~n9873;
  assign n9877 = ~pi14  & ~n9872;
  assign n9878 = ~n39214 & ~n39215;
  assign n9879 = n9189 & n39081;
  assign n9880 = ~n9189 & n39081;
  assign n9881 = n9189 & ~n39081;
  assign n9882 = ~n9880 & ~n9881;
  assign n9883 = ~n9197 & ~n9879;
  assign n9884 = ~n9878 & ~n39216;
  assign n9885 = n9185 & ~n9187;
  assign n9886 = ~n9188 & ~n9885;
  assign n9887 = n563 & n5578;
  assign n9888 = pi97  & n37482;
  assign n9889 = pi99  & n578;
  assign n9890 = pi98  & n580;
  assign n9891 = ~n9889 & ~n9890;
  assign n9892 = ~n9888 & ~n9890;
  assign n9893 = ~n9889 & n9892;
  assign n9894 = ~n9888 & n9891;
  assign n9895 = ~n9887 & n39217;
  assign n9896 = pi14  & ~n9895;
  assign n9897 = pi14  & ~n9896;
  assign n9898 = pi14  & n9895;
  assign n9899 = ~n9895 & ~n9896;
  assign n9900 = ~pi14  & ~n9895;
  assign n9901 = ~n39218 & ~n39219;
  assign n9902 = n9886 & ~n9901;
  assign n9903 = n9181 & ~n9183;
  assign n9904 = ~n9184 & ~n9903;
  assign n9905 = n563 & n5610;
  assign n9906 = pi96  & n37482;
  assign n9907 = pi98  & n578;
  assign n9908 = pi97  & n580;
  assign n9909 = ~n9907 & ~n9908;
  assign n9910 = ~n9906 & ~n9908;
  assign n9911 = ~n9907 & n9910;
  assign n9912 = ~n9906 & n9909;
  assign n9913 = ~n9905 & n39220;
  assign n9914 = pi14  & ~n9913;
  assign n9915 = pi14  & ~n9914;
  assign n9916 = pi14  & n9913;
  assign n9917 = ~n9913 & ~n9914;
  assign n9918 = ~pi14  & ~n9913;
  assign n9919 = ~n39221 & ~n39222;
  assign n9920 = n9904 & ~n9919;
  assign n9921 = n9177 & ~n9179;
  assign n9922 = ~n9180 & ~n9921;
  assign n9923 = n563 & n5630;
  assign n9924 = pi95  & n37482;
  assign n9925 = pi97  & n578;
  assign n9926 = pi96  & n580;
  assign n9927 = ~n9925 & ~n9926;
  assign n9928 = ~n9924 & ~n9926;
  assign n9929 = ~n9925 & n9928;
  assign n9930 = ~n9924 & n9927;
  assign n9931 = ~n9923 & n39223;
  assign n9932 = pi14  & ~n9931;
  assign n9933 = pi14  & ~n9932;
  assign n9934 = pi14  & n9931;
  assign n9935 = ~n9931 & ~n9932;
  assign n9936 = ~pi14  & ~n9931;
  assign n9937 = ~n39224 & ~n39225;
  assign n9938 = n9922 & ~n9937;
  assign n9939 = n563 & n5281;
  assign n9940 = pi94  & n37482;
  assign n9941 = pi96  & n578;
  assign n9942 = pi95  & n580;
  assign n9943 = ~n9941 & ~n9942;
  assign n9944 = ~n9940 & ~n9942;
  assign n9945 = ~n9941 & n9944;
  assign n9946 = ~n9940 & n9943;
  assign n9947 = ~n9939 & n39226;
  assign n9948 = pi14  & ~n9947;
  assign n9949 = pi14  & ~n9948;
  assign n9950 = pi14  & n9947;
  assign n9951 = ~n9947 & ~n9948;
  assign n9952 = ~pi14  & ~n9947;
  assign n9953 = ~n39227 & ~n39228;
  assign n9954 = n9173 & ~n9175;
  assign n9955 = ~n9176 & ~n9954;
  assign n9956 = ~n9953 & n9955;
  assign n9957 = n563 & n4494;
  assign n9958 = pi93  & n37482;
  assign n9959 = pi95  & n578;
  assign n9960 = pi94  & n580;
  assign n9961 = ~n9959 & ~n9960;
  assign n9962 = ~n9958 & ~n9960;
  assign n9963 = ~n9959 & n9962;
  assign n9964 = ~n9958 & n9961;
  assign n9965 = ~n9957 & n39229;
  assign n9966 = pi14  & ~n9965;
  assign n9967 = pi14  & ~n9966;
  assign n9968 = pi14  & n9965;
  assign n9969 = ~n9965 & ~n9966;
  assign n9970 = ~pi14  & ~n9965;
  assign n9971 = ~n39230 & ~n39231;
  assign n9972 = n9164 & n39078;
  assign n9973 = ~n9164 & ~n9172;
  assign n9974 = ~n9164 & n39078;
  assign n9975 = ~n39078 & ~n9172;
  assign n9976 = n9164 & ~n39078;
  assign n9977 = ~n39232 & ~n39233;
  assign n9978 = ~n9172 & ~n9972;
  assign n9979 = ~n9971 & ~n39234;
  assign n9980 = n563 & n4524;
  assign n9981 = pi92  & n37482;
  assign n9982 = pi94  & n578;
  assign n9983 = pi93  & n580;
  assign n9984 = ~n9982 & ~n9983;
  assign n9985 = ~n9981 & ~n9983;
  assign n9986 = ~n9982 & n9985;
  assign n9987 = ~n9981 & n9984;
  assign n9988 = ~n9980 & n39235;
  assign n9989 = pi14  & ~n9988;
  assign n9990 = pi14  & ~n9989;
  assign n9991 = pi14  & n9988;
  assign n9992 = ~n9988 & ~n9989;
  assign n9993 = ~pi14  & ~n9988;
  assign n9994 = ~n39236 & ~n39237;
  assign n9995 = n9155 & n39075;
  assign n9996 = ~n9155 & n39075;
  assign n9997 = n9155 & ~n39075;
  assign n9998 = ~n9996 & ~n9997;
  assign n9999 = ~n9163 & ~n9995;
  assign n10000 = ~n9994 & ~n39238;
  assign n10001 = n563 & n4544;
  assign n10002 = pi91  & n37482;
  assign n10003 = pi93  & n578;
  assign n10004 = pi92  & n580;
  assign n10005 = ~n10003 & ~n10004;
  assign n10006 = ~n10002 & ~n10004;
  assign n10007 = ~n10003 & n10006;
  assign n10008 = ~n10002 & n10005;
  assign n10009 = ~n10001 & n39239;
  assign n10010 = pi14  & ~n10009;
  assign n10011 = pi14  & ~n10010;
  assign n10012 = pi14  & n10009;
  assign n10013 = ~n10009 & ~n10010;
  assign n10014 = ~pi14  & ~n10009;
  assign n10015 = ~n39240 & ~n39241;
  assign n10016 = n9151 & ~n9153;
  assign n10017 = ~n9154 & ~n10016;
  assign n10018 = ~n10015 & n10017;
  assign n10019 = n563 & n4453;
  assign n10020 = pi90  & n37482;
  assign n10021 = pi92  & n578;
  assign n10022 = pi91  & n580;
  assign n10023 = ~n10021 & ~n10022;
  assign n10024 = ~n10020 & ~n10022;
  assign n10025 = ~n10021 & n10024;
  assign n10026 = ~n10020 & n10023;
  assign n10027 = ~n10019 & n39242;
  assign n10028 = pi14  & ~n10027;
  assign n10029 = pi14  & ~n10028;
  assign n10030 = pi14  & n10027;
  assign n10031 = ~n10027 & ~n10028;
  assign n10032 = ~pi14  & ~n10027;
  assign n10033 = ~n39243 & ~n39244;
  assign n10034 = n9142 & n39072;
  assign n10035 = ~n9150 & ~n10034;
  assign n10036 = ~n10033 & n10035;
  assign n10037 = n9138 & ~n9140;
  assign n10038 = ~n9141 & ~n10037;
  assign n10039 = n563 & n594;
  assign n10040 = pi89  & n37482;
  assign n10041 = pi91  & n578;
  assign n10042 = pi90  & n580;
  assign n10043 = ~n10041 & ~n10042;
  assign n10044 = ~n10040 & ~n10042;
  assign n10045 = ~n10041 & n10044;
  assign n10046 = ~n10040 & n10043;
  assign n10047 = ~n10039 & n39245;
  assign n10048 = pi14  & ~n10047;
  assign n10049 = pi14  & ~n10048;
  assign n10050 = pi14  & n10047;
  assign n10051 = ~n10047 & ~n10048;
  assign n10052 = ~pi14  & ~n10047;
  assign n10053 = ~n39246 & ~n39247;
  assign n10054 = n10038 & ~n10053;
  assign n10055 = n563 & n3566;
  assign n10056 = pi88  & n37482;
  assign n10057 = pi90  & n578;
  assign n10058 = pi89  & n580;
  assign n10059 = ~n10057 & ~n10058;
  assign n10060 = ~n10056 & ~n10058;
  assign n10061 = ~n10057 & n10060;
  assign n10062 = ~n10056 & n10059;
  assign n10063 = ~n10055 & n39248;
  assign n10064 = pi14  & ~n10063;
  assign n10065 = pi14  & ~n10064;
  assign n10066 = pi14  & n10063;
  assign n10067 = ~n10063 & ~n10064;
  assign n10068 = ~pi14  & ~n10063;
  assign n10069 = ~n39249 & ~n39250;
  assign n10070 = n9132 & ~n9134;
  assign n10071 = ~n9132 & ~n39069;
  assign n10072 = ~n9133 & n9138;
  assign n10073 = ~n10071 & ~n10072;
  assign n10074 = ~n39069 & ~n10070;
  assign n10075 = ~n10069 & ~n39251;
  assign n10076 = n9123 & n39068;
  assign n10077 = ~n9131 & ~n10076;
  assign n10078 = n563 & n3591;
  assign n10079 = pi87  & n37482;
  assign n10080 = pi89  & n578;
  assign n10081 = pi88  & n580;
  assign n10082 = ~n10080 & ~n10081;
  assign n10083 = ~n10079 & ~n10081;
  assign n10084 = ~n10080 & n10083;
  assign n10085 = ~n10079 & n10082;
  assign n10086 = ~n10078 & n39252;
  assign n10087 = pi14  & ~n10086;
  assign n10088 = pi14  & ~n10087;
  assign n10089 = pi14  & n10086;
  assign n10090 = ~n10086 & ~n10087;
  assign n10091 = ~pi14  & ~n10086;
  assign n10092 = ~n39253 & ~n39254;
  assign n10093 = n10077 & ~n10092;
  assign n10094 = n563 & n3354;
  assign n10095 = pi86  & n37482;
  assign n10096 = pi88  & n578;
  assign n10097 = pi87  & n580;
  assign n10098 = ~n10096 & ~n10097;
  assign n10099 = ~n10095 & ~n10097;
  assign n10100 = ~n10096 & n10099;
  assign n10101 = ~n10095 & n10098;
  assign n10102 = ~n10094 & n39255;
  assign n10103 = pi14  & ~n10102;
  assign n10104 = pi14  & ~n10103;
  assign n10105 = pi14  & n10102;
  assign n10106 = ~n10102 & ~n10103;
  assign n10107 = ~pi14  & ~n10102;
  assign n10108 = ~n39256 & ~n39257;
  assign n10109 = n9114 & n39065;
  assign n10110 = ~n9114 & n39065;
  assign n10111 = n9114 & ~n39065;
  assign n10112 = ~n10110 & ~n10111;
  assign n10113 = ~n9122 & ~n10109;
  assign n10114 = ~n10108 & ~n39258;
  assign n10115 = n563 & n636;
  assign n10116 = pi85  & n37482;
  assign n10117 = pi87  & n578;
  assign n10118 = pi86  & n580;
  assign n10119 = ~n10117 & ~n10118;
  assign n10120 = ~n10116 & ~n10118;
  assign n10121 = ~n10117 & n10120;
  assign n10122 = ~n10116 & n10119;
  assign n10123 = ~n10115 & n39259;
  assign n10124 = pi14  & ~n10123;
  assign n10125 = pi14  & ~n10124;
  assign n10126 = pi14  & n10123;
  assign n10127 = ~n10123 & ~n10124;
  assign n10128 = ~pi14  & ~n10123;
  assign n10129 = ~n39260 & ~n39261;
  assign n10130 = n9108 & ~n9110;
  assign n10131 = ~n9108 & ~n39062;
  assign n10132 = ~n9109 & n9114;
  assign n10133 = ~n10131 & ~n10132;
  assign n10134 = ~n39062 & ~n10130;
  assign n10135 = ~n10129 & ~n39262;
  assign n10136 = n9099 & n39061;
  assign n10137 = ~n9107 & ~n10136;
  assign n10138 = n563 & n2779;
  assign n10139 = pi84  & n37482;
  assign n10140 = pi86  & n578;
  assign n10141 = pi85  & n580;
  assign n10142 = ~n10140 & ~n10141;
  assign n10143 = ~n10139 & ~n10141;
  assign n10144 = ~n10140 & n10143;
  assign n10145 = ~n10139 & n10142;
  assign n10146 = ~n10138 & n39263;
  assign n10147 = pi14  & ~n10146;
  assign n10148 = pi14  & ~n10147;
  assign n10149 = pi14  & n10146;
  assign n10150 = ~n10146 & ~n10147;
  assign n10151 = ~pi14  & ~n10146;
  assign n10152 = ~n39264 & ~n39265;
  assign n10153 = n10137 & ~n10152;
  assign n10154 = n9095 & ~n9097;
  assign n10155 = ~n9098 & ~n10154;
  assign n10156 = n563 & n2804;
  assign n10157 = pi83  & n37482;
  assign n10158 = pi85  & n578;
  assign n10159 = pi84  & n580;
  assign n10160 = ~n10158 & ~n10159;
  assign n10161 = ~n10157 & ~n10159;
  assign n10162 = ~n10158 & n10161;
  assign n10163 = ~n10157 & n10160;
  assign n10164 = ~n10156 & n39266;
  assign n10165 = pi14  & ~n10164;
  assign n10166 = pi14  & ~n10165;
  assign n10167 = pi14  & n10164;
  assign n10168 = ~n10164 & ~n10165;
  assign n10169 = ~pi14  & ~n10164;
  assign n10170 = ~n39267 & ~n39268;
  assign n10171 = n10155 & ~n10170;
  assign n10172 = n9086 & n39058;
  assign n10173 = ~n9094 & ~n10172;
  assign n10174 = n563 & n2591;
  assign n10175 = pi82  & n37482;
  assign n10176 = pi84  & n578;
  assign n10177 = pi83  & n580;
  assign n10178 = ~n10176 & ~n10177;
  assign n10179 = ~n10175 & ~n10177;
  assign n10180 = ~n10176 & n10179;
  assign n10181 = ~n10175 & n10178;
  assign n10182 = ~n10174 & n39269;
  assign n10183 = pi14  & ~n10182;
  assign n10184 = pi14  & ~n10183;
  assign n10185 = pi14  & n10182;
  assign n10186 = ~n10182 & ~n10183;
  assign n10187 = ~pi14  & ~n10182;
  assign n10188 = ~n39270 & ~n39271;
  assign n10189 = n10173 & ~n10188;
  assign n10190 = n9077 & n39055;
  assign n10191 = ~n9085 & ~n10190;
  assign n10192 = n563 & n2091;
  assign n10193 = pi81  & n37482;
  assign n10194 = pi83  & n578;
  assign n10195 = pi82  & n580;
  assign n10196 = ~n10194 & ~n10195;
  assign n10197 = ~n10193 & ~n10195;
  assign n10198 = ~n10194 & n10197;
  assign n10199 = ~n10193 & n10196;
  assign n10200 = ~n10192 & n39272;
  assign n10201 = pi14  & ~n10200;
  assign n10202 = pi14  & ~n10201;
  assign n10203 = pi14  & n10200;
  assign n10204 = ~n10200 & ~n10201;
  assign n10205 = ~pi14  & ~n10200;
  assign n10206 = ~n39273 & ~n39274;
  assign n10207 = n10191 & ~n10206;
  assign n10208 = n9068 & n39052;
  assign n10209 = ~n9076 & ~n10208;
  assign n10210 = n563 & n2134;
  assign n10211 = pi80  & n37482;
  assign n10212 = pi82  & n578;
  assign n10213 = pi81  & n580;
  assign n10214 = ~n10212 & ~n10213;
  assign n10215 = ~n10211 & ~n10213;
  assign n10216 = ~n10212 & n10215;
  assign n10217 = ~n10211 & n10214;
  assign n10218 = ~n10210 & n39275;
  assign n10219 = pi14  & ~n10218;
  assign n10220 = pi14  & ~n10219;
  assign n10221 = pi14  & n10218;
  assign n10222 = ~n10218 & ~n10219;
  assign n10223 = ~pi14  & ~n10218;
  assign n10224 = ~n39276 & ~n39277;
  assign n10225 = n10209 & ~n10224;
  assign n10226 = n9059 & n39049;
  assign n10227 = ~n9067 & ~n10226;
  assign n10228 = n563 & n2154;
  assign n10229 = pi79  & n37482;
  assign n10230 = pi81  & n578;
  assign n10231 = pi80  & n580;
  assign n10232 = ~n10230 & ~n10231;
  assign n10233 = ~n10229 & ~n10231;
  assign n10234 = ~n10230 & n10233;
  assign n10235 = ~n10229 & n10232;
  assign n10236 = ~n10228 & n39278;
  assign n10237 = pi14  & ~n10236;
  assign n10238 = pi14  & ~n10237;
  assign n10239 = pi14  & n10236;
  assign n10240 = ~n10236 & ~n10237;
  assign n10241 = ~pi14  & ~n10236;
  assign n10242 = ~n39279 & ~n39280;
  assign n10243 = n10227 & ~n10242;
  assign n10244 = n563 & n2063;
  assign n10245 = pi78  & n37482;
  assign n10246 = pi80  & n578;
  assign n10247 = pi79  & n580;
  assign n10248 = ~n10246 & ~n10247;
  assign n10249 = ~n10245 & ~n10247;
  assign n10250 = ~n10246 & n10249;
  assign n10251 = ~n10245 & n10248;
  assign n10252 = ~n10244 & n39281;
  assign n10253 = pi14  & ~n10252;
  assign n10254 = pi14  & ~n10253;
  assign n10255 = pi14  & n10252;
  assign n10256 = ~n10252 & ~n10253;
  assign n10257 = ~pi14  & ~n10252;
  assign n10258 = ~n39282 & ~n39283;
  assign n10259 = n9050 & n39046;
  assign n10260 = ~n39046 & ~n9058;
  assign n10261 = n9050 & ~n39046;
  assign n10262 = ~n9050 & ~n9058;
  assign n10263 = ~n9050 & n39046;
  assign n10264 = ~n39284 & ~n39285;
  assign n10265 = ~n9058 & ~n10259;
  assign n10266 = ~n10258 & ~n39286;
  assign n10267 = n9046 & ~n9048;
  assign n10268 = ~n9049 & ~n10267;
  assign n10269 = n563 & n678;
  assign n10270 = pi77  & n37482;
  assign n10271 = pi79  & n578;
  assign n10272 = pi78  & n580;
  assign n10273 = ~n10271 & ~n10272;
  assign n10274 = ~n10270 & ~n10272;
  assign n10275 = ~n10271 & n10274;
  assign n10276 = ~n10270 & n10273;
  assign n10277 = ~n10269 & n39287;
  assign n10278 = pi14  & ~n10277;
  assign n10279 = pi14  & ~n10278;
  assign n10280 = pi14  & n10277;
  assign n10281 = ~n10277 & ~n10278;
  assign n10282 = ~pi14  & ~n10277;
  assign n10283 = ~n39288 & ~n39289;
  assign n10284 = n10268 & ~n10283;
  assign n10285 = n9042 & ~n9044;
  assign n10286 = ~n9045 & ~n10285;
  assign n10287 = n563 & n1578;
  assign n10288 = pi76  & n37482;
  assign n10289 = pi78  & n578;
  assign n10290 = pi77  & n580;
  assign n10291 = ~n10289 & ~n10290;
  assign n10292 = ~n10288 & ~n10290;
  assign n10293 = ~n10289 & n10292;
  assign n10294 = ~n10288 & n10291;
  assign n10295 = ~n10287 & n39290;
  assign n10296 = pi14  & ~n10295;
  assign n10297 = pi14  & ~n10296;
  assign n10298 = pi14  & n10295;
  assign n10299 = ~n10295 & ~n10296;
  assign n10300 = ~pi14  & ~n10295;
  assign n10301 = ~n39291 & ~n39292;
  assign n10302 = n10286 & ~n10301;
  assign n10303 = n9033 & n39043;
  assign n10304 = ~n9041 & ~n10303;
  assign n10305 = n563 & n1596;
  assign n10306 = pi75  & n37482;
  assign n10307 = pi77  & n578;
  assign n10308 = pi76  & n580;
  assign n10309 = ~n10307 & ~n10308;
  assign n10310 = ~n10306 & ~n10308;
  assign n10311 = ~n10307 & n10310;
  assign n10312 = ~n10306 & n10309;
  assign n10313 = ~n10305 & n39293;
  assign n10314 = pi14  & ~n10313;
  assign n10315 = pi14  & ~n10314;
  assign n10316 = pi14  & n10313;
  assign n10317 = ~n10313 & ~n10314;
  assign n10318 = ~pi14  & ~n10313;
  assign n10319 = ~n39294 & ~n39295;
  assign n10320 = n10304 & ~n10319;
  assign n10321 = ~n10304 & n10319;
  assign n10322 = ~n10320 & ~n10321;
  assign n10323 = n563 & n1465;
  assign n10324 = pi74  & n37482;
  assign n10325 = pi76  & n578;
  assign n10326 = pi75  & n580;
  assign n10327 = ~n10325 & ~n10326;
  assign n10328 = ~n10324 & ~n10326;
  assign n10329 = ~n10325 & n10328;
  assign n10330 = ~n10324 & n10327;
  assign n10331 = ~n10323 & n39296;
  assign n10332 = pi14  & ~n10331;
  assign n10333 = pi14  & ~n10332;
  assign n10334 = pi14  & n10331;
  assign n10335 = ~n10331 & ~n10332;
  assign n10336 = ~pi14  & ~n10331;
  assign n10337 = ~n39297 & ~n39298;
  assign n10338 = n9029 & ~n9031;
  assign n10339 = ~n9032 & ~n10338;
  assign n10340 = ~n10337 & n10339;
  assign n10341 = n563 & n720;
  assign n10342 = pi73  & n37482;
  assign n10343 = pi75  & n578;
  assign n10344 = pi74  & n580;
  assign n10345 = ~n10343 & ~n10344;
  assign n10346 = ~n10342 & ~n10344;
  assign n10347 = ~n10343 & n10346;
  assign n10348 = ~n10342 & n10345;
  assign n10349 = ~n10341 & n39299;
  assign n10350 = pi14  & ~n10349;
  assign n10351 = pi14  & ~n10350;
  assign n10352 = pi14  & n10349;
  assign n10353 = ~n10349 & ~n10350;
  assign n10354 = ~pi14  & ~n10349;
  assign n10355 = ~n39300 & ~n39301;
  assign n10356 = n9025 & ~n9027;
  assign n10357 = ~n9028 & ~n10356;
  assign n10358 = ~n10355 & n10357;
  assign n10359 = n9021 & ~n9023;
  assign n10360 = ~n9024 & ~n10359;
  assign n10361 = n563 & n1218;
  assign n10362 = pi72  & n37482;
  assign n10363 = pi74  & n578;
  assign n10364 = pi73  & n580;
  assign n10365 = ~n10363 & ~n10364;
  assign n10366 = ~n10362 & ~n10364;
  assign n10367 = ~n10363 & n10366;
  assign n10368 = ~n10362 & n10365;
  assign n10369 = ~n10361 & n39302;
  assign n10370 = pi14  & ~n10369;
  assign n10371 = pi14  & ~n10370;
  assign n10372 = pi14  & n10369;
  assign n10373 = ~n10369 & ~n10370;
  assign n10374 = ~pi14  & ~n10369;
  assign n10375 = ~n39303 & ~n39304;
  assign n10376 = n10360 & ~n10375;
  assign n10377 = n563 & n1238;
  assign n10378 = pi71  & n37482;
  assign n10379 = pi73  & n578;
  assign n10380 = pi72  & n580;
  assign n10381 = ~n10379 & ~n10380;
  assign n10382 = ~n10378 & ~n10380;
  assign n10383 = ~n10379 & n10382;
  assign n10384 = ~n10378 & n10381;
  assign n10385 = ~n10377 & n39305;
  assign n10386 = pi14  & ~n10385;
  assign n10387 = pi14  & ~n10386;
  assign n10388 = pi14  & n10385;
  assign n10389 = ~n10385 & ~n10386;
  assign n10390 = ~pi14  & ~n10385;
  assign n10391 = ~n39306 & ~n39307;
  assign n10392 = n9012 & n39040;
  assign n10393 = ~n9012 & n39040;
  assign n10394 = n9012 & ~n39040;
  assign n10395 = ~n10393 & ~n10394;
  assign n10396 = ~n9020 & ~n10392;
  assign n10397 = ~n10391 & ~n39308;
  assign n10398 = n563 & n1124;
  assign n10399 = pi70  & n37482;
  assign n10400 = pi72  & n578;
  assign n10401 = pi71  & n580;
  assign n10402 = ~n10400 & ~n10401;
  assign n10403 = ~n10399 & ~n10401;
  assign n10404 = ~n10400 & n10403;
  assign n10405 = ~n10399 & n10402;
  assign n10406 = ~n10398 & n39309;
  assign n10407 = pi14  & ~n10406;
  assign n10408 = pi14  & ~n10407;
  assign n10409 = pi14  & n10406;
  assign n10410 = ~n10406 & ~n10407;
  assign n10411 = ~pi14  & ~n10406;
  assign n10412 = ~n39310 & ~n39311;
  assign n10413 = n9006 & ~n9008;
  assign n10414 = ~n9006 & ~n39037;
  assign n10415 = ~n9007 & n9012;
  assign n10416 = ~n10414 & ~n10415;
  assign n10417 = ~n39037 & ~n10413;
  assign n10418 = ~n10412 & ~n39312;
  assign n10419 = n563 & n927;
  assign n10420 = pi69  & n37482;
  assign n10421 = pi71  & n578;
  assign n10422 = pi70  & n580;
  assign n10423 = ~n10421 & ~n10422;
  assign n10424 = ~n10420 & ~n10422;
  assign n10425 = ~n10421 & n10424;
  assign n10426 = ~n10420 & n10423;
  assign n10427 = ~n10419 & n39313;
  assign n10428 = pi14  & ~n10427;
  assign n10429 = pi14  & ~n10428;
  assign n10430 = pi14  & n10427;
  assign n10431 = ~n10427 & ~n10428;
  assign n10432 = ~pi14  & ~n10427;
  assign n10433 = ~n39314 & ~n39315;
  assign n10434 = n8999 & n39036;
  assign n10435 = ~n9005 & ~n10434;
  assign n10436 = ~n10433 & n10435;
  assign n10437 = n8992 & n39035;
  assign n10438 = ~n8998 & ~n10437;
  assign n10439 = n563 & n972;
  assign n10440 = pi68  & n37482;
  assign n10441 = pi70  & n578;
  assign n10442 = pi69  & n580;
  assign n10443 = ~n10441 & ~n10442;
  assign n10444 = ~n10440 & ~n10442;
  assign n10445 = ~n10441 & n10444;
  assign n10446 = ~n10440 & n10443;
  assign n10447 = ~n10439 & n39316;
  assign n10448 = pi14  & ~n10447;
  assign n10449 = pi14  & ~n10448;
  assign n10450 = pi14  & n10447;
  assign n10451 = ~n10447 & ~n10448;
  assign n10452 = ~pi14  & ~n10447;
  assign n10453 = ~n39317 & ~n39318;
  assign n10454 = n10438 & ~n10453;
  assign n10455 = n563 & n990;
  assign n10456 = pi67  & n37482;
  assign n10457 = pi69  & n578;
  assign n10458 = pi68  & n580;
  assign n10459 = ~n10457 & ~n10458;
  assign n10460 = ~n10456 & ~n10458;
  assign n10461 = ~n10457 & n10460;
  assign n10462 = ~n10456 & n10459;
  assign n10463 = ~n10455 & n39319;
  assign n10464 = pi14  & ~n10463;
  assign n10465 = pi14  & ~n10464;
  assign n10466 = pi14  & n10463;
  assign n10467 = ~n10463 & ~n10464;
  assign n10468 = ~pi14  & ~n10463;
  assign n10469 = ~n39320 & ~n39321;
  assign n10470 = pi17  & ~n39027;
  assign n10471 = n39030 & ~n10470;
  assign n10472 = ~n39030 & n10470;
  assign n10473 = ~n39027 & n8974;
  assign n10474 = ~n39031 & ~n10473;
  assign n10475 = ~n10471 & ~n10472;
  assign n10476 = ~n10469 & n39322;
  assign n10477 = n563 & n871;
  assign n10478 = pi66  & n37482;
  assign n10479 = pi68  & n578;
  assign n10480 = pi67  & n580;
  assign n10481 = ~n10479 & ~n10480;
  assign n10482 = ~n10478 & ~n10480;
  assign n10483 = ~n10479 & n10482;
  assign n10484 = ~n10478 & n10481;
  assign n10485 = ~n10477 & n39323;
  assign n10486 = pi14  & ~n10485;
  assign n10487 = pi14  & ~n10486;
  assign n10488 = pi14  & n10485;
  assign n10489 = ~n10485 & ~n10486;
  assign n10490 = ~pi14  & ~n10485;
  assign n10491 = ~n39324 & ~n39325;
  assign n10492 = pi17  & n8948;
  assign n10493 = ~n8947 & n10492;
  assign n10494 = n8947 & ~n10492;
  assign n10495 = ~n8949 & n8953;
  assign n10496 = ~n39027 & ~n10495;
  assign n10497 = ~n10493 & ~n10494;
  assign n10498 = ~n10491 & n39326;
  assign n10499 = n563 & n37515;
  assign n10500 = pi65  & n578;
  assign n10501 = pi64  & n580;
  assign n10502 = ~n10500 & ~n10501;
  assign n10503 = ~n10499 & n10502;
  assign n10504 = pi64  & n37479;
  assign n10505 = pi14  & ~n10504;
  assign n10506 = pi14  & ~n10503;
  assign n10507 = pi14  & ~n10506;
  assign n10508 = ~n10503 & ~n10506;
  assign n10509 = ~n10507 & ~n10508;
  assign n10510 = n10505 & ~n10509;
  assign n10511 = n10503 & n10505;
  assign n10512 = pi64  & n37482;
  assign n10513 = pi65  & n580;
  assign n10514 = n563 & ~n37521;
  assign n10515 = pi66  & n578;
  assign n10516 = ~n10514 & ~n10515;
  assign n10517 = ~n10513 & ~n10514;
  assign n10518 = ~n10515 & n10517;
  assign n10519 = ~n10513 & ~n10515;
  assign n10520 = ~n10514 & n10519;
  assign n10521 = ~n10513 & n10516;
  assign n10522 = ~n10512 & ~n10513;
  assign n10523 = ~n10515 & n10522;
  assign n10524 = ~n10512 & n10519;
  assign n10525 = ~n10514 & n39329;
  assign n10526 = ~n10512 & n39328;
  assign n10527 = pi14  & ~n39330;
  assign n10528 = pi14  & ~n10527;
  assign n10529 = ~n39330 & ~n10527;
  assign n10530 = ~n10528 & ~n10529;
  assign n10531 = n39327 & ~n10530;
  assign n10532 = n39327 & n39330;
  assign n10533 = n8948 & n39331;
  assign n10534 = n563 & n847;
  assign n10535 = pi65  & n37482;
  assign n10536 = pi67  & n578;
  assign n10537 = pi66  & n580;
  assign n10538 = ~n10536 & ~n10537;
  assign n10539 = ~n10535 & ~n10537;
  assign n10540 = ~n10536 & n10539;
  assign n10541 = ~n10535 & n10538;
  assign n10542 = ~n10534 & n39332;
  assign n10543 = pi14  & ~n10542;
  assign n10544 = pi14  & ~n10543;
  assign n10545 = pi14  & n10542;
  assign n10546 = ~n10542 & ~n10543;
  assign n10547 = ~pi14  & ~n10542;
  assign n10548 = ~n39333 & ~n39334;
  assign n10549 = ~n8948 & ~n39331;
  assign n10550 = n8948 & ~n39331;
  assign n10551 = ~n8948 & n39331;
  assign n10552 = ~n10550 & ~n10551;
  assign n10553 = ~n10533 & ~n10549;
  assign n10554 = ~n10548 & ~n39335;
  assign n10555 = ~n10533 & ~n10554;
  assign n10556 = n10491 & ~n39326;
  assign n10557 = ~n10498 & ~n10556;
  assign n10558 = ~n10555 & n10557;
  assign n10559 = ~n10498 & ~n10558;
  assign n10560 = n10469 & ~n39322;
  assign n10561 = ~n10476 & ~n10560;
  assign n10562 = ~n10559 & ~n10560;
  assign n10563 = ~n10476 & n10562;
  assign n10564 = ~n10559 & n10561;
  assign n10565 = ~n10476 & ~n39336;
  assign n10566 = ~n10438 & n10453;
  assign n10567 = n10438 & ~n10454;
  assign n10568 = n10438 & n10453;
  assign n10569 = ~n10453 & ~n10454;
  assign n10570 = ~n10438 & ~n10453;
  assign n10571 = ~n39337 & ~n39338;
  assign n10572 = ~n10454 & ~n10566;
  assign n10573 = ~n10565 & ~n39339;
  assign n10574 = ~n10454 & ~n10573;
  assign n10575 = n10433 & ~n10435;
  assign n10576 = ~n10436 & ~n10575;
  assign n10577 = ~n10574 & n10576;
  assign n10578 = ~n10436 & ~n10577;
  assign n10579 = n10412 & n39312;
  assign n10580 = ~n10418 & ~n10579;
  assign n10581 = ~n10578 & n10580;
  assign n10582 = ~n10418 & ~n10581;
  assign n10583 = n10391 & n39308;
  assign n10584 = ~n10397 & ~n10583;
  assign n10585 = ~n10582 & n10584;
  assign n10586 = ~n10397 & ~n10585;
  assign n10587 = ~n10360 & n10375;
  assign n10588 = n10360 & ~n10376;
  assign n10589 = n10360 & n10375;
  assign n10590 = ~n10375 & ~n10376;
  assign n10591 = ~n10360 & ~n10375;
  assign n10592 = ~n39340 & ~n39341;
  assign n10593 = ~n10376 & ~n10587;
  assign n10594 = ~n10586 & ~n39342;
  assign n10595 = ~n10376 & ~n10594;
  assign n10596 = n10355 & ~n10357;
  assign n10597 = ~n10358 & ~n10596;
  assign n10598 = ~n10595 & n10597;
  assign n10599 = ~n10358 & ~n10598;
  assign n10600 = n10337 & ~n10339;
  assign n10601 = ~n10340 & ~n10600;
  assign n10602 = ~n10599 & n10601;
  assign n10603 = ~n10340 & ~n10602;
  assign n10604 = n10322 & ~n10603;
  assign n10605 = ~n10320 & ~n10604;
  assign n10606 = ~n10286 & n10301;
  assign n10607 = n10286 & ~n10302;
  assign n10608 = n10286 & n10301;
  assign n10609 = ~n10301 & ~n10302;
  assign n10610 = ~n10286 & ~n10301;
  assign n10611 = ~n39343 & ~n39344;
  assign n10612 = ~n10302 & ~n10606;
  assign n10613 = ~n10605 & ~n39345;
  assign n10614 = ~n10302 & ~n10613;
  assign n10615 = ~n10268 & n10283;
  assign n10616 = n10268 & ~n10284;
  assign n10617 = n10268 & n10283;
  assign n10618 = ~n10283 & ~n10284;
  assign n10619 = ~n10268 & ~n10283;
  assign n10620 = ~n39346 & ~n39347;
  assign n10621 = ~n10284 & ~n10615;
  assign n10622 = ~n10614 & ~n39348;
  assign n10623 = ~n10284 & ~n10622;
  assign n10624 = n10258 & n39286;
  assign n10625 = ~n39286 & ~n10266;
  assign n10626 = ~n10258 & ~n10266;
  assign n10627 = ~n10625 & ~n10626;
  assign n10628 = ~n10266 & ~n10624;
  assign n10629 = ~n10623 & ~n39349;
  assign n10630 = ~n10266 & ~n10629;
  assign n10631 = ~n10227 & n10242;
  assign n10632 = n10227 & ~n10243;
  assign n10633 = n10227 & n10242;
  assign n10634 = ~n10242 & ~n10243;
  assign n10635 = ~n10227 & ~n10242;
  assign n10636 = ~n39350 & ~n39351;
  assign n10637 = ~n10243 & ~n10631;
  assign n10638 = ~n10630 & ~n39352;
  assign n10639 = ~n10243 & ~n10638;
  assign n10640 = ~n10209 & n10224;
  assign n10641 = n10209 & ~n10225;
  assign n10642 = n10209 & n10224;
  assign n10643 = ~n10224 & ~n10225;
  assign n10644 = ~n10209 & ~n10224;
  assign n10645 = ~n39353 & ~n39354;
  assign n10646 = ~n10225 & ~n10640;
  assign n10647 = ~n10639 & ~n39355;
  assign n10648 = ~n10225 & ~n10647;
  assign n10649 = ~n10191 & n10206;
  assign n10650 = n10191 & ~n10207;
  assign n10651 = n10191 & n10206;
  assign n10652 = ~n10206 & ~n10207;
  assign n10653 = ~n10191 & ~n10206;
  assign n10654 = ~n39356 & ~n39357;
  assign n10655 = ~n10207 & ~n10649;
  assign n10656 = ~n10648 & ~n39358;
  assign n10657 = ~n10207 & ~n10656;
  assign n10658 = ~n10173 & n10188;
  assign n10659 = ~n10189 & ~n10658;
  assign n10660 = ~n10657 & ~n10658;
  assign n10661 = ~n10189 & n10660;
  assign n10662 = ~n10657 & n10659;
  assign n10663 = ~n10189 & ~n39359;
  assign n10664 = ~n10155 & n10170;
  assign n10665 = n10155 & ~n10171;
  assign n10666 = n10155 & n10170;
  assign n10667 = ~n10170 & ~n10171;
  assign n10668 = ~n10155 & ~n10170;
  assign n10669 = ~n39360 & ~n39361;
  assign n10670 = ~n10171 & ~n10664;
  assign n10671 = ~n10663 & ~n39362;
  assign n10672 = ~n10171 & ~n10671;
  assign n10673 = ~n10137 & n10152;
  assign n10674 = n10137 & ~n10153;
  assign n10675 = n10137 & n10152;
  assign n10676 = ~n10152 & ~n10153;
  assign n10677 = ~n10137 & ~n10152;
  assign n10678 = ~n39363 & ~n39364;
  assign n10679 = ~n10153 & ~n10673;
  assign n10680 = ~n10672 & ~n39365;
  assign n10681 = ~n10153 & ~n10680;
  assign n10682 = n10129 & n39262;
  assign n10683 = ~n10135 & ~n10682;
  assign n10684 = ~n10681 & n10683;
  assign n10685 = ~n10135 & ~n10684;
  assign n10686 = n10108 & n39258;
  assign n10687 = ~n10114 & ~n10686;
  assign n10688 = ~n10685 & n10687;
  assign n10689 = ~n10114 & ~n10688;
  assign n10690 = ~n10077 & n10092;
  assign n10691 = ~n10093 & ~n10690;
  assign n10692 = ~n10689 & ~n10690;
  assign n10693 = ~n10093 & n10692;
  assign n10694 = ~n10689 & n10691;
  assign n10695 = ~n10093 & ~n39366;
  assign n10696 = n10069 & n39251;
  assign n10697 = ~n10075 & ~n10696;
  assign n10698 = ~n10695 & n10697;
  assign n10699 = ~n10075 & ~n10698;
  assign n10700 = ~n10038 & n10053;
  assign n10701 = n10038 & ~n10054;
  assign n10702 = n10038 & n10053;
  assign n10703 = ~n10053 & ~n10054;
  assign n10704 = ~n10038 & ~n10053;
  assign n10705 = ~n39367 & ~n39368;
  assign n10706 = ~n10054 & ~n10700;
  assign n10707 = ~n10699 & ~n39369;
  assign n10708 = ~n10054 & ~n10707;
  assign n10709 = n10033 & ~n10035;
  assign n10710 = ~n10033 & ~n10036;
  assign n10711 = ~n10033 & ~n10035;
  assign n10712 = n10035 & ~n10036;
  assign n10713 = n10033 & n10035;
  assign n10714 = ~n39370 & ~n39371;
  assign n10715 = ~n10036 & ~n10709;
  assign n10716 = ~n10708 & ~n39372;
  assign n10717 = ~n10036 & ~n10716;
  assign n10718 = n10015 & ~n10017;
  assign n10719 = ~n10018 & ~n10718;
  assign n10720 = ~n10717 & n10719;
  assign n10721 = ~n10018 & ~n10720;
  assign n10722 = n9994 & n39238;
  assign n10723 = ~n10000 & ~n10722;
  assign n10724 = ~n10721 & n10723;
  assign n10725 = ~n10000 & ~n10724;
  assign n10726 = n9971 & n39234;
  assign n10727 = ~n9979 & ~n10726;
  assign n10728 = ~n10725 & n10727;
  assign n10729 = ~n9979 & ~n10728;
  assign n10730 = n9953 & ~n9955;
  assign n10731 = ~n9956 & ~n10730;
  assign n10732 = ~n10729 & n10731;
  assign n10733 = ~n9956 & ~n10732;
  assign n10734 = ~n9922 & n9937;
  assign n10735 = n9922 & ~n9938;
  assign n10736 = n9922 & n9937;
  assign n10737 = ~n9937 & ~n9938;
  assign n10738 = ~n9922 & ~n9937;
  assign n10739 = ~n39373 & ~n39374;
  assign n10740 = ~n9938 & ~n10734;
  assign n10741 = ~n10733 & ~n39375;
  assign n10742 = ~n9938 & ~n10741;
  assign n10743 = ~n9904 & n9919;
  assign n10744 = n9904 & ~n9920;
  assign n10745 = n9904 & n9919;
  assign n10746 = ~n9919 & ~n9920;
  assign n10747 = ~n9904 & ~n9919;
  assign n10748 = ~n39376 & ~n39377;
  assign n10749 = ~n9920 & ~n10743;
  assign n10750 = ~n10742 & ~n39378;
  assign n10751 = ~n9920 & ~n10750;
  assign n10752 = ~n9886 & n9901;
  assign n10753 = n9886 & ~n9902;
  assign n10754 = n9886 & n9901;
  assign n10755 = ~n9901 & ~n9902;
  assign n10756 = ~n9886 & ~n9901;
  assign n10757 = ~n39379 & ~n39380;
  assign n10758 = ~n9902 & ~n10752;
  assign n10759 = ~n10751 & ~n39381;
  assign n10760 = ~n9902 & ~n10759;
  assign n10761 = n9878 & n39216;
  assign n10762 = ~n9884 & ~n10761;
  assign n10763 = ~n10760 & n10762;
  assign n10764 = ~n9884 & ~n10763;
  assign n10765 = ~n9847 & n9862;
  assign n10766 = n9847 & ~n9863;
  assign n10767 = n9847 & n9862;
  assign n10768 = ~n9862 & ~n9863;
  assign n10769 = ~n9847 & ~n9862;
  assign n10770 = ~n39382 & ~n39383;
  assign n10771 = ~n9863 & ~n10765;
  assign n10772 = ~n10764 & ~n39384;
  assign n10773 = ~n9863 & ~n10772;
  assign n10774 = ~n9829 & n9844;
  assign n10775 = n9829 & ~n9845;
  assign n10776 = n9829 & n9844;
  assign n10777 = ~n9844 & ~n9845;
  assign n10778 = ~n9829 & ~n9844;
  assign n10779 = ~n39385 & ~n39386;
  assign n10780 = ~n9845 & ~n10774;
  assign n10781 = ~n10773 & ~n39387;
  assign n10782 = ~n9845 & ~n10781;
  assign n10783 = ~n9811 & n9826;
  assign n10784 = n9811 & ~n9827;
  assign n10785 = n9811 & n9826;
  assign n10786 = ~n9826 & ~n9827;
  assign n10787 = ~n9811 & ~n9826;
  assign n10788 = ~n39388 & ~n39389;
  assign n10789 = ~n9827 & ~n10783;
  assign n10790 = ~n10782 & ~n39390;
  assign n10791 = ~n9827 & ~n10790;
  assign n10792 = ~n9793 & n9808;
  assign n10793 = n9793 & ~n9809;
  assign n10794 = n9793 & n9808;
  assign n10795 = ~n9808 & ~n9809;
  assign n10796 = ~n9793 & ~n9808;
  assign n10797 = ~n39391 & ~n39392;
  assign n10798 = ~n9809 & ~n10792;
  assign n10799 = ~n10791 & ~n39393;
  assign n10800 = ~n9809 & ~n10799;
  assign n10801 = ~n9775 & n9790;
  assign n10802 = n9775 & ~n9791;
  assign n10803 = n9775 & n9790;
  assign n10804 = ~n9790 & ~n9791;
  assign n10805 = ~n9775 & ~n9790;
  assign n10806 = ~n39394 & ~n39395;
  assign n10807 = ~n9791 & ~n10801;
  assign n10808 = ~n10800 & ~n39396;
  assign n10809 = ~n9791 & ~n10808;
  assign n10810 = ~n9757 & n9772;
  assign n10811 = ~n9773 & ~n10810;
  assign n10812 = ~n10809 & n10811;
  assign n10813 = ~n9773 & ~n10812;
  assign n10814 = ~n9739 & n9754;
  assign n10815 = ~n9755 & ~n10814;
  assign n10816 = ~n10813 & ~n10814;
  assign n10817 = ~n9755 & n10816;
  assign n10818 = ~n10813 & n10815;
  assign n10819 = ~n9755 & ~n39397;
  assign n10820 = ~n9721 & n9736;
  assign n10821 = ~n9737 & ~n10820;
  assign n10822 = ~n10819 & ~n10820;
  assign n10823 = ~n9737 & n10822;
  assign n10824 = ~n10819 & n10821;
  assign n10825 = ~n9737 & ~n39398;
  assign n10826 = n9716 & ~n9718;
  assign n10827 = ~n9716 & ~n9719;
  assign n10828 = ~n9716 & ~n9718;
  assign n10829 = n9718 & ~n9719;
  assign n10830 = n9716 & n9718;
  assign n10831 = ~n39399 & ~n39400;
  assign n10832 = ~n9719 & ~n10826;
  assign n10833 = ~n10825 & ~n39401;
  assign n10834 = ~n9719 & ~n10833;
  assign n10835 = n9693 & n39185;
  assign n10836 = ~n9699 & ~n10835;
  assign n10837 = ~n10834 & n10836;
  assign n10838 = ~n9699 & ~n10837;
  assign n10839 = n592 & n39181;
  assign n10840 = ~n9676 & ~n10839;
  assign n10841 = ~n10838 & n10840;
  assign n10842 = ~n9676 & ~n10841;
  assign n10843 = n505 & ~n507;
  assign n10844 = ~n508 & ~n10843;
  assign n10845 = n563 & n10844;
  assign n10846 = pi110  & n37482;
  assign n10847 = pi112  & n578;
  assign n10848 = pi111  & n580;
  assign n10849 = ~n10847 & ~n10848;
  assign n10850 = ~n10846 & ~n10848;
  assign n10851 = ~n10847 & n10850;
  assign n10852 = ~n10846 & n10849;
  assign n10853 = ~n10845 & n39402;
  assign n10854 = pi14  & ~n10853;
  assign n10855 = pi14  & ~n10854;
  assign n10856 = pi14  & n10853;
  assign n10857 = ~n10853 & ~n10854;
  assign n10858 = ~pi14  & ~n10853;
  assign n10859 = ~n39403 & ~n39404;
  assign n10860 = ~n9662 & ~n9670;
  assign n10861 = n8175 & n9701;
  assign n10862 = pi107  & n38895;
  assign n10863 = pi109  & n8190;
  assign n10864 = pi108  & n8192;
  assign n10865 = ~n10863 & ~n10864;
  assign n10866 = ~n10862 & ~n10864;
  assign n10867 = ~n10863 & n10866;
  assign n10868 = ~n10862 & n10865;
  assign n10869 = ~n10861 & n39405;
  assign n10870 = pi17  & ~n10869;
  assign n10871 = pi17  & ~n10870;
  assign n10872 = pi17  & n10869;
  assign n10873 = ~n10869 & ~n10870;
  assign n10874 = ~pi17  & ~n10869;
  assign n10875 = ~n39406 & ~n39407;
  assign n10876 = ~n9624 & ~n9633;
  assign n10877 = ~n9598 & ~n9607;
  assign n10878 = n4492 & n6474;
  assign n10879 = pi98  & n38208;
  assign n10880 = pi100  & n4507;
  assign n10881 = pi99  & n4509;
  assign n10882 = ~n10880 & ~n10881;
  assign n10883 = ~n10879 & ~n10881;
  assign n10884 = ~n10880 & n10883;
  assign n10885 = ~n10879 & n10882;
  assign n10886 = ~n10878 & n39408;
  assign n10887 = pi26  & ~n10886;
  assign n10888 = pi26  & ~n10887;
  assign n10889 = pi26  & n10886;
  assign n10890 = ~n10886 & ~n10887;
  assign n10891 = ~pi26  & ~n10886;
  assign n10892 = ~n39409 & ~n39410;
  assign n10893 = ~n9578 & ~n9580;
  assign n10894 = ~n9539 & ~n9548;
  assign n10895 = ~n9518 & ~n9522;
  assign n10896 = ~n9506 & ~n9512;
  assign n10897 = n733 & n2804;
  assign n10898 = pi83  & n37510;
  assign n10899 = pi85  & n746;
  assign n10900 = pi84  & n748;
  assign n10901 = ~n10899 & ~n10900;
  assign n10902 = ~n10898 & ~n10900;
  assign n10903 = ~n10899 & n10902;
  assign n10904 = ~n10898 & n10901;
  assign n10905 = ~n10897 & n39411;
  assign n10906 = pi41  & ~n10905;
  assign n10907 = pi41  & ~n10906;
  assign n10908 = pi41  & n10905;
  assign n10909 = ~n10905 & ~n10906;
  assign n10910 = ~pi41  & ~n10905;
  assign n10911 = ~n39412 & ~n39413;
  assign n10912 = ~n9490 & ~n9498;
  assign n10913 = n940 & n2134;
  assign n10914 = pi80  & n37541;
  assign n10915 = pi82  & n953;
  assign n10916 = pi81  & n955;
  assign n10917 = ~n10915 & ~n10916;
  assign n10918 = ~n10914 & ~n10916;
  assign n10919 = ~n10915 & n10918;
  assign n10920 = ~n10914 & n10917;
  assign n10921 = ~n10913 & n39414;
  assign n10922 = pi44  & ~n10921;
  assign n10923 = pi44  & ~n10922;
  assign n10924 = pi44  & n10921;
  assign n10925 = ~n10921 & ~n10922;
  assign n10926 = ~pi44  & ~n10921;
  assign n10927 = ~n39415 & ~n39416;
  assign n10928 = ~n9479 & ~n9487;
  assign n10929 = n678 & n785;
  assign n10930 = pi77  & n37520;
  assign n10931 = pi79  & n787;
  assign n10932 = pi78  & n795;
  assign n10933 = ~n10931 & ~n10932;
  assign n10934 = ~n10930 & ~n10932;
  assign n10935 = ~n10931 & n10934;
  assign n10936 = ~n10930 & n10933;
  assign n10937 = ~n10929 & n39417;
  assign n10938 = pi47  & ~n10937;
  assign n10939 = pi47  & ~n10938;
  assign n10940 = pi47  & n10937;
  assign n10941 = ~n10937 & ~n10938;
  assign n10942 = ~pi47  & ~n10937;
  assign n10943 = ~n39418 & ~n39419;
  assign n10944 = ~n9459 & ~n9461;
  assign n10945 = n894 & n1465;
  assign n10946 = pi74  & n37580;
  assign n10947 = pi76  & n896;
  assign n10948 = pi75  & n904;
  assign n10949 = ~n10947 & ~n10948;
  assign n10950 = ~n10946 & ~n10948;
  assign n10951 = ~n10947 & n10950;
  assign n10952 = ~n10946 & n10949;
  assign n10953 = ~n10945 & n39420;
  assign n10954 = pi50  & ~n10953;
  assign n10955 = pi50  & ~n10954;
  assign n10956 = pi50  & n10953;
  assign n10957 = ~n10953 & ~n10954;
  assign n10958 = ~pi50  & ~n10953;
  assign n10959 = ~n39421 & ~n39422;
  assign n10960 = ~n9453 & ~n9455;
  assign n10961 = n1238 & n1971;
  assign n10962 = pi71  & n37864;
  assign n10963 = pi73  & n1973;
  assign n10964 = pi72  & n1981;
  assign n10965 = ~n10963 & ~n10964;
  assign n10966 = ~n10962 & ~n10964;
  assign n10967 = ~n10963 & n10966;
  assign n10968 = ~n10962 & n10965;
  assign n10969 = ~n10961 & n39423;
  assign n10970 = pi53  & ~n10969;
  assign n10971 = pi53  & ~n10970;
  assign n10972 = pi53  & n10969;
  assign n10973 = ~n10969 & ~n10970;
  assign n10974 = ~pi53  & ~n10969;
  assign n10975 = ~n39424 & ~n39425;
  assign n10976 = n847 & n7882;
  assign n10977 = pi65  & n39128;
  assign n10978 = pi67  & n7884;
  assign n10979 = pi66  & n7892;
  assign n10980 = ~n10978 & ~n10979;
  assign n10981 = ~n10977 & ~n10979;
  assign n10982 = ~n10978 & n10981;
  assign n10983 = ~n10977 & n10980;
  assign n10984 = ~n10976 & n39426;
  assign n10985 = pi59  & ~n10984;
  assign n10986 = pi59  & ~n10985;
  assign n10987 = pi59  & n10984;
  assign n10988 = ~n10984 & ~n10985;
  assign n10989 = ~pi59  & ~n10984;
  assign n10990 = ~n39427 & ~n39428;
  assign n10991 = pi59  & ~pi60 ;
  assign n10992 = ~pi59  & pi60 ;
  assign n10993 = ~pi59  & ~pi60 ;
  assign n10994 = pi59  & pi60 ;
  assign n10995 = ~n10993 & ~n10994;
  assign n10996 = ~n10991 & ~n10992;
  assign n10997 = pi64  & n39429;
  assign n10998 = n39132 & n10997;
  assign n10999 = ~n39132 & ~n10997;
  assign n11000 = ~n39132 & n10997;
  assign n11001 = n39132 & ~n10997;
  assign n11002 = ~n11000 & ~n11001;
  assign n11003 = ~n10998 & ~n10999;
  assign n11004 = ~n10990 & ~n39430;
  assign n11005 = n10990 & n39430;
  assign n11006 = ~n11004 & ~n11005;
  assign n11007 = n972 & n4312;
  assign n11008 = pi68  & n38376;
  assign n11009 = pi70  & n4314;
  assign n11010 = pi69  & n4322;
  assign n11011 = ~n11009 & ~n11010;
  assign n11012 = ~n11008 & ~n11010;
  assign n11013 = ~n11009 & n11012;
  assign n11014 = ~n11008 & n11011;
  assign n11015 = ~n11007 & n39431;
  assign n11016 = pi56  & ~n11015;
  assign n11017 = pi56  & ~n11016;
  assign n11018 = pi56  & n11015;
  assign n11019 = ~n11015 & ~n11016;
  assign n11020 = ~pi56  & ~n11015;
  assign n11021 = ~n39432 & ~n39433;
  assign n11022 = n11006 & ~n11021;
  assign n11023 = ~n11006 & n11021;
  assign n11024 = n11006 & ~n11022;
  assign n11025 = n11006 & n11021;
  assign n11026 = ~n11021 & ~n11022;
  assign n11027 = ~n11006 & ~n11021;
  assign n11028 = ~n39434 & ~n39435;
  assign n11029 = ~n11022 & ~n11023;
  assign n11030 = ~n9448 & ~n39436;
  assign n11031 = n9448 & n39436;
  assign n11032 = ~n9448 & n39436;
  assign n11033 = n9448 & ~n39436;
  assign n11034 = ~n11032 & ~n11033;
  assign n11035 = ~n11030 & ~n11031;
  assign n11036 = ~n10975 & ~n39437;
  assign n11037 = n10975 & n39437;
  assign n11038 = ~n11036 & ~n11037;
  assign n11039 = ~n10960 & n11038;
  assign n11040 = n10960 & ~n11038;
  assign n11041 = ~n11039 & ~n11040;
  assign n11042 = n10959 & ~n11041;
  assign n11043 = ~n10959 & n11041;
  assign n11044 = ~n11042 & ~n11043;
  assign n11045 = ~n10944 & n11044;
  assign n11046 = n10944 & ~n11044;
  assign n11047 = ~n11045 & ~n11046;
  assign n11048 = ~n10943 & n11047;
  assign n11049 = n10943 & ~n11047;
  assign n11050 = ~n11048 & ~n11049;
  assign n11051 = ~n10928 & n11050;
  assign n11052 = n10928 & ~n11050;
  assign n11053 = ~n11051 & ~n11052;
  assign n11054 = ~n10927 & n11053;
  assign n11055 = n10927 & ~n11053;
  assign n11056 = ~n10927 & ~n11054;
  assign n11057 = ~n10927 & ~n11053;
  assign n11058 = n11053 & ~n11054;
  assign n11059 = n10927 & n11053;
  assign n11060 = ~n39438 & ~n39439;
  assign n11061 = ~n11054 & ~n11055;
  assign n11062 = ~n10912 & ~n39440;
  assign n11063 = n10912 & ~n39439;
  assign n11064 = ~n39438 & n11063;
  assign n11065 = n10912 & n39440;
  assign n11066 = ~n11062 & ~n39441;
  assign n11067 = ~n10911 & n11066;
  assign n11068 = n10911 & ~n11066;
  assign n11069 = ~n11067 & ~n11068;
  assign n11070 = ~n10896 & n11069;
  assign n11071 = n10896 & ~n11069;
  assign n11072 = ~n11070 & ~n11071;
  assign n11073 = n691 & n3354;
  assign n11074 = pi86  & n37503;
  assign n11075 = pi88  & n704;
  assign n11076 = pi87  & n706;
  assign n11077 = ~n11075 & ~n11076;
  assign n11078 = ~n11074 & ~n11076;
  assign n11079 = ~n11075 & n11078;
  assign n11080 = ~n11074 & n11077;
  assign n11081 = ~n11073 & n39442;
  assign n11082 = pi38  & ~n11081;
  assign n11083 = pi38  & ~n11082;
  assign n11084 = pi38  & n11081;
  assign n11085 = ~n11081 & ~n11082;
  assign n11086 = ~pi38  & ~n11081;
  assign n11087 = ~n39443 & ~n39444;
  assign n11088 = n11072 & ~n11087;
  assign n11089 = ~n11072 & n11087;
  assign n11090 = n11072 & ~n11088;
  assign n11091 = n11072 & n11087;
  assign n11092 = ~n11087 & ~n11088;
  assign n11093 = ~n11072 & ~n11087;
  assign n11094 = ~n39445 & ~n39446;
  assign n11095 = ~n11088 & ~n11089;
  assign n11096 = n10895 & n39447;
  assign n11097 = ~n10895 & ~n39447;
  assign n11098 = ~n11096 & ~n11097;
  assign n11099 = n594 & n2104;
  assign n11100 = pi89  & n37758;
  assign n11101 = pi91  & n2117;
  assign n11102 = pi90  & n2119;
  assign n11103 = ~n11101 & ~n11102;
  assign n11104 = ~n11100 & ~n11102;
  assign n11105 = ~n11101 & n11104;
  assign n11106 = ~n11100 & n11103;
  assign n11107 = ~n11099 & n39448;
  assign n11108 = pi35  & ~n11107;
  assign n11109 = pi35  & ~n11108;
  assign n11110 = pi35  & n11107;
  assign n11111 = ~n11107 & ~n11108;
  assign n11112 = ~pi35  & ~n11107;
  assign n11113 = ~n39449 & ~n39450;
  assign n11114 = n11098 & ~n11113;
  assign n11115 = ~n11098 & n11113;
  assign n11116 = n11098 & ~n11114;
  assign n11117 = n11098 & n11113;
  assign n11118 = ~n11113 & ~n11114;
  assign n11119 = ~n11098 & ~n11113;
  assign n11120 = ~n39451 & ~n39452;
  assign n11121 = ~n11114 & ~n11115;
  assign n11122 = n10894 & n39453;
  assign n11123 = ~n10894 & ~n39453;
  assign n11124 = ~n11122 & ~n11123;
  assign n11125 = n649 & n4524;
  assign n11126 = pi92  & n37496;
  assign n11127 = pi94  & n662;
  assign n11128 = pi93  & n664;
  assign n11129 = ~n11127 & ~n11128;
  assign n11130 = ~n11126 & ~n11128;
  assign n11131 = ~n11127 & n11130;
  assign n11132 = ~n11126 & n11129;
  assign n11133 = ~n11125 & n39454;
  assign n11134 = pi32  & ~n11133;
  assign n11135 = pi32  & ~n11134;
  assign n11136 = pi32  & n11133;
  assign n11137 = ~n11133 & ~n11134;
  assign n11138 = ~pi32  & ~n11133;
  assign n11139 = ~n39455 & ~n39456;
  assign n11140 = ~n11124 & n11139;
  assign n11141 = n11124 & ~n11139;
  assign n11142 = ~n11140 & ~n11141;
  assign n11143 = ~n9573 & n11142;
  assign n11144 = n9573 & ~n11142;
  assign n11145 = ~n11143 & ~n11144;
  assign n11146 = n607 & n5630;
  assign n11147 = pi95  & n37489;
  assign n11148 = pi97  & n620;
  assign n11149 = pi96  & n622;
  assign n11150 = ~n11148 & ~n11149;
  assign n11151 = ~n11147 & ~n11149;
  assign n11152 = ~n11148 & n11151;
  assign n11153 = ~n11147 & n11150;
  assign n11154 = ~n11146 & n39457;
  assign n11155 = pi29  & ~n11154;
  assign n11156 = pi29  & ~n11155;
  assign n11157 = pi29  & n11154;
  assign n11158 = ~n11154 & ~n11155;
  assign n11159 = ~pi29  & ~n11154;
  assign n11160 = ~n39458 & ~n39459;
  assign n11161 = n11145 & ~n11160;
  assign n11162 = ~n11145 & n11160;
  assign n11163 = n11145 & ~n11161;
  assign n11164 = n11145 & n11160;
  assign n11165 = ~n11160 & ~n11161;
  assign n11166 = ~n11145 & ~n11160;
  assign n11167 = ~n39460 & ~n39461;
  assign n11168 = ~n11161 & ~n11162;
  assign n11169 = ~n10893 & ~n39462;
  assign n11170 = n10893 & n39462;
  assign n11171 = ~n10893 & n39462;
  assign n11172 = n10893 & ~n39462;
  assign n11173 = ~n11171 & ~n11172;
  assign n11174 = ~n11169 & ~n11170;
  assign n11175 = ~n10892 & ~n39463;
  assign n11176 = n10892 & n39463;
  assign n11177 = ~n11175 & ~n11176;
  assign n11178 = n10877 & ~n11177;
  assign n11179 = ~n10877 & n11177;
  assign n11180 = ~n11178 & ~n11179;
  assign n11181 = n5576 & n6787;
  assign n11182 = pi101  & n38406;
  assign n11183 = pi103  & n5591;
  assign n11184 = pi102  & n5593;
  assign n11185 = ~n11183 & ~n11184;
  assign n11186 = ~n11182 & ~n11184;
  assign n11187 = ~n11183 & n11186;
  assign n11188 = ~n11182 & n11185;
  assign n11189 = ~n11181 & n39464;
  assign n11190 = pi23  & ~n11189;
  assign n11191 = pi23  & ~n11190;
  assign n11192 = pi23  & n11189;
  assign n11193 = ~n11189 & ~n11190;
  assign n11194 = ~pi23  & ~n11189;
  assign n11195 = ~n39465 & ~n39466;
  assign n11196 = n11180 & ~n11195;
  assign n11197 = ~n11180 & n11195;
  assign n11198 = n11180 & ~n11196;
  assign n11199 = n11180 & n11195;
  assign n11200 = ~n11195 & ~n11196;
  assign n11201 = ~n11180 & ~n11195;
  assign n11202 = ~n39467 & ~n39468;
  assign n11203 = ~n11196 & ~n11197;
  assign n11204 = n10876 & n39469;
  assign n11205 = ~n10876 & ~n39469;
  assign n11206 = ~n11204 & ~n11205;
  assign n11207 = n6785 & n8209;
  assign n11208 = pi104  & n38631;
  assign n11209 = pi106  & n6800;
  assign n11210 = pi105  & n6802;
  assign n11211 = ~n11209 & ~n11210;
  assign n11212 = ~n11208 & ~n11210;
  assign n11213 = ~n11209 & n11212;
  assign n11214 = ~n11208 & n11211;
  assign n11215 = ~n11207 & n39470;
  assign n11216 = pi20  & ~n11215;
  assign n11217 = pi20  & ~n11216;
  assign n11218 = pi20  & n11215;
  assign n11219 = ~n11215 & ~n11216;
  assign n11220 = ~pi20  & ~n11215;
  assign n11221 = ~n39471 & ~n39472;
  assign n11222 = ~n11206 & n11221;
  assign n11223 = n11206 & ~n11221;
  assign n11224 = ~n11222 & ~n11223;
  assign n11225 = ~n9658 & n11224;
  assign n11226 = n9658 & ~n11224;
  assign n11227 = ~n11225 & ~n11226;
  assign n11228 = ~n10875 & n11227;
  assign n11229 = n10875 & ~n11227;
  assign n11230 = ~n10875 & ~n11228;
  assign n11231 = ~n10875 & ~n11227;
  assign n11232 = n11227 & ~n11228;
  assign n11233 = n10875 & n11227;
  assign n11234 = ~n39473 & ~n39474;
  assign n11235 = ~n11228 & ~n11229;
  assign n11236 = ~n10860 & ~n39475;
  assign n11237 = n10860 & ~n39474;
  assign n11238 = ~n39473 & n11237;
  assign n11239 = n10860 & n39475;
  assign n11240 = ~n11236 & ~n39476;
  assign n11241 = ~n10859 & n11240;
  assign n11242 = n10859 & ~n11240;
  assign n11243 = ~n10859 & ~n11241;
  assign n11244 = ~n10859 & ~n11240;
  assign n11245 = n11240 & ~n11241;
  assign n11246 = n10859 & n11240;
  assign n11247 = ~n39477 & ~n39478;
  assign n11248 = ~n11241 & ~n11242;
  assign n11249 = ~n10842 & ~n39479;
  assign n11250 = n10842 & ~n39478;
  assign n11251 = ~n39477 & n11250;
  assign n11252 = n10842 & n39479;
  assign n11253 = ~n11249 & ~n39480;
  assign n11254 = ~n550 & n11253;
  assign n11255 = n10838 & ~n10840;
  assign n11256 = ~n10841 & ~n11255;
  assign n11257 = n513 & ~n515;
  assign n11258 = ~n516 & ~n11257;
  assign n11259 = n269 & n11258;
  assign n11260 = pi112  & n37475;
  assign n11261 = pi114  & n536;
  assign n11262 = pi113  & n538;
  assign n11263 = ~n11261 & ~n11262;
  assign n11264 = ~n11260 & ~n11262;
  assign n11265 = ~n11261 & n11264;
  assign n11266 = ~n11260 & n11263;
  assign n11267 = ~n11259 & n39481;
  assign n11268 = pi11  & ~n11267;
  assign n11269 = pi11  & ~n11268;
  assign n11270 = pi11  & n11267;
  assign n11271 = ~n11267 & ~n11268;
  assign n11272 = ~pi11  & ~n11267;
  assign n11273 = ~n39482 & ~n39483;
  assign n11274 = n11256 & ~n11273;
  assign n11275 = n509 & ~n511;
  assign n11276 = ~n512 & ~n11275;
  assign n11277 = n269 & n11276;
  assign n11278 = pi111  & n37475;
  assign n11279 = pi113  & n536;
  assign n11280 = pi112  & n538;
  assign n11281 = ~n11279 & ~n11280;
  assign n11282 = ~n11278 & ~n11280;
  assign n11283 = ~n11279 & n11282;
  assign n11284 = ~n11278 & n11281;
  assign n11285 = ~n11277 & n39484;
  assign n11286 = pi11  & ~n11285;
  assign n11287 = pi11  & ~n11286;
  assign n11288 = pi11  & n11285;
  assign n11289 = ~n11285 & ~n11286;
  assign n11290 = ~pi11  & ~n11285;
  assign n11291 = ~n39485 & ~n39486;
  assign n11292 = n10834 & ~n10836;
  assign n11293 = ~n10837 & ~n11292;
  assign n11294 = ~n11291 & n11293;
  assign n11295 = n269 & n10844;
  assign n11296 = pi110  & n37475;
  assign n11297 = pi112  & n536;
  assign n11298 = pi111  & n538;
  assign n11299 = ~n11297 & ~n11298;
  assign n11300 = ~n11296 & ~n11298;
  assign n11301 = ~n11297 & n11300;
  assign n11302 = ~n11296 & n11299;
  assign n11303 = ~n11295 & n39487;
  assign n11304 = pi11  & ~n11303;
  assign n11305 = pi11  & ~n11304;
  assign n11306 = pi11  & n11303;
  assign n11307 = ~n11303 & ~n11304;
  assign n11308 = ~pi11  & ~n11303;
  assign n11309 = ~n39488 & ~n39489;
  assign n11310 = n10825 & ~n39400;
  assign n11311 = ~n39399 & n11310;
  assign n11312 = n10825 & n39401;
  assign n11313 = ~n10833 & ~n39490;
  assign n11314 = ~n11309 & n11313;
  assign n11315 = n269 & n565;
  assign n11316 = pi109  & n37475;
  assign n11317 = pi111  & n536;
  assign n11318 = pi110  & n538;
  assign n11319 = ~n11317 & ~n11318;
  assign n11320 = ~n11316 & ~n11318;
  assign n11321 = ~n11317 & n11320;
  assign n11322 = ~n11316 & n11319;
  assign n11323 = ~n11315 & n39491;
  assign n11324 = pi11  & ~n11323;
  assign n11325 = pi11  & ~n11324;
  assign n11326 = pi11  & n11323;
  assign n11327 = ~n11323 & ~n11324;
  assign n11328 = ~pi11  & ~n11323;
  assign n11329 = ~n39492 & ~n39493;
  assign n11330 = n10819 & ~n10821;
  assign n11331 = ~n10819 & ~n39398;
  assign n11332 = ~n10820 & n10825;
  assign n11333 = ~n11331 & ~n11332;
  assign n11334 = ~n39398 & ~n11330;
  assign n11335 = ~n11329 & ~n39494;
  assign n11336 = n269 & n9678;
  assign n11337 = pi108  & n37475;
  assign n11338 = pi110  & n536;
  assign n11339 = pi109  & n538;
  assign n11340 = ~n11338 & ~n11339;
  assign n11341 = ~n11337 & ~n11339;
  assign n11342 = ~n11338 & n11341;
  assign n11343 = ~n11337 & n11340;
  assign n11344 = ~n11336 & n39495;
  assign n11345 = pi11  & ~n11344;
  assign n11346 = pi11  & ~n11345;
  assign n11347 = pi11  & n11344;
  assign n11348 = ~n11344 & ~n11345;
  assign n11349 = ~pi11  & ~n11344;
  assign n11350 = ~n39496 & ~n39497;
  assign n11351 = n10813 & ~n10815;
  assign n11352 = ~n10813 & ~n39397;
  assign n11353 = ~n10814 & n10819;
  assign n11354 = ~n11352 & ~n11353;
  assign n11355 = ~n39397 & ~n11351;
  assign n11356 = ~n11350 & ~n39498;
  assign n11357 = n269 & n9701;
  assign n11358 = pi107  & n37475;
  assign n11359 = pi109  & n536;
  assign n11360 = pi108  & n538;
  assign n11361 = ~n11359 & ~n11360;
  assign n11362 = ~n11358 & ~n11360;
  assign n11363 = ~n11359 & n11362;
  assign n11364 = ~n11358 & n11361;
  assign n11365 = ~n11357 & n39499;
  assign n11366 = pi11  & ~n11365;
  assign n11367 = pi11  & ~n11366;
  assign n11368 = pi11  & n11365;
  assign n11369 = ~n11365 & ~n11366;
  assign n11370 = ~pi11  & ~n11365;
  assign n11371 = ~n39500 & ~n39501;
  assign n11372 = n10809 & ~n10811;
  assign n11373 = ~n10812 & ~n11372;
  assign n11374 = ~n11371 & n11373;
  assign n11375 = n10800 & n39396;
  assign n11376 = ~n10808 & ~n11375;
  assign n11377 = n269 & n9277;
  assign n11378 = pi106  & n37475;
  assign n11379 = pi108  & n536;
  assign n11380 = pi107  & n538;
  assign n11381 = ~n11379 & ~n11380;
  assign n11382 = ~n11378 & ~n11380;
  assign n11383 = ~n11379 & n11382;
  assign n11384 = ~n11378 & n11381;
  assign n11385 = ~n11377 & n39502;
  assign n11386 = pi11  & ~n11385;
  assign n11387 = pi11  & ~n11386;
  assign n11388 = pi11  & n11385;
  assign n11389 = ~n11385 & ~n11386;
  assign n11390 = ~pi11  & ~n11385;
  assign n11391 = ~n39503 & ~n39504;
  assign n11392 = n11376 & ~n11391;
  assign n11393 = n10791 & n39393;
  assign n11394 = ~n10799 & ~n11393;
  assign n11395 = n269 & n8177;
  assign n11396 = pi105  & n37475;
  assign n11397 = pi107  & n536;
  assign n11398 = pi106  & n538;
  assign n11399 = ~n11397 & ~n11398;
  assign n11400 = ~n11396 & ~n11398;
  assign n11401 = ~n11397 & n11400;
  assign n11402 = ~n11396 & n11399;
  assign n11403 = ~n11395 & n39505;
  assign n11404 = pi11  & ~n11403;
  assign n11405 = pi11  & ~n11404;
  assign n11406 = pi11  & n11403;
  assign n11407 = ~n11403 & ~n11404;
  assign n11408 = ~pi11  & ~n11403;
  assign n11409 = ~n39506 & ~n39507;
  assign n11410 = n11394 & ~n11409;
  assign n11411 = n10782 & n39390;
  assign n11412 = ~n10790 & ~n11411;
  assign n11413 = n269 & n8209;
  assign n11414 = pi104  & n37475;
  assign n11415 = pi106  & n536;
  assign n11416 = pi105  & n538;
  assign n11417 = ~n11415 & ~n11416;
  assign n11418 = ~n11414 & ~n11416;
  assign n11419 = ~n11415 & n11418;
  assign n11420 = ~n11414 & n11417;
  assign n11421 = ~n11413 & n39508;
  assign n11422 = pi11  & ~n11421;
  assign n11423 = pi11  & ~n11422;
  assign n11424 = pi11  & n11421;
  assign n11425 = ~n11421 & ~n11422;
  assign n11426 = ~pi11  & ~n11421;
  assign n11427 = ~n39509 & ~n39510;
  assign n11428 = n11412 & ~n11427;
  assign n11429 = ~n11412 & n11427;
  assign n11430 = ~n11428 & ~n11429;
  assign n11431 = n10773 & n39387;
  assign n11432 = ~n10781 & ~n11431;
  assign n11433 = n269 & n8229;
  assign n11434 = pi103  & n37475;
  assign n11435 = pi105  & n536;
  assign n11436 = pi104  & n538;
  assign n11437 = ~n11435 & ~n11436;
  assign n11438 = ~n11434 & ~n11436;
  assign n11439 = ~n11435 & n11438;
  assign n11440 = ~n11434 & n11437;
  assign n11441 = ~n11433 & n39511;
  assign n11442 = pi11  & ~n11441;
  assign n11443 = pi11  & ~n11442;
  assign n11444 = pi11  & n11441;
  assign n11445 = ~n11441 & ~n11442;
  assign n11446 = ~pi11  & ~n11441;
  assign n11447 = ~n39512 & ~n39513;
  assign n11448 = n11432 & ~n11447;
  assign n11449 = n10764 & n39384;
  assign n11450 = ~n10772 & ~n11449;
  assign n11451 = n269 & n8136;
  assign n11452 = pi102  & n37475;
  assign n11453 = pi104  & n536;
  assign n11454 = pi103  & n538;
  assign n11455 = ~n11453 & ~n11454;
  assign n11456 = ~n11452 & ~n11454;
  assign n11457 = ~n11453 & n11456;
  assign n11458 = ~n11452 & n11455;
  assign n11459 = ~n11451 & n39514;
  assign n11460 = pi11  & ~n11459;
  assign n11461 = pi11  & ~n11460;
  assign n11462 = pi11  & n11459;
  assign n11463 = ~n11459 & ~n11460;
  assign n11464 = ~pi11  & ~n11459;
  assign n11465 = ~n39515 & ~n39516;
  assign n11466 = n11450 & ~n11465;
  assign n11467 = n10760 & ~n10762;
  assign n11468 = ~n10763 & ~n11467;
  assign n11469 = n269 & n6787;
  assign n11470 = pi101  & n37475;
  assign n11471 = pi103  & n536;
  assign n11472 = pi102  & n538;
  assign n11473 = ~n11471 & ~n11472;
  assign n11474 = ~n11470 & ~n11472;
  assign n11475 = ~n11471 & n11474;
  assign n11476 = ~n11470 & n11473;
  assign n11477 = ~n11469 & n39517;
  assign n11478 = pi11  & ~n11477;
  assign n11479 = pi11  & ~n11478;
  assign n11480 = pi11  & n11477;
  assign n11481 = ~n11477 & ~n11478;
  assign n11482 = ~pi11  & ~n11477;
  assign n11483 = ~n39518 & ~n39519;
  assign n11484 = n11468 & ~n11483;
  assign n11485 = n10751 & n39381;
  assign n11486 = ~n10759 & ~n11485;
  assign n11487 = n269 & n6819;
  assign n11488 = pi100  & n37475;
  assign n11489 = pi102  & n536;
  assign n11490 = pi101  & n538;
  assign n11491 = ~n11489 & ~n11490;
  assign n11492 = ~n11488 & ~n11490;
  assign n11493 = ~n11489 & n11492;
  assign n11494 = ~n11488 & n11491;
  assign n11495 = ~n11487 & n39520;
  assign n11496 = pi11  & ~n11495;
  assign n11497 = pi11  & ~n11496;
  assign n11498 = pi11  & n11495;
  assign n11499 = ~n11495 & ~n11496;
  assign n11500 = ~pi11  & ~n11495;
  assign n11501 = ~n39521 & ~n39522;
  assign n11502 = n11486 & ~n11501;
  assign n11503 = n10742 & n39378;
  assign n11504 = ~n10750 & ~n11503;
  assign n11505 = n269 & n6839;
  assign n11506 = pi99  & n37475;
  assign n11507 = pi101  & n536;
  assign n11508 = pi100  & n538;
  assign n11509 = ~n11507 & ~n11508;
  assign n11510 = ~n11506 & ~n11508;
  assign n11511 = ~n11507 & n11510;
  assign n11512 = ~n11506 & n11509;
  assign n11513 = ~n11505 & n39523;
  assign n11514 = pi11  & ~n11513;
  assign n11515 = pi11  & ~n11514;
  assign n11516 = pi11  & n11513;
  assign n11517 = ~n11513 & ~n11514;
  assign n11518 = ~pi11  & ~n11513;
  assign n11519 = ~n39524 & ~n39525;
  assign n11520 = n11504 & ~n11519;
  assign n11521 = n269 & n6474;
  assign n11522 = pi98  & n37475;
  assign n11523 = pi100  & n536;
  assign n11524 = pi99  & n538;
  assign n11525 = ~n11523 & ~n11524;
  assign n11526 = ~n11522 & ~n11524;
  assign n11527 = ~n11523 & n11526;
  assign n11528 = ~n11522 & n11525;
  assign n11529 = ~n11521 & n39526;
  assign n11530 = pi11  & ~n11529;
  assign n11531 = pi11  & ~n11530;
  assign n11532 = pi11  & n11529;
  assign n11533 = ~n11529 & ~n11530;
  assign n11534 = ~pi11  & ~n11529;
  assign n11535 = ~n39527 & ~n39528;
  assign n11536 = n10733 & n39375;
  assign n11537 = ~n10733 & n39375;
  assign n11538 = n10733 & ~n39375;
  assign n11539 = ~n11537 & ~n11538;
  assign n11540 = ~n10741 & ~n11536;
  assign n11541 = ~n11535 & ~n39529;
  assign n11542 = n10729 & ~n10731;
  assign n11543 = ~n10732 & ~n11542;
  assign n11544 = n269 & n5578;
  assign n11545 = pi97  & n37475;
  assign n11546 = pi99  & n536;
  assign n11547 = pi98  & n538;
  assign n11548 = ~n11546 & ~n11547;
  assign n11549 = ~n11545 & ~n11547;
  assign n11550 = ~n11546 & n11549;
  assign n11551 = ~n11545 & n11548;
  assign n11552 = ~n11544 & n39530;
  assign n11553 = pi11  & ~n11552;
  assign n11554 = pi11  & ~n11553;
  assign n11555 = pi11  & n11552;
  assign n11556 = ~n11552 & ~n11553;
  assign n11557 = ~pi11  & ~n11552;
  assign n11558 = ~n39531 & ~n39532;
  assign n11559 = n11543 & ~n11558;
  assign n11560 = n10725 & ~n10727;
  assign n11561 = ~n10728 & ~n11560;
  assign n11562 = n269 & n5610;
  assign n11563 = pi96  & n37475;
  assign n11564 = pi98  & n536;
  assign n11565 = pi97  & n538;
  assign n11566 = ~n11564 & ~n11565;
  assign n11567 = ~n11563 & ~n11565;
  assign n11568 = ~n11564 & n11567;
  assign n11569 = ~n11563 & n11566;
  assign n11570 = ~n11562 & n39533;
  assign n11571 = pi11  & ~n11570;
  assign n11572 = pi11  & ~n11571;
  assign n11573 = pi11  & n11570;
  assign n11574 = ~n11570 & ~n11571;
  assign n11575 = ~pi11  & ~n11570;
  assign n11576 = ~n39534 & ~n39535;
  assign n11577 = n11561 & ~n11576;
  assign n11578 = n10721 & ~n10723;
  assign n11579 = ~n10724 & ~n11578;
  assign n11580 = n269 & n5630;
  assign n11581 = pi95  & n37475;
  assign n11582 = pi97  & n536;
  assign n11583 = pi96  & n538;
  assign n11584 = ~n11582 & ~n11583;
  assign n11585 = ~n11581 & ~n11583;
  assign n11586 = ~n11582 & n11585;
  assign n11587 = ~n11581 & n11584;
  assign n11588 = ~n11580 & n39536;
  assign n11589 = pi11  & ~n11588;
  assign n11590 = pi11  & ~n11589;
  assign n11591 = pi11  & n11588;
  assign n11592 = ~n11588 & ~n11589;
  assign n11593 = ~pi11  & ~n11588;
  assign n11594 = ~n39537 & ~n39538;
  assign n11595 = n11579 & ~n11594;
  assign n11596 = n269 & n5281;
  assign n11597 = pi94  & n37475;
  assign n11598 = pi96  & n536;
  assign n11599 = pi95  & n538;
  assign n11600 = ~n11598 & ~n11599;
  assign n11601 = ~n11597 & ~n11599;
  assign n11602 = ~n11598 & n11601;
  assign n11603 = ~n11597 & n11600;
  assign n11604 = ~n11596 & n39539;
  assign n11605 = pi11  & ~n11604;
  assign n11606 = pi11  & ~n11605;
  assign n11607 = pi11  & n11604;
  assign n11608 = ~n11604 & ~n11605;
  assign n11609 = ~pi11  & ~n11604;
  assign n11610 = ~n39540 & ~n39541;
  assign n11611 = n10717 & ~n10719;
  assign n11612 = ~n10720 & ~n11611;
  assign n11613 = ~n11610 & n11612;
  assign n11614 = n269 & n4494;
  assign n11615 = pi93  & n37475;
  assign n11616 = pi95  & n536;
  assign n11617 = pi94  & n538;
  assign n11618 = ~n11616 & ~n11617;
  assign n11619 = ~n11615 & ~n11617;
  assign n11620 = ~n11616 & n11619;
  assign n11621 = ~n11615 & n11618;
  assign n11622 = ~n11614 & n39542;
  assign n11623 = pi11  & ~n11622;
  assign n11624 = pi11  & ~n11623;
  assign n11625 = pi11  & n11622;
  assign n11626 = ~n11622 & ~n11623;
  assign n11627 = ~pi11  & ~n11622;
  assign n11628 = ~n39543 & ~n39544;
  assign n11629 = n10708 & n39372;
  assign n11630 = ~n10708 & ~n10716;
  assign n11631 = ~n10708 & n39372;
  assign n11632 = ~n39372 & ~n10716;
  assign n11633 = n10708 & ~n39372;
  assign n11634 = ~n39545 & ~n39546;
  assign n11635 = ~n10716 & ~n11629;
  assign n11636 = ~n11628 & ~n39547;
  assign n11637 = n269 & n4524;
  assign n11638 = pi92  & n37475;
  assign n11639 = pi94  & n536;
  assign n11640 = pi93  & n538;
  assign n11641 = ~n11639 & ~n11640;
  assign n11642 = ~n11638 & ~n11640;
  assign n11643 = ~n11639 & n11642;
  assign n11644 = ~n11638 & n11641;
  assign n11645 = ~n11637 & n39548;
  assign n11646 = pi11  & ~n11645;
  assign n11647 = pi11  & ~n11646;
  assign n11648 = pi11  & n11645;
  assign n11649 = ~n11645 & ~n11646;
  assign n11650 = ~pi11  & ~n11645;
  assign n11651 = ~n39549 & ~n39550;
  assign n11652 = n10699 & n39369;
  assign n11653 = ~n10699 & n39369;
  assign n11654 = n10699 & ~n39369;
  assign n11655 = ~n11653 & ~n11654;
  assign n11656 = ~n10707 & ~n11652;
  assign n11657 = ~n11651 & ~n39551;
  assign n11658 = n269 & n4544;
  assign n11659 = pi91  & n37475;
  assign n11660 = pi93  & n536;
  assign n11661 = pi92  & n538;
  assign n11662 = ~n11660 & ~n11661;
  assign n11663 = ~n11659 & ~n11661;
  assign n11664 = ~n11660 & n11663;
  assign n11665 = ~n11659 & n11662;
  assign n11666 = ~n11658 & n39552;
  assign n11667 = pi11  & ~n11666;
  assign n11668 = pi11  & ~n11667;
  assign n11669 = pi11  & n11666;
  assign n11670 = ~n11666 & ~n11667;
  assign n11671 = ~pi11  & ~n11666;
  assign n11672 = ~n39553 & ~n39554;
  assign n11673 = n10695 & ~n10697;
  assign n11674 = ~n10698 & ~n11673;
  assign n11675 = ~n11672 & n11674;
  assign n11676 = n269 & n4453;
  assign n11677 = pi90  & n37475;
  assign n11678 = pi92  & n536;
  assign n11679 = pi91  & n538;
  assign n11680 = ~n11678 & ~n11679;
  assign n11681 = ~n11677 & ~n11679;
  assign n11682 = ~n11678 & n11681;
  assign n11683 = ~n11677 & n11680;
  assign n11684 = ~n11676 & n39555;
  assign n11685 = pi11  & ~n11684;
  assign n11686 = pi11  & ~n11685;
  assign n11687 = pi11  & n11684;
  assign n11688 = ~n11684 & ~n11685;
  assign n11689 = ~pi11  & ~n11684;
  assign n11690 = ~n39556 & ~n39557;
  assign n11691 = n10689 & ~n10691;
  assign n11692 = ~n10689 & ~n39366;
  assign n11693 = ~n10690 & n10695;
  assign n11694 = ~n11692 & ~n11693;
  assign n11695 = ~n39366 & ~n11691;
  assign n11696 = ~n11690 & ~n39558;
  assign n11697 = n10685 & ~n10687;
  assign n11698 = ~n10688 & ~n11697;
  assign n11699 = n269 & n594;
  assign n11700 = pi89  & n37475;
  assign n11701 = pi91  & n536;
  assign n11702 = pi90  & n538;
  assign n11703 = ~n11701 & ~n11702;
  assign n11704 = ~n11700 & ~n11702;
  assign n11705 = ~n11701 & n11704;
  assign n11706 = ~n11700 & n11703;
  assign n11707 = ~n11699 & n39559;
  assign n11708 = pi11  & ~n11707;
  assign n11709 = pi11  & ~n11708;
  assign n11710 = pi11  & n11707;
  assign n11711 = ~n11707 & ~n11708;
  assign n11712 = ~pi11  & ~n11707;
  assign n11713 = ~n39560 & ~n39561;
  assign n11714 = n11698 & ~n11713;
  assign n11715 = n269 & n3566;
  assign n11716 = pi88  & n37475;
  assign n11717 = pi90  & n536;
  assign n11718 = pi89  & n538;
  assign n11719 = ~n11717 & ~n11718;
  assign n11720 = ~n11716 & ~n11718;
  assign n11721 = ~n11717 & n11720;
  assign n11722 = ~n11716 & n11719;
  assign n11723 = ~n11715 & n39562;
  assign n11724 = pi11  & ~n11723;
  assign n11725 = pi11  & ~n11724;
  assign n11726 = pi11  & n11723;
  assign n11727 = ~n11723 & ~n11724;
  assign n11728 = ~pi11  & ~n11723;
  assign n11729 = ~n39563 & ~n39564;
  assign n11730 = n10681 & ~n10683;
  assign n11731 = ~n10684 & ~n11730;
  assign n11732 = ~n11729 & n11731;
  assign n11733 = n10672 & n39365;
  assign n11734 = ~n10680 & ~n11733;
  assign n11735 = n269 & n3591;
  assign n11736 = pi87  & n37475;
  assign n11737 = pi89  & n536;
  assign n11738 = pi88  & n538;
  assign n11739 = ~n11737 & ~n11738;
  assign n11740 = ~n11736 & ~n11738;
  assign n11741 = ~n11737 & n11740;
  assign n11742 = ~n11736 & n11739;
  assign n11743 = ~n11735 & n39565;
  assign n11744 = pi11  & ~n11743;
  assign n11745 = pi11  & ~n11744;
  assign n11746 = pi11  & n11743;
  assign n11747 = ~n11743 & ~n11744;
  assign n11748 = ~pi11  & ~n11743;
  assign n11749 = ~n39566 & ~n39567;
  assign n11750 = n11734 & ~n11749;
  assign n11751 = n269 & n3354;
  assign n11752 = pi86  & n37475;
  assign n11753 = pi88  & n536;
  assign n11754 = pi87  & n538;
  assign n11755 = ~n11753 & ~n11754;
  assign n11756 = ~n11752 & ~n11754;
  assign n11757 = ~n11753 & n11756;
  assign n11758 = ~n11752 & n11755;
  assign n11759 = ~n11751 & n39568;
  assign n11760 = pi11  & ~n11759;
  assign n11761 = pi11  & ~n11760;
  assign n11762 = pi11  & n11759;
  assign n11763 = ~n11759 & ~n11760;
  assign n11764 = ~pi11  & ~n11759;
  assign n11765 = ~n39569 & ~n39570;
  assign n11766 = n10663 & n39362;
  assign n11767 = ~n10663 & n39362;
  assign n11768 = n10663 & ~n39362;
  assign n11769 = ~n11767 & ~n11768;
  assign n11770 = ~n10671 & ~n11766;
  assign n11771 = ~n11765 & ~n39571;
  assign n11772 = n269 & n636;
  assign n11773 = pi85  & n37475;
  assign n11774 = pi87  & n536;
  assign n11775 = pi86  & n538;
  assign n11776 = ~n11774 & ~n11775;
  assign n11777 = ~n11773 & ~n11775;
  assign n11778 = ~n11774 & n11777;
  assign n11779 = ~n11773 & n11776;
  assign n11780 = ~n11772 & n39572;
  assign n11781 = pi11  & ~n11780;
  assign n11782 = pi11  & ~n11781;
  assign n11783 = pi11  & n11780;
  assign n11784 = ~n11780 & ~n11781;
  assign n11785 = ~pi11  & ~n11780;
  assign n11786 = ~n39573 & ~n39574;
  assign n11787 = n10657 & ~n10659;
  assign n11788 = ~n10657 & ~n39359;
  assign n11789 = ~n10658 & n10663;
  assign n11790 = ~n11788 & ~n11789;
  assign n11791 = ~n39359 & ~n11787;
  assign n11792 = ~n11786 & ~n39575;
  assign n11793 = n10648 & n39358;
  assign n11794 = ~n10656 & ~n11793;
  assign n11795 = n269 & n2779;
  assign n11796 = pi84  & n37475;
  assign n11797 = pi86  & n536;
  assign n11798 = pi85  & n538;
  assign n11799 = ~n11797 & ~n11798;
  assign n11800 = ~n11796 & ~n11798;
  assign n11801 = ~n11797 & n11800;
  assign n11802 = ~n11796 & n11799;
  assign n11803 = ~n11795 & n39576;
  assign n11804 = pi11  & ~n11803;
  assign n11805 = pi11  & ~n11804;
  assign n11806 = pi11  & n11803;
  assign n11807 = ~n11803 & ~n11804;
  assign n11808 = ~pi11  & ~n11803;
  assign n11809 = ~n39577 & ~n39578;
  assign n11810 = n11794 & ~n11809;
  assign n11811 = n10639 & n39355;
  assign n11812 = ~n10647 & ~n11811;
  assign n11813 = n269 & n2804;
  assign n11814 = pi83  & n37475;
  assign n11815 = pi85  & n536;
  assign n11816 = pi84  & n538;
  assign n11817 = ~n11815 & ~n11816;
  assign n11818 = ~n11814 & ~n11816;
  assign n11819 = ~n11815 & n11818;
  assign n11820 = ~n11814 & n11817;
  assign n11821 = ~n11813 & n39579;
  assign n11822 = pi11  & ~n11821;
  assign n11823 = pi11  & ~n11822;
  assign n11824 = pi11  & n11821;
  assign n11825 = ~n11821 & ~n11822;
  assign n11826 = ~pi11  & ~n11821;
  assign n11827 = ~n39580 & ~n39581;
  assign n11828 = n11812 & ~n11827;
  assign n11829 = n10630 & n39352;
  assign n11830 = ~n10638 & ~n11829;
  assign n11831 = n269 & n2591;
  assign n11832 = pi82  & n37475;
  assign n11833 = pi84  & n536;
  assign n11834 = pi83  & n538;
  assign n11835 = ~n11833 & ~n11834;
  assign n11836 = ~n11832 & ~n11834;
  assign n11837 = ~n11833 & n11836;
  assign n11838 = ~n11832 & n11835;
  assign n11839 = ~n11831 & n39582;
  assign n11840 = pi11  & ~n11839;
  assign n11841 = pi11  & ~n11840;
  assign n11842 = pi11  & n11839;
  assign n11843 = ~n11839 & ~n11840;
  assign n11844 = ~pi11  & ~n11839;
  assign n11845 = ~n39583 & ~n39584;
  assign n11846 = n11830 & ~n11845;
  assign n11847 = n10623 & n39349;
  assign n11848 = ~n10629 & ~n11847;
  assign n11849 = n269 & n2091;
  assign n11850 = pi81  & n37475;
  assign n11851 = pi83  & n536;
  assign n11852 = pi82  & n538;
  assign n11853 = ~n11851 & ~n11852;
  assign n11854 = ~n11850 & ~n11852;
  assign n11855 = ~n11851 & n11854;
  assign n11856 = ~n11850 & n11853;
  assign n11857 = ~n11849 & n39585;
  assign n11858 = pi11  & ~n11857;
  assign n11859 = pi11  & ~n11858;
  assign n11860 = pi11  & n11857;
  assign n11861 = ~n11857 & ~n11858;
  assign n11862 = ~pi11  & ~n11857;
  assign n11863 = ~n39586 & ~n39587;
  assign n11864 = n11848 & ~n11863;
  assign n11865 = n10614 & n39348;
  assign n11866 = ~n10622 & ~n11865;
  assign n11867 = n269 & n2134;
  assign n11868 = pi80  & n37475;
  assign n11869 = pi82  & n536;
  assign n11870 = pi81  & n538;
  assign n11871 = ~n11869 & ~n11870;
  assign n11872 = ~n11868 & ~n11870;
  assign n11873 = ~n11869 & n11872;
  assign n11874 = ~n11868 & n11871;
  assign n11875 = ~n11867 & n39588;
  assign n11876 = pi11  & ~n11875;
  assign n11877 = pi11  & ~n11876;
  assign n11878 = pi11  & n11875;
  assign n11879 = ~n11875 & ~n11876;
  assign n11880 = ~pi11  & ~n11875;
  assign n11881 = ~n39589 & ~n39590;
  assign n11882 = n11866 & ~n11881;
  assign n11883 = n269 & n2154;
  assign n11884 = pi79  & n37475;
  assign n11885 = pi81  & n536;
  assign n11886 = pi80  & n538;
  assign n11887 = ~n11885 & ~n11886;
  assign n11888 = ~n11884 & ~n11886;
  assign n11889 = ~n11885 & n11888;
  assign n11890 = ~n11884 & n11887;
  assign n11891 = ~n11883 & n39591;
  assign n11892 = pi11  & ~n11891;
  assign n11893 = pi11  & ~n11892;
  assign n11894 = pi11  & n11891;
  assign n11895 = ~n11891 & ~n11892;
  assign n11896 = ~pi11  & ~n11891;
  assign n11897 = ~n39592 & ~n39593;
  assign n11898 = n10605 & n39345;
  assign n11899 = ~n10605 & n39345;
  assign n11900 = n10605 & ~n39345;
  assign n11901 = ~n11899 & ~n11900;
  assign n11902 = ~n10613 & ~n11898;
  assign n11903 = ~n11897 & ~n39594;
  assign n11904 = ~n10322 & n10603;
  assign n11905 = ~n10604 & ~n11904;
  assign n11906 = n269 & n2063;
  assign n11907 = pi78  & n37475;
  assign n11908 = pi80  & n536;
  assign n11909 = pi79  & n538;
  assign n11910 = ~n11908 & ~n11909;
  assign n11911 = ~n11907 & ~n11909;
  assign n11912 = ~n11908 & n11911;
  assign n11913 = ~n11907 & n11910;
  assign n11914 = ~n11906 & n39595;
  assign n11915 = pi11  & ~n11914;
  assign n11916 = pi11  & ~n11915;
  assign n11917 = pi11  & n11914;
  assign n11918 = ~n11914 & ~n11915;
  assign n11919 = ~pi11  & ~n11914;
  assign n11920 = ~n39596 & ~n39597;
  assign n11921 = n11905 & ~n11920;
  assign n11922 = n10599 & ~n10601;
  assign n11923 = ~n10602 & ~n11922;
  assign n11924 = n269 & n678;
  assign n11925 = pi77  & n37475;
  assign n11926 = pi79  & n536;
  assign n11927 = pi78  & n538;
  assign n11928 = ~n11926 & ~n11927;
  assign n11929 = ~n11925 & ~n11927;
  assign n11930 = ~n11926 & n11929;
  assign n11931 = ~n11925 & n11928;
  assign n11932 = ~n11924 & n39598;
  assign n11933 = pi11  & ~n11932;
  assign n11934 = pi11  & ~n11933;
  assign n11935 = pi11  & n11932;
  assign n11936 = ~n11932 & ~n11933;
  assign n11937 = ~pi11  & ~n11932;
  assign n11938 = ~n39599 & ~n39600;
  assign n11939 = n11923 & ~n11938;
  assign n11940 = n10595 & ~n10597;
  assign n11941 = ~n10598 & ~n11940;
  assign n11942 = n269 & n1578;
  assign n11943 = pi76  & n37475;
  assign n11944 = pi78  & n536;
  assign n11945 = pi77  & n538;
  assign n11946 = ~n11944 & ~n11945;
  assign n11947 = ~n11943 & ~n11945;
  assign n11948 = ~n11944 & n11947;
  assign n11949 = ~n11943 & n11946;
  assign n11950 = ~n11942 & n39601;
  assign n11951 = pi11  & ~n11950;
  assign n11952 = pi11  & ~n11951;
  assign n11953 = pi11  & n11950;
  assign n11954 = ~n11950 & ~n11951;
  assign n11955 = ~pi11  & ~n11950;
  assign n11956 = ~n39602 & ~n39603;
  assign n11957 = n11941 & ~n11956;
  assign n11958 = n10586 & n39342;
  assign n11959 = ~n10594 & ~n11958;
  assign n11960 = n269 & n1596;
  assign n11961 = pi75  & n37475;
  assign n11962 = pi77  & n536;
  assign n11963 = pi76  & n538;
  assign n11964 = ~n11962 & ~n11963;
  assign n11965 = ~n11961 & ~n11963;
  assign n11966 = ~n11962 & n11965;
  assign n11967 = ~n11961 & n11964;
  assign n11968 = ~n11960 & n39604;
  assign n11969 = pi11  & ~n11968;
  assign n11970 = pi11  & ~n11969;
  assign n11971 = pi11  & n11968;
  assign n11972 = ~n11968 & ~n11969;
  assign n11973 = ~pi11  & ~n11968;
  assign n11974 = ~n39605 & ~n39606;
  assign n11975 = n11959 & ~n11974;
  assign n11976 = n269 & n1465;
  assign n11977 = pi74  & n37475;
  assign n11978 = pi76  & n536;
  assign n11979 = pi75  & n538;
  assign n11980 = ~n11978 & ~n11979;
  assign n11981 = ~n11977 & ~n11979;
  assign n11982 = ~n11978 & n11981;
  assign n11983 = ~n11977 & n11980;
  assign n11984 = ~n11976 & n39607;
  assign n11985 = pi11  & ~n11984;
  assign n11986 = pi11  & ~n11985;
  assign n11987 = pi11  & n11984;
  assign n11988 = ~n11984 & ~n11985;
  assign n11989 = ~pi11  & ~n11984;
  assign n11990 = ~n39608 & ~n39609;
  assign n11991 = n10582 & ~n10584;
  assign n11992 = ~n10585 & ~n11991;
  assign n11993 = ~n11990 & n11992;
  assign n11994 = n269 & n720;
  assign n11995 = pi73  & n37475;
  assign n11996 = pi75  & n536;
  assign n11997 = pi74  & n538;
  assign n11998 = ~n11996 & ~n11997;
  assign n11999 = ~n11995 & ~n11997;
  assign n12000 = ~n11996 & n11999;
  assign n12001 = ~n11995 & n11998;
  assign n12002 = ~n11994 & n39610;
  assign n12003 = pi11  & ~n12002;
  assign n12004 = pi11  & ~n12003;
  assign n12005 = pi11  & n12002;
  assign n12006 = ~n12002 & ~n12003;
  assign n12007 = ~pi11  & ~n12002;
  assign n12008 = ~n39611 & ~n39612;
  assign n12009 = n10578 & ~n10580;
  assign n12010 = ~n10581 & ~n12009;
  assign n12011 = ~n12008 & n12010;
  assign n12012 = n10574 & ~n10576;
  assign n12013 = ~n10577 & ~n12012;
  assign n12014 = n269 & n1218;
  assign n12015 = pi72  & n37475;
  assign n12016 = pi74  & n536;
  assign n12017 = pi73  & n538;
  assign n12018 = ~n12016 & ~n12017;
  assign n12019 = ~n12015 & ~n12017;
  assign n12020 = ~n12016 & n12019;
  assign n12021 = ~n12015 & n12018;
  assign n12022 = ~n12014 & n39613;
  assign n12023 = pi11  & ~n12022;
  assign n12024 = pi11  & ~n12023;
  assign n12025 = pi11  & n12022;
  assign n12026 = ~n12022 & ~n12023;
  assign n12027 = ~pi11  & ~n12022;
  assign n12028 = ~n39614 & ~n39615;
  assign n12029 = n12013 & ~n12028;
  assign n12030 = n269 & n1238;
  assign n12031 = pi71  & n37475;
  assign n12032 = pi73  & n536;
  assign n12033 = pi72  & n538;
  assign n12034 = ~n12032 & ~n12033;
  assign n12035 = ~n12031 & ~n12033;
  assign n12036 = ~n12032 & n12035;
  assign n12037 = ~n12031 & n12034;
  assign n12038 = ~n12030 & n39616;
  assign n12039 = pi11  & ~n12038;
  assign n12040 = pi11  & ~n12039;
  assign n12041 = pi11  & n12038;
  assign n12042 = ~n12038 & ~n12039;
  assign n12043 = ~pi11  & ~n12038;
  assign n12044 = ~n39617 & ~n39618;
  assign n12045 = n10565 & n39339;
  assign n12046 = ~n10565 & n39339;
  assign n12047 = n10565 & ~n39339;
  assign n12048 = ~n12046 & ~n12047;
  assign n12049 = ~n10573 & ~n12045;
  assign n12050 = ~n12044 & ~n39619;
  assign n12051 = n269 & n1124;
  assign n12052 = pi70  & n37475;
  assign n12053 = pi72  & n536;
  assign n12054 = pi71  & n538;
  assign n12055 = ~n12053 & ~n12054;
  assign n12056 = ~n12052 & ~n12054;
  assign n12057 = ~n12053 & n12056;
  assign n12058 = ~n12052 & n12055;
  assign n12059 = ~n12051 & n39620;
  assign n12060 = pi11  & ~n12059;
  assign n12061 = pi11  & ~n12060;
  assign n12062 = pi11  & n12059;
  assign n12063 = ~n12059 & ~n12060;
  assign n12064 = ~pi11  & ~n12059;
  assign n12065 = ~n39621 & ~n39622;
  assign n12066 = n10559 & ~n10561;
  assign n12067 = ~n10559 & ~n39336;
  assign n12068 = ~n10560 & n10565;
  assign n12069 = ~n12067 & ~n12068;
  assign n12070 = ~n39336 & ~n12066;
  assign n12071 = ~n12065 & ~n39623;
  assign n12072 = n269 & n927;
  assign n12073 = pi69  & n37475;
  assign n12074 = pi71  & n536;
  assign n12075 = pi70  & n538;
  assign n12076 = ~n12074 & ~n12075;
  assign n12077 = ~n12073 & ~n12075;
  assign n12078 = ~n12074 & n12077;
  assign n12079 = ~n12073 & n12076;
  assign n12080 = ~n12072 & n39624;
  assign n12081 = pi11  & ~n12080;
  assign n12082 = pi11  & ~n12081;
  assign n12083 = pi11  & n12080;
  assign n12084 = ~n12080 & ~n12081;
  assign n12085 = ~pi11  & ~n12080;
  assign n12086 = ~n39625 & ~n39626;
  assign n12087 = n10555 & ~n10557;
  assign n12088 = ~n10558 & ~n12087;
  assign n12089 = ~n12086 & n12088;
  assign n12090 = n10548 & n39335;
  assign n12091 = ~n10554 & ~n12090;
  assign n12092 = n269 & n972;
  assign n12093 = pi68  & n37475;
  assign n12094 = pi70  & n536;
  assign n12095 = pi69  & n538;
  assign n12096 = ~n12094 & ~n12095;
  assign n12097 = ~n12093 & ~n12095;
  assign n12098 = ~n12094 & n12097;
  assign n12099 = ~n12093 & n12096;
  assign n12100 = ~n12092 & n39627;
  assign n12101 = pi11  & ~n12100;
  assign n12102 = pi11  & ~n12101;
  assign n12103 = pi11  & n12100;
  assign n12104 = ~n12100 & ~n12101;
  assign n12105 = ~pi11  & ~n12100;
  assign n12106 = ~n39628 & ~n39629;
  assign n12107 = n12091 & ~n12106;
  assign n12108 = n269 & n990;
  assign n12109 = pi67  & n37475;
  assign n12110 = pi69  & n536;
  assign n12111 = pi68  & n538;
  assign n12112 = ~n12110 & ~n12111;
  assign n12113 = ~n12109 & ~n12111;
  assign n12114 = ~n12110 & n12113;
  assign n12115 = ~n12109 & n12112;
  assign n12116 = ~n12108 & n39630;
  assign n12117 = pi11  & ~n12116;
  assign n12118 = pi11  & ~n12117;
  assign n12119 = pi11  & n12116;
  assign n12120 = ~n12116 & ~n12117;
  assign n12121 = ~pi11  & ~n12116;
  assign n12122 = ~n39631 & ~n39632;
  assign n12123 = pi14  & ~n39327;
  assign n12124 = n39330 & ~n12123;
  assign n12125 = ~n39330 & n12123;
  assign n12126 = ~n39327 & n10530;
  assign n12127 = ~n39331 & ~n12126;
  assign n12128 = ~n12124 & ~n12125;
  assign n12129 = ~n12122 & n39633;
  assign n12130 = n269 & n871;
  assign n12131 = pi66  & n37475;
  assign n12132 = pi68  & n536;
  assign n12133 = pi67  & n538;
  assign n12134 = ~n12132 & ~n12133;
  assign n12135 = ~n12131 & ~n12133;
  assign n12136 = ~n12132 & n12135;
  assign n12137 = ~n12131 & n12134;
  assign n12138 = ~n12130 & n39634;
  assign n12139 = pi11  & ~n12138;
  assign n12140 = pi11  & ~n12139;
  assign n12141 = pi11  & n12138;
  assign n12142 = ~n12138 & ~n12139;
  assign n12143 = ~pi11  & ~n12138;
  assign n12144 = ~n39635 & ~n39636;
  assign n12145 = pi14  & n10504;
  assign n12146 = ~n10503 & n12145;
  assign n12147 = n10503 & ~n12145;
  assign n12148 = ~n10505 & n10509;
  assign n12149 = ~n39327 & ~n12148;
  assign n12150 = ~n12146 & ~n12147;
  assign n12151 = ~n12144 & n39637;
  assign n12152 = n269 & n37515;
  assign n12153 = pi65  & n536;
  assign n12154 = pi64  & n538;
  assign n12155 = ~n12153 & ~n12154;
  assign n12156 = ~n12152 & n12155;
  assign n12157 = pi64  & n37470;
  assign n12158 = pi11  & ~n12157;
  assign n12159 = pi11  & ~n12156;
  assign n12160 = pi11  & ~n12159;
  assign n12161 = ~n12156 & ~n12159;
  assign n12162 = ~n12160 & ~n12161;
  assign n12163 = n12158 & ~n12162;
  assign n12164 = n12156 & n12158;
  assign n12165 = pi64  & n37475;
  assign n12166 = pi65  & n538;
  assign n12167 = n269 & ~n37521;
  assign n12168 = pi66  & n536;
  assign n12169 = ~n12167 & ~n12168;
  assign n12170 = ~n12166 & ~n12167;
  assign n12171 = ~n12168 & n12170;
  assign n12172 = ~n12166 & ~n12168;
  assign n12173 = ~n12167 & n12172;
  assign n12174 = ~n12166 & n12169;
  assign n12175 = ~n12165 & ~n12166;
  assign n12176 = ~n12168 & n12175;
  assign n12177 = ~n12165 & n12172;
  assign n12178 = ~n12167 & n39640;
  assign n12179 = ~n12165 & n39639;
  assign n12180 = pi11  & ~n39641;
  assign n12181 = pi11  & ~n12180;
  assign n12182 = ~n39641 & ~n12180;
  assign n12183 = ~n12181 & ~n12182;
  assign n12184 = n39638 & ~n12183;
  assign n12185 = n39638 & n39641;
  assign n12186 = n10504 & n39642;
  assign n12187 = n269 & n847;
  assign n12188 = pi65  & n37475;
  assign n12189 = pi67  & n536;
  assign n12190 = pi66  & n538;
  assign n12191 = ~n12189 & ~n12190;
  assign n12192 = ~n12188 & ~n12190;
  assign n12193 = ~n12189 & n12192;
  assign n12194 = ~n12188 & n12191;
  assign n12195 = ~n12187 & n39643;
  assign n12196 = pi11  & ~n12195;
  assign n12197 = pi11  & ~n12196;
  assign n12198 = pi11  & n12195;
  assign n12199 = ~n12195 & ~n12196;
  assign n12200 = ~pi11  & ~n12195;
  assign n12201 = ~n39644 & ~n39645;
  assign n12202 = ~n10504 & ~n39642;
  assign n12203 = n10504 & ~n39642;
  assign n12204 = ~n10504 & n39642;
  assign n12205 = ~n12203 & ~n12204;
  assign n12206 = ~n12186 & ~n12202;
  assign n12207 = ~n12201 & ~n39646;
  assign n12208 = ~n12186 & ~n12207;
  assign n12209 = n12144 & ~n39637;
  assign n12210 = ~n12151 & ~n12209;
  assign n12211 = ~n12208 & n12210;
  assign n12212 = ~n12151 & ~n12211;
  assign n12213 = n12122 & ~n39633;
  assign n12214 = ~n12129 & ~n12213;
  assign n12215 = ~n12212 & ~n12213;
  assign n12216 = ~n12129 & n12215;
  assign n12217 = ~n12212 & n12214;
  assign n12218 = ~n12129 & ~n39647;
  assign n12219 = ~n12091 & n12106;
  assign n12220 = n12091 & ~n12107;
  assign n12221 = n12091 & n12106;
  assign n12222 = ~n12106 & ~n12107;
  assign n12223 = ~n12091 & ~n12106;
  assign n12224 = ~n39648 & ~n39649;
  assign n12225 = ~n12107 & ~n12219;
  assign n12226 = ~n12218 & ~n39650;
  assign n12227 = ~n12107 & ~n12226;
  assign n12228 = n12086 & ~n12088;
  assign n12229 = ~n12089 & ~n12228;
  assign n12230 = ~n12227 & n12229;
  assign n12231 = ~n12089 & ~n12230;
  assign n12232 = n12065 & n39623;
  assign n12233 = ~n12071 & ~n12232;
  assign n12234 = ~n12231 & n12233;
  assign n12235 = ~n12071 & ~n12234;
  assign n12236 = n12044 & n39619;
  assign n12237 = ~n12050 & ~n12236;
  assign n12238 = ~n12235 & n12237;
  assign n12239 = ~n12050 & ~n12238;
  assign n12240 = ~n12013 & n12028;
  assign n12241 = n12013 & ~n12029;
  assign n12242 = n12013 & n12028;
  assign n12243 = ~n12028 & ~n12029;
  assign n12244 = ~n12013 & ~n12028;
  assign n12245 = ~n39651 & ~n39652;
  assign n12246 = ~n12029 & ~n12240;
  assign n12247 = ~n12239 & ~n39653;
  assign n12248 = ~n12029 & ~n12247;
  assign n12249 = n12008 & ~n12010;
  assign n12250 = ~n12011 & ~n12249;
  assign n12251 = ~n12248 & n12250;
  assign n12252 = ~n12011 & ~n12251;
  assign n12253 = n11990 & ~n11992;
  assign n12254 = ~n11993 & ~n12253;
  assign n12255 = ~n12252 & n12254;
  assign n12256 = ~n11993 & ~n12255;
  assign n12257 = ~n11959 & n11974;
  assign n12258 = ~n11975 & ~n12257;
  assign n12259 = ~n12256 & n12258;
  assign n12260 = ~n11975 & ~n12259;
  assign n12261 = ~n11941 & n11956;
  assign n12262 = n11941 & ~n11957;
  assign n12263 = n11941 & n11956;
  assign n12264 = ~n11956 & ~n11957;
  assign n12265 = ~n11941 & ~n11956;
  assign n12266 = ~n39654 & ~n39655;
  assign n12267 = ~n11957 & ~n12261;
  assign n12268 = ~n12260 & ~n39656;
  assign n12269 = ~n11957 & ~n12268;
  assign n12270 = ~n11923 & n11938;
  assign n12271 = n11923 & ~n11939;
  assign n12272 = n11923 & n11938;
  assign n12273 = ~n11938 & ~n11939;
  assign n12274 = ~n11923 & ~n11938;
  assign n12275 = ~n39657 & ~n39658;
  assign n12276 = ~n11939 & ~n12270;
  assign n12277 = ~n12269 & ~n39659;
  assign n12278 = ~n11939 & ~n12277;
  assign n12279 = ~n11905 & n11920;
  assign n12280 = n11905 & ~n11921;
  assign n12281 = n11905 & n11920;
  assign n12282 = ~n11920 & ~n11921;
  assign n12283 = ~n11905 & ~n11920;
  assign n12284 = ~n39660 & ~n39661;
  assign n12285 = ~n11921 & ~n12279;
  assign n12286 = ~n12278 & ~n39662;
  assign n12287 = ~n11921 & ~n12286;
  assign n12288 = n11897 & n39594;
  assign n12289 = ~n11903 & ~n12288;
  assign n12290 = ~n12287 & n12289;
  assign n12291 = ~n11903 & ~n12290;
  assign n12292 = ~n11866 & n11881;
  assign n12293 = n11866 & ~n11882;
  assign n12294 = n11866 & n11881;
  assign n12295 = ~n11881 & ~n11882;
  assign n12296 = ~n11866 & ~n11881;
  assign n12297 = ~n39663 & ~n39664;
  assign n12298 = ~n11882 & ~n12292;
  assign n12299 = ~n12291 & ~n39665;
  assign n12300 = ~n11882 & ~n12299;
  assign n12301 = ~n11848 & n11863;
  assign n12302 = n11848 & ~n11864;
  assign n12303 = n11848 & n11863;
  assign n12304 = ~n11863 & ~n11864;
  assign n12305 = ~n11848 & ~n11863;
  assign n12306 = ~n39666 & ~n39667;
  assign n12307 = ~n11864 & ~n12301;
  assign n12308 = ~n12300 & ~n39668;
  assign n12309 = ~n11864 & ~n12308;
  assign n12310 = ~n11830 & n11845;
  assign n12311 = ~n11846 & ~n12310;
  assign n12312 = ~n12309 & ~n12310;
  assign n12313 = ~n11846 & n12312;
  assign n12314 = ~n12309 & n12311;
  assign n12315 = ~n11846 & ~n39669;
  assign n12316 = ~n11812 & n11827;
  assign n12317 = n11812 & ~n11828;
  assign n12318 = n11812 & n11827;
  assign n12319 = ~n11827 & ~n11828;
  assign n12320 = ~n11812 & ~n11827;
  assign n12321 = ~n39670 & ~n39671;
  assign n12322 = ~n11828 & ~n12316;
  assign n12323 = ~n12315 & ~n39672;
  assign n12324 = ~n11828 & ~n12323;
  assign n12325 = ~n11794 & n11809;
  assign n12326 = n11794 & ~n11810;
  assign n12327 = n11794 & n11809;
  assign n12328 = ~n11809 & ~n11810;
  assign n12329 = ~n11794 & ~n11809;
  assign n12330 = ~n39673 & ~n39674;
  assign n12331 = ~n11810 & ~n12325;
  assign n12332 = ~n12324 & ~n39675;
  assign n12333 = ~n11810 & ~n12332;
  assign n12334 = n11786 & n39575;
  assign n12335 = ~n11792 & ~n12334;
  assign n12336 = ~n12333 & n12335;
  assign n12337 = ~n11792 & ~n12336;
  assign n12338 = n11765 & n39571;
  assign n12339 = ~n11771 & ~n12338;
  assign n12340 = ~n12337 & n12339;
  assign n12341 = ~n11771 & ~n12340;
  assign n12342 = ~n11734 & n11749;
  assign n12343 = ~n11750 & ~n12342;
  assign n12344 = ~n12341 & ~n12342;
  assign n12345 = ~n11750 & n12344;
  assign n12346 = ~n12341 & n12343;
  assign n12347 = ~n11750 & ~n39676;
  assign n12348 = n11729 & ~n11731;
  assign n12349 = ~n11732 & ~n12348;
  assign n12350 = ~n12347 & n12349;
  assign n12351 = ~n11732 & ~n12350;
  assign n12352 = ~n11698 & n11713;
  assign n12353 = n11698 & ~n11714;
  assign n12354 = n11698 & n11713;
  assign n12355 = ~n11713 & ~n11714;
  assign n12356 = ~n11698 & ~n11713;
  assign n12357 = ~n39677 & ~n39678;
  assign n12358 = ~n11714 & ~n12352;
  assign n12359 = ~n12351 & ~n39679;
  assign n12360 = ~n11714 & ~n12359;
  assign n12361 = n11690 & n39558;
  assign n12362 = ~n11696 & ~n12361;
  assign n12363 = ~n12360 & n12362;
  assign n12364 = ~n11696 & ~n12363;
  assign n12365 = n11672 & ~n11674;
  assign n12366 = ~n11675 & ~n12365;
  assign n12367 = ~n12364 & n12366;
  assign n12368 = ~n11675 & ~n12367;
  assign n12369 = n11651 & n39551;
  assign n12370 = ~n11657 & ~n12369;
  assign n12371 = ~n12368 & n12370;
  assign n12372 = ~n11657 & ~n12371;
  assign n12373 = n11628 & n39547;
  assign n12374 = ~n11636 & ~n12373;
  assign n12375 = ~n12372 & n12374;
  assign n12376 = ~n11636 & ~n12375;
  assign n12377 = n11610 & ~n11612;
  assign n12378 = ~n11613 & ~n12377;
  assign n12379 = ~n12376 & n12378;
  assign n12380 = ~n11613 & ~n12379;
  assign n12381 = ~n11579 & n11594;
  assign n12382 = n11579 & ~n11595;
  assign n12383 = n11579 & n11594;
  assign n12384 = ~n11594 & ~n11595;
  assign n12385 = ~n11579 & ~n11594;
  assign n12386 = ~n39680 & ~n39681;
  assign n12387 = ~n11595 & ~n12381;
  assign n12388 = ~n12380 & ~n39682;
  assign n12389 = ~n11595 & ~n12388;
  assign n12390 = ~n11561 & n11576;
  assign n12391 = n11561 & ~n11577;
  assign n12392 = n11561 & n11576;
  assign n12393 = ~n11576 & ~n11577;
  assign n12394 = ~n11561 & ~n11576;
  assign n12395 = ~n39683 & ~n39684;
  assign n12396 = ~n11577 & ~n12390;
  assign n12397 = ~n12389 & ~n39685;
  assign n12398 = ~n11577 & ~n12397;
  assign n12399 = ~n11543 & n11558;
  assign n12400 = n11543 & ~n11559;
  assign n12401 = n11543 & n11558;
  assign n12402 = ~n11558 & ~n11559;
  assign n12403 = ~n11543 & ~n11558;
  assign n12404 = ~n39686 & ~n39687;
  assign n12405 = ~n11559 & ~n12399;
  assign n12406 = ~n12398 & ~n39688;
  assign n12407 = ~n11559 & ~n12406;
  assign n12408 = n11535 & n39529;
  assign n12409 = ~n11541 & ~n12408;
  assign n12410 = ~n12407 & n12409;
  assign n12411 = ~n11541 & ~n12410;
  assign n12412 = ~n11504 & n11519;
  assign n12413 = n11504 & ~n11520;
  assign n12414 = n11504 & n11519;
  assign n12415 = ~n11519 & ~n11520;
  assign n12416 = ~n11504 & ~n11519;
  assign n12417 = ~n39689 & ~n39690;
  assign n12418 = ~n11520 & ~n12412;
  assign n12419 = ~n12411 & ~n39691;
  assign n12420 = ~n11520 & ~n12419;
  assign n12421 = ~n11486 & n11501;
  assign n12422 = n11486 & ~n11502;
  assign n12423 = n11486 & n11501;
  assign n12424 = ~n11501 & ~n11502;
  assign n12425 = ~n11486 & ~n11501;
  assign n12426 = ~n39692 & ~n39693;
  assign n12427 = ~n11502 & ~n12421;
  assign n12428 = ~n12420 & ~n39694;
  assign n12429 = ~n11502 & ~n12428;
  assign n12430 = ~n11468 & n11483;
  assign n12431 = n11468 & ~n11484;
  assign n12432 = n11468 & n11483;
  assign n12433 = ~n11483 & ~n11484;
  assign n12434 = ~n11468 & ~n11483;
  assign n12435 = ~n39695 & ~n39696;
  assign n12436 = ~n11484 & ~n12430;
  assign n12437 = ~n12429 & ~n39697;
  assign n12438 = ~n11484 & ~n12437;
  assign n12439 = ~n11450 & n11465;
  assign n12440 = n11450 & ~n11466;
  assign n12441 = n11450 & n11465;
  assign n12442 = ~n11465 & ~n11466;
  assign n12443 = ~n11450 & ~n11465;
  assign n12444 = ~n39698 & ~n39699;
  assign n12445 = ~n11466 & ~n12439;
  assign n12446 = ~n12438 & ~n39700;
  assign n12447 = ~n11466 & ~n12446;
  assign n12448 = ~n11432 & n11447;
  assign n12449 = n11432 & ~n11448;
  assign n12450 = n11432 & n11447;
  assign n12451 = ~n11447 & ~n11448;
  assign n12452 = ~n11432 & ~n11447;
  assign n12453 = ~n39701 & ~n39702;
  assign n12454 = ~n11448 & ~n12448;
  assign n12455 = ~n12447 & ~n39703;
  assign n12456 = ~n11448 & ~n12455;
  assign n12457 = n11430 & ~n12456;
  assign n12458 = ~n11428 & ~n12457;
  assign n12459 = ~n11394 & n11409;
  assign n12460 = ~n11410 & ~n12459;
  assign n12461 = ~n12458 & ~n12459;
  assign n12462 = ~n11410 & n12461;
  assign n12463 = ~n12458 & n12460;
  assign n12464 = ~n11410 & ~n39704;
  assign n12465 = ~n11376 & n11391;
  assign n12466 = ~n11392 & ~n12465;
  assign n12467 = ~n12464 & ~n12465;
  assign n12468 = ~n11392 & n12467;
  assign n12469 = ~n12464 & n12466;
  assign n12470 = ~n11392 & ~n39705;
  assign n12471 = n11371 & ~n11373;
  assign n12472 = ~n11371 & ~n11374;
  assign n12473 = ~n11371 & ~n11373;
  assign n12474 = n11373 & ~n11374;
  assign n12475 = n11371 & n11373;
  assign n12476 = ~n39706 & ~n39707;
  assign n12477 = ~n11374 & ~n12471;
  assign n12478 = ~n12470 & ~n39708;
  assign n12479 = ~n11374 & ~n12478;
  assign n12480 = n11350 & n39498;
  assign n12481 = ~n11356 & ~n12480;
  assign n12482 = ~n12479 & n12481;
  assign n12483 = ~n11356 & ~n12482;
  assign n12484 = n11329 & n39494;
  assign n12485 = ~n39494 & ~n11335;
  assign n12486 = n11329 & ~n39494;
  assign n12487 = ~n11329 & ~n11335;
  assign n12488 = ~n11329 & n39494;
  assign n12489 = ~n39709 & ~n39710;
  assign n12490 = ~n11335 & ~n12484;
  assign n12491 = ~n12483 & ~n39711;
  assign n12492 = ~n11335 & ~n12491;
  assign n12493 = n11309 & ~n11313;
  assign n12494 = ~n11309 & ~n11314;
  assign n12495 = ~n11309 & ~n11313;
  assign n12496 = n11313 & ~n11314;
  assign n12497 = n11309 & n11313;
  assign n12498 = ~n39712 & ~n39713;
  assign n12499 = ~n11314 & ~n12493;
  assign n12500 = ~n12492 & ~n39714;
  assign n12501 = ~n11314 & ~n12500;
  assign n12502 = n11291 & ~n11293;
  assign n12503 = ~n11294 & ~n12502;
  assign n12504 = ~n12501 & n12503;
  assign n12505 = ~n11294 & ~n12504;
  assign n12506 = ~n11256 & n11273;
  assign n12507 = n11256 & ~n11274;
  assign n12508 = n11256 & n11273;
  assign n12509 = ~n11273 & ~n11274;
  assign n12510 = ~n11256 & ~n11273;
  assign n12511 = ~n39715 & ~n39716;
  assign n12512 = ~n11274 & ~n12506;
  assign n12513 = ~n12505 & ~n39717;
  assign n12514 = ~n11274 & ~n12513;
  assign n12515 = n550 & ~n11253;
  assign n12516 = ~n550 & ~n11254;
  assign n12517 = ~n550 & ~n11253;
  assign n12518 = n11253 & ~n11254;
  assign n12519 = n550 & n11253;
  assign n12520 = ~n39718 & ~n39719;
  assign n12521 = ~n11254 & ~n12515;
  assign n12522 = ~n12514 & ~n39720;
  assign n12523 = ~n11254 & ~n12522;
  assign n12524 = ~n519 & ~n521;
  assign n12525 = ~pi115  & ~pi116 ;
  assign n12526 = pi115  & pi116 ;
  assign n12527 = ~n12525 & ~n12526;
  assign n12528 = ~n12524 & n12527;
  assign n12529 = n12524 & ~n12527;
  assign n12530 = ~n12528 & ~n12529;
  assign n12531 = n269 & n12530;
  assign n12532 = pi114  & n37475;
  assign n12533 = pi116  & n536;
  assign n12534 = pi115  & n538;
  assign n12535 = ~n12533 & ~n12534;
  assign n12536 = ~n12532 & ~n12534;
  assign n12537 = ~n12533 & n12536;
  assign n12538 = ~n12532 & n12535;
  assign n12539 = ~n12531 & n39721;
  assign n12540 = pi11  & ~n12539;
  assign n12541 = pi11  & ~n12540;
  assign n12542 = pi11  & n12539;
  assign n12543 = ~n12539 & ~n12540;
  assign n12544 = ~pi11  & ~n12539;
  assign n12545 = ~n39722 & ~n39723;
  assign n12546 = ~n11241 & ~n11249;
  assign n12547 = n563 & n11276;
  assign n12548 = pi111  & n37482;
  assign n12549 = pi113  & n578;
  assign n12550 = pi112  & n580;
  assign n12551 = ~n12549 & ~n12550;
  assign n12552 = ~n12548 & ~n12550;
  assign n12553 = ~n12549 & n12552;
  assign n12554 = ~n12548 & n12551;
  assign n12555 = ~n12547 & n39724;
  assign n12556 = pi14  & ~n12555;
  assign n12557 = pi14  & ~n12556;
  assign n12558 = pi14  & n12555;
  assign n12559 = ~n12555 & ~n12556;
  assign n12560 = ~pi14  & ~n12555;
  assign n12561 = ~n39725 & ~n39726;
  assign n12562 = ~n11228 & ~n11236;
  assign n12563 = n8175 & n9678;
  assign n12564 = pi108  & n38895;
  assign n12565 = pi110  & n8190;
  assign n12566 = pi109  & n8192;
  assign n12567 = ~n12565 & ~n12566;
  assign n12568 = ~n12564 & ~n12566;
  assign n12569 = ~n12565 & n12568;
  assign n12570 = ~n12564 & n12567;
  assign n12571 = ~n12563 & n39727;
  assign n12572 = pi17  & ~n12571;
  assign n12573 = pi17  & ~n12572;
  assign n12574 = pi17  & n12571;
  assign n12575 = ~n12571 & ~n12572;
  assign n12576 = ~pi17  & ~n12571;
  assign n12577 = ~n39728 & ~n39729;
  assign n12578 = ~n11223 & ~n11225;
  assign n12579 = ~n11196 & ~n11205;
  assign n12580 = ~n11175 & ~n11179;
  assign n12581 = ~n11161 & ~n11169;
  assign n12582 = n607 & n5610;
  assign n12583 = pi96  & n37489;
  assign n12584 = pi98  & n620;
  assign n12585 = pi97  & n622;
  assign n12586 = ~n12584 & ~n12585;
  assign n12587 = ~n12583 & ~n12585;
  assign n12588 = ~n12584 & n12587;
  assign n12589 = ~n12583 & n12586;
  assign n12590 = ~n12582 & n39730;
  assign n12591 = pi29  & ~n12590;
  assign n12592 = pi29  & ~n12591;
  assign n12593 = pi29  & n12590;
  assign n12594 = ~n12590 & ~n12591;
  assign n12595 = ~pi29  & ~n12590;
  assign n12596 = ~n39731 & ~n39732;
  assign n12597 = ~n11141 & ~n11143;
  assign n12598 = ~n11114 & ~n11123;
  assign n12599 = ~n11088 & ~n11097;
  assign n12600 = ~n11067 & ~n11070;
  assign n12601 = n733 & n2779;
  assign n12602 = pi84  & n37510;
  assign n12603 = pi86  & n746;
  assign n12604 = pi85  & n748;
  assign n12605 = ~n12603 & ~n12604;
  assign n12606 = ~n12602 & ~n12604;
  assign n12607 = ~n12603 & n12606;
  assign n12608 = ~n12602 & n12605;
  assign n12609 = ~n12601 & n39733;
  assign n12610 = pi41  & ~n12609;
  assign n12611 = pi41  & ~n12610;
  assign n12612 = pi41  & n12609;
  assign n12613 = ~n12609 & ~n12610;
  assign n12614 = ~pi41  & ~n12609;
  assign n12615 = ~n39734 & ~n39735;
  assign n12616 = ~n11054 & ~n11062;
  assign n12617 = ~n11048 & ~n11051;
  assign n12618 = n785 & n2063;
  assign n12619 = pi78  & n37520;
  assign n12620 = pi80  & n787;
  assign n12621 = pi79  & n795;
  assign n12622 = ~n12620 & ~n12621;
  assign n12623 = ~n12619 & ~n12621;
  assign n12624 = ~n12620 & n12623;
  assign n12625 = ~n12619 & n12622;
  assign n12626 = ~n12618 & n39736;
  assign n12627 = pi47  & ~n12626;
  assign n12628 = pi47  & ~n12627;
  assign n12629 = pi47  & n12626;
  assign n12630 = ~n12626 & ~n12627;
  assign n12631 = ~pi47  & ~n12626;
  assign n12632 = ~n39737 & ~n39738;
  assign n12633 = ~n11043 & ~n11045;
  assign n12634 = ~n11036 & ~n11039;
  assign n12635 = ~n11022 & ~n11030;
  assign n12636 = n927 & n4312;
  assign n12637 = pi69  & n38376;
  assign n12638 = pi71  & n4314;
  assign n12639 = pi70  & n4322;
  assign n12640 = ~n12638 & ~n12639;
  assign n12641 = ~n12637 & ~n12639;
  assign n12642 = ~n12638 & n12641;
  assign n12643 = ~n12637 & n12640;
  assign n12644 = ~n12636 & n39739;
  assign n12645 = pi56  & ~n12644;
  assign n12646 = pi56  & ~n12645;
  assign n12647 = pi56  & n12644;
  assign n12648 = ~n12644 & ~n12645;
  assign n12649 = ~pi56  & ~n12644;
  assign n12650 = ~n39740 & ~n39741;
  assign n12651 = ~n10998 & ~n11004;
  assign n12652 = n871 & n7882;
  assign n12653 = pi66  & n39128;
  assign n12654 = pi68  & n7884;
  assign n12655 = pi67  & n7892;
  assign n12656 = ~n12654 & ~n12655;
  assign n12657 = ~n12653 & ~n12655;
  assign n12658 = ~n12654 & n12657;
  assign n12659 = ~n12653 & n12656;
  assign n12660 = ~n12652 & n39742;
  assign n12661 = pi59  & ~n12660;
  assign n12662 = pi59  & ~n12661;
  assign n12663 = pi59  & n12660;
  assign n12664 = ~n12660 & ~n12661;
  assign n12665 = ~pi59  & ~n12660;
  assign n12666 = ~n39743 & ~n39744;
  assign n12667 = pi62  & n10997;
  assign n12668 = pi61  & ~pi62 ;
  assign n12669 = ~pi61  & pi62 ;
  assign n12670 = ~pi61  & ~pi62 ;
  assign n12671 = pi61  & pi62 ;
  assign n12672 = ~n12670 & ~n12671;
  assign n12673 = ~n12668 & ~n12669;
  assign n12674 = n39429 & n39745;
  assign n12675 = n37515 & n12674;
  assign n12676 = n39429 & ~n39745;
  assign n12677 = pi65  & n12676;
  assign n12678 = pi60  & ~pi61 ;
  assign n12679 = ~pi60  & pi61 ;
  assign n12680 = ~pi60  & ~pi61 ;
  assign n12681 = pi60  & pi61 ;
  assign n12682 = ~n12680 & ~n12681;
  assign n12683 = ~n12678 & ~n12679;
  assign n12684 = ~n39429 & n39746;
  assign n12685 = pi64  & n12684;
  assign n12686 = ~n12677 & ~n12685;
  assign n12687 = ~n12675 & n12686;
  assign n12688 = n12667 & ~n12687;
  assign n12689 = ~n12667 & n12687;
  assign n12690 = pi62  & ~n10997;
  assign n12691 = pi62  & ~n12687;
  assign n12692 = pi62  & ~n12691;
  assign n12693 = ~n12687 & ~n12691;
  assign n12694 = ~n12692 & ~n12693;
  assign n12695 = n12690 & ~n12694;
  assign n12696 = n12687 & n12690;
  assign n12697 = ~n12690 & n12694;
  assign n12698 = ~n39747 & ~n12697;
  assign n12699 = ~n12688 & ~n12689;
  assign n12700 = n12666 & ~n39748;
  assign n12701 = ~n12666 & n39748;
  assign n12702 = ~n12700 & ~n12701;
  assign n12703 = ~n12651 & n12702;
  assign n12704 = n12651 & ~n12702;
  assign n12705 = ~n12703 & ~n12704;
  assign n12706 = n12650 & ~n12705;
  assign n12707 = ~n12650 & n12705;
  assign n12708 = ~n12706 & ~n12707;
  assign n12709 = ~n12635 & n12708;
  assign n12710 = n12635 & ~n12708;
  assign n12711 = ~n12709 & ~n12710;
  assign n12712 = n1218 & n1971;
  assign n12713 = pi72  & n37864;
  assign n12714 = pi74  & n1973;
  assign n12715 = pi73  & n1981;
  assign n12716 = ~n12714 & ~n12715;
  assign n12717 = ~n12713 & ~n12715;
  assign n12718 = ~n12714 & n12717;
  assign n12719 = ~n12713 & n12716;
  assign n12720 = ~n12712 & n39749;
  assign n12721 = pi53  & ~n12720;
  assign n12722 = pi53  & ~n12721;
  assign n12723 = pi53  & n12720;
  assign n12724 = ~n12720 & ~n12721;
  assign n12725 = ~pi53  & ~n12720;
  assign n12726 = ~n39750 & ~n39751;
  assign n12727 = n12711 & ~n12726;
  assign n12728 = ~n12711 & n12726;
  assign n12729 = n12711 & ~n12727;
  assign n12730 = n12711 & n12726;
  assign n12731 = ~n12726 & ~n12727;
  assign n12732 = ~n12711 & ~n12726;
  assign n12733 = ~n39752 & ~n39753;
  assign n12734 = ~n12727 & ~n12728;
  assign n12735 = n12634 & n39754;
  assign n12736 = ~n12634 & ~n39754;
  assign n12737 = ~n12735 & ~n12736;
  assign n12738 = n894 & n1596;
  assign n12739 = pi75  & n37580;
  assign n12740 = pi77  & n896;
  assign n12741 = pi76  & n904;
  assign n12742 = ~n12740 & ~n12741;
  assign n12743 = ~n12739 & ~n12741;
  assign n12744 = ~n12740 & n12743;
  assign n12745 = ~n12739 & n12742;
  assign n12746 = ~n12738 & n39755;
  assign n12747 = pi50  & ~n12746;
  assign n12748 = pi50  & ~n12747;
  assign n12749 = pi50  & n12746;
  assign n12750 = ~n12746 & ~n12747;
  assign n12751 = ~pi50  & ~n12746;
  assign n12752 = ~n39756 & ~n39757;
  assign n12753 = n12737 & ~n12752;
  assign n12754 = ~n12737 & n12752;
  assign n12755 = ~n12753 & ~n12754;
  assign n12756 = ~n12633 & ~n12754;
  assign n12757 = ~n12753 & n12756;
  assign n12758 = ~n12633 & n12755;
  assign n12759 = n12633 & ~n12755;
  assign n12760 = ~n12633 & ~n39758;
  assign n12761 = ~n12753 & ~n39758;
  assign n12762 = ~n12754 & n12761;
  assign n12763 = ~n12760 & ~n12762;
  assign n12764 = ~n39758 & ~n12759;
  assign n12765 = ~n12632 & ~n39759;
  assign n12766 = n12632 & n39759;
  assign n12767 = ~n39759 & ~n12765;
  assign n12768 = n12632 & ~n39759;
  assign n12769 = ~n12632 & ~n12765;
  assign n12770 = ~n12632 & n39759;
  assign n12771 = ~n39760 & ~n39761;
  assign n12772 = ~n12765 & ~n12766;
  assign n12773 = n12617 & n39762;
  assign n12774 = ~n12617 & ~n39762;
  assign n12775 = ~n12773 & ~n12774;
  assign n12776 = n940 & n2091;
  assign n12777 = pi81  & n37541;
  assign n12778 = pi83  & n953;
  assign n12779 = pi82  & n955;
  assign n12780 = ~n12778 & ~n12779;
  assign n12781 = ~n12777 & ~n12779;
  assign n12782 = ~n12778 & n12781;
  assign n12783 = ~n12777 & n12780;
  assign n12784 = ~n12776 & n39763;
  assign n12785 = pi44  & ~n12784;
  assign n12786 = pi44  & ~n12785;
  assign n12787 = pi44  & n12784;
  assign n12788 = ~n12784 & ~n12785;
  assign n12789 = ~pi44  & ~n12784;
  assign n12790 = ~n39764 & ~n39765;
  assign n12791 = n12775 & ~n12790;
  assign n12792 = ~n12775 & n12790;
  assign n12793 = ~n12791 & ~n12792;
  assign n12794 = ~n12616 & ~n12792;
  assign n12795 = ~n12791 & n12794;
  assign n12796 = ~n12616 & n12793;
  assign n12797 = n12616 & ~n12793;
  assign n12798 = ~n12616 & ~n39766;
  assign n12799 = ~n12791 & ~n39766;
  assign n12800 = ~n12792 & n12799;
  assign n12801 = ~n12798 & ~n12800;
  assign n12802 = ~n39766 & ~n12797;
  assign n12803 = ~n12615 & ~n39767;
  assign n12804 = n12615 & n39767;
  assign n12805 = ~n39767 & ~n12803;
  assign n12806 = n12615 & ~n39767;
  assign n12807 = ~n12615 & ~n12803;
  assign n12808 = ~n12615 & n39767;
  assign n12809 = ~n39768 & ~n39769;
  assign n12810 = ~n12803 & ~n12804;
  assign n12811 = n12600 & n39770;
  assign n12812 = ~n12600 & ~n39770;
  assign n12813 = ~n12811 & ~n12812;
  assign n12814 = n691 & n3591;
  assign n12815 = pi87  & n37503;
  assign n12816 = pi89  & n704;
  assign n12817 = pi88  & n706;
  assign n12818 = ~n12816 & ~n12817;
  assign n12819 = ~n12815 & ~n12817;
  assign n12820 = ~n12816 & n12819;
  assign n12821 = ~n12815 & n12818;
  assign n12822 = ~n12814 & n39771;
  assign n12823 = pi38  & ~n12822;
  assign n12824 = pi38  & ~n12823;
  assign n12825 = pi38  & n12822;
  assign n12826 = ~n12822 & ~n12823;
  assign n12827 = ~pi38  & ~n12822;
  assign n12828 = ~n39772 & ~n39773;
  assign n12829 = n12813 & ~n12828;
  assign n12830 = ~n12813 & n12828;
  assign n12831 = n12813 & ~n12829;
  assign n12832 = n12813 & n12828;
  assign n12833 = ~n12828 & ~n12829;
  assign n12834 = ~n12813 & ~n12828;
  assign n12835 = ~n39774 & ~n39775;
  assign n12836 = ~n12829 & ~n12830;
  assign n12837 = n12599 & n39776;
  assign n12838 = ~n12599 & ~n39776;
  assign n12839 = ~n12837 & ~n12838;
  assign n12840 = n2104 & n4453;
  assign n12841 = pi90  & n37758;
  assign n12842 = pi92  & n2117;
  assign n12843 = pi91  & n2119;
  assign n12844 = ~n12842 & ~n12843;
  assign n12845 = ~n12841 & ~n12843;
  assign n12846 = ~n12842 & n12845;
  assign n12847 = ~n12841 & n12844;
  assign n12848 = ~n12840 & n39777;
  assign n12849 = pi35  & ~n12848;
  assign n12850 = pi35  & ~n12849;
  assign n12851 = pi35  & n12848;
  assign n12852 = ~n12848 & ~n12849;
  assign n12853 = ~pi35  & ~n12848;
  assign n12854 = ~n39778 & ~n39779;
  assign n12855 = n12839 & ~n12854;
  assign n12856 = ~n12839 & n12854;
  assign n12857 = n12839 & ~n12855;
  assign n12858 = n12839 & n12854;
  assign n12859 = ~n12854 & ~n12855;
  assign n12860 = ~n12839 & ~n12854;
  assign n12861 = ~n39780 & ~n39781;
  assign n12862 = ~n12855 & ~n12856;
  assign n12863 = n12598 & n39782;
  assign n12864 = ~n12598 & ~n39782;
  assign n12865 = ~n12863 & ~n12864;
  assign n12866 = n649 & n4494;
  assign n12867 = pi93  & n37496;
  assign n12868 = pi95  & n662;
  assign n12869 = pi94  & n664;
  assign n12870 = ~n12868 & ~n12869;
  assign n12871 = ~n12867 & ~n12869;
  assign n12872 = ~n12868 & n12871;
  assign n12873 = ~n12867 & n12870;
  assign n12874 = ~n12866 & n39783;
  assign n12875 = pi32  & ~n12874;
  assign n12876 = pi32  & ~n12875;
  assign n12877 = pi32  & n12874;
  assign n12878 = ~n12874 & ~n12875;
  assign n12879 = ~pi32  & ~n12874;
  assign n12880 = ~n39784 & ~n39785;
  assign n12881 = n12865 & ~n12880;
  assign n12882 = ~n12865 & n12880;
  assign n12883 = n12865 & ~n12881;
  assign n12884 = n12865 & n12880;
  assign n12885 = ~n12880 & ~n12881;
  assign n12886 = ~n12865 & ~n12880;
  assign n12887 = ~n39786 & ~n39787;
  assign n12888 = ~n12881 & ~n12882;
  assign n12889 = ~n12597 & ~n39788;
  assign n12890 = n12597 & n39788;
  assign n12891 = ~n12597 & n39788;
  assign n12892 = n12597 & ~n39788;
  assign n12893 = ~n12891 & ~n12892;
  assign n12894 = ~n12889 & ~n12890;
  assign n12895 = ~n12596 & ~n39789;
  assign n12896 = n12596 & n39789;
  assign n12897 = ~n12895 & ~n12896;
  assign n12898 = n12581 & ~n12897;
  assign n12899 = ~n12581 & n12897;
  assign n12900 = ~n12898 & ~n12899;
  assign n12901 = n4492 & n6839;
  assign n12902 = pi99  & n38208;
  assign n12903 = pi101  & n4507;
  assign n12904 = pi100  & n4509;
  assign n12905 = ~n12903 & ~n12904;
  assign n12906 = ~n12902 & ~n12904;
  assign n12907 = ~n12903 & n12906;
  assign n12908 = ~n12902 & n12905;
  assign n12909 = ~n12901 & n39790;
  assign n12910 = pi26  & ~n12909;
  assign n12911 = pi26  & ~n12910;
  assign n12912 = pi26  & n12909;
  assign n12913 = ~n12909 & ~n12910;
  assign n12914 = ~pi26  & ~n12909;
  assign n12915 = ~n39791 & ~n39792;
  assign n12916 = n12900 & ~n12915;
  assign n12917 = ~n12900 & n12915;
  assign n12918 = n12900 & ~n12916;
  assign n12919 = n12900 & n12915;
  assign n12920 = ~n12915 & ~n12916;
  assign n12921 = ~n12900 & ~n12915;
  assign n12922 = ~n39793 & ~n39794;
  assign n12923 = ~n12916 & ~n12917;
  assign n12924 = n12580 & n39795;
  assign n12925 = ~n12580 & ~n39795;
  assign n12926 = ~n12924 & ~n12925;
  assign n12927 = n5576 & n8136;
  assign n12928 = pi102  & n38406;
  assign n12929 = pi104  & n5591;
  assign n12930 = pi103  & n5593;
  assign n12931 = ~n12929 & ~n12930;
  assign n12932 = ~n12928 & ~n12930;
  assign n12933 = ~n12929 & n12932;
  assign n12934 = ~n12928 & n12931;
  assign n12935 = ~n12927 & n39796;
  assign n12936 = pi23  & ~n12935;
  assign n12937 = pi23  & ~n12936;
  assign n12938 = pi23  & n12935;
  assign n12939 = ~n12935 & ~n12936;
  assign n12940 = ~pi23  & ~n12935;
  assign n12941 = ~n39797 & ~n39798;
  assign n12942 = n12926 & ~n12941;
  assign n12943 = ~n12926 & n12941;
  assign n12944 = n12926 & ~n12942;
  assign n12945 = n12926 & n12941;
  assign n12946 = ~n12941 & ~n12942;
  assign n12947 = ~n12926 & ~n12941;
  assign n12948 = ~n39799 & ~n39800;
  assign n12949 = ~n12942 & ~n12943;
  assign n12950 = n12579 & n39801;
  assign n12951 = ~n12579 & ~n39801;
  assign n12952 = ~n12950 & ~n12951;
  assign n12953 = n6785 & n8177;
  assign n12954 = pi105  & n38631;
  assign n12955 = pi107  & n6800;
  assign n12956 = pi106  & n6802;
  assign n12957 = ~n12955 & ~n12956;
  assign n12958 = ~n12954 & ~n12956;
  assign n12959 = ~n12955 & n12958;
  assign n12960 = ~n12954 & n12957;
  assign n12961 = ~n12953 & n39802;
  assign n12962 = pi20  & ~n12961;
  assign n12963 = pi20  & ~n12962;
  assign n12964 = pi20  & n12961;
  assign n12965 = ~n12961 & ~n12962;
  assign n12966 = ~pi20  & ~n12961;
  assign n12967 = ~n39803 & ~n39804;
  assign n12968 = n12952 & ~n12967;
  assign n12969 = ~n12952 & n12967;
  assign n12970 = ~n12968 & ~n12969;
  assign n12971 = ~n12578 & ~n12969;
  assign n12972 = ~n12968 & n12971;
  assign n12973 = ~n12578 & n12970;
  assign n12974 = n12578 & ~n12970;
  assign n12975 = ~n12578 & ~n39805;
  assign n12976 = ~n12968 & ~n39805;
  assign n12977 = ~n12969 & n12976;
  assign n12978 = ~n12975 & ~n12977;
  assign n12979 = ~n39805 & ~n12974;
  assign n12980 = n12577 & n39806;
  assign n12981 = ~n12577 & ~n39806;
  assign n12982 = ~n12980 & ~n12981;
  assign n12983 = ~n12562 & n12982;
  assign n12984 = n12562 & ~n12982;
  assign n12985 = ~n12983 & ~n12984;
  assign n12986 = n12561 & ~n12985;
  assign n12987 = ~n12561 & n12985;
  assign n12988 = ~n12986 & ~n12987;
  assign n12989 = ~n12546 & n12988;
  assign n12990 = n12546 & ~n12988;
  assign n12991 = ~n12989 & ~n12990;
  assign n12992 = n12545 & ~n12991;
  assign n12993 = ~n12545 & n12991;
  assign n12994 = ~n12992 & ~n12993;
  assign n12995 = ~n12523 & n12994;
  assign n12996 = n12523 & ~n12994;
  assign n12997 = ~n12995 & ~n12996;
  assign n12998 = pi5  & ~pi6 ;
  assign n12999 = ~pi5  & pi6 ;
  assign n13000 = ~pi5  & ~pi6 ;
  assign n13001 = pi5  & pi6 ;
  assign n13002 = ~n13000 & ~n13001;
  assign n13003 = ~n12998 & ~n12999;
  assign n13004 = pi7  & ~pi8 ;
  assign n13005 = ~pi7  & pi8 ;
  assign n13006 = ~pi7  & ~pi8 ;
  assign n13007 = pi7  & pi8 ;
  assign n13008 = ~n13006 & ~n13007;
  assign n13009 = ~n13004 & ~n13005;
  assign n13010 = n39807 & n39808;
  assign n13011 = pi117  & pi118 ;
  assign n13012 = pi116  & pi117 ;
  assign n13013 = ~n12526 & ~n12528;
  assign n13014 = ~pi116  & ~pi117 ;
  assign n13015 = ~n13012 & ~n13014;
  assign n13016 = ~n13013 & n13015;
  assign n13017 = ~n13012 & ~n13016;
  assign n13018 = ~pi117  & ~pi118 ;
  assign n13019 = ~n13011 & ~n13018;
  assign n13020 = ~n13017 & n13019;
  assign n13021 = ~n13011 & ~n13020;
  assign n13022 = ~pi118  & ~pi119 ;
  assign n13023 = pi118  & pi119 ;
  assign n13024 = ~n13022 & ~n13023;
  assign n13025 = ~n13021 & n13024;
  assign n13026 = n13021 & ~n13024;
  assign n13027 = ~n13025 & ~n13026;
  assign n13028 = n13010 & n13027;
  assign n13029 = pi6  & ~pi7 ;
  assign n13030 = ~pi6  & pi7 ;
  assign n13031 = ~pi6  & ~pi7 ;
  assign n13032 = pi6  & pi7 ;
  assign n13033 = ~n13031 & ~n13032;
  assign n13034 = ~n13029 & ~n13030;
  assign n13035 = ~n39807 & n39808;
  assign n13036 = ~n39807 & ~n39809;
  assign n13037 = n39808 & n13036;
  assign n13038 = ~n39809 & n13035;
  assign n13039 = pi117  & n39810;
  assign n13040 = n39807 & ~n39808;
  assign n13041 = pi119  & n13040;
  assign n13042 = ~n39807 & n39809;
  assign n13043 = pi118  & n13042;
  assign n13044 = ~n13041 & ~n13043;
  assign n13045 = ~n13039 & ~n13043;
  assign n13046 = ~n13041 & n13045;
  assign n13047 = ~n13039 & n13044;
  assign n13048 = ~n13028 & n39811;
  assign n13049 = pi8  & ~n13048;
  assign n13050 = pi8  & ~n13049;
  assign n13051 = pi8  & n13048;
  assign n13052 = ~n13048 & ~n13049;
  assign n13053 = ~pi8  & ~n13048;
  assign n13054 = ~n39812 & ~n39813;
  assign n13055 = n12997 & ~n13054;
  assign n13056 = n13017 & ~n13019;
  assign n13057 = ~n13020 & ~n13056;
  assign n13058 = n13010 & n13057;
  assign n13059 = pi116  & n39810;
  assign n13060 = pi118  & n13040;
  assign n13061 = pi117  & n13042;
  assign n13062 = ~n13060 & ~n13061;
  assign n13063 = ~n13059 & ~n13061;
  assign n13064 = ~n13060 & n13063;
  assign n13065 = ~n13059 & n13062;
  assign n13066 = ~n13058 & n39814;
  assign n13067 = pi8  & ~n13066;
  assign n13068 = pi8  & ~n13067;
  assign n13069 = pi8  & n13066;
  assign n13070 = ~n13066 & ~n13067;
  assign n13071 = ~pi8  & ~n13066;
  assign n13072 = ~n39815 & ~n39816;
  assign n13073 = n12514 & ~n39719;
  assign n13074 = ~n39718 & n13073;
  assign n13075 = n12514 & n39720;
  assign n13076 = ~n12522 & ~n39817;
  assign n13077 = ~n13072 & n13076;
  assign n13078 = n13013 & ~n13015;
  assign n13079 = ~n13016 & ~n13078;
  assign n13080 = n13010 & n13079;
  assign n13081 = pi115  & n39810;
  assign n13082 = pi117  & n13040;
  assign n13083 = pi116  & n13042;
  assign n13084 = ~n13082 & ~n13083;
  assign n13085 = ~n13081 & ~n13083;
  assign n13086 = ~n13082 & n13085;
  assign n13087 = ~n13081 & n13084;
  assign n13088 = ~n13080 & n39818;
  assign n13089 = pi8  & ~n13088;
  assign n13090 = pi8  & ~n13089;
  assign n13091 = pi8  & n13088;
  assign n13092 = ~n13088 & ~n13089;
  assign n13093 = ~pi8  & ~n13088;
  assign n13094 = ~n39819 & ~n39820;
  assign n13095 = n12505 & n39717;
  assign n13096 = ~n12513 & ~n13095;
  assign n13097 = ~n13094 & n13096;
  assign n13098 = n12530 & n13010;
  assign n13099 = pi114  & n39810;
  assign n13100 = pi116  & n13040;
  assign n13101 = pi115  & n13042;
  assign n13102 = ~n13100 & ~n13101;
  assign n13103 = ~n13099 & ~n13101;
  assign n13104 = ~n13100 & n13103;
  assign n13105 = ~n13099 & n13102;
  assign n13106 = ~n13098 & n39821;
  assign n13107 = pi8  & ~n13106;
  assign n13108 = pi8  & ~n13107;
  assign n13109 = pi8  & n13106;
  assign n13110 = ~n13106 & ~n13107;
  assign n13111 = ~pi8  & ~n13106;
  assign n13112 = ~n39822 & ~n39823;
  assign n13113 = n12501 & ~n12503;
  assign n13114 = ~n12504 & ~n13113;
  assign n13115 = ~n13112 & n13114;
  assign n13116 = n523 & n13010;
  assign n13117 = pi113  & n39810;
  assign n13118 = pi115  & n13040;
  assign n13119 = pi114  & n13042;
  assign n13120 = ~n13118 & ~n13119;
  assign n13121 = ~n13117 & ~n13119;
  assign n13122 = ~n13118 & n13121;
  assign n13123 = ~n13117 & n13120;
  assign n13124 = ~n13116 & n39824;
  assign n13125 = pi8  & ~n13124;
  assign n13126 = pi8  & ~n13125;
  assign n13127 = pi8  & n13124;
  assign n13128 = ~n13124 & ~n13125;
  assign n13129 = ~pi8  & ~n13124;
  assign n13130 = ~n39825 & ~n39826;
  assign n13131 = n12492 & ~n39713;
  assign n13132 = ~n39712 & n13131;
  assign n13133 = n12492 & n39714;
  assign n13134 = ~n12500 & ~n39827;
  assign n13135 = ~n13130 & n13134;
  assign n13136 = n11258 & n13010;
  assign n13137 = pi112  & n39810;
  assign n13138 = pi114  & n13040;
  assign n13139 = pi113  & n13042;
  assign n13140 = ~n13138 & ~n13139;
  assign n13141 = ~n13137 & ~n13139;
  assign n13142 = ~n13138 & n13141;
  assign n13143 = ~n13137 & n13140;
  assign n13144 = ~n13136 & n39828;
  assign n13145 = pi8  & ~n13144;
  assign n13146 = pi8  & ~n13145;
  assign n13147 = pi8  & n13144;
  assign n13148 = ~n13144 & ~n13145;
  assign n13149 = ~pi8  & ~n13144;
  assign n13150 = ~n39829 & ~n39830;
  assign n13151 = n12483 & n39711;
  assign n13152 = ~n12491 & ~n13151;
  assign n13153 = ~n13150 & n13152;
  assign n13154 = n11276 & n13010;
  assign n13155 = pi111  & n39810;
  assign n13156 = pi113  & n13040;
  assign n13157 = pi112  & n13042;
  assign n13158 = ~n13156 & ~n13157;
  assign n13159 = ~n13155 & ~n13157;
  assign n13160 = ~n13156 & n13159;
  assign n13161 = ~n13155 & n13158;
  assign n13162 = ~n13154 & n39831;
  assign n13163 = pi8  & ~n13162;
  assign n13164 = pi8  & ~n13163;
  assign n13165 = pi8  & n13162;
  assign n13166 = ~n13162 & ~n13163;
  assign n13167 = ~pi8  & ~n13162;
  assign n13168 = ~n39832 & ~n39833;
  assign n13169 = n12479 & ~n12481;
  assign n13170 = ~n12482 & ~n13169;
  assign n13171 = ~n13168 & n13170;
  assign n13172 = n10844 & n13010;
  assign n13173 = pi110  & n39810;
  assign n13174 = pi112  & n13040;
  assign n13175 = pi111  & n13042;
  assign n13176 = ~n13174 & ~n13175;
  assign n13177 = ~n13173 & ~n13175;
  assign n13178 = ~n13174 & n13177;
  assign n13179 = ~n13173 & n13176;
  assign n13180 = ~n13172 & n39834;
  assign n13181 = pi8  & ~n13180;
  assign n13182 = pi8  & ~n13181;
  assign n13183 = pi8  & n13180;
  assign n13184 = ~n13180 & ~n13181;
  assign n13185 = ~pi8  & ~n13180;
  assign n13186 = ~n39835 & ~n39836;
  assign n13187 = n12470 & n39708;
  assign n13188 = ~n12470 & ~n12478;
  assign n13189 = ~n39708 & ~n12478;
  assign n13190 = ~n13188 & ~n13189;
  assign n13191 = ~n12478 & ~n13187;
  assign n13192 = ~n13186 & ~n39837;
  assign n13193 = n565 & n13010;
  assign n13194 = pi109  & n39810;
  assign n13195 = pi111  & n13040;
  assign n13196 = pi110  & n13042;
  assign n13197 = ~n13195 & ~n13196;
  assign n13198 = ~n13194 & ~n13196;
  assign n13199 = ~n13195 & n13198;
  assign n13200 = ~n13194 & n13197;
  assign n13201 = ~n13193 & n39838;
  assign n13202 = pi8  & ~n13201;
  assign n13203 = pi8  & ~n13202;
  assign n13204 = pi8  & n13201;
  assign n13205 = ~n13201 & ~n13202;
  assign n13206 = ~pi8  & ~n13201;
  assign n13207 = ~n39839 & ~n39840;
  assign n13208 = n12464 & ~n12466;
  assign n13209 = ~n12464 & ~n39705;
  assign n13210 = ~n12465 & n12470;
  assign n13211 = ~n13209 & ~n13210;
  assign n13212 = ~n39705 & ~n13208;
  assign n13213 = ~n13207 & ~n39841;
  assign n13214 = n9678 & n13010;
  assign n13215 = pi108  & n39810;
  assign n13216 = pi110  & n13040;
  assign n13217 = pi109  & n13042;
  assign n13218 = ~n13216 & ~n13217;
  assign n13219 = ~n13215 & ~n13217;
  assign n13220 = ~n13216 & n13219;
  assign n13221 = ~n13215 & n13218;
  assign n13222 = ~n13214 & n39842;
  assign n13223 = pi8  & ~n13222;
  assign n13224 = pi8  & ~n13223;
  assign n13225 = pi8  & n13222;
  assign n13226 = ~n13222 & ~n13223;
  assign n13227 = ~pi8  & ~n13222;
  assign n13228 = ~n39843 & ~n39844;
  assign n13229 = n12458 & ~n12460;
  assign n13230 = ~n12458 & ~n39704;
  assign n13231 = ~n12459 & n12464;
  assign n13232 = ~n13230 & ~n13231;
  assign n13233 = ~n39704 & ~n13229;
  assign n13234 = ~n13228 & ~n39845;
  assign n13235 = ~n11430 & n12456;
  assign n13236 = ~n12457 & ~n13235;
  assign n13237 = n9701 & n13010;
  assign n13238 = pi107  & n39810;
  assign n13239 = pi109  & n13040;
  assign n13240 = pi108  & n13042;
  assign n13241 = ~n13239 & ~n13240;
  assign n13242 = ~n13238 & ~n13240;
  assign n13243 = ~n13239 & n13242;
  assign n13244 = ~n13238 & n13241;
  assign n13245 = ~n13237 & n39846;
  assign n13246 = pi8  & ~n13245;
  assign n13247 = pi8  & ~n13246;
  assign n13248 = pi8  & n13245;
  assign n13249 = ~n13245 & ~n13246;
  assign n13250 = ~pi8  & ~n13245;
  assign n13251 = ~n39847 & ~n39848;
  assign n13252 = n13236 & ~n13251;
  assign n13253 = n12447 & n39703;
  assign n13254 = ~n12455 & ~n13253;
  assign n13255 = n9277 & n13010;
  assign n13256 = pi106  & n39810;
  assign n13257 = pi108  & n13040;
  assign n13258 = pi107  & n13042;
  assign n13259 = ~n13257 & ~n13258;
  assign n13260 = ~n13256 & ~n13258;
  assign n13261 = ~n13257 & n13260;
  assign n13262 = ~n13256 & n13259;
  assign n13263 = ~n13255 & n39849;
  assign n13264 = pi8  & ~n13263;
  assign n13265 = pi8  & ~n13264;
  assign n13266 = pi8  & n13263;
  assign n13267 = ~n13263 & ~n13264;
  assign n13268 = ~pi8  & ~n13263;
  assign n13269 = ~n39850 & ~n39851;
  assign n13270 = n13254 & ~n13269;
  assign n13271 = n12438 & n39700;
  assign n13272 = ~n12446 & ~n13271;
  assign n13273 = n8177 & n13010;
  assign n13274 = pi105  & n39810;
  assign n13275 = pi107  & n13040;
  assign n13276 = pi106  & n13042;
  assign n13277 = ~n13275 & ~n13276;
  assign n13278 = ~n13274 & ~n13276;
  assign n13279 = ~n13275 & n13278;
  assign n13280 = ~n13274 & n13277;
  assign n13281 = ~n13273 & n39852;
  assign n13282 = pi8  & ~n13281;
  assign n13283 = pi8  & ~n13282;
  assign n13284 = pi8  & n13281;
  assign n13285 = ~n13281 & ~n13282;
  assign n13286 = ~pi8  & ~n13281;
  assign n13287 = ~n39853 & ~n39854;
  assign n13288 = n13272 & ~n13287;
  assign n13289 = n12429 & n39697;
  assign n13290 = ~n12437 & ~n13289;
  assign n13291 = n8209 & n13010;
  assign n13292 = pi104  & n39810;
  assign n13293 = pi106  & n13040;
  assign n13294 = pi105  & n13042;
  assign n13295 = ~n13293 & ~n13294;
  assign n13296 = ~n13292 & ~n13294;
  assign n13297 = ~n13293 & n13296;
  assign n13298 = ~n13292 & n13295;
  assign n13299 = ~n13291 & n39855;
  assign n13300 = pi8  & ~n13299;
  assign n13301 = pi8  & ~n13300;
  assign n13302 = pi8  & n13299;
  assign n13303 = ~n13299 & ~n13300;
  assign n13304 = ~pi8  & ~n13299;
  assign n13305 = ~n39856 & ~n39857;
  assign n13306 = n13290 & ~n13305;
  assign n13307 = n12420 & n39694;
  assign n13308 = ~n12428 & ~n13307;
  assign n13309 = n8229 & n13010;
  assign n13310 = pi103  & n39810;
  assign n13311 = pi105  & n13040;
  assign n13312 = pi104  & n13042;
  assign n13313 = ~n13311 & ~n13312;
  assign n13314 = ~n13310 & ~n13312;
  assign n13315 = ~n13311 & n13314;
  assign n13316 = ~n13310 & n13313;
  assign n13317 = ~n13309 & n39858;
  assign n13318 = pi8  & ~n13317;
  assign n13319 = pi8  & ~n13318;
  assign n13320 = pi8  & n13317;
  assign n13321 = ~n13317 & ~n13318;
  assign n13322 = ~pi8  & ~n13317;
  assign n13323 = ~n39859 & ~n39860;
  assign n13324 = n13308 & ~n13323;
  assign n13325 = n12411 & n39691;
  assign n13326 = ~n12419 & ~n13325;
  assign n13327 = n8136 & n13010;
  assign n13328 = pi102  & n39810;
  assign n13329 = pi104  & n13040;
  assign n13330 = pi103  & n13042;
  assign n13331 = ~n13329 & ~n13330;
  assign n13332 = ~n13328 & ~n13330;
  assign n13333 = ~n13329 & n13332;
  assign n13334 = ~n13328 & n13331;
  assign n13335 = ~n13327 & n39861;
  assign n13336 = pi8  & ~n13335;
  assign n13337 = pi8  & ~n13336;
  assign n13338 = pi8  & n13335;
  assign n13339 = ~n13335 & ~n13336;
  assign n13340 = ~pi8  & ~n13335;
  assign n13341 = ~n39862 & ~n39863;
  assign n13342 = n13326 & ~n13341;
  assign n13343 = n12407 & ~n12409;
  assign n13344 = ~n12410 & ~n13343;
  assign n13345 = n6787 & n13010;
  assign n13346 = pi101  & n39810;
  assign n13347 = pi103  & n13040;
  assign n13348 = pi102  & n13042;
  assign n13349 = ~n13347 & ~n13348;
  assign n13350 = ~n13346 & ~n13348;
  assign n13351 = ~n13347 & n13350;
  assign n13352 = ~n13346 & n13349;
  assign n13353 = ~n13345 & n39864;
  assign n13354 = pi8  & ~n13353;
  assign n13355 = pi8  & ~n13354;
  assign n13356 = pi8  & n13353;
  assign n13357 = ~n13353 & ~n13354;
  assign n13358 = ~pi8  & ~n13353;
  assign n13359 = ~n39865 & ~n39866;
  assign n13360 = n13344 & ~n13359;
  assign n13361 = n12398 & n39688;
  assign n13362 = ~n12406 & ~n13361;
  assign n13363 = n6819 & n13010;
  assign n13364 = pi100  & n39810;
  assign n13365 = pi102  & n13040;
  assign n13366 = pi101  & n13042;
  assign n13367 = ~n13365 & ~n13366;
  assign n13368 = ~n13364 & ~n13366;
  assign n13369 = ~n13365 & n13368;
  assign n13370 = ~n13364 & n13367;
  assign n13371 = ~n13363 & n39867;
  assign n13372 = pi8  & ~n13371;
  assign n13373 = pi8  & ~n13372;
  assign n13374 = pi8  & n13371;
  assign n13375 = ~n13371 & ~n13372;
  assign n13376 = ~pi8  & ~n13371;
  assign n13377 = ~n39868 & ~n39869;
  assign n13378 = n13362 & ~n13377;
  assign n13379 = n12389 & n39685;
  assign n13380 = ~n12397 & ~n13379;
  assign n13381 = n6839 & n13010;
  assign n13382 = pi99  & n39810;
  assign n13383 = pi101  & n13040;
  assign n13384 = pi100  & n13042;
  assign n13385 = ~n13383 & ~n13384;
  assign n13386 = ~n13382 & ~n13384;
  assign n13387 = ~n13383 & n13386;
  assign n13388 = ~n13382 & n13385;
  assign n13389 = ~n13381 & n39870;
  assign n13390 = pi8  & ~n13389;
  assign n13391 = pi8  & ~n13390;
  assign n13392 = pi8  & n13389;
  assign n13393 = ~n13389 & ~n13390;
  assign n13394 = ~pi8  & ~n13389;
  assign n13395 = ~n39871 & ~n39872;
  assign n13396 = n13380 & ~n13395;
  assign n13397 = n6474 & n13010;
  assign n13398 = pi98  & n39810;
  assign n13399 = pi100  & n13040;
  assign n13400 = pi99  & n13042;
  assign n13401 = ~n13399 & ~n13400;
  assign n13402 = ~n13398 & ~n13400;
  assign n13403 = ~n13399 & n13402;
  assign n13404 = ~n13398 & n13401;
  assign n13405 = ~n13397 & n39873;
  assign n13406 = pi8  & ~n13405;
  assign n13407 = pi8  & ~n13406;
  assign n13408 = pi8  & n13405;
  assign n13409 = ~n13405 & ~n13406;
  assign n13410 = ~pi8  & ~n13405;
  assign n13411 = ~n39874 & ~n39875;
  assign n13412 = n12380 & n39682;
  assign n13413 = ~n12380 & n39682;
  assign n13414 = n12380 & ~n39682;
  assign n13415 = ~n13413 & ~n13414;
  assign n13416 = ~n12388 & ~n13412;
  assign n13417 = ~n13411 & ~n39876;
  assign n13418 = n12376 & ~n12378;
  assign n13419 = ~n12379 & ~n13418;
  assign n13420 = n5578 & n13010;
  assign n13421 = pi97  & n39810;
  assign n13422 = pi99  & n13040;
  assign n13423 = pi98  & n13042;
  assign n13424 = ~n13422 & ~n13423;
  assign n13425 = ~n13421 & ~n13423;
  assign n13426 = ~n13422 & n13425;
  assign n13427 = ~n13421 & n13424;
  assign n13428 = ~n13420 & n39877;
  assign n13429 = pi8  & ~n13428;
  assign n13430 = pi8  & ~n13429;
  assign n13431 = pi8  & n13428;
  assign n13432 = ~n13428 & ~n13429;
  assign n13433 = ~pi8  & ~n13428;
  assign n13434 = ~n39878 & ~n39879;
  assign n13435 = n13419 & ~n13434;
  assign n13436 = n5610 & n13010;
  assign n13437 = pi96  & n39810;
  assign n13438 = pi98  & n13040;
  assign n13439 = pi97  & n13042;
  assign n13440 = ~n13438 & ~n13439;
  assign n13441 = ~n13437 & ~n13439;
  assign n13442 = ~n13438 & n13441;
  assign n13443 = ~n13437 & n13440;
  assign n13444 = ~n13436 & n39880;
  assign n13445 = pi8  & ~n13444;
  assign n13446 = pi8  & ~n13445;
  assign n13447 = pi8  & n13444;
  assign n13448 = ~n13444 & ~n13445;
  assign n13449 = ~pi8  & ~n13444;
  assign n13450 = ~n39881 & ~n39882;
  assign n13451 = n12372 & ~n12374;
  assign n13452 = ~n12375 & ~n13451;
  assign n13453 = ~n13450 & n13452;
  assign n13454 = n12368 & ~n12370;
  assign n13455 = ~n12371 & ~n13454;
  assign n13456 = n5630 & n13010;
  assign n13457 = pi95  & n39810;
  assign n13458 = pi97  & n13040;
  assign n13459 = pi96  & n13042;
  assign n13460 = ~n13458 & ~n13459;
  assign n13461 = ~n13457 & ~n13459;
  assign n13462 = ~n13458 & n13461;
  assign n13463 = ~n13457 & n13460;
  assign n13464 = ~n13456 & n39883;
  assign n13465 = pi8  & ~n13464;
  assign n13466 = pi8  & ~n13465;
  assign n13467 = pi8  & n13464;
  assign n13468 = ~n13464 & ~n13465;
  assign n13469 = ~pi8  & ~n13464;
  assign n13470 = ~n39884 & ~n39885;
  assign n13471 = n13455 & ~n13470;
  assign n13472 = n5281 & n13010;
  assign n13473 = pi94  & n39810;
  assign n13474 = pi96  & n13040;
  assign n13475 = pi95  & n13042;
  assign n13476 = ~n13474 & ~n13475;
  assign n13477 = ~n13473 & ~n13475;
  assign n13478 = ~n13474 & n13477;
  assign n13479 = ~n13473 & n13476;
  assign n13480 = ~n13472 & n39886;
  assign n13481 = pi8  & ~n13480;
  assign n13482 = pi8  & ~n13481;
  assign n13483 = pi8  & n13480;
  assign n13484 = ~n13480 & ~n13481;
  assign n13485 = ~pi8  & ~n13480;
  assign n13486 = ~n39887 & ~n39888;
  assign n13487 = n12364 & ~n12366;
  assign n13488 = ~n12367 & ~n13487;
  assign n13489 = ~n13486 & n13488;
  assign n13490 = n4494 & n13010;
  assign n13491 = pi93  & n39810;
  assign n13492 = pi95  & n13040;
  assign n13493 = pi94  & n13042;
  assign n13494 = ~n13492 & ~n13493;
  assign n13495 = ~n13491 & ~n13493;
  assign n13496 = ~n13492 & n13495;
  assign n13497 = ~n13491 & n13494;
  assign n13498 = ~n13490 & n39889;
  assign n13499 = pi8  & ~n13498;
  assign n13500 = pi8  & ~n13499;
  assign n13501 = pi8  & n13498;
  assign n13502 = ~n13498 & ~n13499;
  assign n13503 = ~pi8  & ~n13498;
  assign n13504 = ~n39890 & ~n39891;
  assign n13505 = n12360 & ~n12362;
  assign n13506 = ~n12363 & ~n13505;
  assign n13507 = ~n13504 & n13506;
  assign n13508 = n4524 & n13010;
  assign n13509 = pi92  & n39810;
  assign n13510 = pi94  & n13040;
  assign n13511 = pi93  & n13042;
  assign n13512 = ~n13510 & ~n13511;
  assign n13513 = ~n13509 & ~n13511;
  assign n13514 = ~n13510 & n13513;
  assign n13515 = ~n13509 & n13512;
  assign n13516 = ~n13508 & n39892;
  assign n13517 = pi8  & ~n13516;
  assign n13518 = pi8  & ~n13517;
  assign n13519 = pi8  & n13516;
  assign n13520 = ~n13516 & ~n13517;
  assign n13521 = ~pi8  & ~n13516;
  assign n13522 = ~n39893 & ~n39894;
  assign n13523 = n12351 & n39679;
  assign n13524 = ~n12351 & n39679;
  assign n13525 = n12351 & ~n39679;
  assign n13526 = ~n13524 & ~n13525;
  assign n13527 = ~n12359 & ~n13523;
  assign n13528 = ~n13522 & ~n39895;
  assign n13529 = n12347 & ~n12349;
  assign n13530 = ~n12350 & ~n13529;
  assign n13531 = n4544 & n13010;
  assign n13532 = pi91  & n39810;
  assign n13533 = pi93  & n13040;
  assign n13534 = pi92  & n13042;
  assign n13535 = ~n13533 & ~n13534;
  assign n13536 = ~n13532 & ~n13534;
  assign n13537 = ~n13533 & n13536;
  assign n13538 = ~n13532 & n13535;
  assign n13539 = ~n13531 & n39896;
  assign n13540 = pi8  & ~n13539;
  assign n13541 = pi8  & ~n13540;
  assign n13542 = pi8  & n13539;
  assign n13543 = ~n13539 & ~n13540;
  assign n13544 = ~pi8  & ~n13539;
  assign n13545 = ~n39897 & ~n39898;
  assign n13546 = n13530 & ~n13545;
  assign n13547 = n4453 & n13010;
  assign n13548 = pi90  & n39810;
  assign n13549 = pi92  & n13040;
  assign n13550 = pi91  & n13042;
  assign n13551 = ~n13549 & ~n13550;
  assign n13552 = ~n13548 & ~n13550;
  assign n13553 = ~n13549 & n13552;
  assign n13554 = ~n13548 & n13551;
  assign n13555 = ~n13547 & n39899;
  assign n13556 = pi8  & ~n13555;
  assign n13557 = pi8  & ~n13556;
  assign n13558 = pi8  & n13555;
  assign n13559 = ~n13555 & ~n13556;
  assign n13560 = ~pi8  & ~n13555;
  assign n13561 = ~n39900 & ~n39901;
  assign n13562 = n12341 & ~n12343;
  assign n13563 = ~n12341 & ~n39676;
  assign n13564 = ~n12342 & n12347;
  assign n13565 = ~n13563 & ~n13564;
  assign n13566 = ~n39676 & ~n13562;
  assign n13567 = ~n13561 & ~n39902;
  assign n13568 = n12337 & ~n12339;
  assign n13569 = ~n12340 & ~n13568;
  assign n13570 = n594 & n13010;
  assign n13571 = pi89  & n39810;
  assign n13572 = pi91  & n13040;
  assign n13573 = pi90  & n13042;
  assign n13574 = ~n13572 & ~n13573;
  assign n13575 = ~n13571 & ~n13573;
  assign n13576 = ~n13572 & n13575;
  assign n13577 = ~n13571 & n13574;
  assign n13578 = ~n13570 & n39903;
  assign n13579 = pi8  & ~n13578;
  assign n13580 = pi8  & ~n13579;
  assign n13581 = pi8  & n13578;
  assign n13582 = ~n13578 & ~n13579;
  assign n13583 = ~pi8  & ~n13578;
  assign n13584 = ~n39904 & ~n39905;
  assign n13585 = n13569 & ~n13584;
  assign n13586 = n12333 & ~n12335;
  assign n13587 = ~n12336 & ~n13586;
  assign n13588 = n3566 & n13010;
  assign n13589 = pi88  & n39810;
  assign n13590 = pi90  & n13040;
  assign n13591 = pi89  & n13042;
  assign n13592 = ~n13590 & ~n13591;
  assign n13593 = ~n13589 & ~n13591;
  assign n13594 = ~n13590 & n13593;
  assign n13595 = ~n13589 & n13592;
  assign n13596 = ~n13588 & n39906;
  assign n13597 = pi8  & ~n13596;
  assign n13598 = pi8  & ~n13597;
  assign n13599 = pi8  & n13596;
  assign n13600 = ~n13596 & ~n13597;
  assign n13601 = ~pi8  & ~n13596;
  assign n13602 = ~n39907 & ~n39908;
  assign n13603 = n13587 & ~n13602;
  assign n13604 = n12324 & n39675;
  assign n13605 = ~n12332 & ~n13604;
  assign n13606 = n3591 & n13010;
  assign n13607 = pi87  & n39810;
  assign n13608 = pi89  & n13040;
  assign n13609 = pi88  & n13042;
  assign n13610 = ~n13608 & ~n13609;
  assign n13611 = ~n13607 & ~n13609;
  assign n13612 = ~n13608 & n13611;
  assign n13613 = ~n13607 & n13610;
  assign n13614 = ~n13606 & n39909;
  assign n13615 = pi8  & ~n13614;
  assign n13616 = pi8  & ~n13615;
  assign n13617 = pi8  & n13614;
  assign n13618 = ~n13614 & ~n13615;
  assign n13619 = ~pi8  & ~n13614;
  assign n13620 = ~n39910 & ~n39911;
  assign n13621 = n13605 & ~n13620;
  assign n13622 = n3354 & n13010;
  assign n13623 = pi86  & n39810;
  assign n13624 = pi88  & n13040;
  assign n13625 = pi87  & n13042;
  assign n13626 = ~n13624 & ~n13625;
  assign n13627 = ~n13623 & ~n13625;
  assign n13628 = ~n13624 & n13627;
  assign n13629 = ~n13623 & n13626;
  assign n13630 = ~n13622 & n39912;
  assign n13631 = pi8  & ~n13630;
  assign n13632 = pi8  & ~n13631;
  assign n13633 = pi8  & n13630;
  assign n13634 = ~n13630 & ~n13631;
  assign n13635 = ~pi8  & ~n13630;
  assign n13636 = ~n39913 & ~n39914;
  assign n13637 = n12315 & n39672;
  assign n13638 = ~n12315 & n39672;
  assign n13639 = n12315 & ~n39672;
  assign n13640 = ~n13638 & ~n13639;
  assign n13641 = ~n12323 & ~n13637;
  assign n13642 = ~n13636 & ~n39915;
  assign n13643 = n636 & n13010;
  assign n13644 = pi85  & n39810;
  assign n13645 = pi87  & n13040;
  assign n13646 = pi86  & n13042;
  assign n13647 = ~n13645 & ~n13646;
  assign n13648 = ~n13644 & ~n13646;
  assign n13649 = ~n13645 & n13648;
  assign n13650 = ~n13644 & n13647;
  assign n13651 = ~n13643 & n39916;
  assign n13652 = pi8  & ~n13651;
  assign n13653 = pi8  & ~n13652;
  assign n13654 = pi8  & n13651;
  assign n13655 = ~n13651 & ~n13652;
  assign n13656 = ~pi8  & ~n13651;
  assign n13657 = ~n39917 & ~n39918;
  assign n13658 = n12309 & ~n12311;
  assign n13659 = ~n12309 & ~n39669;
  assign n13660 = ~n12310 & n12315;
  assign n13661 = ~n13659 & ~n13660;
  assign n13662 = ~n39669 & ~n13658;
  assign n13663 = ~n13657 & ~n39919;
  assign n13664 = n12300 & n39668;
  assign n13665 = ~n12308 & ~n13664;
  assign n13666 = n2779 & n13010;
  assign n13667 = pi84  & n39810;
  assign n13668 = pi86  & n13040;
  assign n13669 = pi85  & n13042;
  assign n13670 = ~n13668 & ~n13669;
  assign n13671 = ~n13667 & ~n13669;
  assign n13672 = ~n13668 & n13671;
  assign n13673 = ~n13667 & n13670;
  assign n13674 = ~n13666 & n39920;
  assign n13675 = pi8  & ~n13674;
  assign n13676 = pi8  & ~n13675;
  assign n13677 = pi8  & n13674;
  assign n13678 = ~n13674 & ~n13675;
  assign n13679 = ~pi8  & ~n13674;
  assign n13680 = ~n39921 & ~n39922;
  assign n13681 = n13665 & ~n13680;
  assign n13682 = ~n13665 & n13680;
  assign n13683 = ~n13681 & ~n13682;
  assign n13684 = n12291 & n39665;
  assign n13685 = ~n12299 & ~n13684;
  assign n13686 = n2804 & n13010;
  assign n13687 = pi83  & n39810;
  assign n13688 = pi85  & n13040;
  assign n13689 = pi84  & n13042;
  assign n13690 = ~n13688 & ~n13689;
  assign n13691 = ~n13687 & ~n13689;
  assign n13692 = ~n13688 & n13691;
  assign n13693 = ~n13687 & n13690;
  assign n13694 = ~n13686 & n39923;
  assign n13695 = pi8  & ~n13694;
  assign n13696 = pi8  & ~n13695;
  assign n13697 = pi8  & n13694;
  assign n13698 = ~n13694 & ~n13695;
  assign n13699 = ~pi8  & ~n13694;
  assign n13700 = ~n39924 & ~n39925;
  assign n13701 = n13685 & ~n13700;
  assign n13702 = ~n13685 & n13700;
  assign n13703 = ~n13701 & ~n13702;
  assign n13704 = n12287 & ~n12289;
  assign n13705 = ~n12290 & ~n13704;
  assign n13706 = n2591 & n13010;
  assign n13707 = pi82  & n39810;
  assign n13708 = pi84  & n13040;
  assign n13709 = pi83  & n13042;
  assign n13710 = ~n13708 & ~n13709;
  assign n13711 = ~n13707 & ~n13709;
  assign n13712 = ~n13708 & n13711;
  assign n13713 = ~n13707 & n13710;
  assign n13714 = ~n13706 & n39926;
  assign n13715 = pi8  & ~n13714;
  assign n13716 = pi8  & ~n13715;
  assign n13717 = pi8  & n13714;
  assign n13718 = ~n13714 & ~n13715;
  assign n13719 = ~pi8  & ~n13714;
  assign n13720 = ~n39927 & ~n39928;
  assign n13721 = n13705 & ~n13720;
  assign n13722 = n12278 & n39662;
  assign n13723 = ~n12286 & ~n13722;
  assign n13724 = n2091 & n13010;
  assign n13725 = pi81  & n39810;
  assign n13726 = pi83  & n13040;
  assign n13727 = pi82  & n13042;
  assign n13728 = ~n13726 & ~n13727;
  assign n13729 = ~n13725 & ~n13727;
  assign n13730 = ~n13726 & n13729;
  assign n13731 = ~n13725 & n13728;
  assign n13732 = ~n13724 & n39929;
  assign n13733 = pi8  & ~n13732;
  assign n13734 = pi8  & ~n13733;
  assign n13735 = pi8  & n13732;
  assign n13736 = ~n13732 & ~n13733;
  assign n13737 = ~pi8  & ~n13732;
  assign n13738 = ~n39930 & ~n39931;
  assign n13739 = n13723 & ~n13738;
  assign n13740 = n12269 & n39659;
  assign n13741 = ~n12277 & ~n13740;
  assign n13742 = n2134 & n13010;
  assign n13743 = pi80  & n39810;
  assign n13744 = pi82  & n13040;
  assign n13745 = pi81  & n13042;
  assign n13746 = ~n13744 & ~n13745;
  assign n13747 = ~n13743 & ~n13745;
  assign n13748 = ~n13744 & n13747;
  assign n13749 = ~n13743 & n13746;
  assign n13750 = ~n13742 & n39932;
  assign n13751 = pi8  & ~n13750;
  assign n13752 = pi8  & ~n13751;
  assign n13753 = pi8  & n13750;
  assign n13754 = ~n13750 & ~n13751;
  assign n13755 = ~pi8  & ~n13750;
  assign n13756 = ~n39933 & ~n39934;
  assign n13757 = n13741 & ~n13756;
  assign n13758 = n2154 & n13010;
  assign n13759 = pi79  & n39810;
  assign n13760 = pi81  & n13040;
  assign n13761 = pi80  & n13042;
  assign n13762 = ~n13760 & ~n13761;
  assign n13763 = ~n13759 & ~n13761;
  assign n13764 = ~n13760 & n13763;
  assign n13765 = ~n13759 & n13762;
  assign n13766 = ~n13758 & n39935;
  assign n13767 = pi8  & ~n13766;
  assign n13768 = pi8  & ~n13767;
  assign n13769 = pi8  & n13766;
  assign n13770 = ~n13766 & ~n13767;
  assign n13771 = ~pi8  & ~n13766;
  assign n13772 = ~n39936 & ~n39937;
  assign n13773 = n12260 & n39656;
  assign n13774 = ~n12268 & ~n13773;
  assign n13775 = ~n13772 & n13774;
  assign n13776 = n2063 & n13010;
  assign n13777 = pi78  & n39810;
  assign n13778 = pi80  & n13040;
  assign n13779 = pi79  & n13042;
  assign n13780 = ~n13778 & ~n13779;
  assign n13781 = ~n13777 & ~n13779;
  assign n13782 = ~n13778 & n13781;
  assign n13783 = ~n13777 & n13780;
  assign n13784 = ~n13776 & n39938;
  assign n13785 = pi8  & ~n13784;
  assign n13786 = pi8  & ~n13785;
  assign n13787 = pi8  & n13784;
  assign n13788 = ~n13784 & ~n13785;
  assign n13789 = ~pi8  & ~n13784;
  assign n13790 = ~n39939 & ~n39940;
  assign n13791 = n12256 & ~n12258;
  assign n13792 = ~n12259 & ~n13791;
  assign n13793 = ~n13790 & n13792;
  assign n13794 = n678 & n13010;
  assign n13795 = pi77  & n39810;
  assign n13796 = pi79  & n13040;
  assign n13797 = pi78  & n13042;
  assign n13798 = ~n13796 & ~n13797;
  assign n13799 = ~n13795 & ~n13797;
  assign n13800 = ~n13796 & n13799;
  assign n13801 = ~n13795 & n13798;
  assign n13802 = ~n13794 & n39941;
  assign n13803 = pi8  & ~n13802;
  assign n13804 = pi8  & ~n13803;
  assign n13805 = pi8  & n13802;
  assign n13806 = ~n13802 & ~n13803;
  assign n13807 = ~pi8  & ~n13802;
  assign n13808 = ~n39942 & ~n39943;
  assign n13809 = n12252 & ~n12254;
  assign n13810 = ~n12255 & ~n13809;
  assign n13811 = ~n13808 & n13810;
  assign n13812 = n12248 & ~n12250;
  assign n13813 = ~n12251 & ~n13812;
  assign n13814 = n1578 & n13010;
  assign n13815 = pi76  & n39810;
  assign n13816 = pi78  & n13040;
  assign n13817 = pi77  & n13042;
  assign n13818 = ~n13816 & ~n13817;
  assign n13819 = ~n13815 & ~n13817;
  assign n13820 = ~n13816 & n13819;
  assign n13821 = ~n13815 & n13818;
  assign n13822 = ~n13814 & n39944;
  assign n13823 = pi8  & ~n13822;
  assign n13824 = pi8  & ~n13823;
  assign n13825 = pi8  & n13822;
  assign n13826 = ~n13822 & ~n13823;
  assign n13827 = ~pi8  & ~n13822;
  assign n13828 = ~n39945 & ~n39946;
  assign n13829 = n13813 & ~n13828;
  assign n13830 = n12239 & n39653;
  assign n13831 = ~n12247 & ~n13830;
  assign n13832 = n1596 & n13010;
  assign n13833 = pi75  & n39810;
  assign n13834 = pi77  & n13040;
  assign n13835 = pi76  & n13042;
  assign n13836 = ~n13834 & ~n13835;
  assign n13837 = ~n13833 & ~n13835;
  assign n13838 = ~n13834 & n13837;
  assign n13839 = ~n13833 & n13836;
  assign n13840 = ~n13832 & n39947;
  assign n13841 = pi8  & ~n13840;
  assign n13842 = pi8  & ~n13841;
  assign n13843 = pi8  & n13840;
  assign n13844 = ~n13840 & ~n13841;
  assign n13845 = ~pi8  & ~n13840;
  assign n13846 = ~n39948 & ~n39949;
  assign n13847 = n13831 & ~n13846;
  assign n13848 = ~n13831 & n13846;
  assign n13849 = ~n13847 & ~n13848;
  assign n13850 = n1465 & n13010;
  assign n13851 = pi74  & n39810;
  assign n13852 = pi76  & n13040;
  assign n13853 = pi75  & n13042;
  assign n13854 = ~n13852 & ~n13853;
  assign n13855 = ~n13851 & ~n13853;
  assign n13856 = ~n13852 & n13855;
  assign n13857 = ~n13851 & n13854;
  assign n13858 = ~n13850 & n39950;
  assign n13859 = pi8  & ~n13858;
  assign n13860 = pi8  & ~n13859;
  assign n13861 = pi8  & n13858;
  assign n13862 = ~n13858 & ~n13859;
  assign n13863 = ~pi8  & ~n13858;
  assign n13864 = ~n39951 & ~n39952;
  assign n13865 = n12235 & ~n12237;
  assign n13866 = ~n12238 & ~n13865;
  assign n13867 = ~n13864 & n13866;
  assign n13868 = n720 & n13010;
  assign n13869 = pi73  & n39810;
  assign n13870 = pi75  & n13040;
  assign n13871 = pi74  & n13042;
  assign n13872 = ~n13870 & ~n13871;
  assign n13873 = ~n13869 & ~n13871;
  assign n13874 = ~n13870 & n13873;
  assign n13875 = ~n13869 & n13872;
  assign n13876 = ~n13868 & n39953;
  assign n13877 = pi8  & ~n13876;
  assign n13878 = pi8  & ~n13877;
  assign n13879 = pi8  & n13876;
  assign n13880 = ~n13876 & ~n13877;
  assign n13881 = ~pi8  & ~n13876;
  assign n13882 = ~n39954 & ~n39955;
  assign n13883 = n12231 & ~n12233;
  assign n13884 = ~n12234 & ~n13883;
  assign n13885 = ~n13882 & n13884;
  assign n13886 = n1218 & n13010;
  assign n13887 = pi72  & n39810;
  assign n13888 = pi74  & n13040;
  assign n13889 = pi73  & n13042;
  assign n13890 = ~n13888 & ~n13889;
  assign n13891 = ~n13887 & ~n13889;
  assign n13892 = ~n13888 & n13891;
  assign n13893 = ~n13887 & n13890;
  assign n13894 = ~n13886 & n39956;
  assign n13895 = pi8  & ~n13894;
  assign n13896 = pi8  & ~n13895;
  assign n13897 = pi8  & n13894;
  assign n13898 = ~n13894 & ~n13895;
  assign n13899 = ~pi8  & ~n13894;
  assign n13900 = ~n39957 & ~n39958;
  assign n13901 = n12227 & ~n12229;
  assign n13902 = ~n12230 & ~n13901;
  assign n13903 = ~n13900 & n13902;
  assign n13904 = n1238 & n13010;
  assign n13905 = pi71  & n39810;
  assign n13906 = pi73  & n13040;
  assign n13907 = pi72  & n13042;
  assign n13908 = ~n13906 & ~n13907;
  assign n13909 = ~n13905 & ~n13907;
  assign n13910 = ~n13906 & n13909;
  assign n13911 = ~n13905 & n13908;
  assign n13912 = ~n13904 & n39959;
  assign n13913 = pi8  & ~n13912;
  assign n13914 = pi8  & ~n13913;
  assign n13915 = pi8  & n13912;
  assign n13916 = ~n13912 & ~n13913;
  assign n13917 = ~pi8  & ~n13912;
  assign n13918 = ~n39960 & ~n39961;
  assign n13919 = n12218 & n39650;
  assign n13920 = ~n12226 & ~n13919;
  assign n13921 = ~n13918 & n13920;
  assign n13922 = n1124 & n13010;
  assign n13923 = pi70  & n39810;
  assign n13924 = pi72  & n13040;
  assign n13925 = pi71  & n13042;
  assign n13926 = ~n13924 & ~n13925;
  assign n13927 = ~n13923 & ~n13925;
  assign n13928 = ~n13924 & n13927;
  assign n13929 = ~n13923 & n13926;
  assign n13930 = ~n13922 & n39962;
  assign n13931 = pi8  & ~n13930;
  assign n13932 = pi8  & ~n13931;
  assign n13933 = pi8  & n13930;
  assign n13934 = ~n13930 & ~n13931;
  assign n13935 = ~pi8  & ~n13930;
  assign n13936 = ~n39963 & ~n39964;
  assign n13937 = n12212 & ~n12214;
  assign n13938 = ~n12212 & ~n39647;
  assign n13939 = ~n12213 & n12218;
  assign n13940 = ~n13938 & ~n13939;
  assign n13941 = ~n39647 & ~n13937;
  assign n13942 = ~n13936 & ~n39965;
  assign n13943 = n12208 & ~n12210;
  assign n13944 = ~n12211 & ~n13943;
  assign n13945 = n927 & n13010;
  assign n13946 = pi69  & n39810;
  assign n13947 = pi71  & n13040;
  assign n13948 = pi70  & n13042;
  assign n13949 = ~n13947 & ~n13948;
  assign n13950 = ~n13946 & ~n13948;
  assign n13951 = ~n13947 & n13950;
  assign n13952 = ~n13946 & n13949;
  assign n13953 = ~n13945 & n39966;
  assign n13954 = pi8  & ~n13953;
  assign n13955 = pi8  & ~n13954;
  assign n13956 = pi8  & n13953;
  assign n13957 = ~n13953 & ~n13954;
  assign n13958 = ~pi8  & ~n13953;
  assign n13959 = ~n39967 & ~n39968;
  assign n13960 = n13944 & ~n13959;
  assign n13961 = n12201 & n39646;
  assign n13962 = ~n12207 & ~n13961;
  assign n13963 = n972 & n13010;
  assign n13964 = pi68  & n39810;
  assign n13965 = pi70  & n13040;
  assign n13966 = pi69  & n13042;
  assign n13967 = ~n13965 & ~n13966;
  assign n13968 = ~n13964 & ~n13966;
  assign n13969 = ~n13965 & n13968;
  assign n13970 = ~n13964 & n13967;
  assign n13971 = ~n13963 & n39969;
  assign n13972 = pi8  & ~n13971;
  assign n13973 = pi8  & ~n13972;
  assign n13974 = pi8  & n13971;
  assign n13975 = ~n13971 & ~n13972;
  assign n13976 = ~pi8  & ~n13971;
  assign n13977 = ~n39970 & ~n39971;
  assign n13978 = n13962 & ~n13977;
  assign n13979 = n990 & n13010;
  assign n13980 = pi67  & n39810;
  assign n13981 = pi69  & n13040;
  assign n13982 = pi68  & n13042;
  assign n13983 = ~n13981 & ~n13982;
  assign n13984 = ~n13980 & ~n13982;
  assign n13985 = ~n13981 & n13984;
  assign n13986 = ~n13980 & n13983;
  assign n13987 = ~n13979 & n39972;
  assign n13988 = pi8  & ~n13987;
  assign n13989 = pi8  & ~n13988;
  assign n13990 = pi8  & n13987;
  assign n13991 = ~n13987 & ~n13988;
  assign n13992 = ~pi8  & ~n13987;
  assign n13993 = ~n39973 & ~n39974;
  assign n13994 = pi11  & ~n39638;
  assign n13995 = n39641 & ~n13994;
  assign n13996 = ~n39641 & n13994;
  assign n13997 = ~n39638 & n12183;
  assign n13998 = ~n39642 & ~n13997;
  assign n13999 = ~n13995 & ~n13996;
  assign n14000 = ~n13993 & n39975;
  assign n14001 = n871 & n13010;
  assign n14002 = pi66  & n39810;
  assign n14003 = pi68  & n13040;
  assign n14004 = pi67  & n13042;
  assign n14005 = ~n14003 & ~n14004;
  assign n14006 = ~n14002 & ~n14004;
  assign n14007 = ~n14003 & n14006;
  assign n14008 = ~n14002 & n14005;
  assign n14009 = ~n14001 & n39976;
  assign n14010 = pi8  & ~n14009;
  assign n14011 = pi8  & ~n14010;
  assign n14012 = pi8  & n14009;
  assign n14013 = ~n14009 & ~n14010;
  assign n14014 = ~pi8  & ~n14009;
  assign n14015 = ~n39977 & ~n39978;
  assign n14016 = pi11  & n12157;
  assign n14017 = ~n12156 & n14016;
  assign n14018 = n12156 & ~n14016;
  assign n14019 = ~n12158 & n12162;
  assign n14020 = ~n39638 & ~n14019;
  assign n14021 = ~n14017 & ~n14018;
  assign n14022 = ~n14015 & n39979;
  assign n14023 = n37515 & n13010;
  assign n14024 = pi65  & n13040;
  assign n14025 = pi64  & n13042;
  assign n14026 = ~n14024 & ~n14025;
  assign n14027 = ~n14023 & n14026;
  assign n14028 = pi64  & n39807;
  assign n14029 = pi8  & ~n14028;
  assign n14030 = pi8  & ~n14027;
  assign n14031 = pi8  & ~n14030;
  assign n14032 = ~n14027 & ~n14030;
  assign n14033 = ~n14031 & ~n14032;
  assign n14034 = n14029 & ~n14033;
  assign n14035 = n14027 & n14029;
  assign n14036 = pi64  & n39810;
  assign n14037 = pi65  & n13042;
  assign n14038 = ~n37521 & n13010;
  assign n14039 = pi66  & n13040;
  assign n14040 = ~n14038 & ~n14039;
  assign n14041 = ~n14037 & ~n14038;
  assign n14042 = ~n14039 & n14041;
  assign n14043 = ~n14037 & ~n14039;
  assign n14044 = ~n14038 & n14043;
  assign n14045 = ~n14037 & n14040;
  assign n14046 = ~n14036 & ~n14037;
  assign n14047 = ~n14039 & n14046;
  assign n14048 = ~n14036 & n14043;
  assign n14049 = ~n14038 & n39982;
  assign n14050 = ~n14036 & n39981;
  assign n14051 = pi8  & ~n39983;
  assign n14052 = pi8  & ~n14051;
  assign n14053 = ~n39983 & ~n14051;
  assign n14054 = ~n14052 & ~n14053;
  assign n14055 = n39980 & ~n14054;
  assign n14056 = n39980 & n39983;
  assign n14057 = n12157 & n39984;
  assign n14058 = n847 & n13010;
  assign n14059 = pi65  & n39810;
  assign n14060 = pi67  & n13040;
  assign n14061 = pi66  & n13042;
  assign n14062 = ~n14060 & ~n14061;
  assign n14063 = ~n14059 & ~n14061;
  assign n14064 = ~n14060 & n14063;
  assign n14065 = ~n14059 & n14062;
  assign n14066 = ~n14058 & n39985;
  assign n14067 = pi8  & ~n14066;
  assign n14068 = pi8  & ~n14067;
  assign n14069 = pi8  & n14066;
  assign n14070 = ~n14066 & ~n14067;
  assign n14071 = ~pi8  & ~n14066;
  assign n14072 = ~n39986 & ~n39987;
  assign n14073 = ~n12157 & ~n39984;
  assign n14074 = n12157 & ~n39984;
  assign n14075 = ~n12157 & n39984;
  assign n14076 = ~n14074 & ~n14075;
  assign n14077 = ~n14057 & ~n14073;
  assign n14078 = ~n14072 & ~n39988;
  assign n14079 = ~n14057 & ~n14078;
  assign n14080 = n14015 & ~n39979;
  assign n14081 = ~n14022 & ~n14080;
  assign n14082 = ~n14079 & n14081;
  assign n14083 = ~n14022 & ~n14082;
  assign n14084 = n13993 & ~n39975;
  assign n14085 = n39975 & ~n14000;
  assign n14086 = n13993 & n39975;
  assign n14087 = ~n13993 & ~n14000;
  assign n14088 = ~n13993 & ~n39975;
  assign n14089 = ~n39989 & ~n39990;
  assign n14090 = ~n14000 & ~n14084;
  assign n14091 = ~n14083 & ~n39991;
  assign n14092 = ~n14000 & ~n14091;
  assign n14093 = ~n13962 & n13977;
  assign n14094 = n13962 & ~n13978;
  assign n14095 = n13962 & n13977;
  assign n14096 = ~n13977 & ~n13978;
  assign n14097 = ~n13962 & ~n13977;
  assign n14098 = ~n39992 & ~n39993;
  assign n14099 = ~n13978 & ~n14093;
  assign n14100 = ~n14092 & ~n39994;
  assign n14101 = ~n13978 & ~n14100;
  assign n14102 = ~n13944 & n13959;
  assign n14103 = n13944 & ~n13960;
  assign n14104 = n13944 & n13959;
  assign n14105 = ~n13959 & ~n13960;
  assign n14106 = ~n13944 & ~n13959;
  assign n14107 = ~n39995 & ~n39996;
  assign n14108 = ~n13960 & ~n14102;
  assign n14109 = ~n14101 & ~n39997;
  assign n14110 = ~n13960 & ~n14109;
  assign n14111 = n13936 & n39965;
  assign n14112 = ~n13942 & ~n14111;
  assign n14113 = ~n14110 & n14112;
  assign n14114 = ~n13942 & ~n14113;
  assign n14115 = n13918 & ~n13920;
  assign n14116 = ~n13918 & ~n13921;
  assign n14117 = ~n13918 & ~n13920;
  assign n14118 = n13920 & ~n13921;
  assign n14119 = n13918 & n13920;
  assign n14120 = ~n39998 & ~n39999;
  assign n14121 = ~n13921 & ~n14115;
  assign n14122 = ~n14114 & ~n40000;
  assign n14123 = ~n13921 & ~n14122;
  assign n14124 = n13900 & ~n13902;
  assign n14125 = ~n13903 & ~n14124;
  assign n14126 = ~n14123 & n14125;
  assign n14127 = ~n13903 & ~n14126;
  assign n14128 = n13882 & ~n13884;
  assign n14129 = ~n13885 & ~n14128;
  assign n14130 = ~n14127 & n14129;
  assign n14131 = ~n13885 & ~n14130;
  assign n14132 = n13864 & ~n13866;
  assign n14133 = ~n13867 & ~n14132;
  assign n14134 = ~n14131 & n14133;
  assign n14135 = ~n13867 & ~n14134;
  assign n14136 = n13849 & ~n14135;
  assign n14137 = ~n13847 & ~n14136;
  assign n14138 = ~n13813 & n13828;
  assign n14139 = n13813 & ~n13829;
  assign n14140 = n13813 & n13828;
  assign n14141 = ~n13828 & ~n13829;
  assign n14142 = ~n13813 & ~n13828;
  assign n14143 = ~n40001 & ~n40002;
  assign n14144 = ~n13829 & ~n14138;
  assign n14145 = ~n14137 & ~n40003;
  assign n14146 = ~n13829 & ~n14145;
  assign n14147 = n13808 & ~n13810;
  assign n14148 = ~n13811 & ~n14147;
  assign n14149 = ~n14146 & n14148;
  assign n14150 = ~n13811 & ~n14149;
  assign n14151 = n13790 & ~n13792;
  assign n14152 = ~n13793 & ~n14151;
  assign n14153 = ~n14150 & n14152;
  assign n14154 = ~n13793 & ~n14153;
  assign n14155 = n13772 & ~n13774;
  assign n14156 = ~n13772 & ~n13775;
  assign n14157 = ~n13772 & ~n13774;
  assign n14158 = n13774 & ~n13775;
  assign n14159 = n13772 & n13774;
  assign n14160 = ~n40004 & ~n40005;
  assign n14161 = ~n13775 & ~n14155;
  assign n14162 = ~n14154 & ~n40006;
  assign n14163 = ~n13775 & ~n14162;
  assign n14164 = ~n13741 & n13756;
  assign n14165 = ~n13757 & ~n14164;
  assign n14166 = ~n14163 & n14165;
  assign n14167 = ~n13757 & ~n14166;
  assign n14168 = ~n13723 & n13738;
  assign n14169 = n13723 & ~n13739;
  assign n14170 = n13723 & n13738;
  assign n14171 = ~n13738 & ~n13739;
  assign n14172 = ~n13723 & ~n13738;
  assign n14173 = ~n40007 & ~n40008;
  assign n14174 = ~n13739 & ~n14168;
  assign n14175 = ~n14167 & ~n40009;
  assign n14176 = ~n13739 & ~n14175;
  assign n14177 = ~n13705 & n13720;
  assign n14178 = n13705 & ~n13721;
  assign n14179 = n13705 & n13720;
  assign n14180 = ~n13720 & ~n13721;
  assign n14181 = ~n13705 & ~n13720;
  assign n14182 = ~n40010 & ~n40011;
  assign n14183 = ~n13721 & ~n14177;
  assign n14184 = ~n14176 & ~n40012;
  assign n14185 = ~n13721 & ~n14184;
  assign n14186 = n13703 & ~n14185;
  assign n14187 = ~n13701 & ~n14186;
  assign n14188 = n13683 & ~n14187;
  assign n14189 = ~n13681 & ~n14188;
  assign n14190 = n13657 & n39919;
  assign n14191 = ~n39919 & ~n13663;
  assign n14192 = n13657 & ~n39919;
  assign n14193 = ~n13657 & ~n13663;
  assign n14194 = ~n13657 & n39919;
  assign n14195 = ~n40013 & ~n40014;
  assign n14196 = ~n13663 & ~n14190;
  assign n14197 = ~n14189 & ~n40015;
  assign n14198 = ~n13663 & ~n14197;
  assign n14199 = n13636 & n39915;
  assign n14200 = ~n13642 & ~n14199;
  assign n14201 = ~n14198 & n14200;
  assign n14202 = ~n13642 & ~n14201;
  assign n14203 = ~n13605 & n13620;
  assign n14204 = n13605 & ~n13621;
  assign n14205 = n13605 & n13620;
  assign n14206 = ~n13620 & ~n13621;
  assign n14207 = ~n13605 & ~n13620;
  assign n14208 = ~n40016 & ~n40017;
  assign n14209 = ~n13621 & ~n14203;
  assign n14210 = ~n14202 & ~n40018;
  assign n14211 = ~n13621 & ~n14210;
  assign n14212 = ~n13587 & n13602;
  assign n14213 = n13587 & ~n13603;
  assign n14214 = n13587 & n13602;
  assign n14215 = ~n13602 & ~n13603;
  assign n14216 = ~n13587 & ~n13602;
  assign n14217 = ~n40019 & ~n40020;
  assign n14218 = ~n13603 & ~n14212;
  assign n14219 = ~n14211 & ~n40021;
  assign n14220 = ~n13603 & ~n14219;
  assign n14221 = ~n13569 & n13584;
  assign n14222 = n13569 & ~n13585;
  assign n14223 = n13569 & n13584;
  assign n14224 = ~n13584 & ~n13585;
  assign n14225 = ~n13569 & ~n13584;
  assign n14226 = ~n40022 & ~n40023;
  assign n14227 = ~n13585 & ~n14221;
  assign n14228 = ~n14220 & ~n40024;
  assign n14229 = ~n13585 & ~n14228;
  assign n14230 = n13561 & n39902;
  assign n14231 = ~n39902 & ~n13567;
  assign n14232 = n13561 & ~n39902;
  assign n14233 = ~n13561 & ~n13567;
  assign n14234 = ~n13561 & n39902;
  assign n14235 = ~n40025 & ~n40026;
  assign n14236 = ~n13567 & ~n14230;
  assign n14237 = ~n14229 & ~n40027;
  assign n14238 = ~n13567 & ~n14237;
  assign n14239 = ~n13530 & n13545;
  assign n14240 = n13530 & ~n13546;
  assign n14241 = n13530 & n13545;
  assign n14242 = ~n13545 & ~n13546;
  assign n14243 = ~n13530 & ~n13545;
  assign n14244 = ~n40028 & ~n40029;
  assign n14245 = ~n13546 & ~n14239;
  assign n14246 = ~n14238 & ~n40030;
  assign n14247 = ~n13546 & ~n14246;
  assign n14248 = n13522 & n39895;
  assign n14249 = ~n13528 & ~n14248;
  assign n14250 = ~n14247 & n14249;
  assign n14251 = ~n13528 & ~n14250;
  assign n14252 = n13504 & ~n13506;
  assign n14253 = ~n13507 & ~n14252;
  assign n14254 = ~n14251 & n14253;
  assign n14255 = ~n13507 & ~n14254;
  assign n14256 = n13486 & ~n13488;
  assign n14257 = ~n13489 & ~n14256;
  assign n14258 = ~n14255 & n14257;
  assign n14259 = ~n13489 & ~n14258;
  assign n14260 = ~n13455 & n13470;
  assign n14261 = n13455 & ~n13471;
  assign n14262 = n13455 & n13470;
  assign n14263 = ~n13470 & ~n13471;
  assign n14264 = ~n13455 & ~n13470;
  assign n14265 = ~n40031 & ~n40032;
  assign n14266 = ~n13471 & ~n14260;
  assign n14267 = ~n14259 & ~n40033;
  assign n14268 = ~n13471 & ~n14267;
  assign n14269 = n13450 & ~n13452;
  assign n14270 = ~n13453 & ~n14269;
  assign n14271 = ~n14268 & n14270;
  assign n14272 = ~n13453 & ~n14271;
  assign n14273 = ~n13419 & n13434;
  assign n14274 = n13419 & ~n13435;
  assign n14275 = n13419 & n13434;
  assign n14276 = ~n13434 & ~n13435;
  assign n14277 = ~n13419 & ~n13434;
  assign n14278 = ~n40034 & ~n40035;
  assign n14279 = ~n13435 & ~n14273;
  assign n14280 = ~n14272 & ~n40036;
  assign n14281 = ~n13435 & ~n14280;
  assign n14282 = n13411 & n39876;
  assign n14283 = ~n13417 & ~n14282;
  assign n14284 = ~n14281 & n14283;
  assign n14285 = ~n13417 & ~n14284;
  assign n14286 = ~n13380 & n13395;
  assign n14287 = ~n13396 & ~n14286;
  assign n14288 = ~n14285 & ~n14286;
  assign n14289 = ~n13396 & n14288;
  assign n14290 = ~n14285 & n14287;
  assign n14291 = ~n13396 & ~n40037;
  assign n14292 = ~n13362 & n13377;
  assign n14293 = n13362 & ~n13378;
  assign n14294 = n13362 & n13377;
  assign n14295 = ~n13377 & ~n13378;
  assign n14296 = ~n13362 & ~n13377;
  assign n14297 = ~n40038 & ~n40039;
  assign n14298 = ~n13378 & ~n14292;
  assign n14299 = ~n14291 & ~n40040;
  assign n14300 = ~n13378 & ~n14299;
  assign n14301 = ~n13344 & n13359;
  assign n14302 = n13344 & ~n13360;
  assign n14303 = n13344 & n13359;
  assign n14304 = ~n13359 & ~n13360;
  assign n14305 = ~n13344 & ~n13359;
  assign n14306 = ~n40041 & ~n40042;
  assign n14307 = ~n13360 & ~n14301;
  assign n14308 = ~n14300 & ~n40043;
  assign n14309 = ~n13360 & ~n14308;
  assign n14310 = ~n13326 & n13341;
  assign n14311 = ~n13342 & ~n14310;
  assign n14312 = ~n14309 & ~n14310;
  assign n14313 = ~n13342 & n14312;
  assign n14314 = ~n14309 & n14311;
  assign n14315 = ~n13342 & ~n40044;
  assign n14316 = ~n13308 & n13323;
  assign n14317 = ~n13324 & ~n14316;
  assign n14318 = ~n14315 & ~n14316;
  assign n14319 = ~n13324 & n14318;
  assign n14320 = ~n14315 & n14317;
  assign n14321 = ~n13324 & ~n40045;
  assign n14322 = ~n13290 & n13305;
  assign n14323 = n13290 & ~n13306;
  assign n14324 = n13290 & n13305;
  assign n14325 = ~n13305 & ~n13306;
  assign n14326 = ~n13290 & ~n13305;
  assign n14327 = ~n40046 & ~n40047;
  assign n14328 = ~n13306 & ~n14322;
  assign n14329 = ~n14321 & ~n40048;
  assign n14330 = ~n13306 & ~n14329;
  assign n14331 = ~n13272 & n13287;
  assign n14332 = n13272 & ~n13288;
  assign n14333 = n13272 & n13287;
  assign n14334 = ~n13287 & ~n13288;
  assign n14335 = ~n13272 & ~n13287;
  assign n14336 = ~n40049 & ~n40050;
  assign n14337 = ~n13288 & ~n14331;
  assign n14338 = ~n14330 & ~n40051;
  assign n14339 = ~n13288 & ~n14338;
  assign n14340 = ~n13254 & n13269;
  assign n14341 = ~n13270 & ~n14340;
  assign n14342 = ~n14339 & ~n14340;
  assign n14343 = ~n13270 & n14342;
  assign n14344 = ~n14339 & n14341;
  assign n14345 = ~n13270 & ~n40052;
  assign n14346 = ~n13236 & n13251;
  assign n14347 = n13236 & ~n13252;
  assign n14348 = n13236 & n13251;
  assign n14349 = ~n13251 & ~n13252;
  assign n14350 = ~n13236 & ~n13251;
  assign n14351 = ~n40053 & ~n40054;
  assign n14352 = ~n13252 & ~n14346;
  assign n14353 = ~n14345 & ~n40055;
  assign n14354 = ~n13252 & ~n14353;
  assign n14355 = n13228 & n39845;
  assign n14356 = ~n39845 & ~n13234;
  assign n14357 = n13228 & ~n39845;
  assign n14358 = ~n13228 & ~n13234;
  assign n14359 = ~n13228 & n39845;
  assign n14360 = ~n40056 & ~n40057;
  assign n14361 = ~n13234 & ~n14355;
  assign n14362 = ~n14354 & ~n40058;
  assign n14363 = ~n13234 & ~n14362;
  assign n14364 = n13207 & n39841;
  assign n14365 = ~n39841 & ~n13213;
  assign n14366 = n13207 & ~n39841;
  assign n14367 = ~n13207 & ~n13213;
  assign n14368 = ~n13207 & n39841;
  assign n14369 = ~n40059 & ~n40060;
  assign n14370 = ~n13213 & ~n14364;
  assign n14371 = ~n14363 & ~n40061;
  assign n14372 = ~n13213 & ~n14371;
  assign n14373 = n13186 & n39837;
  assign n14374 = ~n39837 & ~n13192;
  assign n14375 = n13186 & ~n39837;
  assign n14376 = ~n13186 & ~n13192;
  assign n14377 = ~n13186 & n39837;
  assign n14378 = ~n40062 & ~n40063;
  assign n14379 = ~n13192 & ~n14373;
  assign n14380 = ~n14372 & ~n40064;
  assign n14381 = ~n13192 & ~n14380;
  assign n14382 = n13168 & ~n13170;
  assign n14383 = ~n13171 & ~n14382;
  assign n14384 = ~n14381 & n14383;
  assign n14385 = ~n13171 & ~n14384;
  assign n14386 = n13150 & ~n13152;
  assign n14387 = ~n13150 & ~n13153;
  assign n14388 = ~n13150 & ~n13152;
  assign n14389 = n13152 & ~n13153;
  assign n14390 = n13150 & n13152;
  assign n14391 = ~n40065 & ~n40066;
  assign n14392 = ~n13153 & ~n14386;
  assign n14393 = ~n14385 & ~n40067;
  assign n14394 = ~n13153 & ~n14393;
  assign n14395 = n13130 & ~n13134;
  assign n14396 = ~n13130 & ~n13135;
  assign n14397 = ~n13130 & ~n13134;
  assign n14398 = n13134 & ~n13135;
  assign n14399 = n13130 & n13134;
  assign n14400 = ~n40068 & ~n40069;
  assign n14401 = ~n13135 & ~n14395;
  assign n14402 = ~n14394 & ~n40070;
  assign n14403 = ~n13135 & ~n14402;
  assign n14404 = n13112 & ~n13114;
  assign n14405 = ~n13115 & ~n14404;
  assign n14406 = ~n14403 & n14405;
  assign n14407 = ~n13115 & ~n14406;
  assign n14408 = n13094 & ~n13096;
  assign n14409 = ~n13094 & ~n13097;
  assign n14410 = ~n13094 & ~n13096;
  assign n14411 = n13096 & ~n13097;
  assign n14412 = n13094 & n13096;
  assign n14413 = ~n40071 & ~n40072;
  assign n14414 = ~n13097 & ~n14408;
  assign n14415 = ~n14407 & ~n40073;
  assign n14416 = ~n13097 & ~n14415;
  assign n14417 = n13072 & ~n13076;
  assign n14418 = ~n13077 & ~n14417;
  assign n14419 = ~n14416 & n14418;
  assign n14420 = ~n13077 & ~n14419;
  assign n14421 = ~n12997 & n13054;
  assign n14422 = n12997 & ~n13055;
  assign n14423 = n12997 & n13054;
  assign n14424 = ~n13054 & ~n13055;
  assign n14425 = ~n12997 & ~n13054;
  assign n14426 = ~n40074 & ~n40075;
  assign n14427 = ~n13055 & ~n14421;
  assign n14428 = ~n14420 & ~n40076;
  assign n14429 = ~n13055 & ~n14428;
  assign n14430 = ~n12993 & ~n12995;
  assign n14431 = n269 & n13079;
  assign n14432 = pi115  & n37475;
  assign n14433 = pi117  & n536;
  assign n14434 = pi116  & n538;
  assign n14435 = ~n14433 & ~n14434;
  assign n14436 = ~n14432 & ~n14434;
  assign n14437 = ~n14433 & n14436;
  assign n14438 = ~n14432 & n14435;
  assign n14439 = ~n14431 & n40077;
  assign n14440 = pi11  & ~n14439;
  assign n14441 = pi11  & ~n14440;
  assign n14442 = pi11  & n14439;
  assign n14443 = ~n14439 & ~n14440;
  assign n14444 = ~pi11  & ~n14439;
  assign n14445 = ~n40078 & ~n40079;
  assign n14446 = ~n12987 & ~n12989;
  assign n14447 = ~n12981 & ~n12983;
  assign n14448 = n565 & n8175;
  assign n14449 = pi109  & n38895;
  assign n14450 = pi111  & n8190;
  assign n14451 = pi110  & n8192;
  assign n14452 = ~n14450 & ~n14451;
  assign n14453 = ~n14449 & ~n14451;
  assign n14454 = ~n14450 & n14453;
  assign n14455 = ~n14449 & n14452;
  assign n14456 = ~n14448 & n40080;
  assign n14457 = pi17  & ~n14456;
  assign n14458 = pi17  & ~n14457;
  assign n14459 = pi17  & n14456;
  assign n14460 = ~n14456 & ~n14457;
  assign n14461 = ~pi17  & ~n14456;
  assign n14462 = ~n40081 & ~n40082;
  assign n14463 = n6785 & n9277;
  assign n14464 = pi106  & n38631;
  assign n14465 = pi108  & n6800;
  assign n14466 = pi107  & n6802;
  assign n14467 = ~n14465 & ~n14466;
  assign n14468 = ~n14464 & ~n14466;
  assign n14469 = ~n14465 & n14468;
  assign n14470 = ~n14464 & n14467;
  assign n14471 = ~n14463 & n40083;
  assign n14472 = pi20  & ~n14471;
  assign n14473 = pi20  & ~n14472;
  assign n14474 = pi20  & n14471;
  assign n14475 = ~n14471 & ~n14472;
  assign n14476 = ~pi20  & ~n14471;
  assign n14477 = ~n40084 & ~n40085;
  assign n14478 = ~n12942 & ~n12951;
  assign n14479 = ~n12916 & ~n12925;
  assign n14480 = ~n12895 & ~n12899;
  assign n14481 = n607 & n5578;
  assign n14482 = pi97  & n37489;
  assign n14483 = pi99  & n620;
  assign n14484 = pi98  & n622;
  assign n14485 = ~n14483 & ~n14484;
  assign n14486 = ~n14482 & ~n14484;
  assign n14487 = ~n14483 & n14486;
  assign n14488 = ~n14482 & n14485;
  assign n14489 = ~n14481 & n40086;
  assign n14490 = pi29  & ~n14489;
  assign n14491 = pi29  & ~n14490;
  assign n14492 = pi29  & n14489;
  assign n14493 = ~n14489 & ~n14490;
  assign n14494 = ~pi29  & ~n14489;
  assign n14495 = ~n40087 & ~n40088;
  assign n14496 = ~n12881 & ~n12889;
  assign n14497 = ~n12855 & ~n12864;
  assign n14498 = ~n12829 & ~n12838;
  assign n14499 = ~n12803 & ~n12812;
  assign n14500 = n636 & n733;
  assign n14501 = pi85  & n37510;
  assign n14502 = pi87  & n746;
  assign n14503 = pi86  & n748;
  assign n14504 = ~n14502 & ~n14503;
  assign n14505 = ~n14501 & ~n14503;
  assign n14506 = ~n14502 & n14505;
  assign n14507 = ~n14501 & n14504;
  assign n14508 = ~n14500 & n40089;
  assign n14509 = pi41  & ~n14508;
  assign n14510 = pi41  & ~n14509;
  assign n14511 = pi41  & n14508;
  assign n14512 = ~n14508 & ~n14509;
  assign n14513 = ~pi41  & ~n14508;
  assign n14514 = ~n40090 & ~n40091;
  assign n14515 = n940 & n2591;
  assign n14516 = pi82  & n37541;
  assign n14517 = pi84  & n953;
  assign n14518 = pi83  & n955;
  assign n14519 = ~n14517 & ~n14518;
  assign n14520 = ~n14516 & ~n14518;
  assign n14521 = ~n14517 & n14520;
  assign n14522 = ~n14516 & n14519;
  assign n14523 = ~n14515 & n40092;
  assign n14524 = pi44  & ~n14523;
  assign n14525 = pi44  & ~n14524;
  assign n14526 = pi44  & n14523;
  assign n14527 = ~n14523 & ~n14524;
  assign n14528 = ~pi44  & ~n14523;
  assign n14529 = ~n40093 & ~n40094;
  assign n14530 = ~n12765 & ~n12774;
  assign n14531 = n785 & n2154;
  assign n14532 = pi79  & n37520;
  assign n14533 = pi81  & n787;
  assign n14534 = pi80  & n795;
  assign n14535 = ~n14533 & ~n14534;
  assign n14536 = ~n14532 & ~n14534;
  assign n14537 = ~n14533 & n14536;
  assign n14538 = ~n14532 & n14535;
  assign n14539 = ~n14531 & n40095;
  assign n14540 = pi47  & ~n14539;
  assign n14541 = pi47  & ~n14540;
  assign n14542 = pi47  & n14539;
  assign n14543 = ~n14539 & ~n14540;
  assign n14544 = ~pi47  & ~n14539;
  assign n14545 = ~n40096 & ~n40097;
  assign n14546 = ~n12727 & ~n12736;
  assign n14547 = n720 & n1971;
  assign n14548 = pi73  & n37864;
  assign n14549 = pi75  & n1973;
  assign n14550 = pi74  & n1981;
  assign n14551 = ~n14549 & ~n14550;
  assign n14552 = ~n14548 & ~n14550;
  assign n14553 = ~n14549 & n14552;
  assign n14554 = ~n14548 & n14551;
  assign n14555 = ~n14547 & n40098;
  assign n14556 = pi53  & ~n14555;
  assign n14557 = pi53  & ~n14556;
  assign n14558 = pi53  & n14555;
  assign n14559 = ~n14555 & ~n14556;
  assign n14560 = ~pi53  & ~n14555;
  assign n14561 = ~n40099 & ~n40100;
  assign n14562 = ~n12707 & ~n12709;
  assign n14563 = n1124 & n4312;
  assign n14564 = pi70  & n38376;
  assign n14565 = pi72  & n4314;
  assign n14566 = pi71  & n4322;
  assign n14567 = ~n14565 & ~n14566;
  assign n14568 = ~n14564 & ~n14566;
  assign n14569 = ~n14565 & n14568;
  assign n14570 = ~n14564 & n14567;
  assign n14571 = ~n14563 & n40101;
  assign n14572 = pi56  & ~n14571;
  assign n14573 = pi56  & ~n14572;
  assign n14574 = pi56  & n14571;
  assign n14575 = ~n14571 & ~n14572;
  assign n14576 = ~pi56  & ~n14571;
  assign n14577 = ~n40102 & ~n40103;
  assign n14578 = ~n12701 & ~n12703;
  assign n14579 = n990 & n7882;
  assign n14580 = pi67  & n39128;
  assign n14581 = pi69  & n7884;
  assign n14582 = pi68  & n7892;
  assign n14583 = ~n14581 & ~n14582;
  assign n14584 = ~n14580 & ~n14582;
  assign n14585 = ~n14581 & n14584;
  assign n14586 = ~n14580 & n14583;
  assign n14587 = ~n14579 & n40104;
  assign n14588 = pi59  & ~n14587;
  assign n14589 = pi59  & ~n14588;
  assign n14590 = pi59  & n14587;
  assign n14591 = ~n14587 & ~n14588;
  assign n14592 = ~pi59  & ~n14587;
  assign n14593 = ~n40105 & ~n40106;
  assign n14594 = pi62  & ~n39747;
  assign n14595 = ~n39429 & n39745;
  assign n14596 = ~n39429 & ~n39746;
  assign n14597 = n39745 & n14596;
  assign n14598 = ~n39746 & n14595;
  assign n14599 = pi64  & n40107;
  assign n14600 = pi65  & n12684;
  assign n14601 = ~n37521 & n12674;
  assign n14602 = pi66  & n12676;
  assign n14603 = ~n14601 & ~n14602;
  assign n14604 = ~n14600 & ~n14601;
  assign n14605 = ~n14602 & n14604;
  assign n14606 = ~n14600 & ~n14602;
  assign n14607 = ~n14601 & n14606;
  assign n14608 = ~n14600 & n14603;
  assign n14609 = ~n14599 & ~n14600;
  assign n14610 = ~n14602 & n14609;
  assign n14611 = ~n14599 & n14606;
  assign n14612 = ~n14601 & n40109;
  assign n14613 = ~n14599 & n40108;
  assign n14614 = ~n14594 & n40110;
  assign n14615 = n14594 & ~n40110;
  assign n14616 = pi62  & ~n40110;
  assign n14617 = pi62  & ~n14616;
  assign n14618 = ~n40110 & ~n14616;
  assign n14619 = ~n14617 & ~n14618;
  assign n14620 = n39747 & ~n14619;
  assign n14621 = n39747 & n40110;
  assign n14622 = ~n39747 & n14619;
  assign n14623 = ~n40111 & ~n14622;
  assign n14624 = ~n14614 & ~n14615;
  assign n14625 = ~n14593 & n40112;
  assign n14626 = n14593 & ~n40112;
  assign n14627 = ~n14625 & ~n14626;
  assign n14628 = ~n14578 & ~n14626;
  assign n14629 = ~n14625 & n14628;
  assign n14630 = ~n14578 & n14627;
  assign n14631 = n14578 & ~n14627;
  assign n14632 = ~n14578 & ~n40113;
  assign n14633 = ~n14625 & ~n40113;
  assign n14634 = ~n14626 & n14633;
  assign n14635 = ~n14632 & ~n14634;
  assign n14636 = ~n40113 & ~n14631;
  assign n14637 = n14577 & n40114;
  assign n14638 = ~n14577 & ~n40114;
  assign n14639 = ~n14637 & ~n14638;
  assign n14640 = ~n14562 & n14639;
  assign n14641 = n14562 & ~n14639;
  assign n14642 = ~n14640 & ~n14641;
  assign n14643 = n14561 & ~n14642;
  assign n14644 = ~n14561 & n14642;
  assign n14645 = ~n14643 & ~n14644;
  assign n14646 = ~n14546 & n14645;
  assign n14647 = n14546 & ~n14645;
  assign n14648 = ~n14646 & ~n14647;
  assign n14649 = n894 & n1578;
  assign n14650 = pi76  & n37580;
  assign n14651 = pi78  & n896;
  assign n14652 = pi77  & n904;
  assign n14653 = ~n14651 & ~n14652;
  assign n14654 = ~n14650 & ~n14652;
  assign n14655 = ~n14651 & n14654;
  assign n14656 = ~n14650 & n14653;
  assign n14657 = ~n14649 & n40115;
  assign n14658 = pi50  & ~n14657;
  assign n14659 = pi50  & ~n14658;
  assign n14660 = pi50  & n14657;
  assign n14661 = ~n14657 & ~n14658;
  assign n14662 = ~pi50  & ~n14657;
  assign n14663 = ~n40116 & ~n40117;
  assign n14664 = n14648 & ~n14663;
  assign n14665 = ~n14648 & n14663;
  assign n14666 = n14648 & ~n14664;
  assign n14667 = n14648 & n14663;
  assign n14668 = ~n14663 & ~n14664;
  assign n14669 = ~n14648 & ~n14663;
  assign n14670 = ~n40118 & ~n40119;
  assign n14671 = ~n14664 & ~n14665;
  assign n14672 = ~n12761 & ~n40120;
  assign n14673 = n12761 & n40120;
  assign n14674 = ~n14672 & ~n14673;
  assign n14675 = ~n14545 & n14674;
  assign n14676 = n14545 & ~n14674;
  assign n14677 = ~n14545 & ~n14675;
  assign n14678 = ~n14545 & ~n14674;
  assign n14679 = n14674 & ~n14675;
  assign n14680 = n14545 & n14674;
  assign n14681 = ~n40121 & ~n40122;
  assign n14682 = ~n14675 & ~n14676;
  assign n14683 = ~n14530 & ~n40123;
  assign n14684 = n14530 & n40123;
  assign n14685 = ~n14530 & ~n14683;
  assign n14686 = ~n14530 & n40123;
  assign n14687 = ~n40123 & ~n14683;
  assign n14688 = n14530 & ~n40123;
  assign n14689 = ~n40124 & ~n40125;
  assign n14690 = ~n14683 & ~n14684;
  assign n14691 = ~n14529 & ~n40126;
  assign n14692 = n14529 & n40126;
  assign n14693 = ~n40126 & ~n14691;
  assign n14694 = ~n14529 & ~n14691;
  assign n14695 = ~n14693 & ~n14694;
  assign n14696 = ~n14691 & ~n14692;
  assign n14697 = ~n12799 & ~n40127;
  assign n14698 = n12799 & n40127;
  assign n14699 = ~n12799 & n40127;
  assign n14700 = n12799 & ~n40127;
  assign n14701 = ~n14699 & ~n14700;
  assign n14702 = ~n14697 & ~n14698;
  assign n14703 = ~n14514 & ~n40128;
  assign n14704 = n14514 & n40128;
  assign n14705 = ~n14703 & ~n14704;
  assign n14706 = n14499 & ~n14705;
  assign n14707 = ~n14499 & n14705;
  assign n14708 = ~n14706 & ~n14707;
  assign n14709 = n691 & n3566;
  assign n14710 = pi88  & n37503;
  assign n14711 = pi90  & n704;
  assign n14712 = pi89  & n706;
  assign n14713 = ~n14711 & ~n14712;
  assign n14714 = ~n14710 & ~n14712;
  assign n14715 = ~n14711 & n14714;
  assign n14716 = ~n14710 & n14713;
  assign n14717 = ~n14709 & n40129;
  assign n14718 = pi38  & ~n14717;
  assign n14719 = pi38  & ~n14718;
  assign n14720 = pi38  & n14717;
  assign n14721 = ~n14717 & ~n14718;
  assign n14722 = ~pi38  & ~n14717;
  assign n14723 = ~n40130 & ~n40131;
  assign n14724 = n14708 & ~n14723;
  assign n14725 = ~n14708 & n14723;
  assign n14726 = n14708 & ~n14724;
  assign n14727 = n14708 & n14723;
  assign n14728 = ~n14723 & ~n14724;
  assign n14729 = ~n14708 & ~n14723;
  assign n14730 = ~n40132 & ~n40133;
  assign n14731 = ~n14724 & ~n14725;
  assign n14732 = n14498 & n40134;
  assign n14733 = ~n14498 & ~n40134;
  assign n14734 = ~n14732 & ~n14733;
  assign n14735 = n2104 & n4544;
  assign n14736 = pi91  & n37758;
  assign n14737 = pi93  & n2117;
  assign n14738 = pi92  & n2119;
  assign n14739 = ~n14737 & ~n14738;
  assign n14740 = ~n14736 & ~n14738;
  assign n14741 = ~n14737 & n14740;
  assign n14742 = ~n14736 & n14739;
  assign n14743 = ~n14735 & n40135;
  assign n14744 = pi35  & ~n14743;
  assign n14745 = pi35  & ~n14744;
  assign n14746 = pi35  & n14743;
  assign n14747 = ~n14743 & ~n14744;
  assign n14748 = ~pi35  & ~n14743;
  assign n14749 = ~n40136 & ~n40137;
  assign n14750 = n14734 & ~n14749;
  assign n14751 = ~n14734 & n14749;
  assign n14752 = n14734 & ~n14750;
  assign n14753 = n14734 & n14749;
  assign n14754 = ~n14749 & ~n14750;
  assign n14755 = ~n14734 & ~n14749;
  assign n14756 = ~n40138 & ~n40139;
  assign n14757 = ~n14750 & ~n14751;
  assign n14758 = n14497 & n40140;
  assign n14759 = ~n14497 & ~n40140;
  assign n14760 = ~n14758 & ~n14759;
  assign n14761 = n649 & n5281;
  assign n14762 = pi94  & n37496;
  assign n14763 = pi96  & n662;
  assign n14764 = pi95  & n664;
  assign n14765 = ~n14763 & ~n14764;
  assign n14766 = ~n14762 & ~n14764;
  assign n14767 = ~n14763 & n14766;
  assign n14768 = ~n14762 & n14765;
  assign n14769 = ~n14761 & n40141;
  assign n14770 = pi32  & ~n14769;
  assign n14771 = pi32  & ~n14770;
  assign n14772 = pi32  & n14769;
  assign n14773 = ~n14769 & ~n14770;
  assign n14774 = ~pi32  & ~n14769;
  assign n14775 = ~n40142 & ~n40143;
  assign n14776 = n14760 & ~n14775;
  assign n14777 = ~n14760 & n14775;
  assign n14778 = ~n14776 & ~n14777;
  assign n14779 = ~n14496 & ~n14777;
  assign n14780 = ~n14776 & n14779;
  assign n14781 = ~n14496 & n14778;
  assign n14782 = n14496 & ~n14778;
  assign n14783 = ~n14496 & ~n40144;
  assign n14784 = ~n14776 & ~n40144;
  assign n14785 = ~n14777 & n14784;
  assign n14786 = ~n14783 & ~n14785;
  assign n14787 = ~n40144 & ~n14782;
  assign n14788 = ~n14495 & ~n40145;
  assign n14789 = n14495 & n40145;
  assign n14790 = ~n40145 & ~n14788;
  assign n14791 = n14495 & ~n40145;
  assign n14792 = ~n14495 & ~n14788;
  assign n14793 = ~n14495 & n40145;
  assign n14794 = ~n40146 & ~n40147;
  assign n14795 = ~n14788 & ~n14789;
  assign n14796 = n14480 & n40148;
  assign n14797 = ~n14480 & ~n40148;
  assign n14798 = ~n14796 & ~n14797;
  assign n14799 = n4492 & n6819;
  assign n14800 = pi100  & n38208;
  assign n14801 = pi102  & n4507;
  assign n14802 = pi101  & n4509;
  assign n14803 = ~n14801 & ~n14802;
  assign n14804 = ~n14800 & ~n14802;
  assign n14805 = ~n14801 & n14804;
  assign n14806 = ~n14800 & n14803;
  assign n14807 = ~n14799 & n40149;
  assign n14808 = pi26  & ~n14807;
  assign n14809 = pi26  & ~n14808;
  assign n14810 = pi26  & n14807;
  assign n14811 = ~n14807 & ~n14808;
  assign n14812 = ~pi26  & ~n14807;
  assign n14813 = ~n40150 & ~n40151;
  assign n14814 = n14798 & ~n14813;
  assign n14815 = ~n14798 & n14813;
  assign n14816 = n14798 & ~n14814;
  assign n14817 = n14798 & n14813;
  assign n14818 = ~n14813 & ~n14814;
  assign n14819 = ~n14798 & ~n14813;
  assign n14820 = ~n40152 & ~n40153;
  assign n14821 = ~n14814 & ~n14815;
  assign n14822 = n14479 & n40154;
  assign n14823 = ~n14479 & ~n40154;
  assign n14824 = ~n14822 & ~n14823;
  assign n14825 = n5576 & n8229;
  assign n14826 = pi103  & n38406;
  assign n14827 = pi105  & n5591;
  assign n14828 = pi104  & n5593;
  assign n14829 = ~n14827 & ~n14828;
  assign n14830 = ~n14826 & ~n14828;
  assign n14831 = ~n14827 & n14830;
  assign n14832 = ~n14826 & n14829;
  assign n14833 = ~n14825 & n40155;
  assign n14834 = pi23  & ~n14833;
  assign n14835 = pi23  & ~n14834;
  assign n14836 = pi23  & n14833;
  assign n14837 = ~n14833 & ~n14834;
  assign n14838 = ~pi23  & ~n14833;
  assign n14839 = ~n40156 & ~n40157;
  assign n14840 = n14824 & ~n14839;
  assign n14841 = ~n14824 & n14839;
  assign n14842 = ~n14840 & ~n14841;
  assign n14843 = ~n14478 & ~n14841;
  assign n14844 = ~n14840 & n14843;
  assign n14845 = ~n14478 & n14842;
  assign n14846 = n14478 & ~n14842;
  assign n14847 = ~n14478 & ~n40158;
  assign n14848 = ~n14840 & ~n40158;
  assign n14849 = ~n14841 & n14848;
  assign n14850 = ~n14847 & ~n14849;
  assign n14851 = ~n40158 & ~n14846;
  assign n14852 = ~n14477 & ~n40159;
  assign n14853 = n14477 & n40159;
  assign n14854 = ~n40159 & ~n14852;
  assign n14855 = n14477 & ~n40159;
  assign n14856 = ~n14477 & ~n14852;
  assign n14857 = ~n14477 & n40159;
  assign n14858 = ~n40160 & ~n40161;
  assign n14859 = ~n14852 & ~n14853;
  assign n14860 = ~n12976 & ~n40162;
  assign n14861 = n12976 & n40162;
  assign n14862 = ~n12976 & n40162;
  assign n14863 = n12976 & ~n40162;
  assign n14864 = ~n14862 & ~n14863;
  assign n14865 = ~n14860 & ~n14861;
  assign n14866 = ~n14462 & ~n40163;
  assign n14867 = n14462 & n40163;
  assign n14868 = ~n14866 & ~n14867;
  assign n14869 = ~n14447 & n14868;
  assign n14870 = n14447 & ~n14868;
  assign n14871 = ~n14869 & ~n14870;
  assign n14872 = n563 & n11258;
  assign n14873 = pi112  & n37482;
  assign n14874 = pi114  & n578;
  assign n14875 = pi113  & n580;
  assign n14876 = ~n14874 & ~n14875;
  assign n14877 = ~n14873 & ~n14875;
  assign n14878 = ~n14874 & n14877;
  assign n14879 = ~n14873 & n14876;
  assign n14880 = ~n14872 & n40164;
  assign n14881 = pi14  & ~n14880;
  assign n14882 = pi14  & ~n14881;
  assign n14883 = pi14  & n14880;
  assign n14884 = ~n14880 & ~n14881;
  assign n14885 = ~pi14  & ~n14880;
  assign n14886 = ~n40165 & ~n40166;
  assign n14887 = n14871 & ~n14886;
  assign n14888 = ~n14871 & n14886;
  assign n14889 = n14871 & ~n14887;
  assign n14890 = n14871 & n14886;
  assign n14891 = ~n14886 & ~n14887;
  assign n14892 = ~n14871 & ~n14886;
  assign n14893 = ~n40167 & ~n40168;
  assign n14894 = ~n14887 & ~n14888;
  assign n14895 = ~n14446 & ~n40169;
  assign n14896 = n14446 & n40169;
  assign n14897 = ~n14446 & n40169;
  assign n14898 = n14446 & ~n40169;
  assign n14899 = ~n14897 & ~n14898;
  assign n14900 = ~n14895 & ~n14896;
  assign n14901 = ~n14445 & ~n40170;
  assign n14902 = n14445 & n40170;
  assign n14903 = ~n14901 & ~n14902;
  assign n14904 = ~n14430 & n14903;
  assign n14905 = n14430 & ~n14903;
  assign n14906 = ~n14904 & ~n14905;
  assign n14907 = ~n13023 & ~n13025;
  assign n14908 = ~pi119  & ~pi120 ;
  assign n14909 = pi119  & pi120 ;
  assign n14910 = ~n14908 & ~n14909;
  assign n14911 = ~n14907 & n14910;
  assign n14912 = n14907 & ~n14910;
  assign n14913 = ~n14911 & ~n14912;
  assign n14914 = n13010 & n14913;
  assign n14915 = pi118  & n39810;
  assign n14916 = pi120  & n13040;
  assign n14917 = pi119  & n13042;
  assign n14918 = ~n14916 & ~n14917;
  assign n14919 = ~n14915 & ~n14917;
  assign n14920 = ~n14916 & n14919;
  assign n14921 = ~n14915 & n14918;
  assign n14922 = ~n14914 & n40171;
  assign n14923 = pi8  & ~n14922;
  assign n14924 = pi8  & ~n14923;
  assign n14925 = pi8  & n14922;
  assign n14926 = ~n14922 & ~n14923;
  assign n14927 = ~pi8  & ~n14922;
  assign n14928 = ~n40172 & ~n40173;
  assign n14929 = ~n14906 & n14928;
  assign n14930 = n14906 & ~n14928;
  assign n14931 = ~n14929 & ~n14930;
  assign n14932 = pi2  & ~pi3 ;
  assign n14933 = ~pi2  & pi3 ;
  assign n14934 = ~pi2  & ~pi3 ;
  assign n14935 = pi2  & pi3 ;
  assign n14936 = ~n14934 & ~n14935;
  assign n14937 = ~n14932 & ~n14933;
  assign n14938 = pi4  & ~pi5 ;
  assign n14939 = ~pi4  & pi5 ;
  assign n14940 = ~pi4  & ~pi5 ;
  assign n14941 = pi4  & pi5 ;
  assign n14942 = ~n14940 & ~n14941;
  assign n14943 = ~n14938 & ~n14939;
  assign n14944 = n40174 & n40175;
  assign n14945 = pi121  & pi122 ;
  assign n14946 = pi120  & pi121 ;
  assign n14947 = ~n14909 & ~n14911;
  assign n14948 = ~pi120  & ~pi121 ;
  assign n14949 = ~n14946 & ~n14948;
  assign n14950 = ~n14947 & n14949;
  assign n14951 = ~n14946 & ~n14950;
  assign n14952 = ~pi121  & ~pi122 ;
  assign n14953 = ~n14945 & ~n14952;
  assign n14954 = ~n14951 & n14953;
  assign n14955 = ~n14945 & ~n14954;
  assign n14956 = ~pi122  & ~pi123 ;
  assign n14957 = pi122  & pi123 ;
  assign n14958 = ~n14956 & ~n14957;
  assign n14959 = ~n14955 & n14958;
  assign n14960 = n14955 & ~n14958;
  assign n14961 = ~n14959 & ~n14960;
  assign n14962 = n14944 & n14961;
  assign n14963 = pi3  & ~pi4 ;
  assign n14964 = ~pi3  & pi4 ;
  assign n14965 = ~pi3  & ~pi4 ;
  assign n14966 = pi3  & pi4 ;
  assign n14967 = ~n14965 & ~n14966;
  assign n14968 = ~n14963 & ~n14964;
  assign n14969 = ~n40174 & n40175;
  assign n14970 = ~n40174 & ~n40176;
  assign n14971 = n40175 & n14970;
  assign n14972 = ~n40176 & n14969;
  assign n14973 = pi121  & n40177;
  assign n14974 = n40174 & ~n40175;
  assign n14975 = pi123  & n14974;
  assign n14976 = ~n40174 & n40176;
  assign n14977 = pi122  & n14976;
  assign n14978 = ~n14975 & ~n14977;
  assign n14979 = ~n14973 & ~n14977;
  assign n14980 = ~n14975 & n14979;
  assign n14981 = ~n14973 & n14978;
  assign n14982 = ~n14962 & n40178;
  assign n14983 = pi5  & ~n14982;
  assign n14984 = pi5  & ~n14983;
  assign n14985 = pi5  & n14982;
  assign n14986 = ~n14982 & ~n14983;
  assign n14987 = ~pi5  & ~n14982;
  assign n14988 = ~n40179 & ~n40180;
  assign n14989 = ~n14931 & n14988;
  assign n14990 = n14931 & ~n14988;
  assign n14991 = n14931 & ~n14990;
  assign n14992 = ~n14988 & ~n14990;
  assign n14993 = ~n14991 & ~n14992;
  assign n14994 = ~n14989 & ~n14990;
  assign n14995 = n14429 & n40181;
  assign n14996 = ~n14429 & ~n40181;
  assign n14997 = ~n14995 & ~n14996;
  assign n14998 = pi1  & ~pi2 ;
  assign n14999 = ~pi1  & pi2 ;
  assign n15000 = ~pi1  & ~pi2 ;
  assign n15001 = pi1  & pi2 ;
  assign n15002 = ~n15000 & ~n15001;
  assign n15003 = ~n14998 & ~n14999;
  assign n15004 = pi0  & n40182;
  assign n15005 = pi124  & pi125 ;
  assign n15006 = pi123  & pi124 ;
  assign n15007 = ~n14957 & ~n14959;
  assign n15008 = ~pi123  & ~pi124 ;
  assign n15009 = ~n15006 & ~n15008;
  assign n15010 = ~n15007 & n15009;
  assign n15011 = ~n15006 & ~n15010;
  assign n15012 = ~pi124  & ~pi125 ;
  assign n15013 = ~n15005 & ~n15012;
  assign n15014 = ~n15011 & n15013;
  assign n15015 = ~n15005 & ~n15014;
  assign n15016 = ~pi125  & ~pi126 ;
  assign n15017 = pi125  & pi126 ;
  assign n15018 = ~n15016 & ~n15017;
  assign n15019 = ~n15015 & n15018;
  assign n15020 = n15015 & ~n15018;
  assign n15021 = ~n15019 & ~n15020;
  assign n15022 = n15004 & n15021;
  assign n15023 = pi0  & ~n40182;
  assign n15024 = pi126  & n15023;
  assign n15025 = ~pi0  & ~pi1 ;
  assign n15026 = ~pi0  & n40182;
  assign n15027 = ~pi1  & n15026;
  assign n15028 = n40182 & n15025;
  assign n15029 = pi124  & n40183;
  assign n15030 = ~pi0  & pi1 ;
  assign n15031 = pi125  & n15030;
  assign n15032 = ~n15029 & ~n15031;
  assign n15033 = ~n15024 & ~n15031;
  assign n15034 = ~n15029 & n15033;
  assign n15035 = ~n15024 & n15032;
  assign n15036 = ~n15022 & n40184;
  assign n15037 = pi2  & ~n15036;
  assign n15038 = pi2  & ~n15037;
  assign n15039 = pi2  & n15036;
  assign n15040 = ~n15036 & ~n15037;
  assign n15041 = ~pi2  & ~n15036;
  assign n15042 = ~n40185 & ~n40186;
  assign n15043 = ~n14997 & n15042;
  assign n15044 = n14997 & ~n15042;
  assign n15045 = ~n15043 & ~n15044;
  assign n15046 = n14420 & n40076;
  assign n15047 = ~n14428 & ~n15046;
  assign n15048 = n14951 & ~n14953;
  assign n15049 = ~n14954 & ~n15048;
  assign n15050 = n14944 & n15049;
  assign n15051 = pi120  & n40177;
  assign n15052 = pi122  & n14974;
  assign n15053 = pi121  & n14976;
  assign n15054 = ~n15052 & ~n15053;
  assign n15055 = ~n15051 & ~n15053;
  assign n15056 = ~n15052 & n15055;
  assign n15057 = ~n15051 & n15054;
  assign n15058 = ~n15050 & n40187;
  assign n15059 = pi5  & ~n15058;
  assign n15060 = pi5  & ~n15059;
  assign n15061 = pi5  & n15058;
  assign n15062 = ~n15058 & ~n15059;
  assign n15063 = ~pi5  & ~n15058;
  assign n15064 = ~n40188 & ~n40189;
  assign n15065 = n15047 & ~n15064;
  assign n15066 = ~n15047 & n15064;
  assign n15067 = n15011 & ~n15013;
  assign n15068 = ~n15014 & ~n15067;
  assign n15069 = n15004 & n15068;
  assign n15070 = pi125  & n15023;
  assign n15071 = pi123  & n40183;
  assign n15072 = pi124  & n15030;
  assign n15073 = ~n15071 & ~n15072;
  assign n15074 = ~n15070 & ~n15072;
  assign n15075 = ~n15071 & n15074;
  assign n15076 = ~n15070 & n15073;
  assign n15077 = ~n15069 & n40190;
  assign n15078 = pi2  & ~n15077;
  assign n15079 = pi2  & ~n15078;
  assign n15080 = pi2  & n15077;
  assign n15081 = ~n15077 & ~n15078;
  assign n15082 = ~pi2  & ~n15077;
  assign n15083 = ~n40191 & ~n40192;
  assign n15084 = ~n15066 & ~n15083;
  assign n15085 = ~n15065 & ~n15066;
  assign n15086 = ~n15083 & n15085;
  assign n15087 = ~n15065 & ~n15086;
  assign n15088 = ~n15065 & ~n15084;
  assign n15089 = n15045 & ~n40193;
  assign n15090 = n14947 & ~n14949;
  assign n15091 = ~n14950 & ~n15090;
  assign n15092 = n14944 & n15091;
  assign n15093 = pi119  & n40177;
  assign n15094 = pi121  & n14974;
  assign n15095 = pi120  & n14976;
  assign n15096 = ~n15094 & ~n15095;
  assign n15097 = ~n15093 & ~n15095;
  assign n15098 = ~n15094 & n15097;
  assign n15099 = ~n15093 & n15096;
  assign n15100 = ~n15092 & n40194;
  assign n15101 = pi5  & ~n15100;
  assign n15102 = pi5  & ~n15101;
  assign n15103 = pi5  & n15100;
  assign n15104 = ~n15100 & ~n15101;
  assign n15105 = ~pi5  & ~n15100;
  assign n15106 = ~n40195 & ~n40196;
  assign n15107 = n14416 & ~n14418;
  assign n15108 = ~n14419 & ~n15107;
  assign n15109 = ~n15106 & n15108;
  assign n15110 = n15007 & ~n15009;
  assign n15111 = ~n15010 & ~n15110;
  assign n15112 = n15004 & n15111;
  assign n15113 = pi124  & n15023;
  assign n15114 = pi122  & n40183;
  assign n15115 = pi123  & n15030;
  assign n15116 = ~n15114 & ~n15115;
  assign n15117 = ~n15113 & ~n15115;
  assign n15118 = ~n15114 & n15117;
  assign n15119 = ~n15113 & n15116;
  assign n15120 = ~n15112 & n40197;
  assign n15121 = pi2  & ~n15120;
  assign n15122 = pi2  & ~n15121;
  assign n15123 = pi2  & n15120;
  assign n15124 = ~n15120 & ~n15121;
  assign n15125 = ~pi2  & ~n15120;
  assign n15126 = ~n40198 & ~n40199;
  assign n15127 = n15106 & ~n15108;
  assign n15128 = ~n15109 & ~n15127;
  assign n15129 = ~n15126 & n15128;
  assign n15130 = ~n15109 & ~n15129;
  assign n15131 = n15083 & ~n15085;
  assign n15132 = n15085 & ~n15086;
  assign n15133 = ~n15083 & ~n15086;
  assign n15134 = ~n15132 & ~n15133;
  assign n15135 = ~n15086 & ~n15131;
  assign n15136 = ~n15130 & ~n40200;
  assign n15137 = n15130 & n40200;
  assign n15138 = ~n15136 & ~n15137;
  assign n15139 = n15126 & ~n15128;
  assign n15140 = ~n15129 & ~n15139;
  assign n15141 = n14913 & n14944;
  assign n15142 = pi118  & n40177;
  assign n15143 = pi120  & n14974;
  assign n15144 = pi119  & n14976;
  assign n15145 = ~n15143 & ~n15144;
  assign n15146 = ~n15142 & ~n15144;
  assign n15147 = ~n15143 & n15146;
  assign n15148 = ~n15142 & n15145;
  assign n15149 = ~n15141 & n40201;
  assign n15150 = pi5  & ~n15149;
  assign n15151 = pi5  & ~n15150;
  assign n15152 = pi5  & n15149;
  assign n15153 = ~n15149 & ~n15150;
  assign n15154 = ~pi5  & ~n15149;
  assign n15155 = ~n40202 & ~n40203;
  assign n15156 = n14407 & n40073;
  assign n15157 = ~n14407 & ~n14415;
  assign n15158 = ~n14407 & n40073;
  assign n15159 = ~n40073 & ~n14415;
  assign n15160 = n14407 & ~n40073;
  assign n15161 = ~n40204 & ~n40205;
  assign n15162 = ~n14415 & ~n15156;
  assign n15163 = n15155 & n40206;
  assign n15164 = n14961 & n15004;
  assign n15165 = pi123  & n15023;
  assign n15166 = pi121  & n40183;
  assign n15167 = pi122  & n15030;
  assign n15168 = ~n15166 & ~n15167;
  assign n15169 = ~n15165 & ~n15167;
  assign n15170 = ~n15166 & n15169;
  assign n15171 = ~n15165 & n15168;
  assign n15172 = ~n15164 & n40207;
  assign n15173 = pi2  & ~n15172;
  assign n15174 = pi2  & ~n15173;
  assign n15175 = pi2  & n15172;
  assign n15176 = ~n15172 & ~n15173;
  assign n15177 = ~pi2  & ~n15172;
  assign n15178 = ~n40208 & ~n40209;
  assign n15179 = ~n15155 & ~n40206;
  assign n15180 = n15178 & ~n15179;
  assign n15181 = ~n40206 & ~n15179;
  assign n15182 = ~n15155 & ~n15179;
  assign n15183 = ~n15181 & ~n15182;
  assign n15184 = ~n15163 & ~n15179;
  assign n15185 = ~n15178 & ~n40210;
  assign n15186 = ~n15179 & ~n15185;
  assign n15187 = ~n15163 & ~n15180;
  assign n15188 = n15140 & ~n40211;
  assign n15189 = n13027 & n14944;
  assign n15190 = pi117  & n40177;
  assign n15191 = pi119  & n14974;
  assign n15192 = pi118  & n14976;
  assign n15193 = ~n15191 & ~n15192;
  assign n15194 = ~n15190 & ~n15192;
  assign n15195 = ~n15191 & n15194;
  assign n15196 = ~n15190 & n15193;
  assign n15197 = ~n15189 & n40212;
  assign n15198 = pi5  & ~n15197;
  assign n15199 = pi5  & ~n15198;
  assign n15200 = pi5  & n15197;
  assign n15201 = ~n15197 & ~n15198;
  assign n15202 = ~pi5  & ~n15197;
  assign n15203 = ~n40213 & ~n40214;
  assign n15204 = n14403 & ~n14405;
  assign n15205 = ~n14406 & ~n15204;
  assign n15206 = ~n15203 & n15205;
  assign n15207 = n13057 & n14944;
  assign n15208 = pi116  & n40177;
  assign n15209 = pi118  & n14974;
  assign n15210 = pi117  & n14976;
  assign n15211 = ~n15209 & ~n15210;
  assign n15212 = ~n15208 & ~n15210;
  assign n15213 = ~n15209 & n15212;
  assign n15214 = ~n15208 & n15211;
  assign n15215 = ~n15207 & n40215;
  assign n15216 = pi5  & ~n15215;
  assign n15217 = pi5  & ~n15216;
  assign n15218 = pi5  & n15215;
  assign n15219 = ~n15215 & ~n15216;
  assign n15220 = ~pi5  & ~n15215;
  assign n15221 = ~n40216 & ~n40217;
  assign n15222 = n14394 & ~n40069;
  assign n15223 = ~n40068 & n15222;
  assign n15224 = n14394 & n40070;
  assign n15225 = ~n14402 & ~n40218;
  assign n15226 = ~n15221 & n15225;
  assign n15227 = n13079 & n14944;
  assign n15228 = pi115  & n40177;
  assign n15229 = pi117  & n14974;
  assign n15230 = pi116  & n14976;
  assign n15231 = ~n15229 & ~n15230;
  assign n15232 = ~n15228 & ~n15230;
  assign n15233 = ~n15229 & n15232;
  assign n15234 = ~n15228 & n15231;
  assign n15235 = ~n15227 & n40219;
  assign n15236 = pi5  & ~n15235;
  assign n15237 = pi5  & ~n15236;
  assign n15238 = pi5  & n15235;
  assign n15239 = ~n15235 & ~n15236;
  assign n15240 = ~pi5  & ~n15235;
  assign n15241 = ~n40220 & ~n40221;
  assign n15242 = n14385 & n40067;
  assign n15243 = ~n14385 & ~n14393;
  assign n15244 = ~n14385 & n40067;
  assign n15245 = ~n40067 & ~n14393;
  assign n15246 = n14385 & ~n40067;
  assign n15247 = ~n40222 & ~n40223;
  assign n15248 = ~n14393 & ~n15242;
  assign n15249 = ~n15241 & ~n40224;
  assign n15250 = n14381 & ~n14383;
  assign n15251 = ~n14384 & ~n15250;
  assign n15252 = n12530 & n14944;
  assign n15253 = pi114  & n40177;
  assign n15254 = pi116  & n14974;
  assign n15255 = pi115  & n14976;
  assign n15256 = ~n15254 & ~n15255;
  assign n15257 = ~n15253 & ~n15255;
  assign n15258 = ~n15254 & n15257;
  assign n15259 = ~n15253 & n15256;
  assign n15260 = ~n15252 & n40225;
  assign n15261 = pi5  & ~n15260;
  assign n15262 = pi5  & ~n15261;
  assign n15263 = pi5  & n15260;
  assign n15264 = ~n15260 & ~n15261;
  assign n15265 = ~pi5  & ~n15260;
  assign n15266 = ~n40226 & ~n40227;
  assign n15267 = n15251 & ~n15266;
  assign n15268 = n14372 & n40064;
  assign n15269 = ~n14380 & ~n15268;
  assign n15270 = n523 & n14944;
  assign n15271 = pi113  & n40177;
  assign n15272 = pi115  & n14974;
  assign n15273 = pi114  & n14976;
  assign n15274 = ~n15272 & ~n15273;
  assign n15275 = ~n15271 & ~n15273;
  assign n15276 = ~n15272 & n15275;
  assign n15277 = ~n15271 & n15274;
  assign n15278 = ~n15270 & n40228;
  assign n15279 = pi5  & ~n15278;
  assign n15280 = pi5  & ~n15279;
  assign n15281 = pi5  & n15278;
  assign n15282 = ~n15278 & ~n15279;
  assign n15283 = ~pi5  & ~n15278;
  assign n15284 = ~n40229 & ~n40230;
  assign n15285 = n15269 & ~n15284;
  assign n15286 = n14363 & n40061;
  assign n15287 = ~n14371 & ~n15286;
  assign n15288 = n11258 & n14944;
  assign n15289 = pi112  & n40177;
  assign n15290 = pi114  & n14974;
  assign n15291 = pi113  & n14976;
  assign n15292 = ~n15290 & ~n15291;
  assign n15293 = ~n15289 & ~n15291;
  assign n15294 = ~n15290 & n15293;
  assign n15295 = ~n15289 & n15292;
  assign n15296 = ~n15288 & n40231;
  assign n15297 = pi5  & ~n15296;
  assign n15298 = pi5  & ~n15297;
  assign n15299 = pi5  & n15296;
  assign n15300 = ~n15296 & ~n15297;
  assign n15301 = ~pi5  & ~n15296;
  assign n15302 = ~n40232 & ~n40233;
  assign n15303 = n15287 & ~n15302;
  assign n15304 = n14354 & n40058;
  assign n15305 = ~n14362 & ~n15304;
  assign n15306 = n11276 & n14944;
  assign n15307 = pi111  & n40177;
  assign n15308 = pi113  & n14974;
  assign n15309 = pi112  & n14976;
  assign n15310 = ~n15308 & ~n15309;
  assign n15311 = ~n15307 & ~n15309;
  assign n15312 = ~n15308 & n15311;
  assign n15313 = ~n15307 & n15310;
  assign n15314 = ~n15306 & n40234;
  assign n15315 = pi5  & ~n15314;
  assign n15316 = pi5  & ~n15315;
  assign n15317 = pi5  & n15314;
  assign n15318 = ~n15314 & ~n15315;
  assign n15319 = ~pi5  & ~n15314;
  assign n15320 = ~n40235 & ~n40236;
  assign n15321 = n15305 & ~n15320;
  assign n15322 = n10844 & n14944;
  assign n15323 = pi110  & n40177;
  assign n15324 = pi112  & n14974;
  assign n15325 = pi111  & n14976;
  assign n15326 = ~n15324 & ~n15325;
  assign n15327 = ~n15323 & ~n15325;
  assign n15328 = ~n15324 & n15327;
  assign n15329 = ~n15323 & n15326;
  assign n15330 = ~n15322 & n40237;
  assign n15331 = pi5  & ~n15330;
  assign n15332 = pi5  & ~n15331;
  assign n15333 = pi5  & n15330;
  assign n15334 = ~n15330 & ~n15331;
  assign n15335 = ~pi5  & ~n15330;
  assign n15336 = ~n40238 & ~n40239;
  assign n15337 = n14345 & n40055;
  assign n15338 = ~n14345 & n40055;
  assign n15339 = n14345 & ~n40055;
  assign n15340 = ~n15338 & ~n15339;
  assign n15341 = ~n14353 & ~n15337;
  assign n15342 = ~n15336 & ~n40240;
  assign n15343 = n565 & n14944;
  assign n15344 = pi109  & n40177;
  assign n15345 = pi111  & n14974;
  assign n15346 = pi110  & n14976;
  assign n15347 = ~n15345 & ~n15346;
  assign n15348 = ~n15344 & ~n15346;
  assign n15349 = ~n15345 & n15348;
  assign n15350 = ~n15344 & n15347;
  assign n15351 = ~n15343 & n40241;
  assign n15352 = pi5  & ~n15351;
  assign n15353 = pi5  & ~n15352;
  assign n15354 = pi5  & n15351;
  assign n15355 = ~n15351 & ~n15352;
  assign n15356 = ~pi5  & ~n15351;
  assign n15357 = ~n40242 & ~n40243;
  assign n15358 = n14339 & ~n14341;
  assign n15359 = ~n14339 & ~n40052;
  assign n15360 = ~n14340 & n14345;
  assign n15361 = ~n15359 & ~n15360;
  assign n15362 = ~n40052 & ~n15358;
  assign n15363 = ~n15357 & ~n40244;
  assign n15364 = n14330 & n40051;
  assign n15365 = ~n14338 & ~n15364;
  assign n15366 = n9678 & n14944;
  assign n15367 = pi108  & n40177;
  assign n15368 = pi110  & n14974;
  assign n15369 = pi109  & n14976;
  assign n15370 = ~n15368 & ~n15369;
  assign n15371 = ~n15367 & ~n15369;
  assign n15372 = ~n15368 & n15371;
  assign n15373 = ~n15367 & n15370;
  assign n15374 = ~n15366 & n40245;
  assign n15375 = pi5  & ~n15374;
  assign n15376 = pi5  & ~n15375;
  assign n15377 = pi5  & n15374;
  assign n15378 = ~n15374 & ~n15375;
  assign n15379 = ~pi5  & ~n15374;
  assign n15380 = ~n40246 & ~n40247;
  assign n15381 = n15365 & ~n15380;
  assign n15382 = n9701 & n14944;
  assign n15383 = pi107  & n40177;
  assign n15384 = pi109  & n14974;
  assign n15385 = pi108  & n14976;
  assign n15386 = ~n15384 & ~n15385;
  assign n15387 = ~n15383 & ~n15385;
  assign n15388 = ~n15384 & n15387;
  assign n15389 = ~n15383 & n15386;
  assign n15390 = ~n15382 & n40248;
  assign n15391 = pi5  & ~n15390;
  assign n15392 = pi5  & ~n15391;
  assign n15393 = pi5  & n15390;
  assign n15394 = ~n15390 & ~n15391;
  assign n15395 = ~pi5  & ~n15390;
  assign n15396 = ~n40249 & ~n40250;
  assign n15397 = n14321 & n40048;
  assign n15398 = ~n14321 & n40048;
  assign n15399 = n14321 & ~n40048;
  assign n15400 = ~n15398 & ~n15399;
  assign n15401 = ~n14329 & ~n15397;
  assign n15402 = ~n15396 & ~n40251;
  assign n15403 = n9277 & n14944;
  assign n15404 = pi106  & n40177;
  assign n15405 = pi108  & n14974;
  assign n15406 = pi107  & n14976;
  assign n15407 = ~n15405 & ~n15406;
  assign n15408 = ~n15404 & ~n15406;
  assign n15409 = ~n15405 & n15408;
  assign n15410 = ~n15404 & n15407;
  assign n15411 = ~n15403 & n40252;
  assign n15412 = pi5  & ~n15411;
  assign n15413 = pi5  & ~n15412;
  assign n15414 = pi5  & n15411;
  assign n15415 = ~n15411 & ~n15412;
  assign n15416 = ~pi5  & ~n15411;
  assign n15417 = ~n40253 & ~n40254;
  assign n15418 = n14315 & ~n14317;
  assign n15419 = ~n14315 & ~n40045;
  assign n15420 = ~n14316 & n14321;
  assign n15421 = ~n15419 & ~n15420;
  assign n15422 = ~n40045 & ~n15418;
  assign n15423 = ~n15417 & ~n40255;
  assign n15424 = n8177 & n14944;
  assign n15425 = pi105  & n40177;
  assign n15426 = pi107  & n14974;
  assign n15427 = pi106  & n14976;
  assign n15428 = ~n15426 & ~n15427;
  assign n15429 = ~n15425 & ~n15427;
  assign n15430 = ~n15426 & n15429;
  assign n15431 = ~n15425 & n15428;
  assign n15432 = ~n15424 & n40256;
  assign n15433 = pi5  & ~n15432;
  assign n15434 = pi5  & ~n15433;
  assign n15435 = pi5  & n15432;
  assign n15436 = ~n15432 & ~n15433;
  assign n15437 = ~pi5  & ~n15432;
  assign n15438 = ~n40257 & ~n40258;
  assign n15439 = n14309 & ~n14311;
  assign n15440 = ~n14309 & ~n40044;
  assign n15441 = ~n14310 & n14315;
  assign n15442 = ~n15440 & ~n15441;
  assign n15443 = ~n40044 & ~n15439;
  assign n15444 = ~n15438 & ~n40259;
  assign n15445 = n14300 & n40043;
  assign n15446 = ~n14308 & ~n15445;
  assign n15447 = n8209 & n14944;
  assign n15448 = pi104  & n40177;
  assign n15449 = pi106  & n14974;
  assign n15450 = pi105  & n14976;
  assign n15451 = ~n15449 & ~n15450;
  assign n15452 = ~n15448 & ~n15450;
  assign n15453 = ~n15449 & n15452;
  assign n15454 = ~n15448 & n15451;
  assign n15455 = ~n15447 & n40260;
  assign n15456 = pi5  & ~n15455;
  assign n15457 = pi5  & ~n15456;
  assign n15458 = pi5  & n15455;
  assign n15459 = ~n15455 & ~n15456;
  assign n15460 = ~pi5  & ~n15455;
  assign n15461 = ~n40261 & ~n40262;
  assign n15462 = n15446 & ~n15461;
  assign n15463 = n8229 & n14944;
  assign n15464 = pi103  & n40177;
  assign n15465 = pi105  & n14974;
  assign n15466 = pi104  & n14976;
  assign n15467 = ~n15465 & ~n15466;
  assign n15468 = ~n15464 & ~n15466;
  assign n15469 = ~n15465 & n15468;
  assign n15470 = ~n15464 & n15467;
  assign n15471 = ~n15463 & n40263;
  assign n15472 = pi5  & ~n15471;
  assign n15473 = pi5  & ~n15472;
  assign n15474 = pi5  & n15471;
  assign n15475 = ~n15471 & ~n15472;
  assign n15476 = ~pi5  & ~n15471;
  assign n15477 = ~n40264 & ~n40265;
  assign n15478 = n14291 & n40040;
  assign n15479 = ~n14299 & ~n15478;
  assign n15480 = ~n15477 & n15479;
  assign n15481 = n8136 & n14944;
  assign n15482 = pi102  & n40177;
  assign n15483 = pi104  & n14974;
  assign n15484 = pi103  & n14976;
  assign n15485 = ~n15483 & ~n15484;
  assign n15486 = ~n15482 & ~n15484;
  assign n15487 = ~n15483 & n15486;
  assign n15488 = ~n15482 & n15485;
  assign n15489 = ~n15481 & n40266;
  assign n15490 = pi5  & ~n15489;
  assign n15491 = pi5  & ~n15490;
  assign n15492 = pi5  & n15489;
  assign n15493 = ~n15489 & ~n15490;
  assign n15494 = ~pi5  & ~n15489;
  assign n15495 = ~n40267 & ~n40268;
  assign n15496 = n14285 & ~n14287;
  assign n15497 = ~n14285 & ~n40037;
  assign n15498 = ~n14286 & n14291;
  assign n15499 = ~n15497 & ~n15498;
  assign n15500 = ~n40037 & ~n15496;
  assign n15501 = ~n15495 & ~n40269;
  assign n15502 = n6787 & n14944;
  assign n15503 = pi101  & n40177;
  assign n15504 = pi103  & n14974;
  assign n15505 = pi102  & n14976;
  assign n15506 = ~n15504 & ~n15505;
  assign n15507 = ~n15503 & ~n15505;
  assign n15508 = ~n15504 & n15507;
  assign n15509 = ~n15503 & n15506;
  assign n15510 = ~n15502 & n40270;
  assign n15511 = pi5  & ~n15510;
  assign n15512 = pi5  & ~n15511;
  assign n15513 = pi5  & n15510;
  assign n15514 = ~n15510 & ~n15511;
  assign n15515 = ~pi5  & ~n15510;
  assign n15516 = ~n40271 & ~n40272;
  assign n15517 = n14281 & ~n14283;
  assign n15518 = ~n14284 & ~n15517;
  assign n15519 = ~n15516 & n15518;
  assign n15520 = n6819 & n14944;
  assign n15521 = pi100  & n40177;
  assign n15522 = pi102  & n14974;
  assign n15523 = pi101  & n14976;
  assign n15524 = ~n15522 & ~n15523;
  assign n15525 = ~n15521 & ~n15523;
  assign n15526 = ~n15522 & n15525;
  assign n15527 = ~n15521 & n15524;
  assign n15528 = ~n15520 & n40273;
  assign n15529 = pi5  & ~n15528;
  assign n15530 = pi5  & ~n15529;
  assign n15531 = pi5  & n15528;
  assign n15532 = ~n15528 & ~n15529;
  assign n15533 = ~pi5  & ~n15528;
  assign n15534 = ~n40274 & ~n40275;
  assign n15535 = n14272 & n40036;
  assign n15536 = ~n14272 & n40036;
  assign n15537 = n14272 & ~n40036;
  assign n15538 = ~n15536 & ~n15537;
  assign n15539 = ~n14280 & ~n15535;
  assign n15540 = ~n15534 & ~n40276;
  assign n15541 = n14268 & ~n14270;
  assign n15542 = ~n14271 & ~n15541;
  assign n15543 = n6839 & n14944;
  assign n15544 = pi99  & n40177;
  assign n15545 = pi101  & n14974;
  assign n15546 = pi100  & n14976;
  assign n15547 = ~n15545 & ~n15546;
  assign n15548 = ~n15544 & ~n15546;
  assign n15549 = ~n15545 & n15548;
  assign n15550 = ~n15544 & n15547;
  assign n15551 = ~n15543 & n40277;
  assign n15552 = pi5  & ~n15551;
  assign n15553 = pi5  & ~n15552;
  assign n15554 = pi5  & n15551;
  assign n15555 = ~n15551 & ~n15552;
  assign n15556 = ~pi5  & ~n15551;
  assign n15557 = ~n40278 & ~n40279;
  assign n15558 = n15542 & ~n15557;
  assign n15559 = n6474 & n14944;
  assign n15560 = pi98  & n40177;
  assign n15561 = pi100  & n14974;
  assign n15562 = pi99  & n14976;
  assign n15563 = ~n15561 & ~n15562;
  assign n15564 = ~n15560 & ~n15562;
  assign n15565 = ~n15561 & n15564;
  assign n15566 = ~n15560 & n15563;
  assign n15567 = ~n15559 & n40280;
  assign n15568 = pi5  & ~n15567;
  assign n15569 = pi5  & ~n15568;
  assign n15570 = pi5  & n15567;
  assign n15571 = ~n15567 & ~n15568;
  assign n15572 = ~pi5  & ~n15567;
  assign n15573 = ~n40281 & ~n40282;
  assign n15574 = n14259 & n40033;
  assign n15575 = ~n14259 & n40033;
  assign n15576 = n14259 & ~n40033;
  assign n15577 = ~n15575 & ~n15576;
  assign n15578 = ~n14267 & ~n15574;
  assign n15579 = ~n15573 & ~n40283;
  assign n15580 = n5578 & n14944;
  assign n15581 = pi97  & n40177;
  assign n15582 = pi99  & n14974;
  assign n15583 = pi98  & n14976;
  assign n15584 = ~n15582 & ~n15583;
  assign n15585 = ~n15581 & ~n15583;
  assign n15586 = ~n15582 & n15585;
  assign n15587 = ~n15581 & n15584;
  assign n15588 = ~n15580 & n40284;
  assign n15589 = pi5  & ~n15588;
  assign n15590 = pi5  & ~n15589;
  assign n15591 = pi5  & n15588;
  assign n15592 = ~n15588 & ~n15589;
  assign n15593 = ~pi5  & ~n15588;
  assign n15594 = ~n40285 & ~n40286;
  assign n15595 = n14255 & ~n14257;
  assign n15596 = ~n14258 & ~n15595;
  assign n15597 = ~n15594 & n15596;
  assign n15598 = n14251 & ~n14253;
  assign n15599 = ~n14254 & ~n15598;
  assign n15600 = n5610 & n14944;
  assign n15601 = pi96  & n40177;
  assign n15602 = pi98  & n14974;
  assign n15603 = pi97  & n14976;
  assign n15604 = ~n15602 & ~n15603;
  assign n15605 = ~n15601 & ~n15603;
  assign n15606 = ~n15602 & n15605;
  assign n15607 = ~n15601 & n15604;
  assign n15608 = ~n15600 & n40287;
  assign n15609 = pi5  & ~n15608;
  assign n15610 = pi5  & ~n15609;
  assign n15611 = pi5  & n15608;
  assign n15612 = ~n15608 & ~n15609;
  assign n15613 = ~pi5  & ~n15608;
  assign n15614 = ~n40288 & ~n40289;
  assign n15615 = n15599 & ~n15614;
  assign n15616 = n5630 & n14944;
  assign n15617 = pi95  & n40177;
  assign n15618 = pi97  & n14974;
  assign n15619 = pi96  & n14976;
  assign n15620 = ~n15618 & ~n15619;
  assign n15621 = ~n15617 & ~n15619;
  assign n15622 = ~n15618 & n15621;
  assign n15623 = ~n15617 & n15620;
  assign n15624 = ~n15616 & n40290;
  assign n15625 = pi5  & ~n15624;
  assign n15626 = pi5  & ~n15625;
  assign n15627 = pi5  & n15624;
  assign n15628 = ~n15624 & ~n15625;
  assign n15629 = ~pi5  & ~n15624;
  assign n15630 = ~n40291 & ~n40292;
  assign n15631 = n14247 & ~n14249;
  assign n15632 = ~n14250 & ~n15631;
  assign n15633 = ~n15630 & n15632;
  assign n15634 = n14238 & n40030;
  assign n15635 = ~n14246 & ~n15634;
  assign n15636 = n5281 & n14944;
  assign n15637 = pi94  & n40177;
  assign n15638 = pi96  & n14974;
  assign n15639 = pi95  & n14976;
  assign n15640 = ~n15638 & ~n15639;
  assign n15641 = ~n15637 & ~n15639;
  assign n15642 = ~n15638 & n15641;
  assign n15643 = ~n15637 & n15640;
  assign n15644 = ~n15636 & n40293;
  assign n15645 = pi5  & ~n15644;
  assign n15646 = pi5  & ~n15645;
  assign n15647 = pi5  & n15644;
  assign n15648 = ~n15644 & ~n15645;
  assign n15649 = ~pi5  & ~n15644;
  assign n15650 = ~n40294 & ~n40295;
  assign n15651 = n15635 & ~n15650;
  assign n15652 = n14229 & n40027;
  assign n15653 = ~n14237 & ~n15652;
  assign n15654 = n4494 & n14944;
  assign n15655 = pi93  & n40177;
  assign n15656 = pi95  & n14974;
  assign n15657 = pi94  & n14976;
  assign n15658 = ~n15656 & ~n15657;
  assign n15659 = ~n15655 & ~n15657;
  assign n15660 = ~n15656 & n15659;
  assign n15661 = ~n15655 & n15658;
  assign n15662 = ~n15654 & n40296;
  assign n15663 = pi5  & ~n15662;
  assign n15664 = pi5  & ~n15663;
  assign n15665 = pi5  & n15662;
  assign n15666 = ~n15662 & ~n15663;
  assign n15667 = ~pi5  & ~n15662;
  assign n15668 = ~n40297 & ~n40298;
  assign n15669 = n15653 & ~n15668;
  assign n15670 = n14220 & n40024;
  assign n15671 = ~n14228 & ~n15670;
  assign n15672 = n4524 & n14944;
  assign n15673 = pi92  & n40177;
  assign n15674 = pi94  & n14974;
  assign n15675 = pi93  & n14976;
  assign n15676 = ~n15674 & ~n15675;
  assign n15677 = ~n15673 & ~n15675;
  assign n15678 = ~n15674 & n15677;
  assign n15679 = ~n15673 & n15676;
  assign n15680 = ~n15672 & n40299;
  assign n15681 = pi5  & ~n15680;
  assign n15682 = pi5  & ~n15681;
  assign n15683 = pi5  & n15680;
  assign n15684 = ~n15680 & ~n15681;
  assign n15685 = ~pi5  & ~n15680;
  assign n15686 = ~n40300 & ~n40301;
  assign n15687 = n15671 & ~n15686;
  assign n15688 = n14211 & n40021;
  assign n15689 = ~n14219 & ~n15688;
  assign n15690 = n4544 & n14944;
  assign n15691 = pi91  & n40177;
  assign n15692 = pi93  & n14974;
  assign n15693 = pi92  & n14976;
  assign n15694 = ~n15692 & ~n15693;
  assign n15695 = ~n15691 & ~n15693;
  assign n15696 = ~n15692 & n15695;
  assign n15697 = ~n15691 & n15694;
  assign n15698 = ~n15690 & n40302;
  assign n15699 = pi5  & ~n15698;
  assign n15700 = pi5  & ~n15699;
  assign n15701 = pi5  & n15698;
  assign n15702 = ~n15698 & ~n15699;
  assign n15703 = ~pi5  & ~n15698;
  assign n15704 = ~n40303 & ~n40304;
  assign n15705 = n15689 & ~n15704;
  assign n15706 = n14202 & n40018;
  assign n15707 = ~n14210 & ~n15706;
  assign n15708 = n4453 & n14944;
  assign n15709 = pi90  & n40177;
  assign n15710 = pi92  & n14974;
  assign n15711 = pi91  & n14976;
  assign n15712 = ~n15710 & ~n15711;
  assign n15713 = ~n15709 & ~n15711;
  assign n15714 = ~n15710 & n15713;
  assign n15715 = ~n15709 & n15712;
  assign n15716 = ~n15708 & n40305;
  assign n15717 = pi5  & ~n15716;
  assign n15718 = pi5  & ~n15717;
  assign n15719 = pi5  & n15716;
  assign n15720 = ~n15716 & ~n15717;
  assign n15721 = ~pi5  & ~n15716;
  assign n15722 = ~n40306 & ~n40307;
  assign n15723 = n15707 & ~n15722;
  assign n15724 = n14198 & ~n14200;
  assign n15725 = ~n14201 & ~n15724;
  assign n15726 = n594 & n14944;
  assign n15727 = pi89  & n40177;
  assign n15728 = pi91  & n14974;
  assign n15729 = pi90  & n14976;
  assign n15730 = ~n15728 & ~n15729;
  assign n15731 = ~n15727 & ~n15729;
  assign n15732 = ~n15728 & n15731;
  assign n15733 = ~n15727 & n15730;
  assign n15734 = ~n15726 & n40308;
  assign n15735 = pi5  & ~n15734;
  assign n15736 = pi5  & ~n15735;
  assign n15737 = pi5  & n15734;
  assign n15738 = ~n15734 & ~n15735;
  assign n15739 = ~pi5  & ~n15734;
  assign n15740 = ~n40309 & ~n40310;
  assign n15741 = n15725 & ~n15740;
  assign n15742 = n3566 & n14944;
  assign n15743 = pi88  & n40177;
  assign n15744 = pi90  & n14974;
  assign n15745 = pi89  & n14976;
  assign n15746 = ~n15744 & ~n15745;
  assign n15747 = ~n15743 & ~n15745;
  assign n15748 = ~n15744 & n15747;
  assign n15749 = ~n15743 & n15746;
  assign n15750 = ~n15742 & n40311;
  assign n15751 = pi5  & ~n15750;
  assign n15752 = pi5  & ~n15751;
  assign n15753 = pi5  & n15750;
  assign n15754 = ~n15750 & ~n15751;
  assign n15755 = ~pi5  & ~n15750;
  assign n15756 = ~n40312 & ~n40313;
  assign n15757 = n14189 & n40015;
  assign n15758 = ~n14197 & ~n15757;
  assign n15759 = ~n15756 & n15758;
  assign n15760 = ~n13683 & n14187;
  assign n15761 = ~n14188 & ~n15760;
  assign n15762 = n3591 & n14944;
  assign n15763 = pi87  & n40177;
  assign n15764 = pi89  & n14974;
  assign n15765 = pi88  & n14976;
  assign n15766 = ~n15764 & ~n15765;
  assign n15767 = ~n15763 & ~n15765;
  assign n15768 = ~n15764 & n15767;
  assign n15769 = ~n15763 & n15766;
  assign n15770 = ~n15762 & n40314;
  assign n15771 = pi5  & ~n15770;
  assign n15772 = pi5  & ~n15771;
  assign n15773 = pi5  & n15770;
  assign n15774 = ~n15770 & ~n15771;
  assign n15775 = ~pi5  & ~n15770;
  assign n15776 = ~n40315 & ~n40316;
  assign n15777 = n15761 & ~n15776;
  assign n15778 = ~n13703 & n14185;
  assign n15779 = ~n14186 & ~n15778;
  assign n15780 = n3354 & n14944;
  assign n15781 = pi86  & n40177;
  assign n15782 = pi88  & n14974;
  assign n15783 = pi87  & n14976;
  assign n15784 = ~n15782 & ~n15783;
  assign n15785 = ~n15781 & ~n15783;
  assign n15786 = ~n15782 & n15785;
  assign n15787 = ~n15781 & n15784;
  assign n15788 = ~n15780 & n40317;
  assign n15789 = pi5  & ~n15788;
  assign n15790 = pi5  & ~n15789;
  assign n15791 = pi5  & n15788;
  assign n15792 = ~n15788 & ~n15789;
  assign n15793 = ~pi5  & ~n15788;
  assign n15794 = ~n40318 & ~n40319;
  assign n15795 = n15779 & ~n15794;
  assign n15796 = n14176 & n40012;
  assign n15797 = ~n14184 & ~n15796;
  assign n15798 = n636 & n14944;
  assign n15799 = pi85  & n40177;
  assign n15800 = pi87  & n14974;
  assign n15801 = pi86  & n14976;
  assign n15802 = ~n15800 & ~n15801;
  assign n15803 = ~n15799 & ~n15801;
  assign n15804 = ~n15800 & n15803;
  assign n15805 = ~n15799 & n15802;
  assign n15806 = ~n15798 & n40320;
  assign n15807 = pi5  & ~n15806;
  assign n15808 = pi5  & ~n15807;
  assign n15809 = pi5  & n15806;
  assign n15810 = ~n15806 & ~n15807;
  assign n15811 = ~pi5  & ~n15806;
  assign n15812 = ~n40321 & ~n40322;
  assign n15813 = n15797 & ~n15812;
  assign n15814 = n2779 & n14944;
  assign n15815 = pi84  & n40177;
  assign n15816 = pi86  & n14974;
  assign n15817 = pi85  & n14976;
  assign n15818 = ~n15816 & ~n15817;
  assign n15819 = ~n15815 & ~n15817;
  assign n15820 = ~n15816 & n15819;
  assign n15821 = ~n15815 & n15818;
  assign n15822 = ~n15814 & n40323;
  assign n15823 = pi5  & ~n15822;
  assign n15824 = pi5  & ~n15823;
  assign n15825 = pi5  & n15822;
  assign n15826 = ~n15822 & ~n15823;
  assign n15827 = ~pi5  & ~n15822;
  assign n15828 = ~n40324 & ~n40325;
  assign n15829 = n14167 & n40009;
  assign n15830 = ~n40009 & ~n14175;
  assign n15831 = n14167 & ~n40009;
  assign n15832 = ~n14167 & ~n14175;
  assign n15833 = ~n14167 & n40009;
  assign n15834 = ~n40326 & ~n40327;
  assign n15835 = ~n14175 & ~n15829;
  assign n15836 = ~n15828 & ~n40328;
  assign n15837 = n2804 & n14944;
  assign n15838 = pi83  & n40177;
  assign n15839 = pi85  & n14974;
  assign n15840 = pi84  & n14976;
  assign n15841 = ~n15839 & ~n15840;
  assign n15842 = ~n15838 & ~n15840;
  assign n15843 = ~n15839 & n15842;
  assign n15844 = ~n15838 & n15841;
  assign n15845 = ~n15837 & n40329;
  assign n15846 = pi5  & ~n15845;
  assign n15847 = pi5  & ~n15846;
  assign n15848 = pi5  & n15845;
  assign n15849 = ~n15845 & ~n15846;
  assign n15850 = ~pi5  & ~n15845;
  assign n15851 = ~n40330 & ~n40331;
  assign n15852 = n14163 & ~n14165;
  assign n15853 = ~n14166 & ~n15852;
  assign n15854 = ~n15851 & n15853;
  assign n15855 = n2591 & n14944;
  assign n15856 = pi82  & n40177;
  assign n15857 = pi84  & n14974;
  assign n15858 = pi83  & n14976;
  assign n15859 = ~n15857 & ~n15858;
  assign n15860 = ~n15856 & ~n15858;
  assign n15861 = ~n15857 & n15860;
  assign n15862 = ~n15856 & n15859;
  assign n15863 = ~n15855 & n40332;
  assign n15864 = pi5  & ~n15863;
  assign n15865 = pi5  & ~n15864;
  assign n15866 = pi5  & n15863;
  assign n15867 = ~n15863 & ~n15864;
  assign n15868 = ~pi5  & ~n15863;
  assign n15869 = ~n40333 & ~n40334;
  assign n15870 = n14154 & n40006;
  assign n15871 = ~n14154 & ~n14162;
  assign n15872 = ~n14154 & n40006;
  assign n15873 = ~n40006 & ~n14162;
  assign n15874 = n14154 & ~n40006;
  assign n15875 = ~n40335 & ~n40336;
  assign n15876 = ~n14162 & ~n15870;
  assign n15877 = ~n15869 & ~n40337;
  assign n15878 = n14150 & ~n14152;
  assign n15879 = ~n14153 & ~n15878;
  assign n15880 = n2091 & n14944;
  assign n15881 = pi81  & n40177;
  assign n15882 = pi83  & n14974;
  assign n15883 = pi82  & n14976;
  assign n15884 = ~n15882 & ~n15883;
  assign n15885 = ~n15881 & ~n15883;
  assign n15886 = ~n15882 & n15885;
  assign n15887 = ~n15881 & n15884;
  assign n15888 = ~n15880 & n40338;
  assign n15889 = pi5  & ~n15888;
  assign n15890 = pi5  & ~n15889;
  assign n15891 = pi5  & n15888;
  assign n15892 = ~n15888 & ~n15889;
  assign n15893 = ~pi5  & ~n15888;
  assign n15894 = ~n40339 & ~n40340;
  assign n15895 = n15879 & ~n15894;
  assign n15896 = n14146 & ~n14148;
  assign n15897 = ~n14149 & ~n15896;
  assign n15898 = n2134 & n14944;
  assign n15899 = pi80  & n40177;
  assign n15900 = pi82  & n14974;
  assign n15901 = pi81  & n14976;
  assign n15902 = ~n15900 & ~n15901;
  assign n15903 = ~n15899 & ~n15901;
  assign n15904 = ~n15900 & n15903;
  assign n15905 = ~n15899 & n15902;
  assign n15906 = ~n15898 & n40341;
  assign n15907 = pi5  & ~n15906;
  assign n15908 = pi5  & ~n15907;
  assign n15909 = pi5  & n15906;
  assign n15910 = ~n15906 & ~n15907;
  assign n15911 = ~pi5  & ~n15906;
  assign n15912 = ~n40342 & ~n40343;
  assign n15913 = n15897 & ~n15912;
  assign n15914 = n2154 & n14944;
  assign n15915 = pi79  & n40177;
  assign n15916 = pi81  & n14974;
  assign n15917 = pi80  & n14976;
  assign n15918 = ~n15916 & ~n15917;
  assign n15919 = ~n15915 & ~n15917;
  assign n15920 = ~n15916 & n15919;
  assign n15921 = ~n15915 & n15918;
  assign n15922 = ~n15914 & n40344;
  assign n15923 = pi5  & ~n15922;
  assign n15924 = pi5  & ~n15923;
  assign n15925 = pi5  & n15922;
  assign n15926 = ~n15922 & ~n15923;
  assign n15927 = ~pi5  & ~n15922;
  assign n15928 = ~n40345 & ~n40346;
  assign n15929 = n14137 & n40003;
  assign n15930 = ~n14145 & ~n15929;
  assign n15931 = ~n15928 & n15930;
  assign n15932 = ~n13849 & n14135;
  assign n15933 = ~n14136 & ~n15932;
  assign n15934 = n2063 & n14944;
  assign n15935 = pi78  & n40177;
  assign n15936 = pi80  & n14974;
  assign n15937 = pi79  & n14976;
  assign n15938 = ~n15936 & ~n15937;
  assign n15939 = ~n15935 & ~n15937;
  assign n15940 = ~n15936 & n15939;
  assign n15941 = ~n15935 & n15938;
  assign n15942 = ~n15934 & n40347;
  assign n15943 = pi5  & ~n15942;
  assign n15944 = pi5  & ~n15943;
  assign n15945 = pi5  & n15942;
  assign n15946 = ~n15942 & ~n15943;
  assign n15947 = ~pi5  & ~n15942;
  assign n15948 = ~n40348 & ~n40349;
  assign n15949 = n15933 & ~n15948;
  assign n15950 = n678 & n14944;
  assign n15951 = pi77  & n40177;
  assign n15952 = pi79  & n14974;
  assign n15953 = pi78  & n14976;
  assign n15954 = ~n15952 & ~n15953;
  assign n15955 = ~n15951 & ~n15953;
  assign n15956 = ~n15952 & n15955;
  assign n15957 = ~n15951 & n15954;
  assign n15958 = ~n15950 & n40350;
  assign n15959 = pi5  & ~n15958;
  assign n15960 = pi5  & ~n15959;
  assign n15961 = pi5  & n15958;
  assign n15962 = ~n15958 & ~n15959;
  assign n15963 = ~pi5  & ~n15958;
  assign n15964 = ~n40351 & ~n40352;
  assign n15965 = n14131 & ~n14133;
  assign n15966 = ~n14134 & ~n15965;
  assign n15967 = ~n15964 & n15966;
  assign n15968 = n1578 & n14944;
  assign n15969 = pi76  & n40177;
  assign n15970 = pi78  & n14974;
  assign n15971 = pi77  & n14976;
  assign n15972 = ~n15970 & ~n15971;
  assign n15973 = ~n15969 & ~n15971;
  assign n15974 = ~n15970 & n15973;
  assign n15975 = ~n15969 & n15972;
  assign n15976 = ~n15968 & n40353;
  assign n15977 = pi5  & ~n15976;
  assign n15978 = pi5  & ~n15977;
  assign n15979 = pi5  & n15976;
  assign n15980 = ~n15976 & ~n15977;
  assign n15981 = ~pi5  & ~n15976;
  assign n15982 = ~n40354 & ~n40355;
  assign n15983 = n14127 & ~n14129;
  assign n15984 = ~n14130 & ~n15983;
  assign n15985 = ~n15982 & n15984;
  assign n15986 = n1596 & n14944;
  assign n15987 = pi75  & n40177;
  assign n15988 = pi77  & n14974;
  assign n15989 = pi76  & n14976;
  assign n15990 = ~n15988 & ~n15989;
  assign n15991 = ~n15987 & ~n15989;
  assign n15992 = ~n15988 & n15991;
  assign n15993 = ~n15987 & n15990;
  assign n15994 = ~n15986 & n40356;
  assign n15995 = pi5  & ~n15994;
  assign n15996 = pi5  & ~n15995;
  assign n15997 = pi5  & n15994;
  assign n15998 = ~n15994 & ~n15995;
  assign n15999 = ~pi5  & ~n15994;
  assign n16000 = ~n40357 & ~n40358;
  assign n16001 = n14123 & ~n14125;
  assign n16002 = ~n14126 & ~n16001;
  assign n16003 = ~n16000 & n16002;
  assign n16004 = n1465 & n14944;
  assign n16005 = pi74  & n40177;
  assign n16006 = pi76  & n14974;
  assign n16007 = pi75  & n14976;
  assign n16008 = ~n16006 & ~n16007;
  assign n16009 = ~n16005 & ~n16007;
  assign n16010 = ~n16006 & n16009;
  assign n16011 = ~n16005 & n16008;
  assign n16012 = ~n16004 & n40359;
  assign n16013 = pi5  & ~n16012;
  assign n16014 = pi5  & ~n16013;
  assign n16015 = pi5  & n16012;
  assign n16016 = ~n16012 & ~n16013;
  assign n16017 = ~pi5  & ~n16012;
  assign n16018 = ~n40360 & ~n40361;
  assign n16019 = n14114 & ~n39999;
  assign n16020 = ~n39998 & n16019;
  assign n16021 = n14114 & n40000;
  assign n16022 = ~n14122 & ~n40362;
  assign n16023 = ~n16018 & n16022;
  assign n16024 = n720 & n14944;
  assign n16025 = pi73  & n40177;
  assign n16026 = pi75  & n14974;
  assign n16027 = pi74  & n14976;
  assign n16028 = ~n16026 & ~n16027;
  assign n16029 = ~n16025 & ~n16027;
  assign n16030 = ~n16026 & n16029;
  assign n16031 = ~n16025 & n16028;
  assign n16032 = ~n16024 & n40363;
  assign n16033 = pi5  & ~n16032;
  assign n16034 = pi5  & ~n16033;
  assign n16035 = pi5  & n16032;
  assign n16036 = ~n16032 & ~n16033;
  assign n16037 = ~pi5  & ~n16032;
  assign n16038 = ~n40364 & ~n40365;
  assign n16039 = n14110 & ~n14112;
  assign n16040 = ~n14113 & ~n16039;
  assign n16041 = ~n16038 & n16040;
  assign n16042 = n14101 & n39997;
  assign n16043 = ~n14109 & ~n16042;
  assign n16044 = n1218 & n14944;
  assign n16045 = pi72  & n40177;
  assign n16046 = pi74  & n14974;
  assign n16047 = pi73  & n14976;
  assign n16048 = ~n16046 & ~n16047;
  assign n16049 = ~n16045 & ~n16047;
  assign n16050 = ~n16046 & n16049;
  assign n16051 = ~n16045 & n16048;
  assign n16052 = ~n16044 & n40366;
  assign n16053 = pi5  & ~n16052;
  assign n16054 = pi5  & ~n16053;
  assign n16055 = pi5  & n16052;
  assign n16056 = ~n16052 & ~n16053;
  assign n16057 = ~pi5  & ~n16052;
  assign n16058 = ~n40367 & ~n40368;
  assign n16059 = n16043 & ~n16058;
  assign n16060 = n14092 & n39994;
  assign n16061 = ~n14100 & ~n16060;
  assign n16062 = n1238 & n14944;
  assign n16063 = pi71  & n40177;
  assign n16064 = pi73  & n14974;
  assign n16065 = pi72  & n14976;
  assign n16066 = ~n16064 & ~n16065;
  assign n16067 = ~n16063 & ~n16065;
  assign n16068 = ~n16064 & n16067;
  assign n16069 = ~n16063 & n16066;
  assign n16070 = ~n16062 & n40369;
  assign n16071 = pi5  & ~n16070;
  assign n16072 = pi5  & ~n16071;
  assign n16073 = pi5  & n16070;
  assign n16074 = ~n16070 & ~n16071;
  assign n16075 = ~pi5  & ~n16070;
  assign n16076 = ~n40370 & ~n40371;
  assign n16077 = n16061 & ~n16076;
  assign n16078 = ~n16061 & n16076;
  assign n16079 = ~n16077 & ~n16078;
  assign n16080 = n1124 & n14944;
  assign n16081 = pi70  & n40177;
  assign n16082 = pi72  & n14974;
  assign n16083 = pi71  & n14976;
  assign n16084 = ~n16082 & ~n16083;
  assign n16085 = ~n16081 & ~n16083;
  assign n16086 = ~n16082 & n16085;
  assign n16087 = ~n16081 & n16084;
  assign n16088 = ~n16080 & n40372;
  assign n16089 = pi5  & ~n16088;
  assign n16090 = pi5  & ~n16089;
  assign n16091 = pi5  & n16088;
  assign n16092 = ~n16088 & ~n16089;
  assign n16093 = ~pi5  & ~n16088;
  assign n16094 = ~n40373 & ~n40374;
  assign n16095 = n14083 & n39991;
  assign n16096 = ~n14091 & ~n16095;
  assign n16097 = ~n16094 & n16096;
  assign n16098 = n14079 & ~n14081;
  assign n16099 = ~n14082 & ~n16098;
  assign n16100 = n927 & n14944;
  assign n16101 = pi69  & n40177;
  assign n16102 = pi71  & n14974;
  assign n16103 = pi70  & n14976;
  assign n16104 = ~n16102 & ~n16103;
  assign n16105 = ~n16101 & ~n16103;
  assign n16106 = ~n16102 & n16105;
  assign n16107 = ~n16101 & n16104;
  assign n16108 = ~n16100 & n40375;
  assign n16109 = pi5  & ~n16108;
  assign n16110 = pi5  & ~n16109;
  assign n16111 = pi5  & n16108;
  assign n16112 = ~n16108 & ~n16109;
  assign n16113 = ~pi5  & ~n16108;
  assign n16114 = ~n40376 & ~n40377;
  assign n16115 = n16099 & ~n16114;
  assign n16116 = n14072 & n39988;
  assign n16117 = ~n14078 & ~n16116;
  assign n16118 = n972 & n14944;
  assign n16119 = pi68  & n40177;
  assign n16120 = pi70  & n14974;
  assign n16121 = pi69  & n14976;
  assign n16122 = ~n16120 & ~n16121;
  assign n16123 = ~n16119 & ~n16121;
  assign n16124 = ~n16120 & n16123;
  assign n16125 = ~n16119 & n16122;
  assign n16126 = ~n16118 & n40378;
  assign n16127 = pi5  & ~n16126;
  assign n16128 = pi5  & ~n16127;
  assign n16129 = pi5  & n16126;
  assign n16130 = ~n16126 & ~n16127;
  assign n16131 = ~pi5  & ~n16126;
  assign n16132 = ~n40379 & ~n40380;
  assign n16133 = n16117 & ~n16132;
  assign n16134 = n990 & n14944;
  assign n16135 = pi67  & n40177;
  assign n16136 = pi69  & n14974;
  assign n16137 = pi68  & n14976;
  assign n16138 = ~n16136 & ~n16137;
  assign n16139 = ~n16135 & ~n16137;
  assign n16140 = ~n16136 & n16139;
  assign n16141 = ~n16135 & n16138;
  assign n16142 = ~n16134 & n40381;
  assign n16143 = pi5  & ~n16142;
  assign n16144 = pi5  & ~n16143;
  assign n16145 = pi5  & n16142;
  assign n16146 = ~n16142 & ~n16143;
  assign n16147 = ~pi5  & ~n16142;
  assign n16148 = ~n40382 & ~n40383;
  assign n16149 = pi8  & ~n39980;
  assign n16150 = n39983 & ~n16149;
  assign n16151 = ~n39983 & n16149;
  assign n16152 = ~n39980 & n14054;
  assign n16153 = ~n39984 & ~n16152;
  assign n16154 = ~n16150 & ~n16151;
  assign n16155 = ~n16148 & n40384;
  assign n16156 = n871 & n14944;
  assign n16157 = pi66  & n40177;
  assign n16158 = pi68  & n14974;
  assign n16159 = pi67  & n14976;
  assign n16160 = ~n16158 & ~n16159;
  assign n16161 = ~n16157 & ~n16159;
  assign n16162 = ~n16158 & n16161;
  assign n16163 = ~n16157 & n16160;
  assign n16164 = ~n16156 & n40385;
  assign n16165 = pi5  & ~n16164;
  assign n16166 = pi5  & ~n16165;
  assign n16167 = pi5  & n16164;
  assign n16168 = ~n16164 & ~n16165;
  assign n16169 = ~pi5  & ~n16164;
  assign n16170 = ~n40386 & ~n40387;
  assign n16171 = pi8  & n14028;
  assign n16172 = ~n14027 & n16171;
  assign n16173 = n14027 & ~n16171;
  assign n16174 = ~n14029 & n14033;
  assign n16175 = ~n39980 & ~n16174;
  assign n16176 = ~n16172 & ~n16173;
  assign n16177 = ~n16170 & n40388;
  assign n16178 = n37515 & n14944;
  assign n16179 = pi65  & n14974;
  assign n16180 = pi64  & n14976;
  assign n16181 = ~n16179 & ~n16180;
  assign n16182 = ~n16178 & n16181;
  assign n16183 = pi64  & n40174;
  assign n16184 = pi5  & ~n16183;
  assign n16185 = pi5  & ~n16182;
  assign n16186 = pi5  & ~n16185;
  assign n16187 = ~n16182 & ~n16185;
  assign n16188 = ~n16186 & ~n16187;
  assign n16189 = n16184 & ~n16188;
  assign n16190 = n16182 & n16184;
  assign n16191 = pi64  & n40177;
  assign n16192 = pi65  & n14976;
  assign n16193 = pi66  & n14974;
  assign n16194 = ~n37521 & n14944;
  assign n16195 = ~n16193 & ~n16194;
  assign n16196 = ~n16192 & ~n16193;
  assign n16197 = ~n16194 & n16196;
  assign n16198 = ~n16192 & n16195;
  assign n16199 = ~n16191 & ~n16192;
  assign n16200 = ~n16193 & n16199;
  assign n16201 = ~n16191 & n16196;
  assign n16202 = ~n16194 & n40391;
  assign n16203 = ~n14944 & n40391;
  assign n16204 = n37521 & n40391;
  assign n16205 = ~n16203 & ~n16204;
  assign n16206 = ~n16191 & n40390;
  assign n16207 = pi5  & n40392;
  assign n16208 = ~pi5  & ~n40392;
  assign n16209 = ~n16207 & ~n16208;
  assign n16210 = n40389 & ~n16209;
  assign n16211 = n40389 & n40392;
  assign n16212 = n14028 & n40393;
  assign n16213 = n847 & n14944;
  assign n16214 = pi65  & n40177;
  assign n16215 = pi67  & n14974;
  assign n16216 = pi66  & n14976;
  assign n16217 = ~n16215 & ~n16216;
  assign n16218 = ~n16214 & ~n16216;
  assign n16219 = ~n16215 & n16218;
  assign n16220 = ~n16214 & n16217;
  assign n16221 = ~n16213 & n40394;
  assign n16222 = pi5  & ~n16221;
  assign n16223 = pi5  & ~n16222;
  assign n16224 = pi5  & n16221;
  assign n16225 = ~n16221 & ~n16222;
  assign n16226 = ~pi5  & ~n16221;
  assign n16227 = ~n40395 & ~n40396;
  assign n16228 = ~n14028 & ~n40393;
  assign n16229 = n40393 & ~n16212;
  assign n16230 = ~n14028 & n40393;
  assign n16231 = n14028 & ~n16212;
  assign n16232 = n14028 & ~n40393;
  assign n16233 = ~n40397 & ~n40398;
  assign n16234 = ~n16212 & ~n16228;
  assign n16235 = ~n16227 & ~n40399;
  assign n16236 = ~n16212 & ~n16235;
  assign n16237 = n16170 & ~n40388;
  assign n16238 = n40388 & ~n16177;
  assign n16239 = n16170 & n40388;
  assign n16240 = ~n16170 & ~n16177;
  assign n16241 = ~n16170 & ~n40388;
  assign n16242 = ~n40400 & ~n40401;
  assign n16243 = ~n16177 & ~n16237;
  assign n16244 = ~n16236 & ~n40402;
  assign n16245 = ~n16177 & ~n16244;
  assign n16246 = n16148 & ~n40384;
  assign n16247 = n40384 & ~n16155;
  assign n16248 = n16148 & n40384;
  assign n16249 = ~n16148 & ~n16155;
  assign n16250 = ~n16148 & ~n40384;
  assign n16251 = ~n40403 & ~n40404;
  assign n16252 = ~n16155 & ~n16246;
  assign n16253 = ~n16245 & ~n40405;
  assign n16254 = ~n16155 & ~n16253;
  assign n16255 = ~n16117 & n16132;
  assign n16256 = n16117 & ~n16133;
  assign n16257 = n16117 & n16132;
  assign n16258 = ~n16132 & ~n16133;
  assign n16259 = ~n16117 & ~n16132;
  assign n16260 = ~n40406 & ~n40407;
  assign n16261 = ~n16133 & ~n16255;
  assign n16262 = ~n16254 & ~n40408;
  assign n16263 = ~n16133 & ~n16262;
  assign n16264 = ~n16099 & n16114;
  assign n16265 = n16099 & ~n16115;
  assign n16266 = n16099 & n16114;
  assign n16267 = ~n16114 & ~n16115;
  assign n16268 = ~n16099 & ~n16114;
  assign n16269 = ~n40409 & ~n40410;
  assign n16270 = ~n16115 & ~n16264;
  assign n16271 = ~n16263 & ~n40411;
  assign n16272 = ~n16115 & ~n16271;
  assign n16273 = n16094 & ~n16096;
  assign n16274 = ~n16094 & ~n16097;
  assign n16275 = ~n16094 & ~n16096;
  assign n16276 = n16096 & ~n16097;
  assign n16277 = n16094 & n16096;
  assign n16278 = ~n40412 & ~n40413;
  assign n16279 = ~n16097 & ~n16273;
  assign n16280 = ~n16272 & ~n40414;
  assign n16281 = ~n16097 & ~n16280;
  assign n16282 = n16079 & ~n16281;
  assign n16283 = ~n16077 & ~n16282;
  assign n16284 = ~n16043 & n16058;
  assign n16285 = ~n16059 & ~n16284;
  assign n16286 = ~n16283 & ~n16284;
  assign n16287 = ~n16059 & n16286;
  assign n16288 = ~n16283 & n16285;
  assign n16289 = ~n16059 & ~n40415;
  assign n16290 = n16038 & ~n16040;
  assign n16291 = ~n16041 & ~n16290;
  assign n16292 = ~n16289 & n16291;
  assign n16293 = ~n16041 & ~n16292;
  assign n16294 = n16018 & ~n16022;
  assign n16295 = ~n16018 & ~n16023;
  assign n16296 = ~n16018 & ~n16022;
  assign n16297 = n16022 & ~n16023;
  assign n16298 = n16018 & n16022;
  assign n16299 = ~n40416 & ~n40417;
  assign n16300 = ~n16023 & ~n16294;
  assign n16301 = ~n16293 & ~n40418;
  assign n16302 = ~n16023 & ~n16301;
  assign n16303 = n16000 & ~n16002;
  assign n16304 = ~n16003 & ~n16303;
  assign n16305 = ~n16302 & n16304;
  assign n16306 = ~n16003 & ~n16305;
  assign n16307 = n15982 & ~n15984;
  assign n16308 = ~n15985 & ~n16307;
  assign n16309 = ~n16306 & n16308;
  assign n16310 = ~n15985 & ~n16309;
  assign n16311 = n15964 & ~n15966;
  assign n16312 = ~n15967 & ~n16311;
  assign n16313 = ~n16310 & n16312;
  assign n16314 = ~n15967 & ~n16313;
  assign n16315 = ~n15933 & n15948;
  assign n16316 = n15933 & ~n15949;
  assign n16317 = n15933 & n15948;
  assign n16318 = ~n15948 & ~n15949;
  assign n16319 = ~n15933 & ~n15948;
  assign n16320 = ~n40419 & ~n40420;
  assign n16321 = ~n15949 & ~n16315;
  assign n16322 = ~n16314 & ~n40421;
  assign n16323 = ~n15949 & ~n16322;
  assign n16324 = n15928 & ~n15930;
  assign n16325 = ~n15928 & ~n15931;
  assign n16326 = ~n15928 & ~n15930;
  assign n16327 = n15930 & ~n15931;
  assign n16328 = n15928 & n15930;
  assign n16329 = ~n40422 & ~n40423;
  assign n16330 = ~n15931 & ~n16324;
  assign n16331 = ~n16323 & ~n40424;
  assign n16332 = ~n15931 & ~n16331;
  assign n16333 = ~n15897 & n15912;
  assign n16334 = n15897 & ~n15913;
  assign n16335 = n15897 & n15912;
  assign n16336 = ~n15912 & ~n15913;
  assign n16337 = ~n15897 & ~n15912;
  assign n16338 = ~n40425 & ~n40426;
  assign n16339 = ~n15913 & ~n16333;
  assign n16340 = ~n16332 & ~n40427;
  assign n16341 = ~n15913 & ~n16340;
  assign n16342 = ~n15879 & n15894;
  assign n16343 = n15879 & ~n15895;
  assign n16344 = n15879 & n15894;
  assign n16345 = ~n15894 & ~n15895;
  assign n16346 = ~n15879 & ~n15894;
  assign n16347 = ~n40428 & ~n40429;
  assign n16348 = ~n15895 & ~n16342;
  assign n16349 = ~n16341 & ~n40430;
  assign n16350 = ~n15895 & ~n16349;
  assign n16351 = n15869 & n40337;
  assign n16352 = ~n40337 & ~n15877;
  assign n16353 = ~n15869 & ~n15877;
  assign n16354 = ~n16352 & ~n16353;
  assign n16355 = ~n15877 & ~n16351;
  assign n16356 = ~n16350 & ~n40431;
  assign n16357 = ~n15877 & ~n16356;
  assign n16358 = n15851 & ~n15853;
  assign n16359 = ~n15851 & ~n15854;
  assign n16360 = ~n15851 & ~n15853;
  assign n16361 = n15853 & ~n15854;
  assign n16362 = n15851 & n15853;
  assign n16363 = ~n40432 & ~n40433;
  assign n16364 = ~n15854 & ~n16358;
  assign n16365 = ~n16357 & ~n40434;
  assign n16366 = ~n15854 & ~n16365;
  assign n16367 = n15828 & n40328;
  assign n16368 = n15828 & ~n40328;
  assign n16369 = ~n15828 & n40328;
  assign n16370 = ~n16368 & ~n16369;
  assign n16371 = ~n15836 & ~n16367;
  assign n16372 = ~n16366 & ~n40435;
  assign n16373 = ~n15836 & ~n16372;
  assign n16374 = ~n15797 & n15812;
  assign n16375 = n15797 & ~n15813;
  assign n16376 = n15797 & n15812;
  assign n16377 = ~n15812 & ~n15813;
  assign n16378 = ~n15797 & ~n15812;
  assign n16379 = ~n40436 & ~n40437;
  assign n16380 = ~n15813 & ~n16374;
  assign n16381 = ~n16373 & ~n40438;
  assign n16382 = ~n15813 & ~n16381;
  assign n16383 = ~n15779 & n15794;
  assign n16384 = n15779 & ~n15795;
  assign n16385 = n15779 & n15794;
  assign n16386 = ~n15794 & ~n15795;
  assign n16387 = ~n15779 & ~n15794;
  assign n16388 = ~n40439 & ~n40440;
  assign n16389 = ~n15795 & ~n16383;
  assign n16390 = ~n16382 & ~n40441;
  assign n16391 = ~n15795 & ~n16390;
  assign n16392 = ~n15761 & n15776;
  assign n16393 = n15761 & ~n15777;
  assign n16394 = n15761 & n15776;
  assign n16395 = ~n15776 & ~n15777;
  assign n16396 = ~n15761 & ~n15776;
  assign n16397 = ~n40442 & ~n40443;
  assign n16398 = ~n15777 & ~n16392;
  assign n16399 = ~n16391 & ~n40444;
  assign n16400 = ~n15777 & ~n16399;
  assign n16401 = n15756 & ~n15758;
  assign n16402 = ~n15756 & ~n15759;
  assign n16403 = ~n15756 & ~n15758;
  assign n16404 = n15758 & ~n15759;
  assign n16405 = n15756 & n15758;
  assign n16406 = ~n40445 & ~n40446;
  assign n16407 = ~n15759 & ~n16401;
  assign n16408 = ~n16400 & ~n40447;
  assign n16409 = ~n15759 & ~n16408;
  assign n16410 = ~n15725 & n15740;
  assign n16411 = n15725 & ~n15741;
  assign n16412 = n15725 & n15740;
  assign n16413 = ~n15740 & ~n15741;
  assign n16414 = ~n15725 & ~n15740;
  assign n16415 = ~n40448 & ~n40449;
  assign n16416 = ~n15741 & ~n16410;
  assign n16417 = ~n16409 & ~n40450;
  assign n16418 = ~n15741 & ~n16417;
  assign n16419 = ~n15707 & n15722;
  assign n16420 = n15707 & ~n15723;
  assign n16421 = n15707 & n15722;
  assign n16422 = ~n15722 & ~n15723;
  assign n16423 = ~n15707 & ~n15722;
  assign n16424 = ~n40451 & ~n40452;
  assign n16425 = ~n15723 & ~n16419;
  assign n16426 = ~n16418 & ~n40453;
  assign n16427 = ~n15723 & ~n16426;
  assign n16428 = ~n15689 & n15704;
  assign n16429 = ~n15705 & ~n16428;
  assign n16430 = ~n16427 & ~n16428;
  assign n16431 = ~n15705 & n16430;
  assign n16432 = ~n16427 & n16429;
  assign n16433 = ~n15705 & ~n40454;
  assign n16434 = ~n15671 & n15686;
  assign n16435 = n15671 & ~n15687;
  assign n16436 = n15671 & n15686;
  assign n16437 = ~n15686 & ~n15687;
  assign n16438 = ~n15671 & ~n15686;
  assign n16439 = ~n40455 & ~n40456;
  assign n16440 = ~n15687 & ~n16434;
  assign n16441 = ~n16433 & ~n40457;
  assign n16442 = ~n15687 & ~n16441;
  assign n16443 = ~n15653 & n15668;
  assign n16444 = ~n15669 & ~n16443;
  assign n16445 = ~n16442 & ~n16443;
  assign n16446 = ~n15669 & n16445;
  assign n16447 = ~n16442 & n16444;
  assign n16448 = ~n15669 & ~n40458;
  assign n16449 = ~n15635 & n15650;
  assign n16450 = ~n15651 & ~n16449;
  assign n16451 = ~n16448 & ~n16449;
  assign n16452 = ~n15651 & n16451;
  assign n16453 = ~n16448 & n16450;
  assign n16454 = ~n15651 & ~n40459;
  assign n16455 = n15630 & ~n15632;
  assign n16456 = ~n15633 & ~n16455;
  assign n16457 = ~n16454 & n16456;
  assign n16458 = ~n15633 & ~n16457;
  assign n16459 = ~n15599 & n15614;
  assign n16460 = n15599 & ~n15615;
  assign n16461 = n15599 & n15614;
  assign n16462 = ~n15614 & ~n15615;
  assign n16463 = ~n15599 & ~n15614;
  assign n16464 = ~n40460 & ~n40461;
  assign n16465 = ~n15615 & ~n16459;
  assign n16466 = ~n16458 & ~n40462;
  assign n16467 = ~n15615 & ~n16466;
  assign n16468 = n15594 & ~n15596;
  assign n16469 = ~n15597 & ~n16468;
  assign n16470 = ~n16467 & n16469;
  assign n16471 = ~n15597 & ~n16470;
  assign n16472 = n15573 & n40283;
  assign n16473 = ~n15579 & ~n16472;
  assign n16474 = ~n16471 & n16473;
  assign n16475 = ~n15579 & ~n16474;
  assign n16476 = ~n15542 & n15557;
  assign n16477 = n15542 & ~n15558;
  assign n16478 = n15542 & n15557;
  assign n16479 = ~n15557 & ~n15558;
  assign n16480 = ~n15542 & ~n15557;
  assign n16481 = ~n40463 & ~n40464;
  assign n16482 = ~n15558 & ~n16476;
  assign n16483 = ~n16475 & ~n40465;
  assign n16484 = ~n15558 & ~n16483;
  assign n16485 = n15534 & n40276;
  assign n16486 = ~n15540 & ~n16485;
  assign n16487 = ~n16484 & n16486;
  assign n16488 = ~n15540 & ~n16487;
  assign n16489 = n15516 & ~n15518;
  assign n16490 = ~n15516 & ~n15519;
  assign n16491 = ~n15516 & ~n15518;
  assign n16492 = n15518 & ~n15519;
  assign n16493 = n15516 & n15518;
  assign n16494 = ~n40466 & ~n40467;
  assign n16495 = ~n15519 & ~n16489;
  assign n16496 = ~n16488 & ~n40468;
  assign n16497 = ~n15519 & ~n16496;
  assign n16498 = n15495 & n40269;
  assign n16499 = ~n15501 & ~n16498;
  assign n16500 = ~n16497 & n16499;
  assign n16501 = ~n15501 & ~n16500;
  assign n16502 = n15477 & ~n15479;
  assign n16503 = ~n15477 & ~n15480;
  assign n16504 = ~n15477 & ~n15479;
  assign n16505 = n15479 & ~n15480;
  assign n16506 = n15477 & n15479;
  assign n16507 = ~n40469 & ~n40470;
  assign n16508 = ~n15480 & ~n16502;
  assign n16509 = ~n16501 & ~n40471;
  assign n16510 = ~n15480 & ~n16509;
  assign n16511 = ~n15446 & n15461;
  assign n16512 = n15446 & ~n15462;
  assign n16513 = n15446 & n15461;
  assign n16514 = ~n15461 & ~n15462;
  assign n16515 = ~n15446 & ~n15461;
  assign n16516 = ~n40472 & ~n40473;
  assign n16517 = ~n15462 & ~n16511;
  assign n16518 = ~n16510 & ~n40474;
  assign n16519 = ~n15462 & ~n16518;
  assign n16520 = n15438 & n40259;
  assign n16521 = ~n40259 & ~n15444;
  assign n16522 = n15438 & ~n40259;
  assign n16523 = ~n15438 & ~n15444;
  assign n16524 = ~n15438 & n40259;
  assign n16525 = ~n40475 & ~n40476;
  assign n16526 = ~n15444 & ~n16520;
  assign n16527 = ~n16519 & ~n40477;
  assign n16528 = ~n15444 & ~n16527;
  assign n16529 = n15417 & n40255;
  assign n16530 = ~n15423 & ~n16529;
  assign n16531 = ~n16528 & n16530;
  assign n16532 = ~n15423 & ~n16531;
  assign n16533 = n15396 & n40251;
  assign n16534 = ~n15402 & ~n16533;
  assign n16535 = ~n16532 & n16534;
  assign n16536 = ~n15402 & ~n16535;
  assign n16537 = ~n15365 & n15380;
  assign n16538 = n15365 & ~n15381;
  assign n16539 = n15365 & n15380;
  assign n16540 = ~n15380 & ~n15381;
  assign n16541 = ~n15365 & ~n15380;
  assign n16542 = ~n40478 & ~n40479;
  assign n16543 = ~n15381 & ~n16537;
  assign n16544 = ~n16536 & ~n40480;
  assign n16545 = ~n15381 & ~n16544;
  assign n16546 = n15357 & n40244;
  assign n16547 = ~n40244 & ~n15363;
  assign n16548 = n15357 & ~n40244;
  assign n16549 = ~n15357 & ~n15363;
  assign n16550 = ~n15357 & n40244;
  assign n16551 = ~n40481 & ~n40482;
  assign n16552 = ~n15363 & ~n16546;
  assign n16553 = ~n16545 & ~n40483;
  assign n16554 = ~n15363 & ~n16553;
  assign n16555 = n15336 & n40240;
  assign n16556 = ~n15342 & ~n16555;
  assign n16557 = ~n16554 & n16556;
  assign n16558 = ~n15342 & ~n16557;
  assign n16559 = ~n15305 & n15320;
  assign n16560 = n15305 & ~n15321;
  assign n16561 = n15305 & n15320;
  assign n16562 = ~n15320 & ~n15321;
  assign n16563 = ~n15305 & ~n15320;
  assign n16564 = ~n40484 & ~n40485;
  assign n16565 = ~n15321 & ~n16559;
  assign n16566 = ~n16558 & ~n40486;
  assign n16567 = ~n15321 & ~n16566;
  assign n16568 = ~n15287 & n15302;
  assign n16569 = ~n15303 & ~n16568;
  assign n16570 = ~n16567 & ~n16568;
  assign n16571 = ~n15303 & n16570;
  assign n16572 = ~n16567 & n16569;
  assign n16573 = ~n15303 & ~n40487;
  assign n16574 = ~n15269 & n15284;
  assign n16575 = ~n15285 & ~n16574;
  assign n16576 = ~n16573 & n16575;
  assign n16577 = ~n15285 & ~n16576;
  assign n16578 = ~n15251 & n15266;
  assign n16579 = n15251 & ~n15267;
  assign n16580 = n15251 & n15266;
  assign n16581 = ~n15266 & ~n15267;
  assign n16582 = ~n15251 & ~n15266;
  assign n16583 = ~n40488 & ~n40489;
  assign n16584 = ~n15267 & ~n16578;
  assign n16585 = ~n16577 & ~n40490;
  assign n16586 = ~n15267 & ~n16585;
  assign n16587 = n15241 & n40224;
  assign n16588 = ~n15249 & ~n16587;
  assign n16589 = ~n16586 & n16588;
  assign n16590 = ~n15249 & ~n16589;
  assign n16591 = n15221 & ~n15225;
  assign n16592 = ~n15221 & ~n15226;
  assign n16593 = ~n15221 & ~n15225;
  assign n16594 = n15225 & ~n15226;
  assign n16595 = n15221 & n15225;
  assign n16596 = ~n40491 & ~n40492;
  assign n16597 = ~n15226 & ~n16591;
  assign n16598 = ~n16590 & ~n40493;
  assign n16599 = ~n15226 & ~n16598;
  assign n16600 = n15203 & ~n15205;
  assign n16601 = ~n15206 & ~n16600;
  assign n16602 = ~n16599 & n16601;
  assign n16603 = ~n15206 & ~n16602;
  assign n16604 = n15178 & n40210;
  assign n16605 = n15178 & ~n40210;
  assign n16606 = ~n15178 & n40210;
  assign n16607 = ~n16605 & ~n16606;
  assign n16608 = ~n15185 & ~n16604;
  assign n16609 = ~n16603 & ~n40494;
  assign n16610 = n16599 & ~n16601;
  assign n16611 = ~n16602 & ~n16610;
  assign n16612 = n15004 & n15049;
  assign n16613 = pi120  & n40183;
  assign n16614 = pi122  & n15023;
  assign n16615 = pi121  & n15030;
  assign n16616 = ~n16614 & ~n16615;
  assign n16617 = ~n16613 & ~n16615;
  assign n16618 = ~n16614 & n16617;
  assign n16619 = ~n16613 & n16616;
  assign n16620 = ~n16612 & n40495;
  assign n16621 = pi2  & ~n16620;
  assign n16622 = pi2  & ~n16621;
  assign n16623 = pi2  & n16620;
  assign n16624 = ~n16620 & ~n16621;
  assign n16625 = ~pi2  & ~n16620;
  assign n16626 = ~n40496 & ~n40497;
  assign n16627 = n16611 & ~n16626;
  assign n16628 = n15004 & n15091;
  assign n16629 = pi119  & n40183;
  assign n16630 = pi121  & n15023;
  assign n16631 = pi120  & n15030;
  assign n16632 = ~n16630 & ~n16631;
  assign n16633 = ~n16629 & ~n16631;
  assign n16634 = ~n16630 & n16633;
  assign n16635 = ~n16629 & n16632;
  assign n16636 = ~n16628 & n40498;
  assign n16637 = pi2  & ~n16636;
  assign n16638 = pi2  & ~n16637;
  assign n16639 = pi2  & n16636;
  assign n16640 = ~n16636 & ~n16637;
  assign n16641 = ~pi2  & ~n16636;
  assign n16642 = ~n40499 & ~n40500;
  assign n16643 = n16590 & n40493;
  assign n16644 = ~n16590 & ~n16598;
  assign n16645 = ~n16590 & n40493;
  assign n16646 = ~n40493 & ~n16598;
  assign n16647 = n16590 & ~n40493;
  assign n16648 = ~n40501 & ~n40502;
  assign n16649 = ~n16598 & ~n16643;
  assign n16650 = ~n16642 & ~n40503;
  assign n16651 = n16586 & ~n16588;
  assign n16652 = ~n16589 & ~n16651;
  assign n16653 = n14913 & n15004;
  assign n16654 = pi118  & n40183;
  assign n16655 = pi120  & n15023;
  assign n16656 = pi119  & n15030;
  assign n16657 = ~n16655 & ~n16656;
  assign n16658 = ~n16654 & ~n16656;
  assign n16659 = ~n16655 & n16658;
  assign n16660 = ~n16654 & n16657;
  assign n16661 = ~n16653 & n40504;
  assign n16662 = pi2  & ~n16661;
  assign n16663 = pi2  & ~n16662;
  assign n16664 = pi2  & n16661;
  assign n16665 = ~n16661 & ~n16662;
  assign n16666 = ~pi2  & ~n16661;
  assign n16667 = ~n40505 & ~n40506;
  assign n16668 = n16652 & ~n16667;
  assign n16669 = n13027 & n15004;
  assign n16670 = pi117  & n40183;
  assign n16671 = pi119  & n15023;
  assign n16672 = pi118  & n15030;
  assign n16673 = ~n16671 & ~n16672;
  assign n16674 = ~n16670 & ~n16672;
  assign n16675 = ~n16671 & n16674;
  assign n16676 = ~n16670 & n16673;
  assign n16677 = ~n16669 & n40507;
  assign n16678 = pi2  & ~n16677;
  assign n16679 = pi2  & ~n16678;
  assign n16680 = pi2  & n16677;
  assign n16681 = ~n16677 & ~n16678;
  assign n16682 = ~pi2  & ~n16677;
  assign n16683 = ~n40508 & ~n40509;
  assign n16684 = n16577 & n40490;
  assign n16685 = ~n16577 & n40490;
  assign n16686 = n16577 & ~n40490;
  assign n16687 = ~n16685 & ~n16686;
  assign n16688 = ~n16585 & ~n16684;
  assign n16689 = ~n16683 & ~n40510;
  assign n16690 = n13057 & n15004;
  assign n16691 = pi116  & n40183;
  assign n16692 = pi118  & n15023;
  assign n16693 = pi117  & n15030;
  assign n16694 = ~n16692 & ~n16693;
  assign n16695 = ~n16691 & ~n16693;
  assign n16696 = ~n16692 & n16695;
  assign n16697 = ~n16691 & n16694;
  assign n16698 = ~n16690 & n40511;
  assign n16699 = pi2  & ~n16698;
  assign n16700 = pi2  & ~n16699;
  assign n16701 = pi2  & n16698;
  assign n16702 = ~n16698 & ~n16699;
  assign n16703 = ~pi2  & ~n16698;
  assign n16704 = ~n40512 & ~n40513;
  assign n16705 = n16573 & ~n16575;
  assign n16706 = ~n16576 & ~n16705;
  assign n16707 = ~n16704 & n16706;
  assign n16708 = n13079 & n15004;
  assign n16709 = pi115  & n40183;
  assign n16710 = pi117  & n15023;
  assign n16711 = pi116  & n15030;
  assign n16712 = ~n16710 & ~n16711;
  assign n16713 = ~n16709 & ~n16711;
  assign n16714 = ~n16710 & n16713;
  assign n16715 = ~n16709 & n16712;
  assign n16716 = ~n16708 & n40514;
  assign n16717 = pi2  & ~n16716;
  assign n16718 = pi2  & ~n16717;
  assign n16719 = pi2  & n16716;
  assign n16720 = ~n16716 & ~n16717;
  assign n16721 = ~pi2  & ~n16716;
  assign n16722 = ~n40515 & ~n40516;
  assign n16723 = n16567 & ~n16569;
  assign n16724 = ~n16567 & ~n40487;
  assign n16725 = ~n16568 & n16573;
  assign n16726 = ~n16724 & ~n16725;
  assign n16727 = ~n40487 & ~n16723;
  assign n16728 = ~n16722 & ~n40517;
  assign n16729 = n12530 & n15004;
  assign n16730 = pi114  & n40183;
  assign n16731 = pi116  & n15023;
  assign n16732 = pi115  & n15030;
  assign n16733 = ~n16731 & ~n16732;
  assign n16734 = ~n16730 & ~n16732;
  assign n16735 = ~n16731 & n16734;
  assign n16736 = ~n16730 & n16733;
  assign n16737 = ~n16729 & n40518;
  assign n16738 = pi2  & ~n16737;
  assign n16739 = pi2  & ~n16738;
  assign n16740 = pi2  & n16737;
  assign n16741 = ~n16737 & ~n16738;
  assign n16742 = ~pi2  & ~n16737;
  assign n16743 = ~n40519 & ~n40520;
  assign n16744 = n16558 & n40486;
  assign n16745 = ~n16558 & n40486;
  assign n16746 = n16558 & ~n40486;
  assign n16747 = ~n16745 & ~n16746;
  assign n16748 = ~n16566 & ~n16744;
  assign n16749 = ~n16743 & ~n40521;
  assign n16750 = n523 & n15004;
  assign n16751 = pi113  & n40183;
  assign n16752 = pi115  & n15023;
  assign n16753 = pi114  & n15030;
  assign n16754 = ~n16752 & ~n16753;
  assign n16755 = ~n16751 & ~n16753;
  assign n16756 = ~n16752 & n16755;
  assign n16757 = ~n16751 & n16754;
  assign n16758 = ~n16750 & n40522;
  assign n16759 = pi2  & ~n16758;
  assign n16760 = pi2  & ~n16759;
  assign n16761 = pi2  & n16758;
  assign n16762 = ~n16758 & ~n16759;
  assign n16763 = ~pi2  & ~n16758;
  assign n16764 = ~n40523 & ~n40524;
  assign n16765 = n16554 & ~n16556;
  assign n16766 = ~n16557 & ~n16765;
  assign n16767 = ~n16764 & n16766;
  assign n16768 = n16545 & n40483;
  assign n16769 = ~n16553 & ~n16768;
  assign n16770 = n11258 & n15004;
  assign n16771 = pi112  & n40183;
  assign n16772 = pi114  & n15023;
  assign n16773 = pi113  & n15030;
  assign n16774 = ~n16772 & ~n16773;
  assign n16775 = ~n16771 & ~n16773;
  assign n16776 = ~n16772 & n16775;
  assign n16777 = ~n16771 & n16774;
  assign n16778 = ~n16770 & n40525;
  assign n16779 = pi2  & ~n16778;
  assign n16780 = pi2  & ~n16779;
  assign n16781 = pi2  & n16778;
  assign n16782 = ~n16778 & ~n16779;
  assign n16783 = ~pi2  & ~n16778;
  assign n16784 = ~n40526 & ~n40527;
  assign n16785 = n16769 & ~n16784;
  assign n16786 = n16536 & n40480;
  assign n16787 = ~n16544 & ~n16786;
  assign n16788 = n11276 & n15004;
  assign n16789 = pi111  & n40183;
  assign n16790 = pi113  & n15023;
  assign n16791 = pi112  & n15030;
  assign n16792 = ~n16790 & ~n16791;
  assign n16793 = ~n16789 & ~n16791;
  assign n16794 = ~n16790 & n16793;
  assign n16795 = ~n16789 & n16792;
  assign n16796 = ~n16788 & n40528;
  assign n16797 = pi2  & ~n16796;
  assign n16798 = pi2  & ~n16797;
  assign n16799 = pi2  & n16796;
  assign n16800 = ~n16796 & ~n16797;
  assign n16801 = ~pi2  & ~n16796;
  assign n16802 = ~n40529 & ~n40530;
  assign n16803 = n16787 & ~n16802;
  assign n16804 = n10844 & n15004;
  assign n16805 = pi110  & n40183;
  assign n16806 = pi112  & n15023;
  assign n16807 = pi111  & n15030;
  assign n16808 = ~n16806 & ~n16807;
  assign n16809 = ~n16805 & ~n16807;
  assign n16810 = ~n16806 & n16809;
  assign n16811 = ~n16805 & n16808;
  assign n16812 = ~n16804 & n40531;
  assign n16813 = pi2  & ~n16812;
  assign n16814 = pi2  & ~n16813;
  assign n16815 = pi2  & n16812;
  assign n16816 = ~n16812 & ~n16813;
  assign n16817 = ~pi2  & ~n16812;
  assign n16818 = ~n40532 & ~n40533;
  assign n16819 = n16532 & ~n16534;
  assign n16820 = ~n16535 & ~n16819;
  assign n16821 = ~n16818 & n16820;
  assign n16822 = n16528 & ~n16530;
  assign n16823 = ~n16531 & ~n16822;
  assign n16824 = n565 & n15004;
  assign n16825 = pi109  & n40183;
  assign n16826 = pi111  & n15023;
  assign n16827 = pi110  & n15030;
  assign n16828 = ~n16826 & ~n16827;
  assign n16829 = ~n16825 & ~n16827;
  assign n16830 = ~n16826 & n16829;
  assign n16831 = ~n16825 & n16828;
  assign n16832 = ~n16824 & n40534;
  assign n16833 = pi2  & ~n16832;
  assign n16834 = pi2  & ~n16833;
  assign n16835 = pi2  & n16832;
  assign n16836 = ~n16832 & ~n16833;
  assign n16837 = ~pi2  & ~n16832;
  assign n16838 = ~n40535 & ~n40536;
  assign n16839 = n16823 & ~n16838;
  assign n16840 = n16519 & n40477;
  assign n16841 = ~n16527 & ~n16840;
  assign n16842 = n9678 & n15004;
  assign n16843 = pi108  & n40183;
  assign n16844 = pi110  & n15023;
  assign n16845 = pi109  & n15030;
  assign n16846 = ~n16844 & ~n16845;
  assign n16847 = ~n16843 & ~n16845;
  assign n16848 = ~n16844 & n16847;
  assign n16849 = ~n16843 & n16846;
  assign n16850 = ~n16842 & n40537;
  assign n16851 = pi2  & ~n16850;
  assign n16852 = pi2  & ~n16851;
  assign n16853 = pi2  & n16850;
  assign n16854 = ~n16850 & ~n16851;
  assign n16855 = ~pi2  & ~n16850;
  assign n16856 = ~n40538 & ~n40539;
  assign n16857 = n16841 & ~n16856;
  assign n16858 = n16510 & n40474;
  assign n16859 = ~n16518 & ~n16858;
  assign n16860 = n9701 & n15004;
  assign n16861 = pi107  & n40183;
  assign n16862 = pi109  & n15023;
  assign n16863 = pi108  & n15030;
  assign n16864 = ~n16862 & ~n16863;
  assign n16865 = ~n16861 & ~n16863;
  assign n16866 = ~n16862 & n16865;
  assign n16867 = ~n16861 & n16864;
  assign n16868 = ~n16860 & n40540;
  assign n16869 = pi2  & ~n16868;
  assign n16870 = pi2  & ~n16869;
  assign n16871 = pi2  & n16868;
  assign n16872 = ~n16868 & ~n16869;
  assign n16873 = ~pi2  & ~n16868;
  assign n16874 = ~n40541 & ~n40542;
  assign n16875 = n16859 & ~n16874;
  assign n16876 = n9277 & n15004;
  assign n16877 = pi106  & n40183;
  assign n16878 = pi108  & n15023;
  assign n16879 = pi107  & n15030;
  assign n16880 = ~n16878 & ~n16879;
  assign n16881 = ~n16877 & ~n16879;
  assign n16882 = ~n16878 & n16881;
  assign n16883 = ~n16877 & n16880;
  assign n16884 = ~n16876 & n40543;
  assign n16885 = pi2  & ~n16884;
  assign n16886 = pi2  & ~n16885;
  assign n16887 = pi2  & n16884;
  assign n16888 = ~n16884 & ~n16885;
  assign n16889 = ~pi2  & ~n16884;
  assign n16890 = ~n40544 & ~n40545;
  assign n16891 = n16501 & n40471;
  assign n16892 = ~n16501 & ~n16509;
  assign n16893 = ~n16501 & n40471;
  assign n16894 = ~n40471 & ~n16509;
  assign n16895 = n16501 & ~n40471;
  assign n16896 = ~n40546 & ~n40547;
  assign n16897 = ~n16509 & ~n16891;
  assign n16898 = ~n16890 & ~n40548;
  assign n16899 = n16497 & ~n16499;
  assign n16900 = ~n16500 & ~n16899;
  assign n16901 = n8177 & n15004;
  assign n16902 = pi105  & n40183;
  assign n16903 = pi107  & n15023;
  assign n16904 = pi106  & n15030;
  assign n16905 = ~n16903 & ~n16904;
  assign n16906 = ~n16902 & ~n16904;
  assign n16907 = ~n16903 & n16906;
  assign n16908 = ~n16902 & n16905;
  assign n16909 = ~n16901 & n40549;
  assign n16910 = pi2  & ~n16909;
  assign n16911 = pi2  & ~n16910;
  assign n16912 = pi2  & n16909;
  assign n16913 = ~n16909 & ~n16910;
  assign n16914 = ~pi2  & ~n16909;
  assign n16915 = ~n40550 & ~n40551;
  assign n16916 = n16900 & ~n16915;
  assign n16917 = n8209 & n15004;
  assign n16918 = pi104  & n40183;
  assign n16919 = pi106  & n15023;
  assign n16920 = pi105  & n15030;
  assign n16921 = ~n16919 & ~n16920;
  assign n16922 = ~n16918 & ~n16920;
  assign n16923 = ~n16919 & n16922;
  assign n16924 = ~n16918 & n16921;
  assign n16925 = ~n16917 & n40552;
  assign n16926 = pi2  & ~n16925;
  assign n16927 = pi2  & ~n16926;
  assign n16928 = pi2  & n16925;
  assign n16929 = ~n16925 & ~n16926;
  assign n16930 = ~pi2  & ~n16925;
  assign n16931 = ~n40553 & ~n40554;
  assign n16932 = n16488 & n40468;
  assign n16933 = ~n16488 & ~n16496;
  assign n16934 = ~n40468 & ~n16496;
  assign n16935 = ~n16933 & ~n16934;
  assign n16936 = ~n16496 & ~n16932;
  assign n16937 = ~n16931 & ~n40555;
  assign n16938 = n16484 & ~n16486;
  assign n16939 = ~n16487 & ~n16938;
  assign n16940 = n8229 & n15004;
  assign n16941 = pi103  & n40183;
  assign n16942 = pi105  & n15023;
  assign n16943 = pi104  & n15030;
  assign n16944 = ~n16942 & ~n16943;
  assign n16945 = ~n16941 & ~n16943;
  assign n16946 = ~n16942 & n16945;
  assign n16947 = ~n16941 & n16944;
  assign n16948 = ~n16940 & n40556;
  assign n16949 = pi2  & ~n16948;
  assign n16950 = pi2  & ~n16949;
  assign n16951 = pi2  & n16948;
  assign n16952 = ~n16948 & ~n16949;
  assign n16953 = ~pi2  & ~n16948;
  assign n16954 = ~n40557 & ~n40558;
  assign n16955 = n16939 & ~n16954;
  assign n16956 = n8136 & n15004;
  assign n16957 = pi102  & n40183;
  assign n16958 = pi104  & n15023;
  assign n16959 = pi103  & n15030;
  assign n16960 = ~n16958 & ~n16959;
  assign n16961 = ~n16957 & ~n16959;
  assign n16962 = ~n16958 & n16961;
  assign n16963 = ~n16957 & n16960;
  assign n16964 = ~n16956 & n40559;
  assign n16965 = pi2  & ~n16964;
  assign n16966 = pi2  & ~n16965;
  assign n16967 = pi2  & n16964;
  assign n16968 = ~n16964 & ~n16965;
  assign n16969 = ~pi2  & ~n16964;
  assign n16970 = ~n40560 & ~n40561;
  assign n16971 = n16475 & n40465;
  assign n16972 = ~n16475 & n40465;
  assign n16973 = n16475 & ~n40465;
  assign n16974 = ~n16972 & ~n16973;
  assign n16975 = ~n16483 & ~n16971;
  assign n16976 = ~n16970 & ~n40562;
  assign n16977 = n16471 & ~n16473;
  assign n16978 = ~n16474 & ~n16977;
  assign n16979 = n6787 & n15004;
  assign n16980 = pi101  & n40183;
  assign n16981 = pi103  & n15023;
  assign n16982 = pi102  & n15030;
  assign n16983 = ~n16981 & ~n16982;
  assign n16984 = ~n16980 & ~n16982;
  assign n16985 = ~n16981 & n16984;
  assign n16986 = ~n16980 & n16983;
  assign n16987 = ~n16979 & n40563;
  assign n16988 = pi2  & ~n16987;
  assign n16989 = pi2  & ~n16988;
  assign n16990 = pi2  & n16987;
  assign n16991 = ~n16987 & ~n16988;
  assign n16992 = ~pi2  & ~n16987;
  assign n16993 = ~n40564 & ~n40565;
  assign n16994 = n16978 & ~n16993;
  assign n16995 = n16467 & ~n16469;
  assign n16996 = ~n16470 & ~n16995;
  assign n16997 = n6819 & n15004;
  assign n16998 = pi100  & n40183;
  assign n16999 = pi102  & n15023;
  assign n17000 = pi101  & n15030;
  assign n17001 = ~n16999 & ~n17000;
  assign n17002 = ~n16998 & ~n17000;
  assign n17003 = ~n16999 & n17002;
  assign n17004 = ~n16998 & n17001;
  assign n17005 = ~n16997 & n40566;
  assign n17006 = pi2  & ~n17005;
  assign n17007 = pi2  & ~n17006;
  assign n17008 = pi2  & n17005;
  assign n17009 = ~n17005 & ~n17006;
  assign n17010 = ~pi2  & ~n17005;
  assign n17011 = ~n40567 & ~n40568;
  assign n17012 = n16996 & ~n17011;
  assign n17013 = n16458 & n40462;
  assign n17014 = ~n16466 & ~n17013;
  assign n17015 = n6839 & n15004;
  assign n17016 = pi99  & n40183;
  assign n17017 = pi101  & n15023;
  assign n17018 = pi100  & n15030;
  assign n17019 = ~n17017 & ~n17018;
  assign n17020 = ~n17016 & ~n17018;
  assign n17021 = ~n17017 & n17020;
  assign n17022 = ~n17016 & n17019;
  assign n17023 = ~n17015 & n40569;
  assign n17024 = pi2  & ~n17023;
  assign n17025 = pi2  & ~n17024;
  assign n17026 = pi2  & n17023;
  assign n17027 = ~n17023 & ~n17024;
  assign n17028 = ~pi2  & ~n17023;
  assign n17029 = ~n40570 & ~n40571;
  assign n17030 = n17014 & ~n17029;
  assign n17031 = n16454 & ~n16456;
  assign n17032 = ~n16457 & ~n17031;
  assign n17033 = n6474 & n15004;
  assign n17034 = pi98  & n40183;
  assign n17035 = pi100  & n15023;
  assign n17036 = pi99  & n15030;
  assign n17037 = ~n17035 & ~n17036;
  assign n17038 = ~n17034 & ~n17036;
  assign n17039 = ~n17035 & n17038;
  assign n17040 = ~n17034 & n17037;
  assign n17041 = ~n17033 & n40572;
  assign n17042 = pi2  & ~n17041;
  assign n17043 = pi2  & ~n17042;
  assign n17044 = pi2  & n17041;
  assign n17045 = ~n17041 & ~n17042;
  assign n17046 = ~pi2  & ~n17041;
  assign n17047 = ~n40573 & ~n40574;
  assign n17048 = n17032 & ~n17047;
  assign n17049 = n5578 & n15004;
  assign n17050 = pi97  & n40183;
  assign n17051 = pi99  & n15023;
  assign n17052 = pi98  & n15030;
  assign n17053 = ~n17051 & ~n17052;
  assign n17054 = ~n17050 & ~n17052;
  assign n17055 = ~n17051 & n17054;
  assign n17056 = ~n17050 & n17053;
  assign n17057 = ~n17049 & n40575;
  assign n17058 = pi2  & ~n17057;
  assign n17059 = pi2  & ~n17058;
  assign n17060 = pi2  & n17057;
  assign n17061 = ~n17057 & ~n17058;
  assign n17062 = ~pi2  & ~n17057;
  assign n17063 = ~n40576 & ~n40577;
  assign n17064 = n16448 & ~n16450;
  assign n17065 = ~n16448 & ~n40459;
  assign n17066 = ~n16449 & n16454;
  assign n17067 = ~n17065 & ~n17066;
  assign n17068 = ~n40459 & ~n17064;
  assign n17069 = ~n17063 & ~n40578;
  assign n17070 = n5610 & n15004;
  assign n17071 = pi96  & n40183;
  assign n17072 = pi98  & n15023;
  assign n17073 = pi97  & n15030;
  assign n17074 = ~n17072 & ~n17073;
  assign n17075 = ~n17071 & ~n17073;
  assign n17076 = ~n17072 & n17075;
  assign n17077 = ~n17071 & n17074;
  assign n17078 = ~n17070 & n40579;
  assign n17079 = pi2  & ~n17078;
  assign n17080 = pi2  & ~n17079;
  assign n17081 = pi2  & n17078;
  assign n17082 = ~n17078 & ~n17079;
  assign n17083 = ~pi2  & ~n17078;
  assign n17084 = ~n40580 & ~n40581;
  assign n17085 = n16442 & ~n16444;
  assign n17086 = ~n16442 & ~n40458;
  assign n17087 = ~n16443 & n16448;
  assign n17088 = ~n17086 & ~n17087;
  assign n17089 = ~n40458 & ~n17085;
  assign n17090 = ~n17084 & ~n40582;
  assign n17091 = n5630 & n15004;
  assign n17092 = pi95  & n40183;
  assign n17093 = pi97  & n15023;
  assign n17094 = pi96  & n15030;
  assign n17095 = ~n17093 & ~n17094;
  assign n17096 = ~n17092 & ~n17094;
  assign n17097 = ~n17093 & n17096;
  assign n17098 = ~n17092 & n17095;
  assign n17099 = ~n17091 & n40583;
  assign n17100 = pi2  & ~n17099;
  assign n17101 = pi2  & ~n17100;
  assign n17102 = pi2  & n17099;
  assign n17103 = ~n17099 & ~n17100;
  assign n17104 = ~pi2  & ~n17099;
  assign n17105 = ~n40584 & ~n40585;
  assign n17106 = n16433 & n40457;
  assign n17107 = ~n16433 & n40457;
  assign n17108 = n16433 & ~n40457;
  assign n17109 = ~n17107 & ~n17108;
  assign n17110 = ~n16441 & ~n17106;
  assign n17111 = ~n17105 & ~n40586;
  assign n17112 = n5281 & n15004;
  assign n17113 = pi94  & n40183;
  assign n17114 = pi96  & n15023;
  assign n17115 = pi95  & n15030;
  assign n17116 = ~n17114 & ~n17115;
  assign n17117 = ~n17113 & ~n17115;
  assign n17118 = ~n17114 & n17117;
  assign n17119 = ~n17113 & n17116;
  assign n17120 = ~n17112 & n40587;
  assign n17121 = pi2  & ~n17120;
  assign n17122 = pi2  & ~n17121;
  assign n17123 = pi2  & n17120;
  assign n17124 = ~n17120 & ~n17121;
  assign n17125 = ~pi2  & ~n17120;
  assign n17126 = ~n40588 & ~n40589;
  assign n17127 = n16427 & ~n16429;
  assign n17128 = ~n16427 & ~n40454;
  assign n17129 = ~n16428 & n16433;
  assign n17130 = ~n17128 & ~n17129;
  assign n17131 = ~n40454 & ~n17127;
  assign n17132 = ~n17126 & ~n40590;
  assign n17133 = n16418 & n40453;
  assign n17134 = ~n16426 & ~n17133;
  assign n17135 = n4494 & n15004;
  assign n17136 = pi93  & n40183;
  assign n17137 = pi95  & n15023;
  assign n17138 = pi94  & n15030;
  assign n17139 = ~n17137 & ~n17138;
  assign n17140 = ~n17136 & ~n17138;
  assign n17141 = ~n17137 & n17140;
  assign n17142 = ~n17136 & n17139;
  assign n17143 = ~n17135 & n40591;
  assign n17144 = pi2  & ~n17143;
  assign n17145 = pi2  & ~n17144;
  assign n17146 = pi2  & n17143;
  assign n17147 = ~n17143 & ~n17144;
  assign n17148 = ~pi2  & ~n17143;
  assign n17149 = ~n40592 & ~n40593;
  assign n17150 = n17134 & ~n17149;
  assign n17151 = n16409 & n40450;
  assign n17152 = ~n16417 & ~n17151;
  assign n17153 = n4524 & n15004;
  assign n17154 = pi92  & n40183;
  assign n17155 = pi94  & n15023;
  assign n17156 = pi93  & n15030;
  assign n17157 = ~n17155 & ~n17156;
  assign n17158 = ~n17154 & ~n17156;
  assign n17159 = ~n17155 & n17158;
  assign n17160 = ~n17154 & n17157;
  assign n17161 = ~n17153 & n40594;
  assign n17162 = pi2  & ~n17161;
  assign n17163 = pi2  & ~n17162;
  assign n17164 = pi2  & n17161;
  assign n17165 = ~n17161 & ~n17162;
  assign n17166 = ~pi2  & ~n17161;
  assign n17167 = ~n40595 & ~n40596;
  assign n17168 = n17152 & ~n17167;
  assign n17169 = n4544 & n15004;
  assign n17170 = pi91  & n40183;
  assign n17171 = pi93  & n15023;
  assign n17172 = pi92  & n15030;
  assign n17173 = ~n17171 & ~n17172;
  assign n17174 = ~n17170 & ~n17172;
  assign n17175 = ~n17171 & n17174;
  assign n17176 = ~n17170 & n17173;
  assign n17177 = ~n17169 & n40597;
  assign n17178 = pi2  & ~n17177;
  assign n17179 = pi2  & ~n17178;
  assign n17180 = pi2  & n17177;
  assign n17181 = ~n17177 & ~n17178;
  assign n17182 = ~pi2  & ~n17177;
  assign n17183 = ~n40598 & ~n40599;
  assign n17184 = n16400 & n40447;
  assign n17185 = ~n16400 & ~n16408;
  assign n17186 = ~n16400 & n40447;
  assign n17187 = ~n40447 & ~n16408;
  assign n17188 = n16400 & ~n40447;
  assign n17189 = ~n40600 & ~n40601;
  assign n17190 = ~n16408 & ~n17184;
  assign n17191 = ~n17183 & ~n40602;
  assign n17192 = n16391 & n40444;
  assign n17193 = ~n16399 & ~n17192;
  assign n17194 = n4453 & n15004;
  assign n17195 = pi90  & n40183;
  assign n17196 = pi92  & n15023;
  assign n17197 = pi91  & n15030;
  assign n17198 = ~n17196 & ~n17197;
  assign n17199 = ~n17195 & ~n17197;
  assign n17200 = ~n17196 & n17199;
  assign n17201 = ~n17195 & n17198;
  assign n17202 = ~n17194 & n40603;
  assign n17203 = pi2  & ~n17202;
  assign n17204 = pi2  & ~n17203;
  assign n17205 = pi2  & n17202;
  assign n17206 = ~n17202 & ~n17203;
  assign n17207 = ~pi2  & ~n17202;
  assign n17208 = ~n40604 & ~n40605;
  assign n17209 = n17193 & ~n17208;
  assign n17210 = n16382 & n40441;
  assign n17211 = ~n16390 & ~n17210;
  assign n17212 = n594 & n15004;
  assign n17213 = pi89  & n40183;
  assign n17214 = pi91  & n15023;
  assign n17215 = pi90  & n15030;
  assign n17216 = ~n17214 & ~n17215;
  assign n17217 = ~n17213 & ~n17215;
  assign n17218 = ~n17214 & n17217;
  assign n17219 = ~n17213 & n17216;
  assign n17220 = ~n17212 & n40606;
  assign n17221 = pi2  & ~n17220;
  assign n17222 = pi2  & ~n17221;
  assign n17223 = pi2  & n17220;
  assign n17224 = ~n17220 & ~n17221;
  assign n17225 = ~pi2  & ~n17220;
  assign n17226 = ~n40607 & ~n40608;
  assign n17227 = n17211 & ~n17226;
  assign n17228 = n3566 & n15004;
  assign n17229 = pi88  & n40183;
  assign n17230 = pi90  & n15023;
  assign n17231 = pi89  & n15030;
  assign n17232 = ~n17230 & ~n17231;
  assign n17233 = ~n17229 & ~n17231;
  assign n17234 = ~n17230 & n17233;
  assign n17235 = ~n17229 & n17232;
  assign n17236 = ~n17228 & n40609;
  assign n17237 = pi2  & ~n17236;
  assign n17238 = pi2  & ~n17237;
  assign n17239 = pi2  & n17236;
  assign n17240 = ~n17236 & ~n17237;
  assign n17241 = ~pi2  & ~n17236;
  assign n17242 = ~n40610 & ~n40611;
  assign n17243 = n16373 & n40438;
  assign n17244 = ~n16373 & n40438;
  assign n17245 = n16373 & ~n40438;
  assign n17246 = ~n17244 & ~n17245;
  assign n17247 = ~n16381 & ~n17243;
  assign n17248 = ~n17242 & ~n40612;
  assign n17249 = n3591 & n15004;
  assign n17250 = pi87  & n40183;
  assign n17251 = pi89  & n15023;
  assign n17252 = pi88  & n15030;
  assign n17253 = ~n17251 & ~n17252;
  assign n17254 = ~n17250 & ~n17252;
  assign n17255 = ~n17251 & n17254;
  assign n17256 = ~n17250 & n17253;
  assign n17257 = ~n17249 & n40613;
  assign n17258 = pi2  & ~n17257;
  assign n17259 = pi2  & ~n17258;
  assign n17260 = pi2  & n17257;
  assign n17261 = ~n17257 & ~n17258;
  assign n17262 = ~pi2  & ~n17257;
  assign n17263 = ~n40614 & ~n40615;
  assign n17264 = n16366 & n40435;
  assign n17265 = ~n16372 & ~n17264;
  assign n17266 = ~n17263 & n17265;
  assign n17267 = n3354 & n15004;
  assign n17268 = pi86  & n40183;
  assign n17269 = pi88  & n15023;
  assign n17270 = pi87  & n15030;
  assign n17271 = ~n17269 & ~n17270;
  assign n17272 = ~n17268 & ~n17270;
  assign n17273 = ~n17269 & n17272;
  assign n17274 = ~n17268 & n17271;
  assign n17275 = ~n17267 & n40616;
  assign n17276 = pi2  & ~n17275;
  assign n17277 = pi2  & ~n17276;
  assign n17278 = pi2  & n17275;
  assign n17279 = ~n17275 & ~n17276;
  assign n17280 = ~pi2  & ~n17275;
  assign n17281 = ~n40617 & ~n40618;
  assign n17282 = n16357 & n40434;
  assign n17283 = ~n16357 & ~n16365;
  assign n17284 = ~n40434 & ~n16365;
  assign n17285 = ~n17283 & ~n17284;
  assign n17286 = ~n16365 & ~n17282;
  assign n17287 = ~n17281 & ~n40619;
  assign n17288 = n16350 & n40431;
  assign n17289 = ~n16356 & ~n17288;
  assign n17290 = n636 & n15004;
  assign n17291 = pi85  & n40183;
  assign n17292 = pi87  & n15023;
  assign n17293 = pi86  & n15030;
  assign n17294 = ~n17292 & ~n17293;
  assign n17295 = ~n17291 & ~n17293;
  assign n17296 = ~n17292 & n17295;
  assign n17297 = ~n17291 & n17294;
  assign n17298 = ~n17290 & n40620;
  assign n17299 = pi2  & ~n17298;
  assign n17300 = pi2  & ~n17299;
  assign n17301 = pi2  & n17298;
  assign n17302 = ~n17298 & ~n17299;
  assign n17303 = ~pi2  & ~n17298;
  assign n17304 = ~n40621 & ~n40622;
  assign n17305 = n17289 & ~n17304;
  assign n17306 = n16341 & n40430;
  assign n17307 = ~n16349 & ~n17306;
  assign n17308 = n2779 & n15004;
  assign n17309 = pi84  & n40183;
  assign n17310 = pi86  & n15023;
  assign n17311 = pi85  & n15030;
  assign n17312 = ~n17310 & ~n17311;
  assign n17313 = ~n17309 & ~n17311;
  assign n17314 = ~n17310 & n17313;
  assign n17315 = ~n17309 & n17312;
  assign n17316 = ~n17308 & n40623;
  assign n17317 = pi2  & ~n17316;
  assign n17318 = pi2  & ~n17317;
  assign n17319 = pi2  & n17316;
  assign n17320 = ~n17316 & ~n17317;
  assign n17321 = ~pi2  & ~n17316;
  assign n17322 = ~n40624 & ~n40625;
  assign n17323 = n17307 & ~n17322;
  assign n17324 = n16332 & n40427;
  assign n17325 = ~n16340 & ~n17324;
  assign n17326 = n2804 & n15004;
  assign n17327 = pi83  & n40183;
  assign n17328 = pi85  & n15023;
  assign n17329 = pi84  & n15030;
  assign n17330 = ~n17328 & ~n17329;
  assign n17331 = ~n17327 & ~n17329;
  assign n17332 = ~n17328 & n17331;
  assign n17333 = ~n17327 & n17330;
  assign n17334 = ~n17326 & n40626;
  assign n17335 = pi2  & ~n17334;
  assign n17336 = pi2  & ~n17335;
  assign n17337 = pi2  & n17334;
  assign n17338 = ~n17334 & ~n17335;
  assign n17339 = ~pi2  & ~n17334;
  assign n17340 = ~n40627 & ~n40628;
  assign n17341 = n17325 & ~n17340;
  assign n17342 = n2591 & n15004;
  assign n17343 = pi82  & n40183;
  assign n17344 = pi84  & n15023;
  assign n17345 = pi83  & n15030;
  assign n17346 = ~n17344 & ~n17345;
  assign n17347 = ~n17343 & ~n17345;
  assign n17348 = ~n17344 & n17347;
  assign n17349 = ~n17343 & n17346;
  assign n17350 = ~n17342 & n40629;
  assign n17351 = pi2  & ~n17350;
  assign n17352 = pi2  & ~n17351;
  assign n17353 = pi2  & n17350;
  assign n17354 = ~n17350 & ~n17351;
  assign n17355 = ~pi2  & ~n17350;
  assign n17356 = ~n40630 & ~n40631;
  assign n17357 = n16323 & n40424;
  assign n17358 = ~n16323 & ~n16331;
  assign n17359 = ~n16323 & n40424;
  assign n17360 = ~n40424 & ~n16331;
  assign n17361 = n16323 & ~n40424;
  assign n17362 = ~n40632 & ~n40633;
  assign n17363 = ~n16331 & ~n17357;
  assign n17364 = ~n17356 & ~n40634;
  assign n17365 = n16314 & n40421;
  assign n17366 = ~n16322 & ~n17365;
  assign n17367 = n2091 & n15004;
  assign n17368 = pi81  & n40183;
  assign n17369 = pi83  & n15023;
  assign n17370 = pi82  & n15030;
  assign n17371 = ~n17369 & ~n17370;
  assign n17372 = ~n17368 & ~n17370;
  assign n17373 = ~n17369 & n17372;
  assign n17374 = ~n17368 & n17371;
  assign n17375 = ~n17367 & n40635;
  assign n17376 = pi2  & ~n17375;
  assign n17377 = pi2  & ~n17376;
  assign n17378 = pi2  & n17375;
  assign n17379 = ~n17375 & ~n17376;
  assign n17380 = ~pi2  & ~n17375;
  assign n17381 = ~n40636 & ~n40637;
  assign n17382 = n17366 & ~n17381;
  assign n17383 = n16310 & ~n16312;
  assign n17384 = ~n16313 & ~n17383;
  assign n17385 = n2134 & n15004;
  assign n17386 = pi80  & n40183;
  assign n17387 = pi82  & n15023;
  assign n17388 = pi81  & n15030;
  assign n17389 = ~n17387 & ~n17388;
  assign n17390 = ~n17386 & ~n17388;
  assign n17391 = ~n17387 & n17390;
  assign n17392 = ~n17386 & n17389;
  assign n17393 = ~n17385 & n40638;
  assign n17394 = pi2  & ~n17393;
  assign n17395 = pi2  & ~n17394;
  assign n17396 = pi2  & n17393;
  assign n17397 = ~n17393 & ~n17394;
  assign n17398 = ~pi2  & ~n17393;
  assign n17399 = ~n40639 & ~n40640;
  assign n17400 = n17384 & ~n17399;
  assign n17401 = n16306 & ~n16308;
  assign n17402 = ~n16309 & ~n17401;
  assign n17403 = n2154 & n15004;
  assign n17404 = pi79  & n40183;
  assign n17405 = pi81  & n15023;
  assign n17406 = pi80  & n15030;
  assign n17407 = ~n17405 & ~n17406;
  assign n17408 = ~n17404 & ~n17406;
  assign n17409 = ~n17405 & n17408;
  assign n17410 = ~n17404 & n17407;
  assign n17411 = ~n17403 & n40641;
  assign n17412 = pi2  & ~n17411;
  assign n17413 = pi2  & ~n17412;
  assign n17414 = pi2  & n17411;
  assign n17415 = ~n17411 & ~n17412;
  assign n17416 = ~pi2  & ~n17411;
  assign n17417 = ~n40642 & ~n40643;
  assign n17418 = n17402 & ~n17417;
  assign n17419 = n2063 & n15004;
  assign n17420 = pi78  & n40183;
  assign n17421 = pi80  & n15023;
  assign n17422 = pi79  & n15030;
  assign n17423 = ~n17421 & ~n17422;
  assign n17424 = ~n17420 & ~n17422;
  assign n17425 = ~n17421 & n17424;
  assign n17426 = ~n17420 & n17423;
  assign n17427 = ~n17419 & n40644;
  assign n17428 = pi2  & ~n17427;
  assign n17429 = pi2  & ~n17428;
  assign n17430 = pi2  & n17427;
  assign n17431 = ~n17427 & ~n17428;
  assign n17432 = ~pi2  & ~n17427;
  assign n17433 = ~n40645 & ~n40646;
  assign n17434 = n16302 & ~n16304;
  assign n17435 = ~n16305 & ~n17434;
  assign n17436 = ~n17433 & n17435;
  assign n17437 = n678 & n15004;
  assign n17438 = pi77  & n40183;
  assign n17439 = pi79  & n15023;
  assign n17440 = pi78  & n15030;
  assign n17441 = ~n17439 & ~n17440;
  assign n17442 = ~n17438 & ~n17440;
  assign n17443 = ~n17439 & n17442;
  assign n17444 = ~n17438 & n17441;
  assign n17445 = ~n17437 & n40647;
  assign n17446 = pi2  & ~n17445;
  assign n17447 = pi2  & ~n17446;
  assign n17448 = pi2  & n17445;
  assign n17449 = ~n17445 & ~n17446;
  assign n17450 = ~pi2  & ~n17445;
  assign n17451 = ~n40648 & ~n40649;
  assign n17452 = n16293 & ~n40417;
  assign n17453 = ~n40416 & n17452;
  assign n17454 = n16293 & n40418;
  assign n17455 = ~n16301 & ~n40650;
  assign n17456 = ~n17451 & n17455;
  assign n17457 = n1578 & n15004;
  assign n17458 = pi76  & n40183;
  assign n17459 = pi78  & n15023;
  assign n17460 = pi77  & n15030;
  assign n17461 = ~n17459 & ~n17460;
  assign n17462 = ~n17458 & ~n17460;
  assign n17463 = ~n17459 & n17462;
  assign n17464 = ~n17458 & n17461;
  assign n17465 = ~n17457 & n40651;
  assign n17466 = pi2  & ~n17465;
  assign n17467 = pi2  & ~n17466;
  assign n17468 = pi2  & n17465;
  assign n17469 = ~n17465 & ~n17466;
  assign n17470 = ~pi2  & ~n17465;
  assign n17471 = ~n40652 & ~n40653;
  assign n17472 = n16289 & ~n16291;
  assign n17473 = ~n16292 & ~n17472;
  assign n17474 = ~n17471 & n17473;
  assign n17475 = n1596 & n15004;
  assign n17476 = pi75  & n40183;
  assign n17477 = pi77  & n15023;
  assign n17478 = pi76  & n15030;
  assign n17479 = ~n17477 & ~n17478;
  assign n17480 = ~n17476 & ~n17478;
  assign n17481 = ~n17477 & n17480;
  assign n17482 = ~n17476 & n17479;
  assign n17483 = ~n17475 & n40654;
  assign n17484 = pi2  & ~n17483;
  assign n17485 = pi2  & ~n17484;
  assign n17486 = pi2  & n17483;
  assign n17487 = ~n17483 & ~n17484;
  assign n17488 = ~pi2  & ~n17483;
  assign n17489 = ~n40655 & ~n40656;
  assign n17490 = n16283 & ~n16285;
  assign n17491 = ~n16283 & ~n40415;
  assign n17492 = ~n16284 & n16289;
  assign n17493 = ~n17491 & ~n17492;
  assign n17494 = ~n40415 & ~n17490;
  assign n17495 = ~n17489 & ~n40657;
  assign n17496 = ~n16079 & n16281;
  assign n17497 = ~n16282 & ~n17496;
  assign n17498 = n1465 & n15004;
  assign n17499 = pi74  & n40183;
  assign n17500 = pi76  & n15023;
  assign n17501 = pi75  & n15030;
  assign n17502 = ~n17500 & ~n17501;
  assign n17503 = ~n17499 & ~n17501;
  assign n17504 = ~n17500 & n17503;
  assign n17505 = ~n17499 & n17502;
  assign n17506 = ~n17498 & n40658;
  assign n17507 = pi2  & ~n17506;
  assign n17508 = pi2  & ~n17507;
  assign n17509 = pi2  & n17506;
  assign n17510 = ~n17506 & ~n17507;
  assign n17511 = ~pi2  & ~n17506;
  assign n17512 = ~n40659 & ~n40660;
  assign n17513 = n17497 & ~n17512;
  assign n17514 = n720 & n15004;
  assign n17515 = pi73  & n40183;
  assign n17516 = pi75  & n15023;
  assign n17517 = pi74  & n15030;
  assign n17518 = ~n17516 & ~n17517;
  assign n17519 = ~n17515 & ~n17517;
  assign n17520 = ~n17516 & n17519;
  assign n17521 = ~n17515 & n17518;
  assign n17522 = ~n17514 & n40661;
  assign n17523 = pi2  & ~n17522;
  assign n17524 = pi2  & ~n17523;
  assign n17525 = pi2  & n17522;
  assign n17526 = ~n17522 & ~n17523;
  assign n17527 = ~pi2  & ~n17522;
  assign n17528 = ~n40662 & ~n40663;
  assign n17529 = n16272 & n40414;
  assign n17530 = ~n16272 & ~n16280;
  assign n17531 = ~n16272 & n40414;
  assign n17532 = ~n40414 & ~n16280;
  assign n17533 = n16272 & ~n40414;
  assign n17534 = ~n40664 & ~n40665;
  assign n17535 = ~n16280 & ~n17529;
  assign n17536 = ~n17528 & ~n40666;
  assign n17537 = n16263 & n40411;
  assign n17538 = ~n16271 & ~n17537;
  assign n17539 = n1218 & n15004;
  assign n17540 = pi72  & n40183;
  assign n17541 = pi74  & n15023;
  assign n17542 = pi73  & n15030;
  assign n17543 = ~n17541 & ~n17542;
  assign n17544 = ~n17540 & ~n17542;
  assign n17545 = ~n17541 & n17544;
  assign n17546 = ~n17540 & n17543;
  assign n17547 = ~n17539 & n40667;
  assign n17548 = pi2  & ~n17547;
  assign n17549 = pi2  & ~n17548;
  assign n17550 = pi2  & n17547;
  assign n17551 = ~n17547 & ~n17548;
  assign n17552 = ~pi2  & ~n17547;
  assign n17553 = ~n40668 & ~n40669;
  assign n17554 = n17538 & ~n17553;
  assign n17555 = n16254 & n40408;
  assign n17556 = ~n16262 & ~n17555;
  assign n17557 = n1238 & n15004;
  assign n17558 = pi71  & n40183;
  assign n17559 = pi73  & n15023;
  assign n17560 = pi72  & n15030;
  assign n17561 = ~n17559 & ~n17560;
  assign n17562 = ~n17558 & ~n17560;
  assign n17563 = ~n17559 & n17562;
  assign n17564 = ~n17558 & n17561;
  assign n17565 = ~n17557 & n40670;
  assign n17566 = pi2  & ~n17565;
  assign n17567 = pi2  & ~n17566;
  assign n17568 = pi2  & n17565;
  assign n17569 = ~n17565 & ~n17566;
  assign n17570 = ~pi2  & ~n17565;
  assign n17571 = ~n40671 & ~n40672;
  assign n17572 = n17556 & ~n17571;
  assign n17573 = n16245 & n40405;
  assign n17574 = ~n16253 & ~n17573;
  assign n17575 = n1124 & n15004;
  assign n17576 = pi70  & n40183;
  assign n17577 = pi72  & n15023;
  assign n17578 = pi71  & n15030;
  assign n17579 = ~n17577 & ~n17578;
  assign n17580 = ~n17576 & ~n17578;
  assign n17581 = ~n17577 & n17580;
  assign n17582 = ~n17576 & n17579;
  assign n17583 = ~n17575 & n40673;
  assign n17584 = pi2  & ~n17583;
  assign n17585 = pi2  & ~n17584;
  assign n17586 = pi2  & n17583;
  assign n17587 = ~n17583 & ~n17584;
  assign n17588 = ~pi2  & ~n17583;
  assign n17589 = ~n40674 & ~n40675;
  assign n17590 = n17574 & ~n17589;
  assign n17591 = n927 & n15004;
  assign n17592 = pi69  & n40183;
  assign n17593 = pi71  & n15023;
  assign n17594 = pi70  & n15030;
  assign n17595 = ~n17593 & ~n17594;
  assign n17596 = ~n17592 & ~n17594;
  assign n17597 = ~n17593 & n17596;
  assign n17598 = ~n17592 & n17595;
  assign n17599 = ~n17591 & n40676;
  assign n17600 = pi2  & ~n17599;
  assign n17601 = pi2  & ~n17600;
  assign n17602 = pi2  & n17599;
  assign n17603 = ~n17599 & ~n17600;
  assign n17604 = ~pi2  & ~n17599;
  assign n17605 = ~n40677 & ~n40678;
  assign n17606 = n16236 & n40402;
  assign n17607 = ~n16244 & ~n17606;
  assign n17608 = ~n17605 & n17607;
  assign n17609 = n972 & n15004;
  assign n17610 = pi68  & n40183;
  assign n17611 = pi70  & n15023;
  assign n17612 = pi69  & n15030;
  assign n17613 = ~n17611 & ~n17612;
  assign n17614 = ~n17610 & ~n17612;
  assign n17615 = ~n17611 & n17614;
  assign n17616 = ~n17610 & n17613;
  assign n17617 = ~n17609 & n40679;
  assign n17618 = pi2  & ~n17617;
  assign n17619 = pi2  & ~n17618;
  assign n17620 = pi2  & n17617;
  assign n17621 = ~n17617 & ~n17618;
  assign n17622 = ~pi2  & ~n17617;
  assign n17623 = ~n40680 & ~n40681;
  assign n17624 = n16227 & n40399;
  assign n17625 = n16227 & ~n40399;
  assign n17626 = ~n16227 & n40399;
  assign n17627 = ~n17625 & ~n17626;
  assign n17628 = ~n16235 & ~n17624;
  assign n17629 = ~n17623 & ~n40682;
  assign n17630 = n990 & n15004;
  assign n17631 = pi67  & n40183;
  assign n17632 = pi69  & n15023;
  assign n17633 = pi68  & n15030;
  assign n17634 = ~n17632 & ~n17633;
  assign n17635 = ~n17631 & ~n17633;
  assign n17636 = ~n17632 & n17635;
  assign n17637 = ~n17631 & n17634;
  assign n17638 = ~n17630 & n40683;
  assign n17639 = pi2  & ~n17638;
  assign n17640 = pi2  & ~n17639;
  assign n17641 = pi2  & n17638;
  assign n17642 = ~n17638 & ~n17639;
  assign n17643 = ~pi2  & ~n17638;
  assign n17644 = ~n40684 & ~n40685;
  assign n17645 = pi5  & ~n40389;
  assign n17646 = n40392 & ~n17645;
  assign n17647 = ~n40392 & n17645;
  assign n17648 = ~n40389 & n16209;
  assign n17649 = ~n40393 & ~n17648;
  assign n17650 = ~n17646 & ~n17647;
  assign n17651 = ~n17644 & n40686;
  assign n17652 = n871 & n15004;
  assign n17653 = pi66  & n40183;
  assign n17654 = pi68  & n15023;
  assign n17655 = pi67  & n15030;
  assign n17656 = ~n17654 & ~n17655;
  assign n17657 = ~n17653 & ~n17655;
  assign n17658 = ~n17654 & n17657;
  assign n17659 = ~n17653 & n17656;
  assign n17660 = ~n17652 & n40687;
  assign n17661 = pi2  & ~n17660;
  assign n17662 = pi2  & ~n17661;
  assign n17663 = pi2  & n17660;
  assign n17664 = ~n17660 & ~n17661;
  assign n17665 = ~pi2  & ~n17660;
  assign n17666 = ~n40688 & ~n40689;
  assign n17667 = pi5  & n16183;
  assign n17668 = ~n16182 & n17667;
  assign n17669 = n16182 & ~n17667;
  assign n17670 = ~n16184 & n16188;
  assign n17671 = ~n40389 & ~n17670;
  assign n17672 = ~n17668 & ~n17669;
  assign n17673 = ~n17666 & n40690;
  assign n17674 = n847 & n15004;
  assign n17675 = pi65  & n40183;
  assign n17676 = pi67  & n15023;
  assign n17677 = pi66  & n15030;
  assign n17678 = ~n17676 & ~n17677;
  assign n17679 = ~n17675 & ~n17677;
  assign n17680 = ~n17676 & n17679;
  assign n17681 = ~n17675 & n17678;
  assign n17682 = ~n17674 & n40691;
  assign n17683 = pi2  & ~n17682;
  assign n17684 = pi2  & ~n17683;
  assign n17685 = pi2  & n17682;
  assign n17686 = ~n17682 & ~n17683;
  assign n17687 = ~pi2  & ~n17682;
  assign n17688 = ~n40692 & ~n40693;
  assign n17689 = n16183 & ~n17688;
  assign n17690 = ~n16183 & n17688;
  assign n17691 = ~n17689 & ~n17690;
  assign n17692 = n37515 & n15004;
  assign n17693 = pi65  & n15023;
  assign n17694 = pi64  & n15030;
  assign n17695 = ~n17693 & ~n17694;
  assign n17696 = ~n17692 & n17695;
  assign po0  = pi0  & pi64 ;
  assign n17698 = pi2  & ~po0 ;
  assign n17699 = pi2  & ~n17696;
  assign n17700 = pi2  & ~n17699;
  assign n17701 = ~n17696 & ~n17699;
  assign n17702 = ~n17700 & ~n17701;
  assign n17703 = n17698 & ~n17702;
  assign n17704 = n17696 & n17698;
  assign n17705 = pi64  & n40183;
  assign n17706 = pi65  & n15030;
  assign n17707 = ~n17705 & ~n17706;
  assign n17708 = pi66  & n15023;
  assign n17709 = ~n37521 & n15004;
  assign n17710 = ~n17708 & ~n17709;
  assign n17711 = ~n17706 & ~n17708;
  assign n17712 = n17707 & ~n17708;
  assign n17713 = ~n17705 & n17711;
  assign n17714 = ~n17709 & n40695;
  assign n17715 = n17707 & n17710;
  assign n17716 = pi2  & ~n40696;
  assign n17717 = pi2  & ~n17716;
  assign n17718 = ~n40696 & ~n17716;
  assign n17719 = ~n17717 & ~n17718;
  assign n17720 = n40694 & ~n17719;
  assign n17721 = n40694 & n40696;
  assign n17722 = n17691 & n40697;
  assign n17723 = ~n17689 & ~n17722;
  assign n17724 = n17666 & ~n40690;
  assign n17725 = n40690 & ~n17673;
  assign n17726 = n17666 & n40690;
  assign n17727 = ~n17666 & ~n17673;
  assign n17728 = ~n17666 & ~n40690;
  assign n17729 = ~n40698 & ~n40699;
  assign n17730 = ~n17673 & ~n17724;
  assign n17731 = ~n17723 & ~n40700;
  assign n17732 = ~n17673 & ~n17731;
  assign n17733 = n17644 & ~n40686;
  assign n17734 = n40686 & ~n17651;
  assign n17735 = n17644 & n40686;
  assign n17736 = ~n17644 & ~n17651;
  assign n17737 = ~n17644 & ~n40686;
  assign n17738 = ~n40701 & ~n40702;
  assign n17739 = ~n17651 & ~n17733;
  assign n17740 = ~n17732 & ~n40703;
  assign n17741 = ~n17651 & ~n17740;
  assign n17742 = n17623 & n40682;
  assign n17743 = ~n17629 & ~n17742;
  assign n17744 = ~n17741 & n17743;
  assign n17745 = ~n17629 & ~n17744;
  assign n17746 = n17605 & ~n17607;
  assign n17747 = ~n17608 & ~n17746;
  assign n17748 = ~n17745 & n17747;
  assign n17749 = ~n17608 & ~n17748;
  assign n17750 = ~n17574 & n17589;
  assign n17751 = n17574 & ~n17590;
  assign n17752 = n17574 & n17589;
  assign n17753 = ~n17589 & ~n17590;
  assign n17754 = ~n17574 & ~n17589;
  assign n17755 = ~n40704 & ~n40705;
  assign n17756 = ~n17590 & ~n17750;
  assign n17757 = ~n17749 & ~n40706;
  assign n17758 = ~n17590 & ~n17757;
  assign n17759 = ~n17556 & n17571;
  assign n17760 = n17556 & ~n17572;
  assign n17761 = n17556 & n17571;
  assign n17762 = ~n17571 & ~n17572;
  assign n17763 = ~n17556 & ~n17571;
  assign n17764 = ~n40707 & ~n40708;
  assign n17765 = ~n17572 & ~n17759;
  assign n17766 = ~n17758 & ~n40709;
  assign n17767 = ~n17572 & ~n17766;
  assign n17768 = ~n17538 & n17553;
  assign n17769 = ~n17554 & ~n17768;
  assign n17770 = ~n17767 & n17769;
  assign n17771 = ~n17554 & ~n17770;
  assign n17772 = n17528 & n40666;
  assign n17773 = n17528 & ~n40666;
  assign n17774 = ~n17528 & n40666;
  assign n17775 = ~n17773 & ~n17774;
  assign n17776 = ~n17536 & ~n17772;
  assign n17777 = ~n17771 & ~n40710;
  assign n17778 = ~n17536 & ~n17777;
  assign n17779 = ~n17497 & n17512;
  assign n17780 = n17497 & ~n17513;
  assign n17781 = n17497 & n17512;
  assign n17782 = ~n17512 & ~n17513;
  assign n17783 = ~n17497 & ~n17512;
  assign n17784 = ~n40711 & ~n40712;
  assign n17785 = ~n17513 & ~n17779;
  assign n17786 = ~n17778 & ~n40713;
  assign n17787 = ~n17513 & ~n17786;
  assign n17788 = n17489 & n40657;
  assign n17789 = n17489 & ~n40657;
  assign n17790 = ~n17489 & n40657;
  assign n17791 = ~n17789 & ~n17790;
  assign n17792 = ~n17495 & ~n17788;
  assign n17793 = ~n17787 & ~n40714;
  assign n17794 = ~n17495 & ~n17793;
  assign n17795 = n17471 & ~n17473;
  assign n17796 = n17471 & n17473;
  assign n17797 = ~n17471 & ~n17473;
  assign n17798 = ~n17796 & ~n17797;
  assign n17799 = ~n17474 & ~n17795;
  assign n17800 = ~n17794 & ~n40715;
  assign n17801 = ~n17474 & ~n17800;
  assign n17802 = n17451 & ~n17455;
  assign n17803 = ~n17451 & ~n17456;
  assign n17804 = ~n17451 & ~n17455;
  assign n17805 = n17455 & ~n17456;
  assign n17806 = n17451 & n17455;
  assign n17807 = ~n40716 & ~n40717;
  assign n17808 = ~n17456 & ~n17802;
  assign n17809 = ~n17801 & ~n40718;
  assign n17810 = ~n17456 & ~n17809;
  assign n17811 = n17433 & ~n17435;
  assign n17812 = n17433 & n17435;
  assign n17813 = ~n17433 & ~n17435;
  assign n17814 = ~n17812 & ~n17813;
  assign n17815 = ~n17436 & ~n17811;
  assign n17816 = ~n17810 & ~n40719;
  assign n17817 = ~n17436 & ~n17816;
  assign n17818 = ~n17402 & n17417;
  assign n17819 = n17402 & ~n17418;
  assign n17820 = n17402 & n17417;
  assign n17821 = ~n17417 & ~n17418;
  assign n17822 = ~n17402 & ~n17417;
  assign n17823 = ~n40720 & ~n40721;
  assign n17824 = ~n17418 & ~n17818;
  assign n17825 = ~n17817 & ~n40722;
  assign n17826 = ~n17418 & ~n17825;
  assign n17827 = ~n17384 & n17399;
  assign n17828 = n17384 & ~n17400;
  assign n17829 = n17384 & n17399;
  assign n17830 = ~n17399 & ~n17400;
  assign n17831 = ~n17384 & ~n17399;
  assign n17832 = ~n40723 & ~n40724;
  assign n17833 = ~n17400 & ~n17827;
  assign n17834 = ~n17826 & ~n40725;
  assign n17835 = ~n17400 & ~n17834;
  assign n17836 = ~n17366 & n17381;
  assign n17837 = n17366 & ~n17382;
  assign n17838 = n17366 & n17381;
  assign n17839 = ~n17381 & ~n17382;
  assign n17840 = ~n17366 & ~n17381;
  assign n17841 = ~n40726 & ~n40727;
  assign n17842 = ~n17382 & ~n17836;
  assign n17843 = ~n17835 & ~n40728;
  assign n17844 = ~n17382 & ~n17843;
  assign n17845 = n17356 & n40634;
  assign n17846 = ~n40634 & ~n17364;
  assign n17847 = ~n17356 & ~n17364;
  assign n17848 = ~n17846 & ~n17847;
  assign n17849 = ~n17364 & ~n17845;
  assign n17850 = ~n17844 & ~n40729;
  assign n17851 = ~n17364 & ~n17850;
  assign n17852 = ~n17325 & n17340;
  assign n17853 = n17325 & ~n17341;
  assign n17854 = n17325 & n17340;
  assign n17855 = ~n17340 & ~n17341;
  assign n17856 = ~n17325 & ~n17340;
  assign n17857 = ~n40730 & ~n40731;
  assign n17858 = ~n17341 & ~n17852;
  assign n17859 = ~n17851 & ~n40732;
  assign n17860 = ~n17341 & ~n17859;
  assign n17861 = ~n17307 & n17322;
  assign n17862 = ~n17323 & ~n17861;
  assign n17863 = ~n17860 & n17862;
  assign n17864 = ~n17323 & ~n17863;
  assign n17865 = ~n17289 & n17304;
  assign n17866 = n17289 & ~n17305;
  assign n17867 = n17289 & n17304;
  assign n17868 = ~n17304 & ~n17305;
  assign n17869 = ~n17289 & ~n17304;
  assign n17870 = ~n40733 & ~n40734;
  assign n17871 = ~n17305 & ~n17865;
  assign n17872 = ~n17864 & ~n40735;
  assign n17873 = ~n17305 & ~n17872;
  assign n17874 = n17281 & n40619;
  assign n17875 = ~n40619 & ~n17287;
  assign n17876 = n17281 & ~n40619;
  assign n17877 = ~n17281 & ~n17287;
  assign n17878 = ~n17281 & n40619;
  assign n17879 = ~n40736 & ~n40737;
  assign n17880 = ~n17287 & ~n17874;
  assign n17881 = ~n17873 & ~n40738;
  assign n17882 = ~n17287 & ~n17881;
  assign n17883 = n17263 & ~n17265;
  assign n17884 = ~n17266 & ~n17883;
  assign n17885 = ~n17882 & n17884;
  assign n17886 = ~n17266 & ~n17885;
  assign n17887 = n17242 & n40612;
  assign n17888 = ~n17248 & ~n17887;
  assign n17889 = ~n17886 & n17888;
  assign n17890 = ~n17248 & ~n17889;
  assign n17891 = ~n17211 & n17226;
  assign n17892 = ~n17227 & ~n17891;
  assign n17893 = ~n17890 & n17892;
  assign n17894 = ~n17227 & ~n17893;
  assign n17895 = ~n17193 & n17208;
  assign n17896 = ~n17209 & ~n17895;
  assign n17897 = ~n17894 & n17896;
  assign n17898 = ~n17209 & ~n17897;
  assign n17899 = n17183 & n40602;
  assign n17900 = ~n40602 & ~n17191;
  assign n17901 = ~n17183 & ~n17191;
  assign n17902 = ~n17900 & ~n17901;
  assign n17903 = ~n17191 & ~n17899;
  assign n17904 = ~n17898 & ~n40739;
  assign n17905 = ~n17191 & ~n17904;
  assign n17906 = ~n17152 & n17167;
  assign n17907 = n17152 & ~n17168;
  assign n17908 = n17152 & n17167;
  assign n17909 = ~n17167 & ~n17168;
  assign n17910 = ~n17152 & ~n17167;
  assign n17911 = ~n40740 & ~n40741;
  assign n17912 = ~n17168 & ~n17906;
  assign n17913 = ~n17905 & ~n40742;
  assign n17914 = ~n17168 & ~n17913;
  assign n17915 = ~n17134 & n17149;
  assign n17916 = n17134 & ~n17150;
  assign n17917 = n17134 & n17149;
  assign n17918 = ~n17149 & ~n17150;
  assign n17919 = ~n17134 & ~n17149;
  assign n17920 = ~n40743 & ~n40744;
  assign n17921 = ~n17150 & ~n17915;
  assign n17922 = ~n17914 & ~n40745;
  assign n17923 = ~n17150 & ~n17922;
  assign n17924 = n17126 & n40590;
  assign n17925 = n17126 & ~n40590;
  assign n17926 = ~n17126 & n40590;
  assign n17927 = ~n17925 & ~n17926;
  assign n17928 = ~n17132 & ~n17924;
  assign n17929 = ~n17923 & ~n40746;
  assign n17930 = ~n17132 & ~n17929;
  assign n17931 = n17105 & n40586;
  assign n17932 = ~n17111 & ~n17931;
  assign n17933 = ~n17930 & n17932;
  assign n17934 = ~n17111 & ~n17933;
  assign n17935 = n17084 & n40582;
  assign n17936 = n17084 & ~n40582;
  assign n17937 = ~n17084 & n40582;
  assign n17938 = ~n17936 & ~n17937;
  assign n17939 = ~n17090 & ~n17935;
  assign n17940 = ~n17934 & ~n40747;
  assign n17941 = ~n17090 & ~n17940;
  assign n17942 = n17063 & n40578;
  assign n17943 = n17063 & ~n40578;
  assign n17944 = ~n17063 & n40578;
  assign n17945 = ~n17943 & ~n17944;
  assign n17946 = ~n17069 & ~n17942;
  assign n17947 = ~n17941 & ~n40748;
  assign n17948 = ~n17069 & ~n17947;
  assign n17949 = ~n17032 & n17047;
  assign n17950 = n17032 & ~n17048;
  assign n17951 = n17032 & n17047;
  assign n17952 = ~n17047 & ~n17048;
  assign n17953 = ~n17032 & ~n17047;
  assign n17954 = ~n40749 & ~n40750;
  assign n17955 = ~n17048 & ~n17949;
  assign n17956 = ~n17948 & ~n40751;
  assign n17957 = ~n17048 & ~n17956;
  assign n17958 = ~n17014 & n17029;
  assign n17959 = ~n17030 & ~n17958;
  assign n17960 = ~n17957 & n17959;
  assign n17961 = ~n17030 & ~n17960;
  assign n17962 = ~n16996 & n17011;
  assign n17963 = n16996 & ~n17012;
  assign n17964 = n16996 & n17011;
  assign n17965 = ~n17011 & ~n17012;
  assign n17966 = ~n16996 & ~n17011;
  assign n17967 = ~n40752 & ~n40753;
  assign n17968 = ~n17012 & ~n17962;
  assign n17969 = ~n17961 & ~n40754;
  assign n17970 = ~n17012 & ~n17969;
  assign n17971 = ~n16978 & n16993;
  assign n17972 = n16978 & ~n16994;
  assign n17973 = n16978 & n16993;
  assign n17974 = ~n16993 & ~n16994;
  assign n17975 = ~n16978 & ~n16993;
  assign n17976 = ~n40755 & ~n40756;
  assign n17977 = ~n16994 & ~n17971;
  assign n17978 = ~n17970 & ~n40757;
  assign n17979 = ~n16994 & ~n17978;
  assign n17980 = n16970 & n40562;
  assign n17981 = ~n16976 & ~n17980;
  assign n17982 = ~n17979 & n17981;
  assign n17983 = ~n16976 & ~n17982;
  assign n17984 = ~n16939 & n16954;
  assign n17985 = ~n16955 & ~n17984;
  assign n17986 = ~n17983 & n17985;
  assign n17987 = ~n16955 & ~n17986;
  assign n17988 = n16931 & n40555;
  assign n17989 = ~n40555 & ~n16937;
  assign n17990 = n16931 & ~n40555;
  assign n17991 = ~n16931 & ~n16937;
  assign n17992 = ~n16931 & n40555;
  assign n17993 = ~n40758 & ~n40759;
  assign n17994 = ~n16937 & ~n17988;
  assign n17995 = ~n17987 & ~n40760;
  assign n17996 = ~n16937 & ~n17995;
  assign n17997 = ~n16900 & n16915;
  assign n17998 = n16900 & ~n16916;
  assign n17999 = n16900 & n16915;
  assign n18000 = ~n16915 & ~n16916;
  assign n18001 = ~n16900 & ~n16915;
  assign n18002 = ~n40761 & ~n40762;
  assign n18003 = ~n16916 & ~n17997;
  assign n18004 = ~n17996 & ~n40763;
  assign n18005 = ~n16916 & ~n18004;
  assign n18006 = n16890 & n40548;
  assign n18007 = n16890 & ~n40548;
  assign n18008 = ~n16890 & n40548;
  assign n18009 = ~n18007 & ~n18008;
  assign n18010 = ~n16898 & ~n18006;
  assign n18011 = ~n18005 & ~n40764;
  assign n18012 = ~n16898 & ~n18011;
  assign n18013 = ~n16859 & n16874;
  assign n18014 = ~n16875 & ~n18013;
  assign n18015 = ~n18012 & n18014;
  assign n18016 = ~n16875 & ~n18015;
  assign n18017 = ~n16841 & n16856;
  assign n18018 = n16841 & ~n16857;
  assign n18019 = n16841 & n16856;
  assign n18020 = ~n16856 & ~n16857;
  assign n18021 = ~n16841 & ~n16856;
  assign n18022 = ~n40765 & ~n40766;
  assign n18023 = ~n16857 & ~n18017;
  assign n18024 = ~n18016 & ~n40767;
  assign n18025 = ~n16857 & ~n18024;
  assign n18026 = ~n16823 & n16838;
  assign n18027 = n16823 & ~n16839;
  assign n18028 = n16823 & n16838;
  assign n18029 = ~n16838 & ~n16839;
  assign n18030 = ~n16823 & ~n16838;
  assign n18031 = ~n40768 & ~n40769;
  assign n18032 = ~n16839 & ~n18026;
  assign n18033 = ~n18025 & ~n40770;
  assign n18034 = ~n16839 & ~n18033;
  assign n18035 = n16818 & ~n16820;
  assign n18036 = ~n16821 & ~n18035;
  assign n18037 = ~n18034 & n18036;
  assign n18038 = ~n16821 & ~n18037;
  assign n18039 = ~n16787 & n16802;
  assign n18040 = ~n16803 & ~n18039;
  assign n18041 = ~n18038 & n18040;
  assign n18042 = ~n16803 & ~n18041;
  assign n18043 = ~n16769 & n16784;
  assign n18044 = n16769 & ~n16785;
  assign n18045 = n16769 & n16784;
  assign n18046 = ~n16784 & ~n16785;
  assign n18047 = ~n16769 & ~n16784;
  assign n18048 = ~n40771 & ~n40772;
  assign n18049 = ~n16785 & ~n18043;
  assign n18050 = ~n18042 & ~n40773;
  assign n18051 = ~n16785 & ~n18050;
  assign n18052 = n16764 & ~n16766;
  assign n18053 = ~n16767 & ~n18052;
  assign n18054 = ~n18051 & n18053;
  assign n18055 = ~n16767 & ~n18054;
  assign n18056 = n16743 & n40521;
  assign n18057 = ~n16749 & ~n18056;
  assign n18058 = ~n18055 & n18057;
  assign n18059 = ~n16749 & ~n18058;
  assign n18060 = n16722 & n40517;
  assign n18061 = n16722 & ~n40517;
  assign n18062 = ~n16722 & n40517;
  assign n18063 = ~n18061 & ~n18062;
  assign n18064 = ~n16728 & ~n18060;
  assign n18065 = ~n18059 & ~n40774;
  assign n18066 = ~n16728 & ~n18065;
  assign n18067 = n16704 & ~n16706;
  assign n18068 = ~n16707 & ~n18067;
  assign n18069 = ~n18066 & n18068;
  assign n18070 = ~n16707 & ~n18069;
  assign n18071 = n16683 & n40510;
  assign n18072 = ~n16689 & ~n18071;
  assign n18073 = ~n18070 & n18072;
  assign n18074 = ~n16689 & ~n18073;
  assign n18075 = ~n16652 & n16667;
  assign n18076 = n16652 & ~n16668;
  assign n18077 = n16652 & n16667;
  assign n18078 = ~n16667 & ~n16668;
  assign n18079 = ~n16652 & ~n16667;
  assign n18080 = ~n40775 & ~n40776;
  assign n18081 = ~n16668 & ~n18075;
  assign n18082 = ~n18074 & ~n40777;
  assign n18083 = ~n16668 & ~n18082;
  assign n18084 = n16642 & n40503;
  assign n18085 = ~n40503 & ~n16650;
  assign n18086 = ~n16642 & ~n16650;
  assign n18087 = ~n18085 & ~n18086;
  assign n18088 = ~n16650 & ~n18084;
  assign n18089 = ~n18083 & ~n40778;
  assign n18090 = ~n16650 & ~n18089;
  assign n18091 = ~n16611 & n16626;
  assign n18092 = n16611 & ~n16627;
  assign n18093 = n16611 & n16626;
  assign n18094 = ~n16626 & ~n16627;
  assign n18095 = ~n16611 & ~n16626;
  assign n18096 = ~n40779 & ~n40780;
  assign n18097 = ~n16627 & ~n18091;
  assign n18098 = ~n18090 & ~n40781;
  assign n18099 = ~n16627 & ~n18098;
  assign n18100 = n16603 & n40494;
  assign n18101 = ~n16603 & ~n16609;
  assign n18102 = ~n40494 & ~n16609;
  assign n18103 = ~n18101 & ~n18102;
  assign n18104 = ~n16609 & ~n18100;
  assign n18105 = ~n18099 & ~n40782;
  assign n18106 = ~n16609 & ~n18105;
  assign n18107 = ~n15140 & n40211;
  assign n18108 = ~n15188 & ~n18107;
  assign n18109 = ~n18106 & n18108;
  assign n18110 = ~n15188 & ~n18109;
  assign n18111 = n15138 & ~n18110;
  assign n18112 = ~n15136 & ~n18111;
  assign n18113 = ~n15045 & n40193;
  assign n18114 = ~n15089 & ~n18113;
  assign n18115 = ~n18112 & n18114;
  assign n18116 = ~n15089 & ~n18115;
  assign n18117 = ~n14996 & ~n15044;
  assign n18118 = ~n14929 & ~n14988;
  assign n18119 = ~n14930 & ~n14990;
  assign n18120 = ~n14930 & ~n18118;
  assign n18121 = n14944 & n15111;
  assign n18122 = pi122  & n40177;
  assign n18123 = pi124  & n14974;
  assign n18124 = pi123  & n14976;
  assign n18125 = ~n18123 & ~n18124;
  assign n18126 = ~n18122 & ~n18124;
  assign n18127 = ~n18123 & n18126;
  assign n18128 = ~n18122 & n18125;
  assign n18129 = ~n18121 & n40784;
  assign n18130 = pi5  & ~n18129;
  assign n18131 = pi5  & ~n18130;
  assign n18132 = pi5  & n18129;
  assign n18133 = ~n18129 & ~n18130;
  assign n18134 = ~pi5  & ~n18129;
  assign n18135 = ~n40785 & ~n40786;
  assign n18136 = ~n14901 & ~n14904;
  assign n18137 = ~n14887 & ~n14895;
  assign n18138 = n523 & n563;
  assign n18139 = pi113  & n37482;
  assign n18140 = pi115  & n578;
  assign n18141 = pi114  & n580;
  assign n18142 = ~n18140 & ~n18141;
  assign n18143 = ~n18139 & ~n18141;
  assign n18144 = ~n18140 & n18143;
  assign n18145 = ~n18139 & n18142;
  assign n18146 = ~n18138 & n40787;
  assign n18147 = pi14  & ~n18146;
  assign n18148 = pi14  & ~n18147;
  assign n18149 = pi14  & n18146;
  assign n18150 = ~n18146 & ~n18147;
  assign n18151 = ~pi14  & ~n18146;
  assign n18152 = ~n40788 & ~n40789;
  assign n18153 = ~n14866 & ~n14869;
  assign n18154 = n8175 & n10844;
  assign n18155 = pi110  & n38895;
  assign n18156 = pi112  & n8190;
  assign n18157 = pi111  & n8192;
  assign n18158 = ~n18156 & ~n18157;
  assign n18159 = ~n18155 & ~n18157;
  assign n18160 = ~n18156 & n18159;
  assign n18161 = ~n18155 & n18158;
  assign n18162 = ~n18154 & n40790;
  assign n18163 = pi17  & ~n18162;
  assign n18164 = pi17  & ~n18163;
  assign n18165 = pi17  & n18162;
  assign n18166 = ~n18162 & ~n18163;
  assign n18167 = ~pi17  & ~n18162;
  assign n18168 = ~n40791 & ~n40792;
  assign n18169 = ~n14852 & ~n14860;
  assign n18170 = n6785 & n9701;
  assign n18171 = pi107  & n38631;
  assign n18172 = pi109  & n6800;
  assign n18173 = pi108  & n6802;
  assign n18174 = ~n18172 & ~n18173;
  assign n18175 = ~n18171 & ~n18173;
  assign n18176 = ~n18172 & n18175;
  assign n18177 = ~n18171 & n18174;
  assign n18178 = ~n18170 & n40793;
  assign n18179 = pi20  & ~n18178;
  assign n18180 = pi20  & ~n18179;
  assign n18181 = pi20  & n18178;
  assign n18182 = ~n18178 & ~n18179;
  assign n18183 = ~pi20  & ~n18178;
  assign n18184 = ~n40794 & ~n40795;
  assign n18185 = n5576 & n8209;
  assign n18186 = pi104  & n38406;
  assign n18187 = pi106  & n5591;
  assign n18188 = pi105  & n5593;
  assign n18189 = ~n18187 & ~n18188;
  assign n18190 = ~n18186 & ~n18188;
  assign n18191 = ~n18187 & n18190;
  assign n18192 = ~n18186 & n18189;
  assign n18193 = ~n18185 & n40796;
  assign n18194 = pi23  & ~n18193;
  assign n18195 = pi23  & ~n18194;
  assign n18196 = pi23  & n18193;
  assign n18197 = ~n18193 & ~n18194;
  assign n18198 = ~pi23  & ~n18193;
  assign n18199 = ~n40797 & ~n40798;
  assign n18200 = ~n14814 & ~n14823;
  assign n18201 = ~n14788 & ~n14797;
  assign n18202 = n607 & n6474;
  assign n18203 = pi98  & n37489;
  assign n18204 = pi100  & n620;
  assign n18205 = pi99  & n622;
  assign n18206 = ~n18204 & ~n18205;
  assign n18207 = ~n18203 & ~n18205;
  assign n18208 = ~n18204 & n18207;
  assign n18209 = ~n18203 & n18206;
  assign n18210 = ~n18202 & n40799;
  assign n18211 = pi29  & ~n18210;
  assign n18212 = pi29  & ~n18211;
  assign n18213 = pi29  & n18210;
  assign n18214 = ~n18210 & ~n18211;
  assign n18215 = ~pi29  & ~n18210;
  assign n18216 = ~n40800 & ~n40801;
  assign n18217 = ~n14724 & ~n14733;
  assign n18218 = ~n14703 & ~n14707;
  assign n18219 = ~n14691 & ~n14697;
  assign n18220 = n940 & n2804;
  assign n18221 = pi83  & n37541;
  assign n18222 = pi85  & n953;
  assign n18223 = pi84  & n955;
  assign n18224 = ~n18222 & ~n18223;
  assign n18225 = ~n18221 & ~n18223;
  assign n18226 = ~n18222 & n18225;
  assign n18227 = ~n18221 & n18224;
  assign n18228 = ~n18220 & n40802;
  assign n18229 = pi44  & ~n18228;
  assign n18230 = pi44  & ~n18229;
  assign n18231 = pi44  & n18228;
  assign n18232 = ~n18228 & ~n18229;
  assign n18233 = ~pi44  & ~n18228;
  assign n18234 = ~n40803 & ~n40804;
  assign n18235 = ~n14675 & ~n14683;
  assign n18236 = ~n14664 & ~n14672;
  assign n18237 = ~n14644 & ~n14646;
  assign n18238 = n1465 & n1971;
  assign n18239 = pi74  & n37864;
  assign n18240 = pi76  & n1973;
  assign n18241 = pi75  & n1981;
  assign n18242 = ~n18240 & ~n18241;
  assign n18243 = ~n18239 & ~n18241;
  assign n18244 = ~n18240 & n18243;
  assign n18245 = ~n18239 & n18242;
  assign n18246 = ~n18238 & n40805;
  assign n18247 = pi53  & ~n18246;
  assign n18248 = pi53  & ~n18247;
  assign n18249 = pi53  & n18246;
  assign n18250 = ~n18246 & ~n18247;
  assign n18251 = ~pi53  & ~n18246;
  assign n18252 = ~n40806 & ~n40807;
  assign n18253 = ~n14638 & ~n14640;
  assign n18254 = n972 & n7882;
  assign n18255 = pi68  & n39128;
  assign n18256 = pi70  & n7884;
  assign n18257 = pi69  & n7892;
  assign n18258 = ~n18256 & ~n18257;
  assign n18259 = ~n18255 & ~n18257;
  assign n18260 = ~n18256 & n18259;
  assign n18261 = ~n18255 & n18258;
  assign n18262 = ~n18254 & n40808;
  assign n18263 = pi59  & ~n18262;
  assign n18264 = pi59  & ~n18263;
  assign n18265 = pi59  & n18262;
  assign n18266 = ~n18262 & ~n18263;
  assign n18267 = ~pi59  & ~n18262;
  assign n18268 = ~n40809 & ~n40810;
  assign n18269 = n847 & n12674;
  assign n18270 = pi65  & n40107;
  assign n18271 = pi67  & n12676;
  assign n18272 = pi66  & n12684;
  assign n18273 = ~n18271 & ~n18272;
  assign n18274 = ~n18270 & ~n18272;
  assign n18275 = ~n18271 & n18274;
  assign n18276 = ~n18270 & n18273;
  assign n18277 = ~n18269 & n40811;
  assign n18278 = pi62  & ~n18277;
  assign n18279 = pi62  & ~n18278;
  assign n18280 = pi62  & n18277;
  assign n18281 = ~n18277 & ~n18278;
  assign n18282 = ~pi62  & ~n18277;
  assign n18283 = ~n40812 & ~n40813;
  assign n18284 = ~pi62  & ~pi63 ;
  assign n18285 = pi62  & pi63 ;
  assign n18286 = pi62  & ~pi63 ;
  assign n18287 = ~pi62  & pi63 ;
  assign n18288 = ~n18286 & ~n18287;
  assign n18289 = ~n18284 & ~n18285;
  assign n18290 = pi64  & ~n40814;
  assign n18291 = n40111 & n18290;
  assign n18292 = ~n40111 & ~n18290;
  assign n18293 = n40111 & ~n18291;
  assign n18294 = n40111 & ~n18290;
  assign n18295 = n18290 & ~n18291;
  assign n18296 = ~n40111 & n18290;
  assign n18297 = ~n40815 & ~n40816;
  assign n18298 = ~n18291 & ~n18292;
  assign n18299 = ~n18283 & ~n40817;
  assign n18300 = n18283 & n40817;
  assign n18301 = ~n40817 & ~n18299;
  assign n18302 = ~n18283 & ~n18299;
  assign n18303 = ~n18301 & ~n18302;
  assign n18304 = ~n18299 & ~n18300;
  assign n18305 = n18268 & n40818;
  assign n18306 = ~n18268 & ~n40818;
  assign n18307 = ~n18305 & ~n18306;
  assign n18308 = ~n14633 & n18307;
  assign n18309 = n14633 & ~n18307;
  assign n18310 = ~n18308 & ~n18309;
  assign n18311 = n1238 & n4312;
  assign n18312 = pi71  & n38376;
  assign n18313 = pi73  & n4314;
  assign n18314 = pi72  & n4322;
  assign n18315 = ~n18313 & ~n18314;
  assign n18316 = ~n18312 & ~n18314;
  assign n18317 = ~n18313 & n18316;
  assign n18318 = ~n18312 & n18315;
  assign n18319 = ~n18311 & n40819;
  assign n18320 = pi56  & ~n18319;
  assign n18321 = pi56  & ~n18320;
  assign n18322 = pi56  & n18319;
  assign n18323 = ~n18319 & ~n18320;
  assign n18324 = ~pi56  & ~n18319;
  assign n18325 = ~n40820 & ~n40821;
  assign n18326 = n18310 & ~n18325;
  assign n18327 = ~n18310 & n18325;
  assign n18328 = n18310 & ~n18326;
  assign n18329 = n18310 & n18325;
  assign n18330 = ~n18325 & ~n18326;
  assign n18331 = ~n18310 & ~n18325;
  assign n18332 = ~n40822 & ~n40823;
  assign n18333 = ~n18326 & ~n18327;
  assign n18334 = ~n18253 & ~n40824;
  assign n18335 = n18253 & n40824;
  assign n18336 = ~n18253 & n40824;
  assign n18337 = n18253 & ~n40824;
  assign n18338 = ~n18336 & ~n18337;
  assign n18339 = ~n18334 & ~n18335;
  assign n18340 = n18252 & n40825;
  assign n18341 = ~n18252 & ~n40825;
  assign n18342 = ~n18340 & ~n18341;
  assign n18343 = ~n18237 & n18342;
  assign n18344 = n18237 & ~n18342;
  assign n18345 = ~n18343 & ~n18344;
  assign n18346 = n678 & n894;
  assign n18347 = pi77  & n37580;
  assign n18348 = pi79  & n896;
  assign n18349 = pi78  & n904;
  assign n18350 = ~n18348 & ~n18349;
  assign n18351 = ~n18347 & ~n18349;
  assign n18352 = ~n18348 & n18351;
  assign n18353 = ~n18347 & n18350;
  assign n18354 = ~n18346 & n40826;
  assign n18355 = pi50  & ~n18354;
  assign n18356 = pi50  & ~n18355;
  assign n18357 = pi50  & n18354;
  assign n18358 = ~n18354 & ~n18355;
  assign n18359 = ~pi50  & ~n18354;
  assign n18360 = ~n40827 & ~n40828;
  assign n18361 = n18345 & ~n18360;
  assign n18362 = ~n18345 & n18360;
  assign n18363 = n18345 & ~n18361;
  assign n18364 = n18345 & n18360;
  assign n18365 = ~n18360 & ~n18361;
  assign n18366 = ~n18345 & ~n18360;
  assign n18367 = ~n40829 & ~n40830;
  assign n18368 = ~n18361 & ~n18362;
  assign n18369 = n18236 & n40831;
  assign n18370 = ~n18236 & ~n40831;
  assign n18371 = ~n18369 & ~n18370;
  assign n18372 = n785 & n2134;
  assign n18373 = pi80  & n37520;
  assign n18374 = pi82  & n787;
  assign n18375 = pi81  & n795;
  assign n18376 = ~n18374 & ~n18375;
  assign n18377 = ~n18373 & ~n18375;
  assign n18378 = ~n18374 & n18377;
  assign n18379 = ~n18373 & n18376;
  assign n18380 = ~n18372 & n40832;
  assign n18381 = pi47  & ~n18380;
  assign n18382 = pi47  & ~n18381;
  assign n18383 = pi47  & n18380;
  assign n18384 = ~n18380 & ~n18381;
  assign n18385 = ~pi47  & ~n18380;
  assign n18386 = ~n40833 & ~n40834;
  assign n18387 = ~n18371 & n18386;
  assign n18388 = n18371 & ~n18386;
  assign n18389 = ~n18387 & ~n18388;
  assign n18390 = ~n18235 & n18389;
  assign n18391 = n18235 & ~n18389;
  assign n18392 = ~n18390 & ~n18391;
  assign n18393 = ~n18234 & n18392;
  assign n18394 = n18234 & ~n18392;
  assign n18395 = ~n18393 & ~n18394;
  assign n18396 = ~n18219 & n18395;
  assign n18397 = n18219 & ~n18395;
  assign n18398 = ~n18396 & ~n18397;
  assign n18399 = n733 & n3354;
  assign n18400 = pi86  & n37510;
  assign n18401 = pi88  & n746;
  assign n18402 = pi87  & n748;
  assign n18403 = ~n18401 & ~n18402;
  assign n18404 = ~n18400 & ~n18402;
  assign n18405 = ~n18401 & n18404;
  assign n18406 = ~n18400 & n18403;
  assign n18407 = ~n18399 & n40835;
  assign n18408 = pi41  & ~n18407;
  assign n18409 = pi41  & ~n18408;
  assign n18410 = pi41  & n18407;
  assign n18411 = ~n18407 & ~n18408;
  assign n18412 = ~pi41  & ~n18407;
  assign n18413 = ~n40836 & ~n40837;
  assign n18414 = n18398 & ~n18413;
  assign n18415 = ~n18398 & n18413;
  assign n18416 = n18398 & ~n18414;
  assign n18417 = n18398 & n18413;
  assign n18418 = ~n18413 & ~n18414;
  assign n18419 = ~n18398 & ~n18413;
  assign n18420 = ~n40838 & ~n40839;
  assign n18421 = ~n18414 & ~n18415;
  assign n18422 = n18218 & n40840;
  assign n18423 = ~n18218 & ~n40840;
  assign n18424 = ~n18422 & ~n18423;
  assign n18425 = n594 & n691;
  assign n18426 = pi89  & n37503;
  assign n18427 = pi91  & n704;
  assign n18428 = pi90  & n706;
  assign n18429 = ~n18427 & ~n18428;
  assign n18430 = ~n18426 & ~n18428;
  assign n18431 = ~n18427 & n18430;
  assign n18432 = ~n18426 & n18429;
  assign n18433 = ~n18425 & n40841;
  assign n18434 = pi38  & ~n18433;
  assign n18435 = pi38  & ~n18434;
  assign n18436 = pi38  & n18433;
  assign n18437 = ~n18433 & ~n18434;
  assign n18438 = ~pi38  & ~n18433;
  assign n18439 = ~n40842 & ~n40843;
  assign n18440 = n18424 & ~n18439;
  assign n18441 = ~n18424 & n18439;
  assign n18442 = n18424 & ~n18440;
  assign n18443 = n18424 & n18439;
  assign n18444 = ~n18439 & ~n18440;
  assign n18445 = ~n18424 & ~n18439;
  assign n18446 = ~n40844 & ~n40845;
  assign n18447 = ~n18440 & ~n18441;
  assign n18448 = n18217 & n40846;
  assign n18449 = ~n18217 & ~n40846;
  assign n18450 = ~n18448 & ~n18449;
  assign n18451 = n2104 & n4524;
  assign n18452 = pi92  & n37758;
  assign n18453 = pi94  & n2117;
  assign n18454 = pi93  & n2119;
  assign n18455 = ~n18453 & ~n18454;
  assign n18456 = ~n18452 & ~n18454;
  assign n18457 = ~n18453 & n18456;
  assign n18458 = ~n18452 & n18455;
  assign n18459 = ~n18451 & n40847;
  assign n18460 = pi35  & ~n18459;
  assign n18461 = pi35  & ~n18460;
  assign n18462 = pi35  & n18459;
  assign n18463 = ~n18459 & ~n18460;
  assign n18464 = ~pi35  & ~n18459;
  assign n18465 = ~n40848 & ~n40849;
  assign n18466 = ~n18450 & n18465;
  assign n18467 = n18450 & ~n18465;
  assign n18468 = ~n18466 & ~n18467;
  assign n18469 = ~n14750 & ~n14759;
  assign n18470 = n18468 & ~n18469;
  assign n18471 = ~n18468 & n18469;
  assign n18472 = ~n18470 & ~n18471;
  assign n18473 = n649 & n5630;
  assign n18474 = pi95  & n37496;
  assign n18475 = pi97  & n662;
  assign n18476 = pi96  & n664;
  assign n18477 = ~n18475 & ~n18476;
  assign n18478 = ~n18474 & ~n18476;
  assign n18479 = ~n18475 & n18478;
  assign n18480 = ~n18474 & n18477;
  assign n18481 = ~n18473 & n40850;
  assign n18482 = pi32  & ~n18481;
  assign n18483 = pi32  & ~n18482;
  assign n18484 = pi32  & n18481;
  assign n18485 = ~n18481 & ~n18482;
  assign n18486 = ~pi32  & ~n18481;
  assign n18487 = ~n40851 & ~n40852;
  assign n18488 = n18472 & ~n18487;
  assign n18489 = ~n18472 & n18487;
  assign n18490 = n18472 & ~n18488;
  assign n18491 = n18472 & n18487;
  assign n18492 = ~n18487 & ~n18488;
  assign n18493 = ~n18472 & ~n18487;
  assign n18494 = ~n40853 & ~n40854;
  assign n18495 = ~n18488 & ~n18489;
  assign n18496 = ~n14784 & ~n40855;
  assign n18497 = n14784 & n40855;
  assign n18498 = ~n14784 & n40855;
  assign n18499 = n14784 & ~n40855;
  assign n18500 = ~n18498 & ~n18499;
  assign n18501 = ~n18496 & ~n18497;
  assign n18502 = ~n18216 & ~n40856;
  assign n18503 = n18216 & n40856;
  assign n18504 = ~n18502 & ~n18503;
  assign n18505 = n18201 & ~n18504;
  assign n18506 = ~n18201 & n18504;
  assign n18507 = ~n18505 & ~n18506;
  assign n18508 = n4492 & n6787;
  assign n18509 = pi101  & n38208;
  assign n18510 = pi103  & n4507;
  assign n18511 = pi102  & n4509;
  assign n18512 = ~n18510 & ~n18511;
  assign n18513 = ~n18509 & ~n18511;
  assign n18514 = ~n18510 & n18513;
  assign n18515 = ~n18509 & n18512;
  assign n18516 = ~n18508 & n40857;
  assign n18517 = pi26  & ~n18516;
  assign n18518 = pi26  & ~n18517;
  assign n18519 = pi26  & n18516;
  assign n18520 = ~n18516 & ~n18517;
  assign n18521 = ~pi26  & ~n18516;
  assign n18522 = ~n40858 & ~n40859;
  assign n18523 = ~n18507 & n18522;
  assign n18524 = n18507 & ~n18522;
  assign n18525 = ~n18523 & ~n18524;
  assign n18526 = ~n18200 & n18525;
  assign n18527 = n18200 & ~n18525;
  assign n18528 = ~n18526 & ~n18527;
  assign n18529 = ~n18199 & n18528;
  assign n18530 = n18199 & ~n18528;
  assign n18531 = ~n18199 & ~n18529;
  assign n18532 = ~n18199 & ~n18528;
  assign n18533 = n18528 & ~n18529;
  assign n18534 = n18199 & n18528;
  assign n18535 = ~n40860 & ~n40861;
  assign n18536 = ~n18529 & ~n18530;
  assign n18537 = ~n14848 & ~n40862;
  assign n18538 = n14848 & ~n40861;
  assign n18539 = ~n40860 & n18538;
  assign n18540 = n14848 & n40862;
  assign n18541 = ~n18537 & ~n40863;
  assign n18542 = ~n18184 & n18541;
  assign n18543 = n18184 & ~n18541;
  assign n18544 = ~n18184 & ~n18542;
  assign n18545 = ~n18184 & ~n18541;
  assign n18546 = n18541 & ~n18542;
  assign n18547 = n18184 & n18541;
  assign n18548 = ~n40864 & ~n40865;
  assign n18549 = ~n18542 & ~n18543;
  assign n18550 = ~n18169 & ~n40866;
  assign n18551 = n18169 & ~n40865;
  assign n18552 = ~n40864 & n18551;
  assign n18553 = n18169 & n40866;
  assign n18554 = ~n18550 & ~n40867;
  assign n18555 = ~n18168 & n18554;
  assign n18556 = n18168 & ~n18554;
  assign n18557 = ~n18168 & ~n18555;
  assign n18558 = ~n18168 & ~n18554;
  assign n18559 = n18554 & ~n18555;
  assign n18560 = n18168 & n18554;
  assign n18561 = ~n40868 & ~n40869;
  assign n18562 = ~n18555 & ~n18556;
  assign n18563 = ~n18153 & ~n40870;
  assign n18564 = n18153 & ~n40869;
  assign n18565 = ~n40868 & n18564;
  assign n18566 = n18153 & n40870;
  assign n18567 = ~n18563 & ~n40871;
  assign n18568 = ~n18152 & n18567;
  assign n18569 = n18152 & ~n18567;
  assign n18570 = ~n18568 & ~n18569;
  assign n18571 = ~n18137 & n18570;
  assign n18572 = n18137 & ~n18570;
  assign n18573 = ~n18571 & ~n18572;
  assign n18574 = n269 & n13057;
  assign n18575 = pi116  & n37475;
  assign n18576 = pi118  & n536;
  assign n18577 = pi117  & n538;
  assign n18578 = ~n18576 & ~n18577;
  assign n18579 = ~n18575 & ~n18577;
  assign n18580 = ~n18576 & n18579;
  assign n18581 = ~n18575 & n18578;
  assign n18582 = ~n18574 & n40872;
  assign n18583 = pi11  & ~n18582;
  assign n18584 = pi11  & ~n18583;
  assign n18585 = pi11  & n18582;
  assign n18586 = ~n18582 & ~n18583;
  assign n18587 = ~pi11  & ~n18582;
  assign n18588 = ~n40873 & ~n40874;
  assign n18589 = n18573 & ~n18588;
  assign n18590 = ~n18573 & n18588;
  assign n18591 = n18573 & ~n18589;
  assign n18592 = n18573 & n18588;
  assign n18593 = ~n18588 & ~n18589;
  assign n18594 = ~n18573 & ~n18588;
  assign n18595 = ~n40875 & ~n40876;
  assign n18596 = ~n18589 & ~n18590;
  assign n18597 = n18136 & n40877;
  assign n18598 = ~n18136 & ~n40877;
  assign n18599 = ~n18597 & ~n18598;
  assign n18600 = n13010 & n15091;
  assign n18601 = pi119  & n39810;
  assign n18602 = pi121  & n13040;
  assign n18603 = pi120  & n13042;
  assign n18604 = ~n18602 & ~n18603;
  assign n18605 = ~n18601 & ~n18603;
  assign n18606 = ~n18602 & n18605;
  assign n18607 = ~n18601 & n18604;
  assign n18608 = ~n18600 & n40878;
  assign n18609 = pi8  & ~n18608;
  assign n18610 = pi8  & ~n18609;
  assign n18611 = pi8  & n18608;
  assign n18612 = ~n18608 & ~n18609;
  assign n18613 = ~pi8  & ~n18608;
  assign n18614 = ~n40879 & ~n40880;
  assign n18615 = n18599 & ~n18614;
  assign n18616 = ~n18599 & n18614;
  assign n18617 = n18599 & ~n18615;
  assign n18618 = n18599 & n18614;
  assign n18619 = ~n18614 & ~n18615;
  assign n18620 = ~n18599 & ~n18614;
  assign n18621 = ~n40881 & ~n40882;
  assign n18622 = ~n18615 & ~n18616;
  assign n18623 = ~n18135 & ~n40883;
  assign n18624 = n18135 & n40883;
  assign n18625 = n18135 & ~n40883;
  assign n18626 = ~n18135 & n40883;
  assign n18627 = ~n18625 & ~n18626;
  assign n18628 = ~n18623 & ~n18624;
  assign n18629 = n40783 & n40884;
  assign n18630 = ~n40783 & ~n40884;
  assign n18631 = ~n18629 & ~n18630;
  assign n18632 = ~n15017 & ~n15019;
  assign n18633 = pi126  & ~pi127 ;
  assign n18634 = ~pi126  & pi127 ;
  assign n18635 = ~n18633 & ~n18634;
  assign n18636 = n18632 & ~n18635;
  assign n18637 = ~n18632 & n18635;
  assign n18638 = ~n18632 & ~n18635;
  assign n18639 = n18632 & n18635;
  assign n18640 = ~n18638 & ~n18639;
  assign n18641 = ~n18636 & ~n18637;
  assign n18642 = n15004 & n40885;
  assign n18643 = pi127  & n15023;
  assign n18644 = pi125  & n40183;
  assign n18645 = pi126  & n15030;
  assign n18646 = ~n18644 & ~n18645;
  assign n18647 = ~n18643 & ~n18645;
  assign n18648 = ~n18644 & n18647;
  assign n18649 = ~n18643 & n18646;
  assign n18650 = ~n18642 & n40886;
  assign n18651 = pi2  & ~n18650;
  assign n18652 = pi2  & ~n18651;
  assign n18653 = pi2  & n18650;
  assign n18654 = ~n18650 & ~n18651;
  assign n18655 = ~pi2  & ~n18650;
  assign n18656 = ~n40887 & ~n40888;
  assign n18657 = n18631 & ~n18656;
  assign n18658 = ~n18631 & n18656;
  assign n18659 = n18631 & ~n18657;
  assign n18660 = ~n18656 & ~n18657;
  assign n18661 = ~n18659 & ~n18660;
  assign n18662 = ~n18657 & ~n18658;
  assign n18663 = ~n18117 & ~n40889;
  assign n18664 = n18117 & n40889;
  assign n18665 = ~n40889 & ~n18663;
  assign n18666 = ~n18117 & ~n18663;
  assign n18667 = ~n18665 & ~n18666;
  assign n18668 = ~n18663 & ~n18664;
  assign n18669 = ~n18116 & ~n40890;
  assign n18670 = n18116 & n40890;
  assign po63  = ~n18669 & ~n18670;
  assign n18672 = ~n18663 & ~n18669;
  assign n18673 = n18632 & ~n18634;
  assign n18674 = ~n18632 & ~n18633;
  assign n18675 = ~pi126  & n18632;
  assign n18676 = pi126  & ~n18632;
  assign n18677 = ~n18675 & ~n18676;
  assign n18678 = ~n18635 & ~n18677;
  assign n18679 = ~pi126  & ~n18638;
  assign n18680 = pi127  & ~n18679;
  assign n18681 = pi127  & ~n18680;
  assign n18682 = ~n18632 & n18633;
  assign n18683 = ~n18681 & ~n18682;
  assign n18684 = ~n18673 & ~n18674;
  assign n18685 = n15004 & n40891;
  assign n18686 = pi126  & n40183;
  assign n18687 = pi127  & n15030;
  assign n18688 = ~n18686 & ~n18687;
  assign n18689 = ~n18685 & n18688;
  assign n18690 = pi2  & ~n18689;
  assign n18691 = pi2  & ~n18690;
  assign n18692 = pi2  & n18689;
  assign n18693 = ~n18689 & ~n18690;
  assign n18694 = ~pi2  & ~n18689;
  assign n18695 = ~n40892 & ~n40893;
  assign n18696 = ~n18615 & ~n18623;
  assign n18697 = n14944 & n15068;
  assign n18698 = pi123  & n40177;
  assign n18699 = pi125  & n14974;
  assign n18700 = pi124  & n14976;
  assign n18701 = ~n18699 & ~n18700;
  assign n18702 = ~n18698 & ~n18700;
  assign n18703 = ~n18699 & n18702;
  assign n18704 = ~n18698 & n18701;
  assign n18705 = ~n18697 & n40894;
  assign n18706 = pi5  & ~n18705;
  assign n18707 = pi5  & ~n18706;
  assign n18708 = pi5  & n18705;
  assign n18709 = ~n18705 & ~n18706;
  assign n18710 = ~pi5  & ~n18705;
  assign n18711 = ~n40895 & ~n40896;
  assign n18712 = ~n18589 & ~n18598;
  assign n18713 = n269 & n13027;
  assign n18714 = pi117  & n37475;
  assign n18715 = pi119  & n536;
  assign n18716 = pi118  & n538;
  assign n18717 = ~n18715 & ~n18716;
  assign n18718 = ~n18714 & ~n18716;
  assign n18719 = ~n18715 & n18718;
  assign n18720 = ~n18714 & n18717;
  assign n18721 = ~n18713 & n40897;
  assign n18722 = pi11  & ~n18721;
  assign n18723 = pi11  & ~n18722;
  assign n18724 = pi11  & n18721;
  assign n18725 = ~n18721 & ~n18722;
  assign n18726 = ~pi11  & ~n18721;
  assign n18727 = ~n40898 & ~n40899;
  assign n18728 = ~n18568 & ~n18571;
  assign n18729 = n563 & n12530;
  assign n18730 = pi114  & n37482;
  assign n18731 = pi116  & n578;
  assign n18732 = pi115  & n580;
  assign n18733 = ~n18731 & ~n18732;
  assign n18734 = ~n18730 & ~n18732;
  assign n18735 = ~n18731 & n18734;
  assign n18736 = ~n18730 & n18733;
  assign n18737 = ~n18729 & n40900;
  assign n18738 = pi14  & ~n18737;
  assign n18739 = pi14  & ~n18738;
  assign n18740 = pi14  & n18737;
  assign n18741 = ~n18737 & ~n18738;
  assign n18742 = ~pi14  & ~n18737;
  assign n18743 = ~n40901 & ~n40902;
  assign n18744 = ~n18555 & ~n18563;
  assign n18745 = n8175 & n11276;
  assign n18746 = pi111  & n38895;
  assign n18747 = pi113  & n8190;
  assign n18748 = pi112  & n8192;
  assign n18749 = ~n18747 & ~n18748;
  assign n18750 = ~n18746 & ~n18748;
  assign n18751 = ~n18747 & n18750;
  assign n18752 = ~n18746 & n18749;
  assign n18753 = ~n18745 & n40903;
  assign n18754 = pi17  & ~n18753;
  assign n18755 = pi17  & ~n18754;
  assign n18756 = pi17  & n18753;
  assign n18757 = ~n18753 & ~n18754;
  assign n18758 = ~pi17  & ~n18753;
  assign n18759 = ~n40904 & ~n40905;
  assign n18760 = ~n18542 & ~n18550;
  assign n18761 = n6785 & n9678;
  assign n18762 = pi108  & n38631;
  assign n18763 = pi110  & n6800;
  assign n18764 = pi109  & n6802;
  assign n18765 = ~n18763 & ~n18764;
  assign n18766 = ~n18762 & ~n18764;
  assign n18767 = ~n18763 & n18766;
  assign n18768 = ~n18762 & n18765;
  assign n18769 = ~n18761 & n40906;
  assign n18770 = pi20  & ~n18769;
  assign n18771 = pi20  & ~n18770;
  assign n18772 = pi20  & n18769;
  assign n18773 = ~n18769 & ~n18770;
  assign n18774 = ~pi20  & ~n18769;
  assign n18775 = ~n40907 & ~n40908;
  assign n18776 = ~n18529 & ~n18537;
  assign n18777 = n5576 & n8177;
  assign n18778 = pi105  & n38406;
  assign n18779 = pi107  & n5591;
  assign n18780 = pi106  & n5593;
  assign n18781 = ~n18779 & ~n18780;
  assign n18782 = ~n18778 & ~n18780;
  assign n18783 = ~n18779 & n18782;
  assign n18784 = ~n18778 & n18781;
  assign n18785 = ~n18777 & n40909;
  assign n18786 = pi23  & ~n18785;
  assign n18787 = pi23  & ~n18786;
  assign n18788 = pi23  & n18785;
  assign n18789 = ~n18785 & ~n18786;
  assign n18790 = ~pi23  & ~n18785;
  assign n18791 = ~n40910 & ~n40911;
  assign n18792 = ~n18524 & ~n18526;
  assign n18793 = ~n18502 & ~n18506;
  assign n18794 = ~n18488 & ~n18496;
  assign n18795 = ~n18440 & ~n18449;
  assign n18796 = ~n18414 & ~n18423;
  assign n18797 = ~n18393 & ~n18396;
  assign n18798 = ~n18361 & ~n18370;
  assign n18799 = ~n18326 & ~n18334;
  assign n18800 = ~n18306 & ~n18308;
  assign n18801 = ~n18291 & ~n18299;
  assign n18802 = n871 & n12674;
  assign n18803 = pi66  & n40107;
  assign n18804 = pi68  & n12676;
  assign n18805 = pi67  & n12684;
  assign n18806 = ~n18804 & ~n18805;
  assign n18807 = ~n18803 & ~n18805;
  assign n18808 = ~n18804 & n18807;
  assign n18809 = ~n18803 & n18806;
  assign n18810 = ~n18802 & n40912;
  assign n18811 = pi62  & ~n18810;
  assign n18812 = pi62  & ~n18811;
  assign n18813 = pi62  & n18810;
  assign n18814 = ~n18810 & ~n18811;
  assign n18815 = ~pi62  & ~n18810;
  assign n18816 = ~n40913 & ~n40914;
  assign n18817 = pi65  & ~n40814;
  assign n18818 = pi64  & n18285;
  assign n18819 = ~n18817 & ~n18818;
  assign n18820 = ~n18816 & ~n18819;
  assign n18821 = n18816 & n18819;
  assign n18822 = ~n18819 & ~n18820;
  assign n18823 = n18816 & ~n18819;
  assign n18824 = ~n18816 & ~n18820;
  assign n18825 = ~n18816 & n18819;
  assign n18826 = ~n40915 & ~n40916;
  assign n18827 = ~n18820 & ~n18821;
  assign n18828 = n18801 & n40917;
  assign n18829 = ~n18801 & ~n40917;
  assign n18830 = ~n18828 & ~n18829;
  assign n18831 = n927 & n7882;
  assign n18832 = pi69  & n39128;
  assign n18833 = pi71  & n7884;
  assign n18834 = pi70  & n7892;
  assign n18835 = ~n18833 & ~n18834;
  assign n18836 = ~n18832 & ~n18834;
  assign n18837 = ~n18833 & n18836;
  assign n18838 = ~n18832 & n18835;
  assign n18839 = ~n18831 & n40918;
  assign n18840 = pi59  & ~n18839;
  assign n18841 = pi59  & ~n18840;
  assign n18842 = pi59  & n18839;
  assign n18843 = ~n18839 & ~n18840;
  assign n18844 = ~pi59  & ~n18839;
  assign n18845 = ~n40919 & ~n40920;
  assign n18846 = ~n18830 & n18845;
  assign n18847 = n18830 & ~n18845;
  assign n18848 = ~n18846 & ~n18847;
  assign n18849 = ~n18800 & n18848;
  assign n18850 = n18800 & ~n18848;
  assign n18851 = ~n18849 & ~n18850;
  assign n18852 = n1218 & n4312;
  assign n18853 = pi72  & n38376;
  assign n18854 = pi74  & n4314;
  assign n18855 = pi73  & n4322;
  assign n18856 = ~n18854 & ~n18855;
  assign n18857 = ~n18853 & ~n18855;
  assign n18858 = ~n18854 & n18857;
  assign n18859 = ~n18853 & n18856;
  assign n18860 = ~n18852 & n40921;
  assign n18861 = pi56  & ~n18860;
  assign n18862 = pi56  & ~n18861;
  assign n18863 = pi56  & n18860;
  assign n18864 = ~n18860 & ~n18861;
  assign n18865 = ~pi56  & ~n18860;
  assign n18866 = ~n40922 & ~n40923;
  assign n18867 = n18851 & ~n18866;
  assign n18868 = ~n18851 & n18866;
  assign n18869 = n18851 & ~n18867;
  assign n18870 = n18851 & n18866;
  assign n18871 = ~n18866 & ~n18867;
  assign n18872 = ~n18851 & ~n18866;
  assign n18873 = ~n40924 & ~n40925;
  assign n18874 = ~n18867 & ~n18868;
  assign n18875 = n18799 & n40926;
  assign n18876 = ~n18799 & ~n40926;
  assign n18877 = ~n18875 & ~n18876;
  assign n18878 = n1596 & n1971;
  assign n18879 = pi75  & n37864;
  assign n18880 = pi77  & n1973;
  assign n18881 = pi76  & n1981;
  assign n18882 = ~n18880 & ~n18881;
  assign n18883 = ~n18879 & ~n18881;
  assign n18884 = ~n18880 & n18883;
  assign n18885 = ~n18879 & n18882;
  assign n18886 = ~n18878 & n40927;
  assign n18887 = pi53  & ~n18886;
  assign n18888 = pi53  & ~n18887;
  assign n18889 = pi53  & n18886;
  assign n18890 = ~n18886 & ~n18887;
  assign n18891 = ~pi53  & ~n18886;
  assign n18892 = ~n40928 & ~n40929;
  assign n18893 = ~n18877 & n18892;
  assign n18894 = n18877 & ~n18892;
  assign n18895 = ~n18893 & ~n18894;
  assign n18896 = ~n18341 & ~n18343;
  assign n18897 = n18895 & ~n18896;
  assign n18898 = ~n18895 & n18896;
  assign n18899 = ~n18897 & ~n18898;
  assign n18900 = n894 & n2063;
  assign n18901 = pi78  & n37580;
  assign n18902 = pi80  & n896;
  assign n18903 = pi79  & n904;
  assign n18904 = ~n18902 & ~n18903;
  assign n18905 = ~n18901 & ~n18903;
  assign n18906 = ~n18902 & n18905;
  assign n18907 = ~n18901 & n18904;
  assign n18908 = ~n18900 & n40930;
  assign n18909 = pi50  & ~n18908;
  assign n18910 = pi50  & ~n18909;
  assign n18911 = pi50  & n18908;
  assign n18912 = ~n18908 & ~n18909;
  assign n18913 = ~pi50  & ~n18908;
  assign n18914 = ~n40931 & ~n40932;
  assign n18915 = n18899 & ~n18914;
  assign n18916 = ~n18899 & n18914;
  assign n18917 = n18899 & ~n18915;
  assign n18918 = n18899 & n18914;
  assign n18919 = ~n18914 & ~n18915;
  assign n18920 = ~n18899 & ~n18914;
  assign n18921 = ~n40933 & ~n40934;
  assign n18922 = ~n18915 & ~n18916;
  assign n18923 = n18798 & n40935;
  assign n18924 = ~n18798 & ~n40935;
  assign n18925 = ~n18923 & ~n18924;
  assign n18926 = n785 & n2091;
  assign n18927 = pi81  & n37520;
  assign n18928 = pi83  & n787;
  assign n18929 = pi82  & n795;
  assign n18930 = ~n18928 & ~n18929;
  assign n18931 = ~n18927 & ~n18929;
  assign n18932 = ~n18928 & n18931;
  assign n18933 = ~n18927 & n18930;
  assign n18934 = ~n18926 & n40936;
  assign n18935 = pi47  & ~n18934;
  assign n18936 = pi47  & ~n18935;
  assign n18937 = pi47  & n18934;
  assign n18938 = ~n18934 & ~n18935;
  assign n18939 = ~pi47  & ~n18934;
  assign n18940 = ~n40937 & ~n40938;
  assign n18941 = ~n18925 & n18940;
  assign n18942 = n18925 & ~n18940;
  assign n18943 = ~n18941 & ~n18942;
  assign n18944 = ~n18388 & ~n18390;
  assign n18945 = n18943 & ~n18944;
  assign n18946 = ~n18943 & n18944;
  assign n18947 = ~n18945 & ~n18946;
  assign n18948 = n940 & n2779;
  assign n18949 = pi84  & n37541;
  assign n18950 = pi86  & n953;
  assign n18951 = pi85  & n955;
  assign n18952 = ~n18950 & ~n18951;
  assign n18953 = ~n18949 & ~n18951;
  assign n18954 = ~n18950 & n18953;
  assign n18955 = ~n18949 & n18952;
  assign n18956 = ~n18948 & n40939;
  assign n18957 = pi44  & ~n18956;
  assign n18958 = pi44  & ~n18957;
  assign n18959 = pi44  & n18956;
  assign n18960 = ~n18956 & ~n18957;
  assign n18961 = ~pi44  & ~n18956;
  assign n18962 = ~n40940 & ~n40941;
  assign n18963 = n18947 & ~n18962;
  assign n18964 = ~n18947 & n18962;
  assign n18965 = n18947 & ~n18963;
  assign n18966 = n18947 & n18962;
  assign n18967 = ~n18962 & ~n18963;
  assign n18968 = ~n18947 & ~n18962;
  assign n18969 = ~n40942 & ~n40943;
  assign n18970 = ~n18963 & ~n18964;
  assign n18971 = n18797 & n40944;
  assign n18972 = ~n18797 & ~n40944;
  assign n18973 = ~n18971 & ~n18972;
  assign n18974 = n733 & n3591;
  assign n18975 = pi87  & n37510;
  assign n18976 = pi89  & n746;
  assign n18977 = pi88  & n748;
  assign n18978 = ~n18976 & ~n18977;
  assign n18979 = ~n18975 & ~n18977;
  assign n18980 = ~n18976 & n18979;
  assign n18981 = ~n18975 & n18978;
  assign n18982 = ~n18974 & n40945;
  assign n18983 = pi41  & ~n18982;
  assign n18984 = pi41  & ~n18983;
  assign n18985 = pi41  & n18982;
  assign n18986 = ~n18982 & ~n18983;
  assign n18987 = ~pi41  & ~n18982;
  assign n18988 = ~n40946 & ~n40947;
  assign n18989 = n18973 & ~n18988;
  assign n18990 = ~n18973 & n18988;
  assign n18991 = n18973 & ~n18989;
  assign n18992 = n18973 & n18988;
  assign n18993 = ~n18988 & ~n18989;
  assign n18994 = ~n18973 & ~n18988;
  assign n18995 = ~n40948 & ~n40949;
  assign n18996 = ~n18989 & ~n18990;
  assign n18997 = n18796 & n40950;
  assign n18998 = ~n18796 & ~n40950;
  assign n18999 = ~n18997 & ~n18998;
  assign n19000 = n691 & n4453;
  assign n19001 = pi90  & n37503;
  assign n19002 = pi92  & n704;
  assign n19003 = pi91  & n706;
  assign n19004 = ~n19002 & ~n19003;
  assign n19005 = ~n19001 & ~n19003;
  assign n19006 = ~n19002 & n19005;
  assign n19007 = ~n19001 & n19004;
  assign n19008 = ~n19000 & n40951;
  assign n19009 = pi38  & ~n19008;
  assign n19010 = pi38  & ~n19009;
  assign n19011 = pi38  & n19008;
  assign n19012 = ~n19008 & ~n19009;
  assign n19013 = ~pi38  & ~n19008;
  assign n19014 = ~n40952 & ~n40953;
  assign n19015 = n18999 & ~n19014;
  assign n19016 = ~n18999 & n19014;
  assign n19017 = n18999 & ~n19015;
  assign n19018 = n18999 & n19014;
  assign n19019 = ~n19014 & ~n19015;
  assign n19020 = ~n18999 & ~n19014;
  assign n19021 = ~n40954 & ~n40955;
  assign n19022 = ~n19015 & ~n19016;
  assign n19023 = n18795 & n40956;
  assign n19024 = ~n18795 & ~n40956;
  assign n19025 = ~n19023 & ~n19024;
  assign n19026 = n2104 & n4494;
  assign n19027 = pi93  & n37758;
  assign n19028 = pi95  & n2117;
  assign n19029 = pi94  & n2119;
  assign n19030 = ~n19028 & ~n19029;
  assign n19031 = ~n19027 & ~n19029;
  assign n19032 = ~n19028 & n19031;
  assign n19033 = ~n19027 & n19030;
  assign n19034 = ~n19026 & n40957;
  assign n19035 = pi35  & ~n19034;
  assign n19036 = pi35  & ~n19035;
  assign n19037 = pi35  & n19034;
  assign n19038 = ~n19034 & ~n19035;
  assign n19039 = ~pi35  & ~n19034;
  assign n19040 = ~n40958 & ~n40959;
  assign n19041 = ~n19025 & n19040;
  assign n19042 = n19025 & ~n19040;
  assign n19043 = ~n19041 & ~n19042;
  assign n19044 = ~n18467 & ~n18470;
  assign n19045 = n19043 & ~n19044;
  assign n19046 = ~n19043 & n19044;
  assign n19047 = ~n19045 & ~n19046;
  assign n19048 = n649 & n5610;
  assign n19049 = pi96  & n37496;
  assign n19050 = pi98  & n662;
  assign n19051 = pi97  & n664;
  assign n19052 = ~n19050 & ~n19051;
  assign n19053 = ~n19049 & ~n19051;
  assign n19054 = ~n19050 & n19053;
  assign n19055 = ~n19049 & n19052;
  assign n19056 = ~n19048 & n40960;
  assign n19057 = pi32  & ~n19056;
  assign n19058 = pi32  & ~n19057;
  assign n19059 = pi32  & n19056;
  assign n19060 = ~n19056 & ~n19057;
  assign n19061 = ~pi32  & ~n19056;
  assign n19062 = ~n40961 & ~n40962;
  assign n19063 = n19047 & ~n19062;
  assign n19064 = ~n19047 & n19062;
  assign n19065 = n19047 & ~n19063;
  assign n19066 = n19047 & n19062;
  assign n19067 = ~n19062 & ~n19063;
  assign n19068 = ~n19047 & ~n19062;
  assign n19069 = ~n40963 & ~n40964;
  assign n19070 = ~n19063 & ~n19064;
  assign n19071 = n18794 & n40965;
  assign n19072 = ~n18794 & ~n40965;
  assign n19073 = ~n19071 & ~n19072;
  assign n19074 = n607 & n6839;
  assign n19075 = pi99  & n37489;
  assign n19076 = pi101  & n620;
  assign n19077 = pi100  & n622;
  assign n19078 = ~n19076 & ~n19077;
  assign n19079 = ~n19075 & ~n19077;
  assign n19080 = ~n19076 & n19079;
  assign n19081 = ~n19075 & n19078;
  assign n19082 = ~n19074 & n40966;
  assign n19083 = pi29  & ~n19082;
  assign n19084 = pi29  & ~n19083;
  assign n19085 = pi29  & n19082;
  assign n19086 = ~n19082 & ~n19083;
  assign n19087 = ~pi29  & ~n19082;
  assign n19088 = ~n40967 & ~n40968;
  assign n19089 = n19073 & ~n19088;
  assign n19090 = ~n19073 & n19088;
  assign n19091 = n19073 & ~n19089;
  assign n19092 = n19073 & n19088;
  assign n19093 = ~n19088 & ~n19089;
  assign n19094 = ~n19073 & ~n19088;
  assign n19095 = ~n40969 & ~n40970;
  assign n19096 = ~n19089 & ~n19090;
  assign n19097 = n18793 & n40971;
  assign n19098 = ~n18793 & ~n40971;
  assign n19099 = ~n19097 & ~n19098;
  assign n19100 = n4492 & n8136;
  assign n19101 = pi102  & n38208;
  assign n19102 = pi104  & n4507;
  assign n19103 = pi103  & n4509;
  assign n19104 = ~n19102 & ~n19103;
  assign n19105 = ~n19101 & ~n19103;
  assign n19106 = ~n19102 & n19105;
  assign n19107 = ~n19101 & n19104;
  assign n19108 = ~n19100 & n40972;
  assign n19109 = pi26  & ~n19108;
  assign n19110 = pi26  & ~n19109;
  assign n19111 = pi26  & n19108;
  assign n19112 = ~n19108 & ~n19109;
  assign n19113 = ~pi26  & ~n19108;
  assign n19114 = ~n40973 & ~n40974;
  assign n19115 = n19099 & ~n19114;
  assign n19116 = ~n19099 & n19114;
  assign n19117 = n19099 & ~n19115;
  assign n19118 = n19099 & n19114;
  assign n19119 = ~n19114 & ~n19115;
  assign n19120 = ~n19099 & ~n19114;
  assign n19121 = ~n40975 & ~n40976;
  assign n19122 = ~n19115 & ~n19116;
  assign n19123 = ~n18792 & ~n40977;
  assign n19124 = n18792 & n40977;
  assign n19125 = ~n40977 & ~n19123;
  assign n19126 = n18792 & ~n40977;
  assign n19127 = ~n18792 & ~n19123;
  assign n19128 = ~n18792 & n40977;
  assign n19129 = ~n40978 & ~n40979;
  assign n19130 = ~n19123 & ~n19124;
  assign n19131 = ~n18791 & ~n40980;
  assign n19132 = n18791 & n40980;
  assign n19133 = n18791 & ~n40980;
  assign n19134 = ~n18791 & n40980;
  assign n19135 = ~n19133 & ~n19134;
  assign n19136 = ~n19131 & ~n19132;
  assign n19137 = ~n18776 & ~n40981;
  assign n19138 = n18776 & n40981;
  assign n19139 = ~n19137 & ~n19138;
  assign n19140 = ~n18775 & n19139;
  assign n19141 = n18775 & ~n19139;
  assign n19142 = ~n18775 & ~n19140;
  assign n19143 = ~n18775 & ~n19139;
  assign n19144 = n19139 & ~n19140;
  assign n19145 = n18775 & n19139;
  assign n19146 = ~n40982 & ~n40983;
  assign n19147 = ~n19140 & ~n19141;
  assign n19148 = ~n18760 & ~n40984;
  assign n19149 = n18760 & ~n40983;
  assign n19150 = ~n40982 & n19149;
  assign n19151 = n18760 & n40984;
  assign n19152 = ~n19148 & ~n40985;
  assign n19153 = ~n18759 & n19152;
  assign n19154 = n18759 & ~n19152;
  assign n19155 = ~n18759 & ~n19153;
  assign n19156 = ~n18759 & ~n19152;
  assign n19157 = n19152 & ~n19153;
  assign n19158 = n18759 & n19152;
  assign n19159 = ~n40986 & ~n40987;
  assign n19160 = ~n19153 & ~n19154;
  assign n19161 = ~n18744 & ~n40988;
  assign n19162 = n18744 & ~n40987;
  assign n19163 = ~n40986 & n19162;
  assign n19164 = n18744 & n40988;
  assign n19165 = ~n19161 & ~n40989;
  assign n19166 = ~n18743 & n19165;
  assign n19167 = n18743 & ~n19165;
  assign n19168 = ~n19166 & ~n19167;
  assign n19169 = ~n18728 & n19168;
  assign n19170 = n18728 & ~n19168;
  assign n19171 = ~n19169 & ~n19170;
  assign n19172 = ~n18727 & n19171;
  assign n19173 = n18727 & ~n19171;
  assign n19174 = ~n19172 & ~n19173;
  assign n19175 = ~n18712 & n19174;
  assign n19176 = n18712 & ~n19174;
  assign n19177 = ~n19175 & ~n19176;
  assign n19178 = n13010 & n15049;
  assign n19179 = pi120  & n39810;
  assign n19180 = pi122  & n13040;
  assign n19181 = pi121  & n13042;
  assign n19182 = ~n19180 & ~n19181;
  assign n19183 = ~n19179 & ~n19181;
  assign n19184 = ~n19180 & n19183;
  assign n19185 = ~n19179 & n19182;
  assign n19186 = ~n19178 & n40990;
  assign n19187 = pi8  & ~n19186;
  assign n19188 = pi8  & ~n19187;
  assign n19189 = pi8  & n19186;
  assign n19190 = ~n19186 & ~n19187;
  assign n19191 = ~pi8  & ~n19186;
  assign n19192 = ~n40991 & ~n40992;
  assign n19193 = n19177 & ~n19192;
  assign n19194 = ~n19177 & n19192;
  assign n19195 = n19177 & ~n19193;
  assign n19196 = n19177 & n19192;
  assign n19197 = ~n19192 & ~n19193;
  assign n19198 = ~n19177 & ~n19192;
  assign n19199 = ~n40993 & ~n40994;
  assign n19200 = ~n19193 & ~n19194;
  assign n19201 = ~n18711 & ~n40995;
  assign n19202 = n18711 & n40995;
  assign n19203 = n18711 & ~n40995;
  assign n19204 = ~n18711 & n40995;
  assign n19205 = ~n19203 & ~n19204;
  assign n19206 = ~n19201 & ~n19202;
  assign n19207 = ~n18696 & ~n40996;
  assign n19208 = n18696 & n40996;
  assign n19209 = ~n19207 & ~n19208;
  assign n19210 = ~n18695 & n19209;
  assign n19211 = n18695 & ~n19209;
  assign n19212 = ~n19210 & ~n19211;
  assign n19213 = ~n18630 & n18656;
  assign n19214 = ~n18630 & ~n18657;
  assign n19215 = ~n18629 & ~n19213;
  assign n19216 = n19212 & ~n40997;
  assign n19217 = ~n19212 & n40997;
  assign n19218 = ~n19216 & ~n19217;
  assign n19219 = ~n18672 & n19218;
  assign n19220 = n18672 & ~n19218;
  assign po64  = ~n19219 & ~n19220;
  assign n19222 = ~n19207 & ~n19210;
  assign n19223 = ~n19193 & ~n19201;
  assign n19224 = pi127  & n15004;
  assign n19225 = n15004 & n18680;
  assign n19226 = ~n18675 & n19224;
  assign n19227 = pi127  & n40183;
  assign n19228 = pi2  & ~n19227;
  assign n19229 = ~n40998 & ~n19228;
  assign n19230 = pi2  & n40998;
  assign n19231 = ~n40998 & ~n19227;
  assign n19232 = pi2  & ~n19231;
  assign n19233 = ~pi2  & ~n40998;
  assign n19234 = ~n19232 & ~n19233;
  assign n19235 = ~n40998 & n19228;
  assign n19236 = ~pi2  & n40998;
  assign n19237 = ~n19235 & ~n19236;
  assign n19238 = ~n19229 & ~n19230;
  assign n19239 = ~n19223 & n40999;
  assign n19240 = n19223 & ~n40999;
  assign n19241 = ~n19239 & ~n19240;
  assign n19242 = ~n19172 & ~n19175;
  assign n19243 = ~n19166 & ~n19169;
  assign n19244 = ~n19153 & ~n19161;
  assign n19245 = n8175 & n11258;
  assign n19246 = pi112  & n38895;
  assign n19247 = pi114  & n8190;
  assign n19248 = pi113  & n8192;
  assign n19249 = ~n19247 & ~n19248;
  assign n19250 = ~n19246 & ~n19248;
  assign n19251 = ~n19247 & n19250;
  assign n19252 = ~n19246 & n19249;
  assign n19253 = ~n19245 & n41000;
  assign n19254 = pi17  & ~n19253;
  assign n19255 = pi17  & ~n19254;
  assign n19256 = pi17  & n19253;
  assign n19257 = ~n19253 & ~n19254;
  assign n19258 = ~pi17  & ~n19253;
  assign n19259 = ~n41001 & ~n41002;
  assign n19260 = ~n19140 & ~n19148;
  assign n19261 = n565 & n6785;
  assign n19262 = pi109  & n38631;
  assign n19263 = pi111  & n6800;
  assign n19264 = pi110  & n6802;
  assign n19265 = ~n19263 & ~n19264;
  assign n19266 = ~n19262 & ~n19264;
  assign n19267 = ~n19263 & n19266;
  assign n19268 = ~n19262 & n19265;
  assign n19269 = ~n19261 & n41003;
  assign n19270 = pi20  & ~n19269;
  assign n19271 = pi20  & ~n19270;
  assign n19272 = pi20  & n19269;
  assign n19273 = ~n19269 & ~n19270;
  assign n19274 = ~pi20  & ~n19269;
  assign n19275 = ~n41004 & ~n41005;
  assign n19276 = ~n19131 & ~n19137;
  assign n19277 = n5576 & n9277;
  assign n19278 = pi106  & n38406;
  assign n19279 = pi108  & n5591;
  assign n19280 = pi107  & n5593;
  assign n19281 = ~n19279 & ~n19280;
  assign n19282 = ~n19278 & ~n19280;
  assign n19283 = ~n19279 & n19282;
  assign n19284 = ~n19278 & n19281;
  assign n19285 = ~n19277 & n41006;
  assign n19286 = pi23  & ~n19285;
  assign n19287 = pi23  & ~n19286;
  assign n19288 = pi23  & n19285;
  assign n19289 = ~n19285 & ~n19286;
  assign n19290 = ~pi23  & ~n19285;
  assign n19291 = ~n41007 & ~n41008;
  assign n19292 = ~n19115 & ~n19123;
  assign n19293 = ~n19089 & ~n19098;
  assign n19294 = ~n19063 & ~n19072;
  assign n19295 = n649 & n5578;
  assign n19296 = pi97  & n37496;
  assign n19297 = pi99  & n662;
  assign n19298 = pi98  & n664;
  assign n19299 = ~n19297 & ~n19298;
  assign n19300 = ~n19296 & ~n19298;
  assign n19301 = ~n19297 & n19300;
  assign n19302 = ~n19296 & n19299;
  assign n19303 = ~n19295 & n41009;
  assign n19304 = pi32  & ~n19303;
  assign n19305 = pi32  & ~n19304;
  assign n19306 = pi32  & n19303;
  assign n19307 = ~n19303 & ~n19304;
  assign n19308 = ~pi32  & ~n19303;
  assign n19309 = ~n41010 & ~n41011;
  assign n19310 = ~n19042 & ~n19045;
  assign n19311 = ~n19015 & ~n19024;
  assign n19312 = ~n18989 & ~n18998;
  assign n19313 = ~n18963 & ~n18972;
  assign n19314 = n636 & n940;
  assign n19315 = pi85  & n37541;
  assign n19316 = pi87  & n953;
  assign n19317 = pi86  & n955;
  assign n19318 = ~n19316 & ~n19317;
  assign n19319 = ~n19315 & ~n19317;
  assign n19320 = ~n19316 & n19319;
  assign n19321 = ~n19315 & n19318;
  assign n19322 = ~n19314 & n41012;
  assign n19323 = pi44  & ~n19322;
  assign n19324 = pi44  & ~n19323;
  assign n19325 = pi44  & n19322;
  assign n19326 = ~n19322 & ~n19323;
  assign n19327 = ~pi44  & ~n19322;
  assign n19328 = ~n41013 & ~n41014;
  assign n19329 = ~n18942 & ~n18945;
  assign n19330 = ~n18915 & ~n18924;
  assign n19331 = n894 & n2154;
  assign n19332 = pi79  & n37580;
  assign n19333 = pi81  & n896;
  assign n19334 = pi80  & n904;
  assign n19335 = ~n19333 & ~n19334;
  assign n19336 = ~n19332 & ~n19334;
  assign n19337 = ~n19333 & n19336;
  assign n19338 = ~n19332 & n19335;
  assign n19339 = ~n19331 & n41015;
  assign n19340 = pi50  & ~n19339;
  assign n19341 = pi50  & ~n19340;
  assign n19342 = pi50  & n19339;
  assign n19343 = ~n19339 & ~n19340;
  assign n19344 = ~pi50  & ~n19339;
  assign n19345 = ~n41016 & ~n41017;
  assign n19346 = ~n18894 & ~n18897;
  assign n19347 = ~n18867 & ~n18876;
  assign n19348 = n720 & n4312;
  assign n19349 = pi73  & n38376;
  assign n19350 = pi75  & n4314;
  assign n19351 = pi74  & n4322;
  assign n19352 = ~n19350 & ~n19351;
  assign n19353 = ~n19349 & ~n19351;
  assign n19354 = ~n19350 & n19353;
  assign n19355 = ~n19349 & n19352;
  assign n19356 = ~n19348 & n41018;
  assign n19357 = pi56  & ~n19356;
  assign n19358 = pi56  & ~n19357;
  assign n19359 = pi56  & n19356;
  assign n19360 = ~n19356 & ~n19357;
  assign n19361 = ~pi56  & ~n19356;
  assign n19362 = ~n41019 & ~n41020;
  assign n19363 = ~n18847 & ~n18849;
  assign n19364 = ~n18820 & ~n18829;
  assign n19365 = n990 & n12674;
  assign n19366 = pi67  & n40107;
  assign n19367 = pi69  & n12676;
  assign n19368 = pi68  & n12684;
  assign n19369 = ~n19367 & ~n19368;
  assign n19370 = ~n19366 & ~n19368;
  assign n19371 = ~n19367 & n19370;
  assign n19372 = ~n19366 & n19369;
  assign n19373 = ~n19365 & n41021;
  assign n19374 = pi62  & ~n19373;
  assign n19375 = pi62  & ~n19374;
  assign n19376 = pi62  & n19373;
  assign n19377 = ~n19373 & ~n19374;
  assign n19378 = ~pi62  & ~n19373;
  assign n19379 = ~n41022 & ~n41023;
  assign n19380 = pi66  & ~n40814;
  assign n19381 = pi65  & n18285;
  assign n19382 = ~n19380 & ~n19381;
  assign n19383 = ~n19379 & ~n19382;
  assign n19384 = n19379 & n19382;
  assign n19385 = ~n19382 & ~n19383;
  assign n19386 = n19379 & ~n19382;
  assign n19387 = ~n19379 & ~n19383;
  assign n19388 = ~n19379 & n19382;
  assign n19389 = ~n41024 & ~n41025;
  assign n19390 = ~n19383 & ~n19384;
  assign n19391 = n19364 & n41026;
  assign n19392 = ~n19364 & ~n41026;
  assign n19393 = ~n19391 & ~n19392;
  assign n19394 = n1124 & n7882;
  assign n19395 = pi70  & n39128;
  assign n19396 = pi72  & n7884;
  assign n19397 = pi71  & n7892;
  assign n19398 = ~n19396 & ~n19397;
  assign n19399 = ~n19395 & ~n19397;
  assign n19400 = ~n19396 & n19399;
  assign n19401 = ~n19395 & n19398;
  assign n19402 = ~n19394 & n41027;
  assign n19403 = pi59  & ~n19402;
  assign n19404 = pi59  & ~n19403;
  assign n19405 = pi59  & n19402;
  assign n19406 = ~n19402 & ~n19403;
  assign n19407 = ~pi59  & ~n19402;
  assign n19408 = ~n41028 & ~n41029;
  assign n19409 = n19393 & ~n19408;
  assign n19410 = ~n19393 & n19408;
  assign n19411 = ~n19409 & ~n19410;
  assign n19412 = ~n19363 & ~n19410;
  assign n19413 = ~n19409 & n19412;
  assign n19414 = ~n19363 & n19411;
  assign n19415 = n19363 & ~n19411;
  assign n19416 = ~n19363 & ~n41030;
  assign n19417 = ~n19409 & ~n41030;
  assign n19418 = ~n19410 & n19417;
  assign n19419 = ~n19416 & ~n19418;
  assign n19420 = ~n41030 & ~n19415;
  assign n19421 = n19362 & n41031;
  assign n19422 = ~n19362 & ~n41031;
  assign n19423 = ~n19421 & ~n19422;
  assign n19424 = ~n19347 & n19423;
  assign n19425 = n19347 & ~n19423;
  assign n19426 = ~n19424 & ~n19425;
  assign n19427 = n1578 & n1971;
  assign n19428 = pi76  & n37864;
  assign n19429 = pi78  & n1973;
  assign n19430 = pi77  & n1981;
  assign n19431 = ~n19429 & ~n19430;
  assign n19432 = ~n19428 & ~n19430;
  assign n19433 = ~n19429 & n19432;
  assign n19434 = ~n19428 & n19431;
  assign n19435 = ~n19427 & n41032;
  assign n19436 = pi53  & ~n19435;
  assign n19437 = pi53  & ~n19436;
  assign n19438 = pi53  & n19435;
  assign n19439 = ~n19435 & ~n19436;
  assign n19440 = ~pi53  & ~n19435;
  assign n19441 = ~n41033 & ~n41034;
  assign n19442 = n19426 & ~n19441;
  assign n19443 = ~n19426 & n19441;
  assign n19444 = n19426 & ~n19442;
  assign n19445 = n19426 & n19441;
  assign n19446 = ~n19441 & ~n19442;
  assign n19447 = ~n19426 & ~n19441;
  assign n19448 = ~n41035 & ~n41036;
  assign n19449 = ~n19442 & ~n19443;
  assign n19450 = ~n19346 & ~n41037;
  assign n19451 = n19346 & n41037;
  assign n19452 = ~n19346 & n41037;
  assign n19453 = n19346 & ~n41037;
  assign n19454 = ~n19452 & ~n19453;
  assign n19455 = ~n19450 & ~n19451;
  assign n19456 = ~n19345 & ~n41038;
  assign n19457 = n19345 & n41038;
  assign n19458 = ~n19456 & ~n19457;
  assign n19459 = n19330 & ~n19458;
  assign n19460 = ~n19330 & n19458;
  assign n19461 = ~n19459 & ~n19460;
  assign n19462 = n785 & n2591;
  assign n19463 = pi82  & n37520;
  assign n19464 = pi84  & n787;
  assign n19465 = pi83  & n795;
  assign n19466 = ~n19464 & ~n19465;
  assign n19467 = ~n19463 & ~n19465;
  assign n19468 = ~n19464 & n19467;
  assign n19469 = ~n19463 & n19466;
  assign n19470 = ~n19462 & n41039;
  assign n19471 = pi47  & ~n19470;
  assign n19472 = pi47  & ~n19471;
  assign n19473 = pi47  & n19470;
  assign n19474 = ~n19470 & ~n19471;
  assign n19475 = ~pi47  & ~n19470;
  assign n19476 = ~n41040 & ~n41041;
  assign n19477 = n19461 & ~n19476;
  assign n19478 = ~n19461 & n19476;
  assign n19479 = n19461 & ~n19477;
  assign n19480 = n19461 & n19476;
  assign n19481 = ~n19476 & ~n19477;
  assign n19482 = ~n19461 & ~n19476;
  assign n19483 = ~n41042 & ~n41043;
  assign n19484 = ~n19477 & ~n19478;
  assign n19485 = ~n19329 & ~n41044;
  assign n19486 = n19329 & n41044;
  assign n19487 = ~n19329 & n41044;
  assign n19488 = n19329 & ~n41044;
  assign n19489 = ~n19487 & ~n19488;
  assign n19490 = ~n19485 & ~n19486;
  assign n19491 = ~n19328 & ~n41045;
  assign n19492 = n19328 & n41045;
  assign n19493 = ~n19491 & ~n19492;
  assign n19494 = n19313 & ~n19493;
  assign n19495 = ~n19313 & n19493;
  assign n19496 = ~n19494 & ~n19495;
  assign n19497 = n733 & n3566;
  assign n19498 = pi88  & n37510;
  assign n19499 = pi90  & n746;
  assign n19500 = pi89  & n748;
  assign n19501 = ~n19499 & ~n19500;
  assign n19502 = ~n19498 & ~n19500;
  assign n19503 = ~n19499 & n19502;
  assign n19504 = ~n19498 & n19501;
  assign n19505 = ~n19497 & n41046;
  assign n19506 = pi41  & ~n19505;
  assign n19507 = pi41  & ~n19506;
  assign n19508 = pi41  & n19505;
  assign n19509 = ~n19505 & ~n19506;
  assign n19510 = ~pi41  & ~n19505;
  assign n19511 = ~n41047 & ~n41048;
  assign n19512 = n19496 & ~n19511;
  assign n19513 = ~n19496 & n19511;
  assign n19514 = n19496 & ~n19512;
  assign n19515 = n19496 & n19511;
  assign n19516 = ~n19511 & ~n19512;
  assign n19517 = ~n19496 & ~n19511;
  assign n19518 = ~n41049 & ~n41050;
  assign n19519 = ~n19512 & ~n19513;
  assign n19520 = n19312 & n41051;
  assign n19521 = ~n19312 & ~n41051;
  assign n19522 = ~n19520 & ~n19521;
  assign n19523 = n691 & n4544;
  assign n19524 = pi91  & n37503;
  assign n19525 = pi93  & n704;
  assign n19526 = pi92  & n706;
  assign n19527 = ~n19525 & ~n19526;
  assign n19528 = ~n19524 & ~n19526;
  assign n19529 = ~n19525 & n19528;
  assign n19530 = ~n19524 & n19527;
  assign n19531 = ~n19523 & n41052;
  assign n19532 = pi38  & ~n19531;
  assign n19533 = pi38  & ~n19532;
  assign n19534 = pi38  & n19531;
  assign n19535 = ~n19531 & ~n19532;
  assign n19536 = ~pi38  & ~n19531;
  assign n19537 = ~n41053 & ~n41054;
  assign n19538 = n19522 & ~n19537;
  assign n19539 = ~n19522 & n19537;
  assign n19540 = n19522 & ~n19538;
  assign n19541 = n19522 & n19537;
  assign n19542 = ~n19537 & ~n19538;
  assign n19543 = ~n19522 & ~n19537;
  assign n19544 = ~n41055 & ~n41056;
  assign n19545 = ~n19538 & ~n19539;
  assign n19546 = n19311 & n41057;
  assign n19547 = ~n19311 & ~n41057;
  assign n19548 = ~n19546 & ~n19547;
  assign n19549 = n2104 & n5281;
  assign n19550 = pi94  & n37758;
  assign n19551 = pi96  & n2117;
  assign n19552 = pi95  & n2119;
  assign n19553 = ~n19551 & ~n19552;
  assign n19554 = ~n19550 & ~n19552;
  assign n19555 = ~n19551 & n19554;
  assign n19556 = ~n19550 & n19553;
  assign n19557 = ~n19549 & n41058;
  assign n19558 = pi35  & ~n19557;
  assign n19559 = pi35  & ~n19558;
  assign n19560 = pi35  & n19557;
  assign n19561 = ~n19557 & ~n19558;
  assign n19562 = ~pi35  & ~n19557;
  assign n19563 = ~n41059 & ~n41060;
  assign n19564 = n19548 & ~n19563;
  assign n19565 = ~n19548 & n19563;
  assign n19566 = ~n19564 & ~n19565;
  assign n19567 = ~n19310 & ~n19565;
  assign n19568 = ~n19564 & n19567;
  assign n19569 = ~n19310 & n19566;
  assign n19570 = n19310 & ~n19566;
  assign n19571 = ~n19310 & ~n41061;
  assign n19572 = ~n19564 & ~n41061;
  assign n19573 = ~n19565 & n19572;
  assign n19574 = ~n19571 & ~n19573;
  assign n19575 = ~n41061 & ~n19570;
  assign n19576 = ~n19309 & ~n41062;
  assign n19577 = n19309 & n41062;
  assign n19578 = ~n41062 & ~n19576;
  assign n19579 = n19309 & ~n41062;
  assign n19580 = ~n19309 & ~n19576;
  assign n19581 = ~n19309 & n41062;
  assign n19582 = ~n41063 & ~n41064;
  assign n19583 = ~n19576 & ~n19577;
  assign n19584 = n19294 & n41065;
  assign n19585 = ~n19294 & ~n41065;
  assign n19586 = ~n19584 & ~n19585;
  assign n19587 = n607 & n6819;
  assign n19588 = pi100  & n37489;
  assign n19589 = pi102  & n620;
  assign n19590 = pi101  & n622;
  assign n19591 = ~n19589 & ~n19590;
  assign n19592 = ~n19588 & ~n19590;
  assign n19593 = ~n19589 & n19592;
  assign n19594 = ~n19588 & n19591;
  assign n19595 = ~n19587 & n41066;
  assign n19596 = pi29  & ~n19595;
  assign n19597 = pi29  & ~n19596;
  assign n19598 = pi29  & n19595;
  assign n19599 = ~n19595 & ~n19596;
  assign n19600 = ~pi29  & ~n19595;
  assign n19601 = ~n41067 & ~n41068;
  assign n19602 = n19586 & ~n19601;
  assign n19603 = ~n19586 & n19601;
  assign n19604 = n19586 & ~n19602;
  assign n19605 = n19586 & n19601;
  assign n19606 = ~n19601 & ~n19602;
  assign n19607 = ~n19586 & ~n19601;
  assign n19608 = ~n41069 & ~n41070;
  assign n19609 = ~n19602 & ~n19603;
  assign n19610 = n19293 & n41071;
  assign n19611 = ~n19293 & ~n41071;
  assign n19612 = ~n19610 & ~n19611;
  assign n19613 = n4492 & n8229;
  assign n19614 = pi103  & n38208;
  assign n19615 = pi105  & n4507;
  assign n19616 = pi104  & n4509;
  assign n19617 = ~n19615 & ~n19616;
  assign n19618 = ~n19614 & ~n19616;
  assign n19619 = ~n19615 & n19618;
  assign n19620 = ~n19614 & n19617;
  assign n19621 = ~n19613 & n41072;
  assign n19622 = pi26  & ~n19621;
  assign n19623 = pi26  & ~n19622;
  assign n19624 = pi26  & n19621;
  assign n19625 = ~n19621 & ~n19622;
  assign n19626 = ~pi26  & ~n19621;
  assign n19627 = ~n41073 & ~n41074;
  assign n19628 = n19612 & ~n19627;
  assign n19629 = ~n19612 & n19627;
  assign n19630 = ~n19628 & ~n19629;
  assign n19631 = ~n19292 & ~n19629;
  assign n19632 = ~n19628 & n19631;
  assign n19633 = ~n19292 & n19630;
  assign n19634 = n19292 & ~n19630;
  assign n19635 = ~n19292 & ~n41075;
  assign n19636 = ~n19628 & ~n41075;
  assign n19637 = ~n19629 & n19636;
  assign n19638 = ~n19635 & ~n19637;
  assign n19639 = ~n41075 & ~n19634;
  assign n19640 = ~n19291 & ~n41076;
  assign n19641 = n19291 & n41076;
  assign n19642 = ~n41076 & ~n19640;
  assign n19643 = n19291 & ~n41076;
  assign n19644 = ~n19291 & ~n19640;
  assign n19645 = ~n19291 & n41076;
  assign n19646 = ~n41077 & ~n41078;
  assign n19647 = ~n19640 & ~n19641;
  assign n19648 = ~n19276 & ~n41079;
  assign n19649 = n19276 & n41079;
  assign n19650 = ~n19648 & ~n19649;
  assign n19651 = ~n19275 & n19650;
  assign n19652 = n19275 & ~n19650;
  assign n19653 = ~n19275 & ~n19651;
  assign n19654 = ~n19275 & ~n19650;
  assign n19655 = n19650 & ~n19651;
  assign n19656 = n19275 & n19650;
  assign n19657 = ~n41080 & ~n41081;
  assign n19658 = ~n19651 & ~n19652;
  assign n19659 = ~n19260 & ~n41082;
  assign n19660 = n19260 & n41082;
  assign n19661 = ~n19260 & ~n19659;
  assign n19662 = ~n19260 & n41082;
  assign n19663 = ~n41082 & ~n19659;
  assign n19664 = n19260 & ~n41082;
  assign n19665 = ~n41083 & ~n41084;
  assign n19666 = ~n19659 & ~n19660;
  assign n19667 = n19259 & n41085;
  assign n19668 = ~n19259 & ~n41085;
  assign n19669 = ~n19667 & ~n19668;
  assign n19670 = ~n19244 & n19669;
  assign n19671 = n19244 & ~n19669;
  assign n19672 = ~n19670 & ~n19671;
  assign n19673 = n563 & n13079;
  assign n19674 = pi115  & n37482;
  assign n19675 = pi117  & n578;
  assign n19676 = pi116  & n580;
  assign n19677 = ~n19675 & ~n19676;
  assign n19678 = ~n19674 & ~n19676;
  assign n19679 = ~n19675 & n19678;
  assign n19680 = ~n19674 & n19677;
  assign n19681 = ~n19673 & n41086;
  assign n19682 = pi14  & ~n19681;
  assign n19683 = pi14  & ~n19682;
  assign n19684 = pi14  & n19681;
  assign n19685 = ~n19681 & ~n19682;
  assign n19686 = ~pi14  & ~n19681;
  assign n19687 = ~n41087 & ~n41088;
  assign n19688 = n19672 & ~n19687;
  assign n19689 = ~n19672 & n19687;
  assign n19690 = n19672 & ~n19688;
  assign n19691 = n19672 & n19687;
  assign n19692 = ~n19687 & ~n19688;
  assign n19693 = ~n19672 & ~n19687;
  assign n19694 = ~n41089 & ~n41090;
  assign n19695 = ~n19688 & ~n19689;
  assign n19696 = n19243 & n41091;
  assign n19697 = ~n19243 & ~n41091;
  assign n19698 = ~n19696 & ~n19697;
  assign n19699 = n269 & n14913;
  assign n19700 = pi118  & n37475;
  assign n19701 = pi120  & n536;
  assign n19702 = pi119  & n538;
  assign n19703 = ~n19701 & ~n19702;
  assign n19704 = ~n19700 & ~n19702;
  assign n19705 = ~n19701 & n19704;
  assign n19706 = ~n19700 & n19703;
  assign n19707 = ~n19699 & n41092;
  assign n19708 = pi11  & ~n19707;
  assign n19709 = pi11  & ~n19708;
  assign n19710 = pi11  & n19707;
  assign n19711 = ~n19707 & ~n19708;
  assign n19712 = ~pi11  & ~n19707;
  assign n19713 = ~n41093 & ~n41094;
  assign n19714 = ~n19698 & n19713;
  assign n19715 = n19698 & ~n19713;
  assign n19716 = ~n19714 & ~n19715;
  assign n19717 = n13010 & n14961;
  assign n19718 = pi121  & n39810;
  assign n19719 = pi123  & n13040;
  assign n19720 = pi122  & n13042;
  assign n19721 = ~n19719 & ~n19720;
  assign n19722 = ~n19718 & ~n19720;
  assign n19723 = ~n19719 & n19722;
  assign n19724 = ~n19718 & n19721;
  assign n19725 = ~n19717 & n41095;
  assign n19726 = pi8  & ~n19725;
  assign n19727 = pi8  & ~n19726;
  assign n19728 = pi8  & n19725;
  assign n19729 = ~n19725 & ~n19726;
  assign n19730 = ~pi8  & ~n19725;
  assign n19731 = ~n41096 & ~n41097;
  assign n19732 = ~n19716 & n19731;
  assign n19733 = n19716 & ~n19731;
  assign n19734 = n19716 & ~n19733;
  assign n19735 = ~n19731 & ~n19733;
  assign n19736 = ~n19734 & ~n19735;
  assign n19737 = ~n19732 & ~n19733;
  assign n19738 = n19242 & n41098;
  assign n19739 = ~n19242 & ~n41098;
  assign n19740 = ~n19738 & ~n19739;
  assign n19741 = n14944 & n15021;
  assign n19742 = pi124  & n40177;
  assign n19743 = pi126  & n14974;
  assign n19744 = pi125  & n14976;
  assign n19745 = ~n19743 & ~n19744;
  assign n19746 = ~n19742 & ~n19744;
  assign n19747 = ~n19743 & n19746;
  assign n19748 = ~n19742 & n19745;
  assign n19749 = ~n19741 & n41099;
  assign n19750 = pi5  & ~n19749;
  assign n19751 = pi5  & ~n19750;
  assign n19752 = pi5  & n19749;
  assign n19753 = ~n19749 & ~n19750;
  assign n19754 = ~pi5  & ~n19749;
  assign n19755 = ~n41100 & ~n41101;
  assign n19756 = n19740 & ~n19755;
  assign n19757 = ~n19740 & n19755;
  assign n19758 = n19740 & ~n19756;
  assign n19759 = ~n19755 & ~n19756;
  assign n19760 = ~n19758 & ~n19759;
  assign n19761 = ~n19756 & ~n19757;
  assign n19762 = n19241 & ~n41102;
  assign n19763 = ~n19241 & n41102;
  assign n19764 = ~n41102 & ~n19762;
  assign n19765 = n19241 & ~n19762;
  assign n19766 = ~n19764 & ~n19765;
  assign n19767 = ~n19762 & ~n19763;
  assign n19768 = n19222 & n41103;
  assign n19769 = ~n19222 & ~n41103;
  assign n19770 = ~n19768 & ~n19769;
  assign n19771 = ~n19216 & ~n19219;
  assign n19772 = n19770 & ~n19771;
  assign n19773 = ~n19770 & n19771;
  assign po65  = ~n19772 & ~n19773;
  assign n19775 = n13010 & n15111;
  assign n19776 = pi122  & n39810;
  assign n19777 = pi124  & n13040;
  assign n19778 = pi123  & n13042;
  assign n19779 = ~n19777 & ~n19778;
  assign n19780 = ~n19776 & ~n19778;
  assign n19781 = ~n19777 & n19780;
  assign n19782 = ~n19776 & n19779;
  assign n19783 = ~n19775 & n41104;
  assign n19784 = pi8  & ~n19783;
  assign n19785 = pi8  & ~n19784;
  assign n19786 = pi8  & n19783;
  assign n19787 = ~n19783 & ~n19784;
  assign n19788 = ~pi8  & ~n19783;
  assign n19789 = ~n41105 & ~n41106;
  assign n19790 = ~n19714 & ~n19731;
  assign n19791 = ~n19715 & ~n19733;
  assign n19792 = ~n19715 & ~n19790;
  assign n19793 = ~n19789 & ~n41107;
  assign n19794 = n19789 & n41107;
  assign n19795 = ~n19789 & ~n19793;
  assign n19796 = ~n19789 & n41107;
  assign n19797 = ~n41107 & ~n19793;
  assign n19798 = n19789 & ~n41107;
  assign n19799 = ~n41108 & ~n41109;
  assign n19800 = ~n19793 & ~n19794;
  assign n19801 = n269 & n15091;
  assign n19802 = pi119  & n37475;
  assign n19803 = pi121  & n536;
  assign n19804 = pi120  & n538;
  assign n19805 = ~n19803 & ~n19804;
  assign n19806 = ~n19802 & ~n19804;
  assign n19807 = ~n19803 & n19806;
  assign n19808 = ~n19802 & n19805;
  assign n19809 = ~n19801 & n41111;
  assign n19810 = pi11  & ~n19809;
  assign n19811 = pi11  & ~n19810;
  assign n19812 = pi11  & n19809;
  assign n19813 = ~n19809 & ~n19810;
  assign n19814 = ~pi11  & ~n19809;
  assign n19815 = ~n41112 & ~n41113;
  assign n19816 = ~n19688 & ~n19697;
  assign n19817 = n19815 & n19816;
  assign n19818 = ~n19815 & ~n19816;
  assign n19819 = ~n19817 & ~n19818;
  assign n19820 = n523 & n8175;
  assign n19821 = pi113  & n38895;
  assign n19822 = pi115  & n8190;
  assign n19823 = pi114  & n8192;
  assign n19824 = ~n19822 & ~n19823;
  assign n19825 = ~n19821 & ~n19823;
  assign n19826 = ~n19822 & n19825;
  assign n19827 = ~n19821 & n19824;
  assign n19828 = ~n19820 & n41114;
  assign n19829 = pi17  & ~n19828;
  assign n19830 = pi17  & ~n19829;
  assign n19831 = pi17  & n19828;
  assign n19832 = ~n19828 & ~n19829;
  assign n19833 = ~pi17  & ~n19828;
  assign n19834 = ~n41115 & ~n41116;
  assign n19835 = ~n19651 & ~n19659;
  assign n19836 = n19834 & n19835;
  assign n19837 = ~n19834 & ~n19835;
  assign n19838 = ~n19836 & ~n19837;
  assign n19839 = n6785 & n10844;
  assign n19840 = pi110  & n38631;
  assign n19841 = pi112  & n6800;
  assign n19842 = pi111  & n6802;
  assign n19843 = ~n19841 & ~n19842;
  assign n19844 = ~n19840 & ~n19842;
  assign n19845 = ~n19841 & n19844;
  assign n19846 = ~n19840 & n19843;
  assign n19847 = ~n19839 & n41117;
  assign n19848 = pi20  & ~n19847;
  assign n19849 = pi20  & ~n19848;
  assign n19850 = pi20  & n19847;
  assign n19851 = ~n19847 & ~n19848;
  assign n19852 = ~pi20  & ~n19847;
  assign n19853 = ~n41118 & ~n41119;
  assign n19854 = ~n19640 & ~n19648;
  assign n19855 = n19853 & n19854;
  assign n19856 = ~n19853 & ~n19854;
  assign n19857 = ~n19855 & ~n19856;
  assign n19858 = n4492 & n8209;
  assign n19859 = pi104  & n38208;
  assign n19860 = pi106  & n4507;
  assign n19861 = pi105  & n4509;
  assign n19862 = ~n19860 & ~n19861;
  assign n19863 = ~n19859 & ~n19861;
  assign n19864 = ~n19860 & n19863;
  assign n19865 = ~n19859 & n19862;
  assign n19866 = ~n19858 & n41120;
  assign n19867 = pi26  & ~n19866;
  assign n19868 = pi26  & ~n19867;
  assign n19869 = pi26  & n19866;
  assign n19870 = ~n19866 & ~n19867;
  assign n19871 = ~pi26  & ~n19866;
  assign n19872 = ~n41121 & ~n41122;
  assign n19873 = ~n19602 & ~n19611;
  assign n19874 = n19872 & n19873;
  assign n19875 = ~n19872 & ~n19873;
  assign n19876 = ~n19874 & ~n19875;
  assign n19877 = ~n19576 & ~n19585;
  assign n19878 = n607 & n6787;
  assign n19879 = pi101  & n37489;
  assign n19880 = pi103  & n620;
  assign n19881 = pi102  & n622;
  assign n19882 = ~n19880 & ~n19881;
  assign n19883 = ~n19879 & ~n19881;
  assign n19884 = ~n19880 & n19883;
  assign n19885 = ~n19879 & n19882;
  assign n19886 = ~n607 & n41123;
  assign n19887 = ~n6787 & n41123;
  assign n19888 = ~n19886 & ~n19887;
  assign n19889 = ~n19878 & n41123;
  assign n19890 = pi29  & ~n41124;
  assign n19891 = ~pi29  & n41124;
  assign n19892 = ~n19890 & ~n19891;
  assign n19893 = ~n19877 & ~n19892;
  assign n19894 = n19877 & n19892;
  assign n19895 = ~n19893 & ~n19894;
  assign n19896 = n649 & n6474;
  assign n19897 = pi98  & n37496;
  assign n19898 = pi100  & n662;
  assign n19899 = pi99  & n664;
  assign n19900 = ~n19898 & ~n19899;
  assign n19901 = ~n19897 & ~n19899;
  assign n19902 = ~n19898 & n19901;
  assign n19903 = ~n19897 & n19900;
  assign n19904 = ~n649 & n41125;
  assign n19905 = ~n6474 & n41125;
  assign n19906 = ~n19904 & ~n19905;
  assign n19907 = ~n19896 & n41125;
  assign n19908 = pi32  & ~n41126;
  assign n19909 = ~pi32  & n41126;
  assign n19910 = ~n19908 & ~n19909;
  assign n19911 = ~n19572 & ~n19910;
  assign n19912 = n19572 & n19910;
  assign n19913 = ~n19572 & ~n19911;
  assign n19914 = ~n19572 & n19910;
  assign n19915 = ~n19910 & ~n19911;
  assign n19916 = n19572 & ~n19910;
  assign n19917 = ~n41127 & ~n41128;
  assign n19918 = ~n19911 & ~n19912;
  assign n19919 = ~n19512 & ~n19521;
  assign n19920 = ~n19491 & ~n19495;
  assign n19921 = ~n19456 & ~n19460;
  assign n19922 = ~n19442 & ~n19450;
  assign n19923 = ~n19422 & ~n19424;
  assign n19924 = n1465 & n4312;
  assign n19925 = pi74  & n38376;
  assign n19926 = pi76  & n4314;
  assign n19927 = pi75  & n4322;
  assign n19928 = ~n19926 & ~n19927;
  assign n19929 = ~n19925 & ~n19927;
  assign n19930 = ~n19926 & n19929;
  assign n19931 = ~n19925 & n19928;
  assign n19932 = ~n19924 & n41130;
  assign n19933 = pi56  & ~n19932;
  assign n19934 = pi56  & ~n19933;
  assign n19935 = pi56  & n19932;
  assign n19936 = ~n19932 & ~n19933;
  assign n19937 = ~pi56  & ~n19932;
  assign n19938 = ~n41131 & ~n41132;
  assign n19939 = ~n19383 & ~n19392;
  assign n19940 = pi67  & ~n40814;
  assign n19941 = pi66  & n18285;
  assign n19942 = ~n19940 & ~n19941;
  assign n19943 = pi2  & ~n19942;
  assign n19944 = ~pi2  & n19942;
  assign n19945 = ~n19943 & ~n19944;
  assign n19946 = n972 & n12674;
  assign n19947 = pi68  & n40107;
  assign n19948 = pi70  & n12676;
  assign n19949 = pi69  & n12684;
  assign n19950 = ~n19948 & ~n19949;
  assign n19951 = ~n19947 & ~n19949;
  assign n19952 = ~n19948 & n19951;
  assign n19953 = ~n19947 & n19950;
  assign n19954 = ~n12674 & n41133;
  assign n19955 = ~n972 & n41133;
  assign n19956 = ~n19954 & ~n19955;
  assign n19957 = ~n19946 & n41133;
  assign n19958 = pi62  & ~n41134;
  assign n19959 = ~pi62  & n41134;
  assign n19960 = ~n19958 & ~n19959;
  assign n19961 = n19945 & ~n19960;
  assign n19962 = ~n19945 & n19960;
  assign n19963 = ~n19961 & ~n19962;
  assign n19964 = ~n19939 & n19963;
  assign n19965 = n19939 & ~n19963;
  assign n19966 = ~n19964 & ~n19965;
  assign n19967 = n1238 & n7882;
  assign n19968 = pi71  & n39128;
  assign n19969 = pi73  & n7884;
  assign n19970 = pi72  & n7892;
  assign n19971 = ~n19969 & ~n19970;
  assign n19972 = ~n19968 & ~n19970;
  assign n19973 = ~n19969 & n19972;
  assign n19974 = ~n19968 & n19971;
  assign n19975 = ~n19967 & n41135;
  assign n19976 = pi59  & ~n19975;
  assign n19977 = pi59  & ~n19976;
  assign n19978 = pi59  & n19975;
  assign n19979 = ~n19975 & ~n19976;
  assign n19980 = ~pi59  & ~n19975;
  assign n19981 = ~n41136 & ~n41137;
  assign n19982 = n19966 & ~n19981;
  assign n19983 = ~n19966 & n19981;
  assign n19984 = n19966 & ~n19982;
  assign n19985 = ~n19981 & ~n19982;
  assign n19986 = ~n19984 & ~n19985;
  assign n19987 = ~n19982 & ~n19983;
  assign n19988 = ~n19417 & ~n41138;
  assign n19989 = n19417 & n41138;
  assign n19990 = ~n19417 & n41138;
  assign n19991 = n19417 & ~n41138;
  assign n19992 = ~n19990 & ~n19991;
  assign n19993 = ~n19988 & ~n19989;
  assign n19994 = n19938 & n41139;
  assign n19995 = ~n19938 & ~n41139;
  assign n19996 = ~n19994 & ~n19995;
  assign n19997 = ~n19923 & n19996;
  assign n19998 = n19923 & ~n19996;
  assign n19999 = ~n19997 & ~n19998;
  assign n20000 = n678 & n1971;
  assign n20001 = pi77  & n37864;
  assign n20002 = pi79  & n1973;
  assign n20003 = pi78  & n1981;
  assign n20004 = ~n20002 & ~n20003;
  assign n20005 = ~n20001 & ~n20003;
  assign n20006 = ~n20002 & n20005;
  assign n20007 = ~n20001 & n20004;
  assign n20008 = ~n20000 & n41140;
  assign n20009 = pi53  & ~n20008;
  assign n20010 = pi53  & ~n20009;
  assign n20011 = pi53  & n20008;
  assign n20012 = ~n20008 & ~n20009;
  assign n20013 = ~pi53  & ~n20008;
  assign n20014 = ~n41141 & ~n41142;
  assign n20015 = n19999 & ~n20014;
  assign n20016 = ~n19999 & n20014;
  assign n20017 = n19999 & ~n20015;
  assign n20018 = ~n20014 & ~n20015;
  assign n20019 = ~n20017 & ~n20018;
  assign n20020 = ~n20015 & ~n20016;
  assign n20021 = n19922 & n41143;
  assign n20022 = ~n19922 & ~n41143;
  assign n20023 = ~n20021 & ~n20022;
  assign n20024 = n894 & n2134;
  assign n20025 = pi80  & n37580;
  assign n20026 = pi82  & n896;
  assign n20027 = pi81  & n904;
  assign n20028 = ~n20026 & ~n20027;
  assign n20029 = ~n20025 & ~n20027;
  assign n20030 = ~n20026 & n20029;
  assign n20031 = ~n20025 & n20028;
  assign n20032 = ~n20024 & n41144;
  assign n20033 = pi50  & ~n20032;
  assign n20034 = pi50  & ~n20033;
  assign n20035 = pi50  & n20032;
  assign n20036 = ~n20032 & ~n20033;
  assign n20037 = ~pi50  & ~n20032;
  assign n20038 = ~n41145 & ~n41146;
  assign n20039 = ~n20023 & n20038;
  assign n20040 = n20023 & ~n20038;
  assign n20041 = n20023 & ~n20040;
  assign n20042 = ~n20038 & ~n20040;
  assign n20043 = ~n20041 & ~n20042;
  assign n20044 = ~n20039 & ~n20040;
  assign n20045 = n19921 & n41147;
  assign n20046 = ~n19921 & ~n41147;
  assign n20047 = ~n20045 & ~n20046;
  assign n20048 = n785 & n2804;
  assign n20049 = pi83  & n37520;
  assign n20050 = pi85  & n787;
  assign n20051 = pi84  & n795;
  assign n20052 = ~n20050 & ~n20051;
  assign n20053 = ~n20049 & ~n20051;
  assign n20054 = ~n20050 & n20053;
  assign n20055 = ~n20049 & n20052;
  assign n20056 = ~n20048 & n41148;
  assign n20057 = pi47  & ~n20056;
  assign n20058 = pi47  & ~n20057;
  assign n20059 = pi47  & n20056;
  assign n20060 = ~n20056 & ~n20057;
  assign n20061 = ~pi47  & ~n20056;
  assign n20062 = ~n41149 & ~n41150;
  assign n20063 = ~n20047 & n20062;
  assign n20064 = n20047 & ~n20062;
  assign n20065 = ~n20063 & ~n20064;
  assign n20066 = ~n19477 & ~n19485;
  assign n20067 = n20065 & ~n20066;
  assign n20068 = ~n20065 & n20066;
  assign n20069 = ~n20067 & ~n20068;
  assign n20070 = n940 & n3354;
  assign n20071 = pi86  & n37541;
  assign n20072 = pi88  & n953;
  assign n20073 = pi87  & n955;
  assign n20074 = ~n20072 & ~n20073;
  assign n20075 = ~n20071 & ~n20073;
  assign n20076 = ~n20072 & n20075;
  assign n20077 = ~n20071 & n20074;
  assign n20078 = ~n20070 & n41151;
  assign n20079 = pi44  & ~n20078;
  assign n20080 = pi44  & ~n20079;
  assign n20081 = pi44  & n20078;
  assign n20082 = ~n20078 & ~n20079;
  assign n20083 = ~pi44  & ~n20078;
  assign n20084 = ~n41152 & ~n41153;
  assign n20085 = ~n20069 & n20084;
  assign n20086 = n20069 & ~n20084;
  assign n20087 = n20069 & ~n20086;
  assign n20088 = ~n20084 & ~n20086;
  assign n20089 = ~n20087 & ~n20088;
  assign n20090 = ~n20085 & ~n20086;
  assign n20091 = n19920 & n41154;
  assign n20092 = ~n19920 & ~n41154;
  assign n20093 = ~n20091 & ~n20092;
  assign n20094 = n594 & n733;
  assign n20095 = pi89  & n37510;
  assign n20096 = pi91  & n746;
  assign n20097 = pi90  & n748;
  assign n20098 = ~n20096 & ~n20097;
  assign n20099 = ~n20095 & ~n20097;
  assign n20100 = ~n20096 & n20099;
  assign n20101 = ~n20095 & n20098;
  assign n20102 = ~n20094 & n41155;
  assign n20103 = pi41  & ~n20102;
  assign n20104 = pi41  & ~n20103;
  assign n20105 = pi41  & n20102;
  assign n20106 = ~n20102 & ~n20103;
  assign n20107 = ~pi41  & ~n20102;
  assign n20108 = ~n41156 & ~n41157;
  assign n20109 = n20093 & ~n20108;
  assign n20110 = ~n20093 & n20108;
  assign n20111 = n20093 & ~n20109;
  assign n20112 = ~n20108 & ~n20109;
  assign n20113 = ~n20111 & ~n20112;
  assign n20114 = ~n20109 & ~n20110;
  assign n20115 = n19919 & n41158;
  assign n20116 = ~n19919 & ~n41158;
  assign n20117 = ~n20115 & ~n20116;
  assign n20118 = n691 & n4524;
  assign n20119 = pi92  & n37503;
  assign n20120 = pi94  & n704;
  assign n20121 = pi93  & n706;
  assign n20122 = ~n20120 & ~n20121;
  assign n20123 = ~n20119 & ~n20121;
  assign n20124 = ~n20120 & n20123;
  assign n20125 = ~n20119 & n20122;
  assign n20126 = ~n20118 & n41159;
  assign n20127 = pi38  & ~n20126;
  assign n20128 = pi38  & ~n20127;
  assign n20129 = pi38  & n20126;
  assign n20130 = ~n20126 & ~n20127;
  assign n20131 = ~pi38  & ~n20126;
  assign n20132 = ~n41160 & ~n41161;
  assign n20133 = ~n20117 & n20132;
  assign n20134 = n20117 & ~n20132;
  assign n20135 = ~n20133 & ~n20134;
  assign n20136 = ~n19538 & ~n19547;
  assign n20137 = n20135 & ~n20136;
  assign n20138 = ~n20135 & n20136;
  assign n20139 = ~n20137 & ~n20138;
  assign n20140 = n2104 & n5630;
  assign n20141 = pi95  & n37758;
  assign n20142 = pi97  & n2117;
  assign n20143 = pi96  & n2119;
  assign n20144 = ~n20142 & ~n20143;
  assign n20145 = ~n20141 & ~n20143;
  assign n20146 = ~n20142 & n20145;
  assign n20147 = ~n20141 & n20144;
  assign n20148 = ~n20140 & n41162;
  assign n20149 = pi35  & ~n20148;
  assign n20150 = pi35  & ~n20149;
  assign n20151 = pi35  & n20148;
  assign n20152 = ~n20148 & ~n20149;
  assign n20153 = ~pi35  & ~n20148;
  assign n20154 = ~n41163 & ~n41164;
  assign n20155 = ~n20139 & n20154;
  assign n20156 = n20139 & ~n20154;
  assign n20157 = n20139 & ~n20156;
  assign n20158 = ~n20154 & ~n20156;
  assign n20159 = ~n20157 & ~n20158;
  assign n20160 = ~n20155 & ~n20156;
  assign n20161 = ~n41129 & ~n41165;
  assign n20162 = n41129 & n41165;
  assign n20163 = ~n41165 & ~n20161;
  assign n20164 = ~n41129 & ~n20161;
  assign n20165 = ~n20163 & ~n20164;
  assign n20166 = ~n20161 & ~n20162;
  assign n20167 = n19895 & ~n41166;
  assign n20168 = ~n19895 & n41166;
  assign n20169 = n19895 & ~n20167;
  assign n20170 = ~n41166 & ~n20167;
  assign n20171 = ~n20169 & ~n20170;
  assign n20172 = ~n20167 & ~n20168;
  assign n20173 = n19876 & ~n41167;
  assign n20174 = ~n19876 & n41167;
  assign n20175 = ~n20173 & ~n20174;
  assign n20176 = n5576 & n9701;
  assign n20177 = pi107  & n38406;
  assign n20178 = pi109  & n5591;
  assign n20179 = pi108  & n5593;
  assign n20180 = ~n20178 & ~n20179;
  assign n20181 = ~n20177 & ~n20179;
  assign n20182 = ~n20178 & n20181;
  assign n20183 = ~n20177 & n20180;
  assign n20184 = ~n20176 & n41168;
  assign n20185 = pi23  & ~n20184;
  assign n20186 = pi23  & ~n20185;
  assign n20187 = pi23  & n20184;
  assign n20188 = ~n20184 & ~n20185;
  assign n20189 = ~pi23  & ~n20184;
  assign n20190 = ~n41169 & ~n41170;
  assign n20191 = ~n19636 & ~n20190;
  assign n20192 = n19636 & n20190;
  assign n20193 = ~n19636 & n20190;
  assign n20194 = n19636 & ~n20190;
  assign n20195 = ~n20193 & ~n20194;
  assign n20196 = ~n20191 & ~n20192;
  assign n20197 = ~n20174 & ~n41171;
  assign n20198 = ~n20173 & n20197;
  assign n20199 = n20175 & ~n41171;
  assign n20200 = ~n20175 & n41171;
  assign n20201 = ~n41171 & ~n41172;
  assign n20202 = ~n20174 & ~n41172;
  assign n20203 = ~n20173 & n20202;
  assign n20204 = n20175 & ~n41172;
  assign n20205 = ~n20201 & ~n41173;
  assign n20206 = ~n41172 & ~n20200;
  assign n20207 = n19857 & ~n41174;
  assign n20208 = ~n19857 & n41174;
  assign n20209 = ~n20207 & ~n20208;
  assign n20210 = n19838 & ~n20208;
  assign n20211 = ~n20207 & n20210;
  assign n20212 = n19838 & n20209;
  assign n20213 = ~n19838 & ~n20209;
  assign n20214 = n19838 & ~n41175;
  assign n20215 = ~n20208 & ~n41175;
  assign n20216 = ~n20207 & n20215;
  assign n20217 = n20209 & ~n41175;
  assign n20218 = ~n20214 & ~n41176;
  assign n20219 = ~n41175 & ~n20213;
  assign n20220 = ~n19668 & ~n19670;
  assign n20221 = n563 & n13057;
  assign n20222 = pi116  & n37482;
  assign n20223 = pi118  & n578;
  assign n20224 = pi117  & n580;
  assign n20225 = ~n20223 & ~n20224;
  assign n20226 = ~n20222 & ~n20224;
  assign n20227 = ~n20223 & n20226;
  assign n20228 = ~n20222 & n20225;
  assign n20229 = ~n563 & n41178;
  assign n20230 = ~n13057 & n41178;
  assign n20231 = ~n20229 & ~n20230;
  assign n20232 = ~n20221 & n41178;
  assign n20233 = pi14  & ~n41179;
  assign n20234 = ~pi14  & n41179;
  assign n20235 = ~n20233 & ~n20234;
  assign n20236 = ~n20220 & ~n20235;
  assign n20237 = n20220 & n20235;
  assign n20238 = ~n20220 & ~n20236;
  assign n20239 = ~n20220 & n20235;
  assign n20240 = ~n20235 & ~n20236;
  assign n20241 = n20220 & ~n20235;
  assign n20242 = ~n41180 & ~n41181;
  assign n20243 = ~n20236 & ~n20237;
  assign n20244 = ~n41177 & ~n41182;
  assign n20245 = n41177 & n41182;
  assign n20246 = ~n41177 & ~n20244;
  assign n20247 = ~n41177 & n41182;
  assign n20248 = ~n41182 & ~n20244;
  assign n20249 = n41177 & ~n41182;
  assign n20250 = ~n41183 & ~n41184;
  assign n20251 = ~n20244 & ~n20245;
  assign n20252 = n19819 & ~n41185;
  assign n20253 = ~n41185 & ~n20252;
  assign n20254 = ~n19819 & ~n41185;
  assign n20255 = n19819 & ~n20252;
  assign n20256 = n19819 & n41185;
  assign n20257 = ~n19819 & n41185;
  assign n20258 = ~n20252 & ~n20257;
  assign n20259 = ~n41186 & ~n41187;
  assign n20260 = ~n41110 & n41188;
  assign n20261 = n41110 & ~n41188;
  assign n20262 = n41188 & ~n20260;
  assign n20263 = ~n41110 & ~n20260;
  assign n20264 = ~n20262 & ~n20263;
  assign n20265 = ~n20260 & ~n20261;
  assign n20266 = n14944 & n40885;
  assign n20267 = pi125  & n40177;
  assign n20268 = pi127  & n14974;
  assign n20269 = pi126  & n14976;
  assign n20270 = ~n20268 & ~n20269;
  assign n20271 = ~n20267 & ~n20269;
  assign n20272 = ~n20268 & n20271;
  assign n20273 = ~n20267 & n20270;
  assign n20274 = ~n20266 & n41190;
  assign n20275 = pi5  & ~n20274;
  assign n20276 = pi5  & ~n20275;
  assign n20277 = pi5  & n20274;
  assign n20278 = ~n20274 & ~n20275;
  assign n20279 = ~pi5  & ~n20274;
  assign n20280 = ~n41191 & ~n41192;
  assign n20281 = ~n19739 & n19755;
  assign n20282 = ~n19739 & ~n19756;
  assign n20283 = ~n19738 & ~n20281;
  assign n20284 = ~n20280 & ~n41193;
  assign n20285 = n20280 & n41193;
  assign n20286 = ~n41193 & ~n20284;
  assign n20287 = n20280 & ~n41193;
  assign n20288 = ~n20280 & ~n20284;
  assign n20289 = ~n20280 & n41193;
  assign n20290 = ~n41194 & ~n41195;
  assign n20291 = ~n20284 & ~n20285;
  assign n20292 = ~n41189 & ~n41196;
  assign n20293 = n41189 & n41196;
  assign n20294 = ~n41196 & ~n20292;
  assign n20295 = n41189 & ~n41196;
  assign n20296 = ~n41189 & ~n20292;
  assign n20297 = ~n41189 & n41196;
  assign n20298 = ~n41197 & ~n41198;
  assign n20299 = ~n20292 & ~n20293;
  assign n20300 = ~n19239 & n41102;
  assign n20301 = ~n19239 & ~n19762;
  assign n20302 = ~n19240 & ~n20300;
  assign n20303 = n41199 & n41200;
  assign n20304 = ~n41199 & ~n41200;
  assign n20305 = ~n20303 & ~n20304;
  assign n20306 = ~n19769 & ~n19772;
  assign n20307 = n20305 & ~n20306;
  assign n20308 = ~n20305 & n20306;
  assign po66  = ~n20307 & ~n20308;
  assign n20310 = ~n20304 & ~n20307;
  assign n20311 = ~n20284 & ~n20292;
  assign n20312 = n563 & n13027;
  assign n20313 = pi117  & n37482;
  assign n20314 = pi119  & n578;
  assign n20315 = pi118  & n580;
  assign n20316 = ~n20314 & ~n20315;
  assign n20317 = ~n20313 & ~n20315;
  assign n20318 = ~n20314 & n20317;
  assign n20319 = ~n20313 & n20316;
  assign n20320 = ~n20312 & n41201;
  assign n20321 = pi14  & ~n20320;
  assign n20322 = pi14  & ~n20321;
  assign n20323 = pi14  & n20320;
  assign n20324 = ~n20320 & ~n20321;
  assign n20325 = ~pi14  & ~n20320;
  assign n20326 = ~n41202 & ~n41203;
  assign n20327 = ~n19837 & ~n41175;
  assign n20328 = n20326 & n20327;
  assign n20329 = ~n20326 & ~n20327;
  assign n20330 = ~n20328 & ~n20329;
  assign n20331 = n8175 & n12530;
  assign n20332 = pi114  & n38895;
  assign n20333 = pi116  & n8190;
  assign n20334 = pi115  & n8192;
  assign n20335 = ~n20333 & ~n20334;
  assign n20336 = ~n20332 & ~n20334;
  assign n20337 = ~n20333 & n20336;
  assign n20338 = ~n20332 & n20335;
  assign n20339 = ~n20331 & n41204;
  assign n20340 = pi17  & ~n20339;
  assign n20341 = pi17  & ~n20340;
  assign n20342 = pi17  & n20339;
  assign n20343 = ~n20339 & ~n20340;
  assign n20344 = ~pi17  & ~n20339;
  assign n20345 = ~n41205 & ~n41206;
  assign n20346 = ~n19856 & ~n20207;
  assign n20347 = ~n20345 & ~n20346;
  assign n20348 = n20345 & n20346;
  assign n20349 = ~n20345 & ~n20347;
  assign n20350 = ~n20345 & n20346;
  assign n20351 = ~n20346 & ~n20347;
  assign n20352 = n20345 & ~n20346;
  assign n20353 = ~n41207 & ~n41208;
  assign n20354 = ~n20347 & ~n20348;
  assign n20355 = n6785 & n11276;
  assign n20356 = pi111  & n38631;
  assign n20357 = pi113  & n6800;
  assign n20358 = pi112  & n6802;
  assign n20359 = ~n20357 & ~n20358;
  assign n20360 = ~n20356 & ~n20358;
  assign n20361 = ~n20357 & n20360;
  assign n20362 = ~n20356 & n20359;
  assign n20363 = ~n20355 & n41210;
  assign n20364 = pi20  & ~n20363;
  assign n20365 = pi20  & ~n20364;
  assign n20366 = pi20  & n20363;
  assign n20367 = ~n20363 & ~n20364;
  assign n20368 = ~pi20  & ~n20363;
  assign n20369 = ~n41211 & ~n41212;
  assign n20370 = ~n20191 & ~n41172;
  assign n20371 = n20369 & n20370;
  assign n20372 = ~n20369 & ~n20370;
  assign n20373 = ~n20371 & ~n20372;
  assign n20374 = n4492 & n8177;
  assign n20375 = pi105  & n38208;
  assign n20376 = pi107  & n4507;
  assign n20377 = pi106  & n4509;
  assign n20378 = ~n20376 & ~n20377;
  assign n20379 = ~n20375 & ~n20377;
  assign n20380 = ~n20376 & n20379;
  assign n20381 = ~n20375 & n20378;
  assign n20382 = ~n20374 & n41213;
  assign n20383 = pi26  & ~n20382;
  assign n20384 = pi26  & ~n20383;
  assign n20385 = pi26  & n20382;
  assign n20386 = ~n20382 & ~n20383;
  assign n20387 = ~pi26  & ~n20382;
  assign n20388 = ~n41214 & ~n41215;
  assign n20389 = ~n19893 & ~n20167;
  assign n20390 = n20388 & n20389;
  assign n20391 = ~n20388 & ~n20389;
  assign n20392 = ~n20390 & ~n20391;
  assign n20393 = n649 & n6839;
  assign n20394 = pi99  & n37496;
  assign n20395 = pi101  & n662;
  assign n20396 = pi100  & n664;
  assign n20397 = ~n20395 & ~n20396;
  assign n20398 = ~n20394 & ~n20396;
  assign n20399 = ~n20395 & n20398;
  assign n20400 = ~n20394 & n20397;
  assign n20401 = ~n649 & n41216;
  assign n20402 = ~n6839 & n41216;
  assign n20403 = ~n20401 & ~n20402;
  assign n20404 = ~n20393 & n41216;
  assign n20405 = pi32  & ~n41217;
  assign n20406 = ~pi32  & n41217;
  assign n20407 = ~n20405 & ~n20406;
  assign n20408 = ~n20138 & ~n20154;
  assign n20409 = ~n20137 & ~n20156;
  assign n20410 = ~n20137 & ~n20408;
  assign n20411 = ~n20407 & ~n41218;
  assign n20412 = n20407 & n41218;
  assign n20413 = ~n20411 & ~n20412;
  assign n20414 = n2104 & n5610;
  assign n20415 = pi96  & n37758;
  assign n20416 = pi98  & n2117;
  assign n20417 = pi97  & n2119;
  assign n20418 = ~n20416 & ~n20417;
  assign n20419 = ~n20415 & ~n20417;
  assign n20420 = ~n20416 & n20419;
  assign n20421 = ~n20415 & n20418;
  assign n20422 = ~n20414 & n41219;
  assign n20423 = pi35  & ~n20422;
  assign n20424 = pi35  & ~n20423;
  assign n20425 = pi35  & n20422;
  assign n20426 = ~n20422 & ~n20423;
  assign n20427 = ~pi35  & ~n20422;
  assign n20428 = ~n41220 & ~n41221;
  assign n20429 = ~n20116 & ~n20134;
  assign n20430 = n940 & n3591;
  assign n20431 = pi87  & n37541;
  assign n20432 = pi89  & n953;
  assign n20433 = pi88  & n955;
  assign n20434 = ~n20432 & ~n20433;
  assign n20435 = ~n20431 & ~n20433;
  assign n20436 = ~n20432 & n20435;
  assign n20437 = ~n20431 & n20434;
  assign n20438 = ~n20430 & n41222;
  assign n20439 = pi44  & ~n20438;
  assign n20440 = pi44  & ~n20439;
  assign n20441 = pi44  & n20438;
  assign n20442 = ~n20438 & ~n20439;
  assign n20443 = ~pi44  & ~n20438;
  assign n20444 = ~n41223 & ~n41224;
  assign n20445 = ~n20046 & ~n20064;
  assign n20446 = ~n19943 & ~n19961;
  assign n20447 = n927 & n12674;
  assign n20448 = pi69  & n40107;
  assign n20449 = pi71  & n12676;
  assign n20450 = pi70  & n12684;
  assign n20451 = ~n20449 & ~n20450;
  assign n20452 = ~n20448 & ~n20450;
  assign n20453 = ~n20449 & n20452;
  assign n20454 = ~n20448 & n20451;
  assign n20455 = ~n20447 & n41225;
  assign n20456 = pi62  & ~n20455;
  assign n20457 = pi62  & ~n20456;
  assign n20458 = pi62  & n20455;
  assign n20459 = ~n20455 & ~n20456;
  assign n20460 = ~pi62  & ~n20455;
  assign n20461 = ~n41226 & ~n41227;
  assign n20462 = pi68  & ~n40814;
  assign n20463 = pi67  & n18285;
  assign n20464 = ~n20462 & ~n20463;
  assign n20465 = pi2  & ~n20464;
  assign n20466 = ~pi2  & n20464;
  assign n20467 = pi2  & ~n20465;
  assign n20468 = pi2  & n20464;
  assign n20469 = ~n20464 & ~n20465;
  assign n20470 = ~pi2  & ~n20464;
  assign n20471 = ~n41228 & ~n41229;
  assign n20472 = ~n20465 & ~n20466;
  assign n20473 = ~n20461 & ~n41230;
  assign n20474 = n20461 & n41230;
  assign n20475 = ~n20461 & ~n20473;
  assign n20476 = ~n20461 & n41230;
  assign n20477 = ~n41230 & ~n20473;
  assign n20478 = n20461 & ~n41230;
  assign n20479 = ~n41231 & ~n41232;
  assign n20480 = ~n20473 & ~n20474;
  assign n20481 = n20446 & n41233;
  assign n20482 = ~n20446 & ~n41233;
  assign n20483 = ~n20481 & ~n20482;
  assign n20484 = n1218 & n7882;
  assign n20485 = pi72  & n39128;
  assign n20486 = pi74  & n7884;
  assign n20487 = pi73  & n7892;
  assign n20488 = ~n20486 & ~n20487;
  assign n20489 = ~n20485 & ~n20487;
  assign n20490 = ~n20486 & n20489;
  assign n20491 = ~n20485 & n20488;
  assign n20492 = ~n20484 & n41234;
  assign n20493 = pi59  & ~n20492;
  assign n20494 = pi59  & ~n20493;
  assign n20495 = pi59  & n20492;
  assign n20496 = ~n20492 & ~n20493;
  assign n20497 = ~pi59  & ~n20492;
  assign n20498 = ~n41235 & ~n41236;
  assign n20499 = n20483 & ~n20498;
  assign n20500 = ~n20483 & n20498;
  assign n20501 = n20483 & ~n20499;
  assign n20502 = ~n20498 & ~n20499;
  assign n20503 = ~n20501 & ~n20502;
  assign n20504 = ~n20499 & ~n20500;
  assign n20505 = ~n19964 & n19981;
  assign n20506 = ~n19964 & ~n19982;
  assign n20507 = ~n19965 & ~n20505;
  assign n20508 = n41237 & n41238;
  assign n20509 = ~n41237 & ~n41238;
  assign n20510 = ~n20508 & ~n20509;
  assign n20511 = n1596 & n4312;
  assign n20512 = pi75  & n38376;
  assign n20513 = pi77  & n4314;
  assign n20514 = pi76  & n4322;
  assign n20515 = ~n20513 & ~n20514;
  assign n20516 = ~n20512 & ~n20514;
  assign n20517 = ~n20513 & n20516;
  assign n20518 = ~n20512 & n20515;
  assign n20519 = ~n20511 & n41239;
  assign n20520 = pi56  & ~n20519;
  assign n20521 = pi56  & ~n20520;
  assign n20522 = pi56  & n20519;
  assign n20523 = ~n20519 & ~n20520;
  assign n20524 = ~pi56  & ~n20519;
  assign n20525 = ~n41240 & ~n41241;
  assign n20526 = ~n20510 & n20525;
  assign n20527 = n20510 & ~n20525;
  assign n20528 = ~n20526 & ~n20527;
  assign n20529 = ~n19988 & ~n19995;
  assign n20530 = n20528 & ~n20529;
  assign n20531 = ~n20528 & n20529;
  assign n20532 = ~n20530 & ~n20531;
  assign n20533 = n1971 & n2063;
  assign n20534 = pi78  & n37864;
  assign n20535 = pi80  & n1973;
  assign n20536 = pi79  & n1981;
  assign n20537 = ~n20535 & ~n20536;
  assign n20538 = ~n20534 & ~n20536;
  assign n20539 = ~n20535 & n20538;
  assign n20540 = ~n20534 & n20537;
  assign n20541 = ~n20533 & n41242;
  assign n20542 = pi53  & ~n20541;
  assign n20543 = pi53  & ~n20542;
  assign n20544 = pi53  & n20541;
  assign n20545 = ~n20541 & ~n20542;
  assign n20546 = ~pi53  & ~n20541;
  assign n20547 = ~n41243 & ~n41244;
  assign n20548 = ~n20532 & n20547;
  assign n20549 = n20532 & ~n20547;
  assign n20550 = n20532 & ~n20549;
  assign n20551 = ~n20547 & ~n20549;
  assign n20552 = ~n20550 & ~n20551;
  assign n20553 = ~n20548 & ~n20549;
  assign n20554 = ~n19997 & n20014;
  assign n20555 = ~n19997 & ~n20015;
  assign n20556 = ~n19998 & ~n20554;
  assign n20557 = n41245 & n41246;
  assign n20558 = ~n41245 & ~n41246;
  assign n20559 = ~n20557 & ~n20558;
  assign n20560 = n894 & n2091;
  assign n20561 = pi81  & n37580;
  assign n20562 = pi83  & n896;
  assign n20563 = pi82  & n904;
  assign n20564 = ~n20562 & ~n20563;
  assign n20565 = ~n20561 & ~n20563;
  assign n20566 = ~n20562 & n20565;
  assign n20567 = ~n20561 & n20564;
  assign n20568 = ~n20560 & n41247;
  assign n20569 = pi50  & ~n20568;
  assign n20570 = pi50  & ~n20569;
  assign n20571 = pi50  & n20568;
  assign n20572 = ~n20568 & ~n20569;
  assign n20573 = ~pi50  & ~n20568;
  assign n20574 = ~n41248 & ~n41249;
  assign n20575 = n20559 & ~n20574;
  assign n20576 = ~n20559 & n20574;
  assign n20577 = n20559 & ~n20575;
  assign n20578 = ~n20574 & ~n20575;
  assign n20579 = ~n20577 & ~n20578;
  assign n20580 = ~n20575 & ~n20576;
  assign n20581 = ~n20022 & n20038;
  assign n20582 = ~n20022 & ~n20040;
  assign n20583 = ~n20021 & ~n20581;
  assign n20584 = n41250 & n41251;
  assign n20585 = ~n41250 & ~n41251;
  assign n20586 = ~n20584 & ~n20585;
  assign n20587 = n785 & n2779;
  assign n20588 = pi84  & n37520;
  assign n20589 = pi86  & n787;
  assign n20590 = pi85  & n795;
  assign n20591 = ~n20589 & ~n20590;
  assign n20592 = ~n20588 & ~n20590;
  assign n20593 = ~n20589 & n20592;
  assign n20594 = ~n20588 & n20591;
  assign n20595 = ~n20587 & n41252;
  assign n20596 = pi47  & ~n20595;
  assign n20597 = pi47  & ~n20596;
  assign n20598 = pi47  & n20595;
  assign n20599 = ~n20595 & ~n20596;
  assign n20600 = ~pi47  & ~n20595;
  assign n20601 = ~n41253 & ~n41254;
  assign n20602 = ~n20586 & n20601;
  assign n20603 = n20586 & ~n20601;
  assign n20604 = n20586 & ~n20603;
  assign n20605 = ~n20601 & ~n20603;
  assign n20606 = ~n20604 & ~n20605;
  assign n20607 = ~n20602 & ~n20603;
  assign n20608 = ~n20445 & ~n41255;
  assign n20609 = n20445 & n41255;
  assign n20610 = ~n41255 & ~n20608;
  assign n20611 = ~n20445 & ~n20608;
  assign n20612 = ~n20610 & ~n20611;
  assign n20613 = ~n20608 & ~n20609;
  assign n20614 = ~n20444 & ~n41256;
  assign n20615 = n20444 & n41256;
  assign n20616 = ~n41256 & ~n20614;
  assign n20617 = ~n20444 & ~n20614;
  assign n20618 = ~n20616 & ~n20617;
  assign n20619 = ~n20614 & ~n20615;
  assign n20620 = ~n20068 & ~n20084;
  assign n20621 = ~n20067 & ~n20086;
  assign n20622 = ~n20067 & ~n20620;
  assign n20623 = n41257 & n41258;
  assign n20624 = ~n41257 & ~n41258;
  assign n20625 = ~n20623 & ~n20624;
  assign n20626 = n733 & n4453;
  assign n20627 = pi90  & n37510;
  assign n20628 = pi92  & n746;
  assign n20629 = pi91  & n748;
  assign n20630 = ~n20628 & ~n20629;
  assign n20631 = ~n20627 & ~n20629;
  assign n20632 = ~n20628 & n20631;
  assign n20633 = ~n20627 & n20630;
  assign n20634 = ~n20626 & n41259;
  assign n20635 = pi41  & ~n20634;
  assign n20636 = pi41  & ~n20635;
  assign n20637 = pi41  & n20634;
  assign n20638 = ~n20634 & ~n20635;
  assign n20639 = ~pi41  & ~n20634;
  assign n20640 = ~n41260 & ~n41261;
  assign n20641 = ~n20625 & n20640;
  assign n20642 = n20625 & ~n20640;
  assign n20643 = n20625 & ~n20642;
  assign n20644 = ~n20640 & ~n20642;
  assign n20645 = ~n20643 & ~n20644;
  assign n20646 = ~n20641 & ~n20642;
  assign n20647 = ~n20092 & n20108;
  assign n20648 = ~n20092 & ~n20109;
  assign n20649 = ~n20091 & ~n20647;
  assign n20650 = n41262 & n41263;
  assign n20651 = ~n41262 & ~n41263;
  assign n20652 = ~n20650 & ~n20651;
  assign n20653 = n691 & n4494;
  assign n20654 = pi93  & n37503;
  assign n20655 = pi95  & n704;
  assign n20656 = pi94  & n706;
  assign n20657 = ~n20655 & ~n20656;
  assign n20658 = ~n20654 & ~n20656;
  assign n20659 = ~n20655 & n20658;
  assign n20660 = ~n20654 & n20657;
  assign n20661 = ~n20653 & n41264;
  assign n20662 = pi38  & ~n20661;
  assign n20663 = pi38  & ~n20662;
  assign n20664 = pi38  & n20661;
  assign n20665 = ~n20661 & ~n20662;
  assign n20666 = ~pi38  & ~n20661;
  assign n20667 = ~n41265 & ~n41266;
  assign n20668 = ~n20652 & n20667;
  assign n20669 = n20652 & ~n20667;
  assign n20670 = ~n20668 & ~n20669;
  assign n20671 = ~n20429 & n20670;
  assign n20672 = n20429 & ~n20670;
  assign n20673 = ~n20429 & ~n20671;
  assign n20674 = n20670 & ~n20671;
  assign n20675 = ~n20673 & ~n20674;
  assign n20676 = ~n20671 & ~n20672;
  assign n20677 = n20428 & n41267;
  assign n20678 = ~n20428 & ~n41267;
  assign n20679 = ~n20428 & ~n20678;
  assign n20680 = ~n41267 & ~n20678;
  assign n20681 = ~n20679 & ~n20680;
  assign n20682 = ~n20677 & ~n20678;
  assign n20683 = ~n20413 & n41268;
  assign n20684 = n20413 & ~n41268;
  assign n20685 = ~n20683 & ~n20684;
  assign n20686 = ~n19911 & ~n20161;
  assign n20687 = n607 & n8136;
  assign n20688 = pi102  & n37489;
  assign n20689 = pi104  & n620;
  assign n20690 = pi103  & n622;
  assign n20691 = ~n20689 & ~n20690;
  assign n20692 = ~n20688 & ~n20690;
  assign n20693 = ~n20689 & n20692;
  assign n20694 = ~n20688 & n20691;
  assign n20695 = ~n607 & n41269;
  assign n20696 = ~n8136 & n41269;
  assign n20697 = ~n20695 & ~n20696;
  assign n20698 = ~n20687 & n41269;
  assign n20699 = pi29  & ~n41270;
  assign n20700 = ~pi29  & n41270;
  assign n20701 = ~n20699 & ~n20700;
  assign n20702 = ~n20686 & ~n20701;
  assign n20703 = n20686 & n20701;
  assign n20704 = ~n20686 & ~n20702;
  assign n20705 = ~n20686 & n20701;
  assign n20706 = ~n20701 & ~n20702;
  assign n20707 = n20686 & ~n20701;
  assign n20708 = ~n41271 & ~n41272;
  assign n20709 = ~n20702 & ~n20703;
  assign n20710 = n20685 & ~n41273;
  assign n20711 = ~n20685 & n41273;
  assign n20712 = n20685 & ~n20710;
  assign n20713 = ~n41273 & ~n20710;
  assign n20714 = ~n20712 & ~n20713;
  assign n20715 = ~n20710 & ~n20711;
  assign n20716 = n20392 & ~n41274;
  assign n20717 = ~n20392 & n41274;
  assign n20718 = n20392 & ~n20716;
  assign n20719 = ~n41274 & ~n20716;
  assign n20720 = ~n20718 & ~n20719;
  assign n20721 = ~n20716 & ~n20717;
  assign n20722 = n5576 & n9678;
  assign n20723 = pi108  & n38406;
  assign n20724 = pi110  & n5591;
  assign n20725 = pi109  & n5593;
  assign n20726 = ~n20724 & ~n20725;
  assign n20727 = ~n20723 & ~n20725;
  assign n20728 = ~n20724 & n20727;
  assign n20729 = ~n20723 & n20726;
  assign n20730 = ~n20722 & n41276;
  assign n20731 = pi23  & ~n20730;
  assign n20732 = pi23  & ~n20731;
  assign n20733 = pi23  & n20730;
  assign n20734 = ~n20730 & ~n20731;
  assign n20735 = ~pi23  & ~n20730;
  assign n20736 = ~n41277 & ~n41278;
  assign n20737 = ~n19875 & ~n20173;
  assign n20738 = ~n20736 & ~n20737;
  assign n20739 = n20736 & n20737;
  assign n20740 = ~n20736 & ~n20738;
  assign n20741 = ~n20736 & n20737;
  assign n20742 = ~n20737 & ~n20738;
  assign n20743 = n20736 & ~n20737;
  assign n20744 = ~n41279 & ~n41280;
  assign n20745 = ~n20738 & ~n20739;
  assign n20746 = ~n41275 & ~n41281;
  assign n20747 = n41275 & n41281;
  assign n20748 = ~n41275 & n41281;
  assign n20749 = n41275 & ~n41281;
  assign n20750 = ~n20748 & ~n20749;
  assign n20751 = ~n20746 & ~n20747;
  assign n20752 = n20373 & ~n41282;
  assign n20753 = ~n41282 & ~n20752;
  assign n20754 = ~n20373 & ~n41282;
  assign n20755 = n20373 & ~n20752;
  assign n20756 = n20373 & n41282;
  assign n20757 = ~n20373 & n41282;
  assign n20758 = ~n20752 & ~n20757;
  assign n20759 = ~n41283 & ~n41284;
  assign n20760 = ~n41209 & n41285;
  assign n20761 = n41209 & ~n41285;
  assign n20762 = n41209 & n41285;
  assign n20763 = ~n41209 & ~n41285;
  assign n20764 = ~n20762 & ~n20763;
  assign n20765 = ~n20760 & ~n20761;
  assign n20766 = n20330 & ~n41286;
  assign n20767 = ~n20330 & n41286;
  assign n20768 = n20330 & ~n20766;
  assign n20769 = ~n41286 & ~n20766;
  assign n20770 = ~n20768 & ~n20769;
  assign n20771 = ~n20766 & ~n20767;
  assign n20772 = ~n20236 & ~n20244;
  assign n20773 = n269 & n15049;
  assign n20774 = pi120  & n37475;
  assign n20775 = pi122  & n536;
  assign n20776 = pi121  & n538;
  assign n20777 = ~n20775 & ~n20776;
  assign n20778 = ~n20774 & ~n20776;
  assign n20779 = ~n20775 & n20778;
  assign n20780 = ~n20774 & n20777;
  assign n20781 = ~n269 & n41288;
  assign n20782 = ~n15049 & n41288;
  assign n20783 = ~n20781 & ~n20782;
  assign n20784 = ~n20773 & n41288;
  assign n20785 = pi11  & ~n41289;
  assign n20786 = ~pi11  & n41289;
  assign n20787 = ~n20785 & ~n20786;
  assign n20788 = ~n20772 & ~n20787;
  assign n20789 = n20772 & n20787;
  assign n20790 = ~n20772 & ~n20788;
  assign n20791 = ~n20772 & n20787;
  assign n20792 = ~n20787 & ~n20788;
  assign n20793 = n20772 & ~n20787;
  assign n20794 = ~n41290 & ~n41291;
  assign n20795 = ~n20788 & ~n20789;
  assign n20796 = ~n41287 & ~n41292;
  assign n20797 = n41287 & n41292;
  assign n20798 = ~n41287 & ~n20796;
  assign n20799 = ~n41287 & n41292;
  assign n20800 = ~n41292 & ~n20796;
  assign n20801 = n41287 & ~n41292;
  assign n20802 = ~n41293 & ~n41294;
  assign n20803 = ~n20796 & ~n20797;
  assign n20804 = n13010 & n15068;
  assign n20805 = pi123  & n39810;
  assign n20806 = pi125  & n13040;
  assign n20807 = pi124  & n13042;
  assign n20808 = ~n20806 & ~n20807;
  assign n20809 = ~n20805 & ~n20807;
  assign n20810 = ~n20806 & n20809;
  assign n20811 = ~n20805 & n20808;
  assign n20812 = ~n13010 & n41296;
  assign n20813 = ~n15068 & n41296;
  assign n20814 = ~n20812 & ~n20813;
  assign n20815 = ~n20804 & n41296;
  assign n20816 = pi8  & ~n41297;
  assign n20817 = ~pi8  & n41297;
  assign n20818 = ~n20816 & ~n20817;
  assign n20819 = ~n19818 & n41185;
  assign n20820 = ~n19818 & ~n20252;
  assign n20821 = ~n19817 & ~n20819;
  assign n20822 = ~n20818 & ~n41298;
  assign n20823 = n20818 & n41298;
  assign n20824 = ~n41298 & ~n20822;
  assign n20825 = n20818 & ~n41298;
  assign n20826 = ~n20818 & ~n20822;
  assign n20827 = ~n20818 & n41298;
  assign n20828 = ~n41299 & ~n41300;
  assign n20829 = ~n20822 & ~n20823;
  assign n20830 = ~n41295 & ~n41301;
  assign n20831 = n41295 & n41301;
  assign n20832 = ~n41295 & ~n20830;
  assign n20833 = ~n41301 & ~n20830;
  assign n20834 = ~n20832 & ~n20833;
  assign n20835 = ~n20830 & ~n20831;
  assign n20836 = ~n19793 & ~n20260;
  assign n20837 = n14944 & n40891;
  assign n20838 = pi126  & n40177;
  assign n20839 = pi127  & n14976;
  assign n20840 = ~n20838 & ~n20839;
  assign n20841 = ~n14944 & n20840;
  assign n20842 = ~n40891 & n20840;
  assign n20843 = ~n20841 & ~n20842;
  assign n20844 = ~n20837 & n20840;
  assign n20845 = pi5  & ~n41303;
  assign n20846 = ~pi5  & n41303;
  assign n20847 = ~n20845 & ~n20846;
  assign n20848 = ~n20836 & ~n20847;
  assign n20849 = n20836 & n20847;
  assign n20850 = ~n20836 & ~n20848;
  assign n20851 = ~n20836 & n20847;
  assign n20852 = ~n20847 & ~n20848;
  assign n20853 = n20836 & ~n20847;
  assign n20854 = ~n41304 & ~n41305;
  assign n20855 = ~n20848 & ~n20849;
  assign n20856 = ~n41302 & ~n41306;
  assign n20857 = n41302 & ~n41305;
  assign n20858 = ~n41304 & n20857;
  assign n20859 = n41302 & ~n41304;
  assign n20860 = ~n41305 & n20859;
  assign n20861 = n41302 & n41306;
  assign n20862 = ~n20856 & ~n41307;
  assign n20863 = ~n20311 & n20862;
  assign n20864 = n20311 & ~n20862;
  assign n20865 = ~n20311 & ~n20863;
  assign n20866 = n20862 & ~n20863;
  assign n20867 = ~n20865 & ~n20866;
  assign n20868 = ~n20863 & ~n20864;
  assign n20869 = ~n20310 & ~n41308;
  assign n20870 = n20310 & ~n20866;
  assign n20871 = ~n20865 & n20870;
  assign n20872 = n20310 & n41308;
  assign po67  = ~n20869 & ~n41309;
  assign n20874 = ~n20863 & ~n20869;
  assign n20875 = ~n20848 & ~n20856;
  assign n20876 = n269 & n14961;
  assign n20877 = pi121  & n37475;
  assign n20878 = pi123  & n536;
  assign n20879 = pi122  & n538;
  assign n20880 = ~n20878 & ~n20879;
  assign n20881 = ~n20877 & ~n20879;
  assign n20882 = ~n20878 & n20881;
  assign n20883 = ~n20877 & n20880;
  assign n20884 = ~n20876 & n41310;
  assign n20885 = pi11  & ~n20884;
  assign n20886 = pi11  & ~n20885;
  assign n20887 = pi11  & n20884;
  assign n20888 = ~n20884 & ~n20885;
  assign n20889 = ~pi11  & ~n20884;
  assign n20890 = ~n41311 & ~n41312;
  assign n20891 = ~n20329 & ~n20766;
  assign n20892 = n20890 & n20891;
  assign n20893 = ~n20890 & ~n20891;
  assign n20894 = ~n20892 & ~n20893;
  assign n20895 = n563 & n14913;
  assign n20896 = pi118  & n37482;
  assign n20897 = pi120  & n578;
  assign n20898 = pi119  & n580;
  assign n20899 = ~n20897 & ~n20898;
  assign n20900 = ~n20896 & ~n20898;
  assign n20901 = ~n20897 & n20900;
  assign n20902 = ~n20896 & n20899;
  assign n20903 = ~n20895 & n41313;
  assign n20904 = pi14  & ~n20903;
  assign n20905 = pi14  & ~n20904;
  assign n20906 = pi14  & n20903;
  assign n20907 = ~n20903 & ~n20904;
  assign n20908 = ~pi14  & ~n20903;
  assign n20909 = ~n41314 & ~n41315;
  assign n20910 = ~n20347 & ~n20760;
  assign n20911 = ~n20909 & ~n20910;
  assign n20912 = n20909 & n20910;
  assign n20913 = ~n20909 & ~n20911;
  assign n20914 = ~n20909 & n20910;
  assign n20915 = ~n20910 & ~n20911;
  assign n20916 = n20909 & ~n20910;
  assign n20917 = ~n41316 & ~n41317;
  assign n20918 = ~n20911 & ~n20912;
  assign n20919 = n8175 & n13079;
  assign n20920 = pi115  & n38895;
  assign n20921 = pi117  & n8190;
  assign n20922 = pi116  & n8192;
  assign n20923 = ~n20921 & ~n20922;
  assign n20924 = ~n20920 & ~n20922;
  assign n20925 = ~n20921 & n20924;
  assign n20926 = ~n20920 & n20923;
  assign n20927 = ~n8175 & n41319;
  assign n20928 = ~n13079 & n41319;
  assign n20929 = ~n20927 & ~n20928;
  assign n20930 = ~n20919 & n41319;
  assign n20931 = pi17  & ~n41320;
  assign n20932 = ~pi17  & n41320;
  assign n20933 = ~n20931 & ~n20932;
  assign n20934 = ~n20372 & n41282;
  assign n20935 = ~n20372 & ~n20752;
  assign n20936 = ~n20371 & ~n20934;
  assign n20937 = ~n20933 & ~n41321;
  assign n20938 = n20933 & n41321;
  assign n20939 = ~n20937 & ~n20938;
  assign n20940 = n565 & n5576;
  assign n20941 = pi109  & n38406;
  assign n20942 = pi111  & n5591;
  assign n20943 = pi110  & n5593;
  assign n20944 = ~n20942 & ~n20943;
  assign n20945 = ~n20941 & ~n20943;
  assign n20946 = ~n20942 & n20945;
  assign n20947 = ~n20941 & n20944;
  assign n20948 = ~n20940 & n41322;
  assign n20949 = pi23  & ~n20948;
  assign n20950 = pi23  & ~n20949;
  assign n20951 = pi23  & n20948;
  assign n20952 = ~n20948 & ~n20949;
  assign n20953 = ~pi23  & ~n20948;
  assign n20954 = ~n41323 & ~n41324;
  assign n20955 = ~n20391 & ~n20716;
  assign n20956 = n20954 & n20955;
  assign n20957 = ~n20954 & ~n20955;
  assign n20958 = ~n20956 & ~n20957;
  assign n20959 = ~n20702 & ~n20710;
  assign n20960 = n4492 & n9277;
  assign n20961 = pi106  & n38208;
  assign n20962 = pi108  & n4507;
  assign n20963 = pi107  & n4509;
  assign n20964 = ~n20962 & ~n20963;
  assign n20965 = ~n20961 & ~n20963;
  assign n20966 = ~n20962 & n20965;
  assign n20967 = ~n20961 & n20964;
  assign n20968 = ~n4492 & n41325;
  assign n20969 = ~n9277 & n41325;
  assign n20970 = ~n20968 & ~n20969;
  assign n20971 = ~n20960 & n41325;
  assign n20972 = pi26  & ~n41326;
  assign n20973 = ~pi26  & n41326;
  assign n20974 = ~n20972 & ~n20973;
  assign n20975 = ~n20959 & ~n20974;
  assign n20976 = n20959 & n20974;
  assign n20977 = ~n20959 & ~n20975;
  assign n20978 = ~n20959 & n20974;
  assign n20979 = ~n20974 & ~n20975;
  assign n20980 = n20959 & ~n20974;
  assign n20981 = ~n41327 & ~n41328;
  assign n20982 = ~n20975 & ~n20976;
  assign n20983 = n607 & n8229;
  assign n20984 = pi103  & n37489;
  assign n20985 = pi105  & n620;
  assign n20986 = pi104  & n622;
  assign n20987 = ~n20985 & ~n20986;
  assign n20988 = ~n20984 & ~n20986;
  assign n20989 = ~n20985 & n20988;
  assign n20990 = ~n20984 & n20987;
  assign n20991 = ~n20983 & n41330;
  assign n20992 = pi29  & ~n20991;
  assign n20993 = pi29  & ~n20992;
  assign n20994 = pi29  & n20991;
  assign n20995 = ~n20991 & ~n20992;
  assign n20996 = ~pi29  & ~n20991;
  assign n20997 = ~n41331 & ~n41332;
  assign n20998 = ~n20411 & ~n20684;
  assign n20999 = n20997 & n20998;
  assign n21000 = ~n20997 & ~n20998;
  assign n21001 = ~n20999 & ~n21000;
  assign n21002 = n649 & n6819;
  assign n21003 = pi100  & n37496;
  assign n21004 = pi102  & n662;
  assign n21005 = pi101  & n664;
  assign n21006 = ~n21004 & ~n21005;
  assign n21007 = ~n21003 & ~n21005;
  assign n21008 = ~n21004 & n21007;
  assign n21009 = ~n21003 & n21006;
  assign n21010 = ~n649 & n41333;
  assign n21011 = ~n6819 & n41333;
  assign n21012 = ~n21010 & ~n21011;
  assign n21013 = ~n21002 & n41333;
  assign n21014 = pi32  & ~n41334;
  assign n21015 = ~pi32  & n41334;
  assign n21016 = ~n21014 & ~n21015;
  assign n21017 = n20428 & ~n20671;
  assign n21018 = ~n20671 & ~n20678;
  assign n21019 = ~n20672 & ~n21017;
  assign n21020 = ~n21016 & ~n41335;
  assign n21021 = n21016 & n41335;
  assign n21022 = ~n21020 & ~n21021;
  assign n21023 = ~n20623 & ~n20640;
  assign n21024 = ~n20624 & ~n20642;
  assign n21025 = ~n20624 & ~n21023;
  assign n21026 = ~n20608 & ~n20614;
  assign n21027 = ~n20531 & ~n20547;
  assign n21028 = ~n20530 & ~n20549;
  assign n21029 = ~n20530 & ~n21027;
  assign n21030 = n1971 & n2154;
  assign n21031 = pi79  & n37864;
  assign n21032 = pi81  & n1973;
  assign n21033 = pi80  & n1981;
  assign n21034 = ~n21032 & ~n21033;
  assign n21035 = ~n21031 & ~n21033;
  assign n21036 = ~n21032 & n21035;
  assign n21037 = ~n21031 & n21034;
  assign n21038 = ~n21030 & n41338;
  assign n21039 = pi53  & ~n21038;
  assign n21040 = pi53  & ~n21039;
  assign n21041 = pi53  & n21038;
  assign n21042 = ~n21038 & ~n21039;
  assign n21043 = ~pi53  & ~n21038;
  assign n21044 = ~n41339 & ~n41340;
  assign n21045 = ~n20509 & ~n20527;
  assign n21046 = ~n20465 & ~n20473;
  assign n21047 = n1124 & n12674;
  assign n21048 = pi70  & n40107;
  assign n21049 = pi72  & n12676;
  assign n21050 = pi71  & n12684;
  assign n21051 = ~n21049 & ~n21050;
  assign n21052 = ~n21048 & ~n21050;
  assign n21053 = ~n21049 & n21052;
  assign n21054 = ~n21048 & n21051;
  assign n21055 = ~n21047 & n41341;
  assign n21056 = pi62  & ~n21055;
  assign n21057 = pi62  & ~n21056;
  assign n21058 = pi62  & n21055;
  assign n21059 = ~n21055 & ~n21056;
  assign n21060 = ~pi62  & ~n21055;
  assign n21061 = ~n41342 & ~n41343;
  assign n21062 = pi69  & ~n40814;
  assign n21063 = pi68  & n18285;
  assign n21064 = ~n21062 & ~n21063;
  assign n21065 = pi2  & ~n21064;
  assign n21066 = ~pi2  & n21064;
  assign n21067 = pi2  & ~n21065;
  assign n21068 = pi2  & n21064;
  assign n21069 = ~n21064 & ~n21065;
  assign n21070 = ~pi2  & ~n21064;
  assign n21071 = ~n41344 & ~n41345;
  assign n21072 = ~n21065 & ~n21066;
  assign n21073 = ~n21061 & ~n41346;
  assign n21074 = n21061 & n41346;
  assign n21075 = ~n21061 & ~n21073;
  assign n21076 = ~n21061 & n41346;
  assign n21077 = ~n41346 & ~n21073;
  assign n21078 = n21061 & ~n41346;
  assign n21079 = ~n41347 & ~n41348;
  assign n21080 = ~n21073 & ~n21074;
  assign n21081 = n21046 & n41349;
  assign n21082 = ~n21046 & ~n41349;
  assign n21083 = ~n21081 & ~n21082;
  assign n21084 = n720 & n7882;
  assign n21085 = pi73  & n39128;
  assign n21086 = pi75  & n7884;
  assign n21087 = pi74  & n7892;
  assign n21088 = ~n21086 & ~n21087;
  assign n21089 = ~n21085 & ~n21087;
  assign n21090 = ~n21086 & n21089;
  assign n21091 = ~n21085 & n21088;
  assign n21092 = ~n21084 & n41350;
  assign n21093 = pi59  & ~n21092;
  assign n21094 = pi59  & ~n21093;
  assign n21095 = pi59  & n21092;
  assign n21096 = ~n21092 & ~n21093;
  assign n21097 = ~pi59  & ~n21092;
  assign n21098 = ~n41351 & ~n41352;
  assign n21099 = ~n21083 & n21098;
  assign n21100 = n21083 & ~n21098;
  assign n21101 = ~n21099 & ~n21100;
  assign n21102 = ~n20482 & n20498;
  assign n21103 = ~n20482 & ~n20499;
  assign n21104 = ~n20481 & ~n21102;
  assign n21105 = n21101 & ~n41353;
  assign n21106 = ~n21101 & n41353;
  assign n21107 = ~n21105 & ~n21106;
  assign n21108 = n1578 & n4312;
  assign n21109 = pi76  & n38376;
  assign n21110 = pi78  & n4314;
  assign n21111 = pi77  & n4322;
  assign n21112 = ~n21110 & ~n21111;
  assign n21113 = ~n21109 & ~n21111;
  assign n21114 = ~n21110 & n21113;
  assign n21115 = ~n21109 & n21112;
  assign n21116 = ~n21108 & n41354;
  assign n21117 = pi56  & ~n21116;
  assign n21118 = pi56  & ~n21117;
  assign n21119 = pi56  & n21116;
  assign n21120 = ~n21116 & ~n21117;
  assign n21121 = ~pi56  & ~n21116;
  assign n21122 = ~n41355 & ~n41356;
  assign n21123 = n21107 & ~n21122;
  assign n21124 = ~n21107 & n21122;
  assign n21125 = n21107 & ~n21123;
  assign n21126 = ~n21122 & ~n21123;
  assign n21127 = ~n21125 & ~n21126;
  assign n21128 = ~n21123 & ~n21124;
  assign n21129 = ~n21045 & ~n41357;
  assign n21130 = n21045 & n41357;
  assign n21131 = ~n41357 & ~n21129;
  assign n21132 = ~n21045 & ~n21129;
  assign n21133 = ~n21131 & ~n21132;
  assign n21134 = ~n21129 & ~n21130;
  assign n21135 = ~n21044 & ~n41358;
  assign n21136 = ~n41358 & ~n21135;
  assign n21137 = n21044 & ~n41358;
  assign n21138 = ~n21044 & ~n21135;
  assign n21139 = ~n21044 & n41358;
  assign n21140 = n21044 & n41358;
  assign n21141 = ~n21135 & ~n21140;
  assign n21142 = ~n41359 & ~n41360;
  assign n21143 = n41337 & ~n41361;
  assign n21144 = ~n41337 & n41361;
  assign n21145 = ~n21143 & ~n21144;
  assign n21146 = n894 & n2591;
  assign n21147 = pi82  & n37580;
  assign n21148 = pi84  & n896;
  assign n21149 = pi83  & n904;
  assign n21150 = ~n21148 & ~n21149;
  assign n21151 = ~n21147 & ~n21149;
  assign n21152 = ~n21148 & n21151;
  assign n21153 = ~n21147 & n21150;
  assign n21154 = ~n21146 & n41362;
  assign n21155 = pi50  & ~n21154;
  assign n21156 = pi50  & ~n21155;
  assign n21157 = pi50  & n21154;
  assign n21158 = ~n21154 & ~n21155;
  assign n21159 = ~pi50  & ~n21154;
  assign n21160 = ~n41363 & ~n41364;
  assign n21161 = ~n21145 & n21160;
  assign n21162 = n21145 & ~n21160;
  assign n21163 = ~n21161 & ~n21162;
  assign n21164 = ~n20558 & n20574;
  assign n21165 = ~n20558 & ~n20575;
  assign n21166 = ~n20557 & ~n21164;
  assign n21167 = n21163 & ~n41365;
  assign n21168 = ~n21163 & n41365;
  assign n21169 = ~n21167 & ~n21168;
  assign n21170 = n636 & n785;
  assign n21171 = pi85  & n37520;
  assign n21172 = pi87  & n787;
  assign n21173 = pi86  & n795;
  assign n21174 = ~n21172 & ~n21173;
  assign n21175 = ~n21171 & ~n21173;
  assign n21176 = ~n21172 & n21175;
  assign n21177 = ~n21171 & n21174;
  assign n21178 = ~n21170 & n41366;
  assign n21179 = pi47  & ~n21178;
  assign n21180 = pi47  & ~n21179;
  assign n21181 = pi47  & n21178;
  assign n21182 = ~n21178 & ~n21179;
  assign n21183 = ~pi47  & ~n21178;
  assign n21184 = ~n41367 & ~n41368;
  assign n21185 = n21169 & ~n21184;
  assign n21186 = ~n21169 & n21184;
  assign n21187 = n21169 & ~n21185;
  assign n21188 = ~n21184 & ~n21185;
  assign n21189 = ~n21187 & ~n21188;
  assign n21190 = ~n21185 & ~n21186;
  assign n21191 = ~n20585 & n20601;
  assign n21192 = ~n20585 & ~n20603;
  assign n21193 = ~n20584 & ~n21191;
  assign n21194 = n41369 & n41370;
  assign n21195 = ~n41369 & ~n41370;
  assign n21196 = ~n21194 & ~n21195;
  assign n21197 = n940 & n3566;
  assign n21198 = pi88  & n37541;
  assign n21199 = pi90  & n953;
  assign n21200 = pi89  & n955;
  assign n21201 = ~n21199 & ~n21200;
  assign n21202 = ~n21198 & ~n21200;
  assign n21203 = ~n21199 & n21202;
  assign n21204 = ~n21198 & n21201;
  assign n21205 = ~n21197 & n41371;
  assign n21206 = pi44  & ~n21205;
  assign n21207 = pi44  & ~n21206;
  assign n21208 = pi44  & n21205;
  assign n21209 = ~n21205 & ~n21206;
  assign n21210 = ~pi44  & ~n21205;
  assign n21211 = ~n41372 & ~n41373;
  assign n21212 = ~n21196 & n21211;
  assign n21213 = n21196 & ~n21211;
  assign n21214 = n21196 & ~n21213;
  assign n21215 = ~n21211 & ~n21213;
  assign n21216 = ~n21214 & ~n21215;
  assign n21217 = ~n21212 & ~n21213;
  assign n21218 = n21026 & n41374;
  assign n21219 = ~n21026 & ~n41374;
  assign n21220 = ~n21218 & ~n21219;
  assign n21221 = n733 & n4544;
  assign n21222 = pi91  & n37510;
  assign n21223 = pi93  & n746;
  assign n21224 = pi92  & n748;
  assign n21225 = ~n21223 & ~n21224;
  assign n21226 = ~n21222 & ~n21224;
  assign n21227 = ~n21223 & n21226;
  assign n21228 = ~n21222 & n21225;
  assign n21229 = ~n21221 & n41375;
  assign n21230 = pi41  & ~n21229;
  assign n21231 = pi41  & ~n21230;
  assign n21232 = pi41  & n21229;
  assign n21233 = ~n21229 & ~n21230;
  assign n21234 = ~pi41  & ~n21229;
  assign n21235 = ~n41376 & ~n41377;
  assign n21236 = n21220 & ~n21235;
  assign n21237 = ~n21220 & n21235;
  assign n21238 = n21220 & ~n21236;
  assign n21239 = ~n21235 & ~n21236;
  assign n21240 = ~n21238 & ~n21239;
  assign n21241 = ~n21236 & ~n21237;
  assign n21242 = n41336 & n41378;
  assign n21243 = ~n41336 & ~n41378;
  assign n21244 = ~n21242 & ~n21243;
  assign n21245 = n691 & n5281;
  assign n21246 = pi94  & n37503;
  assign n21247 = pi96  & n704;
  assign n21248 = pi95  & n706;
  assign n21249 = ~n21247 & ~n21248;
  assign n21250 = ~n21246 & ~n21248;
  assign n21251 = ~n21247 & n21250;
  assign n21252 = ~n21246 & n21249;
  assign n21253 = ~n21245 & n41379;
  assign n21254 = pi38  & ~n21253;
  assign n21255 = pi38  & ~n21254;
  assign n21256 = pi38  & n21253;
  assign n21257 = ~n21253 & ~n21254;
  assign n21258 = ~pi38  & ~n21253;
  assign n21259 = ~n41380 & ~n41381;
  assign n21260 = ~n21244 & n21259;
  assign n21261 = n21244 & ~n21259;
  assign n21262 = ~n21260 & ~n21261;
  assign n21263 = ~n20651 & ~n20669;
  assign n21264 = n21262 & ~n21263;
  assign n21265 = ~n21262 & n21263;
  assign n21266 = ~n21264 & ~n21265;
  assign n21267 = n2104 & n5578;
  assign n21268 = pi97  & n37758;
  assign n21269 = pi99  & n2117;
  assign n21270 = pi98  & n2119;
  assign n21271 = ~n21269 & ~n21270;
  assign n21272 = ~n21268 & ~n21270;
  assign n21273 = ~n21269 & n21272;
  assign n21274 = ~n21268 & n21271;
  assign n21275 = ~n21267 & n41382;
  assign n21276 = pi35  & ~n21275;
  assign n21277 = pi35  & ~n21276;
  assign n21278 = pi35  & n21275;
  assign n21279 = ~n21275 & ~n21276;
  assign n21280 = ~pi35  & ~n21275;
  assign n21281 = ~n41383 & ~n41384;
  assign n21282 = ~n21266 & n21281;
  assign n21283 = n21266 & ~n21281;
  assign n21284 = n21266 & ~n21283;
  assign n21285 = ~n21281 & ~n21283;
  assign n21286 = ~n21284 & ~n21285;
  assign n21287 = ~n21282 & ~n21283;
  assign n21288 = n21022 & ~n41385;
  assign n21289 = ~n21022 & n41385;
  assign n21290 = ~n41385 & ~n21288;
  assign n21291 = n21022 & ~n21288;
  assign n21292 = ~n21290 & ~n21291;
  assign n21293 = ~n21288 & ~n21289;
  assign n21294 = n21001 & ~n41386;
  assign n21295 = ~n21001 & n41386;
  assign n21296 = n21001 & ~n21294;
  assign n21297 = ~n41386 & ~n21294;
  assign n21298 = ~n21296 & ~n21297;
  assign n21299 = ~n21294 & ~n21295;
  assign n21300 = ~n41329 & ~n41387;
  assign n21301 = n41329 & n41387;
  assign n21302 = ~n41387 & ~n21300;
  assign n21303 = ~n41329 & ~n21300;
  assign n21304 = ~n21302 & ~n21303;
  assign n21305 = ~n21300 & ~n21301;
  assign n21306 = n20958 & ~n41388;
  assign n21307 = ~n20958 & n41388;
  assign n21308 = n20958 & ~n21306;
  assign n21309 = ~n41388 & ~n21306;
  assign n21310 = ~n21308 & ~n21309;
  assign n21311 = ~n21306 & ~n21307;
  assign n21312 = n6785 & n11258;
  assign n21313 = pi112  & n38631;
  assign n21314 = pi114  & n6800;
  assign n21315 = pi113  & n6802;
  assign n21316 = ~n21314 & ~n21315;
  assign n21317 = ~n21313 & ~n21315;
  assign n21318 = ~n21314 & n21317;
  assign n21319 = ~n21313 & n21316;
  assign n21320 = ~n21312 & n41390;
  assign n21321 = pi20  & ~n21320;
  assign n21322 = pi20  & ~n21321;
  assign n21323 = pi20  & n21320;
  assign n21324 = ~n21320 & ~n21321;
  assign n21325 = ~pi20  & ~n21320;
  assign n21326 = ~n41391 & ~n41392;
  assign n21327 = ~n20738 & ~n20746;
  assign n21328 = ~n21326 & ~n21327;
  assign n21329 = n21326 & n21327;
  assign n21330 = ~n21326 & ~n21328;
  assign n21331 = ~n21326 & n21327;
  assign n21332 = ~n21327 & ~n21328;
  assign n21333 = n21326 & ~n21327;
  assign n21334 = ~n41393 & ~n41394;
  assign n21335 = ~n21328 & ~n21329;
  assign n21336 = ~n41389 & ~n41395;
  assign n21337 = n41389 & n41395;
  assign n21338 = n41389 & ~n41395;
  assign n21339 = ~n41389 & n41395;
  assign n21340 = ~n21338 & ~n21339;
  assign n21341 = ~n21336 & ~n21337;
  assign n21342 = n20939 & ~n41396;
  assign n21343 = ~n20939 & n41396;
  assign n21344 = n20939 & ~n21342;
  assign n21345 = ~n41396 & ~n21342;
  assign n21346 = ~n21344 & ~n21345;
  assign n21347 = ~n21342 & ~n21343;
  assign n21348 = ~n41318 & ~n41397;
  assign n21349 = n41318 & n41397;
  assign n21350 = ~n41318 & n41397;
  assign n21351 = n41318 & ~n41397;
  assign n21352 = ~n21350 & ~n21351;
  assign n21353 = ~n21348 & ~n21349;
  assign n21354 = n20894 & ~n41398;
  assign n21355 = ~n20894 & n41398;
  assign n21356 = n20894 & ~n21354;
  assign n21357 = ~n41398 & ~n21354;
  assign n21358 = ~n21356 & ~n21357;
  assign n21359 = ~n21354 & ~n21355;
  assign n21360 = ~n20788 & ~n20796;
  assign n21361 = n13010 & n15021;
  assign n21362 = pi124  & n39810;
  assign n21363 = pi126  & n13040;
  assign n21364 = pi125  & n13042;
  assign n21365 = ~n21363 & ~n21364;
  assign n21366 = ~n21362 & ~n21364;
  assign n21367 = ~n21363 & n21366;
  assign n21368 = ~n21362 & n21365;
  assign n21369 = ~n13010 & n41400;
  assign n21370 = ~n15021 & n41400;
  assign n21371 = ~n21369 & ~n21370;
  assign n21372 = ~n21361 & n41400;
  assign n21373 = pi8  & ~n41401;
  assign n21374 = ~pi8  & n41401;
  assign n21375 = ~n21373 & ~n21374;
  assign n21376 = ~n21360 & ~n21375;
  assign n21377 = n21360 & n21375;
  assign n21378 = ~n21360 & ~n21376;
  assign n21379 = ~n21360 & n21375;
  assign n21380 = ~n21375 & ~n21376;
  assign n21381 = n21360 & ~n21375;
  assign n21382 = ~n41402 & ~n41403;
  assign n21383 = ~n21376 & ~n21377;
  assign n21384 = ~n41399 & ~n41404;
  assign n21385 = n41399 & ~n41403;
  assign n21386 = ~n41402 & n21385;
  assign n21387 = n41399 & ~n41402;
  assign n21388 = ~n41403 & n21387;
  assign n21389 = n41399 & n41404;
  assign n21390 = ~n21384 & ~n41405;
  assign n21391 = ~n20822 & ~n20830;
  assign n21392 = n14944 & ~n18675;
  assign n21393 = ~n40177 & ~n21392;
  assign n21394 = pi127  & n40177;
  assign n21395 = n14944 & n18680;
  assign n21396 = ~n21394 & ~n21395;
  assign n21397 = pi127  & ~n21393;
  assign n21398 = pi5  & ~n41406;
  assign n21399 = pi5  & ~n21398;
  assign n21400 = pi5  & n41406;
  assign n21401 = ~n41406 & ~n21398;
  assign n21402 = ~pi5  & ~n41406;
  assign n21403 = ~n41407 & ~n41408;
  assign n21404 = ~n21391 & ~n21403;
  assign n21405 = n21391 & n21403;
  assign n21406 = ~n21391 & ~n21404;
  assign n21407 = ~n21403 & ~n21404;
  assign n21408 = ~n21406 & ~n21407;
  assign n21409 = ~n21404 & ~n21405;
  assign n21410 = n21390 & ~n41409;
  assign n21411 = ~n21390 & n41409;
  assign n21412 = ~n21410 & ~n21411;
  assign n21413 = ~n20875 & n21412;
  assign n21414 = n20875 & ~n21412;
  assign n21415 = ~n20875 & ~n21413;
  assign n21416 = n21412 & ~n21413;
  assign n21417 = ~n21415 & ~n21416;
  assign n21418 = ~n21413 & ~n21414;
  assign n21419 = ~n20874 & ~n41410;
  assign n21420 = n20874 & ~n21416;
  assign n21421 = ~n21415 & n21420;
  assign n21422 = n20874 & n41410;
  assign po68  = ~n21419 & ~n41411;
  assign n21424 = ~n21413 & ~n21419;
  assign n21425 = ~n21404 & ~n21410;
  assign n21426 = ~n21376 & ~n21384;
  assign n21427 = n13010 & n40885;
  assign n21428 = pi125  & n39810;
  assign n21429 = pi127  & n13040;
  assign n21430 = pi126  & n13042;
  assign n21431 = ~n21429 & ~n21430;
  assign n21432 = ~n21428 & ~n21430;
  assign n21433 = ~n21429 & n21432;
  assign n21434 = ~n21428 & n21431;
  assign n21435 = ~n21427 & n41412;
  assign n21436 = pi8  & ~n21435;
  assign n21437 = pi8  & ~n21436;
  assign n21438 = pi8  & n21435;
  assign n21439 = ~n21435 & ~n21436;
  assign n21440 = ~pi8  & ~n21435;
  assign n21441 = ~n41413 & ~n41414;
  assign n21442 = ~n21426 & ~n21441;
  assign n21443 = n21426 & n21441;
  assign n21444 = ~n21426 & ~n21442;
  assign n21445 = ~n21426 & n21441;
  assign n21446 = ~n21441 & ~n21442;
  assign n21447 = n21426 & ~n21441;
  assign n21448 = ~n41415 & ~n41416;
  assign n21449 = ~n21442 & ~n21443;
  assign n21450 = n269 & n15111;
  assign n21451 = pi122  & n37475;
  assign n21452 = pi124  & n536;
  assign n21453 = pi123  & n538;
  assign n21454 = ~n21452 & ~n21453;
  assign n21455 = ~n21451 & ~n21453;
  assign n21456 = ~n21452 & n21455;
  assign n21457 = ~n21451 & n21454;
  assign n21458 = ~n21450 & n41418;
  assign n21459 = pi11  & ~n21458;
  assign n21460 = pi11  & ~n21459;
  assign n21461 = pi11  & n21458;
  assign n21462 = ~n21458 & ~n21459;
  assign n21463 = ~pi11  & ~n21458;
  assign n21464 = ~n41419 & ~n41420;
  assign n21465 = ~n20893 & ~n21354;
  assign n21466 = n21464 & n21465;
  assign n21467 = ~n21464 & ~n21465;
  assign n21468 = ~n21466 & ~n21467;
  assign n21469 = n563 & n15091;
  assign n21470 = pi119  & n37482;
  assign n21471 = pi121  & n578;
  assign n21472 = pi120  & n580;
  assign n21473 = ~n21471 & ~n21472;
  assign n21474 = ~n21470 & ~n21472;
  assign n21475 = ~n21471 & n21474;
  assign n21476 = ~n21470 & n21473;
  assign n21477 = ~n21469 & n41421;
  assign n21478 = pi14  & ~n21477;
  assign n21479 = pi14  & ~n21478;
  assign n21480 = pi14  & n21477;
  assign n21481 = ~n21477 & ~n21478;
  assign n21482 = ~pi14  & ~n21477;
  assign n21483 = ~n41422 & ~n41423;
  assign n21484 = ~n20911 & ~n21348;
  assign n21485 = ~n21483 & ~n21484;
  assign n21486 = n21483 & n21484;
  assign n21487 = ~n21485 & ~n21486;
  assign n21488 = n8175 & n13057;
  assign n21489 = pi116  & n38895;
  assign n21490 = pi118  & n8190;
  assign n21491 = pi117  & n8192;
  assign n21492 = ~n21490 & ~n21491;
  assign n21493 = ~n21489 & ~n21491;
  assign n21494 = ~n21490 & n21493;
  assign n21495 = ~n21489 & n21492;
  assign n21496 = ~n21488 & n41424;
  assign n21497 = pi17  & ~n21496;
  assign n21498 = pi17  & ~n21497;
  assign n21499 = pi17  & n21496;
  assign n21500 = ~n21496 & ~n21497;
  assign n21501 = ~pi17  & ~n21496;
  assign n21502 = ~n41425 & ~n41426;
  assign n21503 = ~n20937 & n41396;
  assign n21504 = ~n20937 & ~n21342;
  assign n21505 = ~n20938 & ~n21503;
  assign n21506 = ~n21502 & ~n41427;
  assign n21507 = n21502 & n41427;
  assign n21508 = ~n41427 & ~n21506;
  assign n21509 = n21502 & ~n41427;
  assign n21510 = ~n21502 & ~n21506;
  assign n21511 = ~n21502 & n41427;
  assign n21512 = ~n41428 & ~n41429;
  assign n21513 = ~n21506 & ~n21507;
  assign n21514 = n523 & n6785;
  assign n21515 = pi113  & n38631;
  assign n21516 = pi115  & n6800;
  assign n21517 = pi114  & n6802;
  assign n21518 = ~n21516 & ~n21517;
  assign n21519 = ~n21515 & ~n21517;
  assign n21520 = ~n21516 & n21519;
  assign n21521 = ~n21515 & n21518;
  assign n21522 = ~n21514 & n41431;
  assign n21523 = pi20  & ~n21522;
  assign n21524 = pi20  & ~n21523;
  assign n21525 = pi20  & n21522;
  assign n21526 = ~n21522 & ~n21523;
  assign n21527 = ~pi20  & ~n21522;
  assign n21528 = ~n41432 & ~n41433;
  assign n21529 = ~n21328 & ~n21336;
  assign n21530 = ~n21528 & ~n21529;
  assign n21531 = n21528 & n21529;
  assign n21532 = ~n21530 & ~n21531;
  assign n21533 = n5576 & n10844;
  assign n21534 = pi110  & n38406;
  assign n21535 = pi112  & n5591;
  assign n21536 = pi111  & n5593;
  assign n21537 = ~n21535 & ~n21536;
  assign n21538 = ~n21534 & ~n21536;
  assign n21539 = ~n21535 & n21538;
  assign n21540 = ~n21534 & n21537;
  assign n21541 = ~n21533 & n41434;
  assign n21542 = pi23  & ~n21541;
  assign n21543 = pi23  & ~n21542;
  assign n21544 = pi23  & n21541;
  assign n21545 = ~n21541 & ~n21542;
  assign n21546 = ~pi23  & ~n21541;
  assign n21547 = ~n41435 & ~n41436;
  assign n21548 = ~n20957 & ~n21306;
  assign n21549 = n21547 & n21548;
  assign n21550 = ~n21547 & ~n21548;
  assign n21551 = ~n21549 & ~n21550;
  assign n21552 = n607 & n8209;
  assign n21553 = pi104  & n37489;
  assign n21554 = pi106  & n620;
  assign n21555 = pi105  & n622;
  assign n21556 = ~n21554 & ~n21555;
  assign n21557 = ~n21553 & ~n21555;
  assign n21558 = ~n21554 & n21557;
  assign n21559 = ~n21553 & n21556;
  assign n21560 = ~n21552 & n41437;
  assign n21561 = pi29  & ~n21560;
  assign n21562 = pi29  & ~n21561;
  assign n21563 = pi29  & n21560;
  assign n21564 = ~n21560 & ~n21561;
  assign n21565 = ~pi29  & ~n21560;
  assign n21566 = ~n41438 & ~n41439;
  assign n21567 = ~n21000 & n41386;
  assign n21568 = ~n21000 & ~n21294;
  assign n21569 = ~n20999 & ~n21567;
  assign n21570 = n21566 & n41440;
  assign n21571 = ~n21566 & ~n41440;
  assign n21572 = ~n21570 & ~n21571;
  assign n21573 = n2104 & n6474;
  assign n21574 = pi98  & n37758;
  assign n21575 = pi100  & n2117;
  assign n21576 = pi99  & n2119;
  assign n21577 = ~n21575 & ~n21576;
  assign n21578 = ~n21574 & ~n21576;
  assign n21579 = ~n21575 & n21578;
  assign n21580 = ~n21574 & n21577;
  assign n21581 = ~n21573 & n41441;
  assign n21582 = pi35  & ~n21581;
  assign n21583 = pi35  & ~n21582;
  assign n21584 = pi35  & n21581;
  assign n21585 = ~n21581 & ~n21582;
  assign n21586 = ~pi35  & ~n21581;
  assign n21587 = ~n41442 & ~n41443;
  assign n21588 = ~n21243 & ~n21261;
  assign n21589 = n691 & n5630;
  assign n21590 = pi95  & n37503;
  assign n21591 = pi97  & n704;
  assign n21592 = pi96  & n706;
  assign n21593 = ~n21591 & ~n21592;
  assign n21594 = ~n21590 & ~n21592;
  assign n21595 = ~n21591 & n21594;
  assign n21596 = ~n21590 & n21593;
  assign n21597 = ~n21589 & n41444;
  assign n21598 = pi38  & ~n21597;
  assign n21599 = pi38  & ~n21598;
  assign n21600 = pi38  & n21597;
  assign n21601 = ~n21597 & ~n21598;
  assign n21602 = ~pi38  & ~n21597;
  assign n21603 = ~n41445 & ~n41446;
  assign n21604 = n785 & n3354;
  assign n21605 = pi86  & n37520;
  assign n21606 = pi88  & n787;
  assign n21607 = pi87  & n795;
  assign n21608 = ~n21606 & ~n21607;
  assign n21609 = ~n21605 & ~n21607;
  assign n21610 = ~n21606 & n21609;
  assign n21611 = ~n21605 & n21608;
  assign n21612 = ~n21604 & n41447;
  assign n21613 = pi47  & ~n21612;
  assign n21614 = pi47  & ~n21613;
  assign n21615 = pi47  & n21612;
  assign n21616 = ~n21612 & ~n21613;
  assign n21617 = ~pi47  & ~n21612;
  assign n21618 = ~n41448 & ~n41449;
  assign n21619 = ~n21144 & ~n21162;
  assign n21620 = n678 & n4312;
  assign n21621 = pi77  & n38376;
  assign n21622 = pi79  & n4314;
  assign n21623 = pi78  & n4322;
  assign n21624 = ~n21622 & ~n21623;
  assign n21625 = ~n21621 & ~n21623;
  assign n21626 = ~n21622 & n21625;
  assign n21627 = ~n21621 & n21624;
  assign n21628 = ~n21620 & n41450;
  assign n21629 = pi56  & ~n21628;
  assign n21630 = pi56  & ~n21629;
  assign n21631 = pi56  & n21628;
  assign n21632 = ~n21628 & ~n21629;
  assign n21633 = ~pi56  & ~n21628;
  assign n21634 = ~n41451 & ~n41452;
  assign n21635 = ~n21082 & ~n21100;
  assign n21636 = n1465 & n7882;
  assign n21637 = pi74  & n39128;
  assign n21638 = pi76  & n7884;
  assign n21639 = pi75  & n7892;
  assign n21640 = ~n21638 & ~n21639;
  assign n21641 = ~n21637 & ~n21639;
  assign n21642 = ~n21638 & n21641;
  assign n21643 = ~n21637 & n21640;
  assign n21644 = ~n21636 & n41453;
  assign n21645 = pi59  & ~n21644;
  assign n21646 = pi59  & ~n21645;
  assign n21647 = pi59  & n21644;
  assign n21648 = ~n21644 & ~n21645;
  assign n21649 = ~pi59  & ~n21644;
  assign n21650 = ~n41454 & ~n41455;
  assign n21651 = ~n21065 & ~n21073;
  assign n21652 = ~pi2  & ~pi5 ;
  assign n21653 = pi2  & pi5 ;
  assign n21654 = pi2  & ~pi5 ;
  assign n21655 = ~pi2  & pi5 ;
  assign n21656 = ~n21654 & ~n21655;
  assign n21657 = ~n21652 & ~n21653;
  assign n21658 = pi70  & ~n40814;
  assign n21659 = pi69  & n18285;
  assign n21660 = ~n21658 & ~n21659;
  assign n21661 = ~n41456 & ~n21660;
  assign n21662 = n41456 & n21660;
  assign n21663 = ~n21661 & ~n21662;
  assign n21664 = n21651 & ~n21663;
  assign n21665 = ~n21651 & n21663;
  assign n21666 = ~n21664 & ~n21665;
  assign n21667 = n1238 & n12674;
  assign n21668 = pi71  & n40107;
  assign n21669 = pi73  & n12676;
  assign n21670 = pi72  & n12684;
  assign n21671 = ~n21669 & ~n21670;
  assign n21672 = ~n21668 & ~n21670;
  assign n21673 = ~n21669 & n21672;
  assign n21674 = ~n21668 & n21671;
  assign n21675 = ~n21667 & n41457;
  assign n21676 = pi62  & ~n21675;
  assign n21677 = pi62  & ~n21676;
  assign n21678 = pi62  & n21675;
  assign n21679 = ~n21675 & ~n21676;
  assign n21680 = ~pi62  & ~n21675;
  assign n21681 = ~n41458 & ~n41459;
  assign n21682 = ~n21666 & n21681;
  assign n21683 = n21666 & ~n21681;
  assign n21684 = ~n21682 & ~n21683;
  assign n21685 = ~n21650 & n21684;
  assign n21686 = n21650 & ~n21684;
  assign n21687 = ~n21650 & ~n21685;
  assign n21688 = ~n21650 & ~n21684;
  assign n21689 = n21684 & ~n21685;
  assign n21690 = n21650 & n21684;
  assign n21691 = ~n41460 & ~n41461;
  assign n21692 = ~n21685 & ~n21686;
  assign n21693 = ~n21635 & ~n41462;
  assign n21694 = n21635 & n41462;
  assign n21695 = ~n21635 & ~n21693;
  assign n21696 = ~n41462 & ~n21693;
  assign n21697 = ~n21695 & ~n21696;
  assign n21698 = ~n21693 & ~n21694;
  assign n21699 = ~n21634 & ~n41463;
  assign n21700 = n21634 & n41463;
  assign n21701 = ~n41463 & ~n21699;
  assign n21702 = n21634 & ~n41463;
  assign n21703 = ~n21634 & ~n21699;
  assign n21704 = ~n21634 & n41463;
  assign n21705 = ~n41464 & ~n41465;
  assign n21706 = ~n21699 & ~n21700;
  assign n21707 = ~n21105 & n21122;
  assign n21708 = ~n21105 & ~n21123;
  assign n21709 = ~n21106 & ~n21707;
  assign n21710 = n41466 & n41467;
  assign n21711 = ~n41466 & ~n41467;
  assign n21712 = ~n21710 & ~n21711;
  assign n21713 = n1971 & n2134;
  assign n21714 = pi80  & n37864;
  assign n21715 = pi82  & n1973;
  assign n21716 = pi81  & n1981;
  assign n21717 = ~n21715 & ~n21716;
  assign n21718 = ~n21714 & ~n21716;
  assign n21719 = ~n21715 & n21718;
  assign n21720 = ~n21714 & n21717;
  assign n21721 = ~n21713 & n41468;
  assign n21722 = pi53  & ~n21721;
  assign n21723 = pi53  & ~n21722;
  assign n21724 = pi53  & n21721;
  assign n21725 = ~n21721 & ~n21722;
  assign n21726 = ~pi53  & ~n21721;
  assign n21727 = ~n41469 & ~n41470;
  assign n21728 = n21712 & ~n21727;
  assign n21729 = ~n21712 & n21727;
  assign n21730 = n21712 & ~n21728;
  assign n21731 = n21712 & n21727;
  assign n21732 = ~n21727 & ~n21728;
  assign n21733 = ~n21712 & ~n21727;
  assign n21734 = ~n41471 & ~n41472;
  assign n21735 = ~n21728 & ~n21729;
  assign n21736 = n21044 & ~n21129;
  assign n21737 = ~n21129 & ~n21135;
  assign n21738 = ~n21130 & ~n21736;
  assign n21739 = n41473 & n41474;
  assign n21740 = ~n41473 & ~n41474;
  assign n21741 = ~n21739 & ~n21740;
  assign n21742 = n894 & n2804;
  assign n21743 = pi83  & n37580;
  assign n21744 = pi85  & n896;
  assign n21745 = pi84  & n904;
  assign n21746 = ~n21744 & ~n21745;
  assign n21747 = ~n21743 & ~n21745;
  assign n21748 = ~n21744 & n21747;
  assign n21749 = ~n21743 & n21746;
  assign n21750 = ~n21742 & n41475;
  assign n21751 = pi50  & ~n21750;
  assign n21752 = pi50  & ~n21751;
  assign n21753 = pi50  & n21750;
  assign n21754 = ~n21750 & ~n21751;
  assign n21755 = ~pi50  & ~n21750;
  assign n21756 = ~n41476 & ~n41477;
  assign n21757 = n21741 & ~n21756;
  assign n21758 = ~n21741 & n21756;
  assign n21759 = n21741 & ~n21757;
  assign n21760 = n21741 & n21756;
  assign n21761 = ~n21756 & ~n21757;
  assign n21762 = ~n21741 & ~n21756;
  assign n21763 = ~n41478 & ~n41479;
  assign n21764 = ~n21757 & ~n21758;
  assign n21765 = ~n21619 & ~n41480;
  assign n21766 = n21619 & n41480;
  assign n21767 = ~n21619 & n41480;
  assign n21768 = n21619 & ~n41480;
  assign n21769 = ~n21767 & ~n21768;
  assign n21770 = ~n21765 & ~n21766;
  assign n21771 = ~n21618 & ~n41481;
  assign n21772 = n21618 & n41481;
  assign n21773 = ~n21771 & ~n21772;
  assign n21774 = ~n21167 & n21184;
  assign n21775 = ~n21167 & ~n21185;
  assign n21776 = ~n21168 & ~n21774;
  assign n21777 = ~n21773 & n41482;
  assign n21778 = n21773 & ~n41482;
  assign n21779 = ~n21777 & ~n21778;
  assign n21780 = n594 & n940;
  assign n21781 = pi89  & n37541;
  assign n21782 = pi91  & n953;
  assign n21783 = pi90  & n955;
  assign n21784 = ~n21782 & ~n21783;
  assign n21785 = ~n21781 & ~n21783;
  assign n21786 = ~n21782 & n21785;
  assign n21787 = ~n21781 & n21784;
  assign n21788 = ~n21780 & n41483;
  assign n21789 = pi44  & ~n21788;
  assign n21790 = pi44  & ~n21789;
  assign n21791 = pi44  & n21788;
  assign n21792 = ~n21788 & ~n21789;
  assign n21793 = ~pi44  & ~n21788;
  assign n21794 = ~n41484 & ~n41485;
  assign n21795 = n21779 & ~n21794;
  assign n21796 = ~n21779 & n21794;
  assign n21797 = n21779 & ~n21795;
  assign n21798 = n21779 & n21794;
  assign n21799 = ~n21794 & ~n21795;
  assign n21800 = ~n21779 & ~n21794;
  assign n21801 = ~n41486 & ~n41487;
  assign n21802 = ~n21795 & ~n21796;
  assign n21803 = ~n21195 & n21211;
  assign n21804 = ~n21195 & ~n21213;
  assign n21805 = ~n21194 & ~n21803;
  assign n21806 = n41488 & n41489;
  assign n21807 = ~n41488 & ~n41489;
  assign n21808 = ~n21806 & ~n21807;
  assign n21809 = n733 & n4524;
  assign n21810 = pi92  & n37510;
  assign n21811 = pi94  & n746;
  assign n21812 = pi93  & n748;
  assign n21813 = ~n21811 & ~n21812;
  assign n21814 = ~n21810 & ~n21812;
  assign n21815 = ~n21811 & n21814;
  assign n21816 = ~n21810 & n21813;
  assign n21817 = ~n21809 & n41490;
  assign n21818 = pi41  & ~n21817;
  assign n21819 = pi41  & ~n21818;
  assign n21820 = pi41  & n21817;
  assign n21821 = ~n21817 & ~n21818;
  assign n21822 = ~pi41  & ~n21817;
  assign n21823 = ~n41491 & ~n41492;
  assign n21824 = n21808 & ~n21823;
  assign n21825 = ~n21808 & n21823;
  assign n21826 = ~n21824 & ~n21825;
  assign n21827 = ~n21219 & n21235;
  assign n21828 = ~n21219 & ~n21236;
  assign n21829 = ~n21218 & ~n21827;
  assign n21830 = ~n21824 & n41493;
  assign n21831 = ~n21824 & ~n41493;
  assign n21832 = ~n21825 & ~n41493;
  assign n21833 = ~n21824 & n21832;
  assign n21834 = ~n21825 & n21831;
  assign n21835 = ~n21824 & ~n41494;
  assign n21836 = ~n21825 & ~n21830;
  assign n21837 = ~n21825 & n41495;
  assign n21838 = n21826 & n41493;
  assign n21839 = ~n41493 & ~n41494;
  assign n21840 = ~n21826 & ~n41493;
  assign n21841 = ~n41496 & ~n41497;
  assign n21842 = ~n21603 & ~n21841;
  assign n21843 = n21603 & n21841;
  assign n21844 = ~n21841 & ~n21842;
  assign n21845 = ~n21603 & ~n21842;
  assign n21846 = ~n21844 & ~n21845;
  assign n21847 = ~n21842 & ~n21843;
  assign n21848 = ~n21588 & ~n41498;
  assign n21849 = n21588 & n41498;
  assign n21850 = ~n21588 & n41498;
  assign n21851 = n21588 & ~n41498;
  assign n21852 = ~n21850 & ~n21851;
  assign n21853 = ~n21848 & ~n21849;
  assign n21854 = ~n21587 & ~n41499;
  assign n21855 = n21587 & n41499;
  assign n21856 = ~n21854 & ~n21855;
  assign n21857 = ~n21265 & ~n21281;
  assign n21858 = ~n21264 & ~n21283;
  assign n21859 = ~n21264 & ~n21857;
  assign n21860 = ~n21856 & n41500;
  assign n21861 = n21856 & ~n41500;
  assign n21862 = ~n21860 & ~n21861;
  assign n21863 = n649 & n6787;
  assign n21864 = pi101  & n37496;
  assign n21865 = pi103  & n662;
  assign n21866 = pi102  & n664;
  assign n21867 = ~n21865 & ~n21866;
  assign n21868 = ~n21864 & ~n21866;
  assign n21869 = ~n21865 & n21868;
  assign n21870 = ~n21864 & n21867;
  assign n21871 = ~n21863 & n41501;
  assign n21872 = pi32  & ~n21871;
  assign n21873 = pi32  & ~n21872;
  assign n21874 = pi32  & n21871;
  assign n21875 = ~n21871 & ~n21872;
  assign n21876 = ~pi32  & ~n21871;
  assign n21877 = ~n41502 & ~n41503;
  assign n21878 = ~n21020 & n41385;
  assign n21879 = ~n21020 & ~n21288;
  assign n21880 = ~n21021 & ~n21878;
  assign n21881 = n21877 & n41504;
  assign n21882 = ~n21877 & ~n41504;
  assign n21883 = ~n21881 & ~n21882;
  assign n21884 = n21862 & n21883;
  assign n21885 = ~n21862 & ~n21883;
  assign n21886 = ~n21884 & ~n21885;
  assign n21887 = n21572 & n21886;
  assign n21888 = ~n21572 & ~n21886;
  assign n21889 = ~n21887 & ~n21888;
  assign n21890 = ~n20975 & ~n21300;
  assign n21891 = n4492 & n9701;
  assign n21892 = pi107  & n38208;
  assign n21893 = pi109  & n4507;
  assign n21894 = pi108  & n4509;
  assign n21895 = ~n21893 & ~n21894;
  assign n21896 = ~n21892 & ~n21894;
  assign n21897 = ~n21893 & n21896;
  assign n21898 = ~n21892 & n21895;
  assign n21899 = ~n21891 & n41505;
  assign n21900 = pi26  & ~n21899;
  assign n21901 = pi26  & ~n21900;
  assign n21902 = pi26  & n21899;
  assign n21903 = ~n21899 & ~n21900;
  assign n21904 = ~pi26  & ~n21899;
  assign n21905 = ~n41506 & ~n41507;
  assign n21906 = ~n21890 & ~n21905;
  assign n21907 = n21890 & n21905;
  assign n21908 = ~n21890 & ~n21906;
  assign n21909 = ~n21890 & n21905;
  assign n21910 = ~n21905 & ~n21906;
  assign n21911 = n21890 & ~n21905;
  assign n21912 = ~n41508 & ~n41509;
  assign n21913 = ~n21906 & ~n21907;
  assign n21914 = n21889 & ~n41510;
  assign n21915 = ~n21889 & n41510;
  assign n21916 = ~n21889 & ~n41510;
  assign n21917 = n21889 & n41510;
  assign n21918 = ~n21916 & ~n21917;
  assign n21919 = ~n21914 & ~n21915;
  assign n21920 = n21551 & ~n41511;
  assign n21921 = ~n41511 & ~n21920;
  assign n21922 = ~n21551 & ~n41511;
  assign n21923 = n21551 & ~n21920;
  assign n21924 = n21551 & n41511;
  assign n21925 = ~n21551 & n41511;
  assign n21926 = ~n21920 & ~n21925;
  assign n21927 = ~n41512 & ~n41513;
  assign n21928 = n21532 & n41514;
  assign n21929 = ~n21532 & ~n41514;
  assign n21930 = n41514 & ~n21928;
  assign n21931 = n21532 & ~n21928;
  assign n21932 = ~n21930 & ~n21931;
  assign n21933 = ~n21928 & ~n21929;
  assign n21934 = ~n41430 & ~n41515;
  assign n21935 = n41430 & n41515;
  assign n21936 = ~n41430 & ~n21934;
  assign n21937 = ~n41515 & ~n21934;
  assign n21938 = ~n21936 & ~n21937;
  assign n21939 = ~n21934 & ~n21935;
  assign n21940 = n21487 & ~n41516;
  assign n21941 = ~n21487 & n41516;
  assign n21942 = ~n41516 & ~n21940;
  assign n21943 = n21487 & ~n21940;
  assign n21944 = ~n21942 & ~n21943;
  assign n21945 = ~n21940 & ~n21941;
  assign n21946 = n21468 & ~n41517;
  assign n21947 = ~n41517 & ~n21946;
  assign n21948 = ~n21468 & ~n41517;
  assign n21949 = n21468 & ~n21946;
  assign n21950 = n21468 & n41517;
  assign n21951 = ~n21468 & n41517;
  assign n21952 = ~n21946 & ~n21951;
  assign n21953 = ~n41518 & ~n41519;
  assign n21954 = ~n41417 & n41520;
  assign n21955 = n41417 & ~n41520;
  assign n21956 = ~n41417 & ~n41520;
  assign n21957 = n41417 & n41520;
  assign n21958 = ~n21956 & ~n21957;
  assign n21959 = ~n21954 & ~n21955;
  assign n21960 = ~n21425 & ~n41521;
  assign n21961 = n21425 & n41521;
  assign n21962 = ~n21960 & ~n21961;
  assign n21963 = ~n21424 & n21962;
  assign n21964 = n21424 & ~n21962;
  assign po69  = ~n21963 & ~n21964;
  assign n21966 = ~n21960 & ~n21963;
  assign n21967 = ~n21442 & ~n21954;
  assign n21968 = n13010 & n40891;
  assign n21969 = pi126  & n39810;
  assign n21970 = pi127  & n13042;
  assign n21971 = ~n21969 & ~n21970;
  assign n21972 = ~n13010 & n21971;
  assign n21973 = ~n40891 & n21971;
  assign n21974 = ~n21972 & ~n21973;
  assign n21975 = ~n21968 & n21971;
  assign n21976 = pi8  & ~n41522;
  assign n21977 = ~pi8  & n41522;
  assign n21978 = ~n21976 & ~n21977;
  assign n21979 = ~n21467 & n41517;
  assign n21980 = ~n21467 & ~n21946;
  assign n21981 = ~n21466 & ~n21979;
  assign n21982 = ~n21978 & ~n41523;
  assign n21983 = n21978 & n41523;
  assign n21984 = ~n21982 & ~n21983;
  assign n21985 = n269 & n15068;
  assign n21986 = pi123  & n37475;
  assign n21987 = pi125  & n536;
  assign n21988 = pi124  & n538;
  assign n21989 = ~n21987 & ~n21988;
  assign n21990 = ~n21986 & ~n21988;
  assign n21991 = ~n21987 & n21990;
  assign n21992 = ~n21986 & n21989;
  assign n21993 = ~n21985 & n41524;
  assign n21994 = pi11  & ~n21993;
  assign n21995 = pi11  & ~n21994;
  assign n21996 = pi11  & n21993;
  assign n21997 = ~n21993 & ~n21994;
  assign n21998 = ~pi11  & ~n21993;
  assign n21999 = ~n41525 & ~n41526;
  assign n22000 = ~n21485 & ~n21940;
  assign n22001 = n21999 & n22000;
  assign n22002 = ~n21999 & ~n22000;
  assign n22003 = ~n22001 & ~n22002;
  assign n22004 = ~n21506 & ~n21934;
  assign n22005 = n563 & n15049;
  assign n22006 = pi120  & n37482;
  assign n22007 = pi122  & n578;
  assign n22008 = pi121  & n580;
  assign n22009 = ~n22007 & ~n22008;
  assign n22010 = ~n22006 & ~n22008;
  assign n22011 = ~n22007 & n22010;
  assign n22012 = ~n22006 & n22009;
  assign n22013 = ~n563 & n41527;
  assign n22014 = ~n15049 & n41527;
  assign n22015 = ~n22013 & ~n22014;
  assign n22016 = ~n22005 & n41527;
  assign n22017 = pi14  & ~n41528;
  assign n22018 = ~pi14  & n41528;
  assign n22019 = ~n22017 & ~n22018;
  assign n22020 = ~n22004 & ~n22019;
  assign n22021 = n22004 & n22019;
  assign n22022 = ~n22020 & ~n22021;
  assign n22023 = n8175 & n13027;
  assign n22024 = pi117  & n38895;
  assign n22025 = pi119  & n8190;
  assign n22026 = pi118  & n8192;
  assign n22027 = ~n22025 & ~n22026;
  assign n22028 = ~n22024 & ~n22026;
  assign n22029 = ~n22025 & n22028;
  assign n22030 = ~n22024 & n22027;
  assign n22031 = ~n22023 & n41529;
  assign n22032 = pi17  & ~n22031;
  assign n22033 = pi17  & ~n22032;
  assign n22034 = pi17  & n22031;
  assign n22035 = ~n22031 & ~n22032;
  assign n22036 = ~pi17  & ~n22031;
  assign n22037 = ~n41530 & ~n41531;
  assign n22038 = ~n21530 & ~n41514;
  assign n22039 = ~n21530 & ~n21928;
  assign n22040 = ~n21531 & ~n22038;
  assign n22041 = n22037 & n41532;
  assign n22042 = ~n22037 & ~n41532;
  assign n22043 = ~n22041 & ~n22042;
  assign n22044 = n6785 & n12530;
  assign n22045 = pi114  & n38631;
  assign n22046 = pi116  & n6800;
  assign n22047 = pi115  & n6802;
  assign n22048 = ~n22046 & ~n22047;
  assign n22049 = ~n22045 & ~n22047;
  assign n22050 = ~n22046 & n22049;
  assign n22051 = ~n22045 & n22048;
  assign n22052 = ~n22044 & n41533;
  assign n22053 = pi20  & ~n22052;
  assign n22054 = pi20  & ~n22053;
  assign n22055 = pi20  & n22052;
  assign n22056 = ~n22052 & ~n22053;
  assign n22057 = ~pi20  & ~n22052;
  assign n22058 = ~n41534 & ~n41535;
  assign n22059 = ~n21550 & n41511;
  assign n22060 = ~n21550 & ~n21920;
  assign n22061 = ~n21549 & ~n22059;
  assign n22062 = n22058 & n41536;
  assign n22063 = ~n22058 & ~n41536;
  assign n22064 = ~n22062 & ~n22063;
  assign n22065 = ~n21571 & ~n21887;
  assign n22066 = n4492 & n9678;
  assign n22067 = pi108  & n38208;
  assign n22068 = pi110  & n4507;
  assign n22069 = pi109  & n4509;
  assign n22070 = ~n22068 & ~n22069;
  assign n22071 = ~n22067 & ~n22069;
  assign n22072 = ~n22068 & n22071;
  assign n22073 = ~n22067 & n22070;
  assign n22074 = ~n4492 & n41537;
  assign n22075 = ~n9678 & n41537;
  assign n22076 = ~n22074 & ~n22075;
  assign n22077 = ~n22066 & n41537;
  assign n22078 = pi26  & ~n41538;
  assign n22079 = ~pi26  & n41538;
  assign n22080 = ~n22078 & ~n22079;
  assign n22081 = ~n22065 & ~n22080;
  assign n22082 = n22065 & n22080;
  assign n22083 = ~n22081 & ~n22082;
  assign n22084 = n607 & n8177;
  assign n22085 = pi105  & n37489;
  assign n22086 = pi107  & n620;
  assign n22087 = pi106  & n622;
  assign n22088 = ~n22086 & ~n22087;
  assign n22089 = ~n22085 & ~n22087;
  assign n22090 = ~n22086 & n22089;
  assign n22091 = ~n22085 & n22088;
  assign n22092 = ~n22084 & n41539;
  assign n22093 = pi29  & ~n22092;
  assign n22094 = pi29  & ~n22093;
  assign n22095 = pi29  & n22092;
  assign n22096 = ~n22092 & ~n22093;
  assign n22097 = ~pi29  & ~n22092;
  assign n22098 = ~n41540 & ~n41541;
  assign n22099 = ~n21882 & ~n21884;
  assign n22100 = ~n22098 & ~n22099;
  assign n22101 = n22098 & n22099;
  assign n22102 = ~n22098 & ~n22100;
  assign n22103 = ~n22098 & n22099;
  assign n22104 = ~n22099 & ~n22100;
  assign n22105 = n22098 & ~n22099;
  assign n22106 = ~n41542 & ~n41543;
  assign n22107 = ~n22100 & ~n22101;
  assign n22108 = n649 & n8136;
  assign n22109 = pi102  & n37496;
  assign n22110 = pi104  & n662;
  assign n22111 = pi103  & n664;
  assign n22112 = ~n22110 & ~n22111;
  assign n22113 = ~n22109 & ~n22111;
  assign n22114 = ~n22110 & n22113;
  assign n22115 = ~n22109 & n22112;
  assign n22116 = ~n22108 & n41545;
  assign n22117 = pi32  & ~n22116;
  assign n22118 = pi32  & ~n22117;
  assign n22119 = pi32  & n22116;
  assign n22120 = ~n22116 & ~n22117;
  assign n22121 = ~pi32  & ~n22116;
  assign n22122 = ~n41546 & ~n41547;
  assign n22123 = ~n21854 & ~n21861;
  assign n22124 = n22122 & n22123;
  assign n22125 = ~n22122 & ~n22123;
  assign n22126 = ~n22124 & ~n22125;
  assign n22127 = n2104 & n6839;
  assign n22128 = pi99  & n37758;
  assign n22129 = pi101  & n2117;
  assign n22130 = pi100  & n2119;
  assign n22131 = ~n22129 & ~n22130;
  assign n22132 = ~n22128 & ~n22130;
  assign n22133 = ~n22129 & n22132;
  assign n22134 = ~n22128 & n22131;
  assign n22135 = ~n22127 & n41548;
  assign n22136 = pi35  & ~n22135;
  assign n22137 = pi35  & ~n22136;
  assign n22138 = pi35  & n22135;
  assign n22139 = ~n22135 & ~n22136;
  assign n22140 = ~pi35  & ~n22135;
  assign n22141 = ~n41549 & ~n41550;
  assign n22142 = ~n21842 & ~n21848;
  assign n22143 = n691 & n5610;
  assign n22144 = pi96  & n37503;
  assign n22145 = pi98  & n704;
  assign n22146 = pi97  & n706;
  assign n22147 = ~n22145 & ~n22146;
  assign n22148 = ~n22144 & ~n22146;
  assign n22149 = ~n22145 & n22148;
  assign n22150 = ~n22144 & n22147;
  assign n22151 = ~n22143 & n41551;
  assign n22152 = pi38  & ~n22151;
  assign n22153 = pi38  & ~n22152;
  assign n22154 = pi38  & n22151;
  assign n22155 = ~n22151 & ~n22152;
  assign n22156 = ~pi38  & ~n22151;
  assign n22157 = ~n41552 & ~n41553;
  assign n22158 = ~n21795 & ~n21807;
  assign n22159 = ~n21771 & ~n21778;
  assign n22160 = ~n21757 & ~n21765;
  assign n22161 = ~n21728 & ~n21740;
  assign n22162 = ~n21699 & ~n21711;
  assign n22163 = ~n21685 & ~n21693;
  assign n22164 = ~n21665 & ~n21683;
  assign n22165 = ~n21652 & ~n21661;
  assign n22166 = pi71  & ~n40814;
  assign n22167 = pi70  & n18285;
  assign n22168 = ~n22166 & ~n22167;
  assign n22169 = ~n22165 & n22168;
  assign n22170 = n22165 & ~n22168;
  assign n22171 = ~n22169 & ~n22170;
  assign n22172 = n1218 & n12674;
  assign n22173 = pi72  & n40107;
  assign n22174 = pi74  & n12676;
  assign n22175 = pi73  & n12684;
  assign n22176 = ~n22174 & ~n22175;
  assign n22177 = ~n22173 & ~n22175;
  assign n22178 = ~n22174 & n22177;
  assign n22179 = ~n22173 & n22176;
  assign n22180 = ~n12674 & n41554;
  assign n22181 = ~n1218 & n41554;
  assign n22182 = ~n22180 & ~n22181;
  assign n22183 = ~n22172 & n41554;
  assign n22184 = pi62  & ~n41555;
  assign n22185 = ~pi62  & n41555;
  assign n22186 = ~n22184 & ~n22185;
  assign n22187 = n22171 & ~n22186;
  assign n22188 = ~n22171 & n22186;
  assign n22189 = ~n22187 & ~n22188;
  assign n22190 = ~n22164 & n22189;
  assign n22191 = n22164 & ~n22189;
  assign n22192 = ~n22190 & ~n22191;
  assign n22193 = n1596 & n7882;
  assign n22194 = pi75  & n39128;
  assign n22195 = pi77  & n7884;
  assign n22196 = pi76  & n7892;
  assign n22197 = ~n22195 & ~n22196;
  assign n22198 = ~n22194 & ~n22196;
  assign n22199 = ~n22195 & n22198;
  assign n22200 = ~n22194 & n22197;
  assign n22201 = ~n22193 & n41556;
  assign n22202 = pi59  & ~n22201;
  assign n22203 = pi59  & ~n22202;
  assign n22204 = pi59  & n22201;
  assign n22205 = ~n22201 & ~n22202;
  assign n22206 = ~pi59  & ~n22201;
  assign n22207 = ~n41557 & ~n41558;
  assign n22208 = n22192 & ~n22207;
  assign n22209 = ~n22192 & n22207;
  assign n22210 = n22192 & ~n22208;
  assign n22211 = ~n22207 & ~n22208;
  assign n22212 = ~n22210 & ~n22211;
  assign n22213 = ~n22208 & ~n22209;
  assign n22214 = n22163 & n41559;
  assign n22215 = ~n22163 & ~n41559;
  assign n22216 = ~n22214 & ~n22215;
  assign n22217 = n2063 & n4312;
  assign n22218 = pi78  & n38376;
  assign n22219 = pi80  & n4314;
  assign n22220 = pi79  & n4322;
  assign n22221 = ~n22219 & ~n22220;
  assign n22222 = ~n22218 & ~n22220;
  assign n22223 = ~n22219 & n22222;
  assign n22224 = ~n22218 & n22221;
  assign n22225 = ~n22217 & n41560;
  assign n22226 = pi56  & ~n22225;
  assign n22227 = pi56  & ~n22226;
  assign n22228 = pi56  & n22225;
  assign n22229 = ~n22225 & ~n22226;
  assign n22230 = ~pi56  & ~n22225;
  assign n22231 = ~n41561 & ~n41562;
  assign n22232 = ~n22216 & n22231;
  assign n22233 = n22216 & ~n22231;
  assign n22234 = n22216 & ~n22233;
  assign n22235 = ~n22231 & ~n22233;
  assign n22236 = ~n22234 & ~n22235;
  assign n22237 = ~n22232 & ~n22233;
  assign n22238 = n22162 & n41563;
  assign n22239 = ~n22162 & ~n41563;
  assign n22240 = ~n22238 & ~n22239;
  assign n22241 = n1971 & n2091;
  assign n22242 = pi81  & n37864;
  assign n22243 = pi83  & n1973;
  assign n22244 = pi82  & n1981;
  assign n22245 = ~n22243 & ~n22244;
  assign n22246 = ~n22242 & ~n22244;
  assign n22247 = ~n22243 & n22246;
  assign n22248 = ~n22242 & n22245;
  assign n22249 = ~n22241 & n41564;
  assign n22250 = pi53  & ~n22249;
  assign n22251 = pi53  & ~n22250;
  assign n22252 = pi53  & n22249;
  assign n22253 = ~n22249 & ~n22250;
  assign n22254 = ~pi53  & ~n22249;
  assign n22255 = ~n41565 & ~n41566;
  assign n22256 = n22240 & ~n22255;
  assign n22257 = ~n22240 & n22255;
  assign n22258 = n22240 & ~n22256;
  assign n22259 = ~n22255 & ~n22256;
  assign n22260 = ~n22258 & ~n22259;
  assign n22261 = ~n22256 & ~n22257;
  assign n22262 = n22161 & n41567;
  assign n22263 = ~n22161 & ~n41567;
  assign n22264 = ~n22262 & ~n22263;
  assign n22265 = n894 & n2779;
  assign n22266 = pi84  & n37580;
  assign n22267 = pi86  & n896;
  assign n22268 = pi85  & n904;
  assign n22269 = ~n22267 & ~n22268;
  assign n22270 = ~n22266 & ~n22268;
  assign n22271 = ~n22267 & n22270;
  assign n22272 = ~n22266 & n22269;
  assign n22273 = ~n22265 & n41568;
  assign n22274 = pi50  & ~n22273;
  assign n22275 = pi50  & ~n22274;
  assign n22276 = pi50  & n22273;
  assign n22277 = ~n22273 & ~n22274;
  assign n22278 = ~pi50  & ~n22273;
  assign n22279 = ~n41569 & ~n41570;
  assign n22280 = ~n22264 & n22279;
  assign n22281 = n22264 & ~n22279;
  assign n22282 = n22264 & ~n22281;
  assign n22283 = ~n22279 & ~n22281;
  assign n22284 = ~n22282 & ~n22283;
  assign n22285 = ~n22280 & ~n22281;
  assign n22286 = n22160 & n41571;
  assign n22287 = ~n22160 & ~n41571;
  assign n22288 = ~n22286 & ~n22287;
  assign n22289 = n785 & n3591;
  assign n22290 = pi87  & n37520;
  assign n22291 = pi89  & n787;
  assign n22292 = pi88  & n795;
  assign n22293 = ~n22291 & ~n22292;
  assign n22294 = ~n22290 & ~n22292;
  assign n22295 = ~n22291 & n22294;
  assign n22296 = ~n22290 & n22293;
  assign n22297 = ~n22289 & n41572;
  assign n22298 = pi47  & ~n22297;
  assign n22299 = pi47  & ~n22298;
  assign n22300 = pi47  & n22297;
  assign n22301 = ~n22297 & ~n22298;
  assign n22302 = ~pi47  & ~n22297;
  assign n22303 = ~n41573 & ~n41574;
  assign n22304 = n22288 & ~n22303;
  assign n22305 = ~n22288 & n22303;
  assign n22306 = n22288 & ~n22304;
  assign n22307 = ~n22303 & ~n22304;
  assign n22308 = ~n22306 & ~n22307;
  assign n22309 = ~n22304 & ~n22305;
  assign n22310 = n22159 & n41575;
  assign n22311 = ~n22159 & ~n41575;
  assign n22312 = ~n22310 & ~n22311;
  assign n22313 = n940 & n4453;
  assign n22314 = pi90  & n37541;
  assign n22315 = pi92  & n953;
  assign n22316 = pi91  & n955;
  assign n22317 = ~n22315 & ~n22316;
  assign n22318 = ~n22314 & ~n22316;
  assign n22319 = ~n22315 & n22318;
  assign n22320 = ~n22314 & n22317;
  assign n22321 = ~n22313 & n41576;
  assign n22322 = pi44  & ~n22321;
  assign n22323 = pi44  & ~n22322;
  assign n22324 = pi44  & n22321;
  assign n22325 = ~n22321 & ~n22322;
  assign n22326 = ~pi44  & ~n22321;
  assign n22327 = ~n41577 & ~n41578;
  assign n22328 = ~n22312 & n22327;
  assign n22329 = n22312 & ~n22327;
  assign n22330 = n22312 & ~n22329;
  assign n22331 = ~n22327 & ~n22329;
  assign n22332 = ~n22330 & ~n22331;
  assign n22333 = ~n22328 & ~n22329;
  assign n22334 = n22158 & n41579;
  assign n22335 = ~n22158 & ~n41579;
  assign n22336 = ~n22334 & ~n22335;
  assign n22337 = n733 & n4494;
  assign n22338 = pi93  & n37510;
  assign n22339 = pi95  & n746;
  assign n22340 = pi94  & n748;
  assign n22341 = ~n22339 & ~n22340;
  assign n22342 = ~n22338 & ~n22340;
  assign n22343 = ~n22339 & n22342;
  assign n22344 = ~n22338 & n22341;
  assign n22345 = ~n22337 & n41580;
  assign n22346 = pi41  & ~n22345;
  assign n22347 = pi41  & ~n22346;
  assign n22348 = pi41  & n22345;
  assign n22349 = ~n22345 & ~n22346;
  assign n22350 = ~pi41  & ~n22345;
  assign n22351 = ~n41581 & ~n41582;
  assign n22352 = ~n22336 & n22351;
  assign n22353 = n22336 & ~n22351;
  assign n22354 = ~n22352 & ~n22353;
  assign n22355 = ~n41495 & n22354;
  assign n22356 = n41495 & ~n22354;
  assign n22357 = ~n22355 & ~n22356;
  assign n22358 = ~n22157 & n22357;
  assign n22359 = n22157 & ~n22357;
  assign n22360 = ~n22358 & ~n22359;
  assign n22361 = ~n22142 & n22360;
  assign n22362 = n22142 & ~n22360;
  assign n22363 = ~n22361 & ~n22362;
  assign n22364 = n22141 & ~n22363;
  assign n22365 = ~n22141 & n22363;
  assign n22366 = ~n22141 & ~n22365;
  assign n22367 = n22363 & ~n22365;
  assign n22368 = ~n22366 & ~n22367;
  assign n22369 = ~n22364 & ~n22365;
  assign n22370 = n22126 & ~n41583;
  assign n22371 = ~n22126 & n41583;
  assign n22372 = n22126 & ~n22370;
  assign n22373 = ~n41583 & ~n22370;
  assign n22374 = ~n22372 & ~n22373;
  assign n22375 = ~n22370 & ~n22371;
  assign n22376 = ~n41544 & ~n41584;
  assign n22377 = n41544 & n41584;
  assign n22378 = ~n41544 & n41584;
  assign n22379 = n41544 & ~n41584;
  assign n22380 = ~n22378 & ~n22379;
  assign n22381 = ~n22376 & ~n22377;
  assign n22382 = n22083 & ~n41585;
  assign n22383 = ~n22083 & n41585;
  assign n22384 = n22083 & ~n22382;
  assign n22385 = ~n41585 & ~n22382;
  assign n22386 = ~n22384 & ~n22385;
  assign n22387 = ~n22382 & ~n22383;
  assign n22388 = n5576 & n11276;
  assign n22389 = pi111  & n38406;
  assign n22390 = pi113  & n5591;
  assign n22391 = pi112  & n5593;
  assign n22392 = ~n22390 & ~n22391;
  assign n22393 = ~n22389 & ~n22391;
  assign n22394 = ~n22390 & n22393;
  assign n22395 = ~n22389 & n22392;
  assign n22396 = ~n22388 & n41587;
  assign n22397 = pi23  & ~n22396;
  assign n22398 = pi23  & ~n22397;
  assign n22399 = pi23  & n22396;
  assign n22400 = ~n22396 & ~n22397;
  assign n22401 = ~pi23  & ~n22396;
  assign n22402 = ~n41588 & ~n41589;
  assign n22403 = ~n21906 & ~n21914;
  assign n22404 = ~n22402 & ~n22403;
  assign n22405 = n22402 & n22403;
  assign n22406 = ~n22402 & ~n22404;
  assign n22407 = ~n22402 & n22403;
  assign n22408 = ~n22403 & ~n22404;
  assign n22409 = n22402 & ~n22403;
  assign n22410 = ~n41590 & ~n41591;
  assign n22411 = ~n22404 & ~n22405;
  assign n22412 = ~n41586 & ~n41592;
  assign n22413 = n41586 & n41592;
  assign n22414 = n41586 & ~n41592;
  assign n22415 = ~n41586 & n41592;
  assign n22416 = ~n22414 & ~n22415;
  assign n22417 = ~n22412 & ~n22413;
  assign n22418 = n22064 & ~n41593;
  assign n22419 = ~n22064 & n41593;
  assign n22420 = n22064 & ~n22418;
  assign n22421 = ~n41593 & ~n22418;
  assign n22422 = ~n22420 & ~n22421;
  assign n22423 = ~n22418 & ~n22419;
  assign n22424 = n22043 & ~n41594;
  assign n22425 = ~n22043 & n41594;
  assign n22426 = ~n22424 & ~n22425;
  assign n22427 = n22022 & ~n22425;
  assign n22428 = ~n22424 & n22427;
  assign n22429 = n22022 & n22426;
  assign n22430 = ~n22022 & ~n22426;
  assign n22431 = n22022 & ~n41595;
  assign n22432 = ~n22425 & ~n41595;
  assign n22433 = ~n22424 & n22432;
  assign n22434 = n22426 & ~n41595;
  assign n22435 = ~n22431 & ~n41596;
  assign n22436 = ~n41595 & ~n22430;
  assign n22437 = n22003 & ~n41597;
  assign n22438 = ~n22003 & n41597;
  assign n22439 = ~n22437 & ~n22438;
  assign n22440 = n21984 & ~n22438;
  assign n22441 = ~n22437 & n22440;
  assign n22442 = n21984 & n22439;
  assign n22443 = ~n21984 & ~n22439;
  assign n22444 = n21984 & ~n41598;
  assign n22445 = ~n22438 & ~n41598;
  assign n22446 = ~n22437 & n22445;
  assign n22447 = n22439 & ~n41598;
  assign n22448 = ~n22444 & ~n41599;
  assign n22449 = ~n41598 & ~n22443;
  assign n22450 = ~n21967 & ~n41600;
  assign n22451 = n21967 & n41600;
  assign n22452 = ~n41600 & ~n22450;
  assign n22453 = ~n21967 & ~n22450;
  assign n22454 = ~n22452 & ~n22453;
  assign n22455 = ~n22450 & ~n22451;
  assign n22456 = ~n21966 & ~n41601;
  assign n22457 = n21966 & n41601;
  assign po70  = ~n22456 & ~n22457;
  assign n22459 = ~n22450 & ~n22456;
  assign n22460 = n563 & n14961;
  assign n22461 = pi121  & n37482;
  assign n22462 = pi123  & n578;
  assign n22463 = pi122  & n580;
  assign n22464 = ~n22462 & ~n22463;
  assign n22465 = ~n22461 & ~n22463;
  assign n22466 = ~n22462 & n22465;
  assign n22467 = ~n22461 & n22464;
  assign n22468 = ~n22460 & n41602;
  assign n22469 = pi14  & ~n22468;
  assign n22470 = pi14  & ~n22469;
  assign n22471 = pi14  & n22468;
  assign n22472 = ~n22468 & ~n22469;
  assign n22473 = ~pi14  & ~n22468;
  assign n22474 = ~n41603 & ~n41604;
  assign n22475 = ~n22042 & ~n22424;
  assign n22476 = ~n22474 & ~n22475;
  assign n22477 = n22474 & n22475;
  assign n22478 = ~n22474 & ~n22476;
  assign n22479 = ~n22474 & n22475;
  assign n22480 = ~n22475 & ~n22476;
  assign n22481 = n22474 & ~n22475;
  assign n22482 = ~n41605 & ~n41606;
  assign n22483 = ~n22476 & ~n22477;
  assign n22484 = n8175 & n14913;
  assign n22485 = pi118  & n38895;
  assign n22486 = pi120  & n8190;
  assign n22487 = pi119  & n8192;
  assign n22488 = ~n22486 & ~n22487;
  assign n22489 = ~n22485 & ~n22487;
  assign n22490 = ~n22486 & n22489;
  assign n22491 = ~n22485 & n22488;
  assign n22492 = ~n22484 & n41608;
  assign n22493 = pi17  & ~n22492;
  assign n22494 = pi17  & ~n22493;
  assign n22495 = pi17  & n22492;
  assign n22496 = ~n22492 & ~n22493;
  assign n22497 = ~pi17  & ~n22492;
  assign n22498 = ~n41609 & ~n41610;
  assign n22499 = ~n22063 & n41593;
  assign n22500 = ~n22063 & ~n22418;
  assign n22501 = ~n22062 & ~n22499;
  assign n22502 = n22498 & n41611;
  assign n22503 = ~n22498 & ~n41611;
  assign n22504 = ~n22502 & ~n22503;
  assign n22505 = n5576 & n11258;
  assign n22506 = pi112  & n38406;
  assign n22507 = pi114  & n5591;
  assign n22508 = pi113  & n5593;
  assign n22509 = ~n22507 & ~n22508;
  assign n22510 = ~n22506 & ~n22508;
  assign n22511 = ~n22507 & n22510;
  assign n22512 = ~n22506 & n22509;
  assign n22513 = ~n22505 & n41612;
  assign n22514 = pi23  & ~n22513;
  assign n22515 = pi23  & ~n22514;
  assign n22516 = pi23  & n22513;
  assign n22517 = ~n22513 & ~n22514;
  assign n22518 = ~pi23  & ~n22513;
  assign n22519 = ~n41613 & ~n41614;
  assign n22520 = ~n22081 & ~n22382;
  assign n22521 = n22519 & n22520;
  assign n22522 = ~n22519 & ~n22520;
  assign n22523 = ~n22521 & ~n22522;
  assign n22524 = n565 & n4492;
  assign n22525 = pi109  & n38208;
  assign n22526 = pi111  & n4507;
  assign n22527 = pi110  & n4509;
  assign n22528 = ~n22526 & ~n22527;
  assign n22529 = ~n22525 & ~n22527;
  assign n22530 = ~n22526 & n22529;
  assign n22531 = ~n22525 & n22528;
  assign n22532 = ~n22524 & n41615;
  assign n22533 = pi26  & ~n22532;
  assign n22534 = pi26  & ~n22533;
  assign n22535 = pi26  & n22532;
  assign n22536 = ~n22532 & ~n22533;
  assign n22537 = ~pi26  & ~n22532;
  assign n22538 = ~n41616 & ~n41617;
  assign n22539 = ~n22100 & ~n22376;
  assign n22540 = ~n22538 & ~n22539;
  assign n22541 = n22538 & n22539;
  assign n22542 = ~n22538 & ~n22540;
  assign n22543 = ~n22538 & n22539;
  assign n22544 = ~n22539 & ~n22540;
  assign n22545 = n22538 & ~n22539;
  assign n22546 = ~n41618 & ~n41619;
  assign n22547 = ~n22540 & ~n22541;
  assign n22548 = n649 & n8229;
  assign n22549 = pi103  & n37496;
  assign n22550 = pi105  & n662;
  assign n22551 = pi104  & n664;
  assign n22552 = ~n22550 & ~n22551;
  assign n22553 = ~n22549 & ~n22551;
  assign n22554 = ~n22550 & n22553;
  assign n22555 = ~n22549 & n22552;
  assign n22556 = ~n22548 & n41621;
  assign n22557 = pi32  & ~n22556;
  assign n22558 = pi32  & ~n22557;
  assign n22559 = pi32  & n22556;
  assign n22560 = ~n22556 & ~n22557;
  assign n22561 = ~pi32  & ~n22556;
  assign n22562 = ~n41622 & ~n41623;
  assign n22563 = n22141 & ~n22361;
  assign n22564 = ~n22361 & ~n22365;
  assign n22565 = ~n22362 & ~n22563;
  assign n22566 = n22562 & n41624;
  assign n22567 = ~n22562 & ~n41624;
  assign n22568 = ~n22566 & ~n22567;
  assign n22569 = ~n22355 & ~n22358;
  assign n22570 = n636 & n894;
  assign n22571 = pi85  & n37580;
  assign n22572 = pi87  & n896;
  assign n22573 = pi86  & n904;
  assign n22574 = ~n22572 & ~n22573;
  assign n22575 = ~n22571 & ~n22573;
  assign n22576 = ~n22572 & n22575;
  assign n22577 = ~n22571 & n22574;
  assign n22578 = ~n22570 & n41625;
  assign n22579 = pi50  & ~n22578;
  assign n22580 = pi50  & ~n22579;
  assign n22581 = pi50  & n22578;
  assign n22582 = ~n22578 & ~n22579;
  assign n22583 = ~pi50  & ~n22578;
  assign n22584 = ~n41626 & ~n41627;
  assign n22585 = n1578 & n7882;
  assign n22586 = pi76  & n39128;
  assign n22587 = pi78  & n7884;
  assign n22588 = pi77  & n7892;
  assign n22589 = ~n22587 & ~n22588;
  assign n22590 = ~n22586 & ~n22588;
  assign n22591 = ~n22587 & n22590;
  assign n22592 = ~n22586 & n22589;
  assign n22593 = ~n22585 & n41628;
  assign n22594 = pi59  & ~n22593;
  assign n22595 = pi59  & ~n22594;
  assign n22596 = pi59  & n22593;
  assign n22597 = ~n22593 & ~n22594;
  assign n22598 = ~pi59  & ~n22593;
  assign n22599 = ~n41629 & ~n41630;
  assign n22600 = n720 & n12674;
  assign n22601 = pi73  & n40107;
  assign n22602 = pi75  & n12676;
  assign n22603 = pi74  & n12684;
  assign n22604 = ~n22602 & ~n22603;
  assign n22605 = ~n22601 & ~n22603;
  assign n22606 = ~n22602 & n22605;
  assign n22607 = ~n22601 & n22604;
  assign n22608 = ~n22600 & n41631;
  assign n22609 = pi62  & ~n22608;
  assign n22610 = pi62  & ~n22609;
  assign n22611 = pi62  & n22608;
  assign n22612 = ~n22608 & ~n22609;
  assign n22613 = ~pi62  & ~n22608;
  assign n22614 = ~n41632 & ~n41633;
  assign n22615 = ~n22169 & ~n22187;
  assign n22616 = pi72  & ~n40814;
  assign n22617 = pi71  & n18285;
  assign n22618 = ~n22616 & ~n22617;
  assign n22619 = n22168 & ~n22618;
  assign n22620 = ~n22168 & n22618;
  assign n22621 = ~n22619 & ~n22620;
  assign n22622 = ~n22615 & ~n22620;
  assign n22623 = ~n22619 & n22622;
  assign n22624 = ~n22615 & n22621;
  assign n22625 = n22615 & ~n22621;
  assign n22626 = ~n22615 & ~n41634;
  assign n22627 = ~n22620 & ~n41634;
  assign n22628 = ~n22619 & n22627;
  assign n22629 = ~n22626 & ~n22628;
  assign n22630 = ~n41634 & ~n22625;
  assign n22631 = ~n22614 & ~n41635;
  assign n22632 = n22614 & n41635;
  assign n22633 = n22614 & ~n41635;
  assign n22634 = ~n22614 & n41635;
  assign n22635 = ~n22633 & ~n22634;
  assign n22636 = ~n22631 & ~n22632;
  assign n22637 = ~n22599 & ~n41636;
  assign n22638 = n22599 & n41636;
  assign n22639 = ~n22637 & ~n22638;
  assign n22640 = ~n22190 & n22207;
  assign n22641 = ~n22190 & ~n22208;
  assign n22642 = ~n22191 & ~n22640;
  assign n22643 = ~n22639 & n41637;
  assign n22644 = n22639 & ~n41637;
  assign n22645 = ~n22643 & ~n22644;
  assign n22646 = n2154 & n4312;
  assign n22647 = pi79  & n38376;
  assign n22648 = pi81  & n4314;
  assign n22649 = pi80  & n4322;
  assign n22650 = ~n22648 & ~n22649;
  assign n22651 = ~n22647 & ~n22649;
  assign n22652 = ~n22648 & n22651;
  assign n22653 = ~n22647 & n22650;
  assign n22654 = ~n22646 & n41638;
  assign n22655 = pi56  & ~n22654;
  assign n22656 = pi56  & ~n22655;
  assign n22657 = pi56  & n22654;
  assign n22658 = ~n22654 & ~n22655;
  assign n22659 = ~pi56  & ~n22654;
  assign n22660 = ~n41639 & ~n41640;
  assign n22661 = n22645 & ~n22660;
  assign n22662 = ~n22645 & n22660;
  assign n22663 = n22645 & ~n22661;
  assign n22664 = ~n22660 & ~n22661;
  assign n22665 = ~n22663 & ~n22664;
  assign n22666 = ~n22661 & ~n22662;
  assign n22667 = ~n22215 & n22231;
  assign n22668 = ~n22215 & ~n22233;
  assign n22669 = ~n22214 & ~n22667;
  assign n22670 = n41641 & n41642;
  assign n22671 = ~n41641 & ~n41642;
  assign n22672 = ~n22670 & ~n22671;
  assign n22673 = n1971 & n2591;
  assign n22674 = pi82  & n37864;
  assign n22675 = pi84  & n1973;
  assign n22676 = pi83  & n1981;
  assign n22677 = ~n22675 & ~n22676;
  assign n22678 = ~n22674 & ~n22676;
  assign n22679 = ~n22675 & n22678;
  assign n22680 = ~n22674 & n22677;
  assign n22681 = ~n22673 & n41643;
  assign n22682 = pi53  & ~n22681;
  assign n22683 = pi53  & ~n22682;
  assign n22684 = pi53  & n22681;
  assign n22685 = ~n22681 & ~n22682;
  assign n22686 = ~pi53  & ~n22681;
  assign n22687 = ~n41644 & ~n41645;
  assign n22688 = ~n22672 & n22687;
  assign n22689 = n22672 & ~n22687;
  assign n22690 = ~n22688 & ~n22689;
  assign n22691 = ~n22239 & n22255;
  assign n22692 = ~n22239 & ~n22256;
  assign n22693 = ~n22238 & ~n22691;
  assign n22694 = n22690 & ~n41646;
  assign n22695 = ~n22690 & n41646;
  assign n22696 = ~n41646 & ~n22694;
  assign n22697 = n22690 & ~n22694;
  assign n22698 = ~n22696 & ~n22697;
  assign n22699 = ~n22694 & ~n22695;
  assign n22700 = ~n22584 & ~n41647;
  assign n22701 = n22584 & ~n22697;
  assign n22702 = ~n22696 & n22701;
  assign n22703 = n22584 & n41647;
  assign n22704 = ~n22700 & ~n41648;
  assign n22705 = ~n22263 & n22279;
  assign n22706 = ~n22263 & ~n22281;
  assign n22707 = ~n22262 & ~n22705;
  assign n22708 = n22704 & ~n41649;
  assign n22709 = ~n22704 & n41649;
  assign n22710 = ~n22708 & ~n22709;
  assign n22711 = n785 & n3566;
  assign n22712 = pi88  & n37520;
  assign n22713 = pi90  & n787;
  assign n22714 = pi89  & n795;
  assign n22715 = ~n22713 & ~n22714;
  assign n22716 = ~n22712 & ~n22714;
  assign n22717 = ~n22713 & n22716;
  assign n22718 = ~n22712 & n22715;
  assign n22719 = ~n22711 & n41650;
  assign n22720 = pi47  & ~n22719;
  assign n22721 = pi47  & ~n22720;
  assign n22722 = pi47  & n22719;
  assign n22723 = ~n22719 & ~n22720;
  assign n22724 = ~pi47  & ~n22719;
  assign n22725 = ~n41651 & ~n41652;
  assign n22726 = n22710 & ~n22725;
  assign n22727 = ~n22710 & n22725;
  assign n22728 = n22710 & ~n22726;
  assign n22729 = ~n22725 & ~n22726;
  assign n22730 = ~n22728 & ~n22729;
  assign n22731 = ~n22726 & ~n22727;
  assign n22732 = ~n22287 & n22303;
  assign n22733 = ~n22287 & ~n22304;
  assign n22734 = ~n22286 & ~n22732;
  assign n22735 = n41653 & n41654;
  assign n22736 = ~n41653 & ~n41654;
  assign n22737 = ~n22735 & ~n22736;
  assign n22738 = n940 & n4544;
  assign n22739 = pi91  & n37541;
  assign n22740 = pi93  & n953;
  assign n22741 = pi92  & n955;
  assign n22742 = ~n22740 & ~n22741;
  assign n22743 = ~n22739 & ~n22741;
  assign n22744 = ~n22740 & n22743;
  assign n22745 = ~n22739 & n22742;
  assign n22746 = ~n22738 & n41655;
  assign n22747 = pi44  & ~n22746;
  assign n22748 = pi44  & ~n22747;
  assign n22749 = pi44  & n22746;
  assign n22750 = ~n22746 & ~n22747;
  assign n22751 = ~pi44  & ~n22746;
  assign n22752 = ~n41656 & ~n41657;
  assign n22753 = ~n22737 & n22752;
  assign n22754 = n22737 & ~n22752;
  assign n22755 = n22737 & ~n22754;
  assign n22756 = ~n22752 & ~n22754;
  assign n22757 = ~n22755 & ~n22756;
  assign n22758 = ~n22753 & ~n22754;
  assign n22759 = ~n22311 & n22327;
  assign n22760 = ~n22311 & ~n22329;
  assign n22761 = ~n22310 & ~n22759;
  assign n22762 = n41658 & n41659;
  assign n22763 = ~n41658 & ~n41659;
  assign n22764 = ~n22762 & ~n22763;
  assign n22765 = n733 & n5281;
  assign n22766 = pi94  & n37510;
  assign n22767 = pi96  & n746;
  assign n22768 = pi95  & n748;
  assign n22769 = ~n22767 & ~n22768;
  assign n22770 = ~n22766 & ~n22768;
  assign n22771 = ~n22767 & n22770;
  assign n22772 = ~n22766 & n22769;
  assign n22773 = ~n22765 & n41660;
  assign n22774 = pi41  & ~n22773;
  assign n22775 = pi41  & ~n22774;
  assign n22776 = pi41  & n22773;
  assign n22777 = ~n22773 & ~n22774;
  assign n22778 = ~pi41  & ~n22773;
  assign n22779 = ~n41661 & ~n41662;
  assign n22780 = ~n22764 & n22779;
  assign n22781 = n22764 & ~n22779;
  assign n22782 = ~n22780 & ~n22781;
  assign n22783 = ~n22335 & ~n22353;
  assign n22784 = n22782 & ~n22783;
  assign n22785 = ~n22782 & n22783;
  assign n22786 = ~n22784 & ~n22785;
  assign n22787 = n691 & n5578;
  assign n22788 = pi97  & n37503;
  assign n22789 = pi99  & n704;
  assign n22790 = pi98  & n706;
  assign n22791 = ~n22789 & ~n22790;
  assign n22792 = ~n22788 & ~n22790;
  assign n22793 = ~n22789 & n22792;
  assign n22794 = ~n22788 & n22791;
  assign n22795 = ~n22787 & n41663;
  assign n22796 = pi38  & ~n22795;
  assign n22797 = pi38  & ~n22796;
  assign n22798 = pi38  & n22795;
  assign n22799 = ~n22795 & ~n22796;
  assign n22800 = ~pi38  & ~n22795;
  assign n22801 = ~n41664 & ~n41665;
  assign n22802 = ~n22786 & n22801;
  assign n22803 = n22786 & ~n22801;
  assign n22804 = n22786 & ~n22803;
  assign n22805 = ~n22801 & ~n22803;
  assign n22806 = ~n22804 & ~n22805;
  assign n22807 = ~n22802 & ~n22803;
  assign n22808 = n22569 & n41666;
  assign n22809 = ~n22569 & ~n41666;
  assign n22810 = ~n22808 & ~n22809;
  assign n22811 = n2104 & n6819;
  assign n22812 = pi100  & n37758;
  assign n22813 = pi102  & n2117;
  assign n22814 = pi101  & n2119;
  assign n22815 = ~n22813 & ~n22814;
  assign n22816 = ~n22812 & ~n22814;
  assign n22817 = ~n22813 & n22816;
  assign n22818 = ~n22812 & n22815;
  assign n22819 = ~n22811 & n41667;
  assign n22820 = pi35  & ~n22819;
  assign n22821 = pi35  & ~n22820;
  assign n22822 = pi35  & n22819;
  assign n22823 = ~n22819 & ~n22820;
  assign n22824 = ~pi35  & ~n22819;
  assign n22825 = ~n41668 & ~n41669;
  assign n22826 = n22810 & ~n22825;
  assign n22827 = ~n22810 & n22825;
  assign n22828 = ~n22826 & ~n22827;
  assign n22829 = n22568 & ~n22827;
  assign n22830 = ~n22826 & n22829;
  assign n22831 = n22568 & n22828;
  assign n22832 = ~n22568 & ~n22828;
  assign n22833 = n22568 & ~n41670;
  assign n22834 = ~n22827 & ~n41670;
  assign n22835 = ~n22826 & n22834;
  assign n22836 = n22828 & ~n41670;
  assign n22837 = ~n22833 & ~n41671;
  assign n22838 = ~n41670 & ~n22832;
  assign n22839 = n607 & n9277;
  assign n22840 = pi106  & n37489;
  assign n22841 = pi108  & n620;
  assign n22842 = pi107  & n622;
  assign n22843 = ~n22841 & ~n22842;
  assign n22844 = ~n22840 & ~n22842;
  assign n22845 = ~n22841 & n22844;
  assign n22846 = ~n22840 & n22843;
  assign n22847 = ~n607 & n41673;
  assign n22848 = ~n9277 & n41673;
  assign n22849 = ~n22847 & ~n22848;
  assign n22850 = ~n22839 & n41673;
  assign n22851 = pi29  & ~n41674;
  assign n22852 = ~pi29  & n41674;
  assign n22853 = ~n22851 & ~n22852;
  assign n22854 = ~n22125 & n41583;
  assign n22855 = ~n22125 & ~n22370;
  assign n22856 = ~n22124 & ~n22854;
  assign n22857 = ~n22853 & ~n41675;
  assign n22858 = n22853 & n41675;
  assign n22859 = ~n41675 & ~n22857;
  assign n22860 = n22853 & ~n41675;
  assign n22861 = ~n22853 & ~n22857;
  assign n22862 = ~n22853 & n41675;
  assign n22863 = ~n41676 & ~n41677;
  assign n22864 = ~n22857 & ~n22858;
  assign n22865 = ~n41672 & ~n41678;
  assign n22866 = n41672 & n41678;
  assign n22867 = ~n41672 & ~n22865;
  assign n22868 = ~n41672 & n41678;
  assign n22869 = ~n41678 & ~n22865;
  assign n22870 = n41672 & ~n41678;
  assign n22871 = ~n41679 & ~n41680;
  assign n22872 = ~n22865 & ~n22866;
  assign n22873 = ~n41620 & ~n41681;
  assign n22874 = n41620 & n41681;
  assign n22875 = ~n41620 & ~n22873;
  assign n22876 = ~n41681 & ~n22873;
  assign n22877 = ~n22875 & ~n22876;
  assign n22878 = ~n22873 & ~n22874;
  assign n22879 = ~n22523 & n41682;
  assign n22880 = n22523 & ~n41682;
  assign n22881 = ~n22879 & ~n22880;
  assign n22882 = ~n22404 & ~n22412;
  assign n22883 = n6785 & n13079;
  assign n22884 = pi115  & n38631;
  assign n22885 = pi117  & n6800;
  assign n22886 = pi116  & n6802;
  assign n22887 = ~n22885 & ~n22886;
  assign n22888 = ~n22884 & ~n22886;
  assign n22889 = ~n22885 & n22888;
  assign n22890 = ~n22884 & n22887;
  assign n22891 = ~n6785 & n41683;
  assign n22892 = ~n13079 & n41683;
  assign n22893 = ~n22891 & ~n22892;
  assign n22894 = ~n22883 & n41683;
  assign n22895 = pi20  & ~n41684;
  assign n22896 = ~pi20  & n41684;
  assign n22897 = ~n22895 & ~n22896;
  assign n22898 = ~n22882 & ~n22897;
  assign n22899 = n22882 & n22897;
  assign n22900 = ~n22882 & ~n22898;
  assign n22901 = ~n22882 & n22897;
  assign n22902 = ~n22897 & ~n22898;
  assign n22903 = n22882 & ~n22897;
  assign n22904 = ~n41685 & ~n41686;
  assign n22905 = ~n22898 & ~n22899;
  assign n22906 = n22881 & ~n41687;
  assign n22907 = ~n22881 & n41687;
  assign n22908 = n22881 & ~n22906;
  assign n22909 = n22881 & n41687;
  assign n22910 = ~n41687 & ~n22906;
  assign n22911 = ~n22881 & ~n41687;
  assign n22912 = ~n41688 & ~n41689;
  assign n22913 = ~n22906 & ~n22907;
  assign n22914 = n22504 & ~n41690;
  assign n22915 = ~n22504 & n41690;
  assign n22916 = n22504 & ~n22914;
  assign n22917 = ~n41690 & ~n22914;
  assign n22918 = ~n22916 & ~n22917;
  assign n22919 = ~n22914 & ~n22915;
  assign n22920 = ~n41607 & ~n41691;
  assign n22921 = n41607 & n41691;
  assign n22922 = n41607 & ~n41691;
  assign n22923 = ~n41607 & n41691;
  assign n22924 = ~n22922 & ~n22923;
  assign n22925 = ~n22920 & ~n22921;
  assign n22926 = ~n22020 & ~n41595;
  assign n22927 = n269 & n15021;
  assign n22928 = pi124  & n37475;
  assign n22929 = pi126  & n536;
  assign n22930 = pi125  & n538;
  assign n22931 = ~n22929 & ~n22930;
  assign n22932 = ~n22928 & ~n22930;
  assign n22933 = ~n22929 & n22932;
  assign n22934 = ~n22928 & n22931;
  assign n22935 = ~n269 & n41693;
  assign n22936 = ~n15021 & n41693;
  assign n22937 = ~n22935 & ~n22936;
  assign n22938 = ~n22927 & n41693;
  assign n22939 = pi11  & ~n41694;
  assign n22940 = ~pi11  & n41694;
  assign n22941 = ~n22939 & ~n22940;
  assign n22942 = ~n22926 & ~n22941;
  assign n22943 = n22926 & n22941;
  assign n22944 = ~n22926 & ~n22942;
  assign n22945 = ~n22926 & n22941;
  assign n22946 = ~n22941 & ~n22942;
  assign n22947 = n22926 & ~n22941;
  assign n22948 = ~n41695 & ~n41696;
  assign n22949 = ~n22942 & ~n22943;
  assign n22950 = ~n41692 & ~n41697;
  assign n22951 = n41692 & ~n41696;
  assign n22952 = ~n41695 & n22951;
  assign n22953 = n41692 & ~n41695;
  assign n22954 = ~n41696 & n22953;
  assign n22955 = n41692 & n41697;
  assign n22956 = ~n22950 & ~n41698;
  assign n22957 = ~n22002 & ~n22437;
  assign n22958 = n13010 & ~n18675;
  assign n22959 = ~n39810 & ~n22958;
  assign n22960 = pi127  & n39810;
  assign n22961 = n13010 & n18680;
  assign n22962 = ~n22960 & ~n22961;
  assign n22963 = pi127  & ~n22959;
  assign n22964 = pi8  & ~n41699;
  assign n22965 = pi8  & ~n22964;
  assign n22966 = pi8  & n41699;
  assign n22967 = ~n41699 & ~n22964;
  assign n22968 = ~pi8  & ~n41699;
  assign n22969 = ~n41700 & ~n41701;
  assign n22970 = ~n22957 & ~n22969;
  assign n22971 = n22957 & n22969;
  assign n22972 = ~n22957 & ~n22970;
  assign n22973 = ~n22969 & ~n22970;
  assign n22974 = ~n22972 & ~n22973;
  assign n22975 = ~n22970 & ~n22971;
  assign n22976 = n22956 & ~n41702;
  assign n22977 = ~n22956 & n41702;
  assign n22978 = ~n22976 & ~n22977;
  assign n22979 = ~n21982 & ~n22439;
  assign n22980 = ~n21982 & ~n41598;
  assign n22981 = ~n21983 & ~n22979;
  assign n22982 = n22978 & ~n41703;
  assign n22983 = ~n22978 & n41703;
  assign n22984 = ~n41703 & ~n22982;
  assign n22985 = n22978 & ~n22982;
  assign n22986 = ~n22984 & ~n22985;
  assign n22987 = ~n22982 & ~n22983;
  assign n22988 = ~n22459 & ~n41704;
  assign n22989 = n22459 & ~n22985;
  assign n22990 = ~n22984 & n22989;
  assign n22991 = n22459 & n41704;
  assign po71  = ~n22988 & ~n41705;
  assign n22993 = ~n22982 & ~n22988;
  assign n22994 = ~n22970 & ~n22976;
  assign n22995 = n8175 & n15091;
  assign n22996 = pi119  & n38895;
  assign n22997 = pi121  & n8190;
  assign n22998 = pi120  & n8192;
  assign n22999 = ~n22997 & ~n22998;
  assign n23000 = ~n22996 & ~n22998;
  assign n23001 = ~n22997 & n23000;
  assign n23002 = ~n22996 & n22999;
  assign n23003 = ~n22995 & n41706;
  assign n23004 = pi17  & ~n23003;
  assign n23005 = pi17  & ~n23004;
  assign n23006 = pi17  & n23003;
  assign n23007 = ~n23003 & ~n23004;
  assign n23008 = ~pi17  & ~n23003;
  assign n23009 = ~n41707 & ~n41708;
  assign n23010 = ~n22503 & n41690;
  assign n23011 = ~n22503 & ~n22914;
  assign n23012 = ~n22502 & ~n23010;
  assign n23013 = n23009 & n41709;
  assign n23014 = ~n23009 & ~n41709;
  assign n23015 = ~n23013 & ~n23014;
  assign n23016 = ~n22898 & ~n22906;
  assign n23017 = n6785 & n13057;
  assign n23018 = pi116  & n38631;
  assign n23019 = pi118  & n6800;
  assign n23020 = pi117  & n6802;
  assign n23021 = ~n23019 & ~n23020;
  assign n23022 = ~n23018 & ~n23020;
  assign n23023 = ~n23019 & n23022;
  assign n23024 = ~n23018 & n23021;
  assign n23025 = ~n23017 & n41710;
  assign n23026 = pi20  & ~n23025;
  assign n23027 = pi20  & ~n23026;
  assign n23028 = pi20  & n23025;
  assign n23029 = ~n23025 & ~n23026;
  assign n23030 = ~pi20  & ~n23025;
  assign n23031 = ~n41711 & ~n41712;
  assign n23032 = ~n23016 & ~n23031;
  assign n23033 = n23016 & n23031;
  assign n23034 = ~n23016 & ~n23032;
  assign n23035 = ~n23016 & n23031;
  assign n23036 = ~n23031 & ~n23032;
  assign n23037 = n23016 & ~n23031;
  assign n23038 = ~n41713 & ~n41714;
  assign n23039 = ~n23032 & ~n23033;
  assign n23040 = n523 & n5576;
  assign n23041 = pi113  & n38406;
  assign n23042 = pi115  & n5591;
  assign n23043 = pi114  & n5593;
  assign n23044 = ~n23042 & ~n23043;
  assign n23045 = ~n23041 & ~n23043;
  assign n23046 = ~n23042 & n23045;
  assign n23047 = ~n23041 & n23044;
  assign n23048 = ~n23040 & n41716;
  assign n23049 = pi23  & ~n23048;
  assign n23050 = pi23  & ~n23049;
  assign n23051 = pi23  & n23048;
  assign n23052 = ~n23048 & ~n23049;
  assign n23053 = ~pi23  & ~n23048;
  assign n23054 = ~n41717 & ~n41718;
  assign n23055 = ~n22522 & ~n22880;
  assign n23056 = ~n23054 & ~n23055;
  assign n23057 = n23054 & n23055;
  assign n23058 = ~n23056 & ~n23057;
  assign n23059 = n4492 & n10844;
  assign n23060 = pi110  & n38208;
  assign n23061 = pi112  & n4507;
  assign n23062 = pi111  & n4509;
  assign n23063 = ~n23061 & ~n23062;
  assign n23064 = ~n23060 & ~n23062;
  assign n23065 = ~n23061 & n23064;
  assign n23066 = ~n23060 & n23063;
  assign n23067 = ~n23059 & n41719;
  assign n23068 = pi26  & ~n23067;
  assign n23069 = pi26  & ~n23068;
  assign n23070 = pi26  & n23067;
  assign n23071 = ~n23067 & ~n23068;
  assign n23072 = ~pi26  & ~n23067;
  assign n23073 = ~n41720 & ~n41721;
  assign n23074 = ~n22540 & ~n22873;
  assign n23075 = n23073 & n23074;
  assign n23076 = ~n23073 & ~n23074;
  assign n23077 = ~n23075 & ~n23076;
  assign n23078 = ~n22857 & ~n22865;
  assign n23079 = n607 & n9701;
  assign n23080 = pi107  & n37489;
  assign n23081 = pi109  & n620;
  assign n23082 = pi108  & n622;
  assign n23083 = ~n23081 & ~n23082;
  assign n23084 = ~n23080 & ~n23082;
  assign n23085 = ~n23081 & n23084;
  assign n23086 = ~n23080 & n23083;
  assign n23087 = ~n23079 & n41722;
  assign n23088 = pi29  & ~n23087;
  assign n23089 = pi29  & ~n23088;
  assign n23090 = pi29  & n23087;
  assign n23091 = ~n23087 & ~n23088;
  assign n23092 = ~pi29  & ~n23087;
  assign n23093 = ~n41723 & ~n41724;
  assign n23094 = ~n23078 & ~n23093;
  assign n23095 = n23078 & n23093;
  assign n23096 = ~n23078 & ~n23094;
  assign n23097 = ~n23078 & n23093;
  assign n23098 = ~n23093 & ~n23094;
  assign n23099 = n23078 & ~n23093;
  assign n23100 = ~n41725 & ~n41726;
  assign n23101 = ~n23094 & ~n23095;
  assign n23102 = ~n22809 & ~n22826;
  assign n23103 = n691 & n6474;
  assign n23104 = pi98  & n37503;
  assign n23105 = pi100  & n704;
  assign n23106 = pi99  & n706;
  assign n23107 = ~n23105 & ~n23106;
  assign n23108 = ~n23104 & ~n23106;
  assign n23109 = ~n23105 & n23108;
  assign n23110 = ~n23104 & n23107;
  assign n23111 = ~n23103 & n41728;
  assign n23112 = pi38  & ~n23111;
  assign n23113 = pi38  & ~n23112;
  assign n23114 = pi38  & n23111;
  assign n23115 = ~n23111 & ~n23112;
  assign n23116 = ~pi38  & ~n23111;
  assign n23117 = ~n41729 & ~n41730;
  assign n23118 = ~n22763 & ~n22781;
  assign n23119 = n733 & n5630;
  assign n23120 = pi95  & n37510;
  assign n23121 = pi97  & n746;
  assign n23122 = pi96  & n748;
  assign n23123 = ~n23121 & ~n23122;
  assign n23124 = ~n23120 & ~n23122;
  assign n23125 = ~n23121 & n23124;
  assign n23126 = ~n23120 & n23123;
  assign n23127 = ~n23119 & n41731;
  assign n23128 = pi41  & ~n23127;
  assign n23129 = pi41  & ~n23128;
  assign n23130 = pi41  & n23127;
  assign n23131 = ~n23127 & ~n23128;
  assign n23132 = ~pi41  & ~n23127;
  assign n23133 = ~n41732 & ~n41733;
  assign n23134 = n594 & n785;
  assign n23135 = pi89  & n37520;
  assign n23136 = pi91  & n787;
  assign n23137 = pi90  & n795;
  assign n23138 = ~n23136 & ~n23137;
  assign n23139 = ~n23135 & ~n23137;
  assign n23140 = ~n23136 & n23139;
  assign n23141 = ~n23135 & n23138;
  assign n23142 = ~n23134 & n41734;
  assign n23143 = pi47  & ~n23142;
  assign n23144 = pi47  & ~n23143;
  assign n23145 = pi47  & n23142;
  assign n23146 = ~n23142 & ~n23143;
  assign n23147 = ~pi47  & ~n23142;
  assign n23148 = ~n41735 & ~n41736;
  assign n23149 = ~n22694 & ~n22700;
  assign n23150 = n894 & n3354;
  assign n23151 = pi86  & n37580;
  assign n23152 = pi88  & n896;
  assign n23153 = pi87  & n904;
  assign n23154 = ~n23152 & ~n23153;
  assign n23155 = ~n23151 & ~n23153;
  assign n23156 = ~n23152 & n23155;
  assign n23157 = ~n23151 & n23154;
  assign n23158 = ~n23150 & n41737;
  assign n23159 = pi50  & ~n23158;
  assign n23160 = pi50  & ~n23159;
  assign n23161 = pi50  & n23158;
  assign n23162 = ~n23158 & ~n23159;
  assign n23163 = ~pi50  & ~n23158;
  assign n23164 = ~n41738 & ~n41739;
  assign n23165 = ~n22671 & ~n22689;
  assign n23166 = ~n22631 & ~n22637;
  assign n23167 = n678 & n7882;
  assign n23168 = pi77  & n39128;
  assign n23169 = pi79  & n7884;
  assign n23170 = pi78  & n7892;
  assign n23171 = ~n23169 & ~n23170;
  assign n23172 = ~n23168 & ~n23170;
  assign n23173 = ~n23169 & n23172;
  assign n23174 = ~n23168 & n23171;
  assign n23175 = ~n23167 & n41740;
  assign n23176 = pi59  & ~n23175;
  assign n23177 = pi59  & ~n23176;
  assign n23178 = pi59  & n23175;
  assign n23179 = ~n23175 & ~n23176;
  assign n23180 = ~pi59  & ~n23175;
  assign n23181 = ~n41741 & ~n41742;
  assign n23182 = n1465 & n12674;
  assign n23183 = pi74  & n40107;
  assign n23184 = pi76  & n12676;
  assign n23185 = pi75  & n12684;
  assign n23186 = ~n23184 & ~n23185;
  assign n23187 = ~n23183 & ~n23185;
  assign n23188 = ~n23184 & n23187;
  assign n23189 = ~n23183 & n23186;
  assign n23190 = ~n23182 & n41743;
  assign n23191 = pi62  & ~n23190;
  assign n23192 = pi62  & ~n23191;
  assign n23193 = pi62  & n23190;
  assign n23194 = ~n23190 & ~n23191;
  assign n23195 = ~pi62  & ~n23190;
  assign n23196 = ~n41744 & ~n41745;
  assign n23197 = ~pi8  & ~n22618;
  assign n23198 = pi8  & n22618;
  assign n23199 = pi8  & ~n22618;
  assign n23200 = ~pi8  & n22618;
  assign n23201 = ~n23199 & ~n23200;
  assign n23202 = ~n23197 & ~n23198;
  assign n23203 = pi73  & ~n40814;
  assign n23204 = pi72  & n18285;
  assign n23205 = ~n23203 & ~n23204;
  assign n23206 = ~n41746 & ~n23205;
  assign n23207 = n41746 & n23205;
  assign n23208 = ~n23206 & ~n23207;
  assign n23209 = ~n22627 & n23208;
  assign n23210 = n22627 & ~n23208;
  assign n23211 = ~n23209 & ~n23210;
  assign n23212 = n23196 & ~n23211;
  assign n23213 = ~n23196 & n23211;
  assign n23214 = n23196 & n23211;
  assign n23215 = ~n23196 & ~n23211;
  assign n23216 = ~n23214 & ~n23215;
  assign n23217 = ~n23212 & ~n23213;
  assign n23218 = ~n23181 & ~n41747;
  assign n23219 = n23181 & n41747;
  assign n23220 = ~n23218 & ~n23219;
  assign n23221 = ~n23166 & n23220;
  assign n23222 = n23166 & ~n23220;
  assign n23223 = ~n23221 & ~n23222;
  assign n23224 = n2134 & n4312;
  assign n23225 = pi80  & n38376;
  assign n23226 = pi82  & n4314;
  assign n23227 = pi81  & n4322;
  assign n23228 = ~n23226 & ~n23227;
  assign n23229 = ~n23225 & ~n23227;
  assign n23230 = ~n23226 & n23229;
  assign n23231 = ~n23225 & n23228;
  assign n23232 = ~n23224 & n41748;
  assign n23233 = pi56  & ~n23232;
  assign n23234 = pi56  & ~n23233;
  assign n23235 = pi56  & n23232;
  assign n23236 = ~n23232 & ~n23233;
  assign n23237 = ~pi56  & ~n23232;
  assign n23238 = ~n41749 & ~n41750;
  assign n23239 = n23223 & ~n23238;
  assign n23240 = ~n23223 & n23238;
  assign n23241 = n23223 & ~n23239;
  assign n23242 = n23223 & n23238;
  assign n23243 = ~n23238 & ~n23239;
  assign n23244 = ~n23223 & ~n23238;
  assign n23245 = ~n41751 & ~n41752;
  assign n23246 = ~n23239 & ~n23240;
  assign n23247 = ~n22644 & n22660;
  assign n23248 = ~n22644 & ~n22661;
  assign n23249 = ~n22643 & ~n23247;
  assign n23250 = n41753 & n41754;
  assign n23251 = ~n41753 & ~n41754;
  assign n23252 = ~n23250 & ~n23251;
  assign n23253 = n1971 & n2804;
  assign n23254 = pi83  & n37864;
  assign n23255 = pi85  & n1973;
  assign n23256 = pi84  & n1981;
  assign n23257 = ~n23255 & ~n23256;
  assign n23258 = ~n23254 & ~n23256;
  assign n23259 = ~n23255 & n23258;
  assign n23260 = ~n23254 & n23257;
  assign n23261 = ~n23253 & n41755;
  assign n23262 = pi53  & ~n23261;
  assign n23263 = pi53  & ~n23262;
  assign n23264 = pi53  & n23261;
  assign n23265 = ~n23261 & ~n23262;
  assign n23266 = ~pi53  & ~n23261;
  assign n23267 = ~n41756 & ~n41757;
  assign n23268 = n23252 & ~n23267;
  assign n23269 = ~n23252 & n23267;
  assign n23270 = n23252 & ~n23268;
  assign n23271 = n23252 & n23267;
  assign n23272 = ~n23267 & ~n23268;
  assign n23273 = ~n23252 & ~n23267;
  assign n23274 = ~n41758 & ~n41759;
  assign n23275 = ~n23268 & ~n23269;
  assign n23276 = ~n23165 & ~n41760;
  assign n23277 = n23165 & n41760;
  assign n23278 = ~n23276 & ~n23277;
  assign n23279 = ~n23164 & n23278;
  assign n23280 = n23164 & ~n23278;
  assign n23281 = ~n23164 & ~n23279;
  assign n23282 = ~n23164 & ~n23278;
  assign n23283 = n23278 & ~n23279;
  assign n23284 = n23164 & n23278;
  assign n23285 = ~n41761 & ~n41762;
  assign n23286 = ~n23279 & ~n23280;
  assign n23287 = ~n23149 & ~n41763;
  assign n23288 = n23149 & n41763;
  assign n23289 = ~n23149 & ~n23287;
  assign n23290 = ~n23149 & n41763;
  assign n23291 = ~n41763 & ~n23287;
  assign n23292 = n23149 & ~n41763;
  assign n23293 = ~n41764 & ~n41765;
  assign n23294 = ~n23287 & ~n23288;
  assign n23295 = ~n23148 & ~n41766;
  assign n23296 = n23148 & n41766;
  assign n23297 = ~n41766 & ~n23295;
  assign n23298 = ~n23148 & ~n23295;
  assign n23299 = ~n23297 & ~n23298;
  assign n23300 = ~n23295 & ~n23296;
  assign n23301 = ~n22708 & n22725;
  assign n23302 = ~n22708 & ~n22726;
  assign n23303 = ~n22709 & ~n23301;
  assign n23304 = n41767 & n41768;
  assign n23305 = ~n41767 & ~n41768;
  assign n23306 = ~n23304 & ~n23305;
  assign n23307 = n940 & n4524;
  assign n23308 = pi92  & n37541;
  assign n23309 = pi94  & n953;
  assign n23310 = pi93  & n955;
  assign n23311 = ~n23309 & ~n23310;
  assign n23312 = ~n23308 & ~n23310;
  assign n23313 = ~n23309 & n23312;
  assign n23314 = ~n23308 & n23311;
  assign n23315 = ~n23307 & n41769;
  assign n23316 = pi44  & ~n23315;
  assign n23317 = pi44  & ~n23316;
  assign n23318 = pi44  & n23315;
  assign n23319 = ~n23315 & ~n23316;
  assign n23320 = ~pi44  & ~n23315;
  assign n23321 = ~n41770 & ~n41771;
  assign n23322 = n23306 & ~n23321;
  assign n23323 = ~n23306 & n23321;
  assign n23324 = ~n23322 & ~n23323;
  assign n23325 = ~n22736 & n22752;
  assign n23326 = ~n22736 & ~n22754;
  assign n23327 = ~n22735 & ~n23325;
  assign n23328 = ~n23322 & n41772;
  assign n23329 = ~n23322 & ~n41772;
  assign n23330 = ~n23323 & ~n41772;
  assign n23331 = ~n23322 & n23330;
  assign n23332 = ~n23323 & n23329;
  assign n23333 = ~n23322 & ~n41773;
  assign n23334 = ~n23323 & ~n23328;
  assign n23335 = ~n23323 & n41774;
  assign n23336 = n23324 & n41772;
  assign n23337 = ~n41772 & ~n41773;
  assign n23338 = ~n23324 & ~n41772;
  assign n23339 = ~n41775 & ~n41776;
  assign n23340 = ~n23133 & ~n23339;
  assign n23341 = n23133 & n23339;
  assign n23342 = ~n23339 & ~n23340;
  assign n23343 = ~n23133 & ~n23340;
  assign n23344 = ~n23342 & ~n23343;
  assign n23345 = ~n23340 & ~n23341;
  assign n23346 = ~n23118 & ~n41777;
  assign n23347 = n23118 & n41777;
  assign n23348 = ~n23118 & n41777;
  assign n23349 = n23118 & ~n41777;
  assign n23350 = ~n23348 & ~n23349;
  assign n23351 = ~n23346 & ~n23347;
  assign n23352 = ~n23117 & ~n41778;
  assign n23353 = n23117 & n41778;
  assign n23354 = ~n23352 & ~n23353;
  assign n23355 = ~n22785 & ~n22801;
  assign n23356 = ~n22784 & ~n22803;
  assign n23357 = ~n22784 & ~n23355;
  assign n23358 = ~n23354 & n41779;
  assign n23359 = n23354 & ~n41779;
  assign n23360 = ~n23358 & ~n23359;
  assign n23361 = n2104 & n6787;
  assign n23362 = pi101  & n37758;
  assign n23363 = pi103  & n2117;
  assign n23364 = pi102  & n2119;
  assign n23365 = ~n23363 & ~n23364;
  assign n23366 = ~n23362 & ~n23364;
  assign n23367 = ~n23363 & n23366;
  assign n23368 = ~n23362 & n23365;
  assign n23369 = ~n23361 & n41780;
  assign n23370 = pi35  & ~n23369;
  assign n23371 = pi35  & ~n23370;
  assign n23372 = pi35  & n23369;
  assign n23373 = ~n23369 & ~n23370;
  assign n23374 = ~pi35  & ~n23369;
  assign n23375 = ~n41781 & ~n41782;
  assign n23376 = n23360 & ~n23375;
  assign n23377 = ~n23360 & n23375;
  assign n23378 = n23360 & ~n23376;
  assign n23379 = n23360 & n23375;
  assign n23380 = ~n23375 & ~n23376;
  assign n23381 = ~n23360 & ~n23375;
  assign n23382 = ~n41783 & ~n41784;
  assign n23383 = ~n23376 & ~n23377;
  assign n23384 = ~n23102 & ~n41785;
  assign n23385 = n23102 & n41785;
  assign n23386 = ~n41785 & ~n23384;
  assign n23387 = ~n23102 & ~n23384;
  assign n23388 = ~n23386 & ~n23387;
  assign n23389 = ~n23384 & ~n23385;
  assign n23390 = ~n22567 & ~n41670;
  assign n23391 = n649 & n8209;
  assign n23392 = pi104  & n37496;
  assign n23393 = pi106  & n662;
  assign n23394 = pi105  & n664;
  assign n23395 = ~n23393 & ~n23394;
  assign n23396 = ~n23392 & ~n23394;
  assign n23397 = ~n23393 & n23396;
  assign n23398 = ~n23392 & n23395;
  assign n23399 = ~n23391 & n41787;
  assign n23400 = pi32  & ~n23399;
  assign n23401 = pi32  & ~n23400;
  assign n23402 = pi32  & n23399;
  assign n23403 = ~n23399 & ~n23400;
  assign n23404 = ~pi32  & ~n23399;
  assign n23405 = ~n41788 & ~n41789;
  assign n23406 = ~n23390 & ~n23405;
  assign n23407 = n23390 & n23405;
  assign n23408 = ~n23390 & ~n23406;
  assign n23409 = ~n23390 & n23405;
  assign n23410 = ~n23405 & ~n23406;
  assign n23411 = n23390 & ~n23405;
  assign n23412 = ~n41790 & ~n41791;
  assign n23413 = ~n23406 & ~n23407;
  assign n23414 = ~n41786 & ~n41792;
  assign n23415 = n41786 & n41792;
  assign n23416 = ~n41792 & ~n23414;
  assign n23417 = n41786 & ~n41792;
  assign n23418 = ~n41786 & ~n23414;
  assign n23419 = ~n41786 & n41792;
  assign n23420 = ~n41793 & ~n41794;
  assign n23421 = ~n23414 & ~n23415;
  assign n23422 = ~n41727 & ~n41795;
  assign n23423 = n41727 & n41795;
  assign n23424 = ~n41727 & n41795;
  assign n23425 = n41727 & ~n41795;
  assign n23426 = ~n23424 & ~n23425;
  assign n23427 = ~n23422 & ~n23423;
  assign n23428 = n23077 & ~n41796;
  assign n23429 = ~n23077 & n41796;
  assign n23430 = n23077 & ~n23428;
  assign n23431 = ~n41796 & ~n23428;
  assign n23432 = ~n23430 & ~n23431;
  assign n23433 = ~n23428 & ~n23429;
  assign n23434 = n23058 & ~n41797;
  assign n23435 = ~n41797 & ~n23434;
  assign n23436 = ~n23058 & ~n41797;
  assign n23437 = n23058 & ~n23434;
  assign n23438 = n23058 & n41797;
  assign n23439 = ~n41798 & ~n41799;
  assign n23440 = ~n41715 & ~n23439;
  assign n23441 = n41715 & n23439;
  assign n23442 = ~n41715 & ~n23440;
  assign n23443 = ~n23439 & ~n23440;
  assign n23444 = ~n23442 & ~n23443;
  assign n23445 = ~n23440 & ~n23441;
  assign n23446 = n23015 & ~n41800;
  assign n23447 = ~n23015 & n41800;
  assign n23448 = ~n23446 & ~n23447;
  assign n23449 = ~n22476 & ~n22920;
  assign n23450 = n563 & n15111;
  assign n23451 = pi122  & n37482;
  assign n23452 = pi124  & n578;
  assign n23453 = pi123  & n580;
  assign n23454 = ~n23452 & ~n23453;
  assign n23455 = ~n23451 & ~n23453;
  assign n23456 = ~n23452 & n23455;
  assign n23457 = ~n23451 & n23454;
  assign n23458 = ~n23450 & n41801;
  assign n23459 = pi14  & ~n23458;
  assign n23460 = pi14  & ~n23459;
  assign n23461 = pi14  & n23458;
  assign n23462 = ~n23458 & ~n23459;
  assign n23463 = ~pi14  & ~n23458;
  assign n23464 = ~n41802 & ~n41803;
  assign n23465 = ~n23449 & ~n23464;
  assign n23466 = n23449 & n23464;
  assign n23467 = ~n23449 & n23464;
  assign n23468 = n23449 & ~n23464;
  assign n23469 = ~n23467 & ~n23468;
  assign n23470 = ~n23465 & ~n23466;
  assign n23471 = ~n23447 & ~n41804;
  assign n23472 = ~n23446 & n23471;
  assign n23473 = n23448 & ~n41804;
  assign n23474 = ~n23448 & n41804;
  assign n23475 = ~n41804 & ~n41805;
  assign n23476 = ~n23447 & ~n41805;
  assign n23477 = ~n23446 & n23476;
  assign n23478 = n23448 & ~n41805;
  assign n23479 = ~n23475 & ~n41806;
  assign n23480 = ~n41805 & ~n23474;
  assign n23481 = ~n22942 & ~n22950;
  assign n23482 = n269 & n40885;
  assign n23483 = pi125  & n37475;
  assign n23484 = pi127  & n536;
  assign n23485 = pi126  & n538;
  assign n23486 = ~n23484 & ~n23485;
  assign n23487 = ~n23483 & ~n23485;
  assign n23488 = ~n23484 & n23487;
  assign n23489 = ~n23483 & n23486;
  assign n23490 = ~n23482 & n41808;
  assign n23491 = pi11  & ~n23490;
  assign n23492 = pi11  & ~n23491;
  assign n23493 = pi11  & n23490;
  assign n23494 = ~n23490 & ~n23491;
  assign n23495 = ~pi11  & ~n23490;
  assign n23496 = ~n41809 & ~n41810;
  assign n23497 = ~n23481 & ~n23496;
  assign n23498 = n23481 & n23496;
  assign n23499 = ~n23481 & ~n23497;
  assign n23500 = ~n23481 & n23496;
  assign n23501 = ~n23496 & ~n23497;
  assign n23502 = n23481 & ~n23496;
  assign n23503 = ~n41811 & ~n41812;
  assign n23504 = ~n23497 & ~n23498;
  assign n23505 = ~n41807 & ~n41813;
  assign n23506 = n41807 & n41813;
  assign n23507 = n41807 & ~n41813;
  assign n23508 = ~n41807 & n41813;
  assign n23509 = ~n23507 & ~n23508;
  assign n23510 = ~n23505 & ~n23506;
  assign n23511 = ~n22994 & ~n41814;
  assign n23512 = n22994 & n41814;
  assign n23513 = ~n22994 & ~n23511;
  assign n23514 = ~n41814 & ~n23511;
  assign n23515 = ~n23513 & ~n23514;
  assign n23516 = ~n23511 & ~n23512;
  assign n23517 = ~n22993 & ~n41815;
  assign n23518 = n22993 & ~n23514;
  assign n23519 = ~n23513 & n23518;
  assign n23520 = n22993 & n41815;
  assign po72  = ~n23517 & ~n41816;
  assign n23522 = ~n23511 & ~n23517;
  assign n23523 = ~n23497 & ~n23505;
  assign n23524 = n563 & n15068;
  assign n23525 = pi123  & n37482;
  assign n23526 = pi125  & n578;
  assign n23527 = pi124  & n580;
  assign n23528 = ~n23526 & ~n23527;
  assign n23529 = ~n23525 & ~n23527;
  assign n23530 = ~n23526 & n23529;
  assign n23531 = ~n23525 & n23528;
  assign n23532 = ~n23524 & n41817;
  assign n23533 = pi14  & ~n23532;
  assign n23534 = pi14  & ~n23533;
  assign n23535 = pi14  & n23532;
  assign n23536 = ~n23532 & ~n23533;
  assign n23537 = ~pi14  & ~n23532;
  assign n23538 = ~n41818 & ~n41819;
  assign n23539 = ~n23014 & ~n23446;
  assign n23540 = ~n23538 & ~n23539;
  assign n23541 = n23538 & n23539;
  assign n23542 = ~n23538 & ~n23540;
  assign n23543 = ~n23538 & n23539;
  assign n23544 = ~n23539 & ~n23540;
  assign n23545 = n23538 & ~n23539;
  assign n23546 = ~n41820 & ~n41821;
  assign n23547 = ~n23540 & ~n23541;
  assign n23548 = n6785 & n13027;
  assign n23549 = pi117  & n38631;
  assign n23550 = pi119  & n6800;
  assign n23551 = pi118  & n6802;
  assign n23552 = ~n23550 & ~n23551;
  assign n23553 = ~n23549 & ~n23551;
  assign n23554 = ~n23550 & n23553;
  assign n23555 = ~n23549 & n23552;
  assign n23556 = ~n23548 & n41823;
  assign n23557 = pi20  & ~n23556;
  assign n23558 = pi20  & ~n23557;
  assign n23559 = pi20  & n23556;
  assign n23560 = ~n23556 & ~n23557;
  assign n23561 = ~pi20  & ~n23556;
  assign n23562 = ~n41824 & ~n41825;
  assign n23563 = ~n23056 & n41797;
  assign n23564 = ~n23056 & ~n23434;
  assign n23565 = ~n23057 & ~n23563;
  assign n23566 = n23562 & n41826;
  assign n23567 = ~n23562 & ~n41826;
  assign n23568 = ~n23566 & ~n23567;
  assign n23569 = n5576 & n12530;
  assign n23570 = pi114  & n38406;
  assign n23571 = pi116  & n5591;
  assign n23572 = pi115  & n5593;
  assign n23573 = ~n23571 & ~n23572;
  assign n23574 = ~n23570 & ~n23572;
  assign n23575 = ~n23571 & n23574;
  assign n23576 = ~n23570 & n23573;
  assign n23577 = ~n23569 & n41827;
  assign n23578 = pi23  & ~n23577;
  assign n23579 = pi23  & ~n23578;
  assign n23580 = pi23  & n23577;
  assign n23581 = ~n23577 & ~n23578;
  assign n23582 = ~pi23  & ~n23577;
  assign n23583 = ~n41828 & ~n41829;
  assign n23584 = ~n23076 & ~n23428;
  assign n23585 = n23583 & n23584;
  assign n23586 = ~n23583 & ~n23584;
  assign n23587 = ~n23585 & ~n23586;
  assign n23588 = ~n23406 & ~n23414;
  assign n23589 = n607 & n9678;
  assign n23590 = pi108  & n37489;
  assign n23591 = pi110  & n620;
  assign n23592 = pi109  & n622;
  assign n23593 = ~n23591 & ~n23592;
  assign n23594 = ~n23590 & ~n23592;
  assign n23595 = ~n23591 & n23594;
  assign n23596 = ~n23590 & n23593;
  assign n23597 = ~n607 & n41830;
  assign n23598 = ~n9678 & n41830;
  assign n23599 = ~n23597 & ~n23598;
  assign n23600 = ~n23589 & n41830;
  assign n23601 = pi29  & ~n41831;
  assign n23602 = ~pi29  & n41831;
  assign n23603 = ~n23601 & ~n23602;
  assign n23604 = ~n23588 & ~n23603;
  assign n23605 = n23588 & n23603;
  assign n23606 = ~n23588 & ~n23604;
  assign n23607 = ~n23588 & n23603;
  assign n23608 = ~n23603 & ~n23604;
  assign n23609 = n23588 & ~n23603;
  assign n23610 = ~n41832 & ~n41833;
  assign n23611 = ~n23604 & ~n23605;
  assign n23612 = n649 & n8177;
  assign n23613 = pi105  & n37496;
  assign n23614 = pi107  & n662;
  assign n23615 = pi106  & n664;
  assign n23616 = ~n23614 & ~n23615;
  assign n23617 = ~n23613 & ~n23615;
  assign n23618 = ~n23614 & n23617;
  assign n23619 = ~n23613 & n23616;
  assign n23620 = ~n23612 & n41835;
  assign n23621 = pi32  & ~n23620;
  assign n23622 = pi32  & ~n23621;
  assign n23623 = pi32  & n23620;
  assign n23624 = ~n23620 & ~n23621;
  assign n23625 = ~pi32  & ~n23620;
  assign n23626 = ~n41836 & ~n41837;
  assign n23627 = ~n23376 & ~n23384;
  assign n23628 = n23626 & n23627;
  assign n23629 = ~n23626 & ~n23627;
  assign n23630 = ~n23628 & ~n23629;
  assign n23631 = n2104 & n8136;
  assign n23632 = pi102  & n37758;
  assign n23633 = pi104  & n2117;
  assign n23634 = pi103  & n2119;
  assign n23635 = ~n23633 & ~n23634;
  assign n23636 = ~n23632 & ~n23634;
  assign n23637 = ~n23633 & n23636;
  assign n23638 = ~n23632 & n23635;
  assign n23639 = ~n23631 & n41838;
  assign n23640 = pi35  & ~n23639;
  assign n23641 = pi35  & ~n23640;
  assign n23642 = pi35  & n23639;
  assign n23643 = ~n23639 & ~n23640;
  assign n23644 = ~pi35  & ~n23639;
  assign n23645 = ~n41839 & ~n41840;
  assign n23646 = ~n23352 & ~n23359;
  assign n23647 = n691 & n6839;
  assign n23648 = pi99  & n37503;
  assign n23649 = pi101  & n704;
  assign n23650 = pi100  & n706;
  assign n23651 = ~n23649 & ~n23650;
  assign n23652 = ~n23648 & ~n23650;
  assign n23653 = ~n23649 & n23652;
  assign n23654 = ~n23648 & n23651;
  assign n23655 = ~n23647 & n41841;
  assign n23656 = pi38  & ~n23655;
  assign n23657 = pi38  & ~n23656;
  assign n23658 = pi38  & n23655;
  assign n23659 = ~n23655 & ~n23656;
  assign n23660 = ~pi38  & ~n23655;
  assign n23661 = ~n41842 & ~n41843;
  assign n23662 = ~n23340 & ~n23346;
  assign n23663 = n733 & n5610;
  assign n23664 = pi96  & n37510;
  assign n23665 = pi98  & n746;
  assign n23666 = pi97  & n748;
  assign n23667 = ~n23665 & ~n23666;
  assign n23668 = ~n23664 & ~n23666;
  assign n23669 = ~n23665 & n23668;
  assign n23670 = ~n23664 & n23667;
  assign n23671 = ~n23663 & n41844;
  assign n23672 = pi41  & ~n23671;
  assign n23673 = pi41  & ~n23672;
  assign n23674 = pi41  & n23671;
  assign n23675 = ~n23671 & ~n23672;
  assign n23676 = ~pi41  & ~n23671;
  assign n23677 = ~n41845 & ~n41846;
  assign n23678 = ~n23295 & ~n23305;
  assign n23679 = ~n23279 & ~n23287;
  assign n23680 = ~n23268 & ~n23276;
  assign n23681 = ~n23239 & ~n23251;
  assign n23682 = ~n23218 & ~n23221;
  assign n23683 = n2063 & n7882;
  assign n23684 = pi78  & n39128;
  assign n23685 = pi80  & n7884;
  assign n23686 = pi79  & n7892;
  assign n23687 = ~n23685 & ~n23686;
  assign n23688 = ~n23684 & ~n23686;
  assign n23689 = ~n23685 & n23688;
  assign n23690 = ~n23684 & n23687;
  assign n23691 = ~n23683 & n41847;
  assign n23692 = pi59  & ~n23691;
  assign n23693 = pi59  & ~n23692;
  assign n23694 = pi59  & n23691;
  assign n23695 = ~n23691 & ~n23692;
  assign n23696 = ~pi59  & ~n23691;
  assign n23697 = ~n41848 & ~n41849;
  assign n23698 = n1596 & n12674;
  assign n23699 = pi75  & n40107;
  assign n23700 = pi77  & n12676;
  assign n23701 = pi76  & n12684;
  assign n23702 = ~n23700 & ~n23701;
  assign n23703 = ~n23699 & ~n23701;
  assign n23704 = ~n23700 & n23703;
  assign n23705 = ~n23699 & n23702;
  assign n23706 = ~n23698 & n41850;
  assign n23707 = pi62  & ~n23706;
  assign n23708 = pi62  & ~n23707;
  assign n23709 = pi62  & n23706;
  assign n23710 = ~n23706 & ~n23707;
  assign n23711 = ~pi62  & ~n23706;
  assign n23712 = ~n41851 & ~n41852;
  assign n23713 = ~n23197 & ~n23206;
  assign n23714 = pi74  & ~n40814;
  assign n23715 = pi73  & n18285;
  assign n23716 = ~n23714 & ~n23715;
  assign n23717 = ~n23713 & n23716;
  assign n23718 = n23713 & ~n23716;
  assign n23719 = n23716 & ~n23717;
  assign n23720 = n23713 & n23716;
  assign n23721 = ~n23713 & ~n23717;
  assign n23722 = ~n23713 & ~n23716;
  assign n23723 = ~n41853 & ~n41854;
  assign n23724 = ~n23717 & ~n23718;
  assign n23725 = ~n23712 & ~n41855;
  assign n23726 = n23712 & n41855;
  assign n23727 = ~n23712 & ~n23725;
  assign n23728 = ~n23712 & n41855;
  assign n23729 = ~n41855 & ~n23725;
  assign n23730 = n23712 & ~n41855;
  assign n23731 = ~n41856 & ~n41857;
  assign n23732 = ~n23725 & ~n23726;
  assign n23733 = n23196 & ~n23209;
  assign n23734 = ~n23209 & ~n23213;
  assign n23735 = ~n23210 & ~n23733;
  assign n23736 = ~n41858 & ~n41859;
  assign n23737 = n41858 & n41859;
  assign n23738 = ~n41858 & ~n23736;
  assign n23739 = ~n41859 & ~n23736;
  assign n23740 = ~n23738 & ~n23739;
  assign n23741 = ~n23736 & ~n23737;
  assign n23742 = n23697 & n41860;
  assign n23743 = ~n23697 & ~n41860;
  assign n23744 = ~n41860 & ~n23743;
  assign n23745 = ~n23697 & ~n23743;
  assign n23746 = ~n23744 & ~n23745;
  assign n23747 = ~n23742 & ~n23743;
  assign n23748 = n23682 & n41861;
  assign n23749 = ~n23682 & ~n41861;
  assign n23750 = ~n23748 & ~n23749;
  assign n23751 = n2091 & n4312;
  assign n23752 = pi81  & n38376;
  assign n23753 = pi83  & n4314;
  assign n23754 = pi82  & n4322;
  assign n23755 = ~n23753 & ~n23754;
  assign n23756 = ~n23752 & ~n23754;
  assign n23757 = ~n23753 & n23756;
  assign n23758 = ~n23752 & n23755;
  assign n23759 = ~n23751 & n41862;
  assign n23760 = pi56  & ~n23759;
  assign n23761 = pi56  & ~n23760;
  assign n23762 = pi56  & n23759;
  assign n23763 = ~n23759 & ~n23760;
  assign n23764 = ~pi56  & ~n23759;
  assign n23765 = ~n41863 & ~n41864;
  assign n23766 = ~n23750 & n23765;
  assign n23767 = n23750 & ~n23765;
  assign n23768 = n23750 & ~n23767;
  assign n23769 = ~n23765 & ~n23767;
  assign n23770 = ~n23768 & ~n23769;
  assign n23771 = ~n23766 & ~n23767;
  assign n23772 = n23681 & n41865;
  assign n23773 = ~n23681 & ~n41865;
  assign n23774 = ~n23772 & ~n23773;
  assign n23775 = n1971 & n2779;
  assign n23776 = pi84  & n37864;
  assign n23777 = pi86  & n1973;
  assign n23778 = pi85  & n1981;
  assign n23779 = ~n23777 & ~n23778;
  assign n23780 = ~n23776 & ~n23778;
  assign n23781 = ~n23777 & n23780;
  assign n23782 = ~n23776 & n23779;
  assign n23783 = ~n23775 & n41866;
  assign n23784 = pi53  & ~n23783;
  assign n23785 = pi53  & ~n23784;
  assign n23786 = pi53  & n23783;
  assign n23787 = ~n23783 & ~n23784;
  assign n23788 = ~pi53  & ~n23783;
  assign n23789 = ~n41867 & ~n41868;
  assign n23790 = n23774 & ~n23789;
  assign n23791 = ~n23774 & n23789;
  assign n23792 = n23774 & ~n23790;
  assign n23793 = ~n23789 & ~n23790;
  assign n23794 = ~n23792 & ~n23793;
  assign n23795 = ~n23790 & ~n23791;
  assign n23796 = n23680 & n41869;
  assign n23797 = ~n23680 & ~n41869;
  assign n23798 = ~n23796 & ~n23797;
  assign n23799 = n894 & n3591;
  assign n23800 = pi87  & n37580;
  assign n23801 = pi89  & n896;
  assign n23802 = pi88  & n904;
  assign n23803 = ~n23801 & ~n23802;
  assign n23804 = ~n23800 & ~n23802;
  assign n23805 = ~n23801 & n23804;
  assign n23806 = ~n23800 & n23803;
  assign n23807 = ~n23799 & n41870;
  assign n23808 = pi50  & ~n23807;
  assign n23809 = pi50  & ~n23808;
  assign n23810 = pi50  & n23807;
  assign n23811 = ~n23807 & ~n23808;
  assign n23812 = ~pi50  & ~n23807;
  assign n23813 = ~n41871 & ~n41872;
  assign n23814 = ~n23798 & n23813;
  assign n23815 = n23798 & ~n23813;
  assign n23816 = n23798 & ~n23815;
  assign n23817 = ~n23813 & ~n23815;
  assign n23818 = ~n23816 & ~n23817;
  assign n23819 = ~n23814 & ~n23815;
  assign n23820 = n23679 & n41873;
  assign n23821 = ~n23679 & ~n41873;
  assign n23822 = ~n23820 & ~n23821;
  assign n23823 = n785 & n4453;
  assign n23824 = pi90  & n37520;
  assign n23825 = pi92  & n787;
  assign n23826 = pi91  & n795;
  assign n23827 = ~n23825 & ~n23826;
  assign n23828 = ~n23824 & ~n23826;
  assign n23829 = ~n23825 & n23828;
  assign n23830 = ~n23824 & n23827;
  assign n23831 = ~n23823 & n41874;
  assign n23832 = pi47  & ~n23831;
  assign n23833 = pi47  & ~n23832;
  assign n23834 = pi47  & n23831;
  assign n23835 = ~n23831 & ~n23832;
  assign n23836 = ~pi47  & ~n23831;
  assign n23837 = ~n41875 & ~n41876;
  assign n23838 = n23822 & ~n23837;
  assign n23839 = ~n23822 & n23837;
  assign n23840 = n23822 & ~n23838;
  assign n23841 = ~n23837 & ~n23838;
  assign n23842 = ~n23840 & ~n23841;
  assign n23843 = ~n23838 & ~n23839;
  assign n23844 = n23678 & n41877;
  assign n23845 = ~n23678 & ~n41877;
  assign n23846 = ~n23844 & ~n23845;
  assign n23847 = n940 & n4494;
  assign n23848 = pi93  & n37541;
  assign n23849 = pi95  & n953;
  assign n23850 = pi94  & n955;
  assign n23851 = ~n23849 & ~n23850;
  assign n23852 = ~n23848 & ~n23850;
  assign n23853 = ~n23849 & n23852;
  assign n23854 = ~n23848 & n23851;
  assign n23855 = ~n23847 & n41878;
  assign n23856 = pi44  & ~n23855;
  assign n23857 = pi44  & ~n23856;
  assign n23858 = pi44  & n23855;
  assign n23859 = ~n23855 & ~n23856;
  assign n23860 = ~pi44  & ~n23855;
  assign n23861 = ~n41879 & ~n41880;
  assign n23862 = ~n23846 & n23861;
  assign n23863 = n23846 & ~n23861;
  assign n23864 = ~n23862 & ~n23863;
  assign n23865 = ~n41774 & n23864;
  assign n23866 = n41774 & ~n23864;
  assign n23867 = ~n23865 & ~n23866;
  assign n23868 = ~n23677 & n23867;
  assign n23869 = n23677 & ~n23867;
  assign n23870 = ~n23868 & ~n23869;
  assign n23871 = ~n23662 & n23870;
  assign n23872 = n23662 & ~n23870;
  assign n23873 = ~n23662 & ~n23871;
  assign n23874 = n23870 & ~n23871;
  assign n23875 = ~n23873 & ~n23874;
  assign n23876 = ~n23871 & ~n23872;
  assign n23877 = ~n23661 & ~n41881;
  assign n23878 = n23661 & ~n23874;
  assign n23879 = ~n23873 & n23878;
  assign n23880 = n23661 & n41881;
  assign n23881 = ~n23877 & ~n41882;
  assign n23882 = ~n23646 & n23881;
  assign n23883 = n23646 & ~n23881;
  assign n23884 = ~n23646 & ~n23882;
  assign n23885 = n23881 & ~n23882;
  assign n23886 = ~n23884 & ~n23885;
  assign n23887 = ~n23882 & ~n23883;
  assign n23888 = n23645 & n41883;
  assign n23889 = ~n23645 & ~n41883;
  assign n23890 = ~n23645 & ~n23889;
  assign n23891 = ~n41883 & ~n23889;
  assign n23892 = ~n23890 & ~n23891;
  assign n23893 = ~n23888 & ~n23889;
  assign n23894 = n23630 & ~n41884;
  assign n23895 = ~n23630 & n41884;
  assign n23896 = n23630 & ~n23894;
  assign n23897 = ~n41884 & ~n23894;
  assign n23898 = ~n23896 & ~n23897;
  assign n23899 = ~n23894 & ~n23895;
  assign n23900 = ~n41834 & ~n41885;
  assign n23901 = n41834 & n41885;
  assign n23902 = ~n41885 & ~n23900;
  assign n23903 = ~n41834 & ~n23900;
  assign n23904 = ~n23902 & ~n23903;
  assign n23905 = ~n23900 & ~n23901;
  assign n23906 = n4492 & n11276;
  assign n23907 = pi111  & n38208;
  assign n23908 = pi113  & n4507;
  assign n23909 = pi112  & n4509;
  assign n23910 = ~n23908 & ~n23909;
  assign n23911 = ~n23907 & ~n23909;
  assign n23912 = ~n23908 & n23911;
  assign n23913 = ~n23907 & n23910;
  assign n23914 = ~n23906 & n41887;
  assign n23915 = pi26  & ~n23914;
  assign n23916 = pi26  & ~n23915;
  assign n23917 = pi26  & n23914;
  assign n23918 = ~n23914 & ~n23915;
  assign n23919 = ~pi26  & ~n23914;
  assign n23920 = ~n41888 & ~n41889;
  assign n23921 = ~n23094 & ~n23422;
  assign n23922 = ~n23920 & ~n23921;
  assign n23923 = n23920 & n23921;
  assign n23924 = ~n23920 & ~n23922;
  assign n23925 = ~n23920 & n23921;
  assign n23926 = ~n23921 & ~n23922;
  assign n23927 = n23920 & ~n23921;
  assign n23928 = ~n41890 & ~n41891;
  assign n23929 = ~n23922 & ~n23923;
  assign n23930 = ~n41886 & ~n41892;
  assign n23931 = n41886 & n41892;
  assign n23932 = ~n41892 & ~n23930;
  assign n23933 = ~n41886 & ~n23930;
  assign n23934 = ~n23932 & ~n23933;
  assign n23935 = ~n23930 & ~n23931;
  assign n23936 = n23587 & ~n41893;
  assign n23937 = ~n23587 & n41893;
  assign n23938 = ~n23936 & ~n23937;
  assign n23939 = n23568 & ~n23937;
  assign n23940 = ~n23936 & n23939;
  assign n23941 = n23568 & n23938;
  assign n23942 = ~n23568 & ~n23938;
  assign n23943 = n23568 & ~n41894;
  assign n23944 = ~n23937 & ~n41894;
  assign n23945 = ~n23936 & n23944;
  assign n23946 = n23938 & ~n41894;
  assign n23947 = ~n23943 & ~n41895;
  assign n23948 = ~n41894 & ~n23942;
  assign n23949 = ~n23032 & ~n23440;
  assign n23950 = n8175 & n15049;
  assign n23951 = pi120  & n38895;
  assign n23952 = pi122  & n8190;
  assign n23953 = pi121  & n8192;
  assign n23954 = ~n23952 & ~n23953;
  assign n23955 = ~n23951 & ~n23953;
  assign n23956 = ~n23952 & n23955;
  assign n23957 = ~n23951 & n23954;
  assign n23958 = ~n8175 & n41897;
  assign n23959 = ~n15049 & n41897;
  assign n23960 = ~n23958 & ~n23959;
  assign n23961 = ~n23950 & n41897;
  assign n23962 = pi17  & ~n41898;
  assign n23963 = ~pi17  & n41898;
  assign n23964 = ~n23962 & ~n23963;
  assign n23965 = ~n23949 & ~n23964;
  assign n23966 = n23949 & n23964;
  assign n23967 = ~n23949 & ~n23965;
  assign n23968 = ~n23949 & n23964;
  assign n23969 = ~n23964 & ~n23965;
  assign n23970 = n23949 & ~n23964;
  assign n23971 = ~n41899 & ~n41900;
  assign n23972 = ~n23965 & ~n23966;
  assign n23973 = ~n41896 & ~n41901;
  assign n23974 = n41896 & n41901;
  assign n23975 = ~n41896 & ~n23973;
  assign n23976 = ~n41896 & n41901;
  assign n23977 = ~n41901 & ~n23973;
  assign n23978 = n41896 & ~n41901;
  assign n23979 = ~n41902 & ~n41903;
  assign n23980 = ~n23973 & ~n23974;
  assign n23981 = ~n41822 & ~n41904;
  assign n23982 = n41822 & n41904;
  assign n23983 = ~n41822 & ~n23981;
  assign n23984 = ~n41904 & ~n23981;
  assign n23985 = ~n23983 & ~n23984;
  assign n23986 = ~n23981 & ~n23982;
  assign n23987 = ~n23465 & ~n41805;
  assign n23988 = n269 & n40891;
  assign n23989 = pi126  & n37475;
  assign n23990 = pi127  & n538;
  assign n23991 = ~n23989 & ~n23990;
  assign n23992 = ~n269 & n23991;
  assign n23993 = ~n40891 & n23991;
  assign n23994 = ~n23992 & ~n23993;
  assign n23995 = ~n23988 & n23991;
  assign n23996 = pi11  & ~n41906;
  assign n23997 = ~pi11  & n41906;
  assign n23998 = ~n23996 & ~n23997;
  assign n23999 = ~n23987 & ~n23998;
  assign n24000 = n23987 & n23998;
  assign n24001 = ~n23987 & ~n23999;
  assign n24002 = ~n23987 & n23998;
  assign n24003 = ~n23998 & ~n23999;
  assign n24004 = n23987 & ~n23998;
  assign n24005 = ~n41907 & ~n41908;
  assign n24006 = ~n23999 & ~n24000;
  assign n24007 = ~n41905 & ~n41909;
  assign n24008 = n41905 & ~n41908;
  assign n24009 = ~n41907 & n24008;
  assign n24010 = n41905 & ~n41907;
  assign n24011 = ~n41908 & n24010;
  assign n24012 = n41905 & n41909;
  assign n24013 = ~n24007 & ~n41910;
  assign n24014 = ~n23523 & n24013;
  assign n24015 = n23523 & ~n24013;
  assign n24016 = ~n23523 & ~n24014;
  assign n24017 = n24013 & ~n24014;
  assign n24018 = ~n24016 & ~n24017;
  assign n24019 = ~n24014 & ~n24015;
  assign n24020 = ~n23522 & ~n41911;
  assign n24021 = n23522 & ~n24017;
  assign n24022 = ~n24016 & n24021;
  assign n24023 = n23522 & n41911;
  assign po73  = ~n24020 & ~n41912;
  assign n24025 = ~n24014 & ~n24020;
  assign n24026 = ~n23999 & ~n24007;
  assign n24027 = ~n23965 & ~n23973;
  assign n24028 = n563 & n15021;
  assign n24029 = pi124  & n37482;
  assign n24030 = pi126  & n578;
  assign n24031 = pi125  & n580;
  assign n24032 = ~n24030 & ~n24031;
  assign n24033 = ~n24029 & ~n24031;
  assign n24034 = ~n24030 & n24033;
  assign n24035 = ~n24029 & n24032;
  assign n24036 = ~n563 & n41913;
  assign n24037 = ~n15021 & n41913;
  assign n24038 = ~n24036 & ~n24037;
  assign n24039 = ~n24028 & n41913;
  assign n24040 = pi14  & ~n41914;
  assign n24041 = ~pi14  & n41914;
  assign n24042 = ~n24040 & ~n24041;
  assign n24043 = ~n24027 & ~n24042;
  assign n24044 = n24027 & n24042;
  assign n24045 = ~n24043 & ~n24044;
  assign n24046 = n8175 & n14961;
  assign n24047 = pi121  & n38895;
  assign n24048 = pi123  & n8190;
  assign n24049 = pi122  & n8192;
  assign n24050 = ~n24048 & ~n24049;
  assign n24051 = ~n24047 & ~n24049;
  assign n24052 = ~n24048 & n24051;
  assign n24053 = ~n24047 & n24050;
  assign n24054 = ~n24046 & n41915;
  assign n24055 = pi17  & ~n24054;
  assign n24056 = pi17  & ~n24055;
  assign n24057 = pi17  & n24054;
  assign n24058 = ~n24054 & ~n24055;
  assign n24059 = ~pi17  & ~n24054;
  assign n24060 = ~n41916 & ~n41917;
  assign n24061 = ~n23567 & ~n41894;
  assign n24062 = n24060 & n24061;
  assign n24063 = ~n24060 & ~n24061;
  assign n24064 = ~n24062 & ~n24063;
  assign n24065 = n6785 & n14913;
  assign n24066 = pi118  & n38631;
  assign n24067 = pi120  & n6800;
  assign n24068 = pi119  & n6802;
  assign n24069 = ~n24067 & ~n24068;
  assign n24070 = ~n24066 & ~n24068;
  assign n24071 = ~n24067 & n24070;
  assign n24072 = ~n24066 & n24069;
  assign n24073 = ~n24065 & n41918;
  assign n24074 = pi20  & ~n24073;
  assign n24075 = pi20  & ~n24074;
  assign n24076 = pi20  & n24073;
  assign n24077 = ~n24073 & ~n24074;
  assign n24078 = ~pi20  & ~n24073;
  assign n24079 = ~n41919 & ~n41920;
  assign n24080 = ~n23586 & ~n23936;
  assign n24081 = ~n24079 & ~n24080;
  assign n24082 = n24079 & n24080;
  assign n24083 = ~n24079 & ~n24081;
  assign n24084 = ~n24079 & n24080;
  assign n24085 = ~n24080 & ~n24081;
  assign n24086 = n24079 & ~n24080;
  assign n24087 = ~n41921 & ~n41922;
  assign n24088 = ~n24081 & ~n24082;
  assign n24089 = ~n23604 & ~n23900;
  assign n24090 = n4492 & n11258;
  assign n24091 = pi112  & n38208;
  assign n24092 = pi114  & n4507;
  assign n24093 = pi113  & n4509;
  assign n24094 = ~n24092 & ~n24093;
  assign n24095 = ~n24091 & ~n24093;
  assign n24096 = ~n24092 & n24095;
  assign n24097 = ~n24091 & n24094;
  assign n24098 = ~n4492 & n41924;
  assign n24099 = ~n11258 & n41924;
  assign n24100 = ~n24098 & ~n24099;
  assign n24101 = ~n24090 & n41924;
  assign n24102 = pi26  & ~n41925;
  assign n24103 = ~pi26  & n41925;
  assign n24104 = ~n24102 & ~n24103;
  assign n24105 = ~n24089 & ~n24104;
  assign n24106 = n24089 & n24104;
  assign n24107 = ~n24105 & ~n24106;
  assign n24108 = n565 & n607;
  assign n24109 = pi109  & n37489;
  assign n24110 = pi111  & n620;
  assign n24111 = pi110  & n622;
  assign n24112 = ~n24110 & ~n24111;
  assign n24113 = ~n24109 & ~n24111;
  assign n24114 = ~n24110 & n24113;
  assign n24115 = ~n24109 & n24112;
  assign n24116 = ~n24108 & n41926;
  assign n24117 = pi29  & ~n24116;
  assign n24118 = pi29  & ~n24117;
  assign n24119 = pi29  & n24116;
  assign n24120 = ~n24116 & ~n24117;
  assign n24121 = ~pi29  & ~n24116;
  assign n24122 = ~n41927 & ~n41928;
  assign n24123 = ~n23629 & n41884;
  assign n24124 = ~n23629 & ~n23894;
  assign n24125 = ~n23628 & ~n24123;
  assign n24126 = n24122 & n41929;
  assign n24127 = ~n24122 & ~n41929;
  assign n24128 = ~n24126 & ~n24127;
  assign n24129 = n649 & n9277;
  assign n24130 = pi106  & n37496;
  assign n24131 = pi108  & n662;
  assign n24132 = pi107  & n664;
  assign n24133 = ~n24131 & ~n24132;
  assign n24134 = ~n24130 & ~n24132;
  assign n24135 = ~n24131 & n24134;
  assign n24136 = ~n24130 & n24133;
  assign n24137 = ~n649 & n41930;
  assign n24138 = ~n9277 & n41930;
  assign n24139 = ~n24137 & ~n24138;
  assign n24140 = ~n24129 & n41930;
  assign n24141 = pi32  & ~n41931;
  assign n24142 = ~pi32  & n41931;
  assign n24143 = ~n24141 & ~n24142;
  assign n24144 = n23645 & ~n23882;
  assign n24145 = ~n23882 & ~n23889;
  assign n24146 = ~n23883 & ~n24144;
  assign n24147 = ~n24143 & ~n41932;
  assign n24148 = n24143 & n41932;
  assign n24149 = ~n24147 & ~n24148;
  assign n24150 = n2104 & n8229;
  assign n24151 = pi103  & n37758;
  assign n24152 = pi105  & n2117;
  assign n24153 = pi104  & n2119;
  assign n24154 = ~n24152 & ~n24153;
  assign n24155 = ~n24151 & ~n24153;
  assign n24156 = ~n24152 & n24155;
  assign n24157 = ~n24151 & n24154;
  assign n24158 = ~n24150 & n41933;
  assign n24159 = pi35  & ~n24158;
  assign n24160 = pi35  & ~n24159;
  assign n24161 = pi35  & n24158;
  assign n24162 = ~n24158 & ~n24159;
  assign n24163 = ~pi35  & ~n24158;
  assign n24164 = ~n41934 & ~n41935;
  assign n24165 = ~n23871 & ~n23877;
  assign n24166 = ~n23865 & ~n23868;
  assign n24167 = n894 & n3566;
  assign n24168 = pi88  & n37580;
  assign n24169 = pi90  & n896;
  assign n24170 = pi89  & n904;
  assign n24171 = ~n24169 & ~n24170;
  assign n24172 = ~n24168 & ~n24170;
  assign n24173 = ~n24169 & n24172;
  assign n24174 = ~n24168 & n24171;
  assign n24175 = ~n24167 & n41936;
  assign n24176 = pi50  & ~n24175;
  assign n24177 = pi50  & ~n24176;
  assign n24178 = pi50  & n24175;
  assign n24179 = ~n24175 & ~n24176;
  assign n24180 = ~pi50  & ~n24175;
  assign n24181 = ~n41937 & ~n41938;
  assign n24182 = n636 & n1971;
  assign n24183 = pi85  & n37864;
  assign n24184 = pi87  & n1973;
  assign n24185 = pi86  & n1981;
  assign n24186 = ~n24184 & ~n24185;
  assign n24187 = ~n24183 & ~n24185;
  assign n24188 = ~n24184 & n24187;
  assign n24189 = ~n24183 & n24186;
  assign n24190 = ~n24182 & n41939;
  assign n24191 = pi53  & ~n24190;
  assign n24192 = pi53  & ~n24191;
  assign n24193 = pi53  & n24190;
  assign n24194 = ~n24190 & ~n24191;
  assign n24195 = ~pi53  & ~n24190;
  assign n24196 = ~n41940 & ~n41941;
  assign n24197 = n2154 & n7882;
  assign n24198 = pi79  & n39128;
  assign n24199 = pi81  & n7884;
  assign n24200 = pi80  & n7892;
  assign n24201 = ~n24199 & ~n24200;
  assign n24202 = ~n24198 & ~n24200;
  assign n24203 = ~n24199 & n24202;
  assign n24204 = ~n24198 & n24201;
  assign n24205 = ~n24197 & n41942;
  assign n24206 = pi59  & ~n24205;
  assign n24207 = pi59  & ~n24206;
  assign n24208 = pi59  & n24205;
  assign n24209 = ~n24205 & ~n24206;
  assign n24210 = ~pi59  & ~n24205;
  assign n24211 = ~n41943 & ~n41944;
  assign n24212 = n1578 & n12674;
  assign n24213 = pi76  & n40107;
  assign n24214 = pi78  & n12676;
  assign n24215 = pi77  & n12684;
  assign n24216 = ~n24214 & ~n24215;
  assign n24217 = ~n24213 & ~n24215;
  assign n24218 = ~n24214 & n24217;
  assign n24219 = ~n24213 & n24216;
  assign n24220 = ~n24212 & n41945;
  assign n24221 = pi62  & ~n24220;
  assign n24222 = pi62  & ~n24221;
  assign n24223 = pi62  & n24220;
  assign n24224 = ~n24220 & ~n24221;
  assign n24225 = ~pi62  & ~n24220;
  assign n24226 = ~n41946 & ~n41947;
  assign n24227 = ~n23717 & ~n23725;
  assign n24228 = pi75  & ~n40814;
  assign n24229 = pi74  & n18285;
  assign n24230 = ~n24228 & ~n24229;
  assign n24231 = n23716 & ~n24230;
  assign n24232 = ~n23716 & n24230;
  assign n24233 = n23716 & ~n24231;
  assign n24234 = n23716 & n24230;
  assign n24235 = ~n24230 & ~n24231;
  assign n24236 = ~n23716 & ~n24230;
  assign n24237 = ~n41948 & ~n41949;
  assign n24238 = ~n24231 & ~n24232;
  assign n24239 = ~n24227 & ~n41950;
  assign n24240 = n24227 & n41950;
  assign n24241 = ~n24227 & ~n24239;
  assign n24242 = ~n24227 & n41950;
  assign n24243 = ~n41950 & ~n24239;
  assign n24244 = n24227 & ~n41950;
  assign n24245 = ~n41951 & ~n41952;
  assign n24246 = ~n24239 & ~n24240;
  assign n24247 = ~n24226 & ~n41953;
  assign n24248 = n24226 & n41953;
  assign n24249 = ~n41953 & ~n24247;
  assign n24250 = ~n24226 & ~n24247;
  assign n24251 = ~n24249 & ~n24250;
  assign n24252 = ~n24247 & ~n24248;
  assign n24253 = n24211 & n41954;
  assign n24254 = ~n24211 & ~n41954;
  assign n24255 = ~n41954 & ~n24254;
  assign n24256 = ~n24211 & ~n24254;
  assign n24257 = ~n24255 & ~n24256;
  assign n24258 = ~n24253 & ~n24254;
  assign n24259 = n23697 & ~n23736;
  assign n24260 = ~n23736 & ~n23743;
  assign n24261 = ~n23737 & ~n24259;
  assign n24262 = n41955 & n41956;
  assign n24263 = ~n41955 & ~n41956;
  assign n24264 = ~n24262 & ~n24263;
  assign n24265 = n2591 & n4312;
  assign n24266 = pi82  & n38376;
  assign n24267 = pi84  & n4314;
  assign n24268 = pi83  & n4322;
  assign n24269 = ~n24267 & ~n24268;
  assign n24270 = ~n24266 & ~n24268;
  assign n24271 = ~n24267 & n24270;
  assign n24272 = ~n24266 & n24269;
  assign n24273 = ~n24265 & n41957;
  assign n24274 = pi56  & ~n24273;
  assign n24275 = pi56  & ~n24274;
  assign n24276 = pi56  & n24273;
  assign n24277 = ~n24273 & ~n24274;
  assign n24278 = ~pi56  & ~n24273;
  assign n24279 = ~n41958 & ~n41959;
  assign n24280 = ~n24264 & n24279;
  assign n24281 = n24264 & ~n24279;
  assign n24282 = ~n24280 & ~n24281;
  assign n24283 = ~n23749 & n23765;
  assign n24284 = ~n23749 & ~n23767;
  assign n24285 = ~n23748 & ~n24283;
  assign n24286 = n24282 & ~n41960;
  assign n24287 = ~n24282 & n41960;
  assign n24288 = ~n41960 & ~n24286;
  assign n24289 = n24282 & ~n24286;
  assign n24290 = ~n24288 & ~n24289;
  assign n24291 = ~n24286 & ~n24287;
  assign n24292 = ~n24196 & ~n41961;
  assign n24293 = n24196 & ~n24289;
  assign n24294 = ~n24288 & n24293;
  assign n24295 = n24196 & n41961;
  assign n24296 = ~n24292 & ~n41962;
  assign n24297 = ~n23773 & n23789;
  assign n24298 = ~n23773 & ~n23790;
  assign n24299 = ~n23772 & ~n24297;
  assign n24300 = n24296 & ~n41963;
  assign n24301 = ~n24296 & n41963;
  assign n24302 = ~n24300 & ~n24301;
  assign n24303 = ~n24181 & n24302;
  assign n24304 = n24181 & ~n24302;
  assign n24305 = ~n24303 & ~n24304;
  assign n24306 = ~n23797 & n23813;
  assign n24307 = ~n23797 & ~n23815;
  assign n24308 = ~n23796 & ~n24306;
  assign n24309 = n24305 & ~n41964;
  assign n24310 = ~n24305 & n41964;
  assign n24311 = ~n24309 & ~n24310;
  assign n24312 = n785 & n4544;
  assign n24313 = pi91  & n37520;
  assign n24314 = pi93  & n787;
  assign n24315 = pi92  & n795;
  assign n24316 = ~n24314 & ~n24315;
  assign n24317 = ~n24313 & ~n24315;
  assign n24318 = ~n24314 & n24317;
  assign n24319 = ~n24313 & n24316;
  assign n24320 = ~n24312 & n41965;
  assign n24321 = pi47  & ~n24320;
  assign n24322 = pi47  & ~n24321;
  assign n24323 = pi47  & n24320;
  assign n24324 = ~n24320 & ~n24321;
  assign n24325 = ~pi47  & ~n24320;
  assign n24326 = ~n41966 & ~n41967;
  assign n24327 = n24311 & ~n24326;
  assign n24328 = ~n24311 & n24326;
  assign n24329 = n24311 & ~n24327;
  assign n24330 = ~n24326 & ~n24327;
  assign n24331 = ~n24329 & ~n24330;
  assign n24332 = ~n24327 & ~n24328;
  assign n24333 = ~n23821 & n23837;
  assign n24334 = ~n23821 & ~n23838;
  assign n24335 = ~n23820 & ~n24333;
  assign n24336 = n41968 & n41969;
  assign n24337 = ~n41968 & ~n41969;
  assign n24338 = ~n24336 & ~n24337;
  assign n24339 = n940 & n5281;
  assign n24340 = pi94  & n37541;
  assign n24341 = pi96  & n953;
  assign n24342 = pi95  & n955;
  assign n24343 = ~n24341 & ~n24342;
  assign n24344 = ~n24340 & ~n24342;
  assign n24345 = ~n24341 & n24344;
  assign n24346 = ~n24340 & n24343;
  assign n24347 = ~n24339 & n41970;
  assign n24348 = pi44  & ~n24347;
  assign n24349 = pi44  & ~n24348;
  assign n24350 = pi44  & n24347;
  assign n24351 = ~n24347 & ~n24348;
  assign n24352 = ~pi44  & ~n24347;
  assign n24353 = ~n41971 & ~n41972;
  assign n24354 = ~n24338 & n24353;
  assign n24355 = n24338 & ~n24353;
  assign n24356 = ~n24354 & ~n24355;
  assign n24357 = ~n23845 & ~n23863;
  assign n24358 = n24356 & ~n24357;
  assign n24359 = ~n24356 & n24357;
  assign n24360 = ~n24358 & ~n24359;
  assign n24361 = n733 & n5578;
  assign n24362 = pi97  & n37510;
  assign n24363 = pi99  & n746;
  assign n24364 = pi98  & n748;
  assign n24365 = ~n24363 & ~n24364;
  assign n24366 = ~n24362 & ~n24364;
  assign n24367 = ~n24363 & n24366;
  assign n24368 = ~n24362 & n24365;
  assign n24369 = ~n24361 & n41973;
  assign n24370 = pi41  & ~n24369;
  assign n24371 = pi41  & ~n24370;
  assign n24372 = pi41  & n24369;
  assign n24373 = ~n24369 & ~n24370;
  assign n24374 = ~pi41  & ~n24369;
  assign n24375 = ~n41974 & ~n41975;
  assign n24376 = ~n24360 & n24375;
  assign n24377 = n24360 & ~n24375;
  assign n24378 = n24360 & ~n24377;
  assign n24379 = ~n24375 & ~n24377;
  assign n24380 = ~n24378 & ~n24379;
  assign n24381 = ~n24376 & ~n24377;
  assign n24382 = n24166 & n41976;
  assign n24383 = ~n24166 & ~n41976;
  assign n24384 = ~n24382 & ~n24383;
  assign n24385 = n691 & n6819;
  assign n24386 = pi100  & n37503;
  assign n24387 = pi102  & n704;
  assign n24388 = pi101  & n706;
  assign n24389 = ~n24387 & ~n24388;
  assign n24390 = ~n24386 & ~n24388;
  assign n24391 = ~n24387 & n24390;
  assign n24392 = ~n24386 & n24389;
  assign n24393 = ~n24385 & n41977;
  assign n24394 = pi38  & ~n24393;
  assign n24395 = pi38  & ~n24394;
  assign n24396 = pi38  & n24393;
  assign n24397 = ~n24393 & ~n24394;
  assign n24398 = ~pi38  & ~n24393;
  assign n24399 = ~n41978 & ~n41979;
  assign n24400 = ~n24384 & n24399;
  assign n24401 = n24384 & ~n24399;
  assign n24402 = ~n24400 & ~n24401;
  assign n24403 = ~n24165 & n24402;
  assign n24404 = n24165 & ~n24402;
  assign n24405 = ~n24403 & ~n24404;
  assign n24406 = n24164 & ~n24405;
  assign n24407 = ~n24164 & n24405;
  assign n24408 = ~n24164 & ~n24407;
  assign n24409 = n24405 & ~n24407;
  assign n24410 = ~n24408 & ~n24409;
  assign n24411 = ~n24406 & ~n24407;
  assign n24412 = n24149 & ~n41980;
  assign n24413 = ~n24149 & n41980;
  assign n24414 = n24149 & ~n24412;
  assign n24415 = ~n41980 & ~n24412;
  assign n24416 = ~n24414 & ~n24415;
  assign n24417 = ~n24412 & ~n24413;
  assign n24418 = n24128 & ~n41981;
  assign n24419 = ~n24128 & n41981;
  assign n24420 = ~n24418 & ~n24419;
  assign n24421 = n24107 & ~n24419;
  assign n24422 = ~n24418 & n24421;
  assign n24423 = n24107 & n24420;
  assign n24424 = ~n24107 & ~n24420;
  assign n24425 = n24107 & ~n41982;
  assign n24426 = ~n24419 & ~n41982;
  assign n24427 = ~n24418 & n24426;
  assign n24428 = n24420 & ~n41982;
  assign n24429 = ~n24425 & ~n41983;
  assign n24430 = ~n41982 & ~n24424;
  assign n24431 = ~n23922 & ~n23930;
  assign n24432 = n5576 & n13079;
  assign n24433 = pi115  & n38406;
  assign n24434 = pi117  & n5591;
  assign n24435 = pi116  & n5593;
  assign n24436 = ~n24434 & ~n24435;
  assign n24437 = ~n24433 & ~n24435;
  assign n24438 = ~n24434 & n24437;
  assign n24439 = ~n24433 & n24436;
  assign n24440 = ~n5576 & n41985;
  assign n24441 = ~n13079 & n41985;
  assign n24442 = ~n24440 & ~n24441;
  assign n24443 = ~n24432 & n41985;
  assign n24444 = pi23  & ~n41986;
  assign n24445 = ~pi23  & n41986;
  assign n24446 = ~n24444 & ~n24445;
  assign n24447 = ~n24431 & ~n24446;
  assign n24448 = n24431 & n24446;
  assign n24449 = ~n24431 & ~n24447;
  assign n24450 = ~n24431 & n24446;
  assign n24451 = ~n24446 & ~n24447;
  assign n24452 = n24431 & ~n24446;
  assign n24453 = ~n41987 & ~n41988;
  assign n24454 = ~n24447 & ~n24448;
  assign n24455 = ~n41984 & ~n41989;
  assign n24456 = n41984 & n41989;
  assign n24457 = ~n41984 & ~n24455;
  assign n24458 = ~n41984 & n41989;
  assign n24459 = ~n41989 & ~n24455;
  assign n24460 = n41984 & ~n41989;
  assign n24461 = ~n41990 & ~n41991;
  assign n24462 = ~n24455 & ~n24456;
  assign n24463 = ~n41923 & ~n41992;
  assign n24464 = n41923 & n41992;
  assign n24465 = ~n41923 & ~n24463;
  assign n24466 = ~n41992 & ~n24463;
  assign n24467 = ~n24465 & ~n24466;
  assign n24468 = ~n24463 & ~n24464;
  assign n24469 = n24064 & ~n41993;
  assign n24470 = ~n24064 & n41993;
  assign n24471 = ~n24469 & ~n24470;
  assign n24472 = n24045 & ~n24470;
  assign n24473 = ~n24469 & n24472;
  assign n24474 = n24045 & n24471;
  assign n24475 = ~n24045 & ~n24471;
  assign n24476 = n24045 & ~n41994;
  assign n24477 = ~n24470 & ~n41994;
  assign n24478 = ~n24469 & n24477;
  assign n24479 = n24471 & ~n41994;
  assign n24480 = ~n24476 & ~n41995;
  assign n24481 = ~n41994 & ~n24475;
  assign n24482 = ~n23540 & ~n23981;
  assign n24483 = n269 & ~n18675;
  assign n24484 = ~n37475 & ~n24483;
  assign n24485 = pi127  & n37475;
  assign n24486 = n269 & n18680;
  assign n24487 = ~n24485 & ~n24486;
  assign n24488 = pi127  & ~n24484;
  assign n24489 = pi11  & ~n41997;
  assign n24490 = pi11  & ~n24489;
  assign n24491 = pi11  & n41997;
  assign n24492 = ~n41997 & ~n24489;
  assign n24493 = ~pi11  & ~n41997;
  assign n24494 = ~n41998 & ~n41999;
  assign n24495 = ~n24482 & ~n24494;
  assign n24496 = n24482 & n24494;
  assign n24497 = ~n24482 & ~n24495;
  assign n24498 = ~n24494 & ~n24495;
  assign n24499 = ~n24497 & ~n24498;
  assign n24500 = ~n24495 & ~n24496;
  assign n24501 = ~n41996 & ~n42000;
  assign n24502 = n41996 & n42000;
  assign n24503 = n41996 & ~n42000;
  assign n24504 = ~n41996 & n42000;
  assign n24505 = ~n24503 & ~n24504;
  assign n24506 = ~n24501 & ~n24502;
  assign n24507 = ~n24026 & ~n42001;
  assign n24508 = n24026 & n42001;
  assign n24509 = ~n24026 & ~n24507;
  assign n24510 = ~n42001 & ~n24507;
  assign n24511 = ~n24509 & ~n24510;
  assign n24512 = ~n24507 & ~n24508;
  assign n24513 = ~n24025 & ~n42002;
  assign n24514 = n24025 & ~n24510;
  assign n24515 = ~n24509 & n24514;
  assign n24516 = n24025 & n42002;
  assign po74  = ~n24513 & ~n42003;
  assign n24518 = ~n24507 & ~n24513;
  assign n24519 = ~n24495 & ~n24501;
  assign n24520 = n6785 & n15091;
  assign n24521 = pi119  & n38631;
  assign n24522 = pi121  & n6800;
  assign n24523 = pi120  & n6802;
  assign n24524 = ~n24522 & ~n24523;
  assign n24525 = ~n24521 & ~n24523;
  assign n24526 = ~n24522 & n24525;
  assign n24527 = ~n24521 & n24524;
  assign n24528 = ~n24520 & n42004;
  assign n24529 = pi20  & ~n24528;
  assign n24530 = pi20  & ~n24529;
  assign n24531 = pi20  & n24528;
  assign n24532 = ~n24528 & ~n24529;
  assign n24533 = ~pi20  & ~n24528;
  assign n24534 = ~n42005 & ~n42006;
  assign n24535 = ~n24081 & ~n24463;
  assign n24536 = n24534 & n24535;
  assign n24537 = ~n24534 & ~n24535;
  assign n24538 = ~n24536 & ~n24537;
  assign n24539 = n523 & n4492;
  assign n24540 = pi113  & n38208;
  assign n24541 = pi115  & n4507;
  assign n24542 = pi114  & n4509;
  assign n24543 = ~n24541 & ~n24542;
  assign n24544 = ~n24540 & ~n24542;
  assign n24545 = ~n24541 & n24544;
  assign n24546 = ~n24540 & n24543;
  assign n24547 = ~n24539 & n42007;
  assign n24548 = pi26  & ~n24547;
  assign n24549 = pi26  & ~n24548;
  assign n24550 = pi26  & n24547;
  assign n24551 = ~n24547 & ~n24548;
  assign n24552 = ~pi26  & ~n24547;
  assign n24553 = ~n42008 & ~n42009;
  assign n24554 = ~n24105 & ~n41982;
  assign n24555 = n24553 & n24554;
  assign n24556 = ~n24553 & ~n24554;
  assign n24557 = ~n24555 & ~n24556;
  assign n24558 = n2104 & n8209;
  assign n24559 = pi104  & n37758;
  assign n24560 = pi106  & n2117;
  assign n24561 = pi105  & n2119;
  assign n24562 = ~n24560 & ~n24561;
  assign n24563 = ~n24559 & ~n24561;
  assign n24564 = ~n24560 & n24563;
  assign n24565 = ~n24559 & n24562;
  assign n24566 = ~n24558 & n42010;
  assign n24567 = pi35  & ~n24566;
  assign n24568 = pi35  & ~n24567;
  assign n24569 = pi35  & n24566;
  assign n24570 = ~n24566 & ~n24567;
  assign n24571 = ~pi35  & ~n24566;
  assign n24572 = ~n42011 & ~n42012;
  assign n24573 = ~n24383 & ~n24401;
  assign n24574 = n733 & n6474;
  assign n24575 = pi98  & n37510;
  assign n24576 = pi100  & n746;
  assign n24577 = pi99  & n748;
  assign n24578 = ~n24576 & ~n24577;
  assign n24579 = ~n24575 & ~n24577;
  assign n24580 = ~n24576 & n24579;
  assign n24581 = ~n24575 & n24578;
  assign n24582 = ~n24574 & n42013;
  assign n24583 = pi41  & ~n24582;
  assign n24584 = pi41  & ~n24583;
  assign n24585 = pi41  & n24582;
  assign n24586 = ~n24582 & ~n24583;
  assign n24587 = ~pi41  & ~n24582;
  assign n24588 = ~n42014 & ~n42015;
  assign n24589 = ~n24337 & ~n24355;
  assign n24590 = n940 & n5630;
  assign n24591 = pi95  & n37541;
  assign n24592 = pi97  & n953;
  assign n24593 = pi96  & n955;
  assign n24594 = ~n24592 & ~n24593;
  assign n24595 = ~n24591 & ~n24593;
  assign n24596 = ~n24592 & n24595;
  assign n24597 = ~n24591 & n24594;
  assign n24598 = ~n24590 & n42016;
  assign n24599 = pi44  & ~n24598;
  assign n24600 = pi44  & ~n24599;
  assign n24601 = pi44  & n24598;
  assign n24602 = ~n24598 & ~n24599;
  assign n24603 = ~pi44  & ~n24598;
  assign n24604 = ~n42017 & ~n42018;
  assign n24605 = ~n24300 & ~n24303;
  assign n24606 = n594 & n894;
  assign n24607 = pi89  & n37580;
  assign n24608 = pi91  & n896;
  assign n24609 = pi90  & n904;
  assign n24610 = ~n24608 & ~n24609;
  assign n24611 = ~n24607 & ~n24609;
  assign n24612 = ~n24608 & n24611;
  assign n24613 = ~n24607 & n24610;
  assign n24614 = ~n24606 & n42019;
  assign n24615 = pi50  & ~n24614;
  assign n24616 = pi50  & ~n24615;
  assign n24617 = pi50  & n24614;
  assign n24618 = ~n24614 & ~n24615;
  assign n24619 = ~pi50  & ~n24614;
  assign n24620 = ~n42020 & ~n42021;
  assign n24621 = ~n24286 & ~n24292;
  assign n24622 = n1971 & n3354;
  assign n24623 = pi86  & n37864;
  assign n24624 = pi88  & n1973;
  assign n24625 = pi87  & n1981;
  assign n24626 = ~n24624 & ~n24625;
  assign n24627 = ~n24623 & ~n24625;
  assign n24628 = ~n24624 & n24627;
  assign n24629 = ~n24623 & n24626;
  assign n24630 = ~n24622 & n42022;
  assign n24631 = pi53  & ~n24630;
  assign n24632 = pi53  & ~n24631;
  assign n24633 = pi53  & n24630;
  assign n24634 = ~n24630 & ~n24631;
  assign n24635 = ~pi53  & ~n24630;
  assign n24636 = ~n42023 & ~n42024;
  assign n24637 = ~n24263 & ~n24281;
  assign n24638 = n2134 & n7882;
  assign n24639 = pi80  & n39128;
  assign n24640 = pi82  & n7884;
  assign n24641 = pi81  & n7892;
  assign n24642 = ~n24640 & ~n24641;
  assign n24643 = ~n24639 & ~n24641;
  assign n24644 = ~n24640 & n24643;
  assign n24645 = ~n24639 & n24642;
  assign n24646 = ~n24638 & n42025;
  assign n24647 = pi59  & ~n24646;
  assign n24648 = pi59  & ~n24647;
  assign n24649 = pi59  & n24646;
  assign n24650 = ~n24646 & ~n24647;
  assign n24651 = ~pi59  & ~n24646;
  assign n24652 = ~n42026 & ~n42027;
  assign n24653 = ~n24231 & ~n24239;
  assign n24654 = n678 & n12674;
  assign n24655 = pi77  & n40107;
  assign n24656 = pi79  & n12676;
  assign n24657 = pi78  & n12684;
  assign n24658 = ~n24656 & ~n24657;
  assign n24659 = ~n24655 & ~n24657;
  assign n24660 = ~n24656 & n24659;
  assign n24661 = ~n24655 & n24658;
  assign n24662 = ~n24654 & n42028;
  assign n24663 = pi62  & ~n24662;
  assign n24664 = pi62  & ~n24663;
  assign n24665 = pi62  & n24662;
  assign n24666 = ~n24662 & ~n24663;
  assign n24667 = ~pi62  & ~n24662;
  assign n24668 = ~n42029 & ~n42030;
  assign n24669 = ~pi11  & ~n23716;
  assign n24670 = pi11  & n23716;
  assign n24671 = pi11  & ~n23716;
  assign n24672 = ~pi11  & n23716;
  assign n24673 = ~n24671 & ~n24672;
  assign n24674 = ~n24669 & ~n24670;
  assign n24675 = pi76  & ~n40814;
  assign n24676 = pi75  & n18285;
  assign n24677 = ~n24675 & ~n24676;
  assign n24678 = ~n42031 & ~n24677;
  assign n24679 = n42031 & n24677;
  assign n24680 = ~n24678 & ~n24679;
  assign n24681 = ~n24668 & n24680;
  assign n24682 = n24668 & ~n24680;
  assign n24683 = ~n24668 & ~n24681;
  assign n24684 = ~n24668 & ~n24680;
  assign n24685 = n24680 & ~n24681;
  assign n24686 = n24668 & n24680;
  assign n24687 = ~n42032 & ~n42033;
  assign n24688 = ~n24681 & ~n24682;
  assign n24689 = ~n24653 & ~n42034;
  assign n24690 = n24653 & n42034;
  assign n24691 = ~n24653 & ~n24689;
  assign n24692 = ~n24653 & n42034;
  assign n24693 = ~n42034 & ~n24689;
  assign n24694 = n24653 & ~n42034;
  assign n24695 = ~n42035 & ~n42036;
  assign n24696 = ~n24689 & ~n24690;
  assign n24697 = ~n24652 & ~n42037;
  assign n24698 = n24652 & n42037;
  assign n24699 = ~n42037 & ~n24697;
  assign n24700 = ~n24652 & ~n24697;
  assign n24701 = ~n24699 & ~n24700;
  assign n24702 = ~n24697 & ~n24698;
  assign n24703 = n24211 & ~n24247;
  assign n24704 = ~n24247 & ~n24254;
  assign n24705 = ~n24248 & ~n24703;
  assign n24706 = n42038 & n42039;
  assign n24707 = ~n42038 & ~n42039;
  assign n24708 = ~n24706 & ~n24707;
  assign n24709 = n2804 & n4312;
  assign n24710 = pi83  & n38376;
  assign n24711 = pi85  & n4314;
  assign n24712 = pi84  & n4322;
  assign n24713 = ~n24711 & ~n24712;
  assign n24714 = ~n24710 & ~n24712;
  assign n24715 = ~n24711 & n24714;
  assign n24716 = ~n24710 & n24713;
  assign n24717 = ~n24709 & n42040;
  assign n24718 = pi56  & ~n24717;
  assign n24719 = pi56  & ~n24718;
  assign n24720 = pi56  & n24717;
  assign n24721 = ~n24717 & ~n24718;
  assign n24722 = ~pi56  & ~n24717;
  assign n24723 = ~n42041 & ~n42042;
  assign n24724 = n24708 & ~n24723;
  assign n24725 = ~n24708 & n24723;
  assign n24726 = n24708 & ~n24724;
  assign n24727 = n24708 & n24723;
  assign n24728 = ~n24723 & ~n24724;
  assign n24729 = ~n24708 & ~n24723;
  assign n24730 = ~n42043 & ~n42044;
  assign n24731 = ~n24724 & ~n24725;
  assign n24732 = ~n24637 & ~n42045;
  assign n24733 = n24637 & n42045;
  assign n24734 = ~n24732 & ~n24733;
  assign n24735 = ~n24636 & n24734;
  assign n24736 = n24636 & ~n24734;
  assign n24737 = ~n24636 & ~n24735;
  assign n24738 = ~n24636 & ~n24734;
  assign n24739 = n24734 & ~n24735;
  assign n24740 = n24636 & n24734;
  assign n24741 = ~n42046 & ~n42047;
  assign n24742 = ~n24735 & ~n24736;
  assign n24743 = ~n24621 & ~n42048;
  assign n24744 = n24621 & n42048;
  assign n24745 = ~n24621 & ~n24743;
  assign n24746 = ~n24621 & n42048;
  assign n24747 = ~n42048 & ~n24743;
  assign n24748 = n24621 & ~n42048;
  assign n24749 = ~n42049 & ~n42050;
  assign n24750 = ~n24743 & ~n24744;
  assign n24751 = ~n24620 & ~n42051;
  assign n24752 = n24620 & n42051;
  assign n24753 = ~n42051 & ~n24751;
  assign n24754 = ~n24620 & ~n24751;
  assign n24755 = ~n24753 & ~n24754;
  assign n24756 = ~n24751 & ~n24752;
  assign n24757 = n24605 & n42052;
  assign n24758 = ~n24605 & ~n42052;
  assign n24759 = ~n24757 & ~n24758;
  assign n24760 = n785 & n4524;
  assign n24761 = pi92  & n37520;
  assign n24762 = pi94  & n787;
  assign n24763 = pi93  & n795;
  assign n24764 = ~n24762 & ~n24763;
  assign n24765 = ~n24761 & ~n24763;
  assign n24766 = ~n24762 & n24765;
  assign n24767 = ~n24761 & n24764;
  assign n24768 = ~n24760 & n42053;
  assign n24769 = pi47  & ~n24768;
  assign n24770 = pi47  & ~n24769;
  assign n24771 = pi47  & n24768;
  assign n24772 = ~n24768 & ~n24769;
  assign n24773 = ~pi47  & ~n24768;
  assign n24774 = ~n42054 & ~n42055;
  assign n24775 = n24759 & ~n24774;
  assign n24776 = ~n24759 & n24774;
  assign n24777 = ~n24775 & ~n24776;
  assign n24778 = ~n24309 & n24326;
  assign n24779 = ~n24309 & ~n24327;
  assign n24780 = ~n24310 & ~n24778;
  assign n24781 = ~n24775 & n42056;
  assign n24782 = ~n24775 & ~n42056;
  assign n24783 = ~n24776 & ~n42056;
  assign n24784 = ~n24775 & n24783;
  assign n24785 = ~n24776 & n24782;
  assign n24786 = ~n24775 & ~n42057;
  assign n24787 = ~n24776 & ~n24781;
  assign n24788 = ~n24776 & n42058;
  assign n24789 = n24777 & n42056;
  assign n24790 = ~n42056 & ~n42057;
  assign n24791 = ~n24777 & ~n42056;
  assign n24792 = ~n42059 & ~n42060;
  assign n24793 = ~n24604 & ~n24792;
  assign n24794 = n24604 & n24792;
  assign n24795 = ~n24792 & ~n24793;
  assign n24796 = ~n24604 & ~n24793;
  assign n24797 = ~n24795 & ~n24796;
  assign n24798 = ~n24793 & ~n24794;
  assign n24799 = ~n24589 & ~n42061;
  assign n24800 = n24589 & n42061;
  assign n24801 = ~n24589 & n42061;
  assign n24802 = n24589 & ~n42061;
  assign n24803 = ~n24801 & ~n24802;
  assign n24804 = ~n24799 & ~n24800;
  assign n24805 = ~n24588 & ~n42062;
  assign n24806 = n24588 & n42062;
  assign n24807 = ~n24805 & ~n24806;
  assign n24808 = ~n24359 & ~n24375;
  assign n24809 = ~n24358 & ~n24377;
  assign n24810 = ~n24358 & ~n24808;
  assign n24811 = ~n24807 & n42063;
  assign n24812 = n24807 & ~n42063;
  assign n24813 = ~n24811 & ~n24812;
  assign n24814 = n691 & n6787;
  assign n24815 = pi101  & n37503;
  assign n24816 = pi103  & n704;
  assign n24817 = pi102  & n706;
  assign n24818 = ~n24816 & ~n24817;
  assign n24819 = ~n24815 & ~n24817;
  assign n24820 = ~n24816 & n24819;
  assign n24821 = ~n24815 & n24818;
  assign n24822 = ~n24814 & n42064;
  assign n24823 = pi38  & ~n24822;
  assign n24824 = pi38  & ~n24823;
  assign n24825 = pi38  & n24822;
  assign n24826 = ~n24822 & ~n24823;
  assign n24827 = ~pi38  & ~n24822;
  assign n24828 = ~n42065 & ~n42066;
  assign n24829 = n24813 & ~n24828;
  assign n24830 = ~n24813 & n24828;
  assign n24831 = n24813 & ~n24829;
  assign n24832 = n24813 & n24828;
  assign n24833 = ~n24828 & ~n24829;
  assign n24834 = ~n24813 & ~n24828;
  assign n24835 = ~n42067 & ~n42068;
  assign n24836 = ~n24829 & ~n24830;
  assign n24837 = ~n24573 & ~n42069;
  assign n24838 = n24573 & n42069;
  assign n24839 = ~n24573 & n42069;
  assign n24840 = n24573 & ~n42069;
  assign n24841 = ~n24839 & ~n24840;
  assign n24842 = ~n24837 & ~n24838;
  assign n24843 = ~n24572 & ~n42070;
  assign n24844 = n24572 & n42070;
  assign n24845 = ~n24843 & ~n24844;
  assign n24846 = n24164 & ~n24403;
  assign n24847 = ~n24403 & ~n24407;
  assign n24848 = ~n24404 & ~n24846;
  assign n24849 = ~n24845 & n42071;
  assign n24850 = n24845 & ~n42071;
  assign n24851 = ~n24849 & ~n24850;
  assign n24852 = n649 & n9701;
  assign n24853 = pi107  & n37496;
  assign n24854 = pi109  & n662;
  assign n24855 = pi108  & n664;
  assign n24856 = ~n24854 & ~n24855;
  assign n24857 = ~n24853 & ~n24855;
  assign n24858 = ~n24854 & n24857;
  assign n24859 = ~n24853 & n24856;
  assign n24860 = ~n24852 & n42072;
  assign n24861 = pi32  & ~n24860;
  assign n24862 = pi32  & ~n24861;
  assign n24863 = pi32  & n24860;
  assign n24864 = ~n24860 & ~n24861;
  assign n24865 = ~pi32  & ~n24860;
  assign n24866 = ~n42073 & ~n42074;
  assign n24867 = ~n24147 & n41980;
  assign n24868 = ~n24147 & ~n24412;
  assign n24869 = ~n24148 & ~n24867;
  assign n24870 = ~n24866 & ~n42075;
  assign n24871 = n24866 & n42075;
  assign n24872 = ~n42075 & ~n24870;
  assign n24873 = n24866 & ~n42075;
  assign n24874 = ~n24866 & ~n24870;
  assign n24875 = ~n24866 & n42075;
  assign n24876 = ~n42076 & ~n42077;
  assign n24877 = ~n24870 & ~n24871;
  assign n24878 = n24851 & ~n42078;
  assign n24879 = ~n24851 & n42078;
  assign n24880 = ~n24878 & ~n24879;
  assign n24881 = ~n24127 & ~n24418;
  assign n24882 = n607 & n10844;
  assign n24883 = pi110  & n37489;
  assign n24884 = pi112  & n620;
  assign n24885 = pi111  & n622;
  assign n24886 = ~n24884 & ~n24885;
  assign n24887 = ~n24883 & ~n24885;
  assign n24888 = ~n24884 & n24887;
  assign n24889 = ~n24883 & n24886;
  assign n24890 = ~n24882 & n42079;
  assign n24891 = pi29  & ~n24890;
  assign n24892 = pi29  & ~n24891;
  assign n24893 = pi29  & n24890;
  assign n24894 = ~n24890 & ~n24891;
  assign n24895 = ~pi29  & ~n24890;
  assign n24896 = ~n42080 & ~n42081;
  assign n24897 = ~n24881 & ~n24896;
  assign n24898 = n24881 & n24896;
  assign n24899 = ~n24881 & n24896;
  assign n24900 = n24881 & ~n24896;
  assign n24901 = ~n24899 & ~n24900;
  assign n24902 = ~n24897 & ~n24898;
  assign n24903 = ~n24879 & ~n42082;
  assign n24904 = ~n24878 & n24903;
  assign n24905 = n24880 & ~n42082;
  assign n24906 = ~n24880 & n42082;
  assign n24907 = ~n42082 & ~n42083;
  assign n24908 = ~n24879 & ~n42083;
  assign n24909 = ~n24878 & n24908;
  assign n24910 = n24880 & ~n42083;
  assign n24911 = ~n24907 & ~n42084;
  assign n24912 = ~n42083 & ~n24906;
  assign n24913 = n24557 & ~n42085;
  assign n24914 = ~n24557 & n42085;
  assign n24915 = ~n24913 & ~n24914;
  assign n24916 = ~n24447 & ~n24455;
  assign n24917 = n5576 & n13057;
  assign n24918 = pi116  & n38406;
  assign n24919 = pi118  & n5591;
  assign n24920 = pi117  & n5593;
  assign n24921 = ~n24919 & ~n24920;
  assign n24922 = ~n24918 & ~n24920;
  assign n24923 = ~n24919 & n24922;
  assign n24924 = ~n24918 & n24921;
  assign n24925 = ~n24917 & n42086;
  assign n24926 = pi23  & ~n24925;
  assign n24927 = pi23  & ~n24926;
  assign n24928 = pi23  & n24925;
  assign n24929 = ~n24925 & ~n24926;
  assign n24930 = ~pi23  & ~n24925;
  assign n24931 = ~n42087 & ~n42088;
  assign n24932 = ~n24916 & ~n24931;
  assign n24933 = n24916 & n24931;
  assign n24934 = ~n24916 & ~n24932;
  assign n24935 = ~n24916 & n24931;
  assign n24936 = ~n24931 & ~n24932;
  assign n24937 = n24916 & ~n24931;
  assign n24938 = ~n42089 & ~n42090;
  assign n24939 = ~n24932 & ~n24933;
  assign n24940 = ~n24914 & ~n42091;
  assign n24941 = ~n24913 & n24940;
  assign n24942 = n24915 & ~n42091;
  assign n24943 = ~n24915 & n42091;
  assign n24944 = ~n42091 & ~n42092;
  assign n24945 = ~n24915 & ~n42091;
  assign n24946 = n24915 & ~n42092;
  assign n24947 = ~n24914 & ~n42092;
  assign n24948 = ~n24913 & n24947;
  assign n24949 = n24915 & n42091;
  assign n24950 = ~n42093 & ~n42094;
  assign n24951 = ~n42092 & ~n24943;
  assign n24952 = n24538 & ~n42095;
  assign n24953 = ~n24538 & n42095;
  assign n24954 = ~n24952 & ~n24953;
  assign n24955 = ~n24063 & ~n24469;
  assign n24956 = n8175 & n15111;
  assign n24957 = pi122  & n38895;
  assign n24958 = pi124  & n8190;
  assign n24959 = pi123  & n8192;
  assign n24960 = ~n24958 & ~n24959;
  assign n24961 = ~n24957 & ~n24959;
  assign n24962 = ~n24958 & n24961;
  assign n24963 = ~n24957 & n24960;
  assign n24964 = ~n24956 & n42096;
  assign n24965 = pi17  & ~n24964;
  assign n24966 = pi17  & ~n24965;
  assign n24967 = pi17  & n24964;
  assign n24968 = ~n24964 & ~n24965;
  assign n24969 = ~pi17  & ~n24964;
  assign n24970 = ~n42097 & ~n42098;
  assign n24971 = ~n24955 & ~n24970;
  assign n24972 = n24955 & n24970;
  assign n24973 = ~n24955 & n24970;
  assign n24974 = n24955 & ~n24970;
  assign n24975 = ~n24973 & ~n24974;
  assign n24976 = ~n24971 & ~n24972;
  assign n24977 = ~n24953 & ~n42099;
  assign n24978 = ~n24952 & n24977;
  assign n24979 = n24954 & ~n42099;
  assign n24980 = ~n24954 & n42099;
  assign n24981 = ~n42099 & ~n42100;
  assign n24982 = ~n24953 & ~n42100;
  assign n24983 = ~n24952 & n24982;
  assign n24984 = n24954 & ~n42100;
  assign n24985 = ~n24981 & ~n42101;
  assign n24986 = ~n42100 & ~n24980;
  assign n24987 = ~n24043 & ~n41994;
  assign n24988 = n563 & n40885;
  assign n24989 = pi125  & n37482;
  assign n24990 = pi127  & n578;
  assign n24991 = pi126  & n580;
  assign n24992 = ~n24990 & ~n24991;
  assign n24993 = ~n24989 & ~n24991;
  assign n24994 = ~n24990 & n24993;
  assign n24995 = ~n24989 & n24992;
  assign n24996 = ~n24988 & n42103;
  assign n24997 = pi14  & ~n24996;
  assign n24998 = pi14  & ~n24997;
  assign n24999 = pi14  & n24996;
  assign n25000 = ~n24996 & ~n24997;
  assign n25001 = ~pi14  & ~n24996;
  assign n25002 = ~n42104 & ~n42105;
  assign n25003 = ~n24987 & ~n25002;
  assign n25004 = n24987 & n25002;
  assign n25005 = ~n24987 & ~n25003;
  assign n25006 = ~n24987 & n25002;
  assign n25007 = ~n25002 & ~n25003;
  assign n25008 = n24987 & ~n25002;
  assign n25009 = ~n42106 & ~n42107;
  assign n25010 = ~n25003 & ~n25004;
  assign n25011 = ~n42102 & ~n42108;
  assign n25012 = n42102 & n42108;
  assign n25013 = n42102 & ~n42108;
  assign n25014 = ~n42102 & n42108;
  assign n25015 = ~n25013 & ~n25014;
  assign n25016 = ~n25011 & ~n25012;
  assign n25017 = ~n24519 & ~n42109;
  assign n25018 = n24519 & n42109;
  assign n25019 = ~n24519 & ~n25017;
  assign n25020 = ~n42109 & ~n25017;
  assign n25021 = ~n25019 & ~n25020;
  assign n25022 = ~n25017 & ~n25018;
  assign n25023 = ~n24518 & ~n42110;
  assign n25024 = n24518 & ~n25020;
  assign n25025 = ~n25019 & n25024;
  assign n25026 = n24518 & n42110;
  assign po75  = ~n25023 & ~n42111;
  assign n25028 = ~n25017 & ~n25023;
  assign n25029 = ~n25003 & ~n25011;
  assign n25030 = n5576 & n13027;
  assign n25031 = pi117  & n38406;
  assign n25032 = pi119  & n5591;
  assign n25033 = pi118  & n5593;
  assign n25034 = ~n25032 & ~n25033;
  assign n25035 = ~n25031 & ~n25033;
  assign n25036 = ~n25032 & n25035;
  assign n25037 = ~n25031 & n25034;
  assign n25038 = ~n25030 & n42112;
  assign n25039 = pi23  & ~n25038;
  assign n25040 = pi23  & ~n25039;
  assign n25041 = pi23  & n25038;
  assign n25042 = ~n25038 & ~n25039;
  assign n25043 = ~pi23  & ~n25038;
  assign n25044 = ~n42113 & ~n42114;
  assign n25045 = ~n24556 & ~n24913;
  assign n25046 = ~n25044 & ~n25045;
  assign n25047 = n25044 & n25045;
  assign n25048 = ~n25044 & ~n25046;
  assign n25049 = ~n25044 & n25045;
  assign n25050 = ~n25045 & ~n25046;
  assign n25051 = n25044 & ~n25045;
  assign n25052 = ~n42115 & ~n42116;
  assign n25053 = ~n25046 & ~n25047;
  assign n25054 = ~n24897 & ~n42083;
  assign n25055 = n4492 & n12530;
  assign n25056 = pi114  & n38208;
  assign n25057 = pi116  & n4507;
  assign n25058 = pi115  & n4509;
  assign n25059 = ~n25057 & ~n25058;
  assign n25060 = ~n25056 & ~n25058;
  assign n25061 = ~n25057 & n25060;
  assign n25062 = ~n25056 & n25059;
  assign n25063 = ~n4492 & n42118;
  assign n25064 = ~n12530 & n42118;
  assign n25065 = ~n25063 & ~n25064;
  assign n25066 = ~n25055 & n42118;
  assign n25067 = pi26  & ~n42119;
  assign n25068 = ~pi26  & n42119;
  assign n25069 = ~n25067 & ~n25068;
  assign n25070 = ~n25054 & ~n25069;
  assign n25071 = n25054 & n25069;
  assign n25072 = ~n25070 & ~n25071;
  assign n25073 = ~n24843 & ~n24850;
  assign n25074 = n649 & n9678;
  assign n25075 = pi108  & n37496;
  assign n25076 = pi110  & n662;
  assign n25077 = pi109  & n664;
  assign n25078 = ~n25076 & ~n25077;
  assign n25079 = ~n25075 & ~n25077;
  assign n25080 = ~n25076 & n25079;
  assign n25081 = ~n25075 & n25078;
  assign n25082 = ~n649 & n42120;
  assign n25083 = ~n9678 & n42120;
  assign n25084 = ~n25082 & ~n25083;
  assign n25085 = ~n25074 & n42120;
  assign n25086 = pi32  & ~n42121;
  assign n25087 = ~pi32  & n42121;
  assign n25088 = ~n25086 & ~n25087;
  assign n25089 = ~n25073 & ~n25088;
  assign n25090 = n25073 & n25088;
  assign n25091 = ~n25073 & ~n25089;
  assign n25092 = ~n25073 & n25088;
  assign n25093 = ~n25088 & ~n25089;
  assign n25094 = n25073 & ~n25088;
  assign n25095 = ~n42122 & ~n42123;
  assign n25096 = ~n25089 & ~n25090;
  assign n25097 = ~n24829 & ~n24837;
  assign n25098 = n691 & n8136;
  assign n25099 = pi102  & n37503;
  assign n25100 = pi104  & n704;
  assign n25101 = pi103  & n706;
  assign n25102 = ~n25100 & ~n25101;
  assign n25103 = ~n25099 & ~n25101;
  assign n25104 = ~n25100 & n25103;
  assign n25105 = ~n25099 & n25102;
  assign n25106 = ~n25098 & n42125;
  assign n25107 = pi38  & ~n25106;
  assign n25108 = pi38  & ~n25107;
  assign n25109 = pi38  & n25106;
  assign n25110 = ~n25106 & ~n25107;
  assign n25111 = ~pi38  & ~n25106;
  assign n25112 = ~n42126 & ~n42127;
  assign n25113 = ~n24805 & ~n24812;
  assign n25114 = n733 & n6839;
  assign n25115 = pi99  & n37510;
  assign n25116 = pi101  & n746;
  assign n25117 = pi100  & n748;
  assign n25118 = ~n25116 & ~n25117;
  assign n25119 = ~n25115 & ~n25117;
  assign n25120 = ~n25116 & n25119;
  assign n25121 = ~n25115 & n25118;
  assign n25122 = ~n25114 & n42128;
  assign n25123 = pi41  & ~n25122;
  assign n25124 = pi41  & ~n25123;
  assign n25125 = pi41  & n25122;
  assign n25126 = ~n25122 & ~n25123;
  assign n25127 = ~pi41  & ~n25122;
  assign n25128 = ~n42129 & ~n42130;
  assign n25129 = ~n24793 & ~n24799;
  assign n25130 = n940 & n5610;
  assign n25131 = pi96  & n37541;
  assign n25132 = pi98  & n953;
  assign n25133 = pi97  & n955;
  assign n25134 = ~n25132 & ~n25133;
  assign n25135 = ~n25131 & ~n25133;
  assign n25136 = ~n25132 & n25135;
  assign n25137 = ~n25131 & n25134;
  assign n25138 = ~n25130 & n42131;
  assign n25139 = pi44  & ~n25138;
  assign n25140 = pi44  & ~n25139;
  assign n25141 = pi44  & n25138;
  assign n25142 = ~n25138 & ~n25139;
  assign n25143 = ~pi44  & ~n25138;
  assign n25144 = ~n42132 & ~n42133;
  assign n25145 = n785 & n4494;
  assign n25146 = pi93  & n37520;
  assign n25147 = pi95  & n787;
  assign n25148 = pi94  & n795;
  assign n25149 = ~n25147 & ~n25148;
  assign n25150 = ~n25146 & ~n25148;
  assign n25151 = ~n25147 & n25150;
  assign n25152 = ~n25146 & n25149;
  assign n25153 = ~n25145 & n42134;
  assign n25154 = pi47  & ~n25153;
  assign n25155 = pi47  & ~n25154;
  assign n25156 = pi47  & n25153;
  assign n25157 = ~n25153 & ~n25154;
  assign n25158 = ~pi47  & ~n25153;
  assign n25159 = ~n42135 & ~n42136;
  assign n25160 = ~n24751 & ~n24758;
  assign n25161 = ~n24735 & ~n24743;
  assign n25162 = ~n24724 & ~n24732;
  assign n25163 = ~n24697 & ~n24707;
  assign n25164 = ~n24681 & ~n24689;
  assign n25165 = n2063 & n12674;
  assign n25166 = pi78  & n40107;
  assign n25167 = pi80  & n12676;
  assign n25168 = pi79  & n12684;
  assign n25169 = ~n25167 & ~n25168;
  assign n25170 = ~n25166 & ~n25168;
  assign n25171 = ~n25167 & n25170;
  assign n25172 = ~n25166 & n25169;
  assign n25173 = ~n25165 & n42137;
  assign n25174 = pi62  & ~n25173;
  assign n25175 = pi62  & ~n25174;
  assign n25176 = pi62  & n25173;
  assign n25177 = ~n25173 & ~n25174;
  assign n25178 = ~pi62  & ~n25173;
  assign n25179 = ~n42138 & ~n42139;
  assign n25180 = ~n24669 & ~n24678;
  assign n25181 = pi77  & ~n40814;
  assign n25182 = pi76  & n18285;
  assign n25183 = ~n25181 & ~n25182;
  assign n25184 = ~n25180 & n25183;
  assign n25185 = n25180 & ~n25183;
  assign n25186 = n25183 & ~n25184;
  assign n25187 = n25180 & n25183;
  assign n25188 = ~n25180 & ~n25184;
  assign n25189 = ~n25180 & ~n25183;
  assign n25190 = ~n42140 & ~n42141;
  assign n25191 = ~n25184 & ~n25185;
  assign n25192 = ~n25179 & ~n42142;
  assign n25193 = n25179 & n42142;
  assign n25194 = n25179 & ~n42142;
  assign n25195 = ~n25179 & n42142;
  assign n25196 = ~n25194 & ~n25195;
  assign n25197 = ~n25192 & ~n25193;
  assign n25198 = n25164 & n42143;
  assign n25199 = ~n25164 & ~n42143;
  assign n25200 = ~n25198 & ~n25199;
  assign n25201 = n2091 & n7882;
  assign n25202 = pi81  & n39128;
  assign n25203 = pi83  & n7884;
  assign n25204 = pi82  & n7892;
  assign n25205 = ~n25203 & ~n25204;
  assign n25206 = ~n25202 & ~n25204;
  assign n25207 = ~n25203 & n25206;
  assign n25208 = ~n25202 & n25205;
  assign n25209 = ~n25201 & n42144;
  assign n25210 = pi59  & ~n25209;
  assign n25211 = pi59  & ~n25210;
  assign n25212 = pi59  & n25209;
  assign n25213 = ~n25209 & ~n25210;
  assign n25214 = ~pi59  & ~n25209;
  assign n25215 = ~n42145 & ~n42146;
  assign n25216 = n25200 & ~n25215;
  assign n25217 = ~n25200 & n25215;
  assign n25218 = n25200 & ~n25216;
  assign n25219 = ~n25215 & ~n25216;
  assign n25220 = ~n25218 & ~n25219;
  assign n25221 = ~n25216 & ~n25217;
  assign n25222 = n25163 & n42147;
  assign n25223 = ~n25163 & ~n42147;
  assign n25224 = ~n25222 & ~n25223;
  assign n25225 = n2779 & n4312;
  assign n25226 = pi84  & n38376;
  assign n25227 = pi86  & n4314;
  assign n25228 = pi85  & n4322;
  assign n25229 = ~n25227 & ~n25228;
  assign n25230 = ~n25226 & ~n25228;
  assign n25231 = ~n25227 & n25230;
  assign n25232 = ~n25226 & n25229;
  assign n25233 = ~n25225 & n42148;
  assign n25234 = pi56  & ~n25233;
  assign n25235 = pi56  & ~n25234;
  assign n25236 = pi56  & n25233;
  assign n25237 = ~n25233 & ~n25234;
  assign n25238 = ~pi56  & ~n25233;
  assign n25239 = ~n42149 & ~n42150;
  assign n25240 = ~n25224 & n25239;
  assign n25241 = n25224 & ~n25239;
  assign n25242 = n25224 & ~n25241;
  assign n25243 = ~n25239 & ~n25241;
  assign n25244 = ~n25242 & ~n25243;
  assign n25245 = ~n25240 & ~n25241;
  assign n25246 = n25162 & n42151;
  assign n25247 = ~n25162 & ~n42151;
  assign n25248 = ~n25246 & ~n25247;
  assign n25249 = n1971 & n3591;
  assign n25250 = pi87  & n37864;
  assign n25251 = pi89  & n1973;
  assign n25252 = pi88  & n1981;
  assign n25253 = ~n25251 & ~n25252;
  assign n25254 = ~n25250 & ~n25252;
  assign n25255 = ~n25251 & n25254;
  assign n25256 = ~n25250 & n25253;
  assign n25257 = ~n25249 & n42152;
  assign n25258 = pi53  & ~n25257;
  assign n25259 = pi53  & ~n25258;
  assign n25260 = pi53  & n25257;
  assign n25261 = ~n25257 & ~n25258;
  assign n25262 = ~pi53  & ~n25257;
  assign n25263 = ~n42153 & ~n42154;
  assign n25264 = n25248 & ~n25263;
  assign n25265 = ~n25248 & n25263;
  assign n25266 = n25248 & ~n25264;
  assign n25267 = ~n25263 & ~n25264;
  assign n25268 = ~n25266 & ~n25267;
  assign n25269 = ~n25264 & ~n25265;
  assign n25270 = n25161 & n42155;
  assign n25271 = ~n25161 & ~n42155;
  assign n25272 = ~n25270 & ~n25271;
  assign n25273 = n894 & n4453;
  assign n25274 = pi90  & n37580;
  assign n25275 = pi92  & n896;
  assign n25276 = pi91  & n904;
  assign n25277 = ~n25275 & ~n25276;
  assign n25278 = ~n25274 & ~n25276;
  assign n25279 = ~n25275 & n25278;
  assign n25280 = ~n25274 & n25277;
  assign n25281 = ~n25273 & n42156;
  assign n25282 = pi50  & ~n25281;
  assign n25283 = pi50  & ~n25282;
  assign n25284 = pi50  & n25281;
  assign n25285 = ~n25281 & ~n25282;
  assign n25286 = ~pi50  & ~n25281;
  assign n25287 = ~n42157 & ~n42158;
  assign n25288 = ~n25272 & n25287;
  assign n25289 = n25272 & ~n25287;
  assign n25290 = ~n25288 & ~n25289;
  assign n25291 = ~n25160 & n25290;
  assign n25292 = n25160 & ~n25290;
  assign n25293 = ~n25160 & ~n25291;
  assign n25294 = n25290 & ~n25291;
  assign n25295 = ~n25293 & ~n25294;
  assign n25296 = ~n25291 & ~n25292;
  assign n25297 = ~n25159 & ~n42159;
  assign n25298 = n25159 & ~n25294;
  assign n25299 = ~n25293 & n25298;
  assign n25300 = n25159 & n42159;
  assign n25301 = ~n25297 & ~n42160;
  assign n25302 = ~n42058 & n25301;
  assign n25303 = n42058 & ~n25301;
  assign n25304 = ~n25302 & ~n25303;
  assign n25305 = ~n25144 & n25304;
  assign n25306 = n25144 & ~n25304;
  assign n25307 = ~n25305 & ~n25306;
  assign n25308 = ~n25129 & n25307;
  assign n25309 = n25129 & ~n25307;
  assign n25310 = ~n25129 & ~n25308;
  assign n25311 = n25307 & ~n25308;
  assign n25312 = ~n25310 & ~n25311;
  assign n25313 = ~n25308 & ~n25309;
  assign n25314 = ~n25128 & ~n42161;
  assign n25315 = n25128 & ~n25311;
  assign n25316 = ~n25310 & n25315;
  assign n25317 = n25128 & n42161;
  assign n25318 = ~n25314 & ~n42162;
  assign n25319 = ~n25113 & n25318;
  assign n25320 = n25113 & ~n25318;
  assign n25321 = ~n25113 & ~n25319;
  assign n25322 = n25318 & ~n25319;
  assign n25323 = ~n25321 & ~n25322;
  assign n25324 = ~n25319 & ~n25320;
  assign n25325 = ~n25112 & ~n42163;
  assign n25326 = n25112 & ~n25322;
  assign n25327 = ~n25321 & n25326;
  assign n25328 = n25112 & n42163;
  assign n25329 = ~n25325 & ~n42164;
  assign n25330 = ~n25097 & n25329;
  assign n25331 = n25097 & ~n25329;
  assign n25332 = ~n25330 & ~n25331;
  assign n25333 = n2104 & n8177;
  assign n25334 = pi105  & n37758;
  assign n25335 = pi107  & n2117;
  assign n25336 = pi106  & n2119;
  assign n25337 = ~n25335 & ~n25336;
  assign n25338 = ~n25334 & ~n25336;
  assign n25339 = ~n25335 & n25338;
  assign n25340 = ~n25334 & n25337;
  assign n25341 = ~n25333 & n42165;
  assign n25342 = pi35  & ~n25341;
  assign n25343 = pi35  & ~n25342;
  assign n25344 = pi35  & n25341;
  assign n25345 = ~n25341 & ~n25342;
  assign n25346 = ~pi35  & ~n25341;
  assign n25347 = ~n42166 & ~n42167;
  assign n25348 = n25332 & ~n25347;
  assign n25349 = ~n25332 & n25347;
  assign n25350 = n25332 & ~n25348;
  assign n25351 = ~n25347 & ~n25348;
  assign n25352 = ~n25350 & ~n25351;
  assign n25353 = ~n25348 & ~n25349;
  assign n25354 = ~n42124 & ~n42168;
  assign n25355 = n42124 & n42168;
  assign n25356 = ~n42168 & ~n25354;
  assign n25357 = ~n42124 & ~n25354;
  assign n25358 = ~n25356 & ~n25357;
  assign n25359 = ~n25354 & ~n25355;
  assign n25360 = n607 & n11276;
  assign n25361 = pi111  & n37489;
  assign n25362 = pi113  & n620;
  assign n25363 = pi112  & n622;
  assign n25364 = ~n25362 & ~n25363;
  assign n25365 = ~n25361 & ~n25363;
  assign n25366 = ~n25362 & n25365;
  assign n25367 = ~n25361 & n25364;
  assign n25368 = ~n25360 & n42170;
  assign n25369 = pi29  & ~n25368;
  assign n25370 = pi29  & ~n25369;
  assign n25371 = pi29  & n25368;
  assign n25372 = ~n25368 & ~n25369;
  assign n25373 = ~pi29  & ~n25368;
  assign n25374 = ~n42171 & ~n42172;
  assign n25375 = ~n24870 & ~n24878;
  assign n25376 = ~n25374 & ~n25375;
  assign n25377 = n25374 & n25375;
  assign n25378 = ~n25374 & ~n25376;
  assign n25379 = ~n25374 & n25375;
  assign n25380 = ~n25375 & ~n25376;
  assign n25381 = n25374 & ~n25375;
  assign n25382 = ~n42173 & ~n42174;
  assign n25383 = ~n25376 & ~n25377;
  assign n25384 = ~n42169 & ~n42175;
  assign n25385 = n42169 & n42175;
  assign n25386 = ~n42175 & ~n25384;
  assign n25387 = ~n42169 & ~n25384;
  assign n25388 = ~n25386 & ~n25387;
  assign n25389 = ~n25384 & ~n25385;
  assign n25390 = n25072 & ~n42176;
  assign n25391 = ~n42176 & ~n25390;
  assign n25392 = ~n25072 & ~n42176;
  assign n25393 = n25072 & ~n25390;
  assign n25394 = n25072 & n42176;
  assign n25395 = ~n25072 & n42176;
  assign n25396 = ~n25390 & ~n25395;
  assign n25397 = ~n42177 & ~n42178;
  assign n25398 = ~n42117 & n42179;
  assign n25399 = n42117 & ~n42179;
  assign n25400 = ~n42117 & ~n25398;
  assign n25401 = n42179 & ~n25398;
  assign n25402 = ~n25400 & ~n25401;
  assign n25403 = ~n25398 & ~n25399;
  assign n25404 = ~n24932 & ~n42092;
  assign n25405 = n6785 & n15049;
  assign n25406 = pi120  & n38631;
  assign n25407 = pi122  & n6800;
  assign n25408 = pi121  & n6802;
  assign n25409 = ~n25407 & ~n25408;
  assign n25410 = ~n25406 & ~n25408;
  assign n25411 = ~n25407 & n25410;
  assign n25412 = ~n25406 & n25409;
  assign n25413 = ~n6785 & n42181;
  assign n25414 = ~n15049 & n42181;
  assign n25415 = ~n25413 & ~n25414;
  assign n25416 = ~n25405 & n42181;
  assign n25417 = pi20  & ~n42182;
  assign n25418 = ~pi20  & n42182;
  assign n25419 = ~n25417 & ~n25418;
  assign n25420 = ~n25404 & ~n25419;
  assign n25421 = n25404 & n25419;
  assign n25422 = ~n25404 & ~n25420;
  assign n25423 = ~n25404 & n25419;
  assign n25424 = ~n25419 & ~n25420;
  assign n25425 = n25404 & ~n25419;
  assign n25426 = ~n42183 & ~n42184;
  assign n25427 = ~n25420 & ~n25421;
  assign n25428 = ~n42180 & ~n42185;
  assign n25429 = n42180 & n42185;
  assign n25430 = ~n42180 & ~n25428;
  assign n25431 = ~n42185 & ~n25428;
  assign n25432 = ~n25430 & ~n25431;
  assign n25433 = ~n25428 & ~n25429;
  assign n25434 = n8175 & n15068;
  assign n25435 = pi123  & n38895;
  assign n25436 = pi125  & n8190;
  assign n25437 = pi124  & n8192;
  assign n25438 = ~n25436 & ~n25437;
  assign n25439 = ~n25435 & ~n25437;
  assign n25440 = ~n25436 & n25439;
  assign n25441 = ~n25435 & n25438;
  assign n25442 = ~n25434 & n42187;
  assign n25443 = pi17  & ~n25442;
  assign n25444 = pi17  & ~n25443;
  assign n25445 = pi17  & n25442;
  assign n25446 = ~n25442 & ~n25443;
  assign n25447 = ~pi17  & ~n25442;
  assign n25448 = ~n42188 & ~n42189;
  assign n25449 = ~n24537 & ~n24952;
  assign n25450 = ~n25448 & ~n25449;
  assign n25451 = n25448 & n25449;
  assign n25452 = ~n25448 & ~n25450;
  assign n25453 = ~n25448 & n25449;
  assign n25454 = ~n25449 & ~n25450;
  assign n25455 = n25448 & ~n25449;
  assign n25456 = ~n42190 & ~n42191;
  assign n25457 = ~n25450 & ~n25451;
  assign n25458 = ~n42186 & ~n42192;
  assign n25459 = n42186 & n42192;
  assign n25460 = ~n42192 & ~n25458;
  assign n25461 = ~n42186 & ~n25458;
  assign n25462 = ~n25460 & ~n25461;
  assign n25463 = ~n25458 & ~n25459;
  assign n25464 = ~n24971 & ~n42100;
  assign n25465 = n563 & n40891;
  assign n25466 = pi126  & n37482;
  assign n25467 = pi127  & n580;
  assign n25468 = ~n25466 & ~n25467;
  assign n25469 = ~n563 & n25468;
  assign n25470 = ~n40891 & n25468;
  assign n25471 = ~n25469 & ~n25470;
  assign n25472 = ~n25465 & n25468;
  assign n25473 = pi14  & ~n42194;
  assign n25474 = ~pi14  & n42194;
  assign n25475 = ~n25473 & ~n25474;
  assign n25476 = ~n25464 & ~n25475;
  assign n25477 = n25464 & n25475;
  assign n25478 = ~n25464 & ~n25476;
  assign n25479 = ~n25464 & n25475;
  assign n25480 = ~n25475 & ~n25476;
  assign n25481 = n25464 & ~n25475;
  assign n25482 = ~n42195 & ~n42196;
  assign n25483 = ~n25476 & ~n25477;
  assign n25484 = ~n42193 & ~n42197;
  assign n25485 = n42193 & ~n42196;
  assign n25486 = ~n42195 & n25485;
  assign n25487 = n42193 & ~n42195;
  assign n25488 = ~n42196 & n25487;
  assign n25489 = n42193 & n42197;
  assign n25490 = ~n25484 & ~n42198;
  assign n25491 = ~n25029 & n25490;
  assign n25492 = n25029 & ~n25490;
  assign n25493 = ~n25029 & ~n25491;
  assign n25494 = n25490 & ~n25491;
  assign n25495 = ~n25493 & ~n25494;
  assign n25496 = ~n25491 & ~n25492;
  assign n25497 = ~n25028 & ~n42199;
  assign n25498 = n25028 & ~n25494;
  assign n25499 = ~n25493 & n25498;
  assign n25500 = n25028 & n42199;
  assign po76  = ~n25497 & ~n42200;
  assign n25502 = ~n25491 & ~n25497;
  assign n25503 = ~n25476 & ~n25484;
  assign n25504 = n6785 & n14961;
  assign n25505 = pi121  & n38631;
  assign n25506 = pi123  & n6800;
  assign n25507 = pi122  & n6802;
  assign n25508 = ~n25506 & ~n25507;
  assign n25509 = ~n25505 & ~n25507;
  assign n25510 = ~n25506 & n25509;
  assign n25511 = ~n25505 & n25508;
  assign n25512 = ~n25504 & n42201;
  assign n25513 = pi20  & ~n25512;
  assign n25514 = pi20  & ~n25513;
  assign n25515 = pi20  & n25512;
  assign n25516 = ~n25512 & ~n25513;
  assign n25517 = ~pi20  & ~n25512;
  assign n25518 = ~n42202 & ~n42203;
  assign n25519 = ~n25046 & ~n25398;
  assign n25520 = n25518 & n25519;
  assign n25521 = ~n25518 & ~n25519;
  assign n25522 = ~n25520 & ~n25521;
  assign n25523 = n5576 & n14913;
  assign n25524 = pi118  & n38406;
  assign n25525 = pi120  & n5591;
  assign n25526 = pi119  & n5593;
  assign n25527 = ~n25525 & ~n25526;
  assign n25528 = ~n25524 & ~n25526;
  assign n25529 = ~n25525 & n25528;
  assign n25530 = ~n25524 & n25527;
  assign n25531 = ~n25523 & n42204;
  assign n25532 = pi23  & ~n25531;
  assign n25533 = pi23  & ~n25532;
  assign n25534 = pi23  & n25531;
  assign n25535 = ~n25531 & ~n25532;
  assign n25536 = ~pi23  & ~n25531;
  assign n25537 = ~n42205 & ~n42206;
  assign n25538 = ~n25070 & n42176;
  assign n25539 = ~n25070 & ~n25390;
  assign n25540 = ~n25071 & ~n25538;
  assign n25541 = n25537 & n42207;
  assign n25542 = ~n25537 & ~n42207;
  assign n25543 = ~n25541 & ~n25542;
  assign n25544 = n4492 & n13079;
  assign n25545 = pi115  & n38208;
  assign n25546 = pi117  & n4507;
  assign n25547 = pi116  & n4509;
  assign n25548 = ~n25546 & ~n25547;
  assign n25549 = ~n25545 & ~n25547;
  assign n25550 = ~n25546 & n25549;
  assign n25551 = ~n25545 & n25548;
  assign n25552 = ~n25544 & n42208;
  assign n25553 = pi26  & ~n25552;
  assign n25554 = pi26  & ~n25553;
  assign n25555 = pi26  & n25552;
  assign n25556 = ~n25552 & ~n25553;
  assign n25557 = ~pi26  & ~n25552;
  assign n25558 = ~n42209 & ~n42210;
  assign n25559 = ~n25376 & ~n25384;
  assign n25560 = n25558 & n25559;
  assign n25561 = ~n25558 & ~n25559;
  assign n25562 = ~n25560 & ~n25561;
  assign n25563 = ~n25089 & ~n25354;
  assign n25564 = n607 & n11258;
  assign n25565 = pi112  & n37489;
  assign n25566 = pi114  & n620;
  assign n25567 = pi113  & n622;
  assign n25568 = ~n25566 & ~n25567;
  assign n25569 = ~n25565 & ~n25567;
  assign n25570 = ~n25566 & n25569;
  assign n25571 = ~n25565 & n25568;
  assign n25572 = ~n607 & n42211;
  assign n25573 = ~n11258 & n42211;
  assign n25574 = ~n25572 & ~n25573;
  assign n25575 = ~n25564 & n42211;
  assign n25576 = pi29  & ~n42212;
  assign n25577 = ~pi29  & n42212;
  assign n25578 = ~n25576 & ~n25577;
  assign n25579 = ~n25563 & ~n25578;
  assign n25580 = n25563 & n25578;
  assign n25581 = ~n25579 & ~n25580;
  assign n25582 = n565 & n649;
  assign n25583 = pi109  & n37496;
  assign n25584 = pi111  & n662;
  assign n25585 = pi110  & n664;
  assign n25586 = ~n25584 & ~n25585;
  assign n25587 = ~n25583 & ~n25585;
  assign n25588 = ~n25584 & n25587;
  assign n25589 = ~n25583 & n25586;
  assign n25590 = ~n649 & n42213;
  assign n25591 = ~n565 & n42213;
  assign n25592 = ~n25590 & ~n25591;
  assign n25593 = ~n25582 & n42213;
  assign n25594 = pi32  & ~n42214;
  assign n25595 = ~pi32  & n42214;
  assign n25596 = ~n25594 & ~n25595;
  assign n25597 = ~n25330 & n25347;
  assign n25598 = ~n25330 & ~n25348;
  assign n25599 = ~n25331 & ~n25597;
  assign n25600 = ~n25596 & ~n42215;
  assign n25601 = n25596 & n42215;
  assign n25602 = ~n25600 & ~n25601;
  assign n25603 = n2104 & n9277;
  assign n25604 = pi106  & n37758;
  assign n25605 = pi108  & n2117;
  assign n25606 = pi107  & n2119;
  assign n25607 = ~n25605 & ~n25606;
  assign n25608 = ~n25604 & ~n25606;
  assign n25609 = ~n25605 & n25608;
  assign n25610 = ~n25604 & n25607;
  assign n25611 = ~n25603 & n42216;
  assign n25612 = pi35  & ~n25611;
  assign n25613 = pi35  & ~n25612;
  assign n25614 = pi35  & n25611;
  assign n25615 = ~n25611 & ~n25612;
  assign n25616 = ~pi35  & ~n25611;
  assign n25617 = ~n42217 & ~n42218;
  assign n25618 = ~n25319 & ~n25325;
  assign n25619 = n691 & n8229;
  assign n25620 = pi103  & n37503;
  assign n25621 = pi105  & n704;
  assign n25622 = pi104  & n706;
  assign n25623 = ~n25621 & ~n25622;
  assign n25624 = ~n25620 & ~n25622;
  assign n25625 = ~n25621 & n25624;
  assign n25626 = ~n25620 & n25623;
  assign n25627 = ~n25619 & n42219;
  assign n25628 = pi38  & ~n25627;
  assign n25629 = pi38  & ~n25628;
  assign n25630 = pi38  & n25627;
  assign n25631 = ~n25627 & ~n25628;
  assign n25632 = ~pi38  & ~n25627;
  assign n25633 = ~n42220 & ~n42221;
  assign n25634 = ~n25308 & ~n25314;
  assign n25635 = ~n25302 & ~n25305;
  assign n25636 = ~n25291 & ~n25297;
  assign n25637 = n785 & n5281;
  assign n25638 = pi94  & n37520;
  assign n25639 = pi96  & n787;
  assign n25640 = pi95  & n795;
  assign n25641 = ~n25639 & ~n25640;
  assign n25642 = ~n25638 & ~n25640;
  assign n25643 = ~n25639 & n25642;
  assign n25644 = ~n25638 & n25641;
  assign n25645 = ~n25637 & n42222;
  assign n25646 = pi47  & ~n25645;
  assign n25647 = pi47  & ~n25646;
  assign n25648 = pi47  & n25645;
  assign n25649 = ~n25645 & ~n25646;
  assign n25650 = ~pi47  & ~n25645;
  assign n25651 = ~n42223 & ~n42224;
  assign n25652 = ~n25271 & ~n25289;
  assign n25653 = n1971 & n3566;
  assign n25654 = pi88  & n37864;
  assign n25655 = pi90  & n1973;
  assign n25656 = pi89  & n1981;
  assign n25657 = ~n25655 & ~n25656;
  assign n25658 = ~n25654 & ~n25656;
  assign n25659 = ~n25655 & n25658;
  assign n25660 = ~n25654 & n25657;
  assign n25661 = ~n25653 & n42225;
  assign n25662 = pi53  & ~n25661;
  assign n25663 = pi53  & ~n25662;
  assign n25664 = pi53  & n25661;
  assign n25665 = ~n25661 & ~n25662;
  assign n25666 = ~pi53  & ~n25661;
  assign n25667 = ~n42226 & ~n42227;
  assign n25668 = ~n25184 & ~n25192;
  assign n25669 = pi78  & ~n40814;
  assign n25670 = pi77  & n18285;
  assign n25671 = ~n25669 & ~n25670;
  assign n25672 = n25183 & ~n25671;
  assign n25673 = ~n25183 & n25671;
  assign n25674 = ~n25672 & ~n25673;
  assign n25675 = n2154 & n12674;
  assign n25676 = pi79  & n40107;
  assign n25677 = pi81  & n12676;
  assign n25678 = pi80  & n12684;
  assign n25679 = ~n25677 & ~n25678;
  assign n25680 = ~n25676 & ~n25678;
  assign n25681 = ~n25677 & n25680;
  assign n25682 = ~n25676 & n25679;
  assign n25683 = ~n12674 & n42228;
  assign n25684 = ~n2154 & n42228;
  assign n25685 = ~n25683 & ~n25684;
  assign n25686 = ~n25675 & n42228;
  assign n25687 = pi62  & ~n42229;
  assign n25688 = ~pi62  & n42229;
  assign n25689 = ~n25687 & ~n25688;
  assign n25690 = n25674 & ~n25689;
  assign n25691 = ~n25674 & n25689;
  assign n25692 = ~n25690 & ~n25691;
  assign n25693 = ~n25668 & n25692;
  assign n25694 = n25668 & ~n25692;
  assign n25695 = ~n25693 & ~n25694;
  assign n25696 = n2591 & n7882;
  assign n25697 = pi82  & n39128;
  assign n25698 = pi84  & n7884;
  assign n25699 = pi83  & n7892;
  assign n25700 = ~n25698 & ~n25699;
  assign n25701 = ~n25697 & ~n25699;
  assign n25702 = ~n25698 & n25701;
  assign n25703 = ~n25697 & n25700;
  assign n25704 = ~n25696 & n42230;
  assign n25705 = pi59  & ~n25704;
  assign n25706 = pi59  & ~n25705;
  assign n25707 = pi59  & n25704;
  assign n25708 = ~n25704 & ~n25705;
  assign n25709 = ~pi59  & ~n25704;
  assign n25710 = ~n42231 & ~n42232;
  assign n25711 = n25695 & ~n25710;
  assign n25712 = ~n25695 & n25710;
  assign n25713 = n25695 & ~n25711;
  assign n25714 = ~n25710 & ~n25711;
  assign n25715 = ~n25713 & ~n25714;
  assign n25716 = ~n25711 & ~n25712;
  assign n25717 = ~n25199 & n25215;
  assign n25718 = ~n25199 & ~n25216;
  assign n25719 = ~n25198 & ~n25717;
  assign n25720 = n42233 & n42234;
  assign n25721 = ~n42233 & ~n42234;
  assign n25722 = ~n25720 & ~n25721;
  assign n25723 = n636 & n4312;
  assign n25724 = pi85  & n38376;
  assign n25725 = pi87  & n4314;
  assign n25726 = pi86  & n4322;
  assign n25727 = ~n25725 & ~n25726;
  assign n25728 = ~n25724 & ~n25726;
  assign n25729 = ~n25725 & n25728;
  assign n25730 = ~n25724 & n25727;
  assign n25731 = ~n25723 & n42235;
  assign n25732 = pi56  & ~n25731;
  assign n25733 = pi56  & ~n25732;
  assign n25734 = pi56  & n25731;
  assign n25735 = ~n25731 & ~n25732;
  assign n25736 = ~pi56  & ~n25731;
  assign n25737 = ~n42236 & ~n42237;
  assign n25738 = ~n25722 & n25737;
  assign n25739 = n25722 & ~n25737;
  assign n25740 = ~n25738 & ~n25739;
  assign n25741 = ~n25223 & n25239;
  assign n25742 = ~n25223 & ~n25241;
  assign n25743 = ~n25222 & ~n25741;
  assign n25744 = n25740 & ~n42238;
  assign n25745 = ~n25740 & n42238;
  assign n25746 = ~n25744 & ~n25745;
  assign n25747 = ~n25667 & n25746;
  assign n25748 = n25667 & ~n25746;
  assign n25749 = ~n25747 & ~n25748;
  assign n25750 = ~n25247 & n25263;
  assign n25751 = ~n25247 & ~n25264;
  assign n25752 = ~n25246 & ~n25750;
  assign n25753 = n25749 & ~n42239;
  assign n25754 = ~n25749 & n42239;
  assign n25755 = ~n25753 & ~n25754;
  assign n25756 = n894 & n4544;
  assign n25757 = pi91  & n37580;
  assign n25758 = pi93  & n896;
  assign n25759 = pi92  & n904;
  assign n25760 = ~n25758 & ~n25759;
  assign n25761 = ~n25757 & ~n25759;
  assign n25762 = ~n25758 & n25761;
  assign n25763 = ~n25757 & n25760;
  assign n25764 = ~n25756 & n42240;
  assign n25765 = pi50  & ~n25764;
  assign n25766 = pi50  & ~n25765;
  assign n25767 = pi50  & n25764;
  assign n25768 = ~n25764 & ~n25765;
  assign n25769 = ~pi50  & ~n25764;
  assign n25770 = ~n42241 & ~n42242;
  assign n25771 = n25755 & ~n25770;
  assign n25772 = ~n25755 & n25770;
  assign n25773 = n25755 & ~n25771;
  assign n25774 = ~n25770 & ~n25771;
  assign n25775 = ~n25773 & ~n25774;
  assign n25776 = ~n25771 & ~n25772;
  assign n25777 = ~n25652 & ~n42243;
  assign n25778 = n25652 & n42243;
  assign n25779 = ~n42243 & ~n25777;
  assign n25780 = ~n25652 & ~n25777;
  assign n25781 = ~n25779 & ~n25780;
  assign n25782 = ~n25777 & ~n25778;
  assign n25783 = n25651 & ~n42244;
  assign n25784 = ~n25651 & n42244;
  assign n25785 = ~n25651 & ~n42244;
  assign n25786 = n25651 & n42244;
  assign n25787 = ~n25785 & ~n25786;
  assign n25788 = ~n25783 & ~n25784;
  assign n25789 = n25636 & ~n42245;
  assign n25790 = ~n25636 & n42245;
  assign n25791 = ~n25789 & ~n25790;
  assign n25792 = n940 & n5578;
  assign n25793 = pi97  & n37541;
  assign n25794 = pi99  & n953;
  assign n25795 = pi98  & n955;
  assign n25796 = ~n25794 & ~n25795;
  assign n25797 = ~n25793 & ~n25795;
  assign n25798 = ~n25794 & n25797;
  assign n25799 = ~n25793 & n25796;
  assign n25800 = ~n25792 & n42246;
  assign n25801 = pi44  & ~n25800;
  assign n25802 = pi44  & ~n25801;
  assign n25803 = pi44  & n25800;
  assign n25804 = ~n25800 & ~n25801;
  assign n25805 = ~pi44  & ~n25800;
  assign n25806 = ~n42247 & ~n42248;
  assign n25807 = n25791 & ~n25806;
  assign n25808 = ~n25791 & n25806;
  assign n25809 = n25791 & ~n25807;
  assign n25810 = ~n25806 & ~n25807;
  assign n25811 = ~n25809 & ~n25810;
  assign n25812 = ~n25807 & ~n25808;
  assign n25813 = n25635 & n42249;
  assign n25814 = ~n25635 & ~n42249;
  assign n25815 = ~n25813 & ~n25814;
  assign n25816 = n733 & n6819;
  assign n25817 = pi100  & n37510;
  assign n25818 = pi102  & n746;
  assign n25819 = pi101  & n748;
  assign n25820 = ~n25818 & ~n25819;
  assign n25821 = ~n25817 & ~n25819;
  assign n25822 = ~n25818 & n25821;
  assign n25823 = ~n25817 & n25820;
  assign n25824 = ~n25816 & n42250;
  assign n25825 = pi41  & ~n25824;
  assign n25826 = pi41  & ~n25825;
  assign n25827 = pi41  & n25824;
  assign n25828 = ~n25824 & ~n25825;
  assign n25829 = ~pi41  & ~n25824;
  assign n25830 = ~n42251 & ~n42252;
  assign n25831 = ~n25815 & n25830;
  assign n25832 = n25815 & ~n25830;
  assign n25833 = ~n25831 & ~n25832;
  assign n25834 = ~n25634 & n25833;
  assign n25835 = n25634 & ~n25833;
  assign n25836 = ~n25834 & ~n25835;
  assign n25837 = ~n25633 & n25836;
  assign n25838 = n25633 & ~n25836;
  assign n25839 = ~n25837 & ~n25838;
  assign n25840 = ~n25618 & n25839;
  assign n25841 = n25618 & ~n25839;
  assign n25842 = ~n25840 & ~n25841;
  assign n25843 = n25617 & ~n25842;
  assign n25844 = ~n25617 & n25842;
  assign n25845 = ~n25617 & ~n25844;
  assign n25846 = n25842 & ~n25844;
  assign n25847 = ~n25845 & ~n25846;
  assign n25848 = ~n25843 & ~n25844;
  assign n25849 = n25602 & ~n42253;
  assign n25850 = ~n25602 & n42253;
  assign n25851 = n25602 & ~n25849;
  assign n25852 = ~n42253 & ~n25849;
  assign n25853 = ~n25851 & ~n25852;
  assign n25854 = ~n25849 & ~n25850;
  assign n25855 = n25581 & ~n42254;
  assign n25856 = n25581 & ~n25855;
  assign n25857 = n25581 & n42254;
  assign n25858 = ~n42254 & ~n25855;
  assign n25859 = ~n25581 & ~n42254;
  assign n25860 = ~n25581 & n42254;
  assign n25861 = ~n25855 & ~n25860;
  assign n25862 = ~n42255 & ~n42256;
  assign n25863 = n25562 & n42257;
  assign n25864 = ~n25562 & ~n42257;
  assign n25865 = n25562 & ~n25863;
  assign n25866 = n25562 & ~n42257;
  assign n25867 = n42257 & ~n25863;
  assign n25868 = ~n25562 & n42257;
  assign n25869 = ~n42258 & ~n42259;
  assign n25870 = ~n25863 & ~n25864;
  assign n25871 = n25543 & ~n42260;
  assign n25872 = ~n25543 & n42260;
  assign n25873 = ~n25871 & ~n25872;
  assign n25874 = n25522 & ~n25872;
  assign n25875 = ~n25871 & n25874;
  assign n25876 = n25522 & n25873;
  assign n25877 = ~n25522 & ~n25873;
  assign n25878 = n25522 & ~n42261;
  assign n25879 = ~n25872 & ~n42261;
  assign n25880 = ~n25871 & n25879;
  assign n25881 = n25873 & ~n42261;
  assign n25882 = ~n25878 & ~n42262;
  assign n25883 = ~n42261 & ~n25877;
  assign n25884 = ~n25420 & ~n25428;
  assign n25885 = n8175 & n15021;
  assign n25886 = pi124  & n38895;
  assign n25887 = pi126  & n8190;
  assign n25888 = pi125  & n8192;
  assign n25889 = ~n25887 & ~n25888;
  assign n25890 = ~n25886 & ~n25888;
  assign n25891 = ~n25887 & n25890;
  assign n25892 = ~n25886 & n25889;
  assign n25893 = ~n8175 & n42264;
  assign n25894 = ~n15021 & n42264;
  assign n25895 = ~n25893 & ~n25894;
  assign n25896 = ~n25885 & n42264;
  assign n25897 = pi17  & ~n42265;
  assign n25898 = ~pi17  & n42265;
  assign n25899 = ~n25897 & ~n25898;
  assign n25900 = ~n25884 & ~n25899;
  assign n25901 = n25884 & n25899;
  assign n25902 = ~n25884 & ~n25900;
  assign n25903 = ~n25884 & n25899;
  assign n25904 = ~n25899 & ~n25900;
  assign n25905 = n25884 & ~n25899;
  assign n25906 = ~n42266 & ~n42267;
  assign n25907 = ~n25900 & ~n25901;
  assign n25908 = ~n42263 & ~n42268;
  assign n25909 = n42263 & ~n42267;
  assign n25910 = ~n42266 & n25909;
  assign n25911 = n42263 & ~n42266;
  assign n25912 = ~n42267 & n25911;
  assign n25913 = n42263 & n42268;
  assign n25914 = ~n25908 & ~n42269;
  assign n25915 = ~n25450 & ~n25458;
  assign n25916 = n563 & ~n18675;
  assign n25917 = ~n37482 & ~n25916;
  assign n25918 = pi127  & n37482;
  assign n25919 = n563 & n18680;
  assign n25920 = ~n25918 & ~n25919;
  assign n25921 = pi127  & ~n25917;
  assign n25922 = pi14  & ~n42270;
  assign n25923 = pi14  & ~n25922;
  assign n25924 = pi14  & n42270;
  assign n25925 = ~n42270 & ~n25922;
  assign n25926 = ~pi14  & ~n42270;
  assign n25927 = ~n42271 & ~n42272;
  assign n25928 = ~n25915 & ~n25927;
  assign n25929 = n25915 & n25927;
  assign n25930 = ~n25915 & ~n25928;
  assign n25931 = ~n25927 & ~n25928;
  assign n25932 = ~n25930 & ~n25931;
  assign n25933 = ~n25928 & ~n25929;
  assign n25934 = n25914 & ~n42273;
  assign n25935 = ~n25914 & n42273;
  assign n25936 = ~n25934 & ~n25935;
  assign n25937 = ~n25503 & n25936;
  assign n25938 = n25503 & ~n25936;
  assign n25939 = ~n25937 & ~n25938;
  assign n25940 = ~n25502 & n25939;
  assign n25941 = n25502 & ~n25939;
  assign po77  = ~n25940 & ~n25941;
  assign n25943 = ~n25928 & ~n25934;
  assign n25944 = n6785 & n15111;
  assign n25945 = pi122  & n38631;
  assign n25946 = pi124  & n6800;
  assign n25947 = pi123  & n6802;
  assign n25948 = ~n25946 & ~n25947;
  assign n25949 = ~n25945 & ~n25947;
  assign n25950 = ~n25946 & n25949;
  assign n25951 = ~n25945 & n25948;
  assign n25952 = ~n25944 & n42274;
  assign n25953 = pi20  & ~n25952;
  assign n25954 = pi20  & ~n25953;
  assign n25955 = pi20  & n25952;
  assign n25956 = ~n25952 & ~n25953;
  assign n25957 = ~pi20  & ~n25952;
  assign n25958 = ~n42275 & ~n42276;
  assign n25959 = ~n25521 & ~n42261;
  assign n25960 = n25958 & n25959;
  assign n25961 = ~n25958 & ~n25959;
  assign n25962 = ~n25960 & ~n25961;
  assign n25963 = n4492 & n13057;
  assign n25964 = pi116  & n38208;
  assign n25965 = pi118  & n4507;
  assign n25966 = pi117  & n4509;
  assign n25967 = ~n25965 & ~n25966;
  assign n25968 = ~n25964 & ~n25966;
  assign n25969 = ~n25965 & n25968;
  assign n25970 = ~n25964 & n25967;
  assign n25971 = ~n25963 & n42277;
  assign n25972 = pi26  & ~n25971;
  assign n25973 = pi26  & ~n25972;
  assign n25974 = pi26  & n25971;
  assign n25975 = ~n25971 & ~n25972;
  assign n25976 = ~pi26  & ~n25971;
  assign n25977 = ~n42278 & ~n42279;
  assign n25978 = ~n25561 & ~n42257;
  assign n25979 = ~n25561 & ~n25863;
  assign n25980 = ~n25560 & ~n25978;
  assign n25981 = n25977 & n42280;
  assign n25982 = ~n25977 & ~n42280;
  assign n25983 = ~n25981 & ~n25982;
  assign n25984 = n523 & n607;
  assign n25985 = pi113  & n37489;
  assign n25986 = pi115  & n620;
  assign n25987 = pi114  & n622;
  assign n25988 = ~n25986 & ~n25987;
  assign n25989 = ~n25985 & ~n25987;
  assign n25990 = ~n25986 & n25989;
  assign n25991 = ~n25985 & n25988;
  assign n25992 = ~n25984 & n42281;
  assign n25993 = pi29  & ~n25992;
  assign n25994 = pi29  & ~n25993;
  assign n25995 = pi29  & n25992;
  assign n25996 = ~n25992 & ~n25993;
  assign n25997 = ~pi29  & ~n25992;
  assign n25998 = ~n42282 & ~n42283;
  assign n25999 = ~n25579 & n42254;
  assign n26000 = ~n25579 & ~n25855;
  assign n26001 = ~n25580 & ~n25999;
  assign n26002 = n25998 & n42284;
  assign n26003 = ~n25998 & ~n42284;
  assign n26004 = ~n26002 & ~n26003;
  assign n26005 = ~n25834 & ~n25837;
  assign n26006 = n691 & n8209;
  assign n26007 = pi104  & n37503;
  assign n26008 = pi106  & n704;
  assign n26009 = pi105  & n706;
  assign n26010 = ~n26008 & ~n26009;
  assign n26011 = ~n26007 & ~n26009;
  assign n26012 = ~n26008 & n26011;
  assign n26013 = ~n26007 & n26010;
  assign n26014 = ~n26006 & n42285;
  assign n26015 = pi38  & ~n26014;
  assign n26016 = pi38  & ~n26015;
  assign n26017 = pi38  & n26014;
  assign n26018 = ~n26014 & ~n26015;
  assign n26019 = ~pi38  & ~n26014;
  assign n26020 = ~n42286 & ~n42287;
  assign n26021 = ~n25814 & ~n25832;
  assign n26022 = n940 & n6474;
  assign n26023 = pi98  & n37541;
  assign n26024 = pi100  & n953;
  assign n26025 = pi99  & n955;
  assign n26026 = ~n26024 & ~n26025;
  assign n26027 = ~n26023 & ~n26025;
  assign n26028 = ~n26024 & n26027;
  assign n26029 = ~n26023 & n26026;
  assign n26030 = ~n26022 & n42288;
  assign n26031 = pi44  & ~n26030;
  assign n26032 = pi44  & ~n26031;
  assign n26033 = pi44  & n26030;
  assign n26034 = ~n26030 & ~n26031;
  assign n26035 = ~pi44  & ~n26030;
  assign n26036 = ~n42289 & ~n42290;
  assign n26037 = ~n25744 & ~n25747;
  assign n26038 = n594 & n1971;
  assign n26039 = pi89  & n37864;
  assign n26040 = pi91  & n1973;
  assign n26041 = pi90  & n1981;
  assign n26042 = ~n26040 & ~n26041;
  assign n26043 = ~n26039 & ~n26041;
  assign n26044 = ~n26040 & n26043;
  assign n26045 = ~n26039 & n26042;
  assign n26046 = ~n26038 & n42291;
  assign n26047 = pi53  & ~n26046;
  assign n26048 = pi53  & ~n26047;
  assign n26049 = pi53  & n26046;
  assign n26050 = ~n26046 & ~n26047;
  assign n26051 = ~pi53  & ~n26046;
  assign n26052 = ~n42292 & ~n42293;
  assign n26053 = ~n25721 & ~n25739;
  assign n26054 = ~n25672 & ~n25690;
  assign n26055 = n2134 & n12674;
  assign n26056 = pi80  & n40107;
  assign n26057 = pi82  & n12676;
  assign n26058 = pi81  & n12684;
  assign n26059 = ~n26057 & ~n26058;
  assign n26060 = ~n26056 & ~n26058;
  assign n26061 = ~n26057 & n26060;
  assign n26062 = ~n26056 & n26059;
  assign n26063 = ~n26055 & n42294;
  assign n26064 = pi62  & ~n26063;
  assign n26065 = pi62  & ~n26064;
  assign n26066 = pi62  & n26063;
  assign n26067 = ~n26063 & ~n26064;
  assign n26068 = ~pi62  & ~n26063;
  assign n26069 = ~n42295 & ~n42296;
  assign n26070 = pi79  & ~n40814;
  assign n26071 = pi78  & n18285;
  assign n26072 = ~n26070 & ~n26071;
  assign n26073 = ~pi14  & ~n26072;
  assign n26074 = pi14  & n26072;
  assign n26075 = ~pi14  & ~n26073;
  assign n26076 = ~pi14  & n26072;
  assign n26077 = ~n26072 & ~n26073;
  assign n26078 = pi14  & ~n26072;
  assign n26079 = ~n42297 & ~n42298;
  assign n26080 = ~n26073 & ~n26074;
  assign n26081 = ~n25183 & ~n42299;
  assign n26082 = n25183 & n42299;
  assign n26083 = ~n25183 & ~n26081;
  assign n26084 = ~n42299 & ~n26081;
  assign n26085 = ~n26083 & ~n26084;
  assign n26086 = ~n26081 & ~n26082;
  assign n26087 = ~n26069 & ~n42300;
  assign n26088 = n26069 & n42300;
  assign n26089 = ~n42300 & ~n26087;
  assign n26090 = n26069 & ~n42300;
  assign n26091 = ~n26069 & ~n26087;
  assign n26092 = ~n26069 & n42300;
  assign n26093 = ~n42301 & ~n42302;
  assign n26094 = ~n26087 & ~n26088;
  assign n26095 = n26054 & n42303;
  assign n26096 = ~n26054 & ~n42303;
  assign n26097 = ~n26095 & ~n26096;
  assign n26098 = n2804 & n7882;
  assign n26099 = pi83  & n39128;
  assign n26100 = pi85  & n7884;
  assign n26101 = pi84  & n7892;
  assign n26102 = ~n26100 & ~n26101;
  assign n26103 = ~n26099 & ~n26101;
  assign n26104 = ~n26100 & n26103;
  assign n26105 = ~n26099 & n26102;
  assign n26106 = ~n26098 & n42304;
  assign n26107 = pi59  & ~n26106;
  assign n26108 = pi59  & ~n26107;
  assign n26109 = pi59  & n26106;
  assign n26110 = ~n26106 & ~n26107;
  assign n26111 = ~pi59  & ~n26106;
  assign n26112 = ~n42305 & ~n42306;
  assign n26113 = n26097 & ~n26112;
  assign n26114 = ~n26097 & n26112;
  assign n26115 = n26097 & ~n26113;
  assign n26116 = n26097 & n26112;
  assign n26117 = ~n26112 & ~n26113;
  assign n26118 = ~n26097 & ~n26112;
  assign n26119 = ~n42307 & ~n42308;
  assign n26120 = ~n26113 & ~n26114;
  assign n26121 = ~n25693 & n25710;
  assign n26122 = ~n25693 & ~n25711;
  assign n26123 = ~n25694 & ~n26121;
  assign n26124 = n42309 & n42310;
  assign n26125 = ~n42309 & ~n42310;
  assign n26126 = ~n26124 & ~n26125;
  assign n26127 = n3354 & n4312;
  assign n26128 = pi86  & n38376;
  assign n26129 = pi88  & n4314;
  assign n26130 = pi87  & n4322;
  assign n26131 = ~n26129 & ~n26130;
  assign n26132 = ~n26128 & ~n26130;
  assign n26133 = ~n26129 & n26132;
  assign n26134 = ~n26128 & n26131;
  assign n26135 = ~n26127 & n42311;
  assign n26136 = pi56  & ~n26135;
  assign n26137 = pi56  & ~n26136;
  assign n26138 = pi56  & n26135;
  assign n26139 = ~n26135 & ~n26136;
  assign n26140 = ~pi56  & ~n26135;
  assign n26141 = ~n42312 & ~n42313;
  assign n26142 = n26126 & ~n26141;
  assign n26143 = ~n26126 & n26141;
  assign n26144 = ~n26142 & ~n26143;
  assign n26145 = n26053 & ~n26144;
  assign n26146 = ~n26053 & ~n26143;
  assign n26147 = ~n26142 & n26146;
  assign n26148 = ~n26053 & ~n26142;
  assign n26149 = ~n26143 & n26148;
  assign n26150 = ~n26053 & n26144;
  assign n26151 = ~n26053 & ~n42314;
  assign n26152 = ~n26053 & ~n26144;
  assign n26153 = n26053 & ~n26142;
  assign n26154 = ~n26142 & ~n42314;
  assign n26155 = ~n26143 & ~n26153;
  assign n26156 = ~n26143 & n42316;
  assign n26157 = n26053 & n26144;
  assign n26158 = ~n42315 & ~n42317;
  assign n26159 = ~n26145 & ~n42314;
  assign n26160 = ~n26052 & ~n42318;
  assign n26161 = n26052 & n42318;
  assign n26162 = ~n42318 & ~n26160;
  assign n26163 = ~n26052 & ~n26160;
  assign n26164 = ~n26162 & ~n26163;
  assign n26165 = ~n26160 & ~n26161;
  assign n26166 = n26037 & n42319;
  assign n26167 = ~n26037 & ~n42319;
  assign n26168 = ~n26166 & ~n26167;
  assign n26169 = n894 & n4524;
  assign n26170 = pi92  & n37580;
  assign n26171 = pi94  & n896;
  assign n26172 = pi93  & n904;
  assign n26173 = ~n26171 & ~n26172;
  assign n26174 = ~n26170 & ~n26172;
  assign n26175 = ~n26171 & n26174;
  assign n26176 = ~n26170 & n26173;
  assign n26177 = ~n26169 & n42320;
  assign n26178 = pi50  & ~n26177;
  assign n26179 = pi50  & ~n26178;
  assign n26180 = pi50  & n26177;
  assign n26181 = ~n26177 & ~n26178;
  assign n26182 = ~pi50  & ~n26177;
  assign n26183 = ~n42321 & ~n42322;
  assign n26184 = n26168 & ~n26183;
  assign n26185 = ~n26168 & n26183;
  assign n26186 = n26168 & ~n26184;
  assign n26187 = n26168 & n26183;
  assign n26188 = ~n26183 & ~n26184;
  assign n26189 = ~n26168 & ~n26183;
  assign n26190 = ~n42323 & ~n42324;
  assign n26191 = ~n26184 & ~n26185;
  assign n26192 = ~n25753 & n25770;
  assign n26193 = ~n25753 & ~n25771;
  assign n26194 = ~n25754 & ~n26192;
  assign n26195 = n42325 & n42326;
  assign n26196 = ~n42325 & ~n42326;
  assign n26197 = ~n26195 & ~n26196;
  assign n26198 = n785 & n5630;
  assign n26199 = pi95  & n37520;
  assign n26200 = pi97  & n787;
  assign n26201 = pi96  & n795;
  assign n26202 = ~n26200 & ~n26201;
  assign n26203 = ~n26199 & ~n26201;
  assign n26204 = ~n26200 & n26203;
  assign n26205 = ~n26199 & n26202;
  assign n26206 = ~n26198 & n42327;
  assign n26207 = pi47  & ~n26206;
  assign n26208 = pi47  & ~n26207;
  assign n26209 = pi47  & n26206;
  assign n26210 = ~n26206 & ~n26207;
  assign n26211 = ~pi47  & ~n26206;
  assign n26212 = ~n42328 & ~n42329;
  assign n26213 = n26197 & ~n26212;
  assign n26214 = ~n26197 & n26212;
  assign n26215 = n26197 & ~n26213;
  assign n26216 = n26197 & n26212;
  assign n26217 = ~n26212 & ~n26213;
  assign n26218 = ~n26197 & ~n26212;
  assign n26219 = ~n42330 & ~n42331;
  assign n26220 = ~n26213 & ~n26214;
  assign n26221 = n25651 & ~n25777;
  assign n26222 = ~n25777 & ~n25785;
  assign n26223 = ~n25778 & ~n26221;
  assign n26224 = ~n42332 & ~n42333;
  assign n26225 = n42332 & n42333;
  assign n26226 = n42332 & ~n42333;
  assign n26227 = ~n42332 & n42333;
  assign n26228 = ~n26226 & ~n26227;
  assign n26229 = ~n26224 & ~n26225;
  assign n26230 = ~n26036 & ~n42334;
  assign n26231 = n26036 & n42334;
  assign n26232 = ~n26230 & ~n26231;
  assign n26233 = ~n25790 & n25806;
  assign n26234 = ~n25790 & ~n25807;
  assign n26235 = ~n25789 & ~n26233;
  assign n26236 = ~n26232 & n42335;
  assign n26237 = n26232 & ~n42335;
  assign n26238 = ~n26236 & ~n26237;
  assign n26239 = n733 & n6787;
  assign n26240 = pi101  & n37510;
  assign n26241 = pi103  & n746;
  assign n26242 = pi102  & n748;
  assign n26243 = ~n26241 & ~n26242;
  assign n26244 = ~n26240 & ~n26242;
  assign n26245 = ~n26241 & n26244;
  assign n26246 = ~n26240 & n26243;
  assign n26247 = ~n26239 & n42336;
  assign n26248 = pi41  & ~n26247;
  assign n26249 = pi41  & ~n26248;
  assign n26250 = pi41  & n26247;
  assign n26251 = ~n26247 & ~n26248;
  assign n26252 = ~pi41  & ~n26247;
  assign n26253 = ~n42337 & ~n42338;
  assign n26254 = n26238 & ~n26253;
  assign n26255 = ~n26238 & n26253;
  assign n26256 = n26238 & ~n26254;
  assign n26257 = n26238 & n26253;
  assign n26258 = ~n26253 & ~n26254;
  assign n26259 = ~n26238 & ~n26253;
  assign n26260 = ~n42339 & ~n42340;
  assign n26261 = ~n26254 & ~n26255;
  assign n26262 = ~n26021 & ~n42341;
  assign n26263 = n26021 & n42341;
  assign n26264 = ~n26021 & n42341;
  assign n26265 = n26021 & ~n42341;
  assign n26266 = ~n26264 & ~n26265;
  assign n26267 = ~n26262 & ~n26263;
  assign n26268 = ~n26020 & ~n42342;
  assign n26269 = n26020 & n42342;
  assign n26270 = ~n26268 & ~n26269;
  assign n26271 = n26005 & ~n26270;
  assign n26272 = ~n26005 & n26270;
  assign n26273 = ~n26271 & ~n26272;
  assign n26274 = n2104 & n9701;
  assign n26275 = pi107  & n37758;
  assign n26276 = pi109  & n2117;
  assign n26277 = pi108  & n2119;
  assign n26278 = ~n26276 & ~n26277;
  assign n26279 = ~n26275 & ~n26277;
  assign n26280 = ~n26276 & n26279;
  assign n26281 = ~n26275 & n26278;
  assign n26282 = ~n26274 & n42343;
  assign n26283 = pi35  & ~n26282;
  assign n26284 = pi35  & ~n26283;
  assign n26285 = pi35  & n26282;
  assign n26286 = ~n26282 & ~n26283;
  assign n26287 = ~pi35  & ~n26282;
  assign n26288 = ~n42344 & ~n42345;
  assign n26289 = n26273 & ~n26288;
  assign n26290 = ~n26273 & n26288;
  assign n26291 = n26273 & ~n26289;
  assign n26292 = n26273 & n26288;
  assign n26293 = ~n26288 & ~n26289;
  assign n26294 = ~n26273 & ~n26288;
  assign n26295 = ~n42346 & ~n42347;
  assign n26296 = ~n26289 & ~n26290;
  assign n26297 = n25617 & ~n25840;
  assign n26298 = ~n25840 & ~n25844;
  assign n26299 = ~n25841 & ~n26297;
  assign n26300 = n42348 & n42349;
  assign n26301 = ~n42348 & ~n42349;
  assign n26302 = ~n26300 & ~n26301;
  assign n26303 = n649 & n10844;
  assign n26304 = pi110  & n37496;
  assign n26305 = pi112  & n662;
  assign n26306 = pi111  & n664;
  assign n26307 = ~n26305 & ~n26306;
  assign n26308 = ~n26304 & ~n26306;
  assign n26309 = ~n26305 & n26308;
  assign n26310 = ~n26304 & n26307;
  assign n26311 = ~n26303 & n42350;
  assign n26312 = pi32  & ~n26311;
  assign n26313 = pi32  & ~n26312;
  assign n26314 = pi32  & n26311;
  assign n26315 = ~n26311 & ~n26312;
  assign n26316 = ~pi32  & ~n26311;
  assign n26317 = ~n42351 & ~n42352;
  assign n26318 = ~n25600 & n42253;
  assign n26319 = ~n25600 & ~n25849;
  assign n26320 = ~n25601 & ~n26318;
  assign n26321 = ~n26317 & ~n42353;
  assign n26322 = n26317 & n42353;
  assign n26323 = ~n42353 & ~n26321;
  assign n26324 = n26317 & ~n42353;
  assign n26325 = ~n26317 & ~n26321;
  assign n26326 = ~n26317 & n42353;
  assign n26327 = ~n42354 & ~n42355;
  assign n26328 = ~n26321 & ~n26322;
  assign n26329 = n26302 & ~n42356;
  assign n26330 = ~n26302 & n42356;
  assign n26331 = ~n26329 & ~n26330;
  assign n26332 = n26004 & ~n26330;
  assign n26333 = ~n26329 & n26332;
  assign n26334 = n26004 & n26331;
  assign n26335 = ~n26004 & ~n26331;
  assign n26336 = n26004 & ~n42357;
  assign n26337 = ~n26330 & ~n42357;
  assign n26338 = ~n26329 & n26337;
  assign n26339 = n26331 & ~n42357;
  assign n26340 = ~n26336 & ~n42358;
  assign n26341 = ~n42357 & ~n26335;
  assign n26342 = n25983 & ~n42359;
  assign n26343 = ~n25983 & n42359;
  assign n26344 = ~n26342 & ~n26343;
  assign n26345 = ~n25542 & ~n25871;
  assign n26346 = n5576 & n15091;
  assign n26347 = pi119  & n38406;
  assign n26348 = pi121  & n5591;
  assign n26349 = pi120  & n5593;
  assign n26350 = ~n26348 & ~n26349;
  assign n26351 = ~n26347 & ~n26349;
  assign n26352 = ~n26348 & n26351;
  assign n26353 = ~n26347 & n26350;
  assign n26354 = ~n26346 & n42360;
  assign n26355 = pi23  & ~n26354;
  assign n26356 = pi23  & ~n26355;
  assign n26357 = pi23  & n26354;
  assign n26358 = ~n26354 & ~n26355;
  assign n26359 = ~pi23  & ~n26354;
  assign n26360 = ~n42361 & ~n42362;
  assign n26361 = ~n26345 & ~n26360;
  assign n26362 = n26345 & n26360;
  assign n26363 = ~n26345 & n26360;
  assign n26364 = n26345 & ~n26360;
  assign n26365 = ~n26363 & ~n26364;
  assign n26366 = ~n26361 & ~n26362;
  assign n26367 = ~n26343 & ~n42363;
  assign n26368 = ~n26342 & n26367;
  assign n26369 = n26344 & ~n42363;
  assign n26370 = ~n26344 & n42363;
  assign n26371 = ~n42363 & ~n42364;
  assign n26372 = ~n26344 & ~n42363;
  assign n26373 = n26344 & ~n42364;
  assign n26374 = ~n26343 & ~n42364;
  assign n26375 = ~n26342 & n26374;
  assign n26376 = n26344 & n42363;
  assign n26377 = ~n42365 & ~n42366;
  assign n26378 = ~n42364 & ~n26370;
  assign n26379 = n25962 & ~n42367;
  assign n26380 = ~n25962 & n42367;
  assign n26381 = ~n26379 & ~n26380;
  assign n26382 = ~n25900 & ~n25908;
  assign n26383 = n8175 & n40885;
  assign n26384 = pi125  & n38895;
  assign n26385 = pi127  & n8190;
  assign n26386 = pi126  & n8192;
  assign n26387 = ~n26385 & ~n26386;
  assign n26388 = ~n26384 & ~n26386;
  assign n26389 = ~n26385 & n26388;
  assign n26390 = ~n26384 & n26387;
  assign n26391 = ~n26383 & n42368;
  assign n26392 = pi17  & ~n26391;
  assign n26393 = pi17  & ~n26392;
  assign n26394 = pi17  & n26391;
  assign n26395 = ~n26391 & ~n26392;
  assign n26396 = ~pi17  & ~n26391;
  assign n26397 = ~n42369 & ~n42370;
  assign n26398 = ~n26382 & ~n26397;
  assign n26399 = n26382 & n26397;
  assign n26400 = ~n26382 & ~n26398;
  assign n26401 = ~n26382 & n26397;
  assign n26402 = ~n26397 & ~n26398;
  assign n26403 = n26382 & ~n26397;
  assign n26404 = ~n42371 & ~n42372;
  assign n26405 = ~n26398 & ~n26399;
  assign n26406 = ~n26380 & ~n42373;
  assign n26407 = ~n26379 & n26406;
  assign n26408 = n26381 & ~n42373;
  assign n26409 = ~n26381 & n42373;
  assign n26410 = ~n42373 & ~n42374;
  assign n26411 = ~n26380 & ~n42374;
  assign n26412 = ~n26379 & n26411;
  assign n26413 = n26381 & ~n42374;
  assign n26414 = ~n26410 & ~n42375;
  assign n26415 = ~n42374 & ~n26409;
  assign n26416 = n25943 & n42376;
  assign n26417 = ~n25943 & ~n42376;
  assign n26418 = ~n26416 & ~n26417;
  assign n26419 = ~n25937 & ~n25940;
  assign n26420 = n26418 & ~n26419;
  assign n26421 = ~n26418 & n26419;
  assign po78  = ~n26420 & ~n26421;
  assign n26423 = ~n26398 & ~n42374;
  assign n26424 = ~n25961 & ~n26379;
  assign n26425 = n8175 & n40891;
  assign n26426 = pi126  & n38895;
  assign n26427 = pi127  & n8192;
  assign n26428 = ~n26426 & ~n26427;
  assign n26429 = ~n8175 & n26428;
  assign n26430 = ~n40891 & n26428;
  assign n26431 = ~n26429 & ~n26430;
  assign n26432 = ~n26425 & n26428;
  assign n26433 = pi17  & ~n42377;
  assign n26434 = ~pi17  & n42377;
  assign n26435 = ~n26433 & ~n26434;
  assign n26436 = ~n26424 & ~n26435;
  assign n26437 = n26424 & n26435;
  assign n26438 = ~n26436 & ~n26437;
  assign n26439 = n6785 & n15068;
  assign n26440 = pi123  & n38631;
  assign n26441 = pi125  & n6800;
  assign n26442 = pi124  & n6802;
  assign n26443 = ~n26441 & ~n26442;
  assign n26444 = ~n26440 & ~n26442;
  assign n26445 = ~n26441 & n26444;
  assign n26446 = ~n26440 & n26443;
  assign n26447 = ~n26439 & n42378;
  assign n26448 = pi20  & ~n26447;
  assign n26449 = pi20  & ~n26448;
  assign n26450 = pi20  & n26447;
  assign n26451 = ~n26447 & ~n26448;
  assign n26452 = ~pi20  & ~n26447;
  assign n26453 = ~n42379 & ~n42380;
  assign n26454 = ~n26361 & ~n42364;
  assign n26455 = n26453 & n26454;
  assign n26456 = ~n26453 & ~n26454;
  assign n26457 = ~n26455 & ~n26456;
  assign n26458 = ~n25982 & ~n26342;
  assign n26459 = n5576 & n15049;
  assign n26460 = pi120  & n38406;
  assign n26461 = pi122  & n5591;
  assign n26462 = pi121  & n5593;
  assign n26463 = ~n26461 & ~n26462;
  assign n26464 = ~n26460 & ~n26462;
  assign n26465 = ~n26461 & n26464;
  assign n26466 = ~n26460 & n26463;
  assign n26467 = ~n5576 & n42381;
  assign n26468 = ~n15049 & n42381;
  assign n26469 = ~n26467 & ~n26468;
  assign n26470 = ~n26459 & n42381;
  assign n26471 = pi23  & ~n42382;
  assign n26472 = ~pi23  & n42382;
  assign n26473 = ~n26471 & ~n26472;
  assign n26474 = ~n26458 & ~n26473;
  assign n26475 = n26458 & n26473;
  assign n26476 = ~n26474 & ~n26475;
  assign n26477 = n4492 & n13027;
  assign n26478 = pi117  & n38208;
  assign n26479 = pi119  & n4507;
  assign n26480 = pi118  & n4509;
  assign n26481 = ~n26479 & ~n26480;
  assign n26482 = ~n26478 & ~n26480;
  assign n26483 = ~n26479 & n26482;
  assign n26484 = ~n26478 & n26481;
  assign n26485 = ~n26477 & n42383;
  assign n26486 = pi26  & ~n26485;
  assign n26487 = pi26  & ~n26486;
  assign n26488 = pi26  & n26485;
  assign n26489 = ~n26485 & ~n26486;
  assign n26490 = ~pi26  & ~n26485;
  assign n26491 = ~n42384 & ~n42385;
  assign n26492 = ~n26003 & ~n42357;
  assign n26493 = n26491 & n26492;
  assign n26494 = ~n26491 & ~n26492;
  assign n26495 = ~n26493 & ~n26494;
  assign n26496 = n649 & n11276;
  assign n26497 = pi111  & n37496;
  assign n26498 = pi113  & n662;
  assign n26499 = pi112  & n664;
  assign n26500 = ~n26498 & ~n26499;
  assign n26501 = ~n26497 & ~n26499;
  assign n26502 = ~n26498 & n26501;
  assign n26503 = ~n26497 & n26500;
  assign n26504 = ~n26496 & n42386;
  assign n26505 = pi32  & ~n26504;
  assign n26506 = pi32  & ~n26505;
  assign n26507 = pi32  & n26504;
  assign n26508 = ~n26504 & ~n26505;
  assign n26509 = ~pi32  & ~n26504;
  assign n26510 = ~n42387 & ~n42388;
  assign n26511 = ~n26289 & ~n26301;
  assign n26512 = n26510 & n26511;
  assign n26513 = ~n26510 & ~n26511;
  assign n26514 = ~n26512 & ~n26513;
  assign n26515 = ~n26268 & ~n26272;
  assign n26516 = ~n26254 & ~n26262;
  assign n26517 = n733 & n8136;
  assign n26518 = pi102  & n37510;
  assign n26519 = pi104  & n746;
  assign n26520 = pi103  & n748;
  assign n26521 = ~n26519 & ~n26520;
  assign n26522 = ~n26518 & ~n26520;
  assign n26523 = ~n26519 & n26522;
  assign n26524 = ~n26518 & n26521;
  assign n26525 = ~n26517 & n42389;
  assign n26526 = pi41  & ~n26525;
  assign n26527 = pi41  & ~n26526;
  assign n26528 = pi41  & n26525;
  assign n26529 = ~n26525 & ~n26526;
  assign n26530 = ~pi41  & ~n26525;
  assign n26531 = ~n42390 & ~n42391;
  assign n26532 = ~n26230 & ~n26237;
  assign n26533 = n940 & n6839;
  assign n26534 = pi99  & n37541;
  assign n26535 = pi101  & n953;
  assign n26536 = pi100  & n955;
  assign n26537 = ~n26535 & ~n26536;
  assign n26538 = ~n26534 & ~n26536;
  assign n26539 = ~n26535 & n26538;
  assign n26540 = ~n26534 & n26537;
  assign n26541 = ~n26533 & n42392;
  assign n26542 = pi44  & ~n26541;
  assign n26543 = pi44  & ~n26542;
  assign n26544 = pi44  & n26541;
  assign n26545 = ~n26541 & ~n26542;
  assign n26546 = ~pi44  & ~n26541;
  assign n26547 = ~n42393 & ~n42394;
  assign n26548 = ~n26213 & ~n26224;
  assign n26549 = ~n26184 & ~n26196;
  assign n26550 = n1971 & n4453;
  assign n26551 = pi90  & n37864;
  assign n26552 = pi92  & n1973;
  assign n26553 = pi91  & n1981;
  assign n26554 = ~n26552 & ~n26553;
  assign n26555 = ~n26551 & ~n26553;
  assign n26556 = ~n26552 & n26555;
  assign n26557 = ~n26551 & n26554;
  assign n26558 = ~n26550 & n42395;
  assign n26559 = pi53  & ~n26558;
  assign n26560 = pi53  & ~n26559;
  assign n26561 = pi53  & n26558;
  assign n26562 = ~n26558 & ~n26559;
  assign n26563 = ~pi53  & ~n26558;
  assign n26564 = ~n42396 & ~n42397;
  assign n26565 = ~n26113 & ~n26125;
  assign n26566 = ~n26087 & ~n26096;
  assign n26567 = ~n26073 & ~n26081;
  assign n26568 = pi80  & ~n40814;
  assign n26569 = pi79  & n18285;
  assign n26570 = ~n26568 & ~n26569;
  assign n26571 = n26567 & ~n26570;
  assign n26572 = ~n26567 & n26570;
  assign n26573 = ~n26571 & ~n26572;
  assign n26574 = n2091 & n12674;
  assign n26575 = pi81  & n40107;
  assign n26576 = pi83  & n12676;
  assign n26577 = pi82  & n12684;
  assign n26578 = ~n26576 & ~n26577;
  assign n26579 = ~n26575 & ~n26577;
  assign n26580 = ~n26576 & n26579;
  assign n26581 = ~n26575 & n26578;
  assign n26582 = ~n12674 & n42398;
  assign n26583 = ~n2091 & n42398;
  assign n26584 = ~n26582 & ~n26583;
  assign n26585 = ~n26574 & n42398;
  assign n26586 = pi62  & ~n42399;
  assign n26587 = ~pi62  & n42399;
  assign n26588 = ~n26586 & ~n26587;
  assign n26589 = n26573 & ~n26588;
  assign n26590 = ~n26573 & n26588;
  assign n26591 = ~n26589 & ~n26590;
  assign n26592 = ~n26566 & n26591;
  assign n26593 = n26566 & ~n26591;
  assign n26594 = ~n26592 & ~n26593;
  assign n26595 = n2779 & n7882;
  assign n26596 = pi84  & n39128;
  assign n26597 = pi86  & n7884;
  assign n26598 = pi85  & n7892;
  assign n26599 = ~n26597 & ~n26598;
  assign n26600 = ~n26596 & ~n26598;
  assign n26601 = ~n26597 & n26600;
  assign n26602 = ~n26596 & n26599;
  assign n26603 = ~n26595 & n42400;
  assign n26604 = pi59  & ~n26603;
  assign n26605 = pi59  & ~n26604;
  assign n26606 = pi59  & n26603;
  assign n26607 = ~n26603 & ~n26604;
  assign n26608 = ~pi59  & ~n26603;
  assign n26609 = ~n42401 & ~n42402;
  assign n26610 = n26594 & ~n26609;
  assign n26611 = ~n26594 & n26609;
  assign n26612 = n26594 & ~n26610;
  assign n26613 = ~n26609 & ~n26610;
  assign n26614 = ~n26612 & ~n26613;
  assign n26615 = ~n26610 & ~n26611;
  assign n26616 = n26565 & n42403;
  assign n26617 = ~n26565 & ~n42403;
  assign n26618 = ~n26616 & ~n26617;
  assign n26619 = n3591 & n4312;
  assign n26620 = pi87  & n38376;
  assign n26621 = pi89  & n4314;
  assign n26622 = pi88  & n4322;
  assign n26623 = ~n26621 & ~n26622;
  assign n26624 = ~n26620 & ~n26622;
  assign n26625 = ~n26621 & n26624;
  assign n26626 = ~n26620 & n26623;
  assign n26627 = ~n26619 & n42404;
  assign n26628 = pi56  & ~n26627;
  assign n26629 = pi56  & ~n26628;
  assign n26630 = pi56  & n26627;
  assign n26631 = ~n26627 & ~n26628;
  assign n26632 = ~pi56  & ~n26627;
  assign n26633 = ~n42405 & ~n42406;
  assign n26634 = ~n26618 & n26633;
  assign n26635 = n26618 & ~n26633;
  assign n26636 = n26618 & ~n26635;
  assign n26637 = ~n26633 & ~n26635;
  assign n26638 = ~n26636 & ~n26637;
  assign n26639 = ~n26634 & ~n26635;
  assign n26640 = ~n42316 & ~n42407;
  assign n26641 = n42316 & n42407;
  assign n26642 = ~n42316 & n42407;
  assign n26643 = n42316 & ~n42407;
  assign n26644 = ~n26642 & ~n26643;
  assign n26645 = ~n26640 & ~n26641;
  assign n26646 = n26564 & n42408;
  assign n26647 = ~n26564 & ~n42408;
  assign n26648 = ~n26646 & ~n26647;
  assign n26649 = ~n26160 & ~n26167;
  assign n26650 = n26648 & ~n26649;
  assign n26651 = ~n26648 & n26649;
  assign n26652 = ~n26650 & ~n26651;
  assign n26653 = n894 & n4494;
  assign n26654 = pi93  & n37580;
  assign n26655 = pi95  & n896;
  assign n26656 = pi94  & n904;
  assign n26657 = ~n26655 & ~n26656;
  assign n26658 = ~n26654 & ~n26656;
  assign n26659 = ~n26655 & n26658;
  assign n26660 = ~n26654 & n26657;
  assign n26661 = ~n26653 & n42409;
  assign n26662 = pi50  & ~n26661;
  assign n26663 = pi50  & ~n26662;
  assign n26664 = pi50  & n26661;
  assign n26665 = ~n26661 & ~n26662;
  assign n26666 = ~pi50  & ~n26661;
  assign n26667 = ~n42410 & ~n42411;
  assign n26668 = ~n26652 & n26667;
  assign n26669 = n26652 & ~n26667;
  assign n26670 = n26652 & ~n26669;
  assign n26671 = ~n26667 & ~n26669;
  assign n26672 = ~n26670 & ~n26671;
  assign n26673 = ~n26668 & ~n26669;
  assign n26674 = n26549 & n42412;
  assign n26675 = ~n26549 & ~n42412;
  assign n26676 = ~n26674 & ~n26675;
  assign n26677 = n785 & n5610;
  assign n26678 = pi96  & n37520;
  assign n26679 = pi98  & n787;
  assign n26680 = pi97  & n795;
  assign n26681 = ~n26679 & ~n26680;
  assign n26682 = ~n26678 & ~n26680;
  assign n26683 = ~n26679 & n26682;
  assign n26684 = ~n26678 & n26681;
  assign n26685 = ~n26677 & n42413;
  assign n26686 = pi47  & ~n26685;
  assign n26687 = pi47  & ~n26686;
  assign n26688 = pi47  & n26685;
  assign n26689 = ~n26685 & ~n26686;
  assign n26690 = ~pi47  & ~n26685;
  assign n26691 = ~n42414 & ~n42415;
  assign n26692 = ~n26676 & n26691;
  assign n26693 = n26676 & ~n26691;
  assign n26694 = ~n26692 & ~n26693;
  assign n26695 = ~n26548 & n26694;
  assign n26696 = n26548 & ~n26694;
  assign n26697 = ~n26548 & ~n26695;
  assign n26698 = n26694 & ~n26695;
  assign n26699 = ~n26697 & ~n26698;
  assign n26700 = ~n26695 & ~n26696;
  assign n26701 = ~n26547 & ~n42416;
  assign n26702 = n26547 & ~n26698;
  assign n26703 = ~n26697 & n26702;
  assign n26704 = n26547 & n42416;
  assign n26705 = ~n26701 & ~n42417;
  assign n26706 = ~n26532 & n26705;
  assign n26707 = n26532 & ~n26705;
  assign n26708 = ~n26532 & ~n26706;
  assign n26709 = n26705 & ~n26706;
  assign n26710 = ~n26708 & ~n26709;
  assign n26711 = ~n26706 & ~n26707;
  assign n26712 = ~n26531 & ~n42418;
  assign n26713 = n26531 & ~n26709;
  assign n26714 = ~n26708 & n26713;
  assign n26715 = n26531 & n42418;
  assign n26716 = ~n26712 & ~n42419;
  assign n26717 = ~n26516 & n26716;
  assign n26718 = n26516 & ~n26716;
  assign n26719 = ~n26717 & ~n26718;
  assign n26720 = n691 & n8177;
  assign n26721 = pi105  & n37503;
  assign n26722 = pi107  & n704;
  assign n26723 = pi106  & n706;
  assign n26724 = ~n26722 & ~n26723;
  assign n26725 = ~n26721 & ~n26723;
  assign n26726 = ~n26722 & n26725;
  assign n26727 = ~n26721 & n26724;
  assign n26728 = ~n26720 & n42420;
  assign n26729 = pi38  & ~n26728;
  assign n26730 = pi38  & ~n26729;
  assign n26731 = pi38  & n26728;
  assign n26732 = ~n26728 & ~n26729;
  assign n26733 = ~pi38  & ~n26728;
  assign n26734 = ~n42421 & ~n42422;
  assign n26735 = n26719 & ~n26734;
  assign n26736 = ~n26719 & n26734;
  assign n26737 = n26719 & ~n26735;
  assign n26738 = ~n26734 & ~n26735;
  assign n26739 = ~n26737 & ~n26738;
  assign n26740 = ~n26735 & ~n26736;
  assign n26741 = n26515 & n42423;
  assign n26742 = ~n26515 & ~n42423;
  assign n26743 = ~n26741 & ~n26742;
  assign n26744 = n2104 & n9678;
  assign n26745 = pi108  & n37758;
  assign n26746 = pi110  & n2117;
  assign n26747 = pi109  & n2119;
  assign n26748 = ~n26746 & ~n26747;
  assign n26749 = ~n26745 & ~n26747;
  assign n26750 = ~n26746 & n26749;
  assign n26751 = ~n26745 & n26748;
  assign n26752 = ~n26744 & n42424;
  assign n26753 = pi35  & ~n26752;
  assign n26754 = pi35  & ~n26753;
  assign n26755 = pi35  & n26752;
  assign n26756 = ~n26752 & ~n26753;
  assign n26757 = ~pi35  & ~n26752;
  assign n26758 = ~n42425 & ~n42426;
  assign n26759 = ~n26743 & n26758;
  assign n26760 = n26743 & ~n26758;
  assign n26761 = n26743 & ~n26760;
  assign n26762 = ~n26758 & ~n26760;
  assign n26763 = ~n26761 & ~n26762;
  assign n26764 = ~n26759 & ~n26760;
  assign n26765 = n26514 & ~n42427;
  assign n26766 = ~n26514 & n42427;
  assign n26767 = ~n26765 & ~n26766;
  assign n26768 = n607 & n12530;
  assign n26769 = pi114  & n37489;
  assign n26770 = pi116  & n620;
  assign n26771 = pi115  & n622;
  assign n26772 = ~n26770 & ~n26771;
  assign n26773 = ~n26769 & ~n26771;
  assign n26774 = ~n26770 & n26773;
  assign n26775 = ~n26769 & n26772;
  assign n26776 = ~n26768 & n42428;
  assign n26777 = pi29  & ~n26776;
  assign n26778 = pi29  & ~n26777;
  assign n26779 = pi29  & n26776;
  assign n26780 = ~n26776 & ~n26777;
  assign n26781 = ~pi29  & ~n26776;
  assign n26782 = ~n42429 & ~n42430;
  assign n26783 = ~n26321 & ~n26329;
  assign n26784 = ~n26782 & ~n26783;
  assign n26785 = n26782 & n26783;
  assign n26786 = ~n26782 & ~n26784;
  assign n26787 = ~n26782 & n26783;
  assign n26788 = ~n26783 & ~n26784;
  assign n26789 = n26782 & ~n26783;
  assign n26790 = ~n42431 & ~n42432;
  assign n26791 = ~n26784 & ~n26785;
  assign n26792 = ~n26766 & ~n42433;
  assign n26793 = ~n26765 & n26792;
  assign n26794 = n26767 & ~n42433;
  assign n26795 = ~n26767 & n42433;
  assign n26796 = ~n42433 & ~n42434;
  assign n26797 = ~n26766 & ~n42434;
  assign n26798 = ~n26765 & n26797;
  assign n26799 = n26767 & ~n42434;
  assign n26800 = ~n26796 & ~n42435;
  assign n26801 = ~n42434 & ~n26795;
  assign n26802 = n26495 & ~n42436;
  assign n26803 = ~n26495 & n42436;
  assign n26804 = ~n26802 & ~n26803;
  assign n26805 = n26476 & ~n26803;
  assign n26806 = ~n26802 & n26805;
  assign n26807 = n26476 & n26804;
  assign n26808 = ~n26476 & ~n26804;
  assign n26809 = n26476 & ~n42437;
  assign n26810 = ~n26803 & ~n42437;
  assign n26811 = ~n26802 & n26810;
  assign n26812 = n26804 & ~n42437;
  assign n26813 = ~n26809 & ~n42438;
  assign n26814 = ~n42437 & ~n26808;
  assign n26815 = n26457 & ~n42439;
  assign n26816 = ~n26457 & n42439;
  assign n26817 = ~n26815 & ~n26816;
  assign n26818 = n26438 & ~n26816;
  assign n26819 = ~n26815 & n26818;
  assign n26820 = n26438 & n26817;
  assign n26821 = ~n26816 & ~n42440;
  assign n26822 = ~n26815 & n26821;
  assign n26823 = n26817 & ~n42440;
  assign n26824 = ~n26438 & n26817;
  assign n26825 = n26438 & ~n42440;
  assign n26826 = n26438 & ~n26817;
  assign n26827 = ~n42441 & ~n42442;
  assign n26828 = n26423 & n26827;
  assign n26829 = ~n26423 & ~n26827;
  assign n26830 = ~n26828 & ~n26829;
  assign n26831 = ~n26417 & ~n26420;
  assign n26832 = n26830 & ~n26831;
  assign n26833 = ~n26830 & n26831;
  assign po79  = ~n26832 & ~n26833;
  assign n26835 = ~n26829 & ~n26832;
  assign n26836 = n6785 & n15021;
  assign n26837 = pi124  & n38631;
  assign n26838 = pi126  & n6800;
  assign n26839 = pi125  & n6802;
  assign n26840 = ~n26838 & ~n26839;
  assign n26841 = ~n26837 & ~n26839;
  assign n26842 = ~n26838 & n26841;
  assign n26843 = ~n26837 & n26840;
  assign n26844 = ~n26836 & n42443;
  assign n26845 = pi20  & ~n26844;
  assign n26846 = pi20  & ~n26845;
  assign n26847 = pi20  & n26844;
  assign n26848 = ~n26844 & ~n26845;
  assign n26849 = ~pi20  & ~n26844;
  assign n26850 = ~n42444 & ~n42445;
  assign n26851 = ~n26474 & ~n42437;
  assign n26852 = n26850 & n26851;
  assign n26853 = ~n26850 & ~n26851;
  assign n26854 = ~n26852 & ~n26853;
  assign n26855 = n4492 & n14913;
  assign n26856 = pi118  & n38208;
  assign n26857 = pi120  & n4507;
  assign n26858 = pi119  & n4509;
  assign n26859 = ~n26857 & ~n26858;
  assign n26860 = ~n26856 & ~n26858;
  assign n26861 = ~n26857 & n26860;
  assign n26862 = ~n26856 & n26859;
  assign n26863 = ~n26855 & n42446;
  assign n26864 = pi26  & ~n26863;
  assign n26865 = pi26  & ~n26864;
  assign n26866 = pi26  & n26863;
  assign n26867 = ~n26863 & ~n26864;
  assign n26868 = ~pi26  & ~n26863;
  assign n26869 = ~n42447 & ~n42448;
  assign n26870 = ~n26784 & ~n42434;
  assign n26871 = n26869 & n26870;
  assign n26872 = ~n26869 & ~n26870;
  assign n26873 = ~n26871 & ~n26872;
  assign n26874 = n649 & n11258;
  assign n26875 = pi112  & n37496;
  assign n26876 = pi114  & n662;
  assign n26877 = pi113  & n664;
  assign n26878 = ~n26876 & ~n26877;
  assign n26879 = ~n26875 & ~n26877;
  assign n26880 = ~n26876 & n26879;
  assign n26881 = ~n26875 & n26878;
  assign n26882 = ~n26874 & n42449;
  assign n26883 = pi32  & ~n26882;
  assign n26884 = pi32  & ~n26883;
  assign n26885 = pi32  & n26882;
  assign n26886 = ~n26882 & ~n26883;
  assign n26887 = ~pi32  & ~n26882;
  assign n26888 = ~n42450 & ~n42451;
  assign n26889 = ~n26742 & n26758;
  assign n26890 = ~n26742 & ~n26760;
  assign n26891 = ~n26741 & ~n26889;
  assign n26892 = n26888 & n42452;
  assign n26893 = ~n26888 & ~n42452;
  assign n26894 = ~n26892 & ~n26893;
  assign n26895 = n691 & n9277;
  assign n26896 = pi106  & n37503;
  assign n26897 = pi108  & n704;
  assign n26898 = pi107  & n706;
  assign n26899 = ~n26897 & ~n26898;
  assign n26900 = ~n26896 & ~n26898;
  assign n26901 = ~n26897 & n26900;
  assign n26902 = ~n26896 & n26899;
  assign n26903 = ~n26895 & n42453;
  assign n26904 = pi38  & ~n26903;
  assign n26905 = pi38  & ~n26904;
  assign n26906 = pi38  & n26903;
  assign n26907 = ~n26903 & ~n26904;
  assign n26908 = ~pi38  & ~n26903;
  assign n26909 = ~n42454 & ~n42455;
  assign n26910 = ~n26706 & ~n26712;
  assign n26911 = n733 & n8229;
  assign n26912 = pi103  & n37510;
  assign n26913 = pi105  & n746;
  assign n26914 = pi104  & n748;
  assign n26915 = ~n26913 & ~n26914;
  assign n26916 = ~n26912 & ~n26914;
  assign n26917 = ~n26913 & n26916;
  assign n26918 = ~n26912 & n26915;
  assign n26919 = ~n26911 & n42456;
  assign n26920 = pi41  & ~n26919;
  assign n26921 = pi41  & ~n26920;
  assign n26922 = pi41  & n26919;
  assign n26923 = ~n26919 & ~n26920;
  assign n26924 = ~pi41  & ~n26919;
  assign n26925 = ~n42457 & ~n42458;
  assign n26926 = ~n26695 & ~n26701;
  assign n26927 = n940 & n6819;
  assign n26928 = pi100  & n37541;
  assign n26929 = pi102  & n953;
  assign n26930 = pi101  & n955;
  assign n26931 = ~n26929 & ~n26930;
  assign n26932 = ~n26928 & ~n26930;
  assign n26933 = ~n26929 & n26932;
  assign n26934 = ~n26928 & n26931;
  assign n26935 = ~n26927 & n42459;
  assign n26936 = pi44  & ~n26935;
  assign n26937 = pi44  & ~n26936;
  assign n26938 = pi44  & n26935;
  assign n26939 = ~n26935 & ~n26936;
  assign n26940 = ~pi44  & ~n26935;
  assign n26941 = ~n42460 & ~n42461;
  assign n26942 = ~n26675 & ~n26693;
  assign n26943 = ~n26651 & ~n26667;
  assign n26944 = ~n26650 & ~n26669;
  assign n26945 = ~n26650 & ~n26943;
  assign n26946 = n894 & n5281;
  assign n26947 = pi94  & n37580;
  assign n26948 = pi96  & n896;
  assign n26949 = pi95  & n904;
  assign n26950 = ~n26948 & ~n26949;
  assign n26951 = ~n26947 & ~n26949;
  assign n26952 = ~n26948 & n26951;
  assign n26953 = ~n26947 & n26950;
  assign n26954 = ~n26946 & n42463;
  assign n26955 = pi50  & ~n26954;
  assign n26956 = pi50  & ~n26955;
  assign n26957 = pi50  & n26954;
  assign n26958 = ~n26954 & ~n26955;
  assign n26959 = ~pi50  & ~n26954;
  assign n26960 = ~n42464 & ~n42465;
  assign n26961 = ~n26640 & ~n26647;
  assign n26962 = n3566 & n4312;
  assign n26963 = pi88  & n38376;
  assign n26964 = pi90  & n4314;
  assign n26965 = pi89  & n4322;
  assign n26966 = ~n26964 & ~n26965;
  assign n26967 = ~n26963 & ~n26965;
  assign n26968 = ~n26964 & n26967;
  assign n26969 = ~n26963 & n26966;
  assign n26970 = ~n26962 & n42466;
  assign n26971 = pi56  & ~n26970;
  assign n26972 = pi56  & ~n26971;
  assign n26973 = pi56  & n26970;
  assign n26974 = ~n26970 & ~n26971;
  assign n26975 = ~pi56  & ~n26970;
  assign n26976 = ~n42467 & ~n42468;
  assign n26977 = ~n26572 & ~n26589;
  assign n26978 = n2591 & n12674;
  assign n26979 = pi82  & n40107;
  assign n26980 = pi84  & n12676;
  assign n26981 = pi83  & n12684;
  assign n26982 = ~n26980 & ~n26981;
  assign n26983 = ~n26979 & ~n26981;
  assign n26984 = ~n26980 & n26983;
  assign n26985 = ~n26979 & n26982;
  assign n26986 = ~n26978 & n42469;
  assign n26987 = pi62  & ~n26986;
  assign n26988 = pi62  & ~n26987;
  assign n26989 = pi62  & n26986;
  assign n26990 = ~n26986 & ~n26987;
  assign n26991 = ~pi62  & ~n26986;
  assign n26992 = ~n42470 & ~n42471;
  assign n26993 = pi81  & ~n40814;
  assign n26994 = pi80  & n18285;
  assign n26995 = ~n26993 & ~n26994;
  assign n26996 = n26570 & ~n26995;
  assign n26997 = ~n26570 & n26995;
  assign n26998 = ~n26996 & ~n26997;
  assign n26999 = ~n26992 & ~n26997;
  assign n27000 = ~n26996 & n26999;
  assign n27001 = ~n26992 & n26998;
  assign n27002 = n26992 & ~n26998;
  assign n27003 = ~n26992 & ~n42472;
  assign n27004 = ~n26997 & ~n42472;
  assign n27005 = ~n26996 & n27004;
  assign n27006 = ~n27003 & ~n27005;
  assign n27007 = ~n42472 & ~n27002;
  assign n27008 = n26977 & n42473;
  assign n27009 = ~n26977 & ~n42473;
  assign n27010 = ~n27008 & ~n27009;
  assign n27011 = n636 & n7882;
  assign n27012 = pi85  & n39128;
  assign n27013 = pi87  & n7884;
  assign n27014 = pi86  & n7892;
  assign n27015 = ~n27013 & ~n27014;
  assign n27016 = ~n27012 & ~n27014;
  assign n27017 = ~n27013 & n27016;
  assign n27018 = ~n27012 & n27015;
  assign n27019 = ~n27011 & n42474;
  assign n27020 = pi59  & ~n27019;
  assign n27021 = pi59  & ~n27020;
  assign n27022 = pi59  & n27019;
  assign n27023 = ~n27019 & ~n27020;
  assign n27024 = ~pi59  & ~n27019;
  assign n27025 = ~n42475 & ~n42476;
  assign n27026 = ~n27010 & n27025;
  assign n27027 = n27010 & ~n27025;
  assign n27028 = ~n27026 & ~n27027;
  assign n27029 = ~n26592 & n26609;
  assign n27030 = ~n26592 & ~n26610;
  assign n27031 = ~n26593 & ~n27029;
  assign n27032 = n27028 & ~n42477;
  assign n27033 = ~n27028 & n42477;
  assign n27034 = ~n27032 & ~n27033;
  assign n27035 = ~n26976 & n27034;
  assign n27036 = n26976 & ~n27034;
  assign n27037 = ~n27035 & ~n27036;
  assign n27038 = ~n26617 & n26633;
  assign n27039 = ~n26617 & ~n26635;
  assign n27040 = ~n26616 & ~n27038;
  assign n27041 = n27037 & ~n42478;
  assign n27042 = ~n27037 & n42478;
  assign n27043 = ~n27041 & ~n27042;
  assign n27044 = n1971 & n4544;
  assign n27045 = pi91  & n37864;
  assign n27046 = pi93  & n1973;
  assign n27047 = pi92  & n1981;
  assign n27048 = ~n27046 & ~n27047;
  assign n27049 = ~n27045 & ~n27047;
  assign n27050 = ~n27046 & n27049;
  assign n27051 = ~n27045 & n27048;
  assign n27052 = ~n27044 & n42479;
  assign n27053 = pi53  & ~n27052;
  assign n27054 = pi53  & ~n27053;
  assign n27055 = pi53  & n27052;
  assign n27056 = ~n27052 & ~n27053;
  assign n27057 = ~pi53  & ~n27052;
  assign n27058 = ~n42480 & ~n42481;
  assign n27059 = n27043 & ~n27058;
  assign n27060 = ~n27043 & n27058;
  assign n27061 = n27043 & ~n27059;
  assign n27062 = ~n27058 & ~n27059;
  assign n27063 = ~n27061 & ~n27062;
  assign n27064 = ~n27059 & ~n27060;
  assign n27065 = ~n26961 & ~n42482;
  assign n27066 = n26961 & n42482;
  assign n27067 = ~n42482 & ~n27065;
  assign n27068 = ~n26961 & ~n27065;
  assign n27069 = ~n27067 & ~n27068;
  assign n27070 = ~n27065 & ~n27066;
  assign n27071 = n26960 & ~n42483;
  assign n27072 = ~n26960 & n42483;
  assign n27073 = ~n26960 & ~n42483;
  assign n27074 = n26960 & n42483;
  assign n27075 = ~n27073 & ~n27074;
  assign n27076 = ~n27071 & ~n27072;
  assign n27077 = n42462 & ~n42484;
  assign n27078 = ~n42462 & n42484;
  assign n27079 = ~n27077 & ~n27078;
  assign n27080 = n785 & n5578;
  assign n27081 = pi97  & n37520;
  assign n27082 = pi99  & n787;
  assign n27083 = pi98  & n795;
  assign n27084 = ~n27082 & ~n27083;
  assign n27085 = ~n27081 & ~n27083;
  assign n27086 = ~n27082 & n27085;
  assign n27087 = ~n27081 & n27084;
  assign n27088 = ~n27080 & n42485;
  assign n27089 = pi47  & ~n27088;
  assign n27090 = pi47  & ~n27089;
  assign n27091 = pi47  & n27088;
  assign n27092 = ~n27088 & ~n27089;
  assign n27093 = ~pi47  & ~n27088;
  assign n27094 = ~n42486 & ~n42487;
  assign n27095 = n27079 & ~n27094;
  assign n27096 = ~n27079 & n27094;
  assign n27097 = n27079 & ~n27095;
  assign n27098 = ~n27094 & ~n27095;
  assign n27099 = ~n27097 & ~n27098;
  assign n27100 = ~n27095 & ~n27096;
  assign n27101 = ~n26942 & ~n42488;
  assign n27102 = n26942 & n42488;
  assign n27103 = ~n42488 & ~n27101;
  assign n27104 = ~n26942 & ~n27101;
  assign n27105 = ~n27103 & ~n27104;
  assign n27106 = ~n27101 & ~n27102;
  assign n27107 = ~n26941 & ~n42489;
  assign n27108 = n26941 & n42489;
  assign n27109 = n26941 & ~n42489;
  assign n27110 = ~n26941 & n42489;
  assign n27111 = ~n27109 & ~n27110;
  assign n27112 = ~n27107 & ~n27108;
  assign n27113 = ~n26926 & ~n42490;
  assign n27114 = n26926 & n42490;
  assign n27115 = ~n27113 & ~n27114;
  assign n27116 = ~n26925 & n27115;
  assign n27117 = n26925 & ~n27115;
  assign n27118 = ~n27116 & ~n27117;
  assign n27119 = ~n26910 & n27118;
  assign n27120 = n26910 & ~n27118;
  assign n27121 = ~n27119 & ~n27120;
  assign n27122 = ~n26909 & n27121;
  assign n27123 = n26909 & ~n27121;
  assign n27124 = ~n27122 & ~n27123;
  assign n27125 = ~n26717 & n26734;
  assign n27126 = ~n26717 & ~n26735;
  assign n27127 = ~n26718 & ~n27125;
  assign n27128 = n27124 & ~n42491;
  assign n27129 = ~n27124 & n42491;
  assign n27130 = ~n27128 & ~n27129;
  assign n27131 = n565 & n2104;
  assign n27132 = pi109  & n37758;
  assign n27133 = pi111  & n2117;
  assign n27134 = pi110  & n2119;
  assign n27135 = ~n27133 & ~n27134;
  assign n27136 = ~n27132 & ~n27134;
  assign n27137 = ~n27133 & n27136;
  assign n27138 = ~n27132 & n27135;
  assign n27139 = ~n27131 & n42492;
  assign n27140 = pi35  & ~n27139;
  assign n27141 = pi35  & ~n27140;
  assign n27142 = pi35  & n27139;
  assign n27143 = ~n27139 & ~n27140;
  assign n27144 = ~pi35  & ~n27139;
  assign n27145 = ~n42493 & ~n42494;
  assign n27146 = n27130 & ~n27145;
  assign n27147 = ~n27130 & n27145;
  assign n27148 = n27130 & ~n27146;
  assign n27149 = ~n27145 & ~n27146;
  assign n27150 = ~n27148 & ~n27149;
  assign n27151 = ~n27146 & ~n27147;
  assign n27152 = n26894 & ~n42495;
  assign n27153 = ~n26894 & n42495;
  assign n27154 = ~n27152 & ~n27153;
  assign n27155 = n607 & n13079;
  assign n27156 = pi115  & n37489;
  assign n27157 = pi117  & n620;
  assign n27158 = pi116  & n622;
  assign n27159 = ~n27157 & ~n27158;
  assign n27160 = ~n27156 & ~n27158;
  assign n27161 = ~n27157 & n27160;
  assign n27162 = ~n27156 & n27159;
  assign n27163 = ~n27155 & n42496;
  assign n27164 = pi29  & ~n27163;
  assign n27165 = pi29  & ~n27164;
  assign n27166 = pi29  & n27163;
  assign n27167 = ~n27163 & ~n27164;
  assign n27168 = ~pi29  & ~n27163;
  assign n27169 = ~n42497 & ~n42498;
  assign n27170 = ~n26513 & ~n26765;
  assign n27171 = ~n27169 & ~n27170;
  assign n27172 = n27169 & n27170;
  assign n27173 = ~n27169 & ~n27171;
  assign n27174 = ~n27169 & n27170;
  assign n27175 = ~n27170 & ~n27171;
  assign n27176 = n27169 & ~n27170;
  assign n27177 = ~n42499 & ~n42500;
  assign n27178 = ~n27171 & ~n27172;
  assign n27179 = ~n27153 & ~n42501;
  assign n27180 = ~n27152 & n27179;
  assign n27181 = n27154 & ~n42501;
  assign n27182 = ~n27154 & n42501;
  assign n27183 = ~n42501 & ~n42502;
  assign n27184 = ~n27153 & ~n42502;
  assign n27185 = ~n27152 & n27184;
  assign n27186 = n27154 & ~n42502;
  assign n27187 = ~n27183 & ~n42503;
  assign n27188 = ~n42502 & ~n27182;
  assign n27189 = n26873 & ~n42504;
  assign n27190 = ~n26873 & n42504;
  assign n27191 = ~n27189 & ~n27190;
  assign n27192 = n5576 & n14961;
  assign n27193 = pi121  & n38406;
  assign n27194 = pi123  & n5591;
  assign n27195 = pi122  & n5593;
  assign n27196 = ~n27194 & ~n27195;
  assign n27197 = ~n27193 & ~n27195;
  assign n27198 = ~n27194 & n27197;
  assign n27199 = ~n27193 & n27196;
  assign n27200 = ~n27192 & n42505;
  assign n27201 = pi23  & ~n27200;
  assign n27202 = pi23  & ~n27201;
  assign n27203 = pi23  & n27200;
  assign n27204 = ~n27200 & ~n27201;
  assign n27205 = ~pi23  & ~n27200;
  assign n27206 = ~n42506 & ~n42507;
  assign n27207 = ~n26494 & ~n26802;
  assign n27208 = ~n27206 & ~n27207;
  assign n27209 = n27206 & n27207;
  assign n27210 = ~n27206 & ~n27208;
  assign n27211 = ~n27206 & n27207;
  assign n27212 = ~n27207 & ~n27208;
  assign n27213 = n27206 & ~n27207;
  assign n27214 = ~n42508 & ~n42509;
  assign n27215 = ~n27208 & ~n27209;
  assign n27216 = ~n27190 & ~n42510;
  assign n27217 = ~n27189 & n27216;
  assign n27218 = n27191 & ~n42510;
  assign n27219 = ~n27191 & n42510;
  assign n27220 = ~n42510 & ~n42511;
  assign n27221 = ~n27191 & ~n42510;
  assign n27222 = n27191 & ~n42511;
  assign n27223 = ~n27190 & ~n42511;
  assign n27224 = ~n27189 & n27223;
  assign n27225 = n27191 & n42510;
  assign n27226 = ~n42512 & ~n42513;
  assign n27227 = ~n42511 & ~n27219;
  assign n27228 = ~n26854 & n42514;
  assign n27229 = n26854 & ~n42514;
  assign n27230 = ~n27228 & ~n27229;
  assign n27231 = ~n26456 & ~n26815;
  assign n27232 = n8175 & ~n18675;
  assign n27233 = ~n38895 & ~n27232;
  assign n27234 = pi127  & n38895;
  assign n27235 = n8175 & n18680;
  assign n27236 = ~n27234 & ~n27235;
  assign n27237 = pi127  & ~n27233;
  assign n27238 = pi17  & ~n42515;
  assign n27239 = pi17  & ~n27238;
  assign n27240 = pi17  & n42515;
  assign n27241 = ~n42515 & ~n27238;
  assign n27242 = ~pi17  & ~n42515;
  assign n27243 = ~n42516 & ~n42517;
  assign n27244 = ~n27231 & ~n27243;
  assign n27245 = n27231 & n27243;
  assign n27246 = ~n27231 & ~n27244;
  assign n27247 = ~n27243 & ~n27244;
  assign n27248 = ~n27246 & ~n27247;
  assign n27249 = ~n27244 & ~n27245;
  assign n27250 = n27230 & ~n42518;
  assign n27251 = ~n27230 & n42518;
  assign n27252 = ~n27250 & ~n27251;
  assign n27253 = ~n26436 & ~n26817;
  assign n27254 = ~n26436 & ~n42440;
  assign n27255 = ~n26437 & ~n27253;
  assign n27256 = n27252 & ~n42519;
  assign n27257 = ~n27252 & n42519;
  assign n27258 = ~n42519 & ~n27256;
  assign n27259 = n27252 & ~n27256;
  assign n27260 = ~n27258 & ~n27259;
  assign n27261 = ~n27256 & ~n27257;
  assign n27262 = ~n26835 & ~n42520;
  assign n27263 = n26835 & ~n27259;
  assign n27264 = ~n27258 & n27263;
  assign n27265 = n26835 & n42520;
  assign po80  = ~n27262 & ~n42521;
  assign n27267 = ~n27256 & ~n27262;
  assign n27268 = ~n27244 & ~n27250;
  assign n27269 = ~n26853 & ~n27229;
  assign n27270 = n6785 & n40885;
  assign n27271 = pi125  & n38631;
  assign n27272 = pi127  & n6800;
  assign n27273 = pi126  & n6802;
  assign n27274 = ~n27272 & ~n27273;
  assign n27275 = ~n27271 & ~n27273;
  assign n27276 = ~n27272 & n27275;
  assign n27277 = ~n27271 & n27274;
  assign n27278 = ~n27270 & n42522;
  assign n27279 = pi20  & ~n27278;
  assign n27280 = pi20  & ~n27279;
  assign n27281 = pi20  & n27278;
  assign n27282 = ~n27278 & ~n27279;
  assign n27283 = ~pi20  & ~n27278;
  assign n27284 = ~n42523 & ~n42524;
  assign n27285 = ~n27269 & ~n27284;
  assign n27286 = n27269 & n27284;
  assign n27287 = ~n27269 & ~n27285;
  assign n27288 = ~n27269 & n27284;
  assign n27289 = ~n27284 & ~n27285;
  assign n27290 = n27269 & ~n27284;
  assign n27291 = ~n42525 & ~n42526;
  assign n27292 = ~n27285 & ~n27286;
  assign n27293 = n5576 & n15111;
  assign n27294 = pi122  & n38406;
  assign n27295 = pi124  & n5591;
  assign n27296 = pi123  & n5593;
  assign n27297 = ~n27295 & ~n27296;
  assign n27298 = ~n27294 & ~n27296;
  assign n27299 = ~n27295 & n27298;
  assign n27300 = ~n27294 & n27297;
  assign n27301 = ~n27293 & n42528;
  assign n27302 = pi23  & ~n27301;
  assign n27303 = pi23  & ~n27302;
  assign n27304 = pi23  & n27301;
  assign n27305 = ~n27301 & ~n27302;
  assign n27306 = ~pi23  & ~n27301;
  assign n27307 = ~n42529 & ~n42530;
  assign n27308 = ~n27208 & ~n42511;
  assign n27309 = n27307 & n27308;
  assign n27310 = ~n27307 & ~n27308;
  assign n27311 = ~n27309 & ~n27310;
  assign n27312 = n4492 & n15091;
  assign n27313 = pi119  & n38208;
  assign n27314 = pi121  & n4507;
  assign n27315 = pi120  & n4509;
  assign n27316 = ~n27314 & ~n27315;
  assign n27317 = ~n27313 & ~n27315;
  assign n27318 = ~n27314 & n27317;
  assign n27319 = ~n27313 & n27316;
  assign n27320 = ~n27312 & n42531;
  assign n27321 = pi26  & ~n27320;
  assign n27322 = pi26  & ~n27321;
  assign n27323 = pi26  & n27320;
  assign n27324 = ~n27320 & ~n27321;
  assign n27325 = ~pi26  & ~n27320;
  assign n27326 = ~n42532 & ~n42533;
  assign n27327 = ~n26872 & ~n27189;
  assign n27328 = ~n27326 & ~n27327;
  assign n27329 = n27326 & n27327;
  assign n27330 = ~n27328 & ~n27329;
  assign n27331 = n607 & n13057;
  assign n27332 = pi116  & n37489;
  assign n27333 = pi118  & n620;
  assign n27334 = pi117  & n622;
  assign n27335 = ~n27333 & ~n27334;
  assign n27336 = ~n27332 & ~n27334;
  assign n27337 = ~n27333 & n27336;
  assign n27338 = ~n27332 & n27335;
  assign n27339 = ~n27331 & n42534;
  assign n27340 = pi29  & ~n27339;
  assign n27341 = pi29  & ~n27340;
  assign n27342 = pi29  & n27339;
  assign n27343 = ~n27339 & ~n27340;
  assign n27344 = ~pi29  & ~n27339;
  assign n27345 = ~n42535 & ~n42536;
  assign n27346 = ~n27171 & ~n42502;
  assign n27347 = n27345 & n27346;
  assign n27348 = ~n27345 & ~n27346;
  assign n27349 = ~n27347 & ~n27348;
  assign n27350 = ~n27119 & ~n27122;
  assign n27351 = ~n27113 & ~n27116;
  assign n27352 = n733 & n8209;
  assign n27353 = pi104  & n37510;
  assign n27354 = pi106  & n746;
  assign n27355 = pi105  & n748;
  assign n27356 = ~n27354 & ~n27355;
  assign n27357 = ~n27353 & ~n27355;
  assign n27358 = ~n27354 & n27357;
  assign n27359 = ~n27353 & n27356;
  assign n27360 = ~n27352 & n42537;
  assign n27361 = pi41  & ~n27360;
  assign n27362 = pi41  & ~n27361;
  assign n27363 = pi41  & n27360;
  assign n27364 = ~n27360 & ~n27361;
  assign n27365 = ~pi41  & ~n27360;
  assign n27366 = ~n42538 & ~n42539;
  assign n27367 = ~n27101 & ~n27107;
  assign n27368 = n785 & n6474;
  assign n27369 = pi98  & n37520;
  assign n27370 = pi100  & n787;
  assign n27371 = pi99  & n795;
  assign n27372 = ~n27370 & ~n27371;
  assign n27373 = ~n27369 & ~n27371;
  assign n27374 = ~n27370 & n27373;
  assign n27375 = ~n27369 & n27372;
  assign n27376 = ~n27368 & n42540;
  assign n27377 = pi47  & ~n27376;
  assign n27378 = pi47  & ~n27377;
  assign n27379 = pi47  & n27376;
  assign n27380 = ~n27376 & ~n27377;
  assign n27381 = ~pi47  & ~n27376;
  assign n27382 = ~n42541 & ~n42542;
  assign n27383 = ~n27032 & ~n27035;
  assign n27384 = ~n27009 & ~n27027;
  assign n27385 = n3354 & n7882;
  assign n27386 = pi86  & n39128;
  assign n27387 = pi88  & n7884;
  assign n27388 = pi87  & n7892;
  assign n27389 = ~n27387 & ~n27388;
  assign n27390 = ~n27386 & ~n27388;
  assign n27391 = ~n27387 & n27390;
  assign n27392 = ~n27386 & n27389;
  assign n27393 = ~n27385 & n42543;
  assign n27394 = pi59  & ~n27393;
  assign n27395 = pi59  & ~n27394;
  assign n27396 = pi59  & n27393;
  assign n27397 = ~n27393 & ~n27394;
  assign n27398 = ~pi59  & ~n27393;
  assign n27399 = ~n42544 & ~n42545;
  assign n27400 = n2804 & n12674;
  assign n27401 = pi83  & n40107;
  assign n27402 = pi85  & n12676;
  assign n27403 = pi84  & n12684;
  assign n27404 = ~n27402 & ~n27403;
  assign n27405 = ~n27401 & ~n27403;
  assign n27406 = ~n27402 & n27405;
  assign n27407 = ~n27401 & n27404;
  assign n27408 = ~n27400 & n42546;
  assign n27409 = pi62  & ~n27408;
  assign n27410 = pi62  & ~n27409;
  assign n27411 = pi62  & n27408;
  assign n27412 = ~n27408 & ~n27409;
  assign n27413 = ~pi62  & ~n27408;
  assign n27414 = ~n42547 & ~n42548;
  assign n27415 = pi82  & ~n40814;
  assign n27416 = pi81  & n18285;
  assign n27417 = ~n27415 & ~n27416;
  assign n27418 = ~pi17  & ~n27417;
  assign n27419 = pi17  & n27417;
  assign n27420 = ~n27418 & ~n27419;
  assign n27421 = ~n26995 & n27420;
  assign n27422 = n26995 & ~n27420;
  assign n27423 = ~n27421 & ~n27422;
  assign n27424 = ~n27414 & n27423;
  assign n27425 = n27414 & ~n27423;
  assign n27426 = ~n27414 & ~n27424;
  assign n27427 = ~n27414 & ~n27423;
  assign n27428 = n27423 & ~n27424;
  assign n27429 = n27414 & n27423;
  assign n27430 = ~n42549 & ~n42550;
  assign n27431 = ~n27424 & ~n27425;
  assign n27432 = ~n27004 & ~n42551;
  assign n27433 = n27004 & n42551;
  assign n27434 = ~n27004 & ~n27432;
  assign n27435 = ~n42551 & ~n27432;
  assign n27436 = ~n27434 & ~n27435;
  assign n27437 = ~n27432 & ~n27433;
  assign n27438 = n27399 & n42552;
  assign n27439 = ~n27399 & ~n42552;
  assign n27440 = ~n27438 & ~n27439;
  assign n27441 = ~n27384 & n27440;
  assign n27442 = n27384 & ~n27440;
  assign n27443 = ~n27441 & ~n27442;
  assign n27444 = n594 & n4312;
  assign n27445 = pi89  & n38376;
  assign n27446 = pi91  & n4314;
  assign n27447 = pi90  & n4322;
  assign n27448 = ~n27446 & ~n27447;
  assign n27449 = ~n27445 & ~n27447;
  assign n27450 = ~n27446 & n27449;
  assign n27451 = ~n27445 & n27448;
  assign n27452 = ~n27444 & n42553;
  assign n27453 = pi56  & ~n27452;
  assign n27454 = pi56  & ~n27453;
  assign n27455 = pi56  & n27452;
  assign n27456 = ~n27452 & ~n27453;
  assign n27457 = ~pi56  & ~n27452;
  assign n27458 = ~n42554 & ~n42555;
  assign n27459 = n27443 & ~n27458;
  assign n27460 = ~n27443 & n27458;
  assign n27461 = n27443 & ~n27459;
  assign n27462 = n27443 & n27458;
  assign n27463 = ~n27458 & ~n27459;
  assign n27464 = ~n27443 & ~n27458;
  assign n27465 = ~n42556 & ~n42557;
  assign n27466 = ~n27459 & ~n27460;
  assign n27467 = n27383 & n42558;
  assign n27468 = ~n27383 & ~n42558;
  assign n27469 = ~n27467 & ~n27468;
  assign n27470 = n1971 & n4524;
  assign n27471 = pi92  & n37864;
  assign n27472 = pi94  & n1973;
  assign n27473 = pi93  & n1981;
  assign n27474 = ~n27472 & ~n27473;
  assign n27475 = ~n27471 & ~n27473;
  assign n27476 = ~n27472 & n27475;
  assign n27477 = ~n27471 & n27474;
  assign n27478 = ~n27470 & n42559;
  assign n27479 = pi53  & ~n27478;
  assign n27480 = pi53  & ~n27479;
  assign n27481 = pi53  & n27478;
  assign n27482 = ~n27478 & ~n27479;
  assign n27483 = ~pi53  & ~n27478;
  assign n27484 = ~n42560 & ~n42561;
  assign n27485 = n27469 & ~n27484;
  assign n27486 = ~n27469 & n27484;
  assign n27487 = n27469 & ~n27485;
  assign n27488 = n27469 & n27484;
  assign n27489 = ~n27484 & ~n27485;
  assign n27490 = ~n27469 & ~n27484;
  assign n27491 = ~n42562 & ~n42563;
  assign n27492 = ~n27485 & ~n27486;
  assign n27493 = ~n27041 & n27058;
  assign n27494 = ~n27041 & ~n27059;
  assign n27495 = ~n27042 & ~n27493;
  assign n27496 = n42564 & n42565;
  assign n27497 = ~n42564 & ~n42565;
  assign n27498 = ~n27496 & ~n27497;
  assign n27499 = n894 & n5630;
  assign n27500 = pi95  & n37580;
  assign n27501 = pi97  & n896;
  assign n27502 = pi96  & n904;
  assign n27503 = ~n27501 & ~n27502;
  assign n27504 = ~n27500 & ~n27502;
  assign n27505 = ~n27501 & n27504;
  assign n27506 = ~n27500 & n27503;
  assign n27507 = ~n27499 & n42566;
  assign n27508 = pi50  & ~n27507;
  assign n27509 = pi50  & ~n27508;
  assign n27510 = pi50  & n27507;
  assign n27511 = ~n27507 & ~n27508;
  assign n27512 = ~pi50  & ~n27507;
  assign n27513 = ~n42567 & ~n42568;
  assign n27514 = n26960 & ~n27065;
  assign n27515 = ~n27065 & ~n27073;
  assign n27516 = ~n27066 & ~n27514;
  assign n27517 = ~n27513 & ~n42569;
  assign n27518 = n27513 & n42569;
  assign n27519 = ~n27517 & ~n27518;
  assign n27520 = n27498 & n27519;
  assign n27521 = ~n27498 & ~n27519;
  assign n27522 = ~n27498 & n27519;
  assign n27523 = n27498 & ~n27519;
  assign n27524 = ~n27522 & ~n27523;
  assign n27525 = ~n27520 & ~n27521;
  assign n27526 = ~n27382 & ~n42570;
  assign n27527 = n27382 & n42570;
  assign n27528 = ~n27526 & ~n27527;
  assign n27529 = ~n27078 & n27094;
  assign n27530 = ~n27078 & ~n27095;
  assign n27531 = ~n27077 & ~n27529;
  assign n27532 = ~n27528 & n42571;
  assign n27533 = n27528 & ~n42571;
  assign n27534 = ~n27532 & ~n27533;
  assign n27535 = n940 & n6787;
  assign n27536 = pi101  & n37541;
  assign n27537 = pi103  & n953;
  assign n27538 = pi102  & n955;
  assign n27539 = ~n27537 & ~n27538;
  assign n27540 = ~n27536 & ~n27538;
  assign n27541 = ~n27537 & n27540;
  assign n27542 = ~n27536 & n27539;
  assign n27543 = ~n27535 & n42572;
  assign n27544 = pi44  & ~n27543;
  assign n27545 = pi44  & ~n27544;
  assign n27546 = pi44  & n27543;
  assign n27547 = ~n27543 & ~n27544;
  assign n27548 = ~pi44  & ~n27543;
  assign n27549 = ~n42573 & ~n42574;
  assign n27550 = n27534 & ~n27549;
  assign n27551 = ~n27534 & n27549;
  assign n27552 = n27534 & ~n27550;
  assign n27553 = n27534 & n27549;
  assign n27554 = ~n27549 & ~n27550;
  assign n27555 = ~n27534 & ~n27549;
  assign n27556 = ~n42575 & ~n42576;
  assign n27557 = ~n27550 & ~n27551;
  assign n27558 = ~n27367 & ~n42577;
  assign n27559 = n27367 & n42577;
  assign n27560 = ~n27367 & n42577;
  assign n27561 = n27367 & ~n42577;
  assign n27562 = ~n27560 & ~n27561;
  assign n27563 = ~n27558 & ~n27559;
  assign n27564 = ~n27366 & ~n42578;
  assign n27565 = n27366 & n42578;
  assign n27566 = ~n27564 & ~n27565;
  assign n27567 = n27351 & ~n27566;
  assign n27568 = ~n27351 & n27566;
  assign n27569 = ~n27567 & ~n27568;
  assign n27570 = n691 & n9701;
  assign n27571 = pi107  & n37503;
  assign n27572 = pi109  & n704;
  assign n27573 = pi108  & n706;
  assign n27574 = ~n27572 & ~n27573;
  assign n27575 = ~n27571 & ~n27573;
  assign n27576 = ~n27572 & n27575;
  assign n27577 = ~n27571 & n27574;
  assign n27578 = ~n27570 & n42579;
  assign n27579 = pi38  & ~n27578;
  assign n27580 = pi38  & ~n27579;
  assign n27581 = pi38  & n27578;
  assign n27582 = ~n27578 & ~n27579;
  assign n27583 = ~pi38  & ~n27578;
  assign n27584 = ~n42580 & ~n42581;
  assign n27585 = n27569 & ~n27584;
  assign n27586 = ~n27569 & n27584;
  assign n27587 = n27569 & ~n27585;
  assign n27588 = n27569 & n27584;
  assign n27589 = ~n27584 & ~n27585;
  assign n27590 = ~n27569 & ~n27584;
  assign n27591 = ~n42582 & ~n42583;
  assign n27592 = ~n27585 & ~n27586;
  assign n27593 = n27350 & n42584;
  assign n27594 = ~n27350 & ~n42584;
  assign n27595 = ~n27593 & ~n27594;
  assign n27596 = n2104 & n10844;
  assign n27597 = pi110  & n37758;
  assign n27598 = pi112  & n2117;
  assign n27599 = pi111  & n2119;
  assign n27600 = ~n27598 & ~n27599;
  assign n27601 = ~n27597 & ~n27599;
  assign n27602 = ~n27598 & n27601;
  assign n27603 = ~n27597 & n27600;
  assign n27604 = ~n27596 & n42585;
  assign n27605 = pi35  & ~n27604;
  assign n27606 = pi35  & ~n27605;
  assign n27607 = pi35  & n27604;
  assign n27608 = ~n27604 & ~n27605;
  assign n27609 = ~pi35  & ~n27604;
  assign n27610 = ~n42586 & ~n42587;
  assign n27611 = n27595 & ~n27610;
  assign n27612 = ~n27595 & n27610;
  assign n27613 = n27595 & ~n27611;
  assign n27614 = n27595 & n27610;
  assign n27615 = ~n27610 & ~n27611;
  assign n27616 = ~n27595 & ~n27610;
  assign n27617 = ~n42588 & ~n42589;
  assign n27618 = ~n27611 & ~n27612;
  assign n27619 = ~n27128 & n27145;
  assign n27620 = ~n27128 & ~n27146;
  assign n27621 = ~n27129 & ~n27619;
  assign n27622 = n42590 & n42591;
  assign n27623 = ~n42590 & ~n42591;
  assign n27624 = ~n27622 & ~n27623;
  assign n27625 = n523 & n649;
  assign n27626 = pi113  & n37496;
  assign n27627 = pi115  & n662;
  assign n27628 = pi114  & n664;
  assign n27629 = ~n27627 & ~n27628;
  assign n27630 = ~n27626 & ~n27628;
  assign n27631 = ~n27627 & n27630;
  assign n27632 = ~n27626 & n27629;
  assign n27633 = ~n27625 & n42592;
  assign n27634 = pi32  & ~n27633;
  assign n27635 = pi32  & ~n27634;
  assign n27636 = pi32  & n27633;
  assign n27637 = ~n27633 & ~n27634;
  assign n27638 = ~pi32  & ~n27633;
  assign n27639 = ~n42593 & ~n42594;
  assign n27640 = ~n26893 & ~n27152;
  assign n27641 = ~n27639 & ~n27640;
  assign n27642 = n27639 & n27640;
  assign n27643 = ~n27641 & ~n27642;
  assign n27644 = n27624 & n27643;
  assign n27645 = ~n27624 & ~n27643;
  assign n27646 = n27624 & ~n27644;
  assign n27647 = n27643 & ~n27644;
  assign n27648 = ~n27646 & ~n27647;
  assign n27649 = ~n27644 & ~n27645;
  assign n27650 = n27349 & ~n42595;
  assign n27651 = n27349 & ~n27650;
  assign n27652 = n27349 & n42595;
  assign n27653 = ~n42595 & ~n27650;
  assign n27654 = ~n27349 & ~n42595;
  assign n27655 = ~n27349 & n42595;
  assign n27656 = ~n27650 & ~n27655;
  assign n27657 = ~n42596 & ~n42597;
  assign n27658 = n27330 & n42598;
  assign n27659 = ~n27330 & ~n42598;
  assign n27660 = n42598 & ~n27658;
  assign n27661 = ~n27330 & n42598;
  assign n27662 = n27330 & ~n27658;
  assign n27663 = n27330 & ~n42598;
  assign n27664 = ~n42599 & ~n42600;
  assign n27665 = ~n27658 & ~n27659;
  assign n27666 = n27311 & ~n42601;
  assign n27667 = ~n27311 & n42601;
  assign n27668 = n27311 & ~n27666;
  assign n27669 = ~n42601 & ~n27666;
  assign n27670 = ~n27668 & ~n27669;
  assign n27671 = ~n27666 & ~n27667;
  assign n27672 = ~n42527 & ~n42602;
  assign n27673 = n42527 & n42602;
  assign n27674 = ~n42527 & n42602;
  assign n27675 = n42527 & ~n42602;
  assign n27676 = ~n27674 & ~n27675;
  assign n27677 = ~n27672 & ~n27673;
  assign n27678 = ~n27268 & ~n42603;
  assign n27679 = n27268 & n42603;
  assign n27680 = ~n27268 & ~n27678;
  assign n27681 = ~n42603 & ~n27678;
  assign n27682 = ~n27680 & ~n27681;
  assign n27683 = ~n27678 & ~n27679;
  assign n27684 = ~n27267 & ~n42604;
  assign n27685 = n27267 & ~n27681;
  assign n27686 = ~n27680 & n27685;
  assign n27687 = n27267 & n42604;
  assign po81  = ~n27684 & ~n42605;
  assign n27689 = ~n27678 & ~n27684;
  assign n27690 = ~n27285 & ~n27672;
  assign n27691 = n6785 & n40891;
  assign n27692 = pi126  & n38631;
  assign n27693 = pi127  & n6802;
  assign n27694 = ~n27692 & ~n27693;
  assign n27695 = ~n6785 & n27694;
  assign n27696 = ~n40891 & n27694;
  assign n27697 = ~n27695 & ~n27696;
  assign n27698 = ~n27691 & n27694;
  assign n27699 = pi20  & ~n42606;
  assign n27700 = ~pi20  & n42606;
  assign n27701 = ~n27699 & ~n27700;
  assign n27702 = ~n27310 & n42601;
  assign n27703 = ~n27310 & ~n27666;
  assign n27704 = ~n27309 & ~n27702;
  assign n27705 = ~n27701 & ~n42607;
  assign n27706 = n27701 & n42607;
  assign n27707 = ~n42607 & ~n27705;
  assign n27708 = n27701 & ~n42607;
  assign n27709 = ~n27701 & ~n27705;
  assign n27710 = ~n27701 & n42607;
  assign n27711 = ~n42608 & ~n42609;
  assign n27712 = ~n27705 & ~n27706;
  assign n27713 = n5576 & n15068;
  assign n27714 = pi123  & n38406;
  assign n27715 = pi125  & n5591;
  assign n27716 = pi124  & n5593;
  assign n27717 = ~n27715 & ~n27716;
  assign n27718 = ~n27714 & ~n27716;
  assign n27719 = ~n27715 & n27718;
  assign n27720 = ~n27714 & n27717;
  assign n27721 = ~n27713 & n42611;
  assign n27722 = pi23  & ~n27721;
  assign n27723 = pi23  & ~n27722;
  assign n27724 = pi23  & n27721;
  assign n27725 = ~n27721 & ~n27722;
  assign n27726 = ~pi23  & ~n27721;
  assign n27727 = ~n42612 & ~n42613;
  assign n27728 = ~n27328 & ~n42598;
  assign n27729 = ~n27328 & ~n27658;
  assign n27730 = ~n27329 & ~n27728;
  assign n27731 = n27727 & n42614;
  assign n27732 = ~n27727 & ~n42614;
  assign n27733 = ~n27731 & ~n27732;
  assign n27734 = n4492 & n15049;
  assign n27735 = pi120  & n38208;
  assign n27736 = pi122  & n4507;
  assign n27737 = pi121  & n4509;
  assign n27738 = ~n27736 & ~n27737;
  assign n27739 = ~n27735 & ~n27737;
  assign n27740 = ~n27736 & n27739;
  assign n27741 = ~n27735 & n27738;
  assign n27742 = ~n27734 & n42615;
  assign n27743 = pi26  & ~n27742;
  assign n27744 = pi26  & ~n27743;
  assign n27745 = pi26  & n27742;
  assign n27746 = ~n27742 & ~n27743;
  assign n27747 = ~pi26  & ~n27742;
  assign n27748 = ~n42616 & ~n42617;
  assign n27749 = ~n27348 & n42595;
  assign n27750 = ~n27348 & ~n27650;
  assign n27751 = ~n27347 & ~n27749;
  assign n27752 = n27748 & n42618;
  assign n27753 = ~n27748 & ~n42618;
  assign n27754 = ~n27752 & ~n27753;
  assign n27755 = n607 & n13027;
  assign n27756 = pi117  & n37489;
  assign n27757 = pi119  & n620;
  assign n27758 = pi118  & n622;
  assign n27759 = ~n27757 & ~n27758;
  assign n27760 = ~n27756 & ~n27758;
  assign n27761 = ~n27757 & n27760;
  assign n27762 = ~n27756 & n27759;
  assign n27763 = ~n27755 & n42619;
  assign n27764 = pi29  & ~n27763;
  assign n27765 = pi29  & ~n27764;
  assign n27766 = pi29  & n27763;
  assign n27767 = ~n27763 & ~n27764;
  assign n27768 = ~pi29  & ~n27763;
  assign n27769 = ~n42620 & ~n42621;
  assign n27770 = n27624 & ~n27642;
  assign n27771 = ~n27641 & ~n27644;
  assign n27772 = ~n27641 & ~n27770;
  assign n27773 = n27769 & n42622;
  assign n27774 = ~n27769 & ~n42622;
  assign n27775 = ~n27773 & ~n27774;
  assign n27776 = n649 & n12530;
  assign n27777 = pi114  & n37496;
  assign n27778 = pi116  & n662;
  assign n27779 = pi115  & n664;
  assign n27780 = ~n27778 & ~n27779;
  assign n27781 = ~n27777 & ~n27779;
  assign n27782 = ~n27778 & n27781;
  assign n27783 = ~n27777 & n27780;
  assign n27784 = ~n27776 & n42623;
  assign n27785 = pi32  & ~n27784;
  assign n27786 = pi32  & ~n27785;
  assign n27787 = pi32  & n27784;
  assign n27788 = ~n27784 & ~n27785;
  assign n27789 = ~pi32  & ~n27784;
  assign n27790 = ~n42624 & ~n42625;
  assign n27791 = ~n27611 & ~n27623;
  assign n27792 = n27790 & n27791;
  assign n27793 = ~n27790 & ~n27791;
  assign n27794 = ~n27792 & ~n27793;
  assign n27795 = ~n27585 & ~n27594;
  assign n27796 = ~n27564 & ~n27568;
  assign n27797 = ~n27550 & ~n27558;
  assign n27798 = n940 & n8136;
  assign n27799 = pi102  & n37541;
  assign n27800 = pi104  & n953;
  assign n27801 = pi103  & n955;
  assign n27802 = ~n27800 & ~n27801;
  assign n27803 = ~n27799 & ~n27801;
  assign n27804 = ~n27800 & n27803;
  assign n27805 = ~n27799 & n27802;
  assign n27806 = ~n27798 & n42626;
  assign n27807 = pi44  & ~n27806;
  assign n27808 = pi44  & ~n27807;
  assign n27809 = pi44  & n27806;
  assign n27810 = ~n27806 & ~n27807;
  assign n27811 = ~pi44  & ~n27806;
  assign n27812 = ~n42627 & ~n42628;
  assign n27813 = ~n27526 & ~n27533;
  assign n27814 = ~n27485 & ~n27497;
  assign n27815 = n4312 & n4453;
  assign n27816 = pi90  & n38376;
  assign n27817 = pi92  & n4314;
  assign n27818 = pi91  & n4322;
  assign n27819 = ~n27817 & ~n27818;
  assign n27820 = ~n27816 & ~n27818;
  assign n27821 = ~n27817 & n27820;
  assign n27822 = ~n27816 & n27819;
  assign n27823 = ~n27815 & n42629;
  assign n27824 = pi56  & ~n27823;
  assign n27825 = pi56  & ~n27824;
  assign n27826 = pi56  & n27823;
  assign n27827 = ~n27823 & ~n27824;
  assign n27828 = ~pi56  & ~n27823;
  assign n27829 = ~n42630 & ~n42631;
  assign n27830 = ~n27439 & ~n27441;
  assign n27831 = ~n27418 & ~n27421;
  assign n27832 = pi83  & ~n40814;
  assign n27833 = pi82  & n18285;
  assign n27834 = ~n27832 & ~n27833;
  assign n27835 = n27831 & ~n27834;
  assign n27836 = ~n27831 & n27834;
  assign n27837 = ~n27835 & ~n27836;
  assign n27838 = n2779 & n12674;
  assign n27839 = pi84  & n40107;
  assign n27840 = pi86  & n12676;
  assign n27841 = pi85  & n12684;
  assign n27842 = ~n27840 & ~n27841;
  assign n27843 = ~n27839 & ~n27841;
  assign n27844 = ~n27840 & n27843;
  assign n27845 = ~n27839 & n27842;
  assign n27846 = ~n27838 & n42632;
  assign n27847 = pi62  & ~n27846;
  assign n27848 = pi62  & ~n27847;
  assign n27849 = pi62  & n27846;
  assign n27850 = ~n27846 & ~n27847;
  assign n27851 = ~pi62  & ~n27846;
  assign n27852 = ~n42633 & ~n42634;
  assign n27853 = ~n27837 & n27852;
  assign n27854 = n27837 & ~n27852;
  assign n27855 = ~n27853 & ~n27854;
  assign n27856 = ~n27424 & ~n27432;
  assign n27857 = n27855 & ~n27856;
  assign n27858 = ~n27855 & n27856;
  assign n27859 = ~n27857 & ~n27858;
  assign n27860 = n3591 & n7882;
  assign n27861 = pi87  & n39128;
  assign n27862 = pi89  & n7884;
  assign n27863 = pi88  & n7892;
  assign n27864 = ~n27862 & ~n27863;
  assign n27865 = ~n27861 & ~n27863;
  assign n27866 = ~n27862 & n27865;
  assign n27867 = ~n27861 & n27864;
  assign n27868 = ~n27860 & n42635;
  assign n27869 = pi59  & ~n27868;
  assign n27870 = pi59  & ~n27869;
  assign n27871 = pi59  & n27868;
  assign n27872 = ~n27868 & ~n27869;
  assign n27873 = ~pi59  & ~n27868;
  assign n27874 = ~n42636 & ~n42637;
  assign n27875 = ~n27859 & n27874;
  assign n27876 = n27859 & ~n27874;
  assign n27877 = n27859 & ~n27876;
  assign n27878 = ~n27874 & ~n27876;
  assign n27879 = ~n27877 & ~n27878;
  assign n27880 = ~n27875 & ~n27876;
  assign n27881 = ~n27830 & ~n42638;
  assign n27882 = n27830 & n42638;
  assign n27883 = ~n27830 & n42638;
  assign n27884 = n27830 & ~n42638;
  assign n27885 = ~n27883 & ~n27884;
  assign n27886 = ~n27881 & ~n27882;
  assign n27887 = n27829 & n42639;
  assign n27888 = ~n27829 & ~n42639;
  assign n27889 = ~n27887 & ~n27888;
  assign n27890 = ~n27459 & ~n27468;
  assign n27891 = n27889 & ~n27890;
  assign n27892 = ~n27889 & n27890;
  assign n27893 = ~n27891 & ~n27892;
  assign n27894 = n1971 & n4494;
  assign n27895 = pi93  & n37864;
  assign n27896 = pi95  & n1973;
  assign n27897 = pi94  & n1981;
  assign n27898 = ~n27896 & ~n27897;
  assign n27899 = ~n27895 & ~n27897;
  assign n27900 = ~n27896 & n27899;
  assign n27901 = ~n27895 & n27898;
  assign n27902 = ~n27894 & n42640;
  assign n27903 = pi53  & ~n27902;
  assign n27904 = pi53  & ~n27903;
  assign n27905 = pi53  & n27902;
  assign n27906 = ~n27902 & ~n27903;
  assign n27907 = ~pi53  & ~n27902;
  assign n27908 = ~n42641 & ~n42642;
  assign n27909 = ~n27893 & n27908;
  assign n27910 = n27893 & ~n27908;
  assign n27911 = n27893 & ~n27910;
  assign n27912 = ~n27908 & ~n27910;
  assign n27913 = ~n27911 & ~n27912;
  assign n27914 = ~n27909 & ~n27910;
  assign n27915 = n27814 & n42643;
  assign n27916 = ~n27814 & ~n42643;
  assign n27917 = ~n27915 & ~n27916;
  assign n27918 = n894 & n5610;
  assign n27919 = pi96  & n37580;
  assign n27920 = pi98  & n896;
  assign n27921 = pi97  & n904;
  assign n27922 = ~n27920 & ~n27921;
  assign n27923 = ~n27919 & ~n27921;
  assign n27924 = ~n27920 & n27923;
  assign n27925 = ~n27919 & n27922;
  assign n27926 = ~n27918 & n42644;
  assign n27927 = pi50  & ~n27926;
  assign n27928 = pi50  & ~n27927;
  assign n27929 = pi50  & n27926;
  assign n27930 = ~n27926 & ~n27927;
  assign n27931 = ~pi50  & ~n27926;
  assign n27932 = ~n42645 & ~n42646;
  assign n27933 = n27917 & ~n27932;
  assign n27934 = ~n27917 & n27932;
  assign n27935 = n27917 & ~n27933;
  assign n27936 = ~n27932 & ~n27933;
  assign n27937 = ~n27935 & ~n27936;
  assign n27938 = ~n27933 & ~n27934;
  assign n27939 = ~n27498 & ~n27517;
  assign n27940 = ~n27517 & ~n27520;
  assign n27941 = ~n27518 & ~n27939;
  assign n27942 = n42647 & n42648;
  assign n27943 = ~n42647 & ~n42648;
  assign n27944 = ~n27942 & ~n27943;
  assign n27945 = n785 & n6839;
  assign n27946 = pi99  & n37520;
  assign n27947 = pi101  & n787;
  assign n27948 = pi100  & n795;
  assign n27949 = ~n27947 & ~n27948;
  assign n27950 = ~n27946 & ~n27948;
  assign n27951 = ~n27947 & n27950;
  assign n27952 = ~n27946 & n27949;
  assign n27953 = ~n27945 & n42649;
  assign n27954 = pi47  & ~n27953;
  assign n27955 = pi47  & ~n27954;
  assign n27956 = pi47  & n27953;
  assign n27957 = ~n27953 & ~n27954;
  assign n27958 = ~pi47  & ~n27953;
  assign n27959 = ~n42650 & ~n42651;
  assign n27960 = ~n27944 & n27959;
  assign n27961 = n27944 & ~n27959;
  assign n27962 = ~n27960 & ~n27961;
  assign n27963 = ~n27813 & n27962;
  assign n27964 = n27813 & ~n27962;
  assign n27965 = ~n27813 & ~n27963;
  assign n27966 = n27962 & ~n27963;
  assign n27967 = ~n27965 & ~n27966;
  assign n27968 = ~n27963 & ~n27964;
  assign n27969 = ~n27812 & ~n42652;
  assign n27970 = n27812 & ~n27966;
  assign n27971 = ~n27965 & n27970;
  assign n27972 = n27812 & n42652;
  assign n27973 = ~n27969 & ~n42653;
  assign n27974 = ~n27797 & n27973;
  assign n27975 = n27797 & ~n27973;
  assign n27976 = ~n27974 & ~n27975;
  assign n27977 = n733 & n8177;
  assign n27978 = pi105  & n37510;
  assign n27979 = pi107  & n746;
  assign n27980 = pi106  & n748;
  assign n27981 = ~n27979 & ~n27980;
  assign n27982 = ~n27978 & ~n27980;
  assign n27983 = ~n27979 & n27982;
  assign n27984 = ~n27978 & n27981;
  assign n27985 = ~n27977 & n42654;
  assign n27986 = pi41  & ~n27985;
  assign n27987 = pi41  & ~n27986;
  assign n27988 = pi41  & n27985;
  assign n27989 = ~n27985 & ~n27986;
  assign n27990 = ~pi41  & ~n27985;
  assign n27991 = ~n42655 & ~n42656;
  assign n27992 = n27976 & ~n27991;
  assign n27993 = ~n27976 & n27991;
  assign n27994 = n27976 & ~n27992;
  assign n27995 = ~n27991 & ~n27992;
  assign n27996 = ~n27994 & ~n27995;
  assign n27997 = ~n27992 & ~n27993;
  assign n27998 = n27796 & n42657;
  assign n27999 = ~n27796 & ~n42657;
  assign n28000 = ~n27998 & ~n27999;
  assign n28001 = n691 & n9678;
  assign n28002 = pi108  & n37503;
  assign n28003 = pi110  & n704;
  assign n28004 = pi109  & n706;
  assign n28005 = ~n28003 & ~n28004;
  assign n28006 = ~n28002 & ~n28004;
  assign n28007 = ~n28003 & n28006;
  assign n28008 = ~n28002 & n28005;
  assign n28009 = ~n28001 & n42658;
  assign n28010 = pi38  & ~n28009;
  assign n28011 = pi38  & ~n28010;
  assign n28012 = pi38  & n28009;
  assign n28013 = ~n28009 & ~n28010;
  assign n28014 = ~pi38  & ~n28009;
  assign n28015 = ~n42659 & ~n42660;
  assign n28016 = ~n28000 & n28015;
  assign n28017 = n28000 & ~n28015;
  assign n28018 = n28000 & ~n28017;
  assign n28019 = ~n28015 & ~n28017;
  assign n28020 = ~n28018 & ~n28019;
  assign n28021 = ~n28016 & ~n28017;
  assign n28022 = n27795 & n42661;
  assign n28023 = ~n27795 & ~n42661;
  assign n28024 = ~n28022 & ~n28023;
  assign n28025 = n2104 & n11276;
  assign n28026 = pi111  & n37758;
  assign n28027 = pi113  & n2117;
  assign n28028 = pi112  & n2119;
  assign n28029 = ~n28027 & ~n28028;
  assign n28030 = ~n28026 & ~n28028;
  assign n28031 = ~n28027 & n28030;
  assign n28032 = ~n28026 & n28029;
  assign n28033 = ~n28025 & n42662;
  assign n28034 = pi35  & ~n28033;
  assign n28035 = pi35  & ~n28034;
  assign n28036 = pi35  & n28033;
  assign n28037 = ~n28033 & ~n28034;
  assign n28038 = ~pi35  & ~n28033;
  assign n28039 = ~n42663 & ~n42664;
  assign n28040 = n28024 & ~n28039;
  assign n28041 = ~n28024 & n28039;
  assign n28042 = n28024 & ~n28040;
  assign n28043 = ~n28039 & ~n28040;
  assign n28044 = ~n28042 & ~n28043;
  assign n28045 = ~n28040 & ~n28041;
  assign n28046 = n27794 & ~n42665;
  assign n28047 = ~n27794 & n42665;
  assign n28048 = ~n28046 & ~n28047;
  assign n28049 = n27775 & ~n28047;
  assign n28050 = ~n28046 & n28049;
  assign n28051 = n27775 & n28048;
  assign n28052 = ~n27775 & ~n28048;
  assign n28053 = n27775 & ~n42666;
  assign n28054 = ~n28047 & ~n42666;
  assign n28055 = ~n28046 & n28054;
  assign n28056 = n28048 & ~n42666;
  assign n28057 = ~n28053 & ~n42667;
  assign n28058 = ~n42666 & ~n28052;
  assign n28059 = n27754 & ~n42668;
  assign n28060 = ~n27754 & n42668;
  assign n28061 = ~n28059 & ~n28060;
  assign n28062 = n27733 & ~n28060;
  assign n28063 = ~n28059 & n28062;
  assign n28064 = n27733 & n28061;
  assign n28065 = ~n27733 & ~n28061;
  assign n28066 = n27733 & ~n42669;
  assign n28067 = ~n28060 & ~n42669;
  assign n28068 = ~n28059 & n28067;
  assign n28069 = n28061 & ~n42669;
  assign n28070 = ~n28066 & ~n42670;
  assign n28071 = ~n42669 & ~n28065;
  assign n28072 = ~n42610 & ~n42671;
  assign n28073 = ~n42609 & n42671;
  assign n28074 = ~n42608 & n28073;
  assign n28075 = ~n42608 & n42671;
  assign n28076 = ~n42609 & n28075;
  assign n28077 = n42610 & n42671;
  assign n28078 = ~n28072 & ~n42672;
  assign n28079 = ~n27690 & n28078;
  assign n28080 = n27690 & ~n28078;
  assign n28081 = ~n27690 & ~n28079;
  assign n28082 = n28078 & ~n28079;
  assign n28083 = ~n28081 & ~n28082;
  assign n28084 = ~n28079 & ~n28080;
  assign n28085 = ~n27689 & ~n42673;
  assign n28086 = n27689 & ~n28082;
  assign n28087 = ~n28081 & n28086;
  assign n28088 = n27689 & n42673;
  assign po82  = ~n28085 & ~n42674;
  assign n28090 = ~n28079 & ~n28085;
  assign n28091 = ~n27705 & ~n28072;
  assign n28092 = n6785 & ~n18675;
  assign n28093 = ~n38631 & ~n28092;
  assign n28094 = pi127  & n38631;
  assign n28095 = n6785 & n18680;
  assign n28096 = ~n28094 & ~n28095;
  assign n28097 = pi127  & ~n28093;
  assign n28098 = pi20  & ~n42675;
  assign n28099 = pi20  & ~n28098;
  assign n28100 = pi20  & n42675;
  assign n28101 = ~n42675 & ~n28098;
  assign n28102 = ~pi20  & ~n42675;
  assign n28103 = ~n42676 & ~n42677;
  assign n28104 = ~n27732 & ~n28061;
  assign n28105 = ~n27732 & ~n42669;
  assign n28106 = ~n27731 & ~n28104;
  assign n28107 = ~n28103 & ~n42678;
  assign n28108 = n28103 & n42678;
  assign n28109 = ~n42678 & ~n28107;
  assign n28110 = ~n28103 & ~n28107;
  assign n28111 = ~n28109 & ~n28110;
  assign n28112 = ~n28107 & ~n28108;
  assign n28113 = n5576 & n15021;
  assign n28114 = pi124  & n38406;
  assign n28115 = pi126  & n5591;
  assign n28116 = pi125  & n5593;
  assign n28117 = ~n28115 & ~n28116;
  assign n28118 = ~n28114 & ~n28116;
  assign n28119 = ~n28115 & n28118;
  assign n28120 = ~n28114 & n28117;
  assign n28121 = ~n28113 & n42680;
  assign n28122 = pi23  & ~n28121;
  assign n28123 = pi23  & ~n28122;
  assign n28124 = pi23  & n28121;
  assign n28125 = ~n28121 & ~n28122;
  assign n28126 = ~pi23  & ~n28121;
  assign n28127 = ~n42681 & ~n42682;
  assign n28128 = ~n27753 & ~n28059;
  assign n28129 = ~n28127 & ~n28128;
  assign n28130 = n28127 & n28128;
  assign n28131 = ~n28127 & ~n28129;
  assign n28132 = ~n28127 & n28128;
  assign n28133 = ~n28128 & ~n28129;
  assign n28134 = n28127 & ~n28128;
  assign n28135 = ~n42683 & ~n42684;
  assign n28136 = ~n28129 & ~n28130;
  assign n28137 = n4492 & n14961;
  assign n28138 = pi121  & n38208;
  assign n28139 = pi123  & n4507;
  assign n28140 = pi122  & n4509;
  assign n28141 = ~n28139 & ~n28140;
  assign n28142 = ~n28138 & ~n28140;
  assign n28143 = ~n28139 & n28142;
  assign n28144 = ~n28138 & n28141;
  assign n28145 = ~n28137 & n42686;
  assign n28146 = pi26  & ~n28145;
  assign n28147 = pi26  & ~n28146;
  assign n28148 = pi26  & n28145;
  assign n28149 = ~n28145 & ~n28146;
  assign n28150 = ~pi26  & ~n28145;
  assign n28151 = ~n42687 & ~n42688;
  assign n28152 = ~n27774 & ~n42666;
  assign n28153 = n28151 & n28152;
  assign n28154 = ~n28151 & ~n28152;
  assign n28155 = ~n28153 & ~n28154;
  assign n28156 = n649 & n13079;
  assign n28157 = pi115  & n37496;
  assign n28158 = pi117  & n662;
  assign n28159 = pi116  & n664;
  assign n28160 = ~n28158 & ~n28159;
  assign n28161 = ~n28157 & ~n28159;
  assign n28162 = ~n28158 & n28161;
  assign n28163 = ~n28157 & n28160;
  assign n28164 = ~n28156 & n42689;
  assign n28165 = pi32  & ~n28164;
  assign n28166 = pi32  & ~n28165;
  assign n28167 = pi32  & n28164;
  assign n28168 = ~n28164 & ~n28165;
  assign n28169 = ~pi32  & ~n28164;
  assign n28170 = ~n42690 & ~n42691;
  assign n28171 = ~n28023 & n28039;
  assign n28172 = ~n28023 & ~n28040;
  assign n28173 = ~n28022 & ~n28171;
  assign n28174 = n28170 & n42692;
  assign n28175 = ~n28170 & ~n42692;
  assign n28176 = ~n28174 & ~n28175;
  assign n28177 = n733 & n9277;
  assign n28178 = pi106  & n37510;
  assign n28179 = pi108  & n746;
  assign n28180 = pi107  & n748;
  assign n28181 = ~n28179 & ~n28180;
  assign n28182 = ~n28178 & ~n28180;
  assign n28183 = ~n28179 & n28182;
  assign n28184 = ~n28178 & n28181;
  assign n28185 = ~n28177 & n42693;
  assign n28186 = pi41  & ~n28185;
  assign n28187 = pi41  & ~n28186;
  assign n28188 = pi41  & n28185;
  assign n28189 = ~n28185 & ~n28186;
  assign n28190 = ~pi41  & ~n28185;
  assign n28191 = ~n42694 & ~n42695;
  assign n28192 = ~n27963 & ~n27969;
  assign n28193 = n940 & n8229;
  assign n28194 = pi103  & n37541;
  assign n28195 = pi105  & n953;
  assign n28196 = pi104  & n955;
  assign n28197 = ~n28195 & ~n28196;
  assign n28198 = ~n28194 & ~n28196;
  assign n28199 = ~n28195 & n28198;
  assign n28200 = ~n28194 & n28197;
  assign n28201 = ~n28193 & n42696;
  assign n28202 = pi44  & ~n28201;
  assign n28203 = pi44  & ~n28202;
  assign n28204 = pi44  & n28201;
  assign n28205 = ~n28201 & ~n28202;
  assign n28206 = ~pi44  & ~n28201;
  assign n28207 = ~n42697 & ~n42698;
  assign n28208 = ~n27943 & ~n27961;
  assign n28209 = n785 & n6819;
  assign n28210 = pi100  & n37520;
  assign n28211 = pi102  & n787;
  assign n28212 = pi101  & n795;
  assign n28213 = ~n28211 & ~n28212;
  assign n28214 = ~n28210 & ~n28212;
  assign n28215 = ~n28211 & n28214;
  assign n28216 = ~n28210 & n28213;
  assign n28217 = ~n28209 & n42699;
  assign n28218 = pi47  & ~n28217;
  assign n28219 = pi47  & ~n28218;
  assign n28220 = pi47  & n28217;
  assign n28221 = ~n28217 & ~n28218;
  assign n28222 = ~pi47  & ~n28217;
  assign n28223 = ~n42700 & ~n42701;
  assign n28224 = n894 & n5578;
  assign n28225 = pi97  & n37580;
  assign n28226 = pi99  & n896;
  assign n28227 = pi98  & n904;
  assign n28228 = ~n28226 & ~n28227;
  assign n28229 = ~n28225 & ~n28227;
  assign n28230 = ~n28226 & n28229;
  assign n28231 = ~n28225 & n28228;
  assign n28232 = ~n28224 & n42702;
  assign n28233 = pi50  & ~n28232;
  assign n28234 = pi50  & ~n28233;
  assign n28235 = pi50  & n28232;
  assign n28236 = ~n28232 & ~n28233;
  assign n28237 = ~pi50  & ~n28232;
  assign n28238 = ~n42703 & ~n42704;
  assign n28239 = ~n27892 & ~n27908;
  assign n28240 = ~n27891 & ~n27910;
  assign n28241 = ~n27891 & ~n28239;
  assign n28242 = n1971 & n5281;
  assign n28243 = pi94  & n37864;
  assign n28244 = pi96  & n1973;
  assign n28245 = pi95  & n1981;
  assign n28246 = ~n28244 & ~n28245;
  assign n28247 = ~n28243 & ~n28245;
  assign n28248 = ~n28244 & n28247;
  assign n28249 = ~n28243 & n28246;
  assign n28250 = ~n28242 & n42706;
  assign n28251 = pi53  & ~n28250;
  assign n28252 = pi53  & ~n28251;
  assign n28253 = pi53  & n28250;
  assign n28254 = ~n28250 & ~n28251;
  assign n28255 = ~pi53  & ~n28250;
  assign n28256 = ~n42707 & ~n42708;
  assign n28257 = ~n27881 & ~n27888;
  assign n28258 = n3566 & n7882;
  assign n28259 = pi88  & n39128;
  assign n28260 = pi90  & n7884;
  assign n28261 = pi89  & n7892;
  assign n28262 = ~n28260 & ~n28261;
  assign n28263 = ~n28259 & ~n28261;
  assign n28264 = ~n28260 & n28263;
  assign n28265 = ~n28259 & n28262;
  assign n28266 = ~n28258 & n42709;
  assign n28267 = pi59  & ~n28266;
  assign n28268 = pi59  & ~n28267;
  assign n28269 = pi59  & n28266;
  assign n28270 = ~n28266 & ~n28267;
  assign n28271 = ~pi59  & ~n28266;
  assign n28272 = ~n42710 & ~n42711;
  assign n28273 = ~n27836 & ~n27854;
  assign n28274 = pi84  & ~n40814;
  assign n28275 = pi83  & n18285;
  assign n28276 = ~n28274 & ~n28275;
  assign n28277 = ~n27834 & n28276;
  assign n28278 = n27834 & ~n28276;
  assign n28279 = ~n28277 & ~n28278;
  assign n28280 = n636 & n12674;
  assign n28281 = pi85  & n40107;
  assign n28282 = pi87  & n12676;
  assign n28283 = pi86  & n12684;
  assign n28284 = ~n28282 & ~n28283;
  assign n28285 = ~n28281 & ~n28283;
  assign n28286 = ~n28282 & n28285;
  assign n28287 = ~n28281 & n28284;
  assign n28288 = ~n12674 & n42712;
  assign n28289 = ~n636 & n42712;
  assign n28290 = ~n28288 & ~n28289;
  assign n28291 = ~n28280 & n42712;
  assign n28292 = pi62  & ~n42713;
  assign n28293 = ~pi62  & n42713;
  assign n28294 = ~n28292 & ~n28293;
  assign n28295 = n28279 & ~n28294;
  assign n28296 = ~n28279 & n28294;
  assign n28297 = ~n28295 & ~n28296;
  assign n28298 = ~n28273 & n28297;
  assign n28299 = n28273 & ~n28297;
  assign n28300 = ~n28298 & ~n28299;
  assign n28301 = ~n28272 & n28300;
  assign n28302 = n28272 & ~n28300;
  assign n28303 = ~n28301 & ~n28302;
  assign n28304 = ~n27858 & ~n27874;
  assign n28305 = ~n27857 & ~n27876;
  assign n28306 = ~n27857 & ~n28304;
  assign n28307 = n28303 & ~n42714;
  assign n28308 = ~n28303 & n42714;
  assign n28309 = ~n28307 & ~n28308;
  assign n28310 = n4312 & n4544;
  assign n28311 = pi91  & n38376;
  assign n28312 = pi93  & n4314;
  assign n28313 = pi92  & n4322;
  assign n28314 = ~n28312 & ~n28313;
  assign n28315 = ~n28311 & ~n28313;
  assign n28316 = ~n28312 & n28315;
  assign n28317 = ~n28311 & n28314;
  assign n28318 = ~n28310 & n42715;
  assign n28319 = pi56  & ~n28318;
  assign n28320 = pi56  & ~n28319;
  assign n28321 = pi56  & n28318;
  assign n28322 = ~n28318 & ~n28319;
  assign n28323 = ~pi56  & ~n28318;
  assign n28324 = ~n42716 & ~n42717;
  assign n28325 = ~n28309 & n28324;
  assign n28326 = n28309 & ~n28324;
  assign n28327 = n28309 & ~n28326;
  assign n28328 = ~n28324 & ~n28326;
  assign n28329 = ~n28327 & ~n28328;
  assign n28330 = ~n28325 & ~n28326;
  assign n28331 = ~n28257 & ~n42718;
  assign n28332 = n28257 & n42718;
  assign n28333 = ~n42718 & ~n28331;
  assign n28334 = ~n28257 & ~n28331;
  assign n28335 = ~n28333 & ~n28334;
  assign n28336 = ~n28331 & ~n28332;
  assign n28337 = n28256 & n42719;
  assign n28338 = ~n28256 & ~n42719;
  assign n28339 = n28256 & ~n42719;
  assign n28340 = ~n28256 & n42719;
  assign n28341 = ~n28339 & ~n28340;
  assign n28342 = ~n28337 & ~n28338;
  assign n28343 = ~n42705 & ~n42720;
  assign n28344 = n42705 & n42720;
  assign n28345 = ~n28343 & ~n28344;
  assign n28346 = ~n28238 & n28345;
  assign n28347 = n28238 & ~n28345;
  assign n28348 = ~n28346 & ~n28347;
  assign n28349 = ~n27916 & n27932;
  assign n28350 = ~n27916 & ~n27933;
  assign n28351 = ~n27915 & ~n28349;
  assign n28352 = n28348 & ~n42721;
  assign n28353 = ~n28348 & n42721;
  assign n28354 = ~n28352 & ~n28353;
  assign n28355 = ~n28223 & n28354;
  assign n28356 = n28223 & ~n28354;
  assign n28357 = ~n28355 & ~n28356;
  assign n28358 = ~n28208 & n28357;
  assign n28359 = n28208 & ~n28357;
  assign n28360 = ~n28358 & ~n28359;
  assign n28361 = ~n28207 & n28360;
  assign n28362 = n28207 & ~n28360;
  assign n28363 = ~n28361 & ~n28362;
  assign n28364 = ~n28192 & n28363;
  assign n28365 = n28192 & ~n28363;
  assign n28366 = ~n28364 & ~n28365;
  assign n28367 = ~n28191 & n28366;
  assign n28368 = n28191 & ~n28366;
  assign n28369 = ~n28367 & ~n28368;
  assign n28370 = ~n27974 & n27991;
  assign n28371 = ~n27974 & ~n27992;
  assign n28372 = ~n27975 & ~n28370;
  assign n28373 = n28369 & ~n42722;
  assign n28374 = ~n28369 & n42722;
  assign n28375 = ~n28373 & ~n28374;
  assign n28376 = n565 & n691;
  assign n28377 = pi109  & n37503;
  assign n28378 = pi111  & n704;
  assign n28379 = pi110  & n706;
  assign n28380 = ~n28378 & ~n28379;
  assign n28381 = ~n28377 & ~n28379;
  assign n28382 = ~n28378 & n28381;
  assign n28383 = ~n28377 & n28380;
  assign n28384 = ~n28376 & n42723;
  assign n28385 = pi38  & ~n28384;
  assign n28386 = pi38  & ~n28385;
  assign n28387 = pi38  & n28384;
  assign n28388 = ~n28384 & ~n28385;
  assign n28389 = ~pi38  & ~n28384;
  assign n28390 = ~n42724 & ~n42725;
  assign n28391 = n28375 & ~n28390;
  assign n28392 = ~n28375 & n28390;
  assign n28393 = n28375 & ~n28391;
  assign n28394 = ~n28390 & ~n28391;
  assign n28395 = ~n28393 & ~n28394;
  assign n28396 = ~n28391 & ~n28392;
  assign n28397 = ~n27999 & n28015;
  assign n28398 = ~n27999 & ~n28017;
  assign n28399 = ~n27998 & ~n28397;
  assign n28400 = n42726 & n42727;
  assign n28401 = ~n42726 & ~n42727;
  assign n28402 = ~n28400 & ~n28401;
  assign n28403 = n2104 & n11258;
  assign n28404 = pi112  & n37758;
  assign n28405 = pi114  & n2117;
  assign n28406 = pi113  & n2119;
  assign n28407 = ~n28405 & ~n28406;
  assign n28408 = ~n28404 & ~n28406;
  assign n28409 = ~n28405 & n28408;
  assign n28410 = ~n28404 & n28407;
  assign n28411 = ~n28403 & n42728;
  assign n28412 = pi35  & ~n28411;
  assign n28413 = pi35  & ~n28412;
  assign n28414 = pi35  & n28411;
  assign n28415 = ~n28411 & ~n28412;
  assign n28416 = ~pi35  & ~n28411;
  assign n28417 = ~n42729 & ~n42730;
  assign n28418 = n28402 & ~n28417;
  assign n28419 = ~n28402 & n28417;
  assign n28420 = ~n28418 & ~n28419;
  assign n28421 = n28176 & ~n28419;
  assign n28422 = ~n28418 & n28421;
  assign n28423 = n28176 & n28420;
  assign n28424 = ~n28176 & ~n28420;
  assign n28425 = n28176 & ~n42731;
  assign n28426 = ~n28419 & ~n42731;
  assign n28427 = ~n28418 & n28426;
  assign n28428 = n28420 & ~n42731;
  assign n28429 = ~n28425 & ~n42732;
  assign n28430 = ~n42731 & ~n28424;
  assign n28431 = n607 & n14913;
  assign n28432 = pi118  & n37489;
  assign n28433 = pi120  & n620;
  assign n28434 = pi119  & n622;
  assign n28435 = ~n28433 & ~n28434;
  assign n28436 = ~n28432 & ~n28434;
  assign n28437 = ~n28433 & n28436;
  assign n28438 = ~n28432 & n28435;
  assign n28439 = ~n28431 & n42734;
  assign n28440 = pi29  & ~n28439;
  assign n28441 = pi29  & ~n28440;
  assign n28442 = pi29  & n28439;
  assign n28443 = ~n28439 & ~n28440;
  assign n28444 = ~pi29  & ~n28439;
  assign n28445 = ~n42735 & ~n42736;
  assign n28446 = ~n27793 & ~n28046;
  assign n28447 = ~n28445 & ~n28446;
  assign n28448 = n28445 & n28446;
  assign n28449 = ~n28445 & ~n28447;
  assign n28450 = ~n28445 & n28446;
  assign n28451 = ~n28446 & ~n28447;
  assign n28452 = n28445 & ~n28446;
  assign n28453 = ~n42737 & ~n42738;
  assign n28454 = ~n28447 & ~n28448;
  assign n28455 = ~n42733 & ~n42739;
  assign n28456 = n42733 & n42739;
  assign n28457 = n42733 & ~n42739;
  assign n28458 = ~n42733 & n42739;
  assign n28459 = ~n28457 & ~n28458;
  assign n28460 = ~n28455 & ~n28456;
  assign n28461 = n28155 & ~n42740;
  assign n28462 = ~n42740 & ~n28461;
  assign n28463 = ~n28155 & ~n42740;
  assign n28464 = n28155 & ~n28461;
  assign n28465 = n28155 & n42740;
  assign n28466 = ~n28155 & n42740;
  assign n28467 = ~n28461 & ~n28466;
  assign n28468 = ~n42741 & ~n42742;
  assign n28469 = ~n42685 & n42743;
  assign n28470 = n42685 & ~n42743;
  assign n28471 = ~n42685 & ~n42743;
  assign n28472 = n42685 & n42743;
  assign n28473 = ~n28471 & ~n28472;
  assign n28474 = ~n28469 & ~n28470;
  assign n28475 = ~n42679 & ~n42744;
  assign n28476 = n42679 & n42744;
  assign n28477 = ~n28475 & ~n28476;
  assign n28478 = ~n28091 & n28477;
  assign n28479 = n28091 & ~n28477;
  assign n28480 = ~n28478 & ~n28479;
  assign n28481 = ~n28090 & n28480;
  assign n28482 = n28090 & ~n28480;
  assign po83  = ~n28481 & ~n28482;
  assign n28484 = ~n28107 & ~n28475;
  assign n28485 = n4492 & n15111;
  assign n28486 = pi122  & n38208;
  assign n28487 = pi124  & n4507;
  assign n28488 = pi123  & n4509;
  assign n28489 = ~n28487 & ~n28488;
  assign n28490 = ~n28486 & ~n28488;
  assign n28491 = ~n28487 & n28490;
  assign n28492 = ~n28486 & n28489;
  assign n28493 = ~n28485 & n42745;
  assign n28494 = pi26  & ~n28493;
  assign n28495 = pi26  & ~n28494;
  assign n28496 = pi26  & n28493;
  assign n28497 = ~n28493 & ~n28494;
  assign n28498 = ~pi26  & ~n28493;
  assign n28499 = ~n42746 & ~n42747;
  assign n28500 = ~n28154 & n42740;
  assign n28501 = ~n28154 & ~n28461;
  assign n28502 = ~n28153 & ~n28500;
  assign n28503 = n28499 & n42748;
  assign n28504 = ~n28499 & ~n42748;
  assign n28505 = ~n28503 & ~n28504;
  assign n28506 = n649 & n13057;
  assign n28507 = pi116  & n37496;
  assign n28508 = pi118  & n662;
  assign n28509 = pi117  & n664;
  assign n28510 = ~n28508 & ~n28509;
  assign n28511 = ~n28507 & ~n28509;
  assign n28512 = ~n28508 & n28511;
  assign n28513 = ~n28507 & n28510;
  assign n28514 = ~n28506 & n42749;
  assign n28515 = pi32  & ~n28514;
  assign n28516 = pi32  & ~n28515;
  assign n28517 = pi32  & n28514;
  assign n28518 = ~n28514 & ~n28515;
  assign n28519 = ~pi32  & ~n28514;
  assign n28520 = ~n42750 & ~n42751;
  assign n28521 = ~n28175 & ~n42731;
  assign n28522 = n28520 & n28521;
  assign n28523 = ~n28520 & ~n28521;
  assign n28524 = ~n28522 & ~n28523;
  assign n28525 = ~n28401 & ~n28418;
  assign n28526 = ~n28364 & ~n28367;
  assign n28527 = ~n28358 & ~n28361;
  assign n28528 = ~n28352 & ~n28355;
  assign n28529 = ~n28343 & ~n28346;
  assign n28530 = n894 & n6474;
  assign n28531 = pi98  & n37580;
  assign n28532 = pi100  & n896;
  assign n28533 = pi99  & n904;
  assign n28534 = ~n28532 & ~n28533;
  assign n28535 = ~n28531 & ~n28533;
  assign n28536 = ~n28532 & n28535;
  assign n28537 = ~n28531 & n28534;
  assign n28538 = ~n28530 & n42752;
  assign n28539 = pi50  & ~n28538;
  assign n28540 = pi50  & ~n28539;
  assign n28541 = pi50  & n28538;
  assign n28542 = ~n28538 & ~n28539;
  assign n28543 = ~pi50  & ~n28538;
  assign n28544 = ~n42753 & ~n42754;
  assign n28545 = ~n28308 & ~n28324;
  assign n28546 = ~n28307 & ~n28326;
  assign n28547 = ~n28307 & ~n28545;
  assign n28548 = ~n28298 & ~n28301;
  assign n28549 = n594 & n7882;
  assign n28550 = pi89  & n39128;
  assign n28551 = pi91  & n7884;
  assign n28552 = pi90  & n7892;
  assign n28553 = ~n28551 & ~n28552;
  assign n28554 = ~n28550 & ~n28552;
  assign n28555 = ~n28551 & n28554;
  assign n28556 = ~n28550 & n28553;
  assign n28557 = ~n28549 & n42756;
  assign n28558 = pi59  & ~n28557;
  assign n28559 = pi59  & ~n28558;
  assign n28560 = pi59  & n28557;
  assign n28561 = ~n28557 & ~n28558;
  assign n28562 = ~pi59  & ~n28557;
  assign n28563 = ~n42757 & ~n42758;
  assign n28564 = ~n28277 & ~n28295;
  assign n28565 = pi85  & ~n40814;
  assign n28566 = pi84  & n18285;
  assign n28567 = ~n28565 & ~n28566;
  assign n28568 = ~pi20  & ~n28567;
  assign n28569 = pi20  & n28567;
  assign n28570 = ~n28568 & ~n28569;
  assign n28571 = ~n28276 & n28570;
  assign n28572 = n28276 & ~n28570;
  assign n28573 = ~n28571 & ~n28572;
  assign n28574 = n3354 & n12674;
  assign n28575 = pi86  & n40107;
  assign n28576 = pi88  & n12676;
  assign n28577 = pi87  & n12684;
  assign n28578 = ~n28576 & ~n28577;
  assign n28579 = ~n28575 & ~n28577;
  assign n28580 = ~n28576 & n28579;
  assign n28581 = ~n28575 & n28578;
  assign n28582 = ~n28574 & n42759;
  assign n28583 = pi62  & ~n28582;
  assign n28584 = pi62  & ~n28583;
  assign n28585 = pi62  & n28582;
  assign n28586 = ~n28582 & ~n28583;
  assign n28587 = ~pi62  & ~n28582;
  assign n28588 = ~n42760 & ~n42761;
  assign n28589 = n28573 & ~n28588;
  assign n28590 = ~n28573 & n28588;
  assign n28591 = n28573 & ~n28589;
  assign n28592 = n28573 & n28588;
  assign n28593 = ~n28588 & ~n28589;
  assign n28594 = ~n28573 & ~n28588;
  assign n28595 = ~n42762 & ~n42763;
  assign n28596 = ~n28589 & ~n28590;
  assign n28597 = ~n28564 & ~n42764;
  assign n28598 = n28564 & n42764;
  assign n28599 = ~n42764 & ~n28597;
  assign n28600 = ~n28564 & ~n28597;
  assign n28601 = ~n28599 & ~n28600;
  assign n28602 = ~n28597 & ~n28598;
  assign n28603 = ~n28563 & ~n42765;
  assign n28604 = n28563 & n42765;
  assign n28605 = ~n42765 & ~n28603;
  assign n28606 = n28563 & ~n42765;
  assign n28607 = ~n28563 & ~n28603;
  assign n28608 = ~n28563 & n42765;
  assign n28609 = ~n42766 & ~n42767;
  assign n28610 = ~n28603 & ~n28604;
  assign n28611 = n28548 & n42768;
  assign n28612 = ~n28548 & ~n42768;
  assign n28613 = ~n28611 & ~n28612;
  assign n28614 = n4312 & n4524;
  assign n28615 = pi92  & n38376;
  assign n28616 = pi94  & n4314;
  assign n28617 = pi93  & n4322;
  assign n28618 = ~n28616 & ~n28617;
  assign n28619 = ~n28615 & ~n28617;
  assign n28620 = ~n28616 & n28619;
  assign n28621 = ~n28615 & n28618;
  assign n28622 = ~n28614 & n42769;
  assign n28623 = pi56  & ~n28622;
  assign n28624 = pi56  & ~n28623;
  assign n28625 = pi56  & n28622;
  assign n28626 = ~n28622 & ~n28623;
  assign n28627 = ~pi56  & ~n28622;
  assign n28628 = ~n42770 & ~n42771;
  assign n28629 = n28613 & ~n28628;
  assign n28630 = ~n28613 & n28628;
  assign n28631 = n28613 & ~n28629;
  assign n28632 = n28613 & n28628;
  assign n28633 = ~n28628 & ~n28629;
  assign n28634 = ~n28613 & ~n28628;
  assign n28635 = ~n42772 & ~n42773;
  assign n28636 = ~n28629 & ~n28630;
  assign n28637 = n42755 & n42774;
  assign n28638 = ~n42755 & ~n42774;
  assign n28639 = ~n28637 & ~n28638;
  assign n28640 = n1971 & n5630;
  assign n28641 = pi95  & n37864;
  assign n28642 = pi97  & n1973;
  assign n28643 = pi96  & n1981;
  assign n28644 = ~n28642 & ~n28643;
  assign n28645 = ~n28641 & ~n28643;
  assign n28646 = ~n28642 & n28645;
  assign n28647 = ~n28641 & n28644;
  assign n28648 = ~n28640 & n42775;
  assign n28649 = pi53  & ~n28648;
  assign n28650 = pi53  & ~n28649;
  assign n28651 = pi53  & n28648;
  assign n28652 = ~n28648 & ~n28649;
  assign n28653 = ~pi53  & ~n28648;
  assign n28654 = ~n42776 & ~n42777;
  assign n28655 = n28256 & ~n28331;
  assign n28656 = ~n28331 & ~n28338;
  assign n28657 = ~n28332 & ~n28655;
  assign n28658 = ~n28654 & ~n42778;
  assign n28659 = n28654 & n42778;
  assign n28660 = ~n28658 & ~n28659;
  assign n28661 = n28639 & n28660;
  assign n28662 = ~n28639 & ~n28660;
  assign n28663 = ~n28639 & n28660;
  assign n28664 = n28639 & ~n28660;
  assign n28665 = ~n28663 & ~n28664;
  assign n28666 = ~n28661 & ~n28662;
  assign n28667 = ~n28544 & ~n42779;
  assign n28668 = n28544 & n42779;
  assign n28669 = ~n28667 & ~n28668;
  assign n28670 = n28529 & ~n28669;
  assign n28671 = ~n28529 & n28669;
  assign n28672 = ~n28670 & ~n28671;
  assign n28673 = n785 & n6787;
  assign n28674 = pi101  & n37520;
  assign n28675 = pi103  & n787;
  assign n28676 = pi102  & n795;
  assign n28677 = ~n28675 & ~n28676;
  assign n28678 = ~n28674 & ~n28676;
  assign n28679 = ~n28675 & n28678;
  assign n28680 = ~n28674 & n28677;
  assign n28681 = ~n28673 & n42780;
  assign n28682 = pi47  & ~n28681;
  assign n28683 = pi47  & ~n28682;
  assign n28684 = pi47  & n28681;
  assign n28685 = ~n28681 & ~n28682;
  assign n28686 = ~pi47  & ~n28681;
  assign n28687 = ~n42781 & ~n42782;
  assign n28688 = n28672 & ~n28687;
  assign n28689 = ~n28672 & n28687;
  assign n28690 = n28672 & ~n28688;
  assign n28691 = n28672 & n28687;
  assign n28692 = ~n28687 & ~n28688;
  assign n28693 = ~n28672 & ~n28687;
  assign n28694 = ~n42783 & ~n42784;
  assign n28695 = ~n28688 & ~n28689;
  assign n28696 = n28528 & n42785;
  assign n28697 = ~n28528 & ~n42785;
  assign n28698 = ~n28696 & ~n28697;
  assign n28699 = n940 & n8209;
  assign n28700 = pi104  & n37541;
  assign n28701 = pi106  & n953;
  assign n28702 = pi105  & n955;
  assign n28703 = ~n28701 & ~n28702;
  assign n28704 = ~n28700 & ~n28702;
  assign n28705 = ~n28701 & n28704;
  assign n28706 = ~n28700 & n28703;
  assign n28707 = ~n28699 & n42786;
  assign n28708 = pi44  & ~n28707;
  assign n28709 = pi44  & ~n28708;
  assign n28710 = pi44  & n28707;
  assign n28711 = ~n28707 & ~n28708;
  assign n28712 = ~pi44  & ~n28707;
  assign n28713 = ~n42787 & ~n42788;
  assign n28714 = n28698 & ~n28713;
  assign n28715 = ~n28698 & n28713;
  assign n28716 = n28698 & ~n28714;
  assign n28717 = n28698 & n28713;
  assign n28718 = ~n28713 & ~n28714;
  assign n28719 = ~n28698 & ~n28713;
  assign n28720 = ~n42789 & ~n42790;
  assign n28721 = ~n28714 & ~n28715;
  assign n28722 = n28527 & n42791;
  assign n28723 = ~n28527 & ~n42791;
  assign n28724 = ~n28722 & ~n28723;
  assign n28725 = n733 & n9701;
  assign n28726 = pi107  & n37510;
  assign n28727 = pi109  & n746;
  assign n28728 = pi108  & n748;
  assign n28729 = ~n28727 & ~n28728;
  assign n28730 = ~n28726 & ~n28728;
  assign n28731 = ~n28727 & n28730;
  assign n28732 = ~n28726 & n28729;
  assign n28733 = ~n28725 & n42792;
  assign n28734 = pi41  & ~n28733;
  assign n28735 = pi41  & ~n28734;
  assign n28736 = pi41  & n28733;
  assign n28737 = ~n28733 & ~n28734;
  assign n28738 = ~pi41  & ~n28733;
  assign n28739 = ~n42793 & ~n42794;
  assign n28740 = n28724 & ~n28739;
  assign n28741 = ~n28724 & n28739;
  assign n28742 = n28724 & ~n28740;
  assign n28743 = n28724 & n28739;
  assign n28744 = ~n28739 & ~n28740;
  assign n28745 = ~n28724 & ~n28739;
  assign n28746 = ~n42795 & ~n42796;
  assign n28747 = ~n28740 & ~n28741;
  assign n28748 = n28526 & n42797;
  assign n28749 = ~n28526 & ~n42797;
  assign n28750 = ~n28748 & ~n28749;
  assign n28751 = n691 & n10844;
  assign n28752 = pi110  & n37503;
  assign n28753 = pi112  & n704;
  assign n28754 = pi111  & n706;
  assign n28755 = ~n28753 & ~n28754;
  assign n28756 = ~n28752 & ~n28754;
  assign n28757 = ~n28753 & n28756;
  assign n28758 = ~n28752 & n28755;
  assign n28759 = ~n28751 & n42798;
  assign n28760 = pi38  & ~n28759;
  assign n28761 = pi38  & ~n28760;
  assign n28762 = pi38  & n28759;
  assign n28763 = ~n28759 & ~n28760;
  assign n28764 = ~pi38  & ~n28759;
  assign n28765 = ~n42799 & ~n42800;
  assign n28766 = n28750 & ~n28765;
  assign n28767 = ~n28750 & n28765;
  assign n28768 = n28750 & ~n28766;
  assign n28769 = n28750 & n28765;
  assign n28770 = ~n28765 & ~n28766;
  assign n28771 = ~n28750 & ~n28765;
  assign n28772 = ~n42801 & ~n42802;
  assign n28773 = ~n28766 & ~n28767;
  assign n28774 = ~n28373 & n28390;
  assign n28775 = ~n28373 & ~n28391;
  assign n28776 = ~n28374 & ~n28774;
  assign n28777 = n42803 & n42804;
  assign n28778 = ~n42803 & ~n42804;
  assign n28779 = ~n28777 & ~n28778;
  assign n28780 = n523 & n2104;
  assign n28781 = pi113  & n37758;
  assign n28782 = pi115  & n2117;
  assign n28783 = pi114  & n2119;
  assign n28784 = ~n28782 & ~n28783;
  assign n28785 = ~n28781 & ~n28783;
  assign n28786 = ~n28782 & n28785;
  assign n28787 = ~n28781 & n28784;
  assign n28788 = ~n28780 & n42805;
  assign n28789 = pi35  & ~n28788;
  assign n28790 = pi35  & ~n28789;
  assign n28791 = pi35  & n28788;
  assign n28792 = ~n28788 & ~n28789;
  assign n28793 = ~pi35  & ~n28788;
  assign n28794 = ~n42806 & ~n42807;
  assign n28795 = n28779 & ~n28794;
  assign n28796 = ~n28779 & n28794;
  assign n28797 = ~n28795 & ~n28796;
  assign n28798 = n28525 & ~n28797;
  assign n28799 = ~n28525 & ~n28796;
  assign n28800 = ~n28795 & n28799;
  assign n28801 = ~n28525 & ~n28795;
  assign n28802 = ~n28796 & n28801;
  assign n28803 = ~n28525 & n28797;
  assign n28804 = ~n28525 & ~n42808;
  assign n28805 = ~n28525 & ~n28797;
  assign n28806 = n28525 & ~n28795;
  assign n28807 = ~n28795 & ~n42808;
  assign n28808 = ~n28796 & ~n28806;
  assign n28809 = ~n28796 & n42810;
  assign n28810 = n28525 & n28797;
  assign n28811 = ~n42809 & ~n42811;
  assign n28812 = ~n28798 & ~n42808;
  assign n28813 = n28524 & ~n42812;
  assign n28814 = ~n28524 & n42812;
  assign n28815 = ~n28813 & ~n28814;
  assign n28816 = ~n28447 & ~n28455;
  assign n28817 = n607 & n15091;
  assign n28818 = pi119  & n37489;
  assign n28819 = pi121  & n620;
  assign n28820 = pi120  & n622;
  assign n28821 = ~n28819 & ~n28820;
  assign n28822 = ~n28818 & ~n28820;
  assign n28823 = ~n28819 & n28822;
  assign n28824 = ~n28818 & n28821;
  assign n28825 = ~n28817 & n42813;
  assign n28826 = pi29  & ~n28825;
  assign n28827 = pi29  & ~n28826;
  assign n28828 = pi29  & n28825;
  assign n28829 = ~n28825 & ~n28826;
  assign n28830 = ~pi29  & ~n28825;
  assign n28831 = ~n42814 & ~n42815;
  assign n28832 = ~n28816 & ~n28831;
  assign n28833 = n28816 & n28831;
  assign n28834 = ~n28816 & n28831;
  assign n28835 = n28816 & ~n28831;
  assign n28836 = ~n28834 & ~n28835;
  assign n28837 = ~n28832 & ~n28833;
  assign n28838 = ~n28814 & ~n42816;
  assign n28839 = ~n28813 & n28838;
  assign n28840 = n28815 & ~n42816;
  assign n28841 = ~n28815 & n42816;
  assign n28842 = ~n42816 & ~n42817;
  assign n28843 = ~n28814 & ~n42817;
  assign n28844 = ~n28813 & n28843;
  assign n28845 = n28815 & ~n42817;
  assign n28846 = ~n28842 & ~n42818;
  assign n28847 = ~n42817 & ~n28841;
  assign n28848 = n28505 & ~n42819;
  assign n28849 = ~n28505 & n42819;
  assign n28850 = ~n28848 & ~n28849;
  assign n28851 = ~n28129 & ~n28469;
  assign n28852 = n5576 & n40885;
  assign n28853 = pi125  & n38406;
  assign n28854 = pi127  & n5591;
  assign n28855 = pi126  & n5593;
  assign n28856 = ~n28854 & ~n28855;
  assign n28857 = ~n28853 & ~n28855;
  assign n28858 = ~n28854 & n28857;
  assign n28859 = ~n28853 & n28856;
  assign n28860 = ~n28852 & n42820;
  assign n28861 = pi23  & ~n28860;
  assign n28862 = pi23  & ~n28861;
  assign n28863 = pi23  & n28860;
  assign n28864 = ~n28860 & ~n28861;
  assign n28865 = ~pi23  & ~n28860;
  assign n28866 = ~n42821 & ~n42822;
  assign n28867 = ~n28851 & ~n28866;
  assign n28868 = n28851 & n28866;
  assign n28869 = ~n28851 & ~n28867;
  assign n28870 = ~n28851 & n28866;
  assign n28871 = ~n28866 & ~n28867;
  assign n28872 = n28851 & ~n28866;
  assign n28873 = ~n42823 & ~n42824;
  assign n28874 = ~n28867 & ~n28868;
  assign n28875 = ~n28849 & ~n42825;
  assign n28876 = ~n28848 & n28875;
  assign n28877 = n28850 & ~n42825;
  assign n28878 = ~n28850 & n42825;
  assign n28879 = ~n42825 & ~n42826;
  assign n28880 = ~n28850 & ~n42825;
  assign n28881 = n28850 & ~n42826;
  assign n28882 = ~n28849 & ~n42826;
  assign n28883 = ~n28848 & n28882;
  assign n28884 = n28850 & n42825;
  assign n28885 = ~n42827 & ~n42828;
  assign n28886 = ~n42826 & ~n28878;
  assign n28887 = n28484 & n42829;
  assign n28888 = ~n28484 & ~n42829;
  assign n28889 = ~n28887 & ~n28888;
  assign n28890 = ~n28478 & ~n28481;
  assign n28891 = n28889 & ~n28890;
  assign n28892 = ~n28889 & n28890;
  assign po84  = ~n28891 & ~n28892;
  assign n28894 = ~n28867 & ~n42826;
  assign n28895 = ~n28504 & ~n28848;
  assign n28896 = n5576 & n40891;
  assign n28897 = pi126  & n38406;
  assign n28898 = pi127  & n5593;
  assign n28899 = ~n28897 & ~n28898;
  assign n28900 = ~n5576 & n28899;
  assign n28901 = ~n40891 & n28899;
  assign n28902 = ~n28900 & ~n28901;
  assign n28903 = ~n28896 & n28899;
  assign n28904 = pi23  & ~n42830;
  assign n28905 = ~pi23  & n42830;
  assign n28906 = ~n28904 & ~n28905;
  assign n28907 = ~n28895 & ~n28906;
  assign n28908 = n28895 & n28906;
  assign n28909 = ~n28907 & ~n28908;
  assign n28910 = n4492 & n15068;
  assign n28911 = pi123  & n38208;
  assign n28912 = pi125  & n4507;
  assign n28913 = pi124  & n4509;
  assign n28914 = ~n28912 & ~n28913;
  assign n28915 = ~n28911 & ~n28913;
  assign n28916 = ~n28912 & n28915;
  assign n28917 = ~n28911 & n28914;
  assign n28918 = ~n28910 & n42831;
  assign n28919 = pi26  & ~n28918;
  assign n28920 = pi26  & ~n28919;
  assign n28921 = pi26  & n28918;
  assign n28922 = ~n28918 & ~n28919;
  assign n28923 = ~pi26  & ~n28918;
  assign n28924 = ~n42832 & ~n42833;
  assign n28925 = ~n28832 & ~n42817;
  assign n28926 = n28924 & n28925;
  assign n28927 = ~n28924 & ~n28925;
  assign n28928 = ~n28926 & ~n28927;
  assign n28929 = ~n28523 & ~n28813;
  assign n28930 = n607 & n15049;
  assign n28931 = pi120  & n37489;
  assign n28932 = pi122  & n620;
  assign n28933 = pi121  & n622;
  assign n28934 = ~n28932 & ~n28933;
  assign n28935 = ~n28931 & ~n28933;
  assign n28936 = ~n28932 & n28935;
  assign n28937 = ~n28931 & n28934;
  assign n28938 = ~n607 & n42834;
  assign n28939 = ~n15049 & n42834;
  assign n28940 = ~n28938 & ~n28939;
  assign n28941 = ~n28930 & n42834;
  assign n28942 = pi29  & ~n42835;
  assign n28943 = ~pi29  & n42835;
  assign n28944 = ~n28942 & ~n28943;
  assign n28945 = ~n28929 & ~n28944;
  assign n28946 = n28929 & n28944;
  assign n28947 = ~n28945 & ~n28946;
  assign n28948 = n649 & n13027;
  assign n28949 = pi117  & n37496;
  assign n28950 = pi119  & n662;
  assign n28951 = pi118  & n664;
  assign n28952 = ~n28950 & ~n28951;
  assign n28953 = ~n28949 & ~n28951;
  assign n28954 = ~n28950 & n28953;
  assign n28955 = ~n28949 & n28952;
  assign n28956 = ~n28948 & n42836;
  assign n28957 = pi32  & ~n28956;
  assign n28958 = pi32  & ~n28957;
  assign n28959 = pi32  & n28956;
  assign n28960 = ~n28956 & ~n28957;
  assign n28961 = ~pi32  & ~n28956;
  assign n28962 = ~n42837 & ~n42838;
  assign n28963 = ~n42810 & ~n28962;
  assign n28964 = n42810 & n28962;
  assign n28965 = ~n42810 & n28962;
  assign n28966 = n42810 & ~n28962;
  assign n28967 = ~n28965 & ~n28966;
  assign n28968 = ~n28963 & ~n28964;
  assign n28969 = ~n28766 & ~n28778;
  assign n28970 = ~n28740 & ~n28749;
  assign n28971 = ~n28714 & ~n28723;
  assign n28972 = ~n28688 & ~n28697;
  assign n28973 = n785 & n8136;
  assign n28974 = pi102  & n37520;
  assign n28975 = pi104  & n787;
  assign n28976 = pi103  & n795;
  assign n28977 = ~n28975 & ~n28976;
  assign n28978 = ~n28974 & ~n28976;
  assign n28979 = ~n28975 & n28978;
  assign n28980 = ~n28974 & n28977;
  assign n28981 = ~n28973 & n42840;
  assign n28982 = pi47  & ~n28981;
  assign n28983 = pi47  & ~n28982;
  assign n28984 = pi47  & n28981;
  assign n28985 = ~n28981 & ~n28982;
  assign n28986 = ~pi47  & ~n28981;
  assign n28987 = ~n42841 & ~n42842;
  assign n28988 = ~n28667 & ~n28671;
  assign n28989 = ~n28629 & ~n28638;
  assign n28990 = ~n28603 & ~n28612;
  assign n28991 = n4453 & n7882;
  assign n28992 = pi90  & n39128;
  assign n28993 = pi92  & n7884;
  assign n28994 = pi91  & n7892;
  assign n28995 = ~n28993 & ~n28994;
  assign n28996 = ~n28992 & ~n28994;
  assign n28997 = ~n28993 & n28996;
  assign n28998 = ~n28992 & n28995;
  assign n28999 = ~n28991 & n42843;
  assign n29000 = pi59  & ~n28999;
  assign n29001 = pi59  & ~n29000;
  assign n29002 = pi59  & n28999;
  assign n29003 = ~n28999 & ~n29000;
  assign n29004 = ~pi59  & ~n28999;
  assign n29005 = ~n42844 & ~n42845;
  assign n29006 = ~n28589 & ~n28597;
  assign n29007 = ~n28568 & ~n28571;
  assign n29008 = pi86  & ~n40814;
  assign n29009 = pi85  & n18285;
  assign n29010 = ~n29008 & ~n29009;
  assign n29011 = n29007 & ~n29010;
  assign n29012 = ~n29007 & n29010;
  assign n29013 = ~n29011 & ~n29012;
  assign n29014 = n3591 & n12674;
  assign n29015 = pi87  & n40107;
  assign n29016 = pi89  & n12676;
  assign n29017 = pi88  & n12684;
  assign n29018 = ~n29016 & ~n29017;
  assign n29019 = ~n29015 & ~n29017;
  assign n29020 = ~n29016 & n29019;
  assign n29021 = ~n29015 & n29018;
  assign n29022 = ~n12674 & n42846;
  assign n29023 = ~n3591 & n42846;
  assign n29024 = ~n29022 & ~n29023;
  assign n29025 = ~n29014 & n42846;
  assign n29026 = pi62  & ~n42847;
  assign n29027 = ~pi62  & n42847;
  assign n29028 = ~n29026 & ~n29027;
  assign n29029 = n29013 & ~n29028;
  assign n29030 = ~n29013 & n29028;
  assign n29031 = ~n29029 & ~n29030;
  assign n29032 = ~n29006 & n29031;
  assign n29033 = n29006 & ~n29031;
  assign n29034 = ~n29032 & ~n29033;
  assign n29035 = ~n29005 & n29034;
  assign n29036 = n29005 & ~n29034;
  assign n29037 = ~n29035 & ~n29036;
  assign n29038 = ~n28990 & n29037;
  assign n29039 = n28990 & ~n29037;
  assign n29040 = ~n29038 & ~n29039;
  assign n29041 = n4312 & n4494;
  assign n29042 = pi93  & n38376;
  assign n29043 = pi95  & n4314;
  assign n29044 = pi94  & n4322;
  assign n29045 = ~n29043 & ~n29044;
  assign n29046 = ~n29042 & ~n29044;
  assign n29047 = ~n29043 & n29046;
  assign n29048 = ~n29042 & n29045;
  assign n29049 = ~n29041 & n42848;
  assign n29050 = pi56  & ~n29049;
  assign n29051 = pi56  & ~n29050;
  assign n29052 = pi56  & n29049;
  assign n29053 = ~n29049 & ~n29050;
  assign n29054 = ~pi56  & ~n29049;
  assign n29055 = ~n42849 & ~n42850;
  assign n29056 = n29040 & ~n29055;
  assign n29057 = ~n29040 & n29055;
  assign n29058 = n29040 & ~n29056;
  assign n29059 = ~n29055 & ~n29056;
  assign n29060 = ~n29058 & ~n29059;
  assign n29061 = ~n29056 & ~n29057;
  assign n29062 = n28989 & n42851;
  assign n29063 = ~n28989 & ~n42851;
  assign n29064 = ~n29062 & ~n29063;
  assign n29065 = n1971 & n5610;
  assign n29066 = pi96  & n37864;
  assign n29067 = pi98  & n1973;
  assign n29068 = pi97  & n1981;
  assign n29069 = ~n29067 & ~n29068;
  assign n29070 = ~n29066 & ~n29068;
  assign n29071 = ~n29067 & n29070;
  assign n29072 = ~n29066 & n29069;
  assign n29073 = ~n29065 & n42852;
  assign n29074 = pi53  & ~n29073;
  assign n29075 = pi53  & ~n29074;
  assign n29076 = pi53  & n29073;
  assign n29077 = ~n29073 & ~n29074;
  assign n29078 = ~pi53  & ~n29073;
  assign n29079 = ~n42853 & ~n42854;
  assign n29080 = ~n29064 & n29079;
  assign n29081 = n29064 & ~n29079;
  assign n29082 = n29064 & ~n29081;
  assign n29083 = ~n29079 & ~n29081;
  assign n29084 = ~n29082 & ~n29083;
  assign n29085 = ~n29080 & ~n29081;
  assign n29086 = ~n28639 & ~n28658;
  assign n29087 = ~n28658 & ~n28661;
  assign n29088 = ~n28659 & ~n29086;
  assign n29089 = n42855 & n42856;
  assign n29090 = ~n42855 & ~n42856;
  assign n29091 = ~n29089 & ~n29090;
  assign n29092 = n894 & n6839;
  assign n29093 = pi99  & n37580;
  assign n29094 = pi101  & n896;
  assign n29095 = pi100  & n904;
  assign n29096 = ~n29094 & ~n29095;
  assign n29097 = ~n29093 & ~n29095;
  assign n29098 = ~n29094 & n29097;
  assign n29099 = ~n29093 & n29096;
  assign n29100 = ~n29092 & n42857;
  assign n29101 = pi50  & ~n29100;
  assign n29102 = pi50  & ~n29101;
  assign n29103 = pi50  & n29100;
  assign n29104 = ~n29100 & ~n29101;
  assign n29105 = ~pi50  & ~n29100;
  assign n29106 = ~n42858 & ~n42859;
  assign n29107 = ~n29091 & n29106;
  assign n29108 = n29091 & ~n29106;
  assign n29109 = ~n29107 & ~n29108;
  assign n29110 = ~n28988 & n29109;
  assign n29111 = n28988 & ~n29109;
  assign n29112 = ~n28988 & ~n29110;
  assign n29113 = n29109 & ~n29110;
  assign n29114 = ~n29112 & ~n29113;
  assign n29115 = ~n29110 & ~n29111;
  assign n29116 = ~n28987 & ~n42860;
  assign n29117 = n28987 & ~n29113;
  assign n29118 = ~n29112 & n29117;
  assign n29119 = n28987 & n42860;
  assign n29120 = ~n29116 & ~n42861;
  assign n29121 = ~n28972 & n29120;
  assign n29122 = n28972 & ~n29120;
  assign n29123 = ~n29121 & ~n29122;
  assign n29124 = n940 & n8177;
  assign n29125 = pi105  & n37541;
  assign n29126 = pi107  & n953;
  assign n29127 = pi106  & n955;
  assign n29128 = ~n29126 & ~n29127;
  assign n29129 = ~n29125 & ~n29127;
  assign n29130 = ~n29126 & n29129;
  assign n29131 = ~n29125 & n29128;
  assign n29132 = ~n29124 & n42862;
  assign n29133 = pi44  & ~n29132;
  assign n29134 = pi44  & ~n29133;
  assign n29135 = pi44  & n29132;
  assign n29136 = ~n29132 & ~n29133;
  assign n29137 = ~pi44  & ~n29132;
  assign n29138 = ~n42863 & ~n42864;
  assign n29139 = n29123 & ~n29138;
  assign n29140 = ~n29123 & n29138;
  assign n29141 = n29123 & ~n29139;
  assign n29142 = ~n29138 & ~n29139;
  assign n29143 = ~n29141 & ~n29142;
  assign n29144 = ~n29139 & ~n29140;
  assign n29145 = n28971 & n42865;
  assign n29146 = ~n28971 & ~n42865;
  assign n29147 = ~n29145 & ~n29146;
  assign n29148 = n733 & n9678;
  assign n29149 = pi108  & n37510;
  assign n29150 = pi110  & n746;
  assign n29151 = pi109  & n748;
  assign n29152 = ~n29150 & ~n29151;
  assign n29153 = ~n29149 & ~n29151;
  assign n29154 = ~n29150 & n29153;
  assign n29155 = ~n29149 & n29152;
  assign n29156 = ~n29148 & n42866;
  assign n29157 = pi41  & ~n29156;
  assign n29158 = pi41  & ~n29157;
  assign n29159 = pi41  & n29156;
  assign n29160 = ~n29156 & ~n29157;
  assign n29161 = ~pi41  & ~n29156;
  assign n29162 = ~n42867 & ~n42868;
  assign n29163 = ~n29147 & n29162;
  assign n29164 = n29147 & ~n29162;
  assign n29165 = n29147 & ~n29164;
  assign n29166 = ~n29162 & ~n29164;
  assign n29167 = ~n29165 & ~n29166;
  assign n29168 = ~n29163 & ~n29164;
  assign n29169 = n28970 & n42869;
  assign n29170 = ~n28970 & ~n42869;
  assign n29171 = ~n29169 & ~n29170;
  assign n29172 = n691 & n11276;
  assign n29173 = pi111  & n37503;
  assign n29174 = pi113  & n704;
  assign n29175 = pi112  & n706;
  assign n29176 = ~n29174 & ~n29175;
  assign n29177 = ~n29173 & ~n29175;
  assign n29178 = ~n29174 & n29177;
  assign n29179 = ~n29173 & n29176;
  assign n29180 = ~n29172 & n42870;
  assign n29181 = pi38  & ~n29180;
  assign n29182 = pi38  & ~n29181;
  assign n29183 = pi38  & n29180;
  assign n29184 = ~n29180 & ~n29181;
  assign n29185 = ~pi38  & ~n29180;
  assign n29186 = ~n42871 & ~n42872;
  assign n29187 = n29171 & ~n29186;
  assign n29188 = ~n29171 & n29186;
  assign n29189 = n29171 & ~n29187;
  assign n29190 = ~n29186 & ~n29187;
  assign n29191 = ~n29189 & ~n29190;
  assign n29192 = ~n29187 & ~n29188;
  assign n29193 = n28969 & n42873;
  assign n29194 = ~n28969 & ~n42873;
  assign n29195 = ~n29193 & ~n29194;
  assign n29196 = n2104 & n12530;
  assign n29197 = pi114  & n37758;
  assign n29198 = pi116  & n2117;
  assign n29199 = pi115  & n2119;
  assign n29200 = ~n29198 & ~n29199;
  assign n29201 = ~n29197 & ~n29199;
  assign n29202 = ~n29198 & n29201;
  assign n29203 = ~n29197 & n29200;
  assign n29204 = ~n29196 & n42874;
  assign n29205 = pi35  & ~n29204;
  assign n29206 = pi35  & ~n29205;
  assign n29207 = pi35  & n29204;
  assign n29208 = ~n29204 & ~n29205;
  assign n29209 = ~pi35  & ~n29204;
  assign n29210 = ~n42875 & ~n42876;
  assign n29211 = ~n29195 & n29210;
  assign n29212 = n29195 & ~n29210;
  assign n29213 = n29195 & ~n29212;
  assign n29214 = ~n29210 & ~n29212;
  assign n29215 = ~n29213 & ~n29214;
  assign n29216 = ~n29211 & ~n29212;
  assign n29217 = ~n42839 & ~n42877;
  assign n29218 = n42839 & n42877;
  assign n29219 = ~n29217 & ~n29218;
  assign n29220 = n28947 & ~n29218;
  assign n29221 = ~n29217 & n29220;
  assign n29222 = n28947 & n29219;
  assign n29223 = ~n28947 & ~n29219;
  assign n29224 = n28947 & ~n42878;
  assign n29225 = ~n29218 & ~n42878;
  assign n29226 = ~n29217 & n29225;
  assign n29227 = n29219 & ~n42878;
  assign n29228 = ~n29224 & ~n42879;
  assign n29229 = ~n42878 & ~n29223;
  assign n29230 = n28928 & ~n42880;
  assign n29231 = ~n28928 & n42880;
  assign n29232 = ~n29230 & ~n29231;
  assign n29233 = n28909 & ~n29231;
  assign n29234 = ~n29230 & n29233;
  assign n29235 = n28909 & n29232;
  assign n29236 = ~n29231 & ~n42881;
  assign n29237 = ~n29230 & n29236;
  assign n29238 = n29232 & ~n42881;
  assign n29239 = ~n28909 & n29232;
  assign n29240 = n28909 & ~n42881;
  assign n29241 = n28909 & ~n29232;
  assign n29242 = ~n42882 & ~n42883;
  assign n29243 = n28894 & n29242;
  assign n29244 = ~n28894 & ~n29242;
  assign n29245 = ~n29243 & ~n29244;
  assign n29246 = ~n28888 & ~n28891;
  assign n29247 = n29245 & ~n29246;
  assign n29248 = ~n29245 & n29246;
  assign po85  = ~n29247 & ~n29248;
  assign n29250 = ~n29244 & ~n29247;
  assign n29251 = ~n28927 & ~n29230;
  assign n29252 = n5576 & ~n18675;
  assign n29253 = ~n38406 & ~n29252;
  assign n29254 = pi127  & n38406;
  assign n29255 = n5576 & n18680;
  assign n29256 = ~n29254 & ~n29255;
  assign n29257 = pi127  & ~n29253;
  assign n29258 = pi23  & ~n42884;
  assign n29259 = pi23  & ~n29258;
  assign n29260 = pi23  & n42884;
  assign n29261 = ~n42884 & ~n29258;
  assign n29262 = ~pi23  & ~n42884;
  assign n29263 = ~n42885 & ~n42886;
  assign n29264 = ~n29251 & ~n29263;
  assign n29265 = n29251 & n29263;
  assign n29266 = ~n29251 & ~n29264;
  assign n29267 = ~n29263 & ~n29264;
  assign n29268 = ~n29266 & ~n29267;
  assign n29269 = ~n29264 & ~n29265;
  assign n29270 = n4492 & n15021;
  assign n29271 = pi124  & n38208;
  assign n29272 = pi126  & n4507;
  assign n29273 = pi125  & n4509;
  assign n29274 = ~n29272 & ~n29273;
  assign n29275 = ~n29271 & ~n29273;
  assign n29276 = ~n29272 & n29275;
  assign n29277 = ~n29271 & n29274;
  assign n29278 = ~n29270 & n42888;
  assign n29279 = pi26  & ~n29278;
  assign n29280 = pi26  & ~n29279;
  assign n29281 = pi26  & n29278;
  assign n29282 = ~n29278 & ~n29279;
  assign n29283 = ~pi26  & ~n29278;
  assign n29284 = ~n42889 & ~n42890;
  assign n29285 = ~n28945 & ~n42878;
  assign n29286 = n29284 & n29285;
  assign n29287 = ~n29284 & ~n29285;
  assign n29288 = ~n29286 & ~n29287;
  assign n29289 = n607 & n14961;
  assign n29290 = pi121  & n37489;
  assign n29291 = pi123  & n620;
  assign n29292 = pi122  & n622;
  assign n29293 = ~n29291 & ~n29292;
  assign n29294 = ~n29290 & ~n29292;
  assign n29295 = ~n29291 & n29294;
  assign n29296 = ~n29290 & n29293;
  assign n29297 = ~n29289 & n42891;
  assign n29298 = pi29  & ~n29297;
  assign n29299 = pi29  & ~n29298;
  assign n29300 = pi29  & n29297;
  assign n29301 = ~n29297 & ~n29298;
  assign n29302 = ~pi29  & ~n29297;
  assign n29303 = ~n42892 & ~n42893;
  assign n29304 = ~n28963 & ~n29217;
  assign n29305 = ~n29303 & ~n29304;
  assign n29306 = n29303 & n29304;
  assign n29307 = ~n29303 & ~n29305;
  assign n29308 = ~n29303 & n29304;
  assign n29309 = ~n29304 & ~n29305;
  assign n29310 = n29303 & ~n29304;
  assign n29311 = ~n42894 & ~n42895;
  assign n29312 = ~n29305 & ~n29306;
  assign n29313 = n649 & n14913;
  assign n29314 = pi118  & n37496;
  assign n29315 = pi120  & n662;
  assign n29316 = pi119  & n664;
  assign n29317 = ~n29315 & ~n29316;
  assign n29318 = ~n29314 & ~n29316;
  assign n29319 = ~n29315 & n29318;
  assign n29320 = ~n29314 & n29317;
  assign n29321 = ~n29313 & n42897;
  assign n29322 = pi32  & ~n29321;
  assign n29323 = pi32  & ~n29322;
  assign n29324 = pi32  & n29321;
  assign n29325 = ~n29321 & ~n29322;
  assign n29326 = ~pi32  & ~n29321;
  assign n29327 = ~n42898 & ~n42899;
  assign n29328 = ~n29194 & n29210;
  assign n29329 = ~n29194 & ~n29212;
  assign n29330 = ~n29193 & ~n29328;
  assign n29331 = n29327 & n42900;
  assign n29332 = ~n29327 & ~n42900;
  assign n29333 = ~n29331 & ~n29332;
  assign n29334 = n2104 & n13079;
  assign n29335 = pi115  & n37758;
  assign n29336 = pi117  & n2117;
  assign n29337 = pi116  & n2119;
  assign n29338 = ~n29336 & ~n29337;
  assign n29339 = ~n29335 & ~n29337;
  assign n29340 = ~n29336 & n29339;
  assign n29341 = ~n29335 & n29338;
  assign n29342 = ~n29334 & n42901;
  assign n29343 = pi35  & ~n29342;
  assign n29344 = pi35  & ~n29343;
  assign n29345 = pi35  & n29342;
  assign n29346 = ~n29342 & ~n29343;
  assign n29347 = ~pi35  & ~n29342;
  assign n29348 = ~n42902 & ~n42903;
  assign n29349 = n940 & n9277;
  assign n29350 = pi106  & n37541;
  assign n29351 = pi108  & n953;
  assign n29352 = pi107  & n955;
  assign n29353 = ~n29351 & ~n29352;
  assign n29354 = ~n29350 & ~n29352;
  assign n29355 = ~n29351 & n29354;
  assign n29356 = ~n29350 & n29353;
  assign n29357 = ~n29349 & n42904;
  assign n29358 = pi44  & ~n29357;
  assign n29359 = pi44  & ~n29358;
  assign n29360 = pi44  & n29357;
  assign n29361 = ~n29357 & ~n29358;
  assign n29362 = ~pi44  & ~n29357;
  assign n29363 = ~n42905 & ~n42906;
  assign n29364 = ~n29110 & ~n29116;
  assign n29365 = n785 & n8229;
  assign n29366 = pi103  & n37520;
  assign n29367 = pi105  & n787;
  assign n29368 = pi104  & n795;
  assign n29369 = ~n29367 & ~n29368;
  assign n29370 = ~n29366 & ~n29368;
  assign n29371 = ~n29367 & n29370;
  assign n29372 = ~n29366 & n29369;
  assign n29373 = ~n29365 & n42907;
  assign n29374 = pi47  & ~n29373;
  assign n29375 = pi47  & ~n29374;
  assign n29376 = pi47  & n29373;
  assign n29377 = ~n29373 & ~n29374;
  assign n29378 = ~pi47  & ~n29373;
  assign n29379 = ~n42908 & ~n42909;
  assign n29380 = ~n29090 & ~n29108;
  assign n29381 = n1971 & n5578;
  assign n29382 = pi97  & n37864;
  assign n29383 = pi99  & n1973;
  assign n29384 = pi98  & n1981;
  assign n29385 = ~n29383 & ~n29384;
  assign n29386 = ~n29382 & ~n29384;
  assign n29387 = ~n29383 & n29386;
  assign n29388 = ~n29382 & n29385;
  assign n29389 = ~n29381 & n42910;
  assign n29390 = pi53  & ~n29389;
  assign n29391 = pi53  & ~n29390;
  assign n29392 = pi53  & n29389;
  assign n29393 = ~n29389 & ~n29390;
  assign n29394 = ~pi53  & ~n29389;
  assign n29395 = ~n42911 & ~n42912;
  assign n29396 = ~n29032 & ~n29035;
  assign n29397 = ~n29012 & ~n29029;
  assign n29398 = pi87  & ~n40814;
  assign n29399 = pi86  & n18285;
  assign n29400 = ~n29398 & ~n29399;
  assign n29401 = ~n29010 & n29400;
  assign n29402 = n29010 & ~n29400;
  assign n29403 = ~n29401 & ~n29402;
  assign n29404 = n3566 & n12674;
  assign n29405 = pi88  & n40107;
  assign n29406 = pi90  & n12676;
  assign n29407 = pi89  & n12684;
  assign n29408 = ~n29406 & ~n29407;
  assign n29409 = ~n29405 & ~n29407;
  assign n29410 = ~n29406 & n29409;
  assign n29411 = ~n29405 & n29408;
  assign n29412 = ~n12674 & n42913;
  assign n29413 = ~n3566 & n42913;
  assign n29414 = ~n29412 & ~n29413;
  assign n29415 = ~n29404 & n42913;
  assign n29416 = pi62  & ~n42914;
  assign n29417 = ~pi62  & n42914;
  assign n29418 = ~n29416 & ~n29417;
  assign n29419 = n29403 & ~n29418;
  assign n29420 = ~n29403 & n29418;
  assign n29421 = ~n29419 & ~n29420;
  assign n29422 = ~n29397 & n29421;
  assign n29423 = n29397 & ~n29421;
  assign n29424 = ~n29422 & ~n29423;
  assign n29425 = n4544 & n7882;
  assign n29426 = pi91  & n39128;
  assign n29427 = pi93  & n7884;
  assign n29428 = pi92  & n7892;
  assign n29429 = ~n29427 & ~n29428;
  assign n29430 = ~n29426 & ~n29428;
  assign n29431 = ~n29427 & n29430;
  assign n29432 = ~n29426 & n29429;
  assign n29433 = ~n29425 & n42915;
  assign n29434 = pi59  & ~n29433;
  assign n29435 = pi59  & ~n29434;
  assign n29436 = pi59  & n29433;
  assign n29437 = ~n29433 & ~n29434;
  assign n29438 = ~pi59  & ~n29433;
  assign n29439 = ~n42916 & ~n42917;
  assign n29440 = n29424 & ~n29439;
  assign n29441 = ~n29424 & n29439;
  assign n29442 = n29424 & ~n29440;
  assign n29443 = ~n29439 & ~n29440;
  assign n29444 = ~n29442 & ~n29443;
  assign n29445 = ~n29440 & ~n29441;
  assign n29446 = n29396 & n42918;
  assign n29447 = ~n29396 & ~n42918;
  assign n29448 = ~n29446 & ~n29447;
  assign n29449 = n4312 & n5281;
  assign n29450 = pi94  & n38376;
  assign n29451 = pi96  & n4314;
  assign n29452 = pi95  & n4322;
  assign n29453 = ~n29451 & ~n29452;
  assign n29454 = ~n29450 & ~n29452;
  assign n29455 = ~n29451 & n29454;
  assign n29456 = ~n29450 & n29453;
  assign n29457 = ~n29449 & n42919;
  assign n29458 = pi56  & ~n29457;
  assign n29459 = pi56  & ~n29458;
  assign n29460 = pi56  & n29457;
  assign n29461 = ~n29457 & ~n29458;
  assign n29462 = ~pi56  & ~n29457;
  assign n29463 = ~n42920 & ~n42921;
  assign n29464 = ~n29448 & n29463;
  assign n29465 = n29448 & ~n29463;
  assign n29466 = ~n29464 & ~n29465;
  assign n29467 = ~n29038 & n29055;
  assign n29468 = ~n29038 & ~n29056;
  assign n29469 = ~n29039 & ~n29467;
  assign n29470 = n29466 & ~n42922;
  assign n29471 = ~n29466 & n42922;
  assign n29472 = ~n29470 & ~n29471;
  assign n29473 = ~n29395 & n29472;
  assign n29474 = n29395 & ~n29472;
  assign n29475 = ~n29473 & ~n29474;
  assign n29476 = ~n29063 & n29079;
  assign n29477 = ~n29063 & ~n29081;
  assign n29478 = ~n29062 & ~n29476;
  assign n29479 = n29475 & ~n42923;
  assign n29480 = ~n29475 & n42923;
  assign n29481 = ~n29479 & ~n29480;
  assign n29482 = n894 & n6819;
  assign n29483 = pi100  & n37580;
  assign n29484 = pi102  & n896;
  assign n29485 = pi101  & n904;
  assign n29486 = ~n29484 & ~n29485;
  assign n29487 = ~n29483 & ~n29485;
  assign n29488 = ~n29484 & n29487;
  assign n29489 = ~n29483 & n29486;
  assign n29490 = ~n29482 & n42924;
  assign n29491 = pi50  & ~n29490;
  assign n29492 = pi50  & ~n29491;
  assign n29493 = pi50  & n29490;
  assign n29494 = ~n29490 & ~n29491;
  assign n29495 = ~pi50  & ~n29490;
  assign n29496 = ~n42925 & ~n42926;
  assign n29497 = n29481 & ~n29496;
  assign n29498 = ~n29481 & n29496;
  assign n29499 = n29481 & ~n29497;
  assign n29500 = ~n29496 & ~n29497;
  assign n29501 = ~n29499 & ~n29500;
  assign n29502 = ~n29497 & ~n29498;
  assign n29503 = ~n29380 & ~n42927;
  assign n29504 = n29380 & n42927;
  assign n29505 = ~n42927 & ~n29503;
  assign n29506 = ~n29380 & ~n29503;
  assign n29507 = ~n29505 & ~n29506;
  assign n29508 = ~n29503 & ~n29504;
  assign n29509 = n29379 & ~n42928;
  assign n29510 = ~n29379 & n42928;
  assign n29511 = ~n29379 & ~n42928;
  assign n29512 = n29379 & n42928;
  assign n29513 = ~n29511 & ~n29512;
  assign n29514 = ~n29509 & ~n29510;
  assign n29515 = ~n29364 & n42929;
  assign n29516 = n29364 & ~n42929;
  assign n29517 = ~n29515 & ~n29516;
  assign n29518 = ~n29363 & n29517;
  assign n29519 = n29363 & ~n29517;
  assign n29520 = ~n29518 & ~n29519;
  assign n29521 = ~n29121 & n29138;
  assign n29522 = ~n29121 & ~n29139;
  assign n29523 = ~n29122 & ~n29521;
  assign n29524 = n29520 & ~n42930;
  assign n29525 = ~n29520 & n42930;
  assign n29526 = ~n29524 & ~n29525;
  assign n29527 = n565 & n733;
  assign n29528 = pi109  & n37510;
  assign n29529 = pi111  & n746;
  assign n29530 = pi110  & n748;
  assign n29531 = ~n29529 & ~n29530;
  assign n29532 = ~n29528 & ~n29530;
  assign n29533 = ~n29529 & n29532;
  assign n29534 = ~n29528 & n29531;
  assign n29535 = ~n29527 & n42931;
  assign n29536 = pi41  & ~n29535;
  assign n29537 = pi41  & ~n29536;
  assign n29538 = pi41  & n29535;
  assign n29539 = ~n29535 & ~n29536;
  assign n29540 = ~pi41  & ~n29535;
  assign n29541 = ~n42932 & ~n42933;
  assign n29542 = n29526 & ~n29541;
  assign n29543 = ~n29526 & n29541;
  assign n29544 = n29526 & ~n29542;
  assign n29545 = ~n29541 & ~n29542;
  assign n29546 = ~n29544 & ~n29545;
  assign n29547 = ~n29542 & ~n29543;
  assign n29548 = ~n29146 & n29162;
  assign n29549 = ~n29146 & ~n29164;
  assign n29550 = ~n29145 & ~n29548;
  assign n29551 = n42934 & n42935;
  assign n29552 = ~n42934 & ~n42935;
  assign n29553 = ~n29551 & ~n29552;
  assign n29554 = n691 & n11258;
  assign n29555 = pi112  & n37503;
  assign n29556 = pi114  & n704;
  assign n29557 = pi113  & n706;
  assign n29558 = ~n29556 & ~n29557;
  assign n29559 = ~n29555 & ~n29557;
  assign n29560 = ~n29556 & n29559;
  assign n29561 = ~n29555 & n29558;
  assign n29562 = ~n29554 & n42936;
  assign n29563 = pi38  & ~n29562;
  assign n29564 = pi38  & ~n29563;
  assign n29565 = pi38  & n29562;
  assign n29566 = ~n29562 & ~n29563;
  assign n29567 = ~pi38  & ~n29562;
  assign n29568 = ~n42937 & ~n42938;
  assign n29569 = ~n29553 & n29568;
  assign n29570 = n29553 & ~n29568;
  assign n29571 = ~n29569 & ~n29570;
  assign n29572 = ~n29170 & n29186;
  assign n29573 = ~n29170 & ~n29187;
  assign n29574 = ~n29169 & ~n29572;
  assign n29575 = n29571 & ~n42939;
  assign n29576 = ~n29571 & n42939;
  assign n29577 = ~n42939 & ~n29575;
  assign n29578 = n29571 & ~n29575;
  assign n29579 = ~n29577 & ~n29578;
  assign n29580 = ~n29575 & ~n29576;
  assign n29581 = n29348 & n42940;
  assign n29582 = ~n29348 & ~n42940;
  assign n29583 = ~n29348 & ~n29582;
  assign n29584 = ~n42940 & ~n29582;
  assign n29585 = ~n29583 & ~n29584;
  assign n29586 = ~n29581 & ~n29582;
  assign n29587 = n29333 & ~n42941;
  assign n29588 = ~n29333 & n42941;
  assign n29589 = n29333 & ~n29587;
  assign n29590 = ~n42941 & ~n29587;
  assign n29591 = ~n29589 & ~n29590;
  assign n29592 = ~n29587 & ~n29588;
  assign n29593 = ~n42896 & ~n42942;
  assign n29594 = n42896 & n42942;
  assign n29595 = ~n42896 & n42942;
  assign n29596 = n42896 & ~n42942;
  assign n29597 = ~n29595 & ~n29596;
  assign n29598 = ~n29593 & ~n29594;
  assign n29599 = n29288 & ~n42943;
  assign n29600 = ~n29288 & n42943;
  assign n29601 = n29288 & ~n29599;
  assign n29602 = ~n42943 & ~n29599;
  assign n29603 = ~n29601 & ~n29602;
  assign n29604 = ~n29599 & ~n29600;
  assign n29605 = ~n42887 & ~n42944;
  assign n29606 = n42887 & n42944;
  assign n29607 = ~n42887 & n42944;
  assign n29608 = n42887 & ~n42944;
  assign n29609 = ~n29607 & ~n29608;
  assign n29610 = ~n29605 & ~n29606;
  assign n29611 = ~n28907 & ~n29232;
  assign n29612 = ~n28907 & ~n42881;
  assign n29613 = ~n28908 & ~n29611;
  assign n29614 = ~n42945 & ~n42946;
  assign n29615 = n42945 & n42946;
  assign n29616 = ~n42946 & ~n29614;
  assign n29617 = ~n42945 & ~n29614;
  assign n29618 = ~n29616 & ~n29617;
  assign n29619 = ~n29614 & ~n29615;
  assign n29620 = ~n29250 & ~n42947;
  assign n29621 = n29250 & ~n29617;
  assign n29622 = ~n29616 & n29621;
  assign n29623 = n29250 & n42947;
  assign po86  = ~n29620 & ~n42948;
  assign n29625 = ~n29614 & ~n29620;
  assign n29626 = ~n29264 & ~n29605;
  assign n29627 = ~n29287 & ~n29599;
  assign n29628 = n4492 & n40885;
  assign n29629 = pi125  & n38208;
  assign n29630 = pi127  & n4507;
  assign n29631 = pi126  & n4509;
  assign n29632 = ~n29630 & ~n29631;
  assign n29633 = ~n29629 & ~n29631;
  assign n29634 = ~n29630 & n29633;
  assign n29635 = ~n29629 & n29632;
  assign n29636 = ~n29628 & n42949;
  assign n29637 = pi26  & ~n29636;
  assign n29638 = pi26  & ~n29637;
  assign n29639 = pi26  & n29636;
  assign n29640 = ~n29636 & ~n29637;
  assign n29641 = ~pi26  & ~n29636;
  assign n29642 = ~n42950 & ~n42951;
  assign n29643 = ~n29627 & ~n29642;
  assign n29644 = n29627 & n29642;
  assign n29645 = ~n29627 & ~n29643;
  assign n29646 = ~n29627 & n29642;
  assign n29647 = ~n29642 & ~n29643;
  assign n29648 = n29627 & ~n29642;
  assign n29649 = ~n42952 & ~n42953;
  assign n29650 = ~n29643 & ~n29644;
  assign n29651 = n649 & n15091;
  assign n29652 = pi119  & n37496;
  assign n29653 = pi121  & n662;
  assign n29654 = pi120  & n664;
  assign n29655 = ~n29653 & ~n29654;
  assign n29656 = ~n29652 & ~n29654;
  assign n29657 = ~n29653 & n29656;
  assign n29658 = ~n29652 & n29655;
  assign n29659 = ~n29651 & n42955;
  assign n29660 = pi32  & ~n29659;
  assign n29661 = pi32  & ~n29660;
  assign n29662 = pi32  & n29659;
  assign n29663 = ~n29659 & ~n29660;
  assign n29664 = ~pi32  & ~n29659;
  assign n29665 = ~n42956 & ~n42957;
  assign n29666 = ~n29332 & n42941;
  assign n29667 = ~n29332 & ~n29587;
  assign n29668 = ~n29331 & ~n29666;
  assign n29669 = n29665 & n42958;
  assign n29670 = ~n29665 & ~n42958;
  assign n29671 = ~n29669 & ~n29670;
  assign n29672 = n2104 & n13057;
  assign n29673 = pi116  & n37758;
  assign n29674 = pi118  & n2117;
  assign n29675 = pi117  & n2119;
  assign n29676 = ~n29674 & ~n29675;
  assign n29677 = ~n29673 & ~n29675;
  assign n29678 = ~n29674 & n29677;
  assign n29679 = ~n29673 & n29676;
  assign n29680 = ~n29672 & n42959;
  assign n29681 = pi35  & ~n29680;
  assign n29682 = pi35  & ~n29681;
  assign n29683 = pi35  & n29680;
  assign n29684 = ~n29680 & ~n29681;
  assign n29685 = ~pi35  & ~n29680;
  assign n29686 = ~n42960 & ~n42961;
  assign n29687 = ~n29552 & ~n29570;
  assign n29688 = ~n29515 & ~n29518;
  assign n29689 = n940 & n9701;
  assign n29690 = pi107  & n37541;
  assign n29691 = pi109  & n953;
  assign n29692 = pi108  & n955;
  assign n29693 = ~n29691 & ~n29692;
  assign n29694 = ~n29690 & ~n29692;
  assign n29695 = ~n29691 & n29694;
  assign n29696 = ~n29690 & n29693;
  assign n29697 = ~n29689 & n42962;
  assign n29698 = pi44  & ~n29697;
  assign n29699 = pi44  & ~n29698;
  assign n29700 = pi44  & n29697;
  assign n29701 = ~n29697 & ~n29698;
  assign n29702 = ~pi44  & ~n29697;
  assign n29703 = ~n42963 & ~n42964;
  assign n29704 = ~n29470 & ~n29473;
  assign n29705 = n4524 & n7882;
  assign n29706 = pi92  & n39128;
  assign n29707 = pi94  & n7884;
  assign n29708 = pi93  & n7892;
  assign n29709 = ~n29707 & ~n29708;
  assign n29710 = ~n29706 & ~n29708;
  assign n29711 = ~n29707 & n29710;
  assign n29712 = ~n29706 & n29709;
  assign n29713 = ~n29705 & n42965;
  assign n29714 = pi59  & ~n29713;
  assign n29715 = pi59  & ~n29714;
  assign n29716 = pi59  & n29713;
  assign n29717 = ~n29713 & ~n29714;
  assign n29718 = ~pi59  & ~n29713;
  assign n29719 = ~n42966 & ~n42967;
  assign n29720 = ~n29401 & ~n29419;
  assign n29721 = pi88  & ~n40814;
  assign n29722 = pi87  & n18285;
  assign n29723 = ~n29721 & ~n29722;
  assign n29724 = ~pi23  & ~n29723;
  assign n29725 = pi23  & n29723;
  assign n29726 = ~n29724 & ~n29725;
  assign n29727 = ~n29400 & n29726;
  assign n29728 = n29400 & ~n29726;
  assign n29729 = ~n29727 & ~n29728;
  assign n29730 = n594 & n12674;
  assign n29731 = pi89  & n40107;
  assign n29732 = pi91  & n12676;
  assign n29733 = pi90  & n12684;
  assign n29734 = ~n29732 & ~n29733;
  assign n29735 = ~n29731 & ~n29733;
  assign n29736 = ~n29732 & n29735;
  assign n29737 = ~n29731 & n29734;
  assign n29738 = ~n29730 & n42968;
  assign n29739 = pi62  & ~n29738;
  assign n29740 = pi62  & ~n29739;
  assign n29741 = pi62  & n29738;
  assign n29742 = ~n29738 & ~n29739;
  assign n29743 = ~pi62  & ~n29738;
  assign n29744 = ~n42969 & ~n42970;
  assign n29745 = n29729 & ~n29744;
  assign n29746 = ~n29729 & n29744;
  assign n29747 = n29729 & ~n29745;
  assign n29748 = n29729 & n29744;
  assign n29749 = ~n29744 & ~n29745;
  assign n29750 = ~n29729 & ~n29744;
  assign n29751 = ~n42971 & ~n42972;
  assign n29752 = ~n29745 & ~n29746;
  assign n29753 = ~n29720 & ~n42973;
  assign n29754 = n29720 & n42973;
  assign n29755 = ~n29720 & n42973;
  assign n29756 = n29720 & ~n42973;
  assign n29757 = ~n29755 & ~n29756;
  assign n29758 = ~n29753 & ~n29754;
  assign n29759 = ~n29719 & ~n42974;
  assign n29760 = n29719 & n42974;
  assign n29761 = ~n29759 & ~n29760;
  assign n29762 = ~n29422 & n29439;
  assign n29763 = ~n29422 & ~n29440;
  assign n29764 = ~n29423 & ~n29762;
  assign n29765 = ~n29761 & n42975;
  assign n29766 = n29761 & ~n42975;
  assign n29767 = ~n29765 & ~n29766;
  assign n29768 = n4312 & n5630;
  assign n29769 = pi95  & n38376;
  assign n29770 = pi97  & n4314;
  assign n29771 = pi96  & n4322;
  assign n29772 = ~n29770 & ~n29771;
  assign n29773 = ~n29769 & ~n29771;
  assign n29774 = ~n29770 & n29773;
  assign n29775 = ~n29769 & n29772;
  assign n29776 = ~n29768 & n42976;
  assign n29777 = pi56  & ~n29776;
  assign n29778 = pi56  & ~n29777;
  assign n29779 = pi56  & n29776;
  assign n29780 = ~n29776 & ~n29777;
  assign n29781 = ~pi56  & ~n29776;
  assign n29782 = ~n42977 & ~n42978;
  assign n29783 = ~n29447 & ~n29465;
  assign n29784 = ~n29782 & ~n29783;
  assign n29785 = n29782 & n29783;
  assign n29786 = ~n29784 & ~n29785;
  assign n29787 = n29767 & n29786;
  assign n29788 = ~n29767 & ~n29786;
  assign n29789 = ~n29787 & ~n29788;
  assign n29790 = n1971 & n6474;
  assign n29791 = pi98  & n37864;
  assign n29792 = pi100  & n1973;
  assign n29793 = pi99  & n1981;
  assign n29794 = ~n29792 & ~n29793;
  assign n29795 = ~n29791 & ~n29793;
  assign n29796 = ~n29792 & n29795;
  assign n29797 = ~n29791 & n29794;
  assign n29798 = ~n29790 & n42979;
  assign n29799 = pi53  & ~n29798;
  assign n29800 = pi53  & ~n29799;
  assign n29801 = pi53  & n29798;
  assign n29802 = ~n29798 & ~n29799;
  assign n29803 = ~pi53  & ~n29798;
  assign n29804 = ~n42980 & ~n42981;
  assign n29805 = n29789 & ~n29804;
  assign n29806 = ~n29789 & n29804;
  assign n29807 = n29789 & ~n29805;
  assign n29808 = n29789 & n29804;
  assign n29809 = ~n29804 & ~n29805;
  assign n29810 = ~n29789 & ~n29804;
  assign n29811 = ~n42982 & ~n42983;
  assign n29812 = ~n29805 & ~n29806;
  assign n29813 = n29704 & n42984;
  assign n29814 = ~n29704 & ~n42984;
  assign n29815 = ~n29813 & ~n29814;
  assign n29816 = n894 & n6787;
  assign n29817 = pi101  & n37580;
  assign n29818 = pi103  & n896;
  assign n29819 = pi102  & n904;
  assign n29820 = ~n29818 & ~n29819;
  assign n29821 = ~n29817 & ~n29819;
  assign n29822 = ~n29818 & n29821;
  assign n29823 = ~n29817 & n29820;
  assign n29824 = ~n29816 & n42985;
  assign n29825 = pi50  & ~n29824;
  assign n29826 = pi50  & ~n29825;
  assign n29827 = pi50  & n29824;
  assign n29828 = ~n29824 & ~n29825;
  assign n29829 = ~pi50  & ~n29824;
  assign n29830 = ~n42986 & ~n42987;
  assign n29831 = n29815 & ~n29830;
  assign n29832 = ~n29815 & n29830;
  assign n29833 = n29815 & ~n29831;
  assign n29834 = n29815 & n29830;
  assign n29835 = ~n29830 & ~n29831;
  assign n29836 = ~n29815 & ~n29830;
  assign n29837 = ~n42988 & ~n42989;
  assign n29838 = ~n29831 & ~n29832;
  assign n29839 = ~n29479 & n29496;
  assign n29840 = ~n29479 & ~n29497;
  assign n29841 = ~n29480 & ~n29839;
  assign n29842 = n42990 & n42991;
  assign n29843 = ~n42990 & ~n42991;
  assign n29844 = ~n29842 & ~n29843;
  assign n29845 = n785 & n8209;
  assign n29846 = pi104  & n37520;
  assign n29847 = pi106  & n787;
  assign n29848 = pi105  & n795;
  assign n29849 = ~n29847 & ~n29848;
  assign n29850 = ~n29846 & ~n29848;
  assign n29851 = ~n29847 & n29850;
  assign n29852 = ~n29846 & n29849;
  assign n29853 = ~n29845 & n42992;
  assign n29854 = pi47  & ~n29853;
  assign n29855 = pi47  & ~n29854;
  assign n29856 = pi47  & n29853;
  assign n29857 = ~n29853 & ~n29854;
  assign n29858 = ~pi47  & ~n29853;
  assign n29859 = ~n42993 & ~n42994;
  assign n29860 = n29844 & ~n29859;
  assign n29861 = ~n29844 & n29859;
  assign n29862 = n29844 & ~n29860;
  assign n29863 = n29844 & n29859;
  assign n29864 = ~n29859 & ~n29860;
  assign n29865 = ~n29844 & ~n29859;
  assign n29866 = ~n42995 & ~n42996;
  assign n29867 = ~n29860 & ~n29861;
  assign n29868 = n29379 & ~n29503;
  assign n29869 = ~n29503 & ~n29511;
  assign n29870 = ~n29504 & ~n29868;
  assign n29871 = ~n42997 & ~n42998;
  assign n29872 = n42997 & n42998;
  assign n29873 = n42997 & ~n42998;
  assign n29874 = ~n42997 & n42998;
  assign n29875 = ~n29873 & ~n29874;
  assign n29876 = ~n29871 & ~n29872;
  assign n29877 = ~n29703 & ~n42999;
  assign n29878 = n29703 & n42999;
  assign n29879 = ~n29877 & ~n29878;
  assign n29880 = n29688 & ~n29879;
  assign n29881 = ~n29688 & n29879;
  assign n29882 = ~n29880 & ~n29881;
  assign n29883 = n733 & n10844;
  assign n29884 = pi110  & n37510;
  assign n29885 = pi112  & n746;
  assign n29886 = pi111  & n748;
  assign n29887 = ~n29885 & ~n29886;
  assign n29888 = ~n29884 & ~n29886;
  assign n29889 = ~n29885 & n29888;
  assign n29890 = ~n29884 & n29887;
  assign n29891 = ~n29883 & n43000;
  assign n29892 = pi41  & ~n29891;
  assign n29893 = pi41  & ~n29892;
  assign n29894 = pi41  & n29891;
  assign n29895 = ~n29891 & ~n29892;
  assign n29896 = ~pi41  & ~n29891;
  assign n29897 = ~n43001 & ~n43002;
  assign n29898 = n29882 & ~n29897;
  assign n29899 = ~n29882 & n29897;
  assign n29900 = n29882 & ~n29898;
  assign n29901 = n29882 & n29897;
  assign n29902 = ~n29897 & ~n29898;
  assign n29903 = ~n29882 & ~n29897;
  assign n29904 = ~n43003 & ~n43004;
  assign n29905 = ~n29898 & ~n29899;
  assign n29906 = ~n29524 & n29541;
  assign n29907 = ~n29524 & ~n29542;
  assign n29908 = ~n29525 & ~n29906;
  assign n29909 = n43005 & n43006;
  assign n29910 = ~n43005 & ~n43006;
  assign n29911 = ~n29909 & ~n29910;
  assign n29912 = n523 & n691;
  assign n29913 = pi113  & n37503;
  assign n29914 = pi115  & n704;
  assign n29915 = pi114  & n706;
  assign n29916 = ~n29914 & ~n29915;
  assign n29917 = ~n29913 & ~n29915;
  assign n29918 = ~n29914 & n29917;
  assign n29919 = ~n29913 & n29916;
  assign n29920 = ~n29912 & n43007;
  assign n29921 = pi38  & ~n29920;
  assign n29922 = pi38  & ~n29921;
  assign n29923 = pi38  & n29920;
  assign n29924 = ~n29920 & ~n29921;
  assign n29925 = ~pi38  & ~n29920;
  assign n29926 = ~n43008 & ~n43009;
  assign n29927 = n29911 & ~n29926;
  assign n29928 = ~n29911 & n29926;
  assign n29929 = ~n29927 & ~n29928;
  assign n29930 = n29687 & ~n29929;
  assign n29931 = ~n29687 & ~n29928;
  assign n29932 = ~n29927 & n29931;
  assign n29933 = ~n29687 & ~n29927;
  assign n29934 = ~n29928 & n29933;
  assign n29935 = ~n29687 & n29929;
  assign n29936 = ~n29687 & ~n43010;
  assign n29937 = ~n29687 & ~n29929;
  assign n29938 = n29687 & ~n29927;
  assign n29939 = ~n29927 & ~n43010;
  assign n29940 = ~n29928 & ~n29938;
  assign n29941 = ~n29928 & n43012;
  assign n29942 = n29687 & n29929;
  assign n29943 = ~n43011 & ~n43013;
  assign n29944 = ~n29930 & ~n43010;
  assign n29945 = n29686 & n43014;
  assign n29946 = ~n29686 & ~n43014;
  assign n29947 = ~n29945 & ~n29946;
  assign n29948 = n29348 & ~n29575;
  assign n29949 = ~n29575 & ~n29582;
  assign n29950 = ~n29576 & ~n29948;
  assign n29951 = n29947 & ~n43015;
  assign n29952 = ~n29947 & n43015;
  assign n29953 = ~n29951 & ~n29952;
  assign n29954 = n29671 & n29953;
  assign n29955 = ~n29671 & ~n29953;
  assign n29956 = ~n29954 & ~n29955;
  assign n29957 = ~n29305 & ~n29593;
  assign n29958 = n607 & n15111;
  assign n29959 = pi122  & n37489;
  assign n29960 = pi124  & n620;
  assign n29961 = pi123  & n622;
  assign n29962 = ~n29960 & ~n29961;
  assign n29963 = ~n29959 & ~n29961;
  assign n29964 = ~n29960 & n29963;
  assign n29965 = ~n29959 & n29962;
  assign n29966 = ~n29958 & n43016;
  assign n29967 = pi29  & ~n29966;
  assign n29968 = pi29  & ~n29967;
  assign n29969 = pi29  & n29966;
  assign n29970 = ~n29966 & ~n29967;
  assign n29971 = ~pi29  & ~n29966;
  assign n29972 = ~n43017 & ~n43018;
  assign n29973 = ~n29957 & ~n29972;
  assign n29974 = n29957 & n29972;
  assign n29975 = ~n29957 & n29972;
  assign n29976 = n29957 & ~n29972;
  assign n29977 = ~n29975 & ~n29976;
  assign n29978 = ~n29973 & ~n29974;
  assign n29979 = ~n29955 & ~n43019;
  assign n29980 = ~n29954 & n29979;
  assign n29981 = n29956 & ~n43019;
  assign n29982 = ~n29956 & n43019;
  assign n29983 = ~n43019 & ~n43020;
  assign n29984 = ~n29956 & ~n43019;
  assign n29985 = n29956 & ~n43020;
  assign n29986 = ~n29955 & ~n43020;
  assign n29987 = ~n29954 & n29986;
  assign n29988 = n29956 & n43019;
  assign n29989 = ~n43021 & ~n43022;
  assign n29990 = ~n43020 & ~n29982;
  assign n29991 = ~n42954 & ~n43023;
  assign n29992 = n42954 & n43023;
  assign n29993 = ~n42954 & n43023;
  assign n29994 = n42954 & ~n43023;
  assign n29995 = ~n29993 & ~n29994;
  assign n29996 = ~n29991 & ~n29992;
  assign n29997 = ~n29626 & ~n43024;
  assign n29998 = n29626 & n43024;
  assign n29999 = ~n29626 & ~n29997;
  assign n30000 = ~n43024 & ~n29997;
  assign n30001 = ~n29999 & ~n30000;
  assign n30002 = ~n29997 & ~n29998;
  assign n30003 = ~n29625 & ~n43025;
  assign n30004 = n29625 & ~n30000;
  assign n30005 = ~n29999 & n30004;
  assign n30006 = n29625 & n43025;
  assign po87  = ~n30003 & ~n43026;
  assign n30008 = ~n29997 & ~n30003;
  assign n30009 = ~n29643 & ~n29991;
  assign n30010 = ~n29946 & ~n29951;
  assign n30011 = n649 & n15049;
  assign n30012 = pi120  & n37496;
  assign n30013 = pi122  & n662;
  assign n30014 = pi121  & n664;
  assign n30015 = ~n30013 & ~n30014;
  assign n30016 = ~n30012 & ~n30014;
  assign n30017 = ~n30013 & n30016;
  assign n30018 = ~n30012 & n30015;
  assign n30019 = ~n649 & n43027;
  assign n30020 = ~n15049 & n43027;
  assign n30021 = ~n30019 & ~n30020;
  assign n30022 = ~n30011 & n43027;
  assign n30023 = pi32  & ~n43028;
  assign n30024 = ~pi32  & n43028;
  assign n30025 = ~n30023 & ~n30024;
  assign n30026 = ~n30010 & ~n30025;
  assign n30027 = n30010 & n30025;
  assign n30028 = ~n30026 & ~n30027;
  assign n30029 = n2104 & n13027;
  assign n30030 = pi117  & n37758;
  assign n30031 = pi119  & n2117;
  assign n30032 = pi118  & n2119;
  assign n30033 = ~n30031 & ~n30032;
  assign n30034 = ~n30030 & ~n30032;
  assign n30035 = ~n30031 & n30034;
  assign n30036 = ~n30030 & n30033;
  assign n30037 = ~n30029 & n43029;
  assign n30038 = pi35  & ~n30037;
  assign n30039 = pi35  & ~n30038;
  assign n30040 = pi35  & n30037;
  assign n30041 = ~n30037 & ~n30038;
  assign n30042 = ~pi35  & ~n30037;
  assign n30043 = ~n43030 & ~n43031;
  assign n30044 = ~n29898 & ~n29910;
  assign n30045 = ~n29877 & ~n29881;
  assign n30046 = ~n29860 & ~n29871;
  assign n30047 = ~n29831 & ~n29843;
  assign n30048 = n894 & n8136;
  assign n30049 = pi102  & n37580;
  assign n30050 = pi104  & n896;
  assign n30051 = pi103  & n904;
  assign n30052 = ~n30050 & ~n30051;
  assign n30053 = ~n30049 & ~n30051;
  assign n30054 = ~n30050 & n30053;
  assign n30055 = ~n30049 & n30052;
  assign n30056 = ~n30048 & n43032;
  assign n30057 = pi50  & ~n30056;
  assign n30058 = pi50  & ~n30057;
  assign n30059 = pi50  & n30056;
  assign n30060 = ~n30056 & ~n30057;
  assign n30061 = ~pi50  & ~n30056;
  assign n30062 = ~n43033 & ~n43034;
  assign n30063 = ~n29805 & ~n29814;
  assign n30064 = ~n29784 & ~n29787;
  assign n30065 = ~n29759 & ~n29766;
  assign n30066 = ~n29745 & ~n29753;
  assign n30067 = ~n29724 & ~n29727;
  assign n30068 = pi89  & ~n40814;
  assign n30069 = pi88  & n18285;
  assign n30070 = ~n30068 & ~n30069;
  assign n30071 = n30067 & ~n30070;
  assign n30072 = ~n30067 & n30070;
  assign n30073 = ~n30071 & ~n30072;
  assign n30074 = n4453 & n12674;
  assign n30075 = pi90  & n40107;
  assign n30076 = pi92  & n12676;
  assign n30077 = pi91  & n12684;
  assign n30078 = ~n30076 & ~n30077;
  assign n30079 = ~n30075 & ~n30077;
  assign n30080 = ~n30076 & n30079;
  assign n30081 = ~n30075 & n30078;
  assign n30082 = ~n12674 & n43035;
  assign n30083 = ~n4453 & n43035;
  assign n30084 = ~n30082 & ~n30083;
  assign n30085 = ~n30074 & n43035;
  assign n30086 = pi62  & ~n43036;
  assign n30087 = ~pi62  & n43036;
  assign n30088 = ~n30086 & ~n30087;
  assign n30089 = n30073 & ~n30088;
  assign n30090 = ~n30073 & n30088;
  assign n30091 = ~n30089 & ~n30090;
  assign n30092 = ~n30066 & n30091;
  assign n30093 = n30066 & ~n30091;
  assign n30094 = ~n30092 & ~n30093;
  assign n30095 = n4494 & n7882;
  assign n30096 = pi93  & n39128;
  assign n30097 = pi95  & n7884;
  assign n30098 = pi94  & n7892;
  assign n30099 = ~n30097 & ~n30098;
  assign n30100 = ~n30096 & ~n30098;
  assign n30101 = ~n30097 & n30100;
  assign n30102 = ~n30096 & n30099;
  assign n30103 = ~n30095 & n43037;
  assign n30104 = pi59  & ~n30103;
  assign n30105 = pi59  & ~n30104;
  assign n30106 = pi59  & n30103;
  assign n30107 = ~n30103 & ~n30104;
  assign n30108 = ~pi59  & ~n30103;
  assign n30109 = ~n43038 & ~n43039;
  assign n30110 = n30094 & ~n30109;
  assign n30111 = ~n30094 & n30109;
  assign n30112 = n30094 & ~n30110;
  assign n30113 = ~n30109 & ~n30110;
  assign n30114 = ~n30112 & ~n30113;
  assign n30115 = ~n30110 & ~n30111;
  assign n30116 = n30065 & n43040;
  assign n30117 = ~n30065 & ~n43040;
  assign n30118 = ~n30116 & ~n30117;
  assign n30119 = n4312 & n5610;
  assign n30120 = pi96  & n38376;
  assign n30121 = pi98  & n4314;
  assign n30122 = pi97  & n4322;
  assign n30123 = ~n30121 & ~n30122;
  assign n30124 = ~n30120 & ~n30122;
  assign n30125 = ~n30121 & n30124;
  assign n30126 = ~n30120 & n30123;
  assign n30127 = ~n30119 & n43041;
  assign n30128 = pi56  & ~n30127;
  assign n30129 = pi56  & ~n30128;
  assign n30130 = pi56  & n30127;
  assign n30131 = ~n30127 & ~n30128;
  assign n30132 = ~pi56  & ~n30127;
  assign n30133 = ~n43042 & ~n43043;
  assign n30134 = ~n30118 & n30133;
  assign n30135 = n30118 & ~n30133;
  assign n30136 = n30118 & ~n30135;
  assign n30137 = ~n30133 & ~n30135;
  assign n30138 = ~n30136 & ~n30137;
  assign n30139 = ~n30134 & ~n30135;
  assign n30140 = n30064 & n43044;
  assign n30141 = ~n30064 & ~n43044;
  assign n30142 = ~n30140 & ~n30141;
  assign n30143 = n1971 & n6839;
  assign n30144 = pi99  & n37864;
  assign n30145 = pi101  & n1973;
  assign n30146 = pi100  & n1981;
  assign n30147 = ~n30145 & ~n30146;
  assign n30148 = ~n30144 & ~n30146;
  assign n30149 = ~n30145 & n30148;
  assign n30150 = ~n30144 & n30147;
  assign n30151 = ~n30143 & n43045;
  assign n30152 = pi53  & ~n30151;
  assign n30153 = pi53  & ~n30152;
  assign n30154 = pi53  & n30151;
  assign n30155 = ~n30151 & ~n30152;
  assign n30156 = ~pi53  & ~n30151;
  assign n30157 = ~n43046 & ~n43047;
  assign n30158 = ~n30142 & n30157;
  assign n30159 = n30142 & ~n30157;
  assign n30160 = ~n30158 & ~n30159;
  assign n30161 = ~n30063 & n30160;
  assign n30162 = n30063 & ~n30160;
  assign n30163 = ~n30063 & ~n30161;
  assign n30164 = n30160 & ~n30161;
  assign n30165 = ~n30163 & ~n30164;
  assign n30166 = ~n30161 & ~n30162;
  assign n30167 = ~n30062 & ~n43048;
  assign n30168 = n30062 & ~n30164;
  assign n30169 = ~n30163 & n30168;
  assign n30170 = n30062 & n43048;
  assign n30171 = ~n30167 & ~n43049;
  assign n30172 = ~n30047 & n30171;
  assign n30173 = n30047 & ~n30171;
  assign n30174 = ~n30172 & ~n30173;
  assign n30175 = n785 & n8177;
  assign n30176 = pi105  & n37520;
  assign n30177 = pi107  & n787;
  assign n30178 = pi106  & n795;
  assign n30179 = ~n30177 & ~n30178;
  assign n30180 = ~n30176 & ~n30178;
  assign n30181 = ~n30177 & n30180;
  assign n30182 = ~n30176 & n30179;
  assign n30183 = ~n30175 & n43050;
  assign n30184 = pi47  & ~n30183;
  assign n30185 = pi47  & ~n30184;
  assign n30186 = pi47  & n30183;
  assign n30187 = ~n30183 & ~n30184;
  assign n30188 = ~pi47  & ~n30183;
  assign n30189 = ~n43051 & ~n43052;
  assign n30190 = n30174 & ~n30189;
  assign n30191 = ~n30174 & n30189;
  assign n30192 = n30174 & ~n30190;
  assign n30193 = ~n30189 & ~n30190;
  assign n30194 = ~n30192 & ~n30193;
  assign n30195 = ~n30190 & ~n30191;
  assign n30196 = n30046 & n43053;
  assign n30197 = ~n30046 & ~n43053;
  assign n30198 = ~n30196 & ~n30197;
  assign n30199 = n940 & n9678;
  assign n30200 = pi108  & n37541;
  assign n30201 = pi110  & n953;
  assign n30202 = pi109  & n955;
  assign n30203 = ~n30201 & ~n30202;
  assign n30204 = ~n30200 & ~n30202;
  assign n30205 = ~n30201 & n30204;
  assign n30206 = ~n30200 & n30203;
  assign n30207 = ~n30199 & n43054;
  assign n30208 = pi44  & ~n30207;
  assign n30209 = pi44  & ~n30208;
  assign n30210 = pi44  & n30207;
  assign n30211 = ~n30207 & ~n30208;
  assign n30212 = ~pi44  & ~n30207;
  assign n30213 = ~n43055 & ~n43056;
  assign n30214 = ~n30198 & n30213;
  assign n30215 = n30198 & ~n30213;
  assign n30216 = n30198 & ~n30215;
  assign n30217 = ~n30213 & ~n30215;
  assign n30218 = ~n30216 & ~n30217;
  assign n30219 = ~n30214 & ~n30215;
  assign n30220 = n30045 & n43057;
  assign n30221 = ~n30045 & ~n43057;
  assign n30222 = ~n30220 & ~n30221;
  assign n30223 = n733 & n11276;
  assign n30224 = pi111  & n37510;
  assign n30225 = pi113  & n746;
  assign n30226 = pi112  & n748;
  assign n30227 = ~n30225 & ~n30226;
  assign n30228 = ~n30224 & ~n30226;
  assign n30229 = ~n30225 & n30228;
  assign n30230 = ~n30224 & n30227;
  assign n30231 = ~n30223 & n43058;
  assign n30232 = pi41  & ~n30231;
  assign n30233 = pi41  & ~n30232;
  assign n30234 = pi41  & n30231;
  assign n30235 = ~n30231 & ~n30232;
  assign n30236 = ~pi41  & ~n30231;
  assign n30237 = ~n43059 & ~n43060;
  assign n30238 = n30222 & ~n30237;
  assign n30239 = ~n30222 & n30237;
  assign n30240 = n30222 & ~n30238;
  assign n30241 = ~n30237 & ~n30238;
  assign n30242 = ~n30240 & ~n30241;
  assign n30243 = ~n30238 & ~n30239;
  assign n30244 = n30044 & n43061;
  assign n30245 = ~n30044 & ~n43061;
  assign n30246 = ~n30244 & ~n30245;
  assign n30247 = n691 & n12530;
  assign n30248 = pi114  & n37503;
  assign n30249 = pi116  & n704;
  assign n30250 = pi115  & n706;
  assign n30251 = ~n30249 & ~n30250;
  assign n30252 = ~n30248 & ~n30250;
  assign n30253 = ~n30249 & n30252;
  assign n30254 = ~n30248 & n30251;
  assign n30255 = ~n30247 & n43062;
  assign n30256 = pi38  & ~n30255;
  assign n30257 = pi38  & ~n30256;
  assign n30258 = pi38  & n30255;
  assign n30259 = ~n30255 & ~n30256;
  assign n30260 = ~pi38  & ~n30255;
  assign n30261 = ~n43063 & ~n43064;
  assign n30262 = ~n30246 & n30261;
  assign n30263 = n30246 & ~n30261;
  assign n30264 = n30246 & ~n30263;
  assign n30265 = ~n30261 & ~n30263;
  assign n30266 = ~n30264 & ~n30265;
  assign n30267 = ~n30262 & ~n30263;
  assign n30268 = ~n43012 & ~n43065;
  assign n30269 = n43012 & n43065;
  assign n30270 = ~n43012 & n43065;
  assign n30271 = n43012 & ~n43065;
  assign n30272 = ~n30270 & ~n30271;
  assign n30273 = ~n30268 & ~n30269;
  assign n30274 = ~n30043 & ~n43066;
  assign n30275 = n30043 & n43066;
  assign n30276 = ~n30274 & ~n30275;
  assign n30277 = n30028 & n30276;
  assign n30278 = ~n30028 & ~n30276;
  assign n30279 = ~n30277 & ~n30278;
  assign n30280 = n607 & n15068;
  assign n30281 = pi123  & n37489;
  assign n30282 = pi125  & n620;
  assign n30283 = pi124  & n622;
  assign n30284 = ~n30282 & ~n30283;
  assign n30285 = ~n30281 & ~n30283;
  assign n30286 = ~n30282 & n30285;
  assign n30287 = ~n30281 & n30284;
  assign n30288 = ~n30280 & n43067;
  assign n30289 = pi29  & ~n30288;
  assign n30290 = pi29  & ~n30289;
  assign n30291 = pi29  & n30288;
  assign n30292 = ~n30288 & ~n30289;
  assign n30293 = ~pi29  & ~n30288;
  assign n30294 = ~n43068 & ~n43069;
  assign n30295 = ~n29670 & ~n29954;
  assign n30296 = ~n30294 & ~n30295;
  assign n30297 = n30294 & n30295;
  assign n30298 = ~n30294 & ~n30296;
  assign n30299 = ~n30294 & n30295;
  assign n30300 = ~n30295 & ~n30296;
  assign n30301 = n30294 & ~n30295;
  assign n30302 = ~n43070 & ~n43071;
  assign n30303 = ~n30296 & ~n30297;
  assign n30304 = n30279 & ~n43072;
  assign n30305 = ~n30279 & n43072;
  assign n30306 = ~n43072 & ~n30304;
  assign n30307 = ~n30279 & ~n43072;
  assign n30308 = n30279 & ~n30304;
  assign n30309 = n30279 & n43072;
  assign n30310 = ~n43073 & ~n43074;
  assign n30311 = ~n30304 & ~n30305;
  assign n30312 = ~n29973 & ~n43020;
  assign n30313 = n4492 & n40891;
  assign n30314 = pi126  & n38208;
  assign n30315 = pi127  & n4509;
  assign n30316 = ~n30314 & ~n30315;
  assign n30317 = ~n4492 & n30316;
  assign n30318 = ~n40891 & n30316;
  assign n30319 = ~n30317 & ~n30318;
  assign n30320 = ~n30313 & n30316;
  assign n30321 = pi26  & ~n43076;
  assign n30322 = ~pi26  & n43076;
  assign n30323 = ~n30321 & ~n30322;
  assign n30324 = ~n30312 & ~n30323;
  assign n30325 = n30312 & n30323;
  assign n30326 = ~n30312 & ~n30324;
  assign n30327 = ~n30312 & n30323;
  assign n30328 = ~n30323 & ~n30324;
  assign n30329 = n30312 & ~n30323;
  assign n30330 = ~n43077 & ~n43078;
  assign n30331 = ~n30324 & ~n30325;
  assign n30332 = ~n43075 & ~n43079;
  assign n30333 = n43075 & ~n43078;
  assign n30334 = ~n43077 & n30333;
  assign n30335 = n43075 & ~n43077;
  assign n30336 = ~n43078 & n30335;
  assign n30337 = n43075 & n43079;
  assign n30338 = ~n30332 & ~n43080;
  assign n30339 = ~n30009 & n30338;
  assign n30340 = n30009 & ~n30338;
  assign n30341 = ~n30009 & ~n30339;
  assign n30342 = n30338 & ~n30339;
  assign n30343 = ~n30341 & ~n30342;
  assign n30344 = ~n30339 & ~n30340;
  assign n30345 = ~n30008 & ~n43081;
  assign n30346 = n30008 & ~n30342;
  assign n30347 = ~n30341 & n30346;
  assign n30348 = n30008 & n43081;
  assign po88  = ~n30345 & ~n43082;
  assign n30350 = ~n30339 & ~n30345;
  assign n30351 = ~n30324 & ~n30332;
  assign n30352 = n607 & n15021;
  assign n30353 = pi124  & n37489;
  assign n30354 = pi126  & n620;
  assign n30355 = pi125  & n622;
  assign n30356 = ~n30354 & ~n30355;
  assign n30357 = ~n30353 & ~n30355;
  assign n30358 = ~n30354 & n30357;
  assign n30359 = ~n30353 & n30356;
  assign n30360 = ~n30352 & n43083;
  assign n30361 = pi29  & ~n30360;
  assign n30362 = pi29  & ~n30361;
  assign n30363 = pi29  & n30360;
  assign n30364 = ~n30360 & ~n30361;
  assign n30365 = ~pi29  & ~n30360;
  assign n30366 = ~n43084 & ~n43085;
  assign n30367 = ~n30026 & ~n30277;
  assign n30368 = n30366 & n30367;
  assign n30369 = ~n30366 & ~n30367;
  assign n30370 = ~n30368 & ~n30369;
  assign n30371 = n649 & n14961;
  assign n30372 = pi121  & n37496;
  assign n30373 = pi123  & n662;
  assign n30374 = pi122  & n664;
  assign n30375 = ~n30373 & ~n30374;
  assign n30376 = ~n30372 & ~n30374;
  assign n30377 = ~n30373 & n30376;
  assign n30378 = ~n30372 & n30375;
  assign n30379 = ~n30371 & n43086;
  assign n30380 = pi32  & ~n30379;
  assign n30381 = pi32  & ~n30380;
  assign n30382 = pi32  & n30379;
  assign n30383 = ~n30379 & ~n30380;
  assign n30384 = ~pi32  & ~n30379;
  assign n30385 = ~n43087 & ~n43088;
  assign n30386 = ~n30268 & ~n30274;
  assign n30387 = n30385 & n30386;
  assign n30388 = ~n30385 & ~n30386;
  assign n30389 = ~n30387 & ~n30388;
  assign n30390 = n2104 & n14913;
  assign n30391 = pi118  & n37758;
  assign n30392 = pi120  & n2117;
  assign n30393 = pi119  & n2119;
  assign n30394 = ~n30392 & ~n30393;
  assign n30395 = ~n30391 & ~n30393;
  assign n30396 = ~n30392 & n30395;
  assign n30397 = ~n30391 & n30394;
  assign n30398 = ~n30390 & n43089;
  assign n30399 = pi35  & ~n30398;
  assign n30400 = pi35  & ~n30399;
  assign n30401 = pi35  & n30398;
  assign n30402 = ~n30398 & ~n30399;
  assign n30403 = ~pi35  & ~n30398;
  assign n30404 = ~n43090 & ~n43091;
  assign n30405 = n691 & n13079;
  assign n30406 = pi115  & n37503;
  assign n30407 = pi117  & n704;
  assign n30408 = pi116  & n706;
  assign n30409 = ~n30407 & ~n30408;
  assign n30410 = ~n30406 & ~n30408;
  assign n30411 = ~n30407 & n30410;
  assign n30412 = ~n30406 & n30409;
  assign n30413 = ~n30405 & n43092;
  assign n30414 = pi38  & ~n30413;
  assign n30415 = pi38  & ~n30414;
  assign n30416 = pi38  & n30413;
  assign n30417 = ~n30413 & ~n30414;
  assign n30418 = ~pi38  & ~n30413;
  assign n30419 = ~n43093 & ~n43094;
  assign n30420 = n785 & n9277;
  assign n30421 = pi106  & n37520;
  assign n30422 = pi108  & n787;
  assign n30423 = pi107  & n795;
  assign n30424 = ~n30422 & ~n30423;
  assign n30425 = ~n30421 & ~n30423;
  assign n30426 = ~n30422 & n30425;
  assign n30427 = ~n30421 & n30424;
  assign n30428 = ~n30420 & n43095;
  assign n30429 = pi47  & ~n30428;
  assign n30430 = pi47  & ~n30429;
  assign n30431 = pi47  & n30428;
  assign n30432 = ~n30428 & ~n30429;
  assign n30433 = ~pi47  & ~n30428;
  assign n30434 = ~n43096 & ~n43097;
  assign n30435 = ~n30161 & ~n30167;
  assign n30436 = n894 & n8229;
  assign n30437 = pi103  & n37580;
  assign n30438 = pi105  & n896;
  assign n30439 = pi104  & n904;
  assign n30440 = ~n30438 & ~n30439;
  assign n30441 = ~n30437 & ~n30439;
  assign n30442 = ~n30438 & n30441;
  assign n30443 = ~n30437 & n30440;
  assign n30444 = ~n30436 & n43098;
  assign n30445 = pi50  & ~n30444;
  assign n30446 = pi50  & ~n30445;
  assign n30447 = pi50  & n30444;
  assign n30448 = ~n30444 & ~n30445;
  assign n30449 = ~pi50  & ~n30444;
  assign n30450 = ~n43099 & ~n43100;
  assign n30451 = ~n30141 & ~n30159;
  assign n30452 = n4312 & n5578;
  assign n30453 = pi97  & n38376;
  assign n30454 = pi99  & n4314;
  assign n30455 = pi98  & n4322;
  assign n30456 = ~n30454 & ~n30455;
  assign n30457 = ~n30453 & ~n30455;
  assign n30458 = ~n30454 & n30457;
  assign n30459 = ~n30453 & n30456;
  assign n30460 = ~n30452 & n43101;
  assign n30461 = pi56  & ~n30460;
  assign n30462 = pi56  & ~n30461;
  assign n30463 = pi56  & n30460;
  assign n30464 = ~n30460 & ~n30461;
  assign n30465 = ~pi56  & ~n30460;
  assign n30466 = ~n43102 & ~n43103;
  assign n30467 = n5281 & n7882;
  assign n30468 = pi94  & n39128;
  assign n30469 = pi96  & n7884;
  assign n30470 = pi95  & n7892;
  assign n30471 = ~n30469 & ~n30470;
  assign n30472 = ~n30468 & ~n30470;
  assign n30473 = ~n30469 & n30472;
  assign n30474 = ~n30468 & n30471;
  assign n30475 = ~n30467 & n43104;
  assign n30476 = pi59  & ~n30475;
  assign n30477 = pi59  & ~n30476;
  assign n30478 = pi59  & n30475;
  assign n30479 = ~n30475 & ~n30476;
  assign n30480 = ~pi59  & ~n30475;
  assign n30481 = ~n43105 & ~n43106;
  assign n30482 = ~n30072 & ~n30089;
  assign n30483 = pi90  & ~n40814;
  assign n30484 = pi89  & n18285;
  assign n30485 = ~n30483 & ~n30484;
  assign n30486 = ~n30070 & n30485;
  assign n30487 = n30070 & ~n30485;
  assign n30488 = ~n30486 & ~n30487;
  assign n30489 = n4544 & n12674;
  assign n30490 = pi91  & n40107;
  assign n30491 = pi93  & n12676;
  assign n30492 = pi92  & n12684;
  assign n30493 = ~n30491 & ~n30492;
  assign n30494 = ~n30490 & ~n30492;
  assign n30495 = ~n30491 & n30494;
  assign n30496 = ~n30490 & n30493;
  assign n30497 = ~n12674 & n43107;
  assign n30498 = ~n4544 & n43107;
  assign n30499 = ~n30497 & ~n30498;
  assign n30500 = ~n30489 & n43107;
  assign n30501 = pi62  & ~n43108;
  assign n30502 = ~pi62  & n43108;
  assign n30503 = ~n30501 & ~n30502;
  assign n30504 = n30488 & ~n30503;
  assign n30505 = ~n30488 & n30503;
  assign n30506 = ~n30504 & ~n30505;
  assign n30507 = ~n30482 & n30506;
  assign n30508 = n30482 & ~n30506;
  assign n30509 = ~n30507 & ~n30508;
  assign n30510 = ~n30481 & n30509;
  assign n30511 = n30481 & ~n30509;
  assign n30512 = ~n30510 & ~n30511;
  assign n30513 = ~n30092 & n30109;
  assign n30514 = ~n30092 & ~n30110;
  assign n30515 = ~n30093 & ~n30513;
  assign n30516 = n30512 & ~n43109;
  assign n30517 = ~n30512 & n43109;
  assign n30518 = ~n30516 & ~n30517;
  assign n30519 = ~n30466 & n30518;
  assign n30520 = n30466 & ~n30518;
  assign n30521 = ~n30519 & ~n30520;
  assign n30522 = ~n30117 & n30133;
  assign n30523 = ~n30117 & ~n30135;
  assign n30524 = ~n30116 & ~n30522;
  assign n30525 = n30521 & ~n43110;
  assign n30526 = ~n30521 & n43110;
  assign n30527 = ~n30525 & ~n30526;
  assign n30528 = n1971 & n6819;
  assign n30529 = pi100  & n37864;
  assign n30530 = pi102  & n1973;
  assign n30531 = pi101  & n1981;
  assign n30532 = ~n30530 & ~n30531;
  assign n30533 = ~n30529 & ~n30531;
  assign n30534 = ~n30530 & n30533;
  assign n30535 = ~n30529 & n30532;
  assign n30536 = ~n30528 & n43111;
  assign n30537 = pi53  & ~n30536;
  assign n30538 = pi53  & ~n30537;
  assign n30539 = pi53  & n30536;
  assign n30540 = ~n30536 & ~n30537;
  assign n30541 = ~pi53  & ~n30536;
  assign n30542 = ~n43112 & ~n43113;
  assign n30543 = n30527 & ~n30542;
  assign n30544 = ~n30527 & n30542;
  assign n30545 = n30527 & ~n30543;
  assign n30546 = ~n30542 & ~n30543;
  assign n30547 = ~n30545 & ~n30546;
  assign n30548 = ~n30543 & ~n30544;
  assign n30549 = ~n30451 & ~n43114;
  assign n30550 = n30451 & n43114;
  assign n30551 = ~n43114 & ~n30549;
  assign n30552 = ~n30451 & ~n30549;
  assign n30553 = ~n30551 & ~n30552;
  assign n30554 = ~n30549 & ~n30550;
  assign n30555 = n30450 & ~n43115;
  assign n30556 = ~n30450 & n43115;
  assign n30557 = ~n30450 & ~n43115;
  assign n30558 = n30450 & n43115;
  assign n30559 = ~n30557 & ~n30558;
  assign n30560 = ~n30555 & ~n30556;
  assign n30561 = ~n30435 & n43116;
  assign n30562 = n30435 & ~n43116;
  assign n30563 = ~n30561 & ~n30562;
  assign n30564 = ~n30434 & n30563;
  assign n30565 = n30434 & ~n30563;
  assign n30566 = ~n30564 & ~n30565;
  assign n30567 = ~n30172 & n30189;
  assign n30568 = ~n30172 & ~n30190;
  assign n30569 = ~n30173 & ~n30567;
  assign n30570 = n30566 & ~n43117;
  assign n30571 = ~n30566 & n43117;
  assign n30572 = ~n30570 & ~n30571;
  assign n30573 = n565 & n940;
  assign n30574 = pi109  & n37541;
  assign n30575 = pi111  & n953;
  assign n30576 = pi110  & n955;
  assign n30577 = ~n30575 & ~n30576;
  assign n30578 = ~n30574 & ~n30576;
  assign n30579 = ~n30575 & n30578;
  assign n30580 = ~n30574 & n30577;
  assign n30581 = ~n30573 & n43118;
  assign n30582 = pi44  & ~n30581;
  assign n30583 = pi44  & ~n30582;
  assign n30584 = pi44  & n30581;
  assign n30585 = ~n30581 & ~n30582;
  assign n30586 = ~pi44  & ~n30581;
  assign n30587 = ~n43119 & ~n43120;
  assign n30588 = n30572 & ~n30587;
  assign n30589 = ~n30572 & n30587;
  assign n30590 = n30572 & ~n30588;
  assign n30591 = ~n30587 & ~n30588;
  assign n30592 = ~n30590 & ~n30591;
  assign n30593 = ~n30588 & ~n30589;
  assign n30594 = ~n30197 & n30213;
  assign n30595 = ~n30197 & ~n30215;
  assign n30596 = ~n30196 & ~n30594;
  assign n30597 = n43121 & n43122;
  assign n30598 = ~n43121 & ~n43122;
  assign n30599 = ~n30597 & ~n30598;
  assign n30600 = n733 & n11258;
  assign n30601 = pi112  & n37510;
  assign n30602 = pi114  & n746;
  assign n30603 = pi113  & n748;
  assign n30604 = ~n30602 & ~n30603;
  assign n30605 = ~n30601 & ~n30603;
  assign n30606 = ~n30602 & n30605;
  assign n30607 = ~n30601 & n30604;
  assign n30608 = ~n30600 & n43123;
  assign n30609 = pi41  & ~n30608;
  assign n30610 = pi41  & ~n30609;
  assign n30611 = pi41  & n30608;
  assign n30612 = ~n30608 & ~n30609;
  assign n30613 = ~pi41  & ~n30608;
  assign n30614 = ~n43124 & ~n43125;
  assign n30615 = ~n30599 & n30614;
  assign n30616 = n30599 & ~n30614;
  assign n30617 = ~n30615 & ~n30616;
  assign n30618 = ~n30221 & n30237;
  assign n30619 = ~n30221 & ~n30238;
  assign n30620 = ~n30220 & ~n30618;
  assign n30621 = n30617 & ~n43126;
  assign n30622 = ~n30617 & n43126;
  assign n30623 = ~n43126 & ~n30621;
  assign n30624 = n30617 & ~n30621;
  assign n30625 = ~n30623 & ~n30624;
  assign n30626 = ~n30621 & ~n30622;
  assign n30627 = ~n30419 & ~n43127;
  assign n30628 = n30419 & ~n30624;
  assign n30629 = ~n30623 & n30628;
  assign n30630 = n30419 & n43127;
  assign n30631 = ~n30627 & ~n43128;
  assign n30632 = ~n30245 & n30261;
  assign n30633 = ~n30245 & ~n30263;
  assign n30634 = ~n30244 & ~n30632;
  assign n30635 = n30631 & ~n43129;
  assign n30636 = ~n30631 & n43129;
  assign n30637 = ~n30635 & ~n30636;
  assign n30638 = n30404 & ~n30637;
  assign n30639 = ~n30404 & n30637;
  assign n30640 = ~n30404 & ~n30639;
  assign n30641 = n30637 & ~n30639;
  assign n30642 = ~n30640 & ~n30641;
  assign n30643 = ~n30638 & ~n30639;
  assign n30644 = n30389 & ~n43130;
  assign n30645 = ~n30389 & n43130;
  assign n30646 = n30389 & ~n30644;
  assign n30647 = ~n43130 & ~n30644;
  assign n30648 = ~n30646 & ~n30647;
  assign n30649 = ~n30644 & ~n30645;
  assign n30650 = ~n30370 & n43131;
  assign n30651 = n30370 & ~n43131;
  assign n30652 = ~n30650 & ~n30651;
  assign n30653 = ~n30296 & ~n30304;
  assign n30654 = n4492 & ~n18675;
  assign n30655 = ~n38208 & ~n30654;
  assign n30656 = pi127  & n38208;
  assign n30657 = n4492 & n18680;
  assign n30658 = ~n30656 & ~n30657;
  assign n30659 = pi127  & ~n30655;
  assign n30660 = pi26  & ~n43132;
  assign n30661 = pi26  & ~n30660;
  assign n30662 = pi26  & n43132;
  assign n30663 = ~n43132 & ~n30660;
  assign n30664 = ~pi26  & ~n43132;
  assign n30665 = ~n43133 & ~n43134;
  assign n30666 = ~n30653 & ~n30665;
  assign n30667 = n30653 & n30665;
  assign n30668 = ~n30653 & ~n30666;
  assign n30669 = ~n30665 & ~n30666;
  assign n30670 = ~n30668 & ~n30669;
  assign n30671 = ~n30666 & ~n30667;
  assign n30672 = n30652 & ~n43135;
  assign n30673 = ~n30652 & n43135;
  assign n30674 = ~n30672 & ~n30673;
  assign n30675 = ~n30351 & n30674;
  assign n30676 = n30351 & ~n30674;
  assign n30677 = ~n30675 & ~n30676;
  assign n30678 = ~n30350 & n30677;
  assign n30679 = n30350 & ~n30677;
  assign po89  = ~n30678 & ~n30679;
  assign n30681 = ~n30666 & ~n30672;
  assign n30682 = ~n30369 & ~n30651;
  assign n30683 = n607 & n40885;
  assign n30684 = pi125  & n37489;
  assign n30685 = pi127  & n620;
  assign n30686 = pi126  & n622;
  assign n30687 = ~n30685 & ~n30686;
  assign n30688 = ~n30684 & ~n30686;
  assign n30689 = ~n30685 & n30688;
  assign n30690 = ~n30684 & n30687;
  assign n30691 = ~n30683 & n43136;
  assign n30692 = pi29  & ~n30691;
  assign n30693 = pi29  & ~n30692;
  assign n30694 = pi29  & n30691;
  assign n30695 = ~n30691 & ~n30692;
  assign n30696 = ~pi29  & ~n30691;
  assign n30697 = ~n43137 & ~n43138;
  assign n30698 = ~n30682 & ~n30697;
  assign n30699 = n30682 & n30697;
  assign n30700 = ~n30682 & ~n30698;
  assign n30701 = ~n30682 & n30697;
  assign n30702 = ~n30697 & ~n30698;
  assign n30703 = n30682 & ~n30697;
  assign n30704 = ~n43139 & ~n43140;
  assign n30705 = ~n30698 & ~n30699;
  assign n30706 = ~n30621 & ~n30627;
  assign n30707 = n691 & n13057;
  assign n30708 = pi116  & n37503;
  assign n30709 = pi118  & n704;
  assign n30710 = pi117  & n706;
  assign n30711 = ~n30709 & ~n30710;
  assign n30712 = ~n30708 & ~n30710;
  assign n30713 = ~n30709 & n30712;
  assign n30714 = ~n30708 & n30711;
  assign n30715 = ~n30707 & n43142;
  assign n30716 = pi38  & ~n30715;
  assign n30717 = pi38  & ~n30716;
  assign n30718 = pi38  & n30715;
  assign n30719 = ~n30715 & ~n30716;
  assign n30720 = ~pi38  & ~n30715;
  assign n30721 = ~n43143 & ~n43144;
  assign n30722 = ~n30598 & ~n30616;
  assign n30723 = ~n30561 & ~n30564;
  assign n30724 = n785 & n9701;
  assign n30725 = pi107  & n37520;
  assign n30726 = pi109  & n787;
  assign n30727 = pi108  & n795;
  assign n30728 = ~n30726 & ~n30727;
  assign n30729 = ~n30725 & ~n30727;
  assign n30730 = ~n30726 & n30729;
  assign n30731 = ~n30725 & n30728;
  assign n30732 = ~n30724 & n43145;
  assign n30733 = pi47  & ~n30732;
  assign n30734 = pi47  & ~n30733;
  assign n30735 = pi47  & n30732;
  assign n30736 = ~n30732 & ~n30733;
  assign n30737 = ~pi47  & ~n30732;
  assign n30738 = ~n43146 & ~n43147;
  assign n30739 = ~n30516 & ~n30519;
  assign n30740 = n5630 & n7882;
  assign n30741 = pi95  & n39128;
  assign n30742 = pi97  & n7884;
  assign n30743 = pi96  & n7892;
  assign n30744 = ~n30742 & ~n30743;
  assign n30745 = ~n30741 & ~n30743;
  assign n30746 = ~n30742 & n30745;
  assign n30747 = ~n30741 & n30744;
  assign n30748 = ~n30740 & n43148;
  assign n30749 = pi59  & ~n30748;
  assign n30750 = pi59  & ~n30749;
  assign n30751 = pi59  & n30748;
  assign n30752 = ~n30748 & ~n30749;
  assign n30753 = ~pi59  & ~n30748;
  assign n30754 = ~n43149 & ~n43150;
  assign n30755 = ~n30507 & ~n30510;
  assign n30756 = n30754 & n30755;
  assign n30757 = ~n30754 & ~n30755;
  assign n30758 = ~n30756 & ~n30757;
  assign n30759 = ~n30486 & ~n30504;
  assign n30760 = pi91  & ~n40814;
  assign n30761 = pi90  & n18285;
  assign n30762 = ~n30760 & ~n30761;
  assign n30763 = ~pi26  & ~n30762;
  assign n30764 = pi26  & n30762;
  assign n30765 = ~n30763 & ~n30764;
  assign n30766 = ~n30485 & n30765;
  assign n30767 = n30485 & ~n30765;
  assign n30768 = ~n30766 & ~n30767;
  assign n30769 = ~n30759 & n30768;
  assign n30770 = n30759 & ~n30768;
  assign n30771 = ~n30769 & ~n30770;
  assign n30772 = n4524 & n12674;
  assign n30773 = pi92  & n40107;
  assign n30774 = pi94  & n12676;
  assign n30775 = pi93  & n12684;
  assign n30776 = ~n30774 & ~n30775;
  assign n30777 = ~n30773 & ~n30775;
  assign n30778 = ~n30774 & n30777;
  assign n30779 = ~n30773 & n30776;
  assign n30780 = ~n30772 & n43151;
  assign n30781 = pi62  & ~n30780;
  assign n30782 = pi62  & ~n30781;
  assign n30783 = pi62  & n30780;
  assign n30784 = ~n30780 & ~n30781;
  assign n30785 = ~pi62  & ~n30780;
  assign n30786 = ~n43152 & ~n43153;
  assign n30787 = n30771 & ~n30786;
  assign n30788 = ~n30771 & n30786;
  assign n30789 = n30771 & ~n30787;
  assign n30790 = ~n30786 & ~n30787;
  assign n30791 = ~n30789 & ~n30790;
  assign n30792 = ~n30787 & ~n30788;
  assign n30793 = ~n30758 & n43154;
  assign n30794 = n30758 & ~n43154;
  assign n30795 = ~n30793 & ~n30794;
  assign n30796 = n4312 & n6474;
  assign n30797 = pi98  & n38376;
  assign n30798 = pi100  & n4314;
  assign n30799 = pi99  & n4322;
  assign n30800 = ~n30798 & ~n30799;
  assign n30801 = ~n30797 & ~n30799;
  assign n30802 = ~n30798 & n30801;
  assign n30803 = ~n30797 & n30800;
  assign n30804 = ~n30796 & n43155;
  assign n30805 = pi56  & ~n30804;
  assign n30806 = pi56  & ~n30805;
  assign n30807 = pi56  & n30804;
  assign n30808 = ~n30804 & ~n30805;
  assign n30809 = ~pi56  & ~n30804;
  assign n30810 = ~n43156 & ~n43157;
  assign n30811 = n30795 & ~n30810;
  assign n30812 = ~n30795 & n30810;
  assign n30813 = n30795 & ~n30811;
  assign n30814 = n30795 & n30810;
  assign n30815 = ~n30810 & ~n30811;
  assign n30816 = ~n30795 & ~n30810;
  assign n30817 = ~n43158 & ~n43159;
  assign n30818 = ~n30811 & ~n30812;
  assign n30819 = n30739 & n43160;
  assign n30820 = ~n30739 & ~n43160;
  assign n30821 = ~n30819 & ~n30820;
  assign n30822 = n1971 & n6787;
  assign n30823 = pi101  & n37864;
  assign n30824 = pi103  & n1973;
  assign n30825 = pi102  & n1981;
  assign n30826 = ~n30824 & ~n30825;
  assign n30827 = ~n30823 & ~n30825;
  assign n30828 = ~n30824 & n30827;
  assign n30829 = ~n30823 & n30826;
  assign n30830 = ~n30822 & n43161;
  assign n30831 = pi53  & ~n30830;
  assign n30832 = pi53  & ~n30831;
  assign n30833 = pi53  & n30830;
  assign n30834 = ~n30830 & ~n30831;
  assign n30835 = ~pi53  & ~n30830;
  assign n30836 = ~n43162 & ~n43163;
  assign n30837 = n30821 & ~n30836;
  assign n30838 = ~n30821 & n30836;
  assign n30839 = n30821 & ~n30837;
  assign n30840 = n30821 & n30836;
  assign n30841 = ~n30836 & ~n30837;
  assign n30842 = ~n30821 & ~n30836;
  assign n30843 = ~n43164 & ~n43165;
  assign n30844 = ~n30837 & ~n30838;
  assign n30845 = ~n30525 & n30542;
  assign n30846 = ~n30525 & ~n30543;
  assign n30847 = ~n30526 & ~n30845;
  assign n30848 = n43166 & n43167;
  assign n30849 = ~n43166 & ~n43167;
  assign n30850 = ~n30848 & ~n30849;
  assign n30851 = n894 & n8209;
  assign n30852 = pi104  & n37580;
  assign n30853 = pi106  & n896;
  assign n30854 = pi105  & n904;
  assign n30855 = ~n30853 & ~n30854;
  assign n30856 = ~n30852 & ~n30854;
  assign n30857 = ~n30853 & n30856;
  assign n30858 = ~n30852 & n30855;
  assign n30859 = ~n30851 & n43168;
  assign n30860 = pi50  & ~n30859;
  assign n30861 = pi50  & ~n30860;
  assign n30862 = pi50  & n30859;
  assign n30863 = ~n30859 & ~n30860;
  assign n30864 = ~pi50  & ~n30859;
  assign n30865 = ~n43169 & ~n43170;
  assign n30866 = n30850 & ~n30865;
  assign n30867 = ~n30850 & n30865;
  assign n30868 = n30850 & ~n30866;
  assign n30869 = n30850 & n30865;
  assign n30870 = ~n30865 & ~n30866;
  assign n30871 = ~n30850 & ~n30865;
  assign n30872 = ~n43171 & ~n43172;
  assign n30873 = ~n30866 & ~n30867;
  assign n30874 = n30450 & ~n30549;
  assign n30875 = ~n30549 & ~n30557;
  assign n30876 = ~n30550 & ~n30874;
  assign n30877 = ~n43173 & ~n43174;
  assign n30878 = n43173 & n43174;
  assign n30879 = n43173 & ~n43174;
  assign n30880 = ~n43173 & n43174;
  assign n30881 = ~n30879 & ~n30880;
  assign n30882 = ~n30877 & ~n30878;
  assign n30883 = ~n30738 & ~n43175;
  assign n30884 = n30738 & n43175;
  assign n30885 = ~n30883 & ~n30884;
  assign n30886 = n30723 & ~n30885;
  assign n30887 = ~n30723 & n30885;
  assign n30888 = ~n30886 & ~n30887;
  assign n30889 = n940 & n10844;
  assign n30890 = pi110  & n37541;
  assign n30891 = pi112  & n953;
  assign n30892 = pi111  & n955;
  assign n30893 = ~n30891 & ~n30892;
  assign n30894 = ~n30890 & ~n30892;
  assign n30895 = ~n30891 & n30894;
  assign n30896 = ~n30890 & n30893;
  assign n30897 = ~n30889 & n43176;
  assign n30898 = pi44  & ~n30897;
  assign n30899 = pi44  & ~n30898;
  assign n30900 = pi44  & n30897;
  assign n30901 = ~n30897 & ~n30898;
  assign n30902 = ~pi44  & ~n30897;
  assign n30903 = ~n43177 & ~n43178;
  assign n30904 = n30888 & ~n30903;
  assign n30905 = ~n30888 & n30903;
  assign n30906 = n30888 & ~n30904;
  assign n30907 = n30888 & n30903;
  assign n30908 = ~n30903 & ~n30904;
  assign n30909 = ~n30888 & ~n30903;
  assign n30910 = ~n43179 & ~n43180;
  assign n30911 = ~n30904 & ~n30905;
  assign n30912 = ~n30570 & n30587;
  assign n30913 = ~n30570 & ~n30588;
  assign n30914 = ~n30571 & ~n30912;
  assign n30915 = n43181 & n43182;
  assign n30916 = ~n43181 & ~n43182;
  assign n30917 = ~n30915 & ~n30916;
  assign n30918 = n523 & n733;
  assign n30919 = pi113  & n37510;
  assign n30920 = pi115  & n746;
  assign n30921 = pi114  & n748;
  assign n30922 = ~n30920 & ~n30921;
  assign n30923 = ~n30919 & ~n30921;
  assign n30924 = ~n30920 & n30923;
  assign n30925 = ~n30919 & n30922;
  assign n30926 = ~n30918 & n43183;
  assign n30927 = pi41  & ~n30926;
  assign n30928 = pi41  & ~n30927;
  assign n30929 = pi41  & n30926;
  assign n30930 = ~n30926 & ~n30927;
  assign n30931 = ~pi41  & ~n30926;
  assign n30932 = ~n43184 & ~n43185;
  assign n30933 = n30917 & ~n30932;
  assign n30934 = ~n30917 & n30932;
  assign n30935 = ~n30933 & ~n30934;
  assign n30936 = n30722 & ~n30935;
  assign n30937 = ~n30722 & ~n30934;
  assign n30938 = ~n30933 & n30937;
  assign n30939 = ~n30722 & ~n30933;
  assign n30940 = ~n30934 & n30939;
  assign n30941 = ~n30722 & n30935;
  assign n30942 = ~n30722 & ~n43186;
  assign n30943 = ~n30722 & ~n30935;
  assign n30944 = n30722 & ~n30933;
  assign n30945 = ~n30933 & ~n43186;
  assign n30946 = ~n30934 & ~n30944;
  assign n30947 = ~n30934 & n43188;
  assign n30948 = n30722 & n30935;
  assign n30949 = ~n43187 & ~n43189;
  assign n30950 = ~n30936 & ~n43186;
  assign n30951 = n30721 & n43190;
  assign n30952 = ~n30721 & ~n43190;
  assign n30953 = ~n30951 & ~n30952;
  assign n30954 = ~n30706 & n30953;
  assign n30955 = n30706 & ~n30953;
  assign n30956 = ~n30954 & ~n30955;
  assign n30957 = n2104 & n15091;
  assign n30958 = pi119  & n37758;
  assign n30959 = pi121  & n2117;
  assign n30960 = pi120  & n2119;
  assign n30961 = ~n30959 & ~n30960;
  assign n30962 = ~n30958 & ~n30960;
  assign n30963 = ~n30959 & n30962;
  assign n30964 = ~n30958 & n30961;
  assign n30965 = ~n30957 & n43191;
  assign n30966 = pi35  & ~n30965;
  assign n30967 = pi35  & ~n30966;
  assign n30968 = pi35  & n30965;
  assign n30969 = ~n30965 & ~n30966;
  assign n30970 = ~pi35  & ~n30965;
  assign n30971 = ~n43192 & ~n43193;
  assign n30972 = n30956 & ~n30971;
  assign n30973 = ~n30956 & n30971;
  assign n30974 = n30956 & ~n30972;
  assign n30975 = n30956 & n30971;
  assign n30976 = ~n30971 & ~n30972;
  assign n30977 = ~n30956 & ~n30971;
  assign n30978 = ~n43194 & ~n43195;
  assign n30979 = ~n30972 & ~n30973;
  assign n30980 = n30404 & ~n30635;
  assign n30981 = ~n30635 & ~n30639;
  assign n30982 = ~n30636 & ~n30980;
  assign n30983 = n43196 & n43197;
  assign n30984 = ~n43196 & ~n43197;
  assign n30985 = ~n30983 & ~n30984;
  assign n30986 = n649 & n15111;
  assign n30987 = pi122  & n37496;
  assign n30988 = pi124  & n662;
  assign n30989 = pi123  & n664;
  assign n30990 = ~n30988 & ~n30989;
  assign n30991 = ~n30987 & ~n30989;
  assign n30992 = ~n30988 & n30991;
  assign n30993 = ~n30987 & n30990;
  assign n30994 = ~n30986 & n43198;
  assign n30995 = pi32  & ~n30994;
  assign n30996 = pi32  & ~n30995;
  assign n30997 = pi32  & n30994;
  assign n30998 = ~n30994 & ~n30995;
  assign n30999 = ~pi32  & ~n30994;
  assign n31000 = ~n43199 & ~n43200;
  assign n31001 = ~n30388 & n43130;
  assign n31002 = ~n30388 & ~n30644;
  assign n31003 = ~n30387 & ~n31001;
  assign n31004 = n31000 & n43201;
  assign n31005 = ~n31000 & ~n43201;
  assign n31006 = ~n31004 & ~n31005;
  assign n31007 = n30985 & n31006;
  assign n31008 = ~n30985 & ~n31006;
  assign n31009 = n30985 & ~n31006;
  assign n31010 = ~n30985 & n31006;
  assign n31011 = ~n31009 & ~n31010;
  assign n31012 = ~n31007 & ~n31008;
  assign n31013 = ~n43141 & ~n43202;
  assign n31014 = n43141 & n43202;
  assign n31015 = ~n31013 & ~n31014;
  assign n31016 = n30681 & ~n31015;
  assign n31017 = ~n30681 & n31015;
  assign n31018 = ~n31016 & ~n31017;
  assign n31019 = ~n30675 & ~n30678;
  assign n31020 = n31018 & ~n31019;
  assign n31021 = ~n31018 & n31019;
  assign po90  = ~n31020 & ~n31021;
  assign n31023 = ~n30698 & ~n31013;
  assign n31024 = n607 & n40891;
  assign n31025 = pi126  & n37489;
  assign n31026 = pi127  & n622;
  assign n31027 = ~n31025 & ~n31026;
  assign n31028 = ~n607 & n31027;
  assign n31029 = ~n40891 & n31027;
  assign n31030 = ~n31028 & ~n31029;
  assign n31031 = ~n31024 & n31027;
  assign n31032 = pi29  & ~n43203;
  assign n31033 = ~pi29  & n43203;
  assign n31034 = ~n31032 & ~n31033;
  assign n31035 = ~n30985 & ~n31005;
  assign n31036 = ~n31005 & ~n31007;
  assign n31037 = ~n31004 & ~n31035;
  assign n31038 = ~n31034 & ~n43204;
  assign n31039 = n31034 & n43204;
  assign n31040 = ~n31038 & ~n31039;
  assign n31041 = n649 & n15068;
  assign n31042 = pi123  & n37496;
  assign n31043 = pi125  & n662;
  assign n31044 = pi124  & n664;
  assign n31045 = ~n31043 & ~n31044;
  assign n31046 = ~n31042 & ~n31044;
  assign n31047 = ~n31043 & n31046;
  assign n31048 = ~n31042 & n31045;
  assign n31049 = ~n31041 & n43205;
  assign n31050 = pi32  & ~n31049;
  assign n31051 = pi32  & ~n31050;
  assign n31052 = pi32  & n31049;
  assign n31053 = ~n31049 & ~n31050;
  assign n31054 = ~pi32  & ~n31049;
  assign n31055 = ~n43206 & ~n43207;
  assign n31056 = ~n30972 & ~n30984;
  assign n31057 = n31055 & n31056;
  assign n31058 = ~n31055 & ~n31056;
  assign n31059 = ~n31057 & ~n31058;
  assign n31060 = ~n30952 & ~n30954;
  assign n31061 = n691 & n13027;
  assign n31062 = pi117  & n37503;
  assign n31063 = pi119  & n704;
  assign n31064 = pi118  & n706;
  assign n31065 = ~n31063 & ~n31064;
  assign n31066 = ~n31062 & ~n31064;
  assign n31067 = ~n31063 & n31066;
  assign n31068 = ~n31062 & n31065;
  assign n31069 = ~n31061 & n43208;
  assign n31070 = pi38  & ~n31069;
  assign n31071 = pi38  & ~n31070;
  assign n31072 = pi38  & n31069;
  assign n31073 = ~n31069 & ~n31070;
  assign n31074 = ~pi38  & ~n31069;
  assign n31075 = ~n43209 & ~n43210;
  assign n31076 = ~n30904 & ~n30916;
  assign n31077 = ~n30883 & ~n30887;
  assign n31078 = ~n30866 & ~n30877;
  assign n31079 = ~n30837 & ~n30849;
  assign n31080 = n1971 & n8136;
  assign n31081 = pi102  & n37864;
  assign n31082 = pi104  & n1973;
  assign n31083 = pi103  & n1981;
  assign n31084 = ~n31082 & ~n31083;
  assign n31085 = ~n31081 & ~n31083;
  assign n31086 = ~n31082 & n31085;
  assign n31087 = ~n31081 & n31084;
  assign n31088 = ~n31080 & n43211;
  assign n31089 = pi53  & ~n31088;
  assign n31090 = pi53  & ~n31089;
  assign n31091 = pi53  & n31088;
  assign n31092 = ~n31088 & ~n31089;
  assign n31093 = ~pi53  & ~n31088;
  assign n31094 = ~n43212 & ~n43213;
  assign n31095 = ~n30811 & ~n30820;
  assign n31096 = n4312 & n6839;
  assign n31097 = pi99  & n38376;
  assign n31098 = pi101  & n4314;
  assign n31099 = pi100  & n4322;
  assign n31100 = ~n31098 & ~n31099;
  assign n31101 = ~n31097 & ~n31099;
  assign n31102 = ~n31098 & n31101;
  assign n31103 = ~n31097 & n31100;
  assign n31104 = ~n31096 & n43214;
  assign n31105 = pi56  & ~n31104;
  assign n31106 = pi56  & ~n31105;
  assign n31107 = pi56  & n31104;
  assign n31108 = ~n31104 & ~n31105;
  assign n31109 = ~pi56  & ~n31104;
  assign n31110 = ~n43215 & ~n43216;
  assign n31111 = ~n30757 & ~n30794;
  assign n31112 = ~n30763 & ~n30766;
  assign n31113 = pi92  & ~n40814;
  assign n31114 = pi91  & n18285;
  assign n31115 = ~n31113 & ~n31114;
  assign n31116 = n31112 & ~n31115;
  assign n31117 = ~n31112 & n31115;
  assign n31118 = ~n31116 & ~n31117;
  assign n31119 = n4494 & n12674;
  assign n31120 = pi93  & n40107;
  assign n31121 = pi95  & n12676;
  assign n31122 = pi94  & n12684;
  assign n31123 = ~n31121 & ~n31122;
  assign n31124 = ~n31120 & ~n31122;
  assign n31125 = ~n31121 & n31124;
  assign n31126 = ~n31120 & n31123;
  assign n31127 = ~n31119 & n43217;
  assign n31128 = pi62  & ~n31127;
  assign n31129 = pi62  & ~n31128;
  assign n31130 = pi62  & n31127;
  assign n31131 = ~n31127 & ~n31128;
  assign n31132 = ~pi62  & ~n31127;
  assign n31133 = ~n43218 & ~n43219;
  assign n31134 = ~n31118 & n31133;
  assign n31135 = n31118 & ~n31133;
  assign n31136 = ~n31134 & ~n31135;
  assign n31137 = ~n30769 & n30786;
  assign n31138 = ~n30769 & ~n30787;
  assign n31139 = ~n30770 & ~n31137;
  assign n31140 = n31136 & ~n43220;
  assign n31141 = ~n31136 & n43220;
  assign n31142 = ~n31140 & ~n31141;
  assign n31143 = n5610 & n7882;
  assign n31144 = pi96  & n39128;
  assign n31145 = pi98  & n7884;
  assign n31146 = pi97  & n7892;
  assign n31147 = ~n31145 & ~n31146;
  assign n31148 = ~n31144 & ~n31146;
  assign n31149 = ~n31145 & n31148;
  assign n31150 = ~n31144 & n31147;
  assign n31151 = ~n31143 & n43221;
  assign n31152 = pi59  & ~n31151;
  assign n31153 = pi59  & ~n31152;
  assign n31154 = pi59  & n31151;
  assign n31155 = ~n31151 & ~n31152;
  assign n31156 = ~pi59  & ~n31151;
  assign n31157 = ~n43222 & ~n43223;
  assign n31158 = n31142 & ~n31157;
  assign n31159 = ~n31142 & n31157;
  assign n31160 = n31142 & ~n31158;
  assign n31161 = ~n31157 & ~n31158;
  assign n31162 = ~n31160 & ~n31161;
  assign n31163 = ~n31158 & ~n31159;
  assign n31164 = ~n31111 & ~n43224;
  assign n31165 = n31111 & n43224;
  assign n31166 = ~n43224 & ~n31164;
  assign n31167 = ~n31111 & ~n31164;
  assign n31168 = ~n31166 & ~n31167;
  assign n31169 = ~n31164 & ~n31165;
  assign n31170 = n31110 & ~n43225;
  assign n31171 = ~n31110 & n43225;
  assign n31172 = ~n31110 & ~n43225;
  assign n31173 = n31110 & n43225;
  assign n31174 = ~n31172 & ~n31173;
  assign n31175 = ~n31170 & ~n31171;
  assign n31176 = ~n31095 & n43226;
  assign n31177 = n31095 & ~n43226;
  assign n31178 = ~n31095 & ~n31176;
  assign n31179 = n43226 & ~n31176;
  assign n31180 = ~n31178 & ~n31179;
  assign n31181 = ~n31176 & ~n31177;
  assign n31182 = ~n31094 & ~n43227;
  assign n31183 = n31094 & ~n31179;
  assign n31184 = ~n31178 & n31183;
  assign n31185 = n31094 & n43227;
  assign n31186 = ~n31182 & ~n43228;
  assign n31187 = ~n31079 & n31186;
  assign n31188 = n31079 & ~n31186;
  assign n31189 = ~n31187 & ~n31188;
  assign n31190 = n894 & n8177;
  assign n31191 = pi105  & n37580;
  assign n31192 = pi107  & n896;
  assign n31193 = pi106  & n904;
  assign n31194 = ~n31192 & ~n31193;
  assign n31195 = ~n31191 & ~n31193;
  assign n31196 = ~n31192 & n31195;
  assign n31197 = ~n31191 & n31194;
  assign n31198 = ~n31190 & n43229;
  assign n31199 = pi50  & ~n31198;
  assign n31200 = pi50  & ~n31199;
  assign n31201 = pi50  & n31198;
  assign n31202 = ~n31198 & ~n31199;
  assign n31203 = ~pi50  & ~n31198;
  assign n31204 = ~n43230 & ~n43231;
  assign n31205 = n31189 & ~n31204;
  assign n31206 = ~n31189 & n31204;
  assign n31207 = n31189 & ~n31205;
  assign n31208 = ~n31204 & ~n31205;
  assign n31209 = ~n31207 & ~n31208;
  assign n31210 = ~n31205 & ~n31206;
  assign n31211 = n31078 & n43232;
  assign n31212 = ~n31078 & ~n43232;
  assign n31213 = ~n31211 & ~n31212;
  assign n31214 = n785 & n9678;
  assign n31215 = pi108  & n37520;
  assign n31216 = pi110  & n787;
  assign n31217 = pi109  & n795;
  assign n31218 = ~n31216 & ~n31217;
  assign n31219 = ~n31215 & ~n31217;
  assign n31220 = ~n31216 & n31219;
  assign n31221 = ~n31215 & n31218;
  assign n31222 = ~n31214 & n43233;
  assign n31223 = pi47  & ~n31222;
  assign n31224 = pi47  & ~n31223;
  assign n31225 = pi47  & n31222;
  assign n31226 = ~n31222 & ~n31223;
  assign n31227 = ~pi47  & ~n31222;
  assign n31228 = ~n43234 & ~n43235;
  assign n31229 = ~n31213 & n31228;
  assign n31230 = n31213 & ~n31228;
  assign n31231 = n31213 & ~n31230;
  assign n31232 = ~n31228 & ~n31230;
  assign n31233 = ~n31231 & ~n31232;
  assign n31234 = ~n31229 & ~n31230;
  assign n31235 = n31077 & n43236;
  assign n31236 = ~n31077 & ~n43236;
  assign n31237 = ~n31235 & ~n31236;
  assign n31238 = n940 & n11276;
  assign n31239 = pi111  & n37541;
  assign n31240 = pi113  & n953;
  assign n31241 = pi112  & n955;
  assign n31242 = ~n31240 & ~n31241;
  assign n31243 = ~n31239 & ~n31241;
  assign n31244 = ~n31240 & n31243;
  assign n31245 = ~n31239 & n31242;
  assign n31246 = ~n31238 & n43237;
  assign n31247 = pi44  & ~n31246;
  assign n31248 = pi44  & ~n31247;
  assign n31249 = pi44  & n31246;
  assign n31250 = ~n31246 & ~n31247;
  assign n31251 = ~pi44  & ~n31246;
  assign n31252 = ~n43238 & ~n43239;
  assign n31253 = n31237 & ~n31252;
  assign n31254 = ~n31237 & n31252;
  assign n31255 = n31237 & ~n31253;
  assign n31256 = ~n31252 & ~n31253;
  assign n31257 = ~n31255 & ~n31256;
  assign n31258 = ~n31253 & ~n31254;
  assign n31259 = n31076 & n43240;
  assign n31260 = ~n31076 & ~n43240;
  assign n31261 = ~n31259 & ~n31260;
  assign n31262 = n733 & n12530;
  assign n31263 = pi114  & n37510;
  assign n31264 = pi116  & n746;
  assign n31265 = pi115  & n748;
  assign n31266 = ~n31264 & ~n31265;
  assign n31267 = ~n31263 & ~n31265;
  assign n31268 = ~n31264 & n31267;
  assign n31269 = ~n31263 & n31266;
  assign n31270 = ~n31262 & n43241;
  assign n31271 = pi41  & ~n31270;
  assign n31272 = pi41  & ~n31271;
  assign n31273 = pi41  & n31270;
  assign n31274 = ~n31270 & ~n31271;
  assign n31275 = ~pi41  & ~n31270;
  assign n31276 = ~n43242 & ~n43243;
  assign n31277 = ~n31261 & n31276;
  assign n31278 = n31261 & ~n31276;
  assign n31279 = n31261 & ~n31278;
  assign n31280 = ~n31276 & ~n31278;
  assign n31281 = ~n31279 & ~n31280;
  assign n31282 = ~n31277 & ~n31278;
  assign n31283 = ~n43188 & ~n43244;
  assign n31284 = n43188 & n43244;
  assign n31285 = ~n43188 & n43244;
  assign n31286 = n43188 & ~n43244;
  assign n31287 = ~n31285 & ~n31286;
  assign n31288 = ~n31283 & ~n31284;
  assign n31289 = ~n31075 & ~n43245;
  assign n31290 = n31075 & n43245;
  assign n31291 = ~n31289 & ~n31290;
  assign n31292 = ~n31060 & n31291;
  assign n31293 = n31060 & ~n31291;
  assign n31294 = ~n31292 & ~n31293;
  assign n31295 = n2104 & n15049;
  assign n31296 = pi120  & n37758;
  assign n31297 = pi122  & n2117;
  assign n31298 = pi121  & n2119;
  assign n31299 = ~n31297 & ~n31298;
  assign n31300 = ~n31296 & ~n31298;
  assign n31301 = ~n31297 & n31300;
  assign n31302 = ~n31296 & n31299;
  assign n31303 = ~n31295 & n43246;
  assign n31304 = pi35  & ~n31303;
  assign n31305 = pi35  & ~n31304;
  assign n31306 = pi35  & n31303;
  assign n31307 = ~n31303 & ~n31304;
  assign n31308 = ~pi35  & ~n31303;
  assign n31309 = ~n43247 & ~n43248;
  assign n31310 = n31294 & ~n31309;
  assign n31311 = ~n31294 & n31309;
  assign n31312 = n31294 & ~n31310;
  assign n31313 = ~n31309 & ~n31310;
  assign n31314 = ~n31312 & ~n31313;
  assign n31315 = ~n31310 & ~n31311;
  assign n31316 = n31059 & ~n43249;
  assign n31317 = ~n31059 & n43249;
  assign n31318 = ~n31316 & ~n31317;
  assign n31319 = n31040 & ~n31317;
  assign n31320 = ~n31316 & n31319;
  assign n31321 = n31040 & n31318;
  assign n31322 = ~n31040 & ~n31318;
  assign n31323 = n31040 & ~n43250;
  assign n31324 = ~n31317 & ~n43250;
  assign n31325 = ~n31316 & n31324;
  assign n31326 = n31318 & ~n43250;
  assign n31327 = ~n31323 & ~n43251;
  assign n31328 = ~n43250 & ~n31322;
  assign n31329 = n31023 & n43252;
  assign n31330 = ~n31023 & ~n43252;
  assign n31331 = ~n31329 & ~n31330;
  assign n31332 = ~n31017 & ~n31020;
  assign n31333 = n31331 & ~n31332;
  assign n31334 = ~n31331 & n31332;
  assign po91  = ~n31333 & ~n31334;
  assign n31336 = ~n31330 & ~n31333;
  assign n31337 = ~n31038 & ~n43250;
  assign n31338 = n649 & n15021;
  assign n31339 = pi124  & n37496;
  assign n31340 = pi126  & n662;
  assign n31341 = pi125  & n664;
  assign n31342 = ~n31340 & ~n31341;
  assign n31343 = ~n31339 & ~n31341;
  assign n31344 = ~n31340 & n31343;
  assign n31345 = ~n31339 & n31342;
  assign n31346 = ~n31338 & n43253;
  assign n31347 = pi32  & ~n31346;
  assign n31348 = pi32  & ~n31347;
  assign n31349 = pi32  & n31346;
  assign n31350 = ~n31346 & ~n31347;
  assign n31351 = ~pi32  & ~n31346;
  assign n31352 = ~n43254 & ~n43255;
  assign n31353 = ~n31292 & n31309;
  assign n31354 = ~n31292 & ~n31310;
  assign n31355 = ~n31293 & ~n31353;
  assign n31356 = n31352 & n43256;
  assign n31357 = ~n31352 & ~n43256;
  assign n31358 = ~n31356 & ~n31357;
  assign n31359 = ~n31283 & ~n31289;
  assign n31360 = n691 & n14913;
  assign n31361 = pi118  & n37503;
  assign n31362 = pi120  & n704;
  assign n31363 = pi119  & n706;
  assign n31364 = ~n31362 & ~n31363;
  assign n31365 = ~n31361 & ~n31363;
  assign n31366 = ~n31362 & n31365;
  assign n31367 = ~n31361 & n31364;
  assign n31368 = ~n31360 & n43257;
  assign n31369 = pi38  & ~n31368;
  assign n31370 = pi38  & ~n31369;
  assign n31371 = pi38  & n31368;
  assign n31372 = ~n31368 & ~n31369;
  assign n31373 = ~pi38  & ~n31368;
  assign n31374 = ~n43258 & ~n43259;
  assign n31375 = n733 & n13079;
  assign n31376 = pi115  & n37510;
  assign n31377 = pi117  & n746;
  assign n31378 = pi116  & n748;
  assign n31379 = ~n31377 & ~n31378;
  assign n31380 = ~n31376 & ~n31378;
  assign n31381 = ~n31377 & n31380;
  assign n31382 = ~n31376 & n31379;
  assign n31383 = ~n31375 & n43260;
  assign n31384 = pi41  & ~n31383;
  assign n31385 = pi41  & ~n31384;
  assign n31386 = pi41  & n31383;
  assign n31387 = ~n31383 & ~n31384;
  assign n31388 = ~pi41  & ~n31383;
  assign n31389 = ~n43261 & ~n43262;
  assign n31390 = n894 & n9277;
  assign n31391 = pi106  & n37580;
  assign n31392 = pi108  & n896;
  assign n31393 = pi107  & n904;
  assign n31394 = ~n31392 & ~n31393;
  assign n31395 = ~n31391 & ~n31393;
  assign n31396 = ~n31392 & n31395;
  assign n31397 = ~n31391 & n31394;
  assign n31398 = ~n31390 & n43263;
  assign n31399 = pi50  & ~n31398;
  assign n31400 = pi50  & ~n31399;
  assign n31401 = pi50  & n31398;
  assign n31402 = ~n31398 & ~n31399;
  assign n31403 = ~pi50  & ~n31398;
  assign n31404 = ~n43264 & ~n43265;
  assign n31405 = ~n31176 & ~n31182;
  assign n31406 = n1971 & n8229;
  assign n31407 = pi103  & n37864;
  assign n31408 = pi105  & n1973;
  assign n31409 = pi104  & n1981;
  assign n31410 = ~n31408 & ~n31409;
  assign n31411 = ~n31407 & ~n31409;
  assign n31412 = ~n31408 & n31411;
  assign n31413 = ~n31407 & n31410;
  assign n31414 = ~n31406 & n43266;
  assign n31415 = pi53  & ~n31414;
  assign n31416 = pi53  & ~n31415;
  assign n31417 = pi53  & n31414;
  assign n31418 = ~n31414 & ~n31415;
  assign n31419 = ~pi53  & ~n31414;
  assign n31420 = ~n43267 & ~n43268;
  assign n31421 = n5578 & n7882;
  assign n31422 = pi97  & n39128;
  assign n31423 = pi99  & n7884;
  assign n31424 = pi98  & n7892;
  assign n31425 = ~n31423 & ~n31424;
  assign n31426 = ~n31422 & ~n31424;
  assign n31427 = ~n31423 & n31426;
  assign n31428 = ~n31422 & n31425;
  assign n31429 = ~n31421 & n43269;
  assign n31430 = pi59  & ~n31429;
  assign n31431 = pi59  & ~n31430;
  assign n31432 = pi59  & n31429;
  assign n31433 = ~n31429 & ~n31430;
  assign n31434 = ~pi59  & ~n31429;
  assign n31435 = ~n43270 & ~n43271;
  assign n31436 = n5281 & n12674;
  assign n31437 = pi94  & n40107;
  assign n31438 = pi96  & n12676;
  assign n31439 = pi95  & n12684;
  assign n31440 = ~n31438 & ~n31439;
  assign n31441 = ~n31437 & ~n31439;
  assign n31442 = ~n31438 & n31441;
  assign n31443 = ~n31437 & n31440;
  assign n31444 = ~n31436 & n43272;
  assign n31445 = pi62  & ~n31444;
  assign n31446 = pi62  & ~n31445;
  assign n31447 = pi62  & n31444;
  assign n31448 = ~n31444 & ~n31445;
  assign n31449 = ~pi62  & ~n31444;
  assign n31450 = ~n43273 & ~n43274;
  assign n31451 = ~n31117 & ~n31135;
  assign n31452 = pi93  & ~n40814;
  assign n31453 = pi92  & n18285;
  assign n31454 = ~n31452 & ~n31453;
  assign n31455 = n31115 & ~n31454;
  assign n31456 = ~n31115 & n31454;
  assign n31457 = ~n31455 & ~n31456;
  assign n31458 = ~n31451 & ~n31456;
  assign n31459 = ~n31455 & n31458;
  assign n31460 = ~n31451 & n31457;
  assign n31461 = n31451 & ~n31457;
  assign n31462 = ~n31451 & ~n43275;
  assign n31463 = ~n31456 & ~n43275;
  assign n31464 = ~n31455 & n31463;
  assign n31465 = ~n31462 & ~n31464;
  assign n31466 = ~n43275 & ~n31461;
  assign n31467 = ~n31450 & ~n43276;
  assign n31468 = n31450 & n43276;
  assign n31469 = n31450 & ~n43276;
  assign n31470 = ~n31450 & n43276;
  assign n31471 = ~n31469 & ~n31470;
  assign n31472 = ~n31467 & ~n31468;
  assign n31473 = ~n31435 & ~n43277;
  assign n31474 = n31435 & n43277;
  assign n31475 = ~n31473 & ~n31474;
  assign n31476 = ~n31140 & n31157;
  assign n31477 = ~n31140 & ~n31158;
  assign n31478 = ~n31141 & ~n31476;
  assign n31479 = n31475 & ~n43278;
  assign n31480 = ~n31475 & n43278;
  assign n31481 = ~n31479 & ~n31480;
  assign n31482 = n4312 & n6819;
  assign n31483 = pi100  & n38376;
  assign n31484 = pi102  & n4314;
  assign n31485 = pi101  & n4322;
  assign n31486 = ~n31484 & ~n31485;
  assign n31487 = ~n31483 & ~n31485;
  assign n31488 = ~n31484 & n31487;
  assign n31489 = ~n31483 & n31486;
  assign n31490 = ~n31482 & n43279;
  assign n31491 = pi56  & ~n31490;
  assign n31492 = pi56  & ~n31491;
  assign n31493 = pi56  & n31490;
  assign n31494 = ~n31490 & ~n31491;
  assign n31495 = ~pi56  & ~n31490;
  assign n31496 = ~n43280 & ~n43281;
  assign n31497 = n31481 & ~n31496;
  assign n31498 = ~n31481 & n31496;
  assign n31499 = n31481 & ~n31497;
  assign n31500 = ~n31496 & ~n31497;
  assign n31501 = ~n31499 & ~n31500;
  assign n31502 = ~n31497 & ~n31498;
  assign n31503 = n31110 & ~n31164;
  assign n31504 = ~n31164 & ~n31172;
  assign n31505 = ~n31165 & ~n31503;
  assign n31506 = ~n43282 & ~n43283;
  assign n31507 = n43282 & n43283;
  assign n31508 = ~n43282 & ~n31506;
  assign n31509 = ~n43283 & ~n31506;
  assign n31510 = ~n31508 & ~n31509;
  assign n31511 = ~n31506 & ~n31507;
  assign n31512 = n31420 & ~n43284;
  assign n31513 = ~n31420 & n43284;
  assign n31514 = ~n31420 & ~n43284;
  assign n31515 = n31420 & n43284;
  assign n31516 = ~n31514 & ~n31515;
  assign n31517 = ~n31512 & ~n31513;
  assign n31518 = ~n31405 & n43285;
  assign n31519 = n31405 & ~n43285;
  assign n31520 = ~n31518 & ~n31519;
  assign n31521 = ~n31404 & n31520;
  assign n31522 = n31404 & ~n31520;
  assign n31523 = ~n31521 & ~n31522;
  assign n31524 = ~n31187 & n31204;
  assign n31525 = ~n31187 & ~n31205;
  assign n31526 = ~n31188 & ~n31524;
  assign n31527 = n31523 & ~n43286;
  assign n31528 = ~n31523 & n43286;
  assign n31529 = ~n31527 & ~n31528;
  assign n31530 = n565 & n785;
  assign n31531 = pi109  & n37520;
  assign n31532 = pi111  & n787;
  assign n31533 = pi110  & n795;
  assign n31534 = ~n31532 & ~n31533;
  assign n31535 = ~n31531 & ~n31533;
  assign n31536 = ~n31532 & n31535;
  assign n31537 = ~n31531 & n31534;
  assign n31538 = ~n31530 & n43287;
  assign n31539 = pi47  & ~n31538;
  assign n31540 = pi47  & ~n31539;
  assign n31541 = pi47  & n31538;
  assign n31542 = ~n31538 & ~n31539;
  assign n31543 = ~pi47  & ~n31538;
  assign n31544 = ~n43288 & ~n43289;
  assign n31545 = n31529 & ~n31544;
  assign n31546 = ~n31529 & n31544;
  assign n31547 = n31529 & ~n31545;
  assign n31548 = ~n31544 & ~n31545;
  assign n31549 = ~n31547 & ~n31548;
  assign n31550 = ~n31545 & ~n31546;
  assign n31551 = ~n31212 & n31228;
  assign n31552 = ~n31212 & ~n31230;
  assign n31553 = ~n31211 & ~n31551;
  assign n31554 = n43290 & n43291;
  assign n31555 = ~n43290 & ~n43291;
  assign n31556 = ~n31554 & ~n31555;
  assign n31557 = n940 & n11258;
  assign n31558 = pi112  & n37541;
  assign n31559 = pi114  & n953;
  assign n31560 = pi113  & n955;
  assign n31561 = ~n31559 & ~n31560;
  assign n31562 = ~n31558 & ~n31560;
  assign n31563 = ~n31559 & n31562;
  assign n31564 = ~n31558 & n31561;
  assign n31565 = ~n31557 & n43292;
  assign n31566 = pi44  & ~n31565;
  assign n31567 = pi44  & ~n31566;
  assign n31568 = pi44  & n31565;
  assign n31569 = ~n31565 & ~n31566;
  assign n31570 = ~pi44  & ~n31565;
  assign n31571 = ~n43293 & ~n43294;
  assign n31572 = ~n31556 & n31571;
  assign n31573 = n31556 & ~n31571;
  assign n31574 = ~n31572 & ~n31573;
  assign n31575 = ~n31236 & n31252;
  assign n31576 = ~n31236 & ~n31253;
  assign n31577 = ~n31235 & ~n31575;
  assign n31578 = n31574 & ~n43295;
  assign n31579 = ~n31574 & n43295;
  assign n31580 = ~n43295 & ~n31578;
  assign n31581 = n31574 & ~n31578;
  assign n31582 = ~n31580 & ~n31581;
  assign n31583 = ~n31578 & ~n31579;
  assign n31584 = ~n31389 & ~n43296;
  assign n31585 = n31389 & ~n31581;
  assign n31586 = ~n31580 & n31585;
  assign n31587 = n31389 & n43296;
  assign n31588 = ~n31584 & ~n43297;
  assign n31589 = ~n31260 & n31276;
  assign n31590 = ~n31260 & ~n31278;
  assign n31591 = ~n31259 & ~n31589;
  assign n31592 = n31588 & ~n43298;
  assign n31593 = ~n31588 & n43298;
  assign n31594 = ~n31592 & ~n31593;
  assign n31595 = ~n31374 & n31594;
  assign n31596 = n31374 & ~n31594;
  assign n31597 = ~n31595 & ~n31596;
  assign n31598 = ~n31359 & n31597;
  assign n31599 = n31359 & ~n31597;
  assign n31600 = ~n31598 & ~n31599;
  assign n31601 = n2104 & n14961;
  assign n31602 = pi121  & n37758;
  assign n31603 = pi123  & n2117;
  assign n31604 = pi122  & n2119;
  assign n31605 = ~n31603 & ~n31604;
  assign n31606 = ~n31602 & ~n31604;
  assign n31607 = ~n31603 & n31606;
  assign n31608 = ~n31602 & n31605;
  assign n31609 = ~n31601 & n43299;
  assign n31610 = pi35  & ~n31609;
  assign n31611 = pi35  & ~n31610;
  assign n31612 = pi35  & n31609;
  assign n31613 = ~n31609 & ~n31610;
  assign n31614 = ~pi35  & ~n31609;
  assign n31615 = ~n43300 & ~n43301;
  assign n31616 = n31600 & ~n31615;
  assign n31617 = ~n31600 & n31615;
  assign n31618 = n31600 & ~n31616;
  assign n31619 = ~n31615 & ~n31616;
  assign n31620 = ~n31618 & ~n31619;
  assign n31621 = ~n31616 & ~n31617;
  assign n31622 = ~n31358 & n43302;
  assign n31623 = n31358 & ~n43302;
  assign n31624 = ~n31622 & ~n31623;
  assign n31625 = ~n31058 & ~n31316;
  assign n31626 = n607 & ~n18675;
  assign n31627 = ~n37489 & ~n31626;
  assign n31628 = pi127  & n37489;
  assign n31629 = n607 & n18680;
  assign n31630 = ~n31628 & ~n31629;
  assign n31631 = pi127  & ~n31627;
  assign n31632 = pi29  & ~n43303;
  assign n31633 = pi29  & ~n31632;
  assign n31634 = pi29  & n43303;
  assign n31635 = ~n43303 & ~n31632;
  assign n31636 = ~pi29  & ~n43303;
  assign n31637 = ~n43304 & ~n43305;
  assign n31638 = ~n31625 & ~n31637;
  assign n31639 = n31625 & n31637;
  assign n31640 = ~n31625 & ~n31638;
  assign n31641 = ~n31637 & ~n31638;
  assign n31642 = ~n31640 & ~n31641;
  assign n31643 = ~n31638 & ~n31639;
  assign n31644 = n31624 & ~n43306;
  assign n31645 = ~n31624 & n43306;
  assign n31646 = ~n31644 & ~n31645;
  assign n31647 = ~n31337 & n31646;
  assign n31648 = n31337 & ~n31646;
  assign n31649 = ~n31337 & ~n31647;
  assign n31650 = n31646 & ~n31647;
  assign n31651 = ~n31649 & ~n31650;
  assign n31652 = ~n31647 & ~n31648;
  assign n31653 = ~n31336 & ~n43307;
  assign n31654 = n31336 & ~n31650;
  assign n31655 = ~n31649 & n31654;
  assign n31656 = n31336 & n43307;
  assign po92  = ~n31653 & ~n43308;
  assign n31658 = ~n31647 & ~n31653;
  assign n31659 = ~n31638 & ~n31644;
  assign n31660 = ~n31592 & ~n31595;
  assign n31661 = ~n31578 & ~n31584;
  assign n31662 = n733 & n13057;
  assign n31663 = pi116  & n37510;
  assign n31664 = pi118  & n746;
  assign n31665 = pi117  & n748;
  assign n31666 = ~n31664 & ~n31665;
  assign n31667 = ~n31663 & ~n31665;
  assign n31668 = ~n31664 & n31667;
  assign n31669 = ~n31663 & n31666;
  assign n31670 = ~n31662 & n43309;
  assign n31671 = pi41  & ~n31670;
  assign n31672 = pi41  & ~n31671;
  assign n31673 = pi41  & n31670;
  assign n31674 = ~n31670 & ~n31671;
  assign n31675 = ~pi41  & ~n31670;
  assign n31676 = ~n43310 & ~n43311;
  assign n31677 = ~n31555 & ~n31573;
  assign n31678 = ~n31518 & ~n31521;
  assign n31679 = n894 & n9701;
  assign n31680 = pi107  & n37580;
  assign n31681 = pi109  & n896;
  assign n31682 = pi108  & n904;
  assign n31683 = ~n31681 & ~n31682;
  assign n31684 = ~n31680 & ~n31682;
  assign n31685 = ~n31681 & n31684;
  assign n31686 = ~n31680 & n31683;
  assign n31687 = ~n31679 & n43312;
  assign n31688 = pi50  & ~n31687;
  assign n31689 = pi50  & ~n31688;
  assign n31690 = pi50  & n31687;
  assign n31691 = ~n31687 & ~n31688;
  assign n31692 = ~pi50  & ~n31687;
  assign n31693 = ~n43313 & ~n43314;
  assign n31694 = ~n31467 & ~n31473;
  assign n31695 = n6474 & n7882;
  assign n31696 = pi98  & n39128;
  assign n31697 = pi100  & n7884;
  assign n31698 = pi99  & n7892;
  assign n31699 = ~n31697 & ~n31698;
  assign n31700 = ~n31696 & ~n31698;
  assign n31701 = ~n31697 & n31700;
  assign n31702 = ~n31696 & n31699;
  assign n31703 = ~n31695 & n43315;
  assign n31704 = pi59  & ~n31703;
  assign n31705 = pi59  & ~n31704;
  assign n31706 = pi59  & n31703;
  assign n31707 = ~n31703 & ~n31704;
  assign n31708 = ~pi59  & ~n31703;
  assign n31709 = ~n43316 & ~n43317;
  assign n31710 = n5630 & n12674;
  assign n31711 = pi95  & n40107;
  assign n31712 = pi97  & n12676;
  assign n31713 = pi96  & n12684;
  assign n31714 = ~n31712 & ~n31713;
  assign n31715 = ~n31711 & ~n31713;
  assign n31716 = ~n31712 & n31715;
  assign n31717 = ~n31711 & n31714;
  assign n31718 = ~n31710 & n43318;
  assign n31719 = pi62  & ~n31718;
  assign n31720 = pi62  & ~n31719;
  assign n31721 = pi62  & n31718;
  assign n31722 = ~n31718 & ~n31719;
  assign n31723 = ~pi62  & ~n31718;
  assign n31724 = ~n43319 & ~n43320;
  assign n31725 = pi94  & ~n40814;
  assign n31726 = pi93  & n18285;
  assign n31727 = ~n31725 & ~n31726;
  assign n31728 = ~pi29  & ~n31727;
  assign n31729 = pi29  & n31727;
  assign n31730 = ~n31728 & ~n31729;
  assign n31731 = n31454 & ~n31730;
  assign n31732 = ~n31454 & ~n31729;
  assign n31733 = ~n31728 & n31732;
  assign n31734 = ~n31454 & n31730;
  assign n31735 = ~n31454 & ~n43321;
  assign n31736 = n31730 & ~n43321;
  assign n31737 = ~n31735 & ~n31736;
  assign n31738 = ~n31731 & ~n43321;
  assign n31739 = ~n31463 & ~n43322;
  assign n31740 = n31463 & n43322;
  assign n31741 = ~n31463 & ~n31739;
  assign n31742 = ~n43322 & ~n31739;
  assign n31743 = ~n31741 & ~n31742;
  assign n31744 = ~n31739 & ~n31740;
  assign n31745 = ~n31724 & ~n43323;
  assign n31746 = n31724 & n43323;
  assign n31747 = n31724 & ~n43323;
  assign n31748 = ~n31724 & n43323;
  assign n31749 = ~n31747 & ~n31748;
  assign n31750 = ~n31745 & ~n31746;
  assign n31751 = ~n31709 & ~n43324;
  assign n31752 = n31709 & n43324;
  assign n31753 = ~n31751 & ~n31752;
  assign n31754 = ~n31694 & n31753;
  assign n31755 = n31694 & ~n31753;
  assign n31756 = ~n31754 & ~n31755;
  assign n31757 = n4312 & n6787;
  assign n31758 = pi101  & n38376;
  assign n31759 = pi103  & n4314;
  assign n31760 = pi102  & n4322;
  assign n31761 = ~n31759 & ~n31760;
  assign n31762 = ~n31758 & ~n31760;
  assign n31763 = ~n31759 & n31762;
  assign n31764 = ~n31758 & n31761;
  assign n31765 = ~n31757 & n43325;
  assign n31766 = pi56  & ~n31765;
  assign n31767 = pi56  & ~n31766;
  assign n31768 = pi56  & n31765;
  assign n31769 = ~n31765 & ~n31766;
  assign n31770 = ~pi56  & ~n31765;
  assign n31771 = ~n43326 & ~n43327;
  assign n31772 = n31756 & ~n31771;
  assign n31773 = ~n31756 & n31771;
  assign n31774 = n31756 & ~n31772;
  assign n31775 = n31756 & n31771;
  assign n31776 = ~n31771 & ~n31772;
  assign n31777 = ~n31756 & ~n31771;
  assign n31778 = ~n43328 & ~n43329;
  assign n31779 = ~n31772 & ~n31773;
  assign n31780 = ~n31479 & n31496;
  assign n31781 = ~n31479 & ~n31497;
  assign n31782 = ~n31480 & ~n31780;
  assign n31783 = n43330 & n43331;
  assign n31784 = ~n43330 & ~n43331;
  assign n31785 = ~n31783 & ~n31784;
  assign n31786 = n1971 & n8209;
  assign n31787 = pi104  & n37864;
  assign n31788 = pi106  & n1973;
  assign n31789 = pi105  & n1981;
  assign n31790 = ~n31788 & ~n31789;
  assign n31791 = ~n31787 & ~n31789;
  assign n31792 = ~n31788 & n31791;
  assign n31793 = ~n31787 & n31790;
  assign n31794 = ~n31786 & n43332;
  assign n31795 = pi53  & ~n31794;
  assign n31796 = pi53  & ~n31795;
  assign n31797 = pi53  & n31794;
  assign n31798 = ~n31794 & ~n31795;
  assign n31799 = ~pi53  & ~n31794;
  assign n31800 = ~n43333 & ~n43334;
  assign n31801 = n31785 & ~n31800;
  assign n31802 = ~n31785 & n31800;
  assign n31803 = n31785 & ~n31801;
  assign n31804 = n31785 & n31800;
  assign n31805 = ~n31800 & ~n31801;
  assign n31806 = ~n31785 & ~n31800;
  assign n31807 = ~n43335 & ~n43336;
  assign n31808 = ~n31801 & ~n31802;
  assign n31809 = n31420 & ~n31506;
  assign n31810 = ~n31506 & ~n31514;
  assign n31811 = ~n31507 & ~n31809;
  assign n31812 = ~n43337 & ~n43338;
  assign n31813 = n43337 & n43338;
  assign n31814 = n43337 & ~n43338;
  assign n31815 = ~n43337 & n43338;
  assign n31816 = ~n31814 & ~n31815;
  assign n31817 = ~n31812 & ~n31813;
  assign n31818 = ~n31693 & ~n43339;
  assign n31819 = n31693 & n43339;
  assign n31820 = ~n31818 & ~n31819;
  assign n31821 = n31678 & ~n31820;
  assign n31822 = ~n31678 & n31820;
  assign n31823 = ~n31821 & ~n31822;
  assign n31824 = n785 & n10844;
  assign n31825 = pi110  & n37520;
  assign n31826 = pi112  & n787;
  assign n31827 = pi111  & n795;
  assign n31828 = ~n31826 & ~n31827;
  assign n31829 = ~n31825 & ~n31827;
  assign n31830 = ~n31826 & n31829;
  assign n31831 = ~n31825 & n31828;
  assign n31832 = ~n31824 & n43340;
  assign n31833 = pi47  & ~n31832;
  assign n31834 = pi47  & ~n31833;
  assign n31835 = pi47  & n31832;
  assign n31836 = ~n31832 & ~n31833;
  assign n31837 = ~pi47  & ~n31832;
  assign n31838 = ~n43341 & ~n43342;
  assign n31839 = n31823 & ~n31838;
  assign n31840 = ~n31823 & n31838;
  assign n31841 = n31823 & ~n31839;
  assign n31842 = n31823 & n31838;
  assign n31843 = ~n31838 & ~n31839;
  assign n31844 = ~n31823 & ~n31838;
  assign n31845 = ~n43343 & ~n43344;
  assign n31846 = ~n31839 & ~n31840;
  assign n31847 = ~n31527 & n31544;
  assign n31848 = ~n31527 & ~n31545;
  assign n31849 = ~n31528 & ~n31847;
  assign n31850 = n43345 & n43346;
  assign n31851 = ~n43345 & ~n43346;
  assign n31852 = ~n31850 & ~n31851;
  assign n31853 = n523 & n940;
  assign n31854 = pi113  & n37541;
  assign n31855 = pi115  & n953;
  assign n31856 = pi114  & n955;
  assign n31857 = ~n31855 & ~n31856;
  assign n31858 = ~n31854 & ~n31856;
  assign n31859 = ~n31855 & n31858;
  assign n31860 = ~n31854 & n31857;
  assign n31861 = ~n31853 & n43347;
  assign n31862 = pi44  & ~n31861;
  assign n31863 = pi44  & ~n31862;
  assign n31864 = pi44  & n31861;
  assign n31865 = ~n31861 & ~n31862;
  assign n31866 = ~pi44  & ~n31861;
  assign n31867 = ~n43348 & ~n43349;
  assign n31868 = n31852 & ~n31867;
  assign n31869 = ~n31852 & n31867;
  assign n31870 = ~n31868 & ~n31869;
  assign n31871 = n31677 & ~n31870;
  assign n31872 = ~n31677 & ~n31869;
  assign n31873 = ~n31868 & n31872;
  assign n31874 = ~n31677 & ~n31868;
  assign n31875 = ~n31869 & n31874;
  assign n31876 = ~n31677 & n31870;
  assign n31877 = ~n31677 & ~n43350;
  assign n31878 = ~n31677 & ~n31870;
  assign n31879 = n31677 & ~n31868;
  assign n31880 = ~n31868 & ~n43350;
  assign n31881 = ~n31869 & ~n31879;
  assign n31882 = ~n31869 & n43352;
  assign n31883 = n31677 & n31870;
  assign n31884 = ~n43351 & ~n43353;
  assign n31885 = ~n31871 & ~n43350;
  assign n31886 = n31676 & n43354;
  assign n31887 = ~n31676 & ~n43354;
  assign n31888 = ~n31886 & ~n31887;
  assign n31889 = ~n31661 & n31888;
  assign n31890 = n31661 & ~n31888;
  assign n31891 = ~n31889 & ~n31890;
  assign n31892 = n691 & n15091;
  assign n31893 = pi119  & n37503;
  assign n31894 = pi121  & n704;
  assign n31895 = pi120  & n706;
  assign n31896 = ~n31894 & ~n31895;
  assign n31897 = ~n31893 & ~n31895;
  assign n31898 = ~n31894 & n31897;
  assign n31899 = ~n31893 & n31896;
  assign n31900 = ~n31892 & n43355;
  assign n31901 = pi38  & ~n31900;
  assign n31902 = pi38  & ~n31901;
  assign n31903 = pi38  & n31900;
  assign n31904 = ~n31900 & ~n31901;
  assign n31905 = ~pi38  & ~n31900;
  assign n31906 = ~n43356 & ~n43357;
  assign n31907 = n31891 & ~n31906;
  assign n31908 = ~n31891 & n31906;
  assign n31909 = n31891 & ~n31907;
  assign n31910 = n31891 & n31906;
  assign n31911 = ~n31906 & ~n31907;
  assign n31912 = ~n31891 & ~n31906;
  assign n31913 = ~n43358 & ~n43359;
  assign n31914 = ~n31907 & ~n31908;
  assign n31915 = n31660 & n43360;
  assign n31916 = ~n31660 & ~n43360;
  assign n31917 = ~n31915 & ~n31916;
  assign n31918 = n2104 & n15111;
  assign n31919 = pi122  & n37758;
  assign n31920 = pi124  & n2117;
  assign n31921 = pi123  & n2119;
  assign n31922 = ~n31920 & ~n31921;
  assign n31923 = ~n31919 & ~n31921;
  assign n31924 = ~n31920 & n31923;
  assign n31925 = ~n31919 & n31922;
  assign n31926 = ~n31918 & n43361;
  assign n31927 = pi35  & ~n31926;
  assign n31928 = pi35  & ~n31927;
  assign n31929 = pi35  & n31926;
  assign n31930 = ~n31926 & ~n31927;
  assign n31931 = ~pi35  & ~n31926;
  assign n31932 = ~n43362 & ~n43363;
  assign n31933 = n31917 & ~n31932;
  assign n31934 = ~n31917 & n31932;
  assign n31935 = n31917 & ~n31933;
  assign n31936 = n31917 & n31932;
  assign n31937 = ~n31932 & ~n31933;
  assign n31938 = ~n31917 & ~n31932;
  assign n31939 = ~n43364 & ~n43365;
  assign n31940 = ~n31933 & ~n31934;
  assign n31941 = ~n31598 & n31615;
  assign n31942 = ~n31598 & ~n31616;
  assign n31943 = ~n31599 & ~n31941;
  assign n31944 = n43366 & n43367;
  assign n31945 = ~n43366 & ~n43367;
  assign n31946 = ~n31944 & ~n31945;
  assign n31947 = ~n31357 & ~n31623;
  assign n31948 = n649 & n40885;
  assign n31949 = pi125  & n37496;
  assign n31950 = pi127  & n662;
  assign n31951 = pi126  & n664;
  assign n31952 = ~n31950 & ~n31951;
  assign n31953 = ~n31949 & ~n31951;
  assign n31954 = ~n31950 & n31953;
  assign n31955 = ~n31949 & n31952;
  assign n31956 = ~n31948 & n43368;
  assign n31957 = pi32  & ~n31956;
  assign n31958 = pi32  & ~n31957;
  assign n31959 = pi32  & n31956;
  assign n31960 = ~n31956 & ~n31957;
  assign n31961 = ~pi32  & ~n31956;
  assign n31962 = ~n43369 & ~n43370;
  assign n31963 = ~n31947 & ~n31962;
  assign n31964 = n31947 & n31962;
  assign n31965 = ~n31947 & ~n31963;
  assign n31966 = ~n31947 & n31962;
  assign n31967 = ~n31962 & ~n31963;
  assign n31968 = n31947 & ~n31962;
  assign n31969 = ~n43371 & ~n43372;
  assign n31970 = ~n31963 & ~n31964;
  assign n31971 = ~n31946 & n43373;
  assign n31972 = n31946 & ~n43373;
  assign n31973 = ~n31971 & ~n31972;
  assign n31974 = ~n31659 & n31973;
  assign n31975 = n31659 & ~n31973;
  assign n31976 = ~n31974 & ~n31975;
  assign n31977 = ~n31658 & n31976;
  assign n31978 = n31658 & ~n31976;
  assign po93  = ~n31977 & ~n31978;
  assign n31980 = ~n31974 & ~n31977;
  assign n31981 = ~n31963 & ~n31972;
  assign n31982 = ~n31933 & ~n31945;
  assign n31983 = n649 & n40891;
  assign n31984 = pi126  & n37496;
  assign n31985 = pi127  & n664;
  assign n31986 = ~n31984 & ~n31985;
  assign n31987 = ~n649 & n31986;
  assign n31988 = ~n40891 & n31986;
  assign n31989 = ~n31987 & ~n31988;
  assign n31990 = ~n31983 & n31986;
  assign n31991 = pi32  & ~n43374;
  assign n31992 = ~pi32  & n43374;
  assign n31993 = ~n31991 & ~n31992;
  assign n31994 = ~n31982 & ~n31993;
  assign n31995 = n31982 & n31993;
  assign n31996 = ~n31994 & ~n31995;
  assign n31997 = ~n31907 & ~n31916;
  assign n31998 = ~n31887 & ~n31889;
  assign n31999 = n733 & n13027;
  assign n32000 = pi117  & n37510;
  assign n32001 = pi119  & n746;
  assign n32002 = pi118  & n748;
  assign n32003 = ~n32001 & ~n32002;
  assign n32004 = ~n32000 & ~n32002;
  assign n32005 = ~n32001 & n32004;
  assign n32006 = ~n32000 & n32003;
  assign n32007 = ~n31999 & n43375;
  assign n32008 = pi41  & ~n32007;
  assign n32009 = pi41  & ~n32008;
  assign n32010 = pi41  & n32007;
  assign n32011 = ~n32007 & ~n32008;
  assign n32012 = ~pi41  & ~n32007;
  assign n32013 = ~n43376 & ~n43377;
  assign n32014 = ~n31839 & ~n31851;
  assign n32015 = ~n31818 & ~n31822;
  assign n32016 = ~n31801 & ~n31812;
  assign n32017 = ~n31772 & ~n31784;
  assign n32018 = n4312 & n8136;
  assign n32019 = pi102  & n38376;
  assign n32020 = pi104  & n4314;
  assign n32021 = pi103  & n4322;
  assign n32022 = ~n32020 & ~n32021;
  assign n32023 = ~n32019 & ~n32021;
  assign n32024 = ~n32020 & n32023;
  assign n32025 = ~n32019 & n32022;
  assign n32026 = ~n32018 & n43378;
  assign n32027 = pi56  & ~n32026;
  assign n32028 = pi56  & ~n32027;
  assign n32029 = pi56  & n32026;
  assign n32030 = ~n32026 & ~n32027;
  assign n32031 = ~pi56  & ~n32026;
  assign n32032 = ~n43379 & ~n43380;
  assign n32033 = ~n31751 & ~n31754;
  assign n32034 = n6839 & n7882;
  assign n32035 = pi99  & n39128;
  assign n32036 = pi101  & n7884;
  assign n32037 = pi100  & n7892;
  assign n32038 = ~n32036 & ~n32037;
  assign n32039 = ~n32035 & ~n32037;
  assign n32040 = ~n32036 & n32039;
  assign n32041 = ~n32035 & n32038;
  assign n32042 = ~n32034 & n43381;
  assign n32043 = pi59  & ~n32042;
  assign n32044 = pi59  & ~n32043;
  assign n32045 = pi59  & n32042;
  assign n32046 = ~n32042 & ~n32043;
  assign n32047 = ~pi59  & ~n32042;
  assign n32048 = ~n43382 & ~n43383;
  assign n32049 = ~n31739 & ~n31745;
  assign n32050 = ~n31728 & ~n43321;
  assign n32051 = ~n31728 & ~n31732;
  assign n32052 = pi95  & ~n40814;
  assign n32053 = pi94  & n18285;
  assign n32054 = ~n32052 & ~n32053;
  assign n32055 = n43384 & ~n32054;
  assign n32056 = ~n43384 & n32054;
  assign n32057 = ~n32055 & ~n32056;
  assign n32058 = n5610 & n12674;
  assign n32059 = pi96  & n40107;
  assign n32060 = pi98  & n12676;
  assign n32061 = pi97  & n12684;
  assign n32062 = ~n32060 & ~n32061;
  assign n32063 = ~n32059 & ~n32061;
  assign n32064 = ~n32060 & n32063;
  assign n32065 = ~n32059 & n32062;
  assign n32066 = ~n32058 & n43385;
  assign n32067 = pi62  & ~n32066;
  assign n32068 = pi62  & ~n32067;
  assign n32069 = pi62  & n32066;
  assign n32070 = ~n32066 & ~n32067;
  assign n32071 = ~pi62  & ~n32066;
  assign n32072 = ~n43386 & ~n43387;
  assign n32073 = ~n32057 & n32072;
  assign n32074 = n32057 & ~n32072;
  assign n32075 = ~n32073 & ~n32074;
  assign n32076 = ~n32049 & n32075;
  assign n32077 = n32049 & ~n32075;
  assign n32078 = ~n32049 & ~n32076;
  assign n32079 = n32075 & ~n32076;
  assign n32080 = ~n32078 & ~n32079;
  assign n32081 = ~n32076 & ~n32077;
  assign n32082 = ~n32048 & ~n43388;
  assign n32083 = n32048 & ~n32079;
  assign n32084 = ~n32078 & n32083;
  assign n32085 = n32048 & n43388;
  assign n32086 = ~n32082 & ~n43389;
  assign n32087 = ~n32033 & n32086;
  assign n32088 = n32033 & ~n32086;
  assign n32089 = ~n32033 & ~n32087;
  assign n32090 = n32086 & ~n32087;
  assign n32091 = ~n32089 & ~n32090;
  assign n32092 = ~n32087 & ~n32088;
  assign n32093 = ~n32032 & ~n43390;
  assign n32094 = n32032 & ~n32090;
  assign n32095 = ~n32089 & n32094;
  assign n32096 = n32032 & n43390;
  assign n32097 = ~n32093 & ~n43391;
  assign n32098 = ~n32017 & n32097;
  assign n32099 = n32017 & ~n32097;
  assign n32100 = ~n32098 & ~n32099;
  assign n32101 = n1971 & n8177;
  assign n32102 = pi105  & n37864;
  assign n32103 = pi107  & n1973;
  assign n32104 = pi106  & n1981;
  assign n32105 = ~n32103 & ~n32104;
  assign n32106 = ~n32102 & ~n32104;
  assign n32107 = ~n32103 & n32106;
  assign n32108 = ~n32102 & n32105;
  assign n32109 = ~n32101 & n43392;
  assign n32110 = pi53  & ~n32109;
  assign n32111 = pi53  & ~n32110;
  assign n32112 = pi53  & n32109;
  assign n32113 = ~n32109 & ~n32110;
  assign n32114 = ~pi53  & ~n32109;
  assign n32115 = ~n43393 & ~n43394;
  assign n32116 = n32100 & ~n32115;
  assign n32117 = ~n32100 & n32115;
  assign n32118 = n32100 & ~n32116;
  assign n32119 = ~n32115 & ~n32116;
  assign n32120 = ~n32118 & ~n32119;
  assign n32121 = ~n32116 & ~n32117;
  assign n32122 = n32016 & n43395;
  assign n32123 = ~n32016 & ~n43395;
  assign n32124 = ~n32122 & ~n32123;
  assign n32125 = n894 & n9678;
  assign n32126 = pi108  & n37580;
  assign n32127 = pi110  & n896;
  assign n32128 = pi109  & n904;
  assign n32129 = ~n32127 & ~n32128;
  assign n32130 = ~n32126 & ~n32128;
  assign n32131 = ~n32127 & n32130;
  assign n32132 = ~n32126 & n32129;
  assign n32133 = ~n32125 & n43396;
  assign n32134 = pi50  & ~n32133;
  assign n32135 = pi50  & ~n32134;
  assign n32136 = pi50  & n32133;
  assign n32137 = ~n32133 & ~n32134;
  assign n32138 = ~pi50  & ~n32133;
  assign n32139 = ~n43397 & ~n43398;
  assign n32140 = ~n32124 & n32139;
  assign n32141 = n32124 & ~n32139;
  assign n32142 = n32124 & ~n32141;
  assign n32143 = ~n32139 & ~n32141;
  assign n32144 = ~n32142 & ~n32143;
  assign n32145 = ~n32140 & ~n32141;
  assign n32146 = n32015 & n43399;
  assign n32147 = ~n32015 & ~n43399;
  assign n32148 = ~n32146 & ~n32147;
  assign n32149 = n785 & n11276;
  assign n32150 = pi111  & n37520;
  assign n32151 = pi113  & n787;
  assign n32152 = pi112  & n795;
  assign n32153 = ~n32151 & ~n32152;
  assign n32154 = ~n32150 & ~n32152;
  assign n32155 = ~n32151 & n32154;
  assign n32156 = ~n32150 & n32153;
  assign n32157 = ~n32149 & n43400;
  assign n32158 = pi47  & ~n32157;
  assign n32159 = pi47  & ~n32158;
  assign n32160 = pi47  & n32157;
  assign n32161 = ~n32157 & ~n32158;
  assign n32162 = ~pi47  & ~n32157;
  assign n32163 = ~n43401 & ~n43402;
  assign n32164 = n32148 & ~n32163;
  assign n32165 = ~n32148 & n32163;
  assign n32166 = n32148 & ~n32164;
  assign n32167 = ~n32163 & ~n32164;
  assign n32168 = ~n32166 & ~n32167;
  assign n32169 = ~n32164 & ~n32165;
  assign n32170 = n32014 & n43403;
  assign n32171 = ~n32014 & ~n43403;
  assign n32172 = ~n32170 & ~n32171;
  assign n32173 = n940 & n12530;
  assign n32174 = pi114  & n37541;
  assign n32175 = pi116  & n953;
  assign n32176 = pi115  & n955;
  assign n32177 = ~n32175 & ~n32176;
  assign n32178 = ~n32174 & ~n32176;
  assign n32179 = ~n32175 & n32178;
  assign n32180 = ~n32174 & n32177;
  assign n32181 = ~n32173 & n43404;
  assign n32182 = pi44  & ~n32181;
  assign n32183 = pi44  & ~n32182;
  assign n32184 = pi44  & n32181;
  assign n32185 = ~n32181 & ~n32182;
  assign n32186 = ~pi44  & ~n32181;
  assign n32187 = ~n43405 & ~n43406;
  assign n32188 = ~n32172 & n32187;
  assign n32189 = n32172 & ~n32187;
  assign n32190 = n32172 & ~n32189;
  assign n32191 = ~n32187 & ~n32189;
  assign n32192 = ~n32190 & ~n32191;
  assign n32193 = ~n32188 & ~n32189;
  assign n32194 = ~n43352 & ~n43407;
  assign n32195 = n43352 & n43407;
  assign n32196 = ~n43352 & n43407;
  assign n32197 = n43352 & ~n43407;
  assign n32198 = ~n32196 & ~n32197;
  assign n32199 = ~n32194 & ~n32195;
  assign n32200 = ~n32013 & ~n43408;
  assign n32201 = n32013 & n43408;
  assign n32202 = ~n32200 & ~n32201;
  assign n32203 = ~n31998 & n32202;
  assign n32204 = n31998 & ~n32202;
  assign n32205 = ~n32203 & ~n32204;
  assign n32206 = n691 & n15049;
  assign n32207 = pi120  & n37503;
  assign n32208 = pi122  & n704;
  assign n32209 = pi121  & n706;
  assign n32210 = ~n32208 & ~n32209;
  assign n32211 = ~n32207 & ~n32209;
  assign n32212 = ~n32208 & n32211;
  assign n32213 = ~n32207 & n32210;
  assign n32214 = ~n32206 & n43409;
  assign n32215 = pi38  & ~n32214;
  assign n32216 = pi38  & ~n32215;
  assign n32217 = pi38  & n32214;
  assign n32218 = ~n32214 & ~n32215;
  assign n32219 = ~pi38  & ~n32214;
  assign n32220 = ~n43410 & ~n43411;
  assign n32221 = n32205 & ~n32220;
  assign n32222 = ~n32205 & n32220;
  assign n32223 = n32205 & ~n32221;
  assign n32224 = ~n32220 & ~n32221;
  assign n32225 = ~n32223 & ~n32224;
  assign n32226 = ~n32221 & ~n32222;
  assign n32227 = n31997 & n43412;
  assign n32228 = ~n31997 & ~n43412;
  assign n32229 = ~n32227 & ~n32228;
  assign n32230 = n2104 & n15068;
  assign n32231 = pi123  & n37758;
  assign n32232 = pi125  & n2117;
  assign n32233 = pi124  & n2119;
  assign n32234 = ~n32232 & ~n32233;
  assign n32235 = ~n32231 & ~n32233;
  assign n32236 = ~n32232 & n32235;
  assign n32237 = ~n32231 & n32234;
  assign n32238 = ~n32230 & n43413;
  assign n32239 = pi35  & ~n32238;
  assign n32240 = pi35  & ~n32239;
  assign n32241 = pi35  & n32238;
  assign n32242 = ~n32238 & ~n32239;
  assign n32243 = ~pi35  & ~n32238;
  assign n32244 = ~n43414 & ~n43415;
  assign n32245 = n32229 & ~n32244;
  assign n32246 = ~n32229 & n32244;
  assign n32247 = ~n32245 & ~n32246;
  assign n32248 = n31996 & ~n32246;
  assign n32249 = ~n32245 & n32248;
  assign n32250 = n31996 & n32247;
  assign n32251 = ~n31996 & ~n32247;
  assign n32252 = n31996 & ~n43416;
  assign n32253 = ~n32246 & ~n43416;
  assign n32254 = ~n32245 & n32253;
  assign n32255 = n32247 & ~n43416;
  assign n32256 = ~n32252 & ~n43417;
  assign n32257 = ~n43416 & ~n32251;
  assign n32258 = ~n31981 & ~n43418;
  assign n32259 = n31981 & n43418;
  assign n32260 = ~n43418 & ~n32258;
  assign n32261 = ~n31981 & ~n32258;
  assign n32262 = ~n32260 & ~n32261;
  assign n32263 = ~n32258 & ~n32259;
  assign n32264 = ~n31980 & ~n43419;
  assign n32265 = n31980 & n43419;
  assign po94  = ~n32264 & ~n32265;
  assign n32267 = ~n32258 & ~n32264;
  assign n32268 = ~n31994 & ~n43416;
  assign n32269 = ~n32228 & ~n32245;
  assign n32270 = n649 & ~n18675;
  assign n32271 = ~n37496 & ~n32270;
  assign n32272 = pi127  & n37496;
  assign n32273 = n649 & n18680;
  assign n32274 = ~n32272 & ~n32273;
  assign n32275 = pi127  & ~n32271;
  assign n32276 = pi32  & ~n43420;
  assign n32277 = pi32  & ~n32276;
  assign n32278 = pi32  & n43420;
  assign n32279 = ~n43420 & ~n32276;
  assign n32280 = ~pi32  & ~n43420;
  assign n32281 = ~n43421 & ~n43422;
  assign n32282 = ~n32269 & ~n32281;
  assign n32283 = n32269 & n32281;
  assign n32284 = ~n32269 & ~n32282;
  assign n32285 = ~n32281 & ~n32282;
  assign n32286 = ~n32284 & ~n32285;
  assign n32287 = ~n32282 & ~n32283;
  assign n32288 = ~n32194 & ~n32200;
  assign n32289 = n733 & n14913;
  assign n32290 = pi118  & n37510;
  assign n32291 = pi120  & n746;
  assign n32292 = pi119  & n748;
  assign n32293 = ~n32291 & ~n32292;
  assign n32294 = ~n32290 & ~n32292;
  assign n32295 = ~n32291 & n32294;
  assign n32296 = ~n32290 & n32293;
  assign n32297 = ~n32289 & n43424;
  assign n32298 = pi41  & ~n32297;
  assign n32299 = pi41  & ~n32298;
  assign n32300 = pi41  & n32297;
  assign n32301 = ~n32297 & ~n32298;
  assign n32302 = ~pi41  & ~n32297;
  assign n32303 = ~n43425 & ~n43426;
  assign n32304 = n940 & n13079;
  assign n32305 = pi115  & n37541;
  assign n32306 = pi117  & n953;
  assign n32307 = pi116  & n955;
  assign n32308 = ~n32306 & ~n32307;
  assign n32309 = ~n32305 & ~n32307;
  assign n32310 = ~n32306 & n32309;
  assign n32311 = ~n32305 & n32308;
  assign n32312 = ~n32304 & n43427;
  assign n32313 = pi44  & ~n32312;
  assign n32314 = pi44  & ~n32313;
  assign n32315 = pi44  & n32312;
  assign n32316 = ~n32312 & ~n32313;
  assign n32317 = ~pi44  & ~n32312;
  assign n32318 = ~n43428 & ~n43429;
  assign n32319 = n1971 & n9277;
  assign n32320 = pi106  & n37864;
  assign n32321 = pi108  & n1973;
  assign n32322 = pi107  & n1981;
  assign n32323 = ~n32321 & ~n32322;
  assign n32324 = ~n32320 & ~n32322;
  assign n32325 = ~n32321 & n32324;
  assign n32326 = ~n32320 & n32323;
  assign n32327 = ~n32319 & n43430;
  assign n32328 = pi53  & ~n32327;
  assign n32329 = pi53  & ~n32328;
  assign n32330 = pi53  & n32327;
  assign n32331 = ~n32327 & ~n32328;
  assign n32332 = ~pi53  & ~n32327;
  assign n32333 = ~n43431 & ~n43432;
  assign n32334 = ~n32087 & ~n32093;
  assign n32335 = n4312 & n8229;
  assign n32336 = pi103  & n38376;
  assign n32337 = pi105  & n4314;
  assign n32338 = pi104  & n4322;
  assign n32339 = ~n32337 & ~n32338;
  assign n32340 = ~n32336 & ~n32338;
  assign n32341 = ~n32337 & n32340;
  assign n32342 = ~n32336 & n32339;
  assign n32343 = ~n32335 & n43433;
  assign n32344 = pi56  & ~n32343;
  assign n32345 = pi56  & ~n32344;
  assign n32346 = pi56  & n32343;
  assign n32347 = ~n32343 & ~n32344;
  assign n32348 = ~pi56  & ~n32343;
  assign n32349 = ~n43434 & ~n43435;
  assign n32350 = ~n32076 & ~n32082;
  assign n32351 = n6819 & n7882;
  assign n32352 = pi100  & n39128;
  assign n32353 = pi102  & n7884;
  assign n32354 = pi101  & n7892;
  assign n32355 = ~n32353 & ~n32354;
  assign n32356 = ~n32352 & ~n32354;
  assign n32357 = ~n32353 & n32356;
  assign n32358 = ~n32352 & n32355;
  assign n32359 = ~n32351 & n43436;
  assign n32360 = pi59  & ~n32359;
  assign n32361 = pi59  & ~n32360;
  assign n32362 = pi59  & n32359;
  assign n32363 = ~n32359 & ~n32360;
  assign n32364 = ~pi59  & ~n32359;
  assign n32365 = ~n43437 & ~n43438;
  assign n32366 = n5578 & n12674;
  assign n32367 = pi97  & n40107;
  assign n32368 = pi99  & n12676;
  assign n32369 = pi98  & n12684;
  assign n32370 = ~n32368 & ~n32369;
  assign n32371 = ~n32367 & ~n32369;
  assign n32372 = ~n32368 & n32371;
  assign n32373 = ~n32367 & n32370;
  assign n32374 = ~n32366 & n43439;
  assign n32375 = pi62  & ~n32374;
  assign n32376 = pi62  & ~n32375;
  assign n32377 = pi62  & n32374;
  assign n32378 = ~n32374 & ~n32375;
  assign n32379 = ~pi62  & ~n32374;
  assign n32380 = ~n43440 & ~n43441;
  assign n32381 = ~n32056 & ~n32074;
  assign n32382 = pi96  & ~n40814;
  assign n32383 = pi95  & n18285;
  assign n32384 = ~n32382 & ~n32383;
  assign n32385 = ~n32054 & n32384;
  assign n32386 = n32054 & ~n32384;
  assign n32387 = ~n32385 & ~n32386;
  assign n32388 = ~n32381 & ~n32386;
  assign n32389 = ~n32385 & n32388;
  assign n32390 = ~n32381 & n32387;
  assign n32391 = n32381 & ~n32387;
  assign n32392 = ~n32381 & ~n43442;
  assign n32393 = ~n32385 & ~n43442;
  assign n32394 = ~n32386 & n32393;
  assign n32395 = ~n32392 & ~n32394;
  assign n32396 = ~n43442 & ~n32391;
  assign n32397 = ~n32380 & ~n43443;
  assign n32398 = n32380 & n43443;
  assign n32399 = ~n43443 & ~n32397;
  assign n32400 = n32380 & ~n43443;
  assign n32401 = ~n32380 & ~n32397;
  assign n32402 = ~n32380 & n43443;
  assign n32403 = ~n43444 & ~n43445;
  assign n32404 = ~n32397 & ~n32398;
  assign n32405 = ~n32365 & ~n43446;
  assign n32406 = n32365 & n43446;
  assign n32407 = n32365 & ~n43446;
  assign n32408 = ~n32365 & n43446;
  assign n32409 = ~n32407 & ~n32408;
  assign n32410 = ~n32405 & ~n32406;
  assign n32411 = ~n32350 & ~n43447;
  assign n32412 = n32350 & n43447;
  assign n32413 = ~n32411 & ~n32412;
  assign n32414 = ~n32349 & n32413;
  assign n32415 = n32349 & ~n32413;
  assign n32416 = ~n32414 & ~n32415;
  assign n32417 = ~n32334 & n32416;
  assign n32418 = n32334 & ~n32416;
  assign n32419 = ~n32417 & ~n32418;
  assign n32420 = ~n32333 & n32419;
  assign n32421 = n32333 & ~n32419;
  assign n32422 = ~n32420 & ~n32421;
  assign n32423 = ~n32098 & n32115;
  assign n32424 = ~n32098 & ~n32116;
  assign n32425 = ~n32099 & ~n32423;
  assign n32426 = n32422 & ~n43448;
  assign n32427 = ~n32422 & n43448;
  assign n32428 = ~n32426 & ~n32427;
  assign n32429 = n565 & n894;
  assign n32430 = pi109  & n37580;
  assign n32431 = pi111  & n896;
  assign n32432 = pi110  & n904;
  assign n32433 = ~n32431 & ~n32432;
  assign n32434 = ~n32430 & ~n32432;
  assign n32435 = ~n32431 & n32434;
  assign n32436 = ~n32430 & n32433;
  assign n32437 = ~n32429 & n43449;
  assign n32438 = pi50  & ~n32437;
  assign n32439 = pi50  & ~n32438;
  assign n32440 = pi50  & n32437;
  assign n32441 = ~n32437 & ~n32438;
  assign n32442 = ~pi50  & ~n32437;
  assign n32443 = ~n43450 & ~n43451;
  assign n32444 = n32428 & ~n32443;
  assign n32445 = ~n32428 & n32443;
  assign n32446 = n32428 & ~n32444;
  assign n32447 = ~n32443 & ~n32444;
  assign n32448 = ~n32446 & ~n32447;
  assign n32449 = ~n32444 & ~n32445;
  assign n32450 = ~n32123 & n32139;
  assign n32451 = ~n32123 & ~n32141;
  assign n32452 = ~n32122 & ~n32450;
  assign n32453 = n43452 & n43453;
  assign n32454 = ~n43452 & ~n43453;
  assign n32455 = ~n32453 & ~n32454;
  assign n32456 = n785 & n11258;
  assign n32457 = pi112  & n37520;
  assign n32458 = pi114  & n787;
  assign n32459 = pi113  & n795;
  assign n32460 = ~n32458 & ~n32459;
  assign n32461 = ~n32457 & ~n32459;
  assign n32462 = ~n32458 & n32461;
  assign n32463 = ~n32457 & n32460;
  assign n32464 = ~n32456 & n43454;
  assign n32465 = pi47  & ~n32464;
  assign n32466 = pi47  & ~n32465;
  assign n32467 = pi47  & n32464;
  assign n32468 = ~n32464 & ~n32465;
  assign n32469 = ~pi47  & ~n32464;
  assign n32470 = ~n43455 & ~n43456;
  assign n32471 = ~n32455 & n32470;
  assign n32472 = n32455 & ~n32470;
  assign n32473 = ~n32471 & ~n32472;
  assign n32474 = ~n32147 & n32163;
  assign n32475 = ~n32147 & ~n32164;
  assign n32476 = ~n32146 & ~n32474;
  assign n32477 = n32473 & ~n43457;
  assign n32478 = ~n32473 & n43457;
  assign n32479 = ~n43457 & ~n32477;
  assign n32480 = n32473 & ~n32477;
  assign n32481 = ~n32479 & ~n32480;
  assign n32482 = ~n32477 & ~n32478;
  assign n32483 = ~n32318 & ~n43458;
  assign n32484 = n32318 & ~n32480;
  assign n32485 = ~n32479 & n32484;
  assign n32486 = n32318 & n43458;
  assign n32487 = ~n32483 & ~n43459;
  assign n32488 = ~n32171 & n32187;
  assign n32489 = ~n32171 & ~n32189;
  assign n32490 = ~n32170 & ~n32488;
  assign n32491 = n32487 & ~n43460;
  assign n32492 = ~n32487 & n43460;
  assign n32493 = ~n32491 & ~n32492;
  assign n32494 = ~n32303 & n32493;
  assign n32495 = n32303 & ~n32493;
  assign n32496 = ~n32494 & ~n32495;
  assign n32497 = ~n32288 & n32496;
  assign n32498 = n32288 & ~n32496;
  assign n32499 = ~n32497 & ~n32498;
  assign n32500 = n691 & n14961;
  assign n32501 = pi121  & n37503;
  assign n32502 = pi123  & n704;
  assign n32503 = pi122  & n706;
  assign n32504 = ~n32502 & ~n32503;
  assign n32505 = ~n32501 & ~n32503;
  assign n32506 = ~n32502 & n32505;
  assign n32507 = ~n32501 & n32504;
  assign n32508 = ~n32500 & n43461;
  assign n32509 = pi38  & ~n32508;
  assign n32510 = pi38  & ~n32509;
  assign n32511 = pi38  & n32508;
  assign n32512 = ~n32508 & ~n32509;
  assign n32513 = ~pi38  & ~n32508;
  assign n32514 = ~n43462 & ~n43463;
  assign n32515 = n32499 & ~n32514;
  assign n32516 = ~n32499 & n32514;
  assign n32517 = n32499 & ~n32515;
  assign n32518 = ~n32514 & ~n32515;
  assign n32519 = ~n32517 & ~n32518;
  assign n32520 = ~n32515 & ~n32516;
  assign n32521 = ~n32203 & n32220;
  assign n32522 = ~n32203 & ~n32221;
  assign n32523 = ~n32204 & ~n32521;
  assign n32524 = n43464 & n43465;
  assign n32525 = ~n43464 & ~n43465;
  assign n32526 = ~n32524 & ~n32525;
  assign n32527 = n2104 & n15021;
  assign n32528 = pi124  & n37758;
  assign n32529 = pi126  & n2117;
  assign n32530 = pi125  & n2119;
  assign n32531 = ~n32529 & ~n32530;
  assign n32532 = ~n32528 & ~n32530;
  assign n32533 = ~n32529 & n32532;
  assign n32534 = ~n32528 & n32531;
  assign n32535 = ~n32527 & n43466;
  assign n32536 = pi35  & ~n32535;
  assign n32537 = pi35  & ~n32536;
  assign n32538 = pi35  & n32535;
  assign n32539 = ~n32535 & ~n32536;
  assign n32540 = ~pi35  & ~n32535;
  assign n32541 = ~n43467 & ~n43468;
  assign n32542 = ~n32526 & n32541;
  assign n32543 = n32526 & ~n32541;
  assign n32544 = n32526 & ~n32543;
  assign n32545 = ~n32541 & ~n32543;
  assign n32546 = ~n32544 & ~n32545;
  assign n32547 = ~n32542 & ~n32543;
  assign n32548 = ~n43423 & ~n43469;
  assign n32549 = n43423 & n43469;
  assign n32550 = ~n43423 & n43469;
  assign n32551 = n43423 & ~n43469;
  assign n32552 = ~n32550 & ~n32551;
  assign n32553 = ~n32548 & ~n32549;
  assign n32554 = ~n32268 & ~n43470;
  assign n32555 = n32268 & n43470;
  assign n32556 = ~n32268 & ~n32554;
  assign n32557 = ~n43470 & ~n32554;
  assign n32558 = ~n32556 & ~n32557;
  assign n32559 = ~n32554 & ~n32555;
  assign n32560 = ~n32267 & ~n43471;
  assign n32561 = n32267 & ~n32557;
  assign n32562 = ~n32556 & n32561;
  assign n32563 = n32267 & n43471;
  assign po95  = ~n32560 & ~n43472;
  assign n32565 = ~n32554 & ~n32560;
  assign n32566 = ~n32491 & ~n32494;
  assign n32567 = ~n32477 & ~n32483;
  assign n32568 = n940 & n13057;
  assign n32569 = pi116  & n37541;
  assign n32570 = pi118  & n953;
  assign n32571 = pi117  & n955;
  assign n32572 = ~n32570 & ~n32571;
  assign n32573 = ~n32569 & ~n32571;
  assign n32574 = ~n32570 & n32573;
  assign n32575 = ~n32569 & n32572;
  assign n32576 = ~n32568 & n43473;
  assign n32577 = pi44  & ~n32576;
  assign n32578 = pi44  & ~n32577;
  assign n32579 = pi44  & n32576;
  assign n32580 = ~n32576 & ~n32577;
  assign n32581 = ~pi44  & ~n32576;
  assign n32582 = ~n43474 & ~n43475;
  assign n32583 = ~n32454 & ~n32472;
  assign n32584 = ~n32417 & ~n32420;
  assign n32585 = ~n32411 & ~n32414;
  assign n32586 = ~n32397 & ~n32405;
  assign n32587 = n6787 & n7882;
  assign n32588 = pi101  & n39128;
  assign n32589 = pi103  & n7884;
  assign n32590 = pi102  & n7892;
  assign n32591 = ~n32589 & ~n32590;
  assign n32592 = ~n32588 & ~n32590;
  assign n32593 = ~n32589 & n32592;
  assign n32594 = ~n32588 & n32591;
  assign n32595 = ~n32587 & n43476;
  assign n32596 = pi59  & ~n32595;
  assign n32597 = pi59  & ~n32596;
  assign n32598 = pi59  & n32595;
  assign n32599 = ~n32595 & ~n32596;
  assign n32600 = ~pi59  & ~n32595;
  assign n32601 = ~n43477 & ~n43478;
  assign n32602 = n6474 & n12674;
  assign n32603 = pi98  & n40107;
  assign n32604 = pi100  & n12676;
  assign n32605 = pi99  & n12684;
  assign n32606 = ~n32604 & ~n32605;
  assign n32607 = ~n32603 & ~n32605;
  assign n32608 = ~n32604 & n32607;
  assign n32609 = ~n32603 & n32606;
  assign n32610 = ~n32602 & n43479;
  assign n32611 = pi62  & ~n32610;
  assign n32612 = pi62  & ~n32611;
  assign n32613 = pi62  & n32610;
  assign n32614 = ~n32610 & ~n32611;
  assign n32615 = ~pi62  & ~n32610;
  assign n32616 = ~n43480 & ~n43481;
  assign n32617 = pi97  & ~n40814;
  assign n32618 = pi96  & n18285;
  assign n32619 = ~n32617 & ~n32618;
  assign n32620 = ~pi32  & ~n32619;
  assign n32621 = pi32  & n32619;
  assign n32622 = ~n32620 & ~n32621;
  assign n32623 = n32384 & ~n32622;
  assign n32624 = ~n32384 & ~n32621;
  assign n32625 = ~n32620 & n32624;
  assign n32626 = ~n32384 & n32622;
  assign n32627 = ~n32384 & ~n43482;
  assign n32628 = n32622 & ~n43482;
  assign n32629 = ~n32627 & ~n32628;
  assign n32630 = ~n32623 & ~n43482;
  assign n32631 = ~n32393 & ~n43483;
  assign n32632 = n32393 & n43483;
  assign n32633 = ~n32393 & ~n32631;
  assign n32634 = ~n43483 & ~n32631;
  assign n32635 = ~n32633 & ~n32634;
  assign n32636 = ~n32631 & ~n32632;
  assign n32637 = ~n32616 & ~n43484;
  assign n32638 = n32616 & n43484;
  assign n32639 = n32616 & ~n43484;
  assign n32640 = ~n32616 & n43484;
  assign n32641 = ~n32639 & ~n32640;
  assign n32642 = ~n32637 & ~n32638;
  assign n32643 = ~n32601 & ~n43485;
  assign n32644 = n32601 & n43485;
  assign n32645 = ~n32643 & ~n32644;
  assign n32646 = ~n32586 & n32645;
  assign n32647 = n32586 & ~n32645;
  assign n32648 = ~n32646 & ~n32647;
  assign n32649 = n4312 & n8209;
  assign n32650 = pi104  & n38376;
  assign n32651 = pi106  & n4314;
  assign n32652 = pi105  & n4322;
  assign n32653 = ~n32651 & ~n32652;
  assign n32654 = ~n32650 & ~n32652;
  assign n32655 = ~n32651 & n32654;
  assign n32656 = ~n32650 & n32653;
  assign n32657 = ~n32649 & n43486;
  assign n32658 = pi56  & ~n32657;
  assign n32659 = pi56  & ~n32658;
  assign n32660 = pi56  & n32657;
  assign n32661 = ~n32657 & ~n32658;
  assign n32662 = ~pi56  & ~n32657;
  assign n32663 = ~n43487 & ~n43488;
  assign n32664 = n32648 & ~n32663;
  assign n32665 = ~n32648 & n32663;
  assign n32666 = n32648 & ~n32664;
  assign n32667 = n32648 & n32663;
  assign n32668 = ~n32663 & ~n32664;
  assign n32669 = ~n32648 & ~n32663;
  assign n32670 = ~n43489 & ~n43490;
  assign n32671 = ~n32664 & ~n32665;
  assign n32672 = n32585 & n43491;
  assign n32673 = ~n32585 & ~n43491;
  assign n32674 = ~n32672 & ~n32673;
  assign n32675 = n1971 & n9701;
  assign n32676 = pi107  & n37864;
  assign n32677 = pi109  & n1973;
  assign n32678 = pi108  & n1981;
  assign n32679 = ~n32677 & ~n32678;
  assign n32680 = ~n32676 & ~n32678;
  assign n32681 = ~n32677 & n32680;
  assign n32682 = ~n32676 & n32679;
  assign n32683 = ~n32675 & n43492;
  assign n32684 = pi53  & ~n32683;
  assign n32685 = pi53  & ~n32684;
  assign n32686 = pi53  & n32683;
  assign n32687 = ~n32683 & ~n32684;
  assign n32688 = ~pi53  & ~n32683;
  assign n32689 = ~n43493 & ~n43494;
  assign n32690 = n32674 & ~n32689;
  assign n32691 = ~n32674 & n32689;
  assign n32692 = n32674 & ~n32690;
  assign n32693 = n32674 & n32689;
  assign n32694 = ~n32689 & ~n32690;
  assign n32695 = ~n32674 & ~n32689;
  assign n32696 = ~n43495 & ~n43496;
  assign n32697 = ~n32690 & ~n32691;
  assign n32698 = n32584 & n43497;
  assign n32699 = ~n32584 & ~n43497;
  assign n32700 = ~n32698 & ~n32699;
  assign n32701 = n894 & n10844;
  assign n32702 = pi110  & n37580;
  assign n32703 = pi112  & n896;
  assign n32704 = pi111  & n904;
  assign n32705 = ~n32703 & ~n32704;
  assign n32706 = ~n32702 & ~n32704;
  assign n32707 = ~n32703 & n32706;
  assign n32708 = ~n32702 & n32705;
  assign n32709 = ~n32701 & n43498;
  assign n32710 = pi50  & ~n32709;
  assign n32711 = pi50  & ~n32710;
  assign n32712 = pi50  & n32709;
  assign n32713 = ~n32709 & ~n32710;
  assign n32714 = ~pi50  & ~n32709;
  assign n32715 = ~n43499 & ~n43500;
  assign n32716 = n32700 & ~n32715;
  assign n32717 = ~n32700 & n32715;
  assign n32718 = n32700 & ~n32716;
  assign n32719 = n32700 & n32715;
  assign n32720 = ~n32715 & ~n32716;
  assign n32721 = ~n32700 & ~n32715;
  assign n32722 = ~n43501 & ~n43502;
  assign n32723 = ~n32716 & ~n32717;
  assign n32724 = ~n32426 & n32443;
  assign n32725 = ~n32426 & ~n32444;
  assign n32726 = ~n32427 & ~n32724;
  assign n32727 = n43503 & n43504;
  assign n32728 = ~n43503 & ~n43504;
  assign n32729 = ~n32727 & ~n32728;
  assign n32730 = n523 & n785;
  assign n32731 = pi113  & n37520;
  assign n32732 = pi115  & n787;
  assign n32733 = pi114  & n795;
  assign n32734 = ~n32732 & ~n32733;
  assign n32735 = ~n32731 & ~n32733;
  assign n32736 = ~n32732 & n32735;
  assign n32737 = ~n32731 & n32734;
  assign n32738 = ~n32730 & n43505;
  assign n32739 = pi47  & ~n32738;
  assign n32740 = pi47  & ~n32739;
  assign n32741 = pi47  & n32738;
  assign n32742 = ~n32738 & ~n32739;
  assign n32743 = ~pi47  & ~n32738;
  assign n32744 = ~n43506 & ~n43507;
  assign n32745 = n32729 & ~n32744;
  assign n32746 = ~n32729 & n32744;
  assign n32747 = ~n32745 & ~n32746;
  assign n32748 = n32583 & ~n32747;
  assign n32749 = ~n32583 & ~n32746;
  assign n32750 = ~n32745 & n32749;
  assign n32751 = ~n32583 & ~n32745;
  assign n32752 = ~n32746 & n32751;
  assign n32753 = ~n32583 & n32747;
  assign n32754 = ~n32583 & ~n43508;
  assign n32755 = ~n32583 & ~n32747;
  assign n32756 = n32583 & ~n32745;
  assign n32757 = ~n32745 & ~n43508;
  assign n32758 = ~n32746 & ~n32756;
  assign n32759 = ~n32746 & n43510;
  assign n32760 = n32583 & n32747;
  assign n32761 = ~n43509 & ~n43511;
  assign n32762 = ~n32748 & ~n43508;
  assign n32763 = n32582 & n43512;
  assign n32764 = ~n32582 & ~n43512;
  assign n32765 = ~n32763 & ~n32764;
  assign n32766 = ~n32567 & n32765;
  assign n32767 = n32567 & ~n32765;
  assign n32768 = ~n32766 & ~n32767;
  assign n32769 = n733 & n15091;
  assign n32770 = pi119  & n37510;
  assign n32771 = pi121  & n746;
  assign n32772 = pi120  & n748;
  assign n32773 = ~n32771 & ~n32772;
  assign n32774 = ~n32770 & ~n32772;
  assign n32775 = ~n32771 & n32774;
  assign n32776 = ~n32770 & n32773;
  assign n32777 = ~n32769 & n43513;
  assign n32778 = pi41  & ~n32777;
  assign n32779 = pi41  & ~n32778;
  assign n32780 = pi41  & n32777;
  assign n32781 = ~n32777 & ~n32778;
  assign n32782 = ~pi41  & ~n32777;
  assign n32783 = ~n43514 & ~n43515;
  assign n32784 = n32768 & ~n32783;
  assign n32785 = ~n32768 & n32783;
  assign n32786 = n32768 & ~n32784;
  assign n32787 = n32768 & n32783;
  assign n32788 = ~n32783 & ~n32784;
  assign n32789 = ~n32768 & ~n32783;
  assign n32790 = ~n43516 & ~n43517;
  assign n32791 = ~n32784 & ~n32785;
  assign n32792 = n32566 & n43518;
  assign n32793 = ~n32566 & ~n43518;
  assign n32794 = ~n32792 & ~n32793;
  assign n32795 = n691 & n15111;
  assign n32796 = pi122  & n37503;
  assign n32797 = pi124  & n704;
  assign n32798 = pi123  & n706;
  assign n32799 = ~n32797 & ~n32798;
  assign n32800 = ~n32796 & ~n32798;
  assign n32801 = ~n32797 & n32800;
  assign n32802 = ~n32796 & n32799;
  assign n32803 = ~n32795 & n43519;
  assign n32804 = pi38  & ~n32803;
  assign n32805 = pi38  & ~n32804;
  assign n32806 = pi38  & n32803;
  assign n32807 = ~n32803 & ~n32804;
  assign n32808 = ~pi38  & ~n32803;
  assign n32809 = ~n43520 & ~n43521;
  assign n32810 = n32794 & ~n32809;
  assign n32811 = ~n32794 & n32809;
  assign n32812 = n32794 & ~n32810;
  assign n32813 = n32794 & n32809;
  assign n32814 = ~n32809 & ~n32810;
  assign n32815 = ~n32794 & ~n32809;
  assign n32816 = ~n43522 & ~n43523;
  assign n32817 = ~n32810 & ~n32811;
  assign n32818 = ~n32497 & n32514;
  assign n32819 = ~n32497 & ~n32515;
  assign n32820 = ~n32498 & ~n32818;
  assign n32821 = n43524 & n43525;
  assign n32822 = ~n43524 & ~n43525;
  assign n32823 = ~n32821 & ~n32822;
  assign n32824 = n2104 & n40885;
  assign n32825 = pi125  & n37758;
  assign n32826 = pi127  & n2117;
  assign n32827 = pi126  & n2119;
  assign n32828 = ~n32826 & ~n32827;
  assign n32829 = ~n32825 & ~n32827;
  assign n32830 = ~n32826 & n32829;
  assign n32831 = ~n32825 & n32828;
  assign n32832 = ~n32824 & n43526;
  assign n32833 = pi35  & ~n32832;
  assign n32834 = pi35  & ~n32833;
  assign n32835 = pi35  & n32832;
  assign n32836 = ~n32832 & ~n32833;
  assign n32837 = ~pi35  & ~n32832;
  assign n32838 = ~n43527 & ~n43528;
  assign n32839 = ~n32525 & n32541;
  assign n32840 = ~n32525 & ~n32543;
  assign n32841 = ~n32524 & ~n32839;
  assign n32842 = ~n32838 & ~n43529;
  assign n32843 = n32838 & n43529;
  assign n32844 = ~n43529 & ~n32842;
  assign n32845 = n32838 & ~n43529;
  assign n32846 = ~n32838 & ~n32842;
  assign n32847 = ~n32838 & n43529;
  assign n32848 = ~n43530 & ~n43531;
  assign n32849 = ~n32842 & ~n32843;
  assign n32850 = ~n32823 & n43532;
  assign n32851 = n32823 & ~n43532;
  assign n32852 = ~n32850 & ~n32851;
  assign n32853 = ~n32282 & n43469;
  assign n32854 = ~n32282 & ~n32548;
  assign n32855 = ~n32283 & ~n32853;
  assign n32856 = n32852 & ~n43533;
  assign n32857 = ~n32852 & n43533;
  assign n32858 = ~n32856 & ~n32857;
  assign n32859 = ~n32565 & n32858;
  assign n32860 = n32565 & ~n32858;
  assign po96  = ~n32859 & ~n32860;
  assign n32862 = ~n32856 & ~n32859;
  assign n32863 = ~n32842 & ~n32851;
  assign n32864 = ~n32810 & ~n32822;
  assign n32865 = n2104 & n40891;
  assign n32866 = pi126  & n37758;
  assign n32867 = pi127  & n2119;
  assign n32868 = ~n32866 & ~n32867;
  assign n32869 = ~n2104 & n32868;
  assign n32870 = ~n40891 & n32868;
  assign n32871 = ~n32869 & ~n32870;
  assign n32872 = ~n32865 & n32868;
  assign n32873 = pi35  & ~n43534;
  assign n32874 = ~pi35  & n43534;
  assign n32875 = ~n32873 & ~n32874;
  assign n32876 = ~n32864 & ~n32875;
  assign n32877 = n32864 & n32875;
  assign n32878 = ~n32876 & ~n32877;
  assign n32879 = ~n32784 & ~n32793;
  assign n32880 = ~n32764 & ~n32766;
  assign n32881 = n940 & n13027;
  assign n32882 = pi117  & n37541;
  assign n32883 = pi119  & n953;
  assign n32884 = pi118  & n955;
  assign n32885 = ~n32883 & ~n32884;
  assign n32886 = ~n32882 & ~n32884;
  assign n32887 = ~n32883 & n32886;
  assign n32888 = ~n32882 & n32885;
  assign n32889 = ~n32881 & n43535;
  assign n32890 = pi44  & ~n32889;
  assign n32891 = pi44  & ~n32890;
  assign n32892 = pi44  & n32889;
  assign n32893 = ~n32889 & ~n32890;
  assign n32894 = ~pi44  & ~n32889;
  assign n32895 = ~n43536 & ~n43537;
  assign n32896 = ~n32716 & ~n32728;
  assign n32897 = ~n32690 & ~n32699;
  assign n32898 = ~n32664 & ~n32673;
  assign n32899 = ~n32643 & ~n32646;
  assign n32900 = n7882 & n8136;
  assign n32901 = pi102  & n39128;
  assign n32902 = pi104  & n7884;
  assign n32903 = pi103  & n7892;
  assign n32904 = ~n32902 & ~n32903;
  assign n32905 = ~n32901 & ~n32903;
  assign n32906 = ~n32902 & n32905;
  assign n32907 = ~n32901 & n32904;
  assign n32908 = ~n32900 & n43538;
  assign n32909 = pi59  & ~n32908;
  assign n32910 = pi59  & ~n32909;
  assign n32911 = pi59  & n32908;
  assign n32912 = ~n32908 & ~n32909;
  assign n32913 = ~pi59  & ~n32908;
  assign n32914 = ~n43539 & ~n43540;
  assign n32915 = ~n32631 & ~n32637;
  assign n32916 = ~n32620 & ~n43482;
  assign n32917 = ~n32620 & ~n32624;
  assign n32918 = pi98  & ~n40814;
  assign n32919 = pi97  & n18285;
  assign n32920 = ~n32918 & ~n32919;
  assign n32921 = n43541 & ~n32920;
  assign n32922 = ~n43541 & n32920;
  assign n32923 = ~n32921 & ~n32922;
  assign n32924 = n6839 & n12674;
  assign n32925 = pi99  & n40107;
  assign n32926 = pi101  & n12676;
  assign n32927 = pi100  & n12684;
  assign n32928 = ~n32926 & ~n32927;
  assign n32929 = ~n32925 & ~n32927;
  assign n32930 = ~n32926 & n32929;
  assign n32931 = ~n32925 & n32928;
  assign n32932 = ~n32924 & n43542;
  assign n32933 = pi62  & ~n32932;
  assign n32934 = pi62  & ~n32933;
  assign n32935 = pi62  & n32932;
  assign n32936 = ~n32932 & ~n32933;
  assign n32937 = ~pi62  & ~n32932;
  assign n32938 = ~n43543 & ~n43544;
  assign n32939 = ~n32923 & n32938;
  assign n32940 = n32923 & ~n32938;
  assign n32941 = ~n32939 & ~n32940;
  assign n32942 = ~n32915 & n32941;
  assign n32943 = n32915 & ~n32941;
  assign n32944 = ~n32915 & ~n32942;
  assign n32945 = n32941 & ~n32942;
  assign n32946 = ~n32944 & ~n32945;
  assign n32947 = ~n32942 & ~n32943;
  assign n32948 = ~n32914 & ~n43545;
  assign n32949 = n32914 & ~n32945;
  assign n32950 = ~n32944 & n32949;
  assign n32951 = n32914 & n43545;
  assign n32952 = ~n32948 & ~n43546;
  assign n32953 = ~n32899 & n32952;
  assign n32954 = n32899 & ~n32952;
  assign n32955 = ~n32953 & ~n32954;
  assign n32956 = n4312 & n8177;
  assign n32957 = pi105  & n38376;
  assign n32958 = pi107  & n4314;
  assign n32959 = pi106  & n4322;
  assign n32960 = ~n32958 & ~n32959;
  assign n32961 = ~n32957 & ~n32959;
  assign n32962 = ~n32958 & n32961;
  assign n32963 = ~n32957 & n32960;
  assign n32964 = ~n32956 & n43547;
  assign n32965 = pi56  & ~n32964;
  assign n32966 = pi56  & ~n32965;
  assign n32967 = pi56  & n32964;
  assign n32968 = ~n32964 & ~n32965;
  assign n32969 = ~pi56  & ~n32964;
  assign n32970 = ~n43548 & ~n43549;
  assign n32971 = n32955 & ~n32970;
  assign n32972 = ~n32955 & n32970;
  assign n32973 = n32955 & ~n32971;
  assign n32974 = ~n32970 & ~n32971;
  assign n32975 = ~n32973 & ~n32974;
  assign n32976 = ~n32971 & ~n32972;
  assign n32977 = n32898 & n43550;
  assign n32978 = ~n32898 & ~n43550;
  assign n32979 = ~n32977 & ~n32978;
  assign n32980 = n1971 & n9678;
  assign n32981 = pi108  & n37864;
  assign n32982 = pi110  & n1973;
  assign n32983 = pi109  & n1981;
  assign n32984 = ~n32982 & ~n32983;
  assign n32985 = ~n32981 & ~n32983;
  assign n32986 = ~n32982 & n32985;
  assign n32987 = ~n32981 & n32984;
  assign n32988 = ~n32980 & n43551;
  assign n32989 = pi53  & ~n32988;
  assign n32990 = pi53  & ~n32989;
  assign n32991 = pi53  & n32988;
  assign n32992 = ~n32988 & ~n32989;
  assign n32993 = ~pi53  & ~n32988;
  assign n32994 = ~n43552 & ~n43553;
  assign n32995 = ~n32979 & n32994;
  assign n32996 = n32979 & ~n32994;
  assign n32997 = n32979 & ~n32996;
  assign n32998 = ~n32994 & ~n32996;
  assign n32999 = ~n32997 & ~n32998;
  assign n33000 = ~n32995 & ~n32996;
  assign n33001 = n32897 & n43554;
  assign n33002 = ~n32897 & ~n43554;
  assign n33003 = ~n33001 & ~n33002;
  assign n33004 = n894 & n11276;
  assign n33005 = pi111  & n37580;
  assign n33006 = pi113  & n896;
  assign n33007 = pi112  & n904;
  assign n33008 = ~n33006 & ~n33007;
  assign n33009 = ~n33005 & ~n33007;
  assign n33010 = ~n33006 & n33009;
  assign n33011 = ~n33005 & n33008;
  assign n33012 = ~n33004 & n43555;
  assign n33013 = pi50  & ~n33012;
  assign n33014 = pi50  & ~n33013;
  assign n33015 = pi50  & n33012;
  assign n33016 = ~n33012 & ~n33013;
  assign n33017 = ~pi50  & ~n33012;
  assign n33018 = ~n43556 & ~n43557;
  assign n33019 = n33003 & ~n33018;
  assign n33020 = ~n33003 & n33018;
  assign n33021 = n33003 & ~n33019;
  assign n33022 = ~n33018 & ~n33019;
  assign n33023 = ~n33021 & ~n33022;
  assign n33024 = ~n33019 & ~n33020;
  assign n33025 = n32896 & n43558;
  assign n33026 = ~n32896 & ~n43558;
  assign n33027 = ~n33025 & ~n33026;
  assign n33028 = n785 & n12530;
  assign n33029 = pi114  & n37520;
  assign n33030 = pi116  & n787;
  assign n33031 = pi115  & n795;
  assign n33032 = ~n33030 & ~n33031;
  assign n33033 = ~n33029 & ~n33031;
  assign n33034 = ~n33030 & n33033;
  assign n33035 = ~n33029 & n33032;
  assign n33036 = ~n33028 & n43559;
  assign n33037 = pi47  & ~n33036;
  assign n33038 = pi47  & ~n33037;
  assign n33039 = pi47  & n33036;
  assign n33040 = ~n33036 & ~n33037;
  assign n33041 = ~pi47  & ~n33036;
  assign n33042 = ~n43560 & ~n43561;
  assign n33043 = ~n33027 & n33042;
  assign n33044 = n33027 & ~n33042;
  assign n33045 = n33027 & ~n33044;
  assign n33046 = ~n33042 & ~n33044;
  assign n33047 = ~n33045 & ~n33046;
  assign n33048 = ~n33043 & ~n33044;
  assign n33049 = ~n43510 & ~n43562;
  assign n33050 = n43510 & n43562;
  assign n33051 = ~n43510 & n43562;
  assign n33052 = n43510 & ~n43562;
  assign n33053 = ~n33051 & ~n33052;
  assign n33054 = ~n33049 & ~n33050;
  assign n33055 = ~n32895 & ~n43563;
  assign n33056 = n32895 & n43563;
  assign n33057 = ~n33055 & ~n33056;
  assign n33058 = ~n32880 & n33057;
  assign n33059 = n32880 & ~n33057;
  assign n33060 = ~n33058 & ~n33059;
  assign n33061 = n733 & n15049;
  assign n33062 = pi120  & n37510;
  assign n33063 = pi122  & n746;
  assign n33064 = pi121  & n748;
  assign n33065 = ~n33063 & ~n33064;
  assign n33066 = ~n33062 & ~n33064;
  assign n33067 = ~n33063 & n33066;
  assign n33068 = ~n33062 & n33065;
  assign n33069 = ~n33061 & n43564;
  assign n33070 = pi41  & ~n33069;
  assign n33071 = pi41  & ~n33070;
  assign n33072 = pi41  & n33069;
  assign n33073 = ~n33069 & ~n33070;
  assign n33074 = ~pi41  & ~n33069;
  assign n33075 = ~n43565 & ~n43566;
  assign n33076 = n33060 & ~n33075;
  assign n33077 = ~n33060 & n33075;
  assign n33078 = n33060 & ~n33076;
  assign n33079 = ~n33075 & ~n33076;
  assign n33080 = ~n33078 & ~n33079;
  assign n33081 = ~n33076 & ~n33077;
  assign n33082 = n32879 & n43567;
  assign n33083 = ~n32879 & ~n43567;
  assign n33084 = ~n33082 & ~n33083;
  assign n33085 = n691 & n15068;
  assign n33086 = pi123  & n37503;
  assign n33087 = pi125  & n704;
  assign n33088 = pi124  & n706;
  assign n33089 = ~n33087 & ~n33088;
  assign n33090 = ~n33086 & ~n33088;
  assign n33091 = ~n33087 & n33090;
  assign n33092 = ~n33086 & n33089;
  assign n33093 = ~n33085 & n43568;
  assign n33094 = pi38  & ~n33093;
  assign n33095 = pi38  & ~n33094;
  assign n33096 = pi38  & n33093;
  assign n33097 = ~n33093 & ~n33094;
  assign n33098 = ~pi38  & ~n33093;
  assign n33099 = ~n43569 & ~n43570;
  assign n33100 = n33084 & ~n33099;
  assign n33101 = ~n33084 & n33099;
  assign n33102 = ~n33100 & ~n33101;
  assign n33103 = n32878 & ~n33101;
  assign n33104 = ~n33100 & n33103;
  assign n33105 = n32878 & n33102;
  assign n33106 = ~n32878 & ~n33102;
  assign n33107 = n32878 & ~n43571;
  assign n33108 = ~n33101 & ~n43571;
  assign n33109 = ~n33100 & n33108;
  assign n33110 = n33102 & ~n43571;
  assign n33111 = ~n33107 & ~n43572;
  assign n33112 = ~n43571 & ~n33106;
  assign n33113 = ~n32863 & ~n43573;
  assign n33114 = n32863 & n43573;
  assign n33115 = ~n43573 & ~n33113;
  assign n33116 = ~n32863 & ~n33113;
  assign n33117 = ~n33115 & ~n33116;
  assign n33118 = ~n33113 & ~n33114;
  assign n33119 = ~n32862 & ~n43574;
  assign n33120 = n32862 & n43574;
  assign po97  = ~n33119 & ~n33120;
  assign n33122 = ~n33113 & ~n33119;
  assign n33123 = ~n32876 & ~n43571;
  assign n33124 = ~n33083 & ~n33100;
  assign n33125 = n2104 & ~n18675;
  assign n33126 = ~n37758 & ~n33125;
  assign n33127 = pi127  & n37758;
  assign n33128 = n2104 & n18680;
  assign n33129 = ~n33127 & ~n33128;
  assign n33130 = pi127  & ~n33126;
  assign n33131 = pi35  & ~n43575;
  assign n33132 = pi35  & ~n33131;
  assign n33133 = pi35  & n43575;
  assign n33134 = ~n43575 & ~n33131;
  assign n33135 = ~pi35  & ~n43575;
  assign n33136 = ~n43576 & ~n43577;
  assign n33137 = ~n33124 & ~n33136;
  assign n33138 = n33124 & n33136;
  assign n33139 = ~n33124 & ~n33137;
  assign n33140 = ~n33136 & ~n33137;
  assign n33141 = ~n33139 & ~n33140;
  assign n33142 = ~n33137 & ~n33138;
  assign n33143 = ~n33049 & ~n33055;
  assign n33144 = n940 & n14913;
  assign n33145 = pi118  & n37541;
  assign n33146 = pi120  & n953;
  assign n33147 = pi119  & n955;
  assign n33148 = ~n33146 & ~n33147;
  assign n33149 = ~n33145 & ~n33147;
  assign n33150 = ~n33146 & n33149;
  assign n33151 = ~n33145 & n33148;
  assign n33152 = ~n33144 & n43579;
  assign n33153 = pi44  & ~n33152;
  assign n33154 = pi44  & ~n33153;
  assign n33155 = pi44  & n33152;
  assign n33156 = ~n33152 & ~n33153;
  assign n33157 = ~pi44  & ~n33152;
  assign n33158 = ~n43580 & ~n43581;
  assign n33159 = n785 & n13079;
  assign n33160 = pi115  & n37520;
  assign n33161 = pi117  & n787;
  assign n33162 = pi116  & n795;
  assign n33163 = ~n33161 & ~n33162;
  assign n33164 = ~n33160 & ~n33162;
  assign n33165 = ~n33161 & n33164;
  assign n33166 = ~n33160 & n33163;
  assign n33167 = ~n33159 & n43582;
  assign n33168 = pi47  & ~n33167;
  assign n33169 = pi47  & ~n33168;
  assign n33170 = pi47  & n33167;
  assign n33171 = ~n33167 & ~n33168;
  assign n33172 = ~pi47  & ~n33167;
  assign n33173 = ~n43583 & ~n43584;
  assign n33174 = n4312 & n9277;
  assign n33175 = pi106  & n38376;
  assign n33176 = pi108  & n4314;
  assign n33177 = pi107  & n4322;
  assign n33178 = ~n33176 & ~n33177;
  assign n33179 = ~n33175 & ~n33177;
  assign n33180 = ~n33176 & n33179;
  assign n33181 = ~n33175 & n33178;
  assign n33182 = ~n33174 & n43585;
  assign n33183 = pi56  & ~n33182;
  assign n33184 = pi56  & ~n33183;
  assign n33185 = pi56  & n33182;
  assign n33186 = ~n33182 & ~n33183;
  assign n33187 = ~pi56  & ~n33182;
  assign n33188 = ~n43586 & ~n43587;
  assign n33189 = ~n32942 & ~n32948;
  assign n33190 = n7882 & n8229;
  assign n33191 = pi103  & n39128;
  assign n33192 = pi105  & n7884;
  assign n33193 = pi104  & n7892;
  assign n33194 = ~n33192 & ~n33193;
  assign n33195 = ~n33191 & ~n33193;
  assign n33196 = ~n33192 & n33195;
  assign n33197 = ~n33191 & n33194;
  assign n33198 = ~n33190 & n43588;
  assign n33199 = pi59  & ~n33198;
  assign n33200 = pi59  & ~n33199;
  assign n33201 = pi59  & n33198;
  assign n33202 = ~n33198 & ~n33199;
  assign n33203 = ~pi59  & ~n33198;
  assign n33204 = ~n43589 & ~n43590;
  assign n33205 = n6819 & n12674;
  assign n33206 = pi100  & n40107;
  assign n33207 = pi102  & n12676;
  assign n33208 = pi101  & n12684;
  assign n33209 = ~n33207 & ~n33208;
  assign n33210 = ~n33206 & ~n33208;
  assign n33211 = ~n33207 & n33210;
  assign n33212 = ~n33206 & n33209;
  assign n33213 = ~n33205 & n43591;
  assign n33214 = pi62  & ~n33213;
  assign n33215 = pi62  & ~n33214;
  assign n33216 = pi62  & n33213;
  assign n33217 = ~n33213 & ~n33214;
  assign n33218 = ~pi62  & ~n33213;
  assign n33219 = ~n43592 & ~n43593;
  assign n33220 = ~n32922 & ~n32940;
  assign n33221 = pi99  & ~n40814;
  assign n33222 = pi98  & n18285;
  assign n33223 = ~n33221 & ~n33222;
  assign n33224 = ~n32920 & n33223;
  assign n33225 = n32920 & ~n33223;
  assign n33226 = ~n33224 & ~n33225;
  assign n33227 = ~n33220 & ~n33225;
  assign n33228 = ~n33224 & n33227;
  assign n33229 = ~n33220 & n33226;
  assign n33230 = n33220 & ~n33226;
  assign n33231 = ~n33220 & ~n43594;
  assign n33232 = ~n33224 & ~n43594;
  assign n33233 = ~n33225 & n33232;
  assign n33234 = ~n33231 & ~n33233;
  assign n33235 = ~n43594 & ~n33230;
  assign n33236 = ~n33219 & ~n43595;
  assign n33237 = n33219 & n43595;
  assign n33238 = ~n43595 & ~n33236;
  assign n33239 = n33219 & ~n43595;
  assign n33240 = ~n33219 & ~n33236;
  assign n33241 = ~n33219 & n43595;
  assign n33242 = ~n43596 & ~n43597;
  assign n33243 = ~n33236 & ~n33237;
  assign n33244 = ~n33204 & ~n43598;
  assign n33245 = n33204 & n43598;
  assign n33246 = n33204 & ~n43598;
  assign n33247 = ~n33204 & n43598;
  assign n33248 = ~n33246 & ~n33247;
  assign n33249 = ~n33244 & ~n33245;
  assign n33250 = ~n33189 & ~n43599;
  assign n33251 = n33189 & n43599;
  assign n33252 = ~n33250 & ~n33251;
  assign n33253 = ~n33188 & n33252;
  assign n33254 = n33188 & ~n33252;
  assign n33255 = ~n33253 & ~n33254;
  assign n33256 = ~n32953 & n32970;
  assign n33257 = ~n32953 & ~n32971;
  assign n33258 = ~n32954 & ~n33256;
  assign n33259 = n33255 & ~n43600;
  assign n33260 = ~n33255 & n43600;
  assign n33261 = ~n33259 & ~n33260;
  assign n33262 = n565 & n1971;
  assign n33263 = pi109  & n37864;
  assign n33264 = pi111  & n1973;
  assign n33265 = pi110  & n1981;
  assign n33266 = ~n33264 & ~n33265;
  assign n33267 = ~n33263 & ~n33265;
  assign n33268 = ~n33264 & n33267;
  assign n33269 = ~n33263 & n33266;
  assign n33270 = ~n33262 & n43601;
  assign n33271 = pi53  & ~n33270;
  assign n33272 = pi53  & ~n33271;
  assign n33273 = pi53  & n33270;
  assign n33274 = ~n33270 & ~n33271;
  assign n33275 = ~pi53  & ~n33270;
  assign n33276 = ~n43602 & ~n43603;
  assign n33277 = n33261 & ~n33276;
  assign n33278 = ~n33261 & n33276;
  assign n33279 = n33261 & ~n33277;
  assign n33280 = ~n33276 & ~n33277;
  assign n33281 = ~n33279 & ~n33280;
  assign n33282 = ~n33277 & ~n33278;
  assign n33283 = ~n32978 & n32994;
  assign n33284 = ~n32978 & ~n32996;
  assign n33285 = ~n32977 & ~n33283;
  assign n33286 = n43604 & n43605;
  assign n33287 = ~n43604 & ~n43605;
  assign n33288 = ~n33286 & ~n33287;
  assign n33289 = n894 & n11258;
  assign n33290 = pi112  & n37580;
  assign n33291 = pi114  & n896;
  assign n33292 = pi113  & n904;
  assign n33293 = ~n33291 & ~n33292;
  assign n33294 = ~n33290 & ~n33292;
  assign n33295 = ~n33291 & n33294;
  assign n33296 = ~n33290 & n33293;
  assign n33297 = ~n33289 & n43606;
  assign n33298 = pi50  & ~n33297;
  assign n33299 = pi50  & ~n33298;
  assign n33300 = pi50  & n33297;
  assign n33301 = ~n33297 & ~n33298;
  assign n33302 = ~pi50  & ~n33297;
  assign n33303 = ~n43607 & ~n43608;
  assign n33304 = ~n33288 & n33303;
  assign n33305 = n33288 & ~n33303;
  assign n33306 = ~n33304 & ~n33305;
  assign n33307 = ~n33002 & n33018;
  assign n33308 = ~n33002 & ~n33019;
  assign n33309 = ~n33001 & ~n33307;
  assign n33310 = n33306 & ~n43609;
  assign n33311 = ~n33306 & n43609;
  assign n33312 = ~n43609 & ~n33310;
  assign n33313 = n33306 & ~n33310;
  assign n33314 = ~n33312 & ~n33313;
  assign n33315 = ~n33310 & ~n33311;
  assign n33316 = ~n33173 & ~n43610;
  assign n33317 = n33173 & ~n33313;
  assign n33318 = ~n33312 & n33317;
  assign n33319 = n33173 & n43610;
  assign n33320 = ~n33316 & ~n43611;
  assign n33321 = ~n33026 & n33042;
  assign n33322 = ~n33026 & ~n33044;
  assign n33323 = ~n33025 & ~n33321;
  assign n33324 = n33320 & ~n43612;
  assign n33325 = ~n33320 & n43612;
  assign n33326 = ~n33324 & ~n33325;
  assign n33327 = ~n33158 & n33326;
  assign n33328 = n33158 & ~n33326;
  assign n33329 = ~n33327 & ~n33328;
  assign n33330 = ~n33143 & n33329;
  assign n33331 = n33143 & ~n33329;
  assign n33332 = ~n33330 & ~n33331;
  assign n33333 = n733 & n14961;
  assign n33334 = pi121  & n37510;
  assign n33335 = pi123  & n746;
  assign n33336 = pi122  & n748;
  assign n33337 = ~n33335 & ~n33336;
  assign n33338 = ~n33334 & ~n33336;
  assign n33339 = ~n33335 & n33338;
  assign n33340 = ~n33334 & n33337;
  assign n33341 = ~n33333 & n43613;
  assign n33342 = pi41  & ~n33341;
  assign n33343 = pi41  & ~n33342;
  assign n33344 = pi41  & n33341;
  assign n33345 = ~n33341 & ~n33342;
  assign n33346 = ~pi41  & ~n33341;
  assign n33347 = ~n43614 & ~n43615;
  assign n33348 = n33332 & ~n33347;
  assign n33349 = ~n33332 & n33347;
  assign n33350 = n33332 & ~n33348;
  assign n33351 = ~n33347 & ~n33348;
  assign n33352 = ~n33350 & ~n33351;
  assign n33353 = ~n33348 & ~n33349;
  assign n33354 = ~n33058 & n33075;
  assign n33355 = ~n33058 & ~n33076;
  assign n33356 = ~n33059 & ~n33354;
  assign n33357 = n43616 & n43617;
  assign n33358 = ~n43616 & ~n43617;
  assign n33359 = ~n33357 & ~n33358;
  assign n33360 = n691 & n15021;
  assign n33361 = pi124  & n37503;
  assign n33362 = pi126  & n704;
  assign n33363 = pi125  & n706;
  assign n33364 = ~n33362 & ~n33363;
  assign n33365 = ~n33361 & ~n33363;
  assign n33366 = ~n33362 & n33365;
  assign n33367 = ~n33361 & n33364;
  assign n33368 = ~n33360 & n43618;
  assign n33369 = pi38  & ~n33368;
  assign n33370 = pi38  & ~n33369;
  assign n33371 = pi38  & n33368;
  assign n33372 = ~n33368 & ~n33369;
  assign n33373 = ~pi38  & ~n33368;
  assign n33374 = ~n43619 & ~n43620;
  assign n33375 = ~n33359 & n33374;
  assign n33376 = n33359 & ~n33374;
  assign n33377 = n33359 & ~n33376;
  assign n33378 = ~n33374 & ~n33376;
  assign n33379 = ~n33377 & ~n33378;
  assign n33380 = ~n33375 & ~n33376;
  assign n33381 = ~n43578 & ~n43621;
  assign n33382 = n43578 & n43621;
  assign n33383 = ~n43578 & n43621;
  assign n33384 = n43578 & ~n43621;
  assign n33385 = ~n33383 & ~n33384;
  assign n33386 = ~n33381 & ~n33382;
  assign n33387 = ~n33123 & ~n43622;
  assign n33388 = n33123 & n43622;
  assign n33389 = ~n33387 & ~n33388;
  assign n33390 = ~n33122 & n33389;
  assign n33391 = n33122 & ~n33389;
  assign po98  = ~n33390 & ~n33391;
  assign n33393 = ~n33387 & ~n33390;
  assign n33394 = ~n33324 & ~n33327;
  assign n33395 = ~n33310 & ~n33316;
  assign n33396 = n785 & n13057;
  assign n33397 = pi116  & n37520;
  assign n33398 = pi118  & n787;
  assign n33399 = pi117  & n795;
  assign n33400 = ~n33398 & ~n33399;
  assign n33401 = ~n33397 & ~n33399;
  assign n33402 = ~n33398 & n33401;
  assign n33403 = ~n33397 & n33400;
  assign n33404 = ~n33396 & n43623;
  assign n33405 = pi47  & ~n33404;
  assign n33406 = pi47  & ~n33405;
  assign n33407 = pi47  & n33404;
  assign n33408 = ~n33404 & ~n33405;
  assign n33409 = ~pi47  & ~n33404;
  assign n33410 = ~n43624 & ~n43625;
  assign n33411 = ~n33287 & ~n33305;
  assign n33412 = ~n33250 & ~n33253;
  assign n33413 = n4312 & n9701;
  assign n33414 = pi107  & n38376;
  assign n33415 = pi109  & n4314;
  assign n33416 = pi108  & n4322;
  assign n33417 = ~n33415 & ~n33416;
  assign n33418 = ~n33414 & ~n33416;
  assign n33419 = ~n33415 & n33418;
  assign n33420 = ~n33414 & n33417;
  assign n33421 = ~n33413 & n43626;
  assign n33422 = pi56  & ~n33421;
  assign n33423 = pi56  & ~n33422;
  assign n33424 = pi56  & n33421;
  assign n33425 = ~n33421 & ~n33422;
  assign n33426 = ~pi56  & ~n33421;
  assign n33427 = ~n43627 & ~n43628;
  assign n33428 = ~n33236 & ~n33244;
  assign n33429 = ~pi35  & ~n33223;
  assign n33430 = pi35  & n33223;
  assign n33431 = pi35  & ~n33223;
  assign n33432 = ~pi35  & n33223;
  assign n33433 = ~n33431 & ~n33432;
  assign n33434 = ~n33429 & ~n33430;
  assign n33435 = pi100  & ~n40814;
  assign n33436 = pi99  & n18285;
  assign n33437 = ~n33435 & ~n33436;
  assign n33438 = ~n43629 & ~n33437;
  assign n33439 = n43629 & n33437;
  assign n33440 = ~n33438 & ~n33439;
  assign n33441 = ~n33232 & n33440;
  assign n33442 = n33232 & ~n33440;
  assign n33443 = ~n33441 & ~n33442;
  assign n33444 = n6787 & n12674;
  assign n33445 = pi101  & n40107;
  assign n33446 = pi103  & n12676;
  assign n33447 = pi102  & n12684;
  assign n33448 = ~n33446 & ~n33447;
  assign n33449 = ~n33445 & ~n33447;
  assign n33450 = ~n33446 & n33449;
  assign n33451 = ~n33445 & n33448;
  assign n33452 = ~n33444 & n43630;
  assign n33453 = pi62  & ~n33452;
  assign n33454 = pi62  & ~n33453;
  assign n33455 = pi62  & n33452;
  assign n33456 = ~n33452 & ~n33453;
  assign n33457 = ~pi62  & ~n33452;
  assign n33458 = ~n43631 & ~n43632;
  assign n33459 = ~n33443 & n33458;
  assign n33460 = n33443 & ~n33458;
  assign n33461 = ~n33459 & ~n33460;
  assign n33462 = n7882 & n8209;
  assign n33463 = pi104  & n39128;
  assign n33464 = pi106  & n7884;
  assign n33465 = pi105  & n7892;
  assign n33466 = ~n33464 & ~n33465;
  assign n33467 = ~n33463 & ~n33465;
  assign n33468 = ~n33464 & n33467;
  assign n33469 = ~n33463 & n33466;
  assign n33470 = ~n33462 & n43633;
  assign n33471 = pi59  & ~n33470;
  assign n33472 = pi59  & ~n33471;
  assign n33473 = pi59  & n33470;
  assign n33474 = ~n33470 & ~n33471;
  assign n33475 = ~pi59  & ~n33470;
  assign n33476 = ~n43634 & ~n43635;
  assign n33477 = n33461 & ~n33476;
  assign n33478 = ~n33461 & n33476;
  assign n33479 = n33461 & ~n33477;
  assign n33480 = n33461 & n33476;
  assign n33481 = ~n33476 & ~n33477;
  assign n33482 = ~n33461 & ~n33476;
  assign n33483 = ~n43636 & ~n43637;
  assign n33484 = ~n33477 & ~n33478;
  assign n33485 = ~n33428 & ~n43638;
  assign n33486 = n33428 & n43638;
  assign n33487 = ~n43638 & ~n33485;
  assign n33488 = ~n33428 & ~n33485;
  assign n33489 = ~n33487 & ~n33488;
  assign n33490 = ~n33485 & ~n33486;
  assign n33491 = ~n33427 & ~n43639;
  assign n33492 = n33427 & n43639;
  assign n33493 = ~n43639 & ~n33491;
  assign n33494 = n33427 & ~n43639;
  assign n33495 = ~n33427 & ~n33491;
  assign n33496 = ~n33427 & n43639;
  assign n33497 = ~n43640 & ~n43641;
  assign n33498 = ~n33491 & ~n33492;
  assign n33499 = n33412 & n43642;
  assign n33500 = ~n33412 & ~n43642;
  assign n33501 = ~n33499 & ~n33500;
  assign n33502 = n1971 & n10844;
  assign n33503 = pi110  & n37864;
  assign n33504 = pi112  & n1973;
  assign n33505 = pi111  & n1981;
  assign n33506 = ~n33504 & ~n33505;
  assign n33507 = ~n33503 & ~n33505;
  assign n33508 = ~n33504 & n33507;
  assign n33509 = ~n33503 & n33506;
  assign n33510 = ~n33502 & n43643;
  assign n33511 = pi53  & ~n33510;
  assign n33512 = pi53  & ~n33511;
  assign n33513 = pi53  & n33510;
  assign n33514 = ~n33510 & ~n33511;
  assign n33515 = ~pi53  & ~n33510;
  assign n33516 = ~n43644 & ~n43645;
  assign n33517 = n33501 & ~n33516;
  assign n33518 = ~n33501 & n33516;
  assign n33519 = n33501 & ~n33517;
  assign n33520 = n33501 & n33516;
  assign n33521 = ~n33516 & ~n33517;
  assign n33522 = ~n33501 & ~n33516;
  assign n33523 = ~n43646 & ~n43647;
  assign n33524 = ~n33517 & ~n33518;
  assign n33525 = ~n33259 & n33276;
  assign n33526 = ~n33259 & ~n33277;
  assign n33527 = ~n33260 & ~n33525;
  assign n33528 = n43648 & n43649;
  assign n33529 = ~n43648 & ~n43649;
  assign n33530 = ~n33528 & ~n33529;
  assign n33531 = n523 & n894;
  assign n33532 = pi113  & n37580;
  assign n33533 = pi115  & n896;
  assign n33534 = pi114  & n904;
  assign n33535 = ~n33533 & ~n33534;
  assign n33536 = ~n33532 & ~n33534;
  assign n33537 = ~n33533 & n33536;
  assign n33538 = ~n33532 & n33535;
  assign n33539 = ~n33531 & n43650;
  assign n33540 = pi50  & ~n33539;
  assign n33541 = pi50  & ~n33540;
  assign n33542 = pi50  & n33539;
  assign n33543 = ~n33539 & ~n33540;
  assign n33544 = ~pi50  & ~n33539;
  assign n33545 = ~n43651 & ~n43652;
  assign n33546 = ~n33530 & n33545;
  assign n33547 = n33530 & ~n33545;
  assign n33548 = ~n33546 & ~n33547;
  assign n33549 = ~n33411 & n33548;
  assign n33550 = n33411 & ~n33548;
  assign n33551 = ~n33549 & ~n33550;
  assign n33552 = ~n33410 & n33551;
  assign n33553 = n33410 & ~n33551;
  assign n33554 = ~n33552 & ~n33553;
  assign n33555 = ~n33395 & n33554;
  assign n33556 = n33395 & ~n33554;
  assign n33557 = ~n33555 & ~n33556;
  assign n33558 = n940 & n15091;
  assign n33559 = pi119  & n37541;
  assign n33560 = pi121  & n953;
  assign n33561 = pi120  & n955;
  assign n33562 = ~n33560 & ~n33561;
  assign n33563 = ~n33559 & ~n33561;
  assign n33564 = ~n33560 & n33563;
  assign n33565 = ~n33559 & n33562;
  assign n33566 = ~n33558 & n43653;
  assign n33567 = pi44  & ~n33566;
  assign n33568 = pi44  & ~n33567;
  assign n33569 = pi44  & n33566;
  assign n33570 = ~n33566 & ~n33567;
  assign n33571 = ~pi44  & ~n33566;
  assign n33572 = ~n43654 & ~n43655;
  assign n33573 = n33557 & ~n33572;
  assign n33574 = ~n33557 & n33572;
  assign n33575 = n33557 & ~n33573;
  assign n33576 = n33557 & n33572;
  assign n33577 = ~n33572 & ~n33573;
  assign n33578 = ~n33557 & ~n33572;
  assign n33579 = ~n43656 & ~n43657;
  assign n33580 = ~n33573 & ~n33574;
  assign n33581 = n33394 & n43658;
  assign n33582 = ~n33394 & ~n43658;
  assign n33583 = ~n33581 & ~n33582;
  assign n33584 = n733 & n15111;
  assign n33585 = pi122  & n37510;
  assign n33586 = pi124  & n746;
  assign n33587 = pi123  & n748;
  assign n33588 = ~n33586 & ~n33587;
  assign n33589 = ~n33585 & ~n33587;
  assign n33590 = ~n33586 & n33589;
  assign n33591 = ~n33585 & n33588;
  assign n33592 = ~n33584 & n43659;
  assign n33593 = pi41  & ~n33592;
  assign n33594 = pi41  & ~n33593;
  assign n33595 = pi41  & n33592;
  assign n33596 = ~n33592 & ~n33593;
  assign n33597 = ~pi41  & ~n33592;
  assign n33598 = ~n43660 & ~n43661;
  assign n33599 = n33583 & ~n33598;
  assign n33600 = ~n33583 & n33598;
  assign n33601 = n33583 & ~n33599;
  assign n33602 = n33583 & n33598;
  assign n33603 = ~n33598 & ~n33599;
  assign n33604 = ~n33583 & ~n33598;
  assign n33605 = ~n43662 & ~n43663;
  assign n33606 = ~n33599 & ~n33600;
  assign n33607 = ~n33330 & n33347;
  assign n33608 = ~n33330 & ~n33348;
  assign n33609 = ~n33331 & ~n33607;
  assign n33610 = n43664 & n43665;
  assign n33611 = ~n43664 & ~n43665;
  assign n33612 = ~n33610 & ~n33611;
  assign n33613 = n691 & n40885;
  assign n33614 = pi125  & n37503;
  assign n33615 = pi127  & n704;
  assign n33616 = pi126  & n706;
  assign n33617 = ~n33615 & ~n33616;
  assign n33618 = ~n33614 & ~n33616;
  assign n33619 = ~n33615 & n33618;
  assign n33620 = ~n33614 & n33617;
  assign n33621 = ~n33613 & n43666;
  assign n33622 = pi38  & ~n33621;
  assign n33623 = pi38  & ~n33622;
  assign n33624 = pi38  & n33621;
  assign n33625 = ~n33621 & ~n33622;
  assign n33626 = ~pi38  & ~n33621;
  assign n33627 = ~n43667 & ~n43668;
  assign n33628 = n33612 & ~n33627;
  assign n33629 = ~n33612 & n33627;
  assign n33630 = n33612 & ~n33628;
  assign n33631 = n33612 & n33627;
  assign n33632 = ~n33627 & ~n33628;
  assign n33633 = ~n33612 & ~n33627;
  assign n33634 = ~n43669 & ~n43670;
  assign n33635 = ~n33628 & ~n33629;
  assign n33636 = ~n33358 & n33374;
  assign n33637 = ~n33358 & ~n33376;
  assign n33638 = ~n33357 & ~n33636;
  assign n33639 = n43671 & n43672;
  assign n33640 = ~n43671 & ~n43672;
  assign n33641 = ~n33639 & ~n33640;
  assign n33642 = ~n33137 & n43621;
  assign n33643 = ~n33137 & ~n33381;
  assign n33644 = ~n33138 & ~n33642;
  assign n33645 = n33641 & ~n43673;
  assign n33646 = ~n33641 & n43673;
  assign n33647 = ~n33645 & ~n33646;
  assign n33648 = ~n33393 & n33647;
  assign n33649 = n33393 & ~n33647;
  assign po99  = ~n33648 & ~n33649;
  assign n33651 = ~n33628 & ~n33640;
  assign n33652 = ~n33599 & ~n33611;
  assign n33653 = n691 & n40891;
  assign n33654 = pi126  & n37503;
  assign n33655 = pi127  & n706;
  assign n33656 = ~n33654 & ~n33655;
  assign n33657 = ~n691 & n33656;
  assign n33658 = ~n40891 & n33656;
  assign n33659 = ~n33657 & ~n33658;
  assign n33660 = ~n33653 & n33656;
  assign n33661 = pi38  & ~n43674;
  assign n33662 = ~pi38  & n43674;
  assign n33663 = ~n33661 & ~n33662;
  assign n33664 = ~n33652 & ~n33663;
  assign n33665 = n33652 & n33663;
  assign n33666 = ~n33664 & ~n33665;
  assign n33667 = ~n33573 & ~n33582;
  assign n33668 = ~n33552 & ~n33555;
  assign n33669 = n785 & n13027;
  assign n33670 = pi117  & n37520;
  assign n33671 = pi119  & n787;
  assign n33672 = pi118  & n795;
  assign n33673 = ~n33671 & ~n33672;
  assign n33674 = ~n33670 & ~n33672;
  assign n33675 = ~n33671 & n33674;
  assign n33676 = ~n33670 & n33673;
  assign n33677 = ~n33669 & n43675;
  assign n33678 = pi47  & ~n33677;
  assign n33679 = pi47  & ~n33678;
  assign n33680 = pi47  & n33677;
  assign n33681 = ~n33677 & ~n33678;
  assign n33682 = ~pi47  & ~n33677;
  assign n33683 = ~n43676 & ~n43677;
  assign n33684 = ~n33547 & ~n33549;
  assign n33685 = ~n33517 & ~n33529;
  assign n33686 = ~n33491 & ~n33500;
  assign n33687 = ~n33477 & ~n33485;
  assign n33688 = ~n33441 & ~n33460;
  assign n33689 = n8136 & n12674;
  assign n33690 = pi102  & n40107;
  assign n33691 = pi104  & n12676;
  assign n33692 = pi103  & n12684;
  assign n33693 = ~n33691 & ~n33692;
  assign n33694 = ~n33690 & ~n33692;
  assign n33695 = ~n33691 & n33694;
  assign n33696 = ~n33690 & n33693;
  assign n33697 = ~n33689 & n43678;
  assign n33698 = pi62  & ~n33697;
  assign n33699 = pi62  & ~n33698;
  assign n33700 = pi62  & n33697;
  assign n33701 = ~n33697 & ~n33698;
  assign n33702 = ~pi62  & ~n33697;
  assign n33703 = ~n43679 & ~n43680;
  assign n33704 = ~n33429 & ~n33438;
  assign n33705 = pi101  & ~n40814;
  assign n33706 = pi100  & n18285;
  assign n33707 = ~n33705 & ~n33706;
  assign n33708 = ~n33704 & n33707;
  assign n33709 = n33704 & ~n33707;
  assign n33710 = n33707 & ~n33708;
  assign n33711 = n33704 & n33707;
  assign n33712 = ~n33704 & ~n33708;
  assign n33713 = ~n33704 & ~n33707;
  assign n33714 = ~n43681 & ~n43682;
  assign n33715 = ~n33708 & ~n33709;
  assign n33716 = ~n33703 & ~n43683;
  assign n33717 = n33703 & n43683;
  assign n33718 = ~n33703 & ~n33716;
  assign n33719 = ~n33703 & n43683;
  assign n33720 = ~n43683 & ~n33716;
  assign n33721 = n33703 & ~n43683;
  assign n33722 = ~n43684 & ~n43685;
  assign n33723 = ~n33716 & ~n33717;
  assign n33724 = n33688 & n43686;
  assign n33725 = ~n33688 & ~n43686;
  assign n33726 = ~n33724 & ~n33725;
  assign n33727 = n7882 & n8177;
  assign n33728 = pi105  & n39128;
  assign n33729 = pi107  & n7884;
  assign n33730 = pi106  & n7892;
  assign n33731 = ~n33729 & ~n33730;
  assign n33732 = ~n33728 & ~n33730;
  assign n33733 = ~n33729 & n33732;
  assign n33734 = ~n33728 & n33731;
  assign n33735 = ~n33727 & n43687;
  assign n33736 = pi59  & ~n33735;
  assign n33737 = pi59  & ~n33736;
  assign n33738 = pi59  & n33735;
  assign n33739 = ~n33735 & ~n33736;
  assign n33740 = ~pi59  & ~n33735;
  assign n33741 = ~n43688 & ~n43689;
  assign n33742 = n33726 & ~n33741;
  assign n33743 = ~n33726 & n33741;
  assign n33744 = n33726 & ~n33742;
  assign n33745 = ~n33741 & ~n33742;
  assign n33746 = ~n33744 & ~n33745;
  assign n33747 = ~n33742 & ~n33743;
  assign n33748 = n33687 & n43690;
  assign n33749 = ~n33687 & ~n43690;
  assign n33750 = ~n33748 & ~n33749;
  assign n33751 = n4312 & n9678;
  assign n33752 = pi108  & n38376;
  assign n33753 = pi110  & n4314;
  assign n33754 = pi109  & n4322;
  assign n33755 = ~n33753 & ~n33754;
  assign n33756 = ~n33752 & ~n33754;
  assign n33757 = ~n33753 & n33756;
  assign n33758 = ~n33752 & n33755;
  assign n33759 = ~n33751 & n43691;
  assign n33760 = pi56  & ~n33759;
  assign n33761 = pi56  & ~n33760;
  assign n33762 = pi56  & n33759;
  assign n33763 = ~n33759 & ~n33760;
  assign n33764 = ~pi56  & ~n33759;
  assign n33765 = ~n43692 & ~n43693;
  assign n33766 = ~n33750 & n33765;
  assign n33767 = n33750 & ~n33765;
  assign n33768 = n33750 & ~n33767;
  assign n33769 = ~n33765 & ~n33767;
  assign n33770 = ~n33768 & ~n33769;
  assign n33771 = ~n33766 & ~n33767;
  assign n33772 = n33686 & n43694;
  assign n33773 = ~n33686 & ~n43694;
  assign n33774 = ~n33772 & ~n33773;
  assign n33775 = n1971 & n11276;
  assign n33776 = pi111  & n37864;
  assign n33777 = pi113  & n1973;
  assign n33778 = pi112  & n1981;
  assign n33779 = ~n33777 & ~n33778;
  assign n33780 = ~n33776 & ~n33778;
  assign n33781 = ~n33777 & n33780;
  assign n33782 = ~n33776 & n33779;
  assign n33783 = ~n33775 & n43695;
  assign n33784 = pi53  & ~n33783;
  assign n33785 = pi53  & ~n33784;
  assign n33786 = pi53  & n33783;
  assign n33787 = ~n33783 & ~n33784;
  assign n33788 = ~pi53  & ~n33783;
  assign n33789 = ~n43696 & ~n43697;
  assign n33790 = n33774 & ~n33789;
  assign n33791 = ~n33774 & n33789;
  assign n33792 = n33774 & ~n33790;
  assign n33793 = ~n33789 & ~n33790;
  assign n33794 = ~n33792 & ~n33793;
  assign n33795 = ~n33790 & ~n33791;
  assign n33796 = n33685 & n43698;
  assign n33797 = ~n33685 & ~n43698;
  assign n33798 = ~n33796 & ~n33797;
  assign n33799 = n894 & n12530;
  assign n33800 = pi114  & n37580;
  assign n33801 = pi116  & n896;
  assign n33802 = pi115  & n904;
  assign n33803 = ~n33801 & ~n33802;
  assign n33804 = ~n33800 & ~n33802;
  assign n33805 = ~n33801 & n33804;
  assign n33806 = ~n33800 & n33803;
  assign n33807 = ~n33799 & n43699;
  assign n33808 = pi50  & ~n33807;
  assign n33809 = pi50  & ~n33808;
  assign n33810 = pi50  & n33807;
  assign n33811 = ~n33807 & ~n33808;
  assign n33812 = ~pi50  & ~n33807;
  assign n33813 = ~n43700 & ~n43701;
  assign n33814 = ~n33798 & n33813;
  assign n33815 = n33798 & ~n33813;
  assign n33816 = n33798 & ~n33815;
  assign n33817 = ~n33813 & ~n33815;
  assign n33818 = ~n33816 & ~n33817;
  assign n33819 = ~n33814 & ~n33815;
  assign n33820 = ~n33684 & ~n43702;
  assign n33821 = n33684 & n43702;
  assign n33822 = ~n43702 & ~n33820;
  assign n33823 = ~n33684 & ~n33820;
  assign n33824 = ~n33822 & ~n33823;
  assign n33825 = ~n33820 & ~n33821;
  assign n33826 = ~n33683 & ~n43703;
  assign n33827 = n33683 & n43703;
  assign n33828 = ~n43703 & ~n33826;
  assign n33829 = ~n33683 & ~n33826;
  assign n33830 = ~n33828 & ~n33829;
  assign n33831 = ~n33826 & ~n33827;
  assign n33832 = n33668 & n43704;
  assign n33833 = ~n33668 & ~n43704;
  assign n33834 = ~n33832 & ~n33833;
  assign n33835 = n940 & n15049;
  assign n33836 = pi120  & n37541;
  assign n33837 = pi122  & n953;
  assign n33838 = pi121  & n955;
  assign n33839 = ~n33837 & ~n33838;
  assign n33840 = ~n33836 & ~n33838;
  assign n33841 = ~n33837 & n33840;
  assign n33842 = ~n33836 & n33839;
  assign n33843 = ~n33835 & n43705;
  assign n33844 = pi44  & ~n33843;
  assign n33845 = pi44  & ~n33844;
  assign n33846 = pi44  & n33843;
  assign n33847 = ~n33843 & ~n33844;
  assign n33848 = ~pi44  & ~n33843;
  assign n33849 = ~n43706 & ~n43707;
  assign n33850 = n33834 & ~n33849;
  assign n33851 = ~n33834 & n33849;
  assign n33852 = n33834 & ~n33850;
  assign n33853 = ~n33849 & ~n33850;
  assign n33854 = ~n33852 & ~n33853;
  assign n33855 = ~n33850 & ~n33851;
  assign n33856 = n33667 & n43708;
  assign n33857 = ~n33667 & ~n43708;
  assign n33858 = ~n33856 & ~n33857;
  assign n33859 = n733 & n15068;
  assign n33860 = pi123  & n37510;
  assign n33861 = pi125  & n746;
  assign n33862 = pi124  & n748;
  assign n33863 = ~n33861 & ~n33862;
  assign n33864 = ~n33860 & ~n33862;
  assign n33865 = ~n33861 & n33864;
  assign n33866 = ~n33860 & n33863;
  assign n33867 = ~n33859 & n43709;
  assign n33868 = pi41  & ~n33867;
  assign n33869 = pi41  & ~n33868;
  assign n33870 = pi41  & n33867;
  assign n33871 = ~n33867 & ~n33868;
  assign n33872 = ~pi41  & ~n33867;
  assign n33873 = ~n43710 & ~n43711;
  assign n33874 = n33858 & ~n33873;
  assign n33875 = ~n33858 & n33873;
  assign n33876 = ~n33874 & ~n33875;
  assign n33877 = n33666 & ~n33875;
  assign n33878 = ~n33874 & n33877;
  assign n33879 = n33666 & n33876;
  assign n33880 = ~n33666 & ~n33876;
  assign n33881 = n33666 & ~n43712;
  assign n33882 = ~n33875 & ~n43712;
  assign n33883 = ~n33874 & n33882;
  assign n33884 = n33876 & ~n43712;
  assign n33885 = ~n33881 & ~n43713;
  assign n33886 = ~n43712 & ~n33880;
  assign n33887 = n33651 & n43714;
  assign n33888 = ~n33651 & ~n43714;
  assign n33889 = ~n33887 & ~n33888;
  assign n33890 = ~n33645 & ~n33648;
  assign n33891 = n33889 & ~n33890;
  assign n33892 = ~n33889 & n33890;
  assign po100  = ~n33891 & ~n33892;
  assign n33894 = ~n33888 & ~n33891;
  assign n33895 = ~n33664 & ~n43712;
  assign n33896 = ~n33857 & ~n33874;
  assign n33897 = n691 & ~n18675;
  assign n33898 = ~n37503 & ~n33897;
  assign n33899 = pi127  & n37503;
  assign n33900 = n691 & n18680;
  assign n33901 = ~n33899 & ~n33900;
  assign n33902 = pi127  & ~n33898;
  assign n33903 = pi38  & ~n43715;
  assign n33904 = pi38  & ~n33903;
  assign n33905 = pi38  & n43715;
  assign n33906 = ~n43715 & ~n33903;
  assign n33907 = ~pi38  & ~n43715;
  assign n33908 = ~n43716 & ~n43717;
  assign n33909 = ~n33896 & ~n33908;
  assign n33910 = n33896 & n33908;
  assign n33911 = ~n33896 & ~n33909;
  assign n33912 = ~n33908 & ~n33909;
  assign n33913 = ~n33911 & ~n33912;
  assign n33914 = ~n33909 & ~n33910;
  assign n33915 = ~n33820 & ~n33826;
  assign n33916 = n785 & n14913;
  assign n33917 = pi118  & n37520;
  assign n33918 = pi120  & n787;
  assign n33919 = pi119  & n795;
  assign n33920 = ~n33918 & ~n33919;
  assign n33921 = ~n33917 & ~n33919;
  assign n33922 = ~n33918 & n33921;
  assign n33923 = ~n33917 & n33920;
  assign n33924 = ~n33916 & n43719;
  assign n33925 = pi47  & ~n33924;
  assign n33926 = pi47  & ~n33925;
  assign n33927 = pi47  & n33924;
  assign n33928 = ~n33924 & ~n33925;
  assign n33929 = ~pi47  & ~n33924;
  assign n33930 = ~n43720 & ~n43721;
  assign n33931 = n894 & n13079;
  assign n33932 = pi115  & n37580;
  assign n33933 = pi117  & n896;
  assign n33934 = pi116  & n904;
  assign n33935 = ~n33933 & ~n33934;
  assign n33936 = ~n33932 & ~n33934;
  assign n33937 = ~n33933 & n33936;
  assign n33938 = ~n33932 & n33935;
  assign n33939 = ~n33931 & n43722;
  assign n33940 = pi50  & ~n33939;
  assign n33941 = pi50  & ~n33940;
  assign n33942 = pi50  & n33939;
  assign n33943 = ~n33939 & ~n33940;
  assign n33944 = ~pi50  & ~n33939;
  assign n33945 = ~n43723 & ~n43724;
  assign n33946 = n7882 & n9277;
  assign n33947 = pi106  & n39128;
  assign n33948 = pi108  & n7884;
  assign n33949 = pi107  & n7892;
  assign n33950 = ~n33948 & ~n33949;
  assign n33951 = ~n33947 & ~n33949;
  assign n33952 = ~n33948 & n33951;
  assign n33953 = ~n33947 & n33950;
  assign n33954 = ~n33946 & n43725;
  assign n33955 = pi59  & ~n33954;
  assign n33956 = pi59  & ~n33955;
  assign n33957 = pi59  & n33954;
  assign n33958 = ~n33954 & ~n33955;
  assign n33959 = ~pi59  & ~n33954;
  assign n33960 = ~n43726 & ~n43727;
  assign n33961 = n8229 & n12674;
  assign n33962 = pi103  & n40107;
  assign n33963 = pi105  & n12676;
  assign n33964 = pi104  & n12684;
  assign n33965 = ~n33963 & ~n33964;
  assign n33966 = ~n33962 & ~n33964;
  assign n33967 = ~n33963 & n33966;
  assign n33968 = ~n33962 & n33965;
  assign n33969 = ~n33961 & n43728;
  assign n33970 = pi62  & ~n33969;
  assign n33971 = pi62  & ~n33970;
  assign n33972 = pi62  & n33969;
  assign n33973 = ~n33969 & ~n33970;
  assign n33974 = ~pi62  & ~n33969;
  assign n33975 = ~n43729 & ~n43730;
  assign n33976 = ~n33708 & ~n33716;
  assign n33977 = pi102  & ~n40814;
  assign n33978 = pi101  & n18285;
  assign n33979 = ~n33977 & ~n33978;
  assign n33980 = n33707 & ~n33979;
  assign n33981 = ~n33707 & n33979;
  assign n33982 = n33707 & ~n33980;
  assign n33983 = n33707 & n33979;
  assign n33984 = ~n33979 & ~n33980;
  assign n33985 = ~n33707 & ~n33979;
  assign n33986 = ~n43731 & ~n43732;
  assign n33987 = ~n33980 & ~n33981;
  assign n33988 = ~n33976 & ~n43733;
  assign n33989 = n33976 & n43733;
  assign n33990 = ~n33976 & ~n33988;
  assign n33991 = ~n33976 & n43733;
  assign n33992 = ~n43733 & ~n33988;
  assign n33993 = n33976 & ~n43733;
  assign n33994 = ~n43734 & ~n43735;
  assign n33995 = ~n33988 & ~n33989;
  assign n33996 = ~n33975 & ~n43736;
  assign n33997 = n33975 & n43736;
  assign n33998 = ~n43736 & ~n33996;
  assign n33999 = ~n33975 & ~n33996;
  assign n34000 = ~n33998 & ~n33999;
  assign n34001 = ~n33996 & ~n33997;
  assign n34002 = n33960 & n43737;
  assign n34003 = ~n33960 & ~n43737;
  assign n34004 = n33960 & ~n43737;
  assign n34005 = ~n33960 & n43737;
  assign n34006 = ~n34004 & ~n34005;
  assign n34007 = ~n34002 & ~n34003;
  assign n34008 = ~n33725 & n33741;
  assign n34009 = ~n33725 & ~n33742;
  assign n34010 = ~n33724 & ~n34008;
  assign n34011 = n43738 & n43739;
  assign n34012 = ~n43738 & ~n43739;
  assign n34013 = ~n34011 & ~n34012;
  assign n34014 = n565 & n4312;
  assign n34015 = pi109  & n38376;
  assign n34016 = pi111  & n4314;
  assign n34017 = pi110  & n4322;
  assign n34018 = ~n34016 & ~n34017;
  assign n34019 = ~n34015 & ~n34017;
  assign n34020 = ~n34016 & n34019;
  assign n34021 = ~n34015 & n34018;
  assign n34022 = ~n34014 & n43740;
  assign n34023 = pi56  & ~n34022;
  assign n34024 = pi56  & ~n34023;
  assign n34025 = pi56  & n34022;
  assign n34026 = ~n34022 & ~n34023;
  assign n34027 = ~pi56  & ~n34022;
  assign n34028 = ~n43741 & ~n43742;
  assign n34029 = ~n34013 & n34028;
  assign n34030 = n34013 & ~n34028;
  assign n34031 = n34013 & ~n34030;
  assign n34032 = ~n34028 & ~n34030;
  assign n34033 = ~n34031 & ~n34032;
  assign n34034 = ~n34029 & ~n34030;
  assign n34035 = ~n33749 & n33765;
  assign n34036 = ~n33749 & ~n33767;
  assign n34037 = ~n33748 & ~n34035;
  assign n34038 = n43743 & n43744;
  assign n34039 = ~n43743 & ~n43744;
  assign n34040 = ~n34038 & ~n34039;
  assign n34041 = n1971 & n11258;
  assign n34042 = pi112  & n37864;
  assign n34043 = pi114  & n1973;
  assign n34044 = pi113  & n1981;
  assign n34045 = ~n34043 & ~n34044;
  assign n34046 = ~n34042 & ~n34044;
  assign n34047 = ~n34043 & n34046;
  assign n34048 = ~n34042 & n34045;
  assign n34049 = ~n34041 & n43745;
  assign n34050 = pi53  & ~n34049;
  assign n34051 = pi53  & ~n34050;
  assign n34052 = pi53  & n34049;
  assign n34053 = ~n34049 & ~n34050;
  assign n34054 = ~pi53  & ~n34049;
  assign n34055 = ~n43746 & ~n43747;
  assign n34056 = ~n34040 & n34055;
  assign n34057 = n34040 & ~n34055;
  assign n34058 = ~n34056 & ~n34057;
  assign n34059 = ~n33773 & n33789;
  assign n34060 = ~n33773 & ~n33790;
  assign n34061 = ~n33772 & ~n34059;
  assign n34062 = n34058 & ~n43748;
  assign n34063 = ~n34058 & n43748;
  assign n34064 = ~n43748 & ~n34062;
  assign n34065 = n34058 & ~n34062;
  assign n34066 = ~n34064 & ~n34065;
  assign n34067 = ~n34062 & ~n34063;
  assign n34068 = ~n33945 & ~n43749;
  assign n34069 = n33945 & ~n34065;
  assign n34070 = ~n34064 & n34069;
  assign n34071 = n33945 & n43749;
  assign n34072 = ~n34068 & ~n43750;
  assign n34073 = ~n33797 & n33813;
  assign n34074 = ~n33797 & ~n33815;
  assign n34075 = ~n33796 & ~n34073;
  assign n34076 = n34072 & ~n43751;
  assign n34077 = ~n34072 & n43751;
  assign n34078 = ~n34076 & ~n34077;
  assign n34079 = ~n33930 & n34078;
  assign n34080 = n33930 & ~n34078;
  assign n34081 = ~n34079 & ~n34080;
  assign n34082 = ~n33915 & n34081;
  assign n34083 = n33915 & ~n34081;
  assign n34084 = ~n34082 & ~n34083;
  assign n34085 = n940 & n14961;
  assign n34086 = pi121  & n37541;
  assign n34087 = pi123  & n953;
  assign n34088 = pi122  & n955;
  assign n34089 = ~n34087 & ~n34088;
  assign n34090 = ~n34086 & ~n34088;
  assign n34091 = ~n34087 & n34090;
  assign n34092 = ~n34086 & n34089;
  assign n34093 = ~n34085 & n43752;
  assign n34094 = pi44  & ~n34093;
  assign n34095 = pi44  & ~n34094;
  assign n34096 = pi44  & n34093;
  assign n34097 = ~n34093 & ~n34094;
  assign n34098 = ~pi44  & ~n34093;
  assign n34099 = ~n43753 & ~n43754;
  assign n34100 = n34084 & ~n34099;
  assign n34101 = ~n34084 & n34099;
  assign n34102 = n34084 & ~n34100;
  assign n34103 = ~n34099 & ~n34100;
  assign n34104 = ~n34102 & ~n34103;
  assign n34105 = ~n34100 & ~n34101;
  assign n34106 = ~n33833 & n33849;
  assign n34107 = ~n33833 & ~n33850;
  assign n34108 = ~n33832 & ~n34106;
  assign n34109 = n43755 & n43756;
  assign n34110 = ~n43755 & ~n43756;
  assign n34111 = ~n34109 & ~n34110;
  assign n34112 = n733 & n15021;
  assign n34113 = pi124  & n37510;
  assign n34114 = pi126  & n746;
  assign n34115 = pi125  & n748;
  assign n34116 = ~n34114 & ~n34115;
  assign n34117 = ~n34113 & ~n34115;
  assign n34118 = ~n34114 & n34117;
  assign n34119 = ~n34113 & n34116;
  assign n34120 = ~n34112 & n43757;
  assign n34121 = pi41  & ~n34120;
  assign n34122 = pi41  & ~n34121;
  assign n34123 = pi41  & n34120;
  assign n34124 = ~n34120 & ~n34121;
  assign n34125 = ~pi41  & ~n34120;
  assign n34126 = ~n43758 & ~n43759;
  assign n34127 = ~n34111 & n34126;
  assign n34128 = n34111 & ~n34126;
  assign n34129 = n34111 & ~n34128;
  assign n34130 = ~n34126 & ~n34128;
  assign n34131 = ~n34129 & ~n34130;
  assign n34132 = ~n34127 & ~n34128;
  assign n34133 = ~n43718 & ~n43760;
  assign n34134 = n43718 & n43760;
  assign n34135 = ~n43718 & n43760;
  assign n34136 = n43718 & ~n43760;
  assign n34137 = ~n34135 & ~n34136;
  assign n34138 = ~n34133 & ~n34134;
  assign n34139 = ~n33895 & ~n43761;
  assign n34140 = n33895 & n43761;
  assign n34141 = ~n34139 & ~n34140;
  assign n34142 = ~n33894 & n34141;
  assign n34143 = n33894 & ~n34141;
  assign po101  = ~n34142 & ~n34143;
  assign n34145 = ~n34139 & ~n34142;
  assign n34146 = ~n34076 & ~n34079;
  assign n34147 = ~n34062 & ~n34068;
  assign n34148 = n894 & n13057;
  assign n34149 = pi116  & n37580;
  assign n34150 = pi118  & n896;
  assign n34151 = pi117  & n904;
  assign n34152 = ~n34150 & ~n34151;
  assign n34153 = ~n34149 & ~n34151;
  assign n34154 = ~n34150 & n34153;
  assign n34155 = ~n34149 & n34152;
  assign n34156 = ~n34148 & n43762;
  assign n34157 = pi50  & ~n34156;
  assign n34158 = pi50  & ~n34157;
  assign n34159 = pi50  & n34156;
  assign n34160 = ~n34156 & ~n34157;
  assign n34161 = ~pi50  & ~n34156;
  assign n34162 = ~n43763 & ~n43764;
  assign n34163 = ~n34039 & ~n34057;
  assign n34164 = n4312 & n10844;
  assign n34165 = pi110  & n38376;
  assign n34166 = pi112  & n4314;
  assign n34167 = pi111  & n4322;
  assign n34168 = ~n34166 & ~n34167;
  assign n34169 = ~n34165 & ~n34167;
  assign n34170 = ~n34166 & n34169;
  assign n34171 = ~n34165 & n34168;
  assign n34172 = ~n34164 & n43765;
  assign n34173 = pi56  & ~n34172;
  assign n34174 = pi56  & ~n34173;
  assign n34175 = pi56  & n34172;
  assign n34176 = ~n34172 & ~n34173;
  assign n34177 = ~pi56  & ~n34172;
  assign n34178 = ~n43766 & ~n43767;
  assign n34179 = n7882 & n9701;
  assign n34180 = pi107  & n39128;
  assign n34181 = pi109  & n7884;
  assign n34182 = pi108  & n7892;
  assign n34183 = ~n34181 & ~n34182;
  assign n34184 = ~n34180 & ~n34182;
  assign n34185 = ~n34181 & n34184;
  assign n34186 = ~n34180 & n34183;
  assign n34187 = ~n34179 & n43768;
  assign n34188 = pi59  & ~n34187;
  assign n34189 = pi59  & ~n34188;
  assign n34190 = pi59  & n34187;
  assign n34191 = ~n34187 & ~n34188;
  assign n34192 = ~pi59  & ~n34187;
  assign n34193 = ~n43769 & ~n43770;
  assign n34194 = ~n33980 & ~n33988;
  assign n34195 = ~pi38  & ~n33707;
  assign n34196 = pi38  & n33707;
  assign n34197 = pi38  & ~n33707;
  assign n34198 = ~pi38  & n33707;
  assign n34199 = ~n34197 & ~n34198;
  assign n34200 = ~n34195 & ~n34196;
  assign n34201 = pi103  & ~n40814;
  assign n34202 = pi102  & n18285;
  assign n34203 = ~n34201 & ~n34202;
  assign n34204 = ~n43771 & ~n34203;
  assign n34205 = n43771 & n34203;
  assign n34206 = ~n34204 & ~n34205;
  assign n34207 = ~n34194 & n34206;
  assign n34208 = n34194 & ~n34206;
  assign n34209 = ~n34207 & ~n34208;
  assign n34210 = n8209 & n12674;
  assign n34211 = pi104  & n40107;
  assign n34212 = pi106  & n12676;
  assign n34213 = pi105  & n12684;
  assign n34214 = ~n34212 & ~n34213;
  assign n34215 = ~n34211 & ~n34213;
  assign n34216 = ~n34212 & n34215;
  assign n34217 = ~n34211 & n34214;
  assign n34218 = ~n34210 & n43772;
  assign n34219 = pi62  & ~n34218;
  assign n34220 = pi62  & ~n34219;
  assign n34221 = pi62  & n34218;
  assign n34222 = ~n34218 & ~n34219;
  assign n34223 = ~pi62  & ~n34218;
  assign n34224 = ~n43773 & ~n43774;
  assign n34225 = n34209 & ~n34224;
  assign n34226 = ~n34209 & n34224;
  assign n34227 = n34209 & ~n34225;
  assign n34228 = ~n34224 & ~n34225;
  assign n34229 = ~n34227 & ~n34228;
  assign n34230 = ~n34225 & ~n34226;
  assign n34231 = ~n34193 & ~n43775;
  assign n34232 = n34193 & n43775;
  assign n34233 = ~n43775 & ~n34231;
  assign n34234 = ~n34193 & ~n34231;
  assign n34235 = ~n34233 & ~n34234;
  assign n34236 = ~n34231 & ~n34232;
  assign n34237 = n33960 & ~n33996;
  assign n34238 = ~n33996 & ~n34003;
  assign n34239 = ~n33997 & ~n34237;
  assign n34240 = ~n43776 & ~n43777;
  assign n34241 = n43776 & n43777;
  assign n34242 = ~n43776 & ~n34240;
  assign n34243 = ~n43777 & ~n34240;
  assign n34244 = ~n34242 & ~n34243;
  assign n34245 = ~n34240 & ~n34241;
  assign n34246 = ~n34178 & ~n43778;
  assign n34247 = n34178 & n43778;
  assign n34248 = ~n43778 & ~n34246;
  assign n34249 = n34178 & ~n43778;
  assign n34250 = ~n34178 & ~n34246;
  assign n34251 = ~n34178 & n43778;
  assign n34252 = ~n43779 & ~n43780;
  assign n34253 = ~n34246 & ~n34247;
  assign n34254 = ~n34012 & n34028;
  assign n34255 = ~n34012 & ~n34030;
  assign n34256 = ~n34011 & ~n34254;
  assign n34257 = n43781 & n43782;
  assign n34258 = ~n43781 & ~n43782;
  assign n34259 = ~n34257 & ~n34258;
  assign n34260 = n523 & n1971;
  assign n34261 = pi113  & n37864;
  assign n34262 = pi115  & n1973;
  assign n34263 = pi114  & n1981;
  assign n34264 = ~n34262 & ~n34263;
  assign n34265 = ~n34261 & ~n34263;
  assign n34266 = ~n34262 & n34265;
  assign n34267 = ~n34261 & n34264;
  assign n34268 = ~n34260 & n43783;
  assign n34269 = pi53  & ~n34268;
  assign n34270 = pi53  & ~n34269;
  assign n34271 = pi53  & n34268;
  assign n34272 = ~n34268 & ~n34269;
  assign n34273 = ~pi53  & ~n34268;
  assign n34274 = ~n43784 & ~n43785;
  assign n34275 = ~n34259 & n34274;
  assign n34276 = n34259 & ~n34274;
  assign n34277 = ~n34275 & ~n34276;
  assign n34278 = ~n34163 & n34277;
  assign n34279 = n34163 & ~n34277;
  assign n34280 = ~n34278 & ~n34279;
  assign n34281 = ~n34162 & n34280;
  assign n34282 = n34162 & ~n34280;
  assign n34283 = ~n34281 & ~n34282;
  assign n34284 = ~n34147 & n34283;
  assign n34285 = n34147 & ~n34283;
  assign n34286 = ~n34284 & ~n34285;
  assign n34287 = n785 & n15091;
  assign n34288 = pi119  & n37520;
  assign n34289 = pi121  & n787;
  assign n34290 = pi120  & n795;
  assign n34291 = ~n34289 & ~n34290;
  assign n34292 = ~n34288 & ~n34290;
  assign n34293 = ~n34289 & n34292;
  assign n34294 = ~n34288 & n34291;
  assign n34295 = ~n34287 & n43786;
  assign n34296 = pi47  & ~n34295;
  assign n34297 = pi47  & ~n34296;
  assign n34298 = pi47  & n34295;
  assign n34299 = ~n34295 & ~n34296;
  assign n34300 = ~pi47  & ~n34295;
  assign n34301 = ~n43787 & ~n43788;
  assign n34302 = n34286 & ~n34301;
  assign n34303 = ~n34286 & n34301;
  assign n34304 = n34286 & ~n34302;
  assign n34305 = n34286 & n34301;
  assign n34306 = ~n34301 & ~n34302;
  assign n34307 = ~n34286 & ~n34301;
  assign n34308 = ~n43789 & ~n43790;
  assign n34309 = ~n34302 & ~n34303;
  assign n34310 = n34146 & n43791;
  assign n34311 = ~n34146 & ~n43791;
  assign n34312 = ~n34310 & ~n34311;
  assign n34313 = n940 & n15111;
  assign n34314 = pi122  & n37541;
  assign n34315 = pi124  & n953;
  assign n34316 = pi123  & n955;
  assign n34317 = ~n34315 & ~n34316;
  assign n34318 = ~n34314 & ~n34316;
  assign n34319 = ~n34315 & n34318;
  assign n34320 = ~n34314 & n34317;
  assign n34321 = ~n34313 & n43792;
  assign n34322 = pi44  & ~n34321;
  assign n34323 = pi44  & ~n34322;
  assign n34324 = pi44  & n34321;
  assign n34325 = ~n34321 & ~n34322;
  assign n34326 = ~pi44  & ~n34321;
  assign n34327 = ~n43793 & ~n43794;
  assign n34328 = n34312 & ~n34327;
  assign n34329 = ~n34312 & n34327;
  assign n34330 = n34312 & ~n34328;
  assign n34331 = n34312 & n34327;
  assign n34332 = ~n34327 & ~n34328;
  assign n34333 = ~n34312 & ~n34327;
  assign n34334 = ~n43795 & ~n43796;
  assign n34335 = ~n34328 & ~n34329;
  assign n34336 = ~n34082 & n34099;
  assign n34337 = ~n34082 & ~n34100;
  assign n34338 = ~n34083 & ~n34336;
  assign n34339 = n43797 & n43798;
  assign n34340 = ~n43797 & ~n43798;
  assign n34341 = ~n34339 & ~n34340;
  assign n34342 = n733 & n40885;
  assign n34343 = pi125  & n37510;
  assign n34344 = pi127  & n746;
  assign n34345 = pi126  & n748;
  assign n34346 = ~n34344 & ~n34345;
  assign n34347 = ~n34343 & ~n34345;
  assign n34348 = ~n34344 & n34347;
  assign n34349 = ~n34343 & n34346;
  assign n34350 = ~n34342 & n43799;
  assign n34351 = pi41  & ~n34350;
  assign n34352 = pi41  & ~n34351;
  assign n34353 = pi41  & n34350;
  assign n34354 = ~n34350 & ~n34351;
  assign n34355 = ~pi41  & ~n34350;
  assign n34356 = ~n43800 & ~n43801;
  assign n34357 = n34341 & ~n34356;
  assign n34358 = ~n34341 & n34356;
  assign n34359 = n34341 & ~n34357;
  assign n34360 = n34341 & n34356;
  assign n34361 = ~n34356 & ~n34357;
  assign n34362 = ~n34341 & ~n34356;
  assign n34363 = ~n43802 & ~n43803;
  assign n34364 = ~n34357 & ~n34358;
  assign n34365 = ~n34110 & n34126;
  assign n34366 = ~n34110 & ~n34128;
  assign n34367 = ~n34109 & ~n34365;
  assign n34368 = n43804 & n43805;
  assign n34369 = ~n43804 & ~n43805;
  assign n34370 = ~n34368 & ~n34369;
  assign n34371 = ~n33909 & n43760;
  assign n34372 = ~n33909 & ~n34133;
  assign n34373 = ~n33910 & ~n34371;
  assign n34374 = n34370 & ~n43806;
  assign n34375 = ~n34370 & n43806;
  assign n34376 = ~n34374 & ~n34375;
  assign n34377 = ~n34145 & n34376;
  assign n34378 = n34145 & ~n34376;
  assign po102  = ~n34377 & ~n34378;
  assign n34380 = ~n34357 & ~n34369;
  assign n34381 = ~n34328 & ~n34340;
  assign n34382 = n733 & n40891;
  assign n34383 = pi126  & n37510;
  assign n34384 = pi127  & n748;
  assign n34385 = ~n34383 & ~n34384;
  assign n34386 = ~n733 & n34385;
  assign n34387 = ~n40891 & n34385;
  assign n34388 = ~n34386 & ~n34387;
  assign n34389 = ~n34382 & n34385;
  assign n34390 = pi41  & ~n43807;
  assign n34391 = ~pi41  & n43807;
  assign n34392 = ~n34390 & ~n34391;
  assign n34393 = ~n34381 & ~n34392;
  assign n34394 = n34381 & n34392;
  assign n34395 = ~n34393 & ~n34394;
  assign n34396 = ~n34302 & ~n34311;
  assign n34397 = ~n34281 & ~n34284;
  assign n34398 = n894 & n13027;
  assign n34399 = pi117  & n37580;
  assign n34400 = pi119  & n896;
  assign n34401 = pi118  & n904;
  assign n34402 = ~n34400 & ~n34401;
  assign n34403 = ~n34399 & ~n34401;
  assign n34404 = ~n34400 & n34403;
  assign n34405 = ~n34399 & n34402;
  assign n34406 = ~n34398 & n43808;
  assign n34407 = pi50  & ~n34406;
  assign n34408 = pi50  & ~n34407;
  assign n34409 = pi50  & n34406;
  assign n34410 = ~n34406 & ~n34407;
  assign n34411 = ~pi50  & ~n34406;
  assign n34412 = ~n43809 & ~n43810;
  assign n34413 = ~n34276 & ~n34278;
  assign n34414 = ~n34246 & ~n34258;
  assign n34415 = ~n34231 & ~n34240;
  assign n34416 = ~n34195 & ~n34204;
  assign n34417 = pi104  & ~n40814;
  assign n34418 = pi103  & n18285;
  assign n34419 = ~n34417 & ~n34418;
  assign n34420 = ~n34416 & n34419;
  assign n34421 = n34416 & ~n34419;
  assign n34422 = ~n34420 & ~n34421;
  assign n34423 = n8177 & n12674;
  assign n34424 = pi105  & n40107;
  assign n34425 = pi107  & n12676;
  assign n34426 = pi106  & n12684;
  assign n34427 = ~n34425 & ~n34426;
  assign n34428 = ~n34424 & ~n34426;
  assign n34429 = ~n34425 & n34428;
  assign n34430 = ~n34424 & n34427;
  assign n34431 = ~n12674 & n43811;
  assign n34432 = ~n8177 & n43811;
  assign n34433 = ~n34431 & ~n34432;
  assign n34434 = ~n34423 & n43811;
  assign n34435 = pi62  & ~n43812;
  assign n34436 = ~pi62  & n43812;
  assign n34437 = ~n34435 & ~n34436;
  assign n34438 = n34422 & ~n34437;
  assign n34439 = ~n34422 & n34437;
  assign n34440 = ~n34438 & ~n34439;
  assign n34441 = ~n34207 & n34224;
  assign n34442 = ~n34207 & ~n34225;
  assign n34443 = ~n34208 & ~n34441;
  assign n34444 = n34440 & ~n43813;
  assign n34445 = ~n34440 & n43813;
  assign n34446 = ~n34444 & ~n34445;
  assign n34447 = n7882 & n9678;
  assign n34448 = pi108  & n39128;
  assign n34449 = pi110  & n7884;
  assign n34450 = pi109  & n7892;
  assign n34451 = ~n34449 & ~n34450;
  assign n34452 = ~n34448 & ~n34450;
  assign n34453 = ~n34449 & n34452;
  assign n34454 = ~n34448 & n34451;
  assign n34455 = ~n34447 & n43814;
  assign n34456 = pi59  & ~n34455;
  assign n34457 = pi59  & ~n34456;
  assign n34458 = pi59  & n34455;
  assign n34459 = ~n34455 & ~n34456;
  assign n34460 = ~pi59  & ~n34455;
  assign n34461 = ~n43815 & ~n43816;
  assign n34462 = n34446 & ~n34461;
  assign n34463 = ~n34446 & n34461;
  assign n34464 = n34446 & ~n34462;
  assign n34465 = ~n34461 & ~n34462;
  assign n34466 = ~n34464 & ~n34465;
  assign n34467 = ~n34462 & ~n34463;
  assign n34468 = n34415 & n43817;
  assign n34469 = ~n34415 & ~n43817;
  assign n34470 = ~n34468 & ~n34469;
  assign n34471 = n4312 & n11276;
  assign n34472 = pi111  & n38376;
  assign n34473 = pi113  & n4314;
  assign n34474 = pi112  & n4322;
  assign n34475 = ~n34473 & ~n34474;
  assign n34476 = ~n34472 & ~n34474;
  assign n34477 = ~n34473 & n34476;
  assign n34478 = ~n34472 & n34475;
  assign n34479 = ~n34471 & n43818;
  assign n34480 = pi56  & ~n34479;
  assign n34481 = pi56  & ~n34480;
  assign n34482 = pi56  & n34479;
  assign n34483 = ~n34479 & ~n34480;
  assign n34484 = ~pi56  & ~n34479;
  assign n34485 = ~n43819 & ~n43820;
  assign n34486 = ~n34470 & n34485;
  assign n34487 = n34470 & ~n34485;
  assign n34488 = n34470 & ~n34487;
  assign n34489 = ~n34485 & ~n34487;
  assign n34490 = ~n34488 & ~n34489;
  assign n34491 = ~n34486 & ~n34487;
  assign n34492 = n34414 & n43821;
  assign n34493 = ~n34414 & ~n43821;
  assign n34494 = ~n34492 & ~n34493;
  assign n34495 = n1971 & n12530;
  assign n34496 = pi114  & n37864;
  assign n34497 = pi116  & n1973;
  assign n34498 = pi115  & n1981;
  assign n34499 = ~n34497 & ~n34498;
  assign n34500 = ~n34496 & ~n34498;
  assign n34501 = ~n34497 & n34500;
  assign n34502 = ~n34496 & n34499;
  assign n34503 = ~n34495 & n43822;
  assign n34504 = pi53  & ~n34503;
  assign n34505 = pi53  & ~n34504;
  assign n34506 = pi53  & n34503;
  assign n34507 = ~n34503 & ~n34504;
  assign n34508 = ~pi53  & ~n34503;
  assign n34509 = ~n43823 & ~n43824;
  assign n34510 = n34494 & ~n34509;
  assign n34511 = ~n34494 & n34509;
  assign n34512 = n34494 & ~n34510;
  assign n34513 = ~n34509 & ~n34510;
  assign n34514 = ~n34512 & ~n34513;
  assign n34515 = ~n34510 & ~n34511;
  assign n34516 = ~n34413 & ~n43825;
  assign n34517 = n34413 & n43825;
  assign n34518 = ~n43825 & ~n34516;
  assign n34519 = ~n34413 & ~n34516;
  assign n34520 = ~n34518 & ~n34519;
  assign n34521 = ~n34516 & ~n34517;
  assign n34522 = ~n34412 & ~n43826;
  assign n34523 = n34412 & n43826;
  assign n34524 = ~n43826 & ~n34522;
  assign n34525 = ~n34412 & ~n34522;
  assign n34526 = ~n34524 & ~n34525;
  assign n34527 = ~n34522 & ~n34523;
  assign n34528 = n34397 & n43827;
  assign n34529 = ~n34397 & ~n43827;
  assign n34530 = ~n34528 & ~n34529;
  assign n34531 = n785 & n15049;
  assign n34532 = pi120  & n37520;
  assign n34533 = pi122  & n787;
  assign n34534 = pi121  & n795;
  assign n34535 = ~n34533 & ~n34534;
  assign n34536 = ~n34532 & ~n34534;
  assign n34537 = ~n34533 & n34536;
  assign n34538 = ~n34532 & n34535;
  assign n34539 = ~n34531 & n43828;
  assign n34540 = pi47  & ~n34539;
  assign n34541 = pi47  & ~n34540;
  assign n34542 = pi47  & n34539;
  assign n34543 = ~n34539 & ~n34540;
  assign n34544 = ~pi47  & ~n34539;
  assign n34545 = ~n43829 & ~n43830;
  assign n34546 = n34530 & ~n34545;
  assign n34547 = ~n34530 & n34545;
  assign n34548 = n34530 & ~n34546;
  assign n34549 = ~n34545 & ~n34546;
  assign n34550 = ~n34548 & ~n34549;
  assign n34551 = ~n34546 & ~n34547;
  assign n34552 = n34396 & n43831;
  assign n34553 = ~n34396 & ~n43831;
  assign n34554 = ~n34552 & ~n34553;
  assign n34555 = n940 & n15068;
  assign n34556 = pi123  & n37541;
  assign n34557 = pi125  & n953;
  assign n34558 = pi124  & n955;
  assign n34559 = ~n34557 & ~n34558;
  assign n34560 = ~n34556 & ~n34558;
  assign n34561 = ~n34557 & n34560;
  assign n34562 = ~n34556 & n34559;
  assign n34563 = ~n34555 & n43832;
  assign n34564 = pi44  & ~n34563;
  assign n34565 = pi44  & ~n34564;
  assign n34566 = pi44  & n34563;
  assign n34567 = ~n34563 & ~n34564;
  assign n34568 = ~pi44  & ~n34563;
  assign n34569 = ~n43833 & ~n43834;
  assign n34570 = n34554 & ~n34569;
  assign n34571 = ~n34554 & n34569;
  assign n34572 = ~n34570 & ~n34571;
  assign n34573 = n34395 & ~n34571;
  assign n34574 = ~n34570 & n34573;
  assign n34575 = n34395 & n34572;
  assign n34576 = ~n34395 & ~n34572;
  assign n34577 = n34395 & ~n43835;
  assign n34578 = ~n34571 & ~n43835;
  assign n34579 = ~n34570 & n34578;
  assign n34580 = n34572 & ~n43835;
  assign n34581 = ~n34577 & ~n43836;
  assign n34582 = ~n43835 & ~n34576;
  assign n34583 = n34380 & n43837;
  assign n34584 = ~n34380 & ~n43837;
  assign n34585 = ~n34583 & ~n34584;
  assign n34586 = ~n34374 & ~n34377;
  assign n34587 = n34585 & ~n34586;
  assign n34588 = ~n34585 & n34586;
  assign po103  = ~n34587 & ~n34588;
  assign n34590 = ~n34584 & ~n34587;
  assign n34591 = ~n34393 & ~n43835;
  assign n34592 = ~n34553 & ~n34570;
  assign n34593 = n733 & ~n18675;
  assign n34594 = ~n37510 & ~n34593;
  assign n34595 = pi127  & n37510;
  assign n34596 = n733 & n18680;
  assign n34597 = ~n34595 & ~n34596;
  assign n34598 = pi127  & ~n34594;
  assign n34599 = pi41  & ~n43838;
  assign n34600 = pi41  & ~n34599;
  assign n34601 = pi41  & n43838;
  assign n34602 = ~n43838 & ~n34599;
  assign n34603 = ~pi41  & ~n43838;
  assign n34604 = ~n43839 & ~n43840;
  assign n34605 = ~n34592 & ~n34604;
  assign n34606 = n34592 & n34604;
  assign n34607 = ~n34592 & ~n34605;
  assign n34608 = ~n34604 & ~n34605;
  assign n34609 = ~n34607 & ~n34608;
  assign n34610 = ~n34605 & ~n34606;
  assign n34611 = ~n34516 & ~n34522;
  assign n34612 = n894 & n14913;
  assign n34613 = pi118  & n37580;
  assign n34614 = pi120  & n896;
  assign n34615 = pi119  & n904;
  assign n34616 = ~n34614 & ~n34615;
  assign n34617 = ~n34613 & ~n34615;
  assign n34618 = ~n34614 & n34617;
  assign n34619 = ~n34613 & n34616;
  assign n34620 = ~n34612 & n43842;
  assign n34621 = pi50  & ~n34620;
  assign n34622 = pi50  & ~n34621;
  assign n34623 = pi50  & n34620;
  assign n34624 = ~n34620 & ~n34621;
  assign n34625 = ~pi50  & ~n34620;
  assign n34626 = ~n43843 & ~n43844;
  assign n34627 = n1971 & n13079;
  assign n34628 = pi115  & n37864;
  assign n34629 = pi117  & n1973;
  assign n34630 = pi116  & n1981;
  assign n34631 = ~n34629 & ~n34630;
  assign n34632 = ~n34628 & ~n34630;
  assign n34633 = ~n34629 & n34632;
  assign n34634 = ~n34628 & n34631;
  assign n34635 = ~n34627 & n43845;
  assign n34636 = pi53  & ~n34635;
  assign n34637 = pi53  & ~n34636;
  assign n34638 = pi53  & n34635;
  assign n34639 = ~n34635 & ~n34636;
  assign n34640 = ~pi53  & ~n34635;
  assign n34641 = ~n43846 & ~n43847;
  assign n34642 = n565 & n7882;
  assign n34643 = pi109  & n39128;
  assign n34644 = pi111  & n7884;
  assign n34645 = pi110  & n7892;
  assign n34646 = ~n34644 & ~n34645;
  assign n34647 = ~n34643 & ~n34645;
  assign n34648 = ~n34644 & n34647;
  assign n34649 = ~n34643 & n34646;
  assign n34650 = ~n34642 & n43848;
  assign n34651 = pi59  & ~n34650;
  assign n34652 = pi59  & ~n34651;
  assign n34653 = pi59  & n34650;
  assign n34654 = ~n34650 & ~n34651;
  assign n34655 = ~pi59  & ~n34650;
  assign n34656 = ~n43849 & ~n43850;
  assign n34657 = n9277 & n12674;
  assign n34658 = pi106  & n40107;
  assign n34659 = pi108  & n12676;
  assign n34660 = pi107  & n12684;
  assign n34661 = ~n34659 & ~n34660;
  assign n34662 = ~n34658 & ~n34660;
  assign n34663 = ~n34659 & n34662;
  assign n34664 = ~n34658 & n34661;
  assign n34665 = ~n34657 & n43851;
  assign n34666 = pi62  & ~n34665;
  assign n34667 = pi62  & ~n34666;
  assign n34668 = pi62  & n34665;
  assign n34669 = ~n34665 & ~n34666;
  assign n34670 = ~pi62  & ~n34665;
  assign n34671 = ~n43852 & ~n43853;
  assign n34672 = ~n34420 & ~n34438;
  assign n34673 = pi105  & ~n40814;
  assign n34674 = pi104  & n18285;
  assign n34675 = ~n34673 & ~n34674;
  assign n34676 = n34419 & ~n34675;
  assign n34677 = ~n34419 & n34675;
  assign n34678 = n34419 & ~n34676;
  assign n34679 = n34419 & n34675;
  assign n34680 = ~n34675 & ~n34676;
  assign n34681 = ~n34419 & ~n34675;
  assign n34682 = ~n43854 & ~n43855;
  assign n34683 = ~n34676 & ~n34677;
  assign n34684 = ~n34672 & ~n43856;
  assign n34685 = n34672 & n43856;
  assign n34686 = ~n34672 & ~n34684;
  assign n34687 = ~n34672 & n43856;
  assign n34688 = ~n43856 & ~n34684;
  assign n34689 = n34672 & ~n43856;
  assign n34690 = ~n43857 & ~n43858;
  assign n34691 = ~n34684 & ~n34685;
  assign n34692 = ~n34671 & ~n43859;
  assign n34693 = n34671 & n43859;
  assign n34694 = n34671 & ~n43859;
  assign n34695 = ~n34671 & n43859;
  assign n34696 = ~n34694 & ~n34695;
  assign n34697 = ~n34692 & ~n34693;
  assign n34698 = ~n34656 & ~n43860;
  assign n34699 = n34656 & n43860;
  assign n34700 = ~n34698 & ~n34699;
  assign n34701 = ~n34444 & n34461;
  assign n34702 = ~n34444 & ~n34462;
  assign n34703 = ~n34445 & ~n34701;
  assign n34704 = ~n34700 & n43861;
  assign n34705 = n34700 & ~n43861;
  assign n34706 = ~n34704 & ~n34705;
  assign n34707 = n4312 & n11258;
  assign n34708 = pi112  & n38376;
  assign n34709 = pi114  & n4314;
  assign n34710 = pi113  & n4322;
  assign n34711 = ~n34709 & ~n34710;
  assign n34712 = ~n34708 & ~n34710;
  assign n34713 = ~n34709 & n34712;
  assign n34714 = ~n34708 & n34711;
  assign n34715 = ~n34707 & n43862;
  assign n34716 = pi56  & ~n34715;
  assign n34717 = pi56  & ~n34716;
  assign n34718 = pi56  & n34715;
  assign n34719 = ~n34715 & ~n34716;
  assign n34720 = ~pi56  & ~n34715;
  assign n34721 = ~n43863 & ~n43864;
  assign n34722 = ~n34706 & n34721;
  assign n34723 = n34706 & ~n34721;
  assign n34724 = ~n34722 & ~n34723;
  assign n34725 = ~n34469 & n34485;
  assign n34726 = ~n34469 & ~n34487;
  assign n34727 = ~n34468 & ~n34725;
  assign n34728 = n34724 & ~n43865;
  assign n34729 = ~n34724 & n43865;
  assign n34730 = ~n43865 & ~n34728;
  assign n34731 = n34724 & ~n34728;
  assign n34732 = ~n34730 & ~n34731;
  assign n34733 = ~n34728 & ~n34729;
  assign n34734 = ~n34641 & ~n43866;
  assign n34735 = n34641 & ~n34731;
  assign n34736 = ~n34730 & n34735;
  assign n34737 = n34641 & n43866;
  assign n34738 = ~n34734 & ~n43867;
  assign n34739 = ~n34493 & n34509;
  assign n34740 = ~n34493 & ~n34510;
  assign n34741 = ~n34492 & ~n34739;
  assign n34742 = n34738 & ~n43868;
  assign n34743 = ~n34738 & n43868;
  assign n34744 = ~n43868 & ~n34742;
  assign n34745 = n34738 & ~n34742;
  assign n34746 = ~n34744 & ~n34745;
  assign n34747 = ~n34742 & ~n34743;
  assign n34748 = ~n34626 & ~n43869;
  assign n34749 = n34626 & ~n34745;
  assign n34750 = ~n34744 & n34749;
  assign n34751 = n34626 & n43869;
  assign n34752 = ~n34748 & ~n43870;
  assign n34753 = ~n34611 & n34752;
  assign n34754 = n34611 & ~n34752;
  assign n34755 = ~n34753 & ~n34754;
  assign n34756 = n785 & n14961;
  assign n34757 = pi121  & n37520;
  assign n34758 = pi123  & n787;
  assign n34759 = pi122  & n795;
  assign n34760 = ~n34758 & ~n34759;
  assign n34761 = ~n34757 & ~n34759;
  assign n34762 = ~n34758 & n34761;
  assign n34763 = ~n34757 & n34760;
  assign n34764 = ~n34756 & n43871;
  assign n34765 = pi47  & ~n34764;
  assign n34766 = pi47  & ~n34765;
  assign n34767 = pi47  & n34764;
  assign n34768 = ~n34764 & ~n34765;
  assign n34769 = ~pi47  & ~n34764;
  assign n34770 = ~n43872 & ~n43873;
  assign n34771 = n34755 & ~n34770;
  assign n34772 = ~n34755 & n34770;
  assign n34773 = n34755 & ~n34771;
  assign n34774 = ~n34770 & ~n34771;
  assign n34775 = ~n34773 & ~n34774;
  assign n34776 = ~n34771 & ~n34772;
  assign n34777 = ~n34529 & n34545;
  assign n34778 = ~n34529 & ~n34546;
  assign n34779 = ~n34528 & ~n34777;
  assign n34780 = n43874 & n43875;
  assign n34781 = ~n43874 & ~n43875;
  assign n34782 = ~n34780 & ~n34781;
  assign n34783 = n940 & n15021;
  assign n34784 = pi124  & n37541;
  assign n34785 = pi126  & n953;
  assign n34786 = pi125  & n955;
  assign n34787 = ~n34785 & ~n34786;
  assign n34788 = ~n34784 & ~n34786;
  assign n34789 = ~n34785 & n34788;
  assign n34790 = ~n34784 & n34787;
  assign n34791 = ~n34783 & n43876;
  assign n34792 = pi44  & ~n34791;
  assign n34793 = pi44  & ~n34792;
  assign n34794 = pi44  & n34791;
  assign n34795 = ~n34791 & ~n34792;
  assign n34796 = ~pi44  & ~n34791;
  assign n34797 = ~n43877 & ~n43878;
  assign n34798 = ~n34782 & n34797;
  assign n34799 = n34782 & ~n34797;
  assign n34800 = n34782 & ~n34799;
  assign n34801 = ~n34797 & ~n34799;
  assign n34802 = ~n34800 & ~n34801;
  assign n34803 = ~n34798 & ~n34799;
  assign n34804 = ~n43841 & ~n43879;
  assign n34805 = n43841 & n43879;
  assign n34806 = ~n43841 & n43879;
  assign n34807 = n43841 & ~n43879;
  assign n34808 = ~n34806 & ~n34807;
  assign n34809 = ~n34804 & ~n34805;
  assign n34810 = ~n34591 & ~n43880;
  assign n34811 = n34591 & n43880;
  assign n34812 = ~n34810 & ~n34811;
  assign n34813 = ~n34590 & n34812;
  assign n34814 = n34590 & ~n34812;
  assign po104  = ~n34813 & ~n34814;
  assign n34816 = ~n34810 & ~n34813;
  assign n34817 = ~n34742 & ~n34748;
  assign n34818 = n894 & n15091;
  assign n34819 = pi119  & n37580;
  assign n34820 = pi121  & n896;
  assign n34821 = pi120  & n904;
  assign n34822 = ~n34820 & ~n34821;
  assign n34823 = ~n34819 & ~n34821;
  assign n34824 = ~n34820 & n34823;
  assign n34825 = ~n34819 & n34822;
  assign n34826 = ~n34818 & n43881;
  assign n34827 = pi50  & ~n34826;
  assign n34828 = pi50  & ~n34827;
  assign n34829 = pi50  & n34826;
  assign n34830 = ~n34826 & ~n34827;
  assign n34831 = ~pi50  & ~n34826;
  assign n34832 = ~n43882 & ~n43883;
  assign n34833 = ~n34728 & ~n34734;
  assign n34834 = n1971 & n13057;
  assign n34835 = pi116  & n37864;
  assign n34836 = pi118  & n1973;
  assign n34837 = pi117  & n1981;
  assign n34838 = ~n34836 & ~n34837;
  assign n34839 = ~n34835 & ~n34837;
  assign n34840 = ~n34836 & n34839;
  assign n34841 = ~n34835 & n34838;
  assign n34842 = ~n34834 & n43884;
  assign n34843 = pi53  & ~n34842;
  assign n34844 = pi53  & ~n34843;
  assign n34845 = pi53  & n34842;
  assign n34846 = ~n34842 & ~n34843;
  assign n34847 = ~pi53  & ~n34842;
  assign n34848 = ~n43885 & ~n43886;
  assign n34849 = ~n34705 & ~n34723;
  assign n34850 = n523 & n4312;
  assign n34851 = pi113  & n38376;
  assign n34852 = pi115  & n4314;
  assign n34853 = pi114  & n4322;
  assign n34854 = ~n34852 & ~n34853;
  assign n34855 = ~n34851 & ~n34853;
  assign n34856 = ~n34852 & n34855;
  assign n34857 = ~n34851 & n34854;
  assign n34858 = ~n34850 & n43887;
  assign n34859 = pi56  & ~n34858;
  assign n34860 = pi56  & ~n34859;
  assign n34861 = pi56  & n34858;
  assign n34862 = ~n34858 & ~n34859;
  assign n34863 = ~pi56  & ~n34858;
  assign n34864 = ~n43888 & ~n43889;
  assign n34865 = ~n34692 & ~n34698;
  assign n34866 = ~n34676 & ~n34684;
  assign n34867 = ~pi41  & ~n34419;
  assign n34868 = pi41  & n34419;
  assign n34869 = pi41  & ~n34419;
  assign n34870 = ~pi41  & n34419;
  assign n34871 = ~n34869 & ~n34870;
  assign n34872 = ~n34867 & ~n34868;
  assign n34873 = pi106  & ~n40814;
  assign n34874 = pi105  & n18285;
  assign n34875 = ~n34873 & ~n34874;
  assign n34876 = n43890 & n34875;
  assign n34877 = ~n43890 & ~n34875;
  assign n34878 = ~n34876 & ~n34877;
  assign n34879 = n9701 & n12674;
  assign n34880 = pi107  & n40107;
  assign n34881 = pi109  & n12676;
  assign n34882 = pi108  & n12684;
  assign n34883 = ~n34881 & ~n34882;
  assign n34884 = ~n34880 & ~n34882;
  assign n34885 = ~n34881 & n34884;
  assign n34886 = ~n34880 & n34883;
  assign n34887 = ~n34879 & n43891;
  assign n34888 = pi62  & ~n34887;
  assign n34889 = pi62  & ~n34888;
  assign n34890 = pi62  & n34887;
  assign n34891 = ~n34887 & ~n34888;
  assign n34892 = ~pi62  & ~n34887;
  assign n34893 = ~n43892 & ~n43893;
  assign n34894 = n34878 & ~n34893;
  assign n34895 = ~n34878 & n34893;
  assign n34896 = n34878 & ~n34894;
  assign n34897 = n34878 & n34893;
  assign n34898 = ~n34893 & ~n34894;
  assign n34899 = ~n34878 & ~n34893;
  assign n34900 = ~n43894 & ~n43895;
  assign n34901 = ~n34894 & ~n34895;
  assign n34902 = n34866 & n43896;
  assign n34903 = ~n34866 & ~n43896;
  assign n34904 = ~n34902 & ~n34903;
  assign n34905 = n7882 & n10844;
  assign n34906 = pi110  & n39128;
  assign n34907 = pi112  & n7884;
  assign n34908 = pi111  & n7892;
  assign n34909 = ~n34907 & ~n34908;
  assign n34910 = ~n34906 & ~n34908;
  assign n34911 = ~n34907 & n34910;
  assign n34912 = ~n34906 & n34909;
  assign n34913 = ~n34905 & n43897;
  assign n34914 = pi59  & ~n34913;
  assign n34915 = pi59  & ~n34914;
  assign n34916 = pi59  & n34913;
  assign n34917 = ~n34913 & ~n34914;
  assign n34918 = ~pi59  & ~n34913;
  assign n34919 = ~n43898 & ~n43899;
  assign n34920 = n34904 & ~n34919;
  assign n34921 = ~n34904 & n34919;
  assign n34922 = n34904 & ~n34920;
  assign n34923 = n34904 & n34919;
  assign n34924 = ~n34919 & ~n34920;
  assign n34925 = ~n34904 & ~n34919;
  assign n34926 = ~n43900 & ~n43901;
  assign n34927 = ~n34920 & ~n34921;
  assign n34928 = ~n34865 & ~n43902;
  assign n34929 = n34865 & n43902;
  assign n34930 = ~n34928 & ~n34929;
  assign n34931 = ~n34864 & n34930;
  assign n34932 = n34864 & ~n34930;
  assign n34933 = ~n34864 & ~n34931;
  assign n34934 = ~n34864 & ~n34930;
  assign n34935 = n34930 & ~n34931;
  assign n34936 = n34864 & n34930;
  assign n34937 = ~n43903 & ~n43904;
  assign n34938 = ~n34931 & ~n34932;
  assign n34939 = ~n34849 & ~n43905;
  assign n34940 = n34849 & n43905;
  assign n34941 = ~n34849 & ~n34939;
  assign n34942 = ~n34849 & n43905;
  assign n34943 = ~n43905 & ~n34939;
  assign n34944 = n34849 & ~n43905;
  assign n34945 = ~n43906 & ~n43907;
  assign n34946 = ~n34939 & ~n34940;
  assign n34947 = n34848 & n43908;
  assign n34948 = ~n34848 & ~n43908;
  assign n34949 = ~n34947 & ~n34948;
  assign n34950 = ~n34833 & n34949;
  assign n34951 = n34833 & ~n34949;
  assign n34952 = ~n34950 & ~n34951;
  assign n34953 = n34832 & ~n34952;
  assign n34954 = ~n34832 & n34952;
  assign n34955 = ~n34953 & ~n34954;
  assign n34956 = ~n34817 & n34955;
  assign n34957 = n34817 & ~n34955;
  assign n34958 = ~n34956 & ~n34957;
  assign n34959 = n785 & n15111;
  assign n34960 = pi122  & n37520;
  assign n34961 = pi124  & n787;
  assign n34962 = pi123  & n795;
  assign n34963 = ~n34961 & ~n34962;
  assign n34964 = ~n34960 & ~n34962;
  assign n34965 = ~n34961 & n34964;
  assign n34966 = ~n34960 & n34963;
  assign n34967 = ~n34959 & n43909;
  assign n34968 = pi47  & ~n34967;
  assign n34969 = pi47  & ~n34968;
  assign n34970 = pi47  & n34967;
  assign n34971 = ~n34967 & ~n34968;
  assign n34972 = ~pi47  & ~n34967;
  assign n34973 = ~n43910 & ~n43911;
  assign n34974 = n34958 & ~n34973;
  assign n34975 = ~n34958 & n34973;
  assign n34976 = n34958 & ~n34974;
  assign n34977 = n34958 & n34973;
  assign n34978 = ~n34973 & ~n34974;
  assign n34979 = ~n34958 & ~n34973;
  assign n34980 = ~n43912 & ~n43913;
  assign n34981 = ~n34974 & ~n34975;
  assign n34982 = ~n34753 & n34770;
  assign n34983 = ~n34753 & ~n34771;
  assign n34984 = ~n34754 & ~n34982;
  assign n34985 = n43914 & n43915;
  assign n34986 = ~n43914 & ~n43915;
  assign n34987 = ~n34985 & ~n34986;
  assign n34988 = n940 & n40885;
  assign n34989 = pi125  & n37541;
  assign n34990 = pi127  & n953;
  assign n34991 = pi126  & n955;
  assign n34992 = ~n34990 & ~n34991;
  assign n34993 = ~n34989 & ~n34991;
  assign n34994 = ~n34990 & n34993;
  assign n34995 = ~n34989 & n34992;
  assign n34996 = ~n34988 & n43916;
  assign n34997 = pi44  & ~n34996;
  assign n34998 = pi44  & ~n34997;
  assign n34999 = pi44  & n34996;
  assign n35000 = ~n34996 & ~n34997;
  assign n35001 = ~pi44  & ~n34996;
  assign n35002 = ~n43917 & ~n43918;
  assign n35003 = n34987 & ~n35002;
  assign n35004 = ~n34987 & n35002;
  assign n35005 = n34987 & ~n35003;
  assign n35006 = n34987 & n35002;
  assign n35007 = ~n35002 & ~n35003;
  assign n35008 = ~n34987 & ~n35002;
  assign n35009 = ~n43919 & ~n43920;
  assign n35010 = ~n35003 & ~n35004;
  assign n35011 = ~n34781 & n34797;
  assign n35012 = ~n34781 & ~n34799;
  assign n35013 = ~n34780 & ~n35011;
  assign n35014 = n43921 & n43922;
  assign n35015 = ~n43921 & ~n43922;
  assign n35016 = ~n35014 & ~n35015;
  assign n35017 = ~n34605 & n43879;
  assign n35018 = ~n34605 & ~n34804;
  assign n35019 = ~n34606 & ~n35017;
  assign n35020 = n35016 & ~n43923;
  assign n35021 = ~n35016 & n43923;
  assign n35022 = ~n35020 & ~n35021;
  assign n35023 = ~n34816 & n35022;
  assign n35024 = n34816 & ~n35022;
  assign po105  = ~n35023 & ~n35024;
  assign n35026 = ~n35003 & ~n35015;
  assign n35027 = ~n34974 & ~n34986;
  assign n35028 = n940 & n40891;
  assign n35029 = pi126  & n37541;
  assign n35030 = pi127  & n955;
  assign n35031 = ~n35029 & ~n35030;
  assign n35032 = ~n940 & n35031;
  assign n35033 = ~n40891 & n35031;
  assign n35034 = ~n35032 & ~n35033;
  assign n35035 = ~n35028 & n35031;
  assign n35036 = pi44  & ~n43924;
  assign n35037 = ~pi44  & n43924;
  assign n35038 = ~n35036 & ~n35037;
  assign n35039 = ~n35027 & ~n35038;
  assign n35040 = n35027 & n35038;
  assign n35041 = ~n35039 & ~n35040;
  assign n35042 = n785 & n15068;
  assign n35043 = pi123  & n37520;
  assign n35044 = pi125  & n787;
  assign n35045 = pi124  & n795;
  assign n35046 = ~n35044 & ~n35045;
  assign n35047 = ~n35043 & ~n35045;
  assign n35048 = ~n35044 & n35047;
  assign n35049 = ~n35043 & n35046;
  assign n35050 = ~n35042 & n43925;
  assign n35051 = pi47  & ~n35050;
  assign n35052 = pi47  & ~n35051;
  assign n35053 = pi47  & n35050;
  assign n35054 = ~n35050 & ~n35051;
  assign n35055 = ~pi47  & ~n35050;
  assign n35056 = ~n43926 & ~n43927;
  assign n35057 = ~n34954 & ~n34956;
  assign n35058 = n894 & n15049;
  assign n35059 = pi120  & n37580;
  assign n35060 = pi122  & n896;
  assign n35061 = pi121  & n904;
  assign n35062 = ~n35060 & ~n35061;
  assign n35063 = ~n35059 & ~n35061;
  assign n35064 = ~n35060 & n35063;
  assign n35065 = ~n35059 & n35062;
  assign n35066 = ~n35058 & n43928;
  assign n35067 = pi50  & ~n35066;
  assign n35068 = pi50  & ~n35067;
  assign n35069 = pi50  & n35066;
  assign n35070 = ~n35066 & ~n35067;
  assign n35071 = ~pi50  & ~n35066;
  assign n35072 = ~n43929 & ~n43930;
  assign n35073 = ~n34948 & ~n34950;
  assign n35074 = ~n34931 & ~n34939;
  assign n35075 = ~n34920 & ~n34928;
  assign n35076 = ~n34894 & ~n34903;
  assign n35077 = n9678 & n12674;
  assign n35078 = pi108  & n40107;
  assign n35079 = pi110  & n12676;
  assign n35080 = pi109  & n12684;
  assign n35081 = ~n35079 & ~n35080;
  assign n35082 = ~n35078 & ~n35080;
  assign n35083 = ~n35079 & n35082;
  assign n35084 = ~n35078 & n35081;
  assign n35085 = ~n12674 & n43931;
  assign n35086 = ~n9678 & n43931;
  assign n35087 = ~n35085 & ~n35086;
  assign n35088 = ~n35077 & n43931;
  assign n35089 = pi62  & ~n43932;
  assign n35090 = ~pi62  & n43932;
  assign n35091 = ~n35089 & ~n35090;
  assign n35092 = ~n34867 & ~n34877;
  assign n35093 = pi107  & ~n40814;
  assign n35094 = pi106  & n18285;
  assign n35095 = ~n35093 & ~n35094;
  assign n35096 = ~n35092 & n35095;
  assign n35097 = n35092 & ~n35095;
  assign n35098 = n35095 & ~n35096;
  assign n35099 = n35092 & n35095;
  assign n35100 = ~n35092 & ~n35096;
  assign n35101 = ~n35092 & ~n35095;
  assign n35102 = ~n43933 & ~n43934;
  assign n35103 = ~n35096 & ~n35097;
  assign n35104 = ~n35091 & ~n43935;
  assign n35105 = n35091 & n43935;
  assign n35106 = ~n35104 & ~n35105;
  assign n35107 = ~n35076 & n35106;
  assign n35108 = n35076 & ~n35106;
  assign n35109 = ~n35107 & ~n35108;
  assign n35110 = n7882 & n11276;
  assign n35111 = pi111  & n39128;
  assign n35112 = pi113  & n7884;
  assign n35113 = pi112  & n7892;
  assign n35114 = ~n35112 & ~n35113;
  assign n35115 = ~n35111 & ~n35113;
  assign n35116 = ~n35112 & n35115;
  assign n35117 = ~n35111 & n35114;
  assign n35118 = ~n35110 & n43936;
  assign n35119 = pi59  & ~n35118;
  assign n35120 = pi59  & ~n35119;
  assign n35121 = pi59  & n35118;
  assign n35122 = ~n35118 & ~n35119;
  assign n35123 = ~pi59  & ~n35118;
  assign n35124 = ~n43937 & ~n43938;
  assign n35125 = n35109 & ~n35124;
  assign n35126 = ~n35109 & n35124;
  assign n35127 = n35109 & ~n35125;
  assign n35128 = ~n35124 & ~n35125;
  assign n35129 = ~n35127 & ~n35128;
  assign n35130 = ~n35125 & ~n35126;
  assign n35131 = n35075 & n43939;
  assign n35132 = ~n35075 & ~n43939;
  assign n35133 = ~n35131 & ~n35132;
  assign n35134 = n4312 & n12530;
  assign n35135 = pi114  & n38376;
  assign n35136 = pi116  & n4314;
  assign n35137 = pi115  & n4322;
  assign n35138 = ~n35136 & ~n35137;
  assign n35139 = ~n35135 & ~n35137;
  assign n35140 = ~n35136 & n35139;
  assign n35141 = ~n35135 & n35138;
  assign n35142 = ~n35134 & n43940;
  assign n35143 = pi56  & ~n35142;
  assign n35144 = pi56  & ~n35143;
  assign n35145 = pi56  & n35142;
  assign n35146 = ~n35142 & ~n35143;
  assign n35147 = ~pi56  & ~n35142;
  assign n35148 = ~n43941 & ~n43942;
  assign n35149 = ~n35133 & n35148;
  assign n35150 = n35133 & ~n35148;
  assign n35151 = n35133 & ~n35150;
  assign n35152 = ~n35148 & ~n35150;
  assign n35153 = ~n35151 & ~n35152;
  assign n35154 = ~n35149 & ~n35150;
  assign n35155 = n35074 & n43943;
  assign n35156 = ~n35074 & ~n43943;
  assign n35157 = ~n35155 & ~n35156;
  assign n35158 = n1971 & n13027;
  assign n35159 = pi117  & n37864;
  assign n35160 = pi119  & n1973;
  assign n35161 = pi118  & n1981;
  assign n35162 = ~n35160 & ~n35161;
  assign n35163 = ~n35159 & ~n35161;
  assign n35164 = ~n35160 & n35163;
  assign n35165 = ~n35159 & n35162;
  assign n35166 = ~n35158 & n43944;
  assign n35167 = pi53  & ~n35166;
  assign n35168 = pi53  & ~n35167;
  assign n35169 = pi53  & n35166;
  assign n35170 = ~n35166 & ~n35167;
  assign n35171 = ~pi53  & ~n35166;
  assign n35172 = ~n43945 & ~n43946;
  assign n35173 = n35157 & ~n35172;
  assign n35174 = ~n35157 & n35172;
  assign n35175 = n35157 & ~n35173;
  assign n35176 = ~n35172 & ~n35173;
  assign n35177 = ~n35175 & ~n35176;
  assign n35178 = ~n35173 & ~n35174;
  assign n35179 = ~n35073 & ~n43947;
  assign n35180 = n35073 & n43947;
  assign n35181 = ~n35073 & n43947;
  assign n35182 = n35073 & ~n43947;
  assign n35183 = ~n35181 & ~n35182;
  assign n35184 = ~n35179 & ~n35180;
  assign n35185 = n35072 & n43948;
  assign n35186 = ~n35072 & ~n43948;
  assign n35187 = ~n35185 & ~n35186;
  assign n35188 = ~n35057 & n35187;
  assign n35189 = n35057 & ~n35187;
  assign n35190 = ~n35057 & ~n35188;
  assign n35191 = n35187 & ~n35188;
  assign n35192 = ~n35190 & ~n35191;
  assign n35193 = ~n35188 & ~n35189;
  assign n35194 = n35056 & n43949;
  assign n35195 = ~n35056 & ~n43949;
  assign n35196 = ~n35056 & ~n35195;
  assign n35197 = ~n43949 & ~n35195;
  assign n35198 = ~n35196 & ~n35197;
  assign n35199 = ~n35194 & ~n35195;
  assign n35200 = n35041 & ~n43950;
  assign n35201 = ~n35041 & n43950;
  assign n35202 = n35041 & ~n35200;
  assign n35203 = ~n43950 & ~n35200;
  assign n35204 = ~n35202 & ~n35203;
  assign n35205 = ~n35200 & ~n35201;
  assign n35206 = n35026 & n43951;
  assign n35207 = ~n35026 & ~n43951;
  assign n35208 = ~n35206 & ~n35207;
  assign n35209 = ~n35020 & ~n35023;
  assign n35210 = n35208 & ~n35209;
  assign n35211 = ~n35208 & n35209;
  assign po106  = ~n35210 & ~n35211;
  assign n35213 = ~n35207 & ~n35210;
  assign n35214 = n940 & ~n18675;
  assign n35215 = ~n37541 & ~n35214;
  assign n35216 = pi127  & n37541;
  assign n35217 = n940 & n18680;
  assign n35218 = ~n35216 & ~n35217;
  assign n35219 = pi127  & ~n35215;
  assign n35220 = pi44  & ~n43952;
  assign n35221 = pi44  & ~n35220;
  assign n35222 = pi44  & n43952;
  assign n35223 = ~n43952 & ~n35220;
  assign n35224 = ~pi44  & ~n43952;
  assign n35225 = ~n43953 & ~n43954;
  assign n35226 = n35056 & ~n35188;
  assign n35227 = ~n35188 & ~n35195;
  assign n35228 = ~n35189 & ~n35226;
  assign n35229 = ~n35225 & ~n43955;
  assign n35230 = n35225 & n43955;
  assign n35231 = ~n43955 & ~n35229;
  assign n35232 = ~n35225 & ~n35229;
  assign n35233 = ~n35231 & ~n35232;
  assign n35234 = ~n35229 & ~n35230;
  assign n35235 = n785 & n15021;
  assign n35236 = pi124  & n37520;
  assign n35237 = pi126  & n787;
  assign n35238 = pi125  & n795;
  assign n35239 = ~n35237 & ~n35238;
  assign n35240 = ~n35236 & ~n35238;
  assign n35241 = ~n35237 & n35240;
  assign n35242 = ~n35236 & n35239;
  assign n35243 = ~n35235 & n43957;
  assign n35244 = pi47  & ~n35243;
  assign n35245 = pi47  & ~n35244;
  assign n35246 = pi47  & n35243;
  assign n35247 = ~n35243 & ~n35244;
  assign n35248 = ~pi47  & ~n35243;
  assign n35249 = ~n43958 & ~n43959;
  assign n35250 = ~n35179 & ~n35186;
  assign n35251 = n1971 & n14913;
  assign n35252 = pi118  & n37864;
  assign n35253 = pi120  & n1973;
  assign n35254 = pi119  & n1981;
  assign n35255 = ~n35253 & ~n35254;
  assign n35256 = ~n35252 & ~n35254;
  assign n35257 = ~n35253 & n35256;
  assign n35258 = ~n35252 & n35255;
  assign n35259 = ~n35251 & n43960;
  assign n35260 = pi53  & ~n35259;
  assign n35261 = pi53  & ~n35260;
  assign n35262 = pi53  & n35259;
  assign n35263 = ~n35259 & ~n35260;
  assign n35264 = ~pi53  & ~n35259;
  assign n35265 = ~n43961 & ~n43962;
  assign n35266 = n4312 & n13079;
  assign n35267 = pi115  & n38376;
  assign n35268 = pi117  & n4314;
  assign n35269 = pi116  & n4322;
  assign n35270 = ~n35268 & ~n35269;
  assign n35271 = ~n35267 & ~n35269;
  assign n35272 = ~n35268 & n35271;
  assign n35273 = ~n35267 & n35270;
  assign n35274 = ~n35266 & n43963;
  assign n35275 = pi56  & ~n35274;
  assign n35276 = pi56  & ~n35275;
  assign n35277 = pi56  & n35274;
  assign n35278 = ~n35274 & ~n35275;
  assign n35279 = ~pi56  & ~n35274;
  assign n35280 = ~n43964 & ~n43965;
  assign n35281 = n7882 & n11258;
  assign n35282 = pi112  & n39128;
  assign n35283 = pi114  & n7884;
  assign n35284 = pi113  & n7892;
  assign n35285 = ~n35283 & ~n35284;
  assign n35286 = ~n35282 & ~n35284;
  assign n35287 = ~n35283 & n35286;
  assign n35288 = ~n35282 & n35285;
  assign n35289 = ~n35281 & n43966;
  assign n35290 = pi59  & ~n35289;
  assign n35291 = pi59  & ~n35290;
  assign n35292 = pi59  & n35289;
  assign n35293 = ~n35289 & ~n35290;
  assign n35294 = ~pi59  & ~n35289;
  assign n35295 = ~n43967 & ~n43968;
  assign n35296 = ~n35096 & ~n35104;
  assign n35297 = pi108  & ~n40814;
  assign n35298 = pi107  & n18285;
  assign n35299 = ~n35297 & ~n35298;
  assign n35300 = n35095 & ~n35299;
  assign n35301 = ~n35095 & n35299;
  assign n35302 = ~n35300 & ~n35301;
  assign n35303 = n565 & n12674;
  assign n35304 = pi109  & n40107;
  assign n35305 = pi111  & n12676;
  assign n35306 = pi110  & n12684;
  assign n35307 = ~n35305 & ~n35306;
  assign n35308 = ~n35304 & ~n35306;
  assign n35309 = ~n35305 & n35308;
  assign n35310 = ~n35304 & n35307;
  assign n35311 = ~n12674 & n43969;
  assign n35312 = ~n565 & n43969;
  assign n35313 = ~n35311 & ~n35312;
  assign n35314 = ~n35303 & n43969;
  assign n35315 = pi62  & ~n43970;
  assign n35316 = ~pi62  & n43970;
  assign n35317 = ~n35315 & ~n35316;
  assign n35318 = n35302 & ~n35317;
  assign n35319 = ~n35302 & n35317;
  assign n35320 = ~n35318 & ~n35319;
  assign n35321 = ~n35296 & n35320;
  assign n35322 = n35296 & ~n35320;
  assign n35323 = ~n35296 & ~n35321;
  assign n35324 = n35320 & ~n35321;
  assign n35325 = ~n35323 & ~n35324;
  assign n35326 = ~n35321 & ~n35322;
  assign n35327 = ~n35295 & ~n43971;
  assign n35328 = n35295 & ~n35324;
  assign n35329 = ~n35323 & n35328;
  assign n35330 = n35295 & n43971;
  assign n35331 = ~n35327 & ~n43972;
  assign n35332 = ~n35107 & n35124;
  assign n35333 = ~n35107 & ~n35125;
  assign n35334 = ~n35108 & ~n35332;
  assign n35335 = n35331 & ~n43973;
  assign n35336 = ~n35331 & n43973;
  assign n35337 = ~n43973 & ~n35335;
  assign n35338 = n35331 & ~n35335;
  assign n35339 = ~n35337 & ~n35338;
  assign n35340 = ~n35335 & ~n35336;
  assign n35341 = ~n35280 & ~n43974;
  assign n35342 = n35280 & ~n35338;
  assign n35343 = ~n35337 & n35342;
  assign n35344 = n35280 & n43974;
  assign n35345 = ~n35341 & ~n43975;
  assign n35346 = ~n35132 & n35148;
  assign n35347 = ~n35132 & ~n35150;
  assign n35348 = ~n35131 & ~n35346;
  assign n35349 = n35345 & ~n43976;
  assign n35350 = ~n35345 & n43976;
  assign n35351 = ~n43976 & ~n35349;
  assign n35352 = n35345 & ~n35349;
  assign n35353 = ~n35351 & ~n35352;
  assign n35354 = ~n35349 & ~n35350;
  assign n35355 = ~n35265 & ~n43977;
  assign n35356 = n35265 & ~n35352;
  assign n35357 = ~n35351 & n35356;
  assign n35358 = n35265 & n43977;
  assign n35359 = ~n35355 & ~n43978;
  assign n35360 = ~n35156 & n35172;
  assign n35361 = ~n35156 & ~n35173;
  assign n35362 = ~n35155 & ~n35360;
  assign n35363 = n35359 & ~n43979;
  assign n35364 = ~n35359 & n43979;
  assign n35365 = ~n35363 & ~n35364;
  assign n35366 = n894 & n14961;
  assign n35367 = pi121  & n37580;
  assign n35368 = pi123  & n896;
  assign n35369 = pi122  & n904;
  assign n35370 = ~n35368 & ~n35369;
  assign n35371 = ~n35367 & ~n35369;
  assign n35372 = ~n35368 & n35371;
  assign n35373 = ~n35367 & n35370;
  assign n35374 = ~n35366 & n43980;
  assign n35375 = pi50  & ~n35374;
  assign n35376 = pi50  & ~n35375;
  assign n35377 = pi50  & n35374;
  assign n35378 = ~n35374 & ~n35375;
  assign n35379 = ~pi50  & ~n35374;
  assign n35380 = ~n43981 & ~n43982;
  assign n35381 = n35365 & ~n35380;
  assign n35382 = ~n35365 & n35380;
  assign n35383 = n35365 & ~n35381;
  assign n35384 = ~n35380 & ~n35381;
  assign n35385 = ~n35383 & ~n35384;
  assign n35386 = ~n35381 & ~n35382;
  assign n35387 = ~n35250 & ~n43983;
  assign n35388 = n35250 & n43983;
  assign n35389 = ~n43983 & ~n35387;
  assign n35390 = ~n35250 & ~n35387;
  assign n35391 = ~n35389 & ~n35390;
  assign n35392 = ~n35387 & ~n35388;
  assign n35393 = ~n35249 & ~n43984;
  assign n35394 = ~n43984 & ~n35393;
  assign n35395 = n35249 & ~n43984;
  assign n35396 = ~n35249 & ~n35393;
  assign n35397 = ~n35249 & n43984;
  assign n35398 = n35249 & n43984;
  assign n35399 = ~n35393 & ~n35398;
  assign n35400 = ~n43985 & ~n43986;
  assign n35401 = ~n43956 & n43987;
  assign n35402 = n43956 & ~n43987;
  assign n35403 = ~n43956 & ~n43987;
  assign n35404 = n43956 & n43987;
  assign n35405 = ~n35403 & ~n35404;
  assign n35406 = ~n35401 & ~n35402;
  assign n35407 = ~n35039 & n43950;
  assign n35408 = ~n35039 & ~n35200;
  assign n35409 = ~n35040 & ~n35407;
  assign n35410 = ~n43988 & ~n43989;
  assign n35411 = n43988 & n43989;
  assign n35412 = ~n35410 & ~n35411;
  assign n35413 = ~n35213 & n35412;
  assign n35414 = n35213 & ~n35412;
  assign po107  = ~n35413 & ~n35414;
  assign n35416 = ~n35410 & ~n35413;
  assign n35417 = n894 & n15111;
  assign n35418 = pi122  & n37580;
  assign n35419 = pi124  & n896;
  assign n35420 = pi123  & n904;
  assign n35421 = ~n35419 & ~n35420;
  assign n35422 = ~n35418 & ~n35420;
  assign n35423 = ~n35419 & n35422;
  assign n35424 = ~n35418 & n35421;
  assign n35425 = ~n35417 & n43990;
  assign n35426 = pi50  & ~n35425;
  assign n35427 = pi50  & ~n35426;
  assign n35428 = pi50  & n35425;
  assign n35429 = ~n35425 & ~n35426;
  assign n35430 = ~pi50  & ~n35425;
  assign n35431 = ~n43991 & ~n43992;
  assign n35432 = ~n35349 & ~n35355;
  assign n35433 = n1971 & n15091;
  assign n35434 = pi119  & n37864;
  assign n35435 = pi121  & n1973;
  assign n35436 = pi120  & n1981;
  assign n35437 = ~n35435 & ~n35436;
  assign n35438 = ~n35434 & ~n35436;
  assign n35439 = ~n35435 & n35438;
  assign n35440 = ~n35434 & n35437;
  assign n35441 = ~n35433 & n43993;
  assign n35442 = pi53  & ~n35441;
  assign n35443 = pi53  & ~n35442;
  assign n35444 = pi53  & n35441;
  assign n35445 = ~n35441 & ~n35442;
  assign n35446 = ~pi53  & ~n35441;
  assign n35447 = ~n43994 & ~n43995;
  assign n35448 = ~n35335 & ~n35341;
  assign n35449 = n4312 & n13057;
  assign n35450 = pi116  & n38376;
  assign n35451 = pi118  & n4314;
  assign n35452 = pi117  & n4322;
  assign n35453 = ~n35451 & ~n35452;
  assign n35454 = ~n35450 & ~n35452;
  assign n35455 = ~n35451 & n35454;
  assign n35456 = ~n35450 & n35453;
  assign n35457 = ~n35449 & n43996;
  assign n35458 = pi56  & ~n35457;
  assign n35459 = pi56  & ~n35458;
  assign n35460 = pi56  & n35457;
  assign n35461 = ~n35457 & ~n35458;
  assign n35462 = ~pi56  & ~n35457;
  assign n35463 = ~n43997 & ~n43998;
  assign n35464 = ~n35321 & ~n35327;
  assign n35465 = n523 & n7882;
  assign n35466 = pi113  & n39128;
  assign n35467 = pi115  & n7884;
  assign n35468 = pi114  & n7892;
  assign n35469 = ~n35467 & ~n35468;
  assign n35470 = ~n35466 & ~n35468;
  assign n35471 = ~n35467 & n35470;
  assign n35472 = ~n35466 & n35469;
  assign n35473 = ~n35465 & n43999;
  assign n35474 = pi59  & ~n35473;
  assign n35475 = pi59  & ~n35474;
  assign n35476 = pi59  & n35473;
  assign n35477 = ~n35473 & ~n35474;
  assign n35478 = ~pi59  & ~n35473;
  assign n35479 = ~n44000 & ~n44001;
  assign n35480 = n10844 & n12674;
  assign n35481 = pi110  & n40107;
  assign n35482 = pi112  & n12676;
  assign n35483 = pi111  & n12684;
  assign n35484 = ~n35482 & ~n35483;
  assign n35485 = ~n35481 & ~n35483;
  assign n35486 = ~n35482 & n35485;
  assign n35487 = ~n35481 & n35484;
  assign n35488 = ~n35480 & n44002;
  assign n35489 = pi62  & ~n35488;
  assign n35490 = pi62  & ~n35489;
  assign n35491 = pi62  & n35488;
  assign n35492 = ~n35488 & ~n35489;
  assign n35493 = ~pi62  & ~n35488;
  assign n35494 = ~n44003 & ~n44004;
  assign n35495 = ~n35300 & ~n35318;
  assign n35496 = pi109  & ~n40814;
  assign n35497 = pi108  & n18285;
  assign n35498 = ~n35496 & ~n35497;
  assign n35499 = ~pi44  & ~n35498;
  assign n35500 = pi44  & n35498;
  assign n35501 = ~n35499 & ~n35500;
  assign n35502 = n35095 & ~n35501;
  assign n35503 = ~n35095 & ~n35500;
  assign n35504 = ~n35499 & n35503;
  assign n35505 = ~n35095 & n35501;
  assign n35506 = ~n35095 & ~n44005;
  assign n35507 = n35501 & ~n44005;
  assign n35508 = ~n35506 & ~n35507;
  assign n35509 = ~n35502 & ~n44005;
  assign n35510 = ~n35495 & ~n44006;
  assign n35511 = n35495 & n44006;
  assign n35512 = ~n35495 & ~n35510;
  assign n35513 = ~n44006 & ~n35510;
  assign n35514 = ~n35512 & ~n35513;
  assign n35515 = ~n35510 & ~n35511;
  assign n35516 = ~n35494 & ~n44007;
  assign n35517 = n35494 & n44007;
  assign n35518 = ~n44007 & ~n35516;
  assign n35519 = ~n35494 & ~n35516;
  assign n35520 = ~n35518 & ~n35519;
  assign n35521 = ~n35516 & ~n35517;
  assign n35522 = n35479 & n44008;
  assign n35523 = ~n35479 & ~n44008;
  assign n35524 = ~n35522 & ~n35523;
  assign n35525 = ~n35464 & n35524;
  assign n35526 = n35464 & ~n35524;
  assign n35527 = ~n35525 & ~n35526;
  assign n35528 = n35463 & ~n35527;
  assign n35529 = ~n35463 & n35527;
  assign n35530 = ~n35528 & ~n35529;
  assign n35531 = ~n35448 & n35530;
  assign n35532 = n35448 & ~n35530;
  assign n35533 = ~n35531 & ~n35532;
  assign n35534 = n35447 & ~n35533;
  assign n35535 = ~n35447 & n35533;
  assign n35536 = ~n35534 & ~n35535;
  assign n35537 = ~n35432 & n35536;
  assign n35538 = n35432 & ~n35536;
  assign n35539 = ~n35537 & ~n35538;
  assign n35540 = n35431 & ~n35539;
  assign n35541 = ~n35431 & n35539;
  assign n35542 = ~n35540 & ~n35541;
  assign n35543 = ~n35363 & n35380;
  assign n35544 = ~n35363 & ~n35381;
  assign n35545 = ~n35364 & ~n35543;
  assign n35546 = n35542 & ~n44009;
  assign n35547 = ~n35542 & n44009;
  assign n35548 = ~n35546 & ~n35547;
  assign n35549 = n785 & n40885;
  assign n35550 = pi125  & n37520;
  assign n35551 = pi127  & n787;
  assign n35552 = pi126  & n795;
  assign n35553 = ~n35551 & ~n35552;
  assign n35554 = ~n35550 & ~n35552;
  assign n35555 = ~n35551 & n35554;
  assign n35556 = ~n35550 & n35553;
  assign n35557 = ~n35549 & n44010;
  assign n35558 = pi47  & ~n35557;
  assign n35559 = pi47  & ~n35558;
  assign n35560 = pi47  & n35557;
  assign n35561 = ~n35557 & ~n35558;
  assign n35562 = ~pi47  & ~n35557;
  assign n35563 = ~n44011 & ~n44012;
  assign n35564 = n35548 & ~n35563;
  assign n35565 = ~n35548 & n35563;
  assign n35566 = n35548 & ~n35564;
  assign n35567 = n35548 & n35563;
  assign n35568 = ~n35563 & ~n35564;
  assign n35569 = ~n35548 & ~n35563;
  assign n35570 = ~n44013 & ~n44014;
  assign n35571 = ~n35564 & ~n35565;
  assign n35572 = n35249 & ~n35387;
  assign n35573 = ~n35387 & ~n35393;
  assign n35574 = ~n35388 & ~n35572;
  assign n35575 = n44015 & n44016;
  assign n35576 = ~n44015 & ~n44016;
  assign n35577 = ~n35575 & ~n35576;
  assign n35578 = ~n35229 & ~n43987;
  assign n35579 = ~n35229 & ~n35401;
  assign n35580 = ~n35230 & ~n35578;
  assign n35581 = n35577 & ~n44017;
  assign n35582 = ~n35577 & n44017;
  assign n35583 = ~n35581 & ~n35582;
  assign n35584 = ~n35416 & n35583;
  assign n35585 = n35416 & ~n35583;
  assign po108  = ~n35584 & ~n35585;
  assign n35587 = ~n35564 & ~n35576;
  assign n35588 = ~n35541 & ~n35546;
  assign n35589 = n785 & n40891;
  assign n35590 = pi126  & n37520;
  assign n35591 = pi127  & n795;
  assign n35592 = ~n35590 & ~n35591;
  assign n35593 = ~n785 & n35592;
  assign n35594 = ~n40891 & n35592;
  assign n35595 = ~n35593 & ~n35594;
  assign n35596 = ~n35589 & n35592;
  assign n35597 = pi47  & ~n44018;
  assign n35598 = ~pi47  & n44018;
  assign n35599 = ~n35597 & ~n35598;
  assign n35600 = ~n35588 & ~n35599;
  assign n35601 = n35588 & n35599;
  assign n35602 = ~n35600 & ~n35601;
  assign n35603 = n894 & n15068;
  assign n35604 = pi123  & n37580;
  assign n35605 = pi125  & n896;
  assign n35606 = pi124  & n904;
  assign n35607 = ~n35605 & ~n35606;
  assign n35608 = ~n35604 & ~n35606;
  assign n35609 = ~n35605 & n35608;
  assign n35610 = ~n35604 & n35607;
  assign n35611 = ~n35603 & n44019;
  assign n35612 = pi50  & ~n35611;
  assign n35613 = pi50  & ~n35612;
  assign n35614 = pi50  & n35611;
  assign n35615 = ~n35611 & ~n35612;
  assign n35616 = ~pi50  & ~n35611;
  assign n35617 = ~n44020 & ~n44021;
  assign n35618 = ~n35535 & ~n35537;
  assign n35619 = n1971 & n15049;
  assign n35620 = pi120  & n37864;
  assign n35621 = pi122  & n1973;
  assign n35622 = pi121  & n1981;
  assign n35623 = ~n35621 & ~n35622;
  assign n35624 = ~n35620 & ~n35622;
  assign n35625 = ~n35621 & n35624;
  assign n35626 = ~n35620 & n35623;
  assign n35627 = ~n35619 & n44022;
  assign n35628 = pi53  & ~n35627;
  assign n35629 = pi53  & ~n35628;
  assign n35630 = pi53  & n35627;
  assign n35631 = ~n35627 & ~n35628;
  assign n35632 = ~pi53  & ~n35627;
  assign n35633 = ~n44023 & ~n44024;
  assign n35634 = ~n35529 & ~n35531;
  assign n35635 = ~n35523 & ~n35525;
  assign n35636 = n7882 & n12530;
  assign n35637 = pi114  & n39128;
  assign n35638 = pi116  & n7884;
  assign n35639 = pi115  & n7892;
  assign n35640 = ~n35638 & ~n35639;
  assign n35641 = ~n35637 & ~n35639;
  assign n35642 = ~n35638 & n35641;
  assign n35643 = ~n35637 & n35640;
  assign n35644 = ~n35636 & n44025;
  assign n35645 = pi59  & ~n35644;
  assign n35646 = pi59  & ~n35645;
  assign n35647 = pi59  & n35644;
  assign n35648 = ~n35644 & ~n35645;
  assign n35649 = ~pi59  & ~n35644;
  assign n35650 = ~n44026 & ~n44027;
  assign n35651 = ~n35510 & ~n35516;
  assign n35652 = ~n35499 & ~n44005;
  assign n35653 = ~n35499 & ~n35503;
  assign n35654 = pi110  & ~n40814;
  assign n35655 = pi109  & n18285;
  assign n35656 = ~n35654 & ~n35655;
  assign n35657 = n44028 & ~n35656;
  assign n35658 = ~n44028 & n35656;
  assign n35659 = ~n35657 & ~n35658;
  assign n35660 = n11276 & n12674;
  assign n35661 = pi111  & n40107;
  assign n35662 = pi113  & n12676;
  assign n35663 = pi112  & n12684;
  assign n35664 = ~n35662 & ~n35663;
  assign n35665 = ~n35661 & ~n35663;
  assign n35666 = ~n35662 & n35665;
  assign n35667 = ~n35661 & n35664;
  assign n35668 = ~n35660 & n44029;
  assign n35669 = pi62  & ~n35668;
  assign n35670 = pi62  & ~n35669;
  assign n35671 = pi62  & n35668;
  assign n35672 = ~n35668 & ~n35669;
  assign n35673 = ~pi62  & ~n35668;
  assign n35674 = ~n44030 & ~n44031;
  assign n35675 = ~n35659 & n35674;
  assign n35676 = n35659 & ~n35674;
  assign n35677 = ~n35675 & ~n35676;
  assign n35678 = ~n35651 & n35677;
  assign n35679 = n35651 & ~n35677;
  assign n35680 = ~n35651 & ~n35678;
  assign n35681 = n35677 & ~n35678;
  assign n35682 = ~n35680 & ~n35681;
  assign n35683 = ~n35678 & ~n35679;
  assign n35684 = ~n35650 & ~n44032;
  assign n35685 = n35650 & ~n35681;
  assign n35686 = ~n35680 & n35685;
  assign n35687 = n35650 & n44032;
  assign n35688 = ~n35684 & ~n44033;
  assign n35689 = ~n35635 & n35688;
  assign n35690 = n35635 & ~n35688;
  assign n35691 = ~n35689 & ~n35690;
  assign n35692 = n4312 & n13027;
  assign n35693 = pi117  & n38376;
  assign n35694 = pi119  & n4314;
  assign n35695 = pi118  & n4322;
  assign n35696 = ~n35694 & ~n35695;
  assign n35697 = ~n35693 & ~n35695;
  assign n35698 = ~n35694 & n35697;
  assign n35699 = ~n35693 & n35696;
  assign n35700 = ~n35692 & n44034;
  assign n35701 = pi56  & ~n35700;
  assign n35702 = pi56  & ~n35701;
  assign n35703 = pi56  & n35700;
  assign n35704 = ~n35700 & ~n35701;
  assign n35705 = ~pi56  & ~n35700;
  assign n35706 = ~n44035 & ~n44036;
  assign n35707 = n35691 & ~n35706;
  assign n35708 = ~n35691 & n35706;
  assign n35709 = n35691 & ~n35707;
  assign n35710 = ~n35706 & ~n35707;
  assign n35711 = ~n35709 & ~n35710;
  assign n35712 = ~n35707 & ~n35708;
  assign n35713 = ~n35634 & ~n44037;
  assign n35714 = n35634 & n44037;
  assign n35715 = ~n35634 & n44037;
  assign n35716 = n35634 & ~n44037;
  assign n35717 = ~n35715 & ~n35716;
  assign n35718 = ~n35713 & ~n35714;
  assign n35719 = n35633 & n44038;
  assign n35720 = ~n35633 & ~n44038;
  assign n35721 = ~n35719 & ~n35720;
  assign n35722 = ~n35618 & n35721;
  assign n35723 = n35618 & ~n35721;
  assign n35724 = ~n35618 & ~n35722;
  assign n35725 = n35721 & ~n35722;
  assign n35726 = ~n35724 & ~n35725;
  assign n35727 = ~n35722 & ~n35723;
  assign n35728 = n35617 & n44039;
  assign n35729 = ~n35617 & ~n44039;
  assign n35730 = ~n35617 & ~n35729;
  assign n35731 = ~n44039 & ~n35729;
  assign n35732 = ~n35730 & ~n35731;
  assign n35733 = ~n35728 & ~n35729;
  assign n35734 = n35602 & ~n44040;
  assign n35735 = ~n35602 & n44040;
  assign n35736 = n35602 & ~n35734;
  assign n35737 = ~n44040 & ~n35734;
  assign n35738 = ~n35736 & ~n35737;
  assign n35739 = ~n35734 & ~n35735;
  assign n35740 = n35587 & n44041;
  assign n35741 = ~n35587 & ~n44041;
  assign n35742 = ~n35740 & ~n35741;
  assign n35743 = ~n35581 & ~n35584;
  assign n35744 = n35742 & ~n35743;
  assign n35745 = ~n35742 & n35743;
  assign po109  = ~n35744 & ~n35745;
  assign n35747 = n785 & ~n18675;
  assign n35748 = ~n37520 & ~n35747;
  assign n35749 = pi127  & n37520;
  assign n35750 = ~n785 & ~n35749;
  assign n35751 = ~n18680 & ~n35749;
  assign n35752 = ~n35750 & ~n35751;
  assign n35753 = pi127  & ~n35748;
  assign n35754 = pi47  & ~n44042;
  assign n35755 = ~pi47  & n44042;
  assign n35756 = ~n35754 & ~n35755;
  assign n35757 = n35617 & ~n35722;
  assign n35758 = ~n35722 & ~n35729;
  assign n35759 = ~n35723 & ~n35757;
  assign n35760 = ~n35756 & ~n44043;
  assign n35761 = n35756 & n44043;
  assign n35762 = ~n35760 & ~n35761;
  assign n35763 = n894 & n15021;
  assign n35764 = pi124  & n37580;
  assign n35765 = pi126  & n896;
  assign n35766 = pi125  & n904;
  assign n35767 = ~n35765 & ~n35766;
  assign n35768 = ~n35764 & ~n35766;
  assign n35769 = ~n35765 & n35768;
  assign n35770 = ~n35764 & n35767;
  assign n35771 = ~n35763 & n44044;
  assign n35772 = pi50  & ~n35771;
  assign n35773 = pi50  & ~n35772;
  assign n35774 = pi50  & n35771;
  assign n35775 = ~n35771 & ~n35772;
  assign n35776 = ~pi50  & ~n35771;
  assign n35777 = ~n44045 & ~n44046;
  assign n35778 = ~n35713 & ~n35720;
  assign n35779 = n4312 & n14913;
  assign n35780 = pi118  & n38376;
  assign n35781 = pi120  & n4314;
  assign n35782 = pi119  & n4322;
  assign n35783 = ~n35781 & ~n35782;
  assign n35784 = ~n35780 & ~n35782;
  assign n35785 = ~n35781 & n35784;
  assign n35786 = ~n35780 & n35783;
  assign n35787 = ~n35779 & n44047;
  assign n35788 = pi56  & ~n35787;
  assign n35789 = pi56  & ~n35788;
  assign n35790 = pi56  & n35787;
  assign n35791 = ~n35787 & ~n35788;
  assign n35792 = ~pi56  & ~n35787;
  assign n35793 = ~n44048 & ~n44049;
  assign n35794 = ~n35678 & ~n35684;
  assign n35795 = n7882 & n13079;
  assign n35796 = pi115  & n39128;
  assign n35797 = pi117  & n7884;
  assign n35798 = pi116  & n7892;
  assign n35799 = ~n35797 & ~n35798;
  assign n35800 = ~n35796 & ~n35798;
  assign n35801 = ~n35797 & n35800;
  assign n35802 = ~n35796 & n35799;
  assign n35803 = ~n35795 & n44050;
  assign n35804 = pi59  & ~n35803;
  assign n35805 = pi59  & ~n35804;
  assign n35806 = pi59  & n35803;
  assign n35807 = ~n35803 & ~n35804;
  assign n35808 = ~pi59  & ~n35803;
  assign n35809 = ~n44051 & ~n44052;
  assign n35810 = n11258 & n12674;
  assign n35811 = pi112  & n40107;
  assign n35812 = pi114  & n12676;
  assign n35813 = pi113  & n12684;
  assign n35814 = ~n35812 & ~n35813;
  assign n35815 = ~n35811 & ~n35813;
  assign n35816 = ~n35812 & n35815;
  assign n35817 = ~n35811 & n35814;
  assign n35818 = ~n35810 & n44053;
  assign n35819 = pi62  & ~n35818;
  assign n35820 = pi62  & ~n35819;
  assign n35821 = pi62  & n35818;
  assign n35822 = ~n35818 & ~n35819;
  assign n35823 = ~pi62  & ~n35818;
  assign n35824 = ~n44054 & ~n44055;
  assign n35825 = ~n35658 & ~n35676;
  assign n35826 = pi111  & ~n40814;
  assign n35827 = pi110  & n18285;
  assign n35828 = ~n35826 & ~n35827;
  assign n35829 = n35656 & ~n35828;
  assign n35830 = ~n35656 & n35828;
  assign n35831 = ~n35829 & ~n35830;
  assign n35832 = ~n35825 & ~n35830;
  assign n35833 = ~n35829 & n35832;
  assign n35834 = ~n35825 & n35831;
  assign n35835 = n35825 & ~n35831;
  assign n35836 = ~n35825 & ~n44056;
  assign n35837 = ~n35830 & ~n44056;
  assign n35838 = ~n35829 & n35837;
  assign n35839 = ~n35836 & ~n35838;
  assign n35840 = ~n44056 & ~n35835;
  assign n35841 = ~n35824 & ~n44057;
  assign n35842 = n35824 & n44057;
  assign n35843 = n35824 & ~n44057;
  assign n35844 = ~n35824 & n44057;
  assign n35845 = ~n35843 & ~n35844;
  assign n35846 = ~n35841 & ~n35842;
  assign n35847 = ~n35809 & ~n44058;
  assign n35848 = n35809 & n44058;
  assign n35849 = ~n35847 & ~n35848;
  assign n35850 = ~n35794 & n35849;
  assign n35851 = n35794 & ~n35849;
  assign n35852 = ~n35794 & ~n35850;
  assign n35853 = n35849 & ~n35850;
  assign n35854 = ~n35852 & ~n35853;
  assign n35855 = ~n35850 & ~n35851;
  assign n35856 = ~n35793 & ~n44059;
  assign n35857 = n35793 & ~n35853;
  assign n35858 = ~n35852 & n35857;
  assign n35859 = n35793 & n44059;
  assign n35860 = ~n35856 & ~n44060;
  assign n35861 = ~n35689 & n35706;
  assign n35862 = ~n35689 & ~n35707;
  assign n35863 = ~n35690 & ~n35861;
  assign n35864 = n35860 & ~n44061;
  assign n35865 = ~n35860 & n44061;
  assign n35866 = ~n35864 & ~n35865;
  assign n35867 = n1971 & n14961;
  assign n35868 = pi121  & n37864;
  assign n35869 = pi123  & n1973;
  assign n35870 = pi122  & n1981;
  assign n35871 = ~n35869 & ~n35870;
  assign n35872 = ~n35868 & ~n35870;
  assign n35873 = ~n35869 & n35872;
  assign n35874 = ~n35868 & n35871;
  assign n35875 = ~n35867 & n44062;
  assign n35876 = pi53  & ~n35875;
  assign n35877 = pi53  & ~n35876;
  assign n35878 = pi53  & n35875;
  assign n35879 = ~n35875 & ~n35876;
  assign n35880 = ~pi53  & ~n35875;
  assign n35881 = ~n44063 & ~n44064;
  assign n35882 = n35866 & ~n35881;
  assign n35883 = ~n35866 & n35881;
  assign n35884 = n35866 & ~n35882;
  assign n35885 = ~n35881 & ~n35882;
  assign n35886 = ~n35884 & ~n35885;
  assign n35887 = ~n35882 & ~n35883;
  assign n35888 = ~n35778 & ~n44065;
  assign n35889 = n35778 & n44065;
  assign n35890 = ~n44065 & ~n35888;
  assign n35891 = ~n35778 & ~n35888;
  assign n35892 = ~n35890 & ~n35891;
  assign n35893 = ~n35888 & ~n35889;
  assign n35894 = ~n35777 & ~n44066;
  assign n35895 = ~n44066 & ~n35894;
  assign n35896 = n35777 & ~n44066;
  assign n35897 = ~n35777 & ~n35894;
  assign n35898 = ~n35777 & n44066;
  assign n35899 = n35777 & n44066;
  assign n35900 = ~n35894 & ~n35899;
  assign n35901 = ~n44067 & ~n44068;
  assign n35902 = n35762 & n44069;
  assign n35903 = ~n35762 & ~n44069;
  assign n35904 = n44069 & ~n35902;
  assign n35905 = n35762 & ~n35902;
  assign n35906 = ~n35904 & ~n35905;
  assign n35907 = ~n35902 & ~n35903;
  assign n35908 = ~n35600 & n44040;
  assign n35909 = ~n35600 & ~n35734;
  assign n35910 = ~n35601 & ~n35908;
  assign n35911 = n44070 & n44071;
  assign n35912 = ~n44070 & ~n44071;
  assign n35913 = ~n35911 & ~n35912;
  assign n35914 = ~n35741 & ~n35744;
  assign n35915 = n35913 & ~n35914;
  assign n35916 = ~n35913 & n35914;
  assign po110  = ~n35915 & ~n35916;
  assign n35918 = n1971 & n15111;
  assign n35919 = pi122  & n37864;
  assign n35920 = pi124  & n1973;
  assign n35921 = pi123  & n1981;
  assign n35922 = ~n35920 & ~n35921;
  assign n35923 = ~n35919 & ~n35921;
  assign n35924 = ~n35920 & n35923;
  assign n35925 = ~n35919 & n35922;
  assign n35926 = ~n35918 & n44072;
  assign n35927 = pi53  & ~n35926;
  assign n35928 = pi53  & ~n35927;
  assign n35929 = pi53  & n35926;
  assign n35930 = ~n35926 & ~n35927;
  assign n35931 = ~pi53  & ~n35926;
  assign n35932 = ~n44073 & ~n44074;
  assign n35933 = ~n35850 & ~n35856;
  assign n35934 = n4312 & n15091;
  assign n35935 = pi119  & n38376;
  assign n35936 = pi121  & n4314;
  assign n35937 = pi120  & n4322;
  assign n35938 = ~n35936 & ~n35937;
  assign n35939 = ~n35935 & ~n35937;
  assign n35940 = ~n35936 & n35939;
  assign n35941 = ~n35935 & n35938;
  assign n35942 = ~n35934 & n44075;
  assign n35943 = pi56  & ~n35942;
  assign n35944 = pi56  & ~n35943;
  assign n35945 = pi56  & n35942;
  assign n35946 = ~n35942 & ~n35943;
  assign n35947 = ~pi56  & ~n35942;
  assign n35948 = ~n44076 & ~n44077;
  assign n35949 = ~n35841 & ~n35847;
  assign n35950 = n7882 & n13057;
  assign n35951 = pi116  & n39128;
  assign n35952 = pi118  & n7884;
  assign n35953 = pi117  & n7892;
  assign n35954 = ~n35952 & ~n35953;
  assign n35955 = ~n35951 & ~n35953;
  assign n35956 = ~n35952 & n35955;
  assign n35957 = ~n35951 & n35954;
  assign n35958 = ~n35950 & n44078;
  assign n35959 = pi59  & ~n35958;
  assign n35960 = pi59  & ~n35959;
  assign n35961 = pi59  & n35958;
  assign n35962 = ~n35958 & ~n35959;
  assign n35963 = ~pi59  & ~n35958;
  assign n35964 = ~n44079 & ~n44080;
  assign n35965 = n523 & n12674;
  assign n35966 = pi113  & n40107;
  assign n35967 = pi115  & n12676;
  assign n35968 = pi114  & n12684;
  assign n35969 = ~n35967 & ~n35968;
  assign n35970 = ~n35966 & ~n35968;
  assign n35971 = ~n35967 & n35970;
  assign n35972 = ~n35966 & n35969;
  assign n35973 = ~n35965 & n44081;
  assign n35974 = pi62  & ~n35973;
  assign n35975 = pi62  & ~n35974;
  assign n35976 = pi62  & n35973;
  assign n35977 = ~n35973 & ~n35974;
  assign n35978 = ~pi62  & ~n35973;
  assign n35979 = ~n44082 & ~n44083;
  assign n35980 = ~pi47  & ~n35828;
  assign n35981 = pi47  & n35828;
  assign n35982 = pi47  & ~n35828;
  assign n35983 = ~pi47  & n35828;
  assign n35984 = ~n35982 & ~n35983;
  assign n35985 = ~n35980 & ~n35981;
  assign n35986 = pi112  & ~n40814;
  assign n35987 = pi111  & n18285;
  assign n35988 = ~n35986 & ~n35987;
  assign n35989 = ~n44084 & ~n35988;
  assign n35990 = n44084 & n35988;
  assign n35991 = ~n35989 & ~n35990;
  assign n35992 = ~n35979 & n35991;
  assign n35993 = n35979 & ~n35991;
  assign n35994 = ~n35979 & ~n35992;
  assign n35995 = ~n35979 & ~n35991;
  assign n35996 = n35991 & ~n35992;
  assign n35997 = n35979 & n35991;
  assign n35998 = ~n44085 & ~n44086;
  assign n35999 = ~n35992 & ~n35993;
  assign n36000 = ~n35837 & ~n44087;
  assign n36001 = n35837 & n44087;
  assign n36002 = ~n35837 & ~n36000;
  assign n36003 = ~n35837 & n44087;
  assign n36004 = ~n44087 & ~n36000;
  assign n36005 = n35837 & ~n44087;
  assign n36006 = ~n44088 & ~n44089;
  assign n36007 = ~n36000 & ~n36001;
  assign n36008 = n35964 & n44090;
  assign n36009 = ~n35964 & ~n44090;
  assign n36010 = ~n36008 & ~n36009;
  assign n36011 = ~n35949 & n36010;
  assign n36012 = n35949 & ~n36010;
  assign n36013 = ~n36011 & ~n36012;
  assign n36014 = n35948 & ~n36013;
  assign n36015 = ~n35948 & n36013;
  assign n36016 = ~n36014 & ~n36015;
  assign n36017 = ~n35933 & n36016;
  assign n36018 = n35933 & ~n36016;
  assign n36019 = ~n36017 & ~n36018;
  assign n36020 = n35932 & ~n36019;
  assign n36021 = ~n35932 & n36019;
  assign n36022 = ~n36020 & ~n36021;
  assign n36023 = ~n35864 & n35881;
  assign n36024 = ~n35864 & ~n35882;
  assign n36025 = ~n35865 & ~n36023;
  assign n36026 = n36022 & ~n44091;
  assign n36027 = ~n36022 & n44091;
  assign n36028 = ~n36026 & ~n36027;
  assign n36029 = n894 & n40885;
  assign n36030 = pi125  & n37580;
  assign n36031 = pi127  & n896;
  assign n36032 = pi126  & n904;
  assign n36033 = ~n36031 & ~n36032;
  assign n36034 = ~n36030 & ~n36032;
  assign n36035 = ~n36031 & n36034;
  assign n36036 = ~n36030 & n36033;
  assign n36037 = ~n36029 & n44092;
  assign n36038 = pi50  & ~n36037;
  assign n36039 = pi50  & ~n36038;
  assign n36040 = pi50  & n36037;
  assign n36041 = ~n36037 & ~n36038;
  assign n36042 = ~pi50  & ~n36037;
  assign n36043 = ~n44093 & ~n44094;
  assign n36044 = n36028 & ~n36043;
  assign n36045 = ~n36028 & n36043;
  assign n36046 = n36028 & ~n36044;
  assign n36047 = n36028 & n36043;
  assign n36048 = ~n36043 & ~n36044;
  assign n36049 = ~n36028 & ~n36043;
  assign n36050 = ~n44095 & ~n44096;
  assign n36051 = ~n36044 & ~n36045;
  assign n36052 = n35777 & ~n35888;
  assign n36053 = ~n35888 & ~n35894;
  assign n36054 = ~n35889 & ~n36052;
  assign n36055 = n44097 & n44098;
  assign n36056 = ~n44097 & ~n44098;
  assign n36057 = ~n36055 & ~n36056;
  assign n36058 = ~n35760 & ~n44069;
  assign n36059 = ~n35760 & ~n35902;
  assign n36060 = ~n35761 & ~n36058;
  assign n36061 = ~n36057 & n44099;
  assign n36062 = n36057 & ~n44099;
  assign n36063 = ~n36061 & ~n36062;
  assign n36064 = ~n35912 & ~n35915;
  assign n36065 = n36063 & ~n36064;
  assign n36066 = ~n36063 & n36064;
  assign po111  = ~n36065 & ~n36066;
  assign n36068 = ~n36044 & ~n36056;
  assign n36069 = ~n36021 & ~n36026;
  assign n36070 = n1971 & n15068;
  assign n36071 = pi123  & n37864;
  assign n36072 = pi125  & n1973;
  assign n36073 = pi124  & n1981;
  assign n36074 = ~n36072 & ~n36073;
  assign n36075 = ~n36071 & ~n36073;
  assign n36076 = ~n36072 & n36075;
  assign n36077 = ~n36071 & n36074;
  assign n36078 = ~n36070 & n44100;
  assign n36079 = pi53  & ~n36078;
  assign n36080 = pi53  & ~n36079;
  assign n36081 = pi53  & n36078;
  assign n36082 = ~n36078 & ~n36079;
  assign n36083 = ~pi53  & ~n36078;
  assign n36084 = ~n44101 & ~n44102;
  assign n36085 = ~n36015 & ~n36017;
  assign n36086 = n4312 & n15049;
  assign n36087 = pi120  & n38376;
  assign n36088 = pi122  & n4314;
  assign n36089 = pi121  & n4322;
  assign n36090 = ~n36088 & ~n36089;
  assign n36091 = ~n36087 & ~n36089;
  assign n36092 = ~n36088 & n36091;
  assign n36093 = ~n36087 & n36090;
  assign n36094 = ~n36086 & n44103;
  assign n36095 = pi56  & ~n36094;
  assign n36096 = pi56  & ~n36095;
  assign n36097 = pi56  & n36094;
  assign n36098 = ~n36094 & ~n36095;
  assign n36099 = ~pi56  & ~n36094;
  assign n36100 = ~n44104 & ~n44105;
  assign n36101 = ~n36009 & ~n36011;
  assign n36102 = n7882 & n13027;
  assign n36103 = pi117  & n39128;
  assign n36104 = pi119  & n7884;
  assign n36105 = pi118  & n7892;
  assign n36106 = ~n36104 & ~n36105;
  assign n36107 = ~n36103 & ~n36105;
  assign n36108 = ~n36104 & n36107;
  assign n36109 = ~n36103 & n36106;
  assign n36110 = ~n36102 & n44106;
  assign n36111 = pi59  & ~n36110;
  assign n36112 = pi59  & ~n36111;
  assign n36113 = pi59  & n36110;
  assign n36114 = ~n36110 & ~n36111;
  assign n36115 = ~pi59  & ~n36110;
  assign n36116 = ~n44107 & ~n44108;
  assign n36117 = ~n35992 & ~n36000;
  assign n36118 = ~n35980 & ~n35989;
  assign n36119 = pi113  & ~n40814;
  assign n36120 = pi112  & n18285;
  assign n36121 = ~n36119 & ~n36120;
  assign n36122 = ~n36118 & n36121;
  assign n36123 = n36118 & ~n36121;
  assign n36124 = ~n36122 & ~n36123;
  assign n36125 = n12530 & n12674;
  assign n36126 = pi114  & n40107;
  assign n36127 = pi116  & n12676;
  assign n36128 = pi115  & n12684;
  assign n36129 = ~n36127 & ~n36128;
  assign n36130 = ~n36126 & ~n36128;
  assign n36131 = ~n36127 & n36130;
  assign n36132 = ~n36126 & n36129;
  assign n36133 = ~n12674 & n44109;
  assign n36134 = ~n12530 & n44109;
  assign n36135 = ~n36133 & ~n36134;
  assign n36136 = ~n36125 & n44109;
  assign n36137 = pi62  & ~n44110;
  assign n36138 = ~pi62  & n44110;
  assign n36139 = ~n36137 & ~n36138;
  assign n36140 = n36124 & ~n36139;
  assign n36141 = ~n36124 & n36139;
  assign n36142 = ~n36140 & ~n36141;
  assign n36143 = ~n36117 & n36142;
  assign n36144 = n36117 & ~n36142;
  assign n36145 = ~n36117 & ~n36143;
  assign n36146 = n36142 & ~n36143;
  assign n36147 = ~n36145 & ~n36146;
  assign n36148 = ~n36143 & ~n36144;
  assign n36149 = ~n36116 & ~n44111;
  assign n36150 = n36116 & ~n36146;
  assign n36151 = ~n36145 & n36150;
  assign n36152 = n36116 & n44111;
  assign n36153 = ~n36149 & ~n44112;
  assign n36154 = ~n36101 & n36153;
  assign n36155 = n36101 & ~n36153;
  assign n36156 = ~n36154 & ~n36155;
  assign n36157 = ~n36100 & n36156;
  assign n36158 = n36100 & ~n36156;
  assign n36159 = ~n36157 & ~n36158;
  assign n36160 = ~n36085 & n36159;
  assign n36161 = n36085 & ~n36159;
  assign n36162 = ~n36085 & ~n36160;
  assign n36163 = n36159 & ~n36160;
  assign n36164 = ~n36162 & ~n36163;
  assign n36165 = ~n36160 & ~n36161;
  assign n36166 = ~n36084 & ~n44113;
  assign n36167 = n36084 & ~n36163;
  assign n36168 = ~n36162 & n36167;
  assign n36169 = n36084 & n44113;
  assign n36170 = ~n36166 & ~n44114;
  assign n36171 = ~n36069 & n36170;
  assign n36172 = n36069 & ~n36170;
  assign n36173 = ~n36171 & ~n36172;
  assign n36174 = n894 & n40891;
  assign n36175 = pi126  & n37580;
  assign n36176 = pi127  & n904;
  assign n36177 = ~n36175 & ~n36176;
  assign n36178 = ~n36174 & n36177;
  assign n36179 = pi50  & ~n36178;
  assign n36180 = pi50  & ~n36179;
  assign n36181 = pi50  & n36178;
  assign n36182 = ~n36178 & ~n36179;
  assign n36183 = ~pi50  & ~n36178;
  assign n36184 = ~n44115 & ~n44116;
  assign n36185 = n36173 & ~n36184;
  assign n36186 = ~n36173 & n36184;
  assign n36187 = n36173 & ~n36185;
  assign n36188 = ~n36184 & ~n36185;
  assign n36189 = ~n36187 & ~n36188;
  assign n36190 = ~n36185 & ~n36186;
  assign n36191 = n36068 & n44117;
  assign n36192 = ~n36068 & ~n44117;
  assign n36193 = ~n36191 & ~n36192;
  assign n36194 = ~n36062 & ~n36065;
  assign n36195 = n36193 & ~n36194;
  assign n36196 = ~n36193 & n36194;
  assign po112  = ~n36195 & ~n36196;
  assign n36198 = ~n36160 & ~n36166;
  assign n36199 = n894 & ~n18675;
  assign n36200 = ~n37580 & ~n36199;
  assign n36201 = pi127  & n37580;
  assign n36202 = ~n894 & ~n36201;
  assign n36203 = ~n18680 & ~n36201;
  assign n36204 = ~n36202 & ~n36203;
  assign n36205 = pi127  & ~n36200;
  assign n36206 = pi50  & ~n44118;
  assign n36207 = ~pi50  & n44118;
  assign n36208 = ~n36206 & ~n36207;
  assign n36209 = ~n36198 & ~n36208;
  assign n36210 = n36198 & n36208;
  assign n36211 = ~n36209 & ~n36210;
  assign n36212 = ~n36154 & ~n36157;
  assign n36213 = ~n36143 & ~n36149;
  assign n36214 = ~n36122 & ~n36140;
  assign n36215 = n12674 & n13079;
  assign n36216 = pi115  & n40107;
  assign n36217 = pi117  & n12676;
  assign n36218 = pi116  & n12684;
  assign n36219 = ~n36217 & ~n36218;
  assign n36220 = ~n36216 & ~n36218;
  assign n36221 = ~n36217 & n36220;
  assign n36222 = ~n36216 & n36219;
  assign n36223 = ~n36215 & n44119;
  assign n36224 = pi62  & ~n36223;
  assign n36225 = pi62  & ~n36224;
  assign n36226 = pi62  & n36223;
  assign n36227 = ~n36223 & ~n36224;
  assign n36228 = ~pi62  & ~n36223;
  assign n36229 = ~n44120 & ~n44121;
  assign n36230 = pi114  & ~n40814;
  assign n36231 = pi113  & n18285;
  assign n36232 = ~n36230 & ~n36231;
  assign n36233 = n36121 & ~n36232;
  assign n36234 = ~n36121 & n36232;
  assign n36235 = n36121 & ~n36233;
  assign n36236 = n36121 & n36232;
  assign n36237 = ~n36232 & ~n36233;
  assign n36238 = ~n36121 & ~n36232;
  assign n36239 = ~n44122 & ~n44123;
  assign n36240 = ~n36233 & ~n36234;
  assign n36241 = ~n36229 & ~n44124;
  assign n36242 = n36229 & n44124;
  assign n36243 = ~n36229 & ~n36241;
  assign n36244 = ~n36229 & n44124;
  assign n36245 = ~n44124 & ~n36241;
  assign n36246 = n36229 & ~n44124;
  assign n36247 = ~n44125 & ~n44126;
  assign n36248 = ~n36241 & ~n36242;
  assign n36249 = n36214 & n44127;
  assign n36250 = ~n36214 & ~n44127;
  assign n36251 = ~n36249 & ~n36250;
  assign n36252 = n7882 & n14913;
  assign n36253 = pi118  & n39128;
  assign n36254 = pi120  & n7884;
  assign n36255 = pi119  & n7892;
  assign n36256 = ~n36254 & ~n36255;
  assign n36257 = ~n36253 & ~n36255;
  assign n36258 = ~n36254 & n36257;
  assign n36259 = ~n36253 & n36256;
  assign n36260 = ~n36252 & n44128;
  assign n36261 = pi59  & ~n36260;
  assign n36262 = pi59  & ~n36261;
  assign n36263 = pi59  & n36260;
  assign n36264 = ~n36260 & ~n36261;
  assign n36265 = ~pi59  & ~n36260;
  assign n36266 = ~n44129 & ~n44130;
  assign n36267 = ~n36251 & n36266;
  assign n36268 = n36251 & ~n36266;
  assign n36269 = ~n36267 & ~n36268;
  assign n36270 = ~n36213 & n36269;
  assign n36271 = n36213 & ~n36269;
  assign n36272 = ~n36270 & ~n36271;
  assign n36273 = n4312 & n14961;
  assign n36274 = pi121  & n38376;
  assign n36275 = pi123  & n4314;
  assign n36276 = pi122  & n4322;
  assign n36277 = ~n36275 & ~n36276;
  assign n36278 = ~n36274 & ~n36276;
  assign n36279 = ~n36275 & n36278;
  assign n36280 = ~n36274 & n36277;
  assign n36281 = ~n36273 & n44131;
  assign n36282 = pi56  & ~n36281;
  assign n36283 = pi56  & ~n36282;
  assign n36284 = pi56  & n36281;
  assign n36285 = ~n36281 & ~n36282;
  assign n36286 = ~pi56  & ~n36281;
  assign n36287 = ~n44132 & ~n44133;
  assign n36288 = n36272 & ~n36287;
  assign n36289 = ~n36272 & n36287;
  assign n36290 = n36272 & ~n36288;
  assign n36291 = ~n36287 & ~n36288;
  assign n36292 = ~n36290 & ~n36291;
  assign n36293 = ~n36288 & ~n36289;
  assign n36294 = n36212 & n44134;
  assign n36295 = ~n36212 & ~n44134;
  assign n36296 = ~n36294 & ~n36295;
  assign n36297 = n1971 & n15021;
  assign n36298 = pi124  & n37864;
  assign n36299 = pi126  & n1973;
  assign n36300 = pi125  & n1981;
  assign n36301 = ~n36299 & ~n36300;
  assign n36302 = ~n36298 & ~n36300;
  assign n36303 = ~n36299 & n36302;
  assign n36304 = ~n36298 & n36301;
  assign n36305 = ~n36297 & n44135;
  assign n36306 = pi53  & ~n36305;
  assign n36307 = pi53  & ~n36306;
  assign n36308 = pi53  & n36305;
  assign n36309 = ~n36305 & ~n36306;
  assign n36310 = ~pi53  & ~n36305;
  assign n36311 = ~n44136 & ~n44137;
  assign n36312 = ~n36296 & n36311;
  assign n36313 = n36296 & ~n36311;
  assign n36314 = n36296 & ~n36313;
  assign n36315 = ~n36311 & ~n36313;
  assign n36316 = ~n36314 & ~n36315;
  assign n36317 = ~n36312 & ~n36313;
  assign n36318 = n36211 & ~n44138;
  assign n36319 = ~n36211 & n44138;
  assign n36320 = ~n44138 & ~n36318;
  assign n36321 = n36211 & ~n36318;
  assign n36322 = ~n36320 & ~n36321;
  assign n36323 = ~n36318 & ~n36319;
  assign n36324 = ~n36171 & n36184;
  assign n36325 = ~n36171 & ~n36185;
  assign n36326 = ~n36172 & ~n36324;
  assign n36327 = n44139 & n44140;
  assign n36328 = ~n44139 & ~n44140;
  assign n36329 = ~n36327 & ~n36328;
  assign n36330 = ~n36192 & ~n36195;
  assign n36331 = n36329 & ~n36330;
  assign n36332 = ~n36329 & n36330;
  assign po113  = ~n36331 & ~n36332;
  assign n36334 = n4312 & n15111;
  assign n36335 = pi122  & n38376;
  assign n36336 = pi124  & n4314;
  assign n36337 = pi123  & n4322;
  assign n36338 = ~n36336 & ~n36337;
  assign n36339 = ~n36335 & ~n36337;
  assign n36340 = ~n36336 & n36339;
  assign n36341 = ~n36335 & n36338;
  assign n36342 = ~n36334 & n44141;
  assign n36343 = pi56  & ~n36342;
  assign n36344 = pi56  & ~n36343;
  assign n36345 = pi56  & n36342;
  assign n36346 = ~n36342 & ~n36343;
  assign n36347 = ~pi56  & ~n36342;
  assign n36348 = ~n44142 & ~n44143;
  assign n36349 = ~n36250 & ~n36268;
  assign n36350 = n7882 & n15091;
  assign n36351 = pi119  & n39128;
  assign n36352 = pi121  & n7884;
  assign n36353 = pi120  & n7892;
  assign n36354 = ~n36352 & ~n36353;
  assign n36355 = ~n36351 & ~n36353;
  assign n36356 = ~n36352 & n36355;
  assign n36357 = ~n36351 & n36354;
  assign n36358 = ~n36350 & n44144;
  assign n36359 = pi59  & ~n36358;
  assign n36360 = pi59  & ~n36359;
  assign n36361 = pi59  & n36358;
  assign n36362 = ~n36358 & ~n36359;
  assign n36363 = ~pi59  & ~n36358;
  assign n36364 = ~n44145 & ~n44146;
  assign n36365 = n12674 & n13057;
  assign n36366 = pi116  & n40107;
  assign n36367 = pi118  & n12676;
  assign n36368 = pi117  & n12684;
  assign n36369 = ~n36367 & ~n36368;
  assign n36370 = ~n36366 & ~n36368;
  assign n36371 = ~n36367 & n36370;
  assign n36372 = ~n36366 & n36369;
  assign n36373 = ~n36365 & n44147;
  assign n36374 = pi62  & ~n36373;
  assign n36375 = pi62  & ~n36374;
  assign n36376 = pi62  & n36373;
  assign n36377 = ~n36373 & ~n36374;
  assign n36378 = ~pi62  & ~n36373;
  assign n36379 = ~n44148 & ~n44149;
  assign n36380 = ~n36233 & ~n36241;
  assign n36381 = pi115  & ~n40814;
  assign n36382 = pi114  & n18285;
  assign n36383 = ~n36381 & ~n36382;
  assign n36384 = ~pi50  & ~n36383;
  assign n36385 = pi50  & n36383;
  assign n36386 = ~n36384 & ~n36385;
  assign n36387 = ~n36121 & n36386;
  assign n36388 = n36121 & ~n36386;
  assign n36389 = ~n36387 & ~n36388;
  assign n36390 = ~n36380 & n36389;
  assign n36391 = n36380 & ~n36389;
  assign n36392 = ~n36380 & ~n36390;
  assign n36393 = ~n36380 & ~n36389;
  assign n36394 = n36389 & ~n36390;
  assign n36395 = n36380 & n36389;
  assign n36396 = ~n44150 & ~n44151;
  assign n36397 = ~n36390 & ~n36391;
  assign n36398 = ~n36379 & ~n44152;
  assign n36399 = n36379 & ~n44151;
  assign n36400 = ~n44150 & n36399;
  assign n36401 = n36379 & ~n44150;
  assign n36402 = ~n44151 & n36401;
  assign n36403 = n36379 & n44152;
  assign n36404 = ~n36398 & ~n44153;
  assign n36405 = ~n36364 & n36404;
  assign n36406 = n36364 & ~n36404;
  assign n36407 = ~n36364 & ~n36405;
  assign n36408 = ~n36364 & ~n36404;
  assign n36409 = n36404 & ~n36405;
  assign n36410 = n36364 & n36404;
  assign n36411 = ~n44154 & ~n44155;
  assign n36412 = ~n36405 & ~n36406;
  assign n36413 = ~n36349 & ~n44156;
  assign n36414 = n36349 & ~n44155;
  assign n36415 = ~n44154 & n36414;
  assign n36416 = n36349 & ~n44154;
  assign n36417 = ~n44155 & n36416;
  assign n36418 = n36349 & n44156;
  assign n36419 = ~n36413 & ~n44157;
  assign n36420 = ~n36348 & n36419;
  assign n36421 = n36348 & ~n36419;
  assign n36422 = ~n36420 & ~n36421;
  assign n36423 = ~n36270 & n36287;
  assign n36424 = ~n36270 & ~n36288;
  assign n36425 = ~n36271 & ~n36423;
  assign n36426 = n36422 & ~n44158;
  assign n36427 = ~n36422 & n44158;
  assign n36428 = ~n36426 & ~n36427;
  assign n36429 = n1971 & n40885;
  assign n36430 = pi125  & n37864;
  assign n36431 = pi127  & n1973;
  assign n36432 = pi126  & n1981;
  assign n36433 = ~n36431 & ~n36432;
  assign n36434 = ~n36430 & ~n36432;
  assign n36435 = ~n36431 & n36434;
  assign n36436 = ~n36430 & n36433;
  assign n36437 = ~n36429 & n44159;
  assign n36438 = pi53  & ~n36437;
  assign n36439 = pi53  & ~n36438;
  assign n36440 = pi53  & n36437;
  assign n36441 = ~n36437 & ~n36438;
  assign n36442 = ~pi53  & ~n36437;
  assign n36443 = ~n44160 & ~n44161;
  assign n36444 = n36428 & ~n36443;
  assign n36445 = ~n36428 & n36443;
  assign n36446 = n36428 & ~n36444;
  assign n36447 = n36428 & n36443;
  assign n36448 = ~n36443 & ~n36444;
  assign n36449 = ~n36428 & ~n36443;
  assign n36450 = ~n44162 & ~n44163;
  assign n36451 = ~n36444 & ~n36445;
  assign n36452 = ~n36295 & n36311;
  assign n36453 = ~n36295 & ~n36313;
  assign n36454 = ~n36294 & ~n36452;
  assign n36455 = n44164 & n44165;
  assign n36456 = ~n44164 & ~n44165;
  assign n36457 = ~n36455 & ~n36456;
  assign n36458 = ~n36209 & n44138;
  assign n36459 = ~n36209 & ~n36318;
  assign n36460 = ~n36210 & ~n36458;
  assign n36461 = ~n36457 & n44166;
  assign n36462 = n36457 & ~n44166;
  assign n36463 = ~n36461 & ~n36462;
  assign n36464 = ~n36328 & ~n36331;
  assign n36465 = n36463 & ~n36464;
  assign n36466 = ~n36463 & n36464;
  assign po114  = ~n36465 & ~n36466;
  assign n36468 = ~n36444 & ~n36456;
  assign n36469 = ~n36420 & ~n36426;
  assign n36470 = n4312 & n15068;
  assign n36471 = pi123  & n38376;
  assign n36472 = pi125  & n4314;
  assign n36473 = pi124  & n4322;
  assign n36474 = ~n36472 & ~n36473;
  assign n36475 = ~n36471 & ~n36473;
  assign n36476 = ~n36472 & n36475;
  assign n36477 = ~n36471 & n36474;
  assign n36478 = ~n36470 & n44167;
  assign n36479 = pi56  & ~n36478;
  assign n36480 = pi56  & ~n36479;
  assign n36481 = pi56  & n36478;
  assign n36482 = ~n36478 & ~n36479;
  assign n36483 = ~pi56  & ~n36478;
  assign n36484 = ~n44168 & ~n44169;
  assign n36485 = ~n36405 & ~n36413;
  assign n36486 = n7882 & n15049;
  assign n36487 = pi120  & n39128;
  assign n36488 = pi122  & n7884;
  assign n36489 = pi121  & n7892;
  assign n36490 = ~n36488 & ~n36489;
  assign n36491 = ~n36487 & ~n36489;
  assign n36492 = ~n36488 & n36491;
  assign n36493 = ~n36487 & n36490;
  assign n36494 = ~n36486 & n44170;
  assign n36495 = pi59  & ~n36494;
  assign n36496 = pi59  & ~n36495;
  assign n36497 = pi59  & n36494;
  assign n36498 = ~n36494 & ~n36495;
  assign n36499 = ~pi59  & ~n36494;
  assign n36500 = ~n44171 & ~n44172;
  assign n36501 = ~n36390 & ~n36398;
  assign n36502 = ~n36384 & ~n36387;
  assign n36503 = pi116  & ~n40814;
  assign n36504 = pi115  & n18285;
  assign n36505 = ~n36503 & ~n36504;
  assign n36506 = n36502 & ~n36505;
  assign n36507 = ~n36502 & n36505;
  assign n36508 = ~n36506 & ~n36507;
  assign n36509 = n12674 & n13027;
  assign n36510 = pi117  & n40107;
  assign n36511 = pi119  & n12676;
  assign n36512 = pi118  & n12684;
  assign n36513 = ~n36511 & ~n36512;
  assign n36514 = ~n36510 & ~n36512;
  assign n36515 = ~n36511 & n36514;
  assign n36516 = ~n36510 & n36513;
  assign n36517 = ~n36509 & n44173;
  assign n36518 = pi62  & ~n36517;
  assign n36519 = pi62  & ~n36518;
  assign n36520 = pi62  & n36517;
  assign n36521 = ~n36517 & ~n36518;
  assign n36522 = ~pi62  & ~n36517;
  assign n36523 = ~n44174 & ~n44175;
  assign n36524 = ~n36508 & n36523;
  assign n36525 = n36508 & ~n36523;
  assign n36526 = ~n36524 & ~n36525;
  assign n36527 = ~n36501 & n36526;
  assign n36528 = n36501 & ~n36526;
  assign n36529 = ~n36527 & ~n36528;
  assign n36530 = ~n36500 & n36529;
  assign n36531 = n36500 & ~n36529;
  assign n36532 = ~n36530 & ~n36531;
  assign n36533 = ~n36485 & n36532;
  assign n36534 = n36485 & ~n36532;
  assign n36535 = ~n36485 & ~n36533;
  assign n36536 = n36532 & ~n36533;
  assign n36537 = ~n36535 & ~n36536;
  assign n36538 = ~n36533 & ~n36534;
  assign n36539 = ~n36484 & ~n44176;
  assign n36540 = n36484 & ~n36536;
  assign n36541 = ~n36535 & n36540;
  assign n36542 = n36484 & n44176;
  assign n36543 = ~n36539 & ~n44177;
  assign n36544 = ~n36469 & n36543;
  assign n36545 = n36469 & ~n36543;
  assign n36546 = ~n36544 & ~n36545;
  assign n36547 = n1971 & n40891;
  assign n36548 = pi126  & n37864;
  assign n36549 = pi127  & n1981;
  assign n36550 = ~n36548 & ~n36549;
  assign n36551 = ~n36547 & n36550;
  assign n36552 = pi53  & ~n36551;
  assign n36553 = pi53  & ~n36552;
  assign n36554 = pi53  & n36551;
  assign n36555 = ~n36551 & ~n36552;
  assign n36556 = ~pi53  & ~n36551;
  assign n36557 = ~n44178 & ~n44179;
  assign n36558 = n36546 & ~n36557;
  assign n36559 = ~n36546 & n36557;
  assign n36560 = n36546 & ~n36558;
  assign n36561 = ~n36557 & ~n36558;
  assign n36562 = ~n36560 & ~n36561;
  assign n36563 = ~n36558 & ~n36559;
  assign n36564 = n36468 & n44180;
  assign n36565 = ~n36468 & ~n44180;
  assign n36566 = ~n36564 & ~n36565;
  assign n36567 = ~n36462 & ~n36465;
  assign n36568 = n36566 & ~n36567;
  assign n36569 = ~n36566 & n36567;
  assign po115  = ~n36568 & ~n36569;
  assign n36571 = ~n36533 & ~n36539;
  assign n36572 = n1971 & ~n18675;
  assign n36573 = ~n37864 & ~n36572;
  assign n36574 = pi127  & n37864;
  assign n36575 = ~n1971 & ~n36574;
  assign n36576 = ~n18680 & ~n36574;
  assign n36577 = ~n36575 & ~n36576;
  assign n36578 = pi127  & ~n36573;
  assign n36579 = pi53  & ~n44181;
  assign n36580 = ~pi53  & n44181;
  assign n36581 = ~n36579 & ~n36580;
  assign n36582 = ~n36571 & ~n36581;
  assign n36583 = n36571 & n36581;
  assign n36584 = ~n36582 & ~n36583;
  assign n36585 = ~n36527 & ~n36530;
  assign n36586 = n7882 & n14961;
  assign n36587 = pi121  & n39128;
  assign n36588 = pi123  & n7884;
  assign n36589 = pi122  & n7892;
  assign n36590 = ~n36588 & ~n36589;
  assign n36591 = ~n36587 & ~n36589;
  assign n36592 = ~n36588 & n36591;
  assign n36593 = ~n36587 & n36590;
  assign n36594 = ~n36586 & n44182;
  assign n36595 = pi59  & ~n36594;
  assign n36596 = pi59  & ~n36595;
  assign n36597 = pi59  & n36594;
  assign n36598 = ~n36594 & ~n36595;
  assign n36599 = ~pi59  & ~n36594;
  assign n36600 = ~n44183 & ~n44184;
  assign n36601 = n12674 & n14913;
  assign n36602 = pi118  & n40107;
  assign n36603 = pi120  & n12676;
  assign n36604 = pi119  & n12684;
  assign n36605 = ~n36603 & ~n36604;
  assign n36606 = ~n36602 & ~n36604;
  assign n36607 = ~n36603 & n36606;
  assign n36608 = ~n36602 & n36605;
  assign n36609 = ~n36601 & n44185;
  assign n36610 = pi62  & ~n36609;
  assign n36611 = pi62  & ~n36610;
  assign n36612 = pi62  & n36609;
  assign n36613 = ~n36609 & ~n36610;
  assign n36614 = ~pi62  & ~n36609;
  assign n36615 = ~n44186 & ~n44187;
  assign n36616 = ~n36507 & ~n36525;
  assign n36617 = pi117  & ~n40814;
  assign n36618 = pi116  & n18285;
  assign n36619 = ~n36617 & ~n36618;
  assign n36620 = n36505 & ~n36619;
  assign n36621 = ~n36505 & n36619;
  assign n36622 = ~n36620 & ~n36621;
  assign n36623 = ~n36616 & ~n36621;
  assign n36624 = ~n36620 & n36623;
  assign n36625 = ~n36616 & n36622;
  assign n36626 = n36616 & ~n36622;
  assign n36627 = ~n36616 & ~n44188;
  assign n36628 = ~n36621 & ~n44188;
  assign n36629 = ~n36620 & n36628;
  assign n36630 = ~n36627 & ~n36629;
  assign n36631 = ~n44188 & ~n36626;
  assign n36632 = ~n36615 & ~n44189;
  assign n36633 = n36615 & n44189;
  assign n36634 = n36615 & ~n44189;
  assign n36635 = ~n36615 & n44189;
  assign n36636 = ~n36634 & ~n36635;
  assign n36637 = ~n36632 & ~n36633;
  assign n36638 = ~n36600 & ~n44190;
  assign n36639 = n36600 & n44190;
  assign n36640 = ~n36638 & ~n36639;
  assign n36641 = n36585 & ~n36640;
  assign n36642 = ~n36585 & n36640;
  assign n36643 = ~n36641 & ~n36642;
  assign n36644 = n4312 & n15021;
  assign n36645 = pi124  & n38376;
  assign n36646 = pi126  & n4314;
  assign n36647 = pi125  & n4322;
  assign n36648 = ~n36646 & ~n36647;
  assign n36649 = ~n36645 & ~n36647;
  assign n36650 = ~n36646 & n36649;
  assign n36651 = ~n36645 & n36648;
  assign n36652 = ~n36644 & n44191;
  assign n36653 = pi56  & ~n36652;
  assign n36654 = pi56  & ~n36653;
  assign n36655 = pi56  & n36652;
  assign n36656 = ~n36652 & ~n36653;
  assign n36657 = ~pi56  & ~n36652;
  assign n36658 = ~n44192 & ~n44193;
  assign n36659 = n36643 & ~n36658;
  assign n36660 = ~n36643 & n36658;
  assign n36661 = n36643 & ~n36659;
  assign n36662 = ~n36658 & ~n36659;
  assign n36663 = ~n36661 & ~n36662;
  assign n36664 = ~n36659 & ~n36660;
  assign n36665 = n36584 & ~n44194;
  assign n36666 = ~n36584 & n44194;
  assign n36667 = ~n44194 & ~n36665;
  assign n36668 = n36584 & ~n36665;
  assign n36669 = ~n36667 & ~n36668;
  assign n36670 = ~n36665 & ~n36666;
  assign n36671 = ~n36544 & n36557;
  assign n36672 = ~n36544 & ~n36558;
  assign n36673 = ~n36545 & ~n36671;
  assign n36674 = n44195 & n44196;
  assign n36675 = ~n44195 & ~n44196;
  assign n36676 = ~n36674 & ~n36675;
  assign n36677 = ~n36565 & ~n36568;
  assign n36678 = n36676 & ~n36677;
  assign n36679 = ~n36676 & n36677;
  assign po116  = ~n36678 & ~n36679;
  assign n36681 = ~n36675 & ~n36678;
  assign n36682 = n4312 & n40885;
  assign n36683 = pi125  & n38376;
  assign n36684 = pi127  & n4314;
  assign n36685 = pi126  & n4322;
  assign n36686 = ~n36684 & ~n36685;
  assign n36687 = ~n36683 & ~n36685;
  assign n36688 = ~n36684 & n36687;
  assign n36689 = ~n36683 & n36686;
  assign n36690 = ~n36682 & n44197;
  assign n36691 = pi56  & ~n36690;
  assign n36692 = pi56  & ~n36691;
  assign n36693 = pi56  & n36690;
  assign n36694 = ~n36690 & ~n36691;
  assign n36695 = ~pi56  & ~n36690;
  assign n36696 = ~n44198 & ~n44199;
  assign n36697 = ~n36642 & n36658;
  assign n36698 = ~n36642 & ~n36659;
  assign n36699 = ~n36641 & ~n36697;
  assign n36700 = ~n36696 & ~n44200;
  assign n36701 = n36696 & n44200;
  assign n36702 = ~n44200 & ~n36700;
  assign n36703 = n36696 & ~n44200;
  assign n36704 = ~n36696 & ~n36700;
  assign n36705 = ~n36696 & n44200;
  assign n36706 = ~n44201 & ~n44202;
  assign n36707 = ~n36700 & ~n36701;
  assign n36708 = ~n36632 & ~n36638;
  assign n36709 = n7882 & n15111;
  assign n36710 = pi122  & n39128;
  assign n36711 = pi124  & n7884;
  assign n36712 = pi123  & n7892;
  assign n36713 = ~n36711 & ~n36712;
  assign n36714 = ~n36710 & ~n36712;
  assign n36715 = ~n36711 & n36714;
  assign n36716 = ~n36710 & n36713;
  assign n36717 = ~n36709 & n44204;
  assign n36718 = pi59  & ~n36717;
  assign n36719 = pi59  & ~n36718;
  assign n36720 = pi59  & n36717;
  assign n36721 = ~n36717 & ~n36718;
  assign n36722 = ~pi59  & ~n36717;
  assign n36723 = ~n44205 & ~n44206;
  assign n36724 = ~pi53  & ~n36619;
  assign n36725 = pi53  & n36619;
  assign n36726 = pi53  & ~n36619;
  assign n36727 = ~pi53  & n36619;
  assign n36728 = ~n36726 & ~n36727;
  assign n36729 = ~n36724 & ~n36725;
  assign n36730 = pi118  & ~n40814;
  assign n36731 = pi117  & n18285;
  assign n36732 = ~n36730 & ~n36731;
  assign n36733 = n44207 & n36732;
  assign n36734 = ~n44207 & ~n36732;
  assign n36735 = ~n36733 & ~n36734;
  assign n36736 = n12674 & n15091;
  assign n36737 = pi119  & n40107;
  assign n36738 = pi121  & n12676;
  assign n36739 = pi120  & n12684;
  assign n36740 = ~n36738 & ~n36739;
  assign n36741 = ~n36737 & ~n36739;
  assign n36742 = ~n36738 & n36741;
  assign n36743 = ~n36737 & n36740;
  assign n36744 = ~n36736 & n44208;
  assign n36745 = pi62  & ~n36744;
  assign n36746 = pi62  & ~n36745;
  assign n36747 = pi62  & n36744;
  assign n36748 = ~n36744 & ~n36745;
  assign n36749 = ~pi62  & ~n36744;
  assign n36750 = ~n44209 & ~n44210;
  assign n36751 = n36735 & ~n36750;
  assign n36752 = ~n36735 & n36750;
  assign n36753 = n36735 & ~n36751;
  assign n36754 = n36735 & n36750;
  assign n36755 = ~n36750 & ~n36751;
  assign n36756 = ~n36735 & ~n36750;
  assign n36757 = ~n44211 & ~n44212;
  assign n36758 = ~n36751 & ~n36752;
  assign n36759 = ~n36628 & ~n44213;
  assign n36760 = n36628 & n44213;
  assign n36761 = ~n36759 & ~n36760;
  assign n36762 = ~n36723 & n36761;
  assign n36763 = n36723 & ~n36761;
  assign n36764 = ~n36723 & ~n36762;
  assign n36765 = ~n36723 & ~n36761;
  assign n36766 = n36761 & ~n36762;
  assign n36767 = n36723 & n36761;
  assign n36768 = ~n44214 & ~n44215;
  assign n36769 = ~n36762 & ~n36763;
  assign n36770 = ~n36708 & ~n44216;
  assign n36771 = n36708 & n44216;
  assign n36772 = ~n36708 & ~n36770;
  assign n36773 = ~n36708 & n44216;
  assign n36774 = ~n44216 & ~n36770;
  assign n36775 = n36708 & ~n44216;
  assign n36776 = ~n44217 & ~n44218;
  assign n36777 = ~n36770 & ~n36771;
  assign n36778 = ~n44203 & ~n44219;
  assign n36779 = n44203 & n44219;
  assign n36780 = ~n44203 & n44219;
  assign n36781 = n44203 & ~n44219;
  assign n36782 = ~n36780 & ~n36781;
  assign n36783 = ~n36778 & ~n36779;
  assign n36784 = ~n36582 & n44194;
  assign n36785 = ~n36582 & ~n36665;
  assign n36786 = ~n36583 & ~n36784;
  assign n36787 = ~n44220 & ~n44221;
  assign n36788 = n44220 & n44221;
  assign n36789 = ~n36787 & ~n36788;
  assign n36790 = ~n36681 & n36789;
  assign n36791 = n36681 & ~n36789;
  assign po117  = ~n36790 & ~n36791;
  assign n36793 = ~n36787 & ~n36790;
  assign n36794 = ~n36700 & ~n36778;
  assign n36795 = ~n36762 & ~n36770;
  assign n36796 = n7882 & n15068;
  assign n36797 = pi123  & n39128;
  assign n36798 = pi125  & n7884;
  assign n36799 = pi124  & n7892;
  assign n36800 = ~n36798 & ~n36799;
  assign n36801 = ~n36797 & ~n36799;
  assign n36802 = ~n36798 & n36801;
  assign n36803 = ~n36797 & n36800;
  assign n36804 = ~n36796 & n44222;
  assign n36805 = pi59  & ~n36804;
  assign n36806 = pi59  & ~n36805;
  assign n36807 = pi59  & n36804;
  assign n36808 = ~n36804 & ~n36805;
  assign n36809 = ~pi59  & ~n36804;
  assign n36810 = ~n44223 & ~n44224;
  assign n36811 = ~n36751 & ~n36759;
  assign n36812 = ~n36724 & ~n36734;
  assign n36813 = pi119  & ~n40814;
  assign n36814 = pi118  & n18285;
  assign n36815 = ~n36813 & ~n36814;
  assign n36816 = ~n36812 & n36815;
  assign n36817 = n36812 & ~n36815;
  assign n36818 = ~n36816 & ~n36817;
  assign n36819 = n12674 & n15049;
  assign n36820 = pi120  & n40107;
  assign n36821 = pi122  & n12676;
  assign n36822 = pi121  & n12684;
  assign n36823 = ~n36821 & ~n36822;
  assign n36824 = ~n36820 & ~n36822;
  assign n36825 = ~n36821 & n36824;
  assign n36826 = ~n36820 & n36823;
  assign n36827 = ~n12674 & n44225;
  assign n36828 = ~n15049 & n44225;
  assign n36829 = ~n36827 & ~n36828;
  assign n36830 = ~n36819 & n44225;
  assign n36831 = pi62  & ~n44226;
  assign n36832 = ~pi62  & n44226;
  assign n36833 = ~n36831 & ~n36832;
  assign n36834 = n36818 & ~n36833;
  assign n36835 = ~n36818 & n36833;
  assign n36836 = ~n36834 & ~n36835;
  assign n36837 = ~n36811 & n36836;
  assign n36838 = n36811 & ~n36836;
  assign n36839 = ~n36811 & ~n36837;
  assign n36840 = n36836 & ~n36837;
  assign n36841 = ~n36839 & ~n36840;
  assign n36842 = ~n36837 & ~n36838;
  assign n36843 = ~n36810 & ~n44227;
  assign n36844 = n36810 & ~n36840;
  assign n36845 = ~n36839 & n36844;
  assign n36846 = n36810 & n44227;
  assign n36847 = ~n36843 & ~n44228;
  assign n36848 = ~n36795 & n36847;
  assign n36849 = n36795 & ~n36847;
  assign n36850 = ~n36848 & ~n36849;
  assign n36851 = n4312 & n40891;
  assign n36852 = pi126  & n38376;
  assign n36853 = pi127  & n4322;
  assign n36854 = ~n36852 & ~n36853;
  assign n36855 = ~n36851 & n36854;
  assign n36856 = pi56  & ~n36855;
  assign n36857 = pi56  & ~n36856;
  assign n36858 = pi56  & n36855;
  assign n36859 = ~n36855 & ~n36856;
  assign n36860 = ~pi56  & ~n36855;
  assign n36861 = ~n44229 & ~n44230;
  assign n36862 = n36850 & ~n36861;
  assign n36863 = ~n36850 & n36861;
  assign n36864 = n36850 & ~n36862;
  assign n36865 = ~n36861 & ~n36862;
  assign n36866 = ~n36864 & ~n36865;
  assign n36867 = ~n36862 & ~n36863;
  assign n36868 = ~n36794 & ~n44231;
  assign n36869 = n36794 & n44231;
  assign n36870 = ~n44231 & ~n36868;
  assign n36871 = ~n36794 & ~n36868;
  assign n36872 = ~n36870 & ~n36871;
  assign n36873 = ~n36868 & ~n36869;
  assign n36874 = ~n36793 & ~n44232;
  assign n36875 = n36793 & n44232;
  assign po118  = ~n36874 & ~n36875;
  assign n36877 = ~n36837 & ~n36843;
  assign n36878 = n4312 & ~n18675;
  assign n36879 = ~n38376 & ~n36878;
  assign n36880 = pi127  & n38376;
  assign n36881 = ~n4312 & ~n36880;
  assign n36882 = ~n18680 & ~n36880;
  assign n36883 = ~n36881 & ~n36882;
  assign n36884 = pi127  & ~n36879;
  assign n36885 = pi56  & ~n44233;
  assign n36886 = ~pi56  & n44233;
  assign n36887 = ~n36885 & ~n36886;
  assign n36888 = ~n36877 & ~n36887;
  assign n36889 = n36877 & n36887;
  assign n36890 = ~n36888 & ~n36889;
  assign n36891 = ~n36816 & ~n36834;
  assign n36892 = n12674 & n14961;
  assign n36893 = pi121  & n40107;
  assign n36894 = pi123  & n12676;
  assign n36895 = pi122  & n12684;
  assign n36896 = ~n36894 & ~n36895;
  assign n36897 = ~n36893 & ~n36895;
  assign n36898 = ~n36894 & n36897;
  assign n36899 = ~n36893 & n36896;
  assign n36900 = ~n36892 & n44234;
  assign n36901 = pi62  & ~n36900;
  assign n36902 = pi62  & ~n36901;
  assign n36903 = pi62  & n36900;
  assign n36904 = ~n36900 & ~n36901;
  assign n36905 = ~pi62  & ~n36900;
  assign n36906 = ~n44235 & ~n44236;
  assign n36907 = pi120  & ~n40814;
  assign n36908 = pi119  & n18285;
  assign n36909 = ~n36907 & ~n36908;
  assign n36910 = n36815 & ~n36909;
  assign n36911 = ~n36815 & n36909;
  assign n36912 = n36815 & ~n36910;
  assign n36913 = n36815 & n36909;
  assign n36914 = ~n36909 & ~n36910;
  assign n36915 = ~n36815 & ~n36909;
  assign n36916 = ~n44237 & ~n44238;
  assign n36917 = ~n36910 & ~n36911;
  assign n36918 = ~n36906 & ~n44239;
  assign n36919 = n36906 & n44239;
  assign n36920 = ~n36906 & ~n36918;
  assign n36921 = ~n36906 & n44239;
  assign n36922 = ~n44239 & ~n36918;
  assign n36923 = n36906 & ~n44239;
  assign n36924 = ~n44240 & ~n44241;
  assign n36925 = ~n36918 & ~n36919;
  assign n36926 = n36891 & n44242;
  assign n36927 = ~n36891 & ~n44242;
  assign n36928 = ~n36926 & ~n36927;
  assign n36929 = n7882 & n15021;
  assign n36930 = pi124  & n39128;
  assign n36931 = pi126  & n7884;
  assign n36932 = pi125  & n7892;
  assign n36933 = ~n36931 & ~n36932;
  assign n36934 = ~n36930 & ~n36932;
  assign n36935 = ~n36931 & n36934;
  assign n36936 = ~n36930 & n36933;
  assign n36937 = ~n36929 & n44243;
  assign n36938 = pi59  & ~n36937;
  assign n36939 = pi59  & ~n36938;
  assign n36940 = pi59  & n36937;
  assign n36941 = ~n36937 & ~n36938;
  assign n36942 = ~pi59  & ~n36937;
  assign n36943 = ~n44244 & ~n44245;
  assign n36944 = n36928 & ~n36943;
  assign n36945 = ~n36928 & n36943;
  assign n36946 = n36928 & ~n36944;
  assign n36947 = ~n36943 & ~n36944;
  assign n36948 = ~n36946 & ~n36947;
  assign n36949 = ~n36944 & ~n36945;
  assign n36950 = n36890 & ~n44246;
  assign n36951 = ~n36890 & n44246;
  assign n36952 = ~n44246 & ~n36950;
  assign n36953 = n36890 & ~n36950;
  assign n36954 = ~n36952 & ~n36953;
  assign n36955 = ~n36950 & ~n36951;
  assign n36956 = ~n36848 & n36861;
  assign n36957 = ~n36848 & ~n36862;
  assign n36958 = ~n36849 & ~n36956;
  assign n36959 = n44247 & n44248;
  assign n36960 = ~n44247 & ~n44248;
  assign n36961 = ~n36959 & ~n36960;
  assign n36962 = ~n36868 & ~n36874;
  assign n36963 = n36961 & ~n36962;
  assign n36964 = ~n36961 & n36962;
  assign po119  = ~n36963 & ~n36964;
  assign n36966 = ~n36910 & ~n36918;
  assign n36967 = pi121  & ~n40814;
  assign n36968 = pi120  & n18285;
  assign n36969 = ~n36967 & ~n36968;
  assign n36970 = ~pi56  & ~n36969;
  assign n36971 = pi56  & n36969;
  assign n36972 = ~pi56  & ~n36970;
  assign n36973 = ~pi56  & n36969;
  assign n36974 = ~n36969 & ~n36970;
  assign n36975 = pi56  & ~n36969;
  assign n36976 = ~n44249 & ~n44250;
  assign n36977 = ~n36970 & ~n36971;
  assign n36978 = ~n36815 & ~n44251;
  assign n36979 = n36815 & n44251;
  assign n36980 = ~n36815 & ~n36978;
  assign n36981 = ~n44251 & ~n36978;
  assign n36982 = ~n36980 & ~n36981;
  assign n36983 = ~n36978 & ~n36979;
  assign n36984 = n36966 & n44252;
  assign n36985 = ~n36966 & ~n44252;
  assign n36986 = ~n36984 & ~n36985;
  assign n36987 = n12674 & n15111;
  assign n36988 = pi122  & n40107;
  assign n36989 = pi124  & n12676;
  assign n36990 = pi123  & n12684;
  assign n36991 = ~n36989 & ~n36990;
  assign n36992 = ~n36988 & ~n36990;
  assign n36993 = ~n36989 & n36992;
  assign n36994 = ~n36988 & n36991;
  assign n36995 = ~n36987 & n44253;
  assign n36996 = pi62  & ~n36995;
  assign n36997 = pi62  & ~n36996;
  assign n36998 = pi62  & n36995;
  assign n36999 = ~n36995 & ~n36996;
  assign n37000 = ~pi62  & ~n36995;
  assign n37001 = ~n44254 & ~n44255;
  assign n37002 = n36986 & ~n37001;
  assign n37003 = ~n36986 & n37001;
  assign n37004 = ~n37002 & ~n37003;
  assign n37005 = n7882 & n40885;
  assign n37006 = pi125  & n39128;
  assign n37007 = pi127  & n7884;
  assign n37008 = pi126  & n7892;
  assign n37009 = ~n37007 & ~n37008;
  assign n37010 = ~n37006 & ~n37008;
  assign n37011 = ~n37007 & n37010;
  assign n37012 = ~n37006 & n37009;
  assign n37013 = ~n37005 & n44256;
  assign n37014 = pi59  & ~n37013;
  assign n37015 = pi59  & ~n37014;
  assign n37016 = pi59  & n37013;
  assign n37017 = ~n37013 & ~n37014;
  assign n37018 = ~pi59  & ~n37013;
  assign n37019 = ~n44257 & ~n44258;
  assign n37020 = ~n36927 & n36943;
  assign n37021 = ~n36927 & ~n36944;
  assign n37022 = ~n36926 & ~n37020;
  assign n37023 = ~n37019 & ~n44259;
  assign n37024 = n37019 & n44259;
  assign n37025 = ~n44259 & ~n37023;
  assign n37026 = n37019 & ~n44259;
  assign n37027 = ~n37019 & ~n37023;
  assign n37028 = ~n37019 & n44259;
  assign n37029 = ~n44260 & ~n44261;
  assign n37030 = ~n37023 & ~n37024;
  assign n37031 = ~n37003 & ~n44262;
  assign n37032 = ~n37002 & n37031;
  assign n37033 = n37004 & ~n44262;
  assign n37034 = ~n37004 & n44262;
  assign n37035 = ~n44262 & ~n44263;
  assign n37036 = ~n37003 & ~n44263;
  assign n37037 = ~n37002 & n37036;
  assign n37038 = n37004 & ~n44263;
  assign n37039 = ~n37035 & ~n44264;
  assign n37040 = ~n44263 & ~n37034;
  assign n37041 = ~n36888 & n44246;
  assign n37042 = ~n36888 & ~n36950;
  assign n37043 = ~n36889 & ~n37041;
  assign n37044 = n44265 & n44266;
  assign n37045 = ~n44265 & ~n44266;
  assign n37046 = ~n37044 & ~n37045;
  assign n37047 = ~n36960 & ~n36963;
  assign n37048 = n37046 & ~n37047;
  assign n37049 = ~n37046 & n37047;
  assign po120  = ~n37048 & ~n37049;
  assign n37051 = ~n37023 & ~n44263;
  assign n37052 = ~n36985 & ~n37002;
  assign n37053 = ~n36970 & ~n36978;
  assign n37054 = pi122  & ~n40814;
  assign n37055 = pi121  & n18285;
  assign n37056 = ~n37054 & ~n37055;
  assign n37057 = n37053 & ~n37056;
  assign n37058 = ~n37053 & n37056;
  assign n37059 = ~n37057 & ~n37058;
  assign n37060 = n12674 & n15068;
  assign n37061 = pi123  & n40107;
  assign n37062 = pi125  & n12676;
  assign n37063 = pi124  & n12684;
  assign n37064 = ~n37062 & ~n37063;
  assign n37065 = ~n37061 & ~n37063;
  assign n37066 = ~n37062 & n37065;
  assign n37067 = ~n37061 & n37064;
  assign n37068 = ~n12674 & n44267;
  assign n37069 = ~n15068 & n44267;
  assign n37070 = ~n37068 & ~n37069;
  assign n37071 = ~n37060 & n44267;
  assign n37072 = pi62  & ~n44268;
  assign n37073 = ~pi62  & n44268;
  assign n37074 = ~n37072 & ~n37073;
  assign n37075 = n37059 & ~n37074;
  assign n37076 = ~n37059 & n37074;
  assign n37077 = ~n37075 & ~n37076;
  assign n37078 = ~n37052 & n37077;
  assign n37079 = n37052 & ~n37077;
  assign n37080 = ~n37078 & ~n37079;
  assign n37081 = n7882 & n40891;
  assign n37082 = pi126  & n39128;
  assign n37083 = pi127  & n7892;
  assign n37084 = ~n37082 & ~n37083;
  assign n37085 = ~n37081 & n37084;
  assign n37086 = pi59  & ~n37085;
  assign n37087 = pi59  & ~n37086;
  assign n37088 = pi59  & n37085;
  assign n37089 = ~n37085 & ~n37086;
  assign n37090 = ~pi59  & ~n37085;
  assign n37091 = ~n44269 & ~n44270;
  assign n37092 = n37080 & ~n37091;
  assign n37093 = ~n37080 & n37091;
  assign n37094 = n37080 & ~n37092;
  assign n37095 = ~n37091 & ~n37092;
  assign n37096 = ~n37094 & ~n37095;
  assign n37097 = ~n37092 & ~n37093;
  assign n37098 = n37051 & n44271;
  assign n37099 = ~n37051 & ~n44271;
  assign n37100 = ~n37098 & ~n37099;
  assign n37101 = ~n37045 & ~n37048;
  assign n37102 = n37100 & ~n37101;
  assign n37103 = ~n37100 & n37101;
  assign po121  = ~n37102 & ~n37103;
  assign n37105 = ~n37099 & ~n37102;
  assign n37106 = ~n37058 & ~n37075;
  assign n37107 = pi123  & ~n40814;
  assign n37108 = pi122  & n18285;
  assign n37109 = ~n37107 & ~n37108;
  assign n37110 = n37056 & ~n37109;
  assign n37111 = ~n37056 & n37109;
  assign n37112 = ~n37110 & ~n37111;
  assign n37113 = ~n37106 & ~n37111;
  assign n37114 = ~n37110 & n37113;
  assign n37115 = ~n37106 & n37112;
  assign n37116 = n37106 & ~n37112;
  assign n37117 = ~n37106 & ~n44272;
  assign n37118 = ~n37111 & ~n44272;
  assign n37119 = ~n37110 & n37118;
  assign n37120 = ~n37117 & ~n37119;
  assign n37121 = ~n44272 & ~n37116;
  assign n37122 = n12674 & n15021;
  assign n37123 = pi124  & n40107;
  assign n37124 = pi126  & n12676;
  assign n37125 = pi125  & n12684;
  assign n37126 = ~n37124 & ~n37125;
  assign n37127 = ~n37123 & ~n37125;
  assign n37128 = ~n37124 & n37127;
  assign n37129 = ~n37123 & n37126;
  assign n37130 = ~n37122 & n44274;
  assign n37131 = pi62  & ~n37130;
  assign n37132 = pi62  & ~n37131;
  assign n37133 = pi62  & n37130;
  assign n37134 = ~n37130 & ~n37131;
  assign n37135 = ~pi62  & ~n37130;
  assign n37136 = ~n44275 & ~n44276;
  assign n37137 = n7882 & ~n18675;
  assign n37138 = ~n39128 & ~n37137;
  assign n37139 = pi127  & n39128;
  assign n37140 = n7882 & n18680;
  assign n37141 = ~n37139 & ~n37140;
  assign n37142 = pi127  & ~n37138;
  assign n37143 = pi59  & ~n44277;
  assign n37144 = pi59  & ~n37143;
  assign n37145 = pi59  & n44277;
  assign n37146 = ~n44277 & ~n37143;
  assign n37147 = ~pi59  & ~n44277;
  assign n37148 = ~n44278 & ~n44279;
  assign n37149 = ~n37136 & ~n37148;
  assign n37150 = n37136 & n37148;
  assign n37151 = ~n37136 & ~n37149;
  assign n37152 = ~n37148 & ~n37149;
  assign n37153 = ~n37151 & ~n37152;
  assign n37154 = ~n37149 & ~n37150;
  assign n37155 = ~n44273 & ~n44280;
  assign n37156 = n44273 & n44280;
  assign n37157 = ~n44273 & n44280;
  assign n37158 = n44273 & ~n44280;
  assign n37159 = ~n37157 & ~n37158;
  assign n37160 = ~n37155 & ~n37156;
  assign n37161 = ~n37078 & n37091;
  assign n37162 = ~n37078 & ~n37092;
  assign n37163 = ~n37079 & ~n37161;
  assign n37164 = ~n44281 & ~n44282;
  assign n37165 = n44281 & n44282;
  assign n37166 = ~n44282 & ~n37164;
  assign n37167 = ~n44281 & ~n37164;
  assign n37168 = ~n37166 & ~n37167;
  assign n37169 = ~n37164 & ~n37165;
  assign n37170 = ~n37105 & ~n44283;
  assign n37171 = n37105 & ~n37167;
  assign n37172 = ~n37166 & n37171;
  assign n37173 = n37105 & n44283;
  assign po122  = ~n37170 & ~n44284;
  assign n37175 = ~n37164 & ~n37170;
  assign n37176 = ~n37149 & ~n37155;
  assign n37177 = ~pi59  & ~n37109;
  assign n37178 = pi59  & n37109;
  assign n37179 = pi59  & ~n37109;
  assign n37180 = ~pi59  & n37109;
  assign n37181 = ~n37179 & ~n37180;
  assign n37182 = ~n37177 & ~n37178;
  assign n37183 = pi124  & ~n40814;
  assign n37184 = pi123  & n18285;
  assign n37185 = ~n37183 & ~n37184;
  assign n37186 = n44285 & n37185;
  assign n37187 = ~n44285 & ~n37185;
  assign n37188 = ~n37186 & ~n37187;
  assign n37189 = n12674 & n40885;
  assign n37190 = pi125  & n40107;
  assign n37191 = pi127  & n12676;
  assign n37192 = pi126  & n12684;
  assign n37193 = ~n37191 & ~n37192;
  assign n37194 = ~n37190 & ~n37192;
  assign n37195 = ~n37191 & n37194;
  assign n37196 = ~n37190 & n37193;
  assign n37197 = ~n37189 & n44286;
  assign n37198 = pi62  & ~n37197;
  assign n37199 = pi62  & ~n37198;
  assign n37200 = pi62  & n37197;
  assign n37201 = ~n37197 & ~n37198;
  assign n37202 = ~pi62  & ~n37197;
  assign n37203 = ~n44287 & ~n44288;
  assign n37204 = n37188 & ~n37203;
  assign n37205 = ~n37188 & n37203;
  assign n37206 = n37188 & ~n37204;
  assign n37207 = n37188 & n37203;
  assign n37208 = ~n37203 & ~n37204;
  assign n37209 = ~n37188 & ~n37203;
  assign n37210 = ~n44289 & ~n44290;
  assign n37211 = ~n37204 & ~n37205;
  assign n37212 = ~n37118 & ~n44291;
  assign n37213 = n37118 & n44291;
  assign n37214 = ~n37212 & ~n37213;
  assign n37215 = ~n37176 & n37214;
  assign n37216 = n37176 & ~n37214;
  assign n37217 = ~n37176 & ~n37215;
  assign n37218 = n37214 & ~n37215;
  assign n37219 = ~n37217 & ~n37218;
  assign n37220 = ~n37215 & ~n37216;
  assign n37221 = ~n37175 & ~n44292;
  assign n37222 = n37175 & ~n37218;
  assign n37223 = ~n37217 & n37222;
  assign n37224 = n37175 & n44292;
  assign po123  = ~n37221 & ~n44293;
  assign n37226 = ~n37215 & ~n37221;
  assign n37227 = ~n37204 & ~n37212;
  assign n37228 = ~n37177 & ~n37187;
  assign n37229 = pi125  & ~n40814;
  assign n37230 = pi124  & n18285;
  assign n37231 = ~n37229 & ~n37230;
  assign n37232 = ~n37228 & n37231;
  assign n37233 = n37228 & ~n37231;
  assign n37234 = ~n37232 & ~n37233;
  assign n37235 = n12674 & n40891;
  assign n37236 = pi126  & n40107;
  assign n37237 = pi127  & n12684;
  assign n37238 = ~n37236 & ~n37237;
  assign n37239 = ~n12674 & n37238;
  assign n37240 = ~n40891 & n37238;
  assign n37241 = ~n37239 & ~n37240;
  assign n37242 = ~n37235 & n37238;
  assign n37243 = pi62  & ~n44294;
  assign n37244 = ~pi62  & n44294;
  assign n37245 = ~n37243 & ~n37244;
  assign n37246 = n37234 & ~n37245;
  assign n37247 = ~n37234 & n37245;
  assign n37248 = ~n37246 & ~n37247;
  assign n37249 = ~n37227 & n37248;
  assign n37250 = n37227 & ~n37248;
  assign n37251 = ~n37227 & ~n37249;
  assign n37252 = n37248 & ~n37249;
  assign n37253 = ~n37251 & ~n37252;
  assign n37254 = ~n37249 & ~n37250;
  assign n37255 = ~n37226 & ~n44295;
  assign n37256 = n37226 & ~n37252;
  assign n37257 = ~n37251 & n37256;
  assign n37258 = n37226 & n44295;
  assign po124  = ~n37255 & ~n44296;
  assign n37260 = ~n37249 & ~n37255;
  assign n37261 = ~n37232 & ~n37246;
  assign n37262 = pi126  & ~n40814;
  assign n37263 = pi125  & n18285;
  assign n37264 = ~n37262 & ~n37263;
  assign n37265 = n37231 & ~n37264;
  assign n37266 = ~n37231 & n37264;
  assign n37267 = ~n37265 & ~n37266;
  assign n37268 = n12674 & ~n18675;
  assign n37269 = ~n40107 & ~n37268;
  assign n37270 = pi127  & n40107;
  assign n37271 = ~n12674 & ~n37270;
  assign n37272 = ~n18680 & ~n37270;
  assign n37273 = ~n37271 & ~n37272;
  assign n37274 = pi127  & ~n37269;
  assign n37275 = pi62  & ~n44297;
  assign n37276 = ~pi62  & n44297;
  assign n37277 = ~n37275 & ~n37276;
  assign n37278 = n37267 & ~n37277;
  assign n37279 = ~n37267 & n37277;
  assign n37280 = ~n37278 & ~n37279;
  assign n37281 = ~n37261 & n37280;
  assign n37282 = n37261 & ~n37280;
  assign n37283 = ~n37261 & ~n37281;
  assign n37284 = n37280 & ~n37281;
  assign n37285 = ~n37283 & ~n37284;
  assign n37286 = ~n37281 & ~n37282;
  assign n37287 = ~n37260 & ~n44298;
  assign n37288 = n37260 & ~n37284;
  assign n37289 = ~n37283 & n37288;
  assign n37290 = n37260 & n44298;
  assign po125  = ~n37287 & ~n44299;
  assign n37292 = ~n37281 & ~n37287;
  assign n37293 = ~n37265 & ~n37278;
  assign n37294 = pi63  & pi127 ;
  assign n37295 = pi62  & ~pi127 ;
  assign n37296 = ~n37294 & ~n37295;
  assign n37297 = pi62  & pi126 ;
  assign n37298 = n18285 & n37297;
  assign n37299 = pi126  & n18285;
  assign n37300 = pi127  & ~n40814;
  assign n37301 = ~n44300 & ~n37300;
  assign n37302 = ~pi62  & ~n37301;
  assign n37303 = pi62  & n37301;
  assign n37304 = ~n37302 & ~n37303;
  assign n37305 = ~n37296 & ~n44300;
  assign n37306 = ~n37231 & n44301;
  assign n37307 = n37231 & ~n44301;
  assign n37308 = ~n37306 & ~n37307;
  assign n37309 = ~n37293 & n37308;
  assign n37310 = n37293 & ~n37308;
  assign n37311 = ~n37309 & ~n37310;
  assign n37312 = ~n37292 & n37311;
  assign n37313 = n37292 & ~n37311;
  assign po126  = ~n37312 & ~n37313;
  assign n37315 = ~n37309 & ~n37312;
  assign n37316 = pi127  & n18285;
  assign n37317 = pi62  & n37294;
  assign n37318 = ~n37302 & ~n37306;
  assign n37319 = n44302 & ~n37318;
  assign n37320 = n37306 & n44302;
  assign n37321 = ~n44302 & n37318;
  assign n37322 = ~n37294 & ~n37306;
  assign n37323 = ~n37294 & n37306;
  assign n37324 = pi62  & n37306;
  assign n37325 = n37294 & ~n37324;
  assign n37326 = ~n37323 & ~n37325;
  assign n37327 = ~n44303 & ~n44304;
  assign n37328 = n37315 & n44305;
  assign n37329 = ~n37315 & ~n44305;
  assign n37330 = n37315 & ~n44305;
  assign n37331 = ~n37315 & n44305;
  assign n37332 = ~n37330 & ~n37331;
  assign n37333 = ~n37328 & ~n37329;
  assign n37334 = n18112 & ~n18114;
  assign po62  = ~n18115 & ~n37334;
  assign n37336 = ~n15138 & n18110;
  assign po61  = ~n18111 & ~n37336;
  assign n37338 = n18106 & ~n18108;
  assign po60  = ~n18109 & ~n37338;
  assign n37340 = n18099 & ~n18102;
  assign n37341 = ~n18101 & n37340;
  assign n37342 = n18099 & n40782;
  assign po59  = ~n18105 & ~n44307;
  assign n37344 = n18090 & n40781;
  assign po58  = ~n18098 & ~n37344;
  assign n37346 = n18083 & n40778;
  assign po57  = ~n18089 & ~n37346;
  assign n37348 = n18074 & n40777;
  assign po56  = ~n18082 & ~n37348;
  assign n37350 = n18070 & ~n18072;
  assign po55  = ~n18073 & ~n37350;
  assign n37352 = n18066 & ~n18068;
  assign po54  = ~n18069 & ~n37352;
  assign n37354 = n18059 & n40774;
  assign po53  = ~n18065 & ~n37354;
  assign n37356 = n18055 & ~n18057;
  assign po52  = ~n18058 & ~n37356;
  assign n37358 = n18051 & ~n18053;
  assign po51  = ~n18054 & ~n37358;
  assign n37360 = n18042 & n40773;
  assign po50  = ~n18050 & ~n37360;
  assign n37362 = n18038 & ~n18040;
  assign po49  = ~n18041 & ~n37362;
  assign n37364 = n18034 & ~n18036;
  assign po48  = ~n18037 & ~n37364;
  assign n37366 = n18025 & n40770;
  assign po47  = ~n18033 & ~n37366;
  assign n37368 = n18016 & n40767;
  assign po46  = ~n18024 & ~n37368;
  assign n37370 = n18012 & ~n18014;
  assign po45  = ~n18015 & ~n37370;
  assign n37372 = n18005 & n40764;
  assign po44  = ~n18011 & ~n37372;
  assign n37374 = n17996 & n40763;
  assign po43  = ~n18004 & ~n37374;
  assign n37376 = n17987 & n40760;
  assign po42  = ~n17995 & ~n37376;
  assign n37378 = n17983 & ~n17985;
  assign po41  = ~n17986 & ~n37378;
  assign n37380 = n17979 & ~n17981;
  assign po40  = ~n17982 & ~n37380;
  assign n37382 = n17970 & n40757;
  assign po39  = ~n17978 & ~n37382;
  assign n37384 = n17961 & n40754;
  assign po38  = ~n17969 & ~n37384;
  assign n37386 = n17957 & ~n17959;
  assign po37  = ~n17960 & ~n37386;
  assign n37388 = n17948 & n40751;
  assign po36  = ~n17956 & ~n37388;
  assign n37390 = n17941 & n40748;
  assign po35  = ~n17947 & ~n37390;
  assign n37392 = n17934 & n40747;
  assign po34  = ~n17940 & ~n37392;
  assign n37394 = n17930 & ~n17932;
  assign po33  = ~n17933 & ~n37394;
  assign n37396 = n17923 & n40746;
  assign po32  = ~n17929 & ~n37396;
  assign n37398 = n17914 & n40745;
  assign po31  = ~n17922 & ~n37398;
  assign n37400 = n17905 & n40742;
  assign po30  = ~n17913 & ~n37400;
  assign n37402 = n17898 & n40739;
  assign po29  = ~n17904 & ~n37402;
  assign n37404 = n17894 & ~n17896;
  assign po28  = ~n17897 & ~n37404;
  assign n37406 = n17890 & ~n17892;
  assign po27  = ~n17893 & ~n37406;
  assign n37408 = n17886 & ~n17888;
  assign po26  = ~n17889 & ~n37408;
  assign n37410 = n17882 & ~n17884;
  assign po25  = ~n17885 & ~n37410;
  assign n37412 = n17873 & n40738;
  assign po24  = ~n17881 & ~n37412;
  assign n37414 = n17864 & n40735;
  assign po23  = ~n17872 & ~n37414;
  assign n37416 = n17860 & ~n17862;
  assign po22  = ~n17863 & ~n37416;
  assign n37418 = n17851 & n40732;
  assign po21  = ~n17859 & ~n37418;
  assign n37420 = n17844 & n40729;
  assign po20  = ~n17850 & ~n37420;
  assign n37422 = n17835 & n40728;
  assign po19  = ~n17843 & ~n37422;
  assign n37424 = n17826 & n40725;
  assign po18  = ~n17834 & ~n37424;
  assign n37426 = n17817 & n40722;
  assign po17  = ~n17825 & ~n37426;
  assign n37428 = n17810 & n40719;
  assign po16  = ~n17816 & ~n37428;
  assign n37430 = n17801 & ~n40717;
  assign n37431 = ~n40716 & n37430;
  assign n37432 = n17801 & n40718;
  assign po15  = ~n17809 & ~n44308;
  assign n37434 = n17794 & n40715;
  assign po14  = ~n17800 & ~n37434;
  assign n37436 = n17787 & n40714;
  assign po13  = ~n17793 & ~n37436;
  assign n37438 = n17778 & n40713;
  assign po12  = ~n17786 & ~n37438;
  assign n37440 = n17771 & n40710;
  assign po11  = ~n17777 & ~n37440;
  assign n37442 = n17767 & ~n17769;
  assign po10  = ~n17770 & ~n37442;
  assign n37444 = n17758 & n40709;
  assign po9  = ~n17766 & ~n37444;
  assign n37446 = n17749 & n40706;
  assign po8  = ~n17757 & ~n37446;
  assign n37448 = n17745 & ~n17747;
  assign po7  = ~n17748 & ~n37448;
  assign n37450 = n17741 & ~n17743;
  assign po6  = ~n17744 & ~n37450;
  assign n37452 = n17732 & n40703;
  assign po5  = ~n17740 & ~n37452;
  assign n37454 = n17723 & n40700;
  assign po4  = ~n17731 & ~n37454;
  assign n37456 = ~n17691 & ~n40697;
  assign po3  = ~n17722 & ~n37456;
  assign n37458 = pi2  & ~n40694;
  assign n37459 = n40696 & ~n37458;
  assign n37460 = ~n40696 & n37458;
  assign n37461 = ~n40694 & n17719;
  assign n37462 = ~n40697 & ~n37461;
  assign n37463 = ~n37459 & ~n37460;
  assign n37464 = pi2  & po0 ;
  assign n37465 = ~n17696 & n37464;
  assign n37466 = n17696 & ~n37464;
  assign n37467 = ~n17698 & n17702;
  assign n37468 = ~n40694 & ~n37467;
  assign n37469 = ~n37465 & ~n37466;
  assign n37470 = n261 | ~n262;
  assign n37471 = n267 | ~n268;
  assign n37472 = n323 | n324;
  assign n37473 = n326 | ~n327;
  assign n37474 = n529 | ~n530;
  assign n37475 = n533 | n534;
  assign n37476 = n542 | n543;
  assign n37477 = n546 | n547;
  assign n37478 = n548 | n549;
  assign n37479 = n555 | ~n556;
  assign n37480 = n561 | ~n562;
  assign n37481 = n571 | ~n572;
  assign n37482 = n575 | n576;
  assign n37483 = n584 | n585;
  assign n37484 = n588 | n589;
  assign n37485 = n590 | n591;
  assign n37486 = n599 | ~n600;
  assign n37487 = n605 | ~n606;
  assign n37488 = n613 | ~n614;
  assign n37489 = n617 | n618;
  assign n37490 = n626 | n627;
  assign n37491 = n630 | n631;
  assign n37492 = n632 | n633;
  assign n37493 = n641 | ~n642;
  assign n37494 = n647 | ~n648;
  assign n37495 = n655 | ~n656;
  assign n37496 = n659 | n660;
  assign n37497 = n668 | n669;
  assign n37498 = n672 | n673;
  assign n37499 = n674 | n675;
  assign n37500 = n683 | ~n684;
  assign n37501 = n689 | ~n690;
  assign n37502 = n697 | ~n698;
  assign n37503 = n701 | n702;
  assign n37504 = n710 | n711;
  assign n37505 = n714 | n715;
  assign n37506 = n716 | n717;
  assign n37507 = n725 | ~n726;
  assign n37508 = n731 | ~n732;
  assign n37509 = n739 | ~n740;
  assign n37510 = n743 | n744;
  assign n37511 = n752 | n753;
  assign n37512 = n756 | n757;
  assign n37513 = n758 | n759;
  assign n37514 = n765 | ~n766;
  assign n37515 = n771 | ~n772;
  assign n37516 = n777 | ~n778;
  assign n37517 = n783 | ~n784;
  assign n37518 = n793 | ~n794;
  assign n37519 = n805 | n806;
  assign n37520 = n809 | n810;
  assign n37521 = ~n825 | n817 | ~n824;
  assign n37522 = n822 | n823;
  assign n37523 = n833 | n830 | n832;
  assign n37524 = n835 | n836;
  assign n37525 = n837 | n838;
  assign n37526 = n843 | n844;
  assign n37527 = n854 | n855;
  assign n37528 = n858 | n859;
  assign n37529 = n860 | n861;
  assign n37530 = n866 | ~n867;
  assign n37531 = n878 | n879;
  assign n37532 = n882 | n883;
  assign n37533 = n884 | n885;
  assign n37534 = n892 | ~n893;
  assign n37535 = n902 | ~n903;
  assign n37536 = n915 | n916;
  assign n37537 = n918 | n919;
  assign n37538 = n932 | ~n933;
  assign n37539 = n938 | ~n939;
  assign n37540 = n946 | ~n947;
  assign n37541 = n950 | n951;
  assign n37542 = n959 | n960;
  assign n37543 = n963 | n964;
  assign n37544 = n965 | n966;
  assign n37545 = n979 | n980;
  assign n37546 = n983 | n984;
  assign n37547 = n985 | n986;
  assign n37548 = n997 | n998;
  assign n37549 = n1001 | n1002;
  assign n37550 = n1003 | n1004;
  assign n37551 = n1010 | n1011;
  assign n37552 = n1019 | n1020;
  assign n37553 = n1023 | n1024;
  assign n37554 = n1025 | n1026;
  assign n37555 = n1032 | n1033;
  assign n37556 = n1046 | n1047;
  assign n37557 = n1057 | n1054 | n1056;
  assign n37558 = n1059 | n1060;
  assign n37559 = n1061 | n1062;
  assign n37560 = n1067 | n1068;
  assign n37561 = n1076 | n1077;
  assign n37562 = n1080 | n1081;
  assign n37563 = n1082 | n1083;
  assign n37564 = n1088 | ~n1089;
  assign n37565 = n1097 | n1098;
  assign n37566 = n1099 | n1100;
  assign n37567 = n1101 | ~n1102;
  assign n37568 = n1106 | n1107;
  assign n37569 = n1108 | n1109;
  assign n37570 = n1110 | ~n1111;
  assign n37571 = n1115 | n1116;
  assign n37572 = n1117 | n1118;
  assign n37573 = n1119 | ~n1120;
  assign n37574 = n1131 | n1132;
  assign n37575 = n1135 | n1136;
  assign n37576 = n1137 | n1138;
  assign n37577 = n1147 | n1148;
  assign n37578 = n1151 | n1152;
  assign n37579 = n1153 | n1154;
  assign n37580 = n1159 | n1160;
  assign n37581 = n1170 | n1167 | n1169;
  assign n37582 = n1172 | n1173;
  assign n37583 = n1174 | n1175;
  assign n37584 = n1182 | n1183;
  assign n37585 = n1185 | n1186;
  assign n37586 = n1189 | n1190;
  assign n37587 = n1191 | n1192;
  assign n37588 = n1193 | ~n1194;
  assign n37589 = n1200 | n1201;
  assign n37590 = n1202 | n1203;
  assign n37591 = n1204 | ~n1205;
  assign n37592 = n1208 | n1209;
  assign n37593 = n1210 | n1211;
  assign n37594 = n1212 | ~n1213;
  assign n37595 = n1225 | n1226;
  assign n37596 = n1229 | n1230;
  assign n37597 = n1231 | n1232;
  assign n37598 = n1245 | n1246;
  assign n37599 = n1249 | n1250;
  assign n37600 = n1251 | n1252;
  assign n37601 = n1261 | n1262;
  assign n37602 = n1265 | n1266;
  assign n37603 = n1267 | n1268;
  assign n37604 = n1281 | n1282;
  assign n37605 = n1285 | n1286;
  assign n37606 = n1287 | n1288;
  assign n37607 = n1299 | n1300;
  assign n37608 = n1303 | n1304;
  assign n37609 = n1305 | n1306;
  assign n37610 = n1315 | n1316;
  assign n37611 = n1319 | n1320;
  assign n37612 = n1321 | n1322;
  assign n37613 = n1328 | n1329;
  assign n37614 = n1337 | n1338;
  assign n37615 = n1341 | n1342;
  assign n37616 = n1343 | n1344;
  assign n37617 = n1350 | n1351;
  assign n37618 = n1364 | n1365;
  assign n37619 = n1375 | n1372 | n1374;
  assign n37620 = n1377 | n1378;
  assign n37621 = n1379 | n1380;
  assign n37622 = n1385 | n1386;
  assign n37623 = n1394 | n1395;
  assign n37624 = n1398 | n1399;
  assign n37625 = n1400 | n1401;
  assign n37626 = n1406 | ~n1407;
  assign n37627 = n1415 | n1416;
  assign n37628 = n1417 | n1418;
  assign n37629 = n1419 | ~n1420;
  assign n37630 = n1424 | n1425;
  assign n37631 = n1426 | n1427;
  assign n37632 = n1428 | ~n1429;
  assign n37633 = n1433 | n1434;
  assign n37634 = n1435 | n1436;
  assign n37635 = n1437 | ~n1438;
  assign n37636 = n1442 | n1443;
  assign n37637 = n1444 | n1445;
  assign n37638 = n1446 | ~n1447;
  assign n37639 = n1457 | n1458;
  assign n37640 = n1472 | n1473;
  assign n37641 = n1476 | n1477;
  assign n37642 = n1478 | n1479;
  assign n37643 = n1489 | n1490;
  assign n37644 = n1493 | n1494;
  assign n37645 = n1495 | n1496;
  assign n37646 = n1502 | ~n1503;
  assign n37647 = n1509 | ~n1510;
  assign n37648 = n1520 | n1521;
  assign n37649 = n1524 | n1525;
  assign n37650 = n1526 | n1527;
  assign n37651 = n1531 | n1532;
  assign n37652 = n1533 | n1534;
  assign n37653 = n1535 | ~n1536;
  assign n37654 = n1546 | n1547;
  assign n37655 = n1550 | n1551;
  assign n37656 = n1552 | n1553;
  assign n37657 = n1563 | n1564;
  assign n37658 = n1565 | n1566;
  assign n37659 = n1567 | ~n1568;
  assign n37660 = n1571 | n1572;
  assign n37661 = n1585 | n1586;
  assign n37662 = n1589 | n1590;
  assign n37663 = n1591 | n1592;
  assign n37664 = n1603 | n1604;
  assign n37665 = n1607 | n1608;
  assign n37666 = n1609 | n1610;
  assign n37667 = n1615 | ~n1616;
  assign n37668 = n1624 | n1625;
  assign n37669 = n1628 | n1629;
  assign n37670 = n1630 | n1631;
  assign n37671 = n1642 | n1643;
  assign n37672 = n1646 | n1647;
  assign n37673 = n1648 | n1649;
  assign n37674 = n1652 | n1653;
  assign n37675 = n1654 | n1655;
  assign n37676 = n1656 | ~n1657;
  assign n37677 = n1667 | n1668;
  assign n37678 = n1671 | n1672;
  assign n37679 = n1673 | n1674;
  assign n37680 = n1685 | n1686;
  assign n37681 = n1689 | n1690;
  assign n37682 = n1691 | n1692;
  assign n37683 = n1701 | n1702;
  assign n37684 = n1705 | n1706;
  assign n37685 = n1707 | n1708;
  assign n37686 = n1721 | n1722;
  assign n37687 = n1725 | n1726;
  assign n37688 = n1727 | n1728;
  assign n37689 = n1739 | n1740;
  assign n37690 = n1743 | n1744;
  assign n37691 = n1745 | n1746;
  assign n37692 = n1755 | n1756;
  assign n37693 = n1759 | n1760;
  assign n37694 = n1761 | n1762;
  assign n37695 = n1768 | n1769;
  assign n37696 = n1777 | n1778;
  assign n37697 = n1781 | n1782;
  assign n37698 = n1783 | n1784;
  assign n37699 = n1790 | n1791;
  assign n37700 = n1804 | n1805;
  assign n37701 = n1815 | n1812 | n1814;
  assign n37702 = n1817 | n1818;
  assign n37703 = n1819 | n1820;
  assign n37704 = n1825 | n1826;
  assign n37705 = n1834 | n1835;
  assign n37706 = n1838 | n1839;
  assign n37707 = n1840 | n1841;
  assign n37708 = n1846 | ~n1847;
  assign n37709 = n1855 | n1856;
  assign n37710 = n1857 | n1858;
  assign n37711 = n1859 | ~n1860;
  assign n37712 = n1864 | n1865;
  assign n37713 = n1866 | n1867;
  assign n37714 = n1868 | ~n1869;
  assign n37715 = n1873 | n1874;
  assign n37716 = n1875 | n1876;
  assign n37717 = n1877 | ~n1878;
  assign n37718 = n1882 | n1883;
  assign n37719 = n1884 | n1885;
  assign n37720 = n1886 | ~n1887;
  assign n37721 = n1897 | n1898;
  assign n37722 = n1905 | n1906;
  assign n37723 = n1907 | n1908;
  assign n37724 = n1909 | ~n1910;
  assign n37725 = n1918 | n1919;
  assign n37726 = n1920 | n1921;
  assign n37727 = n1922 | ~n1923;
  assign n37728 = n1937 | n1938;
  assign n37729 = n1941 | n1942;
  assign n37730 = n1943 | n1944;
  assign n37731 = n1955 | n1956;
  assign n37732 = n1959 | n1960;
  assign n37733 = n1961 | n1962;
  assign n37734 = n1969 | ~n1970;
  assign n37735 = n1979 | ~n1980;
  assign n37736 = n1992 | n1993;
  assign n37737 = n1995 | n1996;
  assign n37738 = n2009 | n2010;
  assign n37739 = n2013 | n2014;
  assign n37740 = n2015 | n2016;
  assign n37741 = n2020 | n2021;
  assign n37742 = n2022 | n2023;
  assign n37743 = n2024 | ~n2025;
  assign n37744 = n2035 | n2036;
  assign n37745 = n2039 | n2040;
  assign n37746 = n2041 | n2042;
  assign n37747 = n2048 | n2049;
  assign n37748 = n2054 | ~n2055;
  assign n37749 = n2070 | n2071;
  assign n37750 = n2074 | n2075;
  assign n37751 = n2076 | n2077;
  assign n37752 = n2081 | n2082;
  assign n37753 = n2083 | n2084;
  assign n37754 = n2085 | ~n2086;
  assign n37755 = n2096 | ~n2097;
  assign n37756 = n2102 | ~n2103;
  assign n37757 = n2110 | ~n2111;
  assign n37758 = n2114 | n2115;
  assign n37759 = n2123 | n2124;
  assign n37760 = n2127 | n2128;
  assign n37761 = n2129 | n2130;
  assign n37762 = n2141 | n2142;
  assign n37763 = n2145 | n2146;
  assign n37764 = n2147 | n2148;
  assign n37765 = n2161 | n2162;
  assign n37766 = n2165 | n2166;
  assign n37767 = n2167 | n2168;
  assign n37768 = n2181 | n2182;
  assign n37769 = n2185 | n2186;
  assign n37770 = n2187 | n2188;
  assign n37771 = n2197 | n2198;
  assign n37772 = n2201 | n2202;
  assign n37773 = n2203 | n2204;
  assign n37774 = n2207 | n2208;
  assign n37775 = n2219 | n2220;
  assign n37776 = n2223 | n2224;
  assign n37777 = n2225 | n2226;
  assign n37778 = n2235 | n2236;
  assign n37779 = n2239 | n2240;
  assign n37780 = n2241 | n2242;
  assign n37781 = n2247 | ~n2248;
  assign n37782 = n2256 | n2257;
  assign n37783 = n2260 | n2261;
  assign n37784 = n2262 | n2263;
  assign n37785 = n2274 | n2275;
  assign n37786 = n2278 | n2279;
  assign n37787 = n2280 | n2281;
  assign n37788 = n2284 | n2285;
  assign n37789 = n2286 | n2287;
  assign n37790 = n2288 | ~n2289;
  assign n37791 = n2299 | n2300;
  assign n37792 = n2303 | n2304;
  assign n37793 = n2305 | n2306;
  assign n37794 = n2317 | n2318;
  assign n37795 = n2321 | n2322;
  assign n37796 = n2323 | n2324;
  assign n37797 = n2333 | n2334;
  assign n37798 = n2337 | n2338;
  assign n37799 = n2339 | n2340;
  assign n37800 = n2353 | n2354;
  assign n37801 = n2357 | n2358;
  assign n37802 = n2359 | n2360;
  assign n37803 = n2371 | n2372;
  assign n37804 = n2375 | n2376;
  assign n37805 = n2377 | n2378;
  assign n37806 = n2387 | n2388;
  assign n37807 = n2391 | n2392;
  assign n37808 = n2393 | n2394;
  assign n37809 = n2400 | n2401;
  assign n37810 = n2409 | n2410;
  assign n37811 = n2413 | n2414;
  assign n37812 = n2415 | n2416;
  assign n37813 = n2422 | n2423;
  assign n37814 = n2436 | n2437;
  assign n37815 = n2447 | n2444 | n2446;
  assign n37816 = n2449 | n2450;
  assign n37817 = n2451 | n2452;
  assign n37818 = n2457 | n2458;
  assign n37819 = n2466 | n2467;
  assign n37820 = n2470 | n2471;
  assign n37821 = n2472 | n2473;
  assign n37822 = n2478 | ~n2479;
  assign n37823 = n2487 | n2488;
  assign n37824 = n2489 | n2490;
  assign n37825 = n2491 | ~n2492;
  assign n37826 = n2496 | n2497;
  assign n37827 = n2498 | n2499;
  assign n37828 = n2500 | ~n2501;
  assign n37829 = n2505 | n2506;
  assign n37830 = n2507 | n2508;
  assign n37831 = n2509 | ~n2510;
  assign n37832 = n2514 | n2515;
  assign n37833 = n2516 | n2517;
  assign n37834 = n2518 | ~n2519;
  assign n37835 = n2529 | n2530;
  assign n37836 = n2537 | n2538;
  assign n37837 = n2539 | n2540;
  assign n37838 = n2541 | ~n2542;
  assign n37839 = n2550 | n2551;
  assign n37840 = n2552 | n2553;
  assign n37841 = n2554 | ~n2555;
  assign n37842 = n2563 | n2564;
  assign n37843 = n2565 | n2566;
  assign n37844 = n2567 | ~n2568;
  assign n37845 = n2572 | n2573;
  assign n37846 = n2574 | n2575;
  assign n37847 = n2576 | ~n2577;
  assign n37848 = n2587 | n2588;
  assign n37849 = n2598 | n2599;
  assign n37850 = n2602 | n2603;
  assign n37851 = n2604 | n2605;
  assign n37852 = n2614 | n2615;
  assign n37853 = n2618 | n2619;
  assign n37854 = n2620 | n2621;
  assign n37855 = n2630 | n2631;
  assign n37856 = n2634 | n2635;
  assign n37857 = n2636 | n2637;
  assign n37858 = n2646 | n2647;
  assign n37859 = n2650 | n2651;
  assign n37860 = n2652 | n2653;
  assign n37861 = n2662 | n2663;
  assign n37862 = n2666 | n2667;
  assign n37863 = n2668 | n2669;
  assign n37864 = n2674 | n2675;
  assign n37865 = n2685 | n2682 | n2684;
  assign n37866 = n2687 | n2688;
  assign n37867 = n2689 | n2690;
  assign n37868 = n2697 | n2698;
  assign n37869 = n2700 | n2701;
  assign n37870 = n2706 | n2707;
  assign n37871 = n2712 | ~n2713;
  assign n37872 = n2732 | n2733;
  assign n37873 = n2736 | n2737;
  assign n37874 = n2738 | n2739;
  assign n37875 = n2743 | n2744;
  assign n37876 = n2745 | n2746;
  assign n37877 = n2747 | ~n2748;
  assign n37878 = n2754 | n2755;
  assign n37879 = n2756 | n2757;
  assign n37880 = n2758 | ~n2759;
  assign n37881 = n2762 | n2763;
  assign n37882 = n2764 | n2765;
  assign n37883 = n2766 | ~n2767;
  assign n37884 = n2772 | ~n2773;
  assign n37885 = n2786 | n2787;
  assign n37886 = n2790 | n2791;
  assign n37887 = n2792 | n2793;
  assign n37888 = n2798 | ~n2799;
  assign n37889 = n2811 | n2812;
  assign n37890 = n2815 | n2816;
  assign n37891 = n2817 | n2818;
  assign n37892 = n2827 | n2828;
  assign n37893 = n2831 | n2832;
  assign n37894 = n2833 | n2834;
  assign n37895 = n2837 | n2838;
  assign n37896 = n2839 | n2840;
  assign n37897 = n2841 | ~n2842;
  assign n37898 = n2852 | n2853;
  assign n37899 = n2856 | n2857;
  assign n37900 = n2858 | n2859;
  assign n37901 = n2870 | n2871;
  assign n37902 = n2874 | n2875;
  assign n37903 = n2876 | n2877;
  assign n37904 = n2886 | n2887;
  assign n37905 = n2890 | n2891;
  assign n37906 = n2892 | n2893;
  assign n37907 = n2906 | n2907;
  assign n37908 = n2910 | n2911;
  assign n37909 = n2912 | n2913;
  assign n37910 = n2922 | n2923;
  assign n37911 = n2926 | n2927;
  assign n37912 = n2928 | n2929;
  assign n37913 = n2934 | ~n2935;
  assign n37914 = n2943 | n2944;
  assign n37915 = n2947 | n2948;
  assign n37916 = n2949 | n2950;
  assign n37917 = n2961 | n2962;
  assign n37918 = n2965 | n2966;
  assign n37919 = n2967 | n2968;
  assign n37920 = n2973 | ~n2974;
  assign n37921 = n2982 | n2983;
  assign n37922 = n2986 | n2987;
  assign n37923 = n2988 | n2989;
  assign n37924 = n3000 | n3001;
  assign n37925 = n3004 | n3005;
  assign n37926 = n3006 | n3007;
  assign n37927 = n3010 | n3011;
  assign n37928 = n3012 | n3013;
  assign n37929 = n3014 | ~n3015;
  assign n37930 = n3025 | n3026;
  assign n37931 = n3029 | n3030;
  assign n37932 = n3031 | n3032;
  assign n37933 = n3043 | n3044;
  assign n37934 = n3047 | n3048;
  assign n37935 = n3049 | n3050;
  assign n37936 = n3059 | n3060;
  assign n37937 = n3063 | n3064;
  assign n37938 = n3065 | n3066;
  assign n37939 = n3071 | ~n3072;
  assign n37940 = n3080 | n3081;
  assign n37941 = n3084 | n3085;
  assign n37942 = n3086 | n3087;
  assign n37943 = n3100 | n3101;
  assign n37944 = n3104 | n3105;
  assign n37945 = n3106 | n3107;
  assign n37946 = n3116 | n3117;
  assign n37947 = n3120 | n3121;
  assign n37948 = n3122 | n3123;
  assign n37949 = n3129 | n3130;
  assign n37950 = n3138 | n3139;
  assign n37951 = n3142 | n3143;
  assign n37952 = n3144 | n3145;
  assign n37953 = n3151 | n3152;
  assign n37954 = n3165 | n3166;
  assign n37955 = n3176 | n3173 | n3175;
  assign n37956 = n3178 | n3179;
  assign n37957 = n3180 | n3181;
  assign n37958 = n3186 | n3187;
  assign n37959 = n3195 | n3196;
  assign n37960 = n3199 | n3200;
  assign n37961 = n3201 | n3202;
  assign n37962 = n3207 | ~n3208;
  assign n37963 = n3218 | n3219;
  assign n37964 = n3222 | n3223;
  assign n37965 = n3224 | n3225;
  assign n37966 = n3226 | ~n3227;
  assign n37967 = n3239 | n3240;
  assign n37968 = n3241 | n3242;
  assign n37969 = n3243 | ~n3244;
  assign n37970 = n3250 | n3251;
  assign n37971 = n3258 | n3259;
  assign n37972 = n3260 | n3261;
  assign n37973 = n3262 | ~n3263;
  assign n37974 = n3275 | n3276;
  assign n37975 = n3277 | n3278;
  assign n37976 = n3279 | ~n3280;
  assign n37977 = n3284 | n3285;
  assign n37978 = n3286 | n3287;
  assign n37979 = n3288 | ~n3289;
  assign n37980 = n3293 | n3294;
  assign n37981 = n3295 | n3296;
  assign n37982 = n3297 | ~n3298;
  assign n37983 = n3302 | n3303;
  assign n37984 = n3304 | n3305;
  assign n37985 = n3306 | ~n3307;
  assign n37986 = n3311 | n3312;
  assign n37987 = n3313 | n3314;
  assign n37988 = n3315 | ~n3316;
  assign n37989 = n3322 | ~n3323;
  assign n37990 = n3327 | n3328;
  assign n37991 = n3329 | n3330;
  assign n37992 = n3331 | ~n3332;
  assign n37993 = n3336 | n3337;
  assign n37994 = n3338 | n3339;
  assign n37995 = n3340 | ~n3341;
  assign n37996 = n3345 | n3346;
  assign n37997 = n3347 | n3348;
  assign n37998 = n3349 | ~n3350;
  assign n37999 = n3361 | n3362;
  assign n38000 = n3365 | n3366;
  assign n38001 = n3367 | n3368;
  assign n38002 = n3377 | n3378;
  assign n38003 = n3381 | n3382;
  assign n38004 = n3383 | n3384;
  assign n38005 = n3393 | n3394;
  assign n38006 = n3397 | n3398;
  assign n38007 = n3399 | n3400;
  assign n38008 = n3409 | n3410;
  assign n38009 = n3413 | n3414;
  assign n38010 = n3415 | n3416;
  assign n38011 = n3425 | n3426;
  assign n38012 = n3429 | n3430;
  assign n38013 = n3431 | n3432;
  assign n38014 = n3441 | n3442;
  assign n38015 = n3445 | n3446;
  assign n38016 = n3447 | n3448;
  assign n38017 = n3456 | n3457;
  assign n38018 = n3460 | n3461;
  assign n38019 = n3462 | n3463;
  assign n38020 = n3469 | ~n3470;
  assign n38021 = n3476 | ~n3477;
  assign n38022 = n3487 | n3488;
  assign n38023 = n3491 | n3492;
  assign n38024 = n3493 | n3494;
  assign n38025 = n3498 | n3499;
  assign n38026 = n3500 | n3501;
  assign n38027 = n3502 | ~n3503;
  assign n38028 = n3509 | n3510;
  assign n38029 = n3511 | n3512;
  assign n38030 = n3513 | ~n3514;
  assign n38031 = n3517 | n3518;
  assign n38032 = n3522 | n3523;
  assign n38033 = n3524 | n3525;
  assign n38034 = n3526 | ~n3527;
  assign n38035 = n3530 | n3531;
  assign n38036 = n3541 | n3542;
  assign n38037 = n3543 | n3544;
  assign n38038 = n3545 | ~n3546;
  assign n38039 = n3549 | n3550;
  assign n38040 = n3573 | n3574;
  assign n38041 = n3577 | n3578;
  assign n38042 = n3579 | n3580;
  assign n38043 = n3585 | ~n3586;
  assign n38044 = n3598 | n3599;
  assign n38045 = n3602 | n3603;
  assign n38046 = n3604 | n3605;
  assign n38047 = n3616 | n3617;
  assign n38048 = n3620 | n3621;
  assign n38049 = n3622 | n3623;
  assign n38050 = n3634 | n3635;
  assign n38051 = n3638 | n3639;
  assign n38052 = n3640 | n3641;
  assign n38053 = n3652 | n3653;
  assign n38054 = n3656 | n3657;
  assign n38055 = n3658 | n3659;
  assign n38056 = n3670 | n3671;
  assign n38057 = n3674 | n3675;
  assign n38058 = n3676 | n3677;
  assign n38059 = n3686 | n3687;
  assign n38060 = n3690 | n3691;
  assign n38061 = n3692 | n3693;
  assign n38062 = n3696 | n3697;
  assign n38063 = n3698 | n3699;
  assign n38064 = n3700 | ~n3701;
  assign n38065 = n3711 | n3712;
  assign n38066 = n3715 | n3716;
  assign n38067 = n3717 | n3718;
  assign n38068 = n3727 | n3728;
  assign n38069 = n3731 | n3732;
  assign n38070 = n3733 | n3734;
  assign n38071 = n3739 | ~n3740;
  assign n38072 = n3748 | n3749;
  assign n38073 = n3752 | n3753;
  assign n38074 = n3754 | n3755;
  assign n38075 = n3768 | n3769;
  assign n38076 = n3772 | n3773;
  assign n38077 = n3774 | n3775;
  assign n38078 = n3784 | n3785;
  assign n38079 = n3788 | n3789;
  assign n38080 = n3790 | n3791;
  assign n38081 = n3796 | ~n3797;
  assign n38082 = n3805 | n3806;
  assign n38083 = n3809 | n3810;
  assign n38084 = n3811 | n3812;
  assign n38085 = n3823 | n3824;
  assign n38086 = n3827 | n3828;
  assign n38087 = n3829 | n3830;
  assign n38088 = n3835 | ~n3836;
  assign n38089 = n3846 | n3847;
  assign n38090 = n3850 | n3851;
  assign n38091 = n3852 | n3853;
  assign n38092 = n3864 | n3865;
  assign n38093 = n3868 | n3869;
  assign n38094 = n3870 | n3871;
  assign n38095 = n3882 | n3883;
  assign n38096 = n3886 | n3887;
  assign n38097 = n3888 | n3889;
  assign n38098 = n3900 | n3901;
  assign n38099 = n3904 | n3905;
  assign n38100 = n3906 | n3907;
  assign n38101 = n3912 | ~n3913;
  assign n38102 = n3921 | n3922;
  assign n38103 = n3925 | n3926;
  assign n38104 = n3927 | n3928;
  assign n38105 = n3933 | ~n3934;
  assign n38106 = n3942 | n3943;
  assign n38107 = n3946 | n3947;
  assign n38108 = n3948 | n3949;
  assign n38109 = n3962 | n3963;
  assign n38110 = n3966 | n3967;
  assign n38111 = n3968 | n3969;
  assign n38112 = n3978 | n3979;
  assign n38113 = n3982 | n3983;
  assign n38114 = n3984 | n3985;
  assign n38115 = n3991 | n3992;
  assign n38116 = n4000 | n4001;
  assign n38117 = n4004 | n4005;
  assign n38118 = n4006 | n4007;
  assign n38119 = n4013 | n4014;
  assign n38120 = n4027 | n4028;
  assign n38121 = n4038 | n4035 | n4037;
  assign n38122 = n4040 | n4041;
  assign n38123 = n4042 | n4043;
  assign n38124 = n4048 | n4049;
  assign n38125 = n4057 | n4058;
  assign n38126 = n4061 | n4062;
  assign n38127 = n4063 | n4064;
  assign n38128 = n4069 | ~n4070;
  assign n38129 = n4076 | ~n4077;
  assign n38130 = n4083 | n4084;
  assign n38131 = n4087 | n4088;
  assign n38132 = n4089 | n4090;
  assign n38133 = n4091 | ~n4092;
  assign n38134 = n4100 | n4101;
  assign n38135 = n4102 | n4103;
  assign n38136 = n4104 | ~n4105;
  assign n38137 = n4117 | n4118;
  assign n38138 = n4119 | n4120;
  assign n38139 = n4121 | ~n4122;
  assign n38140 = n4136 | n4137;
  assign n38141 = n4138 | n4139;
  assign n38142 = n4140 | ~n4141;
  assign n38143 = n4145 | n4146;
  assign n38144 = n4147 | n4148;
  assign n38145 = n4149 | ~n4150;
  assign n38146 = n4162 | n4163;
  assign n38147 = n4164 | n4165;
  assign n38148 = n4166 | ~n4167;
  assign n38149 = n4173 | ~n4174;
  assign n38150 = n4178 | n4179;
  assign n38151 = n4180 | n4181;
  assign n38152 = n4182 | ~n4183;
  assign n38153 = n4187 | n4188;
  assign n38154 = n4189 | n4190;
  assign n38155 = n4191 | ~n4192;
  assign n38156 = n4198 | n4199;
  assign n38157 = n4206 | n4207;
  assign n38158 = n4208 | n4209;
  assign n38159 = n4210 | ~n4211;
  assign n38160 = n4230 | n4231;
  assign n38161 = n4234 | n4235;
  assign n38162 = n4236 | n4237;
  assign n38163 = n4248 | n4249;
  assign n38164 = n4252 | n4253;
  assign n38165 = n4254 | n4255;
  assign n38166 = n4264 | n4265;
  assign n38167 = n4268 | n4269;
  assign n38168 = n4270 | n4271;
  assign n38169 = n4280 | n4281;
  assign n38170 = n4284 | n4285;
  assign n38171 = n4286 | n4287;
  assign n38172 = n4296 | n4297;
  assign n38173 = n4300 | n4301;
  assign n38174 = n4302 | n4303;
  assign n38175 = n4310 | ~n4311;
  assign n38176 = n4320 | ~n4321;
  assign n38177 = n4333 | n4334;
  assign n38178 = n4336 | n4337;
  assign n38179 = n4368 | n4369;
  assign n38180 = n4372 | n4373;
  assign n38181 = n4374 | n4375;
  assign n38182 = n4379 | n4380;
  assign n38183 = n4381 | n4382;
  assign n38184 = n4383 | ~n4384;
  assign n38185 = n4394 | n4395;
  assign n38186 = n4398 | n4399;
  assign n38187 = n4400 | n4401;
  assign n38188 = n4407 | n4408;
  assign n38189 = n4413 | ~n4414;
  assign n38190 = n4417 | n4418;
  assign n38191 = n4419 | n4420;
  assign n38192 = n4421 | ~n4422;
  assign n38193 = n4432 | n4433;
  assign n38194 = n4436 | n4437;
  assign n38195 = n4438 | n4439;
  assign n38196 = n4443 | n4444;
  assign n38197 = n4445 | n4446;
  assign n38198 = n4447 | ~n4448;
  assign n38199 = n4460 | n4461;
  assign n38200 = n4464 | n4465;
  assign n38201 = n4466 | n4467;
  assign n38202 = n4471 | n4472;
  assign n38203 = n4473 | n4474;
  assign n38204 = n4475 | ~n4476;
  assign n38205 = n4484 | ~n4485;
  assign n38206 = n4490 | ~n4491;
  assign n38207 = n4500 | ~n4501;
  assign n38208 = n4504 | n4505;
  assign n38209 = n4513 | n4514;
  assign n38210 = n4517 | n4518;
  assign n38211 = n4519 | n4520;
  assign n38212 = n4531 | n4532;
  assign n38213 = n4535 | n4536;
  assign n38214 = n4537 | n4538;
  assign n38215 = n4551 | n4552;
  assign n38216 = n4555 | n4556;
  assign n38217 = n4557 | n4558;
  assign n38218 = n4569 | n4570;
  assign n38219 = n4573 | n4574;
  assign n38220 = n4575 | n4576;
  assign n38221 = n4581 | ~n4582;
  assign n38222 = n4592 | n4593;
  assign n38223 = n4596 | n4597;
  assign n38224 = n4598 | n4599;
  assign n38225 = n4608 | n4609;
  assign n38226 = n4612 | n4613;
  assign n38227 = n4614 | n4615;
  assign n38228 = n4620 | ~n4621;
  assign n38229 = n4631 | n4632;
  assign n38230 = n4635 | n4636;
  assign n38231 = n4637 | n4638;
  assign n38232 = n4649 | n4650;
  assign n38233 = n4653 | n4654;
  assign n38234 = n4655 | n4656;
  assign n38235 = n4667 | n4668;
  assign n38236 = n4671 | n4672;
  assign n38237 = n4673 | n4674;
  assign n38238 = n4685 | n4686;
  assign n38239 = n4689 | n4690;
  assign n38240 = n4691 | n4692;
  assign n38241 = n4703 | n4704;
  assign n38242 = n4707 | n4708;
  assign n38243 = n4709 | n4710;
  assign n38244 = n4721 | n4722;
  assign n38245 = n4725 | n4726;
  assign n38246 = n4727 | n4728;
  assign n38247 = n4739 | n4740;
  assign n38248 = n4743 | n4744;
  assign n38249 = n4745 | n4746;
  assign n38250 = n4755 | n4756;
  assign n38251 = n4759 | n4760;
  assign n38252 = n4761 | n4762;
  assign n38253 = n4767 | ~n4768;
  assign n38254 = n4776 | n4777;
  assign n38255 = n4780 | n4781;
  assign n38256 = n4782 | n4783;
  assign n38257 = n4796 | n4797;
  assign n38258 = n4800 | n4801;
  assign n38259 = n4802 | n4803;
  assign n38260 = n4814 | n4815;
  assign n38261 = n4818 | n4819;
  assign n38262 = n4820 | n4821;
  assign n38263 = n4830 | n4831;
  assign n38264 = n4834 | n4835;
  assign n38265 = n4836 | n4837;
  assign n38266 = n4842 | ~n4843;
  assign n38267 = n4851 | n4852;
  assign n38268 = n4855 | n4856;
  assign n38269 = n4857 | n4858;
  assign n38270 = n4871 | n4872;
  assign n38271 = n4875 | n4876;
  assign n38272 = n4877 | n4878;
  assign n38273 = n4889 | n4890;
  assign n38274 = n4893 | n4894;
  assign n38275 = n4895 | n4896;
  assign n38276 = n4909 | n4910;
  assign n38277 = n4913 | n4914;
  assign n38278 = n4915 | n4916;
  assign n38279 = n4925 | n4926;
  assign n38280 = n4929 | n4930;
  assign n38281 = n4931 | n4932;
  assign n38282 = n4937 | ~n4938;
  assign n38283 = n4946 | n4947;
  assign n38284 = n4950 | n4951;
  assign n38285 = n4952 | n4953;
  assign n38286 = n4958 | ~n4959;
  assign n38287 = n4967 | n4968;
  assign n38288 = n4971 | n4972;
  assign n38289 = n4973 | n4974;
  assign n38290 = n4987 | n4988;
  assign n38291 = n4991 | n4992;
  assign n38292 = n4993 | n4994;
  assign n38293 = n5003 | n5004;
  assign n38294 = n5007 | n5008;
  assign n38295 = n5009 | n5010;
  assign n38296 = n5016 | n5017;
  assign n38297 = n5025 | n5026;
  assign n38298 = n5029 | n5030;
  assign n38299 = n5031 | n5032;
  assign n38300 = n5038 | n5039;
  assign n38301 = n5052 | n5053;
  assign n38302 = n5063 | n5060 | n5062;
  assign n38303 = n5065 | n5066;
  assign n38304 = n5067 | n5068;
  assign n38305 = n5073 | n5074;
  assign n38306 = n5082 | n5083;
  assign n38307 = n5086 | n5087;
  assign n38308 = n5088 | n5089;
  assign n38309 = n5094 | ~n5095;
  assign n38310 = n5101 | ~n5102;
  assign n38311 = n5108 | n5109;
  assign n38312 = n5112 | n5113;
  assign n38313 = n5114 | n5115;
  assign n38314 = n5116 | ~n5117;
  assign n38315 = n5125 | n5126;
  assign n38316 = n5127 | n5128;
  assign n38317 = n5129 | ~n5130;
  assign n38318 = n5138 | n5139;
  assign n38319 = n5140 | n5141;
  assign n38320 = n5142 | ~n5143;
  assign n38321 = n5147 | n5148;
  assign n38322 = n5149 | n5150;
  assign n38323 = n5151 | ~n5152;
  assign n38324 = n5166 | n5167;
  assign n38325 = n5168 | n5169;
  assign n38326 = n5170 | ~n5171;
  assign n38327 = n5175 | n5176;
  assign n38328 = n5177 | n5178;
  assign n38329 = n5179 | ~n5180;
  assign n38330 = n5192 | n5193;
  assign n38331 = n5194 | n5195;
  assign n38332 = n5196 | ~n5197;
  assign n38333 = n5201 | n5202;
  assign n38334 = n5203 | n5204;
  assign n38335 = n5205 | ~n5206;
  assign n38336 = n5210 | n5211;
  assign n38337 = n5212 | n5213;
  assign n38338 = n5214 | ~n5215;
  assign n38339 = n5219 | n5220;
  assign n38340 = n5221 | n5222;
  assign n38341 = n5223 | ~n5224;
  assign n38342 = n5230 | n5231;
  assign n38343 = n5238 | n5239;
  assign n38344 = n5240 | n5241;
  assign n38345 = n5242 | ~n5243;
  assign n38346 = n5251 | n5252;
  assign n38347 = n5253 | n5254;
  assign n38348 = n5255 | ~n5256;
  assign n38349 = n5272 | n5273;
  assign n38350 = n5274 | n5275;
  assign n38351 = n5276 | ~n5277;
  assign n38352 = n5288 | n5289;
  assign n38353 = n5292 | n5293;
  assign n38354 = n5294 | n5295;
  assign n38355 = n5304 | n5305;
  assign n38356 = n5308 | n5309;
  assign n38357 = n5310 | n5311;
  assign n38358 = n5321 | n5322;
  assign n38359 = n5325 | n5326;
  assign n38360 = n5327 | n5328;
  assign n38361 = n5336 | n5337;
  assign n38362 = n5340 | n5341;
  assign n38363 = n5342 | n5343;
  assign n38364 = n5352 | n5353;
  assign n38365 = n5356 | n5357;
  assign n38366 = n5358 | n5359;
  assign n38367 = n5369 | n5370;
  assign n38368 = n5373 | n5374;
  assign n38369 = n5375 | n5376;
  assign n38370 = n5385 | n5386;
  assign n38371 = n5389 | n5390;
  assign n38372 = n5391 | n5392;
  assign n38373 = n5401 | n5402;
  assign n38374 = n5405 | n5406;
  assign n38375 = n5407 | n5408;
  assign n38376 = n5413 | n5414;
  assign n38377 = n5424 | n5421 | n5423;
  assign n38378 = n5426 | n5427;
  assign n38379 = n5428 | n5429;
  assign n38380 = n5436 | n5437;
  assign n38381 = n5439 | n5440;
  assign n38382 = n5445 | n5446;
  assign n38383 = n5451 | ~n5452;
  assign n38384 = n5471 | n5472;
  assign n38385 = n5475 | n5476;
  assign n38386 = n5477 | n5478;
  assign n38387 = n5482 | n5483;
  assign n38388 = n5484 | n5485;
  assign n38389 = n5486 | ~n5487;
  assign n38390 = n5493 | n5494;
  assign n38391 = n5495 | n5496;
  assign n38392 = n5497 | ~n5498;
  assign n38393 = n5501 | n5502;
  assign n38394 = n5503 | n5504;
  assign n38395 = n5505 | ~n5506;
  assign n38396 = n5511 | ~n5512;
  assign n38397 = n5517 | ~n5518;
  assign n38398 = n5531 | n5532;
  assign n38399 = n5535 | n5536;
  assign n38400 = n5537 | n5538;
  assign n38401 = n5544 | n5545;
  assign n38402 = n5550 | ~n5551;
  assign n38403 = n5568 | ~n5569;
  assign n38404 = n5574 | ~n5575;
  assign n38405 = n5584 | ~n5585;
  assign n38406 = n5588 | n5589;
  assign n38407 = n5597 | n5598;
  assign n38408 = n5601 | n5602;
  assign n38409 = n5603 | n5604;
  assign n38410 = n5617 | n5618;
  assign n38411 = n5621 | n5622;
  assign n38412 = n5623 | n5624;
  assign n38413 = n5637 | n5638;
  assign n38414 = n5641 | n5642;
  assign n38415 = n5643 | n5644;
  assign n38416 = n5653 | n5654;
  assign n38417 = n5657 | n5658;
  assign n38418 = n5659 | n5660;
  assign n38419 = n5673 | n5674;
  assign n38420 = n5677 | n5678;
  assign n38421 = n5679 | n5680;
  assign n38422 = n5689 | n5690;
  assign n38423 = n5693 | n5694;
  assign n38424 = n5695 | n5696;
  assign n38425 = n5701 | ~n5702;
  assign n38426 = n5710 | n5711;
  assign n38427 = n5714 | n5715;
  assign n38428 = n5716 | n5717;
  assign n38429 = n5728 | n5729;
  assign n38430 = n5732 | n5733;
  assign n38431 = n5734 | n5735;
  assign n38432 = n5748 | n5749;
  assign n38433 = n5752 | n5753;
  assign n38434 = n5754 | n5755;
  assign n38435 = n5764 | n5765;
  assign n38436 = n5768 | n5769;
  assign n38437 = n5770 | n5771;
  assign n38438 = n5776 | ~n5777;
  assign n38439 = n5787 | n5788;
  assign n38440 = n5791 | n5792;
  assign n38441 = n5793 | n5794;
  assign n38442 = n5805 | n5806;
  assign n38443 = n5809 | n5810;
  assign n38444 = n5811 | n5812;
  assign n38445 = n5823 | n5824;
  assign n38446 = n5827 | n5828;
  assign n38447 = n5829 | n5830;
  assign n38448 = n5841 | n5842;
  assign n38449 = n5845 | n5846;
  assign n38450 = n5847 | n5848;
  assign n38451 = n5859 | n5860;
  assign n38452 = n5863 | n5864;
  assign n38453 = n5865 | n5866;
  assign n38454 = n5877 | n5878;
  assign n38455 = n5881 | n5882;
  assign n38456 = n5883 | n5884;
  assign n38457 = n5895 | n5896;
  assign n38458 = n5899 | n5900;
  assign n38459 = n5901 | n5902;
  assign n38460 = n5911 | n5912;
  assign n38461 = n5915 | n5916;
  assign n38462 = n5917 | n5918;
  assign n38463 = n5923 | ~n5924;
  assign n38464 = n5934 | n5935;
  assign n38465 = n5938 | n5939;
  assign n38466 = n5940 | n5941;
  assign n38467 = n5952 | n5953;
  assign n38468 = n5956 | n5957;
  assign n38469 = n5958 | n5959;
  assign n38470 = n5970 | n5971;
  assign n38471 = n5974 | n5975;
  assign n38472 = n5976 | n5977;
  assign n38473 = n5986 | n5987;
  assign n38474 = n5990 | n5991;
  assign n38475 = n5992 | n5993;
  assign n38476 = n5996 | n5997;
  assign n38477 = n5998 | n5999;
  assign n38478 = n6000 | ~n6001;
  assign n38479 = n6011 | n6012;
  assign n38480 = n6015 | n6016;
  assign n38481 = n6017 | n6018;
  assign n38482 = n6029 | n6030;
  assign n38483 = n6033 | n6034;
  assign n38484 = n6035 | n6036;
  assign n38485 = n6047 | n6048;
  assign n38486 = n6051 | n6052;
  assign n38487 = n6053 | n6054;
  assign n38488 = n6065 | n6066;
  assign n38489 = n6069 | n6070;
  assign n38490 = n6071 | n6072;
  assign n38491 = n6081 | n6082;
  assign n38492 = n6085 | n6086;
  assign n38493 = n6087 | n6088;
  assign n38494 = n6093 | ~n6094;
  assign n38495 = n6102 | n6103;
  assign n38496 = n6106 | n6107;
  assign n38497 = n6108 | n6109;
  assign n38498 = n6114 | ~n6115;
  assign n38499 = n6123 | n6124;
  assign n38500 = n6127 | n6128;
  assign n38501 = n6129 | n6130;
  assign n38502 = n6143 | n6144;
  assign n38503 = n6147 | n6148;
  assign n38504 = n6149 | n6150;
  assign n38505 = n6159 | n6160;
  assign n38506 = n6163 | n6164;
  assign n38507 = n6165 | n6166;
  assign n38508 = n6172 | n6173;
  assign n38509 = n6181 | n6182;
  assign n38510 = n6185 | n6186;
  assign n38511 = n6187 | n6188;
  assign n38512 = n6194 | n6195;
  assign n38513 = n6208 | n6209;
  assign n38514 = n6219 | n6216 | n6218;
  assign n38515 = n6221 | n6222;
  assign n38516 = n6223 | n6224;
  assign n38517 = n6229 | n6230;
  assign n38518 = n6238 | n6239;
  assign n38519 = n6242 | n6243;
  assign n38520 = n6244 | n6245;
  assign n38521 = n6250 | ~n6251;
  assign n38522 = n6257 | ~n6258;
  assign n38523 = n6264 | n6265;
  assign n38524 = n6268 | n6269;
  assign n38525 = n6270 | n6271;
  assign n38526 = n6272 | ~n6273;
  assign n38527 = n6289 | n6290;
  assign n38528 = n6291 | n6292;
  assign n38529 = n6293 | ~n6294;
  assign n38530 = n6300 | n6301;
  assign n38531 = n6310 | n6311;
  assign n38532 = n6318 | n6319;
  assign n38533 = n6320 | n6321;
  assign n38534 = n6322 | ~n6323;
  assign n38535 = n6327 | n6328;
  assign n38536 = n6329 | n6330;
  assign n38537 = n6331 | ~n6332;
  assign n38538 = n6336 | n6337;
  assign n38539 = n6338 | n6339;
  assign n38540 = n6340 | ~n6341;
  assign n38541 = n6349 | n6350;
  assign n38542 = n6351 | n6352;
  assign n38543 = n6353 | ~n6354;
  assign n38544 = n6358 | n6359;
  assign n38545 = n6360 | n6361;
  assign n38546 = n6362 | ~n6363;
  assign n38547 = n6367 | n6368;
  assign n38548 = n6369 | n6370;
  assign n38549 = n6371 | ~n6372;
  assign n38550 = n6376 | n6377;
  assign n38551 = n6378 | n6379;
  assign n38552 = n6380 | ~n6381;
  assign n38553 = n6387 | n6388;
  assign n38554 = n6395 | n6396;
  assign n38555 = n6397 | n6398;
  assign n38556 = n6399 | ~n6400;
  assign n38557 = n6408 | n6409;
  assign n38558 = n6410 | n6411;
  assign n38559 = n6412 | ~n6413;
  assign n38560 = n6417 | n6418;
  assign n38561 = n6419 | n6420;
  assign n38562 = n6421 | ~n6422;
  assign n38563 = n6434 | n6435;
  assign n38564 = n6436 | n6437;
  assign n38565 = n6438 | ~n6439;
  assign n38566 = n6447 | n6448;
  assign n38567 = n6449 | n6450;
  assign n38568 = n6451 | ~n6452;
  assign n38569 = n6456 | n6457;
  assign n38570 = n6458 | n6459;
  assign n38571 = n6460 | ~n6461;
  assign n38572 = n6465 | n6466;
  assign n38573 = n6467 | n6468;
  assign n38574 = n6469 | ~n6470;
  assign n38575 = n6481 | n6482;
  assign n38576 = n6485 | n6486;
  assign n38577 = n6487 | n6488;
  assign n38578 = n6498 | n6499;
  assign n38579 = n6502 | n6503;
  assign n38580 = n6504 | n6505;
  assign n38581 = n6515 | n6516;
  assign n38582 = n6519 | n6520;
  assign n38583 = n6521 | n6522;
  assign n38584 = n6531 | n6532;
  assign n38585 = n6535 | n6536;
  assign n38586 = n6537 | n6538;
  assign n38587 = n6547 | n6548;
  assign n38588 = n6551 | n6552;
  assign n38589 = n6553 | n6554;
  assign n38590 = n6563 | n6564;
  assign n38591 = n6567 | n6568;
  assign n38592 = n6569 | n6570;
  assign n38593 = n6579 | n6580;
  assign n38594 = n6583 | n6584;
  assign n38595 = n6585 | n6586;
  assign n38596 = n6594 | n6595;
  assign n38597 = n6598 | n6599;
  assign n38598 = n6600 | n6601;
  assign n38599 = n6607 | ~n6608;
  assign n38600 = n6614 | ~n6615;
  assign n38601 = n6625 | n6626;
  assign n38602 = n6629 | n6630;
  assign n38603 = n6631 | n6632;
  assign n38604 = n6636 | n6637;
  assign n38605 = n6638 | n6639;
  assign n38606 = n6640 | ~n6641;
  assign n38607 = n6646 | ~n6647;
  assign n38608 = n6668 | n6669;
  assign n38609 = n6670 | n6671;
  assign n38610 = n6672 | ~n6673;
  assign n38611 = n6676 | n6677;
  assign n38612 = n6691 | n6692;
  assign n38613 = n6695 | n6696;
  assign n38614 = n6697 | n6698;
  assign n38615 = n6702 | n6703;
  assign n38616 = n6704 | n6705;
  assign n38617 = n6706 | ~n6707;
  assign n38618 = n6717 | n6718;
  assign n38619 = n6721 | n6722;
  assign n38620 = n6723 | n6724;
  assign n38621 = n6744 | n6745;
  assign n38622 = n6748 | n6749;
  assign n38623 = n6750 | n6751;
  assign n38624 = n6755 | n6756;
  assign n38625 = n6757 | n6758;
  assign n38626 = n6759 | ~n6760;
  assign n38627 = n6765 | ~n6766;
  assign n38628 = n6777 | ~n6778;
  assign n38629 = n6783 | ~n6784;
  assign n38630 = n6793 | ~n6794;
  assign n38631 = n6797 | n6798;
  assign n38632 = n6806 | n6807;
  assign n38633 = n6810 | n6811;
  assign n38634 = n6812 | n6813;
  assign n38635 = n6826 | n6827;
  assign n38636 = n6830 | n6831;
  assign n38637 = n6832 | n6833;
  assign n38638 = n6846 | n6847;
  assign n38639 = n6850 | n6851;
  assign n38640 = n6852 | n6853;
  assign n38641 = n6862 | n6863;
  assign n38642 = n6866 | n6867;
  assign n38643 = n6868 | n6869;
  assign n38644 = n6874 | ~n6875;
  assign n38645 = n6885 | n6886;
  assign n38646 = n6889 | n6890;
  assign n38647 = n6891 | n6892;
  assign n38648 = n6903 | n6904;
  assign n38649 = n6907 | n6908;
  assign n38650 = n6909 | n6910;
  assign n38651 = n6921 | n6922;
  assign n38652 = n6925 | n6926;
  assign n38653 = n6927 | n6928;
  assign n38654 = n6937 | n6938;
  assign n38655 = n6941 | n6942;
  assign n38656 = n6943 | n6944;
  assign n38657 = n6955 | n6956;
  assign n38658 = n6959 | n6960;
  assign n38659 = n6961 | n6962;
  assign n38660 = n6965 | n6966;
  assign n38661 = n6967 | n6968;
  assign n38662 = n6969 | ~n6970;
  assign n38663 = n6978 | n6979;
  assign n38664 = n6982 | n6983;
  assign n38665 = n6984 | n6985;
  assign n38666 = n6990 | ~n6991;
  assign n38667 = n6999 | n7000;
  assign n38668 = n7003 | n7004;
  assign n38669 = n7005 | n7006;
  assign n38670 = n7017 | n7018;
  assign n38671 = n7021 | n7022;
  assign n38672 = n7023 | n7024;
  assign n38673 = n7037 | n7038;
  assign n38674 = n7041 | n7042;
  assign n38675 = n7043 | n7044;
  assign n38676 = n7053 | n7054;
  assign n38677 = n7057 | n7058;
  assign n38678 = n7059 | n7060;
  assign n38679 = n7065 | ~n7066;
  assign n38680 = n7076 | n7077;
  assign n38681 = n7080 | n7081;
  assign n38682 = n7082 | n7083;
  assign n38683 = n7094 | n7095;
  assign n38684 = n7098 | n7099;
  assign n38685 = n7100 | n7101;
  assign n38686 = n7112 | n7113;
  assign n38687 = n7116 | n7117;
  assign n38688 = n7118 | n7119;
  assign n38689 = n7130 | n7131;
  assign n38690 = n7134 | n7135;
  assign n38691 = n7136 | n7137;
  assign n38692 = n7148 | n7149;
  assign n38693 = n7152 | n7153;
  assign n38694 = n7154 | n7155;
  assign n38695 = n7166 | n7167;
  assign n38696 = n7170 | n7171;
  assign n38697 = n7172 | n7173;
  assign n38698 = n7184 | n7185;
  assign n38699 = n7188 | n7189;
  assign n38700 = n7190 | n7191;
  assign n38701 = n7200 | n7201;
  assign n38702 = n7204 | n7205;
  assign n38703 = n7206 | n7207;
  assign n38704 = n7212 | ~n7213;
  assign n38705 = n7223 | n7224;
  assign n38706 = n7227 | n7228;
  assign n38707 = n7229 | n7230;
  assign n38708 = n7239 | n7240;
  assign n38709 = n7243 | n7244;
  assign n38710 = n7245 | n7246;
  assign n38711 = n7251 | ~n7252;
  assign n38712 = n7262 | n7263;
  assign n38713 = n7266 | n7267;
  assign n38714 = n7268 | n7269;
  assign n38715 = n7278 | n7279;
  assign n38716 = n7282 | n7283;
  assign n38717 = n7284 | n7285;
  assign n38718 = n7290 | ~n7291;
  assign n38719 = n7301 | n7302;
  assign n38720 = n7305 | n7306;
  assign n38721 = n7307 | n7308;
  assign n38722 = n7319 | n7320;
  assign n38723 = n7323 | n7324;
  assign n38724 = n7325 | n7326;
  assign n38725 = n7337 | n7338;
  assign n38726 = n7341 | n7342;
  assign n38727 = n7343 | n7344;
  assign n38728 = n7357 | n7358;
  assign n38729 = n7361 | n7362;
  assign n38730 = n7363 | n7364;
  assign n38731 = n7373 | n7374;
  assign n38732 = n7377 | n7378;
  assign n38733 = n7379 | n7380;
  assign n38734 = n7385 | ~n7386;
  assign n38735 = n7394 | n7395;
  assign n38736 = n7398 | n7399;
  assign n38737 = n7400 | n7401;
  assign n38738 = n7406 | ~n7407;
  assign n38739 = n7415 | n7416;
  assign n38740 = n7419 | n7420;
  assign n38741 = n7421 | n7422;
  assign n38742 = n7435 | n7436;
  assign n38743 = n7439 | n7440;
  assign n38744 = n7441 | n7442;
  assign n38745 = n7451 | n7452;
  assign n38746 = n7455 | n7456;
  assign n38747 = n7457 | n7458;
  assign n38748 = n7464 | n7465;
  assign n38749 = n7473 | n7474;
  assign n38750 = n7477 | n7478;
  assign n38751 = n7479 | n7480;
  assign n38752 = n7486 | n7487;
  assign n38753 = n7500 | n7501;
  assign n38754 = n7511 | n7508 | n7510;
  assign n38755 = n7513 | n7514;
  assign n38756 = n7515 | n7516;
  assign n38757 = n7521 | n7522;
  assign n38758 = n7530 | n7531;
  assign n38759 = n7534 | n7535;
  assign n38760 = n7536 | n7537;
  assign n38761 = n7542 | ~n7543;
  assign n38762 = n7549 | ~n7550;
  assign n38763 = n7556 | n7557;
  assign n38764 = n7560 | n7561;
  assign n38765 = n7562 | n7563;
  assign n38766 = n7564 | ~n7565;
  assign n38767 = n7581 | n7582;
  assign n38768 = n7583 | n7584;
  assign n38769 = n7585 | ~n7586;
  assign n38770 = n7604 | n7605;
  assign n38771 = n7606 | n7607;
  assign n38772 = n7608 | ~n7609;
  assign n38773 = n7613 | n7614;
  assign n38774 = n7615 | n7616;
  assign n38775 = n7617 | ~n7618;
  assign n38776 = n7622 | n7623;
  assign n38777 = n7624 | n7625;
  assign n38778 = n7626 | ~n7627;
  assign n38779 = n7635 | n7636;
  assign n38780 = n7637 | n7638;
  assign n38781 = n7639 | ~n7640;
  assign n38782 = n7644 | n7645;
  assign n38783 = n7646 | n7647;
  assign n38784 = n7648 | ~n7649;
  assign n38785 = n7653 | n7654;
  assign n38786 = n7655 | n7656;
  assign n38787 = n7657 | ~n7658;
  assign n38788 = n7662 | n7663;
  assign n38789 = n7664 | n7665;
  assign n38790 = n7666 | ~n7667;
  assign n38791 = n7673 | n7674;
  assign n38792 = n7681 | n7682;
  assign n38793 = n7683 | n7684;
  assign n38794 = n7685 | ~n7686;
  assign n38795 = n7694 | n7695;
  assign n38796 = n7696 | n7697;
  assign n38797 = n7698 | ~n7699;
  assign n38798 = n7703 | n7704;
  assign n38799 = n7705 | n7706;
  assign n38800 = n7707 | ~n7708;
  assign n38801 = n7722 | ~n7723;
  assign n38802 = n7731 | n7732;
  assign n38803 = n7733 | n7734;
  assign n38804 = n7735 | ~n7736;
  assign n38805 = n7740 | n7741;
  assign n38806 = n7742 | n7743;
  assign n38807 = n7744 | ~n7745;
  assign n38808 = n7749 | n7750;
  assign n38809 = n7751 | n7752;
  assign n38810 = n7753 | ~n7754;
  assign n38811 = n7762 | n7763;
  assign n38812 = n7764 | n7765;
  assign n38813 = n7766 | ~n7767;
  assign n38814 = n7771 | n7772;
  assign n38815 = n7773 | n7774;
  assign n38816 = n7775 | ~n7776;
  assign n38817 = n7780 | n7781;
  assign n38818 = n7782 | n7783;
  assign n38819 = n7784 | ~n7785;
  assign n38820 = n7797 | n7798;
  assign n38821 = n7801 | n7802;
  assign n38822 = n7803 | n7804;
  assign n38823 = n7815 | n7816;
  assign n38824 = n7819 | n7820;
  assign n38825 = n7821 | n7822;
  assign n38826 = n7832 | n7833;
  assign n38827 = n7836 | n7837;
  assign n38828 = n7838 | n7839;
  assign n38829 = n7850 | n7851;
  assign n38830 = n7854 | n7855;
  assign n38831 = n7856 | n7857;
  assign n38832 = n7866 | n7867;
  assign n38833 = n7870 | n7871;
  assign n38834 = n7872 | n7873;
  assign n38835 = n7880 | ~n7881;
  assign n38836 = n7890 | ~n7891;
  assign n38837 = n7903 | n7904;
  assign n38838 = n7906 | n7907;
  assign n38839 = n7926 | n7927;
  assign n38840 = n7930 | n7931;
  assign n38841 = n7932 | n7933;
  assign n38842 = n7937 | n7938;
  assign n38843 = n7939 | n7940;
  assign n38844 = n7941 | ~n7942;
  assign n38845 = n7952 | n7953;
  assign n38846 = n7956 | n7957;
  assign n38847 = n7958 | n7959;
  assign n38848 = n7965 | n7966;
  assign n38849 = n7971 | ~n7972;
  assign n38850 = n7975 | n7976;
  assign n38851 = n7977 | n7978;
  assign n38852 = n7979 | ~n7980;
  assign n38853 = n7990 | n7991;
  assign n38854 = n7994 | n7995;
  assign n38855 = n7996 | n7997;
  assign n38856 = n8003 | n8004;
  assign n38857 = n8009 | ~n8010;
  assign n38858 = n8013 | n8014;
  assign n38859 = n8015 | n8016;
  assign n38860 = n8017 | ~n8018;
  assign n38861 = n8028 | n8029;
  assign n38862 = n8032 | n8033;
  assign n38863 = n8034 | n8035;
  assign n38864 = n8039 | n8040;
  assign n38865 = n8041 | n8042;
  assign n38866 = n8043 | ~n8044;
  assign n38867 = n8054 | n8055;
  assign n38868 = n8058 | n8059;
  assign n38869 = n8060 | n8061;
  assign n38870 = n8065 | n8066;
  assign n38871 = n8067 | n8068;
  assign n38872 = n8069 | ~n8070;
  assign n38873 = n8075 | ~n8076;
  assign n38874 = n8089 | n8090;
  assign n38875 = n8093 | n8094;
  assign n38876 = n8095 | n8096;
  assign n38877 = n8100 | n8101;
  assign n38878 = n8102 | n8103;
  assign n38879 = n8104 | ~n8105;
  assign n38880 = n8115 | n8116;
  assign n38881 = n8119 | n8120;
  assign n38882 = n8121 | n8122;
  assign n38883 = n8126 | n8127;
  assign n38884 = n8128 | n8129;
  assign n38885 = n8130 | ~n8131;
  assign n38886 = n8143 | n8144;
  assign n38887 = n8147 | n8148;
  assign n38888 = n8149 | n8150;
  assign n38889 = n8154 | n8155;
  assign n38890 = n8156 | n8157;
  assign n38891 = n8158 | ~n8159;
  assign n38892 = n8167 | ~n8168;
  assign n38893 = n8173 | ~n8174;
  assign n38894 = n8183 | ~n8184;
  assign n38895 = n8187 | n8188;
  assign n38896 = n8196 | n8197;
  assign n38897 = n8200 | n8201;
  assign n38898 = n8202 | n8203;
  assign n38899 = n8216 | n8217;
  assign n38900 = n8220 | n8221;
  assign n38901 = n8222 | n8223;
  assign n38902 = n8236 | n8237;
  assign n38903 = n8240 | n8241;
  assign n38904 = n8242 | n8243;
  assign n38905 = n8254 | n8255;
  assign n38906 = n8258 | n8259;
  assign n38907 = n8260 | n8261;
  assign n38908 = n8272 | n8273;
  assign n38909 = n8276 | n8277;
  assign n38910 = n8278 | n8279;
  assign n38911 = n8290 | n8291;
  assign n38912 = n8294 | n8295;
  assign n38913 = n8296 | n8297;
  assign n38914 = n8308 | n8309;
  assign n38915 = n8312 | n8313;
  assign n38916 = n8314 | n8315;
  assign n38917 = n8324 | n8325;
  assign n38918 = n8328 | n8329;
  assign n38919 = n8330 | n8331;
  assign n38920 = n8336 | ~n8337;
  assign n38921 = n8347 | n8348;
  assign n38922 = n8351 | n8352;
  assign n38923 = n8353 | n8354;
  assign n38924 = n8365 | n8366;
  assign n38925 = n8369 | n8370;
  assign n38926 = n8371 | n8372;
  assign n38927 = n8383 | n8384;
  assign n38928 = n8387 | n8388;
  assign n38929 = n8389 | n8390;
  assign n38930 = n8399 | n8400;
  assign n38931 = n8403 | n8404;
  assign n38932 = n8405 | n8406;
  assign n38933 = n8417 | n8418;
  assign n38934 = n8421 | n8422;
  assign n38935 = n8423 | n8424;
  assign n38936 = n8427 | n8428;
  assign n38937 = n8429 | n8430;
  assign n38938 = n8431 | ~n8432;
  assign n38939 = n8440 | n8441;
  assign n38940 = n8444 | n8445;
  assign n38941 = n8446 | n8447;
  assign n38942 = n8452 | ~n8453;
  assign n38943 = n8461 | n8462;
  assign n38944 = n8465 | n8466;
  assign n38945 = n8467 | n8468;
  assign n38946 = n8479 | n8480;
  assign n38947 = n8483 | n8484;
  assign n38948 = n8485 | n8486;
  assign n38949 = n8499 | n8500;
  assign n38950 = n8503 | n8504;
  assign n38951 = n8505 | n8506;
  assign n38952 = n8515 | n8516;
  assign n38953 = n8519 | n8520;
  assign n38954 = n8521 | n8522;
  assign n38955 = n8527 | ~n8528;
  assign n38956 = n8538 | n8539;
  assign n38957 = n8542 | n8543;
  assign n38958 = n8544 | n8545;
  assign n38959 = n8556 | n8557;
  assign n38960 = n8560 | n8561;
  assign n38961 = n8562 | n8563;
  assign n38962 = n8574 | n8575;
  assign n38963 = n8578 | n8579;
  assign n38964 = n8580 | n8581;
  assign n38965 = n8592 | n8593;
  assign n38966 = n8596 | n8597;
  assign n38967 = n8598 | n8599;
  assign n38968 = n8610 | n8611;
  assign n38969 = n8614 | n8615;
  assign n38970 = n8616 | n8617;
  assign n38971 = n8628 | n8629;
  assign n38972 = n8632 | n8633;
  assign n38973 = n8634 | n8635;
  assign n38974 = n8646 | n8647;
  assign n38975 = n8650 | n8651;
  assign n38976 = n8652 | n8653;
  assign n38977 = n8662 | n8663;
  assign n38978 = n8666 | n8667;
  assign n38979 = n8668 | n8669;
  assign n38980 = n8674 | ~n8675;
  assign n38981 = n8685 | n8686;
  assign n38982 = n8689 | n8690;
  assign n38983 = n8691 | n8692;
  assign n38984 = n8703 | n8704;
  assign n38985 = n8707 | n8708;
  assign n38986 = n8709 | n8710;
  assign n38987 = n8721 | n8722;
  assign n38988 = n8725 | n8726;
  assign n38989 = n8727 | n8728;
  assign n38990 = n8739 | n8740;
  assign n38991 = n8743 | n8744;
  assign n38992 = n8745 | n8746;
  assign n38993 = n8757 | n8758;
  assign n38994 = n8761 | n8762;
  assign n38995 = n8763 | n8764;
  assign n38996 = n8773 | n8774;
  assign n38997 = n8777 | n8778;
  assign n38998 = n8779 | n8780;
  assign n38999 = n8791 | n8792;
  assign n39000 = n8795 | n8796;
  assign n39001 = n8797 | n8798;
  assign n39002 = n8811 | n8812;
  assign n39003 = n8815 | n8816;
  assign n39004 = n8817 | n8818;
  assign n39005 = n8827 | n8828;
  assign n39006 = n8831 | n8832;
  assign n39007 = n8833 | n8834;
  assign n39008 = n8839 | ~n8840;
  assign n39009 = n8848 | n8849;
  assign n39010 = n8852 | n8853;
  assign n39011 = n8854 | n8855;
  assign n39012 = n8860 | ~n8861;
  assign n39013 = n8869 | n8870;
  assign n39014 = n8873 | n8874;
  assign n39015 = n8875 | n8876;
  assign n39016 = n8889 | n8890;
  assign n39017 = n8893 | n8894;
  assign n39018 = n8895 | n8896;
  assign n39019 = n8905 | n8906;
  assign n39020 = n8909 | n8910;
  assign n39021 = n8911 | n8912;
  assign n39022 = n8918 | n8919;
  assign n39023 = n8927 | n8928;
  assign n39024 = n8931 | n8932;
  assign n39025 = n8933 | n8934;
  assign n39026 = n8940 | n8941;
  assign n39027 = n8954 | n8955;
  assign n39028 = n8965 | n8962 | n8964;
  assign n39029 = n8967 | n8968;
  assign n39030 = n8969 | n8970;
  assign n39031 = n8975 | n8976;
  assign n39032 = n8984 | n8985;
  assign n39033 = n8988 | n8989;
  assign n39034 = n8990 | n8991;
  assign n39035 = n8996 | ~n8997;
  assign n39036 = n9003 | ~n9004;
  assign n39037 = n9010 | n9011;
  assign n39038 = n9014 | n9015;
  assign n39039 = n9016 | n9017;
  assign n39040 = n9018 | ~n9019;
  assign n39041 = n9035 | n9036;
  assign n39042 = n9037 | n9038;
  assign n39043 = n9039 | ~n9040;
  assign n39044 = n9052 | n9053;
  assign n39045 = n9054 | n9055;
  assign n39046 = n9056 | ~n9057;
  assign n39047 = n9061 | n9062;
  assign n39048 = n9063 | n9064;
  assign n39049 = n9065 | ~n9066;
  assign n39050 = n9070 | n9071;
  assign n39051 = n9072 | n9073;
  assign n39052 = n9074 | ~n9075;
  assign n39053 = n9079 | n9080;
  assign n39054 = n9081 | n9082;
  assign n39055 = n9083 | ~n9084;
  assign n39056 = n9088 | n9089;
  assign n39057 = n9090 | n9091;
  assign n39058 = n9092 | ~n9093;
  assign n39059 = n9101 | n9102;
  assign n39060 = n9103 | n9104;
  assign n39061 = n9105 | ~n9106;
  assign n39062 = n9112 | n9113;
  assign n39063 = n9116 | n9117;
  assign n39064 = n9118 | n9119;
  assign n39065 = n9120 | ~n9121;
  assign n39066 = n9125 | n9126;
  assign n39067 = n9127 | n9128;
  assign n39068 = n9129 | ~n9130;
  assign n39069 = n9136 | n9137;
  assign n39070 = n9144 | n9145;
  assign n39071 = n9146 | n9147;
  assign n39072 = n9148 | ~n9149;
  assign n39073 = n9157 | n9158;
  assign n39074 = n9159 | n9160;
  assign n39075 = n9161 | ~n9162;
  assign n39076 = n9166 | n9167;
  assign n39077 = n9168 | n9169;
  assign n39078 = n9170 | ~n9171;
  assign n39079 = n9191 | n9192;
  assign n39080 = n9193 | n9194;
  assign n39081 = n9195 | ~n9196;
  assign n39082 = n9200 | n9201;
  assign n39083 = n9202 | n9203;
  assign n39084 = n9204 | ~n9205;
  assign n39085 = n9209 | n9210;
  assign n39086 = n9211 | n9212;
  assign n39087 = n9213 | ~n9214;
  assign n39088 = n9222 | n9223;
  assign n39089 = n9224 | n9225;
  assign n39090 = n9226 | ~n9227;
  assign n39091 = n9231 | n9232;
  assign n39092 = n9233 | n9234;
  assign n39093 = n9235 | ~n9236;
  assign n39094 = n9240 | n9241;
  assign n39095 = n9242 | n9243;
  assign n39096 = n9244 | ~n9245;
  assign n39097 = n9249 | n9250;
  assign n39098 = n9251 | n9252;
  assign n39099 = n9253 | ~n9254;
  assign n39100 = n9258 | n9259;
  assign n39101 = n9260 | n9261;
  assign n39102 = n9262 | ~n9263;
  assign n39103 = n9273 | n9274;
  assign n39104 = n9284 | n9285;
  assign n39105 = n9288 | n9289;
  assign n39106 = n9290 | n9291;
  assign n39107 = n9303 | n9304;
  assign n39108 = n9307 | n9308;
  assign n39109 = n9309 | n9310;
  assign n39110 = n9321 | n9322;
  assign n39111 = n9325 | n9326;
  assign n39112 = n9327 | n9328;
  assign n39113 = n9336 | n9337;
  assign n39114 = n9340 | n9341;
  assign n39115 = n9342 | n9343;
  assign n39116 = n9352 | n9353;
  assign n39117 = n9356 | n9357;
  assign n39118 = n9358 | n9359;
  assign n39119 = n9368 | n9369;
  assign n39120 = n9372 | n9373;
  assign n39121 = n9374 | n9375;
  assign n39122 = n9384 | n9385;
  assign n39123 = n9388 | n9389;
  assign n39124 = n9390 | n9391;
  assign n39125 = n9400 | n9401;
  assign n39126 = n9404 | n9405;
  assign n39127 = n9406 | n9407;
  assign n39128 = n9412 | n9413;
  assign n39129 = n9423 | n9420 | n9422;
  assign n39130 = n9425 | n9426;
  assign n39131 = n9427 | n9428;
  assign n39132 = n9435 | n9436;
  assign n39133 = n9438 | n9439;
  assign n39134 = n9444 | n9445;
  assign n39135 = n9450 | ~n9451;
  assign n39136 = n9470 | n9471;
  assign n39137 = n9474 | n9475;
  assign n39138 = n9476 | n9477;
  assign n39139 = n9481 | n9482;
  assign n39140 = n9483 | n9484;
  assign n39141 = n9485 | ~n9486;
  assign n39142 = n9492 | n9493;
  assign n39143 = n9494 | n9495;
  assign n39144 = n9496 | ~n9497;
  assign n39145 = n9500 | n9501;
  assign n39146 = n9502 | n9503;
  assign n39147 = n9504 | ~n9505;
  assign n39148 = n9510 | ~n9511;
  assign n39149 = n9516 | ~n9517;
  assign n39150 = n9530 | n9531;
  assign n39151 = n9534 | n9535;
  assign n39152 = n9536 | n9537;
  assign n39153 = n9541 | n9542;
  assign n39154 = n9543 | n9544;
  assign n39155 = n9545 | ~n9546;
  assign n39156 = n9556 | n9557;
  assign n39157 = n9560 | n9561;
  assign n39158 = n9562 | n9563;
  assign n39159 = n9569 | n9570;
  assign n39160 = n9575 | ~n9576;
  assign n39161 = n9589 | n9590;
  assign n39162 = n9593 | n9594;
  assign n39163 = n9595 | n9596;
  assign n39164 = n9600 | n9601;
  assign n39165 = n9602 | n9603;
  assign n39166 = n9604 | ~n9605;
  assign n39167 = n9615 | n9616;
  assign n39168 = n9619 | n9620;
  assign n39169 = n9621 | n9622;
  assign n39170 = n9626 | n9627;
  assign n39171 = n9628 | n9629;
  assign n39172 = n9630 | ~n9631;
  assign n39173 = n9641 | n9642;
  assign n39174 = n9645 | n9646;
  assign n39175 = n9647 | n9648;
  assign n39176 = n9654 | n9655;
  assign n39177 = n9660 | ~n9661;
  assign n39178 = n9664 | n9665;
  assign n39179 = n9666 | n9667;
  assign n39180 = n9668 | ~n9669;
  assign n39181 = n9674 | ~n9675;
  assign n39182 = n9685 | n9686;
  assign n39183 = n9689 | n9690;
  assign n39184 = n9691 | n9692;
  assign n39185 = n9697 | ~n9698;
  assign n39186 = n9708 | n9709;
  assign n39187 = n9712 | n9713;
  assign n39188 = n9714 | n9715;
  assign n39189 = n9728 | n9729;
  assign n39190 = n9732 | n9733;
  assign n39191 = n9734 | n9735;
  assign n39192 = n9746 | n9747;
  assign n39193 = n9750 | n9751;
  assign n39194 = n9752 | n9753;
  assign n39195 = n9764 | n9765;
  assign n39196 = n9768 | n9769;
  assign n39197 = n9770 | n9771;
  assign n39198 = n9782 | n9783;
  assign n39199 = n9786 | n9787;
  assign n39200 = n9788 | n9789;
  assign n39201 = n9800 | n9801;
  assign n39202 = n9804 | n9805;
  assign n39203 = n9806 | n9807;
  assign n39204 = n9818 | n9819;
  assign n39205 = n9822 | n9823;
  assign n39206 = n9824 | n9825;
  assign n39207 = n9836 | n9837;
  assign n39208 = n9840 | n9841;
  assign n39209 = n9842 | n9843;
  assign n39210 = n9854 | n9855;
  assign n39211 = n9858 | n9859;
  assign n39212 = n9860 | n9861;
  assign n39213 = n9870 | n9871;
  assign n39214 = n9874 | n9875;
  assign n39215 = n9876 | n9877;
  assign n39216 = n9882 | ~n9883;
  assign n39217 = n9893 | n9894;
  assign n39218 = n9897 | n9898;
  assign n39219 = n9899 | n9900;
  assign n39220 = n9911 | n9912;
  assign n39221 = n9915 | n9916;
  assign n39222 = n9917 | n9918;
  assign n39223 = n9929 | n9930;
  assign n39224 = n9933 | n9934;
  assign n39225 = n9935 | n9936;
  assign n39226 = n9945 | n9946;
  assign n39227 = n9949 | n9950;
  assign n39228 = n9951 | n9952;
  assign n39229 = n9963 | n9964;
  assign n39230 = n9967 | n9968;
  assign n39231 = n9969 | n9970;
  assign n39232 = n9973 | n9974;
  assign n39233 = n9975 | n9976;
  assign n39234 = n9977 | ~n9978;
  assign n39235 = n9986 | n9987;
  assign n39236 = n9990 | n9991;
  assign n39237 = n9992 | n9993;
  assign n39238 = n9998 | ~n9999;
  assign n39239 = n10007 | n10008;
  assign n39240 = n10011 | n10012;
  assign n39241 = n10013 | n10014;
  assign n39242 = n10025 | n10026;
  assign n39243 = n10029 | n10030;
  assign n39244 = n10031 | n10032;
  assign n39245 = n10045 | n10046;
  assign n39246 = n10049 | n10050;
  assign n39247 = n10051 | n10052;
  assign n39248 = n10061 | n10062;
  assign n39249 = n10065 | n10066;
  assign n39250 = n10067 | n10068;
  assign n39251 = n10073 | ~n10074;
  assign n39252 = n10084 | n10085;
  assign n39253 = n10088 | n10089;
  assign n39254 = n10090 | n10091;
  assign n39255 = n10100 | n10101;
  assign n39256 = n10104 | n10105;
  assign n39257 = n10106 | n10107;
  assign n39258 = n10112 | ~n10113;
  assign n39259 = n10121 | n10122;
  assign n39260 = n10125 | n10126;
  assign n39261 = n10127 | n10128;
  assign n39262 = n10133 | ~n10134;
  assign n39263 = n10144 | n10145;
  assign n39264 = n10148 | n10149;
  assign n39265 = n10150 | n10151;
  assign n39266 = n10162 | n10163;
  assign n39267 = n10166 | n10167;
  assign n39268 = n10168 | n10169;
  assign n39269 = n10180 | n10181;
  assign n39270 = n10184 | n10185;
  assign n39271 = n10186 | n10187;
  assign n39272 = n10198 | n10199;
  assign n39273 = n10202 | n10203;
  assign n39274 = n10204 | n10205;
  assign n39275 = n10216 | n10217;
  assign n39276 = n10220 | n10221;
  assign n39277 = n10222 | n10223;
  assign n39278 = n10234 | n10235;
  assign n39279 = n10238 | n10239;
  assign n39280 = n10240 | n10241;
  assign n39281 = n10250 | n10251;
  assign n39282 = n10254 | n10255;
  assign n39283 = n10256 | n10257;
  assign n39284 = n10260 | n10261;
  assign n39285 = n10262 | n10263;
  assign n39286 = n10264 | ~n10265;
  assign n39287 = n10275 | n10276;
  assign n39288 = n10279 | n10280;
  assign n39289 = n10281 | n10282;
  assign n39290 = n10293 | n10294;
  assign n39291 = n10297 | n10298;
  assign n39292 = n10299 | n10300;
  assign n39293 = n10311 | n10312;
  assign n39294 = n10315 | n10316;
  assign n39295 = n10317 | n10318;
  assign n39296 = n10329 | n10330;
  assign n39297 = n10333 | n10334;
  assign n39298 = n10335 | n10336;
  assign n39299 = n10347 | n10348;
  assign n39300 = n10351 | n10352;
  assign n39301 = n10353 | n10354;
  assign n39302 = n10367 | n10368;
  assign n39303 = n10371 | n10372;
  assign n39304 = n10373 | n10374;
  assign n39305 = n10383 | n10384;
  assign n39306 = n10387 | n10388;
  assign n39307 = n10389 | n10390;
  assign n39308 = n10395 | ~n10396;
  assign n39309 = n10404 | n10405;
  assign n39310 = n10408 | n10409;
  assign n39311 = n10410 | n10411;
  assign n39312 = n10416 | ~n10417;
  assign n39313 = n10425 | n10426;
  assign n39314 = n10429 | n10430;
  assign n39315 = n10431 | n10432;
  assign n39316 = n10445 | n10446;
  assign n39317 = n10449 | n10450;
  assign n39318 = n10451 | n10452;
  assign n39319 = n10461 | n10462;
  assign n39320 = n10465 | n10466;
  assign n39321 = n10467 | n10468;
  assign n39322 = n10474 | n10475;
  assign n39323 = n10483 | n10484;
  assign n39324 = n10487 | n10488;
  assign n39325 = n10489 | n10490;
  assign n39326 = n10496 | n10497;
  assign n39327 = n10510 | n10511;
  assign n39328 = n10521 | n10518 | n10520;
  assign n39329 = n10523 | n10524;
  assign n39330 = n10525 | n10526;
  assign n39331 = n10531 | n10532;
  assign n39332 = n10540 | n10541;
  assign n39333 = n10544 | n10545;
  assign n39334 = n10546 | n10547;
  assign n39335 = n10552 | ~n10553;
  assign n39336 = n10563 | n10564;
  assign n39337 = n10567 | n10568;
  assign n39338 = n10569 | n10570;
  assign n39339 = n10571 | ~n10572;
  assign n39340 = n10588 | n10589;
  assign n39341 = n10590 | n10591;
  assign n39342 = n10592 | ~n10593;
  assign n39343 = n10607 | n10608;
  assign n39344 = n10609 | n10610;
  assign n39345 = n10611 | ~n10612;
  assign n39346 = n10616 | n10617;
  assign n39347 = n10618 | n10619;
  assign n39348 = n10620 | ~n10621;
  assign n39349 = n10627 | ~n10628;
  assign n39350 = n10632 | n10633;
  assign n39351 = n10634 | n10635;
  assign n39352 = n10636 | ~n10637;
  assign n39353 = n10641 | n10642;
  assign n39354 = n10643 | n10644;
  assign n39355 = n10645 | ~n10646;
  assign n39356 = n10650 | n10651;
  assign n39357 = n10652 | n10653;
  assign n39358 = n10654 | ~n10655;
  assign n39359 = n10661 | n10662;
  assign n39360 = n10665 | n10666;
  assign n39361 = n10667 | n10668;
  assign n39362 = n10669 | ~n10670;
  assign n39363 = n10674 | n10675;
  assign n39364 = n10676 | n10677;
  assign n39365 = n10678 | ~n10679;
  assign n39366 = n10693 | n10694;
  assign n39367 = n10701 | n10702;
  assign n39368 = n10703 | n10704;
  assign n39369 = n10705 | ~n10706;
  assign n39370 = n10710 | n10711;
  assign n39371 = n10712 | n10713;
  assign n39372 = n10714 | ~n10715;
  assign n39373 = n10735 | n10736;
  assign n39374 = n10737 | n10738;
  assign n39375 = n10739 | ~n10740;
  assign n39376 = n10744 | n10745;
  assign n39377 = n10746 | n10747;
  assign n39378 = n10748 | ~n10749;
  assign n39379 = n10753 | n10754;
  assign n39380 = n10755 | n10756;
  assign n39381 = n10757 | ~n10758;
  assign n39382 = n10766 | n10767;
  assign n39383 = n10768 | n10769;
  assign n39384 = n10770 | ~n10771;
  assign n39385 = n10775 | n10776;
  assign n39386 = n10777 | n10778;
  assign n39387 = n10779 | ~n10780;
  assign n39388 = n10784 | n10785;
  assign n39389 = n10786 | n10787;
  assign n39390 = n10788 | ~n10789;
  assign n39391 = n10793 | n10794;
  assign n39392 = n10795 | n10796;
  assign n39393 = n10797 | ~n10798;
  assign n39394 = n10802 | n10803;
  assign n39395 = n10804 | n10805;
  assign n39396 = n10806 | ~n10807;
  assign n39397 = n10817 | n10818;
  assign n39398 = n10823 | n10824;
  assign n39399 = n10827 | n10828;
  assign n39400 = n10829 | n10830;
  assign n39401 = n10831 | ~n10832;
  assign n39402 = n10851 | n10852;
  assign n39403 = n10855 | n10856;
  assign n39404 = n10857 | n10858;
  assign n39405 = n10867 | n10868;
  assign n39406 = n10871 | n10872;
  assign n39407 = n10873 | n10874;
  assign n39408 = n10884 | n10885;
  assign n39409 = n10888 | n10889;
  assign n39410 = n10890 | n10891;
  assign n39411 = n10903 | n10904;
  assign n39412 = n10907 | n10908;
  assign n39413 = n10909 | n10910;
  assign n39414 = n10919 | n10920;
  assign n39415 = n10923 | n10924;
  assign n39416 = n10925 | n10926;
  assign n39417 = n10935 | n10936;
  assign n39418 = n10939 | n10940;
  assign n39419 = n10941 | n10942;
  assign n39420 = n10951 | n10952;
  assign n39421 = n10955 | n10956;
  assign n39422 = n10957 | n10958;
  assign n39423 = n10967 | n10968;
  assign n39424 = n10971 | n10972;
  assign n39425 = n10973 | n10974;
  assign n39426 = n10982 | n10983;
  assign n39427 = n10986 | n10987;
  assign n39428 = n10988 | n10989;
  assign n39429 = n10995 | ~n10996;
  assign n39430 = n11002 | ~n11003;
  assign n39431 = n11013 | n11014;
  assign n39432 = n11017 | n11018;
  assign n39433 = n11019 | n11020;
  assign n39434 = n11024 | n11025;
  assign n39435 = n11026 | n11027;
  assign n39436 = n11028 | ~n11029;
  assign n39437 = n11034 | ~n11035;
  assign n39438 = n11056 | n11057;
  assign n39439 = n11058 | n11059;
  assign n39440 = n11060 | ~n11061;
  assign n39441 = n11064 | n11065;
  assign n39442 = n11079 | n11080;
  assign n39443 = n11083 | n11084;
  assign n39444 = n11085 | n11086;
  assign n39445 = n11090 | n11091;
  assign n39446 = n11092 | n11093;
  assign n39447 = n11094 | ~n11095;
  assign n39448 = n11105 | n11106;
  assign n39449 = n11109 | n11110;
  assign n39450 = n11111 | n11112;
  assign n39451 = n11116 | n11117;
  assign n39452 = n11118 | n11119;
  assign n39453 = n11120 | ~n11121;
  assign n39454 = n11131 | n11132;
  assign n39455 = n11135 | n11136;
  assign n39456 = n11137 | n11138;
  assign n39457 = n11152 | n11153;
  assign n39458 = n11156 | n11157;
  assign n39459 = n11158 | n11159;
  assign n39460 = n11163 | n11164;
  assign n39461 = n11165 | n11166;
  assign n39462 = n11167 | ~n11168;
  assign n39463 = n11173 | ~n11174;
  assign n39464 = n11187 | n11188;
  assign n39465 = n11191 | n11192;
  assign n39466 = n11193 | n11194;
  assign n39467 = n11198 | n11199;
  assign n39468 = n11200 | n11201;
  assign n39469 = n11202 | ~n11203;
  assign n39470 = n11213 | n11214;
  assign n39471 = n11217 | n11218;
  assign n39472 = n11219 | n11220;
  assign n39473 = n11230 | n11231;
  assign n39474 = n11232 | n11233;
  assign n39475 = n11234 | ~n11235;
  assign n39476 = n11238 | n11239;
  assign n39477 = n11243 | n11244;
  assign n39478 = n11245 | n11246;
  assign n39479 = n11247 | ~n11248;
  assign n39480 = n11251 | n11252;
  assign n39481 = n11265 | n11266;
  assign n39482 = n11269 | n11270;
  assign n39483 = n11271 | n11272;
  assign n39484 = n11283 | n11284;
  assign n39485 = n11287 | n11288;
  assign n39486 = n11289 | n11290;
  assign n39487 = n11301 | n11302;
  assign n39488 = n11305 | n11306;
  assign n39489 = n11307 | n11308;
  assign n39490 = n11311 | n11312;
  assign n39491 = n11321 | n11322;
  assign n39492 = n11325 | n11326;
  assign n39493 = n11327 | n11328;
  assign n39494 = n11333 | ~n11334;
  assign n39495 = n11342 | n11343;
  assign n39496 = n11346 | n11347;
  assign n39497 = n11348 | n11349;
  assign n39498 = n11354 | ~n11355;
  assign n39499 = n11363 | n11364;
  assign n39500 = n11367 | n11368;
  assign n39501 = n11369 | n11370;
  assign n39502 = n11383 | n11384;
  assign n39503 = n11387 | n11388;
  assign n39504 = n11389 | n11390;
  assign n39505 = n11401 | n11402;
  assign n39506 = n11405 | n11406;
  assign n39507 = n11407 | n11408;
  assign n39508 = n11419 | n11420;
  assign n39509 = n11423 | n11424;
  assign n39510 = n11425 | n11426;
  assign n39511 = n11439 | n11440;
  assign n39512 = n11443 | n11444;
  assign n39513 = n11445 | n11446;
  assign n39514 = n11457 | n11458;
  assign n39515 = n11461 | n11462;
  assign n39516 = n11463 | n11464;
  assign n39517 = n11475 | n11476;
  assign n39518 = n11479 | n11480;
  assign n39519 = n11481 | n11482;
  assign n39520 = n11493 | n11494;
  assign n39521 = n11497 | n11498;
  assign n39522 = n11499 | n11500;
  assign n39523 = n11511 | n11512;
  assign n39524 = n11515 | n11516;
  assign n39525 = n11517 | n11518;
  assign n39526 = n11527 | n11528;
  assign n39527 = n11531 | n11532;
  assign n39528 = n11533 | n11534;
  assign n39529 = n11539 | ~n11540;
  assign n39530 = n11550 | n11551;
  assign n39531 = n11554 | n11555;
  assign n39532 = n11556 | n11557;
  assign n39533 = n11568 | n11569;
  assign n39534 = n11572 | n11573;
  assign n39535 = n11574 | n11575;
  assign n39536 = n11586 | n11587;
  assign n39537 = n11590 | n11591;
  assign n39538 = n11592 | n11593;
  assign n39539 = n11602 | n11603;
  assign n39540 = n11606 | n11607;
  assign n39541 = n11608 | n11609;
  assign n39542 = n11620 | n11621;
  assign n39543 = n11624 | n11625;
  assign n39544 = n11626 | n11627;
  assign n39545 = n11630 | n11631;
  assign n39546 = n11632 | n11633;
  assign n39547 = n11634 | ~n11635;
  assign n39548 = n11643 | n11644;
  assign n39549 = n11647 | n11648;
  assign n39550 = n11649 | n11650;
  assign n39551 = n11655 | ~n11656;
  assign n39552 = n11664 | n11665;
  assign n39553 = n11668 | n11669;
  assign n39554 = n11670 | n11671;
  assign n39555 = n11682 | n11683;
  assign n39556 = n11686 | n11687;
  assign n39557 = n11688 | n11689;
  assign n39558 = n11694 | ~n11695;
  assign n39559 = n11705 | n11706;
  assign n39560 = n11709 | n11710;
  assign n39561 = n11711 | n11712;
  assign n39562 = n11721 | n11722;
  assign n39563 = n11725 | n11726;
  assign n39564 = n11727 | n11728;
  assign n39565 = n11741 | n11742;
  assign n39566 = n11745 | n11746;
  assign n39567 = n11747 | n11748;
  assign n39568 = n11757 | n11758;
  assign n39569 = n11761 | n11762;
  assign n39570 = n11763 | n11764;
  assign n39571 = n11769 | ~n11770;
  assign n39572 = n11778 | n11779;
  assign n39573 = n11782 | n11783;
  assign n39574 = n11784 | n11785;
  assign n39575 = n11790 | ~n11791;
  assign n39576 = n11801 | n11802;
  assign n39577 = n11805 | n11806;
  assign n39578 = n11807 | n11808;
  assign n39579 = n11819 | n11820;
  assign n39580 = n11823 | n11824;
  assign n39581 = n11825 | n11826;
  assign n39582 = n11837 | n11838;
  assign n39583 = n11841 | n11842;
  assign n39584 = n11843 | n11844;
  assign n39585 = n11855 | n11856;
  assign n39586 = n11859 | n11860;
  assign n39587 = n11861 | n11862;
  assign n39588 = n11873 | n11874;
  assign n39589 = n11877 | n11878;
  assign n39590 = n11879 | n11880;
  assign n39591 = n11889 | n11890;
  assign n39592 = n11893 | n11894;
  assign n39593 = n11895 | n11896;
  assign n39594 = n11901 | ~n11902;
  assign n39595 = n11912 | n11913;
  assign n39596 = n11916 | n11917;
  assign n39597 = n11918 | n11919;
  assign n39598 = n11930 | n11931;
  assign n39599 = n11934 | n11935;
  assign n39600 = n11936 | n11937;
  assign n39601 = n11948 | n11949;
  assign n39602 = n11952 | n11953;
  assign n39603 = n11954 | n11955;
  assign n39604 = n11966 | n11967;
  assign n39605 = n11970 | n11971;
  assign n39606 = n11972 | n11973;
  assign n39607 = n11982 | n11983;
  assign n39608 = n11986 | n11987;
  assign n39609 = n11988 | n11989;
  assign n39610 = n12000 | n12001;
  assign n39611 = n12004 | n12005;
  assign n39612 = n12006 | n12007;
  assign n39613 = n12020 | n12021;
  assign n39614 = n12024 | n12025;
  assign n39615 = n12026 | n12027;
  assign n39616 = n12036 | n12037;
  assign n39617 = n12040 | n12041;
  assign n39618 = n12042 | n12043;
  assign n39619 = n12048 | ~n12049;
  assign n39620 = n12057 | n12058;
  assign n39621 = n12061 | n12062;
  assign n39622 = n12063 | n12064;
  assign n39623 = n12069 | ~n12070;
  assign n39624 = n12078 | n12079;
  assign n39625 = n12082 | n12083;
  assign n39626 = n12084 | n12085;
  assign n39627 = n12098 | n12099;
  assign n39628 = n12102 | n12103;
  assign n39629 = n12104 | n12105;
  assign n39630 = n12114 | n12115;
  assign n39631 = n12118 | n12119;
  assign n39632 = n12120 | n12121;
  assign n39633 = n12127 | n12128;
  assign n39634 = n12136 | n12137;
  assign n39635 = n12140 | n12141;
  assign n39636 = n12142 | n12143;
  assign n39637 = n12149 | n12150;
  assign n39638 = n12163 | n12164;
  assign n39639 = n12174 | n12171 | n12173;
  assign n39640 = n12176 | n12177;
  assign n39641 = n12178 | n12179;
  assign n39642 = n12184 | n12185;
  assign n39643 = n12193 | n12194;
  assign n39644 = n12197 | n12198;
  assign n39645 = n12199 | n12200;
  assign n39646 = n12205 | ~n12206;
  assign n39647 = n12216 | n12217;
  assign n39648 = n12220 | n12221;
  assign n39649 = n12222 | n12223;
  assign n39650 = n12224 | ~n12225;
  assign n39651 = n12241 | n12242;
  assign n39652 = n12243 | n12244;
  assign n39653 = n12245 | ~n12246;
  assign n39654 = n12262 | n12263;
  assign n39655 = n12264 | n12265;
  assign n39656 = n12266 | ~n12267;
  assign n39657 = n12271 | n12272;
  assign n39658 = n12273 | n12274;
  assign n39659 = n12275 | ~n12276;
  assign n39660 = n12280 | n12281;
  assign n39661 = n12282 | n12283;
  assign n39662 = n12284 | ~n12285;
  assign n39663 = n12293 | n12294;
  assign n39664 = n12295 | n12296;
  assign n39665 = n12297 | ~n12298;
  assign n39666 = n12302 | n12303;
  assign n39667 = n12304 | n12305;
  assign n39668 = n12306 | ~n12307;
  assign n39669 = n12313 | n12314;
  assign n39670 = n12317 | n12318;
  assign n39671 = n12319 | n12320;
  assign n39672 = n12321 | ~n12322;
  assign n39673 = n12326 | n12327;
  assign n39674 = n12328 | n12329;
  assign n39675 = n12330 | ~n12331;
  assign n39676 = n12345 | n12346;
  assign n39677 = n12353 | n12354;
  assign n39678 = n12355 | n12356;
  assign n39679 = n12357 | ~n12358;
  assign n39680 = n12382 | n12383;
  assign n39681 = n12384 | n12385;
  assign n39682 = n12386 | ~n12387;
  assign n39683 = n12391 | n12392;
  assign n39684 = n12393 | n12394;
  assign n39685 = n12395 | ~n12396;
  assign n39686 = n12400 | n12401;
  assign n39687 = n12402 | n12403;
  assign n39688 = n12404 | ~n12405;
  assign n39689 = n12413 | n12414;
  assign n39690 = n12415 | n12416;
  assign n39691 = n12417 | ~n12418;
  assign n39692 = n12422 | n12423;
  assign n39693 = n12424 | n12425;
  assign n39694 = n12426 | ~n12427;
  assign n39695 = n12431 | n12432;
  assign n39696 = n12433 | n12434;
  assign n39697 = n12435 | ~n12436;
  assign n39698 = n12440 | n12441;
  assign n39699 = n12442 | n12443;
  assign n39700 = n12444 | ~n12445;
  assign n39701 = n12449 | n12450;
  assign n39702 = n12451 | n12452;
  assign n39703 = n12453 | ~n12454;
  assign n39704 = n12462 | n12463;
  assign n39705 = n12468 | n12469;
  assign n39706 = n12472 | n12473;
  assign n39707 = n12474 | n12475;
  assign n39708 = n12476 | ~n12477;
  assign n39709 = n12485 | n12486;
  assign n39710 = n12487 | n12488;
  assign n39711 = n12489 | ~n12490;
  assign n39712 = n12494 | n12495;
  assign n39713 = n12496 | n12497;
  assign n39714 = n12498 | ~n12499;
  assign n39715 = n12507 | n12508;
  assign n39716 = n12509 | n12510;
  assign n39717 = n12511 | ~n12512;
  assign n39718 = n12516 | n12517;
  assign n39719 = n12518 | n12519;
  assign n39720 = n12520 | ~n12521;
  assign n39721 = n12537 | n12538;
  assign n39722 = n12541 | n12542;
  assign n39723 = n12543 | n12544;
  assign n39724 = n12553 | n12554;
  assign n39725 = n12557 | n12558;
  assign n39726 = n12559 | n12560;
  assign n39727 = n12569 | n12570;
  assign n39728 = n12573 | n12574;
  assign n39729 = n12575 | n12576;
  assign n39730 = n12588 | n12589;
  assign n39731 = n12592 | n12593;
  assign n39732 = n12594 | n12595;
  assign n39733 = n12607 | n12608;
  assign n39734 = n12611 | n12612;
  assign n39735 = n12613 | n12614;
  assign n39736 = n12624 | n12625;
  assign n39737 = n12628 | n12629;
  assign n39738 = n12630 | n12631;
  assign n39739 = n12642 | n12643;
  assign n39740 = n12646 | n12647;
  assign n39741 = n12648 | n12649;
  assign n39742 = n12658 | n12659;
  assign n39743 = n12662 | n12663;
  assign n39744 = n12664 | n12665;
  assign n39745 = n12672 | ~n12673;
  assign n39746 = n12682 | ~n12683;
  assign n39747 = n12695 | n12696;
  assign n39748 = n12698 | n12699;
  assign n39749 = n12718 | n12719;
  assign n39750 = n12722 | n12723;
  assign n39751 = n12724 | n12725;
  assign n39752 = n12729 | n12730;
  assign n39753 = n12731 | n12732;
  assign n39754 = n12733 | ~n12734;
  assign n39755 = n12744 | n12745;
  assign n39756 = n12748 | n12749;
  assign n39757 = n12750 | n12751;
  assign n39758 = n12757 | n12758;
  assign n39759 = n12763 | ~n12764;
  assign n39760 = n12767 | n12768;
  assign n39761 = n12769 | n12770;
  assign n39762 = n12771 | ~n12772;
  assign n39763 = n12782 | n12783;
  assign n39764 = n12786 | n12787;
  assign n39765 = n12788 | n12789;
  assign n39766 = n12795 | n12796;
  assign n39767 = n12801 | ~n12802;
  assign n39768 = n12805 | n12806;
  assign n39769 = n12807 | n12808;
  assign n39770 = n12809 | ~n12810;
  assign n39771 = n12820 | n12821;
  assign n39772 = n12824 | n12825;
  assign n39773 = n12826 | n12827;
  assign n39774 = n12831 | n12832;
  assign n39775 = n12833 | n12834;
  assign n39776 = n12835 | ~n12836;
  assign n39777 = n12846 | n12847;
  assign n39778 = n12850 | n12851;
  assign n39779 = n12852 | n12853;
  assign n39780 = n12857 | n12858;
  assign n39781 = n12859 | n12860;
  assign n39782 = n12861 | ~n12862;
  assign n39783 = n12872 | n12873;
  assign n39784 = n12876 | n12877;
  assign n39785 = n12878 | n12879;
  assign n39786 = n12883 | n12884;
  assign n39787 = n12885 | n12886;
  assign n39788 = n12887 | ~n12888;
  assign n39789 = n12893 | ~n12894;
  assign n39790 = n12907 | n12908;
  assign n39791 = n12911 | n12912;
  assign n39792 = n12913 | n12914;
  assign n39793 = n12918 | n12919;
  assign n39794 = n12920 | n12921;
  assign n39795 = n12922 | ~n12923;
  assign n39796 = n12933 | n12934;
  assign n39797 = n12937 | n12938;
  assign n39798 = n12939 | n12940;
  assign n39799 = n12944 | n12945;
  assign n39800 = n12946 | n12947;
  assign n39801 = n12948 | ~n12949;
  assign n39802 = n12959 | n12960;
  assign n39803 = n12963 | n12964;
  assign n39804 = n12965 | n12966;
  assign n39805 = n12972 | n12973;
  assign n39806 = n12978 | ~n12979;
  assign n39807 = n13002 | ~n13003;
  assign n39808 = n13008 | ~n13009;
  assign n39809 = n13033 | ~n13034;
  assign n39810 = n13037 | n13038;
  assign n39811 = n13046 | n13047;
  assign n39812 = n13050 | n13051;
  assign n39813 = n13052 | n13053;
  assign n39814 = n13064 | n13065;
  assign n39815 = n13068 | n13069;
  assign n39816 = n13070 | n13071;
  assign n39817 = n13074 | n13075;
  assign n39818 = n13086 | n13087;
  assign n39819 = n13090 | n13091;
  assign n39820 = n13092 | n13093;
  assign n39821 = n13104 | n13105;
  assign n39822 = n13108 | n13109;
  assign n39823 = n13110 | n13111;
  assign n39824 = n13122 | n13123;
  assign n39825 = n13126 | n13127;
  assign n39826 = n13128 | n13129;
  assign n39827 = n13132 | n13133;
  assign n39828 = n13142 | n13143;
  assign n39829 = n13146 | n13147;
  assign n39830 = n13148 | n13149;
  assign n39831 = n13160 | n13161;
  assign n39832 = n13164 | n13165;
  assign n39833 = n13166 | n13167;
  assign n39834 = n13178 | n13179;
  assign n39835 = n13182 | n13183;
  assign n39836 = n13184 | n13185;
  assign n39837 = n13190 | ~n13191;
  assign n39838 = n13199 | n13200;
  assign n39839 = n13203 | n13204;
  assign n39840 = n13205 | n13206;
  assign n39841 = n13211 | ~n13212;
  assign n39842 = n13220 | n13221;
  assign n39843 = n13224 | n13225;
  assign n39844 = n13226 | n13227;
  assign n39845 = n13232 | ~n13233;
  assign n39846 = n13243 | n13244;
  assign n39847 = n13247 | n13248;
  assign n39848 = n13249 | n13250;
  assign n39849 = n13261 | n13262;
  assign n39850 = n13265 | n13266;
  assign n39851 = n13267 | n13268;
  assign n39852 = n13279 | n13280;
  assign n39853 = n13283 | n13284;
  assign n39854 = n13285 | n13286;
  assign n39855 = n13297 | n13298;
  assign n39856 = n13301 | n13302;
  assign n39857 = n13303 | n13304;
  assign n39858 = n13315 | n13316;
  assign n39859 = n13319 | n13320;
  assign n39860 = n13321 | n13322;
  assign n39861 = n13333 | n13334;
  assign n39862 = n13337 | n13338;
  assign n39863 = n13339 | n13340;
  assign n39864 = n13351 | n13352;
  assign n39865 = n13355 | n13356;
  assign n39866 = n13357 | n13358;
  assign n39867 = n13369 | n13370;
  assign n39868 = n13373 | n13374;
  assign n39869 = n13375 | n13376;
  assign n39870 = n13387 | n13388;
  assign n39871 = n13391 | n13392;
  assign n39872 = n13393 | n13394;
  assign n39873 = n13403 | n13404;
  assign n39874 = n13407 | n13408;
  assign n39875 = n13409 | n13410;
  assign n39876 = n13415 | ~n13416;
  assign n39877 = n13426 | n13427;
  assign n39878 = n13430 | n13431;
  assign n39879 = n13432 | n13433;
  assign n39880 = n13442 | n13443;
  assign n39881 = n13446 | n13447;
  assign n39882 = n13448 | n13449;
  assign n39883 = n13462 | n13463;
  assign n39884 = n13466 | n13467;
  assign n39885 = n13468 | n13469;
  assign n39886 = n13478 | n13479;
  assign n39887 = n13482 | n13483;
  assign n39888 = n13484 | n13485;
  assign n39889 = n13496 | n13497;
  assign n39890 = n13500 | n13501;
  assign n39891 = n13502 | n13503;
  assign n39892 = n13514 | n13515;
  assign n39893 = n13518 | n13519;
  assign n39894 = n13520 | n13521;
  assign n39895 = n13526 | ~n13527;
  assign n39896 = n13537 | n13538;
  assign n39897 = n13541 | n13542;
  assign n39898 = n13543 | n13544;
  assign n39899 = n13553 | n13554;
  assign n39900 = n13557 | n13558;
  assign n39901 = n13559 | n13560;
  assign n39902 = n13565 | ~n13566;
  assign n39903 = n13576 | n13577;
  assign n39904 = n13580 | n13581;
  assign n39905 = n13582 | n13583;
  assign n39906 = n13594 | n13595;
  assign n39907 = n13598 | n13599;
  assign n39908 = n13600 | n13601;
  assign n39909 = n13612 | n13613;
  assign n39910 = n13616 | n13617;
  assign n39911 = n13618 | n13619;
  assign n39912 = n13628 | n13629;
  assign n39913 = n13632 | n13633;
  assign n39914 = n13634 | n13635;
  assign n39915 = n13640 | ~n13641;
  assign n39916 = n13649 | n13650;
  assign n39917 = n13653 | n13654;
  assign n39918 = n13655 | n13656;
  assign n39919 = n13661 | ~n13662;
  assign n39920 = n13672 | n13673;
  assign n39921 = n13676 | n13677;
  assign n39922 = n13678 | n13679;
  assign n39923 = n13692 | n13693;
  assign n39924 = n13696 | n13697;
  assign n39925 = n13698 | n13699;
  assign n39926 = n13712 | n13713;
  assign n39927 = n13716 | n13717;
  assign n39928 = n13718 | n13719;
  assign n39929 = n13730 | n13731;
  assign n39930 = n13734 | n13735;
  assign n39931 = n13736 | n13737;
  assign n39932 = n13748 | n13749;
  assign n39933 = n13752 | n13753;
  assign n39934 = n13754 | n13755;
  assign n39935 = n13764 | n13765;
  assign n39936 = n13768 | n13769;
  assign n39937 = n13770 | n13771;
  assign n39938 = n13782 | n13783;
  assign n39939 = n13786 | n13787;
  assign n39940 = n13788 | n13789;
  assign n39941 = n13800 | n13801;
  assign n39942 = n13804 | n13805;
  assign n39943 = n13806 | n13807;
  assign n39944 = n13820 | n13821;
  assign n39945 = n13824 | n13825;
  assign n39946 = n13826 | n13827;
  assign n39947 = n13838 | n13839;
  assign n39948 = n13842 | n13843;
  assign n39949 = n13844 | n13845;
  assign n39950 = n13856 | n13857;
  assign n39951 = n13860 | n13861;
  assign n39952 = n13862 | n13863;
  assign n39953 = n13874 | n13875;
  assign n39954 = n13878 | n13879;
  assign n39955 = n13880 | n13881;
  assign n39956 = n13892 | n13893;
  assign n39957 = n13896 | n13897;
  assign n39958 = n13898 | n13899;
  assign n39959 = n13910 | n13911;
  assign n39960 = n13914 | n13915;
  assign n39961 = n13916 | n13917;
  assign n39962 = n13928 | n13929;
  assign n39963 = n13932 | n13933;
  assign n39964 = n13934 | n13935;
  assign n39965 = n13940 | ~n13941;
  assign n39966 = n13951 | n13952;
  assign n39967 = n13955 | n13956;
  assign n39968 = n13957 | n13958;
  assign n39969 = n13969 | n13970;
  assign n39970 = n13973 | n13974;
  assign n39971 = n13975 | n13976;
  assign n39972 = n13985 | n13986;
  assign n39973 = n13989 | n13990;
  assign n39974 = n13991 | n13992;
  assign n39975 = n13998 | n13999;
  assign n39976 = n14007 | n14008;
  assign n39977 = n14011 | n14012;
  assign n39978 = n14013 | n14014;
  assign n39979 = n14020 | n14021;
  assign n39980 = n14034 | n14035;
  assign n39981 = n14045 | n14042 | n14044;
  assign n39982 = n14047 | n14048;
  assign n39983 = n14049 | n14050;
  assign n39984 = n14055 | n14056;
  assign n39985 = n14064 | n14065;
  assign n39986 = n14068 | n14069;
  assign n39987 = n14070 | n14071;
  assign n39988 = n14076 | ~n14077;
  assign n39989 = n14085 | n14086;
  assign n39990 = n14087 | n14088;
  assign n39991 = n14089 | ~n14090;
  assign n39992 = n14094 | n14095;
  assign n39993 = n14096 | n14097;
  assign n39994 = n14098 | ~n14099;
  assign n39995 = n14103 | n14104;
  assign n39996 = n14105 | n14106;
  assign n39997 = n14107 | ~n14108;
  assign n39998 = n14116 | n14117;
  assign n39999 = n14118 | n14119;
  assign n40000 = n14120 | ~n14121;
  assign n40001 = n14139 | n14140;
  assign n40002 = n14141 | n14142;
  assign n40003 = n14143 | ~n14144;
  assign n40004 = n14156 | n14157;
  assign n40005 = n14158 | n14159;
  assign n40006 = n14160 | ~n14161;
  assign n40007 = n14169 | n14170;
  assign n40008 = n14171 | n14172;
  assign n40009 = n14173 | ~n14174;
  assign n40010 = n14178 | n14179;
  assign n40011 = n14180 | n14181;
  assign n40012 = n14182 | ~n14183;
  assign n40013 = n14191 | n14192;
  assign n40014 = n14193 | n14194;
  assign n40015 = n14195 | ~n14196;
  assign n40016 = n14204 | n14205;
  assign n40017 = n14206 | n14207;
  assign n40018 = n14208 | ~n14209;
  assign n40019 = n14213 | n14214;
  assign n40020 = n14215 | n14216;
  assign n40021 = n14217 | ~n14218;
  assign n40022 = n14222 | n14223;
  assign n40023 = n14224 | n14225;
  assign n40024 = n14226 | ~n14227;
  assign n40025 = n14231 | n14232;
  assign n40026 = n14233 | n14234;
  assign n40027 = n14235 | ~n14236;
  assign n40028 = n14240 | n14241;
  assign n40029 = n14242 | n14243;
  assign n40030 = n14244 | ~n14245;
  assign n40031 = n14261 | n14262;
  assign n40032 = n14263 | n14264;
  assign n40033 = n14265 | ~n14266;
  assign n40034 = n14274 | n14275;
  assign n40035 = n14276 | n14277;
  assign n40036 = n14278 | ~n14279;
  assign n40037 = n14289 | n14290;
  assign n40038 = n14293 | n14294;
  assign n40039 = n14295 | n14296;
  assign n40040 = n14297 | ~n14298;
  assign n40041 = n14302 | n14303;
  assign n40042 = n14304 | n14305;
  assign n40043 = n14306 | ~n14307;
  assign n40044 = n14313 | n14314;
  assign n40045 = n14319 | n14320;
  assign n40046 = n14323 | n14324;
  assign n40047 = n14325 | n14326;
  assign n40048 = n14327 | ~n14328;
  assign n40049 = n14332 | n14333;
  assign n40050 = n14334 | n14335;
  assign n40051 = n14336 | ~n14337;
  assign n40052 = n14343 | n14344;
  assign n40053 = n14347 | n14348;
  assign n40054 = n14349 | n14350;
  assign n40055 = n14351 | ~n14352;
  assign n40056 = n14356 | n14357;
  assign n40057 = n14358 | n14359;
  assign n40058 = n14360 | ~n14361;
  assign n40059 = n14365 | n14366;
  assign n40060 = n14367 | n14368;
  assign n40061 = n14369 | ~n14370;
  assign n40062 = n14374 | n14375;
  assign n40063 = n14376 | n14377;
  assign n40064 = n14378 | ~n14379;
  assign n40065 = n14387 | n14388;
  assign n40066 = n14389 | n14390;
  assign n40067 = n14391 | ~n14392;
  assign n40068 = n14396 | n14397;
  assign n40069 = n14398 | n14399;
  assign n40070 = n14400 | ~n14401;
  assign n40071 = n14409 | n14410;
  assign n40072 = n14411 | n14412;
  assign n40073 = n14413 | ~n14414;
  assign n40074 = n14422 | n14423;
  assign n40075 = n14424 | n14425;
  assign n40076 = n14426 | ~n14427;
  assign n40077 = n14437 | n14438;
  assign n40078 = n14441 | n14442;
  assign n40079 = n14443 | n14444;
  assign n40080 = n14454 | n14455;
  assign n40081 = n14458 | n14459;
  assign n40082 = n14460 | n14461;
  assign n40083 = n14469 | n14470;
  assign n40084 = n14473 | n14474;
  assign n40085 = n14475 | n14476;
  assign n40086 = n14487 | n14488;
  assign n40087 = n14491 | n14492;
  assign n40088 = n14493 | n14494;
  assign n40089 = n14506 | n14507;
  assign n40090 = n14510 | n14511;
  assign n40091 = n14512 | n14513;
  assign n40092 = n14521 | n14522;
  assign n40093 = n14525 | n14526;
  assign n40094 = n14527 | n14528;
  assign n40095 = n14537 | n14538;
  assign n40096 = n14541 | n14542;
  assign n40097 = n14543 | n14544;
  assign n40098 = n14553 | n14554;
  assign n40099 = n14557 | n14558;
  assign n40100 = n14559 | n14560;
  assign n40101 = n14569 | n14570;
  assign n40102 = n14573 | n14574;
  assign n40103 = n14575 | n14576;
  assign n40104 = n14585 | n14586;
  assign n40105 = n14589 | n14590;
  assign n40106 = n14591 | n14592;
  assign n40107 = n14597 | n14598;
  assign n40108 = n14608 | n14605 | n14607;
  assign n40109 = n14610 | n14611;
  assign n40110 = n14612 | n14613;
  assign n40111 = n14620 | n14621;
  assign n40112 = n14623 | n14624;
  assign n40113 = n14629 | n14630;
  assign n40114 = n14635 | ~n14636;
  assign n40115 = n14655 | n14656;
  assign n40116 = n14659 | n14660;
  assign n40117 = n14661 | n14662;
  assign n40118 = n14666 | n14667;
  assign n40119 = n14668 | n14669;
  assign n40120 = n14670 | ~n14671;
  assign n40121 = n14677 | n14678;
  assign n40122 = n14679 | n14680;
  assign n40123 = n14681 | ~n14682;
  assign n40124 = n14685 | n14686;
  assign n40125 = n14687 | n14688;
  assign n40126 = n14689 | ~n14690;
  assign n40127 = n14695 | ~n14696;
  assign n40128 = n14701 | ~n14702;
  assign n40129 = n14715 | n14716;
  assign n40130 = n14719 | n14720;
  assign n40131 = n14721 | n14722;
  assign n40132 = n14726 | n14727;
  assign n40133 = n14728 | n14729;
  assign n40134 = n14730 | ~n14731;
  assign n40135 = n14741 | n14742;
  assign n40136 = n14745 | n14746;
  assign n40137 = n14747 | n14748;
  assign n40138 = n14752 | n14753;
  assign n40139 = n14754 | n14755;
  assign n40140 = n14756 | ~n14757;
  assign n40141 = n14767 | n14768;
  assign n40142 = n14771 | n14772;
  assign n40143 = n14773 | n14774;
  assign n40144 = n14780 | n14781;
  assign n40145 = n14786 | ~n14787;
  assign n40146 = n14790 | n14791;
  assign n40147 = n14792 | n14793;
  assign n40148 = n14794 | ~n14795;
  assign n40149 = n14805 | n14806;
  assign n40150 = n14809 | n14810;
  assign n40151 = n14811 | n14812;
  assign n40152 = n14816 | n14817;
  assign n40153 = n14818 | n14819;
  assign n40154 = n14820 | ~n14821;
  assign n40155 = n14831 | n14832;
  assign n40156 = n14835 | n14836;
  assign n40157 = n14837 | n14838;
  assign n40158 = n14844 | n14845;
  assign n40159 = n14850 | ~n14851;
  assign n40160 = n14854 | n14855;
  assign n40161 = n14856 | n14857;
  assign n40162 = n14858 | ~n14859;
  assign n40163 = n14864 | ~n14865;
  assign n40164 = n14878 | n14879;
  assign n40165 = n14882 | n14883;
  assign n40166 = n14884 | n14885;
  assign n40167 = n14889 | n14890;
  assign n40168 = n14891 | n14892;
  assign n40169 = n14893 | ~n14894;
  assign n40170 = n14899 | ~n14900;
  assign n40171 = n14920 | n14921;
  assign n40172 = n14924 | n14925;
  assign n40173 = n14926 | n14927;
  assign n40174 = n14936 | ~n14937;
  assign n40175 = n14942 | ~n14943;
  assign n40176 = n14967 | ~n14968;
  assign n40177 = n14971 | n14972;
  assign n40178 = n14980 | n14981;
  assign n40179 = n14984 | n14985;
  assign n40180 = n14986 | n14987;
  assign n40181 = n14993 | ~n14994;
  assign n40182 = n15002 | ~n15003;
  assign n40183 = n15027 | n15028;
  assign n40184 = n15034 | n15035;
  assign n40185 = n15038 | n15039;
  assign n40186 = n15040 | n15041;
  assign n40187 = n15056 | n15057;
  assign n40188 = n15060 | n15061;
  assign n40189 = n15062 | n15063;
  assign n40190 = n15075 | n15076;
  assign n40191 = n15079 | n15080;
  assign n40192 = n15081 | n15082;
  assign n40193 = n15087 | n15088;
  assign n40194 = n15098 | n15099;
  assign n40195 = n15102 | n15103;
  assign n40196 = n15104 | n15105;
  assign n40197 = n15118 | n15119;
  assign n40198 = n15122 | n15123;
  assign n40199 = n15124 | n15125;
  assign n40200 = n15134 | ~n15135;
  assign n40201 = n15147 | n15148;
  assign n40202 = n15151 | n15152;
  assign n40203 = n15153 | n15154;
  assign n40204 = n15157 | n15158;
  assign n40205 = n15159 | n15160;
  assign n40206 = n15161 | ~n15162;
  assign n40207 = n15170 | n15171;
  assign n40208 = n15174 | n15175;
  assign n40209 = n15176 | n15177;
  assign n40210 = n15183 | ~n15184;
  assign n40211 = n15186 | ~n15187;
  assign n40212 = n15195 | n15196;
  assign n40213 = n15199 | n15200;
  assign n40214 = n15201 | n15202;
  assign n40215 = n15213 | n15214;
  assign n40216 = n15217 | n15218;
  assign n40217 = n15219 | n15220;
  assign n40218 = n15223 | n15224;
  assign n40219 = n15233 | n15234;
  assign n40220 = n15237 | n15238;
  assign n40221 = n15239 | n15240;
  assign n40222 = n15243 | n15244;
  assign n40223 = n15245 | n15246;
  assign n40224 = n15247 | ~n15248;
  assign n40225 = n15258 | n15259;
  assign n40226 = n15262 | n15263;
  assign n40227 = n15264 | n15265;
  assign n40228 = n15276 | n15277;
  assign n40229 = n15280 | n15281;
  assign n40230 = n15282 | n15283;
  assign n40231 = n15294 | n15295;
  assign n40232 = n15298 | n15299;
  assign n40233 = n15300 | n15301;
  assign n40234 = n15312 | n15313;
  assign n40235 = n15316 | n15317;
  assign n40236 = n15318 | n15319;
  assign n40237 = n15328 | n15329;
  assign n40238 = n15332 | n15333;
  assign n40239 = n15334 | n15335;
  assign n40240 = n15340 | ~n15341;
  assign n40241 = n15349 | n15350;
  assign n40242 = n15353 | n15354;
  assign n40243 = n15355 | n15356;
  assign n40244 = n15361 | ~n15362;
  assign n40245 = n15372 | n15373;
  assign n40246 = n15376 | n15377;
  assign n40247 = n15378 | n15379;
  assign n40248 = n15388 | n15389;
  assign n40249 = n15392 | n15393;
  assign n40250 = n15394 | n15395;
  assign n40251 = n15400 | ~n15401;
  assign n40252 = n15409 | n15410;
  assign n40253 = n15413 | n15414;
  assign n40254 = n15415 | n15416;
  assign n40255 = n15421 | ~n15422;
  assign n40256 = n15430 | n15431;
  assign n40257 = n15434 | n15435;
  assign n40258 = n15436 | n15437;
  assign n40259 = n15442 | ~n15443;
  assign n40260 = n15453 | n15454;
  assign n40261 = n15457 | n15458;
  assign n40262 = n15459 | n15460;
  assign n40263 = n15469 | n15470;
  assign n40264 = n15473 | n15474;
  assign n40265 = n15475 | n15476;
  assign n40266 = n15487 | n15488;
  assign n40267 = n15491 | n15492;
  assign n40268 = n15493 | n15494;
  assign n40269 = n15499 | ~n15500;
  assign n40270 = n15508 | n15509;
  assign n40271 = n15512 | n15513;
  assign n40272 = n15514 | n15515;
  assign n40273 = n15526 | n15527;
  assign n40274 = n15530 | n15531;
  assign n40275 = n15532 | n15533;
  assign n40276 = n15538 | ~n15539;
  assign n40277 = n15549 | n15550;
  assign n40278 = n15553 | n15554;
  assign n40279 = n15555 | n15556;
  assign n40280 = n15565 | n15566;
  assign n40281 = n15569 | n15570;
  assign n40282 = n15571 | n15572;
  assign n40283 = n15577 | ~n15578;
  assign n40284 = n15586 | n15587;
  assign n40285 = n15590 | n15591;
  assign n40286 = n15592 | n15593;
  assign n40287 = n15606 | n15607;
  assign n40288 = n15610 | n15611;
  assign n40289 = n15612 | n15613;
  assign n40290 = n15622 | n15623;
  assign n40291 = n15626 | n15627;
  assign n40292 = n15628 | n15629;
  assign n40293 = n15642 | n15643;
  assign n40294 = n15646 | n15647;
  assign n40295 = n15648 | n15649;
  assign n40296 = n15660 | n15661;
  assign n40297 = n15664 | n15665;
  assign n40298 = n15666 | n15667;
  assign n40299 = n15678 | n15679;
  assign n40300 = n15682 | n15683;
  assign n40301 = n15684 | n15685;
  assign n40302 = n15696 | n15697;
  assign n40303 = n15700 | n15701;
  assign n40304 = n15702 | n15703;
  assign n40305 = n15714 | n15715;
  assign n40306 = n15718 | n15719;
  assign n40307 = n15720 | n15721;
  assign n40308 = n15732 | n15733;
  assign n40309 = n15736 | n15737;
  assign n40310 = n15738 | n15739;
  assign n40311 = n15748 | n15749;
  assign n40312 = n15752 | n15753;
  assign n40313 = n15754 | n15755;
  assign n40314 = n15768 | n15769;
  assign n40315 = n15772 | n15773;
  assign n40316 = n15774 | n15775;
  assign n40317 = n15786 | n15787;
  assign n40318 = n15790 | n15791;
  assign n40319 = n15792 | n15793;
  assign n40320 = n15804 | n15805;
  assign n40321 = n15808 | n15809;
  assign n40322 = n15810 | n15811;
  assign n40323 = n15820 | n15821;
  assign n40324 = n15824 | n15825;
  assign n40325 = n15826 | n15827;
  assign n40326 = n15830 | n15831;
  assign n40327 = n15832 | n15833;
  assign n40328 = n15834 | ~n15835;
  assign n40329 = n15843 | n15844;
  assign n40330 = n15847 | n15848;
  assign n40331 = n15849 | n15850;
  assign n40332 = n15861 | n15862;
  assign n40333 = n15865 | n15866;
  assign n40334 = n15867 | n15868;
  assign n40335 = n15871 | n15872;
  assign n40336 = n15873 | n15874;
  assign n40337 = n15875 | ~n15876;
  assign n40338 = n15886 | n15887;
  assign n40339 = n15890 | n15891;
  assign n40340 = n15892 | n15893;
  assign n40341 = n15904 | n15905;
  assign n40342 = n15908 | n15909;
  assign n40343 = n15910 | n15911;
  assign n40344 = n15920 | n15921;
  assign n40345 = n15924 | n15925;
  assign n40346 = n15926 | n15927;
  assign n40347 = n15940 | n15941;
  assign n40348 = n15944 | n15945;
  assign n40349 = n15946 | n15947;
  assign n40350 = n15956 | n15957;
  assign n40351 = n15960 | n15961;
  assign n40352 = n15962 | n15963;
  assign n40353 = n15974 | n15975;
  assign n40354 = n15978 | n15979;
  assign n40355 = n15980 | n15981;
  assign n40356 = n15992 | n15993;
  assign n40357 = n15996 | n15997;
  assign n40358 = n15998 | n15999;
  assign n40359 = n16010 | n16011;
  assign n40360 = n16014 | n16015;
  assign n40361 = n16016 | n16017;
  assign n40362 = n16020 | n16021;
  assign n40363 = n16030 | n16031;
  assign n40364 = n16034 | n16035;
  assign n40365 = n16036 | n16037;
  assign n40366 = n16050 | n16051;
  assign n40367 = n16054 | n16055;
  assign n40368 = n16056 | n16057;
  assign n40369 = n16068 | n16069;
  assign n40370 = n16072 | n16073;
  assign n40371 = n16074 | n16075;
  assign n40372 = n16086 | n16087;
  assign n40373 = n16090 | n16091;
  assign n40374 = n16092 | n16093;
  assign n40375 = n16106 | n16107;
  assign n40376 = n16110 | n16111;
  assign n40377 = n16112 | n16113;
  assign n40378 = n16124 | n16125;
  assign n40379 = n16128 | n16129;
  assign n40380 = n16130 | n16131;
  assign n40381 = n16140 | n16141;
  assign n40382 = n16144 | n16145;
  assign n40383 = n16146 | n16147;
  assign n40384 = n16153 | n16154;
  assign n40385 = n16162 | n16163;
  assign n40386 = n16166 | n16167;
  assign n40387 = n16168 | n16169;
  assign n40388 = n16175 | n16176;
  assign n40389 = n16189 | n16190;
  assign n40390 = n16197 | n16198;
  assign n40391 = n16200 | n16201;
  assign n40392 = n16206 | n16202 | ~n16205;
  assign n40393 = n16210 | n16211;
  assign n40394 = n16219 | n16220;
  assign n40395 = n16223 | n16224;
  assign n40396 = n16225 | n16226;
  assign n40397 = n16229 | n16230;
  assign n40398 = n16231 | n16232;
  assign n40399 = n16233 | ~n16234;
  assign n40400 = n16238 | n16239;
  assign n40401 = n16240 | n16241;
  assign n40402 = n16242 | ~n16243;
  assign n40403 = n16247 | n16248;
  assign n40404 = n16249 | n16250;
  assign n40405 = n16251 | ~n16252;
  assign n40406 = n16256 | n16257;
  assign n40407 = n16258 | n16259;
  assign n40408 = n16260 | ~n16261;
  assign n40409 = n16265 | n16266;
  assign n40410 = n16267 | n16268;
  assign n40411 = n16269 | ~n16270;
  assign n40412 = n16274 | n16275;
  assign n40413 = n16276 | n16277;
  assign n40414 = n16278 | ~n16279;
  assign n40415 = n16287 | n16288;
  assign n40416 = n16295 | n16296;
  assign n40417 = n16297 | n16298;
  assign n40418 = n16299 | ~n16300;
  assign n40419 = n16316 | n16317;
  assign n40420 = n16318 | n16319;
  assign n40421 = n16320 | ~n16321;
  assign n40422 = n16325 | n16326;
  assign n40423 = n16327 | n16328;
  assign n40424 = n16329 | ~n16330;
  assign n40425 = n16334 | n16335;
  assign n40426 = n16336 | n16337;
  assign n40427 = n16338 | ~n16339;
  assign n40428 = n16343 | n16344;
  assign n40429 = n16345 | n16346;
  assign n40430 = n16347 | ~n16348;
  assign n40431 = n16354 | ~n16355;
  assign n40432 = n16359 | n16360;
  assign n40433 = n16361 | n16362;
  assign n40434 = n16363 | ~n16364;
  assign n40435 = n16370 | ~n16371;
  assign n40436 = n16375 | n16376;
  assign n40437 = n16377 | n16378;
  assign n40438 = n16379 | ~n16380;
  assign n40439 = n16384 | n16385;
  assign n40440 = n16386 | n16387;
  assign n40441 = n16388 | ~n16389;
  assign n40442 = n16393 | n16394;
  assign n40443 = n16395 | n16396;
  assign n40444 = n16397 | ~n16398;
  assign n40445 = n16402 | n16403;
  assign n40446 = n16404 | n16405;
  assign n40447 = n16406 | ~n16407;
  assign n40448 = n16411 | n16412;
  assign n40449 = n16413 | n16414;
  assign n40450 = n16415 | ~n16416;
  assign n40451 = n16420 | n16421;
  assign n40452 = n16422 | n16423;
  assign n40453 = n16424 | ~n16425;
  assign n40454 = n16431 | n16432;
  assign n40455 = n16435 | n16436;
  assign n40456 = n16437 | n16438;
  assign n40457 = n16439 | ~n16440;
  assign n40458 = n16446 | n16447;
  assign n40459 = n16452 | n16453;
  assign n40460 = n16460 | n16461;
  assign n40461 = n16462 | n16463;
  assign n40462 = n16464 | ~n16465;
  assign n40463 = n16477 | n16478;
  assign n40464 = n16479 | n16480;
  assign n40465 = n16481 | ~n16482;
  assign n40466 = n16490 | n16491;
  assign n40467 = n16492 | n16493;
  assign n40468 = n16494 | ~n16495;
  assign n40469 = n16503 | n16504;
  assign n40470 = n16505 | n16506;
  assign n40471 = n16507 | ~n16508;
  assign n40472 = n16512 | n16513;
  assign n40473 = n16514 | n16515;
  assign n40474 = n16516 | ~n16517;
  assign n40475 = n16521 | n16522;
  assign n40476 = n16523 | n16524;
  assign n40477 = n16525 | ~n16526;
  assign n40478 = n16538 | n16539;
  assign n40479 = n16540 | n16541;
  assign n40480 = n16542 | ~n16543;
  assign n40481 = n16547 | n16548;
  assign n40482 = n16549 | n16550;
  assign n40483 = n16551 | ~n16552;
  assign n40484 = n16560 | n16561;
  assign n40485 = n16562 | n16563;
  assign n40486 = n16564 | ~n16565;
  assign n40487 = n16571 | n16572;
  assign n40488 = n16579 | n16580;
  assign n40489 = n16581 | n16582;
  assign n40490 = n16583 | ~n16584;
  assign n40491 = n16592 | n16593;
  assign n40492 = n16594 | n16595;
  assign n40493 = n16596 | ~n16597;
  assign n40494 = n16607 | ~n16608;
  assign n40495 = n16618 | n16619;
  assign n40496 = n16622 | n16623;
  assign n40497 = n16624 | n16625;
  assign n40498 = n16634 | n16635;
  assign n40499 = n16638 | n16639;
  assign n40500 = n16640 | n16641;
  assign n40501 = n16644 | n16645;
  assign n40502 = n16646 | n16647;
  assign n40503 = n16648 | ~n16649;
  assign n40504 = n16659 | n16660;
  assign n40505 = n16663 | n16664;
  assign n40506 = n16665 | n16666;
  assign n40507 = n16675 | n16676;
  assign n40508 = n16679 | n16680;
  assign n40509 = n16681 | n16682;
  assign n40510 = n16687 | ~n16688;
  assign n40511 = n16696 | n16697;
  assign n40512 = n16700 | n16701;
  assign n40513 = n16702 | n16703;
  assign n40514 = n16714 | n16715;
  assign n40515 = n16718 | n16719;
  assign n40516 = n16720 | n16721;
  assign n40517 = n16726 | ~n16727;
  assign n40518 = n16735 | n16736;
  assign n40519 = n16739 | n16740;
  assign n40520 = n16741 | n16742;
  assign n40521 = n16747 | ~n16748;
  assign n40522 = n16756 | n16757;
  assign n40523 = n16760 | n16761;
  assign n40524 = n16762 | n16763;
  assign n40525 = n16776 | n16777;
  assign n40526 = n16780 | n16781;
  assign n40527 = n16782 | n16783;
  assign n40528 = n16794 | n16795;
  assign n40529 = n16798 | n16799;
  assign n40530 = n16800 | n16801;
  assign n40531 = n16810 | n16811;
  assign n40532 = n16814 | n16815;
  assign n40533 = n16816 | n16817;
  assign n40534 = n16830 | n16831;
  assign n40535 = n16834 | n16835;
  assign n40536 = n16836 | n16837;
  assign n40537 = n16848 | n16849;
  assign n40538 = n16852 | n16853;
  assign n40539 = n16854 | n16855;
  assign n40540 = n16866 | n16867;
  assign n40541 = n16870 | n16871;
  assign n40542 = n16872 | n16873;
  assign n40543 = n16882 | n16883;
  assign n40544 = n16886 | n16887;
  assign n40545 = n16888 | n16889;
  assign n40546 = n16892 | n16893;
  assign n40547 = n16894 | n16895;
  assign n40548 = n16896 | ~n16897;
  assign n40549 = n16907 | n16908;
  assign n40550 = n16911 | n16912;
  assign n40551 = n16913 | n16914;
  assign n40552 = n16923 | n16924;
  assign n40553 = n16927 | n16928;
  assign n40554 = n16929 | n16930;
  assign n40555 = n16935 | ~n16936;
  assign n40556 = n16946 | n16947;
  assign n40557 = n16950 | n16951;
  assign n40558 = n16952 | n16953;
  assign n40559 = n16962 | n16963;
  assign n40560 = n16966 | n16967;
  assign n40561 = n16968 | n16969;
  assign n40562 = n16974 | ~n16975;
  assign n40563 = n16985 | n16986;
  assign n40564 = n16989 | n16990;
  assign n40565 = n16991 | n16992;
  assign n40566 = n17003 | n17004;
  assign n40567 = n17007 | n17008;
  assign n40568 = n17009 | n17010;
  assign n40569 = n17021 | n17022;
  assign n40570 = n17025 | n17026;
  assign n40571 = n17027 | n17028;
  assign n40572 = n17039 | n17040;
  assign n40573 = n17043 | n17044;
  assign n40574 = n17045 | n17046;
  assign n40575 = n17055 | n17056;
  assign n40576 = n17059 | n17060;
  assign n40577 = n17061 | n17062;
  assign n40578 = n17067 | ~n17068;
  assign n40579 = n17076 | n17077;
  assign n40580 = n17080 | n17081;
  assign n40581 = n17082 | n17083;
  assign n40582 = n17088 | ~n17089;
  assign n40583 = n17097 | n17098;
  assign n40584 = n17101 | n17102;
  assign n40585 = n17103 | n17104;
  assign n40586 = n17109 | ~n17110;
  assign n40587 = n17118 | n17119;
  assign n40588 = n17122 | n17123;
  assign n40589 = n17124 | n17125;
  assign n40590 = n17130 | ~n17131;
  assign n40591 = n17141 | n17142;
  assign n40592 = n17145 | n17146;
  assign n40593 = n17147 | n17148;
  assign n40594 = n17159 | n17160;
  assign n40595 = n17163 | n17164;
  assign n40596 = n17165 | n17166;
  assign n40597 = n17175 | n17176;
  assign n40598 = n17179 | n17180;
  assign n40599 = n17181 | n17182;
  assign n40600 = n17185 | n17186;
  assign n40601 = n17187 | n17188;
  assign n40602 = n17189 | ~n17190;
  assign n40603 = n17200 | n17201;
  assign n40604 = n17204 | n17205;
  assign n40605 = n17206 | n17207;
  assign n40606 = n17218 | n17219;
  assign n40607 = n17222 | n17223;
  assign n40608 = n17224 | n17225;
  assign n40609 = n17234 | n17235;
  assign n40610 = n17238 | n17239;
  assign n40611 = n17240 | n17241;
  assign n40612 = n17246 | ~n17247;
  assign n40613 = n17255 | n17256;
  assign n40614 = n17259 | n17260;
  assign n40615 = n17261 | n17262;
  assign n40616 = n17273 | n17274;
  assign n40617 = n17277 | n17278;
  assign n40618 = n17279 | n17280;
  assign n40619 = n17285 | ~n17286;
  assign n40620 = n17296 | n17297;
  assign n40621 = n17300 | n17301;
  assign n40622 = n17302 | n17303;
  assign n40623 = n17314 | n17315;
  assign n40624 = n17318 | n17319;
  assign n40625 = n17320 | n17321;
  assign n40626 = n17332 | n17333;
  assign n40627 = n17336 | n17337;
  assign n40628 = n17338 | n17339;
  assign n40629 = n17348 | n17349;
  assign n40630 = n17352 | n17353;
  assign n40631 = n17354 | n17355;
  assign n40632 = n17358 | n17359;
  assign n40633 = n17360 | n17361;
  assign n40634 = n17362 | ~n17363;
  assign n40635 = n17373 | n17374;
  assign n40636 = n17377 | n17378;
  assign n40637 = n17379 | n17380;
  assign n40638 = n17391 | n17392;
  assign n40639 = n17395 | n17396;
  assign n40640 = n17397 | n17398;
  assign n40641 = n17409 | n17410;
  assign n40642 = n17413 | n17414;
  assign n40643 = n17415 | n17416;
  assign n40644 = n17425 | n17426;
  assign n40645 = n17429 | n17430;
  assign n40646 = n17431 | n17432;
  assign n40647 = n17443 | n17444;
  assign n40648 = n17447 | n17448;
  assign n40649 = n17449 | n17450;
  assign n40650 = n17453 | n17454;
  assign n40651 = n17463 | n17464;
  assign n40652 = n17467 | n17468;
  assign n40653 = n17469 | n17470;
  assign n40654 = n17481 | n17482;
  assign n40655 = n17485 | n17486;
  assign n40656 = n17487 | n17488;
  assign n40657 = n17493 | ~n17494;
  assign n40658 = n17504 | n17505;
  assign n40659 = n17508 | n17509;
  assign n40660 = n17510 | n17511;
  assign n40661 = n17520 | n17521;
  assign n40662 = n17524 | n17525;
  assign n40663 = n17526 | n17527;
  assign n40664 = n17530 | n17531;
  assign n40665 = n17532 | n17533;
  assign n40666 = n17534 | ~n17535;
  assign n40667 = n17545 | n17546;
  assign n40668 = n17549 | n17550;
  assign n40669 = n17551 | n17552;
  assign n40670 = n17563 | n17564;
  assign n40671 = n17567 | n17568;
  assign n40672 = n17569 | n17570;
  assign n40673 = n17581 | n17582;
  assign n40674 = n17585 | n17586;
  assign n40675 = n17587 | n17588;
  assign n40676 = n17597 | n17598;
  assign n40677 = n17601 | n17602;
  assign n40678 = n17603 | n17604;
  assign n40679 = n17615 | n17616;
  assign n40680 = n17619 | n17620;
  assign n40681 = n17621 | n17622;
  assign n40682 = n17627 | ~n17628;
  assign n40683 = n17636 | n17637;
  assign n40684 = n17640 | n17641;
  assign n40685 = n17642 | n17643;
  assign n40686 = n17649 | n17650;
  assign n40687 = n17658 | n17659;
  assign n40688 = n17662 | n17663;
  assign n40689 = n17664 | n17665;
  assign n40690 = n17671 | n17672;
  assign n40691 = n17680 | n17681;
  assign n40692 = n17684 | n17685;
  assign n40693 = n17686 | n17687;
  assign n40694 = n17703 | n17704;
  assign n40695 = n17712 | n17713;
  assign n40696 = n17714 | n17715;
  assign n40697 = n17720 | n17721;
  assign n40698 = n17725 | n17726;
  assign n40699 = n17727 | n17728;
  assign n40700 = n17729 | ~n17730;
  assign n40701 = n17734 | n17735;
  assign n40702 = n17736 | n17737;
  assign n40703 = n17738 | ~n17739;
  assign n40704 = n17751 | n17752;
  assign n40705 = n17753 | n17754;
  assign n40706 = n17755 | ~n17756;
  assign n40707 = n17760 | n17761;
  assign n40708 = n17762 | n17763;
  assign n40709 = n17764 | ~n17765;
  assign n40710 = n17775 | ~n17776;
  assign n40711 = n17780 | n17781;
  assign n40712 = n17782 | n17783;
  assign n40713 = n17784 | ~n17785;
  assign n40714 = n17791 | ~n17792;
  assign n40715 = n17798 | ~n17799;
  assign n40716 = n17803 | n17804;
  assign n40717 = n17805 | n17806;
  assign n40718 = n17807 | ~n17808;
  assign n40719 = n17814 | ~n17815;
  assign n40720 = n17819 | n17820;
  assign n40721 = n17821 | n17822;
  assign n40722 = n17823 | ~n17824;
  assign n40723 = n17828 | n17829;
  assign n40724 = n17830 | n17831;
  assign n40725 = n17832 | ~n17833;
  assign n40726 = n17837 | n17838;
  assign n40727 = n17839 | n17840;
  assign n40728 = n17841 | ~n17842;
  assign n40729 = n17848 | ~n17849;
  assign n40730 = n17853 | n17854;
  assign n40731 = n17855 | n17856;
  assign n40732 = n17857 | ~n17858;
  assign n40733 = n17866 | n17867;
  assign n40734 = n17868 | n17869;
  assign n40735 = n17870 | ~n17871;
  assign n40736 = n17875 | n17876;
  assign n40737 = n17877 | n17878;
  assign n40738 = n17879 | ~n17880;
  assign n40739 = n17902 | ~n17903;
  assign n40740 = n17907 | n17908;
  assign n40741 = n17909 | n17910;
  assign n40742 = n17911 | ~n17912;
  assign n40743 = n17916 | n17917;
  assign n40744 = n17918 | n17919;
  assign n40745 = n17920 | ~n17921;
  assign n40746 = n17927 | ~n17928;
  assign n40747 = n17938 | ~n17939;
  assign n40748 = n17945 | ~n17946;
  assign n40749 = n17950 | n17951;
  assign n40750 = n17952 | n17953;
  assign n40751 = n17954 | ~n17955;
  assign n40752 = n17963 | n17964;
  assign n40753 = n17965 | n17966;
  assign n40754 = n17967 | ~n17968;
  assign n40755 = n17972 | n17973;
  assign n40756 = n17974 | n17975;
  assign n40757 = n17976 | ~n17977;
  assign n40758 = n17989 | n17990;
  assign n40759 = n17991 | n17992;
  assign n40760 = n17993 | ~n17994;
  assign n40761 = n17998 | n17999;
  assign n40762 = n18000 | n18001;
  assign n40763 = n18002 | ~n18003;
  assign n40764 = n18009 | ~n18010;
  assign n40765 = n18018 | n18019;
  assign n40766 = n18020 | n18021;
  assign n40767 = n18022 | ~n18023;
  assign n40768 = n18027 | n18028;
  assign n40769 = n18029 | n18030;
  assign n40770 = n18031 | ~n18032;
  assign n40771 = n18044 | n18045;
  assign n40772 = n18046 | n18047;
  assign n40773 = n18048 | ~n18049;
  assign n40774 = n18063 | ~n18064;
  assign n40775 = n18076 | n18077;
  assign n40776 = n18078 | n18079;
  assign n40777 = n18080 | ~n18081;
  assign n40778 = n18087 | ~n18088;
  assign n40779 = n18092 | n18093;
  assign n40780 = n18094 | n18095;
  assign n40781 = n18096 | ~n18097;
  assign n40782 = n18103 | ~n18104;
  assign n40783 = n18119 | n18120;
  assign n40784 = n18127 | n18128;
  assign n40785 = n18131 | n18132;
  assign n40786 = n18133 | n18134;
  assign n40787 = n18144 | n18145;
  assign n40788 = n18148 | n18149;
  assign n40789 = n18150 | n18151;
  assign n40790 = n18160 | n18161;
  assign n40791 = n18164 | n18165;
  assign n40792 = n18166 | n18167;
  assign n40793 = n18176 | n18177;
  assign n40794 = n18180 | n18181;
  assign n40795 = n18182 | n18183;
  assign n40796 = n18191 | n18192;
  assign n40797 = n18195 | n18196;
  assign n40798 = n18197 | n18198;
  assign n40799 = n18208 | n18209;
  assign n40800 = n18212 | n18213;
  assign n40801 = n18214 | n18215;
  assign n40802 = n18226 | n18227;
  assign n40803 = n18230 | n18231;
  assign n40804 = n18232 | n18233;
  assign n40805 = n18244 | n18245;
  assign n40806 = n18248 | n18249;
  assign n40807 = n18250 | n18251;
  assign n40808 = n18260 | n18261;
  assign n40809 = n18264 | n18265;
  assign n40810 = n18266 | n18267;
  assign n40811 = n18275 | n18276;
  assign n40812 = n18279 | n18280;
  assign n40813 = n18281 | n18282;
  assign n40814 = n18288 | ~n18289;
  assign n40815 = n18293 | n18294;
  assign n40816 = n18295 | n18296;
  assign n40817 = n18297 | ~n18298;
  assign n40818 = n18303 | ~n18304;
  assign n40819 = n18317 | n18318;
  assign n40820 = n18321 | n18322;
  assign n40821 = n18323 | n18324;
  assign n40822 = n18328 | n18329;
  assign n40823 = n18330 | n18331;
  assign n40824 = n18332 | ~n18333;
  assign n40825 = n18338 | ~n18339;
  assign n40826 = n18352 | n18353;
  assign n40827 = n18356 | n18357;
  assign n40828 = n18358 | n18359;
  assign n40829 = n18363 | n18364;
  assign n40830 = n18365 | n18366;
  assign n40831 = n18367 | ~n18368;
  assign n40832 = n18378 | n18379;
  assign n40833 = n18382 | n18383;
  assign n40834 = n18384 | n18385;
  assign n40835 = n18405 | n18406;
  assign n40836 = n18409 | n18410;
  assign n40837 = n18411 | n18412;
  assign n40838 = n18416 | n18417;
  assign n40839 = n18418 | n18419;
  assign n40840 = n18420 | ~n18421;
  assign n40841 = n18431 | n18432;
  assign n40842 = n18435 | n18436;
  assign n40843 = n18437 | n18438;
  assign n40844 = n18442 | n18443;
  assign n40845 = n18444 | n18445;
  assign n40846 = n18446 | ~n18447;
  assign n40847 = n18457 | n18458;
  assign n40848 = n18461 | n18462;
  assign n40849 = n18463 | n18464;
  assign n40850 = n18479 | n18480;
  assign n40851 = n18483 | n18484;
  assign n40852 = n18485 | n18486;
  assign n40853 = n18490 | n18491;
  assign n40854 = n18492 | n18493;
  assign n40855 = n18494 | ~n18495;
  assign n40856 = n18500 | ~n18501;
  assign n40857 = n18514 | n18515;
  assign n40858 = n18518 | n18519;
  assign n40859 = n18520 | n18521;
  assign n40860 = n18531 | n18532;
  assign n40861 = n18533 | n18534;
  assign n40862 = n18535 | ~n18536;
  assign n40863 = n18539 | n18540;
  assign n40864 = n18544 | n18545;
  assign n40865 = n18546 | n18547;
  assign n40866 = n18548 | ~n18549;
  assign n40867 = n18552 | n18553;
  assign n40868 = n18557 | n18558;
  assign n40869 = n18559 | n18560;
  assign n40870 = n18561 | ~n18562;
  assign n40871 = n18565 | n18566;
  assign n40872 = n18580 | n18581;
  assign n40873 = n18584 | n18585;
  assign n40874 = n18586 | n18587;
  assign n40875 = n18591 | n18592;
  assign n40876 = n18593 | n18594;
  assign n40877 = n18595 | ~n18596;
  assign n40878 = n18606 | n18607;
  assign n40879 = n18610 | n18611;
  assign n40880 = n18612 | n18613;
  assign n40881 = n18617 | n18618;
  assign n40882 = n18619 | n18620;
  assign n40883 = n18621 | ~n18622;
  assign n40884 = n18627 | ~n18628;
  assign n40885 = n18640 | ~n18641;
  assign n40886 = n18648 | n18649;
  assign n40887 = n18652 | n18653;
  assign n40888 = n18654 | n18655;
  assign n40889 = n18661 | ~n18662;
  assign n40890 = n18667 | ~n18668;
  assign n40891 = n18684 | n18678 | ~n18683;
  assign n40892 = n18691 | n18692;
  assign n40893 = n18693 | n18694;
  assign n40894 = n18703 | n18704;
  assign n40895 = n18707 | n18708;
  assign n40896 = n18709 | n18710;
  assign n40897 = n18719 | n18720;
  assign n40898 = n18723 | n18724;
  assign n40899 = n18725 | n18726;
  assign n40900 = n18735 | n18736;
  assign n40901 = n18739 | n18740;
  assign n40902 = n18741 | n18742;
  assign n40903 = n18751 | n18752;
  assign n40904 = n18755 | n18756;
  assign n40905 = n18757 | n18758;
  assign n40906 = n18767 | n18768;
  assign n40907 = n18771 | n18772;
  assign n40908 = n18773 | n18774;
  assign n40909 = n18783 | n18784;
  assign n40910 = n18787 | n18788;
  assign n40911 = n18789 | n18790;
  assign n40912 = n18808 | n18809;
  assign n40913 = n18812 | n18813;
  assign n40914 = n18814 | n18815;
  assign n40915 = n18822 | n18823;
  assign n40916 = n18824 | n18825;
  assign n40917 = n18826 | ~n18827;
  assign n40918 = n18837 | n18838;
  assign n40919 = n18841 | n18842;
  assign n40920 = n18843 | n18844;
  assign n40921 = n18858 | n18859;
  assign n40922 = n18862 | n18863;
  assign n40923 = n18864 | n18865;
  assign n40924 = n18869 | n18870;
  assign n40925 = n18871 | n18872;
  assign n40926 = n18873 | ~n18874;
  assign n40927 = n18884 | n18885;
  assign n40928 = n18888 | n18889;
  assign n40929 = n18890 | n18891;
  assign n40930 = n18906 | n18907;
  assign n40931 = n18910 | n18911;
  assign n40932 = n18912 | n18913;
  assign n40933 = n18917 | n18918;
  assign n40934 = n18919 | n18920;
  assign n40935 = n18921 | ~n18922;
  assign n40936 = n18932 | n18933;
  assign n40937 = n18936 | n18937;
  assign n40938 = n18938 | n18939;
  assign n40939 = n18954 | n18955;
  assign n40940 = n18958 | n18959;
  assign n40941 = n18960 | n18961;
  assign n40942 = n18965 | n18966;
  assign n40943 = n18967 | n18968;
  assign n40944 = n18969 | ~n18970;
  assign n40945 = n18980 | n18981;
  assign n40946 = n18984 | n18985;
  assign n40947 = n18986 | n18987;
  assign n40948 = n18991 | n18992;
  assign n40949 = n18993 | n18994;
  assign n40950 = n18995 | ~n18996;
  assign n40951 = n19006 | n19007;
  assign n40952 = n19010 | n19011;
  assign n40953 = n19012 | n19013;
  assign n40954 = n19017 | n19018;
  assign n40955 = n19019 | n19020;
  assign n40956 = n19021 | ~n19022;
  assign n40957 = n19032 | n19033;
  assign n40958 = n19036 | n19037;
  assign n40959 = n19038 | n19039;
  assign n40960 = n19054 | n19055;
  assign n40961 = n19058 | n19059;
  assign n40962 = n19060 | n19061;
  assign n40963 = n19065 | n19066;
  assign n40964 = n19067 | n19068;
  assign n40965 = n19069 | ~n19070;
  assign n40966 = n19080 | n19081;
  assign n40967 = n19084 | n19085;
  assign n40968 = n19086 | n19087;
  assign n40969 = n19091 | n19092;
  assign n40970 = n19093 | n19094;
  assign n40971 = n19095 | ~n19096;
  assign n40972 = n19106 | n19107;
  assign n40973 = n19110 | n19111;
  assign n40974 = n19112 | n19113;
  assign n40975 = n19117 | n19118;
  assign n40976 = n19119 | n19120;
  assign n40977 = n19121 | ~n19122;
  assign n40978 = n19125 | n19126;
  assign n40979 = n19127 | n19128;
  assign n40980 = n19129 | ~n19130;
  assign n40981 = n19135 | ~n19136;
  assign n40982 = n19142 | n19143;
  assign n40983 = n19144 | n19145;
  assign n40984 = n19146 | ~n19147;
  assign n40985 = n19150 | n19151;
  assign n40986 = n19155 | n19156;
  assign n40987 = n19157 | n19158;
  assign n40988 = n19159 | ~n19160;
  assign n40989 = n19163 | n19164;
  assign n40990 = n19184 | n19185;
  assign n40991 = n19188 | n19189;
  assign n40992 = n19190 | n19191;
  assign n40993 = n19195 | n19196;
  assign n40994 = n19197 | n19198;
  assign n40995 = n19199 | ~n19200;
  assign n40996 = n19205 | ~n19206;
  assign n40997 = n19214 | ~n19215;
  assign n40998 = n19225 | n19226;
  assign n40999 = n19238 | n19234 | ~n19237;
  assign n41000 = n19251 | n19252;
  assign n41001 = n19255 | n19256;
  assign n41002 = n19257 | n19258;
  assign n41003 = n19267 | n19268;
  assign n41004 = n19271 | n19272;
  assign n41005 = n19273 | n19274;
  assign n41006 = n19283 | n19284;
  assign n41007 = n19287 | n19288;
  assign n41008 = n19289 | n19290;
  assign n41009 = n19301 | n19302;
  assign n41010 = n19305 | n19306;
  assign n41011 = n19307 | n19308;
  assign n41012 = n19320 | n19321;
  assign n41013 = n19324 | n19325;
  assign n41014 = n19326 | n19327;
  assign n41015 = n19337 | n19338;
  assign n41016 = n19341 | n19342;
  assign n41017 = n19343 | n19344;
  assign n41018 = n19354 | n19355;
  assign n41019 = n19358 | n19359;
  assign n41020 = n19360 | n19361;
  assign n41021 = n19371 | n19372;
  assign n41022 = n19375 | n19376;
  assign n41023 = n19377 | n19378;
  assign n41024 = n19385 | n19386;
  assign n41025 = n19387 | n19388;
  assign n41026 = n19389 | ~n19390;
  assign n41027 = n19400 | n19401;
  assign n41028 = n19404 | n19405;
  assign n41029 = n19406 | n19407;
  assign n41030 = n19413 | n19414;
  assign n41031 = n19419 | ~n19420;
  assign n41032 = n19433 | n19434;
  assign n41033 = n19437 | n19438;
  assign n41034 = n19439 | n19440;
  assign n41035 = n19444 | n19445;
  assign n41036 = n19446 | n19447;
  assign n41037 = n19448 | ~n19449;
  assign n41038 = n19454 | ~n19455;
  assign n41039 = n19468 | n19469;
  assign n41040 = n19472 | n19473;
  assign n41041 = n19474 | n19475;
  assign n41042 = n19479 | n19480;
  assign n41043 = n19481 | n19482;
  assign n41044 = n19483 | ~n19484;
  assign n41045 = n19489 | ~n19490;
  assign n41046 = n19503 | n19504;
  assign n41047 = n19507 | n19508;
  assign n41048 = n19509 | n19510;
  assign n41049 = n19514 | n19515;
  assign n41050 = n19516 | n19517;
  assign n41051 = n19518 | ~n19519;
  assign n41052 = n19529 | n19530;
  assign n41053 = n19533 | n19534;
  assign n41054 = n19535 | n19536;
  assign n41055 = n19540 | n19541;
  assign n41056 = n19542 | n19543;
  assign n41057 = n19544 | ~n19545;
  assign n41058 = n19555 | n19556;
  assign n41059 = n19559 | n19560;
  assign n41060 = n19561 | n19562;
  assign n41061 = n19568 | n19569;
  assign n41062 = n19574 | ~n19575;
  assign n41063 = n19578 | n19579;
  assign n41064 = n19580 | n19581;
  assign n41065 = n19582 | ~n19583;
  assign n41066 = n19593 | n19594;
  assign n41067 = n19597 | n19598;
  assign n41068 = n19599 | n19600;
  assign n41069 = n19604 | n19605;
  assign n41070 = n19606 | n19607;
  assign n41071 = n19608 | ~n19609;
  assign n41072 = n19619 | n19620;
  assign n41073 = n19623 | n19624;
  assign n41074 = n19625 | n19626;
  assign n41075 = n19632 | n19633;
  assign n41076 = n19638 | ~n19639;
  assign n41077 = n19642 | n19643;
  assign n41078 = n19644 | n19645;
  assign n41079 = n19646 | ~n19647;
  assign n41080 = n19653 | n19654;
  assign n41081 = n19655 | n19656;
  assign n41082 = n19657 | ~n19658;
  assign n41083 = n19661 | n19662;
  assign n41084 = n19663 | n19664;
  assign n41085 = n19665 | ~n19666;
  assign n41086 = n19679 | n19680;
  assign n41087 = n19683 | n19684;
  assign n41088 = n19685 | n19686;
  assign n41089 = n19690 | n19691;
  assign n41090 = n19692 | n19693;
  assign n41091 = n19694 | ~n19695;
  assign n41092 = n19705 | n19706;
  assign n41093 = n19709 | n19710;
  assign n41094 = n19711 | n19712;
  assign n41095 = n19723 | n19724;
  assign n41096 = n19727 | n19728;
  assign n41097 = n19729 | n19730;
  assign n41098 = n19736 | ~n19737;
  assign n41099 = n19747 | n19748;
  assign n41100 = n19751 | n19752;
  assign n41101 = n19753 | n19754;
  assign n41102 = n19760 | ~n19761;
  assign n41103 = n19766 | ~n19767;
  assign n41104 = n19781 | n19782;
  assign n41105 = n19785 | n19786;
  assign n41106 = n19787 | n19788;
  assign n41107 = n19791 | n19792;
  assign n41108 = n19795 | n19796;
  assign n41109 = n19797 | n19798;
  assign n41110 = n19799 | ~n19800;
  assign n41111 = n19807 | n19808;
  assign n41112 = n19811 | n19812;
  assign n41113 = n19813 | n19814;
  assign n41114 = n19826 | n19827;
  assign n41115 = n19830 | n19831;
  assign n41116 = n19832 | n19833;
  assign n41117 = n19845 | n19846;
  assign n41118 = n19849 | n19850;
  assign n41119 = n19851 | n19852;
  assign n41120 = n19864 | n19865;
  assign n41121 = n19868 | n19869;
  assign n41122 = n19870 | n19871;
  assign n41123 = n19884 | n19885;
  assign n41124 = n19888 | ~n19889;
  assign n41125 = n19902 | n19903;
  assign n41126 = n19906 | ~n19907;
  assign n41127 = n19913 | n19914;
  assign n41128 = n19915 | n19916;
  assign n41129 = n19917 | ~n19918;
  assign n41130 = n19930 | n19931;
  assign n41131 = n19934 | n19935;
  assign n41132 = n19936 | n19937;
  assign n41133 = n19952 | n19953;
  assign n41134 = n19956 | ~n19957;
  assign n41135 = n19973 | n19974;
  assign n41136 = n19977 | n19978;
  assign n41137 = n19979 | n19980;
  assign n41138 = n19986 | ~n19987;
  assign n41139 = n19992 | ~n19993;
  assign n41140 = n20006 | n20007;
  assign n41141 = n20010 | n20011;
  assign n41142 = n20012 | n20013;
  assign n41143 = n20019 | ~n20020;
  assign n41144 = n20030 | n20031;
  assign n41145 = n20034 | n20035;
  assign n41146 = n20036 | n20037;
  assign n41147 = n20043 | ~n20044;
  assign n41148 = n20054 | n20055;
  assign n41149 = n20058 | n20059;
  assign n41150 = n20060 | n20061;
  assign n41151 = n20076 | n20077;
  assign n41152 = n20080 | n20081;
  assign n41153 = n20082 | n20083;
  assign n41154 = n20089 | ~n20090;
  assign n41155 = n20100 | n20101;
  assign n41156 = n20104 | n20105;
  assign n41157 = n20106 | n20107;
  assign n41158 = n20113 | ~n20114;
  assign n41159 = n20124 | n20125;
  assign n41160 = n20128 | n20129;
  assign n41161 = n20130 | n20131;
  assign n41162 = n20146 | n20147;
  assign n41163 = n20150 | n20151;
  assign n41164 = n20152 | n20153;
  assign n41165 = n20159 | ~n20160;
  assign n41166 = n20165 | ~n20166;
  assign n41167 = n20171 | ~n20172;
  assign n41168 = n20182 | n20183;
  assign n41169 = n20186 | n20187;
  assign n41170 = n20188 | n20189;
  assign n41171 = n20195 | ~n20196;
  assign n41172 = n20198 | n20199;
  assign n41173 = n20203 | n20204;
  assign n41174 = n20205 | ~n20206;
  assign n41175 = n20211 | n20212;
  assign n41176 = n20216 | n20217;
  assign n41177 = n20218 | ~n20219;
  assign n41178 = n20227 | n20228;
  assign n41179 = n20231 | ~n20232;
  assign n41180 = n20238 | n20239;
  assign n41181 = n20240 | n20241;
  assign n41182 = n20242 | ~n20243;
  assign n41183 = n20246 | n20247;
  assign n41184 = n20248 | n20249;
  assign n41185 = n20250 | ~n20251;
  assign n41186 = n20253 | n20254;
  assign n41187 = n20255 | n20256;
  assign n41188 = n20258 | ~n20259;
  assign n41189 = n20264 | ~n20265;
  assign n41190 = n20272 | n20273;
  assign n41191 = n20276 | n20277;
  assign n41192 = n20278 | n20279;
  assign n41193 = n20282 | ~n20283;
  assign n41194 = n20286 | n20287;
  assign n41195 = n20288 | n20289;
  assign n41196 = n20290 | ~n20291;
  assign n41197 = n20294 | n20295;
  assign n41198 = n20296 | n20297;
  assign n41199 = n20298 | ~n20299;
  assign n41200 = n20301 | ~n20302;
  assign n41201 = n20318 | n20319;
  assign n41202 = n20322 | n20323;
  assign n41203 = n20324 | n20325;
  assign n41204 = n20337 | n20338;
  assign n41205 = n20341 | n20342;
  assign n41206 = n20343 | n20344;
  assign n41207 = n20349 | n20350;
  assign n41208 = n20351 | n20352;
  assign n41209 = n20353 | ~n20354;
  assign n41210 = n20361 | n20362;
  assign n41211 = n20365 | n20366;
  assign n41212 = n20367 | n20368;
  assign n41213 = n20380 | n20381;
  assign n41214 = n20384 | n20385;
  assign n41215 = n20386 | n20387;
  assign n41216 = n20399 | n20400;
  assign n41217 = n20403 | ~n20404;
  assign n41218 = n20409 | n20410;
  assign n41219 = n20420 | n20421;
  assign n41220 = n20424 | n20425;
  assign n41221 = n20426 | n20427;
  assign n41222 = n20436 | n20437;
  assign n41223 = n20440 | n20441;
  assign n41224 = n20442 | n20443;
  assign n41225 = n20453 | n20454;
  assign n41226 = n20457 | n20458;
  assign n41227 = n20459 | n20460;
  assign n41228 = n20467 | n20468;
  assign n41229 = n20469 | n20470;
  assign n41230 = n20471 | ~n20472;
  assign n41231 = n20475 | n20476;
  assign n41232 = n20477 | n20478;
  assign n41233 = n20479 | ~n20480;
  assign n41234 = n20490 | n20491;
  assign n41235 = n20494 | n20495;
  assign n41236 = n20496 | n20497;
  assign n41237 = n20503 | ~n20504;
  assign n41238 = n20506 | ~n20507;
  assign n41239 = n20517 | n20518;
  assign n41240 = n20521 | n20522;
  assign n41241 = n20523 | n20524;
  assign n41242 = n20539 | n20540;
  assign n41243 = n20543 | n20544;
  assign n41244 = n20545 | n20546;
  assign n41245 = n20552 | ~n20553;
  assign n41246 = n20555 | ~n20556;
  assign n41247 = n20566 | n20567;
  assign n41248 = n20570 | n20571;
  assign n41249 = n20572 | n20573;
  assign n41250 = n20579 | ~n20580;
  assign n41251 = n20582 | ~n20583;
  assign n41252 = n20593 | n20594;
  assign n41253 = n20597 | n20598;
  assign n41254 = n20599 | n20600;
  assign n41255 = n20606 | ~n20607;
  assign n41256 = n20612 | ~n20613;
  assign n41257 = n20618 | ~n20619;
  assign n41258 = n20621 | n20622;
  assign n41259 = n20632 | n20633;
  assign n41260 = n20636 | n20637;
  assign n41261 = n20638 | n20639;
  assign n41262 = n20645 | ~n20646;
  assign n41263 = n20648 | ~n20649;
  assign n41264 = n20659 | n20660;
  assign n41265 = n20663 | n20664;
  assign n41266 = n20665 | n20666;
  assign n41267 = n20675 | ~n20676;
  assign n41268 = n20681 | ~n20682;
  assign n41269 = n20693 | n20694;
  assign n41270 = n20697 | ~n20698;
  assign n41271 = n20704 | n20705;
  assign n41272 = n20706 | n20707;
  assign n41273 = n20708 | ~n20709;
  assign n41274 = n20714 | ~n20715;
  assign n41275 = n20720 | ~n20721;
  assign n41276 = n20728 | n20729;
  assign n41277 = n20732 | n20733;
  assign n41278 = n20734 | n20735;
  assign n41279 = n20740 | n20741;
  assign n41280 = n20742 | n20743;
  assign n41281 = n20744 | ~n20745;
  assign n41282 = n20750 | ~n20751;
  assign n41283 = n20753 | n20754;
  assign n41284 = n20755 | n20756;
  assign n41285 = n20758 | ~n20759;
  assign n41286 = n20764 | ~n20765;
  assign n41287 = n20770 | ~n20771;
  assign n41288 = n20779 | n20780;
  assign n41289 = n20783 | ~n20784;
  assign n41290 = n20790 | n20791;
  assign n41291 = n20792 | n20793;
  assign n41292 = n20794 | ~n20795;
  assign n41293 = n20798 | n20799;
  assign n41294 = n20800 | n20801;
  assign n41295 = n20802 | ~n20803;
  assign n41296 = n20810 | n20811;
  assign n41297 = n20814 | ~n20815;
  assign n41298 = n20820 | ~n20821;
  assign n41299 = n20824 | n20825;
  assign n41300 = n20826 | n20827;
  assign n41301 = n20828 | ~n20829;
  assign n41302 = n20834 | ~n20835;
  assign n41303 = n20843 | ~n20844;
  assign n41304 = n20850 | n20851;
  assign n41305 = n20852 | n20853;
  assign n41306 = n20854 | ~n20855;
  assign n41307 = n20861 | n20858 | n20860;
  assign n41308 = n20867 | ~n20868;
  assign n41309 = n20871 | n20872;
  assign n41310 = n20882 | n20883;
  assign n41311 = n20886 | n20887;
  assign n41312 = n20888 | n20889;
  assign n41313 = n20901 | n20902;
  assign n41314 = n20905 | n20906;
  assign n41315 = n20907 | n20908;
  assign n41316 = n20913 | n20914;
  assign n41317 = n20915 | n20916;
  assign n41318 = n20917 | ~n20918;
  assign n41319 = n20925 | n20926;
  assign n41320 = n20929 | ~n20930;
  assign n41321 = n20935 | ~n20936;
  assign n41322 = n20946 | n20947;
  assign n41323 = n20950 | n20951;
  assign n41324 = n20952 | n20953;
  assign n41325 = n20966 | n20967;
  assign n41326 = n20970 | ~n20971;
  assign n41327 = n20977 | n20978;
  assign n41328 = n20979 | n20980;
  assign n41329 = n20981 | ~n20982;
  assign n41330 = n20989 | n20990;
  assign n41331 = n20993 | n20994;
  assign n41332 = n20995 | n20996;
  assign n41333 = n21008 | n21009;
  assign n41334 = n21012 | ~n21013;
  assign n41335 = n21018 | ~n21019;
  assign n41336 = n21024 | n21025;
  assign n41337 = n21028 | n21029;
  assign n41338 = n21036 | n21037;
  assign n41339 = n21040 | n21041;
  assign n41340 = n21042 | n21043;
  assign n41341 = n21053 | n21054;
  assign n41342 = n21057 | n21058;
  assign n41343 = n21059 | n21060;
  assign n41344 = n21067 | n21068;
  assign n41345 = n21069 | n21070;
  assign n41346 = n21071 | ~n21072;
  assign n41347 = n21075 | n21076;
  assign n41348 = n21077 | n21078;
  assign n41349 = n21079 | ~n21080;
  assign n41350 = n21090 | n21091;
  assign n41351 = n21094 | n21095;
  assign n41352 = n21096 | n21097;
  assign n41353 = n21103 | ~n21104;
  assign n41354 = n21114 | n21115;
  assign n41355 = n21118 | n21119;
  assign n41356 = n21120 | n21121;
  assign n41357 = n21127 | ~n21128;
  assign n41358 = n21133 | ~n21134;
  assign n41359 = n21136 | n21137;
  assign n41360 = n21138 | n21139;
  assign n41361 = n21141 | ~n21142;
  assign n41362 = n21152 | n21153;
  assign n41363 = n21156 | n21157;
  assign n41364 = n21158 | n21159;
  assign n41365 = n21165 | ~n21166;
  assign n41366 = n21176 | n21177;
  assign n41367 = n21180 | n21181;
  assign n41368 = n21182 | n21183;
  assign n41369 = n21189 | ~n21190;
  assign n41370 = n21192 | ~n21193;
  assign n41371 = n21203 | n21204;
  assign n41372 = n21207 | n21208;
  assign n41373 = n21209 | n21210;
  assign n41374 = n21216 | ~n21217;
  assign n41375 = n21227 | n21228;
  assign n41376 = n21231 | n21232;
  assign n41377 = n21233 | n21234;
  assign n41378 = n21240 | ~n21241;
  assign n41379 = n21251 | n21252;
  assign n41380 = n21255 | n21256;
  assign n41381 = n21257 | n21258;
  assign n41382 = n21273 | n21274;
  assign n41383 = n21277 | n21278;
  assign n41384 = n21279 | n21280;
  assign n41385 = n21286 | ~n21287;
  assign n41386 = n21292 | ~n21293;
  assign n41387 = n21298 | ~n21299;
  assign n41388 = n21304 | ~n21305;
  assign n41389 = n21310 | ~n21311;
  assign n41390 = n21318 | n21319;
  assign n41391 = n21322 | n21323;
  assign n41392 = n21324 | n21325;
  assign n41393 = n21330 | n21331;
  assign n41394 = n21332 | n21333;
  assign n41395 = n21334 | ~n21335;
  assign n41396 = n21340 | ~n21341;
  assign n41397 = n21346 | ~n21347;
  assign n41398 = n21352 | ~n21353;
  assign n41399 = n21358 | ~n21359;
  assign n41400 = n21367 | n21368;
  assign n41401 = n21371 | ~n21372;
  assign n41402 = n21378 | n21379;
  assign n41403 = n21380 | n21381;
  assign n41404 = n21382 | ~n21383;
  assign n41405 = n21389 | n21386 | n21388;
  assign n41406 = n21396 | ~n21397;
  assign n41407 = n21399 | n21400;
  assign n41408 = n21401 | n21402;
  assign n41409 = n21408 | ~n21409;
  assign n41410 = n21417 | ~n21418;
  assign n41411 = n21421 | n21422;
  assign n41412 = n21433 | n21434;
  assign n41413 = n21437 | n21438;
  assign n41414 = n21439 | n21440;
  assign n41415 = n21444 | n21445;
  assign n41416 = n21446 | n21447;
  assign n41417 = n21448 | ~n21449;
  assign n41418 = n21456 | n21457;
  assign n41419 = n21460 | n21461;
  assign n41420 = n21462 | n21463;
  assign n41421 = n21475 | n21476;
  assign n41422 = n21479 | n21480;
  assign n41423 = n21481 | n21482;
  assign n41424 = n21494 | n21495;
  assign n41425 = n21498 | n21499;
  assign n41426 = n21500 | n21501;
  assign n41427 = n21504 | ~n21505;
  assign n41428 = n21508 | n21509;
  assign n41429 = n21510 | n21511;
  assign n41430 = n21512 | ~n21513;
  assign n41431 = n21520 | n21521;
  assign n41432 = n21524 | n21525;
  assign n41433 = n21526 | n21527;
  assign n41434 = n21539 | n21540;
  assign n41435 = n21543 | n21544;
  assign n41436 = n21545 | n21546;
  assign n41437 = n21558 | n21559;
  assign n41438 = n21562 | n21563;
  assign n41439 = n21564 | n21565;
  assign n41440 = n21568 | ~n21569;
  assign n41441 = n21579 | n21580;
  assign n41442 = n21583 | n21584;
  assign n41443 = n21585 | n21586;
  assign n41444 = n21595 | n21596;
  assign n41445 = n21599 | n21600;
  assign n41446 = n21601 | n21602;
  assign n41447 = n21610 | n21611;
  assign n41448 = n21614 | n21615;
  assign n41449 = n21616 | n21617;
  assign n41450 = n21626 | n21627;
  assign n41451 = n21630 | n21631;
  assign n41452 = n21632 | n21633;
  assign n41453 = n21642 | n21643;
  assign n41454 = n21646 | n21647;
  assign n41455 = n21648 | n21649;
  assign n41456 = n21656 | ~n21657;
  assign n41457 = n21673 | n21674;
  assign n41458 = n21677 | n21678;
  assign n41459 = n21679 | n21680;
  assign n41460 = n21687 | n21688;
  assign n41461 = n21689 | n21690;
  assign n41462 = n21691 | ~n21692;
  assign n41463 = n21697 | ~n21698;
  assign n41464 = n21701 | n21702;
  assign n41465 = n21703 | n21704;
  assign n41466 = n21705 | ~n21706;
  assign n41467 = n21708 | ~n21709;
  assign n41468 = n21719 | n21720;
  assign n41469 = n21723 | n21724;
  assign n41470 = n21725 | n21726;
  assign n41471 = n21730 | n21731;
  assign n41472 = n21732 | n21733;
  assign n41473 = n21734 | ~n21735;
  assign n41474 = n21737 | ~n21738;
  assign n41475 = n21748 | n21749;
  assign n41476 = n21752 | n21753;
  assign n41477 = n21754 | n21755;
  assign n41478 = n21759 | n21760;
  assign n41479 = n21761 | n21762;
  assign n41480 = n21763 | ~n21764;
  assign n41481 = n21769 | ~n21770;
  assign n41482 = n21775 | ~n21776;
  assign n41483 = n21786 | n21787;
  assign n41484 = n21790 | n21791;
  assign n41485 = n21792 | n21793;
  assign n41486 = n21797 | n21798;
  assign n41487 = n21799 | n21800;
  assign n41488 = n21801 | ~n21802;
  assign n41489 = n21804 | ~n21805;
  assign n41490 = n21815 | n21816;
  assign n41491 = n21819 | n21820;
  assign n41492 = n21821 | n21822;
  assign n41493 = n21828 | ~n21829;
  assign n41494 = n21833 | n21834;
  assign n41495 = n21835 | ~n21836;
  assign n41496 = n21837 | n21838;
  assign n41497 = n21839 | n21840;
  assign n41498 = n21846 | ~n21847;
  assign n41499 = n21852 | ~n21853;
  assign n41500 = n21858 | n21859;
  assign n41501 = n21869 | n21870;
  assign n41502 = n21873 | n21874;
  assign n41503 = n21875 | n21876;
  assign n41504 = n21879 | ~n21880;
  assign n41505 = n21897 | n21898;
  assign n41506 = n21901 | n21902;
  assign n41507 = n21903 | n21904;
  assign n41508 = n21908 | n21909;
  assign n41509 = n21910 | n21911;
  assign n41510 = n21912 | ~n21913;
  assign n41511 = n21918 | ~n21919;
  assign n41512 = n21921 | n21922;
  assign n41513 = n21923 | n21924;
  assign n41514 = n21926 | ~n21927;
  assign n41515 = n21932 | ~n21933;
  assign n41516 = n21938 | ~n21939;
  assign n41517 = n21944 | ~n21945;
  assign n41518 = n21947 | n21948;
  assign n41519 = n21949 | n21950;
  assign n41520 = n21952 | ~n21953;
  assign n41521 = n21958 | ~n21959;
  assign n41522 = n21974 | ~n21975;
  assign n41523 = n21980 | ~n21981;
  assign n41524 = n21991 | n21992;
  assign n41525 = n21995 | n21996;
  assign n41526 = n21997 | n21998;
  assign n41527 = n22011 | n22012;
  assign n41528 = n22015 | ~n22016;
  assign n41529 = n22029 | n22030;
  assign n41530 = n22033 | n22034;
  assign n41531 = n22035 | n22036;
  assign n41532 = n22039 | ~n22040;
  assign n41533 = n22050 | n22051;
  assign n41534 = n22054 | n22055;
  assign n41535 = n22056 | n22057;
  assign n41536 = n22060 | ~n22061;
  assign n41537 = n22072 | n22073;
  assign n41538 = n22076 | ~n22077;
  assign n41539 = n22090 | n22091;
  assign n41540 = n22094 | n22095;
  assign n41541 = n22096 | n22097;
  assign n41542 = n22102 | n22103;
  assign n41543 = n22104 | n22105;
  assign n41544 = n22106 | ~n22107;
  assign n41545 = n22114 | n22115;
  assign n41546 = n22118 | n22119;
  assign n41547 = n22120 | n22121;
  assign n41548 = n22133 | n22134;
  assign n41549 = n22137 | n22138;
  assign n41550 = n22139 | n22140;
  assign n41551 = n22149 | n22150;
  assign n41552 = n22153 | n22154;
  assign n41553 = n22155 | n22156;
  assign n41554 = n22178 | n22179;
  assign n41555 = n22182 | ~n22183;
  assign n41556 = n22199 | n22200;
  assign n41557 = n22203 | n22204;
  assign n41558 = n22205 | n22206;
  assign n41559 = n22212 | ~n22213;
  assign n41560 = n22223 | n22224;
  assign n41561 = n22227 | n22228;
  assign n41562 = n22229 | n22230;
  assign n41563 = n22236 | ~n22237;
  assign n41564 = n22247 | n22248;
  assign n41565 = n22251 | n22252;
  assign n41566 = n22253 | n22254;
  assign n41567 = n22260 | ~n22261;
  assign n41568 = n22271 | n22272;
  assign n41569 = n22275 | n22276;
  assign n41570 = n22277 | n22278;
  assign n41571 = n22284 | ~n22285;
  assign n41572 = n22295 | n22296;
  assign n41573 = n22299 | n22300;
  assign n41574 = n22301 | n22302;
  assign n41575 = n22308 | ~n22309;
  assign n41576 = n22319 | n22320;
  assign n41577 = n22323 | n22324;
  assign n41578 = n22325 | n22326;
  assign n41579 = n22332 | ~n22333;
  assign n41580 = n22343 | n22344;
  assign n41581 = n22347 | n22348;
  assign n41582 = n22349 | n22350;
  assign n41583 = n22368 | ~n22369;
  assign n41584 = n22374 | ~n22375;
  assign n41585 = n22380 | ~n22381;
  assign n41586 = n22386 | ~n22387;
  assign n41587 = n22394 | n22395;
  assign n41588 = n22398 | n22399;
  assign n41589 = n22400 | n22401;
  assign n41590 = n22406 | n22407;
  assign n41591 = n22408 | n22409;
  assign n41592 = n22410 | ~n22411;
  assign n41593 = n22416 | ~n22417;
  assign n41594 = n22422 | ~n22423;
  assign n41595 = n22428 | n22429;
  assign n41596 = n22433 | n22434;
  assign n41597 = n22435 | ~n22436;
  assign n41598 = n22441 | n22442;
  assign n41599 = n22446 | n22447;
  assign n41600 = n22448 | ~n22449;
  assign n41601 = n22454 | ~n22455;
  assign n41602 = n22466 | n22467;
  assign n41603 = n22470 | n22471;
  assign n41604 = n22472 | n22473;
  assign n41605 = n22478 | n22479;
  assign n41606 = n22480 | n22481;
  assign n41607 = n22482 | ~n22483;
  assign n41608 = n22490 | n22491;
  assign n41609 = n22494 | n22495;
  assign n41610 = n22496 | n22497;
  assign n41611 = n22500 | ~n22501;
  assign n41612 = n22511 | n22512;
  assign n41613 = n22515 | n22516;
  assign n41614 = n22517 | n22518;
  assign n41615 = n22530 | n22531;
  assign n41616 = n22534 | n22535;
  assign n41617 = n22536 | n22537;
  assign n41618 = n22542 | n22543;
  assign n41619 = n22544 | n22545;
  assign n41620 = n22546 | ~n22547;
  assign n41621 = n22554 | n22555;
  assign n41622 = n22558 | n22559;
  assign n41623 = n22560 | n22561;
  assign n41624 = n22564 | ~n22565;
  assign n41625 = n22576 | n22577;
  assign n41626 = n22580 | n22581;
  assign n41627 = n22582 | n22583;
  assign n41628 = n22591 | n22592;
  assign n41629 = n22595 | n22596;
  assign n41630 = n22597 | n22598;
  assign n41631 = n22606 | n22607;
  assign n41632 = n22610 | n22611;
  assign n41633 = n22612 | n22613;
  assign n41634 = n22623 | n22624;
  assign n41635 = n22629 | ~n22630;
  assign n41636 = n22635 | ~n22636;
  assign n41637 = n22641 | ~n22642;
  assign n41638 = n22652 | n22653;
  assign n41639 = n22656 | n22657;
  assign n41640 = n22658 | n22659;
  assign n41641 = n22665 | ~n22666;
  assign n41642 = n22668 | ~n22669;
  assign n41643 = n22679 | n22680;
  assign n41644 = n22683 | n22684;
  assign n41645 = n22685 | n22686;
  assign n41646 = n22692 | ~n22693;
  assign n41647 = n22698 | ~n22699;
  assign n41648 = n22702 | n22703;
  assign n41649 = n22706 | ~n22707;
  assign n41650 = n22717 | n22718;
  assign n41651 = n22721 | n22722;
  assign n41652 = n22723 | n22724;
  assign n41653 = n22730 | ~n22731;
  assign n41654 = n22733 | ~n22734;
  assign n41655 = n22744 | n22745;
  assign n41656 = n22748 | n22749;
  assign n41657 = n22750 | n22751;
  assign n41658 = n22757 | ~n22758;
  assign n41659 = n22760 | ~n22761;
  assign n41660 = n22771 | n22772;
  assign n41661 = n22775 | n22776;
  assign n41662 = n22777 | n22778;
  assign n41663 = n22793 | n22794;
  assign n41664 = n22797 | n22798;
  assign n41665 = n22799 | n22800;
  assign n41666 = n22806 | ~n22807;
  assign n41667 = n22817 | n22818;
  assign n41668 = n22821 | n22822;
  assign n41669 = n22823 | n22824;
  assign n41670 = n22830 | n22831;
  assign n41671 = n22835 | n22836;
  assign n41672 = n22837 | ~n22838;
  assign n41673 = n22845 | n22846;
  assign n41674 = n22849 | ~n22850;
  assign n41675 = n22855 | ~n22856;
  assign n41676 = n22859 | n22860;
  assign n41677 = n22861 | n22862;
  assign n41678 = n22863 | ~n22864;
  assign n41679 = n22867 | n22868;
  assign n41680 = n22869 | n22870;
  assign n41681 = n22871 | ~n22872;
  assign n41682 = n22877 | ~n22878;
  assign n41683 = n22889 | n22890;
  assign n41684 = n22893 | ~n22894;
  assign n41685 = n22900 | n22901;
  assign n41686 = n22902 | n22903;
  assign n41687 = n22904 | ~n22905;
  assign n41688 = n22908 | n22909;
  assign n41689 = n22910 | n22911;
  assign n41690 = n22912 | ~n22913;
  assign n41691 = n22918 | ~n22919;
  assign n41692 = n22924 | ~n22925;
  assign n41693 = n22933 | n22934;
  assign n41694 = n22937 | ~n22938;
  assign n41695 = n22944 | n22945;
  assign n41696 = n22946 | n22947;
  assign n41697 = n22948 | ~n22949;
  assign n41698 = n22955 | n22952 | n22954;
  assign n41699 = n22962 | ~n22963;
  assign n41700 = n22965 | n22966;
  assign n41701 = n22967 | n22968;
  assign n41702 = n22974 | ~n22975;
  assign n41703 = n22980 | ~n22981;
  assign n41704 = n22986 | ~n22987;
  assign n41705 = n22990 | n22991;
  assign n41706 = n23001 | n23002;
  assign n41707 = n23005 | n23006;
  assign n41708 = n23007 | n23008;
  assign n41709 = n23011 | ~n23012;
  assign n41710 = n23023 | n23024;
  assign n41711 = n23027 | n23028;
  assign n41712 = n23029 | n23030;
  assign n41713 = n23034 | n23035;
  assign n41714 = n23036 | n23037;
  assign n41715 = n23038 | ~n23039;
  assign n41716 = n23046 | n23047;
  assign n41717 = n23050 | n23051;
  assign n41718 = n23052 | n23053;
  assign n41719 = n23065 | n23066;
  assign n41720 = n23069 | n23070;
  assign n41721 = n23071 | n23072;
  assign n41722 = n23085 | n23086;
  assign n41723 = n23089 | n23090;
  assign n41724 = n23091 | n23092;
  assign n41725 = n23096 | n23097;
  assign n41726 = n23098 | n23099;
  assign n41727 = n23100 | ~n23101;
  assign n41728 = n23109 | n23110;
  assign n41729 = n23113 | n23114;
  assign n41730 = n23115 | n23116;
  assign n41731 = n23125 | n23126;
  assign n41732 = n23129 | n23130;
  assign n41733 = n23131 | n23132;
  assign n41734 = n23140 | n23141;
  assign n41735 = n23144 | n23145;
  assign n41736 = n23146 | n23147;
  assign n41737 = n23156 | n23157;
  assign n41738 = n23160 | n23161;
  assign n41739 = n23162 | n23163;
  assign n41740 = n23173 | n23174;
  assign n41741 = n23177 | n23178;
  assign n41742 = n23179 | n23180;
  assign n41743 = n23188 | n23189;
  assign n41744 = n23192 | n23193;
  assign n41745 = n23194 | n23195;
  assign n41746 = n23201 | ~n23202;
  assign n41747 = n23216 | ~n23217;
  assign n41748 = n23230 | n23231;
  assign n41749 = n23234 | n23235;
  assign n41750 = n23236 | n23237;
  assign n41751 = n23241 | n23242;
  assign n41752 = n23243 | n23244;
  assign n41753 = n23245 | ~n23246;
  assign n41754 = n23248 | ~n23249;
  assign n41755 = n23259 | n23260;
  assign n41756 = n23263 | n23264;
  assign n41757 = n23265 | n23266;
  assign n41758 = n23270 | n23271;
  assign n41759 = n23272 | n23273;
  assign n41760 = n23274 | ~n23275;
  assign n41761 = n23281 | n23282;
  assign n41762 = n23283 | n23284;
  assign n41763 = n23285 | ~n23286;
  assign n41764 = n23289 | n23290;
  assign n41765 = n23291 | n23292;
  assign n41766 = n23293 | ~n23294;
  assign n41767 = n23299 | ~n23300;
  assign n41768 = n23302 | ~n23303;
  assign n41769 = n23313 | n23314;
  assign n41770 = n23317 | n23318;
  assign n41771 = n23319 | n23320;
  assign n41772 = n23326 | ~n23327;
  assign n41773 = n23331 | n23332;
  assign n41774 = n23333 | ~n23334;
  assign n41775 = n23335 | n23336;
  assign n41776 = n23337 | n23338;
  assign n41777 = n23344 | ~n23345;
  assign n41778 = n23350 | ~n23351;
  assign n41779 = n23356 | n23357;
  assign n41780 = n23367 | n23368;
  assign n41781 = n23371 | n23372;
  assign n41782 = n23373 | n23374;
  assign n41783 = n23378 | n23379;
  assign n41784 = n23380 | n23381;
  assign n41785 = n23382 | ~n23383;
  assign n41786 = n23388 | ~n23389;
  assign n41787 = n23397 | n23398;
  assign n41788 = n23401 | n23402;
  assign n41789 = n23403 | n23404;
  assign n41790 = n23408 | n23409;
  assign n41791 = n23410 | n23411;
  assign n41792 = n23412 | ~n23413;
  assign n41793 = n23416 | n23417;
  assign n41794 = n23418 | n23419;
  assign n41795 = n23420 | ~n23421;
  assign n41796 = n23426 | ~n23427;
  assign n41797 = n23432 | ~n23433;
  assign n41798 = n23435 | n23436;
  assign n41799 = n23437 | n23438;
  assign n41800 = n23444 | ~n23445;
  assign n41801 = n23456 | n23457;
  assign n41802 = n23460 | n23461;
  assign n41803 = n23462 | n23463;
  assign n41804 = n23469 | ~n23470;
  assign n41805 = n23472 | n23473;
  assign n41806 = n23477 | n23478;
  assign n41807 = n23479 | ~n23480;
  assign n41808 = n23488 | n23489;
  assign n41809 = n23492 | n23493;
  assign n41810 = n23494 | n23495;
  assign n41811 = n23499 | n23500;
  assign n41812 = n23501 | n23502;
  assign n41813 = n23503 | ~n23504;
  assign n41814 = n23509 | ~n23510;
  assign n41815 = n23515 | ~n23516;
  assign n41816 = n23519 | n23520;
  assign n41817 = n23530 | n23531;
  assign n41818 = n23534 | n23535;
  assign n41819 = n23536 | n23537;
  assign n41820 = n23542 | n23543;
  assign n41821 = n23544 | n23545;
  assign n41822 = n23546 | ~n23547;
  assign n41823 = n23554 | n23555;
  assign n41824 = n23558 | n23559;
  assign n41825 = n23560 | n23561;
  assign n41826 = n23564 | ~n23565;
  assign n41827 = n23575 | n23576;
  assign n41828 = n23579 | n23580;
  assign n41829 = n23581 | n23582;
  assign n41830 = n23595 | n23596;
  assign n41831 = n23599 | ~n23600;
  assign n41832 = n23606 | n23607;
  assign n41833 = n23608 | n23609;
  assign n41834 = n23610 | ~n23611;
  assign n41835 = n23618 | n23619;
  assign n41836 = n23622 | n23623;
  assign n41837 = n23624 | n23625;
  assign n41838 = n23637 | n23638;
  assign n41839 = n23641 | n23642;
  assign n41840 = n23643 | n23644;
  assign n41841 = n23653 | n23654;
  assign n41842 = n23657 | n23658;
  assign n41843 = n23659 | n23660;
  assign n41844 = n23669 | n23670;
  assign n41845 = n23673 | n23674;
  assign n41846 = n23675 | n23676;
  assign n41847 = n23689 | n23690;
  assign n41848 = n23693 | n23694;
  assign n41849 = n23695 | n23696;
  assign n41850 = n23704 | n23705;
  assign n41851 = n23708 | n23709;
  assign n41852 = n23710 | n23711;
  assign n41853 = n23719 | n23720;
  assign n41854 = n23721 | n23722;
  assign n41855 = n23723 | ~n23724;
  assign n41856 = n23727 | n23728;
  assign n41857 = n23729 | n23730;
  assign n41858 = n23731 | ~n23732;
  assign n41859 = n23734 | ~n23735;
  assign n41860 = n23740 | ~n23741;
  assign n41861 = n23746 | ~n23747;
  assign n41862 = n23757 | n23758;
  assign n41863 = n23761 | n23762;
  assign n41864 = n23763 | n23764;
  assign n41865 = n23770 | ~n23771;
  assign n41866 = n23781 | n23782;
  assign n41867 = n23785 | n23786;
  assign n41868 = n23787 | n23788;
  assign n41869 = n23794 | ~n23795;
  assign n41870 = n23805 | n23806;
  assign n41871 = n23809 | n23810;
  assign n41872 = n23811 | n23812;
  assign n41873 = n23818 | ~n23819;
  assign n41874 = n23829 | n23830;
  assign n41875 = n23833 | n23834;
  assign n41876 = n23835 | n23836;
  assign n41877 = n23842 | ~n23843;
  assign n41878 = n23853 | n23854;
  assign n41879 = n23857 | n23858;
  assign n41880 = n23859 | n23860;
  assign n41881 = n23875 | ~n23876;
  assign n41882 = n23879 | n23880;
  assign n41883 = n23886 | ~n23887;
  assign n41884 = n23892 | ~n23893;
  assign n41885 = n23898 | ~n23899;
  assign n41886 = n23904 | ~n23905;
  assign n41887 = n23912 | n23913;
  assign n41888 = n23916 | n23917;
  assign n41889 = n23918 | n23919;
  assign n41890 = n23924 | n23925;
  assign n41891 = n23926 | n23927;
  assign n41892 = n23928 | ~n23929;
  assign n41893 = n23934 | ~n23935;
  assign n41894 = n23940 | n23941;
  assign n41895 = n23945 | n23946;
  assign n41896 = n23947 | ~n23948;
  assign n41897 = n23956 | n23957;
  assign n41898 = n23960 | ~n23961;
  assign n41899 = n23967 | n23968;
  assign n41900 = n23969 | n23970;
  assign n41901 = n23971 | ~n23972;
  assign n41902 = n23975 | n23976;
  assign n41903 = n23977 | n23978;
  assign n41904 = n23979 | ~n23980;
  assign n41905 = n23985 | ~n23986;
  assign n41906 = n23994 | ~n23995;
  assign n41907 = n24001 | n24002;
  assign n41908 = n24003 | n24004;
  assign n41909 = n24005 | ~n24006;
  assign n41910 = n24012 | n24009 | n24011;
  assign n41911 = n24018 | ~n24019;
  assign n41912 = n24022 | n24023;
  assign n41913 = n24034 | n24035;
  assign n41914 = n24038 | ~n24039;
  assign n41915 = n24052 | n24053;
  assign n41916 = n24056 | n24057;
  assign n41917 = n24058 | n24059;
  assign n41918 = n24071 | n24072;
  assign n41919 = n24075 | n24076;
  assign n41920 = n24077 | n24078;
  assign n41921 = n24083 | n24084;
  assign n41922 = n24085 | n24086;
  assign n41923 = n24087 | ~n24088;
  assign n41924 = n24096 | n24097;
  assign n41925 = n24100 | ~n24101;
  assign n41926 = n24114 | n24115;
  assign n41927 = n24118 | n24119;
  assign n41928 = n24120 | n24121;
  assign n41929 = n24124 | ~n24125;
  assign n41930 = n24135 | n24136;
  assign n41931 = n24139 | ~n24140;
  assign n41932 = n24145 | ~n24146;
  assign n41933 = n24156 | n24157;
  assign n41934 = n24160 | n24161;
  assign n41935 = n24162 | n24163;
  assign n41936 = n24173 | n24174;
  assign n41937 = n24177 | n24178;
  assign n41938 = n24179 | n24180;
  assign n41939 = n24188 | n24189;
  assign n41940 = n24192 | n24193;
  assign n41941 = n24194 | n24195;
  assign n41942 = n24203 | n24204;
  assign n41943 = n24207 | n24208;
  assign n41944 = n24209 | n24210;
  assign n41945 = n24218 | n24219;
  assign n41946 = n24222 | n24223;
  assign n41947 = n24224 | n24225;
  assign n41948 = n24233 | n24234;
  assign n41949 = n24235 | n24236;
  assign n41950 = n24237 | ~n24238;
  assign n41951 = n24241 | n24242;
  assign n41952 = n24243 | n24244;
  assign n41953 = n24245 | ~n24246;
  assign n41954 = n24251 | ~n24252;
  assign n41955 = n24257 | ~n24258;
  assign n41956 = n24260 | ~n24261;
  assign n41957 = n24271 | n24272;
  assign n41958 = n24275 | n24276;
  assign n41959 = n24277 | n24278;
  assign n41960 = n24284 | ~n24285;
  assign n41961 = n24290 | ~n24291;
  assign n41962 = n24294 | n24295;
  assign n41963 = n24298 | ~n24299;
  assign n41964 = n24307 | ~n24308;
  assign n41965 = n24318 | n24319;
  assign n41966 = n24322 | n24323;
  assign n41967 = n24324 | n24325;
  assign n41968 = n24331 | ~n24332;
  assign n41969 = n24334 | ~n24335;
  assign n41970 = n24345 | n24346;
  assign n41971 = n24349 | n24350;
  assign n41972 = n24351 | n24352;
  assign n41973 = n24367 | n24368;
  assign n41974 = n24371 | n24372;
  assign n41975 = n24373 | n24374;
  assign n41976 = n24380 | ~n24381;
  assign n41977 = n24391 | n24392;
  assign n41978 = n24395 | n24396;
  assign n41979 = n24397 | n24398;
  assign n41980 = n24410 | ~n24411;
  assign n41981 = n24416 | ~n24417;
  assign n41982 = n24422 | n24423;
  assign n41983 = n24427 | n24428;
  assign n41984 = n24429 | ~n24430;
  assign n41985 = n24438 | n24439;
  assign n41986 = n24442 | ~n24443;
  assign n41987 = n24449 | n24450;
  assign n41988 = n24451 | n24452;
  assign n41989 = n24453 | ~n24454;
  assign n41990 = n24457 | n24458;
  assign n41991 = n24459 | n24460;
  assign n41992 = n24461 | ~n24462;
  assign n41993 = n24467 | ~n24468;
  assign n41994 = n24473 | n24474;
  assign n41995 = n24478 | n24479;
  assign n41996 = n24480 | ~n24481;
  assign n41997 = n24487 | ~n24488;
  assign n41998 = n24490 | n24491;
  assign n41999 = n24492 | n24493;
  assign n42000 = n24499 | ~n24500;
  assign n42001 = n24505 | ~n24506;
  assign n42002 = n24511 | ~n24512;
  assign n42003 = n24515 | n24516;
  assign n42004 = n24526 | n24527;
  assign n42005 = n24530 | n24531;
  assign n42006 = n24532 | n24533;
  assign n42007 = n24545 | n24546;
  assign n42008 = n24549 | n24550;
  assign n42009 = n24551 | n24552;
  assign n42010 = n24564 | n24565;
  assign n42011 = n24568 | n24569;
  assign n42012 = n24570 | n24571;
  assign n42013 = n24580 | n24581;
  assign n42014 = n24584 | n24585;
  assign n42015 = n24586 | n24587;
  assign n42016 = n24596 | n24597;
  assign n42017 = n24600 | n24601;
  assign n42018 = n24602 | n24603;
  assign n42019 = n24612 | n24613;
  assign n42020 = n24616 | n24617;
  assign n42021 = n24618 | n24619;
  assign n42022 = n24628 | n24629;
  assign n42023 = n24632 | n24633;
  assign n42024 = n24634 | n24635;
  assign n42025 = n24644 | n24645;
  assign n42026 = n24648 | n24649;
  assign n42027 = n24650 | n24651;
  assign n42028 = n24660 | n24661;
  assign n42029 = n24664 | n24665;
  assign n42030 = n24666 | n24667;
  assign n42031 = n24673 | ~n24674;
  assign n42032 = n24683 | n24684;
  assign n42033 = n24685 | n24686;
  assign n42034 = n24687 | ~n24688;
  assign n42035 = n24691 | n24692;
  assign n42036 = n24693 | n24694;
  assign n42037 = n24695 | ~n24696;
  assign n42038 = n24701 | ~n24702;
  assign n42039 = n24704 | ~n24705;
  assign n42040 = n24715 | n24716;
  assign n42041 = n24719 | n24720;
  assign n42042 = n24721 | n24722;
  assign n42043 = n24726 | n24727;
  assign n42044 = n24728 | n24729;
  assign n42045 = n24730 | ~n24731;
  assign n42046 = n24737 | n24738;
  assign n42047 = n24739 | n24740;
  assign n42048 = n24741 | ~n24742;
  assign n42049 = n24745 | n24746;
  assign n42050 = n24747 | n24748;
  assign n42051 = n24749 | ~n24750;
  assign n42052 = n24755 | ~n24756;
  assign n42053 = n24766 | n24767;
  assign n42054 = n24770 | n24771;
  assign n42055 = n24772 | n24773;
  assign n42056 = n24779 | ~n24780;
  assign n42057 = n24784 | n24785;
  assign n42058 = n24786 | ~n24787;
  assign n42059 = n24788 | n24789;
  assign n42060 = n24790 | n24791;
  assign n42061 = n24797 | ~n24798;
  assign n42062 = n24803 | ~n24804;
  assign n42063 = n24809 | n24810;
  assign n42064 = n24820 | n24821;
  assign n42065 = n24824 | n24825;
  assign n42066 = n24826 | n24827;
  assign n42067 = n24831 | n24832;
  assign n42068 = n24833 | n24834;
  assign n42069 = n24835 | ~n24836;
  assign n42070 = n24841 | ~n24842;
  assign n42071 = n24847 | ~n24848;
  assign n42072 = n24858 | n24859;
  assign n42073 = n24862 | n24863;
  assign n42074 = n24864 | n24865;
  assign n42075 = n24868 | ~n24869;
  assign n42076 = n24872 | n24873;
  assign n42077 = n24874 | n24875;
  assign n42078 = n24876 | ~n24877;
  assign n42079 = n24888 | n24889;
  assign n42080 = n24892 | n24893;
  assign n42081 = n24894 | n24895;
  assign n42082 = n24901 | ~n24902;
  assign n42083 = n24904 | n24905;
  assign n42084 = n24909 | n24910;
  assign n42085 = n24911 | ~n24912;
  assign n42086 = n24923 | n24924;
  assign n42087 = n24927 | n24928;
  assign n42088 = n24929 | n24930;
  assign n42089 = n24934 | n24935;
  assign n42090 = n24936 | n24937;
  assign n42091 = n24938 | ~n24939;
  assign n42092 = n24941 | n24942;
  assign n42093 = n24944 | n24945;
  assign n42094 = n24949 | n24946 | n24948;
  assign n42095 = n24950 | ~n24951;
  assign n42096 = n24962 | n24963;
  assign n42097 = n24966 | n24967;
  assign n42098 = n24968 | n24969;
  assign n42099 = n24975 | ~n24976;
  assign n42100 = n24978 | n24979;
  assign n42101 = n24983 | n24984;
  assign n42102 = n24985 | ~n24986;
  assign n42103 = n24994 | n24995;
  assign n42104 = n24998 | n24999;
  assign n42105 = n25000 | n25001;
  assign n42106 = n25005 | n25006;
  assign n42107 = n25007 | n25008;
  assign n42108 = n25009 | ~n25010;
  assign n42109 = n25015 | ~n25016;
  assign n42110 = n25021 | ~n25022;
  assign n42111 = n25025 | n25026;
  assign n42112 = n25036 | n25037;
  assign n42113 = n25040 | n25041;
  assign n42114 = n25042 | n25043;
  assign n42115 = n25048 | n25049;
  assign n42116 = n25050 | n25051;
  assign n42117 = n25052 | ~n25053;
  assign n42118 = n25061 | n25062;
  assign n42119 = n25065 | ~n25066;
  assign n42120 = n25080 | n25081;
  assign n42121 = n25084 | ~n25085;
  assign n42122 = n25091 | n25092;
  assign n42123 = n25093 | n25094;
  assign n42124 = n25095 | ~n25096;
  assign n42125 = n25104 | n25105;
  assign n42126 = n25108 | n25109;
  assign n42127 = n25110 | n25111;
  assign n42128 = n25120 | n25121;
  assign n42129 = n25124 | n25125;
  assign n42130 = n25126 | n25127;
  assign n42131 = n25136 | n25137;
  assign n42132 = n25140 | n25141;
  assign n42133 = n25142 | n25143;
  assign n42134 = n25151 | n25152;
  assign n42135 = n25155 | n25156;
  assign n42136 = n25157 | n25158;
  assign n42137 = n25171 | n25172;
  assign n42138 = n25175 | n25176;
  assign n42139 = n25177 | n25178;
  assign n42140 = n25186 | n25187;
  assign n42141 = n25188 | n25189;
  assign n42142 = n25190 | ~n25191;
  assign n42143 = n25196 | ~n25197;
  assign n42144 = n25207 | n25208;
  assign n42145 = n25211 | n25212;
  assign n42146 = n25213 | n25214;
  assign n42147 = n25220 | ~n25221;
  assign n42148 = n25231 | n25232;
  assign n42149 = n25235 | n25236;
  assign n42150 = n25237 | n25238;
  assign n42151 = n25244 | ~n25245;
  assign n42152 = n25255 | n25256;
  assign n42153 = n25259 | n25260;
  assign n42154 = n25261 | n25262;
  assign n42155 = n25268 | ~n25269;
  assign n42156 = n25279 | n25280;
  assign n42157 = n25283 | n25284;
  assign n42158 = n25285 | n25286;
  assign n42159 = n25295 | ~n25296;
  assign n42160 = n25299 | n25300;
  assign n42161 = n25312 | ~n25313;
  assign n42162 = n25316 | n25317;
  assign n42163 = n25323 | ~n25324;
  assign n42164 = n25327 | n25328;
  assign n42165 = n25339 | n25340;
  assign n42166 = n25343 | n25344;
  assign n42167 = n25345 | n25346;
  assign n42168 = n25352 | ~n25353;
  assign n42169 = n25358 | ~n25359;
  assign n42170 = n25366 | n25367;
  assign n42171 = n25370 | n25371;
  assign n42172 = n25372 | n25373;
  assign n42173 = n25378 | n25379;
  assign n42174 = n25380 | n25381;
  assign n42175 = n25382 | ~n25383;
  assign n42176 = n25388 | ~n25389;
  assign n42177 = n25391 | n25392;
  assign n42178 = n25393 | n25394;
  assign n42179 = n25396 | ~n25397;
  assign n42180 = n25402 | ~n25403;
  assign n42181 = n25411 | n25412;
  assign n42182 = n25415 | ~n25416;
  assign n42183 = n25422 | n25423;
  assign n42184 = n25424 | n25425;
  assign n42185 = n25426 | ~n25427;
  assign n42186 = n25432 | ~n25433;
  assign n42187 = n25440 | n25441;
  assign n42188 = n25444 | n25445;
  assign n42189 = n25446 | n25447;
  assign n42190 = n25452 | n25453;
  assign n42191 = n25454 | n25455;
  assign n42192 = n25456 | ~n25457;
  assign n42193 = n25462 | ~n25463;
  assign n42194 = n25471 | ~n25472;
  assign n42195 = n25478 | n25479;
  assign n42196 = n25480 | n25481;
  assign n42197 = n25482 | ~n25483;
  assign n42198 = n25489 | n25486 | n25488;
  assign n42199 = n25495 | ~n25496;
  assign n42200 = n25499 | n25500;
  assign n42201 = n25510 | n25511;
  assign n42202 = n25514 | n25515;
  assign n42203 = n25516 | n25517;
  assign n42204 = n25529 | n25530;
  assign n42205 = n25533 | n25534;
  assign n42206 = n25535 | n25536;
  assign n42207 = n25539 | ~n25540;
  assign n42208 = n25550 | n25551;
  assign n42209 = n25554 | n25555;
  assign n42210 = n25556 | n25557;
  assign n42211 = n25570 | n25571;
  assign n42212 = n25574 | ~n25575;
  assign n42213 = n25588 | n25589;
  assign n42214 = n25592 | ~n25593;
  assign n42215 = n25598 | ~n25599;
  assign n42216 = n25609 | n25610;
  assign n42217 = n25613 | n25614;
  assign n42218 = n25615 | n25616;
  assign n42219 = n25625 | n25626;
  assign n42220 = n25629 | n25630;
  assign n42221 = n25631 | n25632;
  assign n42222 = n25643 | n25644;
  assign n42223 = n25647 | n25648;
  assign n42224 = n25649 | n25650;
  assign n42225 = n25659 | n25660;
  assign n42226 = n25663 | n25664;
  assign n42227 = n25665 | n25666;
  assign n42228 = n25681 | n25682;
  assign n42229 = n25685 | ~n25686;
  assign n42230 = n25702 | n25703;
  assign n42231 = n25706 | n25707;
  assign n42232 = n25708 | n25709;
  assign n42233 = n25715 | ~n25716;
  assign n42234 = n25718 | ~n25719;
  assign n42235 = n25729 | n25730;
  assign n42236 = n25733 | n25734;
  assign n42237 = n25735 | n25736;
  assign n42238 = n25742 | ~n25743;
  assign n42239 = n25751 | ~n25752;
  assign n42240 = n25762 | n25763;
  assign n42241 = n25766 | n25767;
  assign n42242 = n25768 | n25769;
  assign n42243 = n25775 | ~n25776;
  assign n42244 = n25781 | ~n25782;
  assign n42245 = n25787 | ~n25788;
  assign n42246 = n25798 | n25799;
  assign n42247 = n25802 | n25803;
  assign n42248 = n25804 | n25805;
  assign n42249 = n25811 | ~n25812;
  assign n42250 = n25822 | n25823;
  assign n42251 = n25826 | n25827;
  assign n42252 = n25828 | n25829;
  assign n42253 = n25847 | ~n25848;
  assign n42254 = n25853 | ~n25854;
  assign n42255 = n25856 | n25857;
  assign n42256 = n25858 | n25859;
  assign n42257 = n25861 | ~n25862;
  assign n42258 = n25865 | n25866;
  assign n42259 = n25867 | n25868;
  assign n42260 = n25869 | ~n25870;
  assign n42261 = n25875 | n25876;
  assign n42262 = n25880 | n25881;
  assign n42263 = n25882 | ~n25883;
  assign n42264 = n25891 | n25892;
  assign n42265 = n25895 | ~n25896;
  assign n42266 = n25902 | n25903;
  assign n42267 = n25904 | n25905;
  assign n42268 = n25906 | ~n25907;
  assign n42269 = n25913 | n25910 | n25912;
  assign n42270 = n25920 | ~n25921;
  assign n42271 = n25923 | n25924;
  assign n42272 = n25925 | n25926;
  assign n42273 = n25932 | ~n25933;
  assign n42274 = n25950 | n25951;
  assign n42275 = n25954 | n25955;
  assign n42276 = n25956 | n25957;
  assign n42277 = n25969 | n25970;
  assign n42278 = n25973 | n25974;
  assign n42279 = n25975 | n25976;
  assign n42280 = n25979 | ~n25980;
  assign n42281 = n25990 | n25991;
  assign n42282 = n25994 | n25995;
  assign n42283 = n25996 | n25997;
  assign n42284 = n26000 | ~n26001;
  assign n42285 = n26012 | n26013;
  assign n42286 = n26016 | n26017;
  assign n42287 = n26018 | n26019;
  assign n42288 = n26028 | n26029;
  assign n42289 = n26032 | n26033;
  assign n42290 = n26034 | n26035;
  assign n42291 = n26044 | n26045;
  assign n42292 = n26048 | n26049;
  assign n42293 = n26050 | n26051;
  assign n42294 = n26061 | n26062;
  assign n42295 = n26065 | n26066;
  assign n42296 = n26067 | n26068;
  assign n42297 = n26075 | n26076;
  assign n42298 = n26077 | n26078;
  assign n42299 = n26079 | ~n26080;
  assign n42300 = n26085 | ~n26086;
  assign n42301 = n26089 | n26090;
  assign n42302 = n26091 | n26092;
  assign n42303 = n26093 | ~n26094;
  assign n42304 = n26104 | n26105;
  assign n42305 = n26108 | n26109;
  assign n42306 = n26110 | n26111;
  assign n42307 = n26115 | n26116;
  assign n42308 = n26117 | n26118;
  assign n42309 = n26119 | ~n26120;
  assign n42310 = n26122 | ~n26123;
  assign n42311 = n26133 | n26134;
  assign n42312 = n26137 | n26138;
  assign n42313 = n26139 | n26140;
  assign n42314 = n26150 | n26147 | n26149;
  assign n42315 = n26151 | n26152;
  assign n42316 = n26154 | ~n26155;
  assign n42317 = n26156 | n26157;
  assign n42318 = n26158 | ~n26159;
  assign n42319 = n26164 | ~n26165;
  assign n42320 = n26175 | n26176;
  assign n42321 = n26179 | n26180;
  assign n42322 = n26181 | n26182;
  assign n42323 = n26186 | n26187;
  assign n42324 = n26188 | n26189;
  assign n42325 = n26190 | ~n26191;
  assign n42326 = n26193 | ~n26194;
  assign n42327 = n26204 | n26205;
  assign n42328 = n26208 | n26209;
  assign n42329 = n26210 | n26211;
  assign n42330 = n26215 | n26216;
  assign n42331 = n26217 | n26218;
  assign n42332 = n26219 | ~n26220;
  assign n42333 = n26222 | ~n26223;
  assign n42334 = n26228 | ~n26229;
  assign n42335 = n26234 | ~n26235;
  assign n42336 = n26245 | n26246;
  assign n42337 = n26249 | n26250;
  assign n42338 = n26251 | n26252;
  assign n42339 = n26256 | n26257;
  assign n42340 = n26258 | n26259;
  assign n42341 = n26260 | ~n26261;
  assign n42342 = n26266 | ~n26267;
  assign n42343 = n26280 | n26281;
  assign n42344 = n26284 | n26285;
  assign n42345 = n26286 | n26287;
  assign n42346 = n26291 | n26292;
  assign n42347 = n26293 | n26294;
  assign n42348 = n26295 | ~n26296;
  assign n42349 = n26298 | ~n26299;
  assign n42350 = n26309 | n26310;
  assign n42351 = n26313 | n26314;
  assign n42352 = n26315 | n26316;
  assign n42353 = n26319 | ~n26320;
  assign n42354 = n26323 | n26324;
  assign n42355 = n26325 | n26326;
  assign n42356 = n26327 | ~n26328;
  assign n42357 = n26333 | n26334;
  assign n42358 = n26338 | n26339;
  assign n42359 = n26340 | ~n26341;
  assign n42360 = n26352 | n26353;
  assign n42361 = n26356 | n26357;
  assign n42362 = n26358 | n26359;
  assign n42363 = n26365 | ~n26366;
  assign n42364 = n26368 | n26369;
  assign n42365 = n26371 | n26372;
  assign n42366 = n26376 | n26373 | n26375;
  assign n42367 = n26377 | ~n26378;
  assign n42368 = n26389 | n26390;
  assign n42369 = n26393 | n26394;
  assign n42370 = n26395 | n26396;
  assign n42371 = n26400 | n26401;
  assign n42372 = n26402 | n26403;
  assign n42373 = n26404 | ~n26405;
  assign n42374 = n26407 | n26408;
  assign n42375 = n26412 | n26413;
  assign n42376 = n26414 | ~n26415;
  assign n42377 = n26431 | ~n26432;
  assign n42378 = n26445 | n26446;
  assign n42379 = n26449 | n26450;
  assign n42380 = n26451 | n26452;
  assign n42381 = n26465 | n26466;
  assign n42382 = n26469 | ~n26470;
  assign n42383 = n26483 | n26484;
  assign n42384 = n26487 | n26488;
  assign n42385 = n26489 | n26490;
  assign n42386 = n26502 | n26503;
  assign n42387 = n26506 | n26507;
  assign n42388 = n26508 | n26509;
  assign n42389 = n26523 | n26524;
  assign n42390 = n26527 | n26528;
  assign n42391 = n26529 | n26530;
  assign n42392 = n26539 | n26540;
  assign n42393 = n26543 | n26544;
  assign n42394 = n26545 | n26546;
  assign n42395 = n26556 | n26557;
  assign n42396 = n26560 | n26561;
  assign n42397 = n26562 | n26563;
  assign n42398 = n26580 | n26581;
  assign n42399 = n26584 | ~n26585;
  assign n42400 = n26601 | n26602;
  assign n42401 = n26605 | n26606;
  assign n42402 = n26607 | n26608;
  assign n42403 = n26614 | ~n26615;
  assign n42404 = n26625 | n26626;
  assign n42405 = n26629 | n26630;
  assign n42406 = n26631 | n26632;
  assign n42407 = n26638 | ~n26639;
  assign n42408 = n26644 | ~n26645;
  assign n42409 = n26659 | n26660;
  assign n42410 = n26663 | n26664;
  assign n42411 = n26665 | n26666;
  assign n42412 = n26672 | ~n26673;
  assign n42413 = n26683 | n26684;
  assign n42414 = n26687 | n26688;
  assign n42415 = n26689 | n26690;
  assign n42416 = n26699 | ~n26700;
  assign n42417 = n26703 | n26704;
  assign n42418 = n26710 | ~n26711;
  assign n42419 = n26714 | n26715;
  assign n42420 = n26726 | n26727;
  assign n42421 = n26730 | n26731;
  assign n42422 = n26732 | n26733;
  assign n42423 = n26739 | ~n26740;
  assign n42424 = n26750 | n26751;
  assign n42425 = n26754 | n26755;
  assign n42426 = n26756 | n26757;
  assign n42427 = n26763 | ~n26764;
  assign n42428 = n26774 | n26775;
  assign n42429 = n26778 | n26779;
  assign n42430 = n26780 | n26781;
  assign n42431 = n26786 | n26787;
  assign n42432 = n26788 | n26789;
  assign n42433 = n26790 | ~n26791;
  assign n42434 = n26793 | n26794;
  assign n42435 = n26798 | n26799;
  assign n42436 = n26800 | ~n26801;
  assign n42437 = n26806 | n26807;
  assign n42438 = n26811 | n26812;
  assign n42439 = n26813 | ~n26814;
  assign n42440 = n26819 | n26820;
  assign n42441 = n26824 | n26822 | n26823;
  assign n42442 = n26825 | n26826;
  assign n42443 = n26842 | n26843;
  assign n42444 = n26846 | n26847;
  assign n42445 = n26848 | n26849;
  assign n42446 = n26861 | n26862;
  assign n42447 = n26865 | n26866;
  assign n42448 = n26867 | n26868;
  assign n42449 = n26880 | n26881;
  assign n42450 = n26884 | n26885;
  assign n42451 = n26886 | n26887;
  assign n42452 = n26890 | ~n26891;
  assign n42453 = n26901 | n26902;
  assign n42454 = n26905 | n26906;
  assign n42455 = n26907 | n26908;
  assign n42456 = n26917 | n26918;
  assign n42457 = n26921 | n26922;
  assign n42458 = n26923 | n26924;
  assign n42459 = n26933 | n26934;
  assign n42460 = n26937 | n26938;
  assign n42461 = n26939 | n26940;
  assign n42462 = n26944 | n26945;
  assign n42463 = n26952 | n26953;
  assign n42464 = n26956 | n26957;
  assign n42465 = n26958 | n26959;
  assign n42466 = n26968 | n26969;
  assign n42467 = n26972 | n26973;
  assign n42468 = n26974 | n26975;
  assign n42469 = n26984 | n26985;
  assign n42470 = n26988 | n26989;
  assign n42471 = n26990 | n26991;
  assign n42472 = n27000 | n27001;
  assign n42473 = n27006 | ~n27007;
  assign n42474 = n27017 | n27018;
  assign n42475 = n27021 | n27022;
  assign n42476 = n27023 | n27024;
  assign n42477 = n27030 | ~n27031;
  assign n42478 = n27039 | ~n27040;
  assign n42479 = n27050 | n27051;
  assign n42480 = n27054 | n27055;
  assign n42481 = n27056 | n27057;
  assign n42482 = n27063 | ~n27064;
  assign n42483 = n27069 | ~n27070;
  assign n42484 = n27075 | ~n27076;
  assign n42485 = n27086 | n27087;
  assign n42486 = n27090 | n27091;
  assign n42487 = n27092 | n27093;
  assign n42488 = n27099 | ~n27100;
  assign n42489 = n27105 | ~n27106;
  assign n42490 = n27111 | ~n27112;
  assign n42491 = n27126 | ~n27127;
  assign n42492 = n27137 | n27138;
  assign n42493 = n27141 | n27142;
  assign n42494 = n27143 | n27144;
  assign n42495 = n27150 | ~n27151;
  assign n42496 = n27161 | n27162;
  assign n42497 = n27165 | n27166;
  assign n42498 = n27167 | n27168;
  assign n42499 = n27173 | n27174;
  assign n42500 = n27175 | n27176;
  assign n42501 = n27177 | ~n27178;
  assign n42502 = n27180 | n27181;
  assign n42503 = n27185 | n27186;
  assign n42504 = n27187 | ~n27188;
  assign n42505 = n27198 | n27199;
  assign n42506 = n27202 | n27203;
  assign n42507 = n27204 | n27205;
  assign n42508 = n27210 | n27211;
  assign n42509 = n27212 | n27213;
  assign n42510 = n27214 | ~n27215;
  assign n42511 = n27217 | n27218;
  assign n42512 = n27220 | n27221;
  assign n42513 = n27225 | n27222 | n27224;
  assign n42514 = n27226 | ~n27227;
  assign n42515 = n27236 | ~n27237;
  assign n42516 = n27239 | n27240;
  assign n42517 = n27241 | n27242;
  assign n42518 = n27248 | ~n27249;
  assign n42519 = n27254 | ~n27255;
  assign n42520 = n27260 | ~n27261;
  assign n42521 = n27264 | n27265;
  assign n42522 = n27276 | n27277;
  assign n42523 = n27280 | n27281;
  assign n42524 = n27282 | n27283;
  assign n42525 = n27287 | n27288;
  assign n42526 = n27289 | n27290;
  assign n42527 = n27291 | ~n27292;
  assign n42528 = n27299 | n27300;
  assign n42529 = n27303 | n27304;
  assign n42530 = n27305 | n27306;
  assign n42531 = n27318 | n27319;
  assign n42532 = n27322 | n27323;
  assign n42533 = n27324 | n27325;
  assign n42534 = n27337 | n27338;
  assign n42535 = n27341 | n27342;
  assign n42536 = n27343 | n27344;
  assign n42537 = n27358 | n27359;
  assign n42538 = n27362 | n27363;
  assign n42539 = n27364 | n27365;
  assign n42540 = n27374 | n27375;
  assign n42541 = n27378 | n27379;
  assign n42542 = n27380 | n27381;
  assign n42543 = n27391 | n27392;
  assign n42544 = n27395 | n27396;
  assign n42545 = n27397 | n27398;
  assign n42546 = n27406 | n27407;
  assign n42547 = n27410 | n27411;
  assign n42548 = n27412 | n27413;
  assign n42549 = n27426 | n27427;
  assign n42550 = n27428 | n27429;
  assign n42551 = n27430 | ~n27431;
  assign n42552 = n27436 | ~n27437;
  assign n42553 = n27450 | n27451;
  assign n42554 = n27454 | n27455;
  assign n42555 = n27456 | n27457;
  assign n42556 = n27461 | n27462;
  assign n42557 = n27463 | n27464;
  assign n42558 = n27465 | ~n27466;
  assign n42559 = n27476 | n27477;
  assign n42560 = n27480 | n27481;
  assign n42561 = n27482 | n27483;
  assign n42562 = n27487 | n27488;
  assign n42563 = n27489 | n27490;
  assign n42564 = n27491 | ~n27492;
  assign n42565 = n27494 | ~n27495;
  assign n42566 = n27505 | n27506;
  assign n42567 = n27509 | n27510;
  assign n42568 = n27511 | n27512;
  assign n42569 = n27515 | ~n27516;
  assign n42570 = n27524 | ~n27525;
  assign n42571 = n27530 | ~n27531;
  assign n42572 = n27541 | n27542;
  assign n42573 = n27545 | n27546;
  assign n42574 = n27547 | n27548;
  assign n42575 = n27552 | n27553;
  assign n42576 = n27554 | n27555;
  assign n42577 = n27556 | ~n27557;
  assign n42578 = n27562 | ~n27563;
  assign n42579 = n27576 | n27577;
  assign n42580 = n27580 | n27581;
  assign n42581 = n27582 | n27583;
  assign n42582 = n27587 | n27588;
  assign n42583 = n27589 | n27590;
  assign n42584 = n27591 | ~n27592;
  assign n42585 = n27602 | n27603;
  assign n42586 = n27606 | n27607;
  assign n42587 = n27608 | n27609;
  assign n42588 = n27613 | n27614;
  assign n42589 = n27615 | n27616;
  assign n42590 = n27617 | ~n27618;
  assign n42591 = n27620 | ~n27621;
  assign n42592 = n27631 | n27632;
  assign n42593 = n27635 | n27636;
  assign n42594 = n27637 | n27638;
  assign n42595 = n27648 | ~n27649;
  assign n42596 = n27651 | n27652;
  assign n42597 = n27653 | n27654;
  assign n42598 = n27656 | ~n27657;
  assign n42599 = n27660 | n27661;
  assign n42600 = n27662 | n27663;
  assign n42601 = n27664 | ~n27665;
  assign n42602 = n27670 | ~n27671;
  assign n42603 = n27676 | ~n27677;
  assign n42604 = n27682 | ~n27683;
  assign n42605 = n27686 | n27687;
  assign n42606 = n27697 | ~n27698;
  assign n42607 = n27703 | ~n27704;
  assign n42608 = n27707 | n27708;
  assign n42609 = n27709 | n27710;
  assign n42610 = n27711 | ~n27712;
  assign n42611 = n27719 | n27720;
  assign n42612 = n27723 | n27724;
  assign n42613 = n27725 | n27726;
  assign n42614 = n27729 | ~n27730;
  assign n42615 = n27740 | n27741;
  assign n42616 = n27744 | n27745;
  assign n42617 = n27746 | n27747;
  assign n42618 = n27750 | ~n27751;
  assign n42619 = n27761 | n27762;
  assign n42620 = n27765 | n27766;
  assign n42621 = n27767 | n27768;
  assign n42622 = n27771 | n27772;
  assign n42623 = n27782 | n27783;
  assign n42624 = n27786 | n27787;
  assign n42625 = n27788 | n27789;
  assign n42626 = n27804 | n27805;
  assign n42627 = n27808 | n27809;
  assign n42628 = n27810 | n27811;
  assign n42629 = n27821 | n27822;
  assign n42630 = n27825 | n27826;
  assign n42631 = n27827 | n27828;
  assign n42632 = n27844 | n27845;
  assign n42633 = n27848 | n27849;
  assign n42634 = n27850 | n27851;
  assign n42635 = n27866 | n27867;
  assign n42636 = n27870 | n27871;
  assign n42637 = n27872 | n27873;
  assign n42638 = n27879 | ~n27880;
  assign n42639 = n27885 | ~n27886;
  assign n42640 = n27900 | n27901;
  assign n42641 = n27904 | n27905;
  assign n42642 = n27906 | n27907;
  assign n42643 = n27913 | ~n27914;
  assign n42644 = n27924 | n27925;
  assign n42645 = n27928 | n27929;
  assign n42646 = n27930 | n27931;
  assign n42647 = n27937 | ~n27938;
  assign n42648 = n27940 | ~n27941;
  assign n42649 = n27951 | n27952;
  assign n42650 = n27955 | n27956;
  assign n42651 = n27957 | n27958;
  assign n42652 = n27967 | ~n27968;
  assign n42653 = n27971 | n27972;
  assign n42654 = n27983 | n27984;
  assign n42655 = n27987 | n27988;
  assign n42656 = n27989 | n27990;
  assign n42657 = n27996 | ~n27997;
  assign n42658 = n28007 | n28008;
  assign n42659 = n28011 | n28012;
  assign n42660 = n28013 | n28014;
  assign n42661 = n28020 | ~n28021;
  assign n42662 = n28031 | n28032;
  assign n42663 = n28035 | n28036;
  assign n42664 = n28037 | n28038;
  assign n42665 = n28044 | ~n28045;
  assign n42666 = n28050 | n28051;
  assign n42667 = n28055 | n28056;
  assign n42668 = n28057 | ~n28058;
  assign n42669 = n28063 | n28064;
  assign n42670 = n28068 | n28069;
  assign n42671 = n28070 | ~n28071;
  assign n42672 = n28077 | n28074 | n28076;
  assign n42673 = n28083 | ~n28084;
  assign n42674 = n28087 | n28088;
  assign n42675 = n28096 | ~n28097;
  assign n42676 = n28099 | n28100;
  assign n42677 = n28101 | n28102;
  assign n42678 = n28105 | ~n28106;
  assign n42679 = n28111 | ~n28112;
  assign n42680 = n28119 | n28120;
  assign n42681 = n28123 | n28124;
  assign n42682 = n28125 | n28126;
  assign n42683 = n28131 | n28132;
  assign n42684 = n28133 | n28134;
  assign n42685 = n28135 | ~n28136;
  assign n42686 = n28143 | n28144;
  assign n42687 = n28147 | n28148;
  assign n42688 = n28149 | n28150;
  assign n42689 = n28162 | n28163;
  assign n42690 = n28166 | n28167;
  assign n42691 = n28168 | n28169;
  assign n42692 = n28172 | ~n28173;
  assign n42693 = n28183 | n28184;
  assign n42694 = n28187 | n28188;
  assign n42695 = n28189 | n28190;
  assign n42696 = n28199 | n28200;
  assign n42697 = n28203 | n28204;
  assign n42698 = n28205 | n28206;
  assign n42699 = n28215 | n28216;
  assign n42700 = n28219 | n28220;
  assign n42701 = n28221 | n28222;
  assign n42702 = n28230 | n28231;
  assign n42703 = n28234 | n28235;
  assign n42704 = n28236 | n28237;
  assign n42705 = n28240 | n28241;
  assign n42706 = n28248 | n28249;
  assign n42707 = n28252 | n28253;
  assign n42708 = n28254 | n28255;
  assign n42709 = n28264 | n28265;
  assign n42710 = n28268 | n28269;
  assign n42711 = n28270 | n28271;
  assign n42712 = n28286 | n28287;
  assign n42713 = n28290 | ~n28291;
  assign n42714 = n28305 | n28306;
  assign n42715 = n28316 | n28317;
  assign n42716 = n28320 | n28321;
  assign n42717 = n28322 | n28323;
  assign n42718 = n28329 | ~n28330;
  assign n42719 = n28335 | ~n28336;
  assign n42720 = n28341 | ~n28342;
  assign n42721 = n28350 | ~n28351;
  assign n42722 = n28371 | ~n28372;
  assign n42723 = n28382 | n28383;
  assign n42724 = n28386 | n28387;
  assign n42725 = n28388 | n28389;
  assign n42726 = n28395 | ~n28396;
  assign n42727 = n28398 | ~n28399;
  assign n42728 = n28409 | n28410;
  assign n42729 = n28413 | n28414;
  assign n42730 = n28415 | n28416;
  assign n42731 = n28422 | n28423;
  assign n42732 = n28427 | n28428;
  assign n42733 = n28429 | ~n28430;
  assign n42734 = n28437 | n28438;
  assign n42735 = n28441 | n28442;
  assign n42736 = n28443 | n28444;
  assign n42737 = n28449 | n28450;
  assign n42738 = n28451 | n28452;
  assign n42739 = n28453 | ~n28454;
  assign n42740 = n28459 | ~n28460;
  assign n42741 = n28462 | n28463;
  assign n42742 = n28464 | n28465;
  assign n42743 = n28467 | ~n28468;
  assign n42744 = n28473 | ~n28474;
  assign n42745 = n28491 | n28492;
  assign n42746 = n28495 | n28496;
  assign n42747 = n28497 | n28498;
  assign n42748 = n28501 | ~n28502;
  assign n42749 = n28512 | n28513;
  assign n42750 = n28516 | n28517;
  assign n42751 = n28518 | n28519;
  assign n42752 = n28536 | n28537;
  assign n42753 = n28540 | n28541;
  assign n42754 = n28542 | n28543;
  assign n42755 = n28546 | n28547;
  assign n42756 = n28555 | n28556;
  assign n42757 = n28559 | n28560;
  assign n42758 = n28561 | n28562;
  assign n42759 = n28580 | n28581;
  assign n42760 = n28584 | n28585;
  assign n42761 = n28586 | n28587;
  assign n42762 = n28591 | n28592;
  assign n42763 = n28593 | n28594;
  assign n42764 = n28595 | ~n28596;
  assign n42765 = n28601 | ~n28602;
  assign n42766 = n28605 | n28606;
  assign n42767 = n28607 | n28608;
  assign n42768 = n28609 | ~n28610;
  assign n42769 = n28620 | n28621;
  assign n42770 = n28624 | n28625;
  assign n42771 = n28626 | n28627;
  assign n42772 = n28631 | n28632;
  assign n42773 = n28633 | n28634;
  assign n42774 = n28635 | ~n28636;
  assign n42775 = n28646 | n28647;
  assign n42776 = n28650 | n28651;
  assign n42777 = n28652 | n28653;
  assign n42778 = n28656 | ~n28657;
  assign n42779 = n28665 | ~n28666;
  assign n42780 = n28679 | n28680;
  assign n42781 = n28683 | n28684;
  assign n42782 = n28685 | n28686;
  assign n42783 = n28690 | n28691;
  assign n42784 = n28692 | n28693;
  assign n42785 = n28694 | ~n28695;
  assign n42786 = n28705 | n28706;
  assign n42787 = n28709 | n28710;
  assign n42788 = n28711 | n28712;
  assign n42789 = n28716 | n28717;
  assign n42790 = n28718 | n28719;
  assign n42791 = n28720 | ~n28721;
  assign n42792 = n28731 | n28732;
  assign n42793 = n28735 | n28736;
  assign n42794 = n28737 | n28738;
  assign n42795 = n28742 | n28743;
  assign n42796 = n28744 | n28745;
  assign n42797 = n28746 | ~n28747;
  assign n42798 = n28757 | n28758;
  assign n42799 = n28761 | n28762;
  assign n42800 = n28763 | n28764;
  assign n42801 = n28768 | n28769;
  assign n42802 = n28770 | n28771;
  assign n42803 = n28772 | ~n28773;
  assign n42804 = n28775 | ~n28776;
  assign n42805 = n28786 | n28787;
  assign n42806 = n28790 | n28791;
  assign n42807 = n28792 | n28793;
  assign n42808 = n28803 | n28800 | n28802;
  assign n42809 = n28804 | n28805;
  assign n42810 = n28807 | ~n28808;
  assign n42811 = n28809 | n28810;
  assign n42812 = n28811 | ~n28812;
  assign n42813 = n28823 | n28824;
  assign n42814 = n28827 | n28828;
  assign n42815 = n28829 | n28830;
  assign n42816 = n28836 | ~n28837;
  assign n42817 = n28839 | n28840;
  assign n42818 = n28844 | n28845;
  assign n42819 = n28846 | ~n28847;
  assign n42820 = n28858 | n28859;
  assign n42821 = n28862 | n28863;
  assign n42822 = n28864 | n28865;
  assign n42823 = n28869 | n28870;
  assign n42824 = n28871 | n28872;
  assign n42825 = n28873 | ~n28874;
  assign n42826 = n28876 | n28877;
  assign n42827 = n28879 | n28880;
  assign n42828 = n28884 | n28881 | n28883;
  assign n42829 = n28885 | ~n28886;
  assign n42830 = n28902 | ~n28903;
  assign n42831 = n28916 | n28917;
  assign n42832 = n28920 | n28921;
  assign n42833 = n28922 | n28923;
  assign n42834 = n28936 | n28937;
  assign n42835 = n28940 | ~n28941;
  assign n42836 = n28954 | n28955;
  assign n42837 = n28958 | n28959;
  assign n42838 = n28960 | n28961;
  assign n42839 = n28967 | ~n28968;
  assign n42840 = n28979 | n28980;
  assign n42841 = n28983 | n28984;
  assign n42842 = n28985 | n28986;
  assign n42843 = n28997 | n28998;
  assign n42844 = n29001 | n29002;
  assign n42845 = n29003 | n29004;
  assign n42846 = n29020 | n29021;
  assign n42847 = n29024 | ~n29025;
  assign n42848 = n29047 | n29048;
  assign n42849 = n29051 | n29052;
  assign n42850 = n29053 | n29054;
  assign n42851 = n29060 | ~n29061;
  assign n42852 = n29071 | n29072;
  assign n42853 = n29075 | n29076;
  assign n42854 = n29077 | n29078;
  assign n42855 = n29084 | ~n29085;
  assign n42856 = n29087 | ~n29088;
  assign n42857 = n29098 | n29099;
  assign n42858 = n29102 | n29103;
  assign n42859 = n29104 | n29105;
  assign n42860 = n29114 | ~n29115;
  assign n42861 = n29118 | n29119;
  assign n42862 = n29130 | n29131;
  assign n42863 = n29134 | n29135;
  assign n42864 = n29136 | n29137;
  assign n42865 = n29143 | ~n29144;
  assign n42866 = n29154 | n29155;
  assign n42867 = n29158 | n29159;
  assign n42868 = n29160 | n29161;
  assign n42869 = n29167 | ~n29168;
  assign n42870 = n29178 | n29179;
  assign n42871 = n29182 | n29183;
  assign n42872 = n29184 | n29185;
  assign n42873 = n29191 | ~n29192;
  assign n42874 = n29202 | n29203;
  assign n42875 = n29206 | n29207;
  assign n42876 = n29208 | n29209;
  assign n42877 = n29215 | ~n29216;
  assign n42878 = n29221 | n29222;
  assign n42879 = n29226 | n29227;
  assign n42880 = n29228 | ~n29229;
  assign n42881 = n29234 | n29235;
  assign n42882 = n29239 | n29237 | n29238;
  assign n42883 = n29240 | n29241;
  assign n42884 = n29256 | ~n29257;
  assign n42885 = n29259 | n29260;
  assign n42886 = n29261 | n29262;
  assign n42887 = n29268 | ~n29269;
  assign n42888 = n29276 | n29277;
  assign n42889 = n29280 | n29281;
  assign n42890 = n29282 | n29283;
  assign n42891 = n29295 | n29296;
  assign n42892 = n29299 | n29300;
  assign n42893 = n29301 | n29302;
  assign n42894 = n29307 | n29308;
  assign n42895 = n29309 | n29310;
  assign n42896 = n29311 | ~n29312;
  assign n42897 = n29319 | n29320;
  assign n42898 = n29323 | n29324;
  assign n42899 = n29325 | n29326;
  assign n42900 = n29329 | ~n29330;
  assign n42901 = n29340 | n29341;
  assign n42902 = n29344 | n29345;
  assign n42903 = n29346 | n29347;
  assign n42904 = n29355 | n29356;
  assign n42905 = n29359 | n29360;
  assign n42906 = n29361 | n29362;
  assign n42907 = n29371 | n29372;
  assign n42908 = n29375 | n29376;
  assign n42909 = n29377 | n29378;
  assign n42910 = n29387 | n29388;
  assign n42911 = n29391 | n29392;
  assign n42912 = n29393 | n29394;
  assign n42913 = n29410 | n29411;
  assign n42914 = n29414 | ~n29415;
  assign n42915 = n29431 | n29432;
  assign n42916 = n29435 | n29436;
  assign n42917 = n29437 | n29438;
  assign n42918 = n29444 | ~n29445;
  assign n42919 = n29455 | n29456;
  assign n42920 = n29459 | n29460;
  assign n42921 = n29461 | n29462;
  assign n42922 = n29468 | ~n29469;
  assign n42923 = n29477 | ~n29478;
  assign n42924 = n29488 | n29489;
  assign n42925 = n29492 | n29493;
  assign n42926 = n29494 | n29495;
  assign n42927 = n29501 | ~n29502;
  assign n42928 = n29507 | ~n29508;
  assign n42929 = n29513 | ~n29514;
  assign n42930 = n29522 | ~n29523;
  assign n42931 = n29533 | n29534;
  assign n42932 = n29537 | n29538;
  assign n42933 = n29539 | n29540;
  assign n42934 = n29546 | ~n29547;
  assign n42935 = n29549 | ~n29550;
  assign n42936 = n29560 | n29561;
  assign n42937 = n29564 | n29565;
  assign n42938 = n29566 | n29567;
  assign n42939 = n29573 | ~n29574;
  assign n42940 = n29579 | ~n29580;
  assign n42941 = n29585 | ~n29586;
  assign n42942 = n29591 | ~n29592;
  assign n42943 = n29597 | ~n29598;
  assign n42944 = n29603 | ~n29604;
  assign n42945 = n29609 | ~n29610;
  assign n42946 = n29612 | ~n29613;
  assign n42947 = n29618 | ~n29619;
  assign n42948 = n29622 | n29623;
  assign n42949 = n29634 | n29635;
  assign n42950 = n29638 | n29639;
  assign n42951 = n29640 | n29641;
  assign n42952 = n29645 | n29646;
  assign n42953 = n29647 | n29648;
  assign n42954 = n29649 | ~n29650;
  assign n42955 = n29657 | n29658;
  assign n42956 = n29661 | n29662;
  assign n42957 = n29663 | n29664;
  assign n42958 = n29667 | ~n29668;
  assign n42959 = n29678 | n29679;
  assign n42960 = n29682 | n29683;
  assign n42961 = n29684 | n29685;
  assign n42962 = n29695 | n29696;
  assign n42963 = n29699 | n29700;
  assign n42964 = n29701 | n29702;
  assign n42965 = n29711 | n29712;
  assign n42966 = n29715 | n29716;
  assign n42967 = n29717 | n29718;
  assign n42968 = n29736 | n29737;
  assign n42969 = n29740 | n29741;
  assign n42970 = n29742 | n29743;
  assign n42971 = n29747 | n29748;
  assign n42972 = n29749 | n29750;
  assign n42973 = n29751 | ~n29752;
  assign n42974 = n29757 | ~n29758;
  assign n42975 = n29763 | ~n29764;
  assign n42976 = n29774 | n29775;
  assign n42977 = n29778 | n29779;
  assign n42978 = n29780 | n29781;
  assign n42979 = n29796 | n29797;
  assign n42980 = n29800 | n29801;
  assign n42981 = n29802 | n29803;
  assign n42982 = n29807 | n29808;
  assign n42983 = n29809 | n29810;
  assign n42984 = n29811 | ~n29812;
  assign n42985 = n29822 | n29823;
  assign n42986 = n29826 | n29827;
  assign n42987 = n29828 | n29829;
  assign n42988 = n29833 | n29834;
  assign n42989 = n29835 | n29836;
  assign n42990 = n29837 | ~n29838;
  assign n42991 = n29840 | ~n29841;
  assign n42992 = n29851 | n29852;
  assign n42993 = n29855 | n29856;
  assign n42994 = n29857 | n29858;
  assign n42995 = n29862 | n29863;
  assign n42996 = n29864 | n29865;
  assign n42997 = n29866 | ~n29867;
  assign n42998 = n29869 | ~n29870;
  assign n42999 = n29875 | ~n29876;
  assign n43000 = n29889 | n29890;
  assign n43001 = n29893 | n29894;
  assign n43002 = n29895 | n29896;
  assign n43003 = n29900 | n29901;
  assign n43004 = n29902 | n29903;
  assign n43005 = n29904 | ~n29905;
  assign n43006 = n29907 | ~n29908;
  assign n43007 = n29918 | n29919;
  assign n43008 = n29922 | n29923;
  assign n43009 = n29924 | n29925;
  assign n43010 = n29935 | n29932 | n29934;
  assign n43011 = n29936 | n29937;
  assign n43012 = n29939 | ~n29940;
  assign n43013 = n29941 | n29942;
  assign n43014 = n29943 | ~n29944;
  assign n43015 = n29949 | ~n29950;
  assign n43016 = n29964 | n29965;
  assign n43017 = n29968 | n29969;
  assign n43018 = n29970 | n29971;
  assign n43019 = n29977 | ~n29978;
  assign n43020 = n29980 | n29981;
  assign n43021 = n29983 | n29984;
  assign n43022 = n29988 | n29985 | n29987;
  assign n43023 = n29989 | ~n29990;
  assign n43024 = n29995 | ~n29996;
  assign n43025 = n30001 | ~n30002;
  assign n43026 = n30005 | n30006;
  assign n43027 = n30017 | n30018;
  assign n43028 = n30021 | ~n30022;
  assign n43029 = n30035 | n30036;
  assign n43030 = n30039 | n30040;
  assign n43031 = n30041 | n30042;
  assign n43032 = n30054 | n30055;
  assign n43033 = n30058 | n30059;
  assign n43034 = n30060 | n30061;
  assign n43035 = n30080 | n30081;
  assign n43036 = n30084 | ~n30085;
  assign n43037 = n30101 | n30102;
  assign n43038 = n30105 | n30106;
  assign n43039 = n30107 | n30108;
  assign n43040 = n30114 | ~n30115;
  assign n43041 = n30125 | n30126;
  assign n43042 = n30129 | n30130;
  assign n43043 = n30131 | n30132;
  assign n43044 = n30138 | ~n30139;
  assign n43045 = n30149 | n30150;
  assign n43046 = n30153 | n30154;
  assign n43047 = n30155 | n30156;
  assign n43048 = n30165 | ~n30166;
  assign n43049 = n30169 | n30170;
  assign n43050 = n30181 | n30182;
  assign n43051 = n30185 | n30186;
  assign n43052 = n30187 | n30188;
  assign n43053 = n30194 | ~n30195;
  assign n43054 = n30205 | n30206;
  assign n43055 = n30209 | n30210;
  assign n43056 = n30211 | n30212;
  assign n43057 = n30218 | ~n30219;
  assign n43058 = n30229 | n30230;
  assign n43059 = n30233 | n30234;
  assign n43060 = n30235 | n30236;
  assign n43061 = n30242 | ~n30243;
  assign n43062 = n30253 | n30254;
  assign n43063 = n30257 | n30258;
  assign n43064 = n30259 | n30260;
  assign n43065 = n30266 | ~n30267;
  assign n43066 = n30272 | ~n30273;
  assign n43067 = n30286 | n30287;
  assign n43068 = n30290 | n30291;
  assign n43069 = n30292 | n30293;
  assign n43070 = n30298 | n30299;
  assign n43071 = n30300 | n30301;
  assign n43072 = n30302 | ~n30303;
  assign n43073 = n30306 | n30307;
  assign n43074 = n30308 | n30309;
  assign n43075 = n30310 | ~n30311;
  assign n43076 = n30319 | ~n30320;
  assign n43077 = n30326 | n30327;
  assign n43078 = n30328 | n30329;
  assign n43079 = n30330 | ~n30331;
  assign n43080 = n30337 | n30334 | n30336;
  assign n43081 = n30343 | ~n30344;
  assign n43082 = n30347 | n30348;
  assign n43083 = n30358 | n30359;
  assign n43084 = n30362 | n30363;
  assign n43085 = n30364 | n30365;
  assign n43086 = n30377 | n30378;
  assign n43087 = n30381 | n30382;
  assign n43088 = n30383 | n30384;
  assign n43089 = n30396 | n30397;
  assign n43090 = n30400 | n30401;
  assign n43091 = n30402 | n30403;
  assign n43092 = n30411 | n30412;
  assign n43093 = n30415 | n30416;
  assign n43094 = n30417 | n30418;
  assign n43095 = n30426 | n30427;
  assign n43096 = n30430 | n30431;
  assign n43097 = n30432 | n30433;
  assign n43098 = n30442 | n30443;
  assign n43099 = n30446 | n30447;
  assign n43100 = n30448 | n30449;
  assign n43101 = n30458 | n30459;
  assign n43102 = n30462 | n30463;
  assign n43103 = n30464 | n30465;
  assign n43104 = n30473 | n30474;
  assign n43105 = n30477 | n30478;
  assign n43106 = n30479 | n30480;
  assign n43107 = n30495 | n30496;
  assign n43108 = n30499 | ~n30500;
  assign n43109 = n30514 | ~n30515;
  assign n43110 = n30523 | ~n30524;
  assign n43111 = n30534 | n30535;
  assign n43112 = n30538 | n30539;
  assign n43113 = n30540 | n30541;
  assign n43114 = n30547 | ~n30548;
  assign n43115 = n30553 | ~n30554;
  assign n43116 = n30559 | ~n30560;
  assign n43117 = n30568 | ~n30569;
  assign n43118 = n30579 | n30580;
  assign n43119 = n30583 | n30584;
  assign n43120 = n30585 | n30586;
  assign n43121 = n30592 | ~n30593;
  assign n43122 = n30595 | ~n30596;
  assign n43123 = n30606 | n30607;
  assign n43124 = n30610 | n30611;
  assign n43125 = n30612 | n30613;
  assign n43126 = n30619 | ~n30620;
  assign n43127 = n30625 | ~n30626;
  assign n43128 = n30629 | n30630;
  assign n43129 = n30633 | ~n30634;
  assign n43130 = n30642 | ~n30643;
  assign n43131 = n30648 | ~n30649;
  assign n43132 = n30658 | ~n30659;
  assign n43133 = n30661 | n30662;
  assign n43134 = n30663 | n30664;
  assign n43135 = n30670 | ~n30671;
  assign n43136 = n30689 | n30690;
  assign n43137 = n30693 | n30694;
  assign n43138 = n30695 | n30696;
  assign n43139 = n30700 | n30701;
  assign n43140 = n30702 | n30703;
  assign n43141 = n30704 | ~n30705;
  assign n43142 = n30713 | n30714;
  assign n43143 = n30717 | n30718;
  assign n43144 = n30719 | n30720;
  assign n43145 = n30730 | n30731;
  assign n43146 = n30734 | n30735;
  assign n43147 = n30736 | n30737;
  assign n43148 = n30746 | n30747;
  assign n43149 = n30750 | n30751;
  assign n43150 = n30752 | n30753;
  assign n43151 = n30778 | n30779;
  assign n43152 = n30782 | n30783;
  assign n43153 = n30784 | n30785;
  assign n43154 = n30791 | ~n30792;
  assign n43155 = n30802 | n30803;
  assign n43156 = n30806 | n30807;
  assign n43157 = n30808 | n30809;
  assign n43158 = n30813 | n30814;
  assign n43159 = n30815 | n30816;
  assign n43160 = n30817 | ~n30818;
  assign n43161 = n30828 | n30829;
  assign n43162 = n30832 | n30833;
  assign n43163 = n30834 | n30835;
  assign n43164 = n30839 | n30840;
  assign n43165 = n30841 | n30842;
  assign n43166 = n30843 | ~n30844;
  assign n43167 = n30846 | ~n30847;
  assign n43168 = n30857 | n30858;
  assign n43169 = n30861 | n30862;
  assign n43170 = n30863 | n30864;
  assign n43171 = n30868 | n30869;
  assign n43172 = n30870 | n30871;
  assign n43173 = n30872 | ~n30873;
  assign n43174 = n30875 | ~n30876;
  assign n43175 = n30881 | ~n30882;
  assign n43176 = n30895 | n30896;
  assign n43177 = n30899 | n30900;
  assign n43178 = n30901 | n30902;
  assign n43179 = n30906 | n30907;
  assign n43180 = n30908 | n30909;
  assign n43181 = n30910 | ~n30911;
  assign n43182 = n30913 | ~n30914;
  assign n43183 = n30924 | n30925;
  assign n43184 = n30928 | n30929;
  assign n43185 = n30930 | n30931;
  assign n43186 = n30941 | n30938 | n30940;
  assign n43187 = n30942 | n30943;
  assign n43188 = n30945 | ~n30946;
  assign n43189 = n30947 | n30948;
  assign n43190 = n30949 | ~n30950;
  assign n43191 = n30963 | n30964;
  assign n43192 = n30967 | n30968;
  assign n43193 = n30969 | n30970;
  assign n43194 = n30974 | n30975;
  assign n43195 = n30976 | n30977;
  assign n43196 = n30978 | ~n30979;
  assign n43197 = n30981 | ~n30982;
  assign n43198 = n30992 | n30993;
  assign n43199 = n30996 | n30997;
  assign n43200 = n30998 | n30999;
  assign n43201 = n31002 | ~n31003;
  assign n43202 = n31011 | ~n31012;
  assign n43203 = n31030 | ~n31031;
  assign n43204 = n31036 | ~n31037;
  assign n43205 = n31047 | n31048;
  assign n43206 = n31051 | n31052;
  assign n43207 = n31053 | n31054;
  assign n43208 = n31067 | n31068;
  assign n43209 = n31071 | n31072;
  assign n43210 = n31073 | n31074;
  assign n43211 = n31086 | n31087;
  assign n43212 = n31090 | n31091;
  assign n43213 = n31092 | n31093;
  assign n43214 = n31102 | n31103;
  assign n43215 = n31106 | n31107;
  assign n43216 = n31108 | n31109;
  assign n43217 = n31125 | n31126;
  assign n43218 = n31129 | n31130;
  assign n43219 = n31131 | n31132;
  assign n43220 = n31138 | ~n31139;
  assign n43221 = n31149 | n31150;
  assign n43222 = n31153 | n31154;
  assign n43223 = n31155 | n31156;
  assign n43224 = n31162 | ~n31163;
  assign n43225 = n31168 | ~n31169;
  assign n43226 = n31174 | ~n31175;
  assign n43227 = n31180 | ~n31181;
  assign n43228 = n31184 | n31185;
  assign n43229 = n31196 | n31197;
  assign n43230 = n31200 | n31201;
  assign n43231 = n31202 | n31203;
  assign n43232 = n31209 | ~n31210;
  assign n43233 = n31220 | n31221;
  assign n43234 = n31224 | n31225;
  assign n43235 = n31226 | n31227;
  assign n43236 = n31233 | ~n31234;
  assign n43237 = n31244 | n31245;
  assign n43238 = n31248 | n31249;
  assign n43239 = n31250 | n31251;
  assign n43240 = n31257 | ~n31258;
  assign n43241 = n31268 | n31269;
  assign n43242 = n31272 | n31273;
  assign n43243 = n31274 | n31275;
  assign n43244 = n31281 | ~n31282;
  assign n43245 = n31287 | ~n31288;
  assign n43246 = n31301 | n31302;
  assign n43247 = n31305 | n31306;
  assign n43248 = n31307 | n31308;
  assign n43249 = n31314 | ~n31315;
  assign n43250 = n31320 | n31321;
  assign n43251 = n31325 | n31326;
  assign n43252 = n31327 | ~n31328;
  assign n43253 = n31344 | n31345;
  assign n43254 = n31348 | n31349;
  assign n43255 = n31350 | n31351;
  assign n43256 = n31354 | ~n31355;
  assign n43257 = n31366 | n31367;
  assign n43258 = n31370 | n31371;
  assign n43259 = n31372 | n31373;
  assign n43260 = n31381 | n31382;
  assign n43261 = n31385 | n31386;
  assign n43262 = n31387 | n31388;
  assign n43263 = n31396 | n31397;
  assign n43264 = n31400 | n31401;
  assign n43265 = n31402 | n31403;
  assign n43266 = n31412 | n31413;
  assign n43267 = n31416 | n31417;
  assign n43268 = n31418 | n31419;
  assign n43269 = n31427 | n31428;
  assign n43270 = n31431 | n31432;
  assign n43271 = n31433 | n31434;
  assign n43272 = n31442 | n31443;
  assign n43273 = n31446 | n31447;
  assign n43274 = n31448 | n31449;
  assign n43275 = n31459 | n31460;
  assign n43276 = n31465 | ~n31466;
  assign n43277 = n31471 | ~n31472;
  assign n43278 = n31477 | ~n31478;
  assign n43279 = n31488 | n31489;
  assign n43280 = n31492 | n31493;
  assign n43281 = n31494 | n31495;
  assign n43282 = n31501 | ~n31502;
  assign n43283 = n31504 | ~n31505;
  assign n43284 = n31510 | ~n31511;
  assign n43285 = n31516 | ~n31517;
  assign n43286 = n31525 | ~n31526;
  assign n43287 = n31536 | n31537;
  assign n43288 = n31540 | n31541;
  assign n43289 = n31542 | n31543;
  assign n43290 = n31549 | ~n31550;
  assign n43291 = n31552 | ~n31553;
  assign n43292 = n31563 | n31564;
  assign n43293 = n31567 | n31568;
  assign n43294 = n31569 | n31570;
  assign n43295 = n31576 | ~n31577;
  assign n43296 = n31582 | ~n31583;
  assign n43297 = n31586 | n31587;
  assign n43298 = n31590 | ~n31591;
  assign n43299 = n31607 | n31608;
  assign n43300 = n31611 | n31612;
  assign n43301 = n31613 | n31614;
  assign n43302 = n31620 | ~n31621;
  assign n43303 = n31630 | ~n31631;
  assign n43304 = n31633 | n31634;
  assign n43305 = n31635 | n31636;
  assign n43306 = n31642 | ~n31643;
  assign n43307 = n31651 | ~n31652;
  assign n43308 = n31655 | n31656;
  assign n43309 = n31668 | n31669;
  assign n43310 = n31672 | n31673;
  assign n43311 = n31674 | n31675;
  assign n43312 = n31685 | n31686;
  assign n43313 = n31689 | n31690;
  assign n43314 = n31691 | n31692;
  assign n43315 = n31701 | n31702;
  assign n43316 = n31705 | n31706;
  assign n43317 = n31707 | n31708;
  assign n43318 = n31716 | n31717;
  assign n43319 = n31720 | n31721;
  assign n43320 = n31722 | n31723;
  assign n43321 = n31733 | n31734;
  assign n43322 = n31737 | ~n31738;
  assign n43323 = n31743 | ~n31744;
  assign n43324 = n31749 | ~n31750;
  assign n43325 = n31763 | n31764;
  assign n43326 = n31767 | n31768;
  assign n43327 = n31769 | n31770;
  assign n43328 = n31774 | n31775;
  assign n43329 = n31776 | n31777;
  assign n43330 = n31778 | ~n31779;
  assign n43331 = n31781 | ~n31782;
  assign n43332 = n31792 | n31793;
  assign n43333 = n31796 | n31797;
  assign n43334 = n31798 | n31799;
  assign n43335 = n31803 | n31804;
  assign n43336 = n31805 | n31806;
  assign n43337 = n31807 | ~n31808;
  assign n43338 = n31810 | ~n31811;
  assign n43339 = n31816 | ~n31817;
  assign n43340 = n31830 | n31831;
  assign n43341 = n31834 | n31835;
  assign n43342 = n31836 | n31837;
  assign n43343 = n31841 | n31842;
  assign n43344 = n31843 | n31844;
  assign n43345 = n31845 | ~n31846;
  assign n43346 = n31848 | ~n31849;
  assign n43347 = n31859 | n31860;
  assign n43348 = n31863 | n31864;
  assign n43349 = n31865 | n31866;
  assign n43350 = n31876 | n31873 | n31875;
  assign n43351 = n31877 | n31878;
  assign n43352 = n31880 | ~n31881;
  assign n43353 = n31882 | n31883;
  assign n43354 = n31884 | ~n31885;
  assign n43355 = n31898 | n31899;
  assign n43356 = n31902 | n31903;
  assign n43357 = n31904 | n31905;
  assign n43358 = n31909 | n31910;
  assign n43359 = n31911 | n31912;
  assign n43360 = n31913 | ~n31914;
  assign n43361 = n31924 | n31925;
  assign n43362 = n31928 | n31929;
  assign n43363 = n31930 | n31931;
  assign n43364 = n31935 | n31936;
  assign n43365 = n31937 | n31938;
  assign n43366 = n31939 | ~n31940;
  assign n43367 = n31942 | ~n31943;
  assign n43368 = n31954 | n31955;
  assign n43369 = n31958 | n31959;
  assign n43370 = n31960 | n31961;
  assign n43371 = n31965 | n31966;
  assign n43372 = n31967 | n31968;
  assign n43373 = n31969 | ~n31970;
  assign n43374 = n31989 | ~n31990;
  assign n43375 = n32005 | n32006;
  assign n43376 = n32009 | n32010;
  assign n43377 = n32011 | n32012;
  assign n43378 = n32024 | n32025;
  assign n43379 = n32028 | n32029;
  assign n43380 = n32030 | n32031;
  assign n43381 = n32040 | n32041;
  assign n43382 = n32044 | n32045;
  assign n43383 = n32046 | n32047;
  assign n43384 = n32050 | n32051;
  assign n43385 = n32064 | n32065;
  assign n43386 = n32068 | n32069;
  assign n43387 = n32070 | n32071;
  assign n43388 = n32080 | ~n32081;
  assign n43389 = n32084 | n32085;
  assign n43390 = n32091 | ~n32092;
  assign n43391 = n32095 | n32096;
  assign n43392 = n32107 | n32108;
  assign n43393 = n32111 | n32112;
  assign n43394 = n32113 | n32114;
  assign n43395 = n32120 | ~n32121;
  assign n43396 = n32131 | n32132;
  assign n43397 = n32135 | n32136;
  assign n43398 = n32137 | n32138;
  assign n43399 = n32144 | ~n32145;
  assign n43400 = n32155 | n32156;
  assign n43401 = n32159 | n32160;
  assign n43402 = n32161 | n32162;
  assign n43403 = n32168 | ~n32169;
  assign n43404 = n32179 | n32180;
  assign n43405 = n32183 | n32184;
  assign n43406 = n32185 | n32186;
  assign n43407 = n32192 | ~n32193;
  assign n43408 = n32198 | ~n32199;
  assign n43409 = n32212 | n32213;
  assign n43410 = n32216 | n32217;
  assign n43411 = n32218 | n32219;
  assign n43412 = n32225 | ~n32226;
  assign n43413 = n32236 | n32237;
  assign n43414 = n32240 | n32241;
  assign n43415 = n32242 | n32243;
  assign n43416 = n32249 | n32250;
  assign n43417 = n32254 | n32255;
  assign n43418 = n32256 | ~n32257;
  assign n43419 = n32262 | ~n32263;
  assign n43420 = n32274 | ~n32275;
  assign n43421 = n32277 | n32278;
  assign n43422 = n32279 | n32280;
  assign n43423 = n32286 | ~n32287;
  assign n43424 = n32295 | n32296;
  assign n43425 = n32299 | n32300;
  assign n43426 = n32301 | n32302;
  assign n43427 = n32310 | n32311;
  assign n43428 = n32314 | n32315;
  assign n43429 = n32316 | n32317;
  assign n43430 = n32325 | n32326;
  assign n43431 = n32329 | n32330;
  assign n43432 = n32331 | n32332;
  assign n43433 = n32341 | n32342;
  assign n43434 = n32345 | n32346;
  assign n43435 = n32347 | n32348;
  assign n43436 = n32357 | n32358;
  assign n43437 = n32361 | n32362;
  assign n43438 = n32363 | n32364;
  assign n43439 = n32372 | n32373;
  assign n43440 = n32376 | n32377;
  assign n43441 = n32378 | n32379;
  assign n43442 = n32389 | n32390;
  assign n43443 = n32395 | ~n32396;
  assign n43444 = n32399 | n32400;
  assign n43445 = n32401 | n32402;
  assign n43446 = n32403 | ~n32404;
  assign n43447 = n32409 | ~n32410;
  assign n43448 = n32424 | ~n32425;
  assign n43449 = n32435 | n32436;
  assign n43450 = n32439 | n32440;
  assign n43451 = n32441 | n32442;
  assign n43452 = n32448 | ~n32449;
  assign n43453 = n32451 | ~n32452;
  assign n43454 = n32462 | n32463;
  assign n43455 = n32466 | n32467;
  assign n43456 = n32468 | n32469;
  assign n43457 = n32475 | ~n32476;
  assign n43458 = n32481 | ~n32482;
  assign n43459 = n32485 | n32486;
  assign n43460 = n32489 | ~n32490;
  assign n43461 = n32506 | n32507;
  assign n43462 = n32510 | n32511;
  assign n43463 = n32512 | n32513;
  assign n43464 = n32519 | ~n32520;
  assign n43465 = n32522 | ~n32523;
  assign n43466 = n32533 | n32534;
  assign n43467 = n32537 | n32538;
  assign n43468 = n32539 | n32540;
  assign n43469 = n32546 | ~n32547;
  assign n43470 = n32552 | ~n32553;
  assign n43471 = n32558 | ~n32559;
  assign n43472 = n32562 | n32563;
  assign n43473 = n32574 | n32575;
  assign n43474 = n32578 | n32579;
  assign n43475 = n32580 | n32581;
  assign n43476 = n32593 | n32594;
  assign n43477 = n32597 | n32598;
  assign n43478 = n32599 | n32600;
  assign n43479 = n32608 | n32609;
  assign n43480 = n32612 | n32613;
  assign n43481 = n32614 | n32615;
  assign n43482 = n32625 | n32626;
  assign n43483 = n32629 | ~n32630;
  assign n43484 = n32635 | ~n32636;
  assign n43485 = n32641 | ~n32642;
  assign n43486 = n32655 | n32656;
  assign n43487 = n32659 | n32660;
  assign n43488 = n32661 | n32662;
  assign n43489 = n32666 | n32667;
  assign n43490 = n32668 | n32669;
  assign n43491 = n32670 | ~n32671;
  assign n43492 = n32681 | n32682;
  assign n43493 = n32685 | n32686;
  assign n43494 = n32687 | n32688;
  assign n43495 = n32692 | n32693;
  assign n43496 = n32694 | n32695;
  assign n43497 = n32696 | ~n32697;
  assign n43498 = n32707 | n32708;
  assign n43499 = n32711 | n32712;
  assign n43500 = n32713 | n32714;
  assign n43501 = n32718 | n32719;
  assign n43502 = n32720 | n32721;
  assign n43503 = n32722 | ~n32723;
  assign n43504 = n32725 | ~n32726;
  assign n43505 = n32736 | n32737;
  assign n43506 = n32740 | n32741;
  assign n43507 = n32742 | n32743;
  assign n43508 = n32753 | n32750 | n32752;
  assign n43509 = n32754 | n32755;
  assign n43510 = n32757 | ~n32758;
  assign n43511 = n32759 | n32760;
  assign n43512 = n32761 | ~n32762;
  assign n43513 = n32775 | n32776;
  assign n43514 = n32779 | n32780;
  assign n43515 = n32781 | n32782;
  assign n43516 = n32786 | n32787;
  assign n43517 = n32788 | n32789;
  assign n43518 = n32790 | ~n32791;
  assign n43519 = n32801 | n32802;
  assign n43520 = n32805 | n32806;
  assign n43521 = n32807 | n32808;
  assign n43522 = n32812 | n32813;
  assign n43523 = n32814 | n32815;
  assign n43524 = n32816 | ~n32817;
  assign n43525 = n32819 | ~n32820;
  assign n43526 = n32830 | n32831;
  assign n43527 = n32834 | n32835;
  assign n43528 = n32836 | n32837;
  assign n43529 = n32840 | ~n32841;
  assign n43530 = n32844 | n32845;
  assign n43531 = n32846 | n32847;
  assign n43532 = n32848 | ~n32849;
  assign n43533 = n32854 | ~n32855;
  assign n43534 = n32871 | ~n32872;
  assign n43535 = n32887 | n32888;
  assign n43536 = n32891 | n32892;
  assign n43537 = n32893 | n32894;
  assign n43538 = n32906 | n32907;
  assign n43539 = n32910 | n32911;
  assign n43540 = n32912 | n32913;
  assign n43541 = n32916 | n32917;
  assign n43542 = n32930 | n32931;
  assign n43543 = n32934 | n32935;
  assign n43544 = n32936 | n32937;
  assign n43545 = n32946 | ~n32947;
  assign n43546 = n32950 | n32951;
  assign n43547 = n32962 | n32963;
  assign n43548 = n32966 | n32967;
  assign n43549 = n32968 | n32969;
  assign n43550 = n32975 | ~n32976;
  assign n43551 = n32986 | n32987;
  assign n43552 = n32990 | n32991;
  assign n43553 = n32992 | n32993;
  assign n43554 = n32999 | ~n33000;
  assign n43555 = n33010 | n33011;
  assign n43556 = n33014 | n33015;
  assign n43557 = n33016 | n33017;
  assign n43558 = n33023 | ~n33024;
  assign n43559 = n33034 | n33035;
  assign n43560 = n33038 | n33039;
  assign n43561 = n33040 | n33041;
  assign n43562 = n33047 | ~n33048;
  assign n43563 = n33053 | ~n33054;
  assign n43564 = n33067 | n33068;
  assign n43565 = n33071 | n33072;
  assign n43566 = n33073 | n33074;
  assign n43567 = n33080 | ~n33081;
  assign n43568 = n33091 | n33092;
  assign n43569 = n33095 | n33096;
  assign n43570 = n33097 | n33098;
  assign n43571 = n33104 | n33105;
  assign n43572 = n33109 | n33110;
  assign n43573 = n33111 | ~n33112;
  assign n43574 = n33117 | ~n33118;
  assign n43575 = n33129 | ~n33130;
  assign n43576 = n33132 | n33133;
  assign n43577 = n33134 | n33135;
  assign n43578 = n33141 | ~n33142;
  assign n43579 = n33150 | n33151;
  assign n43580 = n33154 | n33155;
  assign n43581 = n33156 | n33157;
  assign n43582 = n33165 | n33166;
  assign n43583 = n33169 | n33170;
  assign n43584 = n33171 | n33172;
  assign n43585 = n33180 | n33181;
  assign n43586 = n33184 | n33185;
  assign n43587 = n33186 | n33187;
  assign n43588 = n33196 | n33197;
  assign n43589 = n33200 | n33201;
  assign n43590 = n33202 | n33203;
  assign n43591 = n33211 | n33212;
  assign n43592 = n33215 | n33216;
  assign n43593 = n33217 | n33218;
  assign n43594 = n33228 | n33229;
  assign n43595 = n33234 | ~n33235;
  assign n43596 = n33238 | n33239;
  assign n43597 = n33240 | n33241;
  assign n43598 = n33242 | ~n33243;
  assign n43599 = n33248 | ~n33249;
  assign n43600 = n33257 | ~n33258;
  assign n43601 = n33268 | n33269;
  assign n43602 = n33272 | n33273;
  assign n43603 = n33274 | n33275;
  assign n43604 = n33281 | ~n33282;
  assign n43605 = n33284 | ~n33285;
  assign n43606 = n33295 | n33296;
  assign n43607 = n33299 | n33300;
  assign n43608 = n33301 | n33302;
  assign n43609 = n33308 | ~n33309;
  assign n43610 = n33314 | ~n33315;
  assign n43611 = n33318 | n33319;
  assign n43612 = n33322 | ~n33323;
  assign n43613 = n33339 | n33340;
  assign n43614 = n33343 | n33344;
  assign n43615 = n33345 | n33346;
  assign n43616 = n33352 | ~n33353;
  assign n43617 = n33355 | ~n33356;
  assign n43618 = n33366 | n33367;
  assign n43619 = n33370 | n33371;
  assign n43620 = n33372 | n33373;
  assign n43621 = n33379 | ~n33380;
  assign n43622 = n33385 | ~n33386;
  assign n43623 = n33402 | n33403;
  assign n43624 = n33406 | n33407;
  assign n43625 = n33408 | n33409;
  assign n43626 = n33419 | n33420;
  assign n43627 = n33423 | n33424;
  assign n43628 = n33425 | n33426;
  assign n43629 = n33433 | ~n33434;
  assign n43630 = n33450 | n33451;
  assign n43631 = n33454 | n33455;
  assign n43632 = n33456 | n33457;
  assign n43633 = n33468 | n33469;
  assign n43634 = n33472 | n33473;
  assign n43635 = n33474 | n33475;
  assign n43636 = n33479 | n33480;
  assign n43637 = n33481 | n33482;
  assign n43638 = n33483 | ~n33484;
  assign n43639 = n33489 | ~n33490;
  assign n43640 = n33493 | n33494;
  assign n43641 = n33495 | n33496;
  assign n43642 = n33497 | ~n33498;
  assign n43643 = n33508 | n33509;
  assign n43644 = n33512 | n33513;
  assign n43645 = n33514 | n33515;
  assign n43646 = n33519 | n33520;
  assign n43647 = n33521 | n33522;
  assign n43648 = n33523 | ~n33524;
  assign n43649 = n33526 | ~n33527;
  assign n43650 = n33537 | n33538;
  assign n43651 = n33541 | n33542;
  assign n43652 = n33543 | n33544;
  assign n43653 = n33564 | n33565;
  assign n43654 = n33568 | n33569;
  assign n43655 = n33570 | n33571;
  assign n43656 = n33575 | n33576;
  assign n43657 = n33577 | n33578;
  assign n43658 = n33579 | ~n33580;
  assign n43659 = n33590 | n33591;
  assign n43660 = n33594 | n33595;
  assign n43661 = n33596 | n33597;
  assign n43662 = n33601 | n33602;
  assign n43663 = n33603 | n33604;
  assign n43664 = n33605 | ~n33606;
  assign n43665 = n33608 | ~n33609;
  assign n43666 = n33619 | n33620;
  assign n43667 = n33623 | n33624;
  assign n43668 = n33625 | n33626;
  assign n43669 = n33630 | n33631;
  assign n43670 = n33632 | n33633;
  assign n43671 = n33634 | ~n33635;
  assign n43672 = n33637 | ~n33638;
  assign n43673 = n33643 | ~n33644;
  assign n43674 = n33659 | ~n33660;
  assign n43675 = n33675 | n33676;
  assign n43676 = n33679 | n33680;
  assign n43677 = n33681 | n33682;
  assign n43678 = n33695 | n33696;
  assign n43679 = n33699 | n33700;
  assign n43680 = n33701 | n33702;
  assign n43681 = n33710 | n33711;
  assign n43682 = n33712 | n33713;
  assign n43683 = n33714 | ~n33715;
  assign n43684 = n33718 | n33719;
  assign n43685 = n33720 | n33721;
  assign n43686 = n33722 | ~n33723;
  assign n43687 = n33733 | n33734;
  assign n43688 = n33737 | n33738;
  assign n43689 = n33739 | n33740;
  assign n43690 = n33746 | ~n33747;
  assign n43691 = n33757 | n33758;
  assign n43692 = n33761 | n33762;
  assign n43693 = n33763 | n33764;
  assign n43694 = n33770 | ~n33771;
  assign n43695 = n33781 | n33782;
  assign n43696 = n33785 | n33786;
  assign n43697 = n33787 | n33788;
  assign n43698 = n33794 | ~n33795;
  assign n43699 = n33805 | n33806;
  assign n43700 = n33809 | n33810;
  assign n43701 = n33811 | n33812;
  assign n43702 = n33818 | ~n33819;
  assign n43703 = n33824 | ~n33825;
  assign n43704 = n33830 | ~n33831;
  assign n43705 = n33841 | n33842;
  assign n43706 = n33845 | n33846;
  assign n43707 = n33847 | n33848;
  assign n43708 = n33854 | ~n33855;
  assign n43709 = n33865 | n33866;
  assign n43710 = n33869 | n33870;
  assign n43711 = n33871 | n33872;
  assign n43712 = n33878 | n33879;
  assign n43713 = n33883 | n33884;
  assign n43714 = n33885 | ~n33886;
  assign n43715 = n33901 | ~n33902;
  assign n43716 = n33904 | n33905;
  assign n43717 = n33906 | n33907;
  assign n43718 = n33913 | ~n33914;
  assign n43719 = n33922 | n33923;
  assign n43720 = n33926 | n33927;
  assign n43721 = n33928 | n33929;
  assign n43722 = n33937 | n33938;
  assign n43723 = n33941 | n33942;
  assign n43724 = n33943 | n33944;
  assign n43725 = n33952 | n33953;
  assign n43726 = n33956 | n33957;
  assign n43727 = n33958 | n33959;
  assign n43728 = n33967 | n33968;
  assign n43729 = n33971 | n33972;
  assign n43730 = n33973 | n33974;
  assign n43731 = n33982 | n33983;
  assign n43732 = n33984 | n33985;
  assign n43733 = n33986 | ~n33987;
  assign n43734 = n33990 | n33991;
  assign n43735 = n33992 | n33993;
  assign n43736 = n33994 | ~n33995;
  assign n43737 = n34000 | ~n34001;
  assign n43738 = n34006 | ~n34007;
  assign n43739 = n34009 | ~n34010;
  assign n43740 = n34020 | n34021;
  assign n43741 = n34024 | n34025;
  assign n43742 = n34026 | n34027;
  assign n43743 = n34033 | ~n34034;
  assign n43744 = n34036 | ~n34037;
  assign n43745 = n34047 | n34048;
  assign n43746 = n34051 | n34052;
  assign n43747 = n34053 | n34054;
  assign n43748 = n34060 | ~n34061;
  assign n43749 = n34066 | ~n34067;
  assign n43750 = n34070 | n34071;
  assign n43751 = n34074 | ~n34075;
  assign n43752 = n34091 | n34092;
  assign n43753 = n34095 | n34096;
  assign n43754 = n34097 | n34098;
  assign n43755 = n34104 | ~n34105;
  assign n43756 = n34107 | ~n34108;
  assign n43757 = n34118 | n34119;
  assign n43758 = n34122 | n34123;
  assign n43759 = n34124 | n34125;
  assign n43760 = n34131 | ~n34132;
  assign n43761 = n34137 | ~n34138;
  assign n43762 = n34154 | n34155;
  assign n43763 = n34158 | n34159;
  assign n43764 = n34160 | n34161;
  assign n43765 = n34170 | n34171;
  assign n43766 = n34174 | n34175;
  assign n43767 = n34176 | n34177;
  assign n43768 = n34185 | n34186;
  assign n43769 = n34189 | n34190;
  assign n43770 = n34191 | n34192;
  assign n43771 = n34199 | ~n34200;
  assign n43772 = n34216 | n34217;
  assign n43773 = n34220 | n34221;
  assign n43774 = n34222 | n34223;
  assign n43775 = n34229 | ~n34230;
  assign n43776 = n34235 | ~n34236;
  assign n43777 = n34238 | ~n34239;
  assign n43778 = n34244 | ~n34245;
  assign n43779 = n34248 | n34249;
  assign n43780 = n34250 | n34251;
  assign n43781 = n34252 | ~n34253;
  assign n43782 = n34255 | ~n34256;
  assign n43783 = n34266 | n34267;
  assign n43784 = n34270 | n34271;
  assign n43785 = n34272 | n34273;
  assign n43786 = n34293 | n34294;
  assign n43787 = n34297 | n34298;
  assign n43788 = n34299 | n34300;
  assign n43789 = n34304 | n34305;
  assign n43790 = n34306 | n34307;
  assign n43791 = n34308 | ~n34309;
  assign n43792 = n34319 | n34320;
  assign n43793 = n34323 | n34324;
  assign n43794 = n34325 | n34326;
  assign n43795 = n34330 | n34331;
  assign n43796 = n34332 | n34333;
  assign n43797 = n34334 | ~n34335;
  assign n43798 = n34337 | ~n34338;
  assign n43799 = n34348 | n34349;
  assign n43800 = n34352 | n34353;
  assign n43801 = n34354 | n34355;
  assign n43802 = n34359 | n34360;
  assign n43803 = n34361 | n34362;
  assign n43804 = n34363 | ~n34364;
  assign n43805 = n34366 | ~n34367;
  assign n43806 = n34372 | ~n34373;
  assign n43807 = n34388 | ~n34389;
  assign n43808 = n34404 | n34405;
  assign n43809 = n34408 | n34409;
  assign n43810 = n34410 | n34411;
  assign n43811 = n34429 | n34430;
  assign n43812 = n34433 | ~n34434;
  assign n43813 = n34442 | ~n34443;
  assign n43814 = n34453 | n34454;
  assign n43815 = n34457 | n34458;
  assign n43816 = n34459 | n34460;
  assign n43817 = n34466 | ~n34467;
  assign n43818 = n34477 | n34478;
  assign n43819 = n34481 | n34482;
  assign n43820 = n34483 | n34484;
  assign n43821 = n34490 | ~n34491;
  assign n43822 = n34501 | n34502;
  assign n43823 = n34505 | n34506;
  assign n43824 = n34507 | n34508;
  assign n43825 = n34514 | ~n34515;
  assign n43826 = n34520 | ~n34521;
  assign n43827 = n34526 | ~n34527;
  assign n43828 = n34537 | n34538;
  assign n43829 = n34541 | n34542;
  assign n43830 = n34543 | n34544;
  assign n43831 = n34550 | ~n34551;
  assign n43832 = n34561 | n34562;
  assign n43833 = n34565 | n34566;
  assign n43834 = n34567 | n34568;
  assign n43835 = n34574 | n34575;
  assign n43836 = n34579 | n34580;
  assign n43837 = n34581 | ~n34582;
  assign n43838 = n34597 | ~n34598;
  assign n43839 = n34600 | n34601;
  assign n43840 = n34602 | n34603;
  assign n43841 = n34609 | ~n34610;
  assign n43842 = n34618 | n34619;
  assign n43843 = n34622 | n34623;
  assign n43844 = n34624 | n34625;
  assign n43845 = n34633 | n34634;
  assign n43846 = n34637 | n34638;
  assign n43847 = n34639 | n34640;
  assign n43848 = n34648 | n34649;
  assign n43849 = n34652 | n34653;
  assign n43850 = n34654 | n34655;
  assign n43851 = n34663 | n34664;
  assign n43852 = n34667 | n34668;
  assign n43853 = n34669 | n34670;
  assign n43854 = n34678 | n34679;
  assign n43855 = n34680 | n34681;
  assign n43856 = n34682 | ~n34683;
  assign n43857 = n34686 | n34687;
  assign n43858 = n34688 | n34689;
  assign n43859 = n34690 | ~n34691;
  assign n43860 = n34696 | ~n34697;
  assign n43861 = n34702 | ~n34703;
  assign n43862 = n34713 | n34714;
  assign n43863 = n34717 | n34718;
  assign n43864 = n34719 | n34720;
  assign n43865 = n34726 | ~n34727;
  assign n43866 = n34732 | ~n34733;
  assign n43867 = n34736 | n34737;
  assign n43868 = n34740 | ~n34741;
  assign n43869 = n34746 | ~n34747;
  assign n43870 = n34750 | n34751;
  assign n43871 = n34762 | n34763;
  assign n43872 = n34766 | n34767;
  assign n43873 = n34768 | n34769;
  assign n43874 = n34775 | ~n34776;
  assign n43875 = n34778 | ~n34779;
  assign n43876 = n34789 | n34790;
  assign n43877 = n34793 | n34794;
  assign n43878 = n34795 | n34796;
  assign n43879 = n34802 | ~n34803;
  assign n43880 = n34808 | ~n34809;
  assign n43881 = n34824 | n34825;
  assign n43882 = n34828 | n34829;
  assign n43883 = n34830 | n34831;
  assign n43884 = n34840 | n34841;
  assign n43885 = n34844 | n34845;
  assign n43886 = n34846 | n34847;
  assign n43887 = n34856 | n34857;
  assign n43888 = n34860 | n34861;
  assign n43889 = n34862 | n34863;
  assign n43890 = n34871 | ~n34872;
  assign n43891 = n34885 | n34886;
  assign n43892 = n34889 | n34890;
  assign n43893 = n34891 | n34892;
  assign n43894 = n34896 | n34897;
  assign n43895 = n34898 | n34899;
  assign n43896 = n34900 | ~n34901;
  assign n43897 = n34911 | n34912;
  assign n43898 = n34915 | n34916;
  assign n43899 = n34917 | n34918;
  assign n43900 = n34922 | n34923;
  assign n43901 = n34924 | n34925;
  assign n43902 = n34926 | ~n34927;
  assign n43903 = n34933 | n34934;
  assign n43904 = n34935 | n34936;
  assign n43905 = n34937 | ~n34938;
  assign n43906 = n34941 | n34942;
  assign n43907 = n34943 | n34944;
  assign n43908 = n34945 | ~n34946;
  assign n43909 = n34965 | n34966;
  assign n43910 = n34969 | n34970;
  assign n43911 = n34971 | n34972;
  assign n43912 = n34976 | n34977;
  assign n43913 = n34978 | n34979;
  assign n43914 = n34980 | ~n34981;
  assign n43915 = n34983 | ~n34984;
  assign n43916 = n34994 | n34995;
  assign n43917 = n34998 | n34999;
  assign n43918 = n35000 | n35001;
  assign n43919 = n35005 | n35006;
  assign n43920 = n35007 | n35008;
  assign n43921 = n35009 | ~n35010;
  assign n43922 = n35012 | ~n35013;
  assign n43923 = n35018 | ~n35019;
  assign n43924 = n35034 | ~n35035;
  assign n43925 = n35048 | n35049;
  assign n43926 = n35052 | n35053;
  assign n43927 = n35054 | n35055;
  assign n43928 = n35064 | n35065;
  assign n43929 = n35068 | n35069;
  assign n43930 = n35070 | n35071;
  assign n43931 = n35083 | n35084;
  assign n43932 = n35087 | ~n35088;
  assign n43933 = n35098 | n35099;
  assign n43934 = n35100 | n35101;
  assign n43935 = n35102 | ~n35103;
  assign n43936 = n35116 | n35117;
  assign n43937 = n35120 | n35121;
  assign n43938 = n35122 | n35123;
  assign n43939 = n35129 | ~n35130;
  assign n43940 = n35140 | n35141;
  assign n43941 = n35144 | n35145;
  assign n43942 = n35146 | n35147;
  assign n43943 = n35153 | ~n35154;
  assign n43944 = n35164 | n35165;
  assign n43945 = n35168 | n35169;
  assign n43946 = n35170 | n35171;
  assign n43947 = n35177 | ~n35178;
  assign n43948 = n35183 | ~n35184;
  assign n43949 = n35192 | ~n35193;
  assign n43950 = n35198 | ~n35199;
  assign n43951 = n35204 | ~n35205;
  assign n43952 = n35218 | ~n35219;
  assign n43953 = n35221 | n35222;
  assign n43954 = n35223 | n35224;
  assign n43955 = n35227 | ~n35228;
  assign n43956 = n35233 | ~n35234;
  assign n43957 = n35241 | n35242;
  assign n43958 = n35245 | n35246;
  assign n43959 = n35247 | n35248;
  assign n43960 = n35257 | n35258;
  assign n43961 = n35261 | n35262;
  assign n43962 = n35263 | n35264;
  assign n43963 = n35272 | n35273;
  assign n43964 = n35276 | n35277;
  assign n43965 = n35278 | n35279;
  assign n43966 = n35287 | n35288;
  assign n43967 = n35291 | n35292;
  assign n43968 = n35293 | n35294;
  assign n43969 = n35309 | n35310;
  assign n43970 = n35313 | ~n35314;
  assign n43971 = n35325 | ~n35326;
  assign n43972 = n35329 | n35330;
  assign n43973 = n35333 | ~n35334;
  assign n43974 = n35339 | ~n35340;
  assign n43975 = n35343 | n35344;
  assign n43976 = n35347 | ~n35348;
  assign n43977 = n35353 | ~n35354;
  assign n43978 = n35357 | n35358;
  assign n43979 = n35361 | ~n35362;
  assign n43980 = n35372 | n35373;
  assign n43981 = n35376 | n35377;
  assign n43982 = n35378 | n35379;
  assign n43983 = n35385 | ~n35386;
  assign n43984 = n35391 | ~n35392;
  assign n43985 = n35394 | n35395;
  assign n43986 = n35396 | n35397;
  assign n43987 = n35399 | ~n35400;
  assign n43988 = n35405 | ~n35406;
  assign n43989 = n35408 | ~n35409;
  assign n43990 = n35423 | n35424;
  assign n43991 = n35427 | n35428;
  assign n43992 = n35429 | n35430;
  assign n43993 = n35439 | n35440;
  assign n43994 = n35443 | n35444;
  assign n43995 = n35445 | n35446;
  assign n43996 = n35455 | n35456;
  assign n43997 = n35459 | n35460;
  assign n43998 = n35461 | n35462;
  assign n43999 = n35471 | n35472;
  assign n44000 = n35475 | n35476;
  assign n44001 = n35477 | n35478;
  assign n44002 = n35486 | n35487;
  assign n44003 = n35490 | n35491;
  assign n44004 = n35492 | n35493;
  assign n44005 = n35504 | n35505;
  assign n44006 = n35508 | ~n35509;
  assign n44007 = n35514 | ~n35515;
  assign n44008 = n35520 | ~n35521;
  assign n44009 = n35544 | ~n35545;
  assign n44010 = n35555 | n35556;
  assign n44011 = n35559 | n35560;
  assign n44012 = n35561 | n35562;
  assign n44013 = n35566 | n35567;
  assign n44014 = n35568 | n35569;
  assign n44015 = n35570 | ~n35571;
  assign n44016 = n35573 | ~n35574;
  assign n44017 = n35579 | ~n35580;
  assign n44018 = n35595 | ~n35596;
  assign n44019 = n35609 | n35610;
  assign n44020 = n35613 | n35614;
  assign n44021 = n35615 | n35616;
  assign n44022 = n35625 | n35626;
  assign n44023 = n35629 | n35630;
  assign n44024 = n35631 | n35632;
  assign n44025 = n35642 | n35643;
  assign n44026 = n35646 | n35647;
  assign n44027 = n35648 | n35649;
  assign n44028 = n35652 | n35653;
  assign n44029 = n35666 | n35667;
  assign n44030 = n35670 | n35671;
  assign n44031 = n35672 | n35673;
  assign n44032 = n35682 | ~n35683;
  assign n44033 = n35686 | n35687;
  assign n44034 = n35698 | n35699;
  assign n44035 = n35702 | n35703;
  assign n44036 = n35704 | n35705;
  assign n44037 = n35711 | ~n35712;
  assign n44038 = n35717 | ~n35718;
  assign n44039 = n35726 | ~n35727;
  assign n44040 = n35732 | ~n35733;
  assign n44041 = n35738 | ~n35739;
  assign n44042 = n35752 | n35753;
  assign n44043 = n35758 | ~n35759;
  assign n44044 = n35769 | n35770;
  assign n44045 = n35773 | n35774;
  assign n44046 = n35775 | n35776;
  assign n44047 = n35785 | n35786;
  assign n44048 = n35789 | n35790;
  assign n44049 = n35791 | n35792;
  assign n44050 = n35801 | n35802;
  assign n44051 = n35805 | n35806;
  assign n44052 = n35807 | n35808;
  assign n44053 = n35816 | n35817;
  assign n44054 = n35820 | n35821;
  assign n44055 = n35822 | n35823;
  assign n44056 = n35833 | n35834;
  assign n44057 = n35839 | ~n35840;
  assign n44058 = n35845 | ~n35846;
  assign n44059 = n35854 | ~n35855;
  assign n44060 = n35858 | n35859;
  assign n44061 = n35862 | ~n35863;
  assign n44062 = n35873 | n35874;
  assign n44063 = n35877 | n35878;
  assign n44064 = n35879 | n35880;
  assign n44065 = n35886 | ~n35887;
  assign n44066 = n35892 | ~n35893;
  assign n44067 = n35895 | n35896;
  assign n44068 = n35897 | n35898;
  assign n44069 = n35900 | ~n35901;
  assign n44070 = n35906 | ~n35907;
  assign n44071 = n35909 | ~n35910;
  assign n44072 = n35924 | n35925;
  assign n44073 = n35928 | n35929;
  assign n44074 = n35930 | n35931;
  assign n44075 = n35940 | n35941;
  assign n44076 = n35944 | n35945;
  assign n44077 = n35946 | n35947;
  assign n44078 = n35956 | n35957;
  assign n44079 = n35960 | n35961;
  assign n44080 = n35962 | n35963;
  assign n44081 = n35971 | n35972;
  assign n44082 = n35975 | n35976;
  assign n44083 = n35977 | n35978;
  assign n44084 = n35984 | ~n35985;
  assign n44085 = n35994 | n35995;
  assign n44086 = n35996 | n35997;
  assign n44087 = n35998 | ~n35999;
  assign n44088 = n36002 | n36003;
  assign n44089 = n36004 | n36005;
  assign n44090 = n36006 | ~n36007;
  assign n44091 = n36024 | ~n36025;
  assign n44092 = n36035 | n36036;
  assign n44093 = n36039 | n36040;
  assign n44094 = n36041 | n36042;
  assign n44095 = n36046 | n36047;
  assign n44096 = n36048 | n36049;
  assign n44097 = n36050 | ~n36051;
  assign n44098 = n36053 | ~n36054;
  assign n44099 = n36059 | ~n36060;
  assign n44100 = n36076 | n36077;
  assign n44101 = n36080 | n36081;
  assign n44102 = n36082 | n36083;
  assign n44103 = n36092 | n36093;
  assign n44104 = n36096 | n36097;
  assign n44105 = n36098 | n36099;
  assign n44106 = n36108 | n36109;
  assign n44107 = n36112 | n36113;
  assign n44108 = n36114 | n36115;
  assign n44109 = n36131 | n36132;
  assign n44110 = n36135 | ~n36136;
  assign n44111 = n36147 | ~n36148;
  assign n44112 = n36151 | n36152;
  assign n44113 = n36164 | ~n36165;
  assign n44114 = n36168 | n36169;
  assign n44115 = n36180 | n36181;
  assign n44116 = n36182 | n36183;
  assign n44117 = n36189 | ~n36190;
  assign n44118 = n36204 | n36205;
  assign n44119 = n36221 | n36222;
  assign n44120 = n36225 | n36226;
  assign n44121 = n36227 | n36228;
  assign n44122 = n36235 | n36236;
  assign n44123 = n36237 | n36238;
  assign n44124 = n36239 | ~n36240;
  assign n44125 = n36243 | n36244;
  assign n44126 = n36245 | n36246;
  assign n44127 = n36247 | ~n36248;
  assign n44128 = n36258 | n36259;
  assign n44129 = n36262 | n36263;
  assign n44130 = n36264 | n36265;
  assign n44131 = n36279 | n36280;
  assign n44132 = n36283 | n36284;
  assign n44133 = n36285 | n36286;
  assign n44134 = n36292 | ~n36293;
  assign n44135 = n36303 | n36304;
  assign n44136 = n36307 | n36308;
  assign n44137 = n36309 | n36310;
  assign n44138 = n36316 | ~n36317;
  assign n44139 = n36322 | ~n36323;
  assign n44140 = n36325 | ~n36326;
  assign n44141 = n36340 | n36341;
  assign n44142 = n36344 | n36345;
  assign n44143 = n36346 | n36347;
  assign n44144 = n36356 | n36357;
  assign n44145 = n36360 | n36361;
  assign n44146 = n36362 | n36363;
  assign n44147 = n36371 | n36372;
  assign n44148 = n36375 | n36376;
  assign n44149 = n36377 | n36378;
  assign n44150 = n36392 | n36393;
  assign n44151 = n36394 | n36395;
  assign n44152 = n36396 | ~n36397;
  assign n44153 = n36403 | n36400 | n36402;
  assign n44154 = n36407 | n36408;
  assign n44155 = n36409 | n36410;
  assign n44156 = n36411 | ~n36412;
  assign n44157 = n36418 | n36415 | n36417;
  assign n44158 = n36424 | ~n36425;
  assign n44159 = n36435 | n36436;
  assign n44160 = n36439 | n36440;
  assign n44161 = n36441 | n36442;
  assign n44162 = n36446 | n36447;
  assign n44163 = n36448 | n36449;
  assign n44164 = n36450 | ~n36451;
  assign n44165 = n36453 | ~n36454;
  assign n44166 = n36459 | ~n36460;
  assign n44167 = n36476 | n36477;
  assign n44168 = n36480 | n36481;
  assign n44169 = n36482 | n36483;
  assign n44170 = n36492 | n36493;
  assign n44171 = n36496 | n36497;
  assign n44172 = n36498 | n36499;
  assign n44173 = n36515 | n36516;
  assign n44174 = n36519 | n36520;
  assign n44175 = n36521 | n36522;
  assign n44176 = n36537 | ~n36538;
  assign n44177 = n36541 | n36542;
  assign n44178 = n36553 | n36554;
  assign n44179 = n36555 | n36556;
  assign n44180 = n36562 | ~n36563;
  assign n44181 = n36577 | n36578;
  assign n44182 = n36592 | n36593;
  assign n44183 = n36596 | n36597;
  assign n44184 = n36598 | n36599;
  assign n44185 = n36607 | n36608;
  assign n44186 = n36611 | n36612;
  assign n44187 = n36613 | n36614;
  assign n44188 = n36624 | n36625;
  assign n44189 = n36630 | ~n36631;
  assign n44190 = n36636 | ~n36637;
  assign n44191 = n36650 | n36651;
  assign n44192 = n36654 | n36655;
  assign n44193 = n36656 | n36657;
  assign n44194 = n36663 | ~n36664;
  assign n44195 = n36669 | ~n36670;
  assign n44196 = n36672 | ~n36673;
  assign n44197 = n36688 | n36689;
  assign n44198 = n36692 | n36693;
  assign n44199 = n36694 | n36695;
  assign n44200 = n36698 | ~n36699;
  assign n44201 = n36702 | n36703;
  assign n44202 = n36704 | n36705;
  assign n44203 = n36706 | ~n36707;
  assign n44204 = n36715 | n36716;
  assign n44205 = n36719 | n36720;
  assign n44206 = n36721 | n36722;
  assign n44207 = n36728 | ~n36729;
  assign n44208 = n36742 | n36743;
  assign n44209 = n36746 | n36747;
  assign n44210 = n36748 | n36749;
  assign n44211 = n36753 | n36754;
  assign n44212 = n36755 | n36756;
  assign n44213 = n36757 | ~n36758;
  assign n44214 = n36764 | n36765;
  assign n44215 = n36766 | n36767;
  assign n44216 = n36768 | ~n36769;
  assign n44217 = n36772 | n36773;
  assign n44218 = n36774 | n36775;
  assign n44219 = n36776 | ~n36777;
  assign n44220 = n36782 | ~n36783;
  assign n44221 = n36785 | ~n36786;
  assign n44222 = n36802 | n36803;
  assign n44223 = n36806 | n36807;
  assign n44224 = n36808 | n36809;
  assign n44225 = n36825 | n36826;
  assign n44226 = n36829 | ~n36830;
  assign n44227 = n36841 | ~n36842;
  assign n44228 = n36845 | n36846;
  assign n44229 = n36857 | n36858;
  assign n44230 = n36859 | n36860;
  assign n44231 = n36866 | ~n36867;
  assign n44232 = n36872 | ~n36873;
  assign n44233 = n36883 | n36884;
  assign n44234 = n36898 | n36899;
  assign n44235 = n36902 | n36903;
  assign n44236 = n36904 | n36905;
  assign n44237 = n36912 | n36913;
  assign n44238 = n36914 | n36915;
  assign n44239 = n36916 | ~n36917;
  assign n44240 = n36920 | n36921;
  assign n44241 = n36922 | n36923;
  assign n44242 = n36924 | ~n36925;
  assign n44243 = n36935 | n36936;
  assign n44244 = n36939 | n36940;
  assign n44245 = n36941 | n36942;
  assign n44246 = n36948 | ~n36949;
  assign n44247 = n36954 | ~n36955;
  assign n44248 = n36957 | ~n36958;
  assign n44249 = n36972 | n36973;
  assign n44250 = n36974 | n36975;
  assign n44251 = n36976 | ~n36977;
  assign n44252 = n36982 | ~n36983;
  assign n44253 = n36993 | n36994;
  assign n44254 = n36997 | n36998;
  assign n44255 = n36999 | n37000;
  assign n44256 = n37011 | n37012;
  assign n44257 = n37015 | n37016;
  assign n44258 = n37017 | n37018;
  assign n44259 = n37021 | ~n37022;
  assign n44260 = n37025 | n37026;
  assign n44261 = n37027 | n37028;
  assign n44262 = n37029 | ~n37030;
  assign n44263 = n37032 | n37033;
  assign n44264 = n37037 | n37038;
  assign n44265 = n37039 | ~n37040;
  assign n44266 = n37042 | ~n37043;
  assign n44267 = n37066 | n37067;
  assign n44268 = n37070 | ~n37071;
  assign n44269 = n37087 | n37088;
  assign n44270 = n37089 | n37090;
  assign n44271 = n37096 | ~n37097;
  assign n44272 = n37114 | n37115;
  assign n44273 = n37120 | ~n37121;
  assign n44274 = n37128 | n37129;
  assign n44275 = n37132 | n37133;
  assign n44276 = n37134 | n37135;
  assign n44277 = n37141 | ~n37142;
  assign n44278 = n37144 | n37145;
  assign n44279 = n37146 | n37147;
  assign n44280 = n37153 | ~n37154;
  assign n44281 = n37159 | ~n37160;
  assign n44282 = n37162 | ~n37163;
  assign n44283 = n37168 | ~n37169;
  assign n44284 = n37172 | n37173;
  assign n44285 = n37181 | ~n37182;
  assign n44286 = n37195 | n37196;
  assign n44287 = n37199 | n37200;
  assign n44288 = n37201 | n37202;
  assign n44289 = n37206 | n37207;
  assign n44290 = n37208 | n37209;
  assign n44291 = n37210 | ~n37211;
  assign n44292 = n37219 | ~n37220;
  assign n44293 = n37223 | n37224;
  assign n44294 = n37241 | ~n37242;
  assign n44295 = n37253 | ~n37254;
  assign n44296 = n37257 | n37258;
  assign n44297 = n37273 | n37274;
  assign n44298 = n37285 | ~n37286;
  assign n44299 = n37289 | n37290;
  assign n44300 = n37298 | n37299;
  assign n44301 = n37304 | ~n37305;
  assign n44302 = n37316 | n37317;
  assign n44303 = n37319 | n37320;
  assign n44304 = n37321 | n37322;
  assign n44305 = n37326 | ~n37327;
  assign po127  = n37332 | ~n37333;
  assign n44307 = n37341 | n37342;
  assign n44308 = n37431 | n37432;
  assign po2  = n37462 | n37463;
  assign po1  = n37468 | n37469;
endmodule
