module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 , pi32 ,
    pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 , pi40 ,
    pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 , pi56 ,
    pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 , pi64 ,
    pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 ,
    pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 ,
    pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 ,
    pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 ,
    pi97 , pi98 , pi99 , pi100 , pi101 , pi102 , pi103 ,
    pi104 , pi105 , pi106 , pi107 , pi108 , pi109 , pi110 ,
    pi111 , pi112 , pi113 , pi114 , pi115 , pi116 , pi117 ,
    pi118 , pi119 , pi120 , pi121 , pi122 , pi123 , pi124 ,
    pi125 , pi126 , pi127 , pi128 , pi129 , pi130 , pi131 , pi132 ,
    pi133 , pi134 , pi135 , pi136 , pi137 , pi138 , pi139 , pi140 ,
    pi141 , pi142 , pi143 , pi144 , pi145 , pi146 , pi147 , pi148 ,
    pi149 , pi150 , pi151 , pi152 , pi153 , pi154 , pi155 , pi156 ,
    pi157 , pi158 , pi159 , pi160 , pi161 , pi162 , pi163 , pi164 ,
    pi165 , pi166 , pi167 , pi168 , pi169 , pi170 , pi171 , pi172 ,
    pi173 , pi174 , pi175 , pi176 , pi177 , pi178 , pi179 , pi180 ,
    pi181 , pi182 , pi183 , pi184 , pi185 , pi186 , pi187 , pi188 ,
    pi189 , pi190 , pi191 , pi192 , pi193 , pi194 , pi195 , pi196 ,
    pi197 , pi198 , pi199 , pi200 , pi201 , pi202 , pi203 , pi204 ,
    pi205 , pi206 , pi207 , pi208 , pi209 , pi210 , pi211 , pi212 ,
    pi213 , pi214 , pi215 , pi216 , pi217 , pi218 , pi219 , pi220 ,
    pi221 , pi222 , pi223 , pi224 , pi225 , pi226 , pi227 ,
    pi228 , pi229 , pi230 , pi231 , pi232 , pi233 , pi234 ,
    pi235 , pi236 , pi237 , pi238 , pi239 , pi240 , pi241 ,
    pi242 , pi243 , pi244 , pi245 , pi246 , pi247 , pi248 ,
    pi249 , pi250 , pi251 , pi252 , pi253 , pi254 , pi255 ,
    po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7 , po8 ,
    po9 , po10 , po11 , po12 , po13 , po14 , po15 , po16 ,
    po17 , po18 , po19 , po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 , po30 , po31 , po32 ,
    po33 , po34 , po35 , po36 , po37 , po38 , po39 , po40 ,
    po41 , po42 , po43 , po44 , po45 , po46 , po47 , po48 ,
    po49 , po50 , po51 , po52 , po53 , po54 , po55 , po56 ,
    po57 , po58 , po59 , po60 , po61 , po62 , po63 , po64 ,
    po65 , po66 , po67 , po68 , po69 , po70 , po71 , po72 ,
    po73 , po74 , po75 , po76 , po77 , po78 , po79 , po80 ,
    po81 , po82 , po83 , po84 , po85 , po86 , po87 , po88 ,
    po89 , po90 , po91 , po92 , po93 , po94 , po95 , po96 ,
    po97 , po98 , po99 , po100 , po101 , po102 , po103 ,
    po104 , po105 , po106 , po107 , po108 , po109 , po110 ,
    po111 , po112 , po113 , po114 , po115 , po116 , po117 ,
    po118 , po119 , po120 , po121 , po122 , po123 , po124 ,
    po125 , po126 , po127 , po128  );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    pi32 , pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 ,
    pi56 , pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 ,
    pi64 , pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 ,
    pi72 , pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 ,
    pi80 , pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 ,
    pi88 , pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 ,
    pi96 , pi97 , pi98 , pi99 , pi100 , pi101 , pi102 ,
    pi103 , pi104 , pi105 , pi106 , pi107 , pi108 , pi109 ,
    pi110 , pi111 , pi112 , pi113 , pi114 , pi115 , pi116 ,
    pi117 , pi118 , pi119 , pi120 , pi121 , pi122 , pi123 ,
    pi124 , pi125 , pi126 , pi127 , pi128 , pi129 , pi130 , pi131 ,
    pi132 , pi133 , pi134 , pi135 , pi136 , pi137 , pi138 , pi139 ,
    pi140 , pi141 , pi142 , pi143 , pi144 , pi145 , pi146 , pi147 ,
    pi148 , pi149 , pi150 , pi151 , pi152 , pi153 , pi154 , pi155 ,
    pi156 , pi157 , pi158 , pi159 , pi160 , pi161 , pi162 , pi163 ,
    pi164 , pi165 , pi166 , pi167 , pi168 , pi169 , pi170 , pi171 ,
    pi172 , pi173 , pi174 , pi175 , pi176 , pi177 , pi178 , pi179 ,
    pi180 , pi181 , pi182 , pi183 , pi184 , pi185 , pi186 , pi187 ,
    pi188 , pi189 , pi190 , pi191 , pi192 , pi193 , pi194 , pi195 ,
    pi196 , pi197 , pi198 , pi199 , pi200 , pi201 , pi202 , pi203 ,
    pi204 , pi205 , pi206 , pi207 , pi208 , pi209 , pi210 , pi211 ,
    pi212 , pi213 , pi214 , pi215 , pi216 , pi217 , pi218 , pi219 ,
    pi220 , pi221 , pi222 , pi223 , pi224 , pi225 , pi226 , pi227 ,
    pi228 , pi229 , pi230 , pi231 , pi232 , pi233 , pi234 ,
    pi235 , pi236 , pi237 , pi238 , pi239 , pi240 , pi241 ,
    pi242 , pi243 , pi244 , pi245 , pi246 , pi247 , pi248 ,
    pi249 , pi250 , pi251 , pi252 , pi253 , pi254 , pi255 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7 ,
    po8 , po9 , po10 , po11 , po12 , po13 , po14 , po15 ,
    po16 , po17 , po18 , po19 , po20 , po21 , po22 , po23 ,
    po24 , po25 , po26 , po27 , po28 , po29 , po30 , po31 ,
    po32 , po33 , po34 , po35 , po36 , po37 , po38 , po39 ,
    po40 , po41 , po42 , po43 , po44 , po45 , po46 , po47 ,
    po48 , po49 , po50 , po51 , po52 , po53 , po54 , po55 ,
    po56 , po57 , po58 , po59 , po60 , po61 , po62 , po63 ,
    po64 , po65 , po66 , po67 , po68 , po69 , po70 , po71 ,
    po72 , po73 , po74 , po75 , po76 , po77 , po78 , po79 ,
    po80 , po81 , po82 , po83 , po84 , po85 , po86 , po87 ,
    po88 , po89 , po90 , po91 , po92 , po93 , po94 , po95 ,
    po96 , po97 , po98 , po99 , po100 , po101 , po102 ,
    po103 , po104 , po105 , po106 , po107 , po108 , po109 ,
    po110 , po111 , po112 , po113 , po114 , po115 , po116 ,
    po117 , po118 , po119 , po120 , po121 , po122 , po123 ,
    po124 , po125 , po126 , po127 , po128;
  wire n386, n387, n389, n390, n391, n392, n393,
    n395, n396, n397, n398, n399, n400, n402,
    n403, n404, n405, n406, n407, n409, n410,
    n411, n412, n413, n414, n416, n417, n418,
    n419, n420, n421, n423, n424, n425, n426,
    n427, n428, n430, n431, n432, n433, n434,
    n435, n437, n438, n439, n440, n441, n442,
    n444, n445, n446, n447, n448, n449, n451,
    n452, n453, n454, n455, n456, n458, n459,
    n460, n461, n462, n463, n465, n466, n467,
    n468, n469, n470, n472, n473, n474, n475,
    n476, n477, n479, n480, n481, n482, n483,
    n484, n486, n487, n488, n489, n490, n491,
    n493, n494, n495, n496, n497, n498, n500,
    n501, n502, n503, n504, n505, n507, n508,
    n509, n510, n511, n512, n514, n515, n516,
    n517, n518, n519, n521, n522, n523, n524,
    n525, n526, n528, n529, n530, n531, n532,
    n533, n535, n536, n537, n538, n539, n540,
    n542, n543, n544, n545, n546, n547, n549,
    n550, n551, n552, n553, n554, n556, n557,
    n558, n559, n560, n561, n563, n564, n565,
    n566, n567, n568, n570, n571, n572, n573,
    n574, n575, n577, n578, n579, n580, n581,
    n582, n584, n585, n586, n587, n588, n589,
    n591, n592, n593, n594, n595, n596, n598,
    n599, n600, n601, n602, n603, n605, n606,
    n607, n608, n609, n610, n612, n613, n614,
    n615, n616, n617, n619, n620, n621, n622,
    n623, n624, n626, n627, n628, n629, n630,
    n631, n633, n634, n635, n636, n637, n638,
    n640, n641, n642, n643, n644, n645, n647,
    n648, n649, n650, n651, n652, n654, n655,
    n656, n657, n658, n659, n661, n662, n663,
    n664, n665, n666, n668, n669, n670, n671,
    n672, n673, n675, n676, n677, n678, n679,
    n680, n682, n683, n684, n685, n686, n687,
    n689, n690, n691, n692, n693, n694, n696,
    n697, n698, n699, n700, n701, n703, n704,
    n705, n706, n707, n708, n710, n711, n712,
    n713, n714, n715, n717, n718, n719, n720,
    n721, n722, n724, n725, n726, n727, n728,
    n729, n731, n732, n733, n734, n735, n736,
    n738, n739, n740, n741, n742, n743, n745,
    n746, n747, n748, n749, n750, n752, n753,
    n754, n755, n756, n757, n759, n760, n761,
    n762, n763, n764, n766, n767, n768, n769,
    n770, n771, n773, n774, n775, n776, n777,
    n778, n780, n781, n782, n783, n784, n785,
    n787, n788, n789, n790, n791, n792, n794,
    n795, n796, n797, n798, n799, n801, n802,
    n803, n804, n805, n806, n808, n809, n810,
    n811, n812, n813, n815, n816, n817, n818,
    n819, n820, n822, n823, n824, n825, n826,
    n827, n829, n830, n831, n832, n833, n834,
    n836, n837, n838, n839, n840, n841, n843,
    n844, n845, n846, n847, n848, n850, n851,
    n852, n853, n854, n855, n857, n858, n859,
    n860, n861, n862, n864, n865, n866, n867,
    n868, n869, n871, n872, n873, n874, n875,
    n876, n878, n879, n880, n881, n882, n883,
    n885, n886, n887, n888, n889, n890, n892,
    n893, n894, n895, n896, n897, n899, n900,
    n901, n902, n903, n904, n906, n907, n908,
    n909, n910, n911, n913, n914, n915, n916,
    n917, n918, n920, n921, n922, n923, n924,
    n925, n927, n928, n929, n930, n931, n932,
    n934, n935, n936, n937, n938, n939, n941,
    n942, n943, n944, n945, n946, n948, n949,
    n950, n951, n952, n953, n955, n956, n957,
    n958, n959, n960, n962, n963, n964, n965,
    n966, n967, n969, n970, n971, n972, n973,
    n974, n976, n977, n978, n979, n980, n981,
    n983, n984, n985, n986, n987, n988, n990,
    n991, n992, n993, n994, n995, n997, n998,
    n999, n1000, n1001, n1002, n1004, n1005,
    n1006, n1007, n1008, n1009, n1011, n1012,
    n1013, n1014, n1015, n1016, n1018, n1019,
    n1020, n1021, n1022, n1023, n1025, n1026,
    n1027, n1028, n1029, n1030, n1032, n1033,
    n1034, n1035, n1036, n1037, n1039, n1040,
    n1041, n1042, n1043, n1044, n1046, n1047,
    n1048, n1049, n1050, n1051, n1053, n1054,
    n1055, n1056, n1057, n1058, n1060, n1061,
    n1062, n1063, n1064, n1065, n1067, n1068,
    n1069, n1070, n1071, n1072, n1074, n1075,
    n1076, n1077, n1078, n1079, n1081, n1082,
    n1083, n1084, n1085, n1086, n1088, n1089,
    n1090, n1091, n1092, n1093, n1095, n1096,
    n1097, n1098, n1099, n1100, n1102, n1103,
    n1104, n1105, n1106, n1107, n1109, n1110,
    n1111, n1112, n1113, n1114, n1116, n1117,
    n1118, n1119, n1120, n1121, n1123, n1124,
    n1125, n1126, n1127, n1128, n1130, n1131,
    n1132, n1133, n1134, n1135, n1137, n1138,
    n1139, n1140, n1141, n1142, n1144, n1145,
    n1146, n1147, n1148, n1149, n1151, n1152,
    n1153, n1154, n1155, n1156, n1158, n1159,
    n1160, n1161, n1162, n1163, n1165, n1166,
    n1167, n1168, n1169, n1170, n1172, n1173,
    n1174, n1175, n1176, n1177, n1179, n1180,
    n1181, n1182, n1183, n1184, n1186, n1187,
    n1188, n1189, n1190, n1191, n1193, n1194,
    n1195, n1196, n1197, n1198, n1200, n1201,
    n1202, n1203, n1204, n1205, n1207, n1208,
    n1209, n1210, n1211, n1212, n1214, n1215,
    n1216, n1217, n1218, n1219, n1221, n1222,
    n1223, n1224, n1225, n1226, n1228, n1229,
    n1230, n1231, n1232, n1233, n1235, n1236,
    n1237, n1238, n1239, n1240, n1242, n1243,
    n1244, n1245, n1246, n1247, n1249, n1250,
    n1251, n1252, n1253, n1254, n1256, n1257,
    n1258, n1259, n1260, n1261, n1263, n1264,
    n1265, n1266, n1267, n1268, n1270, n1271,
    n1272, n1273, n1274, n1275;
  assign n386 = pi0  & pi128 ;
  assign n387 = ~pi0  & ~pi128 ;
  assign po0  = ~n386 & ~n387;
  assign n389 = ~pi1  & ~pi129 ;
  assign n390 = pi1  & pi129 ;
  assign n391 = ~n389 & ~n390;
  assign n392 = n386 & ~n391;
  assign n393 = ~n386 & n391;
  assign po1  = n392 | n393;
  assign n395 = ~pi2  & ~pi130 ;
  assign n396 = pi2  & pi130 ;
  assign n397 = ~n395 & ~n396;
  assign n398 = ~n389 & ~n393;
  assign n399 = ~n397 & ~n398;
  assign n400 = n397 & n398;
  assign po2  = ~n399 & ~n400;
  assign n402 = ~pi3  & ~pi131 ;
  assign n403 = pi3  & pi131 ;
  assign n404 = ~n402 & ~n403;
  assign n405 = ~n396 & ~n400;
  assign n406 = ~n404 & n405;
  assign n407 = n404 & ~n405;
  assign po3  = ~n406 & ~n407;
  assign n409 = ~pi4  & ~pi132 ;
  assign n410 = pi4  & pi132 ;
  assign n411 = ~n409 & ~n410;
  assign n412 = ~n403 & ~n407;
  assign n413 = ~n411 & n412;
  assign n414 = n411 & ~n412;
  assign po4  = ~n413 & ~n414;
  assign n416 = ~pi5  & ~pi133 ;
  assign n417 = pi5  & pi133 ;
  assign n418 = ~n416 & ~n417;
  assign n419 = ~n410 & ~n414;
  assign n420 = ~n418 & n419;
  assign n421 = n418 & ~n419;
  assign po5  = ~n420 & ~n421;
  assign n423 = ~pi6  & ~pi134 ;
  assign n424 = pi6  & pi134 ;
  assign n425 = ~n423 & ~n424;
  assign n426 = ~n417 & ~n421;
  assign n427 = ~n425 & n426;
  assign n428 = n425 & ~n426;
  assign po6  = ~n427 & ~n428;
  assign n430 = ~pi7  & ~pi135 ;
  assign n431 = pi7  & pi135 ;
  assign n432 = ~n430 & ~n431;
  assign n433 = ~n424 & ~n428;
  assign n434 = ~n432 & n433;
  assign n435 = n432 & ~n433;
  assign po7  = ~n434 & ~n435;
  assign n437 = ~pi8  & ~pi136 ;
  assign n438 = pi8  & pi136 ;
  assign n439 = ~n437 & ~n438;
  assign n440 = ~n431 & ~n435;
  assign n441 = ~n439 & n440;
  assign n442 = n439 & ~n440;
  assign po8  = ~n441 & ~n442;
  assign n444 = ~pi9  & ~pi137 ;
  assign n445 = pi9  & pi137 ;
  assign n446 = ~n444 & ~n445;
  assign n447 = ~n438 & ~n442;
  assign n448 = ~n446 & n447;
  assign n449 = n446 & ~n447;
  assign po9  = ~n448 & ~n449;
  assign n451 = ~pi10  & ~pi138 ;
  assign n452 = pi10  & pi138 ;
  assign n453 = ~n451 & ~n452;
  assign n454 = ~n445 & ~n449;
  assign n455 = ~n453 & n454;
  assign n456 = n453 & ~n454;
  assign po10  = ~n455 & ~n456;
  assign n458 = ~pi11  & ~pi139 ;
  assign n459 = pi11  & pi139 ;
  assign n460 = ~n458 & ~n459;
  assign n461 = ~n452 & ~n456;
  assign n462 = ~n460 & n461;
  assign n463 = n460 & ~n461;
  assign po11  = ~n462 & ~n463;
  assign n465 = ~pi12  & ~pi140 ;
  assign n466 = pi12  & pi140 ;
  assign n467 = ~n465 & ~n466;
  assign n468 = ~n459 & ~n463;
  assign n469 = ~n467 & n468;
  assign n470 = n467 & ~n468;
  assign po12  = ~n469 & ~n470;
  assign n472 = ~pi13  & ~pi141 ;
  assign n473 = pi13  & pi141 ;
  assign n474 = ~n472 & ~n473;
  assign n475 = ~n466 & ~n470;
  assign n476 = ~n474 & n475;
  assign n477 = n474 & ~n475;
  assign po13  = ~n476 & ~n477;
  assign n479 = ~pi14  & ~pi142 ;
  assign n480 = pi14  & pi142 ;
  assign n481 = ~n479 & ~n480;
  assign n482 = ~n473 & ~n477;
  assign n483 = ~n481 & n482;
  assign n484 = n481 & ~n482;
  assign po14  = ~n483 & ~n484;
  assign n486 = ~pi15  & ~pi143 ;
  assign n487 = pi15  & pi143 ;
  assign n488 = ~n486 & ~n487;
  assign n489 = ~n480 & ~n484;
  assign n490 = ~n488 & n489;
  assign n491 = n488 & ~n489;
  assign po15  = ~n490 & ~n491;
  assign n493 = ~pi16  & ~pi144 ;
  assign n494 = pi16  & pi144 ;
  assign n495 = ~n493 & ~n494;
  assign n496 = ~n487 & ~n491;
  assign n497 = ~n495 & n496;
  assign n498 = n495 & ~n496;
  assign po16  = ~n497 & ~n498;
  assign n500 = ~pi17  & ~pi145 ;
  assign n501 = pi17  & pi145 ;
  assign n502 = ~n500 & ~n501;
  assign n503 = ~n494 & ~n498;
  assign n504 = ~n502 & n503;
  assign n505 = n502 & ~n503;
  assign po17  = ~n504 & ~n505;
  assign n507 = ~pi18  & ~pi146 ;
  assign n508 = pi18  & pi146 ;
  assign n509 = ~n507 & ~n508;
  assign n510 = ~n501 & ~n505;
  assign n511 = ~n509 & n510;
  assign n512 = n509 & ~n510;
  assign po18  = ~n511 & ~n512;
  assign n514 = ~pi19  & ~pi147 ;
  assign n515 = pi19  & pi147 ;
  assign n516 = ~n514 & ~n515;
  assign n517 = ~n508 & ~n512;
  assign n518 = ~n516 & n517;
  assign n519 = n516 & ~n517;
  assign po19  = ~n518 & ~n519;
  assign n521 = ~pi20  & ~pi148 ;
  assign n522 = pi20  & pi148 ;
  assign n523 = ~n521 & ~n522;
  assign n524 = ~n515 & ~n519;
  assign n525 = ~n523 & n524;
  assign n526 = n523 & ~n524;
  assign po20  = ~n525 & ~n526;
  assign n528 = ~pi21  & ~pi149 ;
  assign n529 = pi21  & pi149 ;
  assign n530 = ~n528 & ~n529;
  assign n531 = ~n522 & ~n526;
  assign n532 = ~n530 & n531;
  assign n533 = n530 & ~n531;
  assign po21  = ~n532 & ~n533;
  assign n535 = ~pi22  & ~pi150 ;
  assign n536 = pi22  & pi150 ;
  assign n537 = ~n535 & ~n536;
  assign n538 = ~n529 & ~n533;
  assign n539 = ~n537 & n538;
  assign n540 = n537 & ~n538;
  assign po22  = ~n539 & ~n540;
  assign n542 = ~pi23  & ~pi151 ;
  assign n543 = pi23  & pi151 ;
  assign n544 = ~n542 & ~n543;
  assign n545 = ~n536 & ~n540;
  assign n546 = ~n544 & n545;
  assign n547 = n544 & ~n545;
  assign po23  = ~n546 & ~n547;
  assign n549 = ~pi24  & ~pi152 ;
  assign n550 = pi24  & pi152 ;
  assign n551 = ~n549 & ~n550;
  assign n552 = ~n543 & ~n547;
  assign n553 = ~n551 & n552;
  assign n554 = n551 & ~n552;
  assign po24  = ~n553 & ~n554;
  assign n556 = ~pi25  & ~pi153 ;
  assign n557 = pi25  & pi153 ;
  assign n558 = ~n556 & ~n557;
  assign n559 = ~n550 & ~n554;
  assign n560 = ~n558 & n559;
  assign n561 = n558 & ~n559;
  assign po25  = ~n560 & ~n561;
  assign n563 = ~pi26  & ~pi154 ;
  assign n564 = pi26  & pi154 ;
  assign n565 = ~n563 & ~n564;
  assign n566 = ~n557 & ~n561;
  assign n567 = ~n565 & n566;
  assign n568 = n565 & ~n566;
  assign po26  = ~n567 & ~n568;
  assign n570 = ~pi27  & ~pi155 ;
  assign n571 = pi27  & pi155 ;
  assign n572 = ~n570 & ~n571;
  assign n573 = ~n564 & ~n568;
  assign n574 = ~n572 & n573;
  assign n575 = n572 & ~n573;
  assign po27  = ~n574 & ~n575;
  assign n577 = ~pi28  & ~pi156 ;
  assign n578 = pi28  & pi156 ;
  assign n579 = ~n577 & ~n578;
  assign n580 = ~n571 & ~n575;
  assign n581 = ~n579 & n580;
  assign n582 = n579 & ~n580;
  assign po28  = ~n581 & ~n582;
  assign n584 = ~pi29  & ~pi157 ;
  assign n585 = pi29  & pi157 ;
  assign n586 = ~n584 & ~n585;
  assign n587 = ~n578 & ~n582;
  assign n588 = ~n586 & n587;
  assign n589 = n586 & ~n587;
  assign po29  = ~n588 & ~n589;
  assign n591 = ~pi30  & ~pi158 ;
  assign n592 = pi30  & pi158 ;
  assign n593 = ~n591 & ~n592;
  assign n594 = ~n585 & ~n589;
  assign n595 = ~n593 & n594;
  assign n596 = n593 & ~n594;
  assign po30  = ~n595 & ~n596;
  assign n598 = ~pi31  & ~pi159 ;
  assign n599 = pi31  & pi159 ;
  assign n600 = ~n598 & ~n599;
  assign n601 = ~n592 & ~n596;
  assign n602 = ~n600 & n601;
  assign n603 = n600 & ~n601;
  assign po31  = ~n602 & ~n603;
  assign n605 = ~pi32  & ~pi160 ;
  assign n606 = pi32  & pi160 ;
  assign n607 = ~n605 & ~n606;
  assign n608 = ~n599 & ~n603;
  assign n609 = ~n607 & n608;
  assign n610 = n607 & ~n608;
  assign po32  = ~n609 & ~n610;
  assign n612 = ~pi33  & ~pi161 ;
  assign n613 = pi33  & pi161 ;
  assign n614 = ~n612 & ~n613;
  assign n615 = ~n606 & ~n610;
  assign n616 = ~n614 & n615;
  assign n617 = n614 & ~n615;
  assign po33  = ~n616 & ~n617;
  assign n619 = ~pi34  & ~pi162 ;
  assign n620 = pi34  & pi162 ;
  assign n621 = ~n619 & ~n620;
  assign n622 = ~n613 & ~n617;
  assign n623 = ~n621 & n622;
  assign n624 = n621 & ~n622;
  assign po34  = ~n623 & ~n624;
  assign n626 = ~pi35  & ~pi163 ;
  assign n627 = pi35  & pi163 ;
  assign n628 = ~n626 & ~n627;
  assign n629 = ~n620 & ~n624;
  assign n630 = ~n628 & n629;
  assign n631 = n628 & ~n629;
  assign po35  = ~n630 & ~n631;
  assign n633 = ~pi36  & ~pi164 ;
  assign n634 = pi36  & pi164 ;
  assign n635 = ~n633 & ~n634;
  assign n636 = ~n627 & ~n631;
  assign n637 = ~n635 & n636;
  assign n638 = n635 & ~n636;
  assign po36  = ~n637 & ~n638;
  assign n640 = ~pi37  & ~pi165 ;
  assign n641 = pi37  & pi165 ;
  assign n642 = ~n640 & ~n641;
  assign n643 = ~n634 & ~n638;
  assign n644 = ~n642 & n643;
  assign n645 = n642 & ~n643;
  assign po37  = ~n644 & ~n645;
  assign n647 = ~pi38  & ~pi166 ;
  assign n648 = pi38  & pi166 ;
  assign n649 = ~n647 & ~n648;
  assign n650 = ~n641 & ~n645;
  assign n651 = ~n649 & n650;
  assign n652 = n649 & ~n650;
  assign po38  = ~n651 & ~n652;
  assign n654 = ~pi39  & ~pi167 ;
  assign n655 = pi39  & pi167 ;
  assign n656 = ~n654 & ~n655;
  assign n657 = ~n648 & ~n652;
  assign n658 = ~n656 & n657;
  assign n659 = n656 & ~n657;
  assign po39  = ~n658 & ~n659;
  assign n661 = ~pi40  & ~pi168 ;
  assign n662 = pi40  & pi168 ;
  assign n663 = ~n661 & ~n662;
  assign n664 = ~n655 & ~n659;
  assign n665 = ~n663 & n664;
  assign n666 = n663 & ~n664;
  assign po40  = ~n665 & ~n666;
  assign n668 = ~pi41  & ~pi169 ;
  assign n669 = pi41  & pi169 ;
  assign n670 = ~n668 & ~n669;
  assign n671 = ~n662 & ~n666;
  assign n672 = ~n670 & n671;
  assign n673 = n670 & ~n671;
  assign po41  = ~n672 & ~n673;
  assign n675 = ~pi42  & ~pi170 ;
  assign n676 = pi42  & pi170 ;
  assign n677 = ~n675 & ~n676;
  assign n678 = ~n669 & ~n673;
  assign n679 = ~n677 & n678;
  assign n680 = n677 & ~n678;
  assign po42  = ~n679 & ~n680;
  assign n682 = ~pi43  & ~pi171 ;
  assign n683 = pi43  & pi171 ;
  assign n684 = ~n682 & ~n683;
  assign n685 = ~n676 & ~n680;
  assign n686 = ~n684 & n685;
  assign n687 = n684 & ~n685;
  assign po43  = ~n686 & ~n687;
  assign n689 = ~pi44  & ~pi172 ;
  assign n690 = pi44  & pi172 ;
  assign n691 = ~n689 & ~n690;
  assign n692 = ~n683 & ~n687;
  assign n693 = ~n691 & n692;
  assign n694 = n691 & ~n692;
  assign po44  = ~n693 & ~n694;
  assign n696 = ~pi45  & ~pi173 ;
  assign n697 = pi45  & pi173 ;
  assign n698 = ~n696 & ~n697;
  assign n699 = ~n690 & ~n694;
  assign n700 = ~n698 & n699;
  assign n701 = n698 & ~n699;
  assign po45  = ~n700 & ~n701;
  assign n703 = ~pi46  & ~pi174 ;
  assign n704 = pi46  & pi174 ;
  assign n705 = ~n703 & ~n704;
  assign n706 = ~n697 & ~n701;
  assign n707 = ~n705 & n706;
  assign n708 = n705 & ~n706;
  assign po46  = ~n707 & ~n708;
  assign n710 = ~pi47  & ~pi175 ;
  assign n711 = pi47  & pi175 ;
  assign n712 = ~n710 & ~n711;
  assign n713 = ~n704 & ~n708;
  assign n714 = ~n712 & n713;
  assign n715 = n712 & ~n713;
  assign po47  = ~n714 & ~n715;
  assign n717 = ~pi48  & ~pi176 ;
  assign n718 = pi48  & pi176 ;
  assign n719 = ~n717 & ~n718;
  assign n720 = ~n711 & ~n715;
  assign n721 = ~n719 & n720;
  assign n722 = n719 & ~n720;
  assign po48  = ~n721 & ~n722;
  assign n724 = ~pi49  & ~pi177 ;
  assign n725 = pi49  & pi177 ;
  assign n726 = ~n724 & ~n725;
  assign n727 = ~n718 & ~n722;
  assign n728 = ~n726 & n727;
  assign n729 = n726 & ~n727;
  assign po49  = ~n728 & ~n729;
  assign n731 = ~pi50  & ~pi178 ;
  assign n732 = pi50  & pi178 ;
  assign n733 = ~n731 & ~n732;
  assign n734 = ~n725 & ~n729;
  assign n735 = ~n733 & n734;
  assign n736 = n733 & ~n734;
  assign po50  = ~n735 & ~n736;
  assign n738 = ~pi51  & ~pi179 ;
  assign n739 = pi51  & pi179 ;
  assign n740 = ~n738 & ~n739;
  assign n741 = ~n732 & ~n736;
  assign n742 = ~n740 & n741;
  assign n743 = n740 & ~n741;
  assign po51  = ~n742 & ~n743;
  assign n745 = ~pi52  & ~pi180 ;
  assign n746 = pi52  & pi180 ;
  assign n747 = ~n745 & ~n746;
  assign n748 = ~n739 & ~n743;
  assign n749 = ~n747 & n748;
  assign n750 = n747 & ~n748;
  assign po52  = ~n749 & ~n750;
  assign n752 = ~pi53  & ~pi181 ;
  assign n753 = pi53  & pi181 ;
  assign n754 = ~n752 & ~n753;
  assign n755 = ~n746 & ~n750;
  assign n756 = ~n754 & n755;
  assign n757 = n754 & ~n755;
  assign po53  = ~n756 & ~n757;
  assign n759 = ~pi54  & ~pi182 ;
  assign n760 = pi54  & pi182 ;
  assign n761 = ~n759 & ~n760;
  assign n762 = ~n753 & ~n757;
  assign n763 = ~n761 & n762;
  assign n764 = n761 & ~n762;
  assign po54  = ~n763 & ~n764;
  assign n766 = ~pi55  & ~pi183 ;
  assign n767 = pi55  & pi183 ;
  assign n768 = ~n766 & ~n767;
  assign n769 = ~n760 & ~n764;
  assign n770 = ~n768 & n769;
  assign n771 = n768 & ~n769;
  assign po55  = ~n770 & ~n771;
  assign n773 = ~pi56  & ~pi184 ;
  assign n774 = pi56  & pi184 ;
  assign n775 = ~n773 & ~n774;
  assign n776 = ~n767 & ~n771;
  assign n777 = ~n775 & n776;
  assign n778 = n775 & ~n776;
  assign po56  = ~n777 & ~n778;
  assign n780 = ~pi57  & ~pi185 ;
  assign n781 = pi57  & pi185 ;
  assign n782 = ~n780 & ~n781;
  assign n783 = ~n774 & ~n778;
  assign n784 = ~n782 & n783;
  assign n785 = n782 & ~n783;
  assign po57  = ~n784 & ~n785;
  assign n787 = ~pi58  & ~pi186 ;
  assign n788 = pi58  & pi186 ;
  assign n789 = ~n787 & ~n788;
  assign n790 = ~n781 & ~n785;
  assign n791 = ~n789 & n790;
  assign n792 = n789 & ~n790;
  assign po58  = ~n791 & ~n792;
  assign n794 = ~pi59  & ~pi187 ;
  assign n795 = pi59  & pi187 ;
  assign n796 = ~n794 & ~n795;
  assign n797 = ~n788 & ~n792;
  assign n798 = ~n796 & n797;
  assign n799 = n796 & ~n797;
  assign po59  = ~n798 & ~n799;
  assign n801 = ~pi60  & ~pi188 ;
  assign n802 = pi60  & pi188 ;
  assign n803 = ~n801 & ~n802;
  assign n804 = ~n795 & ~n799;
  assign n805 = ~n803 & n804;
  assign n806 = n803 & ~n804;
  assign po60  = ~n805 & ~n806;
  assign n808 = ~pi61  & ~pi189 ;
  assign n809 = pi61  & pi189 ;
  assign n810 = ~n808 & ~n809;
  assign n811 = ~n802 & ~n806;
  assign n812 = ~n810 & n811;
  assign n813 = n810 & ~n811;
  assign po61  = ~n812 & ~n813;
  assign n815 = ~pi62  & ~pi190 ;
  assign n816 = pi62  & pi190 ;
  assign n817 = ~n815 & ~n816;
  assign n818 = ~n809 & ~n813;
  assign n819 = ~n817 & n818;
  assign n820 = n817 & ~n818;
  assign po62  = ~n819 & ~n820;
  assign n822 = ~pi63  & ~pi191 ;
  assign n823 = pi63  & pi191 ;
  assign n824 = ~n822 & ~n823;
  assign n825 = ~n816 & ~n820;
  assign n826 = ~n824 & n825;
  assign n827 = n824 & ~n825;
  assign po63  = ~n826 & ~n827;
  assign n829 = ~pi64  & ~pi192 ;
  assign n830 = pi64  & pi192 ;
  assign n831 = ~n829 & ~n830;
  assign n832 = ~n823 & ~n827;
  assign n833 = ~n831 & n832;
  assign n834 = n831 & ~n832;
  assign po64  = ~n833 & ~n834;
  assign n836 = ~pi65  & ~pi193 ;
  assign n837 = pi65  & pi193 ;
  assign n838 = ~n836 & ~n837;
  assign n839 = ~n830 & ~n834;
  assign n840 = ~n838 & n839;
  assign n841 = n838 & ~n839;
  assign po65  = ~n840 & ~n841;
  assign n843 = ~pi66  & ~pi194 ;
  assign n844 = pi66  & pi194 ;
  assign n845 = ~n843 & ~n844;
  assign n846 = ~n837 & ~n841;
  assign n847 = ~n845 & n846;
  assign n848 = n845 & ~n846;
  assign po66  = ~n847 & ~n848;
  assign n850 = ~pi67  & ~pi195 ;
  assign n851 = pi67  & pi195 ;
  assign n852 = ~n850 & ~n851;
  assign n853 = ~n844 & ~n848;
  assign n854 = ~n852 & n853;
  assign n855 = n852 & ~n853;
  assign po67  = ~n854 & ~n855;
  assign n857 = ~pi68  & ~pi196 ;
  assign n858 = pi68  & pi196 ;
  assign n859 = ~n857 & ~n858;
  assign n860 = ~n851 & ~n855;
  assign n861 = ~n859 & n860;
  assign n862 = n859 & ~n860;
  assign po68  = ~n861 & ~n862;
  assign n864 = ~pi69  & ~pi197 ;
  assign n865 = pi69  & pi197 ;
  assign n866 = ~n864 & ~n865;
  assign n867 = ~n858 & ~n862;
  assign n868 = ~n866 & n867;
  assign n869 = n866 & ~n867;
  assign po69  = ~n868 & ~n869;
  assign n871 = ~pi70  & ~pi198 ;
  assign n872 = pi70  & pi198 ;
  assign n873 = ~n871 & ~n872;
  assign n874 = ~n865 & ~n869;
  assign n875 = ~n873 & n874;
  assign n876 = n873 & ~n874;
  assign po70  = ~n875 & ~n876;
  assign n878 = ~pi71  & ~pi199 ;
  assign n879 = pi71  & pi199 ;
  assign n880 = ~n878 & ~n879;
  assign n881 = ~n872 & ~n876;
  assign n882 = ~n880 & n881;
  assign n883 = n880 & ~n881;
  assign po71  = ~n882 & ~n883;
  assign n885 = ~pi72  & ~pi200 ;
  assign n886 = pi72  & pi200 ;
  assign n887 = ~n885 & ~n886;
  assign n888 = ~n879 & ~n883;
  assign n889 = ~n887 & n888;
  assign n890 = n887 & ~n888;
  assign po72  = ~n889 & ~n890;
  assign n892 = ~pi73  & ~pi201 ;
  assign n893 = pi73  & pi201 ;
  assign n894 = ~n892 & ~n893;
  assign n895 = ~n886 & ~n890;
  assign n896 = ~n894 & n895;
  assign n897 = n894 & ~n895;
  assign po73  = ~n896 & ~n897;
  assign n899 = ~pi74  & ~pi202 ;
  assign n900 = pi74  & pi202 ;
  assign n901 = ~n899 & ~n900;
  assign n902 = ~n893 & ~n897;
  assign n903 = ~n901 & n902;
  assign n904 = n901 & ~n902;
  assign po74  = ~n903 & ~n904;
  assign n906 = ~pi75  & ~pi203 ;
  assign n907 = pi75  & pi203 ;
  assign n908 = ~n906 & ~n907;
  assign n909 = ~n900 & ~n904;
  assign n910 = ~n908 & n909;
  assign n911 = n908 & ~n909;
  assign po75  = ~n910 & ~n911;
  assign n913 = ~pi76  & ~pi204 ;
  assign n914 = pi76  & pi204 ;
  assign n915 = ~n913 & ~n914;
  assign n916 = ~n907 & ~n911;
  assign n917 = ~n915 & n916;
  assign n918 = n915 & ~n916;
  assign po76  = ~n917 & ~n918;
  assign n920 = ~pi77  & ~pi205 ;
  assign n921 = pi77  & pi205 ;
  assign n922 = ~n920 & ~n921;
  assign n923 = ~n914 & ~n918;
  assign n924 = ~n922 & n923;
  assign n925 = n922 & ~n923;
  assign po77  = ~n924 & ~n925;
  assign n927 = ~pi78  & ~pi206 ;
  assign n928 = pi78  & pi206 ;
  assign n929 = ~n927 & ~n928;
  assign n930 = ~n921 & ~n925;
  assign n931 = ~n929 & n930;
  assign n932 = n929 & ~n930;
  assign po78  = ~n931 & ~n932;
  assign n934 = ~pi79  & ~pi207 ;
  assign n935 = pi79  & pi207 ;
  assign n936 = ~n934 & ~n935;
  assign n937 = ~n928 & ~n932;
  assign n938 = ~n936 & n937;
  assign n939 = n936 & ~n937;
  assign po79  = ~n938 & ~n939;
  assign n941 = ~pi80  & ~pi208 ;
  assign n942 = pi80  & pi208 ;
  assign n943 = ~n941 & ~n942;
  assign n944 = ~n935 & ~n939;
  assign n945 = ~n943 & n944;
  assign n946 = n943 & ~n944;
  assign po80  = ~n945 & ~n946;
  assign n948 = ~pi81  & ~pi209 ;
  assign n949 = pi81  & pi209 ;
  assign n950 = ~n948 & ~n949;
  assign n951 = ~n942 & ~n946;
  assign n952 = ~n950 & n951;
  assign n953 = n950 & ~n951;
  assign po81  = ~n952 & ~n953;
  assign n955 = ~pi82  & ~pi210 ;
  assign n956 = pi82  & pi210 ;
  assign n957 = ~n955 & ~n956;
  assign n958 = ~n949 & ~n953;
  assign n959 = ~n957 & n958;
  assign n960 = n957 & ~n958;
  assign po82  = ~n959 & ~n960;
  assign n962 = ~pi83  & ~pi211 ;
  assign n963 = pi83  & pi211 ;
  assign n964 = ~n962 & ~n963;
  assign n965 = ~n956 & ~n960;
  assign n966 = ~n964 & n965;
  assign n967 = n964 & ~n965;
  assign po83  = ~n966 & ~n967;
  assign n969 = ~pi84  & ~pi212 ;
  assign n970 = pi84  & pi212 ;
  assign n971 = ~n969 & ~n970;
  assign n972 = ~n963 & ~n967;
  assign n973 = ~n971 & n972;
  assign n974 = n971 & ~n972;
  assign po84  = ~n973 & ~n974;
  assign n976 = ~pi85  & ~pi213 ;
  assign n977 = pi85  & pi213 ;
  assign n978 = ~n976 & ~n977;
  assign n979 = ~n970 & ~n974;
  assign n980 = ~n978 & n979;
  assign n981 = n978 & ~n979;
  assign po85  = ~n980 & ~n981;
  assign n983 = ~pi86  & ~pi214 ;
  assign n984 = pi86  & pi214 ;
  assign n985 = ~n983 & ~n984;
  assign n986 = ~n977 & ~n981;
  assign n987 = ~n985 & n986;
  assign n988 = n985 & ~n986;
  assign po86  = ~n987 & ~n988;
  assign n990 = ~pi87  & ~pi215 ;
  assign n991 = pi87  & pi215 ;
  assign n992 = ~n990 & ~n991;
  assign n993 = ~n984 & ~n988;
  assign n994 = ~n992 & n993;
  assign n995 = n992 & ~n993;
  assign po87  = ~n994 & ~n995;
  assign n997 = ~pi88  & ~pi216 ;
  assign n998 = pi88  & pi216 ;
  assign n999 = ~n997 & ~n998;
  assign n1000 = ~n991 & ~n995;
  assign n1001 = ~n999 & n1000;
  assign n1002 = n999 & ~n1000;
  assign po88  = ~n1001 & ~n1002;
  assign n1004 = ~pi89  & ~pi217 ;
  assign n1005 = pi89  & pi217 ;
  assign n1006 = ~n1004 & ~n1005;
  assign n1007 = ~n998 & ~n1002;
  assign n1008 = ~n1006 & n1007;
  assign n1009 = n1006 & ~n1007;
  assign po89  = ~n1008 & ~n1009;
  assign n1011 = ~pi90  & ~pi218 ;
  assign n1012 = pi90  & pi218 ;
  assign n1013 = ~n1011 & ~n1012;
  assign n1014 = ~n1005 & ~n1009;
  assign n1015 = ~n1013 & n1014;
  assign n1016 = n1013 & ~n1014;
  assign po90  = ~n1015 & ~n1016;
  assign n1018 = ~pi91  & ~pi219 ;
  assign n1019 = pi91  & pi219 ;
  assign n1020 = ~n1018 & ~n1019;
  assign n1021 = ~n1012 & ~n1016;
  assign n1022 = ~n1020 & n1021;
  assign n1023 = n1020 & ~n1021;
  assign po91  = ~n1022 & ~n1023;
  assign n1025 = ~pi92  & ~pi220 ;
  assign n1026 = pi92  & pi220 ;
  assign n1027 = ~n1025 & ~n1026;
  assign n1028 = ~n1019 & ~n1023;
  assign n1029 = ~n1027 & n1028;
  assign n1030 = n1027 & ~n1028;
  assign po92  = ~n1029 & ~n1030;
  assign n1032 = ~pi93  & ~pi221 ;
  assign n1033 = pi93  & pi221 ;
  assign n1034 = ~n1032 & ~n1033;
  assign n1035 = ~n1026 & ~n1030;
  assign n1036 = ~n1034 & n1035;
  assign n1037 = n1034 & ~n1035;
  assign po93  = ~n1036 & ~n1037;
  assign n1039 = ~pi94  & ~pi222 ;
  assign n1040 = pi94  & pi222 ;
  assign n1041 = ~n1039 & ~n1040;
  assign n1042 = ~n1033 & ~n1037;
  assign n1043 = ~n1041 & n1042;
  assign n1044 = n1041 & ~n1042;
  assign po94  = ~n1043 & ~n1044;
  assign n1046 = ~pi95  & ~pi223 ;
  assign n1047 = pi95  & pi223 ;
  assign n1048 = ~n1046 & ~n1047;
  assign n1049 = ~n1040 & ~n1044;
  assign n1050 = ~n1048 & n1049;
  assign n1051 = n1048 & ~n1049;
  assign po95  = ~n1050 & ~n1051;
  assign n1053 = ~pi96  & ~pi224 ;
  assign n1054 = pi96  & pi224 ;
  assign n1055 = ~n1053 & ~n1054;
  assign n1056 = ~n1047 & ~n1051;
  assign n1057 = ~n1055 & n1056;
  assign n1058 = n1055 & ~n1056;
  assign po96  = ~n1057 & ~n1058;
  assign n1060 = ~pi97  & ~pi225 ;
  assign n1061 = pi97  & pi225 ;
  assign n1062 = ~n1060 & ~n1061;
  assign n1063 = ~n1054 & ~n1058;
  assign n1064 = ~n1062 & n1063;
  assign n1065 = n1062 & ~n1063;
  assign po97  = ~n1064 & ~n1065;
  assign n1067 = ~pi98  & ~pi226 ;
  assign n1068 = pi98  & pi226 ;
  assign n1069 = ~n1067 & ~n1068;
  assign n1070 = ~n1061 & ~n1065;
  assign n1071 = ~n1069 & n1070;
  assign n1072 = n1069 & ~n1070;
  assign po98  = ~n1071 & ~n1072;
  assign n1074 = ~pi99  & ~pi227 ;
  assign n1075 = pi99  & pi227 ;
  assign n1076 = ~n1074 & ~n1075;
  assign n1077 = ~n1068 & ~n1072;
  assign n1078 = ~n1076 & n1077;
  assign n1079 = n1076 & ~n1077;
  assign po99  = ~n1078 & ~n1079;
  assign n1081 = ~pi100  & ~pi228 ;
  assign n1082 = pi100  & pi228 ;
  assign n1083 = ~n1081 & ~n1082;
  assign n1084 = ~n1075 & ~n1079;
  assign n1085 = ~n1083 & n1084;
  assign n1086 = n1083 & ~n1084;
  assign po100  = ~n1085 & ~n1086;
  assign n1088 = ~pi101  & ~pi229 ;
  assign n1089 = pi101  & pi229 ;
  assign n1090 = ~n1088 & ~n1089;
  assign n1091 = ~n1082 & ~n1086;
  assign n1092 = ~n1090 & n1091;
  assign n1093 = n1090 & ~n1091;
  assign po101  = ~n1092 & ~n1093;
  assign n1095 = ~pi102  & ~pi230 ;
  assign n1096 = pi102  & pi230 ;
  assign n1097 = ~n1095 & ~n1096;
  assign n1098 = ~n1089 & ~n1093;
  assign n1099 = ~n1097 & n1098;
  assign n1100 = n1097 & ~n1098;
  assign po102  = ~n1099 & ~n1100;
  assign n1102 = ~pi103  & ~pi231 ;
  assign n1103 = pi103  & pi231 ;
  assign n1104 = ~n1102 & ~n1103;
  assign n1105 = ~n1096 & ~n1100;
  assign n1106 = ~n1104 & n1105;
  assign n1107 = n1104 & ~n1105;
  assign po103  = ~n1106 & ~n1107;
  assign n1109 = ~pi104  & ~pi232 ;
  assign n1110 = pi104  & pi232 ;
  assign n1111 = ~n1109 & ~n1110;
  assign n1112 = ~n1103 & ~n1107;
  assign n1113 = ~n1111 & n1112;
  assign n1114 = n1111 & ~n1112;
  assign po104  = ~n1113 & ~n1114;
  assign n1116 = ~pi105  & ~pi233 ;
  assign n1117 = pi105  & pi233 ;
  assign n1118 = ~n1116 & ~n1117;
  assign n1119 = ~n1110 & ~n1114;
  assign n1120 = ~n1118 & n1119;
  assign n1121 = n1118 & ~n1119;
  assign po105  = ~n1120 & ~n1121;
  assign n1123 = ~pi106  & ~pi234 ;
  assign n1124 = pi106  & pi234 ;
  assign n1125 = ~n1123 & ~n1124;
  assign n1126 = ~n1117 & ~n1121;
  assign n1127 = ~n1125 & n1126;
  assign n1128 = n1125 & ~n1126;
  assign po106  = ~n1127 & ~n1128;
  assign n1130 = ~pi107  & ~pi235 ;
  assign n1131 = pi107  & pi235 ;
  assign n1132 = ~n1130 & ~n1131;
  assign n1133 = ~n1124 & ~n1128;
  assign n1134 = ~n1132 & n1133;
  assign n1135 = n1132 & ~n1133;
  assign po107  = ~n1134 & ~n1135;
  assign n1137 = ~pi108  & ~pi236 ;
  assign n1138 = pi108  & pi236 ;
  assign n1139 = ~n1137 & ~n1138;
  assign n1140 = ~n1131 & ~n1135;
  assign n1141 = ~n1139 & n1140;
  assign n1142 = n1139 & ~n1140;
  assign po108  = ~n1141 & ~n1142;
  assign n1144 = ~pi109  & ~pi237 ;
  assign n1145 = pi109  & pi237 ;
  assign n1146 = ~n1144 & ~n1145;
  assign n1147 = ~n1138 & ~n1142;
  assign n1148 = ~n1146 & n1147;
  assign n1149 = n1146 & ~n1147;
  assign po109  = ~n1148 & ~n1149;
  assign n1151 = ~pi110  & ~pi238 ;
  assign n1152 = pi110  & pi238 ;
  assign n1153 = ~n1151 & ~n1152;
  assign n1154 = ~n1145 & ~n1149;
  assign n1155 = ~n1153 & n1154;
  assign n1156 = n1153 & ~n1154;
  assign po110  = ~n1155 & ~n1156;
  assign n1158 = ~pi111  & ~pi239 ;
  assign n1159 = pi111  & pi239 ;
  assign n1160 = ~n1158 & ~n1159;
  assign n1161 = ~n1152 & ~n1156;
  assign n1162 = ~n1160 & n1161;
  assign n1163 = n1160 & ~n1161;
  assign po111  = ~n1162 & ~n1163;
  assign n1165 = ~pi112  & ~pi240 ;
  assign n1166 = pi112  & pi240 ;
  assign n1167 = ~n1165 & ~n1166;
  assign n1168 = ~n1159 & ~n1163;
  assign n1169 = ~n1167 & n1168;
  assign n1170 = n1167 & ~n1168;
  assign po112  = ~n1169 & ~n1170;
  assign n1172 = ~pi113  & ~pi241 ;
  assign n1173 = pi113  & pi241 ;
  assign n1174 = ~n1172 & ~n1173;
  assign n1175 = ~n1166 & ~n1170;
  assign n1176 = ~n1174 & n1175;
  assign n1177 = n1174 & ~n1175;
  assign po113  = ~n1176 & ~n1177;
  assign n1179 = ~pi114  & ~pi242 ;
  assign n1180 = pi114  & pi242 ;
  assign n1181 = ~n1179 & ~n1180;
  assign n1182 = ~n1173 & ~n1177;
  assign n1183 = ~n1181 & n1182;
  assign n1184 = n1181 & ~n1182;
  assign po114  = ~n1183 & ~n1184;
  assign n1186 = ~pi115  & ~pi243 ;
  assign n1187 = pi115  & pi243 ;
  assign n1188 = ~n1186 & ~n1187;
  assign n1189 = ~n1180 & ~n1184;
  assign n1190 = ~n1188 & n1189;
  assign n1191 = n1188 & ~n1189;
  assign po115  = ~n1190 & ~n1191;
  assign n1193 = ~pi116  & ~pi244 ;
  assign n1194 = pi116  & pi244 ;
  assign n1195 = ~n1193 & ~n1194;
  assign n1196 = ~n1187 & ~n1191;
  assign n1197 = ~n1195 & n1196;
  assign n1198 = n1195 & ~n1196;
  assign po116  = ~n1197 & ~n1198;
  assign n1200 = ~pi117  & ~pi245 ;
  assign n1201 = pi117  & pi245 ;
  assign n1202 = ~n1200 & ~n1201;
  assign n1203 = ~n1194 & ~n1198;
  assign n1204 = ~n1202 & n1203;
  assign n1205 = n1202 & ~n1203;
  assign po117  = ~n1204 & ~n1205;
  assign n1207 = ~pi118  & ~pi246 ;
  assign n1208 = pi118  & pi246 ;
  assign n1209 = ~n1207 & ~n1208;
  assign n1210 = ~n1201 & ~n1205;
  assign n1211 = ~n1209 & n1210;
  assign n1212 = n1209 & ~n1210;
  assign po118  = ~n1211 & ~n1212;
  assign n1214 = ~pi119  & ~pi247 ;
  assign n1215 = pi119  & pi247 ;
  assign n1216 = ~n1214 & ~n1215;
  assign n1217 = ~n1208 & ~n1212;
  assign n1218 = ~n1216 & n1217;
  assign n1219 = n1216 & ~n1217;
  assign po119  = ~n1218 & ~n1219;
  assign n1221 = ~pi120  & ~pi248 ;
  assign n1222 = pi120  & pi248 ;
  assign n1223 = ~n1221 & ~n1222;
  assign n1224 = ~n1215 & ~n1219;
  assign n1225 = ~n1223 & n1224;
  assign n1226 = n1223 & ~n1224;
  assign po120  = ~n1225 & ~n1226;
  assign n1228 = ~pi121  & ~pi249 ;
  assign n1229 = pi121  & pi249 ;
  assign n1230 = ~n1228 & ~n1229;
  assign n1231 = ~n1222 & ~n1226;
  assign n1232 = ~n1230 & n1231;
  assign n1233 = n1230 & ~n1231;
  assign po121  = ~n1232 & ~n1233;
  assign n1235 = ~pi122  & ~pi250 ;
  assign n1236 = pi122  & pi250 ;
  assign n1237 = ~n1235 & ~n1236;
  assign n1238 = ~n1229 & ~n1233;
  assign n1239 = ~n1237 & n1238;
  assign n1240 = n1237 & ~n1238;
  assign po122  = ~n1239 & ~n1240;
  assign n1242 = ~pi123  & ~pi251 ;
  assign n1243 = pi123  & pi251 ;
  assign n1244 = ~n1242 & ~n1243;
  assign n1245 = ~n1236 & ~n1240;
  assign n1246 = ~n1244 & n1245;
  assign n1247 = n1244 & ~n1245;
  assign po123  = ~n1246 & ~n1247;
  assign n1249 = ~pi124  & ~pi252 ;
  assign n1250 = pi124  & pi252 ;
  assign n1251 = ~n1249 & ~n1250;
  assign n1252 = ~n1243 & ~n1247;
  assign n1253 = ~n1251 & n1252;
  assign n1254 = n1251 & ~n1252;
  assign po124  = ~n1253 & ~n1254;
  assign n1256 = ~pi125  & ~pi253 ;
  assign n1257 = pi125  & pi253 ;
  assign n1258 = ~n1256 & ~n1257;
  assign n1259 = ~n1250 & ~n1254;
  assign n1260 = ~n1258 & n1259;
  assign n1261 = n1258 & ~n1259;
  assign po125  = ~n1260 & ~n1261;
  assign n1263 = ~pi126  & ~pi254 ;
  assign n1264 = pi126  & pi254 ;
  assign n1265 = ~n1263 & ~n1264;
  assign n1266 = ~n1257 & ~n1261;
  assign n1267 = ~n1265 & n1266;
  assign n1268 = n1265 & ~n1266;
  assign po126  = ~n1267 & ~n1268;
  assign n1270 = ~pi127  & ~pi255 ;
  assign n1271 = pi127  & pi255 ;
  assign n1272 = ~n1270 & ~n1271;
  assign n1273 = ~n1264 & ~n1268;
  assign n1274 = ~n1272 & n1273;
  assign n1275 = n1272 & ~n1273;
  assign po127  = ~n1274 & ~n1275;
  assign po128 = n1271 | n1275;
endmodule
