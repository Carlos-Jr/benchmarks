module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 ,
    pi5 , pi6 , pi7 , pi8 , pi9 ,
    pi10 , pi11 , pi12 , pi13 , pi14 ,
    pi15 , pi16 , pi17 , pi18 , pi19 ,
    pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 ,
    pi30 , pi31 , pi32 , pi33 , pi34 ,
    pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 ,
    pi45 , pi46 , pi47 , pi48 , pi49 ,
    pi50 , pi51 , pi52 , pi53 , pi54 ,
    pi55 , pi56 , pi57 , pi58 , pi59 ,
    po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 ,
    po14 , po15 , po16 , po17 ,
    po18 , po19 , po20 , po21 ,
    po22 , po23 , po24 , po25 ,
    po26 , po27 , po28 , po29   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 ,
    pi5 , pi6 , pi7 , pi8 , pi9 ,
    pi10 , pi11 , pi12 , pi13 , pi14 ,
    pi15 , pi16 , pi17 , pi18 , pi19 ,
    pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 ,
    pi30 , pi31 , pi32 , pi33 , pi34 ,
    pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 ,
    pi45 , pi46 , pi47 , pi48 , pi49 ,
    pi50 , pi51 , pi52 , pi53 , pi54 ,
    pi55 , pi56 , pi57 , pi58 , pi59 ;
  output po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 ,
    po14 , po15 , po16 , po17 ,
    po18 , po19 , po20 , po21 ,
    po22 , po23 , po24 , po25 ,
    po26 , po27 , po28 , po29 ;
  wire n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105,
    n106, n107, n108, n109, n110, n111, n112,
    n113, n114, n115, n116, n117, n118, n119,
    n120, n121, n122, n123, n124, n125, n126,
    n127, n128, n129, n130, n131, n132, n133,
    n134, n135, n136, n137, n138, n139, n140,
    n141, n142, n143, n144, n145, n146, n147,
    n148, n149, n150, n151, n152, n153, n154,
    n155, n156, n157, n158, n159, n160, n161,
    n162, n163, n164, n165, n166, n167, n168,
    n169, n170, n171, n172, n173, n174, n175,
    n176, n177, n179, n180, n181, n182, n183,
    n184, n185, n186, n187, n188, n189, n190,
    n191, n192, n193, n194, n195, n196, n197,
    n198, n199, n200, n201, n202, n203, n204,
    n205, n206, n207, n208, n209, n210, n211,
    n212, n213, n214, n215, n216, n217, n218,
    n219, n220, n221, n222, n223, n224, n225,
    n226, n227, n228, n229, n230, n231, n232,
    n233, n234, n235, n236, n237, n238, n239,
    n240, n241, n242, n243, n244, n245, n246,
    n247, n248, n249, n250, n251, n252, n253,
    n254, n255, n256, n257, n258, n259, n260,
    n261, n262, n263, n264, n265, n266, n267,
    n268, n270, n271, n272;
  assign n92 = pi27  & pi28 ;
  assign n93 = pi29  & n92;
  assign n94 = ~pi9  & ~pi10 ;
  assign n95 = pi11  & ~n94;
  assign n96 = ~pi12  & ~pi13 ;
  assign n97 = ~n95 & n96;
  assign n98 = pi14  & ~n97;
  assign n99 = pi15  & n98;
  assign n100 = ~pi16  & ~n99;
  assign n101 = pi17  & ~n100;
  assign n102 = ~pi18  & ~n101;
  assign n103 = pi19  & ~n102;
  assign n104 = pi20  & n103;
  assign n105 = ~pi21  & ~n104;
  assign n106 = ~pi22  & n105;
  assign n107 = pi24  & pi25 ;
  assign n108 = pi23  & n107;
  assign n109 = ~n106 & n108;
  assign n110 = ~pi26  & ~n109;
  assign n111 = n93 & ~n110;
  assign n112 = pi16  & n99;
  assign n113 = pi21  & n104;
  assign n114 = pi11  & pi12 ;
  assign n115 = ~pi20  & ~n103;
  assign n116 = ~n104 & ~n115;
  assign n117 = pi12  & n94;
  assign n118 = ~n95 & ~n117;
  assign n119 = ~pi15  & ~n98;
  assign n120 = ~n99 & ~n119;
  assign n121 = ~pi1  & ~pi2 ;
  assign n122 = ~pi3  & ~pi4 ;
  assign n123 = ~pi5  & ~pi6 ;
  assign n124 = ~pi7  & ~pi8 ;
  assign n125 = pi9  & ~pi10 ;
  assign n126 = ~pi13  & pi14 ;
  assign n127 = ~pi18  & pi19 ;
  assign n128 = ~pi22  & pi23 ;
  assign n129 = ~pi26  & n128;
  assign n130 = n126 & n127;
  assign n131 = n124 & n125;
  assign n132 = n122 & n123;
  assign n133 = n107 & n121;
  assign n134 = ~n114 & n133;
  assign n135 = n131 & n132;
  assign n136 = n129 & n130;
  assign n137 = n135 & n136;
  assign n138 = ~n118 & n134;
  assign n139 = n137 & n138;
  assign n140 = ~n112 & n139;
  assign n141 = ~n120 & n140;
  assign n142 = n101 & n141;
  assign n143 = ~n105 & n142;
  assign n144 = ~n113 & ~n116;
  assign n145 = n143 & n144;
  assign n146 = n111 & ~n145;
  assign n147 = ~pi19  & n102;
  assign n148 = pi18  & n101;
  assign n149 = ~n102 & ~n148;
  assign n150 = ~pi17  & n100;
  assign n151 = ~pi14  & n97;
  assign n152 = pi0  & pi1 ;
  assign n153 = pi2  & pi3 ;
  assign n154 = pi4  & pi5 ;
  assign n155 = pi6  & pi7 ;
  assign n156 = pi8  & pi11 ;
  assign n157 = pi15  & ~pi16 ;
  assign n158 = pi20  & ~pi21 ;
  assign n159 = n107 & n158;
  assign n160 = n96 & n157;
  assign n161 = n155 & n156;
  assign n162 = n153 & n154;
  assign n163 = n94 & n152;
  assign n164 = n162 & n163;
  assign n165 = n160 & n161;
  assign n166 = n129 & n159;
  assign n167 = n93 & n166;
  assign n168 = n164 & n165;
  assign n169 = n167 & n168;
  assign n170 = ~n98 & ~n151;
  assign n171 = n169 & n170;
  assign n172 = ~n101 & n171;
  assign n173 = ~n150 & n172;
  assign n174 = ~n103 & n173;
  assign n175 = ~n147 & ~n149;
  assign n176 = n174 & n175;
  assign n177 = ~n111 & ~n176;
  assign po0  = n146 | n177;
  assign n179 = pi57  & pi58 ;
  assign n180 = pi54  & pi55 ;
  assign n181 = ~pi39  & ~pi40 ;
  assign n182 = pi41  & ~n181;
  assign n183 = ~pi42  & ~n182;
  assign n184 = ~pi43  & n183;
  assign n185 = pi44  & pi45 ;
  assign n186 = ~n184 & n185;
  assign n187 = ~pi46  & ~n186;
  assign n188 = pi47  & ~n187;
  assign n189 = ~pi48  & ~n188;
  assign n190 = pi49  & pi50 ;
  assign n191 = ~n189 & n190;
  assign n192 = ~pi51  & ~pi52 ;
  assign n193 = ~n191 & n192;
  assign n194 = pi53  & n180;
  assign n195 = ~n193 & n194;
  assign n196 = ~pi56  & ~n195;
  assign n197 = pi59  & n179;
  assign n198 = ~n196 & n197;
  assign n199 = ~pi52  & pi53 ;
  assign n200 = pi47  & pi48 ;
  assign n201 = pi48  & n187;
  assign n202 = ~n188 & ~n201;
  assign n203 = pi42  & n182;
  assign n204 = ~pi31  & ~pi32 ;
  assign n205 = ~pi33  & ~pi34 ;
  assign n206 = ~pi35  & ~pi36 ;
  assign n207 = ~pi37  & ~pi38 ;
  assign n208 = pi39  & ~pi40 ;
  assign n209 = pi41  & ~pi43 ;
  assign n210 = ~pi46  & ~pi51 ;
  assign n211 = ~pi56  & pi57 ;
  assign n212 = n210 & n211;
  assign n213 = n185 & n209;
  assign n214 = n207 & n208;
  assign n215 = n205 & n206;
  assign n216 = n180 & n204;
  assign n217 = n190 & n199;
  assign n218 = ~n200 & n217;
  assign n219 = n215 & n216;
  assign n220 = n213 & n214;
  assign n221 = n212 & n220;
  assign n222 = n218 & n219;
  assign n223 = ~n183 & ~n203;
  assign n224 = n222 & n223;
  assign n225 = n221 & n224;
  assign n226 = ~n202 & n225;
  assign n227 = ~pi0  & ~pi30 ;
  assign n228 = n226 & n227;
  assign n229 = n198 & ~n228;
  assign n230 = ~pi0  & ~pi51 ;
  assign n231 = ~n198 & ~n230;
  assign n232 = pi44  & n184;
  assign n233 = pi43  & ~pi44 ;
  assign n234 = n203 & n233;
  assign n235 = ~n232 & ~n234;
  assign n236 = ~n191 & ~n199;
  assign n237 = ~pi49  & ~n189;
  assign n238 = pi49  & n189;
  assign n239 = ~n237 & ~n238;
  assign n240 = pi52  & ~pi53 ;
  assign n241 = n191 & ~n240;
  assign n242 = pi46  & n186;
  assign n243 = ~pi47  & ~n242;
  assign n244 = pi30  & pi31 ;
  assign n245 = pi32  & pi33 ;
  assign n246 = pi34  & pi35 ;
  assign n247 = pi36  & pi37 ;
  assign n248 = pi38  & pi41 ;
  assign n249 = pi45  & ~pi48 ;
  assign n250 = pi50  & ~pi56 ;
  assign n251 = n248 & n249;
  assign n252 = n246 & n247;
  assign n253 = n244 & n245;
  assign n254 = n180 & n250;
  assign n255 = n181 & n254;
  assign n256 = n252 & n253;
  assign n257 = n197 & n251;
  assign n258 = n256 & n257;
  assign n259 = n255 & n258;
  assign n260 = ~n235 & n259;
  assign n261 = ~n188 & n260;
  assign n262 = ~n243 & n261;
  assign n263 = ~n236 & n262;
  assign n264 = ~n239 & ~n241;
  assign n265 = n263 & n264;
  assign n266 = ~n231 & n265;
  assign n267 = ~n229 & ~n266;
  assign n268 = ~n177 & ~n267;
  assign po1  = ~n146 & ~n268;
  assign n270 = pi0  & pi30 ;
  assign n271 = n226 & ~n270;
  assign n272 = n198 & ~n271;
  assign po2  = ~po0  & n272;
  assign po3  = 1'b0;
  assign po4  = 1'b0;
  assign po5  = 1'b0;
  assign po6  = 1'b0;
  assign po7  = 1'b0;
  assign po8  = 1'b0;
  assign po9  = 1'b0;
  assign po10  = 1'b0;
  assign po11  = 1'b0;
  assign po12  = 1'b0;
  assign po13  = 1'b0;
  assign po14  = 1'b0;
  assign po15  = 1'b0;
  assign po16  = 1'b0;
  assign po17  = 1'b0;
  assign po18  = 1'b0;
  assign po19  = 1'b0;
  assign po20  = 1'b0;
  assign po21  = 1'b0;
  assign po22  = 1'b0;
  assign po23  = 1'b0;
  assign po24  = 1'b0;
  assign po25  = 1'b0;
  assign po26  = 1'b0;
  assign po27  = 1'b0;
  assign po28  = 1'b0;
  assign po29  = 1'b0;
endmodule
