module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 , pi32 ,
    pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 , pi40 ,
    pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 , pi56 ,
    pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 , pi64 ,
    pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 ,
    pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 ,
    pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 ,
    pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 ,
    pi97 , pi98 , pi99 , pi100 , pi101 , pi102 , pi103 ,
    pi104 , pi105 , pi106 , pi107 , pi108 , pi109 , pi110 ,
    pi111 , pi112 , pi113 , pi114 , pi115 , pi116 , pi117 ,
    pi118 , pi119 , pi120 , pi121 , pi122 , pi123 , pi124 ,
    pi125 , pi126 , pi127 ,
    po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7  );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    pi32 , pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 ,
    pi56 , pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 ,
    pi64 , pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 ,
    pi72 , pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 ,
    pi80 , pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 ,
    pi88 , pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 ,
    pi96 , pi97 , pi98 , pi99 , pi100 , pi101 , pi102 ,
    pi103 , pi104 , pi105 , pi106 , pi107 , pi108 , pi109 ,
    pi110 , pi111 , pi112 , pi113 , pi114 , pi115 , pi116 ,
    pi117 , pi118 , pi119 , pi120 , pi121 , pi122 , pi123 ,
    pi124 , pi125 , pi126 , pi127 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7;
  wire n137, n138, n139, n140, n141, n142, n143,
    n144, n145, n146, n147, n148, n149, n150,
    n151, n152, n153, n154, n155, n156, n157,
    n158, n159, n160, n161, n162, n163, n164,
    n165, n166, n167, n168, n169, n170, n171,
    n172, n173, n174, n175, n176, n177, n178,
    n179, n180, n181, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192,
    n193, n194, n195, n196, n197, n198, n199,
    n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213,
    n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227,
    n228, n229, n230, n231, n232, n233, n234,
    n235, n236, n237, n238, n239, n240, n241,
    n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339,
    n340, n341, n342, n343, n344, n345, n346,
    n347, n348, n349, n350, n351, n352, n353,
    n354, n355, n356, n357, n358, n359, n360,
    n361, n362, n363, n364, n365, n366, n367,
    n368, n369, n370, n371, n372, n373, n374,
    n375, n376, n377, n378, n379, n380, n381,
    n382, n383, n384, n385, n386, n387, n388,
    n389, n390, n391, n392, n393, n394, n395,
    n396, n397, n398, n399, n400, n401, n402,
    n403, n404, n405, n406, n407, n408, n409,
    n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423,
    n424, n425, n426, n427, n428, n429, n430,
    n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444,
    n445, n446, n447, n448, n449, n450, n451,
    n452, n453, n454, n455, n456, n457, n458,
    n459, n460, n461, n462, n463, n464, n465,
    n466, n467, n468, n469, n470, n471, n472,
    n473, n474, n475, n476, n477, n478, n479,
    n480, n481, n482, n483, n484, n485, n486,
    n487, n488, n489, n490, n491, n492, n493,
    n494, n495, n496, n497, n498, n499, n500,
    n501, n502, n503, n504, n505, n506, n507,
    n508, n509, n510, n511, n512, n513, n514,
    n515, n516, n517, n518, n519, n520, n521,
    n522, n523, n524, n525, n526, n527, n528,
    n529, n530, n531, n532, n533, n534, n535,
    n536, n537, n538, n539, n540, n541, n542,
    n543, n544, n545, n546, n547, n548, n549,
    n550, n551, n552, n553, n554, n555, n556,
    n557, n558, n559, n560, n561, n562, n563,
    n564, n565, n566, n567, n568, n569, n570,
    n571, n572, n573, n574, n575, n576, n577,
    n578, n579, n580, n581, n582, n583, n584,
    n585, n586, n587, n588, n589, n590, n591,
    n592, n593, n594, n595, n596, n597, n598,
    n599, n600, n601, n602, n603, n604, n605,
    n606, n607, n608, n609, n610, n611, n612,
    n613, n614, n615, n616, n617, n618, n619,
    n620, n621, n622, n623, n624, n625, n626,
    n627, n628, n629, n630, n631, n632, n633,
    n634, n635, n636, n637, n638, n639, n640,
    n641, n642, n643, n644, n645, n646, n647,
    n648, n649, n650, n651, n652, n653, n654,
    n655, n656, n657, n658, n659, n660, n661,
    n662, n663, n664, n665, n666, n667, n668,
    n669, n670, n671, n672, n673, n674, n675,
    n676, n677, n678, n679, n680, n681, n682,
    n683, n684, n685, n686, n687, n688, n689,
    n690, n691, n692, n693, n694, n695, n696,
    n697, n698, n699, n700, n701, n702, n703,
    n704, n705, n706, n707, n708, n709, n710,
    n711, n712, n713, n714, n715, n716, n717,
    n718, n719, n720, n721, n722, n723, n724,
    n725, n726, n727, n728, n729, n730, n731,
    n732, n733, n734, n735, n736, n737, n738,
    n739, n740, n741, n742, n743, n744, n745,
    n746, n747, n748, n749, n750, n751, n752,
    n753, n754, n755, n756, n757, n758, n759,
    n760, n761, n762, n763, n764, n765, n766,
    n767, n768, n769, n770, n771, n772, n773,
    n774, n775, n776, n777, n778, n779, n780,
    n781, n782, n783, n784, n785, n786, n787,
    n788, n789, n790, n791, n792, n793, n794,
    n795, n796, n797, n798, n799, n800, n801,
    n802, n803, n804, n805, n806, n807, n808,
    n809, n810, n811, n812, n813, n814, n815,
    n816, n817, n818, n819, n820, n821, n822,
    n823, n824, n825, n826, n827, n828, n829,
    n830, n831, n832, n833, n834, n835, n836,
    n837, n838, n839, n840, n841, n842, n843,
    n844, n845, n846, n847, n848, n849, n850,
    n851, n852, n853, n854, n855, n856, n857,
    n858, n859, n860, n861, n862, n863, n864,
    n865, n866, n867, n868, n869, n870, n871,
    n872, n873, n874, n875, n876, n877, n878,
    n879, n880, n881, n882, n883, n884, n885,
    n886, n887, n888, n889, n890, n891, n892,
    n893, n894, n895, n896, n897, n898, n899,
    n900, n901, n902, n903, n904, n905, n906,
    n907, n908, n909, n910, n911, n912, n913,
    n914, n915, n916, n917, n918, n919, n920,
    n921, n922, n923, n924, n925, n926, n927,
    n928, n929, n930, n931, n932, n933, n934,
    n935, n936, n937, n938, n939, n940, n941,
    n942, n943, n944, n945, n946, n947, n948,
    n949, n950, n951, n952, n953, n954, n955,
    n956, n957, n958, n959, n960, n961, n962,
    n963, n964, n965, n966, n967, n968, n969,
    n970, n971, n972, n973, n974, n975, n976,
    n977, n978, n979, n980, n981, n982, n983,
    n984, n985, n986, n987, n988, n989, n990,
    n991, n992, n993, n994, n995, n996, n997,
    n998, n999, n1000, n1001, n1002, n1003,
    n1004, n1005, n1006, n1007, n1008, n1009,
    n1010, n1011, n1012, n1013, n1014, n1015,
    n1016, n1017, n1018, n1019, n1020, n1021,
    n1022, n1023, n1024, n1025, n1026, n1027,
    n1028, n1029, n1030, n1031, n1032, n1033,
    n1034, n1035, n1036, n1037, n1038, n1039,
    n1040, n1041, n1042, n1043, n1044, n1045,
    n1046, n1047, n1048, n1049, n1050, n1051,
    n1052, n1053, n1054, n1055, n1056, n1057,
    n1058, n1059, n1060, n1061, n1062, n1063,
    n1064, n1065, n1066, n1067, n1068, n1069,
    n1070, n1071, n1072, n1073, n1074, n1075,
    n1076, n1077, n1078, n1079, n1080, n1081,
    n1082, n1083, n1084, n1085, n1086, n1087,
    n1088, n1089, n1090, n1091, n1092, n1093,
    n1094, n1095, n1096, n1097, n1098, n1099,
    n1100, n1101, n1102, n1103, n1104, n1105,
    n1106, n1107, n1108, n1109, n1110, n1111,
    n1112, n1113, n1114, n1115, n1116, n1117,
    n1118, n1119, n1120, n1121, n1122, n1123,
    n1124, n1125, n1126, n1127, n1128, n1129,
    n1130, n1131, n1132, n1133, n1134, n1135,
    n1136, n1137, n1138, n1139, n1140, n1141,
    n1142, n1143, n1144, n1145, n1146, n1147,
    n1148, n1149, n1150, n1151, n1152, n1153,
    n1154, n1155, n1156, n1157, n1158, n1159,
    n1160, n1161, n1162, n1163, n1164, n1165,
    n1166, n1167, n1168, n1169, n1170, n1171,
    n1172, n1173, n1174, n1175, n1176, n1177,
    n1178, n1179, n1180, n1181, n1182, n1183,
    n1184, n1185, n1186, n1187, n1188, n1189,
    n1190, n1191, n1192, n1193, n1194, n1195,
    n1196, n1197, n1198, n1199, n1200, n1201,
    n1202, n1203, n1204, n1205, n1206, n1207,
    n1208, n1209, n1210, n1211, n1212, n1213,
    n1214, n1215, n1216, n1217, n1218, n1219,
    n1220, n1221, n1222, n1223, n1224, n1225,
    n1226, n1227, n1228, n1229, n1230, n1231,
    n1232, n1233, n1234, n1235, n1236, n1237,
    n1238, n1239, n1240, n1241, n1242, n1243,
    n1244, n1245, n1246, n1247, n1248, n1249,
    n1250, n1251, n1252, n1253, n1254, n1255,
    n1256, n1257, n1258, n1259, n1260, n1261,
    n1262, n1263, n1264, n1265, n1266, n1267,
    n1268, n1269, n1270, n1271, n1272, n1273,
    n1274, n1275, n1276, n1277, n1278, n1279,
    n1280, n1281, n1282, n1283, n1284, n1285,
    n1286, n1287, n1288, n1289, n1290, n1291,
    n1292, n1293, n1294, n1295, n1296, n1297,
    n1298, n1299, n1300, n1301, n1302, n1303,
    n1304, n1305, n1306, n1307, n1308, n1309,
    n1310, n1311, n1312, n1313, n1314, n1315,
    n1316, n1317, n1318, n1319, n1320, n1321,
    n1322, n1323, n1324, n1325, n1326, n1327,
    n1328, n1329, n1330, n1331, n1332, n1333,
    n1334, n1335, n1336, n1337, n1338, n1339,
    n1340, n1341, n1342, n1343, n1344, n1345,
    n1346, n1347, n1348, n1349, n1350, n1351,
    n1352, n1353, n1354, n1355, n1356, n1357,
    n1358, n1359, n1360, n1361, n1362, n1363,
    n1364, n1365, n1366, n1367, n1368, n1369,
    n1370, n1371, n1372, n1373, n1374, n1375,
    n1376, n1377, n1378, n1379, n1380, n1381,
    n1382, n1383, n1384, n1385, n1386, n1387,
    n1388, n1389, n1390, n1391, n1392, n1393,
    n1394, n1395, n1396, n1397, n1398, n1399,
    n1400, n1401, n1402, n1403, n1404, n1405,
    n1406, n1407, n1408, n1409, n1410, n1411,
    n1412, n1413, n1414, n1415, n1416, n1417,
    n1418, n1419, n1420, n1421, n1422, n1423,
    n1424, n1425, n1426, n1427, n1428, n1429,
    n1430, n1431, n1432, n1433, n1434, n1435,
    n1436, n1437, n1438, n1439, n1440, n1441,
    n1442, n1443, n1444, n1445, n1446, n1447,
    n1448, n1449, n1450, n1451, n1452, n1453,
    n1454, n1455, n1456, n1457, n1458, n1459,
    n1460, n1461, n1462, n1463, n1464, n1465,
    n1466, n1467, n1468, n1469, n1470, n1471,
    n1472, n1473, n1474, n1475, n1476, n1477,
    n1478, n1479, n1480, n1481, n1482, n1483,
    n1484, n1485, n1486, n1487, n1488, n1489,
    n1490, n1491, n1492, n1493, n1494, n1495,
    n1496, n1497, n1498, n1499, n1500, n1501,
    n1502, n1503, n1504, n1505, n1506, n1507,
    n1508, n1509, n1510, n1511, n1512, n1513,
    n1514, n1515, n1516, n1517, n1518, n1519,
    n1520, n1521, n1522, n1523, n1524, n1525,
    n1526, n1527, n1528, n1529, n1530, n1531,
    n1532, n1533, n1534, n1535, n1536, n1537,
    n1538, n1539, n1540, n1541, n1542, n1543,
    n1544, n1545, n1546, n1547, n1548, n1549,
    n1550, n1551, n1552, n1553, n1554, n1555,
    n1556, n1557, n1558, n1559, n1560, n1561,
    n1562, n1563, n1564, n1565, n1566, n1567,
    n1568, n1569, n1570, n1571, n1572, n1573,
    n1574, n1575, n1576, n1577, n1578, n1579,
    n1580, n1581, n1582, n1583, n1584, n1585,
    n1586, n1587, n1588, n1589, n1590, n1591,
    n1592, n1593, n1594, n1595, n1596, n1597,
    n1598, n1599, n1600, n1601, n1602, n1603,
    n1604, n1605, n1606, n1607, n1608, n1609,
    n1610, n1611, n1612, n1613, n1614, n1615,
    n1616, n1617, n1618, n1619, n1620, n1621,
    n1622, n1623, n1624, n1625, n1626, n1627,
    n1628, n1629, n1630, n1631, n1632, n1633,
    n1634, n1635, n1636, n1637, n1638, n1639,
    n1640, n1641, n1642, n1643, n1644, n1645,
    n1646, n1647, n1648, n1649, n1650, n1651,
    n1652, n1653, n1654, n1655, n1656, n1657,
    n1658, n1659, n1660, n1661, n1662, n1663,
    n1664, n1665, n1666, n1667, n1668, n1669,
    n1670, n1671, n1672, n1673, n1674, n1675,
    n1676, n1677, n1678, n1679, n1680, n1681,
    n1682, n1683, n1684, n1685, n1686, n1687,
    n1688, n1689, n1690, n1691, n1692, n1693,
    n1694, n1695, n1696, n1697, n1698, n1699,
    n1700, n1701, n1702, n1703, n1704, n1705,
    n1706, n1707, n1708, n1709, n1710, n1711,
    n1712, n1713, n1714, n1715, n1716, n1717,
    n1718, n1719, n1720, n1721, n1722, n1723,
    n1724, n1725, n1726, n1727, n1728, n1729,
    n1730, n1731, n1732, n1733, n1734, n1735,
    n1736, n1737, n1738, n1739, n1740, n1741,
    n1742, n1743, n1744, n1745, n1746, n1747,
    n1748, n1749, n1750, n1751, n1752, n1753,
    n1754, n1755, n1756, n1757, n1758, n1759,
    n1760, n1761, n1762, n1763, n1764, n1765,
    n1766, n1767, n1768, n1769, n1770, n1772,
    n1773, n1774, n1775, n1776, n1777, n1778,
    n1779, n1780, n1781, n1782, n1783, n1784,
    n1785, n1786, n1787, n1788, n1789, n1790,
    n1791, n1792, n1793, n1794, n1795, n1796,
    n1797, n1798, n1799, n1800, n1801, n1803,
    n1804, n1805, n1806, n1808, n1809, n1811,
    n1812, n1813, n1814, n1815, n1816, n1817;
  assign n137 = ~pi118  & ~pi119 ;
  assign n138 = ~pi116  & ~pi117 ;
  assign n139 = ~pi117  & n137;
  assign n140 = ~pi116  & n139;
  assign n141 = n137 & n138;
  assign n142 = ~pi114  & ~pi115 ;
  assign n143 = ~pi112  & ~pi113 ;
  assign n144 = n142 & n143;
  assign n145 = ~pi113  & n142;
  assign n146 = ~pi112  & n1714;
  assign n147 = n145 & n146;
  assign n148 = ~pi113  & ~pi114 ;
  assign n149 = ~pi112  & n148;
  assign n150 = ~pi114  & n143;
  assign n151 = ~pi115  & n1714;
  assign n152 = n1716 & n151;
  assign n153 = n1714 & n144;
  assign n154 = ~pi126  & pi127 ;
  assign n155 = ~pi126  & ~n154;
  assign n156 = ~pi126  & ~pi127 ;
  assign n157 = ~pi124  & ~pi125 ;
  assign n158 = n1717 & n157;
  assign n159 = ~pi122  & ~pi123 ;
  assign n160 = ~pi120  & ~pi121 ;
  assign n161 = n159 & n160;
  assign n162 = n158 & n161;
  assign n163 = n1715 & n162;
  assign n164 = ~pi108  & ~pi109 ;
  assign n165 = ~pi110  & ~pi111 ;
  assign n166 = ~pi109  & n165;
  assign n167 = ~pi108  & n166;
  assign n168 = n164 & n165;
  assign n169 = ~pi106  & ~pi107 ;
  assign n170 = ~pi104  & ~pi105 ;
  assign n171 = ~pi105  & n169;
  assign n172 = ~pi104  & n171;
  assign n173 = n169 & n170;
  assign n174 = ~pi107  & n1718;
  assign n175 = ~pi106  & n174;
  assign n176 = ~pi105  & n175;
  assign n177 = ~pi104  & n176;
  assign n178 = n1718 & n1719;
  assign n179 = ~pi102  & ~pi103 ;
  assign n180 = ~pi100  & ~pi101 ;
  assign n181 = ~pi101  & n179;
  assign n182 = ~pi100  & n181;
  assign n183 = n179 & n180;
  assign n184 = ~pi98  & ~pi99 ;
  assign n185 = ~pi96  & ~pi97 ;
  assign n186 = ~pi97  & n184;
  assign n187 = ~pi96  & n186;
  assign n188 = n184 & n185;
  assign n189 = n1721 & n1722;
  assign n190 = ~pi99  & n1721;
  assign n191 = ~pi98  & n1720;
  assign n192 = ~pi97  & n191;
  assign n193 = ~pi96  & n192;
  assign n194 = n190 & n193;
  assign n195 = ~pi101  & ~pi102 ;
  assign n196 = ~pi100  & n195;
  assign n197 = ~pi102  & n180;
  assign n198 = ~pi99  & n1724;
  assign n199 = ~pi98  & n198;
  assign n200 = ~pi97  & n199;
  assign n201 = ~pi96  & n200;
  assign n202 = n1722 & n1724;
  assign n203 = ~pi103  & n1720;
  assign n204 = n1725 & n203;
  assign n205 = n1720 & n189;
  assign n206 = n163 & n1723;
  assign n207 = ~pi94  & ~pi95 ;
  assign n208 = ~pi92  & ~pi93 ;
  assign n209 = ~pi93  & n207;
  assign n210 = ~pi92  & n209;
  assign n211 = n207 & n208;
  assign n212 = ~pi88  & ~pi89 ;
  assign n213 = ~pi90  & ~pi91 ;
  assign n214 = ~pi89  & n213;
  assign n215 = ~pi88  & n214;
  assign n216 = n212 & n213;
  assign n217 = ~pi91  & n1726;
  assign n218 = ~pi90  & n217;
  assign n219 = ~pi89  & n218;
  assign n220 = ~pi88  & n219;
  assign n221 = n1726 & n1727;
  assign n222 = ~pi84  & ~pi85 ;
  assign n223 = ~pi86  & ~pi87 ;
  assign n224 = ~pi85  & n223;
  assign n225 = ~pi84  & n224;
  assign n226 = n222 & n223;
  assign n227 = ~pi80  & ~pi81 ;
  assign n228 = ~pi82  & ~pi83 ;
  assign n229 = ~pi81  & n228;
  assign n230 = ~pi80  & n229;
  assign n231 = n227 & n228;
  assign n232 = ~pi83  & n1729;
  assign n233 = ~pi82  & n232;
  assign n234 = ~pi81  & n233;
  assign n235 = ~pi80  & n234;
  assign n236 = n1729 & n1730;
  assign n237 = ~pi87  & n1728;
  assign n238 = ~pi86  & n237;
  assign n239 = ~pi85  & n238;
  assign n240 = ~pi84  & n239;
  assign n241 = ~pi83  & n240;
  assign n242 = ~pi82  & n241;
  assign n243 = ~pi81  & n242;
  assign n244 = ~pi80  & n243;
  assign n245 = n1728 & n1731;
  assign n246 = ~pi76  & ~pi77 ;
  assign n247 = ~pi78  & ~pi79 ;
  assign n248 = ~pi77  & n247;
  assign n249 = ~pi76  & n248;
  assign n250 = n246 & n247;
  assign n251 = ~pi72  & ~pi73 ;
  assign n252 = ~pi74  & ~pi75 ;
  assign n253 = ~pi73  & n252;
  assign n254 = ~pi72  & n253;
  assign n255 = n251 & n252;
  assign n256 = ~pi75  & n1733;
  assign n257 = ~pi74  & n256;
  assign n258 = ~pi73  & n257;
  assign n259 = ~pi72  & n258;
  assign n260 = n1733 & n1734;
  assign n261 = ~pi68  & ~pi69 ;
  assign n262 = ~pi70  & ~pi71 ;
  assign n263 = ~pi69  & n262;
  assign n264 = ~pi68  & n263;
  assign n265 = n261 & n262;
  assign n266 = ~pi64  & ~pi65 ;
  assign n267 = ~pi66  & ~pi67 ;
  assign n268 = ~pi65  & n267;
  assign n269 = ~pi64  & n268;
  assign n270 = n266 & n267;
  assign n271 = ~pi67  & n1736;
  assign n272 = ~pi66  & n271;
  assign n273 = ~pi65  & n272;
  assign n274 = ~pi64  & n273;
  assign n275 = n1736 & n1737;
  assign n276 = n1735 & n1738;
  assign n277 = ~pi71  & n1735;
  assign n278 = ~pi70  & n1732;
  assign n279 = ~pi69  & n278;
  assign n280 = ~pi68  & n279;
  assign n281 = ~pi67  & n280;
  assign n282 = ~pi66  & n281;
  assign n283 = ~pi65  & n282;
  assign n284 = ~pi64  & n283;
  assign n285 = n277 & n284;
  assign n286 = n1732 & n276;
  assign n287 = n206 & n1739;
  assign n288 = ~pi60  & ~pi61 ;
  assign n289 = ~pi62  & ~pi63 ;
  assign n290 = ~pi61  & n289;
  assign n291 = ~pi60  & n290;
  assign n292 = n288 & n289;
  assign n293 = ~pi56  & ~pi57 ;
  assign n294 = ~pi58  & ~pi59 ;
  assign n295 = ~pi57  & n294;
  assign n296 = ~pi56  & n295;
  assign n297 = n293 & n294;
  assign n298 = ~pi59  & n1740;
  assign n299 = ~pi58  & n298;
  assign n300 = ~pi57  & n299;
  assign n301 = ~pi56  & n300;
  assign n302 = n1740 & n1741;
  assign n303 = ~pi52  & ~pi53 ;
  assign n304 = ~pi54  & ~pi55 ;
  assign n305 = ~pi53  & n304;
  assign n306 = ~pi52  & n305;
  assign n307 = n303 & n304;
  assign n308 = ~pi48  & ~pi49 ;
  assign n309 = ~pi50  & ~pi51 ;
  assign n310 = ~pi49  & n309;
  assign n311 = ~pi48  & n310;
  assign n312 = n308 & n309;
  assign n313 = ~pi51  & n1743;
  assign n314 = ~pi50  & n313;
  assign n315 = ~pi49  & n314;
  assign n316 = ~pi48  & n315;
  assign n317 = n1743 & n1744;
  assign n318 = ~pi55  & n1742;
  assign n319 = ~pi54  & n318;
  assign n320 = ~pi53  & n319;
  assign n321 = ~pi52  & n320;
  assign n322 = ~pi51  & n321;
  assign n323 = ~pi50  & n322;
  assign n324 = ~pi49  & n323;
  assign n325 = ~pi48  & n324;
  assign n326 = n1742 & n1745;
  assign n327 = ~pi44  & ~pi45 ;
  assign n328 = ~pi46  & ~pi47 ;
  assign n329 = ~pi45  & n328;
  assign n330 = ~pi44  & n329;
  assign n331 = n327 & n328;
  assign n332 = ~pi40  & ~pi41 ;
  assign n333 = ~pi42  & ~pi43 ;
  assign n334 = ~pi41  & n333;
  assign n335 = ~pi40  & n334;
  assign n336 = n332 & n333;
  assign n337 = ~pi43  & n1747;
  assign n338 = ~pi42  & n337;
  assign n339 = ~pi41  & n338;
  assign n340 = ~pi40  & n339;
  assign n341 = n1747 & n1748;
  assign n342 = ~pi38  & ~pi39 ;
  assign n343 = ~pi36  & ~pi37 ;
  assign n344 = ~pi37  & n342;
  assign n345 = ~pi36  & n344;
  assign n346 = n342 & n343;
  assign n347 = ~pi34  & ~pi35 ;
  assign n348 = ~pi32  & ~pi33 ;
  assign n349 = ~pi33  & n347;
  assign n350 = ~pi32  & n349;
  assign n351 = n347 & n348;
  assign n352 = ~pi35  & n1750;
  assign n353 = ~pi34  & n352;
  assign n354 = ~pi33  & n353;
  assign n355 = ~pi32  & n354;
  assign n356 = n1750 & n1751;
  assign n357 = ~pi39  & n1749;
  assign n358 = ~pi38  & n357;
  assign n359 = ~pi37  & n358;
  assign n360 = ~pi36  & n359;
  assign n361 = ~pi35  & n360;
  assign n362 = ~pi34  & n361;
  assign n363 = ~pi33  & n362;
  assign n364 = ~pi32  & n363;
  assign n365 = n1749 & n1752;
  assign n366 = ~pi47  & n1746;
  assign n367 = ~pi46  & n366;
  assign n368 = ~pi45  & n367;
  assign n369 = ~pi44  & n368;
  assign n370 = ~pi43  & n369;
  assign n371 = ~pi42  & n370;
  assign n372 = ~pi41  & n371;
  assign n373 = ~pi40  & n372;
  assign n374 = ~pi39  & n373;
  assign n375 = ~pi38  & n374;
  assign n376 = ~pi37  & n375;
  assign n377 = ~pi36  & n376;
  assign n378 = ~pi35  & n377;
  assign n379 = ~pi34  & n378;
  assign n380 = ~pi33  & n379;
  assign n381 = ~pi32  & n380;
  assign n382 = n1746 & n1753;
  assign n383 = ~pi30  & ~pi31 ;
  assign n384 = ~pi28  & ~pi29 ;
  assign n385 = ~pi29  & n383;
  assign n386 = ~pi28  & n385;
  assign n387 = n383 & n384;
  assign n388 = ~pi26  & ~pi27 ;
  assign n389 = ~pi24  & ~pi25 ;
  assign n390 = ~pi25  & n388;
  assign n391 = ~pi24  & n390;
  assign n392 = n388 & n389;
  assign n393 = ~pi27  & n1755;
  assign n394 = ~pi26  & n393;
  assign n395 = ~pi25  & n394;
  assign n396 = ~pi24  & n395;
  assign n397 = n1755 & n1756;
  assign n398 = ~pi22  & ~pi23 ;
  assign n399 = ~pi20  & ~pi21 ;
  assign n400 = ~pi21  & n398;
  assign n401 = ~pi20  & n400;
  assign n402 = n398 & n399;
  assign n403 = ~pi18  & ~pi19 ;
  assign n404 = ~pi16  & ~pi17 ;
  assign n405 = ~pi17  & n403;
  assign n406 = ~pi16  & n405;
  assign n407 = n403 & n404;
  assign n408 = ~pi19  & n1758;
  assign n409 = ~pi18  & n408;
  assign n410 = ~pi17  & n409;
  assign n411 = ~pi16  & n410;
  assign n412 = n1758 & n1759;
  assign n413 = ~pi23  & n1757;
  assign n414 = ~pi22  & n413;
  assign n415 = ~pi21  & n414;
  assign n416 = ~pi20  & n415;
  assign n417 = ~pi19  & n416;
  assign n418 = ~pi18  & n417;
  assign n419 = ~pi17  & n418;
  assign n420 = ~pi16  & n419;
  assign n421 = n1757 & n1760;
  assign n422 = ~pi14  & ~pi15 ;
  assign n423 = ~pi12  & ~pi13 ;
  assign n424 = ~pi13  & n422;
  assign n425 = ~pi12  & n424;
  assign n426 = n422 & n423;
  assign n427 = ~pi10  & ~pi11 ;
  assign n428 = ~pi8  & ~pi9 ;
  assign n429 = ~pi9  & n427;
  assign n430 = ~pi8  & n429;
  assign n431 = n427 & n428;
  assign n432 = ~pi11  & n1762;
  assign n433 = ~pi10  & n432;
  assign n434 = ~pi9  & n433;
  assign n435 = ~pi8  & n434;
  assign n436 = n1762 & n1763;
  assign n437 = ~pi6  & ~pi7 ;
  assign n438 = ~pi4  & ~pi5 ;
  assign n439 = ~pi5  & n437;
  assign n440 = ~pi4  & n439;
  assign n441 = n437 & n438;
  assign n442 = ~pi2  & ~pi3 ;
  assign n443 = ~pi0  & ~pi1 ;
  assign n444 = n442 & n443;
  assign n445 = n1765 & n444;
  assign n446 = n1764 & n445;
  assign n447 = n1761 & n446;
  assign n448 = n1754 & n447;
  assign n449 = ~pi0  & n287;
  assign n450 = n1764 & n449;
  assign n451 = ~pi3  & n450;
  assign n452 = ~pi2  & n451;
  assign n453 = n1754 & n1761;
  assign n454 = n1765 & n453;
  assign n455 = ~pi1  & n454;
  assign n456 = n452 & n455;
  assign n457 = n287 & n448;
  assign n458 = pi118  & ~pi119 ;
  assign n459 = ~pi120  & ~n458;
  assign n460 = ~pi121  & ~n459;
  assign n461 = ~pi122  & ~n460;
  assign n462 = ~pi123  & ~n461;
  assign n463 = ~pi124  & ~n462;
  assign n464 = ~pi125  & ~n463;
  assign n465 = ~pi126  & ~n464;
  assign n466 = pi117  & n465;
  assign n467 = pi119  & ~pi120 ;
  assign n468 = ~pi121  & ~n467;
  assign n469 = ~pi122  & ~n468;
  assign n470 = ~pi123  & ~n469;
  assign n471 = ~pi124  & ~n470;
  assign n472 = ~pi125  & ~n471;
  assign n473 = ~pi117  & ~pi126 ;
  assign n474 = ~n472 & n473;
  assign n475 = ~pi127  & ~n474;
  assign n476 = pi124  & ~pi125 ;
  assign n477 = ~pi126  & ~n476;
  assign n478 = pi123  & n477;
  assign n479 = ~pi123  & pi125 ;
  assign n480 = ~pi126  & n479;
  assign n481 = ~pi127  & ~n480;
  assign n482 = ~pi125  & pi127 ;
  assign n483 = pi126  & pi127 ;
  assign n484 = pi126  & ~n483;
  assign n485 = pi125  & ~n484;
  assign n486 = ~n482 & ~n485;
  assign n487 = ~pi123  & ~n486;
  assign n488 = ~pi124  & ~n484;
  assign n489 = pi124  & ~n486;
  assign n490 = ~n488 & ~n489;
  assign n491 = ~pi127  & ~n477;
  assign n492 = pi123  & ~n1767;
  assign n493 = ~n487 & ~n492;
  assign n494 = ~n478 & n481;
  assign n495 = ~pi121  & ~n1768;
  assign n496 = ~pi122  & ~n1767;
  assign n497 = pi122  & ~n1768;
  assign n498 = ~n496 & ~n497;
  assign n499 = pi121  & ~n498;
  assign n500 = ~n495 & ~n499;
  assign n501 = ~pi119  & ~n500;
  assign n502 = ~pi120  & ~n498;
  assign n503 = pi120  & ~n500;
  assign n504 = ~n502 & ~n503;
  assign n505 = pi119  & ~n504;
  assign n506 = ~n501 & ~n505;
  assign n507 = ~pi117  & ~n506;
  assign n508 = ~pi118  & ~n504;
  assign n509 = pi118  & ~n506;
  assign n510 = ~n508 & ~n509;
  assign n511 = ~pi127  & ~n465;
  assign n512 = pi117  & ~n1769;
  assign n513 = ~n507 & ~n512;
  assign n514 = ~n466 & n475;
  assign n515 = ~pi115  & ~n1770;
  assign n516 = ~pi116  & ~n1769;
  assign n517 = pi116  & ~n1770;
  assign n518 = ~n516 & ~n517;
  assign n519 = pi115  & ~n518;
  assign n520 = ~n515 & ~n519;
  assign n521 = ~pi113  & ~n520;
  assign n522 = ~pi114  & ~n518;
  assign n523 = pi114  & ~n520;
  assign n524 = ~n522 & ~n523;
  assign n525 = pi113  & ~n524;
  assign n526 = ~n521 & ~n525;
  assign n527 = ~pi111  & ~n526;
  assign n528 = ~pi112  & ~n524;
  assign n529 = pi112  & ~n526;
  assign n530 = ~n528 & ~n529;
  assign n531 = pi111  & ~n530;
  assign n532 = ~n527 & ~n531;
  assign n533 = ~pi109  & ~n532;
  assign n534 = ~pi110  & ~n530;
  assign n535 = pi110  & ~n532;
  assign n536 = ~n534 & ~n535;
  assign n537 = pi109  & ~n536;
  assign n538 = ~n533 & ~n537;
  assign n539 = ~pi107  & ~n538;
  assign n540 = ~pi108  & ~n536;
  assign n541 = pi108  & ~n538;
  assign n542 = ~n540 & ~n541;
  assign n543 = pi107  & ~n542;
  assign n544 = ~n539 & ~n543;
  assign n545 = ~pi105  & ~n544;
  assign n546 = ~pi106  & ~n542;
  assign n547 = pi106  & ~n544;
  assign n548 = ~n546 & ~n547;
  assign n549 = pi105  & ~n548;
  assign n550 = ~n545 & ~n549;
  assign n551 = ~pi103  & ~n550;
  assign n552 = ~pi104  & ~n548;
  assign n553 = pi104  & ~n550;
  assign n554 = ~n552 & ~n553;
  assign n555 = pi103  & ~n554;
  assign n556 = ~n551 & ~n555;
  assign n557 = ~pi101  & ~n556;
  assign n558 = ~pi102  & ~n554;
  assign n559 = pi102  & ~n556;
  assign n560 = ~n558 & ~n559;
  assign n561 = pi101  & ~n560;
  assign n562 = ~n557 & ~n561;
  assign n563 = ~pi99  & ~n562;
  assign n564 = ~pi100  & ~n560;
  assign n565 = pi100  & ~n562;
  assign n566 = ~n564 & ~n565;
  assign n567 = pi99  & ~n566;
  assign n568 = ~n563 & ~n567;
  assign n569 = ~pi97  & ~n568;
  assign n570 = ~pi98  & ~n566;
  assign n571 = pi98  & ~n568;
  assign n572 = ~n570 & ~n571;
  assign n573 = pi97  & ~n572;
  assign n574 = ~n569 & ~n573;
  assign n575 = ~pi95  & ~n574;
  assign n576 = ~pi96  & ~n572;
  assign n577 = pi96  & ~n574;
  assign n578 = ~n576 & ~n577;
  assign n579 = pi95  & ~n578;
  assign n580 = ~n575 & ~n579;
  assign n581 = ~pi93  & ~n580;
  assign n582 = ~pi94  & ~n578;
  assign n583 = pi94  & ~n580;
  assign n584 = ~n582 & ~n583;
  assign n585 = pi93  & ~n584;
  assign n586 = ~n581 & ~n585;
  assign n587 = ~pi91  & ~n586;
  assign n588 = ~pi92  & ~n584;
  assign n589 = pi92  & ~n586;
  assign n590 = ~n588 & ~n589;
  assign n591 = pi91  & ~n590;
  assign n592 = ~n587 & ~n591;
  assign n593 = ~pi89  & ~n592;
  assign n594 = ~pi90  & ~n590;
  assign n595 = pi90  & ~n592;
  assign n596 = ~n594 & ~n595;
  assign n597 = pi89  & ~n596;
  assign n598 = ~n593 & ~n597;
  assign n599 = ~pi87  & ~n598;
  assign n600 = ~pi88  & ~n596;
  assign n601 = pi88  & ~n598;
  assign n602 = ~n600 & ~n601;
  assign n603 = pi87  & ~n602;
  assign n604 = ~n599 & ~n603;
  assign n605 = ~pi85  & ~n604;
  assign n606 = ~pi86  & ~n602;
  assign n607 = pi86  & ~n604;
  assign n608 = ~n606 & ~n607;
  assign n609 = pi85  & ~n608;
  assign n610 = ~n605 & ~n609;
  assign n611 = ~pi83  & ~n610;
  assign n612 = ~pi84  & ~n608;
  assign n613 = pi84  & ~n610;
  assign n614 = ~n612 & ~n613;
  assign n615 = pi83  & ~n614;
  assign n616 = ~n611 & ~n615;
  assign n617 = ~pi81  & ~n616;
  assign n618 = ~pi82  & ~n614;
  assign n619 = pi82  & ~n616;
  assign n620 = ~n618 & ~n619;
  assign n621 = pi81  & ~n620;
  assign n622 = ~n617 & ~n621;
  assign n623 = ~pi79  & ~n622;
  assign n624 = ~pi80  & ~n620;
  assign n625 = pi80  & ~n622;
  assign n626 = ~n624 & ~n625;
  assign n627 = pi79  & ~n626;
  assign n628 = ~n623 & ~n627;
  assign n629 = ~pi77  & ~n628;
  assign n630 = ~pi78  & ~n626;
  assign n631 = pi78  & ~n628;
  assign n632 = ~n630 & ~n631;
  assign n633 = pi77  & ~n632;
  assign n634 = ~n629 & ~n633;
  assign n635 = ~pi75  & ~n634;
  assign n636 = ~pi76  & ~n632;
  assign n637 = pi76  & ~n634;
  assign n638 = ~n636 & ~n637;
  assign n639 = pi75  & ~n638;
  assign n640 = ~n635 & ~n639;
  assign n641 = ~pi73  & ~n640;
  assign n642 = ~pi74  & ~n638;
  assign n643 = pi74  & ~n640;
  assign n644 = ~n642 & ~n643;
  assign n645 = pi73  & ~n644;
  assign n646 = ~n641 & ~n645;
  assign n647 = ~pi71  & ~n646;
  assign n648 = ~pi72  & ~n644;
  assign n649 = pi72  & ~n646;
  assign n650 = ~n648 & ~n649;
  assign n651 = pi71  & ~n650;
  assign n652 = ~n647 & ~n651;
  assign n653 = ~pi69  & ~n652;
  assign n654 = ~pi70  & ~n650;
  assign n655 = pi70  & ~n652;
  assign n656 = ~n654 & ~n655;
  assign n657 = pi69  & ~n656;
  assign n658 = ~n653 & ~n657;
  assign n659 = ~pi67  & ~n658;
  assign n660 = ~pi68  & ~n656;
  assign n661 = pi68  & ~n658;
  assign n662 = ~n660 & ~n661;
  assign n663 = pi67  & ~n662;
  assign n664 = ~n659 & ~n663;
  assign n665 = ~pi65  & ~n664;
  assign n666 = ~pi66  & ~n662;
  assign n667 = pi66  & ~n664;
  assign n668 = ~n666 & ~n667;
  assign n669 = pi65  & ~n668;
  assign n670 = ~n665 & ~n669;
  assign n671 = ~pi63  & ~n670;
  assign n672 = ~pi64  & ~n668;
  assign n673 = pi64  & ~n670;
  assign n674 = ~n672 & ~n673;
  assign n675 = pi63  & ~n674;
  assign n676 = ~n671 & ~n675;
  assign n677 = ~pi61  & ~n676;
  assign n678 = ~pi62  & ~n674;
  assign n679 = pi62  & ~n676;
  assign n680 = ~n678 & ~n679;
  assign n681 = pi61  & ~n680;
  assign n682 = ~n677 & ~n681;
  assign n683 = ~pi59  & ~n682;
  assign n684 = ~pi60  & ~n680;
  assign n685 = pi60  & ~n682;
  assign n686 = ~n684 & ~n685;
  assign n687 = pi59  & ~n686;
  assign n688 = ~n683 & ~n687;
  assign n689 = ~pi57  & ~n688;
  assign n690 = ~pi58  & ~n686;
  assign n691 = pi58  & ~n688;
  assign n692 = ~n690 & ~n691;
  assign n693 = pi57  & ~n692;
  assign n694 = ~n689 & ~n693;
  assign n695 = ~pi55  & ~n694;
  assign n696 = ~pi56  & ~n692;
  assign n697 = pi56  & ~n694;
  assign n698 = ~n696 & ~n697;
  assign n699 = pi55  & ~n698;
  assign n700 = ~n695 & ~n699;
  assign n701 = ~pi53  & ~n700;
  assign n702 = ~pi54  & ~n698;
  assign n703 = pi54  & ~n700;
  assign n704 = ~n702 & ~n703;
  assign n705 = pi53  & ~n704;
  assign n706 = ~n701 & ~n705;
  assign n707 = ~pi51  & ~n706;
  assign n708 = ~pi52  & ~n704;
  assign n709 = pi52  & ~n706;
  assign n710 = ~n708 & ~n709;
  assign n711 = pi51  & ~n710;
  assign n712 = ~n707 & ~n711;
  assign n713 = ~pi49  & ~n712;
  assign n714 = ~pi50  & ~n710;
  assign n715 = pi50  & ~n712;
  assign n716 = ~n714 & ~n715;
  assign n717 = pi49  & ~n716;
  assign n718 = ~n713 & ~n717;
  assign n719 = ~pi47  & ~n718;
  assign n720 = ~pi48  & ~n716;
  assign n721 = pi48  & ~n718;
  assign n722 = ~n720 & ~n721;
  assign n723 = pi47  & ~n722;
  assign n724 = ~n719 & ~n723;
  assign n725 = ~pi45  & ~n724;
  assign n726 = ~pi46  & ~n722;
  assign n727 = pi46  & ~n724;
  assign n728 = ~n726 & ~n727;
  assign n729 = pi45  & ~n728;
  assign n730 = ~n725 & ~n729;
  assign n731 = ~pi43  & ~n730;
  assign n732 = ~pi44  & ~n728;
  assign n733 = pi44  & ~n730;
  assign n734 = ~n732 & ~n733;
  assign n735 = pi43  & ~n734;
  assign n736 = ~n731 & ~n735;
  assign n737 = pi42  & ~n736;
  assign n738 = ~pi42  & ~n734;
  assign n739 = pi1  & ~pi2 ;
  assign n740 = ~pi3  & ~n739;
  assign n741 = ~pi4  & ~n740;
  assign n742 = ~pi5  & ~n741;
  assign n743 = ~pi6  & ~n742;
  assign n744 = ~pi7  & ~n743;
  assign n745 = ~pi8  & ~n744;
  assign n746 = ~pi9  & ~n745;
  assign n747 = ~pi10  & ~n746;
  assign n748 = ~pi11  & ~n747;
  assign n749 = ~pi12  & ~n748;
  assign n750 = ~pi13  & ~n749;
  assign n751 = ~pi14  & ~n750;
  assign n752 = ~pi15  & ~n751;
  assign n753 = ~pi16  & ~n752;
  assign n754 = ~pi17  & ~n753;
  assign n755 = ~pi18  & ~n754;
  assign n756 = ~pi19  & ~n755;
  assign n757 = ~pi20  & ~n756;
  assign n758 = ~pi21  & ~n757;
  assign n759 = ~pi22  & ~n758;
  assign n760 = ~pi23  & ~n759;
  assign n761 = ~pi24  & ~n760;
  assign n762 = ~pi25  & ~n761;
  assign n763 = ~pi26  & ~n762;
  assign n764 = ~pi27  & ~n763;
  assign n765 = ~pi28  & ~n764;
  assign n766 = ~pi29  & ~n765;
  assign n767 = ~pi30  & ~n766;
  assign n768 = ~pi31  & ~n767;
  assign n769 = ~pi32  & ~n768;
  assign n770 = ~pi33  & ~n769;
  assign n771 = ~pi34  & ~n770;
  assign n772 = ~pi35  & ~n771;
  assign n773 = ~pi36  & ~n772;
  assign n774 = ~pi37  & ~n773;
  assign n775 = ~pi38  & ~n774;
  assign n776 = ~pi39  & ~n775;
  assign n777 = ~pi40  & ~n776;
  assign n778 = ~pi41  & ~n777;
  assign n779 = ~n738 & ~n778;
  assign n780 = ~n737 & n779;
  assign n781 = n736 & n778;
  assign n782 = ~pi41  & ~n736;
  assign n783 = ~n737 & ~n738;
  assign n784 = pi41  & ~n783;
  assign n785 = ~n782 & ~n784;
  assign n786 = ~pi39  & ~n785;
  assign n787 = ~pi40  & ~n783;
  assign n788 = pi40  & ~n785;
  assign n789 = ~n787 & ~n788;
  assign n790 = pi39  & ~n789;
  assign n791 = ~n786 & ~n790;
  assign n792 = ~pi37  & ~n791;
  assign n793 = ~pi38  & ~n789;
  assign n794 = pi38  & ~n791;
  assign n795 = ~n793 & ~n794;
  assign n796 = pi37  & ~n795;
  assign n797 = ~n792 & ~n796;
  assign n798 = ~pi35  & ~n797;
  assign n799 = ~pi36  & ~n795;
  assign n800 = pi36  & ~n797;
  assign n801 = ~n799 & ~n800;
  assign n802 = pi35  & ~n801;
  assign n803 = ~n798 & ~n802;
  assign n804 = ~pi33  & ~n803;
  assign n805 = ~pi34  & ~n801;
  assign n806 = pi34  & ~n803;
  assign n807 = ~n805 & ~n806;
  assign n808 = pi33  & ~n807;
  assign n809 = ~n804 & ~n808;
  assign n810 = ~pi31  & ~n809;
  assign n811 = ~pi32  & ~n807;
  assign n812 = pi32  & ~n809;
  assign n813 = ~n811 & ~n812;
  assign n814 = pi31  & ~n813;
  assign n815 = ~n810 & ~n814;
  assign n816 = ~pi29  & ~n815;
  assign n817 = ~pi30  & ~n813;
  assign n818 = pi30  & ~n815;
  assign n819 = ~n817 & ~n818;
  assign n820 = pi29  & ~n819;
  assign n821 = ~n816 & ~n820;
  assign n822 = ~pi27  & ~n821;
  assign n823 = ~pi28  & ~n819;
  assign n824 = pi28  & ~n821;
  assign n825 = ~n823 & ~n824;
  assign n826 = pi27  & ~n825;
  assign n827 = ~n822 & ~n826;
  assign n828 = ~pi25  & ~n827;
  assign n829 = ~pi26  & ~n825;
  assign n830 = pi26  & ~n827;
  assign n831 = ~n829 & ~n830;
  assign n832 = pi25  & ~n831;
  assign n833 = ~n828 & ~n832;
  assign n834 = pi24  & ~n833;
  assign n835 = ~pi24  & ~n831;
  assign n836 = ~n760 & ~n835;
  assign n837 = ~n834 & n836;
  assign n838 = n760 & n833;
  assign n839 = ~n837 & ~n838;
  assign n840 = ~pi23  & ~n833;
  assign n841 = ~n834 & ~n835;
  assign n842 = pi23  & ~n841;
  assign n843 = ~n840 & ~n842;
  assign n844 = ~pi21  & ~n843;
  assign n845 = ~pi22  & ~n841;
  assign n846 = pi22  & ~n843;
  assign n847 = ~n845 & ~n846;
  assign n848 = pi21  & ~n847;
  assign n849 = ~n844 & ~n848;
  assign n850 = ~pi19  & ~n849;
  assign n851 = ~pi20  & ~n847;
  assign n852 = pi20  & ~n849;
  assign n853 = ~n851 & ~n852;
  assign n854 = pi19  & ~n853;
  assign n855 = ~n850 & ~n854;
  assign n856 = ~pi17  & ~n855;
  assign n857 = ~pi18  & ~n853;
  assign n858 = pi18  & ~n855;
  assign n859 = ~n857 & ~n858;
  assign n860 = pi17  & ~n859;
  assign n861 = ~n856 & ~n860;
  assign n862 = ~pi15  & ~n861;
  assign n863 = ~pi16  & ~n859;
  assign n864 = pi16  & ~n861;
  assign n865 = ~n863 & ~n864;
  assign n866 = pi15  & ~n865;
  assign n867 = ~n862 & ~n866;
  assign n868 = ~pi13  & ~n867;
  assign n869 = ~pi14  & ~n865;
  assign n870 = pi14  & ~n867;
  assign n871 = ~n869 & ~n870;
  assign n872 = pi13  & ~n871;
  assign n873 = ~n868 & ~n872;
  assign n874 = ~pi11  & ~n873;
  assign n875 = ~pi12  & ~n871;
  assign n876 = pi12  & ~n873;
  assign n877 = ~n875 & ~n876;
  assign n878 = pi11  & ~n877;
  assign n879 = ~n874 & ~n878;
  assign n880 = ~pi9  & ~n879;
  assign n881 = ~pi10  & ~n877;
  assign n882 = pi10  & ~n879;
  assign n883 = ~n881 & ~n882;
  assign n884 = pi9  & ~n883;
  assign n885 = ~n880 & ~n884;
  assign n886 = ~pi7  & ~n885;
  assign n887 = ~pi8  & ~n883;
  assign n888 = pi8  & ~n885;
  assign n889 = ~n887 & ~n888;
  assign n890 = pi7  & ~n889;
  assign n891 = ~n886 & ~n890;
  assign n892 = pi6  & ~n891;
  assign n893 = ~pi6  & ~n889;
  assign n894 = ~n742 & ~n893;
  assign n895 = ~n892 & n894;
  assign n896 = n742 & n891;
  assign n897 = ~n895 & ~n896;
  assign n898 = ~n892 & ~n893;
  assign n899 = ~pi4  & ~n898;
  assign n900 = ~pi5  & ~n891;
  assign n901 = pi5  & ~n898;
  assign n902 = ~n900 & ~n901;
  assign n903 = pi4  & ~n902;
  assign n904 = ~n899 & ~n903;
  assign n905 = pi3  & ~n904;
  assign n906 = ~pi3  & ~n902;
  assign n907 = ~n739 & ~n906;
  assign n908 = ~n905 & ~n906;
  assign n909 = ~n739 & n908;
  assign n910 = ~n905 & n907;
  assign n911 = n739 & n904;
  assign n912 = ~n1772 & ~n911;
  assign n913 = ~n780 & ~n781;
  assign n914 = n207 & ~n208;
  assign n915 = n185 & ~n914;
  assign n916 = n184 & ~n915;
  assign n917 = n212 & ~n916;
  assign n918 = ~n213 & n915;
  assign n919 = n185 & ~n207;
  assign n920 = n213 & n919;
  assign n921 = n184 & ~n920;
  assign n922 = ~n918 & n921;
  assign n923 = ~n212 & ~n922;
  assign n924 = ~n917 & ~n923;
  assign n925 = ~n223 & n924;
  assign n926 = n223 & n922;
  assign n927 = ~n925 & ~n926;
  assign n928 = ~n222 & ~n927;
  assign n929 = n222 & n924;
  assign n930 = ~n928 & ~n929;
  assign n931 = ~n228 & ~n930;
  assign n932 = n228 & ~n927;
  assign n933 = ~n931 & ~n932;
  assign n934 = ~n227 & ~n933;
  assign n935 = n227 & ~n930;
  assign n936 = ~n934 & ~n935;
  assign n937 = ~n247 & ~n936;
  assign n938 = n247 & ~n933;
  assign n939 = ~n937 & ~n938;
  assign n940 = ~n246 & ~n939;
  assign n941 = n246 & ~n936;
  assign n942 = ~n940 & ~n941;
  assign n943 = ~n252 & ~n942;
  assign n944 = n252 & ~n939;
  assign n945 = ~n943 & ~n944;
  assign n946 = ~n251 & ~n945;
  assign n947 = n251 & ~n942;
  assign n948 = ~n946 & ~n947;
  assign n949 = ~n262 & ~n948;
  assign n950 = n262 & ~n945;
  assign n951 = ~n949 & ~n950;
  assign n952 = ~n261 & ~n951;
  assign n953 = n261 & ~n948;
  assign n954 = ~n952 & ~n953;
  assign n955 = ~n267 & ~n954;
  assign n956 = n267 & ~n951;
  assign n957 = ~n955 & ~n956;
  assign n958 = ~n266 & ~n957;
  assign n959 = n266 & ~n954;
  assign n960 = ~n958 & ~n959;
  assign n961 = ~n289 & ~n960;
  assign n962 = n289 & ~n957;
  assign n963 = ~n961 & ~n962;
  assign n964 = ~n288 & ~n963;
  assign n965 = n288 & ~n960;
  assign n966 = ~n964 & ~n965;
  assign n967 = ~n294 & ~n966;
  assign n968 = n294 & ~n963;
  assign n969 = ~n967 & ~n968;
  assign n970 = ~n293 & ~n969;
  assign n971 = n293 & ~n966;
  assign n972 = ~n970 & ~n971;
  assign n973 = ~n304 & ~n972;
  assign n974 = n304 & ~n969;
  assign n975 = ~n973 & ~n974;
  assign n976 = ~n303 & ~n975;
  assign n977 = n303 & ~n972;
  assign n978 = ~n976 & ~n977;
  assign n979 = ~n309 & ~n978;
  assign n980 = n309 & ~n975;
  assign n981 = ~n979 & ~n980;
  assign n982 = ~n308 & ~n981;
  assign n983 = n308 & ~n978;
  assign n984 = ~n982 & ~n983;
  assign n985 = ~n328 & ~n984;
  assign n986 = n328 & ~n981;
  assign n987 = ~n985 & ~n986;
  assign n988 = ~n327 & ~n987;
  assign n989 = n327 & ~n984;
  assign n990 = ~n988 & ~n989;
  assign n991 = ~n333 & ~n990;
  assign n992 = n333 & ~n987;
  assign n993 = ~n991 & ~n992;
  assign n994 = ~n332 & ~n993;
  assign n995 = n332 & ~n990;
  assign n996 = ~n994 & ~n995;
  assign n997 = ~n342 & ~n996;
  assign n998 = n342 & ~n993;
  assign n999 = ~n997 & ~n998;
  assign n1000 = ~n343 & ~n999;
  assign n1001 = n343 & ~n996;
  assign n1002 = ~n1000 & ~n1001;
  assign n1003 = ~n347 & ~n1002;
  assign n1004 = n347 & ~n999;
  assign n1005 = n180 & ~n1004;
  assign n1006 = ~n1003 & n1005;
  assign n1007 = n179 & ~n1006;
  assign n1008 = n438 & ~n442;
  assign n1009 = n437 & ~n1008;
  assign n1010 = n428 & ~n1009;
  assign n1011 = n427 & ~n1010;
  assign n1012 = n423 & ~n1011;
  assign n1013 = n422 & ~n1012;
  assign n1014 = n404 & ~n1013;
  assign n1015 = n403 & ~n1014;
  assign n1016 = n399 & ~n1015;
  assign n1017 = n398 & ~n1016;
  assign n1018 = n389 & ~n1017;
  assign n1019 = n388 & ~n1018;
  assign n1020 = n384 & ~n1019;
  assign n1021 = n383 & ~n1020;
  assign n1022 = n142 & n1021;
  assign n1023 = n1007 & n1022;
  assign n1024 = ~n348 & n1006;
  assign n1025 = n180 & n348;
  assign n1026 = n1002 & n1025;
  assign n1027 = n179 & ~n1026;
  assign n1028 = ~n1024 & n1027;
  assign n1029 = n170 & ~n1028;
  assign n1030 = ~n1023 & n1029;
  assign n1031 = n169 & ~n1030;
  assign n1032 = n164 & ~n1031;
  assign n1033 = n164 & n170;
  assign n1034 = n1021 & n1033;
  assign n1035 = ~n1007 & n1034;
  assign n1036 = n165 & ~n1035;
  assign n1037 = ~n1032 & n1036;
  assign n1038 = n143 & ~n1037;
  assign n1039 = n142 & ~n1038;
  assign n1040 = n164 & ~n169;
  assign n1041 = n165 & ~n1040;
  assign n1042 = n143 & ~n1041;
  assign n1043 = n179 & ~n1042;
  assign n1044 = ~n170 & n1041;
  assign n1045 = ~n164 & n165;
  assign n1046 = n170 & n1045;
  assign n1047 = n143 & ~n1046;
  assign n1048 = ~n1044 & n1047;
  assign n1049 = ~n179 & ~n1048;
  assign n1050 = ~n1043 & ~n1049;
  assign n1051 = ~n180 & n1050;
  assign n1052 = n180 & n1048;
  assign n1053 = ~n1051 & ~n1052;
  assign n1054 = ~n184 & ~n1053;
  assign n1055 = n184 & n1050;
  assign n1056 = ~n1054 & ~n1055;
  assign n1057 = ~n185 & ~n1056;
  assign n1058 = n185 & ~n1053;
  assign n1059 = ~n1057 & ~n1058;
  assign n1060 = ~n207 & ~n1059;
  assign n1061 = n207 & ~n1056;
  assign n1062 = ~n1060 & ~n1061;
  assign n1063 = ~n208 & ~n1062;
  assign n1064 = n208 & ~n1059;
  assign n1065 = ~n1063 & ~n1064;
  assign n1066 = ~n213 & ~n1065;
  assign n1067 = n213 & ~n1062;
  assign n1068 = ~n1066 & ~n1067;
  assign n1069 = ~n212 & ~n1068;
  assign n1070 = n212 & ~n1065;
  assign n1071 = ~n1069 & ~n1070;
  assign n1072 = ~n223 & ~n1071;
  assign n1073 = n223 & ~n1068;
  assign n1074 = ~n1072 & ~n1073;
  assign n1075 = ~n222 & ~n1074;
  assign n1076 = n222 & ~n1071;
  assign n1077 = ~n1075 & ~n1076;
  assign n1078 = ~n228 & ~n1077;
  assign n1079 = n228 & ~n1074;
  assign n1080 = ~n1078 & ~n1079;
  assign n1081 = ~n227 & ~n1080;
  assign n1082 = n227 & ~n1077;
  assign n1083 = ~n1081 & ~n1082;
  assign n1084 = ~n247 & ~n1083;
  assign n1085 = n247 & ~n1080;
  assign n1086 = ~n1084 & ~n1085;
  assign n1087 = ~n246 & ~n1086;
  assign n1088 = n246 & ~n1083;
  assign n1089 = ~n1087 & ~n1088;
  assign n1090 = ~n252 & ~n1089;
  assign n1091 = n252 & ~n1086;
  assign n1092 = ~n1090 & ~n1091;
  assign n1093 = ~n251 & ~n1092;
  assign n1094 = n251 & ~n1089;
  assign n1095 = ~n1093 & ~n1094;
  assign n1096 = ~n262 & ~n1095;
  assign n1097 = n262 & ~n1092;
  assign n1098 = ~n1096 & ~n1097;
  assign n1099 = ~n261 & ~n1098;
  assign n1100 = n261 & ~n1095;
  assign n1101 = ~n1099 & ~n1100;
  assign n1102 = ~n267 & ~n1101;
  assign n1103 = n267 & ~n1098;
  assign n1104 = ~n1102 & ~n1103;
  assign n1105 = ~n266 & ~n1104;
  assign n1106 = n266 & ~n1101;
  assign n1107 = ~n1105 & ~n1106;
  assign n1108 = ~n289 & ~n1107;
  assign n1109 = n289 & ~n1104;
  assign n1110 = ~n1108 & ~n1109;
  assign n1111 = ~n288 & ~n1110;
  assign n1112 = n288 & ~n1107;
  assign n1113 = ~n1111 & ~n1112;
  assign n1114 = ~n294 & ~n1113;
  assign n1115 = n294 & ~n1110;
  assign n1116 = ~n1114 & ~n1115;
  assign n1117 = ~n293 & ~n1116;
  assign n1118 = n293 & ~n1113;
  assign n1119 = ~n1117 & ~n1118;
  assign n1120 = ~n304 & ~n1119;
  assign n1121 = n304 & ~n1116;
  assign n1122 = ~n1120 & ~n1121;
  assign n1123 = ~n303 & ~n1122;
  assign n1124 = n303 & ~n1119;
  assign n1125 = ~n1123 & ~n1124;
  assign n1126 = ~n309 & ~n1125;
  assign n1127 = n309 & ~n1122;
  assign n1128 = ~n1126 & ~n1127;
  assign n1129 = ~n308 & ~n1128;
  assign n1130 = n308 & ~n1125;
  assign n1131 = ~n1129 & ~n1130;
  assign n1132 = ~n328 & ~n1131;
  assign n1133 = n328 & ~n1128;
  assign n1134 = ~n1132 & ~n1133;
  assign n1135 = ~n327 & ~n1134;
  assign n1136 = n327 & ~n1131;
  assign n1137 = ~n1135 & ~n1136;
  assign n1138 = ~n333 & ~n1137;
  assign n1139 = n333 & ~n1134;
  assign n1140 = ~n1138 & ~n1139;
  assign n1141 = ~n332 & ~n1140;
  assign n1142 = n332 & ~n1137;
  assign n1143 = ~n1141 & ~n1142;
  assign n1144 = ~n342 & ~n1143;
  assign n1145 = n342 & ~n1140;
  assign n1146 = ~n1144 & ~n1145;
  assign n1147 = ~n343 & ~n1146;
  assign n1148 = n343 & ~n1143;
  assign n1149 = ~n1147 & ~n1148;
  assign n1150 = ~n347 & ~n1149;
  assign n1151 = n347 & ~n1146;
  assign n1152 = ~n1150 & ~n1151;
  assign n1153 = ~n348 & ~n1152;
  assign n1154 = n348 & ~n1149;
  assign n1155 = n142 & ~n1021;
  assign n1156 = ~n1154 & n1155;
  assign n1157 = ~n1153 & n1156;
  assign n1158 = n1022 & n1152;
  assign n1159 = n138 & ~n1158;
  assign n1160 = ~n1157 & n1159;
  assign n1161 = n138 & ~n1039;
  assign n1162 = n137 & ~n1773;
  assign n1163 = n160 & ~n1162;
  assign n1164 = n159 & ~n1163;
  assign n1165 = n157 & ~n1164;
  assign n1166 = n157 & ~n159;
  assign n1167 = pi120  & n1166;
  assign n1168 = pi121  & n159;
  assign n1169 = ~pi120  & n157;
  assign n1170 = ~n1168 & n1169;
  assign n1171 = n1717 & ~n1170;
  assign n1172 = n157 & ~n1168;
  assign n1173 = n1717 & ~n1172;
  assign n1174 = ~pi120  & ~n1173;
  assign n1175 = n1717 & ~n1166;
  assign n1176 = pi120  & ~n1175;
  assign n1177 = ~n1174 & ~n1176;
  assign n1178 = ~n1167 & n1171;
  assign n1179 = ~n137 & n1774;
  assign n1180 = n137 & n1717;
  assign n1181 = n137 & n1175;
  assign n1182 = ~n1166 & n1180;
  assign n1183 = ~n1179 & ~n1775;
  assign n1184 = ~n138 & n1183;
  assign n1185 = n138 & ~n1774;
  assign n1186 = ~n1184 & ~n1185;
  assign n1187 = ~n142 & n1186;
  assign n1188 = n142 & ~n1183;
  assign n1189 = ~n142 & ~n1186;
  assign n1190 = n142 & n1183;
  assign n1191 = ~n1189 & ~n1190;
  assign n1192 = ~n1187 & ~n1188;
  assign n1193 = ~n143 & ~n1776;
  assign n1194 = n143 & ~n1186;
  assign n1195 = ~n1193 & ~n1194;
  assign n1196 = ~n165 & n1195;
  assign n1197 = n165 & n1776;
  assign n1198 = n165 & ~n1776;
  assign n1199 = ~n165 & ~n1195;
  assign n1200 = ~n1198 & ~n1199;
  assign n1201 = ~n1196 & ~n1197;
  assign n1202 = ~n164 & ~n1777;
  assign n1203 = n164 & ~n1195;
  assign n1204 = ~n1202 & ~n1203;
  assign n1205 = ~n169 & n1204;
  assign n1206 = n169 & n1777;
  assign n1207 = n169 & ~n1777;
  assign n1208 = ~n169 & ~n1204;
  assign n1209 = ~n1207 & ~n1208;
  assign n1210 = ~n1205 & ~n1206;
  assign n1211 = ~n170 & ~n1778;
  assign n1212 = n170 & ~n1204;
  assign n1213 = ~n1211 & ~n1212;
  assign n1214 = ~n179 & n1213;
  assign n1215 = n179 & n1778;
  assign n1216 = n179 & ~n1778;
  assign n1217 = ~n179 & ~n1213;
  assign n1218 = ~n1216 & ~n1217;
  assign n1219 = ~n1214 & ~n1215;
  assign n1220 = ~n180 & ~n1779;
  assign n1221 = n180 & ~n1213;
  assign n1222 = ~n1220 & ~n1221;
  assign n1223 = ~n184 & n1222;
  assign n1224 = n184 & n1779;
  assign n1225 = n184 & ~n1779;
  assign n1226 = ~n184 & ~n1222;
  assign n1227 = ~n1225 & ~n1226;
  assign n1228 = ~n1223 & ~n1224;
  assign n1229 = ~n185 & ~n1780;
  assign n1230 = n185 & ~n1222;
  assign n1231 = ~n1229 & ~n1230;
  assign n1232 = ~n207 & n1231;
  assign n1233 = n207 & n1780;
  assign n1234 = n207 & ~n1780;
  assign n1235 = ~n207 & ~n1231;
  assign n1236 = ~n1234 & ~n1235;
  assign n1237 = ~n1232 & ~n1233;
  assign n1238 = ~n208 & ~n1781;
  assign n1239 = n208 & ~n1231;
  assign n1240 = ~n1238 & ~n1239;
  assign n1241 = ~n213 & n1240;
  assign n1242 = n213 & n1781;
  assign n1243 = n213 & ~n1781;
  assign n1244 = ~n213 & ~n1240;
  assign n1245 = ~n1243 & ~n1244;
  assign n1246 = ~n1241 & ~n1242;
  assign n1247 = ~n212 & ~n1782;
  assign n1248 = n212 & ~n1240;
  assign n1249 = ~n1247 & ~n1248;
  assign n1250 = ~n223 & n1249;
  assign n1251 = n223 & n1782;
  assign n1252 = n223 & ~n1782;
  assign n1253 = ~n223 & ~n1249;
  assign n1254 = ~n1252 & ~n1253;
  assign n1255 = ~n1250 & ~n1251;
  assign n1256 = ~n222 & ~n1783;
  assign n1257 = n222 & ~n1249;
  assign n1258 = ~n1256 & ~n1257;
  assign n1259 = ~n228 & n1258;
  assign n1260 = n228 & n1783;
  assign n1261 = n228 & ~n1783;
  assign n1262 = ~n228 & ~n1258;
  assign n1263 = ~n1261 & ~n1262;
  assign n1264 = ~n1259 & ~n1260;
  assign n1265 = ~n227 & ~n1784;
  assign n1266 = n227 & ~n1258;
  assign n1267 = ~n1265 & ~n1266;
  assign n1268 = ~n247 & n1267;
  assign n1269 = n247 & n1784;
  assign n1270 = n247 & ~n1784;
  assign n1271 = ~n247 & ~n1267;
  assign n1272 = ~n1270 & ~n1271;
  assign n1273 = ~n1268 & ~n1269;
  assign n1274 = ~n246 & ~n1785;
  assign n1275 = n246 & ~n1267;
  assign n1276 = ~n1274 & ~n1275;
  assign n1277 = ~n252 & n1276;
  assign n1278 = n252 & n1785;
  assign n1279 = n252 & ~n1785;
  assign n1280 = ~n252 & ~n1276;
  assign n1281 = ~n1279 & ~n1280;
  assign n1282 = ~n1277 & ~n1278;
  assign n1283 = ~n251 & ~n1786;
  assign n1284 = n251 & ~n1276;
  assign n1285 = ~n1283 & ~n1284;
  assign n1286 = ~n262 & n1285;
  assign n1287 = n262 & n1786;
  assign n1288 = n262 & ~n1786;
  assign n1289 = ~n262 & ~n1285;
  assign n1290 = ~n1288 & ~n1289;
  assign n1291 = ~n1286 & ~n1287;
  assign n1292 = ~n261 & ~n1787;
  assign n1293 = n261 & ~n1285;
  assign n1294 = ~n1292 & ~n1293;
  assign n1295 = ~n267 & n1294;
  assign n1296 = n267 & n1787;
  assign n1297 = n267 & ~n1787;
  assign n1298 = ~n267 & ~n1294;
  assign n1299 = ~n1297 & ~n1298;
  assign n1300 = ~n1295 & ~n1296;
  assign n1301 = ~n266 & ~n1788;
  assign n1302 = n266 & ~n1294;
  assign n1303 = ~n1301 & ~n1302;
  assign n1304 = ~n289 & n1303;
  assign n1305 = n289 & n1788;
  assign n1306 = n289 & ~n1788;
  assign n1307 = ~n289 & ~n1303;
  assign n1308 = ~n1306 & ~n1307;
  assign n1309 = ~n1304 & ~n1305;
  assign n1310 = ~n288 & ~n1789;
  assign n1311 = n288 & ~n1303;
  assign n1312 = ~n1310 & ~n1311;
  assign n1313 = ~n294 & n1312;
  assign n1314 = n294 & n1789;
  assign n1315 = n294 & ~n1789;
  assign n1316 = ~n294 & ~n1312;
  assign n1317 = ~n1315 & ~n1316;
  assign n1318 = ~n1313 & ~n1314;
  assign n1319 = ~n293 & ~n1790;
  assign n1320 = n293 & ~n1312;
  assign n1321 = ~n1319 & ~n1320;
  assign n1322 = ~n304 & n1321;
  assign n1323 = n304 & n1790;
  assign n1324 = n304 & ~n1790;
  assign n1325 = ~n304 & ~n1321;
  assign n1326 = ~n1324 & ~n1325;
  assign n1327 = ~n1322 & ~n1323;
  assign n1328 = ~n303 & ~n1791;
  assign n1329 = n303 & ~n1321;
  assign n1330 = ~n1328 & ~n1329;
  assign n1331 = ~n309 & n1330;
  assign n1332 = n309 & n1791;
  assign n1333 = n309 & ~n1791;
  assign n1334 = ~n309 & ~n1330;
  assign n1335 = ~n1333 & ~n1334;
  assign n1336 = ~n1331 & ~n1332;
  assign n1337 = ~n308 & ~n1792;
  assign n1338 = n308 & ~n1330;
  assign n1339 = ~n1337 & ~n1338;
  assign n1340 = ~n328 & n1339;
  assign n1341 = n328 & n1792;
  assign n1342 = n328 & ~n1792;
  assign n1343 = ~n328 & ~n1339;
  assign n1344 = ~n1342 & ~n1343;
  assign n1345 = ~n1340 & ~n1341;
  assign n1346 = ~n327 & ~n1793;
  assign n1347 = n327 & ~n1339;
  assign n1348 = ~n1346 & ~n1347;
  assign n1349 = ~n333 & n1348;
  assign n1350 = n333 & n1793;
  assign n1351 = n333 & ~n1793;
  assign n1352 = ~n333 & ~n1348;
  assign n1353 = ~n1351 & ~n1352;
  assign n1354 = ~n1349 & ~n1350;
  assign n1355 = ~n332 & ~n1794;
  assign n1356 = n332 & ~n1348;
  assign n1357 = ~n1355 & ~n1356;
  assign n1358 = ~n342 & n1357;
  assign n1359 = n342 & n1794;
  assign n1360 = n342 & ~n1794;
  assign n1361 = ~n342 & ~n1357;
  assign n1362 = ~n1360 & ~n1361;
  assign n1363 = ~n1358 & ~n1359;
  assign n1364 = ~n343 & ~n1795;
  assign n1365 = n343 & ~n1357;
  assign n1366 = ~n1364 & ~n1365;
  assign n1367 = ~n347 & n1366;
  assign n1368 = n347 & n1795;
  assign n1369 = n347 & ~n1795;
  assign n1370 = ~n347 & ~n1366;
  assign n1371 = ~n1369 & ~n1370;
  assign n1372 = ~n1367 & ~n1368;
  assign n1373 = ~n348 & ~n1796;
  assign n1374 = n348 & ~n1366;
  assign n1375 = ~n1373 & ~n1374;
  assign n1376 = ~n383 & n1375;
  assign n1377 = n383 & n1796;
  assign n1378 = n383 & ~n1796;
  assign n1379 = ~n383 & ~n1375;
  assign n1380 = ~n1378 & ~n1379;
  assign n1381 = ~n1376 & ~n1377;
  assign n1382 = ~n384 & ~n1797;
  assign n1383 = n384 & ~n1375;
  assign n1384 = ~n1382 & ~n1383;
  assign n1385 = ~n388 & n1384;
  assign n1386 = n388 & n1797;
  assign n1387 = n388 & ~n1797;
  assign n1388 = ~n388 & ~n1384;
  assign n1389 = ~n1387 & ~n1388;
  assign n1390 = ~n1385 & ~n1386;
  assign n1391 = ~n389 & ~n1798;
  assign n1392 = n389 & ~n1384;
  assign n1393 = ~n1391 & ~n1392;
  assign n1394 = ~n398 & n1393;
  assign n1395 = n398 & n1798;
  assign n1396 = n398 & ~n1798;
  assign n1397 = ~n398 & ~n1393;
  assign n1398 = ~n1396 & ~n1397;
  assign n1399 = ~n1394 & ~n1395;
  assign n1400 = ~n399 & ~n1799;
  assign n1401 = n399 & ~n1393;
  assign n1402 = ~n1400 & ~n1401;
  assign n1403 = ~n403 & n1402;
  assign n1404 = n403 & n1799;
  assign n1405 = n403 & ~n1799;
  assign n1406 = ~n403 & ~n1402;
  assign n1407 = ~n1405 & ~n1406;
  assign n1408 = ~n1403 & ~n1404;
  assign n1409 = ~n404 & ~n1800;
  assign n1410 = n404 & ~n1402;
  assign n1411 = ~n1409 & ~n1410;
  assign n1412 = ~n422 & n1411;
  assign n1413 = n422 & n1800;
  assign n1414 = n422 & ~n1800;
  assign n1415 = ~n422 & ~n1411;
  assign n1416 = ~n1414 & ~n1415;
  assign n1417 = ~n1412 & ~n1413;
  assign n1418 = ~n423 & ~n1801;
  assign n1419 = n423 & ~n1411;
  assign n1420 = ~n1418 & ~n1419;
  assign n1421 = ~n427 & ~n1420;
  assign n1422 = n427 & ~n1801;
  assign n1423 = ~n1010 & ~n1422;
  assign n1424 = ~n1421 & n1423;
  assign n1425 = n1010 & n1420;
  assign n1426 = ~n1424 & ~n1425;
  assign n1427 = ~n427 & n1420;
  assign n1428 = n427 & n1801;
  assign n1429 = ~n1427 & ~n1428;
  assign n1430 = ~n428 & n1429;
  assign n1431 = n428 & ~n1420;
  assign n1432 = ~n1430 & ~n1431;
  assign n1433 = ~n437 & n1432;
  assign n1434 = n437 & ~n1429;
  assign n1435 = ~n1433 & ~n1434;
  assign n1436 = ~n438 & n1435;
  assign n1437 = n438 & ~n1432;
  assign n1438 = ~n442 & ~n1437;
  assign n1439 = ~n1436 & ~n1437;
  assign n1440 = ~n442 & n1439;
  assign n1441 = ~n1436 & n1438;
  assign n1442 = n442 & ~n1435;
  assign n1443 = ~n1803 & ~n1442;
  assign n1444 = n1717 & ~n1165;
  assign n1445 = n1763 & ~n1765;
  assign n1446 = n1762 & ~n1445;
  assign n1447 = n1759 & ~n1446;
  assign n1448 = n1758 & ~n1447;
  assign n1449 = n1756 & ~n1448;
  assign n1450 = n1755 & ~n1449;
  assign n1451 = n1751 & ~n1450;
  assign n1452 = n1750 & ~n1451;
  assign n1453 = n1748 & ~n1452;
  assign n1454 = n1747 & ~n1453;
  assign n1455 = n1744 & ~n1454;
  assign n1456 = n1743 & ~n1455;
  assign n1457 = n1741 & ~n1456;
  assign n1458 = n1740 & ~n1457;
  assign n1459 = n1737 & ~n1458;
  assign n1460 = n1736 & ~n1459;
  assign n1461 = n1734 & ~n1460;
  assign n1462 = n1733 & ~n1461;
  assign n1463 = n1727 & ~n1729;
  assign n1464 = n1726 & ~n1463;
  assign n1465 = n1722 & ~n1464;
  assign n1466 = n1721 & ~n1465;
  assign n1467 = n1719 & ~n1466;
  assign n1468 = n1722 & ~n1726;
  assign n1469 = n1721 & ~n1468;
  assign n1470 = ~n1727 & n1469;
  assign n1471 = n1721 & n1727;
  assign n1472 = ~n1722 & n1471;
  assign n1473 = n1719 & ~n1472;
  assign n1474 = ~n1470 & n1473;
  assign n1475 = ~n1729 & n1474;
  assign n1476 = n1719 & n1729;
  assign n1477 = ~n1469 & n1476;
  assign n1478 = n1718 & ~n1477;
  assign n1479 = ~n1475 & n1478;
  assign n1480 = n1718 & ~n1467;
  assign n1481 = n144 & ~n1804;
  assign n1482 = n1714 & ~n1481;
  assign n1483 = n1462 & n1482;
  assign n1484 = n1729 & ~n1730;
  assign n1485 = n1727 & ~n1484;
  assign n1486 = n1726 & ~n1485;
  assign n1487 = n1722 & ~n1486;
  assign n1488 = n1721 & ~n1487;
  assign n1489 = n1719 & ~n1488;
  assign n1490 = n1718 & ~n1489;
  assign n1491 = ~n1730 & n1804;
  assign n1492 = n1718 & n1730;
  assign n1493 = ~n1474 & n1492;
  assign n1494 = n144 & ~n1493;
  assign n1495 = ~n1491 & n1494;
  assign n1496 = n144 & ~n1490;
  assign n1497 = n1714 & ~n1805;
  assign n1498 = ~n1462 & n1497;
  assign n1499 = n161 & ~n1498;
  assign n1500 = ~n1483 & n1499;
  assign n1501 = ~n1714 & n161;
  assign n1502 = n158 & ~n1501;
  assign n1503 = ~n1716 & n1502;
  assign n1504 = pi115  & n1714;
  assign n1505 = n161 & ~n1504;
  assign n1506 = n1716 & n158;
  assign n1507 = n158 & ~n1505;
  assign n1508 = n1716 & n1507;
  assign n1509 = ~n1505 & n1506;
  assign n1510 = ~n1503 & ~n1806;
  assign n1511 = ~n1718 & n1510;
  assign n1512 = n1718 & ~n1502;
  assign n1513 = ~n1511 & ~n1512;
  assign n1514 = ~n1719 & n1513;
  assign n1515 = n1719 & ~n1510;
  assign n1516 = ~n1514 & ~n1515;
  assign n1517 = ~n1721 & n1516;
  assign n1518 = n1721 & ~n1513;
  assign n1519 = ~n1517 & ~n1518;
  assign n1520 = ~n1722 & n1519;
  assign n1521 = n1722 & ~n1516;
  assign n1522 = ~n1520 & ~n1521;
  assign n1523 = ~n1726 & n1522;
  assign n1524 = n1726 & ~n1519;
  assign n1525 = ~n1523 & ~n1524;
  assign n1526 = ~n1727 & n1525;
  assign n1527 = n1727 & ~n1522;
  assign n1528 = ~n1526 & ~n1527;
  assign n1529 = ~n1729 & n1528;
  assign n1530 = n1729 & ~n1525;
  assign n1531 = ~n1529 & ~n1530;
  assign n1532 = ~n1730 & n1531;
  assign n1533 = n1730 & ~n1528;
  assign n1534 = ~n1532 & ~n1533;
  assign n1535 = ~n1733 & n1534;
  assign n1536 = n1733 & ~n1531;
  assign n1537 = ~n1535 & ~n1536;
  assign n1538 = ~n1734 & n1537;
  assign n1539 = n1734 & ~n1534;
  assign n1540 = ~n1538 & ~n1539;
  assign n1541 = ~n1736 & n1540;
  assign n1542 = n1736 & ~n1537;
  assign n1543 = ~n1541 & ~n1542;
  assign n1544 = ~n1737 & n1543;
  assign n1545 = n1737 & ~n1540;
  assign n1546 = ~n1544 & ~n1545;
  assign n1547 = ~n1740 & n1546;
  assign n1548 = n1740 & ~n1543;
  assign n1549 = ~n1547 & ~n1548;
  assign n1550 = ~n1741 & n1549;
  assign n1551 = n1741 & ~n1546;
  assign n1552 = ~n1550 & ~n1551;
  assign n1553 = ~n1743 & n1552;
  assign n1554 = n1743 & ~n1549;
  assign n1555 = ~n1553 & ~n1554;
  assign n1556 = ~n1744 & n1555;
  assign n1557 = n1744 & ~n1552;
  assign n1558 = ~n1556 & ~n1557;
  assign n1559 = ~n1747 & n1558;
  assign n1560 = n1747 & ~n1555;
  assign n1561 = ~n1559 & ~n1560;
  assign n1562 = ~n1748 & n1561;
  assign n1563 = n1748 & ~n1558;
  assign n1564 = ~n1562 & ~n1563;
  assign n1565 = ~n1750 & n1564;
  assign n1566 = n1750 & ~n1561;
  assign n1567 = ~n1565 & ~n1566;
  assign n1568 = ~n1751 & n1567;
  assign n1569 = n1751 & ~n1564;
  assign n1570 = ~n1568 & ~n1569;
  assign n1571 = ~n1755 & n1570;
  assign n1572 = n1755 & ~n1567;
  assign n1573 = ~n1571 & ~n1572;
  assign n1574 = ~n1756 & n1573;
  assign n1575 = n1756 & ~n1570;
  assign n1576 = ~n1574 & ~n1575;
  assign n1577 = ~n1758 & n1576;
  assign n1578 = n1758 & ~n1573;
  assign n1579 = ~n1447 & ~n1578;
  assign n1580 = ~n1577 & n1579;
  assign n1581 = n1447 & ~n1576;
  assign n1582 = ~n1580 & ~n1581;
  assign n1583 = ~n1577 & ~n1578;
  assign n1584 = ~n1759 & n1583;
  assign n1585 = n1759 & ~n1576;
  assign n1586 = ~n1584 & ~n1585;
  assign n1587 = ~n1762 & n1586;
  assign n1588 = n1762 & ~n1583;
  assign n1589 = ~n1587 & ~n1588;
  assign n1590 = ~n1763 & n1589;
  assign n1591 = n1763 & ~n1586;
  assign n1592 = ~n1765 & ~n1591;
  assign n1593 = ~n1590 & ~n1591;
  assign n1594 = ~n1765 & n1593;
  assign n1595 = ~n1590 & n1592;
  assign n1596 = n1765 & ~n1589;
  assign n1597 = ~n1808 & ~n1596;
  assign n1598 = n158 & ~n1500;
  assign n1599 = n1760 & ~n1764;
  assign n1600 = n1757 & ~n1599;
  assign n1601 = n1752 & ~n1600;
  assign n1602 = n1749 & ~n1601;
  assign n1603 = n1745 & ~n1602;
  assign n1604 = n1742 & ~n1603;
  assign n1605 = n1738 & ~n1604;
  assign n1606 = n1735 & ~n1605;
  assign n1607 = n1731 & ~n1606;
  assign n1608 = n1728 & ~n1607;
  assign n1609 = n1715 & ~n1720;
  assign n1610 = n1608 & n1609;
  assign n1611 = n1720 & ~n189;
  assign n1612 = n1715 & ~n1611;
  assign n1613 = ~n1608 & n1612;
  assign n1614 = n162 & ~n1613;
  assign n1615 = n162 & ~n1609;
  assign n1616 = ~n1725 & n1615;
  assign n1617 = pi103  & n1720;
  assign n1618 = n1715 & ~n1617;
  assign n1619 = n162 & n1725;
  assign n1620 = n162 & ~n1618;
  assign n1621 = n1725 & n1620;
  assign n1622 = ~n1618 & n1619;
  assign n1623 = ~n1616 & ~n1809;
  assign n1624 = ~n1728 & n1623;
  assign n1625 = n1728 & ~n1615;
  assign n1626 = ~n1624 & ~n1625;
  assign n1627 = ~n1731 & n1626;
  assign n1628 = n1731 & ~n1623;
  assign n1629 = ~n1627 & ~n1628;
  assign n1630 = ~n1735 & n1629;
  assign n1631 = n1735 & ~n1626;
  assign n1632 = ~n1630 & ~n1631;
  assign n1633 = ~n1738 & n1632;
  assign n1634 = n1738 & ~n1629;
  assign n1635 = ~n1633 & ~n1634;
  assign n1636 = ~n1742 & n1635;
  assign n1637 = n1742 & ~n1632;
  assign n1638 = ~n1636 & ~n1637;
  assign n1639 = ~n1745 & n1638;
  assign n1640 = n1745 & ~n1635;
  assign n1641 = ~n1639 & ~n1640;
  assign n1642 = ~n1749 & n1641;
  assign n1643 = n1749 & ~n1638;
  assign n1644 = ~n1601 & ~n1643;
  assign n1645 = ~n1642 & n1644;
  assign n1646 = n1601 & ~n1641;
  assign n1647 = ~n1645 & ~n1646;
  assign n1648 = ~n1642 & ~n1643;
  assign n1649 = ~n1752 & n1648;
  assign n1650 = n1752 & ~n1641;
  assign n1651 = ~n1649 & ~n1650;
  assign n1652 = ~n1757 & n1651;
  assign n1653 = n1757 & ~n1648;
  assign n1654 = ~n1652 & ~n1653;
  assign n1655 = ~n1760 & n1654;
  assign n1656 = n1760 & ~n1651;
  assign n1657 = ~n1764 & ~n1656;
  assign n1658 = ~n1655 & ~n1656;
  assign n1659 = ~n1764 & n1658;
  assign n1660 = ~n1655 & n1657;
  assign n1661 = n1764 & ~n1654;
  assign n1662 = ~n1811 & ~n1661;
  assign n1663 = ~n1610 & n1614;
  assign n1664 = n1723 & ~n1732;
  assign n1665 = n163 & ~n1664;
  assign n1666 = n1753 & ~n1761;
  assign n1667 = n1746 & ~n1666;
  assign n1668 = ~pi77  & ~pi78 ;
  assign n1669 = ~pi76  & n1668;
  assign n1670 = ~pi78  & n246;
  assign n1671 = ~pi75  & n1812;
  assign n1672 = ~pi74  & n1671;
  assign n1673 = ~pi73  & n1672;
  assign n1674 = ~pi72  & n1673;
  assign n1675 = n1734 & n1812;
  assign n1676 = ~pi71  & n1813;
  assign n1677 = ~pi70  & n1676;
  assign n1678 = ~pi69  & n1677;
  assign n1679 = ~pi68  & n1678;
  assign n1680 = ~pi67  & n1679;
  assign n1681 = ~pi66  & n1680;
  assign n1682 = ~pi65  & n1681;
  assign n1683 = ~pi64  & n1682;
  assign n1684 = n1738 & n1813;
  assign n1685 = ~n1667 & n1814;
  assign n1686 = n1665 & ~n1685;
  assign n1687 = pi79  & n1732;
  assign n1688 = n1723 & ~n1687;
  assign n1689 = n163 & ~n1688;
  assign n1690 = n1685 & n1689;
  assign n1691 = n276 & ~n1667;
  assign n1692 = n1732 & ~n1691;
  assign n1693 = n1723 & ~n1692;
  assign n1694 = n163 & ~n1693;
  assign n1695 = n1665 & ~n1814;
  assign n1696 = n163 & n1814;
  assign n1697 = n1814 & n1689;
  assign n1698 = ~n1688 & n1696;
  assign n1699 = ~n1695 & ~n1816;
  assign n1700 = ~n1746 & n1699;
  assign n1701 = n1746 & ~n1665;
  assign n1702 = ~n1700 & ~n1701;
  assign n1703 = ~n1753 & n1702;
  assign n1704 = n1753 & ~n1699;
  assign n1705 = ~n1761 & ~n1704;
  assign n1706 = ~n1703 & ~n1704;
  assign n1707 = ~n1761 & n1706;
  assign n1708 = ~n1703 & n1705;
  assign n1709 = n1761 & ~n1702;
  assign n1710 = ~n1817 & ~n1709;
  assign n1711 = ~n1686 & ~n1690;
  assign n1712 = n1739 & ~n1754;
  assign n1713 = n206 & ~n1712;
  assign n1714 = n140 | n141;
  assign n1715 = n153 | n147 | n152;
  assign n1716 = n149 | n150;
  assign n1717 = n155 | n156;
  assign n1718 = n167 | n168;
  assign n1719 = n172 | n173;
  assign n1720 = n177 | n178;
  assign n1721 = n182 | n183;
  assign n1722 = n187 | n188;
  assign n1723 = n205 | n194 | n204;
  assign n1724 = n196 | n197;
  assign n1725 = n201 | n202;
  assign n1726 = n210 | n211;
  assign n1727 = n215 | n216;
  assign n1728 = n220 | n221;
  assign n1729 = n225 | n226;
  assign n1730 = n230 | n231;
  assign n1731 = n235 | n236;
  assign n1732 = n244 | n245;
  assign n1733 = n249 | n250;
  assign n1734 = n254 | n255;
  assign n1735 = n259 | n260;
  assign n1736 = n264 | n265;
  assign n1737 = n269 | n270;
  assign n1738 = n274 | n275;
  assign n1739 = n285 | n286;
  assign n1740 = n291 | n292;
  assign n1741 = n296 | n297;
  assign n1742 = n301 | n302;
  assign n1743 = n306 | n307;
  assign n1744 = n311 | n312;
  assign n1745 = n316 | n317;
  assign n1746 = n325 | n326;
  assign n1747 = n330 | n331;
  assign n1748 = n335 | n336;
  assign n1749 = n340 | n341;
  assign n1750 = n345 | n346;
  assign n1751 = n350 | n351;
  assign n1752 = n355 | n356;
  assign n1753 = n364 | n365;
  assign n1754 = n381 | n382;
  assign n1755 = n386 | n387;
  assign n1756 = n391 | n392;
  assign n1757 = n396 | n397;
  assign n1758 = n401 | n402;
  assign n1759 = n406 | n407;
  assign n1760 = n411 | n412;
  assign n1761 = n420 | n421;
  assign n1762 = n425 | n426;
  assign n1763 = n430 | n431;
  assign n1764 = n435 | n436;
  assign n1765 = n440 | n441;
  assign n1766 = n456 | n457;
  assign n1767 = n490 | n491;
  assign n1768 = n493 | n494;
  assign n1769 = n510 | n511;
  assign n1770 = n513 | n514;
  assign po0  = n839 | n897 | n912 | n913;
  assign n1772 = n909 | n910;
  assign n1773 = n1160 | n1161;
  assign n1774 = n1177 | n1178;
  assign n1775 = n1181 | n1182;
  assign n1776 = n1191 | ~n1192;
  assign n1777 = n1200 | ~n1201;
  assign n1778 = n1209 | ~n1210;
  assign n1779 = n1218 | ~n1219;
  assign n1780 = n1227 | ~n1228;
  assign n1781 = n1236 | ~n1237;
  assign n1782 = n1245 | ~n1246;
  assign n1783 = n1254 | ~n1255;
  assign n1784 = n1263 | ~n1264;
  assign n1785 = n1272 | ~n1273;
  assign n1786 = n1281 | ~n1282;
  assign n1787 = n1290 | ~n1291;
  assign n1788 = n1299 | ~n1300;
  assign n1789 = n1308 | ~n1309;
  assign n1790 = n1317 | ~n1318;
  assign n1791 = n1326 | ~n1327;
  assign n1792 = n1335 | ~n1336;
  assign n1793 = n1344 | ~n1345;
  assign n1794 = n1353 | ~n1354;
  assign n1795 = n1362 | ~n1363;
  assign n1796 = n1371 | ~n1372;
  assign n1797 = n1380 | ~n1381;
  assign n1798 = n1389 | ~n1390;
  assign n1799 = n1398 | ~n1399;
  assign n1800 = n1407 | ~n1408;
  assign n1801 = n1416 | ~n1417;
  assign po1  = ~n1444 | n1426 | n1443;
  assign n1803 = n1440 | n1441;
  assign n1804 = n1479 | n1480;
  assign n1805 = n1495 | n1496;
  assign n1806 = n1508 | n1509;
  assign po2  = ~n1598 | n1582 | ~n1597;
  assign n1808 = n1594 | n1595;
  assign n1809 = n1621 | n1622;
  assign po3  = ~n1663 | n1647 | ~n1662;
  assign n1811 = n1659 | n1660;
  assign n1812 = n1669 | n1670;
  assign n1813 = n1674 | n1675;
  assign n1814 = n1683 | n1684;
  assign n1815 = ~n1711 | n1694 | n1710;
  assign n1816 = n1697 | n1698;
  assign n1817 = n1707 | n1708;
  assign po4  = ~n1815;
  assign po5  = ~n1713;
  assign po6  = ~n287;
  assign po7 = ~n1766;
endmodule
