module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 , pi32 ,
    pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 , pi40 ,
    pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 , pi56 ,
    pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 , pi64 ,
    pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 ,
    pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 ,
    pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 ,
    pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 ,
    pi97 , pi98 , pi99 , pi100 , pi101 , pi102 , pi103 ,
    pi104 , pi105 , pi106 , pi107 , pi108 , pi109 , pi110 ,
    pi111 , pi112 , pi113 , pi114 , pi115 , pi116 , pi117 ,
    pi118 , pi119 , pi120 , pi121 , pi122 , pi123 , pi124 ,
    pi125 , pi126 , pi127 , pi128 , pi129 , pi130 , pi131 , pi132 ,
    pi133 , pi134 , pi135 , pi136 , pi137 , pi138 , pi139 , pi140 ,
    pi141 , pi142 , pi143 , pi144 , pi145 , pi146 , pi147 , pi148 ,
    pi149 , pi150 , pi151 , pi152 , pi153 , pi154 , pi155 , pi156 ,
    pi157 , pi158 , pi159 , pi160 , pi161 , pi162 , pi163 , pi164 ,
    pi165 , pi166 , pi167 , pi168 , pi169 , pi170 , pi171 , pi172 ,
    pi173 , pi174 , pi175 , pi176 , pi177 , pi178 , pi179 , pi180 ,
    pi181 , pi182 , pi183 , pi184 , pi185 , pi186 , pi187 , pi188 ,
    pi189 , pi190 , pi191 , pi192 , pi193 , pi194 , pi195 , pi196 ,
    pi197 , pi198 , pi199 , pi200 , pi201 , pi202 , pi203 , pi204 ,
    pi205 , pi206 , pi207 , pi208 , pi209 , pi210 , pi211 , pi212 ,
    pi213 , pi214 , pi215 , pi216 , pi217 , pi218 , pi219 , pi220 ,
    pi221 , pi222 , pi223 , pi224 , pi225 , pi226 , pi227 ,
    pi228 , pi229 , pi230 , pi231 , pi232 , pi233 , pi234 ,
    pi235 , pi236 , pi237 , pi238 , pi239 , pi240 , pi241 ,
    pi242 , pi243 , pi244 , pi245 , pi246 , pi247 , pi248 ,
    pi249 , pi250 , pi251 , pi252 , pi253 , pi254 , pi255 ,
    po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7 , po8 ,
    po9 , po10 , po11 , po12 , po13 , po14 , po15 , po16 ,
    po17 , po18 , po19 , po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 , po30 , po31 , po32 ,
    po33 , po34 , po35 , po36 , po37 , po38 , po39 , po40 ,
    po41 , po42 , po43 , po44 , po45 , po46 , po47 , po48 ,
    po49 , po50 , po51 , po52 , po53 , po54 , po55 , po56 ,
    po57 , po58 , po59 , po60 , po61 , po62 , po63 , po64 ,
    po65 , po66 , po67 , po68 , po69 , po70 , po71 , po72 ,
    po73 , po74 , po75 , po76 , po77 , po78 , po79 , po80 ,
    po81 , po82 , po83 , po84 , po85 , po86 , po87 , po88 ,
    po89 , po90 , po91 , po92 , po93 , po94 , po95 , po96 ,
    po97 , po98 , po99 , po100 , po101 , po102 , po103 ,
    po104 , po105 , po106 , po107 , po108 , po109 , po110 ,
    po111 , po112 , po113 , po114 , po115 , po116 , po117 ,
    po118 , po119 , po120 , po121 , po122 , po123 , po124 ,
    po125 , po126 , po127 , po128  );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    pi32 , pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 ,
    pi56 , pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 ,
    pi64 , pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 ,
    pi72 , pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 ,
    pi80 , pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 ,
    pi88 , pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 ,
    pi96 , pi97 , pi98 , pi99 , pi100 , pi101 , pi102 ,
    pi103 , pi104 , pi105 , pi106 , pi107 , pi108 , pi109 ,
    pi110 , pi111 , pi112 , pi113 , pi114 , pi115 , pi116 ,
    pi117 , pi118 , pi119 , pi120 , pi121 , pi122 , pi123 ,
    pi124 , pi125 , pi126 , pi127 , pi128 , pi129 , pi130 , pi131 ,
    pi132 , pi133 , pi134 , pi135 , pi136 , pi137 , pi138 , pi139 ,
    pi140 , pi141 , pi142 , pi143 , pi144 , pi145 , pi146 , pi147 ,
    pi148 , pi149 , pi150 , pi151 , pi152 , pi153 , pi154 , pi155 ,
    pi156 , pi157 , pi158 , pi159 , pi160 , pi161 , pi162 , pi163 ,
    pi164 , pi165 , pi166 , pi167 , pi168 , pi169 , pi170 , pi171 ,
    pi172 , pi173 , pi174 , pi175 , pi176 , pi177 , pi178 , pi179 ,
    pi180 , pi181 , pi182 , pi183 , pi184 , pi185 , pi186 , pi187 ,
    pi188 , pi189 , pi190 , pi191 , pi192 , pi193 , pi194 , pi195 ,
    pi196 , pi197 , pi198 , pi199 , pi200 , pi201 , pi202 , pi203 ,
    pi204 , pi205 , pi206 , pi207 , pi208 , pi209 , pi210 , pi211 ,
    pi212 , pi213 , pi214 , pi215 , pi216 , pi217 , pi218 , pi219 ,
    pi220 , pi221 , pi222 , pi223 , pi224 , pi225 , pi226 , pi227 ,
    pi228 , pi229 , pi230 , pi231 , pi232 , pi233 , pi234 ,
    pi235 , pi236 , pi237 , pi238 , pi239 , pi240 , pi241 ,
    pi242 , pi243 , pi244 , pi245 , pi246 , pi247 , pi248 ,
    pi249 , pi250 , pi251 , pi252 , pi253 , pi254 , pi255 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7 ,
    po8 , po9 , po10 , po11 , po12 , po13 , po14 , po15 ,
    po16 , po17 , po18 , po19 , po20 , po21 , po22 , po23 ,
    po24 , po25 , po26 , po27 , po28 , po29 , po30 , po31 ,
    po32 , po33 , po34 , po35 , po36 , po37 , po38 , po39 ,
    po40 , po41 , po42 , po43 , po44 , po45 , po46 , po47 ,
    po48 , po49 , po50 , po51 , po52 , po53 , po54 , po55 ,
    po56 , po57 , po58 , po59 , po60 , po61 , po62 , po63 ,
    po64 , po65 , po66 , po67 , po68 , po69 , po70 , po71 ,
    po72 , po73 , po74 , po75 , po76 , po77 , po78 , po79 ,
    po80 , po81 , po82 , po83 , po84 , po85 , po86 , po87 ,
    po88 , po89 , po90 , po91 , po92 , po93 , po94 , po95 ,
    po96 , po97 , po98 , po99 , po100 , po101 , po102 ,
    po103 , po104 , po105 , po106 , po107 , po108 , po109 ,
    po110 , po111 , po112 , po113 , po114 , po115 , po116 ,
    po117 , po118 , po119 , po120 , po121 , po122 , po123 ,
    po124 , po125 , po126 , po127 , po128;
  wire n386, n387, n388, n389, n390, n391, n392,
    n393, n394, n395, n396, n397, n398, n399,
    n400, n401, n402, n403, n404, n405, n406,
    n407, n408, n409, n410, n411, n412, n413,
    n414, n415, n416, n417, n418, n419, n420,
    n421, n422, n423, n424, n425, n426, n427,
    n428, n429, n430, n431, n432, n433, n434,
    n435, n436, n437, n438, n439, n440, n441,
    n442, n443, n444, n445, n446, n447, n448,
    n449, n450, n451, n452, n453, n454, n455,
    n456, n457, n458, n459, n460, n461, n462,
    n463, n464, n465, n466, n467, n468, n469,
    n470, n471, n472, n473, n474, n475, n476,
    n477, n478, n479, n480, n481, n482, n483,
    n484, n485, n486, n487, n488, n489, n490,
    n491, n492, n493, n494, n495, n496, n497,
    n498, n499, n500, n501, n502, n503, n504,
    n505, n506, n507, n508, n509, n510, n511,
    n512, n513, n514, n515, n516, n517, n518,
    n519, n520, n521, n522, n523, n524, n525,
    n526, n527, n528, n529, n530, n531, n532,
    n533, n534, n535, n536, n537, n538, n539,
    n540, n541, n542, n543, n544, n545, n546,
    n547, n548, n549, n550, n551, n552, n553,
    n554, n555, n556, n557, n558, n559, n560,
    n561, n562, n563, n564, n565, n566, n567,
    n568, n569, n570, n571, n572, n573, n574,
    n575, n576, n577, n578, n579, n580, n581,
    n582, n583, n584, n585, n586, n587, n588,
    n589, n590, n591, n592, n593, n594, n595,
    n596, n597, n598, n599, n600, n601, n602,
    n603, n604, n605, n606, n607, n608, n609,
    n610, n611, n612, n613, n614, n615, n616,
    n617, n618, n619, n620, n621, n622, n623,
    n624, n625, n626, n627, n628, n629, n630,
    n631, n632, n633, n634, n635, n636, n637,
    n638, n639, n640, n641, n642, n643, n644,
    n645, n646, n647, n648, n649, n650, n651,
    n652, n653, n654, n655, n656, n657, n658,
    n659, n660, n661, n662, n663, n664, n665,
    n666, n667, n668, n669, n670, n671, n672,
    n673, n674, n675, n676, n677, n678, n679,
    n680, n681, n682, n683, n684, n685, n686,
    n687, n688, n689, n690, n691, n692, n693,
    n694, n695, n696, n697, n698, n699, n700,
    n701, n702, n703, n704, n705, n706, n707,
    n708, n709, n710, n711, n712, n713, n714,
    n715, n716, n717, n718, n719, n720, n721,
    n722, n723, n724, n725, n726, n727, n728,
    n729, n730, n731, n732, n733, n734, n735,
    n736, n737, n738, n739, n740, n741, n742,
    n743, n744, n745, n746, n747, n748, n749,
    n750, n751, n752, n753, n754, n755, n756,
    n757, n758, n759, n760, n761, n762, n763,
    n764, n765, n766, n767, n768, n769, n770,
    n771, n772, n773, n774, n775, n776, n777,
    n778, n779, n780, n781, n782, n783, n784,
    n785, n786, n787, n788, n789, n790, n791,
    n792, n793, n794, n795, n796, n797, n798,
    n799, n800, n801, n802, n803, n804, n805,
    n806, n807, n808, n809, n810, n811, n812,
    n813, n814, n815, n816, n817, n818, n819,
    n820, n821, n822, n823, n824, n825, n826,
    n827, n828, n829, n830, n831, n832, n833,
    n834, n835, n836, n837, n838, n839, n840,
    n841, n842, n843, n844, n845, n846, n847,
    n848, n849, n850, n851, n852, n853, n854,
    n855, n856, n857, n858, n859, n860, n861,
    n862, n863, n864, n865, n866, n867, n868,
    n869, n870, n871, n872, n873, n874, n875,
    n876, n877, n878, n879, n880, n881, n882,
    n883, n884, n885, n886, n887, n888, n889,
    n890, n891, n892, n893, n894, n895, n896,
    n897, n898, n899, n900, n901, n902, n903,
    n904, n905, n906, n907, n908, n909, n910,
    n911, n912, n913, n914, n915, n916, n917,
    n918, n919, n920, n921, n922, n923, n924,
    n925, n926, n927, n928, n929, n930, n931,
    n932, n933, n934, n935, n936, n937, n938,
    n939, n940, n941, n942, n943, n944, n945,
    n946, n947, n948, n949, n950, n951, n952,
    n953, n954, n955, n956, n957, n958, n959,
    n960, n961, n962, n963, n964, n965, n966,
    n967, n968, n969, n970, n971, n972, n973,
    n974, n975, n976, n977, n978, n979, n980,
    n981, n982, n983, n984, n985, n986, n987,
    n988, n989, n990, n991, n992, n993, n994,
    n995, n996, n997, n998, n999, n1000, n1001,
    n1002, n1003, n1004, n1005, n1006, n1007,
    n1008, n1009, n1010, n1011, n1012, n1013,
    n1014, n1015, n1016, n1017, n1018, n1019,
    n1020, n1021, n1022, n1023, n1024, n1025,
    n1026, n1027, n1028, n1029, n1030, n1031,
    n1032, n1033, n1034, n1035, n1036, n1037,
    n1038, n1039, n1040, n1041, n1042, n1043,
    n1044, n1045, n1046, n1047, n1048, n1049,
    n1050, n1051, n1052, n1053, n1054, n1055,
    n1056, n1057, n1058, n1059, n1060, n1061,
    n1062, n1063, n1064, n1065, n1066, n1067,
    n1068, n1069, n1070, n1071, n1072, n1073,
    n1074, n1075, n1076, n1077, n1078, n1079,
    n1080, n1081, n1082, n1083, n1084, n1085,
    n1086, n1087, n1088, n1089, n1090, n1091,
    n1092, n1093, n1094, n1095, n1096, n1097,
    n1098, n1099, n1100, n1101, n1102, n1103,
    n1104, n1105, n1106, n1107, n1108, n1109,
    n1110, n1111, n1112, n1113, n1114, n1115,
    n1116, n1117, n1118, n1119, n1120, n1121,
    n1122, n1123, n1124, n1125, n1126, n1127,
    n1128, n1129, n1130, n1131, n1132, n1133,
    n1134, n1135, n1136, n1137, n1138, n1139,
    n1140, n1141, n1142, n1143, n1144, n1145,
    n1146, n1147, n1148, n1149, n1150, n1151,
    n1152, n1153, n1154, n1155, n1156, n1157,
    n1158, n1159, n1160, n1161, n1162, n1163,
    n1164, n1165, n1166, n1167, n1168, n1169,
    n1170, n1171, n1172, n1173, n1174, n1175,
    n1176, n1177, n1178, n1179, n1180, n1181,
    n1182, n1183, n1184, n1185, n1186, n1187,
    n1188, n1189, n1190, n1191, n1192, n1193,
    n1194, n1195, n1196, n1197, n1198, n1199,
    n1200, n1201, n1202, n1203, n1204, n1205,
    n1206, n1207, n1208, n1209, n1210, n1211,
    n1212, n1213, n1214, n1215, n1216, n1217,
    n1218, n1219, n1220, n1221, n1222, n1223,
    n1224, n1225, n1226, n1227, n1228, n1229,
    n1230, n1231, n1232, n1233, n1234, n1235,
    n1236, n1237, n1238, n1239, n1240, n1241,
    n1242, n1243, n1244, n1245, n1246, n1247,
    n1248, n1249, n1250, n1251, n1252, n1253,
    n1254, n1255, n1256, n1257, n1258, n1259,
    n1260, n1261, n1262, n1263, n1264, n1265,
    n1266, n1267, n1268, n1269, n1270, n1271,
    n1272, n1273, n1274, n1275, n1276, n1277,
    n1278, n1279, n1280, n1281, n1282, n1283,
    n1284, n1285, n1286, n1287, n1288, n1289,
    n1290, n1291, n1292, n1293, n1294, n1295,
    n1296, n1297, n1298, n1299, n1300, n1301,
    n1302, n1303, n1304, n1305, n1306, n1307,
    n1308, n1309, n1310, n1311, n1312, n1313,
    n1314, n1315, n1316, n1317, n1318, n1319,
    n1320, n1321, n1322, n1323, n1324, n1325,
    n1326, n1327, n1328, n1329, n1330, n1331,
    n1332, n1333, n1334, n1335, n1336, n1337,
    n1338, n1339, n1340, n1341, n1342, n1343,
    n1344, n1345, n1346, n1347, n1348, n1349,
    n1350, n1351, n1352, n1353, n1354, n1355,
    n1356, n1357, n1358, n1359, n1360, n1361,
    n1362, n1363, n1364, n1365, n1366, n1367,
    n1368, n1369, n1370, n1371, n1372, n1373,
    n1374, n1375, n1376, n1377, n1378, n1379,
    n1380, n1381, n1382, n1383, n1384, n1385,
    n1386, n1387, n1388, n1389, n1390, n1391,
    n1392, n1393, n1394, n1395, n1396, n1397,
    n1398, n1399, n1400, n1401, n1402, n1403,
    n1404, n1405, n1406, n1407, n1408, n1409,
    n1410, n1411, n1412, n1413, n1414, n1415,
    n1416, n1417, n1418, n1419, n1420, n1421,
    n1422, n1423, n1424, n1425, n1426, n1427,
    n1428, n1429, n1430, n1431, n1432, n1433,
    n1434, n1435, n1436, n1437, n1438, n1439,
    n1440, n1441, n1442, n1443, n1444, n1445,
    n1446, n1447, n1448, n1449, n1450, n1451,
    n1452, n1453, n1454, n1455, n1456, n1457,
    n1458, n1459, n1460, n1461, n1462, n1463,
    n1464, n1465, n1466, n1467, n1468, n1469,
    n1470, n1471, n1472, n1473, n1474, n1475,
    n1476, n1477, n1478, n1479, n1480, n1481,
    n1482, n1483, n1484, n1485, n1486, n1487,
    n1488, n1489, n1490, n1491, n1492, n1493,
    n1494, n1495, n1496, n1497, n1498, n1499,
    n1500, n1501, n1502, n1503, n1504, n1505,
    n1506, n1507, n1508, n1509, n1510, n1511,
    n1512, n1513, n1514, n1515, n1516, n1517,
    n1518, n1519, n1520, n1521, n1522, n1523,
    n1524, n1525, n1526, n1527, n1528, n1529,
    n1530, n1531, n1532, n1533, n1534, n1535,
    n1536, n1537, n1538, n1539, n1540, n1541,
    n1542, n1543, n1544, n1545, n1546, n1547,
    n1548, n1549, n1550, n1551, n1552, n1553,
    n1554, n1555, n1556, n1557, n1558, n1559,
    n1560, n1561, n1562, n1563, n1564, n1565,
    n1566, n1567, n1568, n1569, n1570, n1571,
    n1572, n1573, n1574, n1575, n1576, n1577,
    n1578, n1579, n1580, n1581, n1582, n1583,
    n1584, n1585, n1586, n1587, n1588, n1589,
    n1590, n1591, n1592, n1593, n1594, n1595,
    n1596, n1597, n1598, n1599, n1600, n1601,
    n1602, n1603, n1604, n1605, n1606, n1607,
    n1608, n1609, n1610, n1611, n1612, n1613,
    n1614, n1615, n1616, n1617, n1618, n1619,
    n1620, n1621, n1622, n1623, n1624, n1625,
    n1626, n1627, n1628, n1629, n1630, n1631,
    n1632, n1633, n1634, n1635, n1636, n1637,
    n1638, n1639, n1640, n1641, n1642, n1643,
    n1644, n1645, n1646, n1647, n1648, n1649,
    n1650, n1651, n1652, n1653, n1654, n1655,
    n1656, n1657, n1658, n1659, n1660, n1661,
    n1662, n1663, n1664, n1665, n1666, n1667,
    n1668, n1669, n1670, n1671, n1672, n1673,
    n1674, n1675, n1676, n1677, n1678, n1679,
    n1680, n1681, n1682, n1683, n1684, n1685,
    n1686, n1687, n1688, n1689, n1690, n1691,
    n1692, n1693, n1694, n1695, n1696, n1697,
    n1698, n1699, n1700, n1701, n1702, n1703,
    n1704, n1705, n1706, n1707, n1708, n1709,
    n1710, n1711, n1712, n1713, n1714, n1715,
    n1716, n1717, n1718, n1719, n1720, n1721,
    n1722, n1723, n1724, n1725, n1726, n1727,
    n1728, n1729, n1730, n1731, n1732, n1733,
    n1734, n1735, n1736, n1737, n1738, n1739,
    n1740, n1741, n1742, n1743, n1744, n1745,
    n1746, n1747, n1748, n1749, n1750, n1751,
    n1752, n1753, n1754, n1755, n1756, n1757,
    n1758, n1759, n1760, n1761, n1762, n1763,
    n1764, n1765, n1766, n1767, n1768, n1769,
    n1770, n1771, n1772, n1773, n1774, n1775,
    n1776, n1777, n1778, n1779, n1780, n1781,
    n1782, n1783, n1784, n1785, n1786, n1787,
    n1788, n1789, n1790, n1791, n1792, n1793,
    n1794, n1795, n1796, n1797, n1798, n1799,
    n1800, n1801, n1802, n1803, n1804, n1805,
    n1806, n1807, n1808, n1809, n1810, n1811,
    n1812, n1813, n1814, n1815, n1816, n1817,
    n1818, n1819, n1820, n1821, n1822, n1823,
    n1824, n1825, n1826, n1827, n1828, n1829,
    n1830, n1831, n1832, n1833, n1834, n1835,
    n1836, n1837, n1838, n1839, n1840, n1841,
    n1842, n1843, n1844, n1845, n1846, n1847,
    n1848, n1849, n1850, n1851, n1852, n1853,
    n1854, n1855, n1856, n1857, n1858, n1859,
    n1860, n1861, n1862, n1863, n1864, n1865,
    n1866, n1867, n1868, n1869, n1870, n1871,
    n1872, n1873, n1874, n1875, n1876, n1877,
    n1878, n1879, n1880, n1881, n1882, n1883,
    n1884, n1885, n1886, n1887, n1888, n1889,
    n1890, n1891, n1892, n1893, n1894, n1895,
    n1896, n1897, n1898, n1899, n1900, n1901,
    n1902, n1903, n1904, n1905, n1906, n1907,
    n1908, n1909, n1910, n1911, n1912, n1913,
    n1914, n1915, n1916, n1917, n1918, n1919,
    n1920, n1921, n1922, n1923, n1924, n1925,
    n1926, n1927, n1928, n1929, n1930, n1931,
    n1932, n1933, n1934, n1935, n1936, n1937,
    n1938, n1939, n1940, n1941, n1942, n1943,
    n1944, n1945, n1946, n1947, n1948, n1949,
    n1950, n1951, n1952, n1953, n1954, n1955,
    n1956, n1957, n1958, n1959, n1960, n1961,
    n1962, n1963, n1964, n1965, n1966, n1967,
    n1968, n1969, n1970, n1971, n1972, n1973,
    n1974, n1975, n1976, n1977, n1978, n1979,
    n1980, n1981, n1982, n1983, n1984, n1985,
    n1986, n1987, n1988, n1989, n1990, n1991,
    n1992, n1993, n1994, n1995, n1996, n1997,
    n1998, n1999, n2000, n2001, n2002, n2003,
    n2004, n2005, n2006, n2007, n2008, n2009,
    n2010, n2011, n2012, n2013, n2014, n2015,
    n2016, n2017, n2018, n2019, n2020, n2021,
    n2022, n2023, n2024, n2025, n2026, n2027,
    n2028, n2029, n2030, n2031, n2032, n2033,
    n2034, n2035, n2036, n2037, n2038, n2039,
    n2040, n2041, n2042, n2043, n2044, n2045,
    n2046, n2047, n2048, n2049, n2050, n2051,
    n2052, n2053, n2054, n2055, n2056, n2057,
    n2058, n2059, n2060, n2061, n2062, n2063,
    n2064, n2065, n2066, n2067, n2068, n2069,
    n2070, n2071, n2072, n2073, n2074, n2075,
    n2076, n2077, n2078, n2079, n2080, n2081,
    n2082, n2083, n2084, n2085, n2086, n2087,
    n2088, n2089, n2090, n2091, n2092, n2093,
    n2094, n2095, n2096, n2097, n2098, n2099,
    n2100, n2101, n2102, n2103, n2104, n2105,
    n2106, n2107, n2108, n2109, n2110, n2111,
    n2112, n2113, n2114, n2115, n2116, n2117,
    n2118, n2119, n2120, n2121, n2122, n2123,
    n2124, n2125, n2126, n2127, n2128, n2129,
    n2130, n2131, n2132, n2133, n2134, n2135,
    n2136, n2137, n2138, n2139, n2140, n2141,
    n2142, n2143, n2144, n2145, n2146, n2147,
    n2148, n2149, n2150, n2151, n2152, n2153,
    n2154, n2155, n2156, n2157, n2158, n2159,
    n2160, n2161, n2162, n2163, n2164, n2165,
    n2166, n2167, n2168, n2169, n2170, n2171,
    n2172, n2173, n2174, n2175, n2176, n2177,
    n2178, n2179, n2180, n2181, n2182, n2183,
    n2184, n2185, n2186, n2187, n2188, n2189,
    n2190, n2191, n2192, n2193, n2194, n2195,
    n2196, n2197, n2198, n2199, n2200, n2201,
    n2202, n2203, n2204, n2205, n2206, n2207,
    n2208, n2209, n2210, n2211, n2212, n2213,
    n2214, n2215, n2216, n2217, n2218, n2219,
    n2220, n2221, n2222, n2223, n2224, n2225,
    n2226, n2227, n2228, n2229, n2230, n2231,
    n2232, n2233, n2234, n2235, n2236, n2237,
    n2238, n2239, n2240, n2241, n2242, n2243,
    n2244, n2245, n2246, n2247, n2248, n2249,
    n2250, n2251, n2252, n2253, n2254, n2255,
    n2256, n2257, n2258, n2259, n2260, n2261,
    n2262, n2263, n2264, n2265, n2266, n2267,
    n2268, n2269, n2270, n2271, n2272, n2273,
    n2274, n2275, n2276, n2277, n2278, n2279,
    n2280, n2281, n2282, n2283, n2284, n2285,
    n2286, n2287, n2288, n2289, n2290, n2292,
    n2293, n2295, n2297, n2299, n2301, n2303,
    n2305, n2307, n2309, n2311, n2313, n2315,
    n2317, n2319, n2321, n2323, n2325, n2327,
    n2329, n2331, n2333, n2335, n2337, n2339,
    n2341, n2343, n2345, n2347, n2349, n2351,
    n2353, n2355, n2357, n2359, n2361, n2363,
    n2365, n2367, n2369, n2371, n2373, n2375,
    n2377, n2379, n2381, n2383, n2385, n2387,
    n2389, n2391, n2393, n2395, n2397, n2399,
    n2401, n2403, n2405, n2407, n2409, n2411,
    n2413, n2415, n2417, n2419, n2421, n2423,
    n2425, n2427, n2429, n2431, n2433, n2435,
    n2437, n2439, n2441, n2443, n2445, n2447,
    n2449, n2451, n2453, n2455, n2457, n2459,
    n2461, n2463, n2465, n2467, n2469, n2471,
    n2473, n2475, n2477, n2479, n2481, n2483,
    n2485, n2487, n2489, n2491, n2493, n2495,
    n2497, n2499, n2501, n2503, n2505, n2507,
    n2509, n2511, n2513, n2515, n2517, n2519,
    n2521, n2523, n2525, n2527, n2529, n2531,
    n2533, n2535, n2537, n2539, n2541, n2543;
  assign n386 = ~pi127  & ~pi255 ;
  assign n387 = pi127  & pi255 ;
  assign n388 = ~n386 & ~n387;
  assign n389 = ~pi126  & ~pi254 ;
  assign n390 = pi126  & pi254 ;
  assign n391 = ~pi125  & ~pi253 ;
  assign n392 = pi125  & pi253 ;
  assign n393 = ~pi124  & ~pi252 ;
  assign n394 = pi124  & pi252 ;
  assign n395 = ~pi123  & ~pi251 ;
  assign n396 = pi123  & pi251 ;
  assign n397 = ~pi122  & ~pi250 ;
  assign n398 = pi122  & pi250 ;
  assign n399 = ~pi121  & ~pi249 ;
  assign n400 = pi121  & pi249 ;
  assign n401 = ~pi120  & ~pi248 ;
  assign n402 = pi120  & pi248 ;
  assign n403 = ~pi119  & ~pi247 ;
  assign n404 = pi119  & pi247 ;
  assign n405 = ~pi118  & ~pi246 ;
  assign n406 = pi118  & pi246 ;
  assign n407 = ~pi117  & ~pi245 ;
  assign n408 = pi117  & pi245 ;
  assign n409 = ~pi116  & ~pi244 ;
  assign n410 = pi116  & pi244 ;
  assign n411 = ~pi115  & ~pi243 ;
  assign n412 = pi115  & pi243 ;
  assign n413 = ~pi114  & ~pi242 ;
  assign n414 = pi114  & pi242 ;
  assign n415 = ~pi113  & ~pi241 ;
  assign n416 = pi113  & pi241 ;
  assign n417 = ~pi112  & ~pi240 ;
  assign n418 = pi112  & pi240 ;
  assign n419 = ~pi111  & ~pi239 ;
  assign n420 = pi111  & pi239 ;
  assign n421 = ~pi110  & ~pi238 ;
  assign n422 = pi110  & pi238 ;
  assign n423 = ~pi109  & ~pi237 ;
  assign n424 = pi109  & pi237 ;
  assign n425 = ~pi108  & ~pi236 ;
  assign n426 = pi108  & pi236 ;
  assign n427 = ~pi107  & ~pi235 ;
  assign n428 = pi107  & pi235 ;
  assign n429 = ~pi106  & ~pi234 ;
  assign n430 = pi106  & pi234 ;
  assign n431 = ~pi105  & ~pi233 ;
  assign n432 = pi105  & pi233 ;
  assign n433 = ~pi104  & ~pi232 ;
  assign n434 = pi104  & pi232 ;
  assign n435 = ~pi103  & ~pi231 ;
  assign n436 = pi103  & pi231 ;
  assign n437 = ~pi102  & ~pi230 ;
  assign n438 = pi102  & pi230 ;
  assign n439 = ~pi101  & ~pi229 ;
  assign n440 = pi101  & pi229 ;
  assign n441 = ~pi100  & ~pi228 ;
  assign n442 = pi100  & pi228 ;
  assign n443 = ~pi99  & ~pi227 ;
  assign n444 = pi99  & pi227 ;
  assign n445 = ~pi98  & ~pi226 ;
  assign n446 = pi98  & pi226 ;
  assign n447 = ~pi97  & ~pi225 ;
  assign n448 = pi97  & pi225 ;
  assign n449 = ~pi96  & ~pi224 ;
  assign n450 = pi96  & pi224 ;
  assign n451 = ~pi95  & ~pi223 ;
  assign n452 = pi95  & pi223 ;
  assign n453 = ~pi94  & ~pi222 ;
  assign n454 = pi94  & pi222 ;
  assign n455 = ~pi93  & ~pi221 ;
  assign n456 = pi93  & pi221 ;
  assign n457 = ~pi92  & ~pi220 ;
  assign n458 = pi92  & pi220 ;
  assign n459 = ~pi91  & ~pi219 ;
  assign n460 = pi91  & pi219 ;
  assign n461 = ~pi90  & ~pi218 ;
  assign n462 = pi90  & pi218 ;
  assign n463 = ~pi89  & ~pi217 ;
  assign n464 = pi89  & pi217 ;
  assign n465 = ~pi88  & ~pi216 ;
  assign n466 = pi88  & pi216 ;
  assign n467 = ~pi87  & ~pi215 ;
  assign n468 = pi87  & pi215 ;
  assign n469 = ~pi86  & ~pi214 ;
  assign n470 = pi86  & pi214 ;
  assign n471 = ~pi85  & ~pi213 ;
  assign n472 = pi85  & pi213 ;
  assign n473 = ~pi84  & ~pi212 ;
  assign n474 = pi84  & pi212 ;
  assign n475 = ~pi83  & ~pi211 ;
  assign n476 = pi83  & pi211 ;
  assign n477 = ~pi82  & ~pi210 ;
  assign n478 = pi82  & pi210 ;
  assign n479 = ~pi81  & ~pi209 ;
  assign n480 = pi81  & pi209 ;
  assign n481 = ~pi80  & ~pi208 ;
  assign n482 = pi80  & pi208 ;
  assign n483 = ~pi79  & ~pi207 ;
  assign n484 = pi79  & pi207 ;
  assign n485 = ~pi78  & ~pi206 ;
  assign n486 = pi78  & pi206 ;
  assign n487 = ~pi77  & ~pi205 ;
  assign n488 = pi77  & pi205 ;
  assign n489 = ~pi76  & ~pi204 ;
  assign n490 = pi76  & pi204 ;
  assign n491 = ~pi75  & ~pi203 ;
  assign n492 = pi75  & pi203 ;
  assign n493 = ~pi74  & ~pi202 ;
  assign n494 = pi74  & pi202 ;
  assign n495 = ~pi73  & ~pi201 ;
  assign n496 = pi73  & pi201 ;
  assign n497 = ~pi72  & ~pi200 ;
  assign n498 = pi72  & pi200 ;
  assign n499 = ~pi71  & ~pi199 ;
  assign n500 = pi71  & pi199 ;
  assign n501 = ~pi70  & ~pi198 ;
  assign n502 = pi70  & pi198 ;
  assign n503 = ~pi69  & ~pi197 ;
  assign n504 = pi69  & pi197 ;
  assign n505 = ~pi68  & ~pi196 ;
  assign n506 = pi68  & pi196 ;
  assign n507 = ~pi67  & ~pi195 ;
  assign n508 = pi67  & pi195 ;
  assign n509 = ~pi66  & ~pi194 ;
  assign n510 = pi66  & pi194 ;
  assign n511 = ~pi65  & ~pi193 ;
  assign n512 = pi65  & pi193 ;
  assign n513 = ~pi64  & ~pi192 ;
  assign n514 = pi64  & pi192 ;
  assign n515 = ~pi63  & ~pi191 ;
  assign n516 = pi63  & pi191 ;
  assign n517 = ~pi62  & ~pi190 ;
  assign n518 = pi62  & pi190 ;
  assign n519 = ~pi61  & ~pi189 ;
  assign n520 = pi61  & pi189 ;
  assign n521 = ~pi60  & ~pi188 ;
  assign n522 = pi60  & pi188 ;
  assign n523 = ~pi59  & ~pi187 ;
  assign n524 = pi59  & pi187 ;
  assign n525 = ~pi58  & ~pi186 ;
  assign n526 = pi58  & pi186 ;
  assign n527 = ~pi57  & ~pi185 ;
  assign n528 = pi57  & pi185 ;
  assign n529 = ~pi56  & ~pi184 ;
  assign n530 = pi56  & pi184 ;
  assign n531 = ~pi55  & ~pi183 ;
  assign n532 = pi55  & pi183 ;
  assign n533 = ~pi54  & ~pi182 ;
  assign n534 = pi54  & pi182 ;
  assign n535 = ~pi53  & ~pi181 ;
  assign n536 = pi53  & pi181 ;
  assign n537 = ~pi52  & ~pi180 ;
  assign n538 = pi52  & pi180 ;
  assign n539 = ~pi51  & ~pi179 ;
  assign n540 = pi51  & pi179 ;
  assign n541 = ~pi50  & ~pi178 ;
  assign n542 = pi50  & pi178 ;
  assign n543 = ~pi49  & ~pi177 ;
  assign n544 = pi49  & pi177 ;
  assign n545 = ~pi48  & ~pi176 ;
  assign n546 = pi48  & pi176 ;
  assign n547 = ~pi47  & ~pi175 ;
  assign n548 = pi47  & pi175 ;
  assign n549 = ~pi46  & ~pi174 ;
  assign n550 = pi46  & pi174 ;
  assign n551 = ~pi45  & ~pi173 ;
  assign n552 = pi45  & pi173 ;
  assign n553 = ~pi44  & ~pi172 ;
  assign n554 = pi44  & pi172 ;
  assign n555 = ~pi43  & ~pi171 ;
  assign n556 = pi43  & pi171 ;
  assign n557 = ~pi42  & ~pi170 ;
  assign n558 = pi42  & pi170 ;
  assign n559 = ~pi41  & ~pi169 ;
  assign n560 = pi41  & pi169 ;
  assign n561 = ~pi40  & ~pi168 ;
  assign n562 = pi40  & pi168 ;
  assign n563 = ~pi39  & ~pi167 ;
  assign n564 = pi39  & pi167 ;
  assign n565 = ~pi38  & ~pi166 ;
  assign n566 = pi38  & pi166 ;
  assign n567 = ~pi37  & ~pi165 ;
  assign n568 = pi37  & pi165 ;
  assign n569 = ~pi36  & ~pi164 ;
  assign n570 = pi36  & pi164 ;
  assign n571 = ~pi35  & ~pi163 ;
  assign n572 = pi35  & pi163 ;
  assign n573 = ~pi34  & ~pi162 ;
  assign n574 = pi34  & pi162 ;
  assign n575 = ~pi33  & ~pi161 ;
  assign n576 = pi33  & pi161 ;
  assign n577 = ~pi32  & ~pi160 ;
  assign n578 = pi32  & pi160 ;
  assign n579 = ~pi31  & ~pi159 ;
  assign n580 = pi31  & pi159 ;
  assign n581 = ~pi30  & ~pi158 ;
  assign n582 = pi30  & pi158 ;
  assign n583 = ~pi29  & ~pi157 ;
  assign n584 = pi29  & pi157 ;
  assign n585 = ~pi28  & ~pi156 ;
  assign n586 = pi28  & pi156 ;
  assign n587 = ~pi27  & ~pi155 ;
  assign n588 = pi27  & pi155 ;
  assign n589 = ~pi26  & ~pi154 ;
  assign n590 = pi26  & pi154 ;
  assign n591 = ~pi25  & ~pi153 ;
  assign n592 = pi25  & pi153 ;
  assign n593 = ~pi24  & ~pi152 ;
  assign n594 = pi24  & pi152 ;
  assign n595 = ~pi23  & ~pi151 ;
  assign n596 = pi23  & pi151 ;
  assign n597 = ~pi22  & ~pi150 ;
  assign n598 = pi22  & pi150 ;
  assign n599 = ~pi21  & ~pi149 ;
  assign n600 = pi21  & pi149 ;
  assign n601 = ~pi20  & ~pi148 ;
  assign n602 = pi20  & pi148 ;
  assign n603 = ~pi19  & ~pi147 ;
  assign n604 = pi19  & pi147 ;
  assign n605 = ~pi18  & ~pi146 ;
  assign n606 = pi18  & pi146 ;
  assign n607 = ~pi17  & ~pi145 ;
  assign n608 = pi17  & pi145 ;
  assign n609 = ~pi16  & ~pi144 ;
  assign n610 = pi16  & pi144 ;
  assign n611 = ~pi15  & ~pi143 ;
  assign n612 = pi15  & pi143 ;
  assign n613 = ~pi14  & ~pi142 ;
  assign n614 = pi14  & pi142 ;
  assign n615 = ~pi13  & ~pi141 ;
  assign n616 = pi13  & pi141 ;
  assign n617 = ~pi12  & ~pi140 ;
  assign n618 = pi12  & pi140 ;
  assign n619 = ~pi11  & ~pi139 ;
  assign n620 = pi11  & pi139 ;
  assign n621 = ~pi10  & ~pi138 ;
  assign n622 = pi10  & pi138 ;
  assign n623 = ~pi9  & ~pi137 ;
  assign n624 = pi9  & pi137 ;
  assign n625 = ~pi8  & ~pi136 ;
  assign n626 = pi8  & pi136 ;
  assign n627 = ~pi7  & ~pi135 ;
  assign n628 = pi7  & pi135 ;
  assign n629 = ~pi6  & ~pi134 ;
  assign n630 = pi6  & pi134 ;
  assign n631 = ~pi5  & ~pi133 ;
  assign n632 = pi5  & pi133 ;
  assign n633 = ~pi4  & ~pi132 ;
  assign n634 = pi4  & pi132 ;
  assign n635 = ~pi3  & ~pi131 ;
  assign n636 = pi3  & pi131 ;
  assign n637 = ~pi2  & ~pi130 ;
  assign n638 = pi2  & pi130 ;
  assign n639 = ~pi1  & ~pi129 ;
  assign n640 = pi0  & pi128 ;
  assign n641 = pi1  & pi129 ;
  assign n642 = ~n640 & ~n641;
  assign n643 = ~n639 & n640;
  assign n644 = ~n641 & ~n643;
  assign n645 = ~n639 & ~n642;
  assign n646 = ~n638 & n2165;
  assign n647 = ~n637 & ~n2165;
  assign n648 = ~n638 & ~n647;
  assign n649 = ~n637 & ~n646;
  assign n650 = ~n636 & n2166;
  assign n651 = ~n635 & ~n2166;
  assign n652 = ~n636 & ~n651;
  assign n653 = ~n635 & ~n650;
  assign n654 = ~n634 & n2167;
  assign n655 = ~n633 & ~n2167;
  assign n656 = ~n634 & ~n655;
  assign n657 = ~n633 & ~n654;
  assign n658 = ~n632 & n2168;
  assign n659 = ~n631 & ~n2168;
  assign n660 = ~n632 & ~n659;
  assign n661 = ~n631 & ~n658;
  assign n662 = ~n630 & n2169;
  assign n663 = ~n629 & ~n2169;
  assign n664 = ~n630 & ~n663;
  assign n665 = ~n629 & ~n662;
  assign n666 = ~n628 & n2170;
  assign n667 = ~n627 & ~n2170;
  assign n668 = ~n628 & ~n667;
  assign n669 = ~n627 & ~n666;
  assign n670 = ~n626 & n2171;
  assign n671 = ~n625 & ~n2171;
  assign n672 = ~n626 & ~n671;
  assign n673 = ~n625 & ~n670;
  assign n674 = ~n624 & n2172;
  assign n675 = ~n623 & ~n2172;
  assign n676 = ~n624 & ~n675;
  assign n677 = ~n623 & ~n674;
  assign n678 = ~n622 & n2173;
  assign n679 = ~n621 & ~n2173;
  assign n680 = ~n622 & ~n679;
  assign n681 = ~n621 & ~n678;
  assign n682 = ~n620 & n2174;
  assign n683 = ~n619 & ~n2174;
  assign n684 = ~n620 & ~n683;
  assign n685 = ~n619 & ~n682;
  assign n686 = ~n618 & n2175;
  assign n687 = ~n617 & ~n2175;
  assign n688 = ~n618 & ~n687;
  assign n689 = ~n617 & ~n686;
  assign n690 = ~n616 & n2176;
  assign n691 = ~n615 & ~n2176;
  assign n692 = ~n616 & ~n691;
  assign n693 = ~n615 & ~n690;
  assign n694 = ~n614 & n2177;
  assign n695 = ~n613 & ~n2177;
  assign n696 = ~n614 & ~n695;
  assign n697 = ~n613 & ~n694;
  assign n698 = ~n612 & n2178;
  assign n699 = ~n611 & ~n2178;
  assign n700 = ~n612 & ~n699;
  assign n701 = ~n611 & ~n698;
  assign n702 = ~n610 & n2179;
  assign n703 = ~n609 & ~n2179;
  assign n704 = ~n610 & ~n703;
  assign n705 = ~n609 & ~n702;
  assign n706 = ~n608 & n2180;
  assign n707 = ~n607 & ~n2180;
  assign n708 = ~n608 & ~n707;
  assign n709 = ~n607 & ~n706;
  assign n710 = ~n606 & n2181;
  assign n711 = ~n605 & ~n2181;
  assign n712 = ~n606 & ~n711;
  assign n713 = ~n605 & ~n710;
  assign n714 = ~n604 & n2182;
  assign n715 = ~n603 & ~n2182;
  assign n716 = ~n604 & ~n715;
  assign n717 = ~n603 & ~n714;
  assign n718 = ~n602 & n2183;
  assign n719 = ~n601 & ~n2183;
  assign n720 = ~n602 & ~n719;
  assign n721 = ~n601 & ~n718;
  assign n722 = ~n600 & n2184;
  assign n723 = ~n599 & ~n2184;
  assign n724 = ~n600 & ~n723;
  assign n725 = ~n599 & ~n722;
  assign n726 = ~n598 & n2185;
  assign n727 = ~n597 & ~n2185;
  assign n728 = ~n598 & ~n727;
  assign n729 = ~n597 & ~n726;
  assign n730 = ~n596 & n2186;
  assign n731 = ~n595 & ~n2186;
  assign n732 = ~n596 & ~n731;
  assign n733 = ~n595 & ~n730;
  assign n734 = ~n594 & n2187;
  assign n735 = ~n593 & ~n2187;
  assign n736 = ~n594 & ~n735;
  assign n737 = ~n593 & ~n734;
  assign n738 = ~n592 & n2188;
  assign n739 = ~n591 & ~n2188;
  assign n740 = ~n592 & ~n739;
  assign n741 = ~n591 & ~n738;
  assign n742 = ~n590 & n2189;
  assign n743 = ~n589 & ~n2189;
  assign n744 = ~n590 & ~n743;
  assign n745 = ~n589 & ~n742;
  assign n746 = ~n588 & n2190;
  assign n747 = ~n587 & ~n2190;
  assign n748 = ~n588 & ~n747;
  assign n749 = ~n587 & ~n746;
  assign n750 = ~n586 & n2191;
  assign n751 = ~n585 & ~n2191;
  assign n752 = ~n586 & ~n751;
  assign n753 = ~n585 & ~n750;
  assign n754 = ~n584 & n2192;
  assign n755 = ~n583 & ~n2192;
  assign n756 = ~n584 & ~n755;
  assign n757 = ~n583 & ~n754;
  assign n758 = ~n582 & n2193;
  assign n759 = ~n581 & ~n2193;
  assign n760 = ~n582 & ~n759;
  assign n761 = ~n581 & ~n758;
  assign n762 = ~n580 & n2194;
  assign n763 = ~n579 & ~n2194;
  assign n764 = ~n580 & ~n763;
  assign n765 = ~n579 & ~n762;
  assign n766 = ~n578 & n2195;
  assign n767 = ~n577 & ~n2195;
  assign n768 = ~n578 & ~n767;
  assign n769 = ~n577 & ~n766;
  assign n770 = ~n576 & n2196;
  assign n771 = ~n575 & ~n2196;
  assign n772 = ~n576 & ~n771;
  assign n773 = ~n575 & ~n770;
  assign n774 = ~n574 & n2197;
  assign n775 = ~n573 & ~n2197;
  assign n776 = ~n574 & ~n775;
  assign n777 = ~n573 & ~n774;
  assign n778 = ~n572 & n2198;
  assign n779 = ~n571 & ~n2198;
  assign n780 = ~n572 & ~n779;
  assign n781 = ~n571 & ~n778;
  assign n782 = ~n570 & n2199;
  assign n783 = ~n569 & ~n2199;
  assign n784 = ~n570 & ~n783;
  assign n785 = ~n569 & ~n782;
  assign n786 = ~n568 & n2200;
  assign n787 = ~n567 & ~n2200;
  assign n788 = ~n568 & ~n787;
  assign n789 = ~n567 & ~n786;
  assign n790 = ~n566 & n2201;
  assign n791 = ~n565 & ~n2201;
  assign n792 = ~n566 & ~n791;
  assign n793 = ~n565 & ~n790;
  assign n794 = ~n564 & n2202;
  assign n795 = ~n563 & ~n2202;
  assign n796 = ~n564 & ~n795;
  assign n797 = ~n563 & ~n794;
  assign n798 = ~n562 & n2203;
  assign n799 = ~n561 & ~n2203;
  assign n800 = ~n562 & ~n799;
  assign n801 = ~n561 & ~n798;
  assign n802 = ~n560 & n2204;
  assign n803 = ~n559 & ~n2204;
  assign n804 = ~n560 & ~n803;
  assign n805 = ~n559 & ~n802;
  assign n806 = ~n558 & n2205;
  assign n807 = ~n557 & ~n2205;
  assign n808 = ~n558 & ~n807;
  assign n809 = ~n557 & ~n806;
  assign n810 = ~n556 & n2206;
  assign n811 = ~n555 & ~n2206;
  assign n812 = ~n556 & ~n811;
  assign n813 = ~n555 & ~n810;
  assign n814 = ~n554 & n2207;
  assign n815 = ~n553 & ~n2207;
  assign n816 = ~n554 & ~n815;
  assign n817 = ~n553 & ~n814;
  assign n818 = ~n552 & n2208;
  assign n819 = ~n551 & ~n2208;
  assign n820 = ~n552 & ~n819;
  assign n821 = ~n551 & ~n818;
  assign n822 = ~n550 & n2209;
  assign n823 = ~n549 & ~n2209;
  assign n824 = ~n550 & ~n823;
  assign n825 = ~n549 & ~n822;
  assign n826 = ~n548 & n2210;
  assign n827 = ~n547 & ~n2210;
  assign n828 = ~n548 & ~n827;
  assign n829 = ~n547 & ~n826;
  assign n830 = ~n546 & n2211;
  assign n831 = ~n545 & ~n2211;
  assign n832 = ~n546 & ~n831;
  assign n833 = ~n545 & ~n830;
  assign n834 = ~n544 & n2212;
  assign n835 = ~n543 & ~n2212;
  assign n836 = ~n544 & ~n835;
  assign n837 = ~n543 & ~n834;
  assign n838 = ~n542 & n2213;
  assign n839 = ~n541 & ~n2213;
  assign n840 = ~n542 & ~n839;
  assign n841 = ~n541 & ~n838;
  assign n842 = ~n540 & n2214;
  assign n843 = ~n539 & ~n2214;
  assign n844 = ~n540 & ~n843;
  assign n845 = ~n539 & ~n842;
  assign n846 = ~n538 & n2215;
  assign n847 = ~n537 & ~n2215;
  assign n848 = ~n538 & ~n847;
  assign n849 = ~n537 & ~n846;
  assign n850 = ~n536 & n2216;
  assign n851 = ~n535 & ~n2216;
  assign n852 = ~n536 & ~n851;
  assign n853 = ~n535 & ~n850;
  assign n854 = ~n534 & n2217;
  assign n855 = ~n533 & ~n2217;
  assign n856 = ~n534 & ~n855;
  assign n857 = ~n533 & ~n854;
  assign n858 = ~n532 & n2218;
  assign n859 = ~n531 & ~n2218;
  assign n860 = ~n532 & ~n859;
  assign n861 = ~n531 & ~n858;
  assign n862 = ~n530 & n2219;
  assign n863 = ~n529 & ~n2219;
  assign n864 = ~n530 & ~n863;
  assign n865 = ~n529 & ~n862;
  assign n866 = ~n528 & n2220;
  assign n867 = ~n527 & ~n2220;
  assign n868 = ~n528 & ~n867;
  assign n869 = ~n527 & ~n866;
  assign n870 = ~n526 & n2221;
  assign n871 = ~n525 & ~n2221;
  assign n872 = ~n526 & ~n871;
  assign n873 = ~n525 & ~n870;
  assign n874 = ~n524 & n2222;
  assign n875 = ~n523 & ~n2222;
  assign n876 = ~n524 & ~n875;
  assign n877 = ~n523 & ~n874;
  assign n878 = ~n522 & n2223;
  assign n879 = ~n521 & ~n2223;
  assign n880 = ~n522 & ~n879;
  assign n881 = ~n521 & ~n878;
  assign n882 = ~n520 & n2224;
  assign n883 = ~n519 & ~n2224;
  assign n884 = ~n520 & ~n883;
  assign n885 = ~n519 & ~n882;
  assign n886 = ~n518 & n2225;
  assign n887 = ~n517 & ~n2225;
  assign n888 = ~n518 & ~n887;
  assign n889 = ~n517 & ~n886;
  assign n890 = ~n516 & n2226;
  assign n891 = ~n515 & ~n2226;
  assign n892 = ~n516 & ~n891;
  assign n893 = ~n515 & ~n890;
  assign n894 = ~n514 & n2227;
  assign n895 = ~n513 & ~n2227;
  assign n896 = ~n514 & ~n895;
  assign n897 = ~n513 & ~n894;
  assign n898 = ~n512 & n2228;
  assign n899 = ~n511 & ~n2228;
  assign n900 = ~n512 & ~n899;
  assign n901 = ~n511 & ~n898;
  assign n902 = ~n510 & n2229;
  assign n903 = ~n509 & ~n2229;
  assign n904 = ~n510 & ~n903;
  assign n905 = ~n509 & ~n902;
  assign n906 = ~n508 & n2230;
  assign n907 = ~n507 & ~n2230;
  assign n908 = ~n508 & ~n907;
  assign n909 = ~n507 & ~n906;
  assign n910 = ~n506 & n2231;
  assign n911 = ~n505 & ~n2231;
  assign n912 = ~n506 & ~n911;
  assign n913 = ~n505 & ~n910;
  assign n914 = ~n504 & n2232;
  assign n915 = ~n503 & ~n2232;
  assign n916 = ~n504 & ~n915;
  assign n917 = ~n503 & ~n914;
  assign n918 = ~n502 & n2233;
  assign n919 = ~n501 & ~n2233;
  assign n920 = ~n502 & ~n919;
  assign n921 = ~n501 & ~n918;
  assign n922 = ~n500 & n2234;
  assign n923 = ~n499 & ~n2234;
  assign n924 = ~n500 & ~n923;
  assign n925 = ~n499 & ~n922;
  assign n926 = ~n498 & n2235;
  assign n927 = ~n497 & ~n2235;
  assign n928 = ~n498 & ~n927;
  assign n929 = ~n497 & ~n926;
  assign n930 = ~n496 & n2236;
  assign n931 = ~n495 & ~n2236;
  assign n932 = ~n496 & ~n931;
  assign n933 = ~n495 & ~n930;
  assign n934 = ~n494 & n2237;
  assign n935 = ~n493 & ~n2237;
  assign n936 = ~n494 & ~n935;
  assign n937 = ~n493 & ~n934;
  assign n938 = ~n492 & n2238;
  assign n939 = ~n491 & ~n2238;
  assign n940 = ~n492 & ~n939;
  assign n941 = ~n491 & ~n938;
  assign n942 = ~n490 & n2239;
  assign n943 = ~n489 & ~n2239;
  assign n944 = ~n490 & ~n943;
  assign n945 = ~n489 & ~n942;
  assign n946 = ~n488 & n2240;
  assign n947 = ~n487 & ~n2240;
  assign n948 = ~n488 & ~n947;
  assign n949 = ~n487 & ~n946;
  assign n950 = ~n486 & n2241;
  assign n951 = ~n485 & ~n2241;
  assign n952 = ~n486 & ~n951;
  assign n953 = ~n485 & ~n950;
  assign n954 = ~n484 & n2242;
  assign n955 = ~n483 & ~n2242;
  assign n956 = ~n484 & ~n955;
  assign n957 = ~n483 & ~n954;
  assign n958 = ~n482 & n2243;
  assign n959 = ~n481 & ~n2243;
  assign n960 = ~n482 & ~n959;
  assign n961 = ~n481 & ~n958;
  assign n962 = ~n480 & n2244;
  assign n963 = ~n479 & ~n2244;
  assign n964 = ~n480 & ~n963;
  assign n965 = ~n479 & ~n962;
  assign n966 = ~n478 & n2245;
  assign n967 = ~n477 & ~n2245;
  assign n968 = ~n478 & ~n967;
  assign n969 = ~n477 & ~n966;
  assign n970 = ~n476 & n2246;
  assign n971 = ~n475 & ~n2246;
  assign n972 = ~n476 & ~n971;
  assign n973 = ~n475 & ~n970;
  assign n974 = ~n474 & n2247;
  assign n975 = ~n473 & ~n2247;
  assign n976 = ~n474 & ~n975;
  assign n977 = ~n473 & ~n974;
  assign n978 = ~n472 & n2248;
  assign n979 = ~n471 & ~n2248;
  assign n980 = ~n472 & ~n979;
  assign n981 = ~n471 & ~n978;
  assign n982 = ~n470 & n2249;
  assign n983 = ~n469 & ~n2249;
  assign n984 = ~n470 & ~n983;
  assign n985 = ~n469 & ~n982;
  assign n986 = ~n468 & n2250;
  assign n987 = ~n467 & ~n2250;
  assign n988 = ~n468 & ~n987;
  assign n989 = ~n467 & ~n986;
  assign n990 = ~n466 & n2251;
  assign n991 = ~n465 & ~n2251;
  assign n992 = ~n466 & ~n991;
  assign n993 = ~n465 & ~n990;
  assign n994 = ~n464 & n2252;
  assign n995 = ~n463 & ~n2252;
  assign n996 = ~n464 & ~n995;
  assign n997 = ~n463 & ~n994;
  assign n998 = ~n462 & n2253;
  assign n999 = ~n461 & ~n2253;
  assign n1000 = ~n462 & ~n999;
  assign n1001 = ~n461 & ~n998;
  assign n1002 = ~n460 & n2254;
  assign n1003 = ~n459 & ~n2254;
  assign n1004 = ~n460 & ~n1003;
  assign n1005 = ~n459 & ~n1002;
  assign n1006 = ~n458 & n2255;
  assign n1007 = ~n457 & ~n2255;
  assign n1008 = ~n458 & ~n1007;
  assign n1009 = ~n457 & ~n1006;
  assign n1010 = ~n456 & n2256;
  assign n1011 = ~n455 & ~n2256;
  assign n1012 = ~n456 & ~n1011;
  assign n1013 = ~n455 & ~n1010;
  assign n1014 = ~n454 & n2257;
  assign n1015 = ~n453 & ~n2257;
  assign n1016 = ~n454 & ~n1015;
  assign n1017 = ~n453 & ~n1014;
  assign n1018 = ~n452 & n2258;
  assign n1019 = ~n451 & ~n2258;
  assign n1020 = ~n452 & ~n1019;
  assign n1021 = ~n451 & ~n1018;
  assign n1022 = ~n450 & n2259;
  assign n1023 = ~n449 & ~n2259;
  assign n1024 = ~n450 & ~n1023;
  assign n1025 = ~n449 & ~n1022;
  assign n1026 = ~n448 & n2260;
  assign n1027 = ~n447 & ~n2260;
  assign n1028 = ~n448 & ~n1027;
  assign n1029 = ~n447 & ~n1026;
  assign n1030 = ~n446 & n2261;
  assign n1031 = ~n445 & ~n2261;
  assign n1032 = ~n446 & ~n1031;
  assign n1033 = ~n445 & ~n1030;
  assign n1034 = ~n444 & n2262;
  assign n1035 = ~n443 & ~n2262;
  assign n1036 = ~n444 & ~n1035;
  assign n1037 = ~n443 & ~n1034;
  assign n1038 = ~n442 & n2263;
  assign n1039 = ~n441 & ~n2263;
  assign n1040 = ~n442 & ~n1039;
  assign n1041 = ~n441 & ~n1038;
  assign n1042 = ~n440 & n2264;
  assign n1043 = ~n439 & ~n2264;
  assign n1044 = ~n440 & ~n1043;
  assign n1045 = ~n439 & ~n1042;
  assign n1046 = ~n438 & n2265;
  assign n1047 = ~n437 & ~n2265;
  assign n1048 = ~n438 & ~n1047;
  assign n1049 = ~n437 & ~n1046;
  assign n1050 = ~n436 & n2266;
  assign n1051 = ~n435 & ~n2266;
  assign n1052 = ~n436 & ~n1051;
  assign n1053 = ~n435 & ~n1050;
  assign n1054 = ~n434 & n2267;
  assign n1055 = ~n433 & ~n2267;
  assign n1056 = ~n434 & ~n1055;
  assign n1057 = ~n433 & ~n1054;
  assign n1058 = ~n432 & n2268;
  assign n1059 = ~n431 & ~n2268;
  assign n1060 = ~n432 & ~n1059;
  assign n1061 = ~n431 & ~n1058;
  assign n1062 = ~n430 & n2269;
  assign n1063 = ~n429 & ~n2269;
  assign n1064 = ~n430 & ~n1063;
  assign n1065 = ~n429 & ~n1062;
  assign n1066 = ~n428 & n2270;
  assign n1067 = ~n427 & ~n2270;
  assign n1068 = ~n428 & ~n1067;
  assign n1069 = ~n427 & ~n1066;
  assign n1070 = ~n426 & n2271;
  assign n1071 = ~n425 & ~n2271;
  assign n1072 = ~n426 & ~n1071;
  assign n1073 = ~n425 & ~n1070;
  assign n1074 = ~n424 & n2272;
  assign n1075 = ~n423 & ~n2272;
  assign n1076 = ~n424 & ~n1075;
  assign n1077 = ~n423 & ~n1074;
  assign n1078 = ~n422 & n2273;
  assign n1079 = ~n421 & ~n2273;
  assign n1080 = ~n422 & ~n1079;
  assign n1081 = ~n421 & ~n1078;
  assign n1082 = ~n420 & n2274;
  assign n1083 = ~n419 & ~n2274;
  assign n1084 = ~n420 & ~n1083;
  assign n1085 = ~n419 & ~n1082;
  assign n1086 = ~n418 & n2275;
  assign n1087 = ~n417 & ~n2275;
  assign n1088 = ~n418 & ~n1087;
  assign n1089 = ~n417 & ~n1086;
  assign n1090 = ~n416 & n2276;
  assign n1091 = ~n415 & ~n2276;
  assign n1092 = ~n416 & ~n1091;
  assign n1093 = ~n415 & ~n1090;
  assign n1094 = ~n414 & n2277;
  assign n1095 = ~n413 & ~n2277;
  assign n1096 = ~n414 & ~n1095;
  assign n1097 = ~n413 & ~n1094;
  assign n1098 = ~n412 & n2278;
  assign n1099 = ~n411 & ~n2278;
  assign n1100 = ~n412 & ~n1099;
  assign n1101 = ~n411 & ~n1098;
  assign n1102 = ~n410 & n2279;
  assign n1103 = ~n409 & ~n2279;
  assign n1104 = ~n410 & ~n1103;
  assign n1105 = ~n409 & ~n1102;
  assign n1106 = ~n408 & n2280;
  assign n1107 = ~n407 & ~n2280;
  assign n1108 = ~n408 & ~n1107;
  assign n1109 = ~n407 & ~n1106;
  assign n1110 = ~n406 & n2281;
  assign n1111 = ~n405 & ~n2281;
  assign n1112 = ~n406 & ~n1111;
  assign n1113 = ~n405 & ~n1110;
  assign n1114 = ~n404 & n2282;
  assign n1115 = ~n403 & ~n2282;
  assign n1116 = ~n404 & ~n1115;
  assign n1117 = ~n403 & ~n1114;
  assign n1118 = ~n402 & n2283;
  assign n1119 = ~n401 & ~n2283;
  assign n1120 = ~n402 & ~n1119;
  assign n1121 = ~n401 & ~n1118;
  assign n1122 = ~n400 & n2284;
  assign n1123 = ~n399 & ~n2284;
  assign n1124 = ~n400 & ~n1123;
  assign n1125 = ~n399 & ~n1122;
  assign n1126 = ~n398 & n2285;
  assign n1127 = ~n397 & ~n2285;
  assign n1128 = ~n398 & ~n1127;
  assign n1129 = ~n397 & ~n1126;
  assign n1130 = ~n396 & n2286;
  assign n1131 = ~n395 & ~n2286;
  assign n1132 = ~n396 & ~n1131;
  assign n1133 = ~n395 & ~n1130;
  assign n1134 = ~n394 & n2287;
  assign n1135 = ~n393 & ~n2287;
  assign n1136 = ~n394 & ~n1135;
  assign n1137 = ~n393 & ~n1134;
  assign n1138 = ~n392 & n2288;
  assign n1139 = ~n391 & ~n2288;
  assign n1140 = ~n392 & ~n1139;
  assign n1141 = ~n391 & ~n1138;
  assign n1142 = ~n390 & n2289;
  assign n1143 = ~n389 & ~n2289;
  assign n1144 = ~n390 & ~n1143;
  assign n1145 = ~n389 & ~n1142;
  assign n1146 = n388 & n2290;
  assign n1147 = ~n388 & ~n2290;
  assign n1148 = ~n388 & n2290;
  assign n1149 = n388 & ~n2290;
  assign n1150 = ~n1148 & ~n1149;
  assign n1151 = ~n1146 & ~n1147;
  assign n1152 = ~n387 & n2290;
  assign n1153 = ~n386 & ~n2290;
  assign n1154 = ~n387 & ~n1153;
  assign n1155 = ~n386 & ~n1152;
  assign n1156 = ~n389 & ~n390;
  assign n1157 = ~n2289 & ~n1156;
  assign n1158 = ~n389 & n1142;
  assign n1159 = n2289 & n1156;
  assign n1160 = n2289 & ~n1156;
  assign n1161 = ~n2289 & n1156;
  assign n1162 = ~n1160 & ~n1161;
  assign n1163 = ~n1157 & ~n2293;
  assign n1164 = ~n391 & ~n392;
  assign n1165 = ~n2288 & ~n1164;
  assign n1166 = ~n391 & n1138;
  assign n1167 = n2288 & n1164;
  assign n1168 = n2288 & ~n1164;
  assign n1169 = ~n2288 & n1164;
  assign n1170 = ~n1168 & ~n1169;
  assign n1171 = ~n1165 & ~n2295;
  assign n1172 = ~n393 & ~n394;
  assign n1173 = ~n2287 & ~n1172;
  assign n1174 = ~n393 & n1134;
  assign n1175 = n2287 & n1172;
  assign n1176 = n2287 & ~n1172;
  assign n1177 = ~n2287 & n1172;
  assign n1178 = ~n1176 & ~n1177;
  assign n1179 = ~n1173 & ~n2297;
  assign n1180 = ~n395 & ~n396;
  assign n1181 = ~n2286 & ~n1180;
  assign n1182 = ~n395 & n1130;
  assign n1183 = n2286 & n1180;
  assign n1184 = n2286 & ~n1180;
  assign n1185 = ~n2286 & n1180;
  assign n1186 = ~n1184 & ~n1185;
  assign n1187 = ~n1181 & ~n2299;
  assign n1188 = ~n397 & ~n398;
  assign n1189 = ~n2285 & ~n1188;
  assign n1190 = ~n397 & n1126;
  assign n1191 = n2285 & n1188;
  assign n1192 = n2285 & ~n1188;
  assign n1193 = ~n2285 & n1188;
  assign n1194 = ~n1192 & ~n1193;
  assign n1195 = ~n1189 & ~n2301;
  assign n1196 = ~n399 & ~n400;
  assign n1197 = ~n2284 & ~n1196;
  assign n1198 = ~n399 & n1122;
  assign n1199 = n2284 & n1196;
  assign n1200 = n2284 & ~n1196;
  assign n1201 = ~n2284 & n1196;
  assign n1202 = ~n1200 & ~n1201;
  assign n1203 = ~n1197 & ~n2303;
  assign n1204 = ~n401 & ~n402;
  assign n1205 = ~n2283 & ~n1204;
  assign n1206 = ~n401 & n1118;
  assign n1207 = n2283 & n1204;
  assign n1208 = n2283 & ~n1204;
  assign n1209 = ~n2283 & n1204;
  assign n1210 = ~n1208 & ~n1209;
  assign n1211 = ~n1205 & ~n2305;
  assign n1212 = ~n403 & ~n404;
  assign n1213 = ~n2282 & ~n1212;
  assign n1214 = ~n403 & n1114;
  assign n1215 = n2282 & n1212;
  assign n1216 = n2282 & ~n1212;
  assign n1217 = ~n2282 & n1212;
  assign n1218 = ~n1216 & ~n1217;
  assign n1219 = ~n1213 & ~n2307;
  assign n1220 = ~n405 & ~n406;
  assign n1221 = ~n2281 & ~n1220;
  assign n1222 = ~n405 & n1110;
  assign n1223 = n2281 & n1220;
  assign n1224 = n2281 & ~n1220;
  assign n1225 = ~n2281 & n1220;
  assign n1226 = ~n1224 & ~n1225;
  assign n1227 = ~n1221 & ~n2309;
  assign n1228 = ~n407 & ~n408;
  assign n1229 = ~n2280 & ~n1228;
  assign n1230 = ~n407 & n1106;
  assign n1231 = n2280 & n1228;
  assign n1232 = n2280 & ~n1228;
  assign n1233 = ~n2280 & n1228;
  assign n1234 = ~n1232 & ~n1233;
  assign n1235 = ~n1229 & ~n2311;
  assign n1236 = ~n409 & ~n410;
  assign n1237 = ~n2279 & ~n1236;
  assign n1238 = ~n409 & n1102;
  assign n1239 = n2279 & n1236;
  assign n1240 = n2279 & ~n1236;
  assign n1241 = ~n2279 & n1236;
  assign n1242 = ~n1240 & ~n1241;
  assign n1243 = ~n1237 & ~n2313;
  assign n1244 = ~n411 & ~n412;
  assign n1245 = ~n2278 & ~n1244;
  assign n1246 = ~n411 & n1098;
  assign n1247 = n2278 & n1244;
  assign n1248 = n2278 & ~n1244;
  assign n1249 = ~n2278 & n1244;
  assign n1250 = ~n1248 & ~n1249;
  assign n1251 = ~n1245 & ~n2315;
  assign n1252 = ~n413 & ~n414;
  assign n1253 = ~n2277 & ~n1252;
  assign n1254 = ~n413 & n1094;
  assign n1255 = n2277 & n1252;
  assign n1256 = n2277 & ~n1252;
  assign n1257 = ~n2277 & n1252;
  assign n1258 = ~n1256 & ~n1257;
  assign n1259 = ~n1253 & ~n2317;
  assign n1260 = ~n415 & ~n416;
  assign n1261 = ~n2276 & ~n1260;
  assign n1262 = ~n415 & n1090;
  assign n1263 = n2276 & n1260;
  assign n1264 = n2276 & ~n1260;
  assign n1265 = ~n2276 & n1260;
  assign n1266 = ~n1264 & ~n1265;
  assign n1267 = ~n1261 & ~n2319;
  assign n1268 = ~n417 & ~n418;
  assign n1269 = ~n2275 & ~n1268;
  assign n1270 = ~n417 & n1086;
  assign n1271 = n2275 & n1268;
  assign n1272 = n2275 & ~n1268;
  assign n1273 = ~n2275 & n1268;
  assign n1274 = ~n1272 & ~n1273;
  assign n1275 = ~n1269 & ~n2321;
  assign n1276 = ~n419 & ~n420;
  assign n1277 = ~n2274 & ~n1276;
  assign n1278 = ~n419 & n1082;
  assign n1279 = n2274 & n1276;
  assign n1280 = n2274 & ~n1276;
  assign n1281 = ~n2274 & n1276;
  assign n1282 = ~n1280 & ~n1281;
  assign n1283 = ~n1277 & ~n2323;
  assign n1284 = ~n421 & ~n422;
  assign n1285 = ~n2273 & ~n1284;
  assign n1286 = ~n421 & n1078;
  assign n1287 = n2273 & n1284;
  assign n1288 = n2273 & ~n1284;
  assign n1289 = ~n2273 & n1284;
  assign n1290 = ~n1288 & ~n1289;
  assign n1291 = ~n1285 & ~n2325;
  assign n1292 = ~n423 & ~n424;
  assign n1293 = ~n2272 & ~n1292;
  assign n1294 = ~n423 & n1074;
  assign n1295 = n2272 & n1292;
  assign n1296 = n2272 & ~n1292;
  assign n1297 = ~n2272 & n1292;
  assign n1298 = ~n1296 & ~n1297;
  assign n1299 = ~n1293 & ~n2327;
  assign n1300 = ~n425 & ~n426;
  assign n1301 = ~n2271 & ~n1300;
  assign n1302 = ~n425 & n1070;
  assign n1303 = n2271 & n1300;
  assign n1304 = n2271 & ~n1300;
  assign n1305 = ~n2271 & n1300;
  assign n1306 = ~n1304 & ~n1305;
  assign n1307 = ~n1301 & ~n2329;
  assign n1308 = ~n427 & ~n428;
  assign n1309 = ~n2270 & ~n1308;
  assign n1310 = ~n427 & n1066;
  assign n1311 = n2270 & n1308;
  assign n1312 = n2270 & ~n1308;
  assign n1313 = ~n2270 & n1308;
  assign n1314 = ~n1312 & ~n1313;
  assign n1315 = ~n1309 & ~n2331;
  assign n1316 = ~n429 & ~n430;
  assign n1317 = ~n2269 & ~n1316;
  assign n1318 = ~n429 & n1062;
  assign n1319 = n2269 & n1316;
  assign n1320 = n2269 & ~n1316;
  assign n1321 = ~n2269 & n1316;
  assign n1322 = ~n1320 & ~n1321;
  assign n1323 = ~n1317 & ~n2333;
  assign n1324 = ~n431 & ~n432;
  assign n1325 = ~n2268 & ~n1324;
  assign n1326 = ~n431 & n1058;
  assign n1327 = n2268 & n1324;
  assign n1328 = n2268 & ~n1324;
  assign n1329 = ~n2268 & n1324;
  assign n1330 = ~n1328 & ~n1329;
  assign n1331 = ~n1325 & ~n2335;
  assign n1332 = ~n433 & ~n434;
  assign n1333 = ~n2267 & ~n1332;
  assign n1334 = ~n433 & n1054;
  assign n1335 = n2267 & n1332;
  assign n1336 = n2267 & ~n1332;
  assign n1337 = ~n2267 & n1332;
  assign n1338 = ~n1336 & ~n1337;
  assign n1339 = ~n1333 & ~n2337;
  assign n1340 = ~n435 & ~n436;
  assign n1341 = ~n2266 & ~n1340;
  assign n1342 = ~n435 & n1050;
  assign n1343 = n2266 & n1340;
  assign n1344 = n2266 & ~n1340;
  assign n1345 = ~n2266 & n1340;
  assign n1346 = ~n1344 & ~n1345;
  assign n1347 = ~n1341 & ~n2339;
  assign n1348 = ~n437 & ~n438;
  assign n1349 = ~n2265 & ~n1348;
  assign n1350 = ~n437 & n1046;
  assign n1351 = n2265 & n1348;
  assign n1352 = n2265 & ~n1348;
  assign n1353 = ~n2265 & n1348;
  assign n1354 = ~n1352 & ~n1353;
  assign n1355 = ~n1349 & ~n2341;
  assign n1356 = ~n439 & ~n440;
  assign n1357 = ~n2264 & ~n1356;
  assign n1358 = ~n439 & n1042;
  assign n1359 = n2264 & n1356;
  assign n1360 = n2264 & ~n1356;
  assign n1361 = ~n2264 & n1356;
  assign n1362 = ~n1360 & ~n1361;
  assign n1363 = ~n1357 & ~n2343;
  assign n1364 = ~n441 & ~n442;
  assign n1365 = ~n2263 & ~n1364;
  assign n1366 = ~n441 & n1038;
  assign n1367 = n2263 & n1364;
  assign n1368 = n2263 & ~n1364;
  assign n1369 = ~n2263 & n1364;
  assign n1370 = ~n1368 & ~n1369;
  assign n1371 = ~n1365 & ~n2345;
  assign n1372 = ~n443 & ~n444;
  assign n1373 = ~n2262 & ~n1372;
  assign n1374 = ~n443 & n1034;
  assign n1375 = n2262 & n1372;
  assign n1376 = n2262 & ~n1372;
  assign n1377 = ~n2262 & n1372;
  assign n1378 = ~n1376 & ~n1377;
  assign n1379 = ~n1373 & ~n2347;
  assign n1380 = ~n445 & ~n446;
  assign n1381 = ~n2261 & ~n1380;
  assign n1382 = ~n445 & n1030;
  assign n1383 = n2261 & n1380;
  assign n1384 = n2261 & ~n1380;
  assign n1385 = ~n2261 & n1380;
  assign n1386 = ~n1384 & ~n1385;
  assign n1387 = ~n1381 & ~n2349;
  assign n1388 = ~n447 & ~n448;
  assign n1389 = ~n2260 & ~n1388;
  assign n1390 = ~n447 & n1026;
  assign n1391 = n2260 & n1388;
  assign n1392 = n2260 & ~n1388;
  assign n1393 = ~n2260 & n1388;
  assign n1394 = ~n1392 & ~n1393;
  assign n1395 = ~n1389 & ~n2351;
  assign n1396 = ~n449 & ~n450;
  assign n1397 = ~n2259 & ~n1396;
  assign n1398 = ~n449 & n1022;
  assign n1399 = n2259 & n1396;
  assign n1400 = n2259 & ~n1396;
  assign n1401 = ~n2259 & n1396;
  assign n1402 = ~n1400 & ~n1401;
  assign n1403 = ~n1397 & ~n2353;
  assign n1404 = ~n451 & ~n452;
  assign n1405 = ~n2258 & ~n1404;
  assign n1406 = ~n451 & n1018;
  assign n1407 = n2258 & n1404;
  assign n1408 = n2258 & ~n1404;
  assign n1409 = ~n2258 & n1404;
  assign n1410 = ~n1408 & ~n1409;
  assign n1411 = ~n1405 & ~n2355;
  assign n1412 = ~n453 & ~n454;
  assign n1413 = ~n2257 & ~n1412;
  assign n1414 = ~n453 & n1014;
  assign n1415 = n2257 & n1412;
  assign n1416 = n2257 & ~n1412;
  assign n1417 = ~n2257 & n1412;
  assign n1418 = ~n1416 & ~n1417;
  assign n1419 = ~n1413 & ~n2357;
  assign n1420 = ~n455 & ~n456;
  assign n1421 = ~n2256 & ~n1420;
  assign n1422 = ~n455 & n1010;
  assign n1423 = n2256 & n1420;
  assign n1424 = n2256 & ~n1420;
  assign n1425 = ~n2256 & n1420;
  assign n1426 = ~n1424 & ~n1425;
  assign n1427 = ~n1421 & ~n2359;
  assign n1428 = ~n457 & ~n458;
  assign n1429 = ~n2255 & ~n1428;
  assign n1430 = ~n457 & n1006;
  assign n1431 = n2255 & n1428;
  assign n1432 = n2255 & ~n1428;
  assign n1433 = ~n2255 & n1428;
  assign n1434 = ~n1432 & ~n1433;
  assign n1435 = ~n1429 & ~n2361;
  assign n1436 = ~n459 & ~n460;
  assign n1437 = ~n2254 & ~n1436;
  assign n1438 = ~n459 & n1002;
  assign n1439 = n2254 & n1436;
  assign n1440 = n2254 & ~n1436;
  assign n1441 = ~n2254 & n1436;
  assign n1442 = ~n1440 & ~n1441;
  assign n1443 = ~n1437 & ~n2363;
  assign n1444 = ~n461 & ~n462;
  assign n1445 = ~n2253 & ~n1444;
  assign n1446 = ~n461 & n998;
  assign n1447 = n2253 & n1444;
  assign n1448 = n2253 & ~n1444;
  assign n1449 = ~n2253 & n1444;
  assign n1450 = ~n1448 & ~n1449;
  assign n1451 = ~n1445 & ~n2365;
  assign n1452 = ~n463 & ~n464;
  assign n1453 = ~n2252 & ~n1452;
  assign n1454 = ~n463 & n994;
  assign n1455 = n2252 & n1452;
  assign n1456 = n2252 & ~n1452;
  assign n1457 = ~n2252 & n1452;
  assign n1458 = ~n1456 & ~n1457;
  assign n1459 = ~n1453 & ~n2367;
  assign n1460 = ~n465 & ~n466;
  assign n1461 = ~n2251 & ~n1460;
  assign n1462 = ~n465 & n990;
  assign n1463 = n2251 & n1460;
  assign n1464 = n2251 & ~n1460;
  assign n1465 = ~n2251 & n1460;
  assign n1466 = ~n1464 & ~n1465;
  assign n1467 = ~n1461 & ~n2369;
  assign n1468 = ~n467 & ~n468;
  assign n1469 = ~n2250 & ~n1468;
  assign n1470 = ~n467 & n986;
  assign n1471 = n2250 & n1468;
  assign n1472 = n2250 & ~n1468;
  assign n1473 = ~n2250 & n1468;
  assign n1474 = ~n1472 & ~n1473;
  assign n1475 = ~n1469 & ~n2371;
  assign n1476 = ~n469 & ~n470;
  assign n1477 = ~n2249 & ~n1476;
  assign n1478 = ~n469 & n982;
  assign n1479 = n2249 & n1476;
  assign n1480 = n2249 & ~n1476;
  assign n1481 = ~n2249 & n1476;
  assign n1482 = ~n1480 & ~n1481;
  assign n1483 = ~n1477 & ~n2373;
  assign n1484 = ~n471 & ~n472;
  assign n1485 = ~n2248 & ~n1484;
  assign n1486 = ~n471 & n978;
  assign n1487 = n2248 & n1484;
  assign n1488 = n2248 & ~n1484;
  assign n1489 = ~n2248 & n1484;
  assign n1490 = ~n1488 & ~n1489;
  assign n1491 = ~n1485 & ~n2375;
  assign n1492 = ~n473 & ~n474;
  assign n1493 = ~n2247 & ~n1492;
  assign n1494 = ~n473 & n974;
  assign n1495 = n2247 & n1492;
  assign n1496 = n2247 & ~n1492;
  assign n1497 = ~n2247 & n1492;
  assign n1498 = ~n1496 & ~n1497;
  assign n1499 = ~n1493 & ~n2377;
  assign n1500 = ~n475 & ~n476;
  assign n1501 = ~n2246 & ~n1500;
  assign n1502 = ~n475 & n970;
  assign n1503 = n2246 & n1500;
  assign n1504 = n2246 & ~n1500;
  assign n1505 = ~n2246 & n1500;
  assign n1506 = ~n1504 & ~n1505;
  assign n1507 = ~n1501 & ~n2379;
  assign n1508 = ~n477 & ~n478;
  assign n1509 = ~n2245 & ~n1508;
  assign n1510 = ~n477 & n966;
  assign n1511 = n2245 & n1508;
  assign n1512 = n2245 & ~n1508;
  assign n1513 = ~n2245 & n1508;
  assign n1514 = ~n1512 & ~n1513;
  assign n1515 = ~n1509 & ~n2381;
  assign n1516 = ~n479 & ~n480;
  assign n1517 = ~n2244 & ~n1516;
  assign n1518 = ~n479 & n962;
  assign n1519 = n2244 & n1516;
  assign n1520 = n2244 & ~n1516;
  assign n1521 = ~n2244 & n1516;
  assign n1522 = ~n1520 & ~n1521;
  assign n1523 = ~n1517 & ~n2383;
  assign n1524 = ~n481 & ~n482;
  assign n1525 = ~n2243 & ~n1524;
  assign n1526 = ~n481 & n958;
  assign n1527 = n2243 & n1524;
  assign n1528 = n2243 & ~n1524;
  assign n1529 = ~n2243 & n1524;
  assign n1530 = ~n1528 & ~n1529;
  assign n1531 = ~n1525 & ~n2385;
  assign n1532 = ~n483 & ~n484;
  assign n1533 = ~n2242 & ~n1532;
  assign n1534 = ~n483 & n954;
  assign n1535 = n2242 & n1532;
  assign n1536 = n2242 & ~n1532;
  assign n1537 = ~n2242 & n1532;
  assign n1538 = ~n1536 & ~n1537;
  assign n1539 = ~n1533 & ~n2387;
  assign n1540 = ~n485 & ~n486;
  assign n1541 = ~n2241 & ~n1540;
  assign n1542 = ~n485 & n950;
  assign n1543 = n2241 & n1540;
  assign n1544 = n2241 & ~n1540;
  assign n1545 = ~n2241 & n1540;
  assign n1546 = ~n1544 & ~n1545;
  assign n1547 = ~n1541 & ~n2389;
  assign n1548 = ~n487 & ~n488;
  assign n1549 = ~n2240 & ~n1548;
  assign n1550 = ~n487 & n946;
  assign n1551 = n2240 & n1548;
  assign n1552 = n2240 & ~n1548;
  assign n1553 = ~n2240 & n1548;
  assign n1554 = ~n1552 & ~n1553;
  assign n1555 = ~n1549 & ~n2391;
  assign n1556 = ~n489 & ~n490;
  assign n1557 = ~n2239 & ~n1556;
  assign n1558 = ~n489 & n942;
  assign n1559 = n2239 & n1556;
  assign n1560 = n2239 & ~n1556;
  assign n1561 = ~n2239 & n1556;
  assign n1562 = ~n1560 & ~n1561;
  assign n1563 = ~n1557 & ~n2393;
  assign n1564 = ~n491 & ~n492;
  assign n1565 = ~n2238 & ~n1564;
  assign n1566 = ~n491 & n938;
  assign n1567 = n2238 & n1564;
  assign n1568 = n2238 & ~n1564;
  assign n1569 = ~n2238 & n1564;
  assign n1570 = ~n1568 & ~n1569;
  assign n1571 = ~n1565 & ~n2395;
  assign n1572 = ~n493 & ~n494;
  assign n1573 = ~n2237 & ~n1572;
  assign n1574 = ~n493 & n934;
  assign n1575 = n2237 & n1572;
  assign n1576 = n2237 & ~n1572;
  assign n1577 = ~n2237 & n1572;
  assign n1578 = ~n1576 & ~n1577;
  assign n1579 = ~n1573 & ~n2397;
  assign n1580 = ~n495 & ~n496;
  assign n1581 = ~n2236 & ~n1580;
  assign n1582 = ~n495 & n930;
  assign n1583 = n2236 & n1580;
  assign n1584 = n2236 & ~n1580;
  assign n1585 = ~n2236 & n1580;
  assign n1586 = ~n1584 & ~n1585;
  assign n1587 = ~n1581 & ~n2399;
  assign n1588 = ~n497 & ~n498;
  assign n1589 = ~n2235 & ~n1588;
  assign n1590 = ~n497 & n926;
  assign n1591 = n2235 & n1588;
  assign n1592 = n2235 & ~n1588;
  assign n1593 = ~n2235 & n1588;
  assign n1594 = ~n1592 & ~n1593;
  assign n1595 = ~n1589 & ~n2401;
  assign n1596 = ~n499 & ~n500;
  assign n1597 = ~n2234 & ~n1596;
  assign n1598 = ~n499 & n922;
  assign n1599 = n2234 & n1596;
  assign n1600 = n2234 & ~n1596;
  assign n1601 = ~n2234 & n1596;
  assign n1602 = ~n1600 & ~n1601;
  assign n1603 = ~n1597 & ~n2403;
  assign n1604 = ~n501 & ~n502;
  assign n1605 = ~n2233 & ~n1604;
  assign n1606 = ~n501 & n918;
  assign n1607 = n2233 & n1604;
  assign n1608 = n2233 & ~n1604;
  assign n1609 = ~n2233 & n1604;
  assign n1610 = ~n1608 & ~n1609;
  assign n1611 = ~n1605 & ~n2405;
  assign n1612 = ~n503 & ~n504;
  assign n1613 = ~n2232 & ~n1612;
  assign n1614 = ~n503 & n914;
  assign n1615 = n2232 & n1612;
  assign n1616 = n2232 & ~n1612;
  assign n1617 = ~n2232 & n1612;
  assign n1618 = ~n1616 & ~n1617;
  assign n1619 = ~n1613 & ~n2407;
  assign n1620 = ~n505 & ~n506;
  assign n1621 = ~n2231 & ~n1620;
  assign n1622 = ~n505 & n910;
  assign n1623 = n2231 & n1620;
  assign n1624 = n2231 & ~n1620;
  assign n1625 = ~n2231 & n1620;
  assign n1626 = ~n1624 & ~n1625;
  assign n1627 = ~n1621 & ~n2409;
  assign n1628 = ~n507 & ~n508;
  assign n1629 = ~n2230 & ~n1628;
  assign n1630 = ~n507 & n906;
  assign n1631 = n2230 & n1628;
  assign n1632 = n2230 & ~n1628;
  assign n1633 = ~n2230 & n1628;
  assign n1634 = ~n1632 & ~n1633;
  assign n1635 = ~n1629 & ~n2411;
  assign n1636 = ~n509 & ~n510;
  assign n1637 = ~n2229 & ~n1636;
  assign n1638 = ~n509 & n902;
  assign n1639 = n2229 & n1636;
  assign n1640 = n2229 & ~n1636;
  assign n1641 = ~n2229 & n1636;
  assign n1642 = ~n1640 & ~n1641;
  assign n1643 = ~n1637 & ~n2413;
  assign n1644 = ~n511 & ~n512;
  assign n1645 = ~n2228 & ~n1644;
  assign n1646 = ~n511 & n898;
  assign n1647 = n2228 & n1644;
  assign n1648 = n2228 & ~n1644;
  assign n1649 = ~n2228 & n1644;
  assign n1650 = ~n1648 & ~n1649;
  assign n1651 = ~n1645 & ~n2415;
  assign n1652 = ~n513 & ~n514;
  assign n1653 = ~n2227 & ~n1652;
  assign n1654 = ~n513 & n894;
  assign n1655 = n2227 & n1652;
  assign n1656 = n2227 & ~n1652;
  assign n1657 = ~n2227 & n1652;
  assign n1658 = ~n1656 & ~n1657;
  assign n1659 = ~n1653 & ~n2417;
  assign n1660 = ~n515 & ~n516;
  assign n1661 = ~n2226 & ~n1660;
  assign n1662 = ~n515 & n890;
  assign n1663 = n2226 & n1660;
  assign n1664 = n2226 & ~n1660;
  assign n1665 = ~n2226 & n1660;
  assign n1666 = ~n1664 & ~n1665;
  assign n1667 = ~n1661 & ~n2419;
  assign n1668 = ~n517 & ~n518;
  assign n1669 = ~n2225 & ~n1668;
  assign n1670 = ~n517 & n886;
  assign n1671 = n2225 & n1668;
  assign n1672 = n2225 & ~n1668;
  assign n1673 = ~n2225 & n1668;
  assign n1674 = ~n1672 & ~n1673;
  assign n1675 = ~n1669 & ~n2421;
  assign n1676 = ~n519 & ~n520;
  assign n1677 = ~n2224 & ~n1676;
  assign n1678 = ~n519 & n882;
  assign n1679 = n2224 & n1676;
  assign n1680 = n2224 & ~n1676;
  assign n1681 = ~n2224 & n1676;
  assign n1682 = ~n1680 & ~n1681;
  assign n1683 = ~n1677 & ~n2423;
  assign n1684 = ~n521 & ~n522;
  assign n1685 = ~n2223 & ~n1684;
  assign n1686 = ~n521 & n878;
  assign n1687 = n2223 & n1684;
  assign n1688 = n2223 & ~n1684;
  assign n1689 = ~n2223 & n1684;
  assign n1690 = ~n1688 & ~n1689;
  assign n1691 = ~n1685 & ~n2425;
  assign n1692 = ~n523 & ~n524;
  assign n1693 = ~n2222 & ~n1692;
  assign n1694 = ~n523 & n874;
  assign n1695 = n2222 & n1692;
  assign n1696 = n2222 & ~n1692;
  assign n1697 = ~n2222 & n1692;
  assign n1698 = ~n1696 & ~n1697;
  assign n1699 = ~n1693 & ~n2427;
  assign n1700 = ~n525 & ~n526;
  assign n1701 = ~n2221 & ~n1700;
  assign n1702 = ~n525 & n870;
  assign n1703 = n2221 & n1700;
  assign n1704 = n2221 & ~n1700;
  assign n1705 = ~n2221 & n1700;
  assign n1706 = ~n1704 & ~n1705;
  assign n1707 = ~n1701 & ~n2429;
  assign n1708 = ~n527 & ~n528;
  assign n1709 = ~n2220 & ~n1708;
  assign n1710 = ~n527 & n866;
  assign n1711 = n2220 & n1708;
  assign n1712 = n2220 & ~n1708;
  assign n1713 = ~n2220 & n1708;
  assign n1714 = ~n1712 & ~n1713;
  assign n1715 = ~n1709 & ~n2431;
  assign n1716 = ~n529 & ~n530;
  assign n1717 = ~n2219 & ~n1716;
  assign n1718 = ~n529 & n862;
  assign n1719 = n2219 & n1716;
  assign n1720 = n2219 & ~n1716;
  assign n1721 = ~n2219 & n1716;
  assign n1722 = ~n1720 & ~n1721;
  assign n1723 = ~n1717 & ~n2433;
  assign n1724 = ~n531 & ~n532;
  assign n1725 = ~n2218 & ~n1724;
  assign n1726 = ~n531 & n858;
  assign n1727 = n2218 & n1724;
  assign n1728 = n2218 & ~n1724;
  assign n1729 = ~n2218 & n1724;
  assign n1730 = ~n1728 & ~n1729;
  assign n1731 = ~n1725 & ~n2435;
  assign n1732 = ~n533 & ~n534;
  assign n1733 = ~n2217 & ~n1732;
  assign n1734 = ~n533 & n854;
  assign n1735 = n2217 & n1732;
  assign n1736 = n2217 & ~n1732;
  assign n1737 = ~n2217 & n1732;
  assign n1738 = ~n1736 & ~n1737;
  assign n1739 = ~n1733 & ~n2437;
  assign n1740 = ~n535 & ~n536;
  assign n1741 = ~n2216 & ~n1740;
  assign n1742 = ~n535 & n850;
  assign n1743 = n2216 & n1740;
  assign n1744 = n2216 & ~n1740;
  assign n1745 = ~n2216 & n1740;
  assign n1746 = ~n1744 & ~n1745;
  assign n1747 = ~n1741 & ~n2439;
  assign n1748 = ~n537 & ~n538;
  assign n1749 = ~n2215 & ~n1748;
  assign n1750 = ~n537 & n846;
  assign n1751 = n2215 & n1748;
  assign n1752 = n2215 & ~n1748;
  assign n1753 = ~n2215 & n1748;
  assign n1754 = ~n1752 & ~n1753;
  assign n1755 = ~n1749 & ~n2441;
  assign n1756 = ~n539 & ~n540;
  assign n1757 = ~n2214 & ~n1756;
  assign n1758 = ~n539 & n842;
  assign n1759 = n2214 & n1756;
  assign n1760 = n2214 & ~n1756;
  assign n1761 = ~n2214 & n1756;
  assign n1762 = ~n1760 & ~n1761;
  assign n1763 = ~n1757 & ~n2443;
  assign n1764 = ~n541 & ~n542;
  assign n1765 = ~n2213 & ~n1764;
  assign n1766 = ~n541 & n838;
  assign n1767 = n2213 & n1764;
  assign n1768 = n2213 & ~n1764;
  assign n1769 = ~n2213 & n1764;
  assign n1770 = ~n1768 & ~n1769;
  assign n1771 = ~n1765 & ~n2445;
  assign n1772 = ~n543 & ~n544;
  assign n1773 = ~n2212 & ~n1772;
  assign n1774 = ~n543 & n834;
  assign n1775 = n2212 & n1772;
  assign n1776 = n2212 & ~n1772;
  assign n1777 = ~n2212 & n1772;
  assign n1778 = ~n1776 & ~n1777;
  assign n1779 = ~n1773 & ~n2447;
  assign n1780 = ~n545 & ~n546;
  assign n1781 = ~n2211 & ~n1780;
  assign n1782 = ~n545 & n830;
  assign n1783 = n2211 & n1780;
  assign n1784 = n2211 & ~n1780;
  assign n1785 = ~n2211 & n1780;
  assign n1786 = ~n1784 & ~n1785;
  assign n1787 = ~n1781 & ~n2449;
  assign n1788 = ~n547 & ~n548;
  assign n1789 = ~n2210 & ~n1788;
  assign n1790 = ~n547 & n826;
  assign n1791 = n2210 & n1788;
  assign n1792 = n2210 & ~n1788;
  assign n1793 = ~n2210 & n1788;
  assign n1794 = ~n1792 & ~n1793;
  assign n1795 = ~n1789 & ~n2451;
  assign n1796 = ~n549 & ~n550;
  assign n1797 = ~n2209 & ~n1796;
  assign n1798 = ~n549 & n822;
  assign n1799 = n2209 & n1796;
  assign n1800 = n2209 & ~n1796;
  assign n1801 = ~n2209 & n1796;
  assign n1802 = ~n1800 & ~n1801;
  assign n1803 = ~n1797 & ~n2453;
  assign n1804 = ~n551 & ~n552;
  assign n1805 = ~n2208 & ~n1804;
  assign n1806 = ~n551 & n818;
  assign n1807 = n2208 & n1804;
  assign n1808 = n2208 & ~n1804;
  assign n1809 = ~n2208 & n1804;
  assign n1810 = ~n1808 & ~n1809;
  assign n1811 = ~n1805 & ~n2455;
  assign n1812 = ~n553 & ~n554;
  assign n1813 = ~n2207 & ~n1812;
  assign n1814 = ~n553 & n814;
  assign n1815 = n2207 & n1812;
  assign n1816 = n2207 & ~n1812;
  assign n1817 = ~n2207 & n1812;
  assign n1818 = ~n1816 & ~n1817;
  assign n1819 = ~n1813 & ~n2457;
  assign n1820 = ~n555 & ~n556;
  assign n1821 = ~n2206 & ~n1820;
  assign n1822 = ~n555 & n810;
  assign n1823 = n2206 & n1820;
  assign n1824 = n2206 & ~n1820;
  assign n1825 = ~n2206 & n1820;
  assign n1826 = ~n1824 & ~n1825;
  assign n1827 = ~n1821 & ~n2459;
  assign n1828 = ~n557 & ~n558;
  assign n1829 = ~n2205 & ~n1828;
  assign n1830 = ~n557 & n806;
  assign n1831 = n2205 & n1828;
  assign n1832 = n2205 & ~n1828;
  assign n1833 = ~n2205 & n1828;
  assign n1834 = ~n1832 & ~n1833;
  assign n1835 = ~n1829 & ~n2461;
  assign n1836 = ~n559 & ~n560;
  assign n1837 = ~n2204 & ~n1836;
  assign n1838 = ~n559 & n802;
  assign n1839 = n2204 & n1836;
  assign n1840 = n2204 & ~n1836;
  assign n1841 = ~n2204 & n1836;
  assign n1842 = ~n1840 & ~n1841;
  assign n1843 = ~n1837 & ~n2463;
  assign n1844 = ~n561 & ~n562;
  assign n1845 = ~n2203 & ~n1844;
  assign n1846 = ~n561 & n798;
  assign n1847 = n2203 & n1844;
  assign n1848 = n2203 & ~n1844;
  assign n1849 = ~n2203 & n1844;
  assign n1850 = ~n1848 & ~n1849;
  assign n1851 = ~n1845 & ~n2465;
  assign n1852 = ~n563 & ~n564;
  assign n1853 = ~n2202 & ~n1852;
  assign n1854 = ~n563 & n794;
  assign n1855 = n2202 & n1852;
  assign n1856 = n2202 & ~n1852;
  assign n1857 = ~n2202 & n1852;
  assign n1858 = ~n1856 & ~n1857;
  assign n1859 = ~n1853 & ~n2467;
  assign n1860 = ~n565 & ~n566;
  assign n1861 = ~n2201 & ~n1860;
  assign n1862 = ~n565 & n790;
  assign n1863 = n2201 & n1860;
  assign n1864 = n2201 & ~n1860;
  assign n1865 = ~n2201 & n1860;
  assign n1866 = ~n1864 & ~n1865;
  assign n1867 = ~n1861 & ~n2469;
  assign n1868 = ~n567 & ~n568;
  assign n1869 = ~n2200 & ~n1868;
  assign n1870 = ~n567 & n786;
  assign n1871 = n2200 & n1868;
  assign n1872 = n2200 & ~n1868;
  assign n1873 = ~n2200 & n1868;
  assign n1874 = ~n1872 & ~n1873;
  assign n1875 = ~n1869 & ~n2471;
  assign n1876 = ~n569 & ~n570;
  assign n1877 = ~n2199 & ~n1876;
  assign n1878 = ~n569 & n782;
  assign n1879 = n2199 & n1876;
  assign n1880 = n2199 & ~n1876;
  assign n1881 = ~n2199 & n1876;
  assign n1882 = ~n1880 & ~n1881;
  assign n1883 = ~n1877 & ~n2473;
  assign n1884 = ~n571 & ~n572;
  assign n1885 = ~n2198 & ~n1884;
  assign n1886 = ~n571 & n778;
  assign n1887 = n2198 & n1884;
  assign n1888 = n2198 & ~n1884;
  assign n1889 = ~n2198 & n1884;
  assign n1890 = ~n1888 & ~n1889;
  assign n1891 = ~n1885 & ~n2475;
  assign n1892 = ~n573 & ~n574;
  assign n1893 = ~n2197 & ~n1892;
  assign n1894 = ~n573 & n774;
  assign n1895 = n2197 & n1892;
  assign n1896 = n2197 & ~n1892;
  assign n1897 = ~n2197 & n1892;
  assign n1898 = ~n1896 & ~n1897;
  assign n1899 = ~n1893 & ~n2477;
  assign n1900 = ~n575 & ~n576;
  assign n1901 = ~n2196 & ~n1900;
  assign n1902 = ~n575 & n770;
  assign n1903 = n2196 & n1900;
  assign n1904 = n2196 & ~n1900;
  assign n1905 = ~n2196 & n1900;
  assign n1906 = ~n1904 & ~n1905;
  assign n1907 = ~n1901 & ~n2479;
  assign n1908 = ~n577 & ~n578;
  assign n1909 = ~n2195 & ~n1908;
  assign n1910 = ~n577 & n766;
  assign n1911 = n2195 & n1908;
  assign n1912 = n2195 & ~n1908;
  assign n1913 = ~n2195 & n1908;
  assign n1914 = ~n1912 & ~n1913;
  assign n1915 = ~n1909 & ~n2481;
  assign n1916 = ~n579 & ~n580;
  assign n1917 = ~n2194 & ~n1916;
  assign n1918 = ~n579 & n762;
  assign n1919 = n2194 & n1916;
  assign n1920 = n2194 & ~n1916;
  assign n1921 = ~n2194 & n1916;
  assign n1922 = ~n1920 & ~n1921;
  assign n1923 = ~n1917 & ~n2483;
  assign n1924 = ~n581 & ~n582;
  assign n1925 = ~n2193 & ~n1924;
  assign n1926 = ~n581 & n758;
  assign n1927 = n2193 & n1924;
  assign n1928 = n2193 & ~n1924;
  assign n1929 = ~n2193 & n1924;
  assign n1930 = ~n1928 & ~n1929;
  assign n1931 = ~n1925 & ~n2485;
  assign n1932 = ~n583 & ~n584;
  assign n1933 = ~n2192 & ~n1932;
  assign n1934 = ~n583 & n754;
  assign n1935 = n2192 & n1932;
  assign n1936 = n2192 & ~n1932;
  assign n1937 = ~n2192 & n1932;
  assign n1938 = ~n1936 & ~n1937;
  assign n1939 = ~n1933 & ~n2487;
  assign n1940 = ~n585 & ~n586;
  assign n1941 = ~n2191 & ~n1940;
  assign n1942 = ~n585 & n750;
  assign n1943 = n2191 & n1940;
  assign n1944 = n2191 & ~n1940;
  assign n1945 = ~n2191 & n1940;
  assign n1946 = ~n1944 & ~n1945;
  assign n1947 = ~n1941 & ~n2489;
  assign n1948 = ~n587 & ~n588;
  assign n1949 = ~n2190 & ~n1948;
  assign n1950 = ~n587 & n746;
  assign n1951 = n2190 & n1948;
  assign n1952 = n2190 & ~n1948;
  assign n1953 = ~n2190 & n1948;
  assign n1954 = ~n1952 & ~n1953;
  assign n1955 = ~n1949 & ~n2491;
  assign n1956 = ~n589 & ~n590;
  assign n1957 = ~n2189 & ~n1956;
  assign n1958 = ~n589 & n742;
  assign n1959 = n2189 & n1956;
  assign n1960 = n2189 & ~n1956;
  assign n1961 = ~n2189 & n1956;
  assign n1962 = ~n1960 & ~n1961;
  assign n1963 = ~n1957 & ~n2493;
  assign n1964 = ~n591 & ~n592;
  assign n1965 = ~n2188 & ~n1964;
  assign n1966 = ~n591 & n738;
  assign n1967 = n2188 & n1964;
  assign n1968 = n2188 & ~n1964;
  assign n1969 = ~n2188 & n1964;
  assign n1970 = ~n1968 & ~n1969;
  assign n1971 = ~n1965 & ~n2495;
  assign n1972 = ~n593 & ~n594;
  assign n1973 = ~n2187 & ~n1972;
  assign n1974 = ~n593 & n734;
  assign n1975 = n2187 & n1972;
  assign n1976 = n2187 & ~n1972;
  assign n1977 = ~n2187 & n1972;
  assign n1978 = ~n1976 & ~n1977;
  assign n1979 = ~n1973 & ~n2497;
  assign n1980 = ~n595 & ~n596;
  assign n1981 = ~n2186 & ~n1980;
  assign n1982 = ~n595 & n730;
  assign n1983 = n2186 & n1980;
  assign n1984 = n2186 & ~n1980;
  assign n1985 = ~n2186 & n1980;
  assign n1986 = ~n1984 & ~n1985;
  assign n1987 = ~n1981 & ~n2499;
  assign n1988 = ~n597 & ~n598;
  assign n1989 = ~n2185 & ~n1988;
  assign n1990 = ~n597 & n726;
  assign n1991 = n2185 & n1988;
  assign n1992 = n2185 & ~n1988;
  assign n1993 = ~n2185 & n1988;
  assign n1994 = ~n1992 & ~n1993;
  assign n1995 = ~n1989 & ~n2501;
  assign n1996 = ~n599 & ~n600;
  assign n1997 = ~n2184 & ~n1996;
  assign n1998 = ~n599 & n722;
  assign n1999 = n2184 & n1996;
  assign n2000 = n2184 & ~n1996;
  assign n2001 = ~n2184 & n1996;
  assign n2002 = ~n2000 & ~n2001;
  assign n2003 = ~n1997 & ~n2503;
  assign n2004 = ~n601 & ~n602;
  assign n2005 = ~n2183 & ~n2004;
  assign n2006 = ~n601 & n718;
  assign n2007 = n2183 & n2004;
  assign n2008 = n2183 & ~n2004;
  assign n2009 = ~n2183 & n2004;
  assign n2010 = ~n2008 & ~n2009;
  assign n2011 = ~n2005 & ~n2505;
  assign n2012 = ~n603 & ~n604;
  assign n2013 = ~n2182 & ~n2012;
  assign n2014 = ~n603 & n714;
  assign n2015 = n2182 & n2012;
  assign n2016 = n2182 & ~n2012;
  assign n2017 = ~n2182 & n2012;
  assign n2018 = ~n2016 & ~n2017;
  assign n2019 = ~n2013 & ~n2507;
  assign n2020 = ~n605 & ~n606;
  assign n2021 = ~n2181 & ~n2020;
  assign n2022 = ~n605 & n710;
  assign n2023 = n2181 & n2020;
  assign n2024 = n2181 & ~n2020;
  assign n2025 = ~n2181 & n2020;
  assign n2026 = ~n2024 & ~n2025;
  assign n2027 = ~n2021 & ~n2509;
  assign n2028 = ~n607 & ~n608;
  assign n2029 = ~n2180 & ~n2028;
  assign n2030 = ~n607 & n706;
  assign n2031 = n2180 & n2028;
  assign n2032 = n2180 & ~n2028;
  assign n2033 = ~n2180 & n2028;
  assign n2034 = ~n2032 & ~n2033;
  assign n2035 = ~n2029 & ~n2511;
  assign n2036 = ~n609 & ~n610;
  assign n2037 = ~n2179 & ~n2036;
  assign n2038 = ~n609 & n702;
  assign n2039 = n2179 & n2036;
  assign n2040 = n2179 & ~n2036;
  assign n2041 = ~n2179 & n2036;
  assign n2042 = ~n2040 & ~n2041;
  assign n2043 = ~n2037 & ~n2513;
  assign n2044 = ~n611 & ~n612;
  assign n2045 = ~n2178 & ~n2044;
  assign n2046 = ~n611 & n698;
  assign n2047 = n2178 & n2044;
  assign n2048 = n2178 & ~n2044;
  assign n2049 = ~n2178 & n2044;
  assign n2050 = ~n2048 & ~n2049;
  assign n2051 = ~n2045 & ~n2515;
  assign n2052 = ~n613 & ~n614;
  assign n2053 = ~n2177 & ~n2052;
  assign n2054 = ~n613 & n694;
  assign n2055 = n2177 & n2052;
  assign n2056 = n2177 & ~n2052;
  assign n2057 = ~n2177 & n2052;
  assign n2058 = ~n2056 & ~n2057;
  assign n2059 = ~n2053 & ~n2517;
  assign n2060 = ~n615 & ~n616;
  assign n2061 = ~n2176 & ~n2060;
  assign n2062 = ~n615 & n690;
  assign n2063 = n2176 & n2060;
  assign n2064 = n2176 & ~n2060;
  assign n2065 = ~n2176 & n2060;
  assign n2066 = ~n2064 & ~n2065;
  assign n2067 = ~n2061 & ~n2519;
  assign n2068 = ~n617 & ~n618;
  assign n2069 = ~n2175 & ~n2068;
  assign n2070 = ~n617 & n686;
  assign n2071 = n2175 & n2068;
  assign n2072 = n2175 & ~n2068;
  assign n2073 = ~n2175 & n2068;
  assign n2074 = ~n2072 & ~n2073;
  assign n2075 = ~n2069 & ~n2521;
  assign n2076 = ~n619 & ~n620;
  assign n2077 = ~n2174 & ~n2076;
  assign n2078 = ~n619 & n682;
  assign n2079 = n2174 & n2076;
  assign n2080 = n2174 & ~n2076;
  assign n2081 = ~n2174 & n2076;
  assign n2082 = ~n2080 & ~n2081;
  assign n2083 = ~n2077 & ~n2523;
  assign n2084 = ~n621 & ~n622;
  assign n2085 = ~n2173 & ~n2084;
  assign n2086 = ~n621 & n678;
  assign n2087 = n2173 & n2084;
  assign n2088 = n2173 & ~n2084;
  assign n2089 = ~n2173 & n2084;
  assign n2090 = ~n2088 & ~n2089;
  assign n2091 = ~n2085 & ~n2525;
  assign n2092 = ~n623 & ~n624;
  assign n2093 = ~n2172 & ~n2092;
  assign n2094 = ~n623 & n674;
  assign n2095 = n2172 & n2092;
  assign n2096 = n2172 & ~n2092;
  assign n2097 = ~n2172 & n2092;
  assign n2098 = ~n2096 & ~n2097;
  assign n2099 = ~n2093 & ~n2527;
  assign n2100 = ~n625 & ~n626;
  assign n2101 = ~n2171 & ~n2100;
  assign n2102 = ~n625 & n670;
  assign n2103 = n2171 & n2100;
  assign n2104 = n2171 & ~n2100;
  assign n2105 = ~n2171 & n2100;
  assign n2106 = ~n2104 & ~n2105;
  assign n2107 = ~n2101 & ~n2529;
  assign n2108 = ~n627 & ~n628;
  assign n2109 = ~n2170 & ~n2108;
  assign n2110 = ~n627 & n666;
  assign n2111 = n2170 & n2108;
  assign n2112 = n2170 & ~n2108;
  assign n2113 = ~n2170 & n2108;
  assign n2114 = ~n2112 & ~n2113;
  assign n2115 = ~n2109 & ~n2531;
  assign n2116 = ~n629 & ~n630;
  assign n2117 = ~n2169 & ~n2116;
  assign n2118 = ~n629 & n662;
  assign n2119 = n2169 & n2116;
  assign n2120 = n2169 & ~n2116;
  assign n2121 = ~n2169 & n2116;
  assign n2122 = ~n2120 & ~n2121;
  assign n2123 = ~n2117 & ~n2533;
  assign n2124 = ~n631 & ~n632;
  assign n2125 = ~n2168 & ~n2124;
  assign n2126 = ~n631 & n658;
  assign n2127 = n2168 & n2124;
  assign n2128 = n2168 & ~n2124;
  assign n2129 = ~n2168 & n2124;
  assign n2130 = ~n2128 & ~n2129;
  assign n2131 = ~n2125 & ~n2535;
  assign n2132 = ~n633 & ~n634;
  assign n2133 = ~n2167 & ~n2132;
  assign n2134 = ~n633 & n654;
  assign n2135 = n2167 & n2132;
  assign n2136 = n2167 & ~n2132;
  assign n2137 = ~n2167 & n2132;
  assign n2138 = ~n2136 & ~n2137;
  assign n2139 = ~n2133 & ~n2537;
  assign n2140 = ~n635 & ~n636;
  assign n2141 = ~n2166 & ~n2140;
  assign n2142 = ~n635 & n650;
  assign n2143 = n2166 & n2140;
  assign n2144 = n2166 & ~n2140;
  assign n2145 = ~n2166 & n2140;
  assign n2146 = ~n2144 & ~n2145;
  assign n2147 = ~n2141 & ~n2539;
  assign n2148 = ~n637 & ~n638;
  assign n2149 = ~n2165 & ~n2148;
  assign n2150 = ~n637 & n646;
  assign n2151 = n2165 & n2148;
  assign n2152 = n2165 & ~n2148;
  assign n2153 = ~n2165 & n2148;
  assign n2154 = ~n2152 & ~n2153;
  assign n2155 = ~n2149 & ~n2541;
  assign n2156 = ~n639 & ~n641;
  assign n2157 = n640 & ~n2156;
  assign n2158 = ~n640 & n2156;
  assign n2159 = ~n2157 & ~n2158;
  assign n2160 = ~pi0  & ~pi128 ;
  assign n2161 = pi0  & ~pi128 ;
  assign n2162 = ~pi0  & pi128 ;
  assign n2163 = ~n2161 & ~n2162;
  assign n2164 = ~n640 & ~n2160;
  assign n2165 = n644 | ~n645;
  assign n2166 = n648 | ~n649;
  assign n2167 = n652 | ~n653;
  assign n2168 = n656 | ~n657;
  assign n2169 = n660 | ~n661;
  assign n2170 = n664 | ~n665;
  assign n2171 = n668 | ~n669;
  assign n2172 = n672 | ~n673;
  assign n2173 = n676 | ~n677;
  assign n2174 = n680 | ~n681;
  assign n2175 = n684 | ~n685;
  assign n2176 = n688 | ~n689;
  assign n2177 = n692 | ~n693;
  assign n2178 = n696 | ~n697;
  assign n2179 = n700 | ~n701;
  assign n2180 = n704 | ~n705;
  assign n2181 = n708 | ~n709;
  assign n2182 = n712 | ~n713;
  assign n2183 = n716 | ~n717;
  assign n2184 = n720 | ~n721;
  assign n2185 = n724 | ~n725;
  assign n2186 = n728 | ~n729;
  assign n2187 = n732 | ~n733;
  assign n2188 = n736 | ~n737;
  assign n2189 = n740 | ~n741;
  assign n2190 = n744 | ~n745;
  assign n2191 = n748 | ~n749;
  assign n2192 = n752 | ~n753;
  assign n2193 = n756 | ~n757;
  assign n2194 = n760 | ~n761;
  assign n2195 = n764 | ~n765;
  assign n2196 = n768 | ~n769;
  assign n2197 = n772 | ~n773;
  assign n2198 = n776 | ~n777;
  assign n2199 = n780 | ~n781;
  assign n2200 = n784 | ~n785;
  assign n2201 = n788 | ~n789;
  assign n2202 = n792 | ~n793;
  assign n2203 = n796 | ~n797;
  assign n2204 = n800 | ~n801;
  assign n2205 = n804 | ~n805;
  assign n2206 = n808 | ~n809;
  assign n2207 = n812 | ~n813;
  assign n2208 = n816 | ~n817;
  assign n2209 = n820 | ~n821;
  assign n2210 = n824 | ~n825;
  assign n2211 = n828 | ~n829;
  assign n2212 = n832 | ~n833;
  assign n2213 = n836 | ~n837;
  assign n2214 = n840 | ~n841;
  assign n2215 = n844 | ~n845;
  assign n2216 = n848 | ~n849;
  assign n2217 = n852 | ~n853;
  assign n2218 = n856 | ~n857;
  assign n2219 = n860 | ~n861;
  assign n2220 = n864 | ~n865;
  assign n2221 = n868 | ~n869;
  assign n2222 = n872 | ~n873;
  assign n2223 = n876 | ~n877;
  assign n2224 = n880 | ~n881;
  assign n2225 = n884 | ~n885;
  assign n2226 = n888 | ~n889;
  assign n2227 = n892 | ~n893;
  assign n2228 = n896 | ~n897;
  assign n2229 = n900 | ~n901;
  assign n2230 = n904 | ~n905;
  assign n2231 = n908 | ~n909;
  assign n2232 = n912 | ~n913;
  assign n2233 = n916 | ~n917;
  assign n2234 = n920 | ~n921;
  assign n2235 = n924 | ~n925;
  assign n2236 = n928 | ~n929;
  assign n2237 = n932 | ~n933;
  assign n2238 = n936 | ~n937;
  assign n2239 = n940 | ~n941;
  assign n2240 = n944 | ~n945;
  assign n2241 = n948 | ~n949;
  assign n2242 = n952 | ~n953;
  assign n2243 = n956 | ~n957;
  assign n2244 = n960 | ~n961;
  assign n2245 = n964 | ~n965;
  assign n2246 = n968 | ~n969;
  assign n2247 = n972 | ~n973;
  assign n2248 = n976 | ~n977;
  assign n2249 = n980 | ~n981;
  assign n2250 = n984 | ~n985;
  assign n2251 = n988 | ~n989;
  assign n2252 = n992 | ~n993;
  assign n2253 = n996 | ~n997;
  assign n2254 = n1000 | ~n1001;
  assign n2255 = n1004 | ~n1005;
  assign n2256 = n1008 | ~n1009;
  assign n2257 = n1012 | ~n1013;
  assign n2258 = n1016 | ~n1017;
  assign n2259 = n1020 | ~n1021;
  assign n2260 = n1024 | ~n1025;
  assign n2261 = n1028 | ~n1029;
  assign n2262 = n1032 | ~n1033;
  assign n2263 = n1036 | ~n1037;
  assign n2264 = n1040 | ~n1041;
  assign n2265 = n1044 | ~n1045;
  assign n2266 = n1048 | ~n1049;
  assign n2267 = n1052 | ~n1053;
  assign n2268 = n1056 | ~n1057;
  assign n2269 = n1060 | ~n1061;
  assign n2270 = n1064 | ~n1065;
  assign n2271 = n1068 | ~n1069;
  assign n2272 = n1072 | ~n1073;
  assign n2273 = n1076 | ~n1077;
  assign n2274 = n1080 | ~n1081;
  assign n2275 = n1084 | ~n1085;
  assign n2276 = n1088 | ~n1089;
  assign n2277 = n1092 | ~n1093;
  assign n2278 = n1096 | ~n1097;
  assign n2279 = n1100 | ~n1101;
  assign n2280 = n1104 | ~n1105;
  assign n2281 = n1108 | ~n1109;
  assign n2282 = n1112 | ~n1113;
  assign n2283 = n1116 | ~n1117;
  assign n2284 = n1120 | ~n1121;
  assign n2285 = n1124 | ~n1125;
  assign n2286 = n1128 | ~n1129;
  assign n2287 = n1132 | ~n1133;
  assign n2288 = n1136 | ~n1137;
  assign n2289 = n1140 | ~n1141;
  assign n2290 = n1144 | ~n1145;
  assign po127  = n1150 | ~n1151;
  assign n2292 = n1154 | ~n1155;
  assign n2293 = n1158 | n1159;
  assign po126  = n1162 | ~n1163;
  assign n2295 = n1166 | n1167;
  assign po125  = n1170 | ~n1171;
  assign n2297 = n1174 | n1175;
  assign po124  = n1178 | ~n1179;
  assign n2299 = n1182 | n1183;
  assign po123  = n1186 | ~n1187;
  assign n2301 = n1190 | n1191;
  assign po122  = n1194 | ~n1195;
  assign n2303 = n1198 | n1199;
  assign po121  = n1202 | ~n1203;
  assign n2305 = n1206 | n1207;
  assign po120  = n1210 | ~n1211;
  assign n2307 = n1214 | n1215;
  assign po119  = n1218 | ~n1219;
  assign n2309 = n1222 | n1223;
  assign po118  = n1226 | ~n1227;
  assign n2311 = n1230 | n1231;
  assign po117  = n1234 | ~n1235;
  assign n2313 = n1238 | n1239;
  assign po116  = n1242 | ~n1243;
  assign n2315 = n1246 | n1247;
  assign po115  = n1250 | ~n1251;
  assign n2317 = n1254 | n1255;
  assign po114  = n1258 | ~n1259;
  assign n2319 = n1262 | n1263;
  assign po113  = n1266 | ~n1267;
  assign n2321 = n1270 | n1271;
  assign po112  = n1274 | ~n1275;
  assign n2323 = n1278 | n1279;
  assign po111  = n1282 | ~n1283;
  assign n2325 = n1286 | n1287;
  assign po110  = n1290 | ~n1291;
  assign n2327 = n1294 | n1295;
  assign po109  = n1298 | ~n1299;
  assign n2329 = n1302 | n1303;
  assign po108  = n1306 | ~n1307;
  assign n2331 = n1310 | n1311;
  assign po107  = n1314 | ~n1315;
  assign n2333 = n1318 | n1319;
  assign po106  = n1322 | ~n1323;
  assign n2335 = n1326 | n1327;
  assign po105  = n1330 | ~n1331;
  assign n2337 = n1334 | n1335;
  assign po104  = n1338 | ~n1339;
  assign n2339 = n1342 | n1343;
  assign po103  = n1346 | ~n1347;
  assign n2341 = n1350 | n1351;
  assign po102  = n1354 | ~n1355;
  assign n2343 = n1358 | n1359;
  assign po101  = n1362 | ~n1363;
  assign n2345 = n1366 | n1367;
  assign po100  = n1370 | ~n1371;
  assign n2347 = n1374 | n1375;
  assign po99  = n1378 | ~n1379;
  assign n2349 = n1382 | n1383;
  assign po98  = n1386 | ~n1387;
  assign n2351 = n1390 | n1391;
  assign po97  = n1394 | ~n1395;
  assign n2353 = n1398 | n1399;
  assign po96  = n1402 | ~n1403;
  assign n2355 = n1406 | n1407;
  assign po95  = n1410 | ~n1411;
  assign n2357 = n1414 | n1415;
  assign po94  = n1418 | ~n1419;
  assign n2359 = n1422 | n1423;
  assign po93  = n1426 | ~n1427;
  assign n2361 = n1430 | n1431;
  assign po92  = n1434 | ~n1435;
  assign n2363 = n1438 | n1439;
  assign po91  = n1442 | ~n1443;
  assign n2365 = n1446 | n1447;
  assign po90  = n1450 | ~n1451;
  assign n2367 = n1454 | n1455;
  assign po89  = n1458 | ~n1459;
  assign n2369 = n1462 | n1463;
  assign po88  = n1466 | ~n1467;
  assign n2371 = n1470 | n1471;
  assign po87  = n1474 | ~n1475;
  assign n2373 = n1478 | n1479;
  assign po86  = n1482 | ~n1483;
  assign n2375 = n1486 | n1487;
  assign po85  = n1490 | ~n1491;
  assign n2377 = n1494 | n1495;
  assign po84  = n1498 | ~n1499;
  assign n2379 = n1502 | n1503;
  assign po83  = n1506 | ~n1507;
  assign n2381 = n1510 | n1511;
  assign po82  = n1514 | ~n1515;
  assign n2383 = n1518 | n1519;
  assign po81  = n1522 | ~n1523;
  assign n2385 = n1526 | n1527;
  assign po80  = n1530 | ~n1531;
  assign n2387 = n1534 | n1535;
  assign po79  = n1538 | ~n1539;
  assign n2389 = n1542 | n1543;
  assign po78  = n1546 | ~n1547;
  assign n2391 = n1550 | n1551;
  assign po77  = n1554 | ~n1555;
  assign n2393 = n1558 | n1559;
  assign po76  = n1562 | ~n1563;
  assign n2395 = n1566 | n1567;
  assign po75  = n1570 | ~n1571;
  assign n2397 = n1574 | n1575;
  assign po74  = n1578 | ~n1579;
  assign n2399 = n1582 | n1583;
  assign po73  = n1586 | ~n1587;
  assign n2401 = n1590 | n1591;
  assign po72  = n1594 | ~n1595;
  assign n2403 = n1598 | n1599;
  assign po71  = n1602 | ~n1603;
  assign n2405 = n1606 | n1607;
  assign po70  = n1610 | ~n1611;
  assign n2407 = n1614 | n1615;
  assign po69  = n1618 | ~n1619;
  assign n2409 = n1622 | n1623;
  assign po68  = n1626 | ~n1627;
  assign n2411 = n1630 | n1631;
  assign po67  = n1634 | ~n1635;
  assign n2413 = n1638 | n1639;
  assign po66  = n1642 | ~n1643;
  assign n2415 = n1646 | n1647;
  assign po65  = n1650 | ~n1651;
  assign n2417 = n1654 | n1655;
  assign po64  = n1658 | ~n1659;
  assign n2419 = n1662 | n1663;
  assign po63  = n1666 | ~n1667;
  assign n2421 = n1670 | n1671;
  assign po62  = n1674 | ~n1675;
  assign n2423 = n1678 | n1679;
  assign po61  = n1682 | ~n1683;
  assign n2425 = n1686 | n1687;
  assign po60  = n1690 | ~n1691;
  assign n2427 = n1694 | n1695;
  assign po59  = n1698 | ~n1699;
  assign n2429 = n1702 | n1703;
  assign po58  = n1706 | ~n1707;
  assign n2431 = n1710 | n1711;
  assign po57  = n1714 | ~n1715;
  assign n2433 = n1718 | n1719;
  assign po56  = n1722 | ~n1723;
  assign n2435 = n1726 | n1727;
  assign po55  = n1730 | ~n1731;
  assign n2437 = n1734 | n1735;
  assign po54  = n1738 | ~n1739;
  assign n2439 = n1742 | n1743;
  assign po53  = n1746 | ~n1747;
  assign n2441 = n1750 | n1751;
  assign po52  = n1754 | ~n1755;
  assign n2443 = n1758 | n1759;
  assign po51  = n1762 | ~n1763;
  assign n2445 = n1766 | n1767;
  assign po50  = n1770 | ~n1771;
  assign n2447 = n1774 | n1775;
  assign po49  = n1778 | ~n1779;
  assign n2449 = n1782 | n1783;
  assign po48  = n1786 | ~n1787;
  assign n2451 = n1790 | n1791;
  assign po47  = n1794 | ~n1795;
  assign n2453 = n1798 | n1799;
  assign po46  = n1802 | ~n1803;
  assign n2455 = n1806 | n1807;
  assign po45  = n1810 | ~n1811;
  assign n2457 = n1814 | n1815;
  assign po44  = n1818 | ~n1819;
  assign n2459 = n1822 | n1823;
  assign po43  = n1826 | ~n1827;
  assign n2461 = n1830 | n1831;
  assign po42  = n1834 | ~n1835;
  assign n2463 = n1838 | n1839;
  assign po41  = n1842 | ~n1843;
  assign n2465 = n1846 | n1847;
  assign po40  = n1850 | ~n1851;
  assign n2467 = n1854 | n1855;
  assign po39  = n1858 | ~n1859;
  assign n2469 = n1862 | n1863;
  assign po38  = n1866 | ~n1867;
  assign n2471 = n1870 | n1871;
  assign po37  = n1874 | ~n1875;
  assign n2473 = n1878 | n1879;
  assign po36  = n1882 | ~n1883;
  assign n2475 = n1886 | n1887;
  assign po35  = n1890 | ~n1891;
  assign n2477 = n1894 | n1895;
  assign po34  = n1898 | ~n1899;
  assign n2479 = n1902 | n1903;
  assign po33  = n1906 | ~n1907;
  assign n2481 = n1910 | n1911;
  assign po32  = n1914 | ~n1915;
  assign n2483 = n1918 | n1919;
  assign po31  = n1922 | ~n1923;
  assign n2485 = n1926 | n1927;
  assign po30  = n1930 | ~n1931;
  assign n2487 = n1934 | n1935;
  assign po29  = n1938 | ~n1939;
  assign n2489 = n1942 | n1943;
  assign po28  = n1946 | ~n1947;
  assign n2491 = n1950 | n1951;
  assign po27  = n1954 | ~n1955;
  assign n2493 = n1958 | n1959;
  assign po26  = n1962 | ~n1963;
  assign n2495 = n1966 | n1967;
  assign po25  = n1970 | ~n1971;
  assign n2497 = n1974 | n1975;
  assign po24  = n1978 | ~n1979;
  assign n2499 = n1982 | n1983;
  assign po23  = n1986 | ~n1987;
  assign n2501 = n1990 | n1991;
  assign po22  = n1994 | ~n1995;
  assign n2503 = n1998 | n1999;
  assign po21  = n2002 | ~n2003;
  assign n2505 = n2006 | n2007;
  assign po20  = n2010 | ~n2011;
  assign n2507 = n2014 | n2015;
  assign po19  = n2018 | ~n2019;
  assign n2509 = n2022 | n2023;
  assign po18  = n2026 | ~n2027;
  assign n2511 = n2030 | n2031;
  assign po17  = n2034 | ~n2035;
  assign n2513 = n2038 | n2039;
  assign po16  = n2042 | ~n2043;
  assign n2515 = n2046 | n2047;
  assign po15  = n2050 | ~n2051;
  assign n2517 = n2054 | n2055;
  assign po14  = n2058 | ~n2059;
  assign n2519 = n2062 | n2063;
  assign po13  = n2066 | ~n2067;
  assign n2521 = n2070 | n2071;
  assign po12  = n2074 | ~n2075;
  assign n2523 = n2078 | n2079;
  assign po11  = n2082 | ~n2083;
  assign n2525 = n2086 | n2087;
  assign po10  = n2090 | ~n2091;
  assign n2527 = n2094 | n2095;
  assign po9  = n2098 | ~n2099;
  assign n2529 = n2102 | n2103;
  assign po8  = n2106 | ~n2107;
  assign n2531 = n2110 | n2111;
  assign po7  = n2114 | ~n2115;
  assign n2533 = n2118 | n2119;
  assign po6  = n2122 | ~n2123;
  assign n2535 = n2126 | n2127;
  assign po5  = n2130 | ~n2131;
  assign n2537 = n2134 | n2135;
  assign po4  = n2138 | ~n2139;
  assign n2539 = n2142 | n2143;
  assign po3  = n2146 | ~n2147;
  assign n2541 = n2150 | n2151;
  assign po2  = n2154 | ~n2155;
  assign n2543 = n2163 | ~n2164;
  assign po0  = ~n2543;
  assign po1  = ~n2159;
  assign po128 = ~n2292;
endmodule
