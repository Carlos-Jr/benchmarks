module mem_ctrl ( 
    pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8,
    pi9, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17,
    pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26,
    pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35,
    pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44,
    pi45, pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53,
    pi54, pi55, pi56, pi57, pi58, pi59, pi60, pi61, pi62,
    pi63, pi64, pi65, pi66, pi67, pi68, pi69, pi70, pi71,
    pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79, pi80,
    pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88, pi89,
    pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97, pi98,
    pi99, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107,
    pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116,
    pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125,
    pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134,
    pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143,
    pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152,
    pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161,
    pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170,
    pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197,
    pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206,
    pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214, pi215,
    pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223, pi224,
    pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232, pi233,
    pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241, pi242,
    pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250, pi251,
    pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259, pi260,
    pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269,
    pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278,
    pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287,
    pi288, pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296,
    pi297, pi298, pi299, pi300, pi301, pi302, pi303, pi304, pi305,
    pi306, pi307, pi308, pi309, pi310, pi311, pi312, pi313, pi314,
    pi315, pi316, pi317, pi318, pi319, pi320, pi321, pi322, pi323,
    pi324, pi325, pi326, pi327, pi328, pi329, pi330, pi331, pi332,
    pi333, pi334, pi335, pi336, pi337, pi338, pi339, pi340, pi341,
    pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349, pi350,
    pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358, pi359,
    pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368,
    pi369, pi370, pi371, pi372, pi373, pi374, pi375, pi376, pi377,
    pi378, pi379, pi380, pi381, pi382, pi383, pi384, pi385, pi386,
    pi387, pi388, pi389, pi390, pi391, pi392, pi393, pi394, pi395,
    pi396, pi397, pi398, pi399, pi400, pi401, pi402, pi403, pi404,
    pi405, pi406, pi407, pi408, pi409, pi410, pi411, pi412, pi413,
    pi414, pi415, pi416, pi417, pi418, pi419, pi420, pi421, pi422,
    pi423, pi424, pi425, pi426, pi427, pi428, pi429, pi430, pi431,
    pi432, pi433, pi434, pi435, pi436, pi437, pi438, pi439, pi440,
    pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448, pi449,
    pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457, pi458,
    pi459, pi460, pi461, pi462, pi463, pi464, pi465, pi466, pi467,
    pi468, pi469, pi470, pi471, pi472, pi473, pi474, pi475, pi476,
    pi477, pi478, pi479, pi480, pi481, pi482, pi483, pi484, pi485,
    pi486, pi487, pi488, pi489, pi490, pi491, pi492, pi493, pi494,
    pi495, pi496, pi497, pi498, pi499, pi500, pi501, pi502, pi503,
    pi504, pi505, pi506, pi507, pi508, pi509, pi510, pi511, pi512,
    pi513, pi514, pi515, pi516, pi517, pi518, pi519, pi520, pi521,
    pi522, pi523, pi524, pi525, pi526, pi527, pi528, pi529, pi530,
    pi531, pi532, pi533, pi534, pi535, pi536, pi537, pi538, pi539,
    pi540, pi541, pi542, pi543, pi544, pi545, pi546, pi547, pi548,
    pi549, pi550, pi551, pi552, pi553, pi554, pi555, pi556, pi557,
    pi558, pi559, pi560, pi561, pi562, pi563, pi564, pi565, pi566,
    pi567, pi568, pi569, pi570, pi571, pi572, pi573, pi574, pi575,
    pi576, pi577, pi578, pi579, pi580, pi581, pi582, pi583, pi584,
    pi585, pi586, pi587, pi588, pi589, pi590, pi591, pi592, pi593,
    pi594, pi595, pi596, pi597, pi598, pi599, pi600, pi601, pi602,
    pi603, pi604, pi605, pi606, pi607, pi608, pi609, pi610, pi611,
    pi612, pi613, pi614, pi615, pi616, pi617, pi618, pi619, pi620,
    pi621, pi622, pi623, pi624, pi625, pi626, pi627, pi628, pi629,
    pi630, pi631, pi632, pi633, pi634, pi635, pi636, pi637, pi638,
    pi639, pi640, pi641, pi642, pi643, pi644, pi645, pi646, pi647,
    pi648, pi649, pi650, pi651, pi652, pi653, pi654, pi655, pi656,
    pi657, pi658, pi659, pi660, pi661, pi662, pi663, pi664, pi665,
    pi666, pi667, pi668, pi669, pi670, pi671, pi672, pi673, pi674,
    pi675, pi676, pi677, pi678, pi679, pi680, pi681, pi682, pi683,
    pi684, pi685, pi686, pi687, pi688, pi689, pi690, pi691, pi692,
    pi693, pi694, pi695, pi696, pi697, pi698, pi699, pi700, pi701,
    pi702, pi703, pi704, pi705, pi706, pi707, pi708, pi709, pi710,
    pi711, pi712, pi713, pi714, pi715, pi716, pi717, pi718, pi719,
    pi720, pi721, pi722, pi723, pi724, pi725, pi726, pi727, pi728,
    pi729, pi730, pi731, pi732, pi733, pi734, pi735, pi736, pi737,
    pi738, pi739, pi740, pi741, pi742, pi743, pi744, pi745, pi746,
    pi747, pi748, pi749, pi750, pi751, pi752, pi753, pi754, pi755,
    pi756, pi757, pi758, pi759, pi760, pi761, pi762, pi763, pi764,
    pi765, pi766, pi767, pi768, pi769, pi770, pi771, pi772, pi773,
    pi774, pi775, pi776, pi777, pi778, pi779, pi780, pi781, pi782,
    pi783, pi784, pi785, pi786, pi787, pi788, pi789, pi790, pi791,
    pi792, pi793, pi794, pi795, pi796, pi797, pi798, pi799, pi800,
    pi801, pi802, pi803, pi804, pi805, pi806, pi807, pi808, pi809,
    pi810, pi811, pi812, pi813, pi814, pi815, pi816, pi817, pi818,
    pi819, pi820, pi821, pi822, pi823, pi824, pi825, pi826, pi827,
    pi828, pi829, pi830, pi831, pi832, pi833, pi834, pi835, pi836,
    pi837, pi838, pi839, pi840, pi841, pi842, pi843, pi844, pi845,
    pi846, pi847, pi848, pi849, pi850, pi851, pi852, pi853, pi854,
    pi855, pi856, pi857, pi858, pi859, pi860, pi861, pi862, pi863,
    pi864, pi865, pi866, pi867, pi868, pi869, pi870, pi871, pi872,
    pi873, pi874, pi875, pi876, pi877, pi878, pi879, pi880, pi881,
    pi882, pi883, pi884, pi885, pi886, pi887, pi888, pi889, pi890,
    pi891, pi892, pi893, pi894, pi895, pi896, pi897, pi898, pi899,
    pi900, pi901, pi902, pi903, pi904, pi905, pi906, pi907, pi908,
    pi909, pi910, pi911, pi912, pi913, pi914, pi915, pi916, pi917,
    pi918, pi919, pi920, pi921, pi922, pi923, pi924, pi925, pi926,
    pi927, pi928, pi929, pi930, pi931, pi932, pi933, pi934, pi935,
    pi936, pi937, pi938, pi939, pi940, pi941, pi942, pi943, pi944,
    pi945, pi946, pi947, pi948, pi949, pi950, pi951, pi952, pi953,
    pi954, pi955, pi956, pi957, pi958, pi959, pi960, pi961, pi962,
    pi963, pi964, pi965, pi966, pi967, pi968, pi969, pi970, pi971,
    pi972, pi973, pi974, pi975, pi976, pi977, pi978, pi979, pi980,
    pi981, pi982, pi983, pi984, pi985, pi986, pi987, pi988, pi989,
    pi990, pi991, pi992, pi993, pi994, pi995, pi996, pi997, pi998,
    pi999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007,
    pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016,
    pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025,
    pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034,
    pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043,
    pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052,
    pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061,
    pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070,
    pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079,
    pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088,
    pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097,
    pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106,
    pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115,
    pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124,
    pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133,
    pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142,
    pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151,
    pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160,
    pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169,
    pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178,
    pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187,
    pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196,
    pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203,
    po0, po1, po2, po3, po4, po5, po6, po7, po8,
    po9, po10, po11, po12, po13, po14, po15, po16, po17,
    po18, po19, po20, po21, po22, po23, po24, po25, po26,
    po27, po28, po29, po30, po31, po32, po33, po34, po35,
    po36, po37, po38, po39, po40, po41, po42, po43, po44,
    po45, po46, po47, po48, po49, po50, po51, po52, po53,
    po54, po55, po56, po57, po58, po59, po60, po61, po62,
    po63, po64, po65, po66, po67, po68, po69, po70, po71,
    po72, po73, po74, po75, po76, po77, po78, po79, po80,
    po81, po82, po83, po84, po85, po86, po87, po88, po89,
    po90, po91, po92, po93, po94, po95, po96, po97, po98,
    po99, po100, po101, po102, po103, po104, po105, po106, po107,
    po108, po109, po110, po111, po112, po113, po114, po115, po116,
    po117, po118, po119, po120, po121, po122, po123, po124, po125,
    po126, po127, po128, po129, po130, po131, po132, po133, po134,
    po135, po136, po137, po138, po139, po140, po141, po142, po143,
    po144, po145, po146, po147, po148, po149, po150, po151, po152,
    po153, po154, po155, po156, po157, po158, po159, po160, po161,
    po162, po163, po164, po165, po166, po167, po168, po169, po170,
    po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188,
    po189, po190, po191, po192, po193, po194, po195, po196, po197,
    po198, po199, po200, po201, po202, po203, po204, po205, po206,
    po207, po208, po209, po210, po211, po212, po213, po214, po215,
    po216, po217, po218, po219, po220, po221, po222, po223, po224,
    po225, po226, po227, po228, po229, po230, po231, po232, po233,
    po234, po235, po236, po237, po238, po239, po240, po241, po242,
    po243, po244, po245, po246, po247, po248, po249, po250, po251,
    po252, po253, po254, po255, po256, po257, po258, po259, po260,
    po261, po262, po263, po264, po265, po266, po267, po268, po269,
    po270, po271, po272, po273, po274, po275, po276, po277, po278,
    po279, po280, po281, po282, po283, po284, po285, po286, po287,
    po288, po289, po290, po291, po292, po293, po294, po295, po296,
    po297, po298, po299, po300, po301, po302, po303, po304, po305,
    po306, po307, po308, po309, po310, po311, po312, po313, po314,
    po315, po316, po317, po318, po319, po320, po321, po322, po323,
    po324, po325, po326, po327, po328, po329, po330, po331, po332,
    po333, po334, po335, po336, po337, po338, po339, po340, po341,
    po342, po343, po344, po345, po346, po347, po348, po349, po350,
    po351, po352, po353, po354, po355, po356, po357, po358, po359,
    po360, po361, po362, po363, po364, po365, po366, po367, po368,
    po369, po370, po371, po372, po373, po374, po375, po376, po377,
    po378, po379, po380, po381, po382, po383, po384, po385, po386,
    po387, po388, po389, po390, po391, po392, po393, po394, po395,
    po396, po397, po398, po399, po400, po401, po402, po403, po404,
    po405, po406, po407, po408, po409, po410, po411, po412, po413,
    po414, po415, po416, po417, po418, po419, po420, po421, po422,
    po423, po424, po425, po426, po427, po428, po429, po430, po431,
    po432, po433, po434, po435, po436, po437, po438, po439, po440,
    po441, po442, po443, po444, po445, po446, po447, po448, po449,
    po450, po451, po452, po453, po454, po455, po456, po457, po458,
    po459, po460, po461, po462, po463, po464, po465, po466, po467,
    po468, po469, po470, po471, po472, po473, po474, po475, po476,
    po477, po478, po479, po480, po481, po482, po483, po484, po485,
    po486, po487, po488, po489, po490, po491, po492, po493, po494,
    po495, po496, po497, po498, po499, po500, po501, po502, po503,
    po504, po505, po506, po507, po508, po509, po510, po511, po512,
    po513, po514, po515, po516, po517, po518, po519, po520, po521,
    po522, po523, po524, po525, po526, po527, po528, po529, po530,
    po531, po532, po533, po534, po535, po536, po537, po538, po539,
    po540, po541, po542, po543, po544, po545, po546, po547, po548,
    po549, po550, po551, po552, po553, po554, po555, po556, po557,
    po558, po559, po560, po561, po562, po563, po564, po565, po566,
    po567, po568, po569, po570, po571, po572, po573, po574, po575,
    po576, po577, po578, po579, po580, po581, po582, po583, po584,
    po585, po586, po587, po588, po589, po590, po591, po592, po593,
    po594, po595, po596, po597, po598, po599, po600, po601, po602,
    po603, po604, po605, po606, po607, po608, po609, po610, po611,
    po612, po613, po614, po615, po616, po617, po618, po619, po620,
    po621, po622, po623, po624, po625, po626, po627, po628, po629,
    po630, po631, po632, po633, po634, po635, po636, po637, po638,
    po639, po640, po641, po642, po643, po644, po645, po646, po647,
    po648, po649, po650, po651, po652, po653, po654, po655, po656,
    po657, po658, po659, po660, po661, po662, po663, po664, po665,
    po666, po667, po668, po669, po670, po671, po672, po673, po674,
    po675, po676, po677, po678, po679, po680, po681, po682, po683,
    po684, po685, po686, po687, po688, po689, po690, po691, po692,
    po693, po694, po695, po696, po697, po698, po699, po700, po701,
    po702, po703, po704, po705, po706, po707, po708, po709, po710,
    po711, po712, po713, po714, po715, po716, po717, po718, po719,
    po720, po721, po722, po723, po724, po725, po726, po727, po728,
    po729, po730, po731, po732, po733, po734, po735, po736, po737,
    po738, po739, po740, po741, po742, po743, po744, po745, po746,
    po747, po748, po749, po750, po751, po752, po753, po754, po755,
    po756, po757, po758, po759, po760, po761, po762, po763, po764,
    po765, po766, po767, po768, po769, po770, po771, po772, po773,
    po774, po775, po776, po777, po778, po779, po780, po781, po782,
    po783, po784, po785, po786, po787, po788, po789, po790, po791,
    po792, po793, po794, po795, po796, po797, po798, po799, po800,
    po801, po802, po803, po804, po805, po806, po807, po808, po809,
    po810, po811, po812, po813, po814, po815, po816, po817, po818,
    po819, po820, po821, po822, po823, po824, po825, po826, po827,
    po828, po829, po830, po831, po832, po833, po834, po835, po836,
    po837, po838, po839, po840, po841, po842, po843, po844, po845,
    po846, po847, po848, po849, po850, po851, po852, po853, po854,
    po855, po856, po857, po858, po859, po860, po861, po862, po863,
    po864, po865, po866, po867, po868, po869, po870, po871, po872,
    po873, po874, po875, po876, po877, po878, po879, po880, po881,
    po882, po883, po884, po885, po886, po887, po888, po889, po890,
    po891, po892, po893, po894, po895, po896, po897, po898, po899,
    po900, po901, po902, po903, po904, po905, po906, po907, po908,
    po909, po910, po911, po912, po913, po914, po915, po916, po917,
    po918, po919, po920, po921, po922, po923, po924, po925, po926,
    po927, po928, po929, po930, po931, po932, po933, po934, po935,
    po936, po937, po938, po939, po940, po941, po942, po943, po944,
    po945, po946, po947, po948, po949, po950, po951, po952, po953,
    po954, po955, po956, po957, po958, po959, po960, po961, po962,
    po963, po964, po965, po966, po967, po968, po969, po970, po971,
    po972, po973, po974, po975, po976, po977, po978, po979, po980,
    po981, po982, po983, po984, po985, po986, po987, po988, po989,
    po990, po991, po992, po993, po994, po995, po996, po997, po998,
    po999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007,
    po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016,
    po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025,
    po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034,
    po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043,
    po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052,
    po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061,
    po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070,
    po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079,
    po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088,
    po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097,
    po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106,
    po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115,
    po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124,
    po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133,
    po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142,
    po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151,
    po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160,
    po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169,
    po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178,
    po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187,
    po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196,
    po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205,
    po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214,
    po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223,
    po1224, po1225, po1226, po1227, po1228, po1229, po1230  );
  input  pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7,
    pi8, pi9, pi10, pi11, pi12, pi13, pi14, pi15, pi16,
    pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25,
    pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34,
    pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43,
    pi44, pi45, pi46, pi47, pi48, pi49, pi50, pi51, pi52,
    pi53, pi54, pi55, pi56, pi57, pi58, pi59, pi60, pi61,
    pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69, pi70,
    pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79,
    pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88,
    pi89, pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97,
    pi98, pi99, pi100, pi101, pi102, pi103, pi104, pi105, pi106,
    pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115,
    pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124,
    pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133,
    pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142,
    pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151,
    pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160,
    pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187,
    pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196,
    pi197, pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205,
    pi206, pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214,
    pi215, pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223,
    pi224, pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232,
    pi233, pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241,
    pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250,
    pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259,
    pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268,
    pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277,
    pi278, pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286,
    pi287, pi288, pi289, pi290, pi291, pi292, pi293, pi294, pi295,
    pi296, pi297, pi298, pi299, pi300, pi301, pi302, pi303, pi304,
    pi305, pi306, pi307, pi308, pi309, pi310, pi311, pi312, pi313,
    pi314, pi315, pi316, pi317, pi318, pi319, pi320, pi321, pi322,
    pi323, pi324, pi325, pi326, pi327, pi328, pi329, pi330, pi331,
    pi332, pi333, pi334, pi335, pi336, pi337, pi338, pi339, pi340,
    pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349,
    pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358,
    pi359, pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367,
    pi368, pi369, pi370, pi371, pi372, pi373, pi374, pi375, pi376,
    pi377, pi378, pi379, pi380, pi381, pi382, pi383, pi384, pi385,
    pi386, pi387, pi388, pi389, pi390, pi391, pi392, pi393, pi394,
    pi395, pi396, pi397, pi398, pi399, pi400, pi401, pi402, pi403,
    pi404, pi405, pi406, pi407, pi408, pi409, pi410, pi411, pi412,
    pi413, pi414, pi415, pi416, pi417, pi418, pi419, pi420, pi421,
    pi422, pi423, pi424, pi425, pi426, pi427, pi428, pi429, pi430,
    pi431, pi432, pi433, pi434, pi435, pi436, pi437, pi438, pi439,
    pi440, pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448,
    pi449, pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457,
    pi458, pi459, pi460, pi461, pi462, pi463, pi464, pi465, pi466,
    pi467, pi468, pi469, pi470, pi471, pi472, pi473, pi474, pi475,
    pi476, pi477, pi478, pi479, pi480, pi481, pi482, pi483, pi484,
    pi485, pi486, pi487, pi488, pi489, pi490, pi491, pi492, pi493,
    pi494, pi495, pi496, pi497, pi498, pi499, pi500, pi501, pi502,
    pi503, pi504, pi505, pi506, pi507, pi508, pi509, pi510, pi511,
    pi512, pi513, pi514, pi515, pi516, pi517, pi518, pi519, pi520,
    pi521, pi522, pi523, pi524, pi525, pi526, pi527, pi528, pi529,
    pi530, pi531, pi532, pi533, pi534, pi535, pi536, pi537, pi538,
    pi539, pi540, pi541, pi542, pi543, pi544, pi545, pi546, pi547,
    pi548, pi549, pi550, pi551, pi552, pi553, pi554, pi555, pi556,
    pi557, pi558, pi559, pi560, pi561, pi562, pi563, pi564, pi565,
    pi566, pi567, pi568, pi569, pi570, pi571, pi572, pi573, pi574,
    pi575, pi576, pi577, pi578, pi579, pi580, pi581, pi582, pi583,
    pi584, pi585, pi586, pi587, pi588, pi589, pi590, pi591, pi592,
    pi593, pi594, pi595, pi596, pi597, pi598, pi599, pi600, pi601,
    pi602, pi603, pi604, pi605, pi606, pi607, pi608, pi609, pi610,
    pi611, pi612, pi613, pi614, pi615, pi616, pi617, pi618, pi619,
    pi620, pi621, pi622, pi623, pi624, pi625, pi626, pi627, pi628,
    pi629, pi630, pi631, pi632, pi633, pi634, pi635, pi636, pi637,
    pi638, pi639, pi640, pi641, pi642, pi643, pi644, pi645, pi646,
    pi647, pi648, pi649, pi650, pi651, pi652, pi653, pi654, pi655,
    pi656, pi657, pi658, pi659, pi660, pi661, pi662, pi663, pi664,
    pi665, pi666, pi667, pi668, pi669, pi670, pi671, pi672, pi673,
    pi674, pi675, pi676, pi677, pi678, pi679, pi680, pi681, pi682,
    pi683, pi684, pi685, pi686, pi687, pi688, pi689, pi690, pi691,
    pi692, pi693, pi694, pi695, pi696, pi697, pi698, pi699, pi700,
    pi701, pi702, pi703, pi704, pi705, pi706, pi707, pi708, pi709,
    pi710, pi711, pi712, pi713, pi714, pi715, pi716, pi717, pi718,
    pi719, pi720, pi721, pi722, pi723, pi724, pi725, pi726, pi727,
    pi728, pi729, pi730, pi731, pi732, pi733, pi734, pi735, pi736,
    pi737, pi738, pi739, pi740, pi741, pi742, pi743, pi744, pi745,
    pi746, pi747, pi748, pi749, pi750, pi751, pi752, pi753, pi754,
    pi755, pi756, pi757, pi758, pi759, pi760, pi761, pi762, pi763,
    pi764, pi765, pi766, pi767, pi768, pi769, pi770, pi771, pi772,
    pi773, pi774, pi775, pi776, pi777, pi778, pi779, pi780, pi781,
    pi782, pi783, pi784, pi785, pi786, pi787, pi788, pi789, pi790,
    pi791, pi792, pi793, pi794, pi795, pi796, pi797, pi798, pi799,
    pi800, pi801, pi802, pi803, pi804, pi805, pi806, pi807, pi808,
    pi809, pi810, pi811, pi812, pi813, pi814, pi815, pi816, pi817,
    pi818, pi819, pi820, pi821, pi822, pi823, pi824, pi825, pi826,
    pi827, pi828, pi829, pi830, pi831, pi832, pi833, pi834, pi835,
    pi836, pi837, pi838, pi839, pi840, pi841, pi842, pi843, pi844,
    pi845, pi846, pi847, pi848, pi849, pi850, pi851, pi852, pi853,
    pi854, pi855, pi856, pi857, pi858, pi859, pi860, pi861, pi862,
    pi863, pi864, pi865, pi866, pi867, pi868, pi869, pi870, pi871,
    pi872, pi873, pi874, pi875, pi876, pi877, pi878, pi879, pi880,
    pi881, pi882, pi883, pi884, pi885, pi886, pi887, pi888, pi889,
    pi890, pi891, pi892, pi893, pi894, pi895, pi896, pi897, pi898,
    pi899, pi900, pi901, pi902, pi903, pi904, pi905, pi906, pi907,
    pi908, pi909, pi910, pi911, pi912, pi913, pi914, pi915, pi916,
    pi917, pi918, pi919, pi920, pi921, pi922, pi923, pi924, pi925,
    pi926, pi927, pi928, pi929, pi930, pi931, pi932, pi933, pi934,
    pi935, pi936, pi937, pi938, pi939, pi940, pi941, pi942, pi943,
    pi944, pi945, pi946, pi947, pi948, pi949, pi950, pi951, pi952,
    pi953, pi954, pi955, pi956, pi957, pi958, pi959, pi960, pi961,
    pi962, pi963, pi964, pi965, pi966, pi967, pi968, pi969, pi970,
    pi971, pi972, pi973, pi974, pi975, pi976, pi977, pi978, pi979,
    pi980, pi981, pi982, pi983, pi984, pi985, pi986, pi987, pi988,
    pi989, pi990, pi991, pi992, pi993, pi994, pi995, pi996, pi997,
    pi998, pi999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006,
    pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015,
    pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024,
    pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033,
    pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042,
    pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051,
    pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060,
    pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069,
    pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078,
    pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087,
    pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096,
    pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105,
    pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114,
    pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123,
    pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132,
    pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141,
    pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150,
    pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159,
    pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168,
    pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177,
    pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186,
    pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195,
    pi1196, pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203;
  output po0, po1, po2, po3, po4, po5, po6, po7,
    po8, po9, po10, po11, po12, po13, po14, po15, po16,
    po17, po18, po19, po20, po21, po22, po23, po24, po25,
    po26, po27, po28, po29, po30, po31, po32, po33, po34,
    po35, po36, po37, po38, po39, po40, po41, po42, po43,
    po44, po45, po46, po47, po48, po49, po50, po51, po52,
    po53, po54, po55, po56, po57, po58, po59, po60, po61,
    po62, po63, po64, po65, po66, po67, po68, po69, po70,
    po71, po72, po73, po74, po75, po76, po77, po78, po79,
    po80, po81, po82, po83, po84, po85, po86, po87, po88,
    po89, po90, po91, po92, po93, po94, po95, po96, po97,
    po98, po99, po100, po101, po102, po103, po104, po105, po106,
    po107, po108, po109, po110, po111, po112, po113, po114, po115,
    po116, po117, po118, po119, po120, po121, po122, po123, po124,
    po125, po126, po127, po128, po129, po130, po131, po132, po133,
    po134, po135, po136, po137, po138, po139, po140, po141, po142,
    po143, po144, po145, po146, po147, po148, po149, po150, po151,
    po152, po153, po154, po155, po156, po157, po158, po159, po160,
    po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178,
    po179, po180, po181, po182, po183, po184, po185, po186, po187,
    po188, po189, po190, po191, po192, po193, po194, po195, po196,
    po197, po198, po199, po200, po201, po202, po203, po204, po205,
    po206, po207, po208, po209, po210, po211, po212, po213, po214,
    po215, po216, po217, po218, po219, po220, po221, po222, po223,
    po224, po225, po226, po227, po228, po229, po230, po231, po232,
    po233, po234, po235, po236, po237, po238, po239, po240, po241,
    po242, po243, po244, po245, po246, po247, po248, po249, po250,
    po251, po252, po253, po254, po255, po256, po257, po258, po259,
    po260, po261, po262, po263, po264, po265, po266, po267, po268,
    po269, po270, po271, po272, po273, po274, po275, po276, po277,
    po278, po279, po280, po281, po282, po283, po284, po285, po286,
    po287, po288, po289, po290, po291, po292, po293, po294, po295,
    po296, po297, po298, po299, po300, po301, po302, po303, po304,
    po305, po306, po307, po308, po309, po310, po311, po312, po313,
    po314, po315, po316, po317, po318, po319, po320, po321, po322,
    po323, po324, po325, po326, po327, po328, po329, po330, po331,
    po332, po333, po334, po335, po336, po337, po338, po339, po340,
    po341, po342, po343, po344, po345, po346, po347, po348, po349,
    po350, po351, po352, po353, po354, po355, po356, po357, po358,
    po359, po360, po361, po362, po363, po364, po365, po366, po367,
    po368, po369, po370, po371, po372, po373, po374, po375, po376,
    po377, po378, po379, po380, po381, po382, po383, po384, po385,
    po386, po387, po388, po389, po390, po391, po392, po393, po394,
    po395, po396, po397, po398, po399, po400, po401, po402, po403,
    po404, po405, po406, po407, po408, po409, po410, po411, po412,
    po413, po414, po415, po416, po417, po418, po419, po420, po421,
    po422, po423, po424, po425, po426, po427, po428, po429, po430,
    po431, po432, po433, po434, po435, po436, po437, po438, po439,
    po440, po441, po442, po443, po444, po445, po446, po447, po448,
    po449, po450, po451, po452, po453, po454, po455, po456, po457,
    po458, po459, po460, po461, po462, po463, po464, po465, po466,
    po467, po468, po469, po470, po471, po472, po473, po474, po475,
    po476, po477, po478, po479, po480, po481, po482, po483, po484,
    po485, po486, po487, po488, po489, po490, po491, po492, po493,
    po494, po495, po496, po497, po498, po499, po500, po501, po502,
    po503, po504, po505, po506, po507, po508, po509, po510, po511,
    po512, po513, po514, po515, po516, po517, po518, po519, po520,
    po521, po522, po523, po524, po525, po526, po527, po528, po529,
    po530, po531, po532, po533, po534, po535, po536, po537, po538,
    po539, po540, po541, po542, po543, po544, po545, po546, po547,
    po548, po549, po550, po551, po552, po553, po554, po555, po556,
    po557, po558, po559, po560, po561, po562, po563, po564, po565,
    po566, po567, po568, po569, po570, po571, po572, po573, po574,
    po575, po576, po577, po578, po579, po580, po581, po582, po583,
    po584, po585, po586, po587, po588, po589, po590, po591, po592,
    po593, po594, po595, po596, po597, po598, po599, po600, po601,
    po602, po603, po604, po605, po606, po607, po608, po609, po610,
    po611, po612, po613, po614, po615, po616, po617, po618, po619,
    po620, po621, po622, po623, po624, po625, po626, po627, po628,
    po629, po630, po631, po632, po633, po634, po635, po636, po637,
    po638, po639, po640, po641, po642, po643, po644, po645, po646,
    po647, po648, po649, po650, po651, po652, po653, po654, po655,
    po656, po657, po658, po659, po660, po661, po662, po663, po664,
    po665, po666, po667, po668, po669, po670, po671, po672, po673,
    po674, po675, po676, po677, po678, po679, po680, po681, po682,
    po683, po684, po685, po686, po687, po688, po689, po690, po691,
    po692, po693, po694, po695, po696, po697, po698, po699, po700,
    po701, po702, po703, po704, po705, po706, po707, po708, po709,
    po710, po711, po712, po713, po714, po715, po716, po717, po718,
    po719, po720, po721, po722, po723, po724, po725, po726, po727,
    po728, po729, po730, po731, po732, po733, po734, po735, po736,
    po737, po738, po739, po740, po741, po742, po743, po744, po745,
    po746, po747, po748, po749, po750, po751, po752, po753, po754,
    po755, po756, po757, po758, po759, po760, po761, po762, po763,
    po764, po765, po766, po767, po768, po769, po770, po771, po772,
    po773, po774, po775, po776, po777, po778, po779, po780, po781,
    po782, po783, po784, po785, po786, po787, po788, po789, po790,
    po791, po792, po793, po794, po795, po796, po797, po798, po799,
    po800, po801, po802, po803, po804, po805, po806, po807, po808,
    po809, po810, po811, po812, po813, po814, po815, po816, po817,
    po818, po819, po820, po821, po822, po823, po824, po825, po826,
    po827, po828, po829, po830, po831, po832, po833, po834, po835,
    po836, po837, po838, po839, po840, po841, po842, po843, po844,
    po845, po846, po847, po848, po849, po850, po851, po852, po853,
    po854, po855, po856, po857, po858, po859, po860, po861, po862,
    po863, po864, po865, po866, po867, po868, po869, po870, po871,
    po872, po873, po874, po875, po876, po877, po878, po879, po880,
    po881, po882, po883, po884, po885, po886, po887, po888, po889,
    po890, po891, po892, po893, po894, po895, po896, po897, po898,
    po899, po900, po901, po902, po903, po904, po905, po906, po907,
    po908, po909, po910, po911, po912, po913, po914, po915, po916,
    po917, po918, po919, po920, po921, po922, po923, po924, po925,
    po926, po927, po928, po929, po930, po931, po932, po933, po934,
    po935, po936, po937, po938, po939, po940, po941, po942, po943,
    po944, po945, po946, po947, po948, po949, po950, po951, po952,
    po953, po954, po955, po956, po957, po958, po959, po960, po961,
    po962, po963, po964, po965, po966, po967, po968, po969, po970,
    po971, po972, po973, po974, po975, po976, po977, po978, po979,
    po980, po981, po982, po983, po984, po985, po986, po987, po988,
    po989, po990, po991, po992, po993, po994, po995, po996, po997,
    po998, po999, po1000, po1001, po1002, po1003, po1004, po1005, po1006,
    po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015,
    po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024,
    po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033,
    po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042,
    po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051,
    po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060,
    po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069,
    po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078,
    po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087,
    po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096,
    po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105,
    po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114,
    po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123,
    po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132,
    po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141,
    po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150,
    po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159,
    po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168,
    po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177,
    po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186,
    po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195,
    po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204,
    po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213,
    po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222,
    po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230;
  wire n2437, n2438, n2439, n2440, n2441, n2442,
    n2443, n2444, n2445, n2446, n2447, n2448,
    n2449, n2450, n2451, n2452, n2453, n2454,
    n2455, n2456, n2457, n2458, n2459, n2460,
    n2461, n2462, n2463, n2464, n2465, n2466,
    n2467, n2468, n2469, n2470, n2471, n2472,
    n2473, n2474, n2475, n2476, n2477, n2478,
    n2479, n2480, n2481, n2482, n2483, n2484,
    n2485, n2486, n2487, n2488, n2489, n2490,
    n2491, n2492, n2493, n2494, n2495, n2496,
    n2497, n2498, n2499, n2500, n2501, n2502,
    n2503, n2504, n2505, n2506, n2507, n2508,
    n2509, n2510, n2511, n2512, n2513, n2514,
    n2515, n2516, n2517, n2518, n2519, n2520,
    n2521, n2522, n2523, n2524, n2525, n2526,
    n2527, n2528, n2529, n2530, n2531, n2532,
    n2533, n2534, n2535, n2536, n2537, n2538,
    n2539, n2540, n2541, n2542, n2543, n2544,
    n2545, n2546, n2547, n2548, n2549, n2550,
    n2551, n2552, n2553, n2554, n2555, n2556,
    n2557, n2558, n2559, n2560, n2561, n2562,
    n2563, n2564, n2565, n2566, n2567, n2568,
    n2569, n2570, n2571, n2572, n2573, n2574,
    n2575, n2576, n2577, n2578, n2579, n2580,
    n2581, n2582, n2583, n2584, n2585, n2586,
    n2587, n2588, n2589, n2590, n2591, n2592,
    n2593, n2594, n2595, n2596, n2597, n2598,
    n2599, n2600, n2601, n2602, n2603, n2604,
    n2605, n2606, n2607, n2608, n2609, n2610,
    n2611, n2612, n2613, n2614, n2615, n2616,
    n2617, n2618, n2619, n2620, n2621, n2622,
    n2623, n2624, n2625, n2626, n2627, n2628,
    n2629, n2630, n2631, n2632, n2633, n2634,
    n2635, n2636, n2637, n2638, n2639, n2640,
    n2641, n2642, n2643, n2644, n2645, n2646,
    n2647, n2648, n2649, n2650, n2651, n2652,
    n2653, n2654, n2655, n2656, n2657, n2658,
    n2659, n2660, n2661, n2662, n2663, n2664,
    n2665, n2666, n2667, n2668, n2669, n2670,
    n2671, n2672, n2673, n2674, n2675, n2676,
    n2677, n2678, n2679, n2680, n2681, n2682,
    n2683, n2684, n2685, n2686, n2687, n2688,
    n2689, n2690, n2691, n2692, n2693, n2694,
    n2695, n2696, n2697, n2698, n2699, n2700,
    n2701, n2702, n2703, n2704, n2705, n2706,
    n2707, n2708, n2709, n2710, n2711, n2712,
    n2713, n2714, n2715, n2716, n2717, n2718,
    n2719, n2720, n2721, n2722, n2723, n2724,
    n2725, n2726, n2727, n2728, n2729, n2730,
    n2731, n2732, n2733, n2734, n2735, n2736,
    n2737, n2738, n2739, n2740, n2741, n2742,
    n2743, n2744, n2745, n2746, n2747, n2748,
    n2749, n2750, n2751, n2752, n2753, n2754,
    n2755, n2756, n2757, n2758, n2759, n2760,
    n2761, n2762, n2763, n2764, n2765, n2766,
    n2767, n2768, n2769, n2770, n2771, n2772,
    n2773, n2774, n2775, n2776, n2777, n2778,
    n2779, n2780, n2781, n2782, n2783, n2784,
    n2785, n2786, n2787, n2788, n2789, n2790,
    n2791, n2792, n2793, n2794, n2795, n2796,
    n2797, n2798, n2799, n2800, n2801, n2802,
    n2803, n2804, n2805, n2806, n2807, n2808,
    n2809, n2810, n2811, n2812, n2813, n2814,
    n2815, n2816, n2817, n2818, n2819, n2820,
    n2821, n2822, n2823, n2824, n2825, n2826,
    n2827, n2828, n2829, n2830, n2831, n2832,
    n2833, n2834, n2835, n2836, n2837, n2838,
    n2839, n2840, n2841, n2842, n2843, n2844,
    n2845, n2846, n2847, n2848, n2849, n2850,
    n2851, n2852, n2853, n2854, n2855, n2856,
    n2857, n2858, n2859, n2860, n2861, n2862,
    n2863, n2864, n2865, n2866, n2867, n2868,
    n2869, n2870, n2871, n2872, n2873, n2874,
    n2875, n2876, n2877, n2878, n2879, n2880,
    n2881, n2882, n2883, n2884, n2885, n2886,
    n2887, n2888, n2889, n2890, n2891, n2892,
    n2893, n2894, n2895, n2896, n2897, n2898,
    n2899, n2900, n2901, n2902, n2903, n2904,
    n2905, n2906, n2907, n2908, n2909, n2910,
    n2911, n2912, n2913, n2914, n2915, n2916,
    n2917, n2918, n2919, n2920, n2921, n2922,
    n2923, n2924, n2925, n2926, n2927, n2928,
    n2929, n2930, n2931, n2932, n2933, n2934,
    n2935, n2936, n2937, n2938, n2939, n2940,
    n2941, n2942, n2943, n2944, n2945, n2946,
    n2947, n2948, n2949, n2950, n2951, n2952,
    n2953, n2954, n2955, n2956, n2957, n2958,
    n2959, n2960, n2961, n2962, n2963, n2964,
    n2965, n2966, n2967, n2968, n2969, n2970,
    n2971, n2972, n2973, n2974, n2975, n2976,
    n2977, n2978, n2979, n2980, n2981, n2982,
    n2983, n2984, n2985, n2986, n2987, n2988,
    n2989, n2990, n2991, n2992, n2993, n2994,
    n2995, n2996, n2997, n2998, n2999, n3000,
    n3001, n3002, n3003, n3004, n3005, n3006,
    n3007, n3008, n3009, n3010, n3011, n3012,
    n3013, n3014, n3015, n3016, n3017, n3018,
    n3019, n3020, n3021, n3022, n3023, n3024,
    n3025, n3026, n3027, n3028, n3029, n3030,
    n3031, n3032, n3033, n3034, n3035, n3036,
    n3037, n3038, n3039, n3040, n3041, n3042,
    n3043, n3044, n3045, n3046, n3047, n3048,
    n3049, n3050, n3051, n3052, n3053, n3054,
    n3055, n3056, n3057, n3058, n3059, n3060,
    n3061, n3062, n3063, n3064, n3065, n3066,
    n3067, n3068, n3069, n3070, n3071, n3072,
    n3073, n3074, n3075, n3076, n3077, n3078,
    n3079, n3080, n3081, n3082, n3083, n3084,
    n3085, n3086, n3087, n3088, n3089, n3090,
    n3091, n3092, n3093, n3094, n3095, n3096,
    n3097, n3098, n3099, n3100, n3101, n3102,
    n3103, n3104, n3105, n3106, n3107, n3108,
    n3109, n3110, n3111, n3112, n3113, n3114,
    n3115, n3116, n3117, n3118, n3119, n3120,
    n3121, n3122, n3123, n3124, n3125, n3126,
    n3127, n3128, n3129, n3130, n3131, n3132,
    n3133, n3134, n3135, n3136, n3137, n3138,
    n3139, n3140, n3141, n3142, n3143, n3144,
    n3145, n3146, n3147, n3148, n3149, n3150,
    n3151, n3152, n3153, n3154, n3155, n3156,
    n3157, n3158, n3159, n3160, n3161, n3162,
    n3163, n3164, n3165, n3166, n3167, n3168,
    n3169, n3170, n3171, n3172, n3173, n3174,
    n3175, n3176, n3177, n3178, n3179, n3180,
    n3181, n3182, n3183, n3184, n3185, n3186,
    n3187, n3188, n3189, n3190, n3191, n3192,
    n3193, n3194, n3195, n3196, n3197, n3198,
    n3199, n3200, n3201, n3202, n3203, n3204,
    n3205, n3206, n3207, n3208, n3209, n3210,
    n3211, n3212, n3213, n3214, n3215, n3216,
    n3217, n3218, n3219, n3220, n3221, n3222,
    n3223, n3224, n3225, n3226, n3227, n3228,
    n3229, n3230, n3231, n3232, n3233, n3234,
    n3235, n3236, n3237, n3238, n3239, n3240,
    n3241, n3242, n3243, n3244, n3245, n3246,
    n3247, n3248, n3249, n3250, n3251, n3252,
    n3253, n3254, n3255, n3256, n3257, n3258,
    n3259, n3260, n3261, n3262, n3263, n3264,
    n3265, n3266, n3267, n3268, n3269, n3270,
    n3271, n3272, n3273, n3274, n3275, n3276,
    n3277, n3278, n3279, n3280, n3281, n3282,
    n3283, n3284, n3285, n3286, n3287, n3288,
    n3289, n3290, n3291, n3292, n3293, n3294,
    n3295, n3296, n3297, n3299, n3300, n3301,
    n3302, n3303, n3304, n3305, n3306, n3307,
    n3308, n3309, n3310, n3311, n3312, n3313,
    n3314, n3315, n3316, n3317, n3318, n3319,
    n3320, n3321, n3322, n3323, n3324, n3325,
    n3326, n3327, n3328, n3329, n3330, n3331,
    n3332, n3333, n3334, n3335, n3336, n3337,
    n3338, n3339, n3340, n3341, n3342, n3343,
    n3344, n3345, n3346, n3347, n3348, n3349,
    n3350, n3351, n3352, n3353, n3354, n3355,
    n3356, n3357, n3358, n3359, n3360, n3361,
    n3362, n3363, n3364, n3365, n3366, n3367,
    n3368, n3369, n3370, n3371, n3372, n3373,
    n3374, n3375, n3376, n3377, n3378, n3379,
    n3380, n3381, n3382, n3383, n3384, n3385,
    n3386, n3387, n3388, n3389, n3390, n3391,
    n3392, n3393, n3394, n3395, n3396, n3397,
    n3398, n3399, n3400, n3401, n3402, n3403,
    n3404, n3405, n3406, n3407, n3408, n3409,
    n3410, n3411, n3412, n3413, n3414, n3415,
    n3416, n3417, n3418, n3419, n3420, n3421,
    n3422, n3423, n3424, n3425, n3426, n3427,
    n3428, n3429, n3430, n3431, n3432, n3433,
    n3434, n3435, n3436, n3437, n3438, n3439,
    n3440, n3441, n3442, n3443, n3444, n3445,
    n3446, n3447, n3448, n3449, n3450, n3451,
    n3452, n3453, n3454, n3455, n3456, n3457,
    n3458, n3459, n3460, n3461, n3462, n3463,
    n3464, n3465, n3466, n3467, n3468, n3469,
    n3470, n3471, n3472, n3473, n3474, n3475,
    n3476, n3477, n3478, n3479, n3480, n3481,
    n3482, n3483, n3484, n3485, n3486, n3487,
    n3488, n3489, n3490, n3491, n3492, n3493,
    n3494, n3495, n3496, n3497, n3498, n3499,
    n3500, n3501, n3502, n3503, n3504, n3505,
    n3506, n3507, n3508, n3509, n3510, n3511,
    n3512, n3513, n3514, n3515, n3516, n3518,
    n3519, n3520, n3521, n3522, n3523, n3524,
    n3525, n3526, n3527, n3528, n3529, n3530,
    n3531, n3532, n3533, n3534, n3535, n3536,
    n3537, n3538, n3539, n3540, n3541, n3542,
    n3543, n3544, n3545, n3546, n3547, n3548,
    n3549, n3550, n3551, n3552, n3553, n3554,
    n3555, n3556, n3557, n3558, n3559, n3560,
    n3561, n3562, n3563, n3564, n3565, n3566,
    n3567, n3568, n3569, n3570, n3571, n3572,
    n3573, n3574, n3575, n3576, n3577, n3578,
    n3579, n3580, n3581, n3582, n3583, n3584,
    n3585, n3586, n3587, n3588, n3589, n3590,
    n3591, n3592, n3593, n3594, n3595, n3596,
    n3597, n3598, n3599, n3600, n3601, n3602,
    n3603, n3604, n3605, n3606, n3607, n3608,
    n3609, n3610, n3611, n3612, n3613, n3614,
    n3615, n3616, n3617, n3618, n3619, n3620,
    n3621, n3622, n3623, n3624, n3625, n3626,
    n3627, n3628, n3629, n3630, n3631, n3632,
    n3633, n3634, n3635, n3636, n3637, n3638,
    n3639, n3640, n3641, n3642, n3643, n3644,
    n3645, n3646, n3647, n3648, n3649, n3650,
    n3651, n3652, n3653, n3654, n3655, n3656,
    n3657, n3658, n3659, n3660, n3661, n3662,
    n3663, n3664, n3665, n3666, n3667, n3668,
    n3669, n3670, n3671, n3672, n3673, n3674,
    n3675, n3676, n3677, n3678, n3679, n3680,
    n3681, n3682, n3683, n3684, n3685, n3686,
    n3687, n3688, n3689, n3691, n3692, n3693,
    n3694, n3695, n3696, n3697, n3698, n3699,
    n3700, n3701, n3702, n3703, n3704, n3705,
    n3706, n3707, n3708, n3709, n3710, n3711,
    n3712, n3713, n3714, n3715, n3716, n3717,
    n3718, n3719, n3720, n3721, n3722, n3723,
    n3724, n3725, n3726, n3727, n3728, n3729,
    n3730, n3731, n3732, n3733, n3734, n3735,
    n3736, n3737, n3738, n3739, n3740, n3741,
    n3742, n3743, n3744, n3745, n3746, n3747,
    n3748, n3749, n3750, n3751, n3752, n3753,
    n3754, n3755, n3756, n3757, n3758, n3759,
    n3760, n3761, n3762, n3763, n3764, n3765,
    n3766, n3767, n3768, n3769, n3770, n3771,
    n3772, n3773, n3774, n3775, n3776, n3777,
    n3778, n3779, n3780, n3781, n3782, n3783,
    n3784, n3785, n3786, n3787, n3788, n3789,
    n3790, n3791, n3792, n3793, n3794, n3795,
    n3796, n3797, n3798, n3799, n3800, n3801,
    n3802, n3803, n3804, n3805, n3806, n3807,
    n3808, n3809, n3810, n3811, n3812, n3813,
    n3814, n3815, n3816, n3817, n3818, n3819,
    n3820, n3821, n3822, n3823, n3824, n3825,
    n3826, n3827, n3828, n3829, n3830, n3831,
    n3832, n3833, n3834, n3835, n3836, n3837,
    n3838, n3839, n3840, n3841, n3842, n3843,
    n3844, n3845, n3846, n3847, n3848, n3849,
    n3850, n3851, n3852, n3853, n3854, n3855,
    n3856, n3857, n3858, n3859, n3860, n3861,
    n3862, n3863, n3864, n3865, n3866, n3867,
    n3868, n3869, n3870, n3871, n3872, n3873,
    n3874, n3875, n3876, n3877, n3878, n3879,
    n3880, n3881, n3882, n3883, n3884, n3885,
    n3886, n3887, n3888, n3889, n3890, n3891,
    n3892, n3893, n3894, n3895, n3896, n3897,
    n3898, n3899, n3900, n3901, n3902, n3903,
    n3904, n3905, n3906, n3907, n3908, n3909,
    n3910, n3911, n3912, n3913, n3914, n3915,
    n3916, n3917, n3918, n3920, n3921, n3922,
    n3923, n3924, n3925, n3926, n3927, n3928,
    n3929, n3930, n3931, n3932, n3933, n3934,
    n3935, n3936, n3937, n3938, n3939, n3940,
    n3941, n3942, n3943, n3944, n3945, n3946,
    n3947, n3948, n3949, n3950, n3951, n3952,
    n3953, n3954, n3955, n3956, n3957, n3958,
    n3959, n3960, n3961, n3962, n3963, n3964,
    n3965, n3966, n3967, n3968, n3969, n3970,
    n3971, n3972, n3973, n3974, n3975, n3976,
    n3977, n3978, n3979, n3980, n3981, n3982,
    n3983, n3984, n3985, n3986, n3987, n3988,
    n3989, n3990, n3991, n3992, n3993, n3994,
    n3995, n3996, n3997, n3998, n3999, n4000,
    n4001, n4002, n4003, n4004, n4005, n4006,
    n4007, n4008, n4009, n4010, n4011, n4012,
    n4013, n4014, n4015, n4016, n4017, n4018,
    n4019, n4020, n4021, n4022, n4023, n4024,
    n4025, n4026, n4027, n4028, n4029, n4030,
    n4031, n4032, n4033, n4034, n4035, n4036,
    n4037, n4038, n4039, n4040, n4041, n4042,
    n4043, n4044, n4045, n4046, n4047, n4048,
    n4049, n4050, n4051, n4052, n4053, n4054,
    n4055, n4056, n4057, n4058, n4059, n4060,
    n4061, n4062, n4063, n4064, n4065, n4066,
    n4067, n4068, n4069, n4070, n4071, n4072,
    n4073, n4074, n4075, n4076, n4077, n4078,
    n4079, n4080, n4081, n4082, n4083, n4084,
    n4085, n4086, n4087, n4088, n4089, n4090,
    n4091, n4092, n4093, n4094, n4095, n4096,
    n4097, n4098, n4099, n4100, n4101, n4102,
    n4103, n4104, n4105, n4106, n4107, n4108,
    n4109, n4110, n4111, n4112, n4113, n4114,
    n4115, n4116, n4117, n4118, n4119, n4120,
    n4121, n4122, n4123, n4124, n4125, n4126,
    n4127, n4128, n4129, n4130, n4131, n4132,
    n4133, n4134, n4135, n4136, n4137, n4138,
    n4139, n4140, n4141, n4142, n4143, n4144,
    n4145, n4147, n4148, n4149, n4150, n4151,
    n4152, n4153, n4154, n4155, n4156, n4157,
    n4158, n4159, n4160, n4161, n4162, n4163,
    n4164, n4165, n4166, n4167, n4168, n4169,
    n4170, n4171, n4172, n4173, n4174, n4175,
    n4176, n4177, n4178, n4179, n4180, n4181,
    n4182, n4183, n4184, n4185, n4186, n4187,
    n4188, n4189, n4190, n4191, n4192, n4193,
    n4194, n4195, n4196, n4197, n4198, n4199,
    n4200, n4201, n4202, n4203, n4204, n4205,
    n4206, n4207, n4208, n4209, n4210, n4211,
    n4212, n4213, n4214, n4215, n4216, n4217,
    n4218, n4219, n4220, n4221, n4222, n4223,
    n4224, n4225, n4226, n4227, n4228, n4229,
    n4230, n4231, n4232, n4233, n4234, n4235,
    n4236, n4237, n4238, n4239, n4240, n4241,
    n4242, n4243, n4244, n4245, n4246, n4247,
    n4248, n4249, n4250, n4251, n4252, n4253,
    n4254, n4255, n4256, n4257, n4258, n4259,
    n4260, n4261, n4262, n4263, n4264, n4265,
    n4266, n4267, n4268, n4269, n4270, n4271,
    n4272, n4273, n4274, n4275, n4276, n4277,
    n4278, n4279, n4280, n4281, n4282, n4283,
    n4284, n4285, n4286, n4287, n4288, n4289,
    n4290, n4291, n4292, n4293, n4294, n4295,
    n4296, n4297, n4298, n4299, n4300, n4301,
    n4302, n4303, n4304, n4305, n4306, n4307,
    n4308, n4309, n4310, n4311, n4312, n4313,
    n4314, n4315, n4316, n4317, n4318, n4319,
    n4320, n4321, n4322, n4323, n4324, n4325,
    n4326, n4327, n4328, n4329, n4330, n4331,
    n4332, n4333, n4334, n4335, n4336, n4337,
    n4338, n4339, n4340, n4341, n4342, n4343,
    n4344, n4345, n4346, n4347, n4348, n4349,
    n4350, n4351, n4352, n4353, n4354, n4355,
    n4356, n4357, n4358, n4359, n4360, n4361,
    n4362, n4363, n4364, n4365, n4366, n4367,
    n4369, n4370, n4371, n4372, n4373, n4374,
    n4375, n4376, n4377, n4378, n4379, n4380,
    n4381, n4382, n4383, n4384, n4385, n4386,
    n4387, n4388, n4389, n4390, n4391, n4392,
    n4393, n4394, n4395, n4396, n4397, n4398,
    n4399, n4400, n4401, n4402, n4403, n4404,
    n4405, n4406, n4407, n4408, n4409, n4410,
    n4411, n4412, n4413, n4414, n4415, n4416,
    n4417, n4418, n4419, n4420, n4421, n4422,
    n4423, n4424, n4425, n4426, n4427, n4428,
    n4429, n4430, n4431, n4432, n4433, n4434,
    n4435, n4436, n4437, n4438, n4439, n4440,
    n4441, n4442, n4443, n4444, n4445, n4446,
    n4447, n4448, n4449, n4450, n4451, n4452,
    n4453, n4454, n4455, n4456, n4457, n4458,
    n4459, n4460, n4461, n4462, n4463, n4464,
    n4465, n4466, n4467, n4468, n4469, n4470,
    n4471, n4472, n4473, n4474, n4475, n4476,
    n4477, n4478, n4479, n4480, n4481, n4482,
    n4483, n4484, n4485, n4486, n4487, n4488,
    n4489, n4490, n4491, n4492, n4493, n4494,
    n4495, n4496, n4497, n4498, n4499, n4500,
    n4501, n4502, n4503, n4504, n4505, n4506,
    n4507, n4508, n4509, n4510, n4511, n4512,
    n4513, n4514, n4515, n4516, n4517, n4518,
    n4519, n4520, n4521, n4522, n4523, n4524,
    n4525, n4526, n4527, n4528, n4529, n4530,
    n4531, n4532, n4533, n4534, n4535, n4536,
    n4537, n4538, n4539, n4540, n4541, n4542,
    n4543, n4544, n4545, n4546, n4547, n4548,
    n4549, n4550, n4551, n4552, n4553, n4554,
    n4555, n4556, n4557, n4558, n4559, n4560,
    n4561, n4562, n4563, n4564, n4565, n4566,
    n4567, n4568, n4569, n4570, n4571, n4572,
    n4573, n4574, n4575, n4576, n4577, n4578,
    n4579, n4580, n4581, n4582, n4583, n4584,
    n4585, n4586, n4587, n4588, n4589, n4591,
    n4592, n4593, n4594, n4595, n4596, n4597,
    n4598, n4599, n4600, n4601, n4602, n4603,
    n4604, n4605, n4606, n4607, n4608, n4609,
    n4610, n4611, n4612, n4613, n4614, n4615,
    n4616, n4617, n4618, n4619, n4620, n4621,
    n4622, n4623, n4624, n4625, n4626, n4627,
    n4628, n4629, n4630, n4631, n4632, n4633,
    n4634, n4635, n4636, n4637, n4638, n4639,
    n4640, n4641, n4642, n4643, n4644, n4645,
    n4646, n4647, n4648, n4649, n4650, n4651,
    n4652, n4653, n4654, n4655, n4656, n4657,
    n4658, n4659, n4660, n4661, n4662, n4663,
    n4664, n4665, n4666, n4667, n4668, n4669,
    n4670, n4671, n4672, n4673, n4674, n4675,
    n4676, n4677, n4678, n4679, n4680, n4681,
    n4682, n4683, n4684, n4685, n4686, n4687,
    n4688, n4689, n4690, n4691, n4692, n4693,
    n4694, n4695, n4696, n4697, n4698, n4699,
    n4700, n4701, n4702, n4703, n4704, n4705,
    n4706, n4707, n4708, n4709, n4710, n4711,
    n4712, n4713, n4714, n4715, n4716, n4717,
    n4718, n4719, n4720, n4721, n4722, n4723,
    n4724, n4725, n4726, n4727, n4728, n4729,
    n4730, n4731, n4732, n4733, n4734, n4735,
    n4736, n4737, n4738, n4739, n4740, n4741,
    n4742, n4743, n4744, n4745, n4746, n4747,
    n4748, n4749, n4750, n4751, n4752, n4753,
    n4754, n4755, n4756, n4757, n4758, n4759,
    n4760, n4761, n4762, n4763, n4764, n4765,
    n4766, n4767, n4768, n4769, n4770, n4771,
    n4772, n4773, n4774, n4775, n4776, n4777,
    n4778, n4779, n4780, n4781, n4782, n4783,
    n4784, n4785, n4786, n4787, n4788, n4789,
    n4790, n4791, n4792, n4793, n4794, n4795,
    n4796, n4797, n4798, n4799, n4800, n4801,
    n4802, n4803, n4804, n4805, n4806, n4807,
    n4808, n4809, n4810, n4811, n4812, n4813,
    n4814, n4815, n4816, n4817, n4819, n4820,
    n4821, n4822, n4823, n4824, n4825, n4826,
    n4827, n4828, n4829, n4830, n4831, n4832,
    n4833, n4834, n4835, n4836, n4837, n4838,
    n4839, n4840, n4841, n4842, n4843, n4844,
    n4845, n4846, n4847, n4848, n4849, n4850,
    n4851, n4852, n4853, n4854, n4855, n4856,
    n4857, n4858, n4859, n4860, n4861, n4862,
    n4863, n4864, n4865, n4866, n4867, n4868,
    n4869, n4870, n4871, n4872, n4873, n4874,
    n4875, n4876, n4877, n4878, n4879, n4880,
    n4881, n4882, n4883, n4884, n4885, n4886,
    n4887, n4888, n4889, n4890, n4891, n4892,
    n4893, n4894, n4895, n4896, n4897, n4898,
    n4899, n4900, n4901, n4902, n4903, n4904,
    n4905, n4906, n4907, n4908, n4909, n4910,
    n4911, n4912, n4913, n4914, n4915, n4916,
    n4917, n4918, n4919, n4920, n4921, n4922,
    n4923, n4924, n4925, n4926, n4927, n4928,
    n4929, n4930, n4931, n4932, n4933, n4934,
    n4935, n4936, n4937, n4938, n4939, n4940,
    n4941, n4942, n4943, n4944, n4945, n4946,
    n4947, n4948, n4949, n4950, n4951, n4952,
    n4953, n4954, n4955, n4956, n4957, n4958,
    n4959, n4960, n4961, n4962, n4963, n4964,
    n4965, n4966, n4967, n4968, n4969, n4970,
    n4971, n4972, n4973, n4974, n4975, n4976,
    n4977, n4978, n4979, n4980, n4981, n4982,
    n4983, n4984, n4985, n4986, n4987, n4988,
    n4989, n4990, n4991, n4992, n4993, n4994,
    n4995, n4996, n4997, n4998, n4999, n5000,
    n5001, n5002, n5003, n5004, n5005, n5006,
    n5007, n5008, n5009, n5010, n5011, n5012,
    n5013, n5014, n5015, n5016, n5017, n5018,
    n5019, n5020, n5021, n5022, n5023, n5024,
    n5025, n5026, n5027, n5028, n5029, n5030,
    n5031, n5032, n5033, n5034, n5035, n5036,
    n5037, n5038, n5039, n5041, n5042, n5043,
    n5044, n5045, n5046, n5047, n5048, n5049,
    n5050, n5051, n5052, n5053, n5054, n5055,
    n5056, n5057, n5058, n5059, n5060, n5061,
    n5062, n5063, n5064, n5065, n5066, n5067,
    n5068, n5069, n5070, n5071, n5072, n5073,
    n5074, n5075, n5076, n5077, n5078, n5079,
    n5080, n5081, n5082, n5083, n5084, n5085,
    n5086, n5087, n5088, n5089, n5090, n5091,
    n5092, n5093, n5094, n5095, n5096, n5097,
    n5098, n5099, n5100, n5101, n5102, n5103,
    n5104, n5105, n5106, n5107, n5108, n5109,
    n5110, n5111, n5112, n5113, n5114, n5115,
    n5116, n5117, n5118, n5119, n5120, n5121,
    n5122, n5123, n5124, n5125, n5126, n5127,
    n5128, n5129, n5130, n5131, n5132, n5133,
    n5134, n5135, n5136, n5137, n5138, n5139,
    n5140, n5141, n5142, n5143, n5144, n5145,
    n5146, n5147, n5148, n5149, n5150, n5151,
    n5152, n5153, n5154, n5155, n5156, n5157,
    n5158, n5159, n5160, n5161, n5162, n5163,
    n5164, n5165, n5166, n5167, n5168, n5169,
    n5170, n5171, n5172, n5173, n5174, n5175,
    n5176, n5177, n5178, n5179, n5180, n5181,
    n5182, n5183, n5184, n5185, n5186, n5187,
    n5188, n5189, n5190, n5191, n5192, n5193,
    n5194, n5195, n5196, n5197, n5198, n5199,
    n5200, n5201, n5202, n5203, n5204, n5205,
    n5206, n5207, n5208, n5209, n5210, n5211,
    n5212, n5213, n5214, n5215, n5216, n5217,
    n5218, n5219, n5220, n5221, n5222, n5223,
    n5224, n5225, n5226, n5227, n5228, n5229,
    n5230, n5231, n5232, n5233, n5234, n5235,
    n5236, n5237, n5238, n5239, n5240, n5241,
    n5242, n5243, n5244, n5245, n5246, n5247,
    n5248, n5249, n5250, n5251, n5252, n5253,
    n5254, n5255, n5256, n5257, n5258, n5259,
    n5260, n5262, n5263, n5264, n5265, n5266,
    n5267, n5268, n5269, n5270, n5271, n5272,
    n5273, n5274, n5275, n5276, n5277, n5278,
    n5279, n5280, n5281, n5282, n5283, n5284,
    n5285, n5286, n5287, n5288, n5289, n5290,
    n5291, n5292, n5293, n5294, n5295, n5296,
    n5297, n5298, n5299, n5300, n5301, n5302,
    n5303, n5304, n5305, n5306, n5307, n5308,
    n5309, n5310, n5311, n5312, n5313, n5314,
    n5315, n5316, n5317, n5318, n5319, n5320,
    n5321, n5322, n5323, n5324, n5325, n5326,
    n5327, n5328, n5329, n5330, n5331, n5332,
    n5333, n5334, n5335, n5336, n5337, n5338,
    n5339, n5340, n5341, n5342, n5343, n5344,
    n5345, n5346, n5347, n5348, n5349, n5350,
    n5351, n5352, n5353, n5354, n5355, n5356,
    n5357, n5358, n5359, n5360, n5361, n5362,
    n5363, n5364, n5365, n5366, n5367, n5368,
    n5369, n5370, n5371, n5372, n5373, n5374,
    n5375, n5376, n5377, n5378, n5379, n5380,
    n5381, n5382, n5383, n5384, n5385, n5386,
    n5387, n5388, n5389, n5390, n5391, n5392,
    n5393, n5394, n5395, n5396, n5397, n5398,
    n5399, n5400, n5401, n5402, n5403, n5404,
    n5405, n5406, n5407, n5408, n5409, n5410,
    n5411, n5412, n5413, n5414, n5415, n5416,
    n5417, n5418, n5419, n5420, n5421, n5422,
    n5423, n5424, n5425, n5426, n5427, n5428,
    n5429, n5430, n5431, n5432, n5433, n5434,
    n5435, n5436, n5437, n5438, n5439, n5440,
    n5441, n5442, n5443, n5444, n5445, n5446,
    n5447, n5448, n5449, n5450, n5451, n5452,
    n5453, n5454, n5455, n5456, n5457, n5458,
    n5459, n5460, n5461, n5462, n5463, n5464,
    n5465, n5466, n5467, n5468, n5469, n5470,
    n5471, n5472, n5473, n5474, n5475, n5476,
    n5477, n5478, n5479, n5480, n5481, n5482,
    n5483, n5484, n5485, n5486, n5487, n5488,
    n5489, n5490, n5491, n5492, n5493, n5494,
    n5496, n5497, n5498, n5499, n5500, n5501,
    n5502, n5503, n5504, n5505, n5506, n5507,
    n5508, n5509, n5510, n5511, n5512, n5513,
    n5514, n5515, n5516, n5517, n5518, n5519,
    n5520, n5521, n5522, n5523, n5524, n5525,
    n5526, n5527, n5528, n5529, n5530, n5531,
    n5532, n5533, n5534, n5535, n5536, n5537,
    n5538, n5539, n5540, n5541, n5542, n5543,
    n5544, n5545, n5546, n5547, n5548, n5549,
    n5550, n5551, n5552, n5553, n5554, n5555,
    n5556, n5557, n5558, n5559, n5560, n5561,
    n5562, n5563, n5564, n5565, n5566, n5567,
    n5568, n5569, n5570, n5571, n5572, n5573,
    n5574, n5575, n5576, n5577, n5578, n5579,
    n5580, n5581, n5582, n5583, n5584, n5585,
    n5586, n5587, n5588, n5589, n5590, n5591,
    n5592, n5593, n5594, n5595, n5596, n5597,
    n5598, n5599, n5600, n5601, n5602, n5603,
    n5604, n5605, n5606, n5607, n5608, n5609,
    n5610, n5611, n5612, n5613, n5614, n5615,
    n5616, n5617, n5618, n5619, n5620, n5621,
    n5622, n5623, n5624, n5625, n5626, n5627,
    n5628, n5629, n5630, n5631, n5632, n5633,
    n5634, n5635, n5636, n5637, n5638, n5639,
    n5640, n5641, n5642, n5643, n5644, n5645,
    n5646, n5647, n5648, n5649, n5650, n5651,
    n5652, n5653, n5654, n5655, n5656, n5657,
    n5658, n5659, n5660, n5661, n5662, n5663,
    n5664, n5665, n5666, n5667, n5668, n5669,
    n5670, n5671, n5672, n5673, n5674, n5675,
    n5676, n5677, n5678, n5679, n5680, n5681,
    n5682, n5683, n5684, n5685, n5686, n5687,
    n5688, n5689, n5690, n5691, n5692, n5693,
    n5694, n5695, n5696, n5697, n5698, n5699,
    n5700, n5701, n5702, n5703, n5704, n5705,
    n5706, n5707, n5708, n5709, n5710, n5711,
    n5712, n5713, n5714, n5715, n5716, n5717,
    n5718, n5719, n5720, n5721, n5722, n5723,
    n5724, n5725, n5726, n5727, n5728, n5730,
    n5731, n5732, n5733, n5734, n5735, n5736,
    n5737, n5738, n5739, n5740, n5741, n5742,
    n5743, n5744, n5745, n5746, n5747, n5748,
    n5749, n5750, n5751, n5752, n5753, n5754,
    n5755, n5756, n5757, n5758, n5759, n5760,
    n5761, n5762, n5763, n5764, n5765, n5766,
    n5767, n5768, n5769, n5770, n5771, n5772,
    n5773, n5774, n5775, n5776, n5777, n5778,
    n5779, n5780, n5781, n5782, n5783, n5784,
    n5785, n5786, n5787, n5788, n5789, n5790,
    n5791, n5792, n5793, n5794, n5795, n5796,
    n5797, n5798, n5799, n5800, n5801, n5802,
    n5803, n5804, n5805, n5806, n5807, n5808,
    n5809, n5810, n5811, n5812, n5813, n5814,
    n5815, n5816, n5817, n5818, n5819, n5820,
    n5821, n5822, n5823, n5824, n5825, n5826,
    n5827, n5828, n5829, n5830, n5831, n5832,
    n5833, n5834, n5835, n5836, n5837, n5838,
    n5839, n5840, n5841, n5842, n5843, n5844,
    n5845, n5846, n5847, n5848, n5849, n5850,
    n5851, n5852, n5853, n5854, n5855, n5856,
    n5857, n5858, n5859, n5860, n5861, n5862,
    n5863, n5864, n5865, n5866, n5867, n5868,
    n5869, n5870, n5871, n5872, n5873, n5874,
    n5875, n5876, n5877, n5878, n5879, n5880,
    n5881, n5882, n5883, n5884, n5885, n5886,
    n5887, n5888, n5889, n5890, n5891, n5892,
    n5893, n5894, n5895, n5896, n5897, n5898,
    n5899, n5900, n5901, n5902, n5903, n5904,
    n5905, n5906, n5907, n5908, n5909, n5910,
    n5911, n5912, n5913, n5914, n5915, n5916,
    n5917, n5918, n5919, n5920, n5921, n5922,
    n5923, n5924, n5925, n5926, n5927, n5928,
    n5929, n5930, n5931, n5932, n5933, n5934,
    n5935, n5936, n5937, n5938, n5939, n5940,
    n5941, n5942, n5943, n5944, n5945, n5946,
    n5947, n5948, n5949, n5950, n5951, n5952,
    n5953, n5954, n5955, n5956, n5957, n5958,
    n5959, n5960, n5961, n5962, n5963, n5964,
    n5965, n5966, n5967, n5968, n5969, n5970,
    n5971, n5972, n5973, n5974, n5975, n5976,
    n5977, n5978, n5979, n5980, n5981, n5982,
    n5983, n5984, n5985, n5986, n5987, n5988,
    n5989, n5990, n5991, n5992, n5993, n5994,
    n5995, n5996, n5997, n5998, n5999, n6000,
    n6001, n6002, n6003, n6004, n6005, n6006,
    n6007, n6008, n6009, n6010, n6011, n6012,
    n6013, n6014, n6015, n6016, n6017, n6018,
    n6019, n6020, n6021, n6022, n6023, n6024,
    n6025, n6026, n6027, n6028, n6029, n6030,
    n6031, n6032, n6033, n6034, n6035, n6036,
    n6037, n6038, n6039, n6040, n6041, n6042,
    n6043, n6044, n6045, n6046, n6047, n6048,
    n6049, n6050, n6051, n6052, n6053, n6054,
    n6055, n6056, n6057, n6058, n6059, n6060,
    n6061, n6062, n6063, n6064, n6065, n6066,
    n6067, n6068, n6069, n6070, n6071, n6072,
    n6073, n6074, n6075, n6076, n6077, n6078,
    n6079, n6080, n6081, n6082, n6084, n6085,
    n6086, n6087, n6088, n6089, n6090, n6091,
    n6092, n6093, n6094, n6095, n6096, n6097,
    n6098, n6099, n6100, n6101, n6102, n6103,
    n6104, n6105, n6106, n6107, n6108, n6109,
    n6110, n6111, n6112, n6113, n6114, n6115,
    n6116, n6118, n6119, n6120, n6121, n6122,
    n6124, n6125, n6126, n6127, n6128, n6129,
    n6130, n6131, n6132, n6133, n6134, n6135,
    n6136, n6137, n6138, n6139, n6140, n6141,
    n6142, n6143, n6144, n6145, n6146, n6147,
    n6148, n6149, n6150, n6151, n6152, n6153,
    n6154, n6155, n6156, n6157, n6158, n6159,
    n6160, n6161, n6162, n6163, n6164, n6165,
    n6166, n6167, n6168, n6169, n6170, n6171,
    n6172, n6173, n6174, n6175, n6176, n6177,
    n6178, n6179, n6180, n6181, n6182, n6183,
    n6184, n6185, n6186, n6187, n6188, n6190,
    n6191, n6192, n6193, n6194, n6195, n6196,
    n6197, n6198, n6199, n6200, n6201, n6202,
    n6203, n6204, n6205, n6206, n6207, n6208,
    n6209, n6210, n6211, n6212, n6213, n6214,
    n6215, n6216, n6217, n6218, n6219, n6220,
    n6221, n6222, n6223, n6224, n6225, n6226,
    n6227, n6228, n6229, n6230, n6231, n6232,
    n6233, n6234, n6235, n6236, n6237, n6238,
    n6239, n6240, n6241, n6242, n6243, n6244,
    n6245, n6246, n6247, n6248, n6249, n6250,
    n6251, n6252, n6253, n6254, n6255, n6256,
    n6257, n6258, n6259, n6260, n6261, n6262,
    n6263, n6264, n6265, n6266, n6267, n6268,
    n6269, n6270, n6271, n6273, n6274, n6275,
    n6276, n6277, n6278, n6279, n6280, n6281,
    n6282, n6283, n6284, n6285, n6286, n6287,
    n6288, n6289, n6290, n6291, n6292, n6293,
    n6294, n6295, n6296, n6297, n6298, n6299,
    n6300, n6301, n6302, n6303, n6304, n6305,
    n6306, n6307, n6308, n6309, n6310, n6311,
    n6312, n6313, n6314, n6315, n6316, n6317,
    n6318, n6319, n6320, n6321, n6322, n6324,
    n6325, n6326, n6327, n6328, n6329, n6330,
    n6331, n6332, n6333, n6334, n6335, n6336,
    n6337, n6338, n6339, n6340, n6341, n6342,
    n6343, n6344, n6345, n6346, n6347, n6348,
    n6349, n6350, n6351, n6352, n6353, n6354,
    n6355, n6356, n6357, n6358, n6359, n6360,
    n6361, n6362, n6363, n6364, n6365, n6366,
    n6367, n6368, n6369, n6370, n6371, n6372,
    n6373, n6374, n6375, n6376, n6377, n6378,
    n6379, n6380, n6381, n6382, n6383, n6384,
    n6385, n6386, n6387, n6388, n6389, n6390,
    n6391, n6392, n6393, n6394, n6395, n6396,
    n6397, n6398, n6399, n6400, n6401, n6402,
    n6403, n6404, n6405, n6406, n6407, n6408,
    n6409, n6410, n6411, n6412, n6413, n6414,
    n6415, n6416, n6417, n6418, n6419, n6420,
    n6421, n6422, n6423, n6424, n6425, n6426,
    n6427, n6428, n6429, n6430, n6431, n6432,
    n6433, n6434, n6435, n6436, n6437, n6438,
    n6439, n6440, n6441, n6442, n6443, n6444,
    n6445, n6446, n6447, n6448, n6449, n6450,
    n6451, n6452, n6453, n6454, n6455, n6456,
    n6457, n6458, n6459, n6460, n6461, n6462,
    n6463, n6464, n6465, n6466, n6467, n6468,
    n6469, n6470, n6471, n6472, n6473, n6474,
    n6475, n6476, n6477, n6478, n6479, n6480,
    n6481, n6482, n6483, n6484, n6485, n6486,
    n6487, n6488, n6489, n6490, n6491, n6492,
    n6493, n6494, n6495, n6496, n6497, n6498,
    n6499, n6500, n6501, n6502, n6503, n6504,
    n6505, n6506, n6507, n6508, n6509, n6510,
    n6511, n6512, n6513, n6514, n6515, n6516,
    n6517, n6518, n6519, n6520, n6521, n6522,
    n6523, n6524, n6525, n6526, n6527, n6528,
    n6529, n6530, n6531, n6532, n6533, n6534,
    n6535, n6536, n6537, n6538, n6539, n6541,
    n6542, n6543, n6544, n6545, n6546, n6547,
    n6548, n6549, n6550, n6551, n6552, n6553,
    n6554, n6555, n6556, n6557, n6558, n6559,
    n6560, n6561, n6562, n6563, n6564, n6565,
    n6566, n6567, n6568, n6569, n6570, n6571,
    n6572, n6573, n6574, n6575, n6576, n6577,
    n6578, n6579, n6580, n6581, n6582, n6583,
    n6584, n6585, n6586, n6587, n6588, n6589,
    n6590, n6591, n6592, n6593, n6594, n6595,
    n6596, n6597, n6598, n6599, n6600, n6601,
    n6602, n6603, n6604, n6605, n6606, n6607,
    n6608, n6609, n6610, n6611, n6612, n6613,
    n6614, n6615, n6616, n6617, n6618, n6619,
    n6620, n6621, n6622, n6623, n6624, n6625,
    n6626, n6627, n6628, n6629, n6630, n6631,
    n6632, n6633, n6634, n6635, n6636, n6637,
    n6638, n6639, n6640, n6641, n6642, n6643,
    n6644, n6645, n6646, n6647, n6648, n6649,
    n6650, n6651, n6652, n6653, n6654, n6655,
    n6656, n6657, n6658, n6659, n6660, n6661,
    n6662, n6664, n6665, n6666, n6667, n6668,
    n6669, n6670, n6671, n6672, n6673, n6674,
    n6675, n6676, n6677, n6678, n6679, n6680,
    n6681, n6682, n6683, n6684, n6685, n6686,
    n6687, n6688, n6689, n6690, n6691, n6692,
    n6693, n6694, n6695, n6696, n6697, n6698,
    n6699, n6700, n6701, n6702, n6703, n6704,
    n6705, n6706, n6707, n6708, n6709, n6710,
    n6711, n6712, n6713, n6714, n6715, n6716,
    n6717, n6718, n6719, n6720, n6721, n6722,
    n6723, n6724, n6725, n6726, n6727, n6728,
    n6729, n6730, n6731, n6732, n6733, n6734,
    n6735, n6736, n6737, n6738, n6739, n6740,
    n6741, n6742, n6743, n6744, n6745, n6746,
    n6747, n6748, n6749, n6750, n6751, n6752,
    n6753, n6754, n6755, n6756, n6757, n6758,
    n6759, n6760, n6761, n6762, n6763, n6764,
    n6765, n6766, n6767, n6768, n6769, n6770,
    n6771, n6772, n6773, n6774, n6775, n6776,
    n6777, n6778, n6779, n6780, n6781, n6782,
    n6783, n6784, n6785, n6786, n6787, n6788,
    n6790, n6791, n6792, n6793, n6794, n6795,
    n6796, n6797, n6798, n6799, n6800, n6801,
    n6802, n6803, n6804, n6805, n6806, n6807,
    n6808, n6809, n6810, n6811, n6812, n6813,
    n6814, n6815, n6816, n6817, n6818, n6819,
    n6820, n6821, n6822, n6823, n6824, n6825,
    n6826, n6827, n6828, n6829, n6830, n6831,
    n6832, n6833, n6834, n6835, n6836, n6837,
    n6838, n6839, n6840, n6841, n6842, n6843,
    n6844, n6845, n6846, n6847, n6848, n6849,
    n6850, n6851, n6852, n6853, n6854, n6855,
    n6856, n6857, n6858, n6859, n6860, n6861,
    n6862, n6863, n6864, n6865, n6866, n6867,
    n6868, n6869, n6870, n6871, n6872, n6873,
    n6874, n6875, n6876, n6877, n6878, n6879,
    n6880, n6882, n6883, n6884, n6885, n6886,
    n6887, n6888, n6889, n6890, n6891, n6892,
    n6893, n6894, n6895, n6896, n6897, n6898,
    n6899, n6900, n6901, n6902, n6903, n6904,
    n6905, n6906, n6907, n6908, n6909, n6910,
    n6911, n6912, n6913, n6914, n6915, n6916,
    n6917, n6918, n6919, n6920, n6921, n6922,
    n6923, n6924, n6925, n6926, n6927, n6928,
    n6929, n6930, n6931, n6932, n6933, n6934,
    n6935, n6936, n6937, n6938, n6939, n6940,
    n6941, n6942, n6943, n6944, n6945, n6946,
    n6947, n6948, n6949, n6950, n6951, n6952,
    n6953, n6954, n6955, n6956, n6957, n6958,
    n6959, n6960, n6961, n6962, n6963, n6964,
    n6965, n6966, n6967, n6968, n6969, n6970,
    n6971, n6972, n6974, n6975, n6976, n6977,
    n6978, n6979, n6980, n6981, n6982, n6983,
    n6984, n6985, n6986, n6987, n6988, n6989,
    n6990, n6991, n6992, n6993, n6994, n6995,
    n6996, n6997, n6998, n6999, n7000, n7001,
    n7002, n7003, n7004, n7005, n7006, n7007,
    n7008, n7009, n7010, n7011, n7012, n7013,
    n7014, n7015, n7016, n7017, n7018, n7019,
    n7020, n7021, n7022, n7023, n7024, n7025,
    n7026, n7027, n7028, n7029, n7030, n7031,
    n7032, n7033, n7034, n7035, n7036, n7037,
    n7038, n7039, n7040, n7041, n7042, n7043,
    n7044, n7045, n7046, n7047, n7048, n7049,
    n7050, n7051, n7052, n7053, n7054, n7055,
    n7056, n7057, n7058, n7059, n7060, n7061,
    n7062, n7063, n7064, n7066, n7067, n7068,
    n7069, n7070, n7071, n7072, n7073, n7074,
    n7075, n7076, n7077, n7078, n7079, n7080,
    n7081, n7082, n7083, n7084, n7085, n7086,
    n7087, n7088, n7089, n7090, n7091, n7092,
    n7093, n7094, n7095, n7096, n7097, n7098,
    n7099, n7100, n7101, n7102, n7103, n7104,
    n7105, n7106, n7107, n7108, n7109, n7110,
    n7111, n7112, n7113, n7114, n7115, n7116,
    n7117, n7118, n7119, n7120, n7121, n7122,
    n7123, n7124, n7125, n7126, n7127, n7128,
    n7129, n7130, n7131, n7132, n7133, n7134,
    n7135, n7136, n7137, n7138, n7139, n7140,
    n7141, n7142, n7143, n7144, n7145, n7146,
    n7147, n7148, n7149, n7150, n7151, n7152,
    n7153, n7154, n7155, n7156, n7158, n7159,
    n7160, n7161, n7162, n7163, n7164, n7165,
    n7166, n7167, n7168, n7169, n7170, n7171,
    n7172, n7173, n7174, n7175, n7176, n7177,
    n7178, n7179, n7180, n7181, n7182, n7183,
    n7184, n7185, n7186, n7187, n7188, n7189,
    n7190, n7191, n7192, n7193, n7194, n7195,
    n7196, n7197, n7198, n7199, n7200, n7201,
    n7202, n7203, n7204, n7205, n7206, n7207,
    n7208, n7209, n7210, n7211, n7212, n7213,
    n7214, n7215, n7216, n7217, n7218, n7219,
    n7220, n7221, n7222, n7223, n7224, n7225,
    n7226, n7227, n7228, n7229, n7230, n7231,
    n7232, n7233, n7234, n7235, n7236, n7237,
    n7238, n7239, n7240, n7241, n7242, n7243,
    n7244, n7245, n7246, n7247, n7249, n7250,
    n7251, n7252, n7253, n7254, n7255, n7256,
    n7257, n7258, n7259, n7260, n7261, n7262,
    n7263, n7264, n7265, n7266, n7267, n7268,
    n7269, n7270, n7271, n7272, n7273, n7274,
    n7275, n7276, n7277, n7278, n7279, n7280,
    n7281, n7282, n7283, n7284, n7285, n7286,
    n7287, n7288, n7289, n7290, n7291, n7292,
    n7293, n7294, n7295, n7296, n7297, n7298,
    n7299, n7300, n7301, n7303, n7304, n7306,
    n7307, n7308, n7309, n7310, n7311, n7312,
    n7313, n7314, n7315, n7316, n7317, n7318,
    n7319, n7320, n7321, n7322, n7323, n7324,
    n7325, n7326, n7327, n7328, n7329, n7330,
    n7331, n7332, n7333, n7334, n7335, n7336,
    n7337, n7338, n7339, n7340, n7341, n7342,
    n7343, n7344, n7345, n7346, n7347, n7348,
    n7349, n7350, n7351, n7352, n7353, n7354,
    n7355, n7357, n7358, n7359, n7360, n7362,
    n7364, n7366, n7368, n7369, n7370, n7371,
    n7372, n7373, n7374, n7375, n7376, n7378,
    n7379, n7380, n7381, n7382, n7383, n7384,
    n7385, n7386, n7387, n7388, n7389, n7390,
    n7391, n7392, n7393, n7394, n7395, n7396,
    n7397, n7398, n7399, n7400, n7401, n7402,
    n7403, n7404, n7405, n7406, n7407, n7408,
    n7409, n7410, n7411, n7412, n7413, n7414,
    n7415, n7416, n7417, n7418, n7419, n7420,
    n7421, n7422, n7423, n7424, n7425, n7426,
    n7427, n7428, n7429, n7430, n7431, n7432,
    n7433, n7434, n7435, n7436, n7437, n7438,
    n7439, n7440, n7441, n7442, n7443, n7444,
    n7445, n7446, n7447, n7448, n7449, n7450,
    n7451, n7452, n7453, n7454, n7455, n7456,
    n7457, n7458, n7459, n7460, n7461, n7462,
    n7463, n7464, n7465, n7466, n7467, n7468,
    n7469, n7470, n7471, n7472, n7473, n7474,
    n7475, n7476, n7477, n7478, n7479, n7480,
    n7481, n7482, n7483, n7484, n7485, n7486,
    n7487, n7488, n7489, n7490, n7491, n7492,
    n7493, n7494, n7495, n7496, n7497, n7498,
    n7499, n7500, n7501, n7502, n7503, n7504,
    n7505, n7506, n7507, n7508, n7509, n7510,
    n7511, n7512, n7513, n7514, n7515, n7516,
    n7517, n7518, n7519, n7520, n7521, n7522,
    n7523, n7524, n7525, n7526, n7527, n7528,
    n7529, n7530, n7531, n7532, n7533, n7534,
    n7535, n7536, n7537, n7538, n7539, n7540,
    n7541, n7542, n7543, n7544, n7545, n7546,
    n7547, n7548, n7549, n7550, n7551, n7552,
    n7553, n7554, n7555, n7556, n7557, n7558,
    n7559, n7560, n7561, n7562, n7563, n7564,
    n7565, n7566, n7567, n7568, n7569, n7570,
    n7571, n7572, n7573, n7574, n7575, n7576,
    n7577, n7578, n7579, n7580, n7581, n7582,
    n7583, n7584, n7585, n7586, n7587, n7588,
    n7589, n7590, n7591, n7592, n7593, n7594,
    n7595, n7596, n7597, n7598, n7599, n7600,
    n7601, n7602, n7603, n7604, n7605, n7606,
    n7607, n7608, n7609, n7610, n7611, n7612,
    n7613, n7614, n7615, n7616, n7617, n7618,
    n7619, n7620, n7621, n7622, n7623, n7624,
    n7625, n7626, n7627, n7628, n7629, n7630,
    n7631, n7632, n7633, n7634, n7635, n7636,
    n7637, n7638, n7639, n7640, n7641, n7642,
    n7643, n7644, n7645, n7646, n7647, n7648,
    n7649, n7650, n7651, n7652, n7653, n7654,
    n7655, n7656, n7657, n7658, n7659, n7660,
    n7661, n7662, n7663, n7664, n7665, n7666,
    n7667, n7668, n7669, n7670, n7671, n7672,
    n7673, n7674, n7675, n7676, n7677, n7678,
    n7679, n7680, n7681, n7682, n7683, n7684,
    n7685, n7686, n7687, n7688, n7689, n7690,
    n7691, n7692, n7693, n7694, n7695, n7696,
    n7697, n7698, n7699, n7700, n7701, n7702,
    n7703, n7704, n7705, n7706, n7707, n7708,
    n7709, n7710, n7711, n7712, n7713, n7714,
    n7715, n7716, n7717, n7718, n7719, n7720,
    n7721, n7722, n7723, n7724, n7725, n7726,
    n7727, n7728, n7729, n7730, n7731, n7732,
    n7733, n7734, n7735, n7736, n7737, n7738,
    n7739, n7740, n7741, n7742, n7743, n7744,
    n7745, n7746, n7747, n7748, n7749, n7750,
    n7751, n7752, n7753, n7754, n7755, n7756,
    n7757, n7758, n7759, n7760, n7761, n7762,
    n7763, n7764, n7765, n7766, n7767, n7768,
    n7769, n7770, n7771, n7772, n7773, n7774,
    n7775, n7776, n7777, n7778, n7779, n7780,
    n7781, n7782, n7783, n7784, n7785, n7786,
    n7787, n7788, n7789, n7790, n7791, n7792,
    n7793, n7794, n7795, n7796, n7797, n7798,
    n7799, n7800, n7801, n7802, n7803, n7804,
    n7805, n7806, n7807, n7808, n7809, n7810,
    n7811, n7812, n7813, n7814, n7815, n7816,
    n7817, n7818, n7819, n7820, n7821, n7822,
    n7823, n7824, n7825, n7826, n7827, n7828,
    n7829, n7830, n7831, n7832, n7833, n7834,
    n7835, n7836, n7837, n7838, n7839, n7840,
    n7841, n7842, n7843, n7844, n7845, n7846,
    n7847, n7848, n7849, n7850, n7851, n7852,
    n7853, n7854, n7855, n7856, n7857, n7858,
    n7859, n7860, n7861, n7862, n7863, n7864,
    n7865, n7866, n7867, n7868, n7869, n7870,
    n7871, n7872, n7873, n7874, n7875, n7876,
    n7877, n7878, n7879, n7880, n7881, n7882,
    n7883, n7884, n7885, n7886, n7887, n7888,
    n7889, n7890, n7891, n7892, n7893, n7894,
    n7895, n7896, n7897, n7898, n7899, n7900,
    n7901, n7902, n7903, n7904, n7905, n7906,
    n7907, n7908, n7909, n7910, n7911, n7912,
    n7913, n7914, n7915, n7916, n7917, n7918,
    n7919, n7920, n7921, n7922, n7923, n7924,
    n7925, n7926, n7927, n7928, n7929, n7930,
    n7931, n7932, n7933, n7934, n7935, n7936,
    n7937, n7938, n7939, n7940, n7941, n7942,
    n7943, n7944, n7945, n7946, n7947, n7948,
    n7949, n7950, n7951, n7952, n7953, n7954,
    n7955, n7956, n7957, n7958, n7959, n7960,
    n7961, n7962, n7963, n7964, n7965, n7966,
    n7967, n7968, n7969, n7970, n7971, n7972,
    n7973, n7974, n7975, n7976, n7977, n7978,
    n7979, n7980, n7981, n7982, n7983, n7984,
    n7985, n7986, n7987, n7988, n7989, n7990,
    n7991, n7992, n7993, n7994, n7995, n7996,
    n7997, n7998, n7999, n8000, n8001, n8002,
    n8003, n8004, n8005, n8006, n8007, n8008,
    n8009, n8010, n8011, n8012, n8013, n8014,
    n8015, n8016, n8017, n8018, n8019, n8020,
    n8021, n8022, n8023, n8024, n8025, n8026,
    n8027, n8028, n8029, n8030, n8031, n8032,
    n8033, n8034, n8035, n8036, n8037, n8038,
    n8039, n8040, n8041, n8042, n8043, n8044,
    n8045, n8046, n8047, n8048, n8049, n8050,
    n8051, n8052, n8053, n8054, n8055, n8056,
    n8057, n8058, n8059, n8060, n8061, n8062,
    n8063, n8064, n8065, n8066, n8067, n8068,
    n8069, n8070, n8071, n8072, n8073, n8074,
    n8075, n8076, n8077, n8078, n8079, n8080,
    n8081, n8082, n8083, n8084, n8085, n8086,
    n8087, n8088, n8089, n8090, n8091, n8092,
    n8093, n8094, n8095, n8096, n8097, n8098,
    n8099, n8100, n8101, n8102, n8103, n8104,
    n8105, n8106, n8107, n8108, n8109, n8110,
    n8111, n8112, n8113, n8114, n8115, n8116,
    n8117, n8118, n8119, n8120, n8121, n8122,
    n8123, n8124, n8125, n8126, n8127, n8128,
    n8129, n8130, n8131, n8132, n8133, n8134,
    n8135, n8136, n8137, n8138, n8139, n8140,
    n8141, n8142, n8143, n8144, n8145, n8146,
    n8147, n8148, n8149, n8150, n8151, n8152,
    n8153, n8154, n8155, n8156, n8157, n8158,
    n8159, n8160, n8161, n8162, n8163, n8164,
    n8165, n8166, n8167, n8168, n8169, n8170,
    n8171, n8172, n8173, n8174, n8175, n8176,
    n8177, n8178, n8179, n8180, n8181, n8182,
    n8183, n8184, n8185, n8186, n8187, n8188,
    n8189, n8190, n8191, n8192, n8193, n8194,
    n8195, n8196, n8197, n8198, n8199, n8200,
    n8201, n8202, n8203, n8204, n8205, n8206,
    n8207, n8208, n8209, n8210, n8211, n8212,
    n8213, n8214, n8215, n8216, n8217, n8218,
    n8219, n8220, n8221, n8222, n8223, n8224,
    n8225, n8226, n8227, n8228, n8229, n8230,
    n8231, n8232, n8233, n8234, n8235, n8236,
    n8237, n8238, n8239, n8240, n8241, n8242,
    n8243, n8244, n8245, n8246, n8247, n8248,
    n8249, n8250, n8251, n8252, n8253, n8254,
    n8255, n8256, n8257, n8258, n8259, n8260,
    n8261, n8262, n8263, n8264, n8265, n8266,
    n8267, n8268, n8269, n8270, n8271, n8272,
    n8273, n8274, n8275, n8276, n8277, n8278,
    n8279, n8280, n8281, n8282, n8283, n8284,
    n8285, n8286, n8287, n8288, n8289, n8290,
    n8291, n8292, n8293, n8294, n8295, n8296,
    n8297, n8298, n8299, n8300, n8301, n8302,
    n8303, n8304, n8305, n8306, n8307, n8308,
    n8309, n8310, n8311, n8312, n8313, n8314,
    n8315, n8316, n8317, n8318, n8319, n8320,
    n8321, n8322, n8323, n8324, n8325, n8326,
    n8327, n8328, n8329, n8330, n8331, n8332,
    n8333, n8334, n8335, n8336, n8337, n8338,
    n8339, n8340, n8341, n8342, n8343, n8344,
    n8345, n8346, n8347, n8348, n8349, n8350,
    n8351, n8352, n8353, n8354, n8355, n8356,
    n8357, n8358, n8359, n8360, n8361, n8362,
    n8363, n8364, n8365, n8366, n8367, n8368,
    n8369, n8370, n8371, n8372, n8373, n8374,
    n8375, n8376, n8377, n8378, n8379, n8380,
    n8381, n8382, n8383, n8384, n8385, n8386,
    n8387, n8388, n8389, n8390, n8391, n8392,
    n8393, n8394, n8395, n8396, n8397, n8398,
    n8399, n8400, n8401, n8402, n8403, n8404,
    n8405, n8406, n8407, n8408, n8409, n8410,
    n8411, n8412, n8413, n8414, n8415, n8416,
    n8417, n8418, n8419, n8420, n8421, n8422,
    n8423, n8424, n8425, n8426, n8427, n8428,
    n8429, n8430, n8431, n8432, n8433, n8434,
    n8435, n8436, n8437, n8438, n8439, n8440,
    n8441, n8442, n8443, n8444, n8445, n8446,
    n8447, n8448, n8449, n8450, n8451, n8452,
    n8453, n8454, n8455, n8456, n8457, n8458,
    n8459, n8460, n8461, n8462, n8463, n8464,
    n8465, n8466, n8467, n8468, n8469, n8470,
    n8471, n8472, n8473, n8474, n8475, n8476,
    n8477, n8478, n8479, n8480, n8481, n8482,
    n8483, n8484, n8485, n8486, n8487, n8488,
    n8489, n8490, n8491, n8492, n8493, n8494,
    n8495, n8496, n8497, n8498, n8499, n8500,
    n8501, n8502, n8503, n8504, n8505, n8506,
    n8507, n8508, n8509, n8510, n8511, n8512,
    n8513, n8514, n8515, n8516, n8517, n8518,
    n8519, n8520, n8521, n8522, n8523, n8524,
    n8525, n8526, n8527, n8528, n8529, n8530,
    n8531, n8532, n8533, n8534, n8535, n8536,
    n8537, n8538, n8539, n8540, n8541, n8542,
    n8543, n8544, n8545, n8546, n8547, n8548,
    n8549, n8550, n8551, n8552, n8553, n8554,
    n8555, n8556, n8557, n8558, n8559, n8560,
    n8561, n8562, n8563, n8564, n8565, n8566,
    n8567, n8568, n8569, n8570, n8571, n8572,
    n8573, n8574, n8575, n8576, n8577, n8578,
    n8579, n8580, n8581, n8582, n8583, n8584,
    n8585, n8586, n8587, n8588, n8589, n8590,
    n8591, n8592, n8593, n8594, n8595, n8596,
    n8597, n8598, n8599, n8600, n8601, n8602,
    n8603, n8604, n8605, n8606, n8607, n8608,
    n8609, n8610, n8611, n8612, n8613, n8614,
    n8615, n8616, n8617, n8618, n8619, n8620,
    n8621, n8622, n8623, n8624, n8625, n8626,
    n8627, n8628, n8629, n8630, n8631, n8632,
    n8633, n8634, n8635, n8636, n8637, n8638,
    n8639, n8640, n8641, n8642, n8643, n8644,
    n8645, n8646, n8647, n8648, n8649, n8650,
    n8651, n8652, n8653, n8654, n8655, n8656,
    n8657, n8658, n8659, n8660, n8661, n8662,
    n8663, n8664, n8665, n8666, n8667, n8668,
    n8669, n8670, n8671, n8672, n8673, n8674,
    n8675, n8676, n8677, n8678, n8679, n8680,
    n8681, n8682, n8683, n8684, n8685, n8686,
    n8687, n8688, n8689, n8690, n8691, n8692,
    n8693, n8694, n8695, n8696, n8697, n8698,
    n8699, n8700, n8701, n8702, n8703, n8704,
    n8705, n8706, n8707, n8708, n8709, n8710,
    n8711, n8712, n8713, n8714, n8715, n8716,
    n8717, n8718, n8719, n8720, n8721, n8722,
    n8723, n8724, n8725, n8726, n8727, n8728,
    n8729, n8730, n8731, n8732, n8733, n8734,
    n8735, n8736, n8738, n8739, n8740, n8741,
    n8742, n8743, n8744, n8745, n8746, n8747,
    n8748, n8749, n8750, n8751, n8752, n8754,
    n8755, n8756, n8757, n8758, n8759, n8760,
    n8761, n8762, n8763, n8764, n8765, n8766,
    n8767, n8768, n8769, n8770, n8771, n8772,
    n8773, n8774, n8775, n8776, n8777, n8778,
    n8779, n8780, n8781, n8782, n8783, n8784,
    n8785, n8786, n8787, n8788, n8789, n8790,
    n8791, n8792, n8793, n8794, n8795, n8796,
    n8797, n8798, n8799, n8800, n8801, n8802,
    n8803, n8804, n8805, n8806, n8807, n8808,
    n8809, n8810, n8811, n8812, n8813, n8814,
    n8815, n8816, n8817, n8818, n8819, n8820,
    n8821, n8822, n8823, n8824, n8825, n8826,
    n8827, n8829, n8830, n8831, n8832, n8833,
    n8834, n8835, n8836, n8837, n8838, n8839,
    n8840, n8841, n8842, n8843, n8844, n8845,
    n8846, n8847, n8848, n8849, n8850, n8851,
    n8852, n8853, n8854, n8855, n8856, n8857,
    n8858, n8859, n8860, n8861, n8862, n8863,
    n8864, n8865, n8866, n8867, n8868, n8869,
    n8870, n8871, n8872, n8873, n8874, n8875,
    n8876, n8877, n8878, n8879, n8880, n8881,
    n8882, n8883, n8884, n8885, n8886, n8887,
    n8888, n8889, n8890, n8891, n8892, n8893,
    n8894, n8895, n8896, n8897, n8898, n8899,
    n8900, n8901, n8902, n8903, n8904, n8905,
    n8906, n8907, n8908, n8909, n8910, n8911,
    n8912, n8913, n8914, n8915, n8916, n8917,
    n8918, n8919, n8920, n8921, n8922, n8923,
    n8924, n8925, n8926, n8927, n8928, n8929,
    n8930, n8931, n8932, n8933, n8934, n8935,
    n8936, n8937, n8938, n8939, n8940, n8941,
    n8942, n8943, n8944, n8945, n8946, n8947,
    n8948, n8949, n8950, n8951, n8952, n8953,
    n8954, n8955, n8956, n8957, n8958, n8959,
    n8960, n8961, n8962, n8963, n8964, n8965,
    n8966, n8967, n8968, n8969, n8970, n8971,
    n8972, n8973, n8974, n8975, n8976, n8977,
    n8978, n8979, n8980, n8981, n8982, n8983,
    n8984, n8985, n8986, n8987, n8988, n8989,
    n8990, n8991, n8992, n8993, n8994, n8995,
    n8996, n8997, n8998, n8999, n9000, n9001,
    n9002, n9003, n9004, n9005, n9006, n9007,
    n9008, n9009, n9010, n9011, n9012, n9013,
    n9014, n9015, n9016, n9017, n9018, n9019,
    n9020, n9021, n9022, n9023, n9024, n9025,
    n9026, n9027, n9028, n9029, n9030, n9031,
    n9032, n9033, n9034, n9035, n9036, n9037,
    n9038, n9039, n9040, n9041, n9042, n9043,
    n9044, n9045, n9046, n9047, n9048, n9049,
    n9050, n9051, n9052, n9053, n9054, n9055,
    n9056, n9057, n9058, n9059, n9060, n9061,
    n9062, n9063, n9064, n9065, n9066, n9067,
    n9068, n9069, n9070, n9071, n9072, n9073,
    n9074, n9075, n9076, n9077, n9078, n9079,
    n9080, n9081, n9082, n9083, n9084, n9085,
    n9086, n9087, n9088, n9089, n9090, n9091,
    n9092, n9093, n9094, n9095, n9096, n9097,
    n9098, n9099, n9100, n9101, n9102, n9103,
    n9104, n9105, n9106, n9107, n9108, n9109,
    n9110, n9111, n9112, n9113, n9114, n9115,
    n9116, n9117, n9118, n9119, n9120, n9121,
    n9122, n9123, n9124, n9125, n9126, n9127,
    n9128, n9129, n9130, n9131, n9132, n9133,
    n9134, n9135, n9136, n9137, n9138, n9139,
    n9140, n9141, n9142, n9143, n9144, n9145,
    n9146, n9147, n9148, n9149, n9150, n9151,
    n9152, n9153, n9154, n9155, n9156, n9157,
    n9158, n9159, n9160, n9161, n9162, n9163,
    n9164, n9165, n9166, n9167, n9168, n9169,
    n9170, n9171, n9172, n9173, n9174, n9175,
    n9176, n9177, n9178, n9179, n9180, n9181,
    n9182, n9183, n9184, n9185, n9186, n9187,
    n9188, n9189, n9190, n9191, n9192, n9193,
    n9194, n9195, n9196, n9197, n9198, n9199,
    n9200, n9201, n9202, n9203, n9204, n9205,
    n9206, n9207, n9208, n9209, n9210, n9211,
    n9212, n9213, n9214, n9215, n9216, n9217,
    n9218, n9219, n9220, n9221, n9222, n9223,
    n9224, n9225, n9226, n9227, n9228, n9229,
    n9230, n9231, n9232, n9233, n9234, n9235,
    n9236, n9237, n9238, n9239, n9240, n9241,
    n9242, n9243, n9244, n9245, n9246, n9247,
    n9248, n9249, n9250, n9251, n9252, n9253,
    n9254, n9255, n9256, n9257, n9258, n9259,
    n9260, n9261, n9262, n9263, n9264, n9265,
    n9266, n9267, n9268, n9269, n9270, n9271,
    n9272, n9273, n9274, n9275, n9276, n9277,
    n9278, n9279, n9280, n9281, n9282, n9283,
    n9284, n9285, n9286, n9287, n9288, n9289,
    n9290, n9291, n9292, n9293, n9294, n9295,
    n9296, n9297, n9298, n9299, n9300, n9301,
    n9302, n9303, n9304, n9305, n9306, n9307,
    n9308, n9309, n9310, n9311, n9312, n9313,
    n9314, n9315, n9316, n9317, n9318, n9319,
    n9320, n9321, n9322, n9323, n9324, n9325,
    n9326, n9327, n9328, n9329, n9330, n9331,
    n9332, n9333, n9334, n9335, n9336, n9337,
    n9338, n9339, n9340, n9341, n9342, n9343,
    n9344, n9345, n9346, n9347, n9348, n9349,
    n9350, n9351, n9352, n9353, n9354, n9355,
    n9356, n9357, n9358, n9359, n9360, n9361,
    n9362, n9363, n9364, n9365, n9366, n9367,
    n9368, n9369, n9370, n9371, n9372, n9373,
    n9374, n9375, n9376, n9377, n9378, n9379,
    n9380, n9381, n9382, n9383, n9384, n9385,
    n9386, n9387, n9388, n9389, n9390, n9391,
    n9392, n9393, n9394, n9395, n9396, n9397,
    n9398, n9399, n9400, n9401, n9402, n9403,
    n9404, n9405, n9406, n9407, n9408, n9409,
    n9410, n9411, n9412, n9413, n9414, n9415,
    n9416, n9417, n9418, n9419, n9420, n9421,
    n9422, n9423, n9424, n9425, n9426, n9427,
    n9428, n9429, n9430, n9431, n9432, n9433,
    n9434, n9435, n9436, n9437, n9438, n9439,
    n9440, n9441, n9442, n9443, n9444, n9445,
    n9446, n9447, n9448, n9449, n9450, n9451,
    n9452, n9453, n9454, n9455, n9456, n9457,
    n9458, n9459, n9460, n9461, n9462, n9463,
    n9464, n9465, n9466, n9467, n9468, n9469,
    n9470, n9471, n9472, n9473, n9474, n9475,
    n9476, n9477, n9478, n9479, n9480, n9481,
    n9482, n9483, n9484, n9485, n9486, n9487,
    n9488, n9489, n9490, n9491, n9492, n9493,
    n9494, n9495, n9496, n9497, n9498, n9499,
    n9500, n9501, n9502, n9503, n9504, n9505,
    n9506, n9507, n9508, n9509, n9510, n9511,
    n9512, n9513, n9514, n9515, n9516, n9517,
    n9518, n9519, n9520, n9521, n9522, n9523,
    n9524, n9525, n9526, n9527, n9528, n9529,
    n9530, n9531, n9533, n9534, n9535, n9536,
    n9537, n9538, n9539, n9540, n9541, n9542,
    n9543, n9544, n9545, n9546, n9547, n9548,
    n9549, n9550, n9551, n9552, n9553, n9554,
    n9555, n9556, n9557, n9558, n9559, n9560,
    n9561, n9562, n9563, n9564, n9565, n9566,
    n9567, n9568, n9569, n9570, n9571, n9572,
    n9573, n9574, n9575, n9576, n9577, n9578,
    n9579, n9580, n9581, n9582, n9583, n9584,
    n9585, n9586, n9587, n9588, n9589, n9590,
    n9591, n9592, n9593, n9594, n9595, n9596,
    n9597, n9598, n9599, n9600, n9601, n9602,
    n9603, n9604, n9605, n9606, n9607, n9608,
    n9609, n9610, n9611, n9612, n9613, n9614,
    n9615, n9616, n9617, n9618, n9619, n9620,
    n9621, n9622, n9623, n9624, n9625, n9626,
    n9627, n9628, n9629, n9630, n9631, n9632,
    n9633, n9634, n9635, n9636, n9637, n9638,
    n9639, n9640, n9641, n9642, n9643, n9644,
    n9645, n9646, n9647, n9648, n9649, n9650,
    n9651, n9652, n9653, n9654, n9655, n9656,
    n9657, n9658, n9659, n9660, n9661, n9662,
    n9663, n9664, n9665, n9666, n9667, n9668,
    n9669, n9670, n9671, n9672, n9673, n9674,
    n9675, n9676, n9677, n9678, n9679, n9680,
    n9681, n9682, n9683, n9684, n9685, n9686,
    n9687, n9688, n9689, n9690, n9691, n9692,
    n9693, n9694, n9695, n9696, n9697, n9698,
    n9699, n9700, n9701, n9702, n9703, n9704,
    n9705, n9706, n9707, n9708, n9709, n9710,
    n9711, n9712, n9713, n9714, n9715, n9716,
    n9717, n9718, n9719, n9720, n9721, n9722,
    n9723, n9724, n9725, n9726, n9727, n9728,
    n9729, n9730, n9731, n9732, n9733, n9734,
    n9735, n9736, n9737, n9738, n9739, n9740,
    n9741, n9742, n9743, n9744, n9745, n9746,
    n9747, n9748, n9749, n9750, n9751, n9752,
    n9753, n9754, n9755, n9756, n9757, n9758,
    n9759, n9760, n9761, n9762, n9763, n9764,
    n9765, n9766, n9767, n9768, n9769, n9770,
    n9771, n9772, n9773, n9774, n9775, n9776,
    n9777, n9778, n9779, n9780, n9781, n9782,
    n9783, n9784, n9785, n9786, n9787, n9788,
    n9789, n9790, n9791, n9792, n9793, n9794,
    n9795, n9796, n9797, n9798, n9799, n9800,
    n9801, n9802, n9803, n9804, n9805, n9806,
    n9807, n9808, n9809, n9810, n9811, n9812,
    n9813, n9814, n9815, n9816, n9817, n9818,
    n9819, n9820, n9821, n9822, n9823, n9824,
    n9825, n9826, n9827, n9828, n9829, n9830,
    n9831, n9832, n9833, n9834, n9835, n9836,
    n9837, n9838, n9839, n9840, n9841, n9842,
    n9843, n9844, n9845, n9846, n9847, n9848,
    n9849, n9850, n9851, n9852, n9853, n9854,
    n9855, n9856, n9857, n9858, n9859, n9860,
    n9861, n9862, n9863, n9864, n9865, n9866,
    n9867, n9868, n9869, n9870, n9871, n9872,
    n9873, n9874, n9875, n9876, n9877, n9878,
    n9879, n9880, n9881, n9882, n9883, n9884,
    n9885, n9886, n9887, n9888, n9889, n9890,
    n9891, n9892, n9893, n9894, n9895, n9896,
    n9897, n9898, n9899, n9900, n9902, n9903,
    n9904, n9905, n9906, n9907, n9908, n9909,
    n9910, n9911, n9912, n9913, n9914, n9915,
    n9916, n9917, n9918, n9919, n9920, n9921,
    n9922, n9923, n9924, n9925, n9926, n9927,
    n9928, n9929, n9930, n9931, n9932, n9933,
    n9934, n9935, n9936, n9937, n9938, n9939,
    n9940, n9941, n9942, n9943, n9944, n9945,
    n9946, n9947, n9948, n9949, n9950, n9951,
    n9952, n9953, n9954, n9955, n9956, n9957,
    n9958, n9959, n9960, n9961, n9962, n9963,
    n9964, n9965, n9966, n9967, n9968, n9969,
    n9971, n9972, n9973, n9974, n9975, n9976,
    n9977, n9978, n9979, n9980, n9981, n9982,
    n9983, n9984, n9985, n9986, n9987, n9988,
    n9989, n9991, n9992, n9993, n9994, n9995,
    n9996, n9997, n9998, n9999, n10000, n10001,
    n10002, n10003, n10004, n10005, n10006, n10007,
    n10008, n10009, n10010, n10011, n10012, n10013,
    n10014, n10015, n10016, n10017, n10018, n10019,
    n10020, n10021, n10022, n10024, n10025, n10026,
    n10027, n10028, n10029, n10030, n10031, n10032,
    n10033, n10034, n10035, n10036, n10037, n10038,
    n10039, n10040, n10041, n10042, n10043, n10044,
    n10045, n10046, n10047, n10048, n10049, n10050,
    n10051, n10052, n10053, n10054, n10055, n10056,
    n10057, n10058, n10059, n10060, n10061, n10062,
    n10063, n10064, n10065, n10066, n10067, n10068,
    n10069, n10070, n10071, n10072, n10073, n10074,
    n10075, n10076, n10077, n10078, n10079, n10080,
    n10081, n10082, n10083, n10084, n10085, n10086,
    n10087, n10088, n10089, n10090, n10091, n10092,
    n10093, n10094, n10095, n10096, n10097, n10098,
    n10099, n10100, n10101, n10102, n10103, n10105,
    n10106, n10107, n10108, n10109, n10110, n10111,
    n10112, n10113, n10114, n10115, n10116, n10118,
    n10119, n10120, n10121, n10122, n10123, n10124,
    n10125, n10126, n10127, n10128, n10129, n10130,
    n10131, n10132, n10133, n10134, n10135, n10136,
    n10137, n10138, n10139, n10140, n10141, n10142,
    n10143, n10144, n10145, n10146, n10147, n10148,
    n10149, n10150, n10151, n10152, n10153, n10154,
    n10155, n10156, n10157, n10158, n10159, n10160,
    n10161, n10162, n10163, n10164, n10165, n10166,
    n10167, n10168, n10169, n10170, n10171, n10172,
    n10173, n10174, n10175, n10176, n10177, n10178,
    n10179, n10180, n10181, n10182, n10183, n10184,
    n10185, n10186, n10187, n10188, n10189, n10190,
    n10191, n10192, n10193, n10194, n10195, n10196,
    n10197, n10198, n10199, n10200, n10201, n10202,
    n10203, n10204, n10205, n10206, n10207, n10208,
    n10209, n10210, n10211, n10212, n10213, n10214,
    n10215, n10216, n10217, n10218, n10219, n10220,
    n10221, n10222, n10223, n10224, n10225, n10226,
    n10227, n10228, n10229, n10230, n10231, n10232,
    n10233, n10234, n10235, n10236, n10237, n10238,
    n10239, n10240, n10241, n10242, n10243, n10244,
    n10245, n10246, n10247, n10248, n10249, n10250,
    n10251, n10252, n10253, n10254, n10255, n10256,
    n10257, n10258, n10259, n10260, n10261, n10262,
    n10263, n10264, n10265, n10266, n10267, n10268,
    n10269, n10270, n10271, n10272, n10273, n10274,
    n10275, n10276, n10277, n10278, n10279, n10280,
    n10281, n10282, n10283, n10284, n10286, n10287,
    n10288, n10289, n10290, n10291, n10292, n10293,
    n10294, n10295, n10296, n10297, n10298, n10299,
    n10300, n10301, n10302, n10303, n10304, n10305,
    n10306, n10307, n10308, n10309, n10310, n10311,
    n10312, n10313, n10314, n10315, n10316, n10317,
    n10318, n10319, n10320, n10321, n10322, n10323,
    n10324, n10325, n10326, n10327, n10328, n10329,
    n10330, n10331, n10332, n10333, n10334, n10335,
    n10336, n10337, n10338, n10339, n10340, n10341,
    n10342, n10343, n10344, n10345, n10346, n10347,
    n10348, n10349, n10350, n10351, n10352, n10353,
    n10354, n10355, n10356, n10357, n10358, n10359,
    n10360, n10361, n10362, n10363, n10364, n10365,
    n10366, n10367, n10368, n10369, n10370, n10371,
    n10372, n10373, n10374, n10375, n10376, n10377,
    n10378, n10379, n10380, n10381, n10382, n10383,
    n10384, n10385, n10386, n10387, n10388, n10389,
    n10390, n10391, n10392, n10393, n10394, n10395,
    n10396, n10397, n10398, n10399, n10400, n10401,
    n10402, n10403, n10404, n10405, n10406, n10407,
    n10408, n10409, n10410, n10411, n10412, n10413,
    n10414, n10415, n10416, n10417, n10418, n10419,
    n10420, n10421, n10422, n10423, n10424, n10425,
    n10426, n10427, n10428, n10429, n10430, n10431,
    n10432, n10433, n10434, n10435, n10436, n10437,
    n10438, n10439, n10440, n10441, n10442, n10443,
    n10444, n10445, n10446, n10447, n10448, n10449,
    n10450, n10451, n10452, n10453, n10454, n10455,
    n10456, n10457, n10458, n10459, n10460, n10461,
    n10462, n10463, n10464, n10465, n10466, n10467,
    n10468, n10469, n10470, n10471, n10472, n10473,
    n10474, n10475, n10476, n10477, n10478, n10479,
    n10480, n10481, n10482, n10483, n10484, n10485,
    n10486, n10487, n10488, n10489, n10490, n10491,
    n10492, n10493, n10494, n10495, n10496, n10497,
    n10498, n10499, n10500, n10501, n10502, n10503,
    n10504, n10505, n10506, n10507, n10508, n10509,
    n10510, n10511, n10512, n10513, n10514, n10515,
    n10516, n10517, n10518, n10519, n10520, n10522,
    n10523, n10524, n10525, n10526, n10527, n10528,
    n10529, n10530, n10531, n10532, n10533, n10534,
    n10535, n10536, n10537, n10538, n10539, n10540,
    n10541, n10542, n10543, n10544, n10545, n10546,
    n10547, n10548, n10549, n10550, n10551, n10552,
    n10553, n10554, n10555, n10556, n10557, n10558,
    n10559, n10560, n10561, n10562, n10563, n10564,
    n10565, n10566, n10567, n10568, n10569, n10570,
    n10571, n10572, n10573, n10574, n10575, n10576,
    n10577, n10578, n10579, n10580, n10581, n10582,
    n10583, n10584, n10585, n10586, n10587, n10588,
    n10589, n10590, n10591, n10592, n10593, n10594,
    n10595, n10596, n10597, n10598, n10599, n10600,
    n10601, n10602, n10603, n10604, n10605, n10606,
    n10607, n10608, n10609, n10610, n10611, n10612,
    n10613, n10614, n10615, n10616, n10617, n10618,
    n10619, n10620, n10621, n10622, n10623, n10624,
    n10625, n10626, n10627, n10628, n10629, n10630,
    n10631, n10632, n10633, n10634, n10635, n10636,
    n10637, n10638, n10639, n10640, n10641, n10642,
    n10643, n10644, n10645, n10646, n10647, n10648,
    n10649, n10650, n10651, n10652, n10653, n10654,
    n10655, n10656, n10657, n10658, n10659, n10660,
    n10661, n10662, n10663, n10664, n10665, n10666,
    n10667, n10668, n10669, n10670, n10671, n10672,
    n10673, n10674, n10675, n10676, n10677, n10678,
    n10679, n10680, n10681, n10682, n10683, n10684,
    n10685, n10686, n10687, n10688, n10689, n10690,
    n10691, n10692, n10693, n10694, n10695, n10696,
    n10697, n10698, n10699, n10700, n10701, n10702,
    n10703, n10704, n10706, n10707, n10708, n10709,
    n10710, n10711, n10712, n10713, n10714, n10715,
    n10716, n10717, n10718, n10719, n10720, n10721,
    n10722, n10723, n10724, n10725, n10726, n10727,
    n10728, n10729, n10730, n10731, n10732, n10733,
    n10734, n10735, n10736, n10737, n10738, n10739,
    n10740, n10741, n10742, n10743, n10744, n10745,
    n10746, n10747, n10748, n10749, n10750, n10751,
    n10752, n10753, n10754, n10755, n10756, n10757,
    n10758, n10759, n10760, n10761, n10762, n10763,
    n10764, n10765, n10766, n10767, n10768, n10769,
    n10770, n10771, n10772, n10773, n10774, n10775,
    n10776, n10777, n10779, n10780, n10781, n10783,
    n10784, n10785, n10786, n10787, n10788, n10789,
    n10790, n10791, n10792, n10793, n10794, n10795,
    n10796, n10797, n10798, n10799, n10800, n10802,
    n10803, n10804, n10805, n10806, n10807, n10808,
    n10809, n10810, n10811, n10812, n10813, n10814,
    n10815, n10816, n10817, n10818, n10819, n10820,
    n10821, n10822, n10823, n10824, n10825, n10826,
    n10827, n10828, n10829, n10830, n10831, n10832,
    n10833, n10834, n10835, n10836, n10837, n10838,
    n10839, n10840, n10841, n10842, n10843, n10844,
    n10846, n10847, n10849, n10850, n10851, n10852,
    n10853, n10854, n10855, n10856, n10857, n10858,
    n10859, n10860, n10861, n10862, n10863, n10864,
    n10865, n10866, n10867, n10869, n10870, n10871,
    n10872, n10873, n10874, n10875, n10876, n10877,
    n10878, n10879, n10880, n10881, n10882, n10883,
    n10884, n10885, n10886, n10887, n10888, n10889,
    n10890, n10891, n10892, n10893, n10895, n10896,
    n10897, n10898, n10899, n10900, n10901, n10903,
    n10904, n10905, n10906, n10907, n10908, n10909,
    n10910, n10911, n10912, n10913, n10914, n10915,
    n10916, n10917, n10918, n10919, n10920, n10921,
    n10922, n10923, n10924, n10925, n10926, n10927,
    n10928, n10929, n10930, n10931, n10932, n10933,
    n10934, n10935, n10936, n10937, n10938, n10939,
    n10940, n10941, n10942, n10943, n10944, n10945,
    n10946, n10947, n10948, n10949, n10950, n10951,
    n10952, n10953, n10954, n10955, n10956, n10957,
    n10958, n10959, n10960, n10961, n10962, n10963,
    n10964, n10965, n10966, n10967, n10968, n10969,
    n10970, n10971, n10972, n10973, n10974, n10975,
    n10976, n10977, n10978, n10979, n10980, n10981,
    n10982, n10983, n10984, n10985, n10986, n10987,
    n10988, n10989, n10990, n10991, n10992, n10993,
    n10994, n10995, n10996, n10997, n10998, n10999,
    n11000, n11001, n11002, n11003, n11004, n11005,
    n11006, n11007, n11008, n11009, n11010, n11011,
    n11012, n11013, n11014, n11015, n11016, n11017,
    n11018, n11019, n11020, n11021, n11022, n11023,
    n11024, n11025, n11026, n11027, n11028, n11029,
    n11030, n11031, n11032, n11033, n11034, n11035,
    n11036, n11037, n11038, n11039, n11040, n11041,
    n11042, n11043, n11044, n11046, n11047, n11048,
    n11049, n11050, n11051, n11052, n11053, n11054,
    n11055, n11056, n11058, n11059, n11060, n11061,
    n11062, n11063, n11064, n11065, n11066, n11067,
    n11068, n11069, n11070, n11071, n11072, n11073,
    n11074, n11075, n11076, n11078, n11079, n11080,
    n11081, n11082, n11083, n11084, n11085, n11086,
    n11087, n11088, n11089, n11090, n11092, n11093,
    n11094, n11095, n11096, n11097, n11098, n11100,
    n11101, n11102, n11103, n11104, n11105, n11106,
    n11107, n11108, n11110, n11111, n11113, n11114,
    n11115, n11116, n11117, n11119, n11120, n11121,
    n11122, n11123, n11124, n11125, n11126, n11128,
    n11129, n11130, n11131, n11133, n11134, n11135,
    n11136, n11138, n11139, n11140, n11141, n11142,
    n11144, n11145, n11146, n11147, n11148, n11149,
    n11150, n11152, n11153, n11154, n11156, n11157,
    n11158, n11159, n11160, n11161, n11162, n11163,
    n11164, n11165, n11166, n11167, n11168, n11169,
    n11170, n11172, n11173, n11174, n11175, n11176,
    n11178, n11179, n11180, n11181, n11182, n11183,
    n11184, n11186, n11187, n11188, n11189, n11190,
    n11191, n11192, n11193, n11194, n11195, n11196,
    n11197, n11199, n11200, n11201, n11202, n11203,
    n11204, n11205, n11206, n11207, n11208, n11209,
    n11210, n11211, n11212, n11213, n11214, n11215,
    n11216, n11217, n11218, n11219, n11221, n11222,
    n11223, n11224, n11225, n11226, n11227, n11228,
    n11229, n11230, n11231, n11232, n11233, n11234,
    n11235, n11236, n11237, n11238, n11239, n11240,
    n11241, n11243, n11244, n11245, n11246, n11247,
    n11248, n11249, n11250, n11251, n11252, n11253,
    n11254, n11255, n11257, n11258, n11259, n11260,
    n11261, n11262, n11263, n11264, n11265, n11266,
    n11267, n11269, n11270, n11271, n11272, n11273,
    n11274, n11275, n11276, n11277, n11278, n11279,
    n11280, n11281, n11282, n11283, n11284, n11286,
    n11287, n11288, n11289, n11290, n11291, n11292,
    n11293, n11295, n11296, n11297, n11298, n11299,
    n11300, n11301, n11302, n11303, n11304, n11305,
    n11306, n11307, n11308, n11309, n11310, n11311,
    n11312, n11313, n11314, n11315, n11316, n11317,
    n11318, n11319, n11320, n11321, n11322, n11323,
    n11324, n11325, n11326, n11327, n11328, n11329,
    n11330, n11331, n11332, n11333, n11334, n11335,
    n11336, n11337, n11338, n11339, n11340, n11341,
    n11342, n11343, n11344, n11345, n11346, n11347,
    n11348, n11349, n11350, n11351, n11352, n11353,
    n11354, n11355, n11356, n11357, n11358, n11359,
    n11360, n11361, n11362, n11363, n11364, n11365,
    n11366, n11367, n11368, n11369, n11370, n11371,
    n11372, n11373, n11374, n11375, n11376, n11377,
    n11378, n11379, n11380, n11381, n11382, n11383,
    n11384, n11385, n11386, n11387, n11388, n11389,
    n11390, n11391, n11392, n11393, n11394, n11395,
    n11396, n11397, n11398, n11399, n11400, n11401,
    n11402, n11403, n11404, n11405, n11406, n11407,
    n11408, n11409, n11410, n11411, n11412, n11413,
    n11414, n11415, n11416, n11417, n11418, n11419,
    n11420, n11421, n11422, n11423, n11424, n11425,
    n11426, n11427, n11428, n11429, n11430, n11431,
    n11432, n11433, n11434, n11435, n11436, n11437,
    n11438, n11439, n11440, n11441, n11442, n11443,
    n11444, n11446, n11447, n11448, n11449, n11450,
    n11451, n11452, n11453, n11454, n11456, n11458,
    n11459, n11460, n11461, n11462, n11463, n11464,
    n11465, n11466, n11467, n11468, n11469, n11470,
    n11471, n11472, n11473, n11474, n11475, n11476,
    n11477, n11478, n11479, n11480, n11481, n11482,
    n11483, n11484, n11485, n11486, n11487, n11488,
    n11489, n11490, n11491, n11492, n11493, n11494,
    n11495, n11496, n11497, n11498, n11499, n11500,
    n11501, n11502, n11503, n11504, n11505, n11506,
    n11507, n11508, n11509, n11510, n11511, n11512,
    n11513, n11514, n11515, n11516, n11517, n11518,
    n11519, n11520, n11521, n11522, n11523, n11524,
    n11525, n11526, n11527, n11528, n11529, n11530,
    n11531, n11532, n11533, n11534, n11535, n11536,
    n11537, n11538, n11539, n11540, n11541, n11542,
    n11543, n11544, n11545, n11546, n11547, n11548,
    n11549, n11550, n11551, n11552, n11553, n11554,
    n11555, n11556, n11557, n11558, n11559, n11560,
    n11561, n11562, n11563, n11564, n11565, n11566,
    n11567, n11568, n11569, n11570, n11571, n11572,
    n11573, n11574, n11575, n11576, n11577, n11578,
    n11579, n11580, n11581, n11582, n11583, n11584,
    n11585, n11586, n11587, n11588, n11589, n11590,
    n11591, n11592, n11593, n11594, n11595, n11596,
    n11597, n11598, n11599, n11600, n11601, n11602,
    n11603, n11604, n11605, n11606, n11607, n11608,
    n11609, n11610, n11611, n11612, n11613, n11614,
    n11615, n11616, n11617, n11618, n11619, n11620,
    n11621, n11622, n11623, n11624, n11625, n11626,
    n11627, n11628, n11629, n11630, n11631, n11632,
    n11633, n11634, n11635, n11636, n11637, n11638,
    n11639, n11640, n11641, n11642, n11643, n11644,
    n11645, n11646, n11647, n11648, n11649, n11650,
    n11651, n11652, n11653, n11654, n11655, n11656,
    n11657, n11658, n11659, n11660, n11661, n11662,
    n11663, n11664, n11665, n11666, n11667, n11668,
    n11669, n11670, n11671, n11672, n11673, n11674,
    n11675, n11676, n11677, n11678, n11679, n11680,
    n11681, n11682, n11683, n11684, n11685, n11686,
    n11687, n11688, n11689, n11690, n11691, n11692,
    n11693, n11694, n11695, n11696, n11697, n11698,
    n11699, n11700, n11701, n11702, n11703, n11704,
    n11705, n11706, n11707, n11708, n11709, n11710,
    n11711, n11712, n11713, n11714, n11715, n11716,
    n11717, n11718, n11719, n11720, n11721, n11722,
    n11723, n11724, n11725, n11726, n11727, n11728,
    n11729, n11730, n11731, n11732, n11733, n11734,
    n11735, n11736, n11737, n11738, n11739, n11740,
    n11741, n11742, n11743, n11744, n11745, n11746,
    n11747, n11748, n11749, n11750, n11751, n11752,
    n11753, n11754, n11755, n11756, n11757, n11758,
    n11759, n11760, n11761, n11762, n11763, n11764,
    n11765, n11766, n11767, n11768, n11769, n11770,
    n11771, n11772, n11773, n11774, n11775, n11776,
    n11777, n11778, n11779, n11780, n11781, n11782,
    n11783, n11784, n11785, n11786, n11787, n11788,
    n11789, n11790, n11791, n11792, n11793, n11794,
    n11795, n11796, n11797, n11798, n11799, n11800,
    n11801, n11802, n11803, n11804, n11805, n11806,
    n11807, n11808, n11809, n11810, n11811, n11812,
    n11813, n11814, n11815, n11816, n11817, n11818,
    n11819, n11820, n11821, n11822, n11823, n11824,
    n11825, n11826, n11827, n11828, n11829, n11830,
    n11831, n11832, n11833, n11834, n11835, n11836,
    n11837, n11838, n11839, n11840, n11841, n11842,
    n11843, n11844, n11845, n11846, n11847, n11848,
    n11849, n11850, n11851, n11852, n11853, n11854,
    n11855, n11856, n11857, n11858, n11859, n11860,
    n11861, n11862, n11863, n11864, n11865, n11866,
    n11867, n11868, n11869, n11870, n11871, n11872,
    n11873, n11874, n11875, n11876, n11877, n11878,
    n11879, n11880, n11881, n11882, n11883, n11884,
    n11885, n11886, n11887, n11888, n11889, n11890,
    n11891, n11892, n11893, n11894, n11895, n11896,
    n11897, n11898, n11899, n11900, n11901, n11902,
    n11903, n11904, n11905, n11906, n11907, n11908,
    n11909, n11910, n11911, n11912, n11913, n11914,
    n11915, n11916, n11917, n11918, n11919, n11920,
    n11921, n11922, n11923, n11924, n11925, n11926,
    n11927, n11928, n11929, n11930, n11931, n11932,
    n11933, n11934, n11935, n11936, n11937, n11938,
    n11939, n11940, n11941, n11942, n11943, n11944,
    n11945, n11947, n11948, n11949, n11950, n11951,
    n11952, n11953, n11954, n11955, n11956, n11957,
    n11958, n11959, n11960, n11961, n11962, n11963,
    n11964, n11965, n11966, n11967, n11968, n11969,
    n11970, n11971, n11972, n11973, n11974, n11975,
    n11976, n11977, n11978, n11979, n11980, n11981,
    n11982, n11983, n11984, n11985, n11986, n11987,
    n11988, n11989, n11990, n11991, n11992, n11993,
    n11994, n11995, n11996, n11997, n11998, n11999,
    n12000, n12001, n12002, n12003, n12004, n12005,
    n12006, n12007, n12008, n12009, n12010, n12011,
    n12012, n12013, n12014, n12015, n12016, n12017,
    n12018, n12019, n12020, n12021, n12022, n12023,
    n12024, n12025, n12026, n12027, n12028, n12029,
    n12030, n12031, n12032, n12033, n12034, n12035,
    n12036, n12037, n12038, n12039, n12040, n12041,
    n12042, n12043, n12044, n12045, n12046, n12047,
    n12048, n12049, n12050, n12051, n12052, n12053,
    n12054, n12055, n12056, n12057, n12058, n12059,
    n12060, n12061, n12062, n12063, n12064, n12065,
    n12066, n12067, n12068, n12069, n12070, n12071,
    n12072, n12073, n12074, n12075, n12076, n12077,
    n12078, n12079, n12080, n12081, n12082, n12083,
    n12084, n12085, n12086, n12087, n12088, n12089,
    n12090, n12091, n12092, n12093, n12094, n12095,
    n12096, n12097, n12098, n12099, n12100, n12101,
    n12102, n12103, n12104, n12105, n12106, n12107,
    n12108, n12109, n12110, n12111, n12112, n12113,
    n12114, n12115, n12116, n12117, n12118, n12119,
    n12120, n12121, n12122, n12123, n12124, n12125,
    n12126, n12127, n12128, n12129, n12130, n12131,
    n12132, n12133, n12134, n12135, n12136, n12137,
    n12138, n12139, n12140, n12141, n12142, n12143,
    n12144, n12145, n12146, n12147, n12148, n12149,
    n12150, n12151, n12152, n12153, n12154, n12155,
    n12156, n12157, n12158, n12159, n12160, n12161,
    n12162, n12163, n12164, n12165, n12166, n12167,
    n12168, n12169, n12170, n12171, n12172, n12173,
    n12174, n12175, n12176, n12177, n12178, n12179,
    n12180, n12181, n12182, n12183, n12184, n12185,
    n12186, n12187, n12188, n12189, n12190, n12191,
    n12192, n12193, n12194, n12195, n12196, n12197,
    n12198, n12199, n12200, n12201, n12202, n12203,
    n12204, n12205, n12206, n12207, n12208, n12209,
    n12210, n12211, n12212, n12213, n12214, n12215,
    n12216, n12217, n12218, n12219, n12220, n12221,
    n12222, n12223, n12224, n12225, n12226, n12227,
    n12228, n12229, n12230, n12231, n12232, n12233,
    n12234, n12235, n12236, n12237, n12238, n12239,
    n12240, n12241, n12242, n12243, n12244, n12245,
    n12246, n12247, n12248, n12249, n12250, n12251,
    n12252, n12253, n12254, n12255, n12256, n12257,
    n12258, n12259, n12260, n12261, n12262, n12263,
    n12264, n12265, n12266, n12267, n12268, n12269,
    n12270, n12271, n12272, n12273, n12274, n12275,
    n12276, n12277, n12278, n12279, n12280, n12281,
    n12282, n12283, n12284, n12285, n12286, n12287,
    n12288, n12289, n12290, n12291, n12292, n12293,
    n12294, n12295, n12296, n12297, n12298, n12299,
    n12300, n12301, n12302, n12303, n12304, n12305,
    n12306, n12307, n12308, n12309, n12310, n12311,
    n12312, n12313, n12314, n12315, n12316, n12317,
    n12318, n12319, n12320, n12321, n12322, n12323,
    n12324, n12325, n12326, n12327, n12328, n12329,
    n12330, n12331, n12332, n12333, n12334, n12335,
    n12336, n12337, n12338, n12339, n12340, n12341,
    n12342, n12343, n12344, n12345, n12346, n12347,
    n12348, n12349, n12350, n12351, n12352, n12353,
    n12354, n12355, n12356, n12357, n12358, n12359,
    n12360, n12361, n12362, n12363, n12364, n12365,
    n12366, n12367, n12368, n12369, n12370, n12371,
    n12372, n12373, n12374, n12375, n12376, n12377,
    n12378, n12379, n12380, n12381, n12382, n12383,
    n12384, n12385, n12386, n12387, n12388, n12389,
    n12390, n12391, n12392, n12393, n12394, n12395,
    n12396, n12397, n12398, n12399, n12400, n12401,
    n12402, n12403, n12404, n12405, n12406, n12407,
    n12408, n12409, n12410, n12411, n12412, n12413,
    n12414, n12415, n12416, n12417, n12418, n12419,
    n12420, n12421, n12422, n12423, n12424, n12425,
    n12426, n12427, n12428, n12429, n12430, n12431,
    n12432, n12433, n12434, n12435, n12436, n12437,
    n12438, n12439, n12440, n12441, n12442, n12443,
    n12444, n12445, n12446, n12447, n12448, n12449,
    n12450, n12451, n12452, n12453, n12454, n12455,
    n12456, n12457, n12458, n12459, n12460, n12461,
    n12462, n12463, n12464, n12465, n12466, n12467,
    n12468, n12469, n12470, n12471, n12472, n12473,
    n12474, n12475, n12476, n12477, n12478, n12479,
    n12480, n12481, n12482, n12483, n12484, n12485,
    n12486, n12487, n12488, n12489, n12490, n12491,
    n12492, n12493, n12494, n12495, n12496, n12497,
    n12498, n12499, n12500, n12501, n12502, n12503,
    n12504, n12505, n12506, n12507, n12508, n12509,
    n12510, n12511, n12512, n12513, n12514, n12515,
    n12516, n12517, n12518, n12519, n12520, n12521,
    n12522, n12523, n12524, n12525, n12526, n12527,
    n12528, n12529, n12530, n12531, n12532, n12533,
    n12534, n12535, n12536, n12537, n12538, n12539,
    n12540, n12541, n12542, n12543, n12544, n12545,
    n12546, n12547, n12548, n12549, n12550, n12551,
    n12552, n12553, n12554, n12555, n12556, n12557,
    n12558, n12559, n12560, n12561, n12562, n12563,
    n12564, n12565, n12566, n12567, n12568, n12569,
    n12570, n12571, n12572, n12573, n12574, n12575,
    n12576, n12577, n12578, n12579, n12580, n12581,
    n12582, n12583, n12584, n12585, n12586, n12587,
    n12588, n12589, n12590, n12591, n12592, n12593,
    n12594, n12595, n12596, n12597, n12598, n12599,
    n12600, n12601, n12602, n12603, n12604, n12605,
    n12606, n12607, n12608, n12609, n12610, n12611,
    n12612, n12613, n12614, n12615, n12616, n12617,
    n12618, n12619, n12620, n12621, n12622, n12623,
    n12624, n12625, n12626, n12627, n12628, n12629,
    n12630, n12631, n12632, n12633, n12634, n12635,
    n12636, n12637, n12638, n12639, n12640, n12641,
    n12642, n12643, n12644, n12645, n12646, n12647,
    n12648, n12649, n12650, n12651, n12652, n12653,
    n12654, n12655, n12656, n12657, n12658, n12659,
    n12660, n12661, n12662, n12663, n12664, n12665,
    n12666, n12667, n12668, n12669, n12670, n12671,
    n12672, n12673, n12674, n12675, n12676, n12677,
    n12678, n12679, n12680, n12681, n12682, n12683,
    n12684, n12685, n12686, n12687, n12688, n12689,
    n12690, n12691, n12692, n12693, n12694, n12695,
    n12696, n12697, n12698, n12699, n12700, n12701,
    n12702, n12703, n12704, n12705, n12706, n12707,
    n12708, n12709, n12710, n12711, n12713, n12714,
    n12715, n12716, n12717, n12718, n12719, n12720,
    n12722, n12723, n12724, n12725, n12726, n12727,
    n12728, n12730, n12731, n12732, n12733, n12734,
    n12735, n12736, n12737, n12738, n12739, n12740,
    n12741, n12743, n12744, n12745, n12746, n12747,
    n12749, n12750, n12751, n12752, n12754, n12755,
    n12756, n12758, n12759, n12760, n12761, n12763,
    n12764, n12765, n12766, n12767, n12768, n12769,
    n12770, n12771, n12772, n12773, n12774, n12775,
    n12776, n12777, n12778, n12779, n12780, n12782,
    n12783, n12784, n12785, n12786, n12787, n12788,
    n12790, n12791, n12792, n12793, n12795, n12796,
    n12797, n12798, n12799, n12800, n12801, n12802,
    n12803, n12804, n12806, n12807, n12808, n12809,
    n12810, n12811, n12812, n12813, n12814, n12815,
    n12816, n12817, n12819, n12820, n12821, n12822,
    n12823, n12824, n12825, n12827, n12828, n12829,
    n12830, n12831, n12832, n12833, n12834, n12835,
    n12836, n12837, n12838, n12839, n12840, n12841,
    n12842, n12844, n12845, n12846, n12847, n12848,
    n12849, n12850, n12851, n12852, n12853, n12854,
    n12855, n12856, n12857, n12858, n12859, n12860,
    n12862, n12863, n12864, n12865, n12866, n12867,
    n12868, n12869, n12870, n12871, n12872, n12873,
    n12874, n12876, n12877, n12878, n12879, n12880,
    n12881, n12882, n12883, n12884, n12886, n12887,
    n12888, n12889, n12891, n12892, n12893, n12894,
    n12895, n12896, n12897, n12898, n12899, n12900,
    n12901, n12902, n12903, n12904, n12905, n12906,
    n12907, n12908, n12909, n12910, n12911, n12912,
    n12913, n12914, n12915, n12916, n12917, n12918,
    n12919, n12920, n12921, n12922, n12923, n12924,
    n12925, n12926, n12927, n12928, n12929, n12930,
    n12931, n12932, n12933, n12934, n12935, n12936,
    n12937, n12938, n12939, n12940, n12941, n12942,
    n12943, n12944, n12945, n12946, n12947, n12948,
    n12949, n12950, n12951, n12952, n12953, n12954,
    n12955, n12956, n12957, n12958, n12959, n12960,
    n12961, n12962, n12963, n12964, n12966, n12967,
    n12968, n12969, n12970, n12971, n12972, n12973,
    n12974, n12975, n12976, n12977, n12978, n12979,
    n12981, n12982, n12983, n12984, n12985, n12986,
    n12987, n12988, n12989, n12990, n12991, n12992,
    n12993, n12994, n12995, n12996, n12997, n12998,
    n12999, n13000, n13001, n13002, n13003, n13004,
    n13005, n13006, n13007, n13008, n13009, n13010,
    n13011, n13012, n13013, n13014, n13015, n13016,
    n13017, n13018, n13019, n13020, n13021, n13022,
    n13023, n13024, n13025, n13026, n13027, n13028,
    n13029, n13030, n13031, n13032, n13033, n13034,
    n13035, n13036, n13037, n13038, n13039, n13040,
    n13041, n13042, n13043, n13044, n13045, n13046,
    n13047, n13048, n13049, n13050, n13051, n13052,
    n13053, n13054, n13055, n13056, n13058, n13060,
    n13061, n13062, n13063, n13064, n13065, n13066,
    n13068, n13069, n13070, n13071, n13072, n13073,
    n13074, n13075, n13076, n13077, n13078, n13080,
    n13081, n13082, n13083, n13084, n13085, n13086,
    n13087, n13088, n13090, n13092, n13093, n13094,
    n13095, n13096, n13097, n13098, n13099, n13100,
    n13101, n13102, n13103, n13104, n13105, n13106,
    n13107, n13108, n13110, n13112, n13113, n13114,
    n13115, n13116, n13117, n13118, n13119, n13121,
    n13122, n13123, n13124, n13125, n13128, n13129,
    n13130, n13131, n13132, n13133, n13134, n13135,
    n13136, n13137, n13138, n13139, n13140, n13141,
    n13142, n13143, n13144, n13145, n13146, n13147,
    n13148, n13149, n13150, n13151, n13152, n13153,
    n13154, n13155, n13156, n13157, n13158, n13159,
    n13160, n13161, n13162, n13163, n13164, n13165,
    n13166, n13167, n13168, n13169, n13170, n13171,
    n13172, n13173, n13174, n13175, n13176, n13177,
    n13179, n13180, n13181, n13182, n13183, n13184,
    n13185, n13186, n13187, n13188, n13189, n13190,
    n13191, n13192, n13193, n13194, n13195, n13196,
    n13197, n13198, n13199, n13200, n13201, n13202,
    n13203, n13204, n13205, n13206, n13207, n13208,
    n13209, n13210, n13211, n13212, n13213, n13214,
    n13215, n13216, n13217, n13218, n13219, n13220,
    n13222, n13223, n13224, n13225, n13226, n13227,
    n13228, n13229, n13230, n13231, n13232, n13233,
    n13234, n13235, n13236, n13237, n13238, n13239,
    n13240, n13241, n13242, n13243, n13244, n13245,
    n13246, n13247, n13248, n13249, n13250, n13251,
    n13252, n13253, n13254, n13255, n13256, n13257,
    n13258, n13259, n13260, n13261, n13262, n13264,
    n13265, n13266, n13267, n13268, n13269, n13270,
    n13271, n13272, n13273, n13274, n13275, n13276,
    n13277, n13278, n13279, n13280, n13281, n13282,
    n13283, n13284, n13285, n13286, n13287, n13288,
    n13289, n13290, n13291, n13292, n13293, n13294,
    n13295, n13296, n13297, n13298, n13299, n13300,
    n13301, n13302, n13303, n13304, n13306, n13307,
    n13308, n13309, n13310, n13311, n13312, n13313,
    n13314, n13315, n13316, n13317, n13318, n13319,
    n13321, n13322, n13323, n13324, n13325, n13326,
    n13327, n13328, n13329, n13330, n13331, n13332,
    n13333, n13334, n13335, n13336, n13337, n13338,
    n13339, n13340, n13341, n13342, n13343, n13344,
    n13345, n13346, n13347, n13348, n13349, n13350,
    n13351, n13352, n13353, n13354, n13355, n13356,
    n13357, n13358, n13359, n13360, n13361, n13362,
    n13363, n13364, n13365, n13366, n13367, n13368,
    n13369, n13370, n13371, n13372, n13373, n13374,
    n13375, n13376, n13377, n13378, n13379, n13380,
    n13381, n13382, n13383, n13384, n13385, n13386,
    n13387, n13388, n13389, n13390, n13391, n13392,
    n13393, n13394, n13395, n13396, n13397, n13398,
    n13399, n13400, n13401, n13402, n13403, n13404,
    n13405, n13406, n13407, n13408, n13409, n13410,
    n13411, n13412, n13413, n13414, n13415, n13416,
    n13417, n13418, n13419, n13420, n13421, n13422,
    n13423, n13424, n13425, n13426, n13427, n13428,
    n13429, n13430, n13431, n13432, n13433, n13434,
    n13435, n13436, n13437, n13438, n13439, n13440,
    n13441, n13442, n13443, n13444, n13445, n13446,
    n13447, n13448, n13449, n13450, n13451, n13452,
    n13453, n13454, n13455, n13456, n13457, n13458,
    n13459, n13460, n13461, n13462, n13463, n13464,
    n13465, n13466, n13467, n13468, n13469, n13470,
    n13471, n13472, n13473, n13474, n13475, n13476,
    n13477, n13478, n13479, n13480, n13481, n13482,
    n13483, n13484, n13485, n13486, n13487, n13488,
    n13489, n13490, n13491, n13492, n13493, n13494,
    n13495, n13496, n13497, n13498, n13499, n13500,
    n13501, n13502, n13503, n13504, n13505, n13506,
    n13507, n13508, n13509, n13510, n13511, n13512,
    n13513, n13514, n13515, n13516, n13517, n13518,
    n13519, n13520, n13521, n13522, n13523, n13524,
    n13525, n13526, n13527, n13528, n13529, n13530,
    n13531, n13532, n13533, n13534, n13535, n13536,
    n13537, n13538, n13539, n13540, n13541, n13542,
    n13543, n13544, n13545, n13546, n13547, n13548,
    n13549, n13550, n13551, n13552, n13553, n13554,
    n13555, n13556, n13557, n13558, n13559, n13560,
    n13561, n13562, n13563, n13564, n13565, n13566,
    n13567, n13568, n13569, n13570, n13571, n13572,
    n13573, n13574, n13575, n13576, n13577, n13578,
    n13579, n13580, n13581, n13582, n13583, n13584,
    n13585, n13586, n13587, n13588, n13589, n13590,
    n13591, n13592, n13593, n13594, n13595, n13596,
    n13597, n13598, n13599, n13600, n13601, n13602,
    n13603, n13604, n13605, n13606, n13607, n13608,
    n13609, n13610, n13611, n13612, n13613, n13615,
    n13616, n13617, n13618, n13619, n13620, n13621,
    n13622, n13623, n13624, n13625, n13626, n13627,
    n13628, n13629, n13630, n13631, n13632, n13633,
    n13634, n13635, n13636, n13637, n13638, n13639,
    n13640, n13641, n13642, n13643, n13644, n13645,
    n13646, n13647, n13648, n13649, n13650, n13651,
    n13652, n13653, n13654, n13655, n13656, n13657,
    n13658, n13659, n13660, n13661, n13662, n13663,
    n13664, n13665, n13666, n13668, n13669, n13670,
    n13671, n13672, n13673, n13674, n13675, n13676,
    n13677, n13678, n13679, n13680, n13681, n13682,
    n13683, n13684, n13685, n13686, n13687, n13688,
    n13689, n13690, n13691, n13692, n13693, n13694,
    n13695, n13696, n13697, n13698, n13699, n13700,
    n13701, n13702, n13703, n13704, n13705, n13706,
    n13707, n13708, n13709, n13710, n13711, n13712,
    n13713, n13714, n13715, n13716, n13717, n13718,
    n13719, n13720, n13721, n13722, n13723, n13724,
    n13725, n13726, n13727, n13728, n13729, n13730,
    n13731, n13732, n13733, n13734, n13735, n13736,
    n13737, n13738, n13739, n13740, n13741, n13742,
    n13743, n13744, n13745, n13746, n13747, n13748,
    n13749, n13750, n13751, n13752, n13753, n13754,
    n13755, n13756, n13757, n13758, n13759, n13760,
    n13761, n13762, n13763, n13764, n13765, n13766,
    n13767, n13768, n13769, n13770, n13771, n13772,
    n13773, n13774, n13775, n13776, n13777, n13778,
    n13779, n13780, n13781, n13782, n13783, n13784,
    n13785, n13786, n13787, n13788, n13789, n13790,
    n13791, n13792, n13793, n13794, n13795, n13796,
    n13797, n13798, n13799, n13800, n13801, n13802,
    n13803, n13804, n13805, n13806, n13807, n13808,
    n13809, n13810, n13811, n13812, n13813, n13814,
    n13815, n13816, n13817, n13818, n13819, n13820,
    n13821, n13822, n13823, n13824, n13825, n13826,
    n13827, n13828, n13829, n13830, n13831, n13832,
    n13833, n13834, n13835, n13836, n13837, n13838,
    n13839, n13840, n13841, n13842, n13843, n13844,
    n13845, n13846, n13847, n13848, n13849, n13850,
    n13851, n13852, n13853, n13854, n13855, n13856,
    n13857, n13858, n13859, n13860, n13861, n13862,
    n13863, n13864, n13865, n13866, n13867, n13868,
    n13869, n13870, n13871, n13872, n13873, n13874,
    n13875, n13876, n13877, n13878, n13879, n13880,
    n13881, n13882, n13883, n13884, n13885, n13886,
    n13887, n13888, n13889, n13890, n13891, n13892,
    n13893, n13894, n13895, n13896, n13897, n13898,
    n13899, n13900, n13901, n13902, n13903, n13904,
    n13905, n13906, n13907, n13908, n13909, n13910,
    n13911, n13912, n13913, n13914, n13915, n13916,
    n13917, n13918, n13919, n13920, n13921, n13922,
    n13923, n13924, n13925, n13926, n13927, n13928,
    n13929, n13930, n13931, n13932, n13933, n13934,
    n13935, n13936, n13937, n13938, n13939, n13940,
    n13941, n13942, n13943, n13944, n13945, n13946,
    n13947, n13948, n13949, n13950, n13951, n13952,
    n13953, n13954, n13955, n13956, n13957, n13958,
    n13959, n13960, n13961, n13962, n13963, n13964,
    n13965, n13966, n13967, n13968, n13969, n13970,
    n13971, n13972, n13973, n13974, n13975, n13976,
    n13977, n13978, n13979, n13980, n13981, n13982,
    n13983, n13984, n13985, n13986, n13988, n13989,
    n13990, n13991, n13992, n13993, n13994, n13995,
    n13996, n13997, n13998, n13999, n14000, n14001,
    n14002, n14003, n14004, n14005, n14006, n14007,
    n14008, n14009, n14010, n14011, n14012, n14013,
    n14014, n14015, n14016, n14017, n14018, n14019,
    n14020, n14021, n14022, n14023, n14024, n14025,
    n14026, n14027, n14028, n14029, n14030, n14031,
    n14032, n14033, n14034, n14035, n14036, n14037,
    n14038, n14039, n14040, n14041, n14042, n14043,
    n14044, n14045, n14046, n14047, n14048, n14049,
    n14050, n14051, n14052, n14053, n14054, n14055,
    n14056, n14057, n14058, n14059, n14060, n14061,
    n14062, n14063, n14064, n14065, n14066, n14067,
    n14068, n14069, n14070, n14071, n14072, n14073,
    n14074, n14075, n14076, n14077, n14078, n14079,
    n14080, n14081, n14082, n14083, n14084, n14085,
    n14086, n14087, n14088, n14089, n14090, n14091,
    n14092, n14093, n14094, n14095, n14096, n14097,
    n14098, n14099, n14100, n14101, n14102, n14103,
    n14104, n14105, n14106, n14107, n14108, n14109,
    n14110, n14111, n14112, n14113, n14114, n14115,
    n14116, n14117, n14118, n14119, n14120, n14121,
    n14122, n14123, n14124, n14125, n14126, n14127,
    n14128, n14129, n14130, n14131, n14132, n14133,
    n14134, n14135, n14136, n14137, n14138, n14139,
    n14140, n14141, n14142, n14143, n14144, n14145,
    n14146, n14147, n14148, n14149, n14150, n14151,
    n14152, n14153, n14154, n14155, n14156, n14157,
    n14158, n14159, n14160, n14161, n14162, n14163,
    n14164, n14165, n14166, n14167, n14168, n14169,
    n14170, n14171, n14172, n14173, n14174, n14175,
    n14176, n14177, n14178, n14179, n14180, n14181,
    n14182, n14183, n14184, n14185, n14186, n14187,
    n14188, n14189, n14190, n14191, n14192, n14193,
    n14194, n14195, n14196, n14197, n14198, n14199,
    n14200, n14201, n14202, n14203, n14204, n14205,
    n14206, n14207, n14208, n14209, n14210, n14211,
    n14212, n14213, n14214, n14215, n14216, n14217,
    n14218, n14219, n14220, n14221, n14222, n14223,
    n14224, n14225, n14226, n14227, n14228, n14229,
    n14230, n14231, n14232, n14233, n14234, n14235,
    n14236, n14237, n14238, n14239, n14240, n14241,
    n14242, n14243, n14244, n14245, n14246, n14247,
    n14248, n14249, n14250, n14251, n14252, n14253,
    n14254, n14255, n14256, n14257, n14258, n14259,
    n14260, n14261, n14262, n14263, n14264, n14265,
    n14266, n14267, n14268, n14269, n14270, n14271,
    n14272, n14273, n14274, n14275, n14276, n14277,
    n14278, n14279, n14280, n14281, n14282, n14283,
    n14284, n14285, n14286, n14287, n14288, n14289,
    n14290, n14291, n14292, n14293, n14294, n14295,
    n14296, n14297, n14298, n14299, n14300, n14301,
    n14302, n14303, n14304, n14305, n14306, n14307,
    n14308, n14309, n14310, n14311, n14312, n14313,
    n14314, n14315, n14316, n14317, n14318, n14319,
    n14320, n14321, n14322, n14323, n14324, n14325,
    n14326, n14327, n14328, n14329, n14330, n14331,
    n14332, n14333, n14334, n14335, n14336, n14337,
    n14338, n14339, n14340, n14341, n14342, n14343,
    n14344, n14345, n14346, n14347, n14348, n14349,
    n14350, n14351, n14352, n14353, n14354, n14355,
    n14356, n14357, n14358, n14359, n14360, n14361,
    n14362, n14363, n14364, n14365, n14366, n14367,
    n14368, n14369, n14370, n14371, n14372, n14373,
    n14374, n14375, n14376, n14377, n14378, n14379,
    n14380, n14381, n14382, n14383, n14384, n14386,
    n14387, n14388, n14389, n14390, n14391, n14392,
    n14394, n14395, n14396, n14397, n14398, n14399,
    n14400, n14401, n14402, n14403, n14404, n14405,
    n14406, n14407, n14408, n14409, n14410, n14411,
    n14412, n14413, n14414, n14415, n14416, n14417,
    n14418, n14419, n14420, n14421, n14422, n14423,
    n14424, n14425, n14426, n14427, n14428, n14429,
    n14430, n14431, n14432, n14433, n14434, n14435,
    n14436, n14437, n14438, n14439, n14440, n14441,
    n14442, n14443, n14444, n14446, n14447, n14448,
    n14449, n14450, n14451, n14452, n14453, n14454,
    n14455, n14456, n14457, n14458, n14459, n14460,
    n14461, n14462, n14463, n14464, n14465, n14466,
    n14467, n14468, n14469, n14470, n14471, n14472,
    n14473, n14474, n14475, n14476, n14477, n14478,
    n14479, n14480, n14481, n14482, n14483, n14484,
    n14485, n14486, n14487, n14488, n14489, n14490,
    n14491, n14492, n14493, n14494, n14495, n14496,
    n14497, n14498, n14499, n14500, n14501, n14502,
    n14503, n14504, n14505, n14506, n14507, n14508,
    n14509, n14510, n14511, n14512, n14513, n14514,
    n14515, n14516, n14517, n14518, n14519, n14520,
    n14521, n14522, n14523, n14524, n14525, n14526,
    n14527, n14528, n14529, n14530, n14531, n14532,
    n14533, n14534, n14535, n14536, n14537, n14538,
    n14539, n14540, n14541, n14542, n14543, n14544,
    n14545, n14546, n14547, n14548, n14549, n14550,
    n14551, n14552, n14553, n14554, n14555, n14556,
    n14557, n14558, n14559, n14560, n14561, n14562,
    n14563, n14564, n14565, n14566, n14567, n14568,
    n14569, n14570, n14571, n14572, n14573, n14574,
    n14575, n14576, n14577, n14578, n14579, n14580,
    n14581, n14582, n14583, n14584, n14585, n14586,
    n14587, n14588, n14589, n14590, n14591, n14592,
    n14593, n14594, n14595, n14596, n14597, n14598,
    n14599, n14600, n14601, n14602, n14603, n14604,
    n14605, n14606, n14607, n14608, n14609, n14610,
    n14611, n14612, n14613, n14614, n14615, n14616,
    n14617, n14618, n14619, n14620, n14621, n14622,
    n14623, n14624, n14625, n14626, n14627, n14628,
    n14629, n14630, n14631, n14632, n14633, n14634,
    n14635, n14636, n14637, n14638, n14639, n14640,
    n14641, n14642, n14643, n14644, n14645, n14646,
    n14647, n14648, n14649, n14650, n14651, n14652,
    n14653, n14654, n14655, n14656, n14657, n14658,
    n14659, n14660, n14661, n14662, n14663, n14664,
    n14665, n14666, n14667, n14668, n14669, n14670,
    n14671, n14672, n14673, n14674, n14675, n14676,
    n14677, n14678, n14679, n14680, n14681, n14682,
    n14683, n14684, n14685, n14686, n14687, n14688,
    n14689, n14690, n14691, n14692, n14693, n14694,
    n14695, n14696, n14697, n14698, n14699, n14700,
    n14701, n14702, n14703, n14704, n14705, n14706,
    n14707, n14708, n14709, n14710, n14711, n14712,
    n14713, n14714, n14715, n14716, n14717, n14718,
    n14719, n14720, n14721, n14722, n14723, n14724,
    n14725, n14726, n14727, n14728, n14729, n14730,
    n14731, n14732, n14733, n14734, n14735, n14736,
    n14737, n14738, n14739, n14740, n14741, n14742,
    n14743, n14744, n14745, n14746, n14747, n14748,
    n14749, n14750, n14751, n14752, n14753, n14754,
    n14755, n14756, n14757, n14758, n14759, n14760,
    n14761, n14762, n14763, n14764, n14765, n14766,
    n14767, n14768, n14769, n14770, n14771, n14772,
    n14773, n14774, n14775, n14776, n14777, n14778,
    n14779, n14780, n14781, n14782, n14783, n14784,
    n14785, n14786, n14787, n14788, n14789, n14790,
    n14791, n14792, n14793, n14794, n14795, n14796,
    n14797, n14798, n14799, n14800, n14801, n14802,
    n14803, n14804, n14805, n14806, n14807, n14808,
    n14809, n14810, n14811, n14812, n14813, n14814,
    n14815, n14816, n14817, n14818, n14819, n14820,
    n14821, n14822, n14823, n14824, n14825, n14826,
    n14827, n14828, n14829, n14830, n14831, n14832,
    n14833, n14834, n14835, n14836, n14838, n14839,
    n14840, n14841, n14842, n14843, n14844, n14845,
    n14846, n14847, n14848, n14849, n14850, n14851,
    n14852, n14853, n14854, n14855, n14856, n14857,
    n14858, n14859, n14860, n14861, n14862, n14863,
    n14864, n14865, n14866, n14867, n14868, n14869,
    n14870, n14871, n14872, n14873, n14874, n14875,
    n14876, n14877, n14878, n14879, n14880, n14881,
    n14882, n14883, n14884, n14885, n14886, n14887,
    n14888, n14889, n14890, n14891, n14892, n14893,
    n14894, n14895, n14896, n14897, n14898, n14899,
    n14900, n14901, n14902, n14903, n14904, n14905,
    n14906, n14907, n14908, n14909, n14910, n14911,
    n14912, n14913, n14914, n14915, n14916, n14917,
    n14918, n14919, n14920, n14921, n14922, n14923,
    n14924, n14925, n14926, n14927, n14928, n14929,
    n14930, n14931, n14932, n14933, n14934, n14935,
    n14936, n14937, n14938, n14939, n14940, n14941,
    n14942, n14943, n14944, n14945, n14946, n14947,
    n14948, n14949, n14950, n14951, n14952, n14953,
    n14954, n14955, n14956, n14957, n14958, n14959,
    n14960, n14961, n14962, n14963, n14964, n14965,
    n14966, n14967, n14968, n14969, n14970, n14971,
    n14972, n14973, n14974, n14975, n14976, n14977,
    n14978, n14979, n14980, n14981, n14982, n14983,
    n14984, n14985, n14986, n14987, n14988, n14989,
    n14990, n14991, n14992, n14993, n14994, n14995,
    n14996, n14997, n14998, n14999, n15000, n15001,
    n15002, n15003, n15004, n15005, n15006, n15007,
    n15008, n15009, n15010, n15011, n15012, n15013,
    n15014, n15015, n15016, n15017, n15018, n15019,
    n15020, n15021, n15022, n15023, n15024, n15025,
    n15026, n15027, n15028, n15029, n15030, n15031,
    n15032, n15033, n15034, n15035, n15036, n15037,
    n15038, n15039, n15040, n15041, n15042, n15043,
    n15044, n15045, n15046, n15047, n15048, n15049,
    n15050, n15051, n15052, n15053, n15054, n15055,
    n15056, n15057, n15058, n15059, n15060, n15061,
    n15062, n15063, n15064, n15065, n15066, n15067,
    n15068, n15069, n15070, n15071, n15072, n15073,
    n15074, n15075, n15076, n15077, n15078, n15079,
    n15080, n15081, n15082, n15083, n15084, n15085,
    n15086, n15087, n15088, n15089, n15090, n15091,
    n15092, n15093, n15094, n15095, n15096, n15097,
    n15098, n15099, n15100, n15101, n15102, n15103,
    n15104, n15105, n15106, n15107, n15108, n15109,
    n15110, n15111, n15112, n15113, n15114, n15115,
    n15116, n15117, n15118, n15119, n15120, n15121,
    n15122, n15123, n15124, n15125, n15126, n15127,
    n15128, n15129, n15130, n15131, n15133, n15134,
    n15135, n15136, n15137, n15138, n15139, n15140,
    n15141, n15142, n15143, n15144, n15145, n15146,
    n15147, n15148, n15149, n15150, n15151, n15152,
    n15153, n15154, n15155, n15156, n15157, n15158,
    n15159, n15160, n15161, n15162, n15163, n15164,
    n15165, n15166, n15167, n15168, n15169, n15170,
    n15171, n15172, n15173, n15174, n15175, n15176,
    n15177, n15178, n15179, n15180, n15181, n15182,
    n15183, n15184, n15185, n15186, n15187, n15188,
    n15189, n15190, n15191, n15192, n15193, n15194,
    n15195, n15196, n15197, n15198, n15199, n15200,
    n15201, n15202, n15203, n15204, n15205, n15206,
    n15207, n15208, n15209, n15210, n15211, n15212,
    n15213, n15214, n15215, n15216, n15217, n15218,
    n15219, n15220, n15221, n15222, n15223, n15224,
    n15225, n15227, n15228, n15229, n15230, n15231,
    n15232, n15233, n15234, n15235, n15236, n15237,
    n15238, n15239, n15240, n15241, n15242, n15243,
    n15244, n15245, n15246, n15247, n15248, n15249,
    n15251, n15252, n15253, n15254, n15255, n15256,
    n15257, n15258, n15259, n15260, n15261, n15262,
    n15263, n15264, n15265, n15266, n15267, n15268,
    n15269, n15270, n15271, n15272, n15273, n15274,
    n15275, n15276, n15277, n15278, n15279, n15280,
    n15281, n15282, n15283, n15284, n15285, n15286,
    n15287, n15288, n15289, n15290, n15291, n15292,
    n15293, n15294, n15295, n15296, n15297, n15298,
    n15299, n15300, n15301, n15302, n15303, n15304,
    n15305, n15306, n15307, n15308, n15309, n15310,
    n15311, n15312, n15313, n15314, n15315, n15316,
    n15317, n15318, n15319, n15320, n15321, n15322,
    n15323, n15324, n15325, n15326, n15327, n15328,
    n15329, n15330, n15331, n15332, n15333, n15334,
    n15335, n15336, n15337, n15338, n15339, n15340,
    n15341, n15342, n15343, n15344, n15345, n15346,
    n15347, n15348, n15349, n15350, n15351, n15352,
    n15353, n15354, n15355, n15356, n15357, n15358,
    n15359, n15360, n15361, n15362, n15363, n15364,
    n15365, n15366, n15367, n15368, n15369, n15370,
    n15372, n15373, n15374, n15375, n15376, n15377,
    n15379, n15380, n15381, n15382, n15383, n15384,
    n15385, n15386, n15387, n15388, n15389, n15390,
    n15391, n15392, n15393, n15394, n15395, n15396,
    n15397, n15398, n15399, n15400, n15401, n15402,
    n15403, n15404, n15405, n15406, n15407, n15408,
    n15409, n15410, n15411, n15412, n15413, n15414,
    n15415, n15416, n15417, n15418, n15419, n15420,
    n15421, n15422, n15423, n15424, n15425, n15426,
    n15427, n15428, n15429, n15430, n15431, n15432,
    n15433, n15434, n15435, n15436, n15437, n15438,
    n15439, n15440, n15441, n15442, n15443, n15444,
    n15445, n15446, n15447, n15448, n15449, n15450,
    n15451, n15452, n15453, n15454, n15455, n15456,
    n15457, n15458, n15459, n15460, n15461, n15462,
    n15463, n15464, n15465, n15466, n15467, n15468,
    n15469, n15470, n15471, n15472, n15473, n15474,
    n15475, n15476, n15477, n15478, n15479, n15480,
    n15481, n15482, n15483, n15484, n15485, n15486,
    n15487, n15488, n15489, n15490, n15491, n15492,
    n15493, n15494, n15495, n15496, n15497, n15498,
    n15499, n15500, n15501, n15502, n15503, n15504,
    n15505, n15506, n15507, n15508, n15509, n15510,
    n15511, n15512, n15513, n15514, n15515, n15516,
    n15517, n15518, n15519, n15520, n15521, n15522,
    n15523, n15524, n15525, n15526, n15527, n15528,
    n15529, n15530, n15531, n15532, n15533, n15534,
    n15535, n15536, n15537, n15538, n15539, n15540,
    n15541, n15542, n15543, n15544, n15545, n15546,
    n15547, n15548, n15549, n15550, n15551, n15552,
    n15553, n15554, n15555, n15556, n15557, n15558,
    n15559, n15560, n15561, n15562, n15563, n15564,
    n15565, n15566, n15567, n15568, n15569, n15570,
    n15571, n15572, n15573, n15574, n15575, n15576,
    n15577, n15578, n15579, n15580, n15581, n15582,
    n15583, n15584, n15585, n15586, n15587, n15588,
    n15589, n15591, n15592, n15593, n15594, n15595,
    n15596, n15597, n15598, n15599, n15600, n15601,
    n15602, n15603, n15604, n15605, n15606, n15607,
    n15608, n15609, n15610, n15611, n15612, n15613,
    n15614, n15615, n15616, n15617, n15618, n15619,
    n15620, n15621, n15622, n15623, n15624, n15625,
    n15626, n15627, n15628, n15629, n15630, n15631,
    n15632, n15633, n15634, n15635, n15636, n15637,
    n15638, n15639, n15640, n15641, n15642, n15643,
    n15644, n15645, n15646, n15647, n15648, n15649,
    n15650, n15652, n15653, n15654, n15655, n15656,
    n15657, n15658, n15659, n15660, n15661, n15662,
    n15663, n15664, n15665, n15666, n15667, n15668,
    n15669, n15670, n15671, n15672, n15673, n15674,
    n15675, n15676, n15677, n15678, n15679, n15680,
    n15681, n15682, n15683, n15684, n15685, n15686,
    n15687, n15688, n15689, n15690, n15691, n15692,
    n15693, n15694, n15695, n15696, n15697, n15698,
    n15699, n15700, n15701, n15702, n15703, n15704,
    n15705, n15706, n15707, n15708, n15709, n15710,
    n15711, n15712, n15713, n15714, n15715, n15716,
    n15717, n15718, n15719, n15720, n15721, n15722,
    n15723, n15724, n15725, n15726, n15727, n15728,
    n15729, n15730, n15731, n15732, n15733, n15734,
    n15735, n15736, n15737, n15738, n15739, n15740,
    n15741, n15742, n15743, n15744, n15745, n15746,
    n15747, n15748, n15749, n15750, n15751, n15752,
    n15753, n15754, n15755, n15756, n15757, n15758,
    n15759, n15760, n15761, n15762, n15763, n15764,
    n15766, n15767, n15768, n15769, n15770, n15771,
    n15772, n15773, n15774, n15775, n15776, n15777,
    n15778, n15779, n15780, n15781, n15782, n15783,
    n15784, n15785, n15786, n15787, n15788, n15789,
    n15790, n15791, n15792, n15793, n15794, n15795,
    n15796, n15797, n15798, n15799, n15800, n15801,
    n15802, n15803, n15804, n15805, n15806, n15807,
    n15808, n15809, n15810, n15811, n15812, n15813,
    n15814, n15815, n15816, n15817, n15818, n15819,
    n15820, n15821, n15822, n15823, n15824, n15825,
    n15826, n15827, n15828, n15829, n15830, n15831,
    n15832, n15833, n15834, n15835, n15836, n15837,
    n15838, n15839, n15840, n15841, n15842, n15843,
    n15844, n15845, n15846, n15847, n15848, n15849,
    n15850, n15851, n15852, n15853, n15854, n15855,
    n15856, n15857, n15858, n15859, n15860, n15861,
    n15862, n15863, n15864, n15865, n15866, n15867,
    n15868, n15869, n15870, n15871, n15872, n15873,
    n15874, n15875, n15876, n15877, n15878, n15879,
    n15880, n15881, n15882, n15883, n15885, n15886,
    n15887, n15888, n15889, n15890, n15891, n15892,
    n15893, n15894, n15895, n15896, n15897, n15898,
    n15899, n15900, n15901, n15902, n15903, n15904,
    n15905, n15906, n15907, n15908, n15909, n15910,
    n15911, n15912, n15913, n15914, n15915, n15916,
    n15917, n15918, n15919, n15920, n15921, n15922,
    n15923, n15924, n15925, n15926, n15927, n15928,
    n15929, n15930, n15931, n15932, n15933, n15934,
    n15935, n15936, n15937, n15938, n15939, n15940,
    n15941, n15942, n15943, n15944, n15945, n15946,
    n15947, n15948, n15949, n15950, n15951, n15952,
    n15953, n15954, n15955, n15956, n15957, n15958,
    n15959, n15960, n15961, n15962, n15963, n15964,
    n15965, n15966, n15967, n15968, n15970, n15971,
    n15972, n15973, n15974, n15975, n15976, n15977,
    n15978, n15979, n15980, n15981, n15983, n15984,
    n15985, n15986, n15987, n15988, n15989, n15990,
    n15991, n15992, n15993, n15994, n15995, n15996,
    n15997, n15998, n15999, n16000, n16001, n16002,
    n16003, n16004, n16005, n16006, n16007, n16008,
    n16009, n16010, n16011, n16012, n16013, n16014,
    n16015, n16016, n16017, n16018, n16019, n16020,
    n16021, n16022, n16023, n16024, n16025, n16026,
    n16027, n16028, n16029, n16030, n16031, n16032,
    n16033, n16034, n16035, n16036, n16037, n16038,
    n16039, n16040, n16041, n16042, n16043, n16044,
    n16045, n16046, n16047, n16048, n16049, n16050,
    n16051, n16052, n16053, n16054, n16055, n16056,
    n16057, n16058, n16059, n16060, n16061, n16062,
    n16063, n16064, n16065, n16067, n16068, n16069,
    n16070, n16071, n16072, n16073, n16074, n16075,
    n16076, n16077, n16078, n16079, n16080, n16081,
    n16082, n16083, n16084, n16085, n16086, n16087,
    n16088, n16089, n16090, n16091, n16092, n16093,
    n16094, n16095, n16096, n16097, n16098, n16099,
    n16100, n16101, n16102, n16103, n16104, n16105,
    n16106, n16107, n16108, n16109, n16110, n16111,
    n16112, n16113, n16114, n16115, n16116, n16117,
    n16118, n16119, n16121, n16122, n16123, n16124,
    n16125, n16126, n16127, n16128, n16129, n16130,
    n16131, n16132, n16133, n16134, n16135, n16136,
    n16137, n16138, n16139, n16140, n16141, n16142,
    n16143, n16144, n16145, n16146, n16147, n16148,
    n16149, n16150, n16151, n16152, n16153, n16154,
    n16155, n16156, n16157, n16158, n16159, n16160,
    n16161, n16162, n16163, n16164, n16165, n16166,
    n16167, n16168, n16169, n16171, n16172, n16173,
    n16174, n16175, n16176, n16177, n16178, n16179,
    n16180, n16181, n16182, n16183, n16184, n16185,
    n16186, n16187, n16188, n16189, n16190, n16191,
    n16192, n16193, n16194, n16195, n16196, n16197,
    n16198, n16199, n16200, n16201, n16202, n16203,
    n16204, n16205, n16206, n16207, n16208, n16209,
    n16210, n16211, n16212, n16213, n16214, n16215,
    n16216, n16217, n16218, n16219, n16220, n16221,
    n16222, n16223, n16224, n16225, n16226, n16227,
    n16228, n16229, n16230, n16231, n16232, n16233,
    n16234, n16235, n16236, n16237, n16238, n16239,
    n16240, n16241, n16242, n16243, n16244, n16245,
    n16246, n16247, n16248, n16249, n16250, n16251,
    n16252, n16253, n16254, n16255, n16256, n16257,
    n16258, n16259, n16260, n16261, n16262, n16263,
    n16264, n16265, n16266, n16267, n16268, n16269,
    n16270, n16271, n16272, n16273, n16274, n16275,
    n16276, n16277, n16278, n16279, n16280, n16281,
    n16282, n16283, n16284, n16285, n16286, n16287,
    n16288, n16289, n16290, n16291, n16292, n16293,
    n16294, n16295, n16296, n16297, n16298, n16299,
    n16300, n16301, n16302, n16303, n16304, n16305,
    n16306, n16307, n16308, n16309, n16310, n16311,
    n16312, n16313, n16314, n16315, n16316, n16317,
    n16318, n16319, n16320, n16321, n16322, n16323,
    n16324, n16325, n16326, n16327, n16328, n16329,
    n16330, n16331, n16332, n16333, n16334, n16335,
    n16336, n16337, n16338, n16339, n16340, n16341,
    n16342, n16343, n16344, n16345, n16346, n16347,
    n16348, n16349, n16350, n16351, n16352, n16353,
    n16354, n16355, n16356, n16357, n16358, n16359,
    n16360, n16361, n16362, n16363, n16364, n16365,
    n16366, n16367, n16368, n16369, n16370, n16371,
    n16372, n16373, n16374, n16375, n16376, n16377,
    n16378, n16379, n16380, n16381, n16382, n16383,
    n16384, n16385, n16386, n16387, n16388, n16389,
    n16390, n16391, n16392, n16393, n16394, n16395,
    n16396, n16397, n16398, n16399, n16400, n16401,
    n16402, n16403, n16404, n16405, n16406, n16407,
    n16408, n16409, n16410, n16411, n16412, n16413,
    n16414, n16415, n16416, n16417, n16418, n16419,
    n16420, n16421, n16422, n16423, n16424, n16425,
    n16426, n16427, n16428, n16429, n16430, n16431,
    n16432, n16433, n16434, n16435, n16436, n16437,
    n16438, n16439, n16440, n16441, n16442, n16443,
    n16444, n16445, n16446, n16447, n16448, n16449,
    n16450, n16451, n16452, n16453, n16454, n16455,
    n16456, n16457, n16458, n16459, n16460, n16461,
    n16462, n16463, n16464, n16465, n16466, n16467,
    n16468, n16469, n16470, n16471, n16472, n16473,
    n16474, n16475, n16476, n16477, n16478, n16479,
    n16480, n16481, n16482, n16483, n16484, n16485,
    n16486, n16487, n16488, n16489, n16490, n16491,
    n16492, n16493, n16494, n16495, n16496, n16497,
    n16498, n16499, n16500, n16501, n16502, n16503,
    n16504, n16505, n16506, n16507, n16508, n16509,
    n16510, n16511, n16512, n16513, n16514, n16515,
    n16516, n16517, n16518, n16519, n16520, n16521,
    n16522, n16523, n16524, n16525, n16526, n16527,
    n16528, n16529, n16530, n16531, n16532, n16533,
    n16534, n16535, n16536, n16537, n16538, n16539,
    n16540, n16541, n16542, n16543, n16544, n16545,
    n16546, n16547, n16548, n16549, n16550, n16551,
    n16552, n16553, n16554, n16555, n16556, n16557,
    n16558, n16559, n16560, n16561, n16562, n16563,
    n16564, n16565, n16566, n16567, n16568, n16569,
    n16570, n16571, n16572, n16573, n16574, n16575,
    n16576, n16577, n16578, n16579, n16580, n16581,
    n16582, n16583, n16584, n16585, n16586, n16587,
    n16588, n16589, n16590, n16591, n16592, n16593,
    n16594, n16595, n16596, n16597, n16598, n16599,
    n16600, n16601, n16602, n16603, n16604, n16605,
    n16606, n16607, n16608, n16609, n16610, n16611,
    n16612, n16613, n16614, n16615, n16616, n16617,
    n16618, n16619, n16620, n16621, n16622, n16623,
    n16624, n16625, n16626, n16627, n16628, n16629,
    n16630, n16631, n16632, n16633, n16634, n16635,
    n16636, n16637, n16638, n16639, n16640, n16641,
    n16642, n16643, n16644, n16645, n16646, n16647,
    n16648, n16649, n16650, n16651, n16652, n16653,
    n16654, n16655, n16656, n16657, n16658, n16659,
    n16660, n16661, n16662, n16663, n16664, n16665,
    n16666, n16667, n16668, n16669, n16670, n16671,
    n16672, n16673, n16674, n16675, n16676, n16677,
    n16678, n16679, n16680, n16681, n16682, n16683,
    n16684, n16685, n16686, n16687, n16688, n16689,
    n16690, n16691, n16692, n16693, n16694, n16695,
    n16696, n16697, n16698, n16699, n16700, n16701,
    n16702, n16703, n16704, n16705, n16706, n16707,
    n16708, n16709, n16710, n16711, n16712, n16713,
    n16714, n16715, n16716, n16717, n16718, n16719,
    n16720, n16721, n16722, n16723, n16724, n16725,
    n16726, n16727, n16728, n16729, n16730, n16731,
    n16732, n16733, n16734, n16735, n16736, n16737,
    n16738, n16739, n16740, n16741, n16742, n16743,
    n16744, n16745, n16746, n16747, n16748, n16749,
    n16750, n16751, n16752, n16753, n16754, n16755,
    n16756, n16757, n16758, n16759, n16760, n16761,
    n16762, n16763, n16764, n16765, n16766, n16767,
    n16768, n16769, n16770, n16771, n16772, n16773,
    n16774, n16775, n16776, n16777, n16778, n16779,
    n16780, n16781, n16782, n16783, n16784, n16785,
    n16786, n16787, n16788, n16789, n16790, n16791,
    n16792, n16793, n16794, n16795, n16796, n16797,
    n16798, n16799, n16800, n16801, n16802, n16803,
    n16804, n16805, n16806, n16807, n16808, n16809,
    n16810, n16811, n16812, n16813, n16814, n16815,
    n16816, n16817, n16818, n16819, n16820, n16821,
    n16822, n16823, n16824, n16825, n16826, n16827,
    n16828, n16829, n16830, n16831, n16832, n16833,
    n16834, n16835, n16836, n16837, n16838, n16839,
    n16840, n16841, n16842, n16843, n16844, n16845,
    n16846, n16847, n16848, n16849, n16850, n16851,
    n16852, n16853, n16854, n16855, n16856, n16857,
    n16858, n16859, n16860, n16861, n16862, n16863,
    n16864, n16865, n16866, n16867, n16868, n16869,
    n16870, n16871, n16872, n16873, n16874, n16875,
    n16876, n16877, n16878, n16879, n16880, n16881,
    n16882, n16883, n16884, n16885, n16886, n16887,
    n16888, n16889, n16890, n16891, n16892, n16893,
    n16894, n16895, n16896, n16897, n16898, n16899,
    n16900, n16901, n16902, n16903, n16904, n16905,
    n16906, n16907, n16908, n16909, n16910, n16911,
    n16912, n16913, n16914, n16915, n16916, n16917,
    n16918, n16919, n16920, n16921, n16922, n16923,
    n16924, n16925, n16926, n16927, n16928, n16929,
    n16930, n16931, n16932, n16933, n16934, n16935,
    n16936, n16937, n16938, n16939, n16940, n16941,
    n16942, n16943, n16944, n16945, n16946, n16947,
    n16948, n16949, n16950, n16951, n16952, n16953,
    n16954, n16955, n16956, n16957, n16958, n16959,
    n16960, n16961, n16962, n16963, n16964, n16965,
    n16966, n16967, n16968, n16969, n16970, n16971,
    n16972, n16973, n16974, n16975, n16976, n16977,
    n16978, n16979, n16980, n16981, n16982, n16983,
    n16984, n16985, n16986, n16987, n16988, n16989,
    n16990, n16991, n16992, n16993, n16994, n16995,
    n16996, n16997, n16998, n16999, n17000, n17001,
    n17002, n17003, n17004, n17005, n17006, n17007,
    n17008, n17009, n17010, n17011, n17012, n17013,
    n17014, n17015, n17016, n17017, n17018, n17019,
    n17020, n17021, n17022, n17023, n17024, n17025,
    n17026, n17027, n17028, n17029, n17030, n17031,
    n17032, n17033, n17034, n17035, n17036, n17037,
    n17038, n17039, n17040, n17041, n17042, n17043,
    n17044, n17045, n17046, n17047, n17048, n17049,
    n17050, n17051, n17052, n17053, n17054, n17055,
    n17056, n17057, n17058, n17059, n17060, n17061,
    n17062, n17063, n17064, n17065, n17066, n17067,
    n17068, n17069, n17070, n17071, n17072, n17073,
    n17074, n17075, n17076, n17077, n17078, n17079,
    n17080, n17081, n17082, n17083, n17084, n17085,
    n17086, n17087, n17088, n17089, n17090, n17091,
    n17092, n17093, n17094, n17095, n17096, n17097,
    n17098, n17099, n17100, n17101, n17102, n17103,
    n17104, n17105, n17106, n17107, n17108, n17109,
    n17110, n17111, n17112, n17113, n17114, n17115,
    n17116, n17117, n17118, n17119, n17120, n17121,
    n17122, n17123, n17124, n17125, n17126, n17127,
    n17128, n17129, n17130, n17131, n17132, n17133,
    n17134, n17135, n17136, n17137, n17138, n17139,
    n17140, n17141, n17142, n17143, n17144, n17145,
    n17146, n17147, n17148, n17149, n17150, n17151,
    n17152, n17153, n17154, n17155, n17156, n17157,
    n17158, n17159, n17160, n17161, n17162, n17163,
    n17164, n17165, n17166, n17167, n17168, n17169,
    n17170, n17171, n17172, n17173, n17174, n17175,
    n17176, n17177, n17178, n17179, n17180, n17181,
    n17182, n17183, n17184, n17185, n17186, n17187,
    n17188, n17189, n17190, n17191, n17192, n17193,
    n17194, n17195, n17196, n17197, n17198, n17199,
    n17200, n17201, n17202, n17203, n17204, n17205,
    n17206, n17207, n17208, n17209, n17210, n17211,
    n17212, n17213, n17214, n17215, n17216, n17217,
    n17218, n17219, n17220, n17221, n17222, n17223,
    n17224, n17225, n17226, n17227, n17228, n17229,
    n17230, n17231, n17232, n17233, n17234, n17235,
    n17236, n17237, n17238, n17239, n17240, n17241,
    n17242, n17243, n17244, n17245, n17246, n17247,
    n17248, n17249, n17250, n17251, n17252, n17253,
    n17254, n17255, n17256, n17257, n17258, n17259,
    n17260, n17261, n17262, n17263, n17264, n17265,
    n17266, n17267, n17268, n17269, n17270, n17271,
    n17272, n17273, n17274, n17275, n17276, n17277,
    n17278, n17279, n17280, n17281, n17282, n17283,
    n17284, n17285, n17286, n17287, n17288, n17289,
    n17290, n17291, n17292, n17293, n17294, n17295,
    n17296, n17297, n17298, n17299, n17300, n17301,
    n17302, n17303, n17304, n17305, n17306, n17307,
    n17308, n17309, n17310, n17311, n17312, n17313,
    n17314, n17315, n17316, n17317, n17318, n17319,
    n17320, n17321, n17322, n17323, n17324, n17325,
    n17326, n17327, n17328, n17329, n17330, n17331,
    n17332, n17333, n17334, n17335, n17336, n17337,
    n17338, n17339, n17340, n17341, n17342, n17343,
    n17344, n17345, n17346, n17347, n17348, n17349,
    n17350, n17351, n17352, n17353, n17354, n17355,
    n17356, n17357, n17358, n17359, n17360, n17361,
    n17362, n17363, n17364, n17365, n17366, n17367,
    n17368, n17369, n17370, n17371, n17372, n17373,
    n17374, n17375, n17376, n17377, n17378, n17379,
    n17380, n17381, n17382, n17383, n17384, n17385,
    n17386, n17387, n17388, n17389, n17390, n17391,
    n17392, n17393, n17394, n17395, n17396, n17397,
    n17398, n17399, n17400, n17401, n17402, n17403,
    n17404, n17405, n17406, n17407, n17408, n17409,
    n17410, n17411, n17412, n17413, n17414, n17415,
    n17416, n17417, n17418, n17419, n17420, n17421,
    n17422, n17423, n17424, n17425, n17426, n17427,
    n17428, n17429, n17430, n17431, n17432, n17433,
    n17434, n17435, n17436, n17437, n17438, n17439,
    n17440, n17441, n17442, n17443, n17444, n17445,
    n17446, n17447, n17448, n17449, n17450, n17451,
    n17452, n17453, n17454, n17455, n17456, n17457,
    n17458, n17459, n17460, n17461, n17462, n17463,
    n17464, n17465, n17466, n17467, n17468, n17469,
    n17470, n17471, n17472, n17473, n17474, n17475,
    n17476, n17477, n17478, n17479, n17480, n17481,
    n17482, n17483, n17484, n17485, n17486, n17487,
    n17488, n17489, n17490, n17491, n17492, n17493,
    n17494, n17495, n17496, n17497, n17498, n17499,
    n17500, n17501, n17502, n17503, n17504, n17505,
    n17507, n17508, n17509, n17510, n17511, n17512,
    n17513, n17514, n17515, n17516, n17517, n17518,
    n17519, n17520, n17521, n17522, n17523, n17524,
    n17525, n17526, n17527, n17528, n17529, n17530,
    n17531, n17532, n17533, n17534, n17535, n17536,
    n17537, n17538, n17539, n17540, n17541, n17542,
    n17543, n17544, n17545, n17546, n17547, n17548,
    n17549, n17550, n17551, n17552, n17553, n17554,
    n17555, n17556, n17557, n17558, n17559, n17560,
    n17561, n17562, n17563, n17564, n17565, n17566,
    n17567, n17568, n17569, n17570, n17571, n17572,
    n17573, n17574, n17575, n17576, n17577, n17578,
    n17579, n17580, n17581, n17582, n17583, n17584,
    n17585, n17586, n17587, n17588, n17589, n17590,
    n17591, n17592, n17593, n17594, n17595, n17596,
    n17597, n17598, n17599, n17600, n17601, n17602,
    n17603, n17604, n17605, n17606, n17607, n17608,
    n17609, n17610, n17611, n17612, n17613, n17614,
    n17615, n17616, n17617, n17618, n17619, n17620,
    n17621, n17622, n17623, n17624, n17625, n17626,
    n17627, n17628, n17629, n17630, n17631, n17632,
    n17633, n17634, n17635, n17636, n17637, n17638,
    n17639, n17640, n17641, n17642, n17643, n17644,
    n17645, n17646, n17647, n17648, n17649, n17650,
    n17651, n17652, n17653, n17654, n17655, n17656,
    n17657, n17658, n17659, n17660, n17661, n17662,
    n17663, n17664, n17665, n17666, n17667, n17668,
    n17669, n17670, n17671, n17672, n17673, n17674,
    n17675, n17676, n17677, n17678, n17679, n17680,
    n17681, n17682, n17683, n17684, n17685, n17686,
    n17687, n17688, n17689, n17690, n17691, n17692,
    n17693, n17694, n17695, n17696, n17697, n17698,
    n17699, n17700, n17701, n17702, n17703, n17704,
    n17705, n17706, n17707, n17708, n17709, n17710,
    n17711, n17712, n17713, n17714, n17715, n17716,
    n17717, n17718, n17719, n17720, n17721, n17722,
    n17723, n17724, n17725, n17726, n17727, n17728,
    n17729, n17730, n17731, n17732, n17733, n17734,
    n17735, n17736, n17737, n17738, n17739, n17740,
    n17741, n17742, n17743, n17744, n17745, n17746,
    n17747, n17748, n17749, n17750, n17751, n17752,
    n17753, n17754, n17755, n17756, n17757, n17758,
    n17759, n17760, n17761, n17762, n17763, n17764,
    n17765, n17766, n17767, n17768, n17769, n17770,
    n17771, n17772, n17773, n17774, n17775, n17776,
    n17777, n17778, n17779, n17780, n17781, n17782,
    n17783, n17784, n17785, n17786, n17787, n17788,
    n17789, n17790, n17791, n17792, n17793, n17794,
    n17795, n17796, n17797, n17798, n17799, n17800,
    n17801, n17802, n17803, n17804, n17805, n17806,
    n17807, n17808, n17809, n17810, n17811, n17812,
    n17813, n17814, n17815, n17816, n17817, n17818,
    n17819, n17820, n17821, n17822, n17823, n17824,
    n17825, n17826, n17827, n17828, n17829, n17830,
    n17831, n17832, n17833, n17834, n17835, n17836,
    n17837, n17838, n17839, n17840, n17841, n17842,
    n17843, n17844, n17845, n17846, n17847, n17848,
    n17849, n17850, n17851, n17852, n17853, n17854,
    n17855, n17856, n17857, n17858, n17859, n17860,
    n17861, n17862, n17863, n17864, n17865, n17866,
    n17867, n17868, n17869, n17870, n17871, n17872,
    n17873, n17874, n17875, n17876, n17877, n17878,
    n17879, n17880, n17881, n17882, n17883, n17884,
    n17885, n17886, n17887, n17888, n17889, n17890,
    n17891, n17892, n17893, n17894, n17895, n17896,
    n17897, n17898, n17899, n17900, n17901, n17902,
    n17903, n17904, n17905, n17906, n17907, n17908,
    n17909, n17910, n17911, n17912, n17913, n17914,
    n17915, n17916, n17917, n17918, n17919, n17920,
    n17921, n17922, n17923, n17924, n17925, n17926,
    n17927, n17928, n17929, n17930, n17931, n17932,
    n17933, n17934, n17935, n17936, n17937, n17938,
    n17939, n17940, n17941, n17942, n17943, n17944,
    n17945, n17946, n17947, n17948, n17949, n17950,
    n17951, n17952, n17953, n17954, n17955, n17956,
    n17957, n17958, n17959, n17960, n17961, n17962,
    n17963, n17964, n17965, n17966, n17967, n17968,
    n17969, n17970, n17971, n17972, n17973, n17974,
    n17975, n17976, n17977, n17978, n17979, n17980,
    n17981, n17982, n17983, n17984, n17985, n17986,
    n17987, n17988, n17989, n17990, n17991, n17992,
    n17993, n17994, n17995, n17996, n17997, n17998,
    n17999, n18000, n18001, n18002, n18003, n18004,
    n18005, n18006, n18007, n18008, n18009, n18010,
    n18011, n18012, n18013, n18014, n18015, n18016,
    n18017, n18018, n18019, n18020, n18021, n18022,
    n18023, n18024, n18025, n18026, n18027, n18028,
    n18029, n18030, n18032, n18033, n18034, n18035,
    n18036, n18037, n18038, n18039, n18040, n18041,
    n18042, n18043, n18044, n18045, n18046, n18047,
    n18048, n18049, n18050, n18051, n18052, n18053,
    n18054, n18055, n18056, n18057, n18058, n18059,
    n18060, n18061, n18062, n18063, n18064, n18065,
    n18066, n18067, n18068, n18069, n18070, n18071,
    n18072, n18073, n18074, n18075, n18076, n18077,
    n18078, n18079, n18080, n18081, n18082, n18083,
    n18084, n18085, n18086, n18087, n18088, n18089,
    n18090, n18091, n18092, n18093, n18094, n18095,
    n18096, n18097, n18098, n18099, n18100, n18101,
    n18102, n18103, n18104, n18105, n18106, n18107,
    n18108, n18109, n18110, n18111, n18112, n18113,
    n18114, n18115, n18116, n18117, n18118, n18119,
    n18120, n18121, n18122, n18123, n18124, n18125,
    n18126, n18127, n18128, n18129, n18130, n18131,
    n18132, n18133, n18134, n18135, n18136, n18137,
    n18138, n18139, n18140, n18141, n18142, n18143,
    n18144, n18145, n18146, n18147, n18148, n18149,
    n18150, n18151, n18152, n18153, n18154, n18155,
    n18156, n18157, n18158, n18159, n18160, n18161,
    n18162, n18163, n18164, n18165, n18166, n18167,
    n18168, n18169, n18170, n18171, n18172, n18173,
    n18174, n18175, n18176, n18177, n18178, n18179,
    n18180, n18181, n18182, n18183, n18184, n18185,
    n18186, n18187, n18188, n18189, n18190, n18191,
    n18192, n18193, n18194, n18195, n18196, n18197,
    n18198, n18199, n18200, n18201, n18202, n18203,
    n18204, n18205, n18206, n18207, n18208, n18209,
    n18210, n18211, n18212, n18213, n18214, n18215,
    n18216, n18217, n18218, n18219, n18220, n18221,
    n18222, n18223, n18224, n18225, n18226, n18227,
    n18228, n18229, n18230, n18231, n18232, n18233,
    n18234, n18235, n18236, n18237, n18238, n18239,
    n18240, n18241, n18242, n18243, n18244, n18245,
    n18246, n18247, n18248, n18249, n18250, n18251,
    n18252, n18253, n18254, n18255, n18256, n18257,
    n18258, n18259, n18260, n18261, n18262, n18263,
    n18264, n18265, n18266, n18267, n18268, n18269,
    n18270, n18271, n18272, n18273, n18274, n18275,
    n18276, n18277, n18278, n18279, n18280, n18281,
    n18282, n18283, n18284, n18285, n18286, n18287,
    n18288, n18289, n18290, n18291, n18292, n18293,
    n18294, n18295, n18296, n18297, n18298, n18299,
    n18300, n18301, n18302, n18303, n18304, n18305,
    n18306, n18307, n18308, n18309, n18310, n18311,
    n18312, n18313, n18314, n18315, n18316, n18317,
    n18318, n18319, n18320, n18321, n18322, n18323,
    n18324, n18325, n18326, n18327, n18328, n18329,
    n18330, n18331, n18332, n18333, n18334, n18335,
    n18336, n18337, n18338, n18339, n18340, n18341,
    n18342, n18343, n18344, n18345, n18346, n18347,
    n18348, n18349, n18350, n18351, n18352, n18353,
    n18354, n18355, n18356, n18357, n18358, n18359,
    n18360, n18361, n18362, n18363, n18364, n18365,
    n18366, n18367, n18368, n18369, n18370, n18371,
    n18372, n18373, n18374, n18375, n18376, n18377,
    n18378, n18379, n18380, n18381, n18382, n18383,
    n18384, n18385, n18386, n18387, n18388, n18389,
    n18390, n18391, n18392, n18393, n18394, n18395,
    n18396, n18397, n18398, n18399, n18400, n18401,
    n18402, n18403, n18404, n18405, n18406, n18407,
    n18408, n18409, n18410, n18411, n18412, n18413,
    n18414, n18415, n18416, n18417, n18418, n18419,
    n18420, n18421, n18422, n18423, n18424, n18425,
    n18426, n18427, n18428, n18429, n18430, n18431,
    n18432, n18433, n18434, n18435, n18436, n18437,
    n18438, n18439, n18440, n18441, n18442, n18443,
    n18444, n18445, n18446, n18447, n18448, n18449,
    n18450, n18451, n18452, n18453, n18454, n18455,
    n18456, n18457, n18458, n18459, n18460, n18461,
    n18462, n18463, n18464, n18465, n18466, n18467,
    n18468, n18469, n18470, n18471, n18472, n18473,
    n18474, n18475, n18476, n18477, n18478, n18479,
    n18480, n18481, n18482, n18483, n18484, n18485,
    n18486, n18487, n18488, n18489, n18490, n18491,
    n18492, n18493, n18494, n18495, n18496, n18497,
    n18498, n18499, n18500, n18501, n18502, n18503,
    n18504, n18505, n18506, n18507, n18508, n18509,
    n18510, n18511, n18512, n18513, n18514, n18515,
    n18516, n18517, n18518, n18519, n18520, n18521,
    n18522, n18523, n18524, n18525, n18526, n18527,
    n18528, n18529, n18530, n18531, n18532, n18533,
    n18534, n18535, n18536, n18537, n18538, n18539,
    n18540, n18541, n18542, n18543, n18544, n18545,
    n18546, n18547, n18548, n18549, n18550, n18551,
    n18552, n18553, n18554, n18555, n18556, n18557,
    n18558, n18559, n18560, n18561, n18562, n18563,
    n18564, n18565, n18566, n18567, n18568, n18569,
    n18570, n18571, n18572, n18573, n18574, n18575,
    n18576, n18577, n18578, n18579, n18580, n18581,
    n18582, n18583, n18584, n18585, n18586, n18587,
    n18588, n18589, n18590, n18591, n18592, n18593,
    n18594, n18595, n18596, n18597, n18598, n18599,
    n18600, n18601, n18602, n18603, n18604, n18605,
    n18606, n18607, n18608, n18609, n18610, n18611,
    n18612, n18613, n18614, n18615, n18616, n18617,
    n18618, n18619, n18620, n18621, n18622, n18623,
    n18624, n18625, n18626, n18627, n18628, n18629,
    n18630, n18631, n18632, n18633, n18634, n18635,
    n18636, n18637, n18638, n18639, n18640, n18641,
    n18642, n18643, n18644, n18645, n18646, n18647,
    n18648, n18649, n18650, n18651, n18652, n18653,
    n18654, n18655, n18656, n18657, n18658, n18659,
    n18660, n18661, n18662, n18663, n18664, n18665,
    n18666, n18667, n18668, n18669, n18670, n18671,
    n18672, n18673, n18674, n18675, n18676, n18677,
    n18678, n18679, n18680, n18681, n18682, n18683,
    n18684, n18685, n18686, n18687, n18688, n18689,
    n18690, n18691, n18692, n18693, n18694, n18695,
    n18696, n18697, n18698, n18699, n18700, n18701,
    n18702, n18703, n18704, n18705, n18706, n18707,
    n18708, n18709, n18710, n18711, n18712, n18713,
    n18714, n18715, n18716, n18717, n18718, n18719,
    n18720, n18721, n18722, n18723, n18724, n18725,
    n18726, n18727, n18728, n18729, n18730, n18731,
    n18732, n18733, n18734, n18735, n18736, n18737,
    n18738, n18739, n18740, n18741, n18742, n18743,
    n18744, n18745, n18746, n18747, n18748, n18749,
    n18750, n18751, n18752, n18753, n18754, n18755,
    n18756, n18757, n18758, n18759, n18760, n18761,
    n18762, n18763, n18764, n18765, n18766, n18767,
    n18768, n18769, n18770, n18771, n18772, n18773,
    n18774, n18775, n18776, n18777, n18778, n18779,
    n18780, n18781, n18782, n18783, n18784, n18785,
    n18786, n18787, n18788, n18789, n18790, n18791,
    n18792, n18793, n18794, n18795, n18796, n18798,
    n18799, n18800, n18801, n18802, n18803, n18804,
    n18805, n18806, n18807, n18808, n18809, n18810,
    n18811, n18812, n18813, n18814, n18815, n18816,
    n18817, n18818, n18819, n18820, n18821, n18822,
    n18823, n18824, n18825, n18826, n18827, n18828,
    n18829, n18830, n18831, n18832, n18833, n18834,
    n18835, n18836, n18837, n18838, n18839, n18840,
    n18841, n18842, n18843, n18844, n18845, n18846,
    n18847, n18848, n18849, n18850, n18851, n18852,
    n18853, n18854, n18855, n18856, n18857, n18858,
    n18859, n18860, n18861, n18862, n18863, n18864,
    n18865, n18866, n18867, n18868, n18869, n18870,
    n18871, n18872, n18873, n18874, n18875, n18876,
    n18877, n18878, n18879, n18880, n18881, n18882,
    n18883, n18884, n18885, n18886, n18887, n18888,
    n18889, n18890, n18891, n18892, n18893, n18894,
    n18895, n18896, n18897, n18898, n18899, n18900,
    n18901, n18902, n18903, n18904, n18905, n18906,
    n18907, n18908, n18909, n18910, n18911, n18912,
    n18913, n18914, n18915, n18916, n18917, n18918,
    n18919, n18920, n18921, n18922, n18923, n18924,
    n18925, n18926, n18927, n18928, n18929, n18930,
    n18931, n18932, n18933, n18934, n18935, n18936,
    n18937, n18938, n18939, n18940, n18941, n18942,
    n18943, n18944, n18945, n18946, n18947, n18948,
    n18949, n18950, n18951, n18952, n18953, n18954,
    n18955, n18956, n18957, n18958, n18959, n18960,
    n18961, n18962, n18963, n18964, n18965, n18966,
    n18967, n18968, n18969, n18970, n18971, n18972,
    n18973, n18974, n18975, n18976, n18977, n18978,
    n18979, n18980, n18981, n18982, n18983, n18984,
    n18985, n18986, n18987, n18988, n18989, n18990,
    n18991, n18992, n18993, n18994, n18995, n18996,
    n18997, n18998, n18999, n19000, n19001, n19002,
    n19003, n19004, n19005, n19006, n19007, n19008,
    n19009, n19010, n19011, n19012, n19013, n19014,
    n19015, n19016, n19017, n19018, n19019, n19020,
    n19021, n19022, n19023, n19024, n19025, n19026,
    n19027, n19028, n19029, n19030, n19031, n19032,
    n19033, n19034, n19035, n19036, n19037, n19038,
    n19039, n19040, n19041, n19042, n19043, n19044,
    n19045, n19046, n19047, n19048, n19049, n19050,
    n19051, n19052, n19053, n19054, n19055, n19056,
    n19057, n19058, n19059, n19060, n19061, n19062,
    n19063, n19064, n19065, n19066, n19067, n19068,
    n19069, n19070, n19071, n19072, n19073, n19074,
    n19075, n19076, n19077, n19078, n19079, n19080,
    n19081, n19082, n19083, n19084, n19085, n19086,
    n19087, n19088, n19089, n19090, n19091, n19092,
    n19093, n19094, n19095, n19096, n19097, n19098,
    n19099, n19100, n19101, n19102, n19103, n19104,
    n19105, n19106, n19107, n19108, n19109, n19110,
    n19111, n19112, n19113, n19114, n19115, n19116,
    n19117, n19118, n19119, n19120, n19121, n19122,
    n19123, n19124, n19125, n19126, n19127, n19128,
    n19129, n19130, n19131, n19132, n19133, n19134,
    n19135, n19136, n19137, n19138, n19139, n19140,
    n19141, n19142, n19143, n19144, n19145, n19146,
    n19147, n19148, n19149, n19150, n19151, n19152,
    n19153, n19154, n19155, n19156, n19157, n19158,
    n19159, n19160, n19161, n19162, n19163, n19164,
    n19165, n19166, n19167, n19168, n19169, n19170,
    n19171, n19172, n19173, n19174, n19175, n19176,
    n19177, n19178, n19179, n19180, n19181, n19182,
    n19183, n19184, n19185, n19186, n19187, n19188,
    n19189, n19190, n19191, n19192, n19193, n19194,
    n19195, n19196, n19197, n19198, n19199, n19200,
    n19201, n19202, n19203, n19204, n19205, n19206,
    n19207, n19208, n19209, n19210, n19211, n19212,
    n19213, n19214, n19215, n19216, n19217, n19218,
    n19219, n19220, n19221, n19222, n19223, n19224,
    n19225, n19226, n19227, n19228, n19229, n19230,
    n19231, n19232, n19233, n19234, n19235, n19236,
    n19237, n19238, n19239, n19240, n19241, n19242,
    n19243, n19244, n19245, n19246, n19247, n19248,
    n19249, n19250, n19251, n19252, n19253, n19254,
    n19255, n19256, n19257, n19258, n19259, n19260,
    n19261, n19262, n19263, n19264, n19265, n19266,
    n19267, n19268, n19269, n19270, n19271, n19272,
    n19273, n19274, n19275, n19276, n19277, n19278,
    n19279, n19280, n19281, n19282, n19283, n19284,
    n19285, n19286, n19287, n19288, n19289, n19290,
    n19291, n19292, n19293, n19294, n19295, n19296,
    n19297, n19298, n19299, n19300, n19301, n19302,
    n19303, n19304, n19305, n19306, n19307, n19308,
    n19309, n19310, n19311, n19312, n19313, n19314,
    n19315, n19316, n19317, n19318, n19319, n19320,
    n19321, n19322, n19323, n19325, n19326, n19327,
    n19328, n19329, n19330, n19331, n19332, n19333,
    n19334, n19335, n19336, n19337, n19338, n19339,
    n19340, n19341, n19342, n19343, n19344, n19345,
    n19346, n19347, n19348, n19349, n19350, n19351,
    n19352, n19353, n19354, n19355, n19356, n19357,
    n19358, n19359, n19360, n19361, n19362, n19363,
    n19364, n19365, n19366, n19367, n19368, n19369,
    n19370, n19371, n19372, n19373, n19374, n19375,
    n19376, n19377, n19378, n19379, n19380, n19381,
    n19382, n19383, n19384, n19385, n19386, n19387,
    n19388, n19389, n19390, n19391, n19392, n19393,
    n19394, n19395, n19396, n19397, n19398, n19399,
    n19400, n19401, n19402, n19403, n19404, n19405,
    n19406, n19407, n19408, n19409, n19410, n19411,
    n19412, n19413, n19414, n19415, n19416, n19417,
    n19418, n19419, n19420, n19421, n19422, n19423,
    n19424, n19425, n19426, n19427, n19428, n19429,
    n19430, n19431, n19432, n19433, n19434, n19435,
    n19436, n19437, n19438, n19439, n19440, n19441,
    n19442, n19443, n19444, n19445, n19446, n19447,
    n19448, n19449, n19450, n19451, n19452, n19453,
    n19454, n19455, n19456, n19457, n19458, n19459,
    n19460, n19461, n19462, n19463, n19464, n19465,
    n19466, n19467, n19468, n19469, n19470, n19471,
    n19472, n19473, n19474, n19475, n19476, n19477,
    n19478, n19479, n19480, n19481, n19482, n19483,
    n19484, n19485, n19486, n19487, n19488, n19489,
    n19490, n19491, n19492, n19493, n19494, n19495,
    n19496, n19497, n19498, n19499, n19500, n19501,
    n19502, n19503, n19504, n19505, n19506, n19507,
    n19508, n19509, n19510, n19511, n19512, n19513,
    n19514, n19515, n19516, n19517, n19518, n19519,
    n19520, n19521, n19522, n19523, n19524, n19525,
    n19526, n19527, n19528, n19529, n19530, n19531,
    n19532, n19533, n19534, n19535, n19536, n19537,
    n19538, n19539, n19540, n19541, n19542, n19543,
    n19544, n19545, n19546, n19547, n19548, n19549,
    n19550, n19551, n19552, n19553, n19554, n19555,
    n19556, n19557, n19558, n19559, n19560, n19561,
    n19562, n19563, n19564, n19565, n19566, n19567,
    n19568, n19569, n19570, n19571, n19572, n19573,
    n19574, n19575, n19576, n19577, n19578, n19579,
    n19580, n19581, n19582, n19583, n19584, n19585,
    n19586, n19587, n19588, n19589, n19590, n19591,
    n19592, n19593, n19594, n19595, n19596, n19597,
    n19598, n19599, n19600, n19601, n19602, n19603,
    n19604, n19605, n19606, n19607, n19608, n19609,
    n19610, n19611, n19612, n19613, n19614, n19615,
    n19616, n19617, n19618, n19619, n19620, n19621,
    n19622, n19623, n19624, n19625, n19626, n19627,
    n19628, n19629, n19630, n19631, n19632, n19633,
    n19634, n19635, n19636, n19637, n19638, n19639,
    n19640, n19641, n19642, n19643, n19644, n19645,
    n19646, n19647, n19648, n19649, n19650, n19651,
    n19652, n19653, n19654, n19655, n19656, n19657,
    n19658, n19659, n19660, n19661, n19662, n19663,
    n19664, n19665, n19666, n19667, n19668, n19669,
    n19670, n19671, n19672, n19673, n19674, n19675,
    n19676, n19677, n19678, n19679, n19680, n19681,
    n19682, n19683, n19684, n19685, n19686, n19687,
    n19688, n19689, n19690, n19691, n19692, n19693,
    n19694, n19695, n19696, n19697, n19698, n19699,
    n19700, n19701, n19702, n19703, n19704, n19705,
    n19706, n19707, n19708, n19709, n19710, n19711,
    n19712, n19713, n19714, n19715, n19716, n19717,
    n19718, n19719, n19720, n19721, n19722, n19723,
    n19724, n19725, n19726, n19727, n19728, n19729,
    n19730, n19731, n19732, n19733, n19734, n19735,
    n19736, n19737, n19738, n19739, n19740, n19741,
    n19742, n19743, n19744, n19745, n19746, n19747,
    n19748, n19749, n19750, n19751, n19752, n19753,
    n19754, n19755, n19756, n19757, n19758, n19759,
    n19760, n19761, n19762, n19763, n19764, n19765,
    n19766, n19767, n19768, n19769, n19770, n19771,
    n19772, n19773, n19774, n19775, n19776, n19777,
    n19778, n19779, n19780, n19781, n19782, n19783,
    n19784, n19785, n19786, n19787, n19788, n19789,
    n19790, n19791, n19792, n19793, n19794, n19795,
    n19796, n19797, n19798, n19799, n19800, n19801,
    n19802, n19803, n19804, n19805, n19806, n19807,
    n19808, n19809, n19810, n19811, n19812, n19813,
    n19814, n19815, n19816, n19817, n19818, n19819,
    n19820, n19821, n19822, n19823, n19824, n19825,
    n19826, n19827, n19828, n19829, n19830, n19831,
    n19832, n19833, n19834, n19836, n19837, n19838,
    n19839, n19840, n19841, n19842, n19843, n19844,
    n19845, n19846, n19847, n19848, n19849, n19850,
    n19851, n19852, n19853, n19854, n19855, n19856,
    n19857, n19858, n19859, n19860, n19861, n19862,
    n19863, n19864, n19865, n19866, n19867, n19868,
    n19869, n19870, n19871, n19872, n19873, n19874,
    n19875, n19876, n19877, n19878, n19879, n19880,
    n19881, n19882, n19883, n19884, n19885, n19886,
    n19887, n19888, n19889, n19890, n19891, n19892,
    n19893, n19894, n19895, n19896, n19897, n19898,
    n19899, n19900, n19901, n19902, n19903, n19904,
    n19905, n19906, n19907, n19908, n19909, n19910,
    n19911, n19912, n19913, n19914, n19915, n19916,
    n19917, n19918, n19919, n19920, n19921, n19922,
    n19923, n19924, n19925, n19926, n19927, n19928,
    n19929, n19930, n19931, n19932, n19933, n19934,
    n19935, n19936, n19937, n19938, n19939, n19940,
    n19941, n19942, n19943, n19944, n19945, n19946,
    n19947, n19948, n19949, n19950, n19951, n19952,
    n19953, n19954, n19955, n19956, n19957, n19958,
    n19959, n19960, n19961, n19962, n19963, n19964,
    n19965, n19966, n19967, n19968, n19969, n19970,
    n19971, n19972, n19973, n19974, n19975, n19976,
    n19977, n19978, n19979, n19980, n19981, n19982,
    n19983, n19984, n19985, n19986, n19987, n19988,
    n19989, n19990, n19991, n19992, n19993, n19994,
    n19995, n19996, n19997, n19998, n19999, n20000,
    n20001, n20002, n20003, n20004, n20005, n20006,
    n20007, n20008, n20009, n20010, n20011, n20012,
    n20013, n20014, n20015, n20016, n20017, n20018,
    n20019, n20020, n20021, n20022, n20023, n20024,
    n20025, n20026, n20027, n20028, n20029, n20030,
    n20031, n20032, n20033, n20034, n20035, n20036,
    n20037, n20038, n20039, n20040, n20041, n20042,
    n20043, n20044, n20045, n20046, n20047, n20048,
    n20049, n20050, n20051, n20052, n20053, n20054,
    n20055, n20056, n20057, n20058, n20059, n20060,
    n20061, n20062, n20063, n20064, n20065, n20066,
    n20067, n20068, n20069, n20070, n20071, n20072,
    n20073, n20074, n20075, n20076, n20077, n20078,
    n20079, n20080, n20081, n20082, n20083, n20084,
    n20085, n20086, n20087, n20088, n20089, n20090,
    n20091, n20092, n20093, n20094, n20095, n20096,
    n20097, n20098, n20099, n20100, n20101, n20102,
    n20103, n20104, n20105, n20106, n20107, n20108,
    n20109, n20110, n20111, n20112, n20113, n20114,
    n20115, n20116, n20117, n20118, n20119, n20120,
    n20121, n20122, n20123, n20124, n20125, n20126,
    n20127, n20128, n20129, n20130, n20131, n20132,
    n20133, n20134, n20135, n20136, n20137, n20138,
    n20139, n20140, n20141, n20142, n20143, n20144,
    n20145, n20146, n20147, n20148, n20149, n20150,
    n20151, n20152, n20153, n20154, n20155, n20156,
    n20157, n20158, n20159, n20160, n20161, n20162,
    n20163, n20164, n20165, n20166, n20167, n20168,
    n20169, n20170, n20171, n20172, n20173, n20174,
    n20175, n20176, n20177, n20178, n20179, n20180,
    n20181, n20182, n20183, n20184, n20185, n20186,
    n20187, n20188, n20189, n20190, n20191, n20192,
    n20193, n20194, n20195, n20196, n20197, n20198,
    n20199, n20200, n20201, n20202, n20203, n20204,
    n20205, n20206, n20207, n20208, n20209, n20210,
    n20211, n20212, n20213, n20214, n20215, n20216,
    n20217, n20218, n20219, n20220, n20221, n20222,
    n20223, n20224, n20225, n20226, n20227, n20228,
    n20229, n20230, n20231, n20232, n20233, n20234,
    n20235, n20236, n20237, n20238, n20239, n20240,
    n20241, n20242, n20243, n20244, n20245, n20246,
    n20247, n20248, n20249, n20250, n20251, n20252,
    n20253, n20254, n20255, n20256, n20257, n20258,
    n20259, n20260, n20261, n20262, n20263, n20264,
    n20265, n20266, n20267, n20268, n20269, n20270,
    n20271, n20272, n20273, n20274, n20275, n20276,
    n20277, n20278, n20279, n20280, n20281, n20282,
    n20283, n20284, n20285, n20286, n20287, n20288,
    n20289, n20290, n20291, n20292, n20293, n20294,
    n20295, n20296, n20297, n20298, n20299, n20300,
    n20301, n20302, n20303, n20304, n20305, n20306,
    n20307, n20308, n20309, n20310, n20311, n20312,
    n20313, n20314, n20315, n20316, n20317, n20318,
    n20319, n20320, n20322, n20323, n20324, n20325,
    n20326, n20327, n20328, n20329, n20330, n20331,
    n20332, n20333, n20334, n20335, n20336, n20337,
    n20338, n20339, n20340, n20341, n20342, n20343,
    n20344, n20345, n20346, n20347, n20348, n20349,
    n20350, n20351, n20352, n20353, n20354, n20355,
    n20356, n20357, n20358, n20359, n20360, n20361,
    n20362, n20363, n20364, n20365, n20366, n20367,
    n20368, n20369, n20370, n20371, n20372, n20373,
    n20374, n20375, n20376, n20377, n20378, n20379,
    n20380, n20381, n20382, n20383, n20384, n20385,
    n20386, n20387, n20388, n20389, n20390, n20391,
    n20392, n20393, n20394, n20395, n20396, n20397,
    n20398, n20399, n20400, n20401, n20403, n20404,
    n20405, n20406, n20407, n20408, n20409, n20410,
    n20411, n20412, n20413, n20414, n20415, n20416,
    n20417, n20418, n20419, n20420, n20421, n20422,
    n20423, n20424, n20425, n20426, n20427, n20428,
    n20429, n20430, n20431, n20432, n20433, n20434,
    n20435, n20436, n20437, n20438, n20439, n20440,
    n20441, n20442, n20443, n20444, n20445, n20446,
    n20447, n20448, n20449, n20450, n20451, n20452,
    n20453, n20454, n20455, n20456, n20457, n20458,
    n20459, n20460, n20461, n20462, n20463, n20464,
    n20465, n20466, n20467, n20468, n20469, n20470,
    n20471, n20472, n20473, n20474, n20475, n20476,
    n20477, n20478, n20479, n20480, n20481, n20482,
    n20483, n20484, n20485, n20486, n20487, n20488,
    n20489, n20490, n20491, n20492, n20493, n20494,
    n20495, n20496, n20497, n20498, n20499, n20500,
    n20501, n20502, n20503, n20504, n20505, n20506,
    n20507, n20508, n20509, n20510, n20511, n20512,
    n20513, n20514, n20515, n20516, n20517, n20518,
    n20519, n20520, n20521, n20522, n20523, n20524,
    n20525, n20526, n20527, n20528, n20529, n20530,
    n20531, n20532, n20533, n20534, n20535, n20537,
    n20538, n20539, n20540, n20541, n20542, n20543,
    n20544, n20545, n20546, n20547, n20548, n20549,
    n20550, n20551, n20552, n20553, n20554, n20555,
    n20556, n20557, n20558, n20559, n20560, n20561,
    n20562, n20563, n20564, n20565, n20566, n20567,
    n20568, n20569, n20570, n20571, n20572, n20573,
    n20574, n20575, n20576, n20577, n20578, n20579,
    n20580, n20581, n20582, n20583, n20584, n20585,
    n20586, n20587, n20588, n20589, n20590, n20591,
    n20592, n20593, n20594, n20595, n20596, n20597,
    n20598, n20599, n20601, n20602, n20603, n20604,
    n20605, n20606, n20607, n20608, n20609, n20610,
    n20611, n20612, n20613, n20614, n20615, n20616,
    n20617, n20618, n20619, n20620, n20621, n20622,
    n20623, n20624, n20625, n20626, n20627, n20628,
    n20629, n20630, n20631, n20632, n20633, n20634,
    n20635, n20636, n20637, n20638, n20639, n20640,
    n20641, n20642, n20643, n20644, n20645, n20646,
    n20647, n20648, n20649, n20650, n20651, n20652,
    n20653, n20654, n20656, n20657, n20658, n20659,
    n20660, n20661, n20662, n20663, n20664, n20665,
    n20666, n20667, n20668, n20669, n20670, n20671,
    n20672, n20673, n20674, n20675, n20676, n20677,
    n20678, n20679, n20680, n20681, n20682, n20683,
    n20684, n20685, n20686, n20687, n20688, n20689,
    n20690, n20691, n20692, n20693, n20694, n20695,
    n20696, n20697, n20698, n20699, n20700, n20701,
    n20702, n20703, n20704, n20705, n20706, n20707,
    n20709, n20710, n20711, n20712, n20713, n20714,
    n20715, n20716, n20717, n20718, n20719, n20720,
    n20721, n20722, n20723, n20724, n20725, n20726,
    n20727, n20728, n20729, n20730, n20731, n20732,
    n20733, n20734, n20735, n20736, n20737, n20738,
    n20739, n20740, n20741, n20742, n20743, n20744,
    n20745, n20746, n20747, n20748, n20749, n20750,
    n20751, n20752, n20753, n20754, n20755, n20756,
    n20757, n20758, n20759, n20760, n20761, n20762,
    n20763, n20764, n20765, n20766, n20767, n20768,
    n20769, n20770, n20771, n20772, n20773, n20774,
    n20775, n20776, n20777, n20778, n20779, n20780,
    n20781, n20782, n20783, n20784, n20786, n20787,
    n20788, n20789, n20790, n20791, n20792, n20793,
    n20794, n20795, n20796, n20797, n20798, n20799,
    n20800, n20801, n20802, n20803, n20804, n20805,
    n20806, n20807, n20808, n20809, n20810, n20811,
    n20812, n20813, n20814, n20815, n20816, n20817,
    n20818, n20819, n20820, n20821, n20822, n20823,
    n20824, n20825, n20826, n20827, n20828, n20829,
    n20830, n20831, n20832, n20833, n20834, n20835,
    n20836, n20837, n20838, n20839, n20840, n20841,
    n20842, n20843, n20844, n20845, n20846, n20847,
    n20848, n20849, n20850, n20851, n20852, n20853,
    n20854, n20855, n20856, n20857, n20858, n20859,
    n20860, n20861, n20862, n20863, n20864, n20865,
    n20866, n20867, n20868, n20869, n20870, n20871,
    n20872, n20873, n20874, n20875, n20876, n20877,
    n20878, n20879, n20880, n20881, n20882, n20883,
    n20884, n20885, n20886, n20887, n20888, n20890,
    n20891, n20892, n20893, n20894, n20895, n20896,
    n20897, n20898, n20899, n20900, n20901, n20902,
    n20903, n20904, n20905, n20906, n20907, n20908,
    n20909, n20910, n20911, n20912, n20913, n20914,
    n20915, n20916, n20917, n20918, n20919, n20920,
    n20921, n20922, n20923, n20924, n20925, n20926,
    n20927, n20928, n20929, n20930, n20931, n20932,
    n20933, n20934, n20935, n20936, n20937, n20938,
    n20939, n20940, n20941, n20942, n20943, n20944,
    n20945, n20946, n20947, n20948, n20949, n20950,
    n20951, n20952, n20953, n20954, n20955, n20956,
    n20957, n20958, n20959, n20960, n20961, n20962,
    n20963, n20964, n20965, n20966, n20967, n20969,
    n20970, n20971, n20972, n20973, n20974, n20975,
    n20976, n20977, n20978, n20979, n20980, n20981,
    n20982, n20983, n20984, n20985, n20986, n20987,
    n20988, n20989, n20990, n20991, n20992, n20993,
    n20994, n20995, n20996, n20997, n20998, n20999,
    n21000, n21001, n21002, n21003, n21004, n21005,
    n21006, n21007, n21008, n21009, n21010, n21011,
    n21012, n21013, n21014, n21015, n21016, n21017,
    n21018, n21019, n21021, n21022, n21023, n21024,
    n21025, n21026, n21027, n21028, n21029, n21030,
    n21031, n21032, n21033, n21034, n21035, n21036,
    n21037, n21038, n21039, n21040, n21041, n21042,
    n21043, n21044, n21045, n21046, n21047, n21048,
    n21049, n21050, n21051, n21052, n21053, n21054,
    n21055, n21056, n21057, n21058, n21059, n21060,
    n21062, n21063, n21064, n21065, n21066, n21067,
    n21068, n21069, n21070, n21071, n21072, n21073,
    n21074, n21075, n21076, n21077, n21078, n21079,
    n21080, n21081, n21082, n21083, n21084, n21085,
    n21086, n21087, n21088, n21089, n21090, n21092,
    n21093, n21094, n21095, n21096, n21097, n21098,
    n21099, n21100, n21101, n21102, n21103, n21104,
    n21105, n21106, n21107, n21108, n21109, n21110,
    n21111, n21112, n21113, n21114, n21115, n21116,
    n21117, n21118, n21119, n21120, n21121, n21122,
    n21123, n21124, n21125, n21126, n21127, n21128,
    n21129, n21130, n21131, n21132, n21133, n21134,
    n21135, n21136, n21137, n21138, n21139, n21140,
    n21141, n21142, n21143, n21144, n21146, n21147,
    n21148, n21149, n21150, n21151, n21152, n21153,
    n21154, n21155, n21156, n21157, n21158, n21159,
    n21160, n21161, n21162, n21163, n21164, n21165,
    n21166, n21167, n21168, n21169, n21170, n21171,
    n21172, n21173, n21174, n21175, n21176, n21177,
    n21178, n21179, n21180, n21181, n21182, n21183,
    n21184, n21185, n21186, n21187, n21188, n21189,
    n21190, n21191, n21192, n21193, n21194, n21195,
    n21196, n21197, n21199, n21200, n21201, n21202,
    n21203, n21204, n21205, n21206, n21207, n21208,
    n21209, n21210, n21211, n21212, n21213, n21214,
    n21215, n21216, n21217, n21218, n21219, n21220,
    n21221, n21222, n21223, n21224, n21225, n21226,
    n21227, n21228, n21229, n21230, n21231, n21232,
    n21233, n21234, n21235, n21236, n21237, n21238,
    n21239, n21240, n21241, n21242, n21243, n21244,
    n21245, n21246, n21247, n21248, n21249, n21250,
    n21252, n21253, n21254, n21255, n21256, n21257,
    n21258, n21259, n21260, n21261, n21262, n21263,
    n21264, n21265, n21266, n21267, n21268, n21269,
    n21270, n21271, n21272, n21273, n21274, n21275,
    n21276, n21277, n21278, n21279, n21280, n21281,
    n21282, n21283, n21284, n21285, n21286, n21287,
    n21288, n21289, n21290, n21291, n21292, n21293,
    n21294, n21295, n21296, n21297, n21298, n21299,
    n21300, n21301, n21302, n21303, n21304, n21305,
    n21306, n21308, n21309, n21310, n21311, n21312,
    n21313, n21314, n21315, n21316, n21317, n21318,
    n21319, n21320, n21321, n21322, n21323, n21324,
    n21325, n21326, n21327, n21328, n21329, n21330,
    n21331, n21332, n21333, n21334, n21335, n21336,
    n21337, n21338, n21339, n21340, n21341, n21342,
    n21343, n21344, n21345, n21346, n21347, n21348,
    n21349, n21350, n21351, n21352, n21353, n21354,
    n21355, n21356, n21357, n21358, n21359, n21360,
    n21361, n21362, n21363, n21364, n21365, n21366,
    n21367, n21368, n21369, n21370, n21371, n21372,
    n21373, n21374, n21375, n21376, n21377, n21378,
    n21379, n21380, n21381, n21382, n21383, n21384,
    n21385, n21386, n21387, n21388, n21389, n21390,
    n21391, n21392, n21393, n21394, n21395, n21396,
    n21397, n21398, n21400, n21401, n21402, n21403,
    n21404, n21405, n21406, n21407, n21408, n21409,
    n21410, n21411, n21412, n21413, n21414, n21415,
    n21416, n21417, n21418, n21419, n21420, n21421,
    n21422, n21423, n21424, n21425, n21426, n21427,
    n21428, n21429, n21430, n21431, n21432, n21433,
    n21434, n21435, n21436, n21437, n21438, n21439,
    n21440, n21441, n21442, n21443, n21444, n21445,
    n21446, n21447, n21448, n21449, n21450, n21452,
    n21453, n21454, n21455, n21456, n21457, n21458,
    n21459, n21460, n21461, n21462, n21463, n21464,
    n21465, n21466, n21467, n21468, n21469, n21470,
    n21471, n21472, n21473, n21474, n21475, n21476,
    n21477, n21478, n21479, n21480, n21481, n21482,
    n21483, n21484, n21485, n21486, n21487, n21488,
    n21489, n21490, n21491, n21492, n21493, n21494,
    n21495, n21496, n21497, n21498, n21499, n21500,
    n21501, n21502, n21503, n21504, n21505, n21507,
    n21508, n21509, n21510, n21511, n21512, n21513,
    n21514, n21515, n21516, n21517, n21518, n21519,
    n21520, n21521, n21522, n21523, n21524, n21525,
    n21526, n21527, n21528, n21529, n21530, n21531,
    n21532, n21533, n21534, n21535, n21536, n21537,
    n21538, n21539, n21540, n21541, n21542, n21543,
    n21544, n21545, n21547, n21548, n21549, n21550,
    n21551, n21552, n21553, n21554, n21555, n21556,
    n21557, n21558, n21559, n21560, n21561, n21562,
    n21563, n21564, n21565, n21566, n21567, n21568,
    n21569, n21570, n21571, n21572, n21573, n21574,
    n21575, n21576, n21577, n21578, n21579, n21580,
    n21581, n21582, n21583, n21584, n21585, n21587,
    n21588, n21589, n21590, n21591, n21592, n21593,
    n21594, n21595, n21596, n21597, n21598, n21599,
    n21600, n21601, n21602, n21603, n21604, n21605,
    n21606, n21607, n21608, n21609, n21610, n21611,
    n21612, n21613, n21614, n21615, n21616, n21617,
    n21618, n21619, n21620, n21621, n21622, n21623,
    n21624, n21625, n21626, n21627, n21628, n21629,
    n21630, n21631, n21632, n21633, n21634, n21635,
    n21636, n21637, n21638, n21639, n21640, n21641,
    n21642, n21643, n21644, n21645, n21646, n21647,
    n21648, n21649, n21650, n21651, n21652, n21653,
    n21654, n21655, n21656, n21657, n21658, n21659,
    n21660, n21661, n21662, n21663, n21664, n21665,
    n21666, n21667, n21668, n21669, n21670, n21671,
    n21672, n21673, n21674, n21675, n21676, n21677,
    n21678, n21679, n21680, n21682, n21683, n21684,
    n21685, n21686, n21687, n21688, n21689, n21690,
    n21691, n21692, n21693, n21694, n21695, n21696,
    n21697, n21698, n21699, n21700, n21701, n21702,
    n21703, n21704, n21705, n21706, n21707, n21708,
    n21709, n21710, n21711, n21712, n21713, n21714,
    n21715, n21716, n21717, n21718, n21719, n21720,
    n21721, n21722, n21723, n21725, n21726, n21727,
    n21728, n21729, n21730, n21731, n21732, n21733,
    n21734, n21735, n21736, n21737, n21738, n21739,
    n21740, n21741, n21742, n21743, n21744, n21745,
    n21746, n21747, n21748, n21749, n21750, n21751,
    n21752, n21753, n21754, n21755, n21756, n21757,
    n21758, n21759, n21760, n21761, n21762, n21763,
    n21764, n21765, n21766, n21767, n21768, n21769,
    n21770, n21771, n21772, n21773, n21774, n21775,
    n21776, n21777, n21778, n21779, n21780, n21781,
    n21782, n21783, n21784, n21785, n21786, n21787,
    n21788, n21789, n21790, n21791, n21792, n21793,
    n21794, n21795, n21796, n21797, n21798, n21799,
    n21800, n21801, n21802, n21804, n21805, n21806,
    n21807, n21808, n21809, n21810, n21811, n21812,
    n21813, n21814, n21815, n21816, n21817, n21818,
    n21819, n21820, n21821, n21822, n21823, n21824,
    n21825, n21826, n21827, n21828, n21829, n21830,
    n21831, n21832, n21833, n21834, n21835, n21836,
    n21837, n21838, n21839, n21840, n21841, n21842,
    n21843, n21844, n21845, n21846, n21847, n21848,
    n21849, n21850, n21851, n21852, n21853, n21854,
    n21855, n21856, n21857, n21858, n21859, n21860,
    n21861, n21862, n21863, n21864, n21865, n21866,
    n21867, n21868, n21869, n21870, n21871, n21872,
    n21873, n21874, n21875, n21876, n21877, n21878,
    n21879, n21880, n21881, n21883, n21884, n21885,
    n21886, n21887, n21888, n21889, n21890, n21891,
    n21892, n21893, n21894, n21895, n21896, n21897,
    n21898, n21899, n21900, n21901, n21902, n21903,
    n21904, n21905, n21906, n21907, n21908, n21909,
    n21910, n21911, n21912, n21913, n21914, n21915,
    n21916, n21917, n21918, n21919, n21920, n21921,
    n21922, n21923, n21924, n21925, n21926, n21927,
    n21928, n21929, n21930, n21931, n21932, n21933,
    n21934, n21935, n21936, n21937, n21938, n21939,
    n21940, n21941, n21942, n21943, n21944, n21945,
    n21946, n21947, n21948, n21949, n21950, n21951,
    n21952, n21953, n21954, n21955, n21956, n21957,
    n21958, n21959, n21960, n21962, n21963, n21964,
    n21965, n21966, n21967, n21968, n21969, n21970,
    n21971, n21972, n21973, n21974, n21975, n21976,
    n21977, n21978, n21979, n21980, n21981, n21982,
    n21983, n21984, n21985, n21986, n21987, n21988,
    n21989, n21990, n21991, n21992, n21993, n21994,
    n21995, n21996, n21997, n21998, n21999, n22000,
    n22001, n22002, n22003, n22004, n22005, n22006,
    n22007, n22008, n22009, n22010, n22011, n22012,
    n22013, n22014, n22015, n22016, n22017, n22018,
    n22019, n22020, n22021, n22022, n22023, n22024,
    n22025, n22026, n22027, n22028, n22029, n22030,
    n22031, n22032, n22033, n22034, n22035, n22036,
    n22037, n22038, n22039, n22041, n22042, n22043,
    n22044, n22045, n22046, n22047, n22048, n22049,
    n22050, n22051, n22052, n22053, n22054, n22055,
    n22056, n22057, n22058, n22059, n22060, n22061,
    n22062, n22063, n22064, n22065, n22066, n22067,
    n22068, n22069, n22070, n22071, n22072, n22073,
    n22074, n22075, n22076, n22077, n22078, n22079,
    n22080, n22081, n22082, n22083, n22084, n22085,
    n22086, n22087, n22088, n22089, n22090, n22091,
    n22092, n22093, n22094, n22095, n22096, n22097,
    n22098, n22099, n22100, n22101, n22102, n22103,
    n22104, n22105, n22106, n22107, n22108, n22109,
    n22110, n22111, n22112, n22113, n22114, n22115,
    n22116, n22117, n22118, n22120, n22121, n22122,
    n22123, n22124, n22125, n22126, n22127, n22128,
    n22129, n22130, n22131, n22132, n22133, n22134,
    n22135, n22136, n22137, n22138, n22139, n22140,
    n22141, n22142, n22143, n22144, n22145, n22146,
    n22147, n22148, n22149, n22150, n22151, n22152,
    n22153, n22154, n22155, n22156, n22157, n22158,
    n22159, n22160, n22161, n22162, n22163, n22164,
    n22165, n22166, n22167, n22168, n22169, n22170,
    n22171, n22172, n22173, n22174, n22175, n22176,
    n22177, n22178, n22179, n22180, n22181, n22182,
    n22183, n22184, n22185, n22186, n22187, n22188,
    n22189, n22190, n22191, n22192, n22193, n22194,
    n22195, n22196, n22197, n22198, n22199, n22200,
    n22201, n22202, n22203, n22204, n22205, n22206,
    n22207, n22208, n22209, n22210, n22211, n22212,
    n22213, n22214, n22215, n22216, n22217, n22218,
    n22219, n22220, n22221, n22222, n22223, n22224,
    n22225, n22226, n22227, n22228, n22229, n22230,
    n22231, n22232, n22233, n22234, n22235, n22236,
    n22237, n22238, n22239, n22240, n22241, n22242,
    n22243, n22244, n22245, n22246, n22247, n22248,
    n22249, n22250, n22251, n22252, n22253, n22254,
    n22255, n22256, n22257, n22258, n22259, n22260,
    n22261, n22262, n22263, n22264, n22265, n22266,
    n22267, n22268, n22269, n22270, n22271, n22272,
    n22273, n22274, n22275, n22276, n22277, n22278,
    n22279, n22280, n22281, n22282, n22283, n22284,
    n22285, n22286, n22287, n22288, n22289, n22290,
    n22291, n22292, n22293, n22294, n22295, n22296,
    n22297, n22298, n22299, n22300, n22301, n22302,
    n22303, n22304, n22305, n22306, n22307, n22308,
    n22309, n22310, n22311, n22312, n22313, n22314,
    n22315, n22316, n22317, n22318, n22319, n22320,
    n22321, n22322, n22323, n22324, n22325, n22326,
    n22327, n22328, n22329, n22330, n22331, n22332,
    n22333, n22334, n22335, n22336, n22337, n22338,
    n22339, n22340, n22341, n22342, n22343, n22344,
    n22345, n22346, n22347, n22348, n22349, n22350,
    n22351, n22352, n22353, n22354, n22355, n22356,
    n22357, n22358, n22359, n22360, n22361, n22362,
    n22363, n22364, n22365, n22366, n22367, n22368,
    n22369, n22370, n22371, n22372, n22373, n22374,
    n22375, n22376, n22377, n22378, n22379, n22380,
    n22381, n22382, n22383, n22384, n22385, n22386,
    n22387, n22388, n22389, n22390, n22391, n22392,
    n22393, n22394, n22395, n22396, n22397, n22398,
    n22399, n22400, n22401, n22402, n22403, n22404,
    n22405, n22406, n22407, n22408, n22409, n22410,
    n22411, n22412, n22413, n22414, n22415, n22416,
    n22417, n22418, n22419, n22420, n22421, n22422,
    n22423, n22424, n22425, n22426, n22427, n22428,
    n22429, n22430, n22431, n22432, n22433, n22434,
    n22435, n22436, n22437, n22438, n22439, n22440,
    n22441, n22442, n22443, n22444, n22445, n22446,
    n22447, n22448, n22449, n22450, n22451, n22452,
    n22453, n22454, n22455, n22456, n22457, n22458,
    n22459, n22460, n22461, n22462, n22463, n22464,
    n22465, n22466, n22467, n22468, n22469, n22470,
    n22471, n22472, n22473, n22474, n22475, n22476,
    n22477, n22478, n22479, n22480, n22481, n22482,
    n22483, n22484, n22485, n22486, n22487, n22488,
    n22489, n22490, n22491, n22492, n22493, n22494,
    n22495, n22496, n22497, n22498, n22499, n22500,
    n22501, n22502, n22503, n22504, n22505, n22506,
    n22507, n22508, n22509, n22510, n22511, n22512,
    n22513, n22514, n22515, n22516, n22517, n22518,
    n22519, n22520, n22521, n22522, n22523, n22524,
    n22525, n22526, n22527, n22528, n22529, n22530,
    n22531, n22532, n22533, n22534, n22535, n22536,
    n22537, n22538, n22539, n22540, n22541, n22542,
    n22543, n22544, n22545, n22546, n22547, n22548,
    n22549, n22550, n22551, n22552, n22553, n22554,
    n22555, n22556, n22557, n22558, n22559, n22560,
    n22561, n22562, n22563, n22564, n22565, n22566,
    n22567, n22568, n22569, n22570, n22571, n22572,
    n22573, n22574, n22575, n22576, n22577, n22578,
    n22579, n22580, n22581, n22582, n22583, n22584,
    n22585, n22586, n22587, n22588, n22589, n22591,
    n22592, n22593, n22594, n22595, n22596, n22597,
    n22598, n22599, n22600, n22601, n22602, n22603,
    n22604, n22605, n22606, n22607, n22608, n22609,
    n22610, n22611, n22612, n22613, n22614, n22615,
    n22616, n22617, n22618, n22619, n22620, n22621,
    n22622, n22623, n22624, n22625, n22626, n22627,
    n22628, n22629, n22630, n22631, n22632, n22633,
    n22634, n22635, n22636, n22637, n22638, n22639,
    n22640, n22641, n22642, n22643, n22644, n22645,
    n22646, n22647, n22648, n22649, n22650, n22651,
    n22652, n22653, n22654, n22655, n22656, n22657,
    n22658, n22659, n22660, n22661, n22662, n22663,
    n22664, n22665, n22666, n22667, n22668, n22669,
    n22670, n22671, n22672, n22673, n22674, n22675,
    n22676, n22677, n22678, n22679, n22680, n22681,
    n22682, n22683, n22684, n22685, n22686, n22687,
    n22688, n22689, n22690, n22691, n22692, n22693,
    n22694, n22695, n22696, n22697, n22698, n22699,
    n22700, n22701, n22702, n22703, n22704, n22705,
    n22706, n22707, n22708, n22709, n22710, n22711,
    n22712, n22713, n22714, n22715, n22716, n22717,
    n22718, n22719, n22720, n22721, n22722, n22723,
    n22724, n22725, n22726, n22727, n22728, n22729,
    n22730, n22731, n22732, n22733, n22734, n22735,
    n22736, n22737, n22738, n22739, n22740, n22741,
    n22742, n22743, n22744, n22745, n22746, n22747,
    n22748, n22749, n22750, n22751, n22752, n22753,
    n22754, n22755, n22756, n22757, n22758, n22759,
    n22760, n22761, n22762, n22763, n22764, n22765,
    n22766, n22767, n22768, n22769, n22770, n22771,
    n22772, n22773, n22774, n22775, n22776, n22777,
    n22778, n22779, n22780, n22781, n22782, n22783,
    n22784, n22785, n22786, n22787, n22788, n22789,
    n22790, n22791, n22792, n22793, n22794, n22795,
    n22796, n22797, n22798, n22799, n22800, n22801,
    n22802, n22803, n22804, n22805, n22806, n22807,
    n22808, n22809, n22810, n22811, n22812, n22813,
    n22814, n22815, n22816, n22817, n22818, n22819,
    n22820, n22821, n22822, n22823, n22824, n22825,
    n22826, n22827, n22828, n22829, n22830, n22831,
    n22832, n22833, n22834, n22835, n22836, n22837,
    n22838, n22839, n22840, n22841, n22842, n22843,
    n22844, n22845, n22846, n22847, n22848, n22849,
    n22850, n22851, n22852, n22853, n22854, n22855,
    n22856, n22857, n22858, n22859, n22860, n22861,
    n22862, n22863, n22864, n22865, n22866, n22867,
    n22868, n22869, n22870, n22871, n22872, n22873,
    n22874, n22875, n22876, n22877, n22878, n22879,
    n22880, n22881, n22882, n22883, n22884, n22885,
    n22886, n22887, n22888, n22889, n22890, n22891,
    n22892, n22893, n22894, n22895, n22896, n22897,
    n22898, n22899, n22900, n22901, n22902, n22903,
    n22904, n22905, n22906, n22907, n22908, n22909,
    n22910, n22911, n22912, n22913, n22914, n22915,
    n22916, n22917, n22918, n22919, n22920, n22921,
    n22922, n22923, n22924, n22925, n22926, n22927,
    n22928, n22929, n22930, n22931, n22932, n22933,
    n22934, n22935, n22936, n22937, n22938, n22939,
    n22940, n22941, n22942, n22943, n22944, n22945,
    n22946, n22947, n22948, n22949, n22950, n22951,
    n22952, n22953, n22954, n22955, n22956, n22957,
    n22958, n22959, n22960, n22961, n22962, n22963,
    n22964, n22965, n22966, n22967, n22968, n22969,
    n22970, n22971, n22972, n22973, n22974, n22975,
    n22976, n22977, n22978, n22979, n22980, n22981,
    n22982, n22983, n22984, n22985, n22986, n22987,
    n22988, n22989, n22990, n22991, n22992, n22993,
    n22994, n22995, n22996, n22997, n22998, n22999,
    n23000, n23001, n23002, n23003, n23004, n23005,
    n23006, n23007, n23008, n23009, n23010, n23011,
    n23012, n23013, n23014, n23015, n23016, n23017,
    n23018, n23019, n23020, n23021, n23022, n23023,
    n23024, n23025, n23026, n23027, n23028, n23029,
    n23030, n23031, n23032, n23033, n23034, n23035,
    n23036, n23037, n23038, n23039, n23040, n23041,
    n23042, n23043, n23044, n23045, n23046, n23047,
    n23048, n23049, n23050, n23051, n23052, n23053,
    n23054, n23055, n23056, n23057, n23058, n23059,
    n23060, n23061, n23062, n23063, n23064, n23065,
    n23066, n23067, n23068, n23069, n23071, n23072,
    n23073, n23074, n23075, n23076, n23077, n23078,
    n23079, n23080, n23081, n23082, n23083, n23084,
    n23085, n23086, n23087, n23088, n23089, n23090,
    n23091, n23092, n23093, n23094, n23095, n23096,
    n23097, n23098, n23099, n23100, n23101, n23102,
    n23103, n23104, n23105, n23106, n23107, n23108,
    n23109, n23110, n23111, n23112, n23113, n23114,
    n23115, n23116, n23117, n23118, n23119, n23120,
    n23121, n23122, n23123, n23124, n23125, n23126,
    n23127, n23128, n23129, n23130, n23131, n23132,
    n23133, n23134, n23135, n23136, n23137, n23138,
    n23139, n23140, n23141, n23142, n23143, n23144,
    n23145, n23146, n23147, n23148, n23149, n23150,
    n23151, n23152, n23153, n23154, n23155, n23156,
    n23157, n23158, n23159, n23160, n23161, n23162,
    n23163, n23164, n23165, n23166, n23167, n23168,
    n23169, n23170, n23171, n23172, n23173, n23174,
    n23175, n23176, n23177, n23178, n23179, n23180,
    n23181, n23182, n23183, n23184, n23185, n23186,
    n23187, n23188, n23189, n23190, n23191, n23192,
    n23193, n23194, n23195, n23196, n23197, n23198,
    n23199, n23200, n23201, n23202, n23203, n23204,
    n23205, n23206, n23207, n23208, n23209, n23210,
    n23211, n23212, n23213, n23214, n23215, n23216,
    n23217, n23218, n23219, n23220, n23221, n23222,
    n23223, n23224, n23225, n23226, n23227, n23228,
    n23229, n23230, n23231, n23232, n23233, n23234,
    n23235, n23236, n23237, n23238, n23239, n23240,
    n23241, n23242, n23243, n23244, n23245, n23246,
    n23247, n23248, n23249, n23250, n23251, n23252,
    n23253, n23254, n23255, n23256, n23257, n23258,
    n23259, n23260, n23261, n23262, n23263, n23264,
    n23265, n23266, n23267, n23268, n23269, n23270,
    n23271, n23272, n23273, n23274, n23275, n23276,
    n23277, n23278, n23279, n23280, n23281, n23282,
    n23283, n23284, n23285, n23286, n23287, n23288,
    n23289, n23290, n23291, n23292, n23293, n23294,
    n23295, n23296, n23297, n23298, n23299, n23300,
    n23301, n23302, n23303, n23304, n23305, n23306,
    n23307, n23308, n23309, n23310, n23311, n23312,
    n23313, n23314, n23315, n23316, n23317, n23318,
    n23319, n23320, n23321, n23322, n23323, n23324,
    n23325, n23326, n23327, n23328, n23329, n23330,
    n23331, n23332, n23333, n23334, n23335, n23336,
    n23337, n23338, n23339, n23340, n23341, n23342,
    n23343, n23344, n23345, n23346, n23347, n23348,
    n23349, n23350, n23351, n23352, n23353, n23354,
    n23355, n23356, n23357, n23358, n23359, n23360,
    n23361, n23362, n23363, n23364, n23365, n23366,
    n23367, n23368, n23369, n23370, n23371, n23372,
    n23373, n23374, n23375, n23376, n23377, n23378,
    n23379, n23380, n23381, n23382, n23383, n23384,
    n23385, n23386, n23387, n23388, n23389, n23390,
    n23391, n23392, n23393, n23394, n23395, n23396,
    n23397, n23398, n23399, n23400, n23401, n23402,
    n23403, n23404, n23405, n23406, n23407, n23408,
    n23409, n23410, n23411, n23412, n23413, n23414,
    n23415, n23416, n23417, n23418, n23419, n23420,
    n23421, n23422, n23423, n23424, n23425, n23426,
    n23427, n23428, n23429, n23430, n23431, n23432,
    n23433, n23434, n23435, n23436, n23437, n23438,
    n23439, n23440, n23441, n23442, n23443, n23444,
    n23445, n23446, n23447, n23448, n23449, n23450,
    n23451, n23452, n23453, n23454, n23455, n23456,
    n23457, n23458, n23459, n23460, n23461, n23462,
    n23463, n23464, n23465, n23466, n23467, n23468,
    n23469, n23470, n23471, n23472, n23473, n23474,
    n23475, n23476, n23477, n23478, n23479, n23480,
    n23481, n23482, n23483, n23484, n23485, n23486,
    n23487, n23488, n23489, n23490, n23491, n23492,
    n23493, n23494, n23495, n23496, n23497, n23498,
    n23499, n23500, n23501, n23502, n23503, n23504,
    n23505, n23506, n23507, n23508, n23509, n23510,
    n23511, n23512, n23513, n23514, n23515, n23516,
    n23517, n23518, n23519, n23520, n23521, n23522,
    n23523, n23524, n23525, n23526, n23527, n23528,
    n23529, n23530, n23531, n23532, n23533, n23534,
    n23535, n23536, n23537, n23538, n23539, n23541,
    n23542, n23543, n23544, n23545, n23546, n23547,
    n23548, n23549, n23550, n23551, n23552, n23553,
    n23554, n23555, n23556, n23557, n23558, n23559,
    n23560, n23561, n23562, n23563, n23564, n23565,
    n23566, n23567, n23568, n23569, n23570, n23571,
    n23572, n23573, n23574, n23575, n23576, n23577,
    n23578, n23579, n23580, n23581, n23582, n23583,
    n23584, n23585, n23586, n23587, n23588, n23589,
    n23590, n23591, n23592, n23593, n23594, n23595,
    n23596, n23597, n23598, n23599, n23600, n23601,
    n23602, n23603, n23604, n23605, n23606, n23607,
    n23608, n23609, n23610, n23611, n23612, n23613,
    n23614, n23615, n23616, n23617, n23618, n23619,
    n23620, n23621, n23622, n23623, n23624, n23625,
    n23626, n23627, n23628, n23629, n23630, n23631,
    n23632, n23633, n23634, n23635, n23636, n23637,
    n23638, n23639, n23640, n23641, n23642, n23643,
    n23644, n23645, n23646, n23647, n23648, n23649,
    n23650, n23651, n23652, n23653, n23654, n23655,
    n23656, n23657, n23658, n23659, n23660, n23661,
    n23662, n23663, n23664, n23665, n23666, n23667,
    n23668, n23669, n23670, n23671, n23672, n23673,
    n23674, n23675, n23676, n23677, n23678, n23679,
    n23680, n23681, n23682, n23683, n23684, n23685,
    n23686, n23687, n23688, n23689, n23690, n23691,
    n23692, n23693, n23694, n23695, n23696, n23697,
    n23698, n23699, n23700, n23701, n23702, n23703,
    n23704, n23705, n23706, n23707, n23708, n23709,
    n23710, n23711, n23712, n23713, n23714, n23715,
    n23716, n23717, n23718, n23719, n23720, n23721,
    n23722, n23723, n23724, n23725, n23726, n23727,
    n23728, n23729, n23730, n23731, n23732, n23733,
    n23734, n23735, n23736, n23737, n23738, n23739,
    n23740, n23741, n23742, n23743, n23744, n23745,
    n23746, n23747, n23748, n23749, n23750, n23751,
    n23752, n23753, n23754, n23755, n23756, n23757,
    n23758, n23759, n23760, n23761, n23762, n23763,
    n23764, n23765, n23766, n23767, n23768, n23769,
    n23770, n23771, n23772, n23773, n23774, n23775,
    n23776, n23777, n23778, n23779, n23780, n23781,
    n23782, n23783, n23784, n23785, n23786, n23787,
    n23788, n23789, n23790, n23791, n23792, n23793,
    n23794, n23795, n23796, n23797, n23798, n23799,
    n23800, n23801, n23802, n23803, n23804, n23805,
    n23806, n23807, n23808, n23809, n23810, n23811,
    n23812, n23813, n23814, n23815, n23816, n23817,
    n23818, n23819, n23820, n23821, n23822, n23823,
    n23824, n23825, n23826, n23827, n23828, n23829,
    n23830, n23831, n23832, n23833, n23834, n23835,
    n23836, n23837, n23838, n23839, n23840, n23841,
    n23842, n23843, n23844, n23845, n23846, n23847,
    n23848, n23849, n23850, n23851, n23852, n23853,
    n23854, n23855, n23856, n23857, n23858, n23859,
    n23860, n23861, n23862, n23863, n23864, n23865,
    n23866, n23867, n23868, n23869, n23870, n23871,
    n23872, n23873, n23874, n23875, n23876, n23877,
    n23878, n23879, n23880, n23881, n23882, n23883,
    n23884, n23885, n23886, n23887, n23888, n23889,
    n23890, n23891, n23892, n23893, n23894, n23895,
    n23896, n23897, n23898, n23899, n23900, n23901,
    n23902, n23903, n23904, n23905, n23906, n23907,
    n23908, n23909, n23910, n23911, n23912, n23913,
    n23914, n23915, n23916, n23917, n23918, n23919,
    n23920, n23921, n23922, n23923, n23924, n23925,
    n23926, n23927, n23928, n23929, n23930, n23931,
    n23932, n23933, n23934, n23935, n23936, n23937,
    n23938, n23939, n23940, n23941, n23942, n23943,
    n23944, n23945, n23946, n23947, n23948, n23949,
    n23950, n23951, n23952, n23953, n23954, n23955,
    n23956, n23957, n23958, n23959, n23960, n23961,
    n23962, n23963, n23964, n23965, n23966, n23967,
    n23968, n23969, n23970, n23971, n23972, n23973,
    n23974, n23975, n23976, n23977, n23978, n23979,
    n23981, n23982, n23983, n23984, n23985, n23986,
    n23987, n23988, n23989, n23990, n23991, n23992,
    n23993, n23994, n23995, n23996, n23997, n23998,
    n23999, n24000, n24001, n24002, n24003, n24004,
    n24005, n24006, n24007, n24008, n24009, n24010,
    n24011, n24012, n24013, n24014, n24015, n24016,
    n24017, n24018, n24019, n24020, n24021, n24022,
    n24023, n24024, n24025, n24026, n24027, n24028,
    n24029, n24030, n24031, n24032, n24033, n24034,
    n24035, n24036, n24037, n24038, n24039, n24040,
    n24041, n24042, n24043, n24044, n24045, n24046,
    n24047, n24048, n24049, n24050, n24051, n24052,
    n24053, n24054, n24055, n24056, n24057, n24058,
    n24059, n24060, n24061, n24062, n24063, n24064,
    n24065, n24066, n24067, n24068, n24069, n24070,
    n24071, n24072, n24073, n24074, n24075, n24076,
    n24077, n24078, n24079, n24080, n24081, n24082,
    n24083, n24084, n24085, n24086, n24087, n24088,
    n24089, n24090, n24091, n24092, n24093, n24094,
    n24095, n24096, n24097, n24098, n24099, n24100,
    n24101, n24102, n24103, n24104, n24105, n24106,
    n24107, n24108, n24109, n24110, n24111, n24112,
    n24113, n24114, n24115, n24116, n24117, n24118,
    n24119, n24120, n24121, n24122, n24123, n24124,
    n24125, n24126, n24127, n24128, n24129, n24130,
    n24131, n24132, n24133, n24134, n24135, n24136,
    n24137, n24138, n24139, n24140, n24141, n24142,
    n24143, n24144, n24145, n24146, n24147, n24148,
    n24149, n24150, n24151, n24152, n24153, n24154,
    n24155, n24156, n24157, n24158, n24159, n24160,
    n24161, n24162, n24163, n24164, n24165, n24166,
    n24167, n24168, n24169, n24170, n24171, n24172,
    n24173, n24174, n24175, n24176, n24177, n24178,
    n24179, n24180, n24181, n24182, n24183, n24184,
    n24185, n24186, n24187, n24188, n24189, n24190,
    n24191, n24192, n24193, n24194, n24195, n24196,
    n24197, n24198, n24199, n24200, n24201, n24202,
    n24203, n24204, n24205, n24206, n24207, n24208,
    n24209, n24210, n24211, n24212, n24213, n24214,
    n24215, n24216, n24217, n24218, n24219, n24220,
    n24221, n24222, n24223, n24224, n24225, n24226,
    n24227, n24228, n24229, n24230, n24231, n24232,
    n24233, n24234, n24235, n24236, n24237, n24238,
    n24239, n24240, n24241, n24242, n24243, n24244,
    n24245, n24246, n24247, n24248, n24249, n24250,
    n24251, n24252, n24253, n24254, n24255, n24256,
    n24257, n24258, n24259, n24260, n24261, n24262,
    n24263, n24264, n24265, n24266, n24267, n24268,
    n24269, n24270, n24271, n24272, n24273, n24274,
    n24275, n24276, n24277, n24278, n24279, n24280,
    n24281, n24282, n24283, n24284, n24285, n24286,
    n24287, n24288, n24289, n24290, n24291, n24292,
    n24293, n24294, n24295, n24296, n24297, n24298,
    n24299, n24300, n24301, n24302, n24303, n24304,
    n24305, n24306, n24307, n24308, n24309, n24310,
    n24311, n24312, n24313, n24314, n24315, n24316,
    n24317, n24318, n24319, n24320, n24321, n24322,
    n24323, n24324, n24325, n24326, n24327, n24328,
    n24329, n24330, n24331, n24332, n24333, n24334,
    n24335, n24336, n24337, n24338, n24339, n24340,
    n24341, n24342, n24343, n24344, n24345, n24346,
    n24347, n24348, n24349, n24350, n24351, n24352,
    n24353, n24354, n24355, n24356, n24357, n24358,
    n24359, n24360, n24361, n24362, n24363, n24364,
    n24365, n24366, n24367, n24368, n24369, n24370,
    n24371, n24372, n24373, n24374, n24375, n24376,
    n24377, n24378, n24379, n24380, n24381, n24382,
    n24383, n24384, n24385, n24386, n24387, n24388,
    n24389, n24390, n24391, n24392, n24393, n24394,
    n24395, n24396, n24397, n24398, n24399, n24400,
    n24401, n24402, n24403, n24404, n24405, n24406,
    n24407, n24408, n24409, n24410, n24411, n24412,
    n24413, n24414, n24415, n24416, n24417, n24418,
    n24419, n24420, n24421, n24422, n24423, n24424,
    n24425, n24426, n24427, n24428, n24429, n24430,
    n24431, n24432, n24433, n24434, n24435, n24436,
    n24437, n24438, n24439, n24440, n24441, n24442,
    n24443, n24444, n24445, n24446, n24447, n24448,
    n24449, n24450, n24451, n24452, n24453, n24454,
    n24455, n24456, n24457, n24458, n24460, n24461,
    n24462, n24463, n24464, n24465, n24466, n24467,
    n24468, n24469, n24470, n24471, n24472, n24473,
    n24474, n24475, n24476, n24477, n24478, n24479,
    n24480, n24481, n24482, n24483, n24484, n24485,
    n24486, n24487, n24488, n24489, n24490, n24491,
    n24492, n24493, n24494, n24495, n24496, n24497,
    n24498, n24499, n24500, n24501, n24502, n24503,
    n24504, n24505, n24506, n24507, n24508, n24509,
    n24510, n24511, n24512, n24513, n24514, n24515,
    n24516, n24517, n24518, n24519, n24520, n24521,
    n24522, n24523, n24524, n24525, n24526, n24527,
    n24528, n24529, n24530, n24531, n24532, n24533,
    n24534, n24535, n24536, n24537, n24538, n24539,
    n24540, n24541, n24542, n24543, n24544, n24545,
    n24546, n24547, n24548, n24549, n24550, n24551,
    n24552, n24553, n24554, n24555, n24556, n24557,
    n24558, n24559, n24560, n24561, n24562, n24563,
    n24564, n24565, n24566, n24567, n24568, n24569,
    n24570, n24571, n24572, n24573, n24574, n24575,
    n24576, n24577, n24578, n24579, n24580, n24581,
    n24582, n24583, n24584, n24585, n24586, n24587,
    n24588, n24589, n24590, n24591, n24592, n24593,
    n24594, n24595, n24596, n24597, n24598, n24599,
    n24600, n24601, n24602, n24603, n24604, n24605,
    n24606, n24607, n24608, n24609, n24610, n24611,
    n24612, n24613, n24614, n24615, n24616, n24617,
    n24618, n24619, n24620, n24621, n24622, n24623,
    n24624, n24625, n24626, n24627, n24628, n24629,
    n24630, n24631, n24632, n24633, n24634, n24635,
    n24636, n24637, n24638, n24639, n24640, n24641,
    n24642, n24643, n24644, n24645, n24646, n24647,
    n24648, n24649, n24650, n24651, n24652, n24653,
    n24654, n24655, n24656, n24657, n24658, n24659,
    n24660, n24661, n24662, n24663, n24664, n24665,
    n24666, n24667, n24668, n24669, n24670, n24671,
    n24672, n24673, n24674, n24675, n24676, n24677,
    n24678, n24679, n24680, n24681, n24682, n24683,
    n24684, n24685, n24686, n24687, n24688, n24689,
    n24690, n24691, n24692, n24693, n24694, n24695,
    n24696, n24697, n24698, n24699, n24700, n24701,
    n24702, n24703, n24704, n24705, n24706, n24707,
    n24708, n24709, n24710, n24711, n24712, n24713,
    n24714, n24715, n24716, n24717, n24718, n24719,
    n24720, n24721, n24722, n24723, n24724, n24725,
    n24726, n24727, n24728, n24729, n24730, n24731,
    n24732, n24733, n24734, n24735, n24736, n24737,
    n24738, n24739, n24740, n24741, n24742, n24743,
    n24744, n24745, n24746, n24747, n24748, n24749,
    n24750, n24751, n24752, n24753, n24754, n24755,
    n24756, n24757, n24758, n24759, n24760, n24761,
    n24762, n24763, n24764, n24765, n24766, n24767,
    n24768, n24769, n24770, n24771, n24772, n24773,
    n24774, n24775, n24776, n24777, n24778, n24779,
    n24780, n24781, n24782, n24783, n24784, n24785,
    n24786, n24787, n24788, n24789, n24790, n24791,
    n24792, n24793, n24794, n24795, n24796, n24797,
    n24798, n24799, n24800, n24801, n24802, n24803,
    n24804, n24805, n24806, n24807, n24808, n24809,
    n24810, n24811, n24812, n24813, n24814, n24815,
    n24816, n24817, n24818, n24819, n24820, n24821,
    n24822, n24823, n24824, n24825, n24826, n24827,
    n24828, n24829, n24830, n24831, n24832, n24833,
    n24834, n24835, n24836, n24837, n24838, n24839,
    n24840, n24841, n24842, n24843, n24844, n24845,
    n24846, n24847, n24848, n24849, n24850, n24851,
    n24852, n24853, n24854, n24855, n24856, n24857,
    n24858, n24859, n24860, n24861, n24862, n24863,
    n24864, n24865, n24866, n24867, n24868, n24869,
    n24870, n24871, n24872, n24873, n24874, n24875,
    n24876, n24877, n24878, n24879, n24880, n24881,
    n24882, n24883, n24884, n24885, n24886, n24887,
    n24888, n24889, n24890, n24891, n24892, n24893,
    n24894, n24895, n24896, n24897, n24898, n24899,
    n24900, n24901, n24902, n24903, n24904, n24905,
    n24906, n24907, n24908, n24909, n24910, n24911,
    n24912, n24913, n24914, n24915, n24916, n24917,
    n24918, n24919, n24920, n24921, n24922, n24923,
    n24924, n24925, n24927, n24928, n24929, n24930,
    n24931, n24932, n24933, n24934, n24935, n24936,
    n24937, n24938, n24939, n24940, n24941, n24942,
    n24943, n24944, n24945, n24946, n24947, n24948,
    n24949, n24950, n24951, n24952, n24953, n24954,
    n24955, n24956, n24957, n24958, n24959, n24960,
    n24961, n24962, n24963, n24964, n24965, n24966,
    n24967, n24968, n24969, n24970, n24971, n24972,
    n24973, n24974, n24975, n24976, n24977, n24978,
    n24979, n24980, n24981, n24982, n24983, n24984,
    n24985, n24986, n24987, n24988, n24989, n24990,
    n24991, n24992, n24993, n24994, n24995, n24996,
    n24997, n24998, n24999, n25000, n25001, n25002,
    n25003, n25004, n25005, n25006, n25007, n25008,
    n25009, n25010, n25011, n25012, n25013, n25014,
    n25015, n25016, n25017, n25018, n25019, n25020,
    n25021, n25022, n25023, n25024, n25025, n25026,
    n25027, n25028, n25029, n25030, n25031, n25032,
    n25033, n25034, n25035, n25036, n25037, n25038,
    n25039, n25040, n25041, n25042, n25043, n25044,
    n25045, n25046, n25047, n25048, n25049, n25050,
    n25051, n25052, n25053, n25054, n25055, n25056,
    n25057, n25058, n25059, n25060, n25061, n25062,
    n25063, n25064, n25065, n25066, n25067, n25068,
    n25069, n25070, n25071, n25072, n25073, n25074,
    n25075, n25076, n25077, n25078, n25079, n25080,
    n25081, n25082, n25083, n25084, n25085, n25086,
    n25087, n25088, n25089, n25090, n25091, n25092,
    n25093, n25094, n25095, n25096, n25097, n25098,
    n25099, n25100, n25101, n25102, n25103, n25104,
    n25105, n25106, n25107, n25108, n25109, n25110,
    n25111, n25112, n25113, n25114, n25115, n25116,
    n25117, n25118, n25119, n25120, n25121, n25122,
    n25123, n25124, n25125, n25126, n25127, n25128,
    n25129, n25130, n25131, n25132, n25133, n25134,
    n25135, n25136, n25137, n25138, n25139, n25140,
    n25141, n25142, n25143, n25144, n25145, n25146,
    n25147, n25148, n25149, n25150, n25151, n25152,
    n25153, n25154, n25155, n25156, n25157, n25158,
    n25159, n25160, n25161, n25162, n25163, n25164,
    n25165, n25166, n25167, n25168, n25169, n25170,
    n25171, n25172, n25173, n25174, n25175, n25176,
    n25177, n25178, n25179, n25180, n25181, n25182,
    n25183, n25184, n25185, n25186, n25187, n25188,
    n25189, n25190, n25191, n25192, n25193, n25194,
    n25195, n25196, n25197, n25198, n25199, n25200,
    n25201, n25202, n25203, n25204, n25205, n25206,
    n25207, n25208, n25209, n25210, n25211, n25212,
    n25213, n25214, n25215, n25216, n25217, n25218,
    n25219, n25220, n25221, n25222, n25223, n25224,
    n25225, n25226, n25227, n25228, n25229, n25230,
    n25231, n25232, n25233, n25234, n25235, n25236,
    n25237, n25238, n25239, n25240, n25241, n25242,
    n25243, n25244, n25245, n25246, n25247, n25248,
    n25249, n25250, n25251, n25252, n25253, n25254,
    n25255, n25256, n25257, n25258, n25259, n25260,
    n25261, n25262, n25263, n25264, n25265, n25266,
    n25267, n25268, n25269, n25270, n25271, n25272,
    n25273, n25274, n25275, n25276, n25277, n25278,
    n25279, n25280, n25281, n25282, n25283, n25284,
    n25285, n25286, n25287, n25288, n25289, n25290,
    n25291, n25292, n25293, n25294, n25295, n25296,
    n25297, n25298, n25299, n25300, n25301, n25302,
    n25303, n25304, n25305, n25306, n25307, n25308,
    n25309, n25310, n25311, n25312, n25313, n25314,
    n25315, n25316, n25317, n25318, n25319, n25320,
    n25321, n25322, n25323, n25324, n25325, n25326,
    n25327, n25328, n25329, n25330, n25331, n25332,
    n25333, n25334, n25335, n25336, n25337, n25338,
    n25339, n25340, n25341, n25342, n25343, n25344,
    n25345, n25346, n25347, n25348, n25349, n25350,
    n25351, n25352, n25353, n25354, n25355, n25356,
    n25357, n25358, n25359, n25360, n25361, n25362,
    n25363, n25364, n25365, n25366, n25367, n25368,
    n25369, n25370, n25371, n25372, n25373, n25374,
    n25375, n25376, n25377, n25378, n25379, n25380,
    n25381, n25382, n25383, n25384, n25385, n25386,
    n25387, n25388, n25389, n25390, n25391, n25392,
    n25393, n25394, n25395, n25396, n25397, n25398,
    n25399, n25400, n25401, n25402, n25403, n25405,
    n25406, n25407, n25408, n25409, n25410, n25411,
    n25412, n25413, n25414, n25415, n25416, n25417,
    n25418, n25419, n25420, n25421, n25422, n25423,
    n25424, n25425, n25426, n25427, n25428, n25429,
    n25430, n25431, n25432, n25433, n25434, n25435,
    n25436, n25437, n25438, n25439, n25440, n25441,
    n25442, n25443, n25444, n25445, n25446, n25447,
    n25448, n25449, n25450, n25451, n25452, n25453,
    n25454, n25455, n25456, n25457, n25458, n25459,
    n25460, n25461, n25462, n25463, n25464, n25465,
    n25466, n25467, n25468, n25469, n25470, n25471,
    n25472, n25473, n25474, n25475, n25476, n25477,
    n25478, n25479, n25480, n25481, n25482, n25483,
    n25484, n25485, n25486, n25487, n25488, n25489,
    n25490, n25491, n25492, n25493, n25494, n25495,
    n25496, n25497, n25498, n25499, n25500, n25501,
    n25502, n25503, n25504, n25505, n25506, n25507,
    n25508, n25509, n25510, n25511, n25512, n25513,
    n25514, n25515, n25516, n25517, n25518, n25519,
    n25520, n25521, n25522, n25523, n25524, n25525,
    n25526, n25527, n25528, n25529, n25530, n25531,
    n25532, n25533, n25534, n25535, n25536, n25537,
    n25538, n25539, n25540, n25541, n25542, n25543,
    n25544, n25545, n25546, n25547, n25548, n25549,
    n25550, n25551, n25552, n25553, n25554, n25555,
    n25556, n25557, n25558, n25559, n25560, n25561,
    n25562, n25563, n25564, n25565, n25566, n25567,
    n25568, n25569, n25570, n25571, n25572, n25573,
    n25574, n25575, n25576, n25577, n25578, n25579,
    n25580, n25581, n25582, n25583, n25584, n25585,
    n25586, n25587, n25588, n25589, n25590, n25591,
    n25592, n25593, n25594, n25595, n25596, n25597,
    n25598, n25599, n25600, n25601, n25602, n25603,
    n25604, n25605, n25606, n25607, n25608, n25609,
    n25610, n25611, n25612, n25613, n25614, n25615,
    n25616, n25617, n25618, n25619, n25620, n25621,
    n25622, n25623, n25624, n25625, n25626, n25627,
    n25628, n25629, n25630, n25631, n25632, n25633,
    n25634, n25635, n25636, n25637, n25638, n25639,
    n25640, n25641, n25642, n25643, n25644, n25645,
    n25646, n25647, n25648, n25649, n25650, n25651,
    n25652, n25653, n25654, n25655, n25656, n25657,
    n25658, n25659, n25660, n25661, n25662, n25663,
    n25664, n25665, n25666, n25667, n25668, n25669,
    n25670, n25671, n25672, n25673, n25674, n25675,
    n25676, n25677, n25678, n25679, n25680, n25681,
    n25682, n25683, n25684, n25685, n25686, n25687,
    n25688, n25689, n25690, n25691, n25692, n25693,
    n25694, n25695, n25696, n25697, n25698, n25699,
    n25700, n25701, n25702, n25703, n25704, n25705,
    n25706, n25707, n25708, n25709, n25710, n25711,
    n25712, n25713, n25714, n25715, n25716, n25717,
    n25718, n25719, n25720, n25721, n25722, n25723,
    n25724, n25725, n25726, n25727, n25728, n25729,
    n25730, n25731, n25732, n25733, n25734, n25735,
    n25736, n25737, n25738, n25739, n25740, n25741,
    n25742, n25743, n25744, n25745, n25746, n25747,
    n25748, n25749, n25750, n25751, n25752, n25753,
    n25754, n25755, n25756, n25757, n25758, n25759,
    n25760, n25761, n25762, n25763, n25764, n25765,
    n25766, n25767, n25768, n25769, n25770, n25771,
    n25772, n25773, n25774, n25775, n25776, n25777,
    n25778, n25779, n25780, n25781, n25782, n25783,
    n25784, n25785, n25786, n25787, n25788, n25789,
    n25790, n25791, n25792, n25793, n25794, n25795,
    n25796, n25797, n25798, n25799, n25800, n25801,
    n25802, n25803, n25804, n25805, n25806, n25807,
    n25808, n25809, n25810, n25811, n25812, n25813,
    n25814, n25815, n25816, n25817, n25818, n25819,
    n25820, n25821, n25822, n25823, n25824, n25825,
    n25826, n25827, n25828, n25829, n25830, n25831,
    n25832, n25833, n25834, n25835, n25836, n25837,
    n25838, n25839, n25840, n25841, n25842, n25843,
    n25844, n25845, n25846, n25847, n25848, n25849,
    n25850, n25851, n25852, n25853, n25854, n25855,
    n25856, n25857, n25858, n25859, n25860, n25861,
    n25862, n25863, n25864, n25865, n25866, n25867,
    n25868, n25869, n25870, n25871, n25872, n25873,
    n25874, n25875, n25876, n25878, n25879, n25880,
    n25881, n25882, n25883, n25884, n25885, n25886,
    n25887, n25888, n25889, n25890, n25891, n25892,
    n25893, n25894, n25895, n25896, n25897, n25898,
    n25899, n25900, n25901, n25902, n25903, n25904,
    n25905, n25906, n25907, n25908, n25909, n25910,
    n25911, n25912, n25913, n25914, n25915, n25916,
    n25917, n25918, n25919, n25920, n25921, n25922,
    n25923, n25924, n25925, n25926, n25927, n25928,
    n25929, n25930, n25931, n25932, n25933, n25934,
    n25935, n25936, n25937, n25938, n25939, n25940,
    n25941, n25942, n25943, n25944, n25945, n25946,
    n25947, n25948, n25949, n25950, n25951, n25952,
    n25953, n25954, n25955, n25956, n25957, n25958,
    n25959, n25960, n25961, n25962, n25963, n25964,
    n25965, n25966, n25967, n25968, n25969, n25970,
    n25971, n25972, n25973, n25974, n25975, n25976,
    n25977, n25978, n25979, n25980, n25981, n25982,
    n25983, n25984, n25985, n25986, n25987, n25988,
    n25989, n25990, n25991, n25992, n25993, n25994,
    n25995, n25996, n25997, n25998, n25999, n26000,
    n26001, n26002, n26003, n26004, n26005, n26006,
    n26007, n26008, n26009, n26010, n26011, n26012,
    n26013, n26014, n26015, n26016, n26017, n26018,
    n26019, n26020, n26021, n26022, n26023, n26024,
    n26025, n26026, n26027, n26028, n26029, n26030,
    n26031, n26032, n26033, n26034, n26035, n26036,
    n26037, n26038, n26039, n26040, n26041, n26042,
    n26043, n26044, n26045, n26046, n26047, n26048,
    n26049, n26050, n26051, n26052, n26053, n26054,
    n26055, n26056, n26057, n26058, n26059, n26060,
    n26061, n26062, n26063, n26064, n26065, n26066,
    n26067, n26068, n26069, n26070, n26071, n26072,
    n26073, n26074, n26075, n26076, n26077, n26078,
    n26079, n26080, n26081, n26082, n26083, n26084,
    n26085, n26086, n26087, n26088, n26089, n26090,
    n26091, n26092, n26093, n26094, n26095, n26096,
    n26097, n26098, n26099, n26100, n26101, n26102,
    n26103, n26104, n26105, n26106, n26107, n26108,
    n26109, n26110, n26111, n26112, n26113, n26114,
    n26115, n26116, n26117, n26118, n26119, n26120,
    n26121, n26122, n26123, n26124, n26125, n26126,
    n26127, n26128, n26129, n26130, n26131, n26132,
    n26133, n26134, n26135, n26136, n26137, n26138,
    n26139, n26140, n26141, n26142, n26143, n26144,
    n26145, n26146, n26147, n26148, n26149, n26150,
    n26151, n26152, n26153, n26154, n26155, n26156,
    n26157, n26158, n26159, n26160, n26161, n26162,
    n26163, n26164, n26165, n26166, n26167, n26168,
    n26169, n26170, n26171, n26172, n26173, n26174,
    n26175, n26176, n26177, n26178, n26179, n26180,
    n26181, n26182, n26183, n26184, n26185, n26186,
    n26187, n26188, n26189, n26190, n26191, n26192,
    n26193, n26194, n26195, n26196, n26197, n26198,
    n26199, n26200, n26201, n26202, n26203, n26204,
    n26205, n26206, n26207, n26208, n26209, n26210,
    n26211, n26212, n26213, n26214, n26215, n26216,
    n26217, n26218, n26219, n26220, n26221, n26222,
    n26223, n26224, n26225, n26226, n26227, n26228,
    n26229, n26230, n26231, n26232, n26233, n26234,
    n26235, n26236, n26237, n26238, n26239, n26240,
    n26241, n26242, n26243, n26244, n26245, n26246,
    n26247, n26248, n26249, n26250, n26251, n26252,
    n26253, n26254, n26255, n26256, n26257, n26258,
    n26259, n26260, n26261, n26262, n26263, n26264,
    n26265, n26266, n26267, n26268, n26269, n26270,
    n26271, n26272, n26273, n26274, n26275, n26276,
    n26277, n26278, n26279, n26280, n26281, n26282,
    n26283, n26284, n26285, n26286, n26287, n26288,
    n26289, n26290, n26291, n26292, n26293, n26294,
    n26295, n26296, n26297, n26298, n26299, n26300,
    n26301, n26302, n26303, n26304, n26305, n26306,
    n26307, n26308, n26309, n26310, n26311, n26312,
    n26313, n26314, n26315, n26316, n26317, n26318,
    n26319, n26320, n26321, n26322, n26323, n26324,
    n26325, n26326, n26327, n26328, n26329, n26330,
    n26331, n26332, n26333, n26334, n26335, n26336,
    n26337, n26338, n26339, n26340, n26341, n26342,
    n26343, n26344, n26345, n26346, n26347, n26348,
    n26349, n26351, n26352, n26353, n26354, n26355,
    n26356, n26357, n26358, n26359, n26360, n26361,
    n26362, n26363, n26364, n26365, n26366, n26367,
    n26368, n26369, n26370, n26371, n26372, n26373,
    n26374, n26375, n26376, n26377, n26378, n26379,
    n26380, n26381, n26382, n26383, n26384, n26385,
    n26386, n26387, n26388, n26389, n26390, n26391,
    n26392, n26393, n26394, n26395, n26396, n26397,
    n26398, n26399, n26400, n26401, n26402, n26403,
    n26404, n26405, n26406, n26407, n26408, n26409,
    n26410, n26411, n26412, n26413, n26414, n26415,
    n26416, n26417, n26418, n26419, n26420, n26421,
    n26422, n26423, n26424, n26425, n26426, n26427,
    n26428, n26429, n26430, n26431, n26432, n26433,
    n26434, n26435, n26436, n26437, n26438, n26439,
    n26440, n26441, n26442, n26443, n26444, n26445,
    n26446, n26447, n26448, n26449, n26450, n26451,
    n26452, n26453, n26454, n26455, n26456, n26457,
    n26458, n26459, n26460, n26461, n26462, n26463,
    n26464, n26465, n26466, n26467, n26468, n26469,
    n26470, n26471, n26472, n26473, n26474, n26475,
    n26476, n26477, n26478, n26479, n26480, n26481,
    n26482, n26483, n26484, n26485, n26486, n26487,
    n26488, n26489, n26490, n26491, n26492, n26493,
    n26494, n26495, n26496, n26497, n26498, n26499,
    n26500, n26501, n26502, n26503, n26504, n26505,
    n26506, n26507, n26508, n26509, n26510, n26511,
    n26512, n26513, n26514, n26515, n26516, n26517,
    n26518, n26519, n26520, n26521, n26522, n26523,
    n26524, n26525, n26526, n26527, n26528, n26529,
    n26530, n26531, n26532, n26533, n26534, n26535,
    n26536, n26537, n26538, n26539, n26540, n26541,
    n26542, n26543, n26544, n26545, n26546, n26547,
    n26548, n26549, n26550, n26551, n26552, n26553,
    n26554, n26555, n26556, n26557, n26558, n26559,
    n26560, n26561, n26562, n26563, n26564, n26565,
    n26566, n26567, n26568, n26569, n26570, n26571,
    n26572, n26573, n26574, n26575, n26576, n26577,
    n26578, n26579, n26580, n26581, n26582, n26583,
    n26584, n26585, n26586, n26587, n26588, n26589,
    n26590, n26591, n26592, n26593, n26594, n26595,
    n26596, n26597, n26598, n26599, n26600, n26601,
    n26602, n26603, n26604, n26605, n26606, n26607,
    n26608, n26609, n26610, n26611, n26612, n26613,
    n26614, n26615, n26616, n26617, n26618, n26619,
    n26620, n26621, n26622, n26623, n26624, n26625,
    n26626, n26627, n26628, n26629, n26630, n26631,
    n26632, n26633, n26634, n26635, n26636, n26637,
    n26638, n26639, n26640, n26641, n26642, n26643,
    n26644, n26645, n26646, n26647, n26648, n26649,
    n26650, n26651, n26652, n26653, n26654, n26655,
    n26656, n26657, n26658, n26659, n26660, n26661,
    n26662, n26663, n26664, n26665, n26666, n26667,
    n26668, n26669, n26670, n26671, n26672, n26673,
    n26674, n26675, n26676, n26677, n26678, n26679,
    n26680, n26681, n26682, n26683, n26684, n26685,
    n26686, n26687, n26688, n26689, n26690, n26691,
    n26692, n26693, n26694, n26695, n26696, n26697,
    n26698, n26699, n26700, n26701, n26702, n26703,
    n26704, n26705, n26706, n26707, n26708, n26709,
    n26710, n26711, n26712, n26713, n26714, n26715,
    n26716, n26717, n26718, n26719, n26720, n26721,
    n26722, n26723, n26724, n26725, n26726, n26727,
    n26728, n26729, n26730, n26731, n26732, n26733,
    n26734, n26735, n26736, n26737, n26738, n26739,
    n26740, n26741, n26742, n26743, n26744, n26745,
    n26746, n26747, n26748, n26749, n26750, n26751,
    n26752, n26753, n26754, n26755, n26756, n26757,
    n26758, n26759, n26760, n26761, n26762, n26763,
    n26764, n26765, n26766, n26767, n26768, n26769,
    n26770, n26771, n26772, n26773, n26774, n26775,
    n26776, n26777, n26778, n26779, n26780, n26781,
    n26782, n26783, n26784, n26785, n26786, n26787,
    n26788, n26789, n26790, n26791, n26792, n26793,
    n26794, n26795, n26796, n26797, n26798, n26799,
    n26800, n26801, n26802, n26803, n26804, n26805,
    n26806, n26807, n26808, n26809, n26810, n26811,
    n26812, n26813, n26814, n26815, n26816, n26818,
    n26819, n26820, n26821, n26822, n26823, n26824,
    n26825, n26826, n26827, n26828, n26829, n26830,
    n26831, n26832, n26833, n26834, n26835, n26836,
    n26837, n26838, n26839, n26840, n26841, n26842,
    n26843, n26844, n26845, n26846, n26847, n26848,
    n26849, n26850, n26851, n26852, n26853, n26854,
    n26855, n26856, n26857, n26858, n26859, n26860,
    n26861, n26862, n26863, n26864, n26865, n26866,
    n26867, n26868, n26869, n26870, n26871, n26872,
    n26873, n26874, n26875, n26876, n26877, n26878,
    n26879, n26880, n26881, n26882, n26883, n26884,
    n26885, n26886, n26887, n26888, n26889, n26890,
    n26891, n26892, n26893, n26894, n26895, n26896,
    n26897, n26898, n26899, n26900, n26901, n26902,
    n26903, n26904, n26905, n26906, n26907, n26908,
    n26909, n26910, n26911, n26912, n26913, n26914,
    n26915, n26916, n26917, n26918, n26919, n26920,
    n26921, n26922, n26923, n26924, n26925, n26926,
    n26927, n26928, n26929, n26930, n26931, n26932,
    n26933, n26934, n26935, n26936, n26937, n26938,
    n26939, n26940, n26941, n26942, n26943, n26944,
    n26945, n26946, n26947, n26948, n26949, n26950,
    n26951, n26952, n26953, n26954, n26955, n26956,
    n26957, n26958, n26959, n26960, n26961, n26962,
    n26963, n26964, n26965, n26966, n26967, n26968,
    n26969, n26970, n26971, n26972, n26973, n26974,
    n26975, n26976, n26977, n26978, n26979, n26980,
    n26981, n26982, n26983, n26984, n26985, n26986,
    n26987, n26988, n26989, n26990, n26991, n26992,
    n26993, n26994, n26995, n26996, n26997, n26998,
    n26999, n27000, n27001, n27002, n27003, n27004,
    n27005, n27006, n27007, n27008, n27009, n27010,
    n27011, n27012, n27013, n27014, n27015, n27016,
    n27017, n27018, n27019, n27020, n27021, n27022,
    n27023, n27024, n27025, n27026, n27027, n27028,
    n27029, n27030, n27031, n27032, n27033, n27034,
    n27035, n27036, n27037, n27038, n27039, n27040,
    n27041, n27042, n27043, n27044, n27045, n27046,
    n27047, n27048, n27049, n27050, n27051, n27052,
    n27053, n27054, n27055, n27056, n27057, n27058,
    n27059, n27060, n27061, n27062, n27063, n27064,
    n27065, n27066, n27067, n27068, n27069, n27070,
    n27071, n27072, n27073, n27074, n27075, n27076,
    n27077, n27078, n27079, n27080, n27081, n27082,
    n27083, n27084, n27085, n27086, n27087, n27088,
    n27089, n27090, n27091, n27092, n27093, n27094,
    n27095, n27096, n27097, n27098, n27099, n27100,
    n27101, n27102, n27103, n27104, n27105, n27106,
    n27107, n27108, n27109, n27110, n27111, n27112,
    n27113, n27114, n27115, n27116, n27117, n27118,
    n27119, n27120, n27121, n27122, n27123, n27124,
    n27125, n27126, n27127, n27128, n27129, n27130,
    n27131, n27132, n27133, n27134, n27135, n27136,
    n27137, n27138, n27139, n27140, n27141, n27142,
    n27143, n27144, n27145, n27146, n27147, n27148,
    n27149, n27150, n27151, n27152, n27153, n27154,
    n27155, n27156, n27157, n27158, n27159, n27160,
    n27161, n27162, n27163, n27164, n27165, n27166,
    n27167, n27168, n27169, n27170, n27171, n27172,
    n27173, n27174, n27175, n27176, n27177, n27178,
    n27179, n27180, n27181, n27182, n27183, n27184,
    n27185, n27186, n27187, n27188, n27189, n27190,
    n27191, n27192, n27193, n27194, n27195, n27196,
    n27197, n27198, n27199, n27200, n27201, n27202,
    n27203, n27204, n27205, n27206, n27207, n27208,
    n27209, n27210, n27211, n27212, n27213, n27214,
    n27215, n27216, n27217, n27218, n27219, n27220,
    n27221, n27222, n27223, n27224, n27225, n27226,
    n27227, n27228, n27229, n27230, n27231, n27232,
    n27233, n27234, n27235, n27236, n27237, n27238,
    n27239, n27240, n27241, n27242, n27243, n27244,
    n27245, n27246, n27247, n27248, n27249, n27250,
    n27251, n27252, n27253, n27254, n27255, n27256,
    n27257, n27258, n27259, n27260, n27261, n27262,
    n27263, n27264, n27265, n27266, n27267, n27268,
    n27269, n27270, n27271, n27272, n27273, n27274,
    n27275, n27276, n27277, n27278, n27279, n27280,
    n27281, n27282, n27283, n27285, n27286, n27287,
    n27288, n27289, n27290, n27291, n27292, n27293,
    n27294, n27295, n27296, n27297, n27298, n27299,
    n27300, n27301, n27302, n27303, n27304, n27305,
    n27306, n27307, n27308, n27309, n27310, n27311,
    n27312, n27313, n27314, n27315, n27316, n27317,
    n27318, n27319, n27320, n27321, n27322, n27323,
    n27324, n27325, n27326, n27327, n27328, n27329,
    n27330, n27331, n27332, n27333, n27334, n27335,
    n27336, n27337, n27338, n27339, n27340, n27341,
    n27342, n27343, n27344, n27345, n27346, n27347,
    n27348, n27349, n27350, n27351, n27352, n27353,
    n27354, n27355, n27356, n27357, n27358, n27359,
    n27360, n27361, n27362, n27363, n27364, n27365,
    n27366, n27367, n27368, n27369, n27370, n27371,
    n27372, n27373, n27374, n27375, n27376, n27377,
    n27378, n27379, n27380, n27381, n27382, n27383,
    n27384, n27385, n27386, n27387, n27388, n27389,
    n27390, n27391, n27392, n27393, n27394, n27395,
    n27396, n27397, n27398, n27399, n27400, n27401,
    n27402, n27403, n27404, n27405, n27406, n27407,
    n27408, n27409, n27410, n27411, n27412, n27413,
    n27414, n27415, n27416, n27417, n27418, n27419,
    n27420, n27421, n27422, n27423, n27424, n27425,
    n27426, n27427, n27428, n27429, n27430, n27431,
    n27432, n27433, n27434, n27435, n27436, n27437,
    n27438, n27439, n27440, n27441, n27442, n27443,
    n27444, n27445, n27446, n27447, n27448, n27449,
    n27450, n27451, n27452, n27453, n27454, n27455,
    n27456, n27457, n27458, n27459, n27460, n27461,
    n27462, n27463, n27464, n27465, n27466, n27467,
    n27468, n27469, n27470, n27471, n27472, n27473,
    n27474, n27475, n27476, n27477, n27478, n27479,
    n27480, n27481, n27482, n27483, n27484, n27485,
    n27486, n27487, n27488, n27489, n27490, n27491,
    n27492, n27493, n27494, n27495, n27496, n27497,
    n27498, n27499, n27500, n27501, n27502, n27503,
    n27504, n27505, n27506, n27507, n27508, n27509,
    n27510, n27511, n27512, n27513, n27514, n27515,
    n27516, n27517, n27518, n27519, n27520, n27521,
    n27522, n27523, n27524, n27525, n27526, n27527,
    n27528, n27529, n27530, n27531, n27532, n27533,
    n27534, n27535, n27536, n27537, n27538, n27539,
    n27540, n27541, n27542, n27543, n27544, n27545,
    n27546, n27547, n27548, n27549, n27550, n27551,
    n27552, n27553, n27554, n27555, n27556, n27557,
    n27558, n27559, n27560, n27561, n27562, n27563,
    n27564, n27565, n27566, n27567, n27568, n27569,
    n27570, n27571, n27572, n27573, n27574, n27575,
    n27576, n27577, n27578, n27579, n27580, n27581,
    n27582, n27583, n27584, n27585, n27586, n27587,
    n27588, n27589, n27590, n27591, n27592, n27593,
    n27594, n27595, n27596, n27597, n27598, n27599,
    n27600, n27601, n27602, n27603, n27604, n27605,
    n27606, n27607, n27608, n27609, n27610, n27611,
    n27612, n27613, n27614, n27615, n27616, n27617,
    n27618, n27619, n27620, n27621, n27622, n27623,
    n27624, n27625, n27626, n27627, n27628, n27629,
    n27630, n27631, n27632, n27633, n27634, n27635,
    n27636, n27637, n27638, n27639, n27640, n27641,
    n27642, n27643, n27644, n27645, n27646, n27647,
    n27648, n27649, n27650, n27651, n27652, n27653,
    n27654, n27655, n27656, n27657, n27658, n27659,
    n27660, n27661, n27662, n27663, n27664, n27665,
    n27666, n27667, n27668, n27669, n27670, n27671,
    n27672, n27673, n27674, n27675, n27676, n27677,
    n27678, n27679, n27680, n27681, n27682, n27683,
    n27684, n27685, n27686, n27687, n27688, n27689,
    n27690, n27691, n27692, n27693, n27694, n27695,
    n27696, n27697, n27698, n27699, n27700, n27701,
    n27702, n27703, n27704, n27705, n27706, n27707,
    n27708, n27709, n27710, n27711, n27712, n27713,
    n27714, n27715, n27716, n27717, n27718, n27719,
    n27720, n27721, n27722, n27723, n27724, n27725,
    n27726, n27727, n27728, n27729, n27730, n27731,
    n27732, n27733, n27734, n27735, n27736, n27737,
    n27738, n27739, n27740, n27741, n27742, n27743,
    n27744, n27745, n27746, n27747, n27748, n27749,
    n27750, n27752, n27753, n27754, n27755, n27756,
    n27757, n27758, n27759, n27760, n27761, n27762,
    n27763, n27764, n27765, n27766, n27767, n27768,
    n27769, n27770, n27771, n27772, n27773, n27774,
    n27775, n27776, n27777, n27778, n27779, n27780,
    n27781, n27782, n27783, n27784, n27785, n27786,
    n27787, n27788, n27789, n27790, n27791, n27792,
    n27793, n27794, n27795, n27796, n27797, n27798,
    n27799, n27800, n27801, n27802, n27803, n27804,
    n27805, n27806, n27807, n27808, n27809, n27810,
    n27811, n27812, n27813, n27814, n27815, n27816,
    n27817, n27818, n27819, n27820, n27821, n27822,
    n27823, n27824, n27825, n27826, n27827, n27828,
    n27829, n27830, n27831, n27832, n27833, n27834,
    n27835, n27836, n27837, n27838, n27839, n27840,
    n27841, n27842, n27843, n27844, n27845, n27846,
    n27847, n27848, n27849, n27850, n27851, n27852,
    n27853, n27854, n27855, n27856, n27857, n27858,
    n27859, n27860, n27861, n27862, n27863, n27864,
    n27865, n27866, n27867, n27868, n27869, n27870,
    n27871, n27872, n27873, n27874, n27875, n27876,
    n27877, n27878, n27879, n27880, n27881, n27882,
    n27883, n27884, n27885, n27886, n27887, n27888,
    n27889, n27890, n27891, n27892, n27893, n27894,
    n27895, n27896, n27897, n27898, n27899, n27900,
    n27901, n27902, n27903, n27904, n27905, n27906,
    n27907, n27908, n27909, n27910, n27911, n27912,
    n27913, n27914, n27915, n27916, n27917, n27918,
    n27919, n27920, n27921, n27922, n27923, n27924,
    n27925, n27926, n27927, n27928, n27929, n27930,
    n27931, n27932, n27933, n27934, n27935, n27936,
    n27937, n27938, n27939, n27940, n27941, n27942,
    n27943, n27944, n27945, n27946, n27947, n27948,
    n27949, n27950, n27951, n27952, n27953, n27954,
    n27955, n27956, n27957, n27958, n27959, n27960,
    n27961, n27962, n27963, n27964, n27965, n27966,
    n27967, n27968, n27969, n27970, n27971, n27972,
    n27973, n27974, n27975, n27976, n27977, n27978,
    n27979, n27980, n27981, n27982, n27983, n27984,
    n27985, n27986, n27987, n27988, n27989, n27990,
    n27991, n27992, n27993, n27994, n27995, n27996,
    n27997, n27998, n27999, n28000, n28001, n28002,
    n28003, n28004, n28005, n28006, n28007, n28008,
    n28009, n28010, n28011, n28012, n28013, n28014,
    n28015, n28016, n28017, n28018, n28019, n28020,
    n28021, n28022, n28023, n28024, n28025, n28026,
    n28027, n28028, n28029, n28030, n28031, n28032,
    n28033, n28034, n28035, n28036, n28037, n28038,
    n28039, n28040, n28041, n28042, n28043, n28044,
    n28045, n28046, n28047, n28048, n28049, n28050,
    n28051, n28052, n28053, n28054, n28055, n28056,
    n28057, n28058, n28059, n28060, n28061, n28062,
    n28063, n28064, n28065, n28066, n28067, n28068,
    n28069, n28070, n28071, n28072, n28073, n28074,
    n28075, n28076, n28077, n28078, n28079, n28080,
    n28081, n28082, n28083, n28084, n28085, n28086,
    n28087, n28088, n28089, n28090, n28091, n28092,
    n28093, n28094, n28095, n28096, n28097, n28098,
    n28099, n28100, n28101, n28102, n28103, n28104,
    n28105, n28106, n28107, n28108, n28109, n28110,
    n28111, n28112, n28113, n28114, n28115, n28116,
    n28117, n28118, n28119, n28120, n28121, n28122,
    n28123, n28124, n28125, n28126, n28127, n28128,
    n28129, n28130, n28131, n28132, n28133, n28134,
    n28135, n28136, n28137, n28138, n28139, n28140,
    n28141, n28142, n28143, n28144, n28145, n28146,
    n28147, n28148, n28149, n28150, n28151, n28152,
    n28153, n28154, n28155, n28156, n28157, n28158,
    n28159, n28160, n28161, n28162, n28163, n28164,
    n28165, n28166, n28167, n28168, n28169, n28170,
    n28171, n28172, n28173, n28174, n28175, n28176,
    n28177, n28178, n28179, n28180, n28181, n28182,
    n28183, n28184, n28185, n28186, n28187, n28188,
    n28189, n28190, n28191, n28192, n28193, n28194,
    n28195, n28196, n28197, n28198, n28199, n28200,
    n28201, n28202, n28203, n28204, n28205, n28206,
    n28207, n28208, n28209, n28210, n28211, n28212,
    n28213, n28214, n28215, n28216, n28217, n28218,
    n28219, n28220, n28221, n28222, n28223, n28225,
    n28226, n28227, n28228, n28229, n28230, n28231,
    n28232, n28233, n28234, n28235, n28236, n28237,
    n28238, n28239, n28240, n28241, n28242, n28243,
    n28244, n28245, n28246, n28247, n28248, n28249,
    n28250, n28251, n28252, n28253, n28254, n28255,
    n28256, n28257, n28258, n28259, n28260, n28261,
    n28262, n28263, n28264, n28265, n28266, n28267,
    n28268, n28269, n28270, n28271, n28272, n28273,
    n28274, n28275, n28276, n28277, n28278, n28279,
    n28280, n28281, n28282, n28283, n28284, n28285,
    n28286, n28287, n28288, n28289, n28290, n28291,
    n28292, n28293, n28294, n28295, n28296, n28297,
    n28298, n28299, n28300, n28301, n28302, n28303,
    n28304, n28305, n28306, n28307, n28308, n28309,
    n28310, n28311, n28312, n28313, n28314, n28315,
    n28316, n28317, n28318, n28319, n28320, n28321,
    n28322, n28323, n28324, n28325, n28326, n28327,
    n28328, n28329, n28330, n28331, n28332, n28333,
    n28334, n28335, n28336, n28337, n28338, n28339,
    n28340, n28341, n28342, n28343, n28344, n28345,
    n28346, n28347, n28348, n28349, n28350, n28351,
    n28352, n28353, n28354, n28355, n28356, n28357,
    n28358, n28359, n28360, n28361, n28362, n28363,
    n28364, n28365, n28366, n28367, n28368, n28369,
    n28370, n28371, n28372, n28373, n28374, n28375,
    n28376, n28377, n28378, n28379, n28380, n28381,
    n28382, n28383, n28384, n28385, n28386, n28387,
    n28388, n28389, n28390, n28391, n28392, n28393,
    n28394, n28395, n28396, n28397, n28398, n28399,
    n28400, n28401, n28402, n28403, n28404, n28405,
    n28406, n28407, n28408, n28409, n28410, n28411,
    n28412, n28413, n28414, n28415, n28416, n28417,
    n28418, n28419, n28420, n28421, n28422, n28423,
    n28424, n28425, n28426, n28427, n28428, n28429,
    n28430, n28431, n28432, n28433, n28434, n28435,
    n28436, n28437, n28438, n28439, n28440, n28441,
    n28442, n28443, n28444, n28445, n28446, n28447,
    n28448, n28449, n28450, n28451, n28452, n28453,
    n28454, n28455, n28456, n28457, n28458, n28459,
    n28460, n28461, n28462, n28463, n28464, n28465,
    n28466, n28467, n28468, n28469, n28470, n28471,
    n28472, n28473, n28474, n28475, n28476, n28477,
    n28478, n28479, n28480, n28481, n28482, n28483,
    n28484, n28485, n28486, n28487, n28488, n28489,
    n28490, n28491, n28492, n28493, n28494, n28495,
    n28496, n28497, n28498, n28499, n28500, n28501,
    n28502, n28503, n28504, n28505, n28506, n28507,
    n28508, n28509, n28510, n28511, n28512, n28513,
    n28514, n28515, n28516, n28517, n28518, n28519,
    n28520, n28521, n28522, n28523, n28524, n28525,
    n28526, n28527, n28528, n28529, n28530, n28531,
    n28532, n28533, n28534, n28535, n28536, n28537,
    n28538, n28539, n28540, n28541, n28542, n28543,
    n28544, n28545, n28546, n28547, n28548, n28549,
    n28550, n28551, n28552, n28553, n28554, n28555,
    n28556, n28557, n28558, n28559, n28560, n28561,
    n28562, n28563, n28564, n28565, n28566, n28567,
    n28568, n28569, n28570, n28571, n28572, n28573,
    n28574, n28575, n28576, n28577, n28578, n28579,
    n28580, n28581, n28582, n28583, n28584, n28585,
    n28586, n28587, n28588, n28589, n28590, n28591,
    n28592, n28593, n28594, n28595, n28596, n28597,
    n28598, n28599, n28600, n28601, n28602, n28603,
    n28604, n28605, n28606, n28607, n28608, n28609,
    n28610, n28611, n28612, n28613, n28614, n28615,
    n28616, n28617, n28618, n28619, n28620, n28621,
    n28622, n28623, n28624, n28625, n28626, n28627,
    n28628, n28629, n28630, n28631, n28632, n28633,
    n28634, n28635, n28636, n28637, n28638, n28639,
    n28640, n28641, n28642, n28643, n28644, n28645,
    n28646, n28647, n28648, n28649, n28650, n28651,
    n28652, n28653, n28654, n28655, n28656, n28657,
    n28658, n28659, n28660, n28661, n28662, n28663,
    n28664, n28665, n28666, n28667, n28668, n28669,
    n28670, n28671, n28672, n28673, n28674, n28675,
    n28676, n28677, n28678, n28679, n28680, n28681,
    n28682, n28683, n28684, n28685, n28686, n28687,
    n28688, n28689, n28690, n28691, n28692, n28693,
    n28694, n28695, n28696, n28698, n28699, n28700,
    n28701, n28702, n28703, n28704, n28705, n28706,
    n28707, n28708, n28709, n28710, n28711, n28712,
    n28713, n28714, n28715, n28716, n28717, n28718,
    n28719, n28720, n28721, n28722, n28723, n28724,
    n28725, n28726, n28727, n28728, n28729, n28730,
    n28731, n28732, n28733, n28734, n28735, n28736,
    n28737, n28738, n28739, n28740, n28741, n28742,
    n28743, n28744, n28745, n28746, n28747, n28748,
    n28749, n28750, n28751, n28752, n28753, n28754,
    n28755, n28756, n28757, n28758, n28759, n28760,
    n28761, n28762, n28763, n28764, n28765, n28766,
    n28767, n28768, n28769, n28770, n28771, n28772,
    n28773, n28774, n28775, n28776, n28777, n28778,
    n28779, n28780, n28781, n28782, n28783, n28784,
    n28785, n28786, n28787, n28788, n28789, n28790,
    n28791, n28792, n28793, n28794, n28795, n28796,
    n28797, n28798, n28799, n28800, n28801, n28802,
    n28803, n28804, n28805, n28806, n28807, n28808,
    n28809, n28810, n28811, n28812, n28813, n28814,
    n28815, n28816, n28817, n28818, n28819, n28820,
    n28821, n28822, n28823, n28824, n28825, n28826,
    n28827, n28828, n28829, n28830, n28831, n28832,
    n28833, n28834, n28835, n28836, n28837, n28838,
    n28839, n28840, n28841, n28842, n28843, n28844,
    n28845, n28846, n28847, n28848, n28849, n28850,
    n28851, n28852, n28853, n28854, n28855, n28856,
    n28857, n28858, n28859, n28860, n28861, n28862,
    n28863, n28864, n28865, n28866, n28867, n28868,
    n28869, n28870, n28871, n28872, n28873, n28874,
    n28875, n28876, n28877, n28878, n28879, n28880,
    n28881, n28882, n28883, n28884, n28885, n28886,
    n28887, n28888, n28889, n28890, n28891, n28892,
    n28893, n28894, n28895, n28896, n28897, n28898,
    n28899, n28900, n28901, n28902, n28903, n28904,
    n28905, n28906, n28907, n28908, n28909, n28910,
    n28911, n28912, n28913, n28914, n28915, n28916,
    n28917, n28918, n28919, n28920, n28921, n28922,
    n28923, n28924, n28925, n28926, n28927, n28928,
    n28929, n28930, n28931, n28932, n28933, n28934,
    n28935, n28936, n28937, n28938, n28939, n28940,
    n28941, n28942, n28943, n28944, n28945, n28946,
    n28947, n28948, n28949, n28950, n28951, n28952,
    n28953, n28954, n28955, n28956, n28957, n28958,
    n28959, n28960, n28961, n28962, n28963, n28964,
    n28965, n28966, n28967, n28968, n28969, n28970,
    n28971, n28972, n28973, n28974, n28975, n28976,
    n28977, n28978, n28979, n28980, n28981, n28982,
    n28983, n28984, n28985, n28986, n28987, n28988,
    n28989, n28990, n28991, n28992, n28993, n28994,
    n28995, n28996, n28997, n28998, n28999, n29000,
    n29001, n29002, n29003, n29004, n29005, n29006,
    n29007, n29008, n29009, n29010, n29011, n29012,
    n29013, n29014, n29015, n29016, n29017, n29018,
    n29019, n29020, n29021, n29022, n29023, n29024,
    n29025, n29026, n29027, n29028, n29029, n29030,
    n29031, n29032, n29033, n29034, n29035, n29036,
    n29037, n29038, n29039, n29040, n29041, n29042,
    n29043, n29044, n29045, n29046, n29047, n29048,
    n29049, n29050, n29051, n29052, n29053, n29054,
    n29055, n29056, n29057, n29058, n29059, n29060,
    n29061, n29062, n29063, n29064, n29065, n29066,
    n29067, n29068, n29069, n29070, n29071, n29072,
    n29073, n29074, n29075, n29076, n29077, n29078,
    n29079, n29080, n29081, n29082, n29083, n29084,
    n29085, n29086, n29087, n29088, n29089, n29090,
    n29091, n29092, n29093, n29094, n29095, n29096,
    n29097, n29098, n29099, n29100, n29101, n29102,
    n29103, n29104, n29105, n29106, n29107, n29108,
    n29109, n29110, n29111, n29112, n29113, n29114,
    n29115, n29116, n29117, n29118, n29119, n29120,
    n29121, n29122, n29123, n29124, n29125, n29126,
    n29127, n29128, n29129, n29130, n29131, n29132,
    n29133, n29134, n29135, n29136, n29137, n29138,
    n29139, n29140, n29141, n29142, n29143, n29144,
    n29145, n29146, n29147, n29148, n29149, n29150,
    n29151, n29152, n29153, n29154, n29155, n29156,
    n29157, n29158, n29159, n29160, n29161, n29162,
    n29163, n29164, n29165, n29166, n29167, n29168,
    n29169, n29171, n29172, n29173, n29174, n29175,
    n29176, n29177, n29178, n29179, n29180, n29181,
    n29182, n29183, n29184, n29185, n29186, n29187,
    n29188, n29189, n29190, n29191, n29192, n29193,
    n29194, n29195, n29196, n29197, n29198, n29199,
    n29200, n29201, n29202, n29203, n29204, n29205,
    n29206, n29207, n29208, n29209, n29210, n29211,
    n29212, n29213, n29214, n29215, n29216, n29217,
    n29218, n29219, n29220, n29221, n29222, n29223,
    n29224, n29225, n29226, n29227, n29228, n29229,
    n29230, n29231, n29232, n29233, n29234, n29235,
    n29236, n29237, n29238, n29239, n29240, n29241,
    n29242, n29243, n29244, n29245, n29246, n29247,
    n29248, n29249, n29250, n29251, n29252, n29253,
    n29254, n29255, n29256, n29257, n29258, n29259,
    n29260, n29261, n29262, n29263, n29264, n29265,
    n29266, n29267, n29268, n29269, n29270, n29271,
    n29272, n29273, n29274, n29275, n29276, n29277,
    n29278, n29279, n29280, n29281, n29282, n29283,
    n29284, n29285, n29286, n29287, n29288, n29289,
    n29290, n29291, n29292, n29293, n29294, n29295,
    n29296, n29297, n29298, n29299, n29300, n29301,
    n29302, n29303, n29304, n29305, n29306, n29307,
    n29308, n29309, n29310, n29311, n29312, n29313,
    n29314, n29315, n29316, n29317, n29318, n29319,
    n29320, n29321, n29322, n29323, n29324, n29325,
    n29326, n29327, n29328, n29329, n29330, n29331,
    n29332, n29333, n29334, n29335, n29336, n29337,
    n29338, n29339, n29340, n29341, n29342, n29343,
    n29344, n29345, n29346, n29347, n29348, n29349,
    n29350, n29351, n29352, n29353, n29354, n29355,
    n29356, n29357, n29358, n29359, n29360, n29361,
    n29362, n29363, n29364, n29365, n29366, n29367,
    n29368, n29369, n29370, n29371, n29372, n29373,
    n29374, n29375, n29376, n29377, n29378, n29379,
    n29380, n29381, n29382, n29383, n29384, n29385,
    n29386, n29387, n29388, n29389, n29390, n29391,
    n29392, n29393, n29394, n29395, n29396, n29397,
    n29398, n29399, n29400, n29401, n29402, n29403,
    n29404, n29405, n29406, n29407, n29408, n29409,
    n29410, n29411, n29412, n29413, n29414, n29415,
    n29416, n29417, n29418, n29419, n29420, n29421,
    n29422, n29423, n29424, n29425, n29426, n29427,
    n29428, n29429, n29430, n29431, n29432, n29433,
    n29434, n29435, n29436, n29437, n29438, n29439,
    n29440, n29441, n29442, n29443, n29444, n29445,
    n29446, n29447, n29448, n29449, n29450, n29451,
    n29452, n29453, n29454, n29455, n29456, n29457,
    n29458, n29459, n29460, n29461, n29462, n29463,
    n29464, n29465, n29466, n29467, n29468, n29469,
    n29470, n29471, n29472, n29473, n29474, n29475,
    n29476, n29477, n29478, n29479, n29480, n29481,
    n29482, n29483, n29484, n29485, n29486, n29487,
    n29488, n29489, n29490, n29491, n29492, n29493,
    n29494, n29495, n29496, n29497, n29498, n29499,
    n29500, n29501, n29502, n29503, n29504, n29505,
    n29506, n29507, n29508, n29509, n29510, n29511,
    n29512, n29513, n29514, n29515, n29516, n29517,
    n29518, n29519, n29520, n29521, n29522, n29523,
    n29524, n29525, n29526, n29527, n29528, n29529,
    n29530, n29531, n29532, n29533, n29534, n29535,
    n29536, n29537, n29538, n29539, n29540, n29541,
    n29542, n29543, n29544, n29545, n29546, n29547,
    n29548, n29549, n29550, n29551, n29552, n29553,
    n29554, n29555, n29556, n29557, n29558, n29559,
    n29560, n29561, n29562, n29563, n29564, n29565,
    n29566, n29567, n29568, n29569, n29570, n29571,
    n29572, n29573, n29574, n29575, n29576, n29577,
    n29578, n29579, n29580, n29581, n29582, n29583,
    n29584, n29585, n29586, n29587, n29588, n29589,
    n29590, n29591, n29592, n29593, n29594, n29595,
    n29596, n29597, n29598, n29599, n29600, n29601,
    n29602, n29603, n29604, n29605, n29606, n29607,
    n29608, n29609, n29610, n29611, n29612, n29613,
    n29614, n29615, n29616, n29617, n29618, n29619,
    n29620, n29621, n29622, n29623, n29624, n29625,
    n29626, n29627, n29628, n29629, n29630, n29631,
    n29632, n29633, n29634, n29635, n29636, n29637,
    n29638, n29639, n29640, n29641, n29642, n29644,
    n29645, n29646, n29647, n29648, n29649, n29650,
    n29651, n29652, n29653, n29654, n29655, n29656,
    n29657, n29658, n29659, n29660, n29661, n29662,
    n29663, n29664, n29665, n29666, n29667, n29668,
    n29669, n29670, n29671, n29672, n29673, n29674,
    n29675, n29676, n29677, n29678, n29679, n29680,
    n29681, n29682, n29683, n29684, n29685, n29686,
    n29687, n29688, n29689, n29690, n29691, n29692,
    n29693, n29694, n29695, n29696, n29697, n29698,
    n29699, n29700, n29701, n29702, n29703, n29704,
    n29705, n29706, n29707, n29708, n29709, n29710,
    n29711, n29712, n29713, n29714, n29715, n29716,
    n29717, n29718, n29719, n29720, n29721, n29722,
    n29723, n29724, n29725, n29726, n29727, n29728,
    n29729, n29730, n29731, n29732, n29733, n29734,
    n29735, n29736, n29737, n29738, n29739, n29740,
    n29741, n29742, n29743, n29744, n29745, n29746,
    n29747, n29748, n29749, n29750, n29751, n29752,
    n29753, n29754, n29755, n29756, n29757, n29758,
    n29759, n29760, n29761, n29762, n29763, n29764,
    n29765, n29766, n29767, n29768, n29769, n29770,
    n29771, n29772, n29773, n29774, n29775, n29776,
    n29777, n29778, n29779, n29780, n29781, n29782,
    n29783, n29784, n29785, n29786, n29787, n29788,
    n29789, n29790, n29791, n29792, n29793, n29794,
    n29795, n29796, n29797, n29798, n29799, n29800,
    n29801, n29802, n29803, n29804, n29805, n29806,
    n29807, n29808, n29809, n29810, n29811, n29812,
    n29813, n29814, n29815, n29816, n29817, n29818,
    n29819, n29820, n29821, n29822, n29823, n29824,
    n29825, n29826, n29827, n29828, n29829, n29830,
    n29831, n29832, n29833, n29834, n29835, n29836,
    n29837, n29838, n29839, n29840, n29841, n29842,
    n29843, n29844, n29845, n29846, n29847, n29848,
    n29849, n29850, n29851, n29852, n29853, n29854,
    n29855, n29856, n29857, n29858, n29859, n29860,
    n29861, n29862, n29863, n29864, n29865, n29866,
    n29867, n29868, n29869, n29870, n29871, n29872,
    n29873, n29874, n29875, n29876, n29877, n29878,
    n29879, n29880, n29881, n29882, n29883, n29884,
    n29885, n29886, n29887, n29888, n29889, n29890,
    n29891, n29892, n29893, n29894, n29895, n29896,
    n29897, n29898, n29899, n29900, n29901, n29902,
    n29903, n29904, n29905, n29906, n29907, n29908,
    n29909, n29910, n29911, n29912, n29913, n29914,
    n29915, n29916, n29917, n29918, n29919, n29920,
    n29921, n29922, n29923, n29924, n29925, n29926,
    n29927, n29928, n29929, n29930, n29931, n29932,
    n29933, n29934, n29935, n29936, n29937, n29938,
    n29939, n29940, n29941, n29942, n29943, n29944,
    n29945, n29946, n29947, n29948, n29949, n29950,
    n29951, n29952, n29953, n29954, n29955, n29956,
    n29957, n29958, n29959, n29960, n29961, n29962,
    n29963, n29964, n29965, n29966, n29967, n29968,
    n29969, n29970, n29971, n29972, n29973, n29974,
    n29975, n29976, n29977, n29978, n29979, n29980,
    n29981, n29982, n29983, n29984, n29985, n29986,
    n29987, n29988, n29989, n29990, n29991, n29992,
    n29993, n29994, n29995, n29996, n29997, n29998,
    n29999, n30000, n30001, n30002, n30003, n30004,
    n30005, n30006, n30007, n30008, n30009, n30010,
    n30011, n30012, n30013, n30014, n30015, n30016,
    n30017, n30018, n30019, n30020, n30021, n30022,
    n30023, n30024, n30025, n30026, n30027, n30028,
    n30029, n30030, n30031, n30032, n30033, n30034,
    n30035, n30036, n30037, n30038, n30039, n30040,
    n30041, n30042, n30043, n30044, n30045, n30046,
    n30047, n30048, n30049, n30050, n30051, n30052,
    n30053, n30054, n30055, n30056, n30057, n30058,
    n30059, n30060, n30061, n30062, n30063, n30064,
    n30065, n30066, n30067, n30068, n30069, n30070,
    n30071, n30072, n30073, n30074, n30075, n30076,
    n30077, n30078, n30079, n30080, n30081, n30082,
    n30083, n30084, n30085, n30086, n30087, n30088,
    n30089, n30090, n30091, n30092, n30093, n30094,
    n30095, n30096, n30097, n30098, n30099, n30100,
    n30101, n30102, n30103, n30104, n30105, n30106,
    n30107, n30108, n30109, n30110, n30111, n30112,
    n30113, n30114, n30115, n30116, n30117, n30118,
    n30120, n30121, n30122, n30123, n30124, n30125,
    n30126, n30127, n30128, n30129, n30130, n30131,
    n30132, n30133, n30134, n30135, n30136, n30137,
    n30138, n30139, n30140, n30141, n30142, n30143,
    n30144, n30145, n30146, n30147, n30148, n30149,
    n30150, n30151, n30152, n30153, n30154, n30155,
    n30156, n30157, n30158, n30159, n30160, n30161,
    n30162, n30163, n30164, n30165, n30166, n30167,
    n30168, n30169, n30170, n30171, n30172, n30173,
    n30174, n30175, n30176, n30177, n30178, n30179,
    n30180, n30181, n30182, n30183, n30184, n30185,
    n30186, n30187, n30188, n30189, n30190, n30191,
    n30192, n30193, n30194, n30195, n30196, n30197,
    n30198, n30199, n30200, n30201, n30202, n30203,
    n30204, n30205, n30206, n30207, n30208, n30209,
    n30210, n30211, n30212, n30213, n30214, n30215,
    n30216, n30217, n30218, n30219, n30220, n30221,
    n30222, n30223, n30224, n30225, n30226, n30227,
    n30228, n30229, n30230, n30231, n30232, n30233,
    n30234, n30235, n30236, n30237, n30238, n30239,
    n30240, n30241, n30242, n30243, n30244, n30245,
    n30246, n30247, n30248, n30249, n30250, n30251,
    n30252, n30253, n30254, n30255, n30256, n30257,
    n30258, n30259, n30260, n30261, n30262, n30263,
    n30264, n30265, n30266, n30267, n30268, n30269,
    n30270, n30271, n30272, n30273, n30274, n30275,
    n30276, n30277, n30278, n30279, n30280, n30281,
    n30282, n30283, n30284, n30285, n30286, n30287,
    n30288, n30289, n30290, n30291, n30292, n30293,
    n30294, n30295, n30296, n30297, n30298, n30299,
    n30300, n30301, n30302, n30303, n30304, n30305,
    n30306, n30307, n30308, n30309, n30310, n30311,
    n30312, n30313, n30314, n30315, n30316, n30317,
    n30318, n30319, n30320, n30321, n30322, n30323,
    n30324, n30325, n30326, n30327, n30328, n30329,
    n30330, n30331, n30332, n30333, n30334, n30335,
    n30336, n30337, n30338, n30339, n30340, n30341,
    n30342, n30343, n30344, n30345, n30346, n30347,
    n30348, n30349, n30350, n30351, n30352, n30353,
    n30354, n30355, n30356, n30357, n30358, n30359,
    n30360, n30361, n30362, n30363, n30364, n30365,
    n30366, n30367, n30368, n30369, n30370, n30371,
    n30372, n30373, n30374, n30375, n30376, n30377,
    n30378, n30379, n30380, n30381, n30382, n30383,
    n30384, n30385, n30386, n30387, n30388, n30389,
    n30390, n30391, n30392, n30393, n30394, n30395,
    n30396, n30397, n30398, n30399, n30400, n30401,
    n30402, n30403, n30404, n30405, n30406, n30407,
    n30408, n30409, n30410, n30411, n30412, n30413,
    n30414, n30415, n30416, n30417, n30418, n30419,
    n30420, n30421, n30422, n30423, n30424, n30425,
    n30426, n30427, n30428, n30429, n30430, n30431,
    n30432, n30433, n30434, n30435, n30436, n30437,
    n30438, n30439, n30440, n30441, n30442, n30443,
    n30444, n30445, n30446, n30447, n30448, n30449,
    n30450, n30451, n30452, n30453, n30454, n30455,
    n30456, n30457, n30458, n30459, n30460, n30461,
    n30462, n30463, n30464, n30465, n30466, n30467,
    n30468, n30469, n30470, n30471, n30472, n30473,
    n30474, n30475, n30476, n30477, n30478, n30479,
    n30480, n30481, n30482, n30483, n30484, n30485,
    n30486, n30487, n30488, n30489, n30490, n30491,
    n30492, n30493, n30494, n30495, n30496, n30497,
    n30498, n30499, n30500, n30501, n30502, n30503,
    n30504, n30505, n30506, n30507, n30508, n30509,
    n30510, n30511, n30512, n30513, n30514, n30515,
    n30516, n30517, n30518, n30519, n30520, n30521,
    n30522, n30523, n30524, n30525, n30526, n30527,
    n30528, n30529, n30530, n30531, n30532, n30533,
    n30534, n30535, n30536, n30537, n30538, n30539,
    n30540, n30541, n30542, n30543, n30544, n30545,
    n30546, n30547, n30548, n30549, n30550, n30551,
    n30552, n30553, n30554, n30555, n30556, n30557,
    n30558, n30559, n30560, n30561, n30562, n30563,
    n30564, n30565, n30566, n30567, n30568, n30569,
    n30570, n30571, n30572, n30573, n30574, n30575,
    n30576, n30577, n30578, n30579, n30580, n30581,
    n30582, n30583, n30584, n30585, n30586, n30587,
    n30589, n30590, n30591, n30592, n30593, n30594,
    n30595, n30596, n30597, n30598, n30599, n30600,
    n30601, n30602, n30603, n30604, n30605, n30606,
    n30607, n30608, n30609, n30610, n30611, n30612,
    n30613, n30614, n30615, n30616, n30617, n30618,
    n30619, n30620, n30621, n30622, n30623, n30624,
    n30625, n30626, n30627, n30628, n30629, n30630,
    n30631, n30632, n30633, n30634, n30635, n30636,
    n30637, n30638, n30639, n30640, n30641, n30642,
    n30643, n30644, n30645, n30646, n30647, n30648,
    n30649, n30650, n30651, n30652, n30653, n30654,
    n30655, n30656, n30657, n30658, n30659, n30660,
    n30661, n30662, n30663, n30664, n30665, n30666,
    n30667, n30668, n30669, n30670, n30671, n30672,
    n30673, n30674, n30675, n30676, n30677, n30678,
    n30679, n30680, n30681, n30682, n30683, n30684,
    n30685, n30686, n30687, n30688, n30689, n30690,
    n30691, n30692, n30693, n30694, n30695, n30696,
    n30697, n30698, n30699, n30700, n30701, n30702,
    n30703, n30704, n30705, n30706, n30707, n30708,
    n30709, n30710, n30711, n30712, n30713, n30714,
    n30715, n30716, n30717, n30718, n30719, n30720,
    n30721, n30722, n30723, n30724, n30725, n30726,
    n30727, n30728, n30729, n30730, n30731, n30732,
    n30733, n30734, n30735, n30736, n30737, n30738,
    n30739, n30740, n30741, n30742, n30743, n30744,
    n30745, n30746, n30747, n30748, n30749, n30750,
    n30751, n30752, n30753, n30754, n30755, n30756,
    n30757, n30758, n30759, n30760, n30761, n30762,
    n30763, n30764, n30765, n30766, n30767, n30768,
    n30769, n30770, n30771, n30772, n30773, n30774,
    n30775, n30776, n30777, n30778, n30779, n30780,
    n30781, n30782, n30783, n30784, n30785, n30786,
    n30787, n30788, n30789, n30790, n30791, n30792,
    n30793, n30794, n30795, n30796, n30797, n30798,
    n30799, n30800, n30801, n30802, n30803, n30804,
    n30805, n30806, n30807, n30808, n30809, n30810,
    n30811, n30812, n30813, n30814, n30815, n30816,
    n30817, n30818, n30819, n30820, n30821, n30822,
    n30823, n30824, n30825, n30826, n30827, n30828,
    n30829, n30830, n30831, n30832, n30833, n30834,
    n30835, n30836, n30837, n30838, n30839, n30840,
    n30841, n30842, n30843, n30844, n30845, n30846,
    n30847, n30848, n30849, n30850, n30851, n30852,
    n30853, n30854, n30855, n30856, n30857, n30858,
    n30859, n30860, n30861, n30862, n30863, n30864,
    n30865, n30866, n30867, n30868, n30869, n30870,
    n30871, n30872, n30873, n30874, n30875, n30876,
    n30877, n30878, n30879, n30880, n30881, n30882,
    n30883, n30884, n30885, n30886, n30887, n30888,
    n30889, n30890, n30891, n30892, n30893, n30894,
    n30895, n30896, n30897, n30898, n30899, n30900,
    n30901, n30902, n30903, n30904, n30905, n30906,
    n30907, n30908, n30909, n30910, n30911, n30912,
    n30913, n30914, n30915, n30916, n30917, n30918,
    n30919, n30920, n30921, n30922, n30923, n30924,
    n30925, n30926, n30927, n30928, n30929, n30930,
    n30931, n30932, n30933, n30934, n30935, n30936,
    n30937, n30938, n30939, n30940, n30941, n30942,
    n30943, n30944, n30945, n30946, n30947, n30948,
    n30949, n30950, n30951, n30952, n30953, n30954,
    n30955, n30956, n30957, n30958, n30959, n30960,
    n30961, n30962, n30963, n30964, n30965, n30966,
    n30967, n30968, n30969, n30970, n30971, n30972,
    n30973, n30974, n30975, n30976, n30977, n30978,
    n30979, n30980, n30981, n30982, n30983, n30984,
    n30985, n30986, n30987, n30988, n30989, n30990,
    n30991, n30992, n30993, n30994, n30995, n30996,
    n30997, n30998, n30999, n31000, n31001, n31002,
    n31003, n31004, n31005, n31006, n31007, n31008,
    n31009, n31010, n31011, n31012, n31013, n31014,
    n31015, n31016, n31017, n31018, n31019, n31020,
    n31021, n31022, n31023, n31024, n31025, n31026,
    n31027, n31028, n31029, n31030, n31031, n31032,
    n31033, n31034, n31035, n31036, n31037, n31038,
    n31039, n31040, n31041, n31042, n31043, n31044,
    n31045, n31046, n31047, n31048, n31049, n31050,
    n31051, n31052, n31053, n31054, n31055, n31056,
    n31058, n31059, n31060, n31061, n31062, n31063,
    n31064, n31065, n31066, n31067, n31068, n31069,
    n31070, n31071, n31072, n31073, n31074, n31075,
    n31076, n31077, n31078, n31079, n31080, n31081,
    n31082, n31083, n31084, n31085, n31086, n31087,
    n31088, n31089, n31090, n31091, n31092, n31093,
    n31094, n31095, n31096, n31097, n31098, n31099,
    n31100, n31101, n31102, n31103, n31104, n31105,
    n31106, n31107, n31108, n31109, n31110, n31111,
    n31112, n31113, n31114, n31115, n31116, n31117,
    n31118, n31119, n31120, n31121, n31122, n31123,
    n31124, n31125, n31126, n31127, n31128, n31129,
    n31130, n31131, n31132, n31133, n31134, n31135,
    n31136, n31137, n31138, n31139, n31140, n31141,
    n31142, n31143, n31144, n31145, n31146, n31147,
    n31148, n31149, n31150, n31151, n31152, n31153,
    n31154, n31155, n31156, n31157, n31158, n31159,
    n31160, n31161, n31162, n31163, n31164, n31165,
    n31166, n31167, n31168, n31169, n31170, n31171,
    n31172, n31173, n31174, n31175, n31176, n31177,
    n31178, n31179, n31180, n31181, n31182, n31183,
    n31184, n31185, n31186, n31187, n31188, n31189,
    n31190, n31191, n31192, n31193, n31194, n31195,
    n31196, n31197, n31198, n31199, n31200, n31201,
    n31202, n31203, n31204, n31205, n31206, n31207,
    n31208, n31209, n31210, n31211, n31212, n31213,
    n31214, n31215, n31216, n31217, n31218, n31219,
    n31220, n31221, n31222, n31223, n31224, n31225,
    n31226, n31227, n31228, n31229, n31230, n31231,
    n31232, n31233, n31234, n31235, n31236, n31237,
    n31238, n31239, n31240, n31241, n31242, n31243,
    n31244, n31245, n31246, n31247, n31248, n31249,
    n31250, n31251, n31252, n31253, n31254, n31255,
    n31256, n31257, n31258, n31259, n31260, n31261,
    n31262, n31263, n31264, n31265, n31266, n31267,
    n31268, n31269, n31270, n31271, n31272, n31273,
    n31274, n31275, n31276, n31277, n31278, n31279,
    n31280, n31281, n31282, n31283, n31284, n31285,
    n31286, n31287, n31288, n31289, n31290, n31291,
    n31292, n31293, n31294, n31295, n31296, n31297,
    n31298, n31299, n31300, n31301, n31302, n31303,
    n31304, n31305, n31306, n31307, n31308, n31309,
    n31310, n31311, n31312, n31313, n31314, n31315,
    n31316, n31317, n31318, n31319, n31320, n31321,
    n31322, n31323, n31324, n31325, n31326, n31327,
    n31328, n31329, n31330, n31331, n31332, n31333,
    n31334, n31335, n31336, n31337, n31338, n31339,
    n31340, n31341, n31342, n31343, n31344, n31345,
    n31346, n31347, n31348, n31349, n31350, n31351,
    n31352, n31353, n31354, n31355, n31356, n31357,
    n31358, n31359, n31360, n31361, n31362, n31363,
    n31364, n31365, n31366, n31367, n31368, n31369,
    n31370, n31371, n31372, n31373, n31374, n31375,
    n31376, n31377, n31378, n31379, n31380, n31381,
    n31382, n31383, n31384, n31385, n31386, n31387,
    n31388, n31389, n31390, n31391, n31392, n31393,
    n31394, n31395, n31396, n31397, n31398, n31399,
    n31400, n31401, n31402, n31403, n31404, n31405,
    n31406, n31407, n31408, n31409, n31410, n31411,
    n31412, n31413, n31414, n31415, n31416, n31417,
    n31418, n31419, n31420, n31421, n31422, n31423,
    n31424, n31425, n31426, n31427, n31428, n31429,
    n31430, n31431, n31432, n31433, n31434, n31435,
    n31436, n31437, n31438, n31439, n31440, n31441,
    n31442, n31443, n31444, n31445, n31446, n31447,
    n31448, n31449, n31450, n31451, n31452, n31453,
    n31454, n31455, n31456, n31457, n31458, n31459,
    n31460, n31461, n31462, n31463, n31464, n31465,
    n31466, n31467, n31468, n31469, n31470, n31471,
    n31472, n31473, n31474, n31475, n31476, n31477,
    n31478, n31479, n31480, n31481, n31482, n31483,
    n31484, n31485, n31486, n31487, n31488, n31489,
    n31490, n31491, n31492, n31493, n31494, n31495,
    n31496, n31497, n31498, n31499, n31500, n31501,
    n31502, n31503, n31504, n31505, n31506, n31507,
    n31508, n31509, n31510, n31511, n31512, n31513,
    n31514, n31515, n31516, n31517, n31518, n31519,
    n31520, n31521, n31522, n31523, n31524, n31525,
    n31527, n31528, n31529, n31530, n31531, n31532,
    n31533, n31534, n31535, n31536, n31537, n31538,
    n31539, n31540, n31541, n31542, n31543, n31544,
    n31545, n31546, n31547, n31548, n31549, n31550,
    n31551, n31552, n31553, n31554, n31555, n31556,
    n31557, n31558, n31559, n31560, n31561, n31562,
    n31563, n31564, n31565, n31566, n31567, n31568,
    n31569, n31570, n31571, n31572, n31573, n31574,
    n31575, n31576, n31577, n31578, n31579, n31580,
    n31581, n31582, n31583, n31584, n31585, n31586,
    n31587, n31588, n31589, n31590, n31591, n31592,
    n31593, n31594, n31595, n31596, n31597, n31598,
    n31599, n31600, n31601, n31602, n31603, n31604,
    n31605, n31606, n31607, n31608, n31609, n31610,
    n31611, n31612, n31613, n31614, n31615, n31616,
    n31617, n31618, n31619, n31620, n31621, n31622,
    n31623, n31624, n31625, n31626, n31627, n31628,
    n31629, n31630, n31631, n31632, n31633, n31634,
    n31635, n31636, n31637, n31638, n31639, n31640,
    n31641, n31642, n31643, n31644, n31645, n31646,
    n31647, n31648, n31649, n31650, n31651, n31652,
    n31653, n31654, n31655, n31656, n31657, n31658,
    n31659, n31660, n31661, n31662, n31663, n31664,
    n31665, n31666, n31667, n31668, n31669, n31670,
    n31671, n31672, n31673, n31674, n31675, n31676,
    n31677, n31678, n31679, n31680, n31681, n31682,
    n31683, n31684, n31685, n31686, n31687, n31688,
    n31689, n31690, n31691, n31692, n31693, n31694,
    n31695, n31696, n31697, n31698, n31699, n31700,
    n31701, n31702, n31703, n31704, n31705, n31706,
    n31707, n31708, n31709, n31710, n31711, n31712,
    n31713, n31714, n31715, n31716, n31717, n31718,
    n31719, n31720, n31721, n31722, n31723, n31724,
    n31725, n31726, n31727, n31728, n31729, n31730,
    n31731, n31732, n31733, n31734, n31735, n31736,
    n31737, n31738, n31739, n31740, n31741, n31742,
    n31743, n31744, n31745, n31746, n31747, n31748,
    n31749, n31750, n31751, n31752, n31753, n31754,
    n31755, n31756, n31757, n31758, n31759, n31760,
    n31761, n31762, n31763, n31764, n31765, n31766,
    n31767, n31768, n31769, n31770, n31771, n31772,
    n31773, n31774, n31775, n31776, n31777, n31778,
    n31779, n31780, n31781, n31782, n31783, n31784,
    n31785, n31786, n31787, n31788, n31789, n31790,
    n31791, n31792, n31793, n31794, n31795, n31796,
    n31797, n31798, n31799, n31800, n31801, n31802,
    n31803, n31804, n31805, n31806, n31807, n31808,
    n31809, n31810, n31811, n31812, n31813, n31814,
    n31815, n31816, n31817, n31818, n31819, n31820,
    n31821, n31822, n31823, n31824, n31825, n31826,
    n31827, n31828, n31829, n31830, n31831, n31832,
    n31833, n31834, n31835, n31836, n31837, n31838,
    n31839, n31840, n31841, n31842, n31843, n31844,
    n31845, n31846, n31847, n31848, n31849, n31850,
    n31851, n31852, n31853, n31854, n31855, n31856,
    n31857, n31858, n31859, n31860, n31861, n31862,
    n31863, n31864, n31865, n31866, n31867, n31868,
    n31869, n31870, n31871, n31872, n31873, n31874,
    n31875, n31876, n31877, n31878, n31879, n31880,
    n31881, n31882, n31883, n31884, n31885, n31886,
    n31887, n31888, n31889, n31890, n31891, n31892,
    n31893, n31894, n31895, n31896, n31897, n31898,
    n31899, n31900, n31901, n31902, n31903, n31904,
    n31905, n31906, n31907, n31908, n31909, n31910,
    n31911, n31912, n31913, n31914, n31915, n31916,
    n31917, n31918, n31919, n31920, n31921, n31922,
    n31923, n31924, n31925, n31926, n31927, n31928,
    n31929, n31930, n31931, n31932, n31933, n31934,
    n31935, n31936, n31937, n31938, n31939, n31940,
    n31941, n31942, n31943, n31944, n31945, n31946,
    n31947, n31948, n31949, n31950, n31951, n31952,
    n31953, n31954, n31955, n31956, n31957, n31958,
    n31959, n31960, n31961, n31962, n31963, n31964,
    n31965, n31966, n31967, n31968, n31969, n31970,
    n31971, n31972, n31973, n31974, n31975, n31976,
    n31977, n31978, n31979, n31980, n31981, n31982,
    n31983, n31984, n31985, n31986, n31987, n31988,
    n31989, n31990, n31991, n31992, n31993, n31994,
    n31996, n31997, n31998, n31999, n32000, n32001,
    n32002, n32003, n32004, n32005, n32006, n32007,
    n32008, n32009, n32010, n32011, n32012, n32013,
    n32014, n32015, n32016, n32017, n32018, n32019,
    n32020, n32021, n32022, n32023, n32024, n32025,
    n32026, n32027, n32028, n32029, n32030, n32031,
    n32032, n32033, n32034, n32035, n32036, n32037,
    n32038, n32039, n32040, n32041, n32042, n32043,
    n32044, n32045, n32046, n32047, n32048, n32049,
    n32050, n32051, n32052, n32053, n32054, n32055,
    n32056, n32057, n32058, n32059, n32060, n32061,
    n32062, n32063, n32064, n32065, n32066, n32067,
    n32068, n32069, n32070, n32071, n32072, n32073,
    n32074, n32075, n32076, n32077, n32078, n32079,
    n32080, n32081, n32082, n32083, n32084, n32085,
    n32086, n32087, n32088, n32089, n32090, n32091,
    n32092, n32093, n32094, n32095, n32096, n32097,
    n32098, n32099, n32100, n32101, n32102, n32103,
    n32104, n32105, n32106, n32107, n32108, n32109,
    n32110, n32111, n32112, n32113, n32114, n32115,
    n32116, n32117, n32118, n32119, n32120, n32121,
    n32122, n32123, n32124, n32125, n32126, n32127,
    n32128, n32129, n32130, n32131, n32132, n32133,
    n32134, n32135, n32136, n32137, n32138, n32139,
    n32140, n32141, n32142, n32143, n32144, n32145,
    n32146, n32147, n32148, n32149, n32150, n32151,
    n32152, n32153, n32154, n32155, n32156, n32157,
    n32158, n32159, n32160, n32161, n32162, n32163,
    n32164, n32165, n32166, n32167, n32168, n32169,
    n32170, n32171, n32172, n32173, n32174, n32175,
    n32176, n32177, n32178, n32179, n32180, n32181,
    n32182, n32183, n32184, n32185, n32186, n32187,
    n32188, n32189, n32190, n32191, n32192, n32193,
    n32194, n32195, n32196, n32197, n32198, n32199,
    n32200, n32201, n32202, n32203, n32204, n32205,
    n32206, n32207, n32208, n32209, n32210, n32211,
    n32212, n32213, n32214, n32215, n32216, n32217,
    n32218, n32219, n32220, n32221, n32222, n32223,
    n32224, n32225, n32226, n32227, n32228, n32229,
    n32230, n32231, n32232, n32233, n32234, n32235,
    n32236, n32237, n32238, n32239, n32240, n32241,
    n32242, n32243, n32244, n32245, n32246, n32247,
    n32248, n32249, n32250, n32251, n32252, n32253,
    n32254, n32255, n32256, n32257, n32258, n32259,
    n32260, n32261, n32262, n32263, n32264, n32265,
    n32266, n32267, n32268, n32269, n32270, n32271,
    n32272, n32273, n32274, n32275, n32276, n32277,
    n32278, n32279, n32280, n32281, n32282, n32283,
    n32284, n32285, n32286, n32287, n32288, n32289,
    n32290, n32291, n32292, n32293, n32294, n32295,
    n32296, n32297, n32298, n32299, n32300, n32301,
    n32302, n32303, n32304, n32305, n32306, n32307,
    n32308, n32309, n32310, n32311, n32312, n32313,
    n32314, n32315, n32316, n32317, n32318, n32319,
    n32320, n32321, n32322, n32323, n32324, n32325,
    n32326, n32327, n32328, n32329, n32330, n32331,
    n32332, n32333, n32334, n32335, n32336, n32337,
    n32338, n32339, n32340, n32341, n32342, n32343,
    n32344, n32345, n32346, n32347, n32348, n32349,
    n32350, n32351, n32352, n32353, n32354, n32355,
    n32356, n32357, n32358, n32359, n32360, n32361,
    n32362, n32363, n32364, n32365, n32366, n32367,
    n32368, n32369, n32370, n32371, n32372, n32373,
    n32374, n32375, n32376, n32377, n32378, n32379,
    n32380, n32381, n32382, n32383, n32384, n32385,
    n32386, n32387, n32388, n32389, n32390, n32391,
    n32392, n32393, n32394, n32395, n32396, n32397,
    n32398, n32399, n32400, n32401, n32402, n32403,
    n32404, n32405, n32406, n32407, n32408, n32409,
    n32410, n32411, n32412, n32413, n32414, n32415,
    n32416, n32417, n32418, n32419, n32420, n32421,
    n32422, n32423, n32424, n32425, n32426, n32427,
    n32428, n32429, n32430, n32431, n32432, n32433,
    n32434, n32435, n32436, n32437, n32438, n32439,
    n32440, n32441, n32442, n32443, n32444, n32445,
    n32446, n32447, n32448, n32449, n32450, n32451,
    n32452, n32453, n32454, n32455, n32456, n32457,
    n32458, n32459, n32460, n32462, n32463, n32464,
    n32465, n32466, n32467, n32468, n32469, n32470,
    n32471, n32472, n32473, n32474, n32475, n32476,
    n32477, n32478, n32479, n32480, n32481, n32482,
    n32483, n32484, n32485, n32486, n32487, n32488,
    n32489, n32490, n32491, n32492, n32493, n32494,
    n32495, n32496, n32497, n32498, n32499, n32500,
    n32501, n32502, n32503, n32504, n32505, n32506,
    n32507, n32508, n32509, n32510, n32512, n32513,
    n32514, n32515, n32516, n32517, n32518, n32519,
    n32520, n32521, n32522, n32523, n32524, n32525,
    n32526, n32527, n32528, n32529, n32530, n32531,
    n32532, n32533, n32534, n32535, n32536, n32537,
    n32538, n32539, n32540, n32541, n32542, n32543,
    n32544, n32545, n32546, n32547, n32548, n32549,
    n32550, n32551, n32552, n32553, n32554, n32555,
    n32556, n32557, n32558, n32559, n32560, n32561,
    n32562, n32563, n32564, n32565, n32566, n32567,
    n32568, n32569, n32570, n32571, n32572, n32573,
    n32574, n32575, n32576, n32577, n32578, n32579,
    n32580, n32582, n32583, n32584, n32585, n32586,
    n32587, n32588, n32589, n32590, n32591, n32592,
    n32593, n32594, n32595, n32596, n32597, n32598,
    n32599, n32600, n32601, n32602, n32603, n32604,
    n32605, n32606, n32607, n32608, n32609, n32610,
    n32611, n32612, n32613, n32614, n32615, n32616,
    n32617, n32618, n32619, n32620, n32621, n32622,
    n32623, n32624, n32625, n32626, n32627, n32628,
    n32629, n32630, n32631, n32632, n32633, n32634,
    n32635, n32636, n32637, n32638, n32640, n32641,
    n32642, n32643, n32644, n32645, n32646, n32647,
    n32648, n32649, n32650, n32651, n32652, n32653,
    n32654, n32655, n32656, n32657, n32658, n32659,
    n32660, n32661, n32662, n32663, n32664, n32665,
    n32666, n32667, n32668, n32669, n32670, n32671,
    n32672, n32673, n32674, n32675, n32676, n32677,
    n32678, n32679, n32680, n32681, n32682, n32683,
    n32684, n32685, n32686, n32687, n32688, n32689,
    n32690, n32691, n32692, n32693, n32694, n32695,
    n32696, n32697, n32698, n32699, n32700, n32701,
    n32702, n32703, n32704, n32705, n32706, n32707,
    n32708, n32709, n32710, n32711, n32712, n32713,
    n32714, n32715, n32716, n32717, n32718, n32719,
    n32720, n32721, n32722, n32723, n32724, n32725,
    n32726, n32727, n32728, n32729, n32730, n32731,
    n32732, n32733, n32734, n32735, n32736, n32737,
    n32738, n32739, n32740, n32741, n32742, n32743,
    n32744, n32745, n32746, n32747, n32748, n32749,
    n32750, n32751, n32752, n32753, n32754, n32755,
    n32756, n32757, n32758, n32759, n32760, n32761,
    n32762, n32763, n32764, n32765, n32766, n32767,
    n32768, n32769, n32770, n32771, n32772, n32773,
    n32774, n32775, n32776, n32777, n32778, n32779,
    n32780, n32781, n32782, n32783, n32784, n32785,
    n32786, n32787, n32788, n32789, n32790, n32791,
    n32792, n32793, n32794, n32795, n32796, n32797,
    n32798, n32799, n32800, n32801, n32802, n32803,
    n32804, n32805, n32806, n32807, n32808, n32809,
    n32810, n32811, n32812, n32813, n32814, n32815,
    n32816, n32817, n32818, n32819, n32820, n32821,
    n32822, n32823, n32824, n32825, n32826, n32827,
    n32828, n32829, n32830, n32831, n32832, n32833,
    n32834, n32835, n32836, n32837, n32838, n32839,
    n32840, n32841, n32842, n32843, n32844, n32845,
    n32846, n32847, n32848, n32849, n32850, n32851,
    n32852, n32853, n32854, n32855, n32856, n32857,
    n32858, n32859, n32860, n32861, n32862, n32863,
    n32864, n32865, n32866, n32867, n32868, n32869,
    n32870, n32871, n32872, n32873, n32874, n32875,
    n32876, n32877, n32878, n32879, n32880, n32881,
    n32882, n32883, n32884, n32885, n32886, n32887,
    n32888, n32889, n32890, n32891, n32892, n32893,
    n32894, n32895, n32896, n32897, n32898, n32899,
    n32900, n32901, n32902, n32903, n32904, n32905,
    n32906, n32907, n32908, n32909, n32910, n32911,
    n32912, n32913, n32914, n32915, n32916, n32917,
    n32918, n32919, n32920, n32921, n32922, n32923,
    n32924, n32925, n32926, n32927, n32928, n32929,
    n32930, n32931, n32932, n32933, n32934, n32935,
    n32936, n32937, n32938, n32939, n32940, n32941,
    n32942, n32943, n32944, n32945, n32946, n32947,
    n32948, n32949, n32950, n32951, n32952, n32953,
    n32954, n32955, n32956, n32957, n32958, n32959,
    n32960, n32961, n32962, n32963, n32964, n32965,
    n32966, n32967, n32968, n32969, n32970, n32971,
    n32972, n32973, n32974, n32975, n32976, n32977,
    n32978, n32979, n32980, n32981, n32982, n32983,
    n32984, n32985, n32986, n32987, n32988, n32989,
    n32990, n32991, n32992, n32993, n32994, n32995,
    n32996, n32997, n32998, n32999, n33000, n33001,
    n33002, n33003, n33004, n33005, n33006, n33007,
    n33008, n33009, n33010, n33011, n33012, n33013,
    n33014, n33015, n33016, n33017, n33018, n33019,
    n33020, n33021, n33022, n33023, n33024, n33025,
    n33026, n33027, n33028, n33029, n33030, n33031,
    n33032, n33033, n33034, n33035, n33036, n33037,
    n33038, n33039, n33040, n33041, n33042, n33043,
    n33044, n33045, n33046, n33047, n33048, n33049,
    n33050, n33051, n33052, n33053, n33054, n33055,
    n33056, n33057, n33058, n33059, n33060, n33061,
    n33062, n33063, n33064, n33065, n33066, n33067,
    n33068, n33069, n33070, n33071, n33072, n33073,
    n33074, n33075, n33076, n33077, n33078, n33079,
    n33080, n33081, n33082, n33083, n33084, n33085,
    n33086, n33087, n33088, n33089, n33090, n33091,
    n33092, n33093, n33094, n33095, n33096, n33097,
    n33098, n33099, n33100, n33101, n33102, n33103,
    n33104, n33105, n33106, n33107, n33108, n33109,
    n33110, n33111, n33112, n33113, n33114, n33115,
    n33116, n33117, n33118, n33119, n33120, n33121,
    n33122, n33123, n33124, n33125, n33126, n33127,
    n33128, n33129, n33130, n33131, n33132, n33133,
    n33134, n33135, n33136, n33137, n33138, n33139,
    n33140, n33141, n33142, n33143, n33144, n33145,
    n33146, n33147, n33148, n33149, n33150, n33151,
    n33152, n33153, n33154, n33155, n33156, n33157,
    n33158, n33159, n33160, n33161, n33162, n33163,
    n33164, n33165, n33166, n33167, n33168, n33169,
    n33170, n33171, n33172, n33173, n33174, n33175,
    n33176, n33177, n33178, n33179, n33180, n33181,
    n33182, n33183, n33184, n33185, n33186, n33187,
    n33188, n33189, n33190, n33191, n33192, n33193,
    n33194, n33195, n33196, n33197, n33198, n33199,
    n33200, n33201, n33202, n33203, n33204, n33205,
    n33206, n33207, n33208, n33209, n33210, n33211,
    n33212, n33213, n33214, n33215, n33216, n33217,
    n33218, n33219, n33220, n33221, n33222, n33223,
    n33224, n33225, n33226, n33227, n33228, n33229,
    n33230, n33231, n33232, n33233, n33234, n33235,
    n33236, n33237, n33238, n33239, n33240, n33241,
    n33242, n33243, n33244, n33245, n33246, n33247,
    n33248, n33249, n33250, n33251, n33252, n33253,
    n33254, n33255, n33256, n33258, n33259, n33260,
    n33261, n33262, n33263, n33264, n33265, n33266,
    n33267, n33268, n33269, n33270, n33271, n33272,
    n33273, n33274, n33275, n33276, n33277, n33278,
    n33279, n33280, n33281, n33282, n33283, n33284,
    n33285, n33286, n33287, n33288, n33289, n33290,
    n33291, n33292, n33293, n33294, n33295, n33296,
    n33297, n33298, n33299, n33300, n33301, n33302,
    n33303, n33304, n33305, n33306, n33307, n33308,
    n33309, n33310, n33311, n33312, n33313, n33314,
    n33315, n33316, n33317, n33318, n33319, n33320,
    n33321, n33322, n33323, n33324, n33325, n33326,
    n33327, n33328, n33329, n33330, n33331, n33332,
    n33333, n33334, n33335, n33336, n33337, n33338,
    n33339, n33340, n33341, n33342, n33343, n33344,
    n33345, n33346, n33347, n33348, n33349, n33350,
    n33351, n33352, n33353, n33354, n33355, n33356,
    n33357, n33358, n33359, n33360, n33361, n33362,
    n33363, n33364, n33365, n33366, n33367, n33368,
    n33369, n33370, n33371, n33372, n33373, n33374,
    n33375, n33376, n33377, n33378, n33379, n33380,
    n33381, n33382, n33383, n33384, n33385, n33386,
    n33387, n33388, n33389, n33390, n33391, n33392,
    n33393, n33394, n33395, n33396, n33397, n33398,
    n33399, n33400, n33401, n33402, n33403, n33404,
    n33405, n33406, n33407, n33408, n33409, n33410,
    n33411, n33412, n33413, n33414, n33415, n33416,
    n33417, n33418, n33419, n33420, n33421, n33422,
    n33423, n33424, n33425, n33426, n33427, n33428,
    n33429, n33430, n33431, n33432, n33433, n33434,
    n33435, n33436, n33437, n33438, n33439, n33440,
    n33441, n33442, n33443, n33444, n33445, n33446,
    n33447, n33448, n33449, n33450, n33451, n33452,
    n33453, n33454, n33455, n33456, n33457, n33458,
    n33459, n33460, n33461, n33462, n33463, n33464,
    n33465, n33466, n33467, n33468, n33469, n33470,
    n33471, n33472, n33473, n33474, n33475, n33476,
    n33477, n33478, n33479, n33480, n33481, n33482,
    n33483, n33484, n33485, n33486, n33487, n33488,
    n33489, n33490, n33491, n33492, n33493, n33494,
    n33495, n33496, n33497, n33498, n33499, n33500,
    n33501, n33502, n33503, n33504, n33505, n33506,
    n33507, n33508, n33509, n33510, n33511, n33512,
    n33513, n33514, n33515, n33516, n33517, n33518,
    n33519, n33520, n33521, n33522, n33523, n33524,
    n33525, n33526, n33527, n33528, n33529, n33530,
    n33531, n33532, n33533, n33534, n33535, n33536,
    n33537, n33538, n33539, n33540, n33541, n33542,
    n33543, n33544, n33545, n33546, n33547, n33548,
    n33550, n33551, n33552, n33553, n33554, n33555,
    n33556, n33557, n33558, n33559, n33560, n33561,
    n33562, n33563, n33564, n33565, n33566, n33567,
    n33568, n33569, n33570, n33571, n33572, n33573,
    n33574, n33575, n33576, n33577, n33578, n33579,
    n33580, n33581, n33582, n33583, n33584, n33585,
    n33586, n33587, n33588, n33589, n33590, n33591,
    n33592, n33593, n33594, n33595, n33596, n33597,
    n33598, n33599, n33600, n33601, n33602, n33603,
    n33604, n33605, n33606, n33607, n33608, n33609,
    n33610, n33611, n33612, n33613, n33614, n33615,
    n33616, n33617, n33618, n33619, n33620, n33621,
    n33622, n33623, n33624, n33625, n33626, n33627,
    n33628, n33629, n33630, n33631, n33632, n33633,
    n33634, n33635, n33636, n33637, n33638, n33639,
    n33640, n33641, n33642, n33643, n33644, n33645,
    n33646, n33647, n33648, n33649, n33650, n33651,
    n33652, n33653, n33654, n33655, n33656, n33657,
    n33658, n33659, n33660, n33661, n33662, n33663,
    n33664, n33665, n33666, n33667, n33668, n33669,
    n33670, n33671, n33672, n33673, n33674, n33675,
    n33676, n33677, n33678, n33679, n33680, n33681,
    n33682, n33683, n33684, n33685, n33686, n33687,
    n33688, n33689, n33690, n33691, n33692, n33693,
    n33694, n33695, n33696, n33697, n33698, n33699,
    n33700, n33701, n33702, n33703, n33704, n33705,
    n33706, n33707, n33708, n33709, n33710, n33711,
    n33712, n33713, n33714, n33715, n33716, n33717,
    n33718, n33719, n33720, n33721, n33722, n33723,
    n33724, n33725, n33726, n33727, n33728, n33729,
    n33730, n33731, n33732, n33733, n33734, n33735,
    n33736, n33737, n33738, n33739, n33740, n33741,
    n33742, n33743, n33744, n33745, n33746, n33747,
    n33748, n33749, n33750, n33751, n33752, n33753,
    n33754, n33755, n33756, n33757, n33758, n33759,
    n33760, n33761, n33762, n33763, n33764, n33765,
    n33766, n33767, n33768, n33769, n33770, n33771,
    n33772, n33773, n33774, n33775, n33776, n33777,
    n33778, n33779, n33780, n33781, n33782, n33783,
    n33784, n33785, n33786, n33787, n33788, n33789,
    n33790, n33791, n33792, n33793, n33794, n33795,
    n33796, n33797, n33798, n33799, n33800, n33801,
    n33802, n33803, n33804, n33805, n33806, n33807,
    n33808, n33809, n33810, n33811, n33812, n33813,
    n33814, n33815, n33816, n33817, n33818, n33819,
    n33820, n33821, n33822, n33823, n33824, n33825,
    n33826, n33827, n33828, n33830, n33831, n33832,
    n33833, n33834, n33835, n33836, n33837, n33838,
    n33839, n33840, n33841, n33842, n33843, n33844,
    n33845, n33846, n33847, n33848, n33849, n33850,
    n33851, n33852, n33853, n33854, n33855, n33856,
    n33857, n33858, n33859, n33860, n33861, n33862,
    n33863, n33864, n33865, n33866, n33867, n33868,
    n33869, n33870, n33871, n33872, n33873, n33874,
    n33875, n33876, n33877, n33878, n33879, n33880,
    n33881, n33882, n33883, n33884, n33885, n33886,
    n33887, n33888, n33889, n33890, n33891, n33892,
    n33893, n33894, n33895, n33896, n33897, n33898,
    n33899, n33900, n33901, n33902, n33903, n33904,
    n33905, n33906, n33907, n33908, n33909, n33910,
    n33911, n33912, n33913, n33914, n33915, n33916,
    n33917, n33918, n33919, n33920, n33921, n33922,
    n33923, n33924, n33925, n33926, n33927, n33928,
    n33929, n33930, n33931, n33932, n33933, n33934,
    n33935, n33936, n33937, n33938, n33939, n33940,
    n33941, n33942, n33943, n33944, n33945, n33946,
    n33947, n33948, n33949, n33950, n33951, n33952,
    n33953, n33954, n33955, n33956, n33957, n33958,
    n33959, n33960, n33961, n33962, n33963, n33964,
    n33965, n33966, n33967, n33968, n33969, n33970,
    n33971, n33972, n33973, n33974, n33975, n33976,
    n33977, n33978, n33979, n33980, n33981, n33982,
    n33983, n33984, n33985, n33986, n33987, n33988,
    n33989, n33990, n33991, n33992, n33993, n33994,
    n33995, n33996, n33997, n33998, n33999, n34000,
    n34001, n34002, n34003, n34004, n34005, n34006,
    n34007, n34008, n34009, n34010, n34011, n34012,
    n34013, n34014, n34015, n34016, n34017, n34018,
    n34019, n34020, n34021, n34022, n34023, n34025,
    n34026, n34027, n34028, n34029, n34030, n34031,
    n34033, n34034, n34035, n34036, n34037, n34038,
    n34039, n34041, n34042, n34043, n34044, n34045,
    n34046, n34047, n34048, n34049, n34050, n34051,
    n34052, n34053, n34054, n34055, n34056, n34057,
    n34058, n34059, n34060, n34061, n34062, n34063,
    n34064, n34065, n34066, n34067, n34068, n34069,
    n34070, n34071, n34072, n34073, n34074, n34075,
    n34076, n34077, n34078, n34079, n34080, n34081,
    n34082, n34083, n34084, n34085, n34086, n34087,
    n34088, n34089, n34090, n34091, n34092, n34093,
    n34094, n34095, n34096, n34097, n34098, n34099,
    n34100, n34101, n34102, n34103, n34104, n34105,
    n34106, n34107, n34108, n34109, n34110, n34111,
    n34112, n34113, n34114, n34115, n34116, n34117,
    n34118, n34119, n34120, n34121, n34122, n34123,
    n34124, n34125, n34126, n34127, n34128, n34129,
    n34130, n34131, n34132, n34133, n34134, n34135,
    n34136, n34137, n34138, n34139, n34140, n34141,
    n34142, n34143, n34144, n34145, n34146, n34147,
    n34149, n34150, n34151, n34152, n34153, n34154,
    n34156, n34157, n34158, n34159, n34160, n34161,
    n34162, n34164, n34165, n34166, n34167, n34168,
    n34169, n34170, n34171, n34172, n34173, n34174,
    n34175, n34176, n34177, n34178, n34179, n34180,
    n34181, n34182, n34183, n34184, n34185, n34186,
    n34187, n34188, n34189, n34190, n34191, n34192,
    n34193, n34194, n34195, n34196, n34197, n34198,
    n34199, n34200, n34201, n34202, n34203, n34204,
    n34205, n34206, n34207, n34208, n34209, n34210,
    n34211, n34212, n34213, n34214, n34215, n34216,
    n34217, n34218, n34219, n34220, n34221, n34222,
    n34223, n34224, n34225, n34226, n34227, n34228,
    n34229, n34230, n34231, n34232, n34233, n34234,
    n34235, n34236, n34237, n34238, n34239, n34240,
    n34241, n34242, n34243, n34244, n34245, n34246,
    n34247, n34248, n34249, n34250, n34251, n34252,
    n34253, n34254, n34255, n34256, n34257, n34258,
    n34259, n34260, n34261, n34262, n34263, n34264,
    n34265, n34266, n34267, n34268, n34269, n34270,
    n34271, n34272, n34273, n34274, n34275, n34276,
    n34277, n34278, n34279, n34280, n34281, n34282,
    n34283, n34284, n34285, n34286, n34287, n34288,
    n34289, n34290, n34291, n34292, n34293, n34294,
    n34295, n34296, n34297, n34298, n34299, n34300,
    n34301, n34302, n34303, n34304, n34305, n34306,
    n34307, n34308, n34309, n34310, n34311, n34312,
    n34313, n34314, n34315, n34316, n34317, n34318,
    n34319, n34320, n34321, n34322, n34323, n34324,
    n34325, n34326, n34327, n34328, n34329, n34330,
    n34331, n34332, n34333, n34334, n34335, n34336,
    n34337, n34338, n34339, n34340, n34341, n34342,
    n34343, n34344, n34345, n34346, n34347, n34348,
    n34349, n34350, n34351, n34352, n34353, n34354,
    n34355, n34356, n34357, n34358, n34359, n34360,
    n34361, n34362, n34363, n34364, n34365, n34366,
    n34367, n34368, n34369, n34370, n34371, n34372,
    n34373, n34374, n34375, n34376, n34377, n34378,
    n34379, n34380, n34381, n34382, n34383, n34384,
    n34385, n34386, n34387, n34388, n34389, n34390,
    n34391, n34392, n34393, n34394, n34395, n34396,
    n34397, n34398, n34399, n34400, n34401, n34402,
    n34403, n34404, n34405, n34406, n34407, n34408,
    n34409, n34410, n34411, n34412, n34413, n34414,
    n34415, n34416, n34417, n34418, n34419, n34420,
    n34421, n34422, n34423, n34424, n34425, n34426,
    n34427, n34428, n34429, n34430, n34431, n34432,
    n34433, n34434, n34435, n34436, n34437, n34438,
    n34439, n34440, n34441, n34442, n34443, n34444,
    n34445, n34446, n34447, n34448, n34449, n34450,
    n34451, n34452, n34453, n34454, n34455, n34456,
    n34457, n34458, n34459, n34460, n34461, n34462,
    n34463, n34464, n34465, n34466, n34467, n34468,
    n34469, n34470, n34471, n34472, n34473, n34474,
    n34475, n34476, n34477, n34478, n34479, n34480,
    n34481, n34482, n34483, n34484, n34485, n34486,
    n34487, n34488, n34489, n34490, n34491, n34492,
    n34493, n34494, n34495, n34496, n34497, n34498,
    n34499, n34500, n34501, n34502, n34503, n34504,
    n34505, n34506, n34507, n34508, n34509, n34510,
    n34511, n34512, n34513, n34514, n34515, n34516,
    n34517, n34518, n34519, n34520, n34521, n34522,
    n34523, n34524, n34525, n34526, n34527, n34528,
    n34529, n34530, n34531, n34532, n34533, n34534,
    n34535, n34536, n34537, n34538, n34539, n34540,
    n34541, n34542, n34543, n34544, n34545, n34546,
    n34547, n34548, n34549, n34550, n34551, n34552,
    n34553, n34554, n34555, n34556, n34557, n34558,
    n34559, n34560, n34561, n34562, n34563, n34564,
    n34565, n34566, n34567, n34568, n34569, n34570,
    n34571, n34572, n34573, n34574, n34575, n34576,
    n34577, n34578, n34579, n34580, n34581, n34582,
    n34583, n34584, n34585, n34586, n34587, n34588,
    n34589, n34590, n34591, n34592, n34593, n34594,
    n34595, n34596, n34597, n34598, n34599, n34600,
    n34601, n34602, n34603, n34604, n34605, n34606,
    n34607, n34608, n34609, n34610, n34611, n34612,
    n34613, n34614, n34615, n34616, n34617, n34618,
    n34619, n34620, n34621, n34622, n34623, n34624,
    n34625, n34626, n34627, n34628, n34629, n34630,
    n34631, n34632, n34633, n34634, n34635, n34636,
    n34637, n34638, n34639, n34640, n34641, n34642,
    n34643, n34644, n34645, n34646, n34647, n34648,
    n34649, n34650, n34652, n34653, n34654, n34655,
    n34656, n34657, n34658, n34659, n34660, n34661,
    n34662, n34663, n34664, n34665, n34666, n34667,
    n34668, n34669, n34670, n34671, n34672, n34673,
    n34674, n34675, n34676, n34677, n34678, n34679,
    n34680, n34681, n34682, n34683, n34684, n34685,
    n34686, n34687, n34688, n34689, n34690, n34691,
    n34692, n34693, n34694, n34695, n34696, n34697,
    n34698, n34699, n34700, n34701, n34702, n34703,
    n34704, n34705, n34706, n34707, n34708, n34709,
    n34710, n34711, n34712, n34713, n34714, n34715,
    n34716, n34717, n34718, n34719, n34720, n34721,
    n34722, n34723, n34725, n34726, n34727, n34728,
    n34729, n34730, n34731, n34732, n34733, n34734,
    n34735, n34736, n34737, n34738, n34739, n34740,
    n34741, n34742, n34743, n34744, n34745, n34746,
    n34747, n34748, n34749, n34750, n34751, n34752,
    n34753, n34754, n34755, n34756, n34757, n34758,
    n34759, n34760, n34761, n34762, n34763, n34764,
    n34765, n34766, n34767, n34768, n34769, n34770,
    n34771, n34772, n34773, n34774, n34775, n34776,
    n34777, n34778, n34779, n34780, n34781, n34782,
    n34783, n34784, n34785, n34786, n34787, n34788,
    n34789, n34790, n34791, n34792, n34793, n34794,
    n34795, n34796, n34797, n34798, n34799, n34800,
    n34801, n34802, n34803, n34804, n34805, n34806,
    n34807, n34808, n34809, n34810, n34811, n34812,
    n34813, n34814, n34815, n34816, n34817, n34818,
    n34819, n34820, n34821, n34822, n34823, n34824,
    n34825, n34826, n34827, n34828, n34829, n34830,
    n34831, n34832, n34833, n34834, n34835, n34836,
    n34837, n34838, n34839, n34840, n34841, n34842,
    n34843, n34844, n34845, n34846, n34847, n34848,
    n34849, n34850, n34851, n34852, n34853, n34854,
    n34855, n34856, n34857, n34858, n34859, n34860,
    n34861, n34862, n34863, n34864, n34865, n34866,
    n34867, n34868, n34869, n34870, n34871, n34872,
    n34873, n34874, n34875, n34876, n34877, n34878,
    n34879, n34880, n34881, n34882, n34883, n34885,
    n34886, n34887, n34888, n34889, n34890, n34891,
    n34892, n34893, n34894, n34895, n34896, n34897,
    n34898, n34899, n34900, n34901, n34902, n34903,
    n34904, n34905, n34906, n34907, n34908, n34909,
    n34910, n34911, n34912, n34913, n34914, n34915,
    n34916, n34917, n34918, n34919, n34920, n34921,
    n34922, n34923, n34924, n34925, n34926, n34927,
    n34928, n34929, n34930, n34931, n34932, n34933,
    n34934, n34935, n34936, n34937, n34938, n34939,
    n34940, n34941, n34942, n34943, n34944, n34945,
    n34946, n34947, n34948, n34949, n34950, n34951,
    n34952, n34953, n34954, n34955, n34956, n34957,
    n34958, n34959, n34960, n34961, n34962, n34963,
    n34964, n34965, n34966, n34967, n34968, n34969,
    n34970, n34971, n34972, n34973, n34974, n34975,
    n34976, n34977, n34978, n34979, n34980, n34981,
    n34982, n34983, n34984, n34985, n34986, n34987,
    n34988, n34989, n34990, n34991, n34992, n34993,
    n34994, n34995, n34996, n34997, n34998, n34999,
    n35000, n35001, n35002, n35003, n35004, n35005,
    n35006, n35007, n35008, n35009, n35011, n35012,
    n35013, n35014, n35015, n35016, n35017, n35018,
    n35019, n35020, n35021, n35022, n35023, n35024,
    n35025, n35026, n35027, n35028, n35029, n35030,
    n35031, n35032, n35033, n35034, n35035, n35036,
    n35038, n35039, n35040, n35041, n35042, n35043,
    n35044, n35045, n35046, n35047, n35048, n35049,
    n35050, n35051, n35052, n35053, n35054, n35055,
    n35056, n35057, n35059, n35060, n35061, n35062,
    n35063, n35064, n35065, n35066, n35067, n35068,
    n35069, n35070, n35071, n35072, n35073, n35074,
    n35075, n35076, n35077, n35078, n35080, n35081,
    n35082, n35083, n35084, n35085, n35086, n35087,
    n35088, n35089, n35090, n35091, n35092, n35093,
    n35094, n35095, n35096, n35097, n35098, n35099,
    n35101, n35102, n35103, n35104, n35105, n35106,
    n35107, n35108, n35109, n35110, n35111, n35112,
    n35113, n35114, n35115, n35116, n35117, n35118,
    n35119, n35120, n35121, n35122, n35123, n35124,
    n35125, n35126, n35127, n35128, n35129, n35130,
    n35131, n35132, n35133, n35134, n35135, n35136,
    n35137, n35138, n35139, n35140, n35141, n35142,
    n35143, n35144, n35145, n35146, n35147, n35148,
    n35149, n35150, n35151, n35152, n35153, n35154,
    n35155, n35156, n35157, n35158, n35159, n35160,
    n35161, n35162, n35163, n35164, n35165, n35166,
    n35167, n35168, n35169, n35170, n35171, n35172,
    n35173, n35174, n35175, n35176, n35177, n35178,
    n35179, n35180, n35181, n35182, n35183, n35184,
    n35185, n35186, n35187, n35188, n35189, n35190,
    n35191, n35192, n35193, n35194, n35195, n35196,
    n35197, n35198, n35199, n35200, n35201, n35202,
    n35203, n35204, n35205, n35206, n35207, n35208,
    n35209, n35211, n35212, n35213, n35214, n35215,
    n35216, n35217, n35218, n35219, n35220, n35221,
    n35222, n35223, n35224, n35225, n35226, n35227,
    n35228, n35229, n35230, n35231, n35232, n35233,
    n35234, n35235, n35236, n35237, n35238, n35239,
    n35240, n35241, n35242, n35243, n35244, n35245,
    n35246, n35247, n35248, n35249, n35250, n35251,
    n35252, n35253, n35254, n35255, n35256, n35257,
    n35258, n35259, n35260, n35261, n35262, n35263,
    n35264, n35265, n35266, n35267, n35268, n35269,
    n35270, n35271, n35272, n35273, n35274, n35275,
    n35276, n35277, n35278, n35279, n35280, n35281,
    n35282, n35283, n35284, n35285, n35286, n35287,
    n35288, n35289, n35290, n35291, n35292, n35293,
    n35294, n35295, n35296, n35297, n35298, n35299,
    n35300, n35301, n35302, n35303, n35304, n35305,
    n35306, n35307, n35309, n35310, n35311, n35312,
    n35313, n35314, n35315, n35316, n35317, n35318,
    n35319, n35320, n35321, n35322, n35323, n35324,
    n35325, n35326, n35328, n35329, n35330, n35331,
    n35332, n35333, n35335, n35336, n35337, n35338,
    n35339, n35340, n35341, n35342, n35343, n35344,
    n35345, n35346, n35347, n35348, n35349, n35350,
    n35351, n35352, n35353, n35354, n35356, n35357,
    n35358, n35359, n35360, n35361, n35363, n35364,
    n35365, n35366, n35367, n35368, n35369, n35370,
    n35371, n35372, n35373, n35374, n35375, n35376,
    n35377, n35378, n35379, n35380, n35381, n35382,
    n35383, n35384, n35385, n35386, n35387, n35388,
    n35389, n35390, n35391, n35392, n35393, n35394,
    n35395, n35396, n35397, n35398, n35399, n35400,
    n35401, n35402, n35403, n35404, n35405, n35406,
    n35407, n35408, n35409, n35410, n35411, n35412,
    n35413, n35414, n35415, n35416, n35417, n35418,
    n35419, n35420, n35421, n35422, n35423, n35424,
    n35425, n35426, n35427, n35428, n35429, n35430,
    n35431, n35432, n35433, n35434, n35435, n35436,
    n35437, n35438, n35439, n35440, n35441, n35442,
    n35443, n35444, n35445, n35446, n35447, n35448,
    n35449, n35450, n35451, n35452, n35453, n35454,
    n35455, n35456, n35457, n35458, n35459, n35460,
    n35461, n35462, n35463, n35464, n35465, n35466,
    n35468, n35469, n35470, n35471, n35472, n35473,
    n35474, n35475, n35476, n35477, n35478, n35479,
    n35480, n35481, n35482, n35483, n35484, n35485,
    n35486, n35487, n35488, n35489, n35490, n35491,
    n35492, n35493, n35494, n35495, n35496, n35497,
    n35498, n35499, n35500, n35501, n35502, n35503,
    n35504, n35505, n35506, n35507, n35508, n35509,
    n35510, n35511, n35512, n35513, n35514, n35515,
    n35516, n35517, n35518, n35519, n35520, n35521,
    n35522, n35523, n35524, n35525, n35526, n35527,
    n35528, n35529, n35530, n35531, n35532, n35533,
    n35534, n35535, n35536, n35537, n35538, n35539,
    n35540, n35541, n35542, n35543, n35544, n35545,
    n35546, n35547, n35548, n35549, n35550, n35551,
    n35552, n35553, n35554, n35555, n35556, n35557,
    n35558, n35559, n35560, n35561, n35562, n35563,
    n35564, n35565, n35566, n35567, n35568, n35569,
    n35570, n35571, n35572, n35573, n35574, n35575,
    n35576, n35577, n35578, n35579, n35580, n35581,
    n35582, n35583, n35584, n35585, n35586, n35587,
    n35588, n35589, n35590, n35591, n35592, n35593,
    n35594, n35595, n35596, n35597, n35598, n35599,
    n35600, n35601, n35602, n35603, n35604, n35605,
    n35606, n35607, n35608, n35609, n35610, n35611,
    n35612, n35613, n35614, n35615, n35616, n35617,
    n35618, n35619, n35620, n35621, n35622, n35623,
    n35624, n35625, n35626, n35627, n35628, n35629,
    n35630, n35631, n35632, n35633, n35634, n35635,
    n35636, n35637, n35638, n35639, n35640, n35641,
    n35642, n35643, n35644, n35645, n35646, n35647,
    n35648, n35649, n35650, n35651, n35652, n35653,
    n35654, n35655, n35656, n35657, n35658, n35659,
    n35660, n35661, n35662, n35663, n35664, n35665,
    n35666, n35667, n35668, n35669, n35670, n35671,
    n35672, n35673, n35674, n35675, n35676, n35677,
    n35678, n35679, n35680, n35681, n35682, n35683,
    n35684, n35685, n35686, n35687, n35688, n35689,
    n35690, n35691, n35692, n35693, n35694, n35695,
    n35696, n35697, n35698, n35699, n35700, n35701,
    n35702, n35703, n35704, n35705, n35706, n35707,
    n35708, n35709, n35710, n35711, n35712, n35713,
    n35714, n35715, n35716, n35717, n35718, n35719,
    n35720, n35721, n35722, n35723, n35724, n35725,
    n35726, n35727, n35728, n35729, n35730, n35731,
    n35732, n35733, n35734, n35735, n35736, n35737,
    n35738, n35739, n35740, n35741, n35742, n35743,
    n35744, n35745, n35746, n35747, n35748, n35749,
    n35750, n35751, n35752, n35753, n35754, n35755,
    n35756, n35757, n35758, n35759, n35760, n35761,
    n35762, n35763, n35764, n35765, n35766, n35767,
    n35768, n35769, n35770, n35771, n35772, n35773,
    n35774, n35775, n35776, n35777, n35778, n35779,
    n35780, n35781, n35782, n35783, n35784, n35785,
    n35786, n35787, n35788, n35789, n35790, n35791,
    n35792, n35793, n35794, n35795, n35796, n35797,
    n35798, n35799, n35800, n35801, n35802, n35803,
    n35804, n35805, n35806, n35807, n35808, n35809,
    n35810, n35811, n35812, n35813, n35814, n35815,
    n35816, n35817, n35818, n35819, n35820, n35821,
    n35822, n35823, n35824, n35825, n35826, n35827,
    n35828, n35829, n35830, n35831, n35832, n35833,
    n35834, n35835, n35836, n35837, n35838, n35839,
    n35840, n35841, n35842, n35843, n35844, n35845,
    n35846, n35847, n35848, n35849, n35850, n35851,
    n35852, n35853, n35854, n35855, n35856, n35857,
    n35858, n35859, n35860, n35861, n35862, n35863,
    n35864, n35865, n35866, n35867, n35868, n35869,
    n35870, n35871, n35872, n35873, n35874, n35875,
    n35876, n35877, n35878, n35879, n35880, n35881,
    n35882, n35883, n35884, n35885, n35886, n35887,
    n35888, n35889, n35890, n35891, n35892, n35893,
    n35894, n35895, n35896, n35897, n35898, n35899,
    n35900, n35901, n35902, n35903, n35904, n35905,
    n35906, n35907, n35908, n35909, n35910, n35911,
    n35912, n35913, n35914, n35915, n35916, n35917,
    n35918, n35919, n35920, n35921, n35922, n35923,
    n35924, n35925, n35926, n35927, n35928, n35929,
    n35930, n35931, n35932, n35933, n35934, n35935,
    n35936, n35937, n35938, n35939, n35940, n35941,
    n35942, n35943, n35944, n35945, n35946, n35947,
    n35948, n35949, n35950, n35951, n35952, n35953,
    n35954, n35955, n35956, n35957, n35958, n35959,
    n35960, n35961, n35962, n35963, n35964, n35965,
    n35966, n35967, n35968, n35969, n35970, n35971,
    n35972, n35973, n35974, n35975, n35976, n35977,
    n35978, n35979, n35980, n35981, n35982, n35983,
    n35984, n35985, n35986, n35987, n35988, n35989,
    n35990, n35991, n35992, n35993, n35994, n35995,
    n35996, n35997, n35998, n35999, n36000, n36001,
    n36002, n36003, n36004, n36005, n36006, n36007,
    n36008, n36009, n36010, n36011, n36012, n36013,
    n36014, n36015, n36016, n36017, n36018, n36019,
    n36020, n36021, n36022, n36023, n36024, n36025,
    n36026, n36027, n36028, n36029, n36030, n36031,
    n36032, n36033, n36034, n36035, n36036, n36037,
    n36038, n36039, n36040, n36041, n36042, n36043,
    n36044, n36045, n36046, n36047, n36048, n36049,
    n36050, n36051, n36052, n36053, n36054, n36055,
    n36056, n36057, n36058, n36059, n36060, n36061,
    n36062, n36063, n36064, n36065, n36066, n36067,
    n36068, n36069, n36070, n36071, n36072, n36073,
    n36074, n36075, n36076, n36077, n36078, n36079,
    n36080, n36081, n36082, n36083, n36084, n36085,
    n36086, n36087, n36088, n36090, n36091, n36092,
    n36093, n36094, n36095, n36096, n36097, n36098,
    n36099, n36100, n36101, n36102, n36103, n36104,
    n36105, n36106, n36107, n36108, n36109, n36110,
    n36111, n36112, n36113, n36114, n36115, n36116,
    n36117, n36118, n36119, n36120, n36121, n36122,
    n36123, n36124, n36125, n36126, n36127, n36128,
    n36129, n36130, n36131, n36132, n36133, n36134,
    n36135, n36136, n36137, n36138, n36139, n36140,
    n36141, n36142, n36143, n36144, n36145, n36146,
    n36147, n36148, n36149, n36150, n36151, n36152,
    n36153, n36154, n36155, n36156, n36157, n36158,
    n36159, n36160, n36161, n36162, n36163, n36164,
    n36165, n36166, n36167, n36168, n36169, n36170,
    n36171, n36172, n36173, n36174, n36175, n36176,
    n36177, n36178, n36179, n36180, n36181, n36182,
    n36183, n36184, n36185, n36186, n36187, n36188,
    n36189, n36190, n36191, n36192, n36193, n36194,
    n36195, n36196, n36197, n36198, n36199, n36200,
    n36201, n36202, n36203, n36204, n36205, n36206,
    n36207, n36208, n36209, n36210, n36211, n36212,
    n36213, n36214, n36215, n36216, n36217, n36218,
    n36219, n36220, n36221, n36222, n36223, n36224,
    n36225, n36226, n36227, n36228, n36229, n36230,
    n36231, n36232, n36233, n36234, n36235, n36236,
    n36237, n36238, n36239, n36240, n36241, n36242,
    n36243, n36244, n36245, n36246, n36247, n36248,
    n36249, n36250, n36251, n36252, n36253, n36254,
    n36255, n36256, n36257, n36258, n36259, n36260,
    n36261, n36262, n36263, n36264, n36265, n36266,
    n36267, n36268, n36269, n36270, n36271, n36272,
    n36273, n36274, n36275, n36276, n36277, n36278,
    n36279, n36280, n36281, n36282, n36283, n36284,
    n36285, n36286, n36287, n36288, n36289, n36290,
    n36291, n36292, n36293, n36294, n36295, n36296,
    n36297, n36298, n36299, n36300, n36301, n36302,
    n36303, n36304, n36305, n36306, n36307, n36308,
    n36309, n36310, n36311, n36312, n36313, n36314,
    n36315, n36316, n36317, n36318, n36319, n36320,
    n36321, n36322, n36323, n36324, n36325, n36326,
    n36327, n36328, n36329, n36330, n36331, n36332,
    n36333, n36334, n36335, n36336, n36337, n36338,
    n36339, n36340, n36341, n36342, n36343, n36344,
    n36345, n36346, n36347, n36348, n36349, n36350,
    n36351, n36352, n36353, n36354, n36355, n36356,
    n36357, n36358, n36359, n36360, n36361, n36362,
    n36363, n36364, n36365, n36366, n36367, n36368,
    n36369, n36370, n36371, n36372, n36373, n36374,
    n36375, n36376, n36377, n36378, n36379, n36380,
    n36381, n36382, n36383, n36384, n36385, n36386,
    n36387, n36388, n36389, n36390, n36391, n36392,
    n36393, n36394, n36395, n36396, n36397, n36398,
    n36399, n36400, n36401, n36402, n36403, n36404,
    n36405, n36406, n36407, n36408, n36409, n36410,
    n36411, n36412, n36413, n36414, n36415, n36416,
    n36417, n36418, n36419, n36420, n36421, n36422,
    n36423, n36424, n36425, n36426, n36427, n36428,
    n36429, n36430, n36431, n36432, n36433, n36434,
    n36435, n36436, n36437, n36438, n36439, n36440,
    n36441, n36442, n36443, n36444, n36445, n36446,
    n36447, n36448, n36449, n36450, n36451, n36452,
    n36453, n36454, n36455, n36456, n36457, n36458,
    n36459, n36460, n36461, n36462, n36463, n36464,
    n36465, n36466, n36467, n36468, n36469, n36470,
    n36471, n36472, n36473, n36474, n36475, n36476,
    n36477, n36478, n36479, n36480, n36481, n36482,
    n36483, n36484, n36485, n36486, n36487, n36488,
    n36489, n36490, n36491, n36492, n36493, n36494,
    n36495, n36496, n36497, n36498, n36499, n36500,
    n36501, n36502, n36503, n36504, n36505, n36506,
    n36507, n36508, n36509, n36510, n36511, n36512,
    n36513, n36514, n36515, n36516, n36517, n36518,
    n36519, n36520, n36521, n36522, n36523, n36524,
    n36525, n36526, n36527, n36528, n36529, n36530,
    n36531, n36532, n36533, n36534, n36535, n36536,
    n36537, n36538, n36539, n36540, n36541, n36542,
    n36543, n36544, n36545, n36546, n36547, n36548,
    n36549, n36550, n36551, n36552, n36553, n36554,
    n36555, n36556, n36557, n36558, n36559, n36560,
    n36561, n36562, n36563, n36564, n36565, n36566,
    n36567, n36568, n36569, n36570, n36571, n36572,
    n36573, n36574, n36575, n36576, n36577, n36578,
    n36579, n36580, n36581, n36582, n36583, n36584,
    n36585, n36586, n36587, n36588, n36589, n36590,
    n36591, n36592, n36593, n36594, n36595, n36596,
    n36597, n36598, n36599, n36600, n36601, n36602,
    n36603, n36604, n36605, n36606, n36607, n36608,
    n36609, n36610, n36611, n36612, n36613, n36614,
    n36615, n36616, n36617, n36618, n36619, n36620,
    n36621, n36622, n36623, n36624, n36625, n36626,
    n36627, n36628, n36629, n36630, n36631, n36632,
    n36633, n36634, n36635, n36636, n36637, n36638,
    n36639, n36640, n36641, n36642, n36643, n36644,
    n36645, n36646, n36647, n36648, n36649, n36650,
    n36651, n36652, n36653, n36654, n36655, n36656,
    n36657, n36658, n36659, n36660, n36662, n36663,
    n36664, n36665, n36666, n36667, n36668, n36669,
    n36670, n36671, n36672, n36673, n36674, n36675,
    n36676, n36677, n36678, n36679, n36680, n36681,
    n36682, n36683, n36684, n36685, n36686, n36687,
    n36688, n36689, n36690, n36691, n36692, n36693,
    n36694, n36695, n36696, n36697, n36698, n36699,
    n36700, n36701, n36702, n36703, n36704, n36705,
    n36706, n36707, n36708, n36709, n36710, n36711,
    n36712, n36713, n36714, n36715, n36716, n36717,
    n36718, n36719, n36720, n36721, n36722, n36723,
    n36724, n36725, n36726, n36727, n36728, n36729,
    n36730, n36731, n36732, n36733, n36734, n36735,
    n36736, n36737, n36738, n36739, n36740, n36741,
    n36742, n36743, n36744, n36745, n36746, n36747,
    n36748, n36749, n36750, n36751, n36752, n36753,
    n36754, n36755, n36756, n36757, n36758, n36759,
    n36760, n36761, n36762, n36763, n36764, n36765,
    n36766, n36767, n36768, n36769, n36770, n36771,
    n36772, n36773, n36774, n36775, n36776, n36777,
    n36778, n36779, n36780, n36781, n36782, n36783,
    n36784, n36785, n36786, n36787, n36788, n36789,
    n36790, n36791, n36792, n36793, n36794, n36795,
    n36796, n36797, n36798, n36799, n36800, n36801,
    n36802, n36803, n36804, n36805, n36806, n36807,
    n36808, n36809, n36810, n36811, n36812, n36813,
    n36814, n36815, n36816, n36817, n36818, n36819,
    n36820, n36821, n36822, n36823, n36824, n36825,
    n36826, n36827, n36828, n36829, n36830, n36831,
    n36832, n36833, n36834, n36835, n36836, n36837,
    n36838, n36839, n36840, n36841, n36842, n36843,
    n36844, n36845, n36846, n36847, n36848, n36849,
    n36850, n36851, n36852, n36853, n36854, n36855,
    n36856, n36857, n36858, n36859, n36860, n36861,
    n36862, n36863, n36864, n36865, n36866, n36867,
    n36868, n36869, n36870, n36871, n36872, n36873,
    n36874, n36875, n36876, n36877, n36878, n36879,
    n36880, n36881, n36882, n36883, n36884, n36885,
    n36886, n36887, n36888, n36889, n36890, n36891,
    n36892, n36893, n36894, n36895, n36896, n36897,
    n36898, n36899, n36900, n36901, n36902, n36903,
    n36904, n36905, n36906, n36907, n36908, n36909,
    n36910, n36911, n36912, n36913, n36914, n36915,
    n36916, n36917, n36918, n36919, n36920, n36921,
    n36922, n36923, n36924, n36925, n36926, n36927,
    n36928, n36929, n36930, n36931, n36932, n36933,
    n36934, n36935, n36936, n36937, n36938, n36939,
    n36940, n36941, n36942, n36943, n36944, n36945,
    n36946, n36947, n36948, n36949, n36950, n36951,
    n36952, n36953, n36954, n36955, n36956, n36957,
    n36958, n36959, n36960, n36961, n36962, n36963,
    n36964, n36965, n36966, n36967, n36968, n36969,
    n36970, n36971, n36972, n36973, n36974, n36975,
    n36976, n36977, n36978, n36979, n36980, n36981,
    n36982, n36983, n36984, n36985, n36986, n36987,
    n36988, n36989, n36990, n36991, n36992, n36993,
    n36994, n36995, n36996, n36997, n36998, n36999,
    n37000, n37001, n37002, n37003, n37004, n37005,
    n37006, n37007, n37008, n37009, n37010, n37011,
    n37012, n37013, n37014, n37015, n37016, n37017,
    n37018, n37019, n37020, n37021, n37022, n37023,
    n37024, n37025, n37026, n37027, n37028, n37029,
    n37030, n37031, n37032, n37033, n37034, n37035,
    n37036, n37037, n37038, n37039, n37040, n37041,
    n37042, n37043, n37044, n37045, n37046, n37047,
    n37048, n37049, n37050, n37051, n37052, n37053,
    n37054, n37055, n37056, n37057, n37058, n37059,
    n37060, n37061, n37062, n37063, n37064, n37065,
    n37066, n37067, n37068, n37069, n37070, n37071,
    n37072, n37073, n37074, n37075, n37076, n37077,
    n37078, n37079, n37080, n37081, n37082, n37083,
    n37084, n37085, n37086, n37087, n37088, n37089,
    n37090, n37091, n37092, n37093, n37094, n37095,
    n37096, n37097, n37098, n37099, n37100, n37101,
    n37102, n37103, n37104, n37105, n37106, n37107,
    n37108, n37109, n37110, n37111, n37112, n37113,
    n37114, n37115, n37116, n37117, n37118, n37119,
    n37120, n37121, n37122, n37123, n37124, n37125,
    n37126, n37127, n37128, n37129, n37130, n37131,
    n37132, n37133, n37134, n37135, n37136, n37137,
    n37138, n37139, n37140, n37141, n37142, n37143,
    n37144, n37145, n37146, n37147, n37148, n37149,
    n37150, n37151, n37152, n37153, n37154, n37155,
    n37156, n37157, n37158, n37159, n37160, n37161,
    n37162, n37163, n37164, n37165, n37166, n37167,
    n37168, n37169, n37170, n37171, n37172, n37173,
    n37174, n37175, n37176, n37177, n37178, n37179,
    n37180, n37181, n37182, n37183, n37184, n37185,
    n37186, n37187, n37188, n37189, n37190, n37191,
    n37192, n37193, n37194, n37195, n37196, n37197,
    n37198, n37199, n37200, n37201, n37202, n37203,
    n37204, n37205, n37206, n37207, n37208, n37209,
    n37210, n37211, n37212, n37213, n37214, n37215,
    n37216, n37217, n37218, n37219, n37220, n37221,
    n37222, n37223, n37224, n37225, n37226, n37227,
    n37228, n37229, n37231, n37232, n37233, n37234,
    n37235, n37236, n37237, n37238, n37239, n37240,
    n37241, n37242, n37243, n37244, n37245, n37246,
    n37247, n37248, n37249, n37250, n37251, n37252,
    n37253, n37254, n37255, n37256, n37257, n37258,
    n37259, n37260, n37261, n37262, n37263, n37264,
    n37265, n37266, n37267, n37268, n37269, n37270,
    n37271, n37272, n37273, n37274, n37275, n37276,
    n37277, n37278, n37279, n37280, n37281, n37282,
    n37283, n37284, n37285, n37286, n37287, n37288,
    n37289, n37290, n37291, n37292, n37293, n37294,
    n37295, n37296, n37297, n37298, n37299, n37300,
    n37301, n37302, n37303, n37304, n37305, n37306,
    n37307, n37308, n37309, n37310, n37311, n37312,
    n37313, n37314, n37315, n37316, n37317, n37318,
    n37319, n37320, n37321, n37322, n37323, n37324,
    n37325, n37326, n37327, n37328, n37329, n37330,
    n37331, n37332, n37333, n37334, n37335, n37336,
    n37337, n37338, n37339, n37340, n37341, n37342,
    n37343, n37344, n37345, n37346, n37347, n37348,
    n37349, n37350, n37351, n37352, n37353, n37354,
    n37356, n37357, n37358, n37359, n37360, n37361,
    n37362, n37363, n37364, n37365, n37366, n37367,
    n37368, n37369, n37370, n37371, n37372, n37373,
    n37374, n37375, n37376, n37377, n37378, n37379,
    n37380, n37381, n37382, n37383, n37384, n37385,
    n37386, n37387, n37388, n37389, n37390, n37391,
    n37392, n37393, n37394, n37395, n37396, n37397,
    n37398, n37399, n37400, n37401, n37402, n37403,
    n37404, n37405, n37406, n37407, n37408, n37410,
    n37411, n37412, n37413, n37414, n37415, n37416,
    n37417, n37418, n37419, n37420, n37421, n37422,
    n37423, n37424, n37425, n37426, n37427, n37428,
    n37429, n37430, n37431, n37432, n37433, n37434,
    n37435, n37436, n37437, n37438, n37440, n37441,
    n37442, n37443, n37444, n37445, n37446, n37447,
    n37448, n37449, n37451, n37452, n37453, n37454,
    n37455, n37456, n37457, n37458, n37459, n37460,
    n37461, n37462, n37463, n37464, n37465, n37466,
    n37467, n37468, n37469, n37470, n37471, n37472,
    n37473, n37474, n37475, n37476, n37477, n37478,
    n37479, n37480, n37481, n37482, n37483, n37484,
    n37485, n37486, n37487, n37488, n37489, n37490,
    n37491, n37492, n37493, n37494, n37495, n37496,
    n37497, n37498, n37499, n37500, n37501, n37502,
    n37503, n37504, n37505, n37506, n37507, n37508,
    n37509, n37510, n37511, n37512, n37513, n37514,
    n37515, n37516, n37517, n37518, n37519, n37520,
    n37521, n37522, n37523, n37524, n37525, n37526,
    n37527, n37528, n37529, n37530, n37531, n37533,
    n37534, n37535, n37536, n37537, n37538, n37539,
    n37540, n37541, n37542, n37543, n37544, n37545,
    n37546, n37547, n37548, n37549, n37550, n37551,
    n37552, n37553, n37554, n37555, n37556, n37557,
    n37558, n37559, n37560, n37561, n37562, n37563,
    n37564, n37565, n37566, n37567, n37568, n37570,
    n37571, n37572, n37573, n37574, n37575, n37576,
    n37577, n37578, n37579, n37580, n37581, n37582,
    n37583, n37584, n37585, n37586, n37587, n37588,
    n37589, n37590, n37591, n37593, n37594, n37595,
    n37596, n37597, n37598, n37599, n37600, n37601,
    n37602, n37603, n37604, n37605, n37606, n37607,
    n37608, n37609, n37610, n37611, n37612, n37613,
    n37614, n37615, n37616, n37617, n37618, n37619,
    n37620, n37621, n37622, n37623, n37624, n37625,
    n37626, n37627, n37628, n37629, n37630, n37631,
    n37632, n37633, n37634, n37635, n37636, n37637,
    n37638, n37639, n37640, n37641, n37642, n37643,
    n37644, n37645, n37646, n37647, n37648, n37649,
    n37650, n37651, n37652, n37653, n37654, n37655,
    n37656, n37657, n37658, n37659, n37660, n37661,
    n37662, n37663, n37664, n37665, n37666, n37667,
    n37668, n37669, n37670, n37671, n37672, n37673,
    n37674, n37675, n37676, n37677, n37678, n37679,
    n37680, n37681, n37682, n37683, n37684, n37685,
    n37686, n37687, n37688, n37689, n37690, n37691,
    n37692, n37693, n37694, n37695, n37696, n37697,
    n37698, n37699, n37700, n37701, n37702, n37703,
    n37704, n37705, n37706, n37707, n37708, n37709,
    n37710, n37711, n37712, n37713, n37714, n37715,
    n37716, n37717, n37718, n37719, n37720, n37721,
    n37722, n37723, n37724, n37725, n37726, n37727,
    n37728, n37729, n37730, n37731, n37732, n37733,
    n37734, n37735, n37736, n37737, n37738, n37739,
    n37740, n37741, n37742, n37743, n37744, n37745,
    n37746, n37747, n37748, n37749, n37750, n37751,
    n37752, n37753, n37754, n37755, n37756, n37757,
    n37758, n37759, n37760, n37761, n37762, n37763,
    n37764, n37765, n37766, n37767, n37768, n37769,
    n37770, n37771, n37772, n37773, n37774, n37775,
    n37776, n37777, n37778, n37779, n37780, n37781,
    n37782, n37783, n37784, n37785, n37786, n37787,
    n37788, n37789, n37790, n37791, n37792, n37793,
    n37794, n37795, n37796, n37797, n37798, n37799,
    n37800, n37801, n37802, n37803, n37804, n37805,
    n37806, n37807, n37808, n37809, n37810, n37811,
    n37812, n37813, n37814, n37815, n37816, n37817,
    n37818, n37819, n37820, n37821, n37822, n37823,
    n37824, n37825, n37826, n37827, n37828, n37829,
    n37830, n37831, n37832, n37833, n37834, n37835,
    n37836, n37837, n37838, n37839, n37840, n37841,
    n37842, n37843, n37844, n37845, n37846, n37847,
    n37848, n37849, n37850, n37851, n37852, n37853,
    n37854, n37855, n37856, n37857, n37858, n37859,
    n37860, n37861, n37862, n37863, n37864, n37865,
    n37866, n37867, n37868, n37869, n37870, n37871,
    n37872, n37873, n37874, n37875, n37876, n37877,
    n37878, n37879, n37880, n37881, n37882, n37883,
    n37884, n37885, n37886, n37887, n37888, n37889,
    n37890, n37891, n37892, n37893, n37894, n37895,
    n37896, n37897, n37898, n37899, n37900, n37901,
    n37902, n37903, n37904, n37905, n37906, n37907,
    n37908, n37909, n37910, n37911, n37912, n37913,
    n37914, n37915, n37916, n37917, n37918, n37919,
    n37920, n37921, n37922, n37923, n37924, n37925,
    n37926, n37927, n37928, n37929, n37930, n37931,
    n37932, n37933, n37934, n37935, n37936, n37937,
    n37938, n37939, n37940, n37941, n37942, n37943,
    n37944, n37945, n37946, n37947, n37948, n37949,
    n37950, n37951, n37952, n37953, n37954, n37956,
    n37957, n37958, n37959, n37960, n37961, n37962,
    n37963, n37964, n37965, n37966, n37967, n37968,
    n37969, n37970, n37971, n37972, n37973, n37974,
    n37975, n37976, n37977, n37978, n37979, n37980,
    n37981, n37982, n37983, n37984, n37985, n37986,
    n37987, n37988, n37989, n37990, n37991, n37992,
    n37993, n37994, n37995, n37996, n37997, n37998,
    n37999, n38000, n38001, n38002, n38003, n38004,
    n38005, n38006, n38007, n38008, n38009, n38010,
    n38011, n38012, n38013, n38014, n38015, n38016,
    n38017, n38018, n38019, n38020, n38021, n38022,
    n38023, n38024, n38025, n38026, n38027, n38028,
    n38029, n38030, n38031, n38032, n38033, n38034,
    n38035, n38036, n38037, n38038, n38039, n38040,
    n38041, n38042, n38043, n38044, n38045, n38046,
    n38047, n38048, n38049, n38050, n38051, n38052,
    n38053, n38054, n38055, n38056, n38057, n38058,
    n38059, n38060, n38061, n38062, n38063, n38064,
    n38065, n38066, n38067, n38068, n38069, n38070,
    n38071, n38072, n38073, n38074, n38075, n38076,
    n38077, n38078, n38079, n38080, n38081, n38082,
    n38083, n38084, n38085, n38086, n38087, n38088,
    n38089, n38090, n38091, n38092, n38093, n38094,
    n38095, n38096, n38097, n38098, n38099, n38100,
    n38101, n38102, n38103, n38104, n38105, n38106,
    n38107, n38108, n38109, n38110, n38111, n38112,
    n38113, n38114, n38115, n38116, n38117, n38118,
    n38119, n38120, n38121, n38122, n38123, n38124,
    n38125, n38126, n38127, n38128, n38129, n38130,
    n38131, n38132, n38133, n38134, n38135, n38136,
    n38137, n38138, n38139, n38140, n38141, n38142,
    n38143, n38144, n38145, n38146, n38147, n38148,
    n38149, n38150, n38151, n38152, n38153, n38154,
    n38155, n38156, n38157, n38158, n38159, n38160,
    n38161, n38162, n38163, n38164, n38165, n38166,
    n38167, n38168, n38169, n38170, n38171, n38172,
    n38173, n38174, n38175, n38176, n38177, n38178,
    n38179, n38180, n38181, n38182, n38183, n38184,
    n38185, n38186, n38187, n38188, n38189, n38190,
    n38191, n38192, n38193, n38194, n38195, n38196,
    n38197, n38198, n38199, n38200, n38201, n38202,
    n38203, n38204, n38205, n38206, n38207, n38208,
    n38209, n38210, n38211, n38212, n38213, n38214,
    n38215, n38216, n38217, n38218, n38219, n38220,
    n38221, n38222, n38223, n38224, n38225, n38226,
    n38227, n38228, n38229, n38230, n38231, n38232,
    n38233, n38234, n38235, n38236, n38237, n38238,
    n38240, n38241, n38242, n38243, n38244, n38245,
    n38246, n38247, n38248, n38249, n38250, n38251,
    n38252, n38253, n38254, n38255, n38256, n38257,
    n38258, n38259, n38260, n38261, n38262, n38263,
    n38264, n38265, n38266, n38267, n38268, n38269,
    n38270, n38271, n38272, n38273, n38274, n38275,
    n38276, n38277, n38278, n38279, n38280, n38281,
    n38282, n38283, n38284, n38285, n38286, n38287,
    n38288, n38289, n38290, n38291, n38292, n38293,
    n38294, n38295, n38296, n38297, n38298, n38299,
    n38300, n38301, n38302, n38303, n38304, n38305,
    n38306, n38307, n38308, n38309, n38310, n38311,
    n38312, n38313, n38314, n38315, n38316, n38317,
    n38318, n38319, n38320, n38321, n38322, n38323,
    n38324, n38325, n38326, n38327, n38328, n38329,
    n38330, n38331, n38332, n38333, n38334, n38335,
    n38336, n38337, n38338, n38339, n38340, n38341,
    n38342, n38343, n38344, n38345, n38346, n38347,
    n38348, n38349, n38350, n38351, n38352, n38353,
    n38354, n38355, n38356, n38357, n38358, n38359,
    n38360, n38361, n38362, n38363, n38364, n38365,
    n38366, n38367, n38368, n38369, n38370, n38371,
    n38372, n38373, n38374, n38375, n38376, n38377,
    n38378, n38379, n38380, n38381, n38382, n38383,
    n38384, n38385, n38386, n38387, n38388, n38389,
    n38390, n38391, n38392, n38393, n38394, n38395,
    n38396, n38397, n38398, n38399, n38400, n38401,
    n38402, n38403, n38404, n38405, n38406, n38407,
    n38408, n38409, n38410, n38411, n38412, n38413,
    n38414, n38415, n38416, n38417, n38418, n38419,
    n38420, n38421, n38422, n38423, n38424, n38425,
    n38426, n38427, n38428, n38429, n38430, n38431,
    n38432, n38433, n38434, n38436, n38437, n38438,
    n38439, n38440, n38441, n38442, n38443, n38444,
    n38445, n38446, n38447, n38449, n38450, n38451,
    n38452, n38453, n38454, n38455, n38456, n38457,
    n38458, n38459, n38460, n38461, n38462, n38463,
    n38464, n38465, n38466, n38467, n38468, n38469,
    n38470, n38471, n38472, n38473, n38474, n38475,
    n38476, n38477, n38478, n38479, n38480, n38481,
    n38482, n38483, n38484, n38485, n38486, n38487,
    n38488, n38489, n38490, n38491, n38492, n38493,
    n38494, n38495, n38496, n38497, n38498, n38499,
    n38500, n38501, n38502, n38503, n38504, n38505,
    n38506, n38507, n38508, n38509, n38510, n38511,
    n38512, n38513, n38514, n38515, n38516, n38517,
    n38518, n38519, n38520, n38521, n38522, n38523,
    n38524, n38525, n38526, n38527, n38528, n38529,
    n38530, n38531, n38532, n38533, n38534, n38535,
    n38536, n38537, n38538, n38539, n38540, n38541,
    n38542, n38543, n38544, n38545, n38546, n38547,
    n38548, n38549, n38550, n38551, n38552, n38553,
    n38554, n38555, n38556, n38557, n38558, n38559,
    n38560, n38561, n38562, n38563, n38564, n38565,
    n38566, n38567, n38568, n38569, n38570, n38571,
    n38572, n38573, n38574, n38575, n38576, n38577,
    n38578, n38579, n38580, n38581, n38582, n38583,
    n38584, n38585, n38586, n38587, n38588, n38589,
    n38590, n38591, n38592, n38593, n38594, n38595,
    n38596, n38597, n38598, n38599, n38600, n38601,
    n38602, n38603, n38604, n38605, n38606, n38607,
    n38608, n38609, n38610, n38611, n38612, n38613,
    n38614, n38615, n38616, n38617, n38618, n38619,
    n38620, n38621, n38622, n38623, n38624, n38625,
    n38626, n38627, n38628, n38629, n38630, n38631,
    n38632, n38633, n38634, n38635, n38636, n38637,
    n38638, n38639, n38640, n38641, n38642, n38643,
    n38644, n38645, n38646, n38647, n38648, n38649,
    n38650, n38651, n38652, n38653, n38654, n38655,
    n38656, n38657, n38658, n38659, n38660, n38661,
    n38662, n38663, n38664, n38665, n38666, n38667,
    n38668, n38669, n38670, n38671, n38672, n38673,
    n38674, n38675, n38676, n38677, n38678, n38679,
    n38680, n38681, n38682, n38683, n38684, n38685,
    n38686, n38687, n38688, n38689, n38690, n38691,
    n38692, n38693, n38694, n38695, n38697, n38698,
    n38699, n38700, n38701, n38702, n38703, n38704,
    n38705, n38706, n38707, n38708, n38709, n38710,
    n38711, n38712, n38713, n38714, n38715, n38716,
    n38717, n38718, n38719, n38720, n38721, n38722,
    n38723, n38724, n38725, n38726, n38727, n38728,
    n38729, n38730, n38731, n38732, n38733, n38734,
    n38735, n38736, n38737, n38738, n38739, n38740,
    n38741, n38742, n38743, n38744, n38745, n38746,
    n38747, n38748, n38749, n38750, n38751, n38752,
    n38753, n38754, n38755, n38756, n38757, n38758,
    n38759, n38760, n38761, n38762, n38763, n38764,
    n38765, n38766, n38767, n38768, n38769, n38770,
    n38771, n38772, n38773, n38774, n38775, n38776,
    n38777, n38778, n38779, n38780, n38781, n38782,
    n38783, n38784, n38785, n38786, n38787, n38788,
    n38789, n38790, n38791, n38792, n38793, n38794,
    n38795, n38796, n38797, n38798, n38799, n38800,
    n38801, n38802, n38803, n38804, n38805, n38806,
    n38807, n38808, n38809, n38810, n38811, n38812,
    n38813, n38814, n38815, n38816, n38817, n38818,
    n38819, n38820, n38821, n38822, n38823, n38824,
    n38825, n38826, n38827, n38828, n38829, n38830,
    n38831, n38832, n38833, n38834, n38835, n38836,
    n38837, n38838, n38839, n38840, n38841, n38842,
    n38843, n38844, n38845, n38846, n38847, n38848,
    n38849, n38850, n38851, n38852, n38853, n38854,
    n38855, n38856, n38857, n38858, n38859, n38860,
    n38861, n38862, n38863, n38864, n38865, n38866,
    n38867, n38868, n38869, n38870, n38871, n38872,
    n38873, n38874, n38875, n38876, n38877, n38878,
    n38879, n38880, n38881, n38882, n38883, n38884,
    n38885, n38886, n38887, n38888, n38889, n38890,
    n38891, n38892, n38893, n38894, n38895, n38896,
    n38897, n38898, n38899, n38900, n38901, n38902,
    n38903, n38904, n38905, n38906, n38907, n38908,
    n38909, n38910, n38911, n38912, n38913, n38914,
    n38915, n38916, n38917, n38918, n38919, n38920,
    n38921, n38922, n38923, n38924, n38925, n38926,
    n38927, n38928, n38929, n38930, n38931, n38932,
    n38933, n38934, n38935, n38936, n38937, n38938,
    n38939, n38940, n38941, n38942, n38943, n38944,
    n38945, n38946, n38947, n38948, n38949, n38950,
    n38951, n38952, n38953, n38954, n38955, n38956,
    n38957, n38958, n38959, n38960, n38961, n38962,
    n38963, n38964, n38965, n38966, n38967, n38968,
    n38969, n38970, n38971, n38972, n38973, n38974,
    n38975, n38976, n38977, n38978, n38979, n38980,
    n38981, n38982, n38983, n38984, n38985, n38986,
    n38987, n38988, n38989, n38990, n38991, n38992,
    n38993, n38995, n38996, n38997, n38998, n38999,
    n39000, n39001, n39002, n39003, n39004, n39005,
    n39006, n39007, n39008, n39009, n39010, n39011,
    n39012, n39013, n39014, n39015, n39016, n39017,
    n39018, n39019, n39020, n39021, n39022, n39023,
    n39024, n39025, n39026, n39027, n39028, n39029,
    n39030, n39031, n39032, n39033, n39034, n39035,
    n39036, n39037, n39038, n39039, n39040, n39041,
    n39042, n39043, n39044, n39045, n39046, n39047,
    n39048, n39049, n39050, n39051, n39052, n39053,
    n39054, n39055, n39056, n39057, n39058, n39059,
    n39060, n39061, n39062, n39063, n39064, n39065,
    n39066, n39067, n39068, n39069, n39070, n39071,
    n39072, n39073, n39074, n39075, n39076, n39077,
    n39079, n39080, n39081, n39082, n39083, n39084,
    n39085, n39086, n39087, n39088, n39089, n39090,
    n39091, n39092, n39093, n39094, n39095, n39096,
    n39097, n39098, n39099, n39100, n39101, n39102,
    n39103, n39104, n39105, n39106, n39107, n39108,
    n39109, n39110, n39111, n39112, n39113, n39114,
    n39115, n39116, n39117, n39118, n39119, n39120,
    n39121, n39122, n39123, n39124, n39125, n39126,
    n39127, n39128, n39129, n39130, n39131, n39132,
    n39133, n39134, n39135, n39136, n39137, n39138,
    n39139, n39140, n39141, n39142, n39143, n39144,
    n39145, n39146, n39147, n39148, n39149, n39150,
    n39151, n39152, n39153, n39154, n39155, n39156,
    n39157, n39158, n39159, n39160, n39161, n39162,
    n39163, n39164, n39165, n39166, n39167, n39168,
    n39169, n39170, n39171, n39172, n39173, n39174,
    n39175, n39176, n39177, n39178, n39179, n39180,
    n39181, n39182, n39183, n39184, n39185, n39186,
    n39187, n39188, n39189, n39190, n39191, n39192,
    n39193, n39194, n39195, n39196, n39197, n39198,
    n39199, n39200, n39201, n39202, n39203, n39204,
    n39205, n39206, n39207, n39208, n39209, n39210,
    n39211, n39212, n39213, n39214, n39215, n39216,
    n39217, n39218, n39219, n39220, n39221, n39222,
    n39223, n39224, n39225, n39226, n39227, n39228,
    n39229, n39230, n39231, n39232, n39233, n39234,
    n39235, n39236, n39237, n39238, n39239, n39240,
    n39241, n39242, n39243, n39244, n39245, n39246,
    n39247, n39248, n39249, n39250, n39251, n39252,
    n39253, n39254, n39255, n39256, n39257, n39258,
    n39259, n39260, n39261, n39262, n39263, n39264,
    n39265, n39266, n39267, n39268, n39269, n39270,
    n39271, n39272, n39273, n39274, n39275, n39276,
    n39277, n39278, n39279, n39280, n39281, n39282,
    n39283, n39284, n39285, n39286, n39287, n39288,
    n39289, n39290, n39291, n39292, n39293, n39294,
    n39295, n39296, n39297, n39298, n39299, n39300,
    n39301, n39302, n39303, n39304, n39305, n39306,
    n39307, n39308, n39309, n39310, n39311, n39312,
    n39313, n39314, n39315, n39316, n39317, n39318,
    n39319, n39320, n39321, n39322, n39323, n39324,
    n39325, n39326, n39327, n39328, n39329, n39330,
    n39331, n39332, n39333, n39334, n39335, n39336,
    n39337, n39338, n39339, n39340, n39341, n39342,
    n39343, n39344, n39345, n39346, n39347, n39348,
    n39349, n39350, n39351, n39352, n39353, n39354,
    n39355, n39356, n39357, n39358, n39359, n39360,
    n39361, n39362, n39363, n39364, n39365, n39366,
    n39367, n39368, n39369, n39370, n39371, n39372,
    n39373, n39374, n39375, n39376, n39377, n39378,
    n39379, n39380, n39381, n39382, n39383, n39384,
    n39385, n39386, n39387, n39388, n39389, n39390,
    n39391, n39392, n39393, n39394, n39395, n39396,
    n39397, n39398, n39399, n39400, n39401, n39402,
    n39403, n39404, n39405, n39406, n39407, n39408,
    n39409, n39410, n39411, n39412, n39413, n39414,
    n39415, n39416, n39417, n39418, n39419, n39420,
    n39421, n39422, n39423, n39424, n39425, n39426,
    n39427, n39428, n39429, n39430, n39431, n39432,
    n39433, n39434, n39435, n39436, n39437, n39438,
    n39439, n39440, n39441, n39442, n39443, n39444,
    n39445, n39446, n39447, n39448, n39450, n39451,
    n39452, n39453, n39454, n39455, n39456, n39457,
    n39458, n39459, n39460, n39461, n39462, n39463,
    n39464, n39465, n39466, n39467, n39468, n39469,
    n39470, n39471, n39472, n39473, n39474, n39475,
    n39476, n39477, n39478, n39479, n39480, n39481,
    n39482, n39483, n39484, n39485, n39486, n39487,
    n39488, n39489, n39490, n39491, n39492, n39493,
    n39494, n39495, n39496, n39497, n39498, n39499,
    n39500, n39501, n39502, n39503, n39504, n39505,
    n39506, n39507, n39508, n39509, n39510, n39511,
    n39512, n39513, n39514, n39515, n39516, n39517,
    n39518, n39519, n39520, n39521, n39522, n39523,
    n39524, n39525, n39526, n39527, n39528, n39529,
    n39530, n39531, n39532, n39533, n39534, n39535,
    n39536, n39537, n39538, n39539, n39540, n39541,
    n39542, n39543, n39544, n39545, n39546, n39547,
    n39548, n39549, n39550, n39551, n39552, n39553,
    n39554, n39555, n39556, n39557, n39558, n39559,
    n39560, n39561, n39562, n39563, n39564, n39565,
    n39566, n39567, n39568, n39569, n39570, n39571,
    n39572, n39573, n39574, n39575, n39576, n39577,
    n39578, n39579, n39580, n39581, n39582, n39583,
    n39584, n39585, n39586, n39587, n39588, n39589,
    n39590, n39591, n39592, n39593, n39594, n39595,
    n39596, n39597, n39598, n39599, n39600, n39601,
    n39602, n39603, n39604, n39605, n39606, n39607,
    n39608, n39609, n39610, n39611, n39612, n39613,
    n39614, n39615, n39616, n39617, n39618, n39619,
    n39620, n39621, n39622, n39623, n39624, n39625,
    n39626, n39627, n39628, n39629, n39630, n39631,
    n39632, n39633, n39634, n39635, n39636, n39637,
    n39638, n39639, n39640, n39641, n39642, n39643,
    n39644, n39645, n39646, n39647, n39648, n39649,
    n39650, n39651, n39652, n39653, n39654, n39655,
    n39656, n39657, n39658, n39659, n39660, n39661,
    n39662, n39663, n39664, n39665, n39666, n39667,
    n39668, n39669, n39670, n39671, n39672, n39673,
    n39674, n39675, n39676, n39677, n39678, n39679,
    n39680, n39681, n39682, n39683, n39684, n39685,
    n39686, n39687, n39688, n39689, n39690, n39691,
    n39692, n39693, n39694, n39695, n39696, n39697,
    n39698, n39699, n39700, n39701, n39702, n39703,
    n39704, n39705, n39706, n39707, n39708, n39709,
    n39710, n39711, n39712, n39714, n39715, n39716,
    n39717, n39718, n39719, n39720, n39721, n39722,
    n39723, n39724, n39725, n39726, n39727, n39728,
    n39729, n39730, n39731, n39732, n39733, n39734,
    n39735, n39736, n39737, n39738, n39739, n39740,
    n39741, n39742, n39743, n39744, n39745, n39746,
    n39747, n39748, n39749, n39750, n39751, n39752,
    n39753, n39754, n39755, n39756, n39757, n39758,
    n39759, n39760, n39761, n39762, n39763, n39764,
    n39765, n39766, n39767, n39768, n39769, n39770,
    n39771, n39772, n39773, n39774, n39775, n39776,
    n39777, n39778, n39779, n39780, n39781, n39782,
    n39783, n39784, n39785, n39786, n39788, n39789,
    n39790, n39791, n39792, n39793, n39794, n39795,
    n39796, n39797, n39798, n39799, n39800, n39801,
    n39802, n39803, n39804, n39805, n39806, n39807,
    n39808, n39809, n39810, n39811, n39812, n39813,
    n39814, n39815, n39816, n39817, n39818, n39819,
    n39820, n39821, n39822, n39823, n39824, n39825,
    n39826, n39827, n39828, n39829, n39830, n39831,
    n39832, n39833, n39834, n39835, n39836, n39837,
    n39838, n39839, n39840, n39841, n39842, n39843,
    n39844, n39845, n39846, n39847, n39848, n39849,
    n39850, n39851, n39852, n39853, n39854, n39855,
    n39856, n39857, n39858, n39859, n39860, n39861,
    n39862, n39863, n39864, n39865, n39866, n39867,
    n39868, n39869, n39870, n39871, n39872, n39873,
    n39874, n39875, n39876, n39877, n39878, n39879,
    n39880, n39881, n39882, n39883, n39884, n39885,
    n39886, n39887, n39888, n39889, n39890, n39891,
    n39892, n39893, n39894, n39895, n39896, n39897,
    n39898, n39899, n39900, n39901, n39902, n39903,
    n39904, n39905, n39906, n39907, n39908, n39909,
    n39910, n39911, n39912, n39913, n39914, n39915,
    n39916, n39917, n39918, n39919, n39920, n39921,
    n39922, n39923, n39924, n39925, n39926, n39927,
    n39928, n39929, n39930, n39931, n39932, n39933,
    n39934, n39935, n39936, n39937, n39938, n39939,
    n39940, n39941, n39942, n39943, n39944, n39945,
    n39946, n39947, n39948, n39949, n39950, n39951,
    n39952, n39953, n39954, n39955, n39956, n39957,
    n39958, n39959, n39960, n39961, n39962, n39963,
    n39964, n39965, n39966, n39967, n39968, n39969,
    n39970, n39971, n39972, n39973, n39974, n39975,
    n39976, n39977, n39978, n39979, n39980, n39981,
    n39982, n39983, n39984, n39985, n39986, n39987,
    n39988, n39989, n39990, n39991, n39992, n39993,
    n39994, n39995, n39996, n39997, n39998, n39999,
    n40000, n40001, n40002, n40003, n40004, n40005,
    n40006, n40007, n40008, n40009, n40010, n40011,
    n40012, n40013, n40014, n40015, n40016, n40017,
    n40018, n40019, n40020, n40021, n40022, n40023,
    n40024, n40025, n40026, n40027, n40028, n40029,
    n40030, n40031, n40032, n40033, n40034, n40035,
    n40036, n40037, n40038, n40039, n40040, n40041,
    n40042, n40043, n40044, n40045, n40046, n40047,
    n40048, n40049, n40050, n40051, n40052, n40053,
    n40054, n40055, n40056, n40057, n40058, n40059,
    n40060, n40061, n40062, n40063, n40064, n40065,
    n40066, n40067, n40068, n40069, n40070, n40071,
    n40072, n40073, n40074, n40075, n40076, n40077,
    n40078, n40079, n40080, n40081, n40082, n40083,
    n40084, n40085, n40086, n40087, n40089, n40090,
    n40091, n40092, n40093, n40094, n40095, n40096,
    n40097, n40098, n40099, n40100, n40101, n40102,
    n40103, n40104, n40105, n40106, n40107, n40108,
    n40109, n40110, n40111, n40112, n40113, n40114,
    n40115, n40116, n40117, n40118, n40119, n40120,
    n40121, n40122, n40123, n40124, n40125, n40126,
    n40127, n40128, n40129, n40130, n40131, n40132,
    n40133, n40134, n40136, n40137, n40138, n40139,
    n40140, n40141, n40142, n40143, n40144, n40145,
    n40146, n40147, n40148, n40149, n40150, n40151,
    n40152, n40153, n40154, n40155, n40156, n40157,
    n40158, n40159, n40160, n40161, n40162, n40163,
    n40164, n40165, n40166, n40167, n40168, n40169,
    n40170, n40171, n40172, n40173, n40174, n40175,
    n40176, n40177, n40178, n40179, n40180, n40181,
    n40182, n40183, n40184, n40185, n40186, n40187,
    n40188, n40189, n40190, n40191, n40192, n40193,
    n40194, n40195, n40196, n40197, n40198, n40199,
    n40200, n40201, n40202, n40203, n40204, n40205,
    n40206, n40207, n40208, n40209, n40210, n40211,
    n40212, n40213, n40214, n40215, n40216, n40217,
    n40218, n40219, n40220, n40221, n40222, n40223,
    n40224, n40225, n40226, n40227, n40228, n40229,
    n40230, n40231, n40232, n40233, n40234, n40235,
    n40236, n40237, n40238, n40239, n40240, n40241,
    n40242, n40243, n40244, n40245, n40246, n40247,
    n40248, n40249, n40250, n40251, n40252, n40253,
    n40254, n40255, n40256, n40257, n40258, n40259,
    n40260, n40261, n40262, n40263, n40264, n40265,
    n40266, n40267, n40268, n40269, n40270, n40271,
    n40272, n40273, n40274, n40275, n40276, n40277,
    n40278, n40279, n40280, n40281, n40282, n40283,
    n40284, n40285, n40286, n40287, n40288, n40289,
    n40290, n40291, n40292, n40293, n40294, n40295,
    n40296, n40297, n40298, n40299, n40300, n40301,
    n40302, n40303, n40304, n40305, n40306, n40307,
    n40308, n40309, n40310, n40311, n40312, n40313,
    n40314, n40315, n40316, n40317, n40318, n40319,
    n40320, n40321, n40322, n40323, n40324, n40325,
    n40326, n40327, n40328, n40329, n40330, n40331,
    n40332, n40333, n40334, n40335, n40336, n40337,
    n40338, n40339, n40340, n40341, n40342, n40344,
    n40345, n40346, n40347, n40348, n40349, n40350,
    n40351, n40352, n40353, n40354, n40355, n40356,
    n40357, n40358, n40359, n40360, n40361, n40362,
    n40363, n40364, n40365, n40366, n40367, n40368,
    n40369, n40370, n40371, n40372, n40373, n40374,
    n40375, n40376, n40377, n40378, n40379, n40380,
    n40381, n40382, n40383, n40384, n40385, n40386,
    n40387, n40388, n40389, n40390, n40391, n40392,
    n40393, n40394, n40395, n40396, n40397, n40398,
    n40399, n40400, n40401, n40402, n40403, n40404,
    n40405, n40406, n40407, n40408, n40409, n40410,
    n40411, n40412, n40413, n40414, n40415, n40416,
    n40417, n40418, n40419, n40420, n40421, n40422,
    n40423, n40424, n40425, n40426, n40427, n40428,
    n40429, n40430, n40431, n40432, n40433, n40434,
    n40435, n40436, n40437, n40438, n40439, n40440,
    n40441, n40442, n40443, n40444, n40445, n40446,
    n40447, n40448, n40449, n40450, n40451, n40452,
    n40453, n40454, n40455, n40456, n40457, n40458,
    n40459, n40460, n40461, n40462, n40463, n40464,
    n40465, n40466, n40467, n40468, n40469, n40470,
    n40471, n40472, n40473, n40474, n40475, n40476,
    n40477, n40478, n40479, n40480, n40481, n40482,
    n40483, n40484, n40485, n40486, n40487, n40488,
    n40489, n40490, n40491, n40492, n40493, n40494,
    n40495, n40496, n40497, n40498, n40499, n40500,
    n40501, n40502, n40503, n40504, n40505, n40506,
    n40507, n40508, n40509, n40510, n40511, n40512,
    n40513, n40514, n40515, n40516, n40517, n40518,
    n40519, n40520, n40521, n40522, n40523, n40524,
    n40525, n40526, n40527, n40528, n40529, n40530,
    n40531, n40532, n40533, n40534, n40535, n40536,
    n40537, n40538, n40539, n40540, n40541, n40542,
    n40543, n40544, n40545, n40546, n40547, n40548,
    n40549, n40550, n40551, n40552, n40553, n40554,
    n40555, n40556, n40557, n40558, n40559, n40560,
    n40561, n40562, n40563, n40564, n40565, n40566,
    n40567, n40568, n40569, n40570, n40571, n40572,
    n40573, n40574, n40575, n40576, n40577, n40578,
    n40579, n40580, n40581, n40582, n40583, n40584,
    n40586, n40587, n40588, n40589, n40590, n40591,
    n40592, n40593, n40594, n40595, n40596, n40597,
    n40598, n40599, n40600, n40601, n40602, n40603,
    n40604, n40605, n40606, n40607, n40608, n40609,
    n40610, n40611, n40612, n40613, n40614, n40615,
    n40616, n40617, n40618, n40619, n40620, n40621,
    n40622, n40623, n40624, n40625, n40626, n40627,
    n40628, n40629, n40630, n40631, n40632, n40633,
    n40634, n40635, n40636, n40637, n40638, n40639,
    n40640, n40641, n40642, n40643, n40644, n40645,
    n40646, n40647, n40648, n40649, n40650, n40651,
    n40652, n40653, n40654, n40655, n40656, n40657,
    n40658, n40659, n40660, n40661, n40662, n40663,
    n40664, n40665, n40666, n40667, n40668, n40669,
    n40670, n40671, n40672, n40673, n40674, n40675,
    n40676, n40677, n40678, n40679, n40680, n40681,
    n40682, n40683, n40684, n40685, n40686, n40687,
    n40688, n40689, n40690, n40691, n40692, n40693,
    n40694, n40695, n40696, n40697, n40698, n40699,
    n40700, n40701, n40702, n40703, n40704, n40705,
    n40706, n40707, n40708, n40709, n40710, n40711,
    n40712, n40713, n40714, n40715, n40716, n40717,
    n40718, n40719, n40720, n40721, n40722, n40723,
    n40724, n40725, n40726, n40727, n40728, n40729,
    n40730, n40731, n40732, n40733, n40734, n40735,
    n40736, n40737, n40738, n40739, n40740, n40741,
    n40742, n40743, n40744, n40745, n40746, n40747,
    n40748, n40749, n40750, n40751, n40752, n40753,
    n40754, n40755, n40756, n40757, n40758, n40759,
    n40760, n40761, n40762, n40763, n40764, n40765,
    n40766, n40767, n40768, n40769, n40770, n40771,
    n40772, n40773, n40774, n40775, n40776, n40777,
    n40778, n40779, n40780, n40781, n40782, n40783,
    n40784, n40785, n40786, n40787, n40788, n40789,
    n40790, n40791, n40792, n40793, n40794, n40795,
    n40796, n40797, n40798, n40799, n40800, n40801,
    n40802, n40803, n40804, n40806, n40807, n40808,
    n40809, n40810, n40811, n40812, n40813, n40814,
    n40815, n40816, n40817, n40818, n40819, n40820,
    n40821, n40822, n40823, n40824, n40825, n40826,
    n40827, n40828, n40829, n40830, n40831, n40832,
    n40833, n40834, n40835, n40836, n40837, n40838,
    n40839, n40840, n40841, n40842, n40843, n40844,
    n40845, n40846, n40847, n40848, n40849, n40850,
    n40851, n40852, n40853, n40854, n40855, n40856,
    n40857, n40858, n40859, n40860, n40861, n40862,
    n40863, n40864, n40865, n40866, n40867, n40868,
    n40869, n40870, n40871, n40872, n40873, n40874,
    n40875, n40876, n40877, n40878, n40879, n40880,
    n40881, n40882, n40883, n40884, n40885, n40886,
    n40887, n40888, n40889, n40890, n40891, n40892,
    n40893, n40894, n40895, n40896, n40897, n40898,
    n40899, n40900, n40901, n40902, n40903, n40904,
    n40905, n40906, n40907, n40908, n40909, n40910,
    n40911, n40912, n40913, n40914, n40915, n40916,
    n40917, n40918, n40919, n40920, n40921, n40922,
    n40923, n40924, n40925, n40926, n40927, n40928,
    n40929, n40930, n40931, n40932, n40933, n40934,
    n40935, n40936, n40937, n40938, n40939, n40940,
    n40941, n40942, n40943, n40944, n40945, n40946,
    n40947, n40948, n40949, n40950, n40951, n40952,
    n40953, n40954, n40955, n40956, n40957, n40958,
    n40959, n40960, n40961, n40962, n40963, n40964,
    n40965, n40966, n40968, n40969, n40970, n40971,
    n40972, n40973, n40974, n40975, n40976, n40977,
    n40978, n40979, n40980, n40981, n40982, n40983,
    n40984, n40985, n40986, n40987, n40988, n40989,
    n40990, n40991, n40992, n40993, n40994, n40995,
    n40996, n40997, n40998, n40999, n41000, n41001,
    n41002, n41003, n41004, n41005, n41006, n41007,
    n41008, n41009, n41010, n41011, n41012, n41013,
    n41014, n41015, n41016, n41017, n41018, n41019,
    n41020, n41021, n41022, n41023, n41024, n41025,
    n41026, n41027, n41028, n41029, n41030, n41031,
    n41032, n41033, n41034, n41035, n41036, n41037,
    n41038, n41039, n41040, n41041, n41042, n41043,
    n41044, n41045, n41046, n41047, n41048, n41049,
    n41050, n41051, n41052, n41053, n41054, n41055,
    n41056, n41057, n41058, n41059, n41060, n41061,
    n41062, n41063, n41064, n41065, n41066, n41067,
    n41068, n41069, n41070, n41071, n41072, n41073,
    n41074, n41075, n41076, n41077, n41078, n41079,
    n41080, n41081, n41082, n41083, n41084, n41085,
    n41086, n41087, n41088, n41089, n41090, n41091,
    n41092, n41093, n41094, n41095, n41096, n41097,
    n41098, n41099, n41100, n41101, n41102, n41103,
    n41104, n41105, n41106, n41107, n41108, n41109,
    n41110, n41111, n41112, n41113, n41114, n41115,
    n41116, n41117, n41118, n41119, n41120, n41121,
    n41122, n41123, n41124, n41125, n41126, n41127,
    n41128, n41129, n41130, n41131, n41132, n41133,
    n41134, n41135, n41136, n41137, n41138, n41139,
    n41140, n41141, n41142, n41143, n41144, n41145,
    n41146, n41147, n41148, n41149, n41150, n41151,
    n41153, n41154, n41155, n41156, n41157, n41158,
    n41159, n41161, n41162, n41163, n41164, n41165,
    n41166, n41167, n41168, n41169, n41171, n41172,
    n41173, n41174, n41175, n41176, n41177, n41178,
    n41179, n41180, n41181, n41182, n41183, n41184,
    n41185, n41186, n41187, n41188, n41189, n41190,
    n41191, n41192, n41193, n41194, n41195, n41196,
    n41197, n41198, n41199, n41200, n41201, n41202,
    n41203, n41204, n41205, n41206, n41207, n41208,
    n41209, n41210, n41211, n41213, n41214, n41215,
    n41216, n41217, n41218, n41219, n41220, n41221,
    n41222, n41223, n41224, n41225, n41226, n41227,
    n41228, n41229, n41230, n41231, n41232, n41233,
    n41234, n41235, n41236, n41237, n41238, n41239,
    n41240, n41241, n41242, n41243, n41244, n41245,
    n41246, n41247, n41248, n41249, n41250, n41251,
    n41252, n41253, n41254, n41255, n41256, n41257,
    n41258, n41259, n41260, n41261, n41262, n41263,
    n41264, n41265, n41266, n41267, n41268, n41269,
    n41270, n41271, n41272, n41273, n41274, n41275,
    n41276, n41277, n41278, n41279, n41280, n41281,
    n41282, n41283, n41284, n41285, n41286, n41287,
    n41288, n41289, n41290, n41291, n41292, n41293,
    n41294, n41295, n41296, n41297, n41298, n41299,
    n41300, n41301, n41302, n41303, n41304, n41305,
    n41306, n41307, n41308, n41309, n41310, n41311,
    n41312, n41313, n41314, n41315, n41316, n41317,
    n41318, n41319, n41320, n41321, n41322, n41323,
    n41324, n41325, n41326, n41327, n41328, n41329,
    n41330, n41331, n41332, n41333, n41334, n41335,
    n41336, n41337, n41338, n41339, n41340, n41341,
    n41342, n41343, n41344, n41345, n41346, n41347,
    n41348, n41349, n41350, n41351, n41352, n41353,
    n41354, n41355, n41356, n41357, n41358, n41359,
    n41360, n41361, n41362, n41363, n41364, n41365,
    n41366, n41367, n41368, n41369, n41370, n41371,
    n41372, n41373, n41374, n41375, n41376, n41377,
    n41378, n41379, n41380, n41381, n41382, n41383,
    n41384, n41385, n41386, n41387, n41388, n41389,
    n41390, n41391, n41392, n41393, n41394, n41395,
    n41396, n41397, n41398, n41399, n41400, n41401,
    n41402, n41403, n41404, n41405, n41406, n41407,
    n41408, n41409, n41410, n41411, n41412, n41413,
    n41414, n41415, n41416, n41417, n41418, n41419,
    n41420, n41421, n41422, n41423, n41424, n41425,
    n41426, n41427, n41428, n41429, n41430, n41431,
    n41432, n41433, n41434, n41435, n41436, n41437,
    n41439, n41440, n41441, n41442, n41443, n41444,
    n41445, n41446, n41447, n41448, n41449, n41450,
    n41451, n41452, n41453, n41454, n41455, n41456,
    n41457, n41458, n41459, n41460, n41461, n41462,
    n41463, n41464, n41465, n41466, n41467, n41468,
    n41469, n41470, n41471, n41472, n41473, n41474,
    n41475, n41476, n41477, n41478, n41479, n41480,
    n41481, n41482, n41483, n41484, n41485, n41486,
    n41487, n41488, n41489, n41490, n41491, n41492,
    n41493, n41494, n41495, n41496, n41497, n41498,
    n41499, n41500, n41501, n41502, n41503, n41504,
    n41505, n41506, n41507, n41508, n41509, n41510,
    n41511, n41512, n41513, n41514, n41515, n41516,
    n41517, n41518, n41519, n41520, n41521, n41522,
    n41523, n41524, n41525, n41526, n41527, n41528,
    n41529, n41530, n41531, n41532, n41533, n41534,
    n41535, n41536, n41537, n41538, n41539, n41540,
    n41541, n41542, n41543, n41544, n41545, n41546,
    n41547, n41548, n41549, n41550, n41551, n41552,
    n41553, n41554, n41555, n41556, n41557, n41558,
    n41559, n41560, n41561, n41562, n41563, n41564,
    n41565, n41566, n41567, n41568, n41569, n41570,
    n41571, n41572, n41573, n41574, n41575, n41576,
    n41577, n41578, n41579, n41580, n41581, n41582,
    n41583, n41584, n41585, n41586, n41587, n41588,
    n41589, n41590, n41591, n41592, n41593, n41594,
    n41595, n41596, n41597, n41598, n41599, n41600,
    n41601, n41602, n41603, n41604, n41605, n41606,
    n41607, n41608, n41609, n41610, n41611, n41612,
    n41613, n41614, n41615, n41616, n41617, n41618,
    n41619, n41620, n41621, n41622, n41623, n41624,
    n41625, n41626, n41627, n41628, n41629, n41630,
    n41631, n41632, n41633, n41634, n41635, n41636,
    n41637, n41638, n41639, n41640, n41641, n41642,
    n41643, n41644, n41645, n41646, n41647, n41648,
    n41649, n41650, n41651, n41652, n41653, n41654,
    n41656, n41657, n41658, n41659, n41660, n41662,
    n41663, n41664, n41665, n41666, n41668, n41669,
    n41670, n41671, n41672, n41674, n41675, n41676,
    n41677, n41678, n41680, n41681, n41682, n41683,
    n41684, n41686, n41687, n41688, n41689, n41690,
    n41691, n41693, n41694, n41695, n41696, n41697,
    n41698, n41700, n41701, n41702, n41703, n41704,
    n41705, n41706, n41707, n41708, n41709, n41710,
    n41711, n41712, n41713, n41714, n41715, n41716,
    n41717, n41718, n41719, n41720, n41721, n41722,
    n41723, n41724, n41725, n41726, n41727, n41728,
    n41729, n41730, n41731, n41732, n41734, n41735,
    n41736, n41737, n41738, n41739, n41740, n41741,
    n41742, n41743, n41744, n41745, n41746, n41747,
    n41748, n41749, n41750, n41751, n41752, n41753,
    n41754, n41755, n41756, n41757, n41758, n41759,
    n41760, n41761, n41762, n41763, n41764, n41765,
    n41766, n41767, n41768, n41769, n41770, n41771,
    n41772, n41773, n41774, n41775, n41776, n41777,
    n41778, n41779, n41780, n41781, n41782, n41783,
    n41784, n41785, n41786, n41787, n41788, n41789,
    n41790, n41791, n41792, n41793, n41794, n41795,
    n41796, n41797, n41798, n41799, n41800, n41801,
    n41802, n41803, n41804, n41805, n41806, n41807,
    n41808, n41809, n41810, n41811, n41812, n41813,
    n41814, n41815, n41816, n41817, n41818, n41819,
    n41820, n41821, n41822, n41823, n41824, n41825,
    n41826, n41827, n41828, n41829, n41830, n41831,
    n41832, n41833, n41834, n41835, n41836, n41837,
    n41838, n41839, n41840, n41841, n41842, n41843,
    n41844, n41845, n41846, n41847, n41848, n41849,
    n41850, n41851, n41852, n41853, n41854, n41855,
    n41856, n41857, n41858, n41859, n41860, n41861,
    n41862, n41863, n41864, n41865, n41866, n41867,
    n41868, n41869, n41870, n41871, n41872, n41873,
    n41874, n41875, n41876, n41877, n41878, n41879,
    n41880, n41881, n41882, n41883, n41884, n41885,
    n41886, n41887, n41888, n41889, n41890, n41891,
    n41892, n41893, n41894, n41895, n41896, n41897,
    n41898, n41899, n41900, n41901, n41902, n41903,
    n41904, n41905, n41906, n41907, n41908, n41909,
    n41910, n41911, n41912, n41913, n41914, n41915,
    n41916, n41917, n41918, n41919, n41920, n41921,
    n41922, n41923, n41924, n41925, n41926, n41927,
    n41928, n41929, n41930, n41931, n41932, n41933,
    n41934, n41935, n41936, n41937, n41938, n41940,
    n41941, n41942, n41943, n41944, n41945, n41946,
    n41947, n41948, n41949, n41950, n41951, n41952,
    n41953, n41954, n41955, n41956, n41957, n41958,
    n41959, n41960, n41961, n41962, n41963, n41964,
    n41965, n41966, n41967, n41968, n41969, n41970,
    n41971, n41972, n41973, n41974, n41975, n41976,
    n41977, n41978, n41979, n41980, n41981, n41982,
    n41983, n41985, n41986, n41987, n41988, n41989,
    n41990, n41991, n41992, n41993, n41994, n41995,
    n41996, n41997, n41998, n41999, n42000, n42001,
    n42002, n42003, n42004, n42005, n42006, n42007,
    n42008, n42009, n42010, n42011, n42012, n42013,
    n42014, n42015, n42016, n42017, n42018, n42019,
    n42020, n42021, n42022, n42023, n42025, n42026,
    n42027, n42028, n42029, n42030, n42031, n42032,
    n42033, n42034, n42035, n42036, n42037, n42038,
    n42039, n42040, n42041, n42042, n42043, n42044,
    n42045, n42046, n42047, n42048, n42049, n42050,
    n42051, n42052, n42053, n42054, n42055, n42056,
    n42057, n42058, n42059, n42060, n42061, n42062,
    n42063, n42064, n42065, n42066, n42067, n42068,
    n42069, n42070, n42071, n42072, n42073, n42074,
    n42075, n42076, n42077, n42078, n42079, n42080,
    n42081, n42082, n42083, n42084, n42085, n42086,
    n42087, n42088, n42089, n42090, n42092, n42093,
    n42094, n42095, n42096, n42097, n42098, n42099,
    n42100, n42101, n42102, n42103, n42104, n42105,
    n42106, n42107, n42108, n42109, n42110, n42111,
    n42112, n42113, n42114, n42115, n42116, n42117,
    n42118, n42119, n42120, n42121, n42122, n42123,
    n42124, n42125, n42126, n42127, n42128, n42129,
    n42130, n42131, n42132, n42133, n42134, n42135,
    n42136, n42137, n42138, n42139, n42140, n42141,
    n42142, n42143, n42144, n42145, n42146, n42147,
    n42148, n42149, n42150, n42151, n42152, n42153,
    n42154, n42155, n42156, n42157, n42158, n42159,
    n42160, n42161, n42162, n42163, n42164, n42165,
    n42166, n42167, n42168, n42169, n42170, n42171,
    n42172, n42173, n42174, n42175, n42176, n42177,
    n42178, n42179, n42180, n42181, n42182, n42183,
    n42184, n42185, n42186, n42187, n42188, n42189,
    n42190, n42191, n42192, n42193, n42194, n42195,
    n42196, n42197, n42198, n42199, n42200, n42201,
    n42202, n42203, n42204, n42205, n42206, n42207,
    n42208, n42209, n42210, n42211, n42212, n42213,
    n42214, n42215, n42216, n42217, n42218, n42219,
    n42220, n42221, n42222, n42223, n42224, n42225,
    n42226, n42227, n42228, n42229, n42230, n42231,
    n42232, n42233, n42234, n42235, n42236, n42237,
    n42238, n42239, n42240, n42241, n42242, n42243,
    n42244, n42245, n42246, n42247, n42248, n42249,
    n42250, n42251, n42252, n42253, n42254, n42255,
    n42256, n42257, n42258, n42259, n42260, n42261,
    n42262, n42263, n42264, n42265, n42266, n42267,
    n42268, n42269, n42270, n42271, n42272, n42273,
    n42274, n42275, n42276, n42277, n42278, n42279,
    n42280, n42281, n42282, n42283, n42284, n42285,
    n42286, n42287, n42289, n42290, n42291, n42292,
    n42293, n42294, n42295, n42296, n42297, n42298,
    n42299, n42300, n42301, n42302, n42303, n42304,
    n42305, n42306, n42307, n42308, n42309, n42310,
    n42311, n42312, n42313, n42314, n42315, n42316,
    n42317, n42318, n42319, n42320, n42321, n42322,
    n42323, n42324, n42325, n42326, n42327, n42328,
    n42329, n42330, n42331, n42332, n42333, n42334,
    n42335, n42336, n42337, n42338, n42339, n42340,
    n42341, n42342, n42343, n42344, n42345, n42346,
    n42347, n42348, n42349, n42350, n42351, n42352,
    n42353, n42354, n42355, n42356, n42357, n42358,
    n42359, n42360, n42361, n42362, n42363, n42364,
    n42365, n42366, n42367, n42368, n42369, n42370,
    n42371, n42372, n42373, n42374, n42375, n42376,
    n42377, n42378, n42379, n42380, n42381, n42382,
    n42383, n42384, n42385, n42386, n42387, n42388,
    n42389, n42390, n42391, n42392, n42393, n42394,
    n42395, n42396, n42397, n42398, n42399, n42400,
    n42401, n42402, n42403, n42404, n42405, n42406,
    n42407, n42408, n42409, n42410, n42411, n42412,
    n42413, n42414, n42415, n42416, n42417, n42418,
    n42419, n42420, n42421, n42422, n42423, n42424,
    n42425, n42426, n42427, n42428, n42429, n42430,
    n42431, n42432, n42433, n42434, n42435, n42436,
    n42437, n42438, n42440, n42441, n42442, n42443,
    n42444, n42445, n42446, n42447, n42448, n42449,
    n42450, n42451, n42452, n42453, n42454, n42455,
    n42456, n42457, n42458, n42459, n42460, n42461,
    n42462, n42463, n42464, n42465, n42466, n42467,
    n42468, n42469, n42470, n42471, n42472, n42473,
    n42474, n42475, n42476, n42477, n42478, n42479,
    n42480, n42481, n42482, n42484, n42485, n42486,
    n42487, n42488, n42489, n42490, n42491, n42492,
    n42493, n42494, n42495, n42496, n42497, n42498,
    n42499, n42500, n42501, n42502, n42503, n42504,
    n42505, n42506, n42507, n42508, n42509, n42510,
    n42511, n42512, n42513, n42514, n42515, n42516,
    n42517, n42518, n42519, n42520, n42521, n42522,
    n42523, n42524, n42525, n42526, n42528, n42529,
    n42530, n42531, n42532, n42533, n42534, n42535,
    n42536, n42537, n42538, n42539, n42540, n42541,
    n42542, n42543, n42544, n42545, n42546, n42547,
    n42548, n42549, n42550, n42551, n42552, n42553,
    n42554, n42555, n42556, n42557, n42558, n42559,
    n42560, n42561, n42562, n42563, n42564, n42565,
    n42566, n42567, n42568, n42569, n42570, n42571,
    n42572, n42573, n42575, n42576, n42577, n42578,
    n42579, n42580, n42581, n42582, n42583, n42584,
    n42585, n42586, n42587, n42588, n42589, n42590,
    n42591, n42592, n42593, n42594, n42595, n42596,
    n42597, n42598, n42599, n42600, n42601, n42602,
    n42603, n42604, n42605, n42606, n42607, n42608,
    n42609, n42610, n42611, n42612, n42613, n42614,
    n42615, n42616, n42617, n42618, n42619, n42620,
    n42621, n42622, n42623, n42624, n42625, n42626,
    n42627, n42628, n42629, n42630, n42631, n42632,
    n42633, n42634, n42635, n42636, n42637, n42638,
    n42639, n42640, n42641, n42642, n42643, n42644,
    n42645, n42646, n42647, n42649, n42650, n42651,
    n42652, n42653, n42654, n42655, n42656, n42657,
    n42658, n42659, n42660, n42661, n42662, n42663,
    n42664, n42665, n42666, n42667, n42668, n42669,
    n42670, n42671, n42672, n42673, n42674, n42675,
    n42676, n42677, n42678, n42679, n42680, n42681,
    n42682, n42683, n42684, n42685, n42686, n42687,
    n42688, n42689, n42690, n42691, n42692, n42693,
    n42694, n42695, n42696, n42697, n42698, n42699,
    n42700, n42701, n42702, n42703, n42704, n42705,
    n42706, n42707, n42708, n42709, n42711, n42712,
    n42713, n42714, n42715, n42716, n42717, n42718,
    n42719, n42720, n42721, n42722, n42723, n42724,
    n42725, n42726, n42727, n42728, n42729, n42730,
    n42731, n42732, n42733, n42734, n42735, n42736,
    n42737, n42738, n42739, n42740, n42741, n42742,
    n42743, n42744, n42745, n42746, n42747, n42748,
    n42749, n42750, n42752, n42753, n42754, n42755,
    n42756, n42757, n42758, n42759, n42760, n42761,
    n42762, n42763, n42764, n42765, n42766, n42767,
    n42768, n42769, n42770, n42771, n42772, n42773,
    n42774, n42775, n42776, n42777, n42778, n42779,
    n42780, n42781, n42782, n42783, n42784, n42785,
    n42786, n42787, n42788, n42789, n42790, n42791,
    n42792, n42793, n42794, n42795, n42796, n42797,
    n42798, n42799, n42800, n42801, n42802, n42803,
    n42804, n42805, n42806, n42807, n42808, n42809,
    n42810, n42811, n42812, n42813, n42814, n42815,
    n42816, n42817, n42818, n42819, n42820, n42821,
    n42822, n42824, n42825, n42826, n42827, n42828,
    n42829, n42830, n42831, n42832, n42833, n42834,
    n42835, n42836, n42837, n42838, n42839, n42840,
    n42841, n42842, n42843, n42844, n42845, n42846,
    n42847, n42848, n42849, n42850, n42851, n42852,
    n42854, n42855, n42856, n42857, n42858, n42859,
    n42860, n42861, n42862, n42863, n42864, n42865,
    n42866, n42867, n42868, n42869, n42870, n42871,
    n42872, n42873, n42874, n42875, n42876, n42877,
    n42878, n42879, n42880, n42881, n42882, n42883,
    n42884, n42885, n42886, n42887, n42888, n42889,
    n42890, n42891, n42892, n42893, n42894, n42895,
    n42897, n42898, n42899, n42900, n42901, n42902,
    n42903, n42904, n42905, n42906, n42907, n42908,
    n42909, n42910, n42911, n42912, n42913, n42914,
    n42915, n42916, n42917, n42918, n42919, n42920,
    n42921, n42922, n42923, n42924, n42925, n42926,
    n42927, n42928, n42929, n42930, n42931, n42932,
    n42933, n42934, n42935, n42936, n42937, n42938,
    n42939, n42940, n42941, n42942, n42943, n42944,
    n42945, n42946, n42947, n42948, n42949, n42950,
    n42951, n42952, n42953, n42954, n42955, n42956,
    n42957, n42958, n42959, n42960, n42961, n42962,
    n42963, n42965, n42966, n42967, n42968, n42969,
    n42970, n42971, n42972, n42973, n42974, n42975,
    n42976, n42977, n42978, n42979, n42980, n42981,
    n42982, n42983, n42984, n42985, n42986, n42987,
    n42988, n42989, n42990, n42991, n42992, n42993,
    n42994, n42995, n42996, n42997, n42998, n42999,
    n43000, n43001, n43002, n43003, n43004, n43005,
    n43006, n43007, n43008, n43009, n43010, n43011,
    n43012, n43013, n43014, n43015, n43016, n43017,
    n43018, n43019, n43020, n43021, n43022, n43024,
    n43025, n43026, n43027, n43028, n43029, n43030,
    n43031, n43032, n43033, n43034, n43035, n43036,
    n43037, n43038, n43039, n43040, n43041, n43042,
    n43043, n43044, n43045, n43046, n43047, n43048,
    n43049, n43050, n43051, n43052, n43053, n43054,
    n43055, n43056, n43057, n43058, n43059, n43060,
    n43061, n43062, n43063, n43064, n43065, n43066,
    n43068, n43069, n43070, n43071, n43072, n43073,
    n43074, n43075, n43076, n43077, n43078, n43079,
    n43080, n43081, n43082, n43083, n43084, n43085,
    n43086, n43087, n43088, n43089, n43090, n43091,
    n43092, n43093, n43094, n43095, n43096, n43097,
    n43098, n43099, n43100, n43101, n43102, n43103,
    n43104, n43105, n43107, n43108, n43109, n43110,
    n43111, n43112, n43113, n43114, n43115, n43116,
    n43117, n43118, n43119, n43120, n43121, n43122,
    n43123, n43124, n43125, n43126, n43127, n43128,
    n43129, n43130, n43131, n43132, n43133, n43134,
    n43135, n43136, n43137, n43138, n43139, n43140,
    n43141, n43142, n43143, n43144, n43145, n43147,
    n43148, n43149, n43150, n43151, n43152, n43153,
    n43154, n43155, n43156, n43157, n43158, n43159,
    n43160, n43161, n43162, n43163, n43164, n43165,
    n43166, n43167, n43168, n43169, n43170, n43171,
    n43172, n43173, n43174, n43175, n43176, n43177,
    n43178, n43179, n43180, n43181, n43182, n43183,
    n43184, n43185, n43186, n43187, n43188, n43189,
    n43190, n43191, n43192, n43193, n43194, n43195,
    n43196, n43197, n43198, n43199, n43200, n43201,
    n43202, n43203, n43204, n43206, n43207, n43208,
    n43210, n43211, n43212, n43213, n43214, n43215,
    n43217, n43218, n43219, n43220, n43221, n43222,
    n43223, n43224, n43225, n43226, n43227, n43229,
    n43230, n43231, n43232, n43233, n43234, n43235,
    n43236, n43237, n43238, n43239, n43240, n43241,
    n43242, n43243, n43244, n43245, n43247, n43249,
    n43250, n43251, n43252, n43253, n43255, n43256,
    n43257, n43258, n43259, n43260, n43261, n43262,
    n43263, n43264, n43265, n43266, n43268, n43269,
    n43271, n43272, n43274, n43275, n43277, n43278,
    n43280, n43281, n43283, n43284, n43286, n43287,
    n43289, n43290, n43292, n43293, n43295, n43296,
    n43297, n43298, n43299, n43300, n43301, n43303,
    n43304, n43305, n43306, n43307, n43308, n43310,
    n43311, n43312, n43313, n43315, n43316, n43317,
    n43318, n43319, n43320, n43321, n43322, n43323,
    n43324, n43325, n43326, n43327, n43328, n43329,
    n43330, n43331, n43332, n43333, n43334, n43335,
    n43336, n43338, n43339, n43341, n43342, n43344,
    n43345, n43347, n43348, n43350, n43351, n43353,
    n43354, n43356, n43357, n43359, n43360, n43361,
    n43362, n43363, n43364, n43365, n43366, n43367,
    n43368, n43369, n43370, n43371, n43372, n43373,
    n43374, n43375, n43376, n43377, n43378, n43379,
    n43380, n43381, n43382, n43384, n43385, n43386,
    n43388, n43389, n43391, n43392, n43393, n43395,
    n43396, n43398, n43399, n43400, n43401, n43402,
    n43403, n43404, n43405, n43406, n43407, n43408,
    n43410, n43411, n43412, n43414, n43415, n43417,
    n43418, n43419, n43421, n43422, n43423, n43425,
    n43426, n43428, n43429, n43431, n43432, n43434,
    n43435, n43437, n43438, n43440, n43441, n43443,
    n43444, n43446, n43447, n43449, n43450, n43452,
    n43453, n43455, n43456, n43458, n43459, n43460,
    n43461, n43462, n43463, n43464, n43465, n43467,
    n43468, n43469, n43470, n43471, n43473, n43474,
    n43475, n43476, n43477, n43478, n43479, n43480,
    n43481, n43482, n43483, n43485, n43486, n43488,
    n43489, n43491, n43492, n43494, n43495, n43497,
    n43498, n43500, n43501, n43503, n43504, n43506,
    n43507, n43508, n43509, n43510, n43512, n43513,
    n43515, n43516, n43518, n43519, n43521, n43522,
    n43524, n43525, n43527, n43528, n43530, n43531,
    n43533, n43534, n43536, n43537, n43539, n43540,
    n43542, n43543, n43545, n43546, n43548, n43549,
    n43551, n43552, n43554, n43555, n43557, n43558,
    n43560, n43561, n43563, n43564, n43566, n43567,
    n43569, n43570, n43572, n43573, n43575, n43576,
    n43578, n43579, n43581, n43582, n43584, n43585,
    n43587, n43588, n43590, n43591, n43593, n43594,
    n43596, n43597, n43599, n43600, n43602, n43603,
    n43605, n43606, n43608, n43609, n43611, n43612,
    n43614, n43615, n43617, n43618, n43620, n43621,
    n43623, n43624, n43626, n43627, n43629, n43630,
    n43632, n43633, n43635, n43636, n43638, n43639,
    n43641, n43642, n43644, n43645, n43647, n43648,
    n43650, n43651, n43653, n43654, n43656, n43657,
    n43659, n43660, n43662, n43663, n43665, n43666,
    n43668, n43669, n43671, n43672, n43674, n43675,
    n43677, n43678, n43680, n43681, n43683, n43684,
    n43686, n43687, n43689, n43690, n43692, n43693,
    n43695, n43696, n43698, n43699, n43701, n43702,
    n43704, n43705, n43707, n43708, n43710, n43711,
    n43713, n43714, n43716, n43717, n43719, n43720,
    n43722, n43723, n43725, n43726, n43728, n43729,
    n43731, n43732, n43733, n43735, n43736, n43738,
    n43739, n43741, n43742, n43744, n43745, n43747,
    n43748, n43750, n43751, n43753, n43754, n43756,
    n43757, n43759, n43760, n43762, n43763, n43765,
    n43766, n43768, n43769, n43771, n43772, n43774,
    n43775, n43777, n43778, n43780, n43781, n43783,
    n43784, n43786, n43787, n43789, n43790, n43792,
    n43793, n43795, n43796, n43798, n43799, n43801,
    n43802, n43804, n43805, n43807, n43808, n43810,
    n43811, n43813, n43814, n43816, n43817, n43819,
    n43820, n43822, n43823, n43825, n43826, n43828,
    n43829, n43831, n43832, n43834, n43835, n43837,
    n43838, n43840, n43841, n43843, n43844, n43846,
    n43847, n43849, n43850, n43852, n43853, n43855,
    n43856, n43858, n43859, n43861, n43862, n43863,
    n43864, n43865, n43866, n43867, n43868, n43869,
    n43870, n43871, n43872, n43873, n43874, n43875,
    n43876, n43877, n43878, n43879, n43880, n43881,
    n43882, n43883, n43885, n43886, n43888, n43889,
    n43891, n43892, n43894, n43895, n43897, n43898,
    n43900, n43901, n43903, n43904, n43906, n43907,
    n43908, n43909, n43910, n43911, n43912, n43913,
    n43914, n43915, n43916, n43917, n43918, n43919,
    n43920, n43921, n43922, n43923, n43924, n43925,
    n43926, n43927, n43928, n43929, n43930, n43932,
    n43933, n43934, n43935, n43936, n43937, n43938,
    n43939, n43940, n43941, n43942, n43943, n43944,
    n43945, n43946, n43947, n43949, n43950, n43951,
    n43952, n43953, n43954, n43955, n43956, n43957,
    n43958, n43959, n43960, n43961, n43962, n43963,
    n43964, n43965, n43966, n43967, n43968, n43969,
    n43970, n43971, n43972, n43973, n43974, n43975,
    n43976, n43978, n43979, n43980, n43981, n43983,
    n43984, n43985, n43986, n43987, n43988, n43989,
    n43990, n43991, n43992, n43993, n43994, n43995,
    n43996, n43997, n43998, n43999, n44000, n44001,
    n44003, n44004, n44005, n44006, n44007, n44008,
    n44009, n44010, n44011, n44012, n44013, n44014,
    n44015, n44016, n44017, n44018, n44019, n44020,
    n44021, n44023, n44024, n44025, n44026, n44027,
    n44028, n44029, n44030, n44031, n44032, n44033,
    n44034, n44035, n44036, n44037, n44038, n44039,
    n44040, n44041, n44043, n44044, n44045, n44046,
    n44047, n44048, n44049, n44050, n44051, n44052,
    n44053, n44054, n44055, n44056, n44057, n44058,
    n44059, n44060, n44061, n44063, n44064, n44065,
    n44066, n44067, n44068, n44069, n44070, n44071,
    n44072, n44074, n44075, n44076, n44077, n44078,
    n44079, n44080, n44081, n44082, n44083, n44085,
    n44086, n44087, n44088, n44089, n44090, n44091,
    n44092, n44093, n44094, n44096, n44097, n44098,
    n44099, n44100, n44101, n44102, n44103, n44104,
    n44105, n44106, n44109, n44110, n44112, n44113,
    n44115, n44116, n44118, n44119, n44121, n44122,
    n44124, n44125, n44127, n44128, n44130, n44131,
    n44133, n44134, n44136, n44137, n44139, n44140,
    n44142, n44143, n44145, n44146, n44148, n44149,
    n44151, n44152, n44154, n44155, n44157, n44158,
    n44160, n44161, n44163, n44164, n44166, n44167,
    n44169, n44170, n44172, n44173, n44175, n44176,
    n44178, n44179, n44181, n44182, n44184, n44185,
    n44187, n44188, n44190, n44191, n44193, n44194,
    n44196, n44197, n44199, n44200, n44202, n44203,
    n44205, n44206, n44208, n44209, n44211, n44212,
    n44214, n44215, n44217, n44218, n44220, n44221,
    n44223, n44224, n44226, n44227, n44229, n44230,
    n44232, n44233, n44235, n44236, n44238, n44239,
    n44241, n44242, n44244, n44245, n44247, n44248,
    n44250, n44251, n44253, n44254, n44256, n44257,
    n44259, n44260, n44262, n44263, n44265, n44266,
    n44268, n44269, n44271, n44272, n44274, n44275,
    n44277, n44278, n44280, n44281, n44283, n44284,
    n44286, n44287, n44289, n44290, n44292, n44293,
    n44295, n44296, n44298, n44299, n44301, n44302,
    n44304, n44305, n44307, n44308, n44310, n44311,
    n44313, n44314, n44316, n44317, n44319, n44320,
    n44322, n44323, n44325, n44326, n44328, n44329,
    n44331, n44332, n44334, n44335, n44337, n44338,
    n44340, n44341, n44343, n44344, n44346, n44347,
    n44349, n44350, n44352, n44353, n44355, n44356,
    n44358, n44359, n44361, n44362, n44364, n44365,
    n44367, n44368, n44369, n44370, n44371, n44372,
    n44373, n44374, n44375, n44376, n44377, n44378,
    n44379, n44380, n44381, n44382, n44383, n44384,
    n44385, n44386, n44387, n44388, n44389, n44390,
    n44391, n44392, n44393, n44394, n44395, n44396,
    n44397, n44398, n44399, n44400, n44401, n44402,
    n44403, n44404, n44405, n44406, n44407, n44408,
    n44409, n44410, n44411, n44412, n44413, n44414,
    n44415, n44416, n44417, n44418, n44419, n44420,
    n44421, n44422, n44423, n44424, n44425, n44426,
    n44427, n44428, n44429, n44430, n44431, n44432,
    n44433, n44434, n44435, n44436, n44437, n44438,
    n44439, n44440, n44441, n44442, n44443, n44444,
    n44445, n44446, n44447, n44448, n44449, n44450,
    n44451, n44452, n44453, n44454, n44455, n44456,
    n44457, n44458, n44459, n44460, n44461, n44462,
    n44463, n44464, n44465, n44466, n44467, n44468,
    n44469, n44470, n44471, n44473, n44474, n44476,
    n44477, n44479, n44480, n44482, n44483, n44485,
    n44486, n44488, n44489, n44491, n44492, n44494,
    n44495, n44497, n44498, n44500, n44501, n44503,
    n44504, n44506, n44507, n44509, n44510, n44512,
    n44513, n44515, n44516, n44518, n44519, n44521,
    n44522, n44524, n44525, n44527, n44528, n44529,
    n44530, n44531, n44532, n44533, n44535, n44536,
    n44537, n44538, n44540, n44541, n44542, n44543,
    n44544, n44545, n44546, n44547, n44548, n44549,
    n44550, n44551, n44552, n44553, n44554, n44555,
    n44556, n44557, n44558, n44559, n44561, n44562,
    n44563, n44565, n44566, n44567, n44569, n44570,
    n44571, n44573, n44574, n44575, n44576, n44577,
    n44578, n44579, n44580, n44581, n44582, n44583,
    n44584, n44585, n44586, n44587, n44588, n44589,
    n44590, n44591, n44592, n44593, n44594, n44595,
    n44596, n44597, n44598, n44599, n44600, n44601,
    n44602, n44603, n44604, n44605, n44606, n44607,
    n44608, n44609, n44610, n44611, n44612, n44613,
    n44614, n44615, n44616, n44617, n44618, n44619,
    n44620, n44621, n44622, n44623, n44624, n44625,
    n44626, n44627, n44628, n44629, n44630, n44631,
    n44632, n44633, n44634, n44635, n44636, n44637,
    n44638, n44639, n44640, n44641, n44642, n44643,
    n44644, n44645, n44646, n44647, n44648, n44649,
    n44650, n44651, n44652, n44653, n44654, n44655,
    n44656, n44657, n44658, n44659, n44660, n44661,
    n44662, n44663, n44664, n44665, n44666, n44667,
    n44668, n44669, n44670, n44671, n44672, n44673,
    n44674, n44675, n44676, n44677, n44678, n44679,
    n44680, n44681, n44682, n44683, n44684, n44685,
    n44686, n44687, n44688, n44689, n44690, n44691,
    n44692, n44693, n44694, n44695, n44696, n44697,
    n44698, n44699, n44700, n44701, n44702, n44703,
    n44704, n44705, n44706, n44707, n44708, n44709,
    n44710, n44711, n44712, n44713, n44714, n44715,
    n44716, n44717, n44718, n44719, n44720, n44721,
    n44722, n44723, n44724, n44725, n44726, n44727,
    n44728, n44729, n44730, n44731, n44732, n44733,
    n44734, n44735, n44736, n44737, n44738, n44739,
    n44740, n44741, n44742, n44743, n44744, n44745,
    n44746, n44747, n44748, n44749, n44750, n44751,
    n44752, n44753, n44754, n44755, n44756, n44757,
    n44758, n44759, n44760, n44761, n44762, n44763,
    n44764, n44765, n44766, n44767, n44768, n44769,
    n44770, n44771, n44772, n44773, n44774, n44775,
    n44776, n44777, n44778, n44779, n44780, n44781,
    n44782, n44783, n44784, n44785, n44786, n44787,
    n44788, n44789, n44790, n44791, n44792, n44793,
    n44794, n44795, n44796, n44797, n44798, n44799,
    n44800, n44801, n44802, n44803, n44804, n44805,
    n44806, n44807, n44808, n44809, n44810, n44811,
    n44812, n44813, n44814, n44815, n44816, n44817,
    n44818, n44819, n44820, n44821, n44822, n44823,
    n44824, n44825, n44826, n44827, n44828, n44829,
    n44830, n44831, n44832, n44833, n44834, n44835,
    n44836, n44837, n44838, n44839, n44840, n44841,
    n44842, n44843, n44844, n44845, n44846, n44847,
    n44848, n44849, n44850, n44851, n44852, n44853,
    n44854, n44855, n44856, n44857, n44858, n44859,
    n44860, n44861, n44862, n44863, n44864, n44865,
    n44866, n44867, n44868, n44869, n44870, n44871,
    n44872, n44873, n44874, n44875, n44876, n44877,
    n44878, n44879, n44880, n44881, n44882, n44883,
    n44884, n44885, n44886, n44887, n44888, n44889,
    n44890, n44891, n44892, n44893, n44894, n44895,
    n44896, n44897, n44898, n44899, n44900, n44901,
    n44902, n44903, n44904, n44905, n44906, n44907,
    n44908, n44909, n44910, n44911, n44912, n44913,
    n44914, n44915, n44916, n44917, n44918, n44919,
    n44920, n44921, n44922, n44923, n44924, n44925,
    n44926, n44927, n44928, n44929, n44930, n44931,
    n44932, n44933, n44934, n44935, n44936, n44937,
    n44938, n44939, n44940, n44941, n44942, n44943,
    n44944, n44945, n44946, n44947, n44948, n44949,
    n44950, n44951, n44952, n44953, n44954, n44955,
    n44956, n44957, n44958, n44959, n44960, n44961,
    n44962, n44963, n44964, n44965, n44966, n44967,
    n44968, n44969, n44970, n44971, n44972, n44973,
    n44974, n44975, n44976, n44977, n44978, n44979,
    n44980, n44981, n44982, n44983, n44984, n44985,
    n44986, n44987, n44988, n44989, n44990, n44991,
    n44992, n44993, n44994, n44995, n44996, n44997,
    n44998, n44999, n45000, n45001, n45002, n45003,
    n45004, n45005, n45006, n45007, n45008, n45009,
    n45010, n45011, n45012, n45013, n45014, n45015,
    n45016, n45017, n45018, n45019, n45020, n45021,
    n45022, n45023, n45024, n45026, n45027, n45028,
    n45029, n45030, n45031, n45033, n45034, n45035,
    n45036, n45037, n45039, n45040, n45041, n45042,
    n45043, n45045, n45046, n45047, n45049, n45050,
    n45051, n45052, n45053, n45055, n45056, n45057,
    n45059, n45060, n45062, n45063, n45064, n45066,
    n45067, n45068, n45069, n45070, n45071, n45072,
    n45073, n45074, n45075, n45076, n45078, n45079,
    n45080, n45081, n45083, n45084, n45085, n45086,
    n45087, n45088, n45089, n45091, n45092, n45093,
    n45094, n45095, n45096, n45098, n45099, n45101,
    n45102, n45103, n45104, n45105, n45107, n45108,
    n45109, n45111, n45112, n45113, n45115, n45116,
    n45117, n45119, n45120, n45121, n45123, n45124,
    n45125, n45127, n45128, n45129, n45131, n45132,
    n45133, n45135, n45136, n45137, n45138, n45140,
    n45141, n45142, n45143, n45145, n45146, n45147,
    n45148, n45150, n45151, n45152, n45153, n45154,
    n45156, n45157, n45158, n45160, n45161, n45162,
    n45164, n45165, n45166, n45168, n45169, n45170,
    n45172, n45173, n45174, n45176, n45177, n45178,
    n45180, n45181, n45182, n45183, n45184, n45186,
    n45187, n45188, n45189, n45191, n45192, n45193,
    n45195, n45196, n45197, n45199, n45200, n45201,
    n45203, n45204, n45205, n45207, n45208, n45209,
    n45211, n45212, n45213, n45215, n45216, n45217,
    n45219, n45220, n45221, n45223, n45224, n45225,
    n45227, n45228, n45229, n45231, n45232, n45233,
    n45235, n45236, n45237, n45239, n45240, n45241,
    n45243, n45244, n45245, n45247, n45248, n45249,
    n45251, n45252, n45253, n45255, n45256, n45257,
    n45259, n45260, n45261, n45263, n45264, n45265,
    n45267, n45268, n45269, n45271, n45272, n45273,
    n45275, n45276, n45277, n45279, n45280, n45281,
    n45283, n45284, n45285, n45287, n45288, n45289,
    n45291, n45292, n45293, n45295, n45296, n45297,
    n45299, n45300, n45301, n45303, n45304, n45305,
    n45307, n45308, n45309, n45311, n45312, n45313,
    n45315, n45316, n45317, n45319, n45320, n45321,
    n45323, n45324, n45325, n45327, n45328, n45329,
    n45330, n45331, n45332, n45333, n45334, n45335,
    n45337, n45339, n45340, n45341, n45343, n45344,
    n45345, n45347, n45348, n45349, n45351, n45352,
    n45353, n45354, n45355, n45356, n45357, n45358,
    n45359, n45360, n45361, n45362, n45363, n45364,
    n45365, n45366, n45367, n45368, n45369, n45370,
    n45371, n45372, n45373, n45374, n45375, n45376,
    n45377, n45378, n45379, n45380, n45381, n45382,
    n45383, n45384, n45385, n45386, n45387, n45388,
    n45389, n45390, n45391, n45392, n45393, n45394,
    n45395, n45396, n45397, n45398, n45400, n45401,
    n45402, n45403, n45404, n45405, n45406, n45407,
    n45408, n45409, n45410, n45411, n45412, n45413,
    n45414, n45415, n45416, n45417, n45418, n45419,
    n45420, n45421, n45422, n45423, n45424, n45425,
    n45426, n45427, n45428, n45429, n45430, n45431,
    n45432, n45433, n45434, n45435, n45436, n45437,
    n45438, n45439, n45440, n45442, n45443, n45444,
    n45446, n45447, n45448, n45449, n45450, n45451,
    n45452, n45453, n45454, n45455, n45456, n45457,
    n45458, n45459, n45460, n45461, n45462, n45463,
    n45464, n45465, n45466, n45467, n45468, n45469,
    n45470, n45471, n45472, n45473, n45474, n45475,
    n45476, n45477, n45478, n45479, n45480, n45482,
    n45483, n45484, n45485, n45486, n45487, n45488,
    n45489, n45490, n45491, n45492, n45493, n45494,
    n45495, n45496, n45497, n45498, n45499, n45500,
    n45501, n45502, n45503, n45504, n45505, n45506,
    n45507, n45508, n45509, n45510, n45511, n45512,
    n45513, n45514, n45515, n45516, n45517, n45519,
    n45520, n45521, n45522, n45523, n45524, n45525,
    n45526, n45527, n45528, n45529, n45530, n45531,
    n45532, n45533, n45534, n45535, n45536, n45537,
    n45538, n45539, n45540, n45541, n45542, n45543,
    n45544, n45545, n45546, n45547, n45548, n45549,
    n45550, n45551, n45552, n45553, n45555, n45556,
    n45557, n45559, n45560, n45561, n45562, n45563,
    n45564, n45565, n45566, n45567, n45568, n45569,
    n45570, n45571, n45572, n45573, n45574, n45575,
    n45576, n45577, n45578, n45579, n45580, n45581,
    n45582, n45583, n45584, n45585, n45586, n45587,
    n45588, n45589, n45591, n45592, n45593, n45594,
    n45595, n45596, n45597, n45598, n45599, n45600,
    n45601, n45602, n45603, n45604, n45605, n45606,
    n45607, n45608, n45609, n45610, n45611, n45612,
    n45613, n45614, n45615, n45616, n45617, n45618,
    n45619, n45620, n45622, n45623, n45624, n45625,
    n45626, n45627, n45628, n45629, n45630, n45631,
    n45632, n45633, n45634, n45635, n45636, n45637,
    n45638, n45639, n45640, n45641, n45642, n45643,
    n45644, n45645, n45646, n45647, n45648, n45649,
    n45650, n45651, n45652, n45653, n45654, n45655,
    n45656, n45658, n45659, n45660, n45661, n45662,
    n45663, n45664, n45665, n45666, n45667, n45668,
    n45669, n45670, n45671, n45672, n45673, n45674,
    n45675, n45676, n45677, n45678, n45679, n45680,
    n45681, n45682, n45683, n45684, n45685, n45686,
    n45687, n45688, n45689, n45690, n45691, n45692,
    n45694, n45695, n45696, n45697, n45698, n45699,
    n45700, n45701, n45702, n45703, n45704, n45705,
    n45706, n45707, n45708, n45709, n45710, n45711,
    n45712, n45713, n45714, n45715, n45716, n45717,
    n45718, n45719, n45720, n45721, n45722, n45723,
    n45724, n45725, n45726, n45727, n45728, n45729,
    n45731, n45732, n45733, n45734, n45735, n45736,
    n45737, n45738, n45739, n45740, n45741, n45742,
    n45743, n45744, n45745, n45746, n45747, n45748,
    n45749, n45750, n45751, n45752, n45753, n45754,
    n45755, n45756, n45757, n45758, n45759, n45760,
    n45761, n45762, n45763, n45764, n45765, n45767,
    n45768, n45769, n45770, n45771, n45772, n45773,
    n45774, n45775, n45776, n45777, n45778, n45779,
    n45780, n45781, n45782, n45783, n45784, n45785,
    n45786, n45787, n45788, n45789, n45790, n45791,
    n45792, n45793, n45794, n45795, n45796, n45797,
    n45798, n45799, n45800, n45801, n45803, n45804,
    n45805, n45806, n45807, n45808, n45809, n45810,
    n45811, n45812, n45813, n45814, n45815, n45816,
    n45817, n45818, n45819, n45820, n45821, n45822,
    n45823, n45824, n45825, n45826, n45827, n45828,
    n45829, n45830, n45831, n45832, n45834, n45835,
    n45836, n45837, n45838, n45839, n45840, n45841,
    n45842, n45843, n45844, n45845, n45846, n45847,
    n45848, n45849, n45850, n45851, n45852, n45853,
    n45854, n45855, n45856, n45857, n45858, n45859,
    n45860, n45861, n45862, n45863, n45865, n45866,
    n45867, n45868, n45869, n45870, n45871, n45872,
    n45873, n45874, n45875, n45876, n45877, n45878,
    n45879, n45880, n45881, n45882, n45883, n45884,
    n45885, n45886, n45887, n45888, n45889, n45890,
    n45891, n45892, n45893, n45894, n45895, n45896,
    n45897, n45898, n45899, n45901, n45902, n45903,
    n45905, n45906, n45907, n45909, n45910, n45911,
    n45912, n45913, n45914, n45915, n45916, n45917,
    n45918, n45919, n45920, n45921, n45922, n45923,
    n45924, n45925, n45926, n45927, n45928, n45929,
    n45930, n45931, n45932, n45933, n45934, n45935,
    n45936, n45937, n45938, n45941, n45942, n45943,
    n45945, n45946, n45947, n45948, n45949, n45950,
    n45951, n45952, n45953, n45954, n45955, n45956,
    n45957, n45958, n45959, n45960, n45961, n45962,
    n45963, n45964, n45965, n45966, n45967, n45968,
    n45969, n45970, n45971, n45972, n45973, n45974,
    n45975, n45976, n45977, n45978, n45979, n45980,
    n45981, n45982, n45984, n45985, n45986, n45988,
    n45989, n45990, n45992, n45993, n45994, n45996,
    n45997, n45998, n45999, n46000, n46001, n46002,
    n46003, n46004, n46005, n46006, n46007, n46008,
    n46009, n46010, n46011, n46012, n46013, n46014,
    n46015, n46016, n46017, n46018, n46019, n46020,
    n46021, n46022, n46023, n46024, n46025, n46026,
    n46027, n46029, n46030, n46031, n46033, n46034,
    n46035, n46037, n46038, n46039, n46040, n46041,
    n46042, n46043, n46044, n46045, n46046, n46047,
    n46048, n46049, n46050, n46051, n46052, n46053,
    n46054, n46055, n46056, n46057, n46058, n46059,
    n46060, n46061, n46062, n46063, n46064, n46065,
    n46066, n46067, n46068, n46069, n46071, n46072,
    n46073, n46075, n46076, n46077, n46079, n46080,
    n46081, n46083, n46084, n46085, n46087, n46088,
    n46089, n46091, n46092, n46093, n46095, n46096,
    n46097, n46099, n46100, n46101, n46103, n46104,
    n46105, n46107, n46108, n46109, n46111, n46112,
    n46113, n46115, n46116, n46117, n46119, n46120,
    n46121, n46123, n46124, n46125, n46127, n46128,
    n46129, n46130, n46131, n46132, n46133, n46134,
    n46135, n46136, n46137, n46138, n46139, n46140,
    n46141, n46142, n46143, n46144, n46145, n46146,
    n46147, n46148, n46149, n46150, n46151, n46152,
    n46153, n46154, n46155, n46156, n46157, n46158,
    n46159, n46160, n46162, n46163, n46164, n46165,
    n46166, n46167, n46168, n46169, n46170, n46171,
    n46172, n46173, n46174, n46175, n46176, n46177,
    n46178, n46179, n46180, n46181, n46182, n46183,
    n46184, n46185, n46186, n46187, n46188, n46189,
    n46190, n46191, n46192, n46193, n46194, n46195,
    n46196, n46197, n46199, n46200, n46201, n46203,
    n46204, n46205, n46207, n46208, n46209, n46210,
    n46211, n46212, n46213, n46214, n46215, n46216,
    n46217, n46218, n46219, n46220, n46221, n46222,
    n46223, n46224, n46225, n46226, n46227, n46228,
    n46229, n46230, n46231, n46232, n46233, n46234,
    n46235, n46236, n46237, n46238, n46240, n46241,
    n46242, n46243, n46244, n46245, n46246, n46247,
    n46248, n46249, n46250, n46251, n46252, n46253,
    n46254, n46255, n46256, n46257, n46258, n46259,
    n46260, n46261, n46262, n46263, n46264, n46265,
    n46266, n46267, n46268, n46269, n46270, n46271,
    n46273, n46274, n46275, n46276, n46277, n46278,
    n46279, n46280, n46281, n46282, n46283, n46284,
    n46285, n46286, n46287, n46288, n46289, n46290,
    n46291, n46292, n46293, n46294, n46295, n46296,
    n46297, n46298, n46299, n46300, n46301, n46302,
    n46303, n46304, n46306, n46307, n46308, n46309,
    n46310, n46311, n46312, n46313, n46314, n46315,
    n46316, n46317, n46318, n46319, n46320, n46321,
    n46322, n46323, n46324, n46325, n46326, n46327,
    n46328, n46329, n46330, n46331, n46332, n46333,
    n46334, n46335, n46336, n46337, n46338, n46340,
    n46341, n46342, n46344, n46345, n46346, n46347,
    n46348, n46349, n46350, n46351, n46352, n46353,
    n46354, n46355, n46356, n46357, n46358, n46359,
    n46360, n46361, n46362, n46363, n46364, n46365,
    n46366, n46367, n46368, n46369, n46370, n46371,
    n46372, n46373, n46374, n46375, n46376, n46377,
    n46379, n46380, n46381, n46382, n46383, n46384,
    n46385, n46386, n46387, n46388, n46389, n46390,
    n46391, n46392, n46393, n46394, n46395, n46396,
    n46397, n46398, n46399, n46400, n46401, n46402,
    n46403, n46404, n46405, n46406, n46407, n46408,
    n46409, n46411, n46412, n46413, n46414, n46415,
    n46416, n46417, n46418, n46419, n46420, n46421,
    n46422, n46423, n46424, n46425, n46426, n46427,
    n46428, n46429, n46430, n46431, n46432, n46433,
    n46434, n46435, n46436, n46437, n46438, n46439,
    n46440, n46441, n46442, n46443, n46444, n46446,
    n46447, n46448, n46449, n46450, n46451, n46452,
    n46453, n46454, n46455, n46456, n46457, n46458,
    n46459, n46460, n46461, n46462, n46463, n46464,
    n46465, n46466, n46467, n46468, n46469, n46470,
    n46471, n46472, n46473, n46474, n46475, n46476,
    n46478, n46479, n46480, n46481, n46482, n46483,
    n46484, n46485, n46486, n46487, n46488, n46489,
    n46490, n46491, n46492, n46493, n46494, n46495,
    n46496, n46497, n46498, n46499, n46500, n46501,
    n46502, n46503, n46504, n46505, n46506, n46507,
    n46508, n46509, n46510, n46512, n46513, n46514,
    n46515, n46516, n46517, n46518, n46519, n46520,
    n46521, n46522, n46523, n46524, n46525, n46526,
    n46527, n46528, n46529, n46530, n46531, n46532,
    n46533, n46534, n46535, n46536, n46537, n46538,
    n46539, n46540, n46541, n46542, n46543, n46544,
    n46545, n46546, n46547, n46548, n46549, n46550,
    n46551, n46552, n46553, n46554, n46555, n46556,
    n46557, n46558, n46559, n46560, n46561, n46562,
    n46563, n46564, n46565, n46567, n46568, n46569,
    n46571, n46572, n46573, n46574, n46575, n46576,
    n46577, n46578, n46579, n46580, n46581, n46582,
    n46583, n46584, n46585, n46586, n46587, n46588,
    n46589, n46590, n46591, n46592, n46593, n46594,
    n46595, n46596, n46597, n46598, n46599, n46600,
    n46601, n46602, n46603, n46605, n46606, n46607,
    n46609, n46610, n46611, n46613, n46614, n46615,
    n46617, n46618, n46619, n46621, n46622, n46623,
    n46625, n46626, n46627, n46629, n46630, n46631,
    n46633, n46634, n46635, n46637, n46638, n46639,
    n46640, n46641, n46642, n46643, n46644, n46645,
    n46646, n46647, n46648, n46649, n46650, n46652,
    n46653, n46654, n46656, n46657, n46658, n46659,
    n46660, n46661, n46662, n46663, n46664, n46665,
    n46666, n46667, n46668, n46669, n46670, n46671,
    n46672, n46673, n46674, n46675, n46676, n46677,
    n46678, n46679, n46680, n46681, n46682, n46683,
    n46684, n46685, n46686, n46687, n46688, n46689,
    n46691, n46692, n46693, n46695, n46696, n46697,
    n46699, n46700, n46701, n46703, n46704, n46705,
    n46707, n46708, n46709, n46711, n46713, n46714,
    n46715, n46717, n46718, n46719, n46721, n46722,
    n46723, n46725, n46726, n46727, n46729, n46730,
    n46731, n46733, n46734, n46735, n46737, n46738,
    n46739, n46741, n46742, n46743, n46744, n46745,
    n46746, n46747, n46748, n46749, n46750, n46751,
    n46753, n46754, n46755, n46757, n46758, n46759,
    n46761, n46762, n46763, n46765, n46766, n46767,
    n46769, n46770, n46771, n46773, n46774, n46775,
    n46777, n46778, n46779, n46781, n46782, n46783,
    n46785, n46786, n46787, n46789, n46790, n46791,
    n46793, n46794, n46795, n46797, n46798, n46799,
    n46801, n46802, n46803, n46805, n46806, n46807,
    n46809, n46810, n46811, n46813, n46814, n46815,
    n46817, n46818, n46819, n46821, n46822, n46823,
    n46824, n46825, n46826, n46827, n46828, n46829,
    n46830, n46831, n46833, n46834, n46835, n46836,
    n46838, n46839, n46840, n46842, n46843, n46844,
    n46846, n46847, n46848, n46850, n46851, n46852,
    n46853, n46854, n46855, n46856, n46857, n46858,
    n46859, n46860, n46861, n46862, n46863, n46864,
    n46866, n46867, n46868, n46870, n46871, n46872,
    n46873, n46875, n46876, n46877, n46879, n46880,
    n46881, n46882, n46883, n46885, n46886, n46887,
    n46889, n46890, n46891, n46892, n46893, n46894,
    n46895, n46896, n46897, n46898, n46899, n46900,
    n46901, n46902, n46903, n46905, n46906, n46907,
    n46909, n46910, n46911, n46913, n46914, n46915,
    n46916, n46917, n46918, n46919, n46923, n46924,
    n46926, n46928, n46929, n46931, n46932, n46934,
    n46935, n46937, n46938, n46940, n46941, n46943,
    n46944, n46946, n46947, n46949, n46950, n46952,
    n46953, n46955, n46956, n46958, n46959, n46960,
    n46962, n46963, n46965, n46966, n46967, n46968,
    n46969, n46970, n46971, n46972, n46973, n46974,
    n46976, n46977, n46979, n46980, n46982, n46983,
    n46985, n46986, n46988, n46989, n46991, n46992,
    n46994, n46996, n46997, n46999, n47000, n47002,
    n47003, n47005, n47006, n47008, n47009, n47011,
    n47012, n47014, n47015, n47017, n47018, n47020,
    n47021, n47023, n47024, n47026, n47028, n47030,
    n47032, n47035, n47036, n47037, n47039, n47040,
    n47041, n47042, n47043, n47044, n47045, n47046,
    n47047, n47048, n47049, n47050, n47051, n47052,
    n47053, n47054, n47055, n47056, n47057, n47058,
    n47059, n47060, n47061, n47062, n47063, n47064,
    n47065, n47067, n47068, n47069, n47070, n47071,
    n47072, n47073, n47074, n47075, n47076, n47077,
    n47078, n47079, n47080, n47081, n47082, n47083,
    n47084, n47085, n47086, n47087, n47088, n47089,
    n47090, n47091, n47092, n47094, n47095, n47096,
    n47097, n47098, n47099, n47100, n47101, n47102,
    n47103, n47104, n47105, n47106, n47107, n47108,
    n47109, n47110, n47111, n47112, n47113, n47114,
    n47115, n47116, n47117, n47118, n47119, n47121,
    n47122, n47123, n47124, n47125, n47126, n47127,
    n47128, n47129, n47130, n47131, n47132, n47133,
    n47134, n47135, n47136, n47137, n47138, n47139,
    n47140, n47141, n47142, n47143, n47144, n47145,
    n47146, n47148, n47149, n47151, n47153, n47155,
    n47158, n47160, n47161, n47163, n47164, n47166,
    n47167, n47169, n47170, n47173, n47174, n47176,
    n47177, n47179, n47180, n47182, n47183, n47185,
    n47186, n47188, n47189, n47191, n47192, n47194,
    n47195, n47197, n47198, n47200, n47201, n47203,
    n47204, n47206, n47207, n47209, n47210, n47212,
    n47213, n47215, n47216, n47218, n47219, n47221,
    n47222, n47224, n47225, n47227, n47228, n47230,
    n47231, n47232, n47233, n47234, n47235, n47236,
    n47237, n47239, n47240, n47242, n47243, n47245,
    n47246, n47248, n47249, n47251, n47252, n47254,
    n47255, n47257, n47258, n47260, n47261, n47262,
    n47263, n47264, n47265, n47266, n47267, n47269,
    n47270, n47272, n47273, n47275, n47276, n47278,
    n47279, n47281, n47282, n47284, n47285, n47286,
    n47287, n47288, n47289, n47290, n47291, n47293,
    n47294, n47296, n47297, n47298, n47299, n47300,
    n47301, n47302, n47303, n47305, n47306, n47307,
    n47308, n47309, n47310, n47311, n47312, n47314,
    n47315, n47316, n47317, n47318, n47319, n47320,
    n47321, n47323, n47324, n47326, n47327, n47329,
    n47331, n47332, n47334, n47335, n47337, n47338,
    n47340, n47342, n47343, n47345, n47346, n47348,
    n47349, n47351, n47352, n47354, n47355, n47357,
    n47358, n47360, n47361, n47363, n47364, n47366,
    n47367, n47369, n47371, n47372, n47374, n47375,
    n47377, n47378, n47380, n47382, n47384, n47385,
    n47387, n47388, n47389, n47390, n47391, n47392,
    n47393, n47394, n47395, n47396, n47398, n47400,
    n47401, n47403, n47404, n47406, n47407, n47409,
    n47411, n47412, n47414, n47416, n47417, n47419,
    n47421, n47422, n47424, n47425, n47427, n47428,
    n47430, n47431, n47433, n47435, n47436, n47438,
    n47439, n47441, n47443, n47444, n47446, n47447,
    n47449, n47450, n47452, n47454, n47455, n47457,
    n47458, n47460, n47461, n47463, n47465, n47467,
    n47468, n47470, n47472, n47473, n47475, n47476,
    n47478, n47480, n47481, n47483, n47485, n47486,
    n47488, n47489, n47491, n47492, n47494, n47495,
    n47498, n47500, n47502, n47503, n47506;
  assign n2437 = ~pi332 & ~pi1144;
  assign n2438 = pi215 & ~n2437;
  assign n2439 = pi265 & ~pi332;
  assign n2440 = pi216 & ~n2439;
  assign n2441 = pi105 & pi228;
  assign n2442 = pi95 & ~pi479;
  assign n2443 = pi234 & n2442;
  assign n2444 = ~pi332 & ~n2443;
  assign n2445 = n2441 & n2444;
  assign n2446 = pi153 & ~pi332;
  assign n2447 = ~n2441 & n2446;
  assign n2448 = ~pi216 & ~n2447;
  assign n2449 = ~n2445 & n2448;
  assign n2450 = ~n2440 & ~n2449;
  assign n2451 = ~pi221 & ~n2450;
  assign n2452 = ~pi216 & pi833;
  assign n2453 = pi929 & n2452;
  assign n2454 = pi1144 & ~n2452;
  assign n2455 = ~pi332 & ~n2454;
  assign n2456 = ~n2453 & n2455;
  assign n2457 = pi221 & ~n2456;
  assign n2458 = ~n2451 & ~n2457;
  assign n2459 = ~pi215 & ~n2458;
  assign n2460 = ~n2438 & ~n2459;
  assign n2461 = ~pi32 & ~pi40;
  assign n2462 = ~pi58 & ~pi90;
  assign n2463 = ~pi88 & ~pi98;
  assign n2464 = ~pi50 & ~pi77;
  assign n2465 = n2463 & n2464;
  assign n2466 = ~pi102 & n2465;
  assign n2467 = ~pi65 & ~pi71;
  assign n2468 = ~pi83 & ~pi103;
  assign n2469 = ~pi67 & ~pi69;
  assign n2470 = ~pi66 & ~pi73;
  assign n2471 = ~pi68 & ~pi84;
  assign n2472 = ~pi82 & ~pi111;
  assign n2473 = ~pi36 & n2472;
  assign n2474 = n2471 & n2473;
  assign n2475 = ~pi61 & ~pi76;
  assign n2476 = ~pi85 & ~pi106;
  assign n2477 = n2475 & n2476;
  assign n2478 = ~pi48 & n2477;
  assign n2479 = ~pi89 & n2478;
  assign n2480 = ~pi49 & n2479;
  assign n2481 = ~pi104 & n2480;
  assign n2482 = ~pi45 & n2481;
  assign n2483 = n2474 & n2482;
  assign n2484 = n2470 & n2483;
  assign n2485 = n2469 & n2484;
  assign n2486 = n2468 & n2485;
  assign n2487 = n2467 & n2486;
  assign n2488 = ~pi63 & ~pi107;
  assign n2489 = n2487 & n2488;
  assign n2490 = ~pi64 & n2489;
  assign n2491 = ~pi81 & n2490;
  assign n2492 = n2466 & n2491;
  assign n2493 = ~pi53 & ~pi60;
  assign n2494 = ~pi86 & n2493;
  assign n2495 = ~pi97 & ~pi108;
  assign n2496 = ~pi46 & ~pi109;
  assign n2497 = n2495 & n2496;
  assign n2498 = ~pi110 & n2497;
  assign n2499 = ~pi94 & n2498;
  assign n2500 = n2494 & n2499;
  assign n2501 = ~pi47 & ~pi91;
  assign n2502 = n2500 & n2501;
  assign n2503 = n2492 & n2502;
  assign n2504 = n2462 & n2503;
  assign n2505 = ~pi93 & n2504;
  assign n2506 = ~pi72 & ~pi96;
  assign n2507 = ~pi35 & ~pi70;
  assign n2508 = ~pi51 & n2507;
  assign n2509 = n2506 & n2508;
  assign n2510 = n2505 & n2509;
  assign n2511 = n2461 & n2510;
  assign n2512 = ~pi95 & n2511;
  assign n2513 = ~n2442 & ~n2512;
  assign n2514 = pi234 & ~n2513;
  assign n2515 = ~pi40 & n2506;
  assign n2516 = ~pi32 & ~pi95;
  assign n2517 = n2515 & n2516;
  assign n2518 = ~pi70 & n2517;
  assign n2519 = ~pi35 & ~pi93;
  assign n2520 = n2504 & n2519;
  assign n2521 = n2518 & n2520;
  assign n2522 = ~pi51 & n2521;
  assign n2523 = ~pi234 & n2522;
  assign n2524 = ~n2514 & ~n2523;
  assign n2525 = pi137 & ~n2524;
  assign n2526 = n2444 & ~n2525;
  assign n2527 = ~pi216 & ~pi221;
  assign n2528 = ~pi215 & n2527;
  assign n2529 = ~n2447 & n2528;
  assign n2530 = ~n2526 & n2529;
  assign n2531 = ~pi56 & ~pi62;
  assign n2532 = ~pi38 & ~pi39;
  assign n2533 = ~pi100 & n2532;
  assign n2534 = ~pi54 & ~pi74;
  assign n2535 = ~pi75 & ~pi87;
  assign n2536 = ~pi92 & n2535;
  assign n2537 = n2534 & n2536;
  assign n2538 = ~pi55 & n2537;
  assign n2539 = n2533 & n2538;
  assign n2540 = n2531 & n2539;
  assign n2541 = n2530 & n2540;
  assign n2542 = ~pi59 & n2541;
  assign n2543 = n2460 & ~n2542;
  assign n2544 = pi57 & ~n2543;
  assign n2545 = n2460 & ~n2539;
  assign n2546 = ~pi105 & ~n2446;
  assign n2547 = pi105 & ~n2526;
  assign n2548 = ~n2546 & ~n2547;
  assign n2549 = pi228 & ~n2548;
  assign n2550 = ~pi332 & n2512;
  assign n2551 = ~pi137 & ~pi153;
  assign n2552 = n2550 & n2551;
  assign n2553 = pi137 & n2522;
  assign n2554 = n2446 & ~n2553;
  assign n2555 = ~pi228 & ~n2554;
  assign n2556 = ~n2552 & n2555;
  assign n2557 = ~n2549 & ~n2556;
  assign n2558 = ~pi216 & ~n2557;
  assign n2559 = ~n2440 & ~n2558;
  assign n2560 = ~pi221 & ~n2559;
  assign n2561 = ~n2457 & ~n2560;
  assign n2562 = ~pi215 & ~n2561;
  assign n2563 = ~n2438 & ~n2562;
  assign n2564 = n2539 & n2563;
  assign n2565 = ~n2545 & ~n2564;
  assign n2566 = ~pi56 & ~n2565;
  assign n2567 = pi62 & ~n2566;
  assign n2568 = pi56 & n2460;
  assign n2569 = n2567 & ~n2568;
  assign n2570 = pi56 & ~n2565;
  assign n2571 = ~pi87 & ~pi100;
  assign n2572 = ~pi38 & n2571;
  assign n2573 = ~pi75 & ~pi92;
  assign n2574 = n2572 & n2573;
  assign n2575 = n2534 & n2574;
  assign n2576 = ~pi39 & n2575;
  assign n2577 = n2460 & ~n2576;
  assign n2578 = pi228 & ~n2546;
  assign n2579 = ~pi332 & n2524;
  assign n2580 = pi105 & ~n2579;
  assign n2581 = n2578 & ~n2580;
  assign n2582 = ~pi228 & ~n2522;
  assign n2583 = n2446 & n2582;
  assign n2584 = ~pi216 & ~n2583;
  assign n2585 = ~n2581 & n2584;
  assign n2586 = ~n2440 & ~n2585;
  assign n2587 = ~pi221 & ~n2586;
  assign n2588 = ~n2457 & ~n2587;
  assign n2589 = ~pi215 & ~n2588;
  assign n2590 = ~n2438 & n2576;
  assign n2591 = ~n2589 & n2590;
  assign n2592 = pi55 & ~n2591;
  assign n2593 = ~n2577 & n2592;
  assign n2594 = pi299 & n2460;
  assign n2595 = ~pi224 & pi833;
  assign n2596 = pi222 & ~n2595;
  assign n2597 = ~pi223 & ~n2596;
  assign n2598 = n2437 & ~n2597;
  assign n2599 = pi224 & ~n2439;
  assign n2600 = ~pi222 & ~n2599;
  assign n2601 = ~pi332 & ~pi929;
  assign n2602 = n2595 & n2601;
  assign n2603 = ~n2600 & ~n2602;
  assign n2604 = ~pi223 & ~n2603;
  assign n2605 = ~n2598 & ~n2604;
  assign n2606 = ~pi299 & ~n2605;
  assign n2607 = ~pi222 & ~pi224;
  assign n2608 = ~pi223 & n2607;
  assign n2609 = ~n2444 & n2608;
  assign n2610 = n2606 & ~n2609;
  assign n2611 = ~n2594 & ~n2610;
  assign n2612 = ~n2535 & ~n2611;
  assign n2613 = pi92 & ~n2612;
  assign n2614 = ~pi38 & ~pi100;
  assign n2615 = ~pi39 & n2614;
  assign n2616 = ~n2611 & ~n2615;
  assign n2617 = ~n2526 & n2608;
  assign n2618 = ~n2605 & ~n2617;
  assign n2619 = ~pi299 & ~n2618;
  assign n2620 = pi299 & ~n2563;
  assign n2621 = ~n2619 & ~n2620;
  assign n2622 = n2615 & n2621;
  assign n2623 = ~n2616 & ~n2622;
  assign n2624 = n2535 & ~n2623;
  assign n2625 = n2613 & ~n2624;
  assign n2626 = ~pi152 & ~pi161;
  assign n2627 = ~pi166 & n2626;
  assign n2628 = ~pi146 & ~n2627;
  assign n2629 = ~pi210 & ~n2628;
  assign n2630 = pi95 & pi234;
  assign n2631 = ~pi137 & ~n2630;
  assign n2632 = ~n2629 & n2631;
  assign n2633 = ~n2524 & ~n2632;
  assign n2634 = ~pi332 & ~n2633;
  assign n2635 = pi105 & ~n2634;
  assign n2636 = n2578 & ~n2635;
  assign n2637 = n2553 & n2628;
  assign n2638 = n2446 & ~n2637;
  assign n2639 = ~pi137 & pi210;
  assign n2640 = n2550 & ~n2639;
  assign n2641 = ~pi252 & n2640;
  assign n2642 = ~n2628 & n2641;
  assign n2643 = n2638 & ~n2642;
  assign n2644 = pi252 & ~n2628;
  assign n2645 = ~n2629 & ~n2644;
  assign n2646 = n2552 & n2645;
  assign n2647 = ~n2643 & ~n2646;
  assign n2648 = ~pi228 & ~n2647;
  assign n2649 = ~pi216 & ~n2648;
  assign n2650 = ~n2636 & n2649;
  assign n2651 = ~n2440 & ~n2650;
  assign n2652 = ~pi221 & ~n2651;
  assign n2653 = ~n2457 & ~n2652;
  assign n2654 = ~pi215 & ~n2653;
  assign n2655 = ~n2438 & ~n2654;
  assign n2656 = pi299 & ~n2655;
  assign n2657 = ~pi144 & ~pi174;
  assign n2658 = ~pi189 & n2657;
  assign n2659 = ~pi223 & ~n2658;
  assign n2660 = pi142 & ~pi198;
  assign n2661 = ~pi137 & ~n2660;
  assign n2662 = ~n2524 & ~n2661;
  assign n2663 = n2444 & ~n2662;
  assign n2664 = n2659 & ~n2663;
  assign n2665 = pi234 & ~pi332;
  assign n2666 = ~pi137 & pi198;
  assign n2667 = ~pi95 & n2666;
  assign n2668 = ~n2513 & ~n2667;
  assign n2669 = n2665 & ~n2668;
  assign n2670 = ~pi234 & ~pi332;
  assign n2671 = n2522 & ~n2666;
  assign n2672 = n2670 & ~n2671;
  assign n2673 = ~pi223 & n2658;
  assign n2674 = ~n2672 & n2673;
  assign n2675 = ~n2669 & n2674;
  assign n2676 = ~n2664 & ~n2675;
  assign n2677 = n2607 & ~n2676;
  assign n2678 = ~n2605 & ~n2677;
  assign n2679 = ~pi299 & ~n2678;
  assign n2680 = ~n2656 & ~n2679;
  assign n2681 = n2532 & n2680;
  assign n2682 = ~n2532 & ~n2611;
  assign n2683 = pi100 & ~n2682;
  assign n2684 = ~n2681 & n2683;
  assign n2685 = pi39 & ~n2621;
  assign n2686 = ~pi40 & ~pi72;
  assign n2687 = ~pi46 & ~pi94;
  assign n2688 = n2495 & n2687;
  assign n2689 = n2494 & n2688;
  assign n2690 = n2492 & n2689;
  assign n2691 = ~pi109 & ~pi110;
  assign n2692 = ~pi58 & ~pi91;
  assign n2693 = ~pi47 & n2692;
  assign n2694 = n2691 & n2693;
  assign n2695 = n2690 & n2694;
  assign n2696 = ~pi90 & ~pi93;
  assign n2697 = ~pi96 & n2508;
  assign n2698 = n2696 & n2697;
  assign n2699 = n2695 & n2698;
  assign n2700 = n2686 & n2699;
  assign n2701 = pi225 & n2700;
  assign n2702 = pi32 & ~n2701;
  assign n2703 = ~pi95 & ~n2702;
  assign n2704 = pi60 & n2492;
  assign n2705 = ~pi53 & ~n2704;
  assign n2706 = ~pi86 & ~pi94;
  assign n2707 = ~pi60 & n2492;
  assign n2708 = pi53 & ~n2707;
  assign n2709 = n2706 & ~n2708;
  assign n2710 = ~n2705 & n2709;
  assign n2711 = ~pi110 & n2693;
  assign n2712 = n2497 & n2711;
  assign n2713 = ~pi90 & n2712;
  assign n2714 = ~pi93 & n2713;
  assign n2715 = n2710 & n2714;
  assign n2716 = ~pi35 & ~n2715;
  assign n2717 = pi35 & ~n2505;
  assign n2718 = pi35 & n2505;
  assign n2719 = ~pi225 & n2718;
  assign n2720 = ~pi70 & ~n2719;
  assign n2721 = ~pi51 & n2720;
  assign n2722 = ~n2717 & n2721;
  assign n2723 = ~n2716 & n2722;
  assign n2724 = ~pi96 & ~n2723;
  assign n2725 = ~pi47 & n2500;
  assign n2726 = n2492 & n2725;
  assign n2727 = n2692 & n2696;
  assign n2728 = n2508 & n2727;
  assign n2729 = n2726 & n2728;
  assign n2730 = pi96 & ~n2729;
  assign n2731 = n2686 & ~n2730;
  assign n2732 = ~n2724 & n2731;
  assign n2733 = ~pi32 & ~n2732;
  assign n2734 = n2703 & ~n2733;
  assign n2735 = ~n2442 & ~n2734;
  assign n2736 = ~pi137 & n2735;
  assign n2737 = pi40 & n2510;
  assign n2738 = ~pi32 & ~n2737;
  assign n2739 = pi72 & ~n2699;
  assign n2740 = ~pi40 & ~n2739;
  assign n2741 = ~pi70 & n2520;
  assign n2742 = pi51 & ~n2741;
  assign n2743 = ~pi96 & ~n2742;
  assign n2744 = ~pi51 & pi70;
  assign n2745 = n2743 & ~n2744;
  assign n2746 = ~n2717 & ~n2719;
  assign n2747 = pi93 & n2504;
  assign n2748 = ~pi35 & ~n2747;
  assign n2749 = pi91 & n2726;
  assign n2750 = n2462 & ~n2749;
  assign n2751 = ~pi109 & n2690;
  assign n2752 = pi110 & ~n2751;
  assign n2753 = pi47 & n2492;
  assign n2754 = n2500 & n2753;
  assign n2755 = pi47 & ~n2754;
  assign n2756 = ~pi91 & ~n2755;
  assign n2757 = ~n2752 & n2756;
  assign n2758 = ~pi47 & ~pi110;
  assign n2759 = pi109 & ~n2690;
  assign n2760 = ~pi50 & n2493;
  assign n2761 = ~pi102 & n2491;
  assign n2762 = n2463 & n2761;
  assign n2763 = ~pi77 & n2762;
  assign n2764 = n2760 & n2763;
  assign n2765 = n2706 & n2764;
  assign n2766 = ~pi97 & n2765;
  assign n2767 = pi108 & ~n2766;
  assign n2768 = ~pi46 & ~n2767;
  assign n2769 = pi97 & ~n2765;
  assign n2770 = ~pi86 & pi94;
  assign n2771 = n2764 & n2770;
  assign n2772 = ~pi97 & ~n2771;
  assign n2773 = pi86 & ~n2764;
  assign n2774 = ~pi94 & ~n2773;
  assign n2775 = pi77 & n2762;
  assign n2776 = ~pi50 & ~n2775;
  assign n2777 = pi81 & ~n2490;
  assign n2778 = pi102 & ~n2491;
  assign n2779 = ~n2777 & ~n2778;
  assign n2780 = pi64 & ~n2489;
  assign n2781 = pi71 & ~n2486;
  assign n2782 = ~pi65 & ~n2781;
  assign n2783 = ~pi67 & n2484;
  assign n2784 = pi69 & ~n2783;
  assign n2785 = pi83 & ~n2485;
  assign n2786 = ~pi103 & ~n2785;
  assign n2787 = ~n2784 & n2786;
  assign n2788 = ~pi69 & ~pi83;
  assign n2789 = pi67 & ~n2484;
  assign n2790 = n2470 & n2482;
  assign n2791 = ~pi84 & n2790;
  assign n2792 = ~pi68 & n2791;
  assign n2793 = n2472 & n2792;
  assign n2794 = pi36 & ~n2793;
  assign n2795 = ~pi36 & ~pi67;
  assign n2796 = ~pi68 & ~pi111;
  assign n2797 = pi82 & n2796;
  assign n2798 = n2791 & n2797;
  assign n2799 = pi111 & ~n2792;
  assign n2800 = ~pi82 & ~n2799;
  assign n2801 = pi84 & ~n2790;
  assign n2802 = pi85 & pi106;
  assign n2803 = n2475 & ~n2802;
  assign n2804 = pi61 & pi76;
  assign n2805 = n2476 & ~n2804;
  assign n2806 = ~n2803 & ~n2805;
  assign n2807 = ~pi48 & ~n2806;
  assign n2808 = ~n2477 & ~n2807;
  assign n2809 = pi89 & ~n2478;
  assign n2810 = ~pi49 & ~n2809;
  assign n2811 = ~n2808 & n2810;
  assign n2812 = ~n2479 & ~n2811;
  assign n2813 = ~pi45 & ~n2812;
  assign n2814 = ~n2481 & ~n2813;
  assign n2815 = pi104 & ~n2480;
  assign n2816 = ~n2482 & ~n2815;
  assign n2817 = ~n2814 & n2816;
  assign n2818 = n2470 & ~n2817;
  assign n2819 = pi66 & pi73;
  assign n2820 = ~n2470 & ~n2482;
  assign n2821 = ~n2819 & ~n2820;
  assign n2822 = ~n2818 & n2821;
  assign n2823 = ~pi84 & ~n2822;
  assign n2824 = ~n2801 & ~n2823;
  assign n2825 = n2796 & ~n2824;
  assign n2826 = pi68 & ~n2791;
  assign n2827 = ~n2825 & ~n2826;
  assign n2828 = n2800 & n2827;
  assign n2829 = ~n2798 & ~n2828;
  assign n2830 = n2795 & n2829;
  assign n2831 = ~n2794 & ~n2830;
  assign n2832 = ~n2789 & n2831;
  assign n2833 = n2788 & ~n2832;
  assign n2834 = n2787 & ~n2833;
  assign n2835 = pi103 & n2485;
  assign n2836 = ~pi83 & n2835;
  assign n2837 = ~pi71 & ~n2836;
  assign n2838 = ~n2834 & n2837;
  assign n2839 = n2782 & ~n2838;
  assign n2840 = ~pi107 & ~n2839;
  assign n2841 = ~pi63 & pi107;
  assign n2842 = n2487 & n2841;
  assign n2843 = ~n2488 & ~n2842;
  assign n2844 = ~n2840 & ~n2843;
  assign n2845 = pi65 & ~pi71;
  assign n2846 = n2486 & n2845;
  assign n2847 = ~n2843 & n2846;
  assign n2848 = ~pi64 & ~n2847;
  assign n2849 = ~n2844 & n2848;
  assign n2850 = ~n2780 & ~n2849;
  assign n2851 = ~pi81 & ~pi102;
  assign n2852 = ~n2850 & n2851;
  assign n2853 = pi63 & n2487;
  assign n2854 = ~pi107 & n2853;
  assign n2855 = ~pi64 & ~n2854;
  assign n2856 = ~n2844 & n2855;
  assign n2857 = ~n2780 & ~n2856;
  assign n2858 = n2852 & ~n2857;
  assign n2859 = n2779 & ~n2858;
  assign n2860 = n2463 & ~n2859;
  assign n2861 = pi98 & ~n2761;
  assign n2862 = ~pi98 & n2761;
  assign n2863 = pi88 & ~n2862;
  assign n2864 = ~pi77 & ~n2863;
  assign n2865 = ~n2861 & n2864;
  assign n2866 = ~n2860 & n2865;
  assign n2867 = n2776 & ~n2866;
  assign n2868 = pi50 & ~n2763;
  assign n2869 = ~pi60 & ~n2868;
  assign n2870 = ~n2867 & n2869;
  assign n2871 = n2705 & ~n2870;
  assign n2872 = ~n2708 & ~n2871;
  assign n2873 = ~pi86 & ~n2872;
  assign n2874 = n2774 & ~n2873;
  assign n2875 = n2772 & ~n2874;
  assign n2876 = ~n2769 & ~n2875;
  assign n2877 = ~pi108 & ~n2876;
  assign n2878 = n2768 & ~n2877;
  assign n2879 = pi46 & n2765;
  assign n2880 = n2495 & n2879;
  assign n2881 = ~pi109 & ~n2880;
  assign n2882 = ~n2878 & n2881;
  assign n2883 = ~n2759 & ~n2882;
  assign n2884 = n2758 & ~n2883;
  assign n2885 = n2757 & ~n2884;
  assign n2886 = n2750 & ~n2885;
  assign n2887 = pi58 & ~n2503;
  assign n2888 = pi90 & ~n2695;
  assign n2889 = ~pi93 & ~n2888;
  assign n2890 = ~n2887 & n2889;
  assign n2891 = ~n2886 & n2890;
  assign n2892 = n2748 & ~n2891;
  assign n2893 = n2746 & ~n2892;
  assign n2894 = ~pi51 & ~n2893;
  assign n2895 = n2745 & ~n2894;
  assign n2896 = ~pi72 & ~n2895;
  assign n2897 = n2740 & ~n2896;
  assign n2898 = n2738 & ~n2897;
  assign n2899 = pi96 & n2729;
  assign n2900 = ~pi51 & ~pi72;
  assign n2901 = n2520 & n2900;
  assign n2902 = ~pi40 & n2901;
  assign n2903 = n2899 & n2902;
  assign n2904 = n2898 & ~n2903;
  assign n2905 = ~n2702 & ~n2904;
  assign n2906 = ~pi95 & ~n2905;
  assign n2907 = pi95 & ~n2511;
  assign n2908 = pi479 & n2907;
  assign n2909 = ~n2906 & ~n2908;
  assign n2910 = pi137 & ~n2909;
  assign n2911 = ~n2736 & ~n2910;
  assign n2912 = pi198 & ~n2911;
  assign n2913 = ~pi833 & pi957;
  assign n2914 = pi1091 & ~n2913;
  assign n2915 = pi841 & n2504;
  assign n2916 = ~pi93 & n2915;
  assign n2917 = ~pi51 & ~pi70;
  assign n2918 = n2506 & n2917;
  assign n2919 = ~pi40 & n2918;
  assign n2920 = ~pi35 & n2919;
  assign n2921 = n2916 & n2920;
  assign n2922 = pi225 & n2921;
  assign n2923 = pi32 & ~n2922;
  assign n2924 = ~n2904 & ~n2923;
  assign n2925 = ~pi95 & ~n2924;
  assign n2926 = ~n2908 & ~n2925;
  assign n2927 = pi137 & ~n2926;
  assign n2928 = ~pi95 & ~n2923;
  assign n2929 = ~n2733 & n2928;
  assign n2930 = ~n2442 & ~n2929;
  assign n2931 = ~pi137 & n2930;
  assign n2932 = ~n2927 & ~n2931;
  assign n2933 = ~n2914 & n2932;
  assign n2934 = pi1092 & pi1093;
  assign n2935 = pi829 & pi950;
  assign n2936 = n2934 & n2935;
  assign n2937 = ~n2930 & ~n2936;
  assign n2938 = n2496 & n2501;
  assign n2939 = ~pi108 & ~n2769;
  assign n2940 = ~pi110 & n2939;
  assign n2941 = ~pi93 & n2462;
  assign n2942 = ~pi97 & ~n2710;
  assign n2943 = n2941 & ~n2942;
  assign n2944 = n2940 & n2943;
  assign n2945 = n2938 & n2944;
  assign n2946 = ~pi35 & ~n2945;
  assign n2947 = n2722 & ~n2946;
  assign n2948 = ~pi96 & ~n2947;
  assign n2949 = n2731 & ~n2948;
  assign n2950 = ~pi32 & ~n2949;
  assign n2951 = n2928 & ~n2950;
  assign n2952 = ~n2442 & ~n2951;
  assign n2953 = n2936 & ~n2952;
  assign n2954 = ~pi137 & ~n2953;
  assign n2955 = ~n2937 & n2954;
  assign n2956 = ~n2927 & ~n2955;
  assign n2957 = n2914 & n2956;
  assign n2958 = ~n2933 & ~n2957;
  assign n2959 = ~pi198 & n2958;
  assign n2960 = ~n2912 & ~n2959;
  assign n2961 = pi142 & n2960;
  assign n2962 = ~pi198 & ~n2932;
  assign n2963 = ~pi142 & ~n2912;
  assign n2964 = ~n2962 & n2963;
  assign n2965 = ~n2961 & ~n2964;
  assign n2966 = n2665 & n2965;
  assign n2967 = n2515 & n2723;
  assign n2968 = ~pi32 & ~n2967;
  assign n2969 = n2703 & ~n2968;
  assign n2970 = ~pi137 & ~n2969;
  assign n2971 = ~n2442 & ~n2907;
  assign n2972 = ~n2702 & ~n2898;
  assign n2973 = ~pi95 & ~n2972;
  assign n2974 = n2971 & ~n2973;
  assign n2975 = pi137 & ~n2974;
  assign n2976 = ~n2970 & ~n2975;
  assign n2977 = pi198 & ~n2976;
  assign n2978 = n2914 & n2936;
  assign n2979 = n2716 & ~n2978;
  assign n2980 = n2919 & ~n2979;
  assign n2981 = n2946 & n2978;
  assign n2982 = n2746 & ~n2981;
  assign n2983 = n2980 & n2982;
  assign n2984 = ~pi32 & ~n2983;
  assign n2985 = n2928 & ~n2984;
  assign n2986 = ~pi137 & ~n2985;
  assign n2987 = ~n2898 & ~n2923;
  assign n2988 = ~pi95 & ~n2987;
  assign n2989 = n2971 & ~n2988;
  assign n2990 = pi137 & ~n2989;
  assign n2991 = ~n2986 & ~n2990;
  assign n2992 = ~pi198 & ~n2991;
  assign n2993 = ~n2977 & ~n2992;
  assign n2994 = pi142 & n2993;
  assign n2995 = n2928 & ~n2968;
  assign n2996 = ~pi137 & ~n2995;
  assign n2997 = ~n2990 & ~n2996;
  assign n2998 = ~pi198 & ~n2997;
  assign n2999 = ~pi142 & ~n2977;
  assign n3000 = ~n2998 & n2999;
  assign n3001 = n2670 & ~n3000;
  assign n3002 = ~n2994 & n3001;
  assign n3003 = n2659 & ~n3002;
  assign n3004 = ~n2966 & n3003;
  assign n3005 = pi234 & n2960;
  assign n3006 = ~pi234 & n2993;
  assign n3007 = ~pi332 & ~n3006;
  assign n3008 = ~n3005 & n3007;
  assign n3009 = n2673 & ~n3008;
  assign n3010 = ~n3004 & ~n3009;
  assign n3011 = n2607 & ~n3010;
  assign n3012 = n2606 & ~n3011;
  assign n3013 = pi210 & ~n2911;
  assign n3014 = ~pi210 & n2958;
  assign n3015 = ~n3013 & ~n3014;
  assign n3016 = pi234 & n3015;
  assign n3017 = pi210 & ~n2976;
  assign n3018 = ~pi210 & ~n2991;
  assign n3019 = ~n3017 & ~n3018;
  assign n3020 = ~pi234 & n3019;
  assign n3021 = ~pi332 & ~n3020;
  assign n3022 = ~n3016 & n3021;
  assign n3023 = n2627 & ~n3022;
  assign n3024 = pi146 & n3015;
  assign n3025 = ~pi210 & ~n2932;
  assign n3026 = ~pi146 & ~n3013;
  assign n3027 = ~n3025 & n3026;
  assign n3028 = ~n3024 & ~n3027;
  assign n3029 = n2665 & n3028;
  assign n3030 = pi146 & n3019;
  assign n3031 = ~pi210 & ~n2997;
  assign n3032 = ~pi146 & ~n3017;
  assign n3033 = ~n3031 & n3032;
  assign n3034 = n2670 & ~n3033;
  assign n3035 = ~n3030 & n3034;
  assign n3036 = ~n2627 & ~n3035;
  assign n3037 = ~n3029 & n3036;
  assign n3038 = ~n3023 & ~n3037;
  assign n3039 = pi105 & ~n3038;
  assign n3040 = ~n2546 & ~n3039;
  assign n3041 = pi228 & ~n3040;
  assign n3042 = ~pi146 & ~pi210;
  assign n3043 = pi93 & ~n2504;
  assign n3044 = ~pi35 & ~n3043;
  assign n3045 = ~n2887 & ~n2888;
  assign n3046 = ~pi53 & n2870;
  assign n3047 = ~pi86 & ~n3046;
  assign n3048 = n2774 & ~n3047;
  assign n3049 = n2772 & ~n3048;
  assign n3050 = ~n2769 & ~n3049;
  assign n3051 = ~pi108 & ~n3050;
  assign n3052 = n2768 & ~n3051;
  assign n3053 = ~pi109 & ~n3052;
  assign n3054 = ~n2759 & ~n3053;
  assign n3055 = n2758 & ~n3054;
  assign n3056 = n2757 & ~n3055;
  assign n3057 = n2750 & ~n3056;
  assign n3058 = n3045 & ~n3057;
  assign n3059 = ~pi93 & ~n3058;
  assign n3060 = n3044 & ~n3059;
  assign n3061 = n2721 & ~n3060;
  assign n3062 = pi70 & ~n2520;
  assign n3063 = n2743 & ~n3062;
  assign n3064 = ~n3061 & n3063;
  assign n3065 = ~pi72 & ~n2899;
  assign n3066 = ~n3064 & n3065;
  assign n3067 = n2740 & ~n3066;
  assign n3068 = n2738 & ~n3067;
  assign n3069 = pi225 & pi841;
  assign n3070 = n2700 & ~n3069;
  assign n3071 = pi32 & ~n3070;
  assign n3072 = ~n3068 & ~n3071;
  assign n3073 = ~pi95 & ~n3072;
  assign n3074 = ~n2907 & ~n3073;
  assign n3075 = ~pi137 & ~n3074;
  assign n3076 = ~pi95 & ~n3071;
  assign n3077 = ~pi51 & ~pi96;
  assign n3078 = ~n3062 & n3077;
  assign n3079 = ~n2720 & n3078;
  assign n3080 = n2686 & n3079;
  assign n3081 = ~pi32 & ~n3080;
  assign n3082 = n3076 & ~n3081;
  assign n3083 = pi137 & ~n3082;
  assign n3084 = ~pi95 & n2461;
  assign n3085 = ~pi72 & n3084;
  assign n3086 = n2899 & n3085;
  assign n3087 = ~n2442 & ~n3086;
  assign n3088 = ~n2907 & ~n3087;
  assign n3089 = n3083 & ~n3088;
  assign n3090 = ~n3075 & ~n3089;
  assign n3091 = n3042 & ~n3090;
  assign n3092 = ~n2978 & n3068;
  assign n3093 = n2738 & n2978;
  assign n3094 = ~pi97 & ~n3049;
  assign n3095 = ~pi108 & ~n3094;
  assign n3096 = n2768 & ~n3095;
  assign n3097 = ~pi109 & ~n3096;
  assign n3098 = ~n2759 & ~n3097;
  assign n3099 = n2758 & ~n3098;
  assign n3100 = n2757 & ~n3099;
  assign n3101 = n2750 & ~n3100;
  assign n3102 = n3045 & ~n3101;
  assign n3103 = ~pi93 & ~n3102;
  assign n3104 = n3044 & ~n3103;
  assign n3105 = n2721 & ~n3104;
  assign n3106 = n3063 & ~n3105;
  assign n3107 = n3065 & ~n3106;
  assign n3108 = n2740 & ~n3107;
  assign n3109 = n3093 & ~n3108;
  assign n3110 = ~n3092 & ~n3109;
  assign n3111 = ~n3071 & n3110;
  assign n3112 = ~pi95 & ~n3111;
  assign n3113 = ~n2907 & ~n3112;
  assign n3114 = ~pi137 & ~n3113;
  assign n3115 = ~n3089 & ~n3114;
  assign n3116 = ~pi210 & ~n3115;
  assign n3117 = pi146 & n3116;
  assign n3118 = ~pi137 & ~n2907;
  assign n3119 = ~pi225 & n2700;
  assign n3120 = pi32 & ~n3119;
  assign n3121 = ~n3068 & ~n3120;
  assign n3122 = ~pi95 & ~n3121;
  assign n3123 = n3118 & ~n3122;
  assign n3124 = ~pi95 & ~n3120;
  assign n3125 = ~n3081 & n3124;
  assign n3126 = ~n3088 & ~n3125;
  assign n3127 = pi137 & ~n3126;
  assign n3128 = ~n3123 & ~n3127;
  assign n3129 = pi210 & n3128;
  assign n3130 = n2670 & ~n3129;
  assign n3131 = ~n3117 & n3130;
  assign n3132 = ~n3091 & n3131;
  assign n3133 = ~pi72 & ~n3064;
  assign n3134 = n2740 & ~n3133;
  assign n3135 = n2738 & ~n3134;
  assign n3136 = ~n3120 & ~n3135;
  assign n3137 = ~pi95 & ~n3136;
  assign n3138 = ~pi137 & n2971;
  assign n3139 = ~n3137 & n3138;
  assign n3140 = pi137 & n3125;
  assign n3141 = ~n3139 & ~n3140;
  assign n3142 = pi210 & n3141;
  assign n3143 = n2665 & ~n3142;
  assign n3144 = ~n3071 & ~n3135;
  assign n3145 = ~pi95 & ~n3144;
  assign n3146 = n2971 & ~n3145;
  assign n3147 = ~pi137 & ~n3146;
  assign n3148 = ~n3083 & ~n3147;
  assign n3149 = n3042 & ~n3148;
  assign n3150 = ~n2978 & n3135;
  assign n3151 = ~pi72 & ~n3106;
  assign n3152 = n2740 & ~n3151;
  assign n3153 = n3093 & ~n3152;
  assign n3154 = ~n3071 & ~n3153;
  assign n3155 = ~n3150 & n3154;
  assign n3156 = ~pi95 & ~n3155;
  assign n3157 = n2971 & ~n3156;
  assign n3158 = ~pi137 & ~n3157;
  assign n3159 = ~n3083 & ~n3158;
  assign n3160 = ~pi210 & ~n3159;
  assign n3161 = pi146 & n3160;
  assign n3162 = ~n3149 & ~n3161;
  assign n3163 = n3143 & n3162;
  assign n3164 = ~n2627 & ~n3163;
  assign n3165 = ~n3132 & n3164;
  assign n3166 = n3143 & ~n3160;
  assign n3167 = ~n3116 & n3130;
  assign n3168 = n2627 & ~n3167;
  assign n3169 = ~n3166 & n3168;
  assign n3170 = ~pi153 & ~n3169;
  assign n3171 = ~n3165 & n3170;
  assign n3172 = ~pi109 & ~n2878;
  assign n3173 = ~n2759 & ~n3172;
  assign n3174 = n2758 & ~n3173;
  assign n3175 = n2757 & ~n3174;
  assign n3176 = n2750 & ~n3175;
  assign n3177 = n2890 & ~n3176;
  assign n3178 = n2748 & ~n3177;
  assign n3179 = n2746 & ~n3178;
  assign n3180 = ~pi51 & ~n3179;
  assign n3181 = n2745 & ~n3180;
  assign n3182 = ~pi72 & ~n3181;
  assign n3183 = n2740 & ~n3182;
  assign n3184 = n2738 & ~n3183;
  assign n3185 = ~n2903 & n3184;
  assign n3186 = ~n2923 & ~n3185;
  assign n3187 = ~pi95 & ~n3186;
  assign n3188 = ~n2907 & ~n3187;
  assign n3189 = pi137 & ~n3188;
  assign n3190 = ~n2628 & n2914;
  assign n3191 = ~n2937 & n3190;
  assign n3192 = ~n2907 & ~n3191;
  assign n3193 = ~n2930 & n3192;
  assign n3194 = ~n2907 & n3190;
  assign n3195 = n2953 & n3194;
  assign n3196 = ~pi137 & ~n3195;
  assign n3197 = ~n3193 & n3196;
  assign n3198 = ~n3189 & ~n3197;
  assign n3199 = ~pi210 & ~n3198;
  assign n3200 = pi234 & ~n3199;
  assign n3201 = ~n2628 & n2986;
  assign n3202 = ~n2923 & ~n3184;
  assign n3203 = ~pi95 & ~n3202;
  assign n3204 = n2971 & ~n3203;
  assign n3205 = pi137 & ~n3204;
  assign n3206 = n2628 & n2996;
  assign n3207 = ~pi210 & ~n3206;
  assign n3208 = ~pi234 & n3207;
  assign n3209 = ~n3205 & n3208;
  assign n3210 = ~n3201 & n3209;
  assign n3211 = ~n2702 & ~n3184;
  assign n3212 = ~pi95 & ~n3211;
  assign n3213 = n2971 & ~n3212;
  assign n3214 = pi137 & ~n3213;
  assign n3215 = ~n2970 & ~n3214;
  assign n3216 = pi210 & n3215;
  assign n3217 = ~n3210 & ~n3216;
  assign n3218 = ~n3200 & n3217;
  assign n3219 = ~n2702 & ~n3185;
  assign n3220 = ~pi95 & ~n3219;
  assign n3221 = pi137 & ~n2907;
  assign n3222 = ~n3220 & n3221;
  assign n3223 = ~n2735 & n3118;
  assign n3224 = pi210 & ~n3223;
  assign n3225 = pi234 & n3224;
  assign n3226 = ~n3222 & n3225;
  assign n3227 = ~n3218 & ~n3226;
  assign n3228 = n2446 & ~n3227;
  assign n3229 = ~pi228 & ~n3228;
  assign n3230 = ~n3171 & n3229;
  assign n3231 = ~n3041 & ~n3230;
  assign n3232 = ~pi216 & ~n3231;
  assign n3233 = ~n2440 & ~n3232;
  assign n3234 = ~pi221 & ~n3233;
  assign n3235 = ~n2457 & ~n3234;
  assign n3236 = ~pi215 & ~n3235;
  assign n3237 = ~n2438 & ~n3236;
  assign n3238 = pi299 & n3237;
  assign n3239 = ~pi39 & ~n3238;
  assign n3240 = ~n3012 & n3239;
  assign n3241 = ~pi38 & ~n3240;
  assign n3242 = ~n2685 & n3241;
  assign n3243 = n2460 & ~n2530;
  assign n3244 = pi299 & ~n3243;
  assign n3245 = ~n2619 & ~n3244;
  assign n3246 = ~pi39 & ~n3245;
  assign n3247 = pi39 & n2611;
  assign n3248 = ~n3246 & ~n3247;
  assign n3249 = pi38 & n3248;
  assign n3250 = ~pi100 & ~n3249;
  assign n3251 = ~n3242 & n3250;
  assign n3252 = ~n2684 & ~n3251;
  assign n3253 = ~pi87 & n3252;
  assign n3254 = pi87 & ~n2623;
  assign n3255 = ~pi75 & ~n3254;
  assign n3256 = ~n3253 & n3255;
  assign n3257 = ~pi39 & ~pi87;
  assign n3258 = n2614 & n3257;
  assign n3259 = ~n2611 & ~n3258;
  assign n3260 = pi75 & ~n3259;
  assign n3261 = n2448 & ~n2636;
  assign n3262 = ~n2440 & ~n3261;
  assign n3263 = ~pi221 & ~n3262;
  assign n3264 = ~n2457 & ~n3263;
  assign n3265 = ~pi215 & ~n3264;
  assign n3266 = ~n2438 & ~n3265;
  assign n3267 = pi299 & ~n3266;
  assign n3268 = ~n2679 & n3258;
  assign n3269 = ~n3267 & n3268;
  assign n3270 = n3260 & ~n3269;
  assign n3271 = ~n3256 & ~n3270;
  assign n3272 = ~pi92 & ~n3271;
  assign n3273 = ~pi54 & ~n3272;
  assign n3274 = ~n2625 & n3273;
  assign n3275 = n2573 & n3258;
  assign n3276 = n2611 & ~n3275;
  assign n3277 = n2574 & n3246;
  assign n3278 = ~n3276 & ~n3277;
  assign n3279 = pi54 & n3278;
  assign n3280 = ~pi74 & ~n3279;
  assign n3281 = ~n3274 & n3280;
  assign n3282 = ~pi54 & n3278;
  assign n3283 = pi54 & ~n2611;
  assign n3284 = pi74 & ~n3283;
  assign n3285 = ~n3282 & n3284;
  assign n3286 = ~n3281 & ~n3285;
  assign n3287 = ~pi55 & ~n3286;
  assign n3288 = ~pi56 & ~n3287;
  assign n3289 = ~n2593 & n3288;
  assign n3290 = ~pi62 & ~n3289;
  assign n3291 = ~n2570 & n3290;
  assign n3292 = ~n2569 & ~n3291;
  assign n3293 = ~pi59 & n3292;
  assign n3294 = pi59 & n2460;
  assign n3295 = ~n2541 & n3294;
  assign n3296 = ~pi57 & ~n3295;
  assign n3297 = ~n3293 & n3296;
  assign po153 = n2544 | n3297;
  assign n3299 = pi215 & pi1146;
  assign n3300 = pi216 & ~pi221;
  assign n3301 = pi276 & n3300;
  assign n3302 = ~pi939 & n2452;
  assign n3303 = ~pi1146 & ~n2452;
  assign n3304 = pi221 & ~n3303;
  assign n3305 = ~n3302 & n3304;
  assign n3306 = ~n3301 & ~n3305;
  assign n3307 = ~pi215 & ~n3306;
  assign n3308 = ~n3299 & ~n3307;
  assign n3309 = pi154 & ~n3308;
  assign n3310 = ~n2441 & n2528;
  assign n3311 = n3308 & ~n3310;
  assign n3312 = ~pi154 & ~n3311;
  assign n3313 = ~n3309 & ~n3312;
  assign n3314 = ~pi56 & n2538;
  assign n3315 = n2533 & n3314;
  assign n3316 = ~n3313 & ~n3315;
  assign n3317 = ~n3299 & ~n3305;
  assign n3318 = ~pi216 & ~pi228;
  assign n3319 = n3317 & n3318;
  assign n3320 = n2522 & n3319;
  assign n3321 = ~n3309 & n3320;
  assign n3322 = ~pi55 & n2576;
  assign n3323 = ~n3313 & n3322;
  assign n3324 = ~n3321 & n3323;
  assign n3325 = ~n3316 & ~n3324;
  assign n3326 = pi62 & ~n3325;
  assign n3327 = ~pi57 & ~pi59;
  assign n3328 = ~n2539 & ~n3313;
  assign n3329 = pi56 & ~n3328;
  assign n3330 = ~n3324 & n3329;
  assign n3331 = pi299 & ~n3313;
  assign n3332 = ~pi222 & pi224;
  assign n3333 = pi276 & n3332;
  assign n3334 = ~pi1146 & ~n2595;
  assign n3335 = ~pi939 & n2595;
  assign n3336 = ~n3334 & ~n3335;
  assign n3337 = pi222 & n3336;
  assign n3338 = ~pi223 & ~n3337;
  assign n3339 = ~n3333 & n3338;
  assign n3340 = pi223 & ~pi1146;
  assign n3341 = ~pi299 & ~n3340;
  assign n3342 = ~n3339 & n3341;
  assign n3343 = ~n3331 & ~n3342;
  assign n3344 = ~n2534 & n3343;
  assign n3345 = n2533 & n2535;
  assign n3346 = n3343 & ~n3345;
  assign n3347 = pi299 & ~n3308;
  assign n3348 = ~n3342 & ~n3347;
  assign n3349 = pi154 & ~n3348;
  assign n3350 = ~pi38 & ~n3349;
  assign n3351 = ~pi39 & ~pi100;
  assign n3352 = pi299 & ~n3311;
  assign n3353 = ~n3320 & n3352;
  assign n3354 = ~n3342 & ~n3353;
  assign n3355 = ~pi154 & ~n3354;
  assign n3356 = n3351 & ~n3355;
  assign n3357 = n3350 & n3356;
  assign n3358 = n2535 & n3357;
  assign n3359 = pi92 & ~n3358;
  assign n3360 = ~n3346 & n3359;
  assign n3361 = pi75 & n3343;
  assign n3362 = ~n2615 & n3343;
  assign n3363 = ~n3357 & ~n3362;
  assign n3364 = pi87 & ~n3363;
  assign n3365 = pi38 & n3343;
  assign n3366 = pi39 & ~n2522;
  assign n3367 = ~pi70 & n3178;
  assign n3368 = ~n2717 & ~n3367;
  assign n3369 = ~n3062 & n3368;
  assign n3370 = ~pi51 & ~n3369;
  assign n3371 = n2743 & ~n3370;
  assign n3372 = n3065 & ~n3371;
  assign n3373 = ~n2739 & ~n3372;
  assign n3374 = n2461 & ~n3373;
  assign n3375 = pi40 & ~n2510;
  assign n3376 = pi32 & ~n2700;
  assign n3377 = ~n3375 & ~n3376;
  assign n3378 = ~n3374 & n3377;
  assign n3379 = ~pi95 & ~n3378;
  assign n3380 = ~n2907 & ~n3379;
  assign n3381 = ~pi39 & ~n3380;
  assign n3382 = ~n3366 & ~n3381;
  assign n3383 = n3319 & n3382;
  assign n3384 = n3352 & ~n3383;
  assign n3385 = ~n3342 & ~n3384;
  assign n3386 = ~pi154 & ~n3385;
  assign n3387 = n3350 & ~n3386;
  assign n3388 = ~pi100 & ~n3387;
  assign n3389 = ~n3365 & n3388;
  assign n3390 = ~pi146 & ~n2522;
  assign n3391 = ~pi252 & n2522;
  assign n3392 = pi146 & ~n3391;
  assign n3393 = ~n3390 & ~n3392;
  assign n3394 = pi152 & ~n3393;
  assign n3395 = ~pi161 & ~pi166;
  assign n3396 = n3393 & ~n3395;
  assign n3397 = n3391 & n3395;
  assign n3398 = ~pi152 & ~n3397;
  assign n3399 = ~n3396 & n3398;
  assign n3400 = ~n3394 & ~n3399;
  assign n3401 = ~pi228 & n3400;
  assign n3402 = ~pi38 & ~pi216;
  assign n3403 = ~pi154 & pi299;
  assign n3404 = ~pi39 & n3317;
  assign n3405 = n3403 & n3404;
  assign n3406 = n3402 & n3405;
  assign n3407 = n3401 & n3406;
  assign n3408 = pi100 & ~n3343;
  assign n3409 = ~n3407 & n3408;
  assign n3410 = ~pi87 & ~n3409;
  assign n3411 = ~n3389 & n3410;
  assign n3412 = ~n3364 & ~n3411;
  assign n3413 = ~pi75 & ~n3412;
  assign n3414 = ~pi92 & ~n3413;
  assign n3415 = ~n3361 & n3414;
  assign n3416 = n2534 & ~n3415;
  assign n3417 = ~n3360 & n3416;
  assign n3418 = ~pi55 & ~n3417;
  assign n3419 = ~n3344 & n3418;
  assign n3420 = n2576 & n3321;
  assign n3421 = ~n3313 & ~n3420;
  assign n3422 = pi55 & n3421;
  assign n3423 = ~pi56 & ~n3422;
  assign n3424 = ~n3419 & n3423;
  assign n3425 = ~pi62 & ~n3424;
  assign n3426 = ~n3330 & n3425;
  assign n3427 = n3327 & ~n3426;
  assign n3428 = ~n3326 & n3427;
  assign n3429 = n3313 & ~n3327;
  assign n3430 = ~pi239 & ~n3429;
  assign n3431 = ~n3428 & n3430;
  assign n3432 = n2441 & n2442;
  assign n3433 = n2528 & n3432;
  assign n3434 = ~n3299 & ~n3433;
  assign n3435 = n3313 & n3434;
  assign n3436 = ~n3315 & ~n3435;
  assign n3437 = n3308 & ~n3433;
  assign n3438 = pi154 & ~n3437;
  assign n3439 = n3320 & ~n3438;
  assign n3440 = ~n3435 & ~n3439;
  assign n3441 = n3322 & n3440;
  assign n3442 = ~pi56 & n3441;
  assign n3443 = ~n3436 & ~n3442;
  assign n3444 = pi62 & ~n3443;
  assign n3445 = n2442 & n2608;
  assign n3446 = ~pi299 & n3445;
  assign n3447 = pi299 & ~n3435;
  assign n3448 = ~n3342 & ~n3447;
  assign n3449 = ~n3446 & n3448;
  assign n3450 = ~n2534 & n3449;
  assign n3451 = pi92 & ~n3449;
  assign n3452 = pi299 & ~n3440;
  assign n3453 = n2615 & n3452;
  assign n3454 = n2535 & n3453;
  assign n3455 = n3451 & ~n3454;
  assign n3456 = pi75 & n3449;
  assign n3457 = ~n3449 & ~n3452;
  assign n3458 = pi39 & ~n3457;
  assign n3459 = ~pi224 & n3087;
  assign n3460 = ~n2607 & ~n3333;
  assign n3461 = ~n3459 & ~n3460;
  assign n3462 = n3338 & ~n3461;
  assign n3463 = n3341 & ~n3462;
  assign n3464 = pi105 & ~n3087;
  assign n3465 = pi228 & ~n3464;
  assign n3466 = ~pi228 & ~n3088;
  assign n3467 = ~n3465 & ~n3466;
  assign n3468 = pi154 & ~n3467;
  assign n3469 = ~pi72 & ~n3371;
  assign n3470 = ~n2739 & ~n3469;
  assign n3471 = n2461 & ~n3470;
  assign n3472 = n3377 & ~n3471;
  assign n3473 = ~pi95 & ~n3472;
  assign n3474 = n2971 & ~n3473;
  assign n3475 = ~pi228 & n3474;
  assign n3476 = n2441 & n3087;
  assign n3477 = ~n3475 & ~n3476;
  assign n3478 = ~pi154 & ~n3477;
  assign n3479 = ~n3468 & ~n3478;
  assign n3480 = n2528 & n3479;
  assign n3481 = n3308 & ~n3480;
  assign n3482 = pi299 & ~n3481;
  assign n3483 = ~pi39 & ~n3482;
  assign n3484 = ~n3463 & n3483;
  assign n3485 = ~n3458 & ~n3484;
  assign n3486 = n2614 & n3485;
  assign n3487 = pi100 & n3407;
  assign n3488 = ~n2614 & ~n3449;
  assign n3489 = ~n3487 & n3488;
  assign n3490 = ~n3486 & ~n3489;
  assign n3491 = ~pi87 & ~n3490;
  assign n3492 = ~n3449 & ~n3453;
  assign n3493 = pi87 & n3492;
  assign n3494 = ~pi75 & ~n3493;
  assign n3495 = ~n3491 & n3494;
  assign n3496 = ~pi92 & ~n3495;
  assign n3497 = ~n3456 & n3496;
  assign n3498 = n2534 & ~n3497;
  assign n3499 = ~n3455 & n3498;
  assign n3500 = ~pi55 & ~n3499;
  assign n3501 = ~n3450 & n3500;
  assign n3502 = n2576 & n3439;
  assign n3503 = ~n3435 & ~n3502;
  assign n3504 = pi55 & n3503;
  assign n3505 = ~pi56 & ~n3504;
  assign n3506 = ~n3501 & n3505;
  assign n3507 = ~n2539 & ~n3435;
  assign n3508 = ~n3441 & ~n3507;
  assign n3509 = pi56 & n3508;
  assign n3510 = ~pi62 & ~n3509;
  assign n3511 = ~n3506 & n3510;
  assign n3512 = n3327 & ~n3511;
  assign n3513 = ~n3444 & n3512;
  assign n3514 = ~n3327 & n3435;
  assign n3515 = pi239 & ~n3514;
  assign n3516 = ~n3513 & n3515;
  assign po154 = n3431 | n3516;
  assign n3518 = pi215 & pi1145;
  assign n3519 = pi216 & pi274;
  assign n3520 = ~pi221 & ~n3519;
  assign n3521 = ~pi151 & ~n2441;
  assign n3522 = ~pi216 & ~n3521;
  assign n3523 = n3520 & ~n3522;
  assign n3524 = ~pi927 & n2452;
  assign n3525 = ~pi1145 & ~n2452;
  assign n3526 = pi221 & ~n3525;
  assign n3527 = ~n3524 & n3526;
  assign n3528 = ~n3523 & ~n3527;
  assign n3529 = ~pi215 & ~n3528;
  assign n3530 = ~n3518 & ~n3529;
  assign n3531 = ~pi215 & ~pi221;
  assign n3532 = n3432 & n3531;
  assign n3533 = ~n3519 & n3532;
  assign n3534 = n3530 & ~n3533;
  assign n3535 = ~n3315 & n3534;
  assign n3536 = ~n3432 & ~n3521;
  assign n3537 = ~pi228 & n2522;
  assign n3538 = ~pi151 & n3537;
  assign n3539 = ~n3536 & ~n3538;
  assign n3540 = ~pi216 & ~n3539;
  assign n3541 = n3520 & ~n3540;
  assign n3542 = ~n3527 & ~n3541;
  assign n3543 = ~pi215 & ~n3542;
  assign n3544 = ~n3518 & ~n3543;
  assign n3545 = n3315 & n3544;
  assign n3546 = ~n3535 & ~n3545;
  assign n3547 = pi62 & n3546;
  assign n3548 = pi235 & ~n3547;
  assign n3549 = pi223 & pi1145;
  assign n3550 = ~pi927 & n2595;
  assign n3551 = ~pi1145 & ~n2595;
  assign n3552 = pi222 & ~n3551;
  assign n3553 = ~n3550 & n3552;
  assign n3554 = pi224 & pi274;
  assign n3555 = n3332 & ~n3554;
  assign n3556 = ~n3553 & ~n3555;
  assign n3557 = ~pi223 & ~n3556;
  assign n3558 = ~n3549 & ~n3557;
  assign n3559 = ~pi299 & ~n3558;
  assign n3560 = ~n3446 & ~n3559;
  assign n3561 = pi299 & ~n3534;
  assign n3562 = n3560 & ~n3561;
  assign n3563 = ~n2534 & n3562;
  assign n3564 = ~n2615 & n3562;
  assign n3565 = pi299 & ~n3544;
  assign n3566 = n3560 & ~n3565;
  assign n3567 = n2615 & n3566;
  assign n3568 = ~n3564 & ~n3567;
  assign n3569 = n2535 & ~n3568;
  assign n3570 = pi92 & ~n3569;
  assign n3571 = ~n2535 & n3562;
  assign n3572 = n3570 & ~n3571;
  assign n3573 = pi75 & n3562;
  assign n3574 = pi87 & n3568;
  assign n3575 = pi39 & ~n3566;
  assign n3576 = ~pi222 & ~n3554;
  assign n3577 = ~n3459 & n3576;
  assign n3578 = ~n3553 & ~n3577;
  assign n3579 = ~pi223 & ~n3578;
  assign n3580 = ~pi299 & ~n3579;
  assign n3581 = ~n3549 & n3580;
  assign n3582 = ~pi151 & n3477;
  assign n3583 = pi151 & n3467;
  assign n3584 = ~pi216 & ~n3583;
  assign n3585 = ~n3582 & n3584;
  assign n3586 = n3520 & ~n3585;
  assign n3587 = ~n3527 & ~n3586;
  assign n3588 = ~pi215 & ~n3587;
  assign n3589 = ~n3518 & ~n3588;
  assign n3590 = pi299 & n3589;
  assign n3591 = ~pi39 & ~n3590;
  assign n3592 = ~n3581 & n3591;
  assign n3593 = ~pi38 & ~n3592;
  assign n3594 = ~n3575 & n3593;
  assign n3595 = pi38 & n3562;
  assign n3596 = ~pi100 & ~n3595;
  assign n3597 = ~n3594 & n3596;
  assign n3598 = ~n2532 & n3562;
  assign n3599 = pi100 & ~n3598;
  assign n3600 = n2441 & ~n2442;
  assign n3601 = ~n3401 & ~n3600;
  assign n3602 = ~pi151 & n3601;
  assign n3603 = n3540 & ~n3602;
  assign n3604 = n3520 & ~n3603;
  assign n3605 = ~n3527 & ~n3604;
  assign n3606 = ~pi215 & ~n3605;
  assign n3607 = ~n3518 & ~n3606;
  assign n3608 = pi299 & ~n3607;
  assign n3609 = n2532 & ~n3608;
  assign n3610 = n3560 & n3609;
  assign n3611 = n3599 & ~n3610;
  assign n3612 = ~n3597 & ~n3611;
  assign n3613 = ~pi87 & ~n3612;
  assign n3614 = ~pi75 & ~n3613;
  assign n3615 = ~n3574 & n3614;
  assign n3616 = ~pi92 & ~n3615;
  assign n3617 = ~n3573 & n3616;
  assign n3618 = n2534 & ~n3617;
  assign n3619 = ~n3572 & n3618;
  assign n3620 = ~pi55 & ~n3619;
  assign n3621 = ~n3563 & n3620;
  assign n3622 = ~n2576 & n3534;
  assign n3623 = pi55 & ~n3622;
  assign n3624 = n2576 & n3544;
  assign n3625 = n3623 & ~n3624;
  assign n3626 = ~pi56 & ~n3625;
  assign n3627 = ~n3621 & n3626;
  assign n3628 = ~n2539 & ~n3534;
  assign n3629 = pi56 & ~n3628;
  assign n3630 = n2539 & ~n3544;
  assign n3631 = n3629 & ~n3630;
  assign n3632 = ~pi62 & ~n3631;
  assign n3633 = ~n3627 & n3632;
  assign n3634 = n3548 & ~n3633;
  assign n3635 = n3327 & n3634;
  assign n3636 = n3318 & ~n3518;
  assign n3637 = ~n3527 & n3636;
  assign n3638 = n2522 & n3637;
  assign n3639 = n2539 & n3638;
  assign n3640 = ~n3530 & ~n3639;
  assign n3641 = pi56 & ~n3640;
  assign n3642 = pi299 & ~n3530;
  assign n3643 = ~n3559 & ~n3642;
  assign n3644 = ~n2534 & n3643;
  assign n3645 = ~n3345 & n3643;
  assign n3646 = ~n3638 & n3642;
  assign n3647 = n2533 & ~n3559;
  assign n3648 = ~n3646 & n3647;
  assign n3649 = n2535 & n3648;
  assign n3650 = pi92 & ~n3649;
  assign n3651 = ~n3645 & n3650;
  assign n3652 = pi75 & n3643;
  assign n3653 = ~n2615 & n3643;
  assign n3654 = ~n3648 & ~n3653;
  assign n3655 = pi87 & ~n3654;
  assign n3656 = ~pi100 & n3382;
  assign n3657 = ~pi39 & pi100;
  assign n3658 = n3400 & n3657;
  assign n3659 = ~n3656 & ~n3658;
  assign n3660 = ~pi38 & n3637;
  assign n3661 = ~n3659 & n3660;
  assign n3662 = n3642 & ~n3661;
  assign n3663 = ~pi87 & ~n3559;
  assign n3664 = ~n3662 & n3663;
  assign n3665 = ~n3655 & ~n3664;
  assign n3666 = ~pi75 & ~n3665;
  assign n3667 = ~pi92 & ~n3666;
  assign n3668 = ~n3652 & n3667;
  assign n3669 = n2534 & ~n3668;
  assign n3670 = ~n3651 & n3669;
  assign n3671 = ~pi55 & ~n3670;
  assign n3672 = ~n3644 & n3671;
  assign n3673 = n2576 & n3638;
  assign n3674 = ~n3530 & ~n3673;
  assign n3675 = pi55 & n3674;
  assign n3676 = ~pi56 & ~n3675;
  assign n3677 = ~n3672 & n3676;
  assign n3678 = ~pi62 & ~n3677;
  assign n3679 = ~n3641 & n3678;
  assign n3680 = n3327 & ~n3679;
  assign n3681 = n3315 & n3638;
  assign n3682 = ~n3530 & ~n3681;
  assign n3683 = pi62 & n3682;
  assign n3684 = ~pi235 & ~n3683;
  assign n3685 = n3680 & n3684;
  assign n3686 = pi235 & n3533;
  assign n3687 = ~n3327 & ~n3686;
  assign n3688 = n3530 & n3687;
  assign n3689 = ~n3685 & ~n3688;
  assign po155 = ~n3635 & n3689;
  assign n3691 = pi215 & pi1143;
  assign n3692 = pi216 & pi264;
  assign n3693 = ~pi221 & ~n3692;
  assign n3694 = pi284 & n2522;
  assign n3695 = ~n3390 & ~n3694;
  assign n3696 = ~pi228 & ~n3695;
  assign n3697 = pi284 & ~n2442;
  assign n3698 = pi105 & ~n3697;
  assign n3699 = ~pi105 & pi146;
  assign n3700 = pi228 & ~n3699;
  assign n3701 = ~n3698 & n3700;
  assign n3702 = ~n3696 & ~n3701;
  assign n3703 = ~pi216 & ~n3702;
  assign n3704 = n3693 & ~n3703;
  assign n3705 = ~pi944 & n2452;
  assign n3706 = ~pi1143 & ~n2452;
  assign n3707 = pi221 & ~n3706;
  assign n3708 = ~n3705 & n3707;
  assign n3709 = ~n3704 & ~n3708;
  assign n3710 = ~pi215 & ~n3709;
  assign n3711 = ~n3691 & ~n3710;
  assign n3712 = n3315 & n3711;
  assign n3713 = ~n3432 & ~n3701;
  assign n3714 = ~pi146 & ~pi228;
  assign n3715 = n3713 & ~n3714;
  assign n3716 = ~pi216 & ~n3715;
  assign n3717 = n3693 & ~n3716;
  assign n3718 = ~n3708 & ~n3717;
  assign n3719 = ~pi215 & ~n3718;
  assign n3720 = ~n3691 & ~n3719;
  assign n3721 = n3532 & ~n3692;
  assign n3722 = n3720 & ~n3721;
  assign n3723 = ~n3315 & n3722;
  assign n3724 = ~n3712 & ~n3723;
  assign n3725 = pi62 & n3724;
  assign n3726 = pi238 & ~n3725;
  assign n3727 = pi223 & pi1143;
  assign n3728 = pi224 & pi264;
  assign n3729 = ~pi222 & ~n3728;
  assign n3730 = ~pi224 & n3697;
  assign n3731 = n3729 & ~n3730;
  assign n3732 = ~pi944 & n2595;
  assign n3733 = ~pi1143 & ~n2595;
  assign n3734 = pi222 & ~n3733;
  assign n3735 = ~n3732 & n3734;
  assign n3736 = ~n3731 & ~n3735;
  assign n3737 = ~pi223 & ~n3736;
  assign n3738 = ~n3727 & ~n3737;
  assign n3739 = ~pi299 & ~n3738;
  assign n3740 = pi299 & ~n3722;
  assign n3741 = ~n3739 & ~n3740;
  assign n3742 = ~n2534 & n3741;
  assign n3743 = ~n2535 & n3741;
  assign n3744 = ~n2615 & n3741;
  assign n3745 = pi299 & ~n3711;
  assign n3746 = ~n3739 & ~n3745;
  assign n3747 = n2615 & n3746;
  assign n3748 = ~n3744 & ~n3747;
  assign n3749 = n2535 & ~n3748;
  assign n3750 = pi92 & ~n3749;
  assign n3751 = ~n3743 & n3750;
  assign n3752 = pi75 & n3741;
  assign n3753 = pi87 & n3748;
  assign n3754 = pi39 & ~n3746;
  assign n3755 = ~pi299 & ~n3727;
  assign n3756 = ~pi284 & n3087;
  assign n3757 = ~pi224 & ~n3756;
  assign n3758 = n3729 & ~n3757;
  assign n3759 = ~n3735 & ~n3758;
  assign n3760 = ~n3087 & n3729;
  assign n3761 = n3759 & ~n3760;
  assign n3762 = ~pi223 & ~n3761;
  assign n3763 = n3755 & ~n3762;
  assign n3764 = ~pi39 & ~n3763;
  assign n3765 = pi299 & ~n3691;
  assign n3766 = ~n3464 & n3701;
  assign n3767 = pi146 & ~n3474;
  assign n3768 = ~pi146 & n3088;
  assign n3769 = pi284 & ~n3768;
  assign n3770 = ~n3767 & n3769;
  assign n3771 = ~pi146 & ~pi284;
  assign n3772 = ~n3380 & n3771;
  assign n3773 = ~n3770 & ~n3772;
  assign n3774 = ~pi228 & ~n3773;
  assign n3775 = ~n3766 & ~n3774;
  assign n3776 = ~pi216 & ~n3775;
  assign n3777 = n3693 & ~n3776;
  assign n3778 = ~n3708 & ~n3777;
  assign n3779 = ~pi215 & ~n3778;
  assign n3780 = n3765 & ~n3779;
  assign n3781 = n3764 & ~n3780;
  assign n3782 = ~pi38 & ~n3781;
  assign n3783 = ~n3754 & n3782;
  assign n3784 = pi38 & n3741;
  assign n3785 = ~pi100 & ~n3784;
  assign n3786 = ~n3783 & n3785;
  assign n3787 = ~n2532 & n3741;
  assign n3788 = pi100 & ~n3787;
  assign n3789 = ~pi228 & ~n3392;
  assign n3790 = pi252 & n2627;
  assign n3791 = ~pi284 & ~n3790;
  assign n3792 = n2522 & n3791;
  assign n3793 = n3789 & ~n3792;
  assign n3794 = ~n3701 & ~n3793;
  assign n3795 = ~pi216 & ~n3794;
  assign n3796 = n3693 & ~n3795;
  assign n3797 = ~n3708 & ~n3796;
  assign n3798 = ~pi215 & ~n3797;
  assign n3799 = ~n3691 & ~n3798;
  assign n3800 = pi299 & ~n3799;
  assign n3801 = ~n3739 & ~n3800;
  assign n3802 = n2532 & n3801;
  assign n3803 = n3788 & ~n3802;
  assign n3804 = ~n3786 & ~n3803;
  assign n3805 = ~pi87 & ~n3804;
  assign n3806 = ~pi75 & ~n3805;
  assign n3807 = ~n3753 & n3806;
  assign n3808 = ~pi92 & ~n3807;
  assign n3809 = ~n3752 & n3808;
  assign n3810 = n2534 & ~n3809;
  assign n3811 = ~n3751 & n3810;
  assign n3812 = ~pi55 & ~n3811;
  assign n3813 = ~n3742 & n3812;
  assign n3814 = ~n2576 & n3722;
  assign n3815 = n2576 & n3711;
  assign n3816 = pi55 & ~n3815;
  assign n3817 = ~n3814 & n3816;
  assign n3818 = ~pi56 & ~n3817;
  assign n3819 = ~n3813 & n3818;
  assign n3820 = ~n2539 & ~n3722;
  assign n3821 = pi56 & ~n3820;
  assign n3822 = n2539 & ~n3711;
  assign n3823 = n3821 & ~n3822;
  assign n3824 = ~pi62 & ~n3823;
  assign n3825 = ~n3819 & n3824;
  assign n3826 = n3726 & ~n3825;
  assign n3827 = n3327 & n3826;
  assign n3828 = ~n3445 & n3739;
  assign n3829 = pi299 & ~n3720;
  assign n3830 = ~n3828 & ~n3829;
  assign n3831 = ~n2534 & n3830;
  assign n3832 = ~n2535 & n3830;
  assign n3833 = ~n2615 & n3830;
  assign n3834 = ~n3696 & n3713;
  assign n3835 = ~pi216 & ~n3834;
  assign n3836 = n3693 & ~n3835;
  assign n3837 = ~n3708 & ~n3836;
  assign n3838 = ~pi215 & ~n3837;
  assign n3839 = ~n3691 & ~n3838;
  assign n3840 = pi299 & ~n3839;
  assign n3841 = ~n3828 & ~n3840;
  assign n3842 = n2615 & n3841;
  assign n3843 = ~n3833 & ~n3842;
  assign n3844 = n2535 & ~n3843;
  assign n3845 = pi92 & ~n3844;
  assign n3846 = ~n3832 & n3845;
  assign n3847 = pi75 & n3830;
  assign n3848 = pi87 & n3843;
  assign n3849 = pi39 & ~n3841;
  assign n3850 = n3755 & n3759;
  assign n3851 = ~pi146 & ~n3474;
  assign n3852 = pi146 & n3088;
  assign n3853 = ~pi284 & ~n3852;
  assign n3854 = ~n3851 & n3853;
  assign n3855 = pi146 & pi284;
  assign n3856 = ~n3380 & n3855;
  assign n3857 = ~pi228 & ~n3856;
  assign n3858 = ~n3854 & n3857;
  assign n3859 = n2441 & ~n3087;
  assign n3860 = ~n3701 & ~n3859;
  assign n3861 = ~n3858 & n3860;
  assign n3862 = ~pi216 & ~n3861;
  assign n3863 = n3693 & ~n3862;
  assign n3864 = ~n3708 & ~n3863;
  assign n3865 = ~pi215 & ~n3864;
  assign n3866 = n3765 & ~n3865;
  assign n3867 = ~n3850 & ~n3866;
  assign n3868 = n3764 & n3867;
  assign n3869 = ~pi38 & ~n3868;
  assign n3870 = ~n3849 & n3869;
  assign n3871 = pi38 & n3830;
  assign n3872 = ~pi100 & ~n3871;
  assign n3873 = ~n3870 & n3872;
  assign n3874 = ~n2532 & n3830;
  assign n3875 = pi100 & ~n3874;
  assign n3876 = n3713 & ~n3793;
  assign n3877 = ~pi216 & ~n3876;
  assign n3878 = n3693 & ~n3877;
  assign n3879 = ~n3708 & ~n3878;
  assign n3880 = ~pi215 & ~n3879;
  assign n3881 = ~n3691 & ~n3880;
  assign n3882 = pi299 & ~n3881;
  assign n3883 = ~n3828 & ~n3882;
  assign n3884 = n2532 & n3883;
  assign n3885 = n3875 & ~n3884;
  assign n3886 = ~n3873 & ~n3885;
  assign n3887 = ~pi87 & ~n3886;
  assign n3888 = ~pi75 & ~n3887;
  assign n3889 = ~n3848 & n3888;
  assign n3890 = ~pi92 & ~n3889;
  assign n3891 = ~n3847 & n3890;
  assign n3892 = n2534 & ~n3891;
  assign n3893 = ~n3846 & n3892;
  assign n3894 = ~pi55 & ~n3893;
  assign n3895 = ~n3831 & n3894;
  assign n3896 = ~n2576 & n3720;
  assign n3897 = pi55 & ~n3896;
  assign n3898 = n2576 & n3839;
  assign n3899 = n3897 & ~n3898;
  assign n3900 = ~pi56 & ~n3899;
  assign n3901 = ~n3895 & n3900;
  assign n3902 = ~n2539 & ~n3720;
  assign n3903 = pi56 & ~n3902;
  assign n3904 = n2539 & ~n3839;
  assign n3905 = n3903 & ~n3904;
  assign n3906 = ~pi62 & ~n3905;
  assign n3907 = ~n3901 & n3906;
  assign n3908 = n3327 & ~n3907;
  assign n3909 = ~n3315 & n3720;
  assign n3910 = n3315 & n3839;
  assign n3911 = ~n3909 & ~n3910;
  assign n3912 = pi62 & n3911;
  assign n3913 = ~pi238 & ~n3912;
  assign n3914 = n3908 & n3913;
  assign n3915 = pi238 & n3721;
  assign n3916 = ~n3327 & ~n3915;
  assign n3917 = n3720 & n3916;
  assign n3918 = ~n3914 & ~n3917;
  assign po156 = ~n3827 & n3918;
  assign n3920 = pi215 & pi1142;
  assign n3921 = pi216 & pi277;
  assign n3922 = ~pi221 & ~n3921;
  assign n3923 = pi172 & ~pi228;
  assign n3924 = pi262 & ~n2442;
  assign n3925 = pi105 & n3924;
  assign n3926 = ~pi105 & pi172;
  assign n3927 = ~n3925 & ~n3926;
  assign n3928 = pi228 & ~n3927;
  assign n3929 = ~n3923 & ~n3928;
  assign n3930 = ~pi216 & ~n3929;
  assign n3931 = n3922 & ~n3930;
  assign n3932 = ~pi932 & n2452;
  assign n3933 = ~pi1142 & ~n2452;
  assign n3934 = pi221 & ~n3933;
  assign n3935 = ~n3932 & n3934;
  assign n3936 = ~n3931 & ~n3935;
  assign n3937 = ~pi215 & ~n3936;
  assign n3938 = ~n3920 & ~n3937;
  assign n3939 = ~n3433 & ~n3938;
  assign n3940 = ~n3315 & ~n3939;
  assign n3941 = pi62 & ~n3940;
  assign n3942 = ~pi262 & n2522;
  assign n3943 = ~n3537 & ~n3923;
  assign n3944 = ~n3942 & ~n3943;
  assign n3945 = ~n3432 & ~n3928;
  assign n3946 = ~n3944 & n3945;
  assign n3947 = ~pi216 & ~n3946;
  assign n3948 = n3922 & ~n3947;
  assign n3949 = ~n3935 & ~n3948;
  assign n3950 = ~pi215 & ~n3949;
  assign n3951 = ~n3920 & ~n3950;
  assign n3952 = n3315 & n3951;
  assign n3953 = n3941 & ~n3952;
  assign n3954 = pi223 & pi1142;
  assign n3955 = pi224 & pi277;
  assign n3956 = ~pi222 & ~n3955;
  assign n3957 = ~pi224 & n3924;
  assign n3958 = n3956 & ~n3957;
  assign n3959 = ~pi932 & n2595;
  assign n3960 = ~pi1142 & ~n2595;
  assign n3961 = pi222 & ~n3960;
  assign n3962 = ~n3959 & n3961;
  assign n3963 = ~n3958 & ~n3962;
  assign n3964 = ~pi223 & ~n3963;
  assign n3965 = ~n3954 & ~n3964;
  assign n3966 = ~pi299 & ~n3965;
  assign n3967 = ~n3445 & n3966;
  assign n3968 = pi299 & n3939;
  assign n3969 = ~n3967 & ~n3968;
  assign n3970 = ~n2534 & n3969;
  assign n3971 = ~n2535 & n3969;
  assign n3972 = ~n2615 & n3969;
  assign n3973 = pi299 & ~n3951;
  assign n3974 = ~n3967 & ~n3973;
  assign n3975 = n2615 & n3974;
  assign n3976 = ~n3972 & ~n3975;
  assign n3977 = n2535 & ~n3976;
  assign n3978 = pi92 & ~n3977;
  assign n3979 = ~n3971 & n3978;
  assign n3980 = pi75 & n3969;
  assign n3981 = pi87 & n3976;
  assign n3982 = pi39 & ~n3974;
  assign n3983 = ~pi299 & ~n3954;
  assign n3984 = ~pi262 & n3087;
  assign n3985 = ~pi224 & ~n3984;
  assign n3986 = n3956 & ~n3985;
  assign n3987 = ~n3962 & ~n3986;
  assign n3988 = ~n3087 & n3956;
  assign n3989 = n3987 & ~n3988;
  assign n3990 = ~pi223 & ~n3989;
  assign n3991 = n3983 & ~n3990;
  assign n3992 = ~pi39 & ~n3991;
  assign n3993 = n3983 & n3987;
  assign n3994 = pi299 & ~n3920;
  assign n3995 = ~pi262 & n3088;
  assign n3996 = ~pi172 & ~n3995;
  assign n3997 = pi172 & ~pi262;
  assign n3998 = n3474 & n3997;
  assign n3999 = ~n3996 & ~n3998;
  assign n4000 = pi262 & n3380;
  assign n4001 = ~pi228 & ~n4000;
  assign n4002 = ~n3999 & n4001;
  assign n4003 = ~n3086 & n3925;
  assign n4004 = pi228 & ~n3926;
  assign n4005 = ~n4003 & n4004;
  assign n4006 = ~n3464 & n4005;
  assign n4007 = ~pi216 & ~n4006;
  assign n4008 = ~n4002 & n4007;
  assign n4009 = n3922 & ~n4008;
  assign n4010 = ~n3935 & ~n4009;
  assign n4011 = ~pi215 & ~n4010;
  assign n4012 = n3994 & ~n4011;
  assign n4013 = ~n3993 & ~n4012;
  assign n4014 = n3992 & n4013;
  assign n4015 = ~pi38 & ~n4014;
  assign n4016 = ~n3982 & n4015;
  assign n4017 = pi38 & n3969;
  assign n4018 = ~pi100 & ~n4017;
  assign n4019 = ~n4016 & n4018;
  assign n4020 = ~n2532 & n3969;
  assign n4021 = pi100 & ~n4020;
  assign n4022 = ~pi262 & n3400;
  assign n4023 = ~n3401 & ~n3923;
  assign n4024 = ~n4022 & ~n4023;
  assign n4025 = n3945 & ~n4024;
  assign n4026 = ~pi216 & ~n4025;
  assign n4027 = n3922 & ~n4026;
  assign n4028 = ~n3935 & ~n4027;
  assign n4029 = ~pi215 & ~n4028;
  assign n4030 = ~n3920 & ~n4029;
  assign n4031 = pi299 & ~n4030;
  assign n4032 = ~n3967 & ~n4031;
  assign n4033 = n2532 & n4032;
  assign n4034 = n4021 & ~n4033;
  assign n4035 = ~n4019 & ~n4034;
  assign n4036 = ~pi87 & ~n4035;
  assign n4037 = ~pi75 & ~n4036;
  assign n4038 = ~n3981 & n4037;
  assign n4039 = ~pi92 & ~n4038;
  assign n4040 = ~n3980 & n4039;
  assign n4041 = n2534 & ~n4040;
  assign n4042 = ~n3979 & n4041;
  assign n4043 = ~pi55 & ~n4042;
  assign n4044 = ~n3970 & n4043;
  assign n4045 = ~n2576 & ~n3939;
  assign n4046 = pi55 & ~n4045;
  assign n4047 = n2576 & n3951;
  assign n4048 = n4046 & ~n4047;
  assign n4049 = ~pi56 & ~n4048;
  assign n4050 = ~n4044 & n4049;
  assign n4051 = ~n2539 & n3939;
  assign n4052 = n2539 & ~n3951;
  assign n4053 = pi56 & ~n4052;
  assign n4054 = ~n4051 & n4053;
  assign n4055 = ~pi62 & ~n4054;
  assign n4056 = ~n4050 & n4055;
  assign n4057 = n3327 & ~n4056;
  assign n4058 = ~n3953 & n4057;
  assign n4059 = ~n3327 & ~n3939;
  assign n4060 = ~pi249 & ~n4059;
  assign n4061 = ~n4058 & n4060;
  assign n4062 = ~n3315 & n3938;
  assign n4063 = pi62 & ~n4062;
  assign n4064 = ~n3928 & ~n3944;
  assign n4065 = ~pi216 & ~n4064;
  assign n4066 = n3922 & ~n4065;
  assign n4067 = ~n3935 & ~n4066;
  assign n4068 = ~pi215 & ~n4067;
  assign n4069 = ~n3920 & ~n4068;
  assign n4070 = n3315 & n4069;
  assign n4071 = n4063 & ~n4070;
  assign n4072 = pi299 & ~n3938;
  assign n4073 = ~n3966 & ~n4072;
  assign n4074 = ~n2534 & n4073;
  assign n4075 = ~n2535 & n4073;
  assign n4076 = ~n2615 & n4073;
  assign n4077 = pi299 & ~n4069;
  assign n4078 = ~n3966 & ~n4077;
  assign n4079 = n2615 & n4078;
  assign n4080 = ~n4076 & ~n4079;
  assign n4081 = n2535 & ~n4080;
  assign n4082 = pi92 & ~n4081;
  assign n4083 = ~n4075 & n4082;
  assign n4084 = pi75 & n4073;
  assign n4085 = pi87 & n4080;
  assign n4086 = pi39 & ~n4078;
  assign n4087 = pi262 & n3474;
  assign n4088 = ~pi172 & ~n4087;
  assign n4089 = ~pi262 & ~n3380;
  assign n4090 = pi262 & ~n3088;
  assign n4091 = pi172 & ~n4090;
  assign n4092 = ~n4089 & n4091;
  assign n4093 = ~n4088 & ~n4092;
  assign n4094 = ~pi228 & ~n4093;
  assign n4095 = ~pi216 & ~n4005;
  assign n4096 = ~n4094 & n4095;
  assign n4097 = n3922 & ~n4096;
  assign n4098 = ~n3935 & ~n4097;
  assign n4099 = ~pi215 & ~n4098;
  assign n4100 = n3994 & ~n4099;
  assign n4101 = n3992 & ~n4100;
  assign n4102 = ~pi38 & ~n4101;
  assign n4103 = ~n4086 & n4102;
  assign n4104 = pi38 & n4073;
  assign n4105 = ~pi100 & ~n4104;
  assign n4106 = ~n4103 & n4105;
  assign n4107 = ~n2532 & n4073;
  assign n4108 = pi100 & ~n4107;
  assign n4109 = ~n3928 & ~n4024;
  assign n4110 = ~pi216 & ~n4109;
  assign n4111 = n3922 & ~n4110;
  assign n4112 = ~n3935 & ~n4111;
  assign n4113 = ~pi215 & ~n4112;
  assign n4114 = ~n3920 & ~n4113;
  assign n4115 = pi299 & ~n4114;
  assign n4116 = ~n3966 & ~n4115;
  assign n4117 = n2532 & n4116;
  assign n4118 = n4108 & ~n4117;
  assign n4119 = ~n4106 & ~n4118;
  assign n4120 = ~pi87 & ~n4119;
  assign n4121 = ~pi75 & ~n4120;
  assign n4122 = ~n4085 & n4121;
  assign n4123 = ~pi92 & ~n4122;
  assign n4124 = ~n4084 & n4123;
  assign n4125 = n2534 & ~n4124;
  assign n4126 = ~n4083 & n4125;
  assign n4127 = ~pi55 & ~n4126;
  assign n4128 = ~n4074 & n4127;
  assign n4129 = ~n2576 & n3938;
  assign n4130 = pi55 & ~n4129;
  assign n4131 = n2576 & n4069;
  assign n4132 = n4130 & ~n4131;
  assign n4133 = ~pi56 & ~n4132;
  assign n4134 = ~n4128 & n4133;
  assign n4135 = ~n2539 & ~n3938;
  assign n4136 = pi56 & ~n4135;
  assign n4137 = n2539 & ~n4069;
  assign n4138 = n4136 & ~n4137;
  assign n4139 = ~pi62 & ~n4138;
  assign n4140 = ~n4134 & n4139;
  assign n4141 = n3327 & ~n4140;
  assign n4142 = ~n4071 & n4141;
  assign n4143 = ~n3327 & n3938;
  assign n4144 = pi249 & ~n4143;
  assign n4145 = ~n4142 & n4144;
  assign po157 = n4061 | n4145;
  assign n4147 = pi223 & pi1141;
  assign n4148 = pi224 & pi270;
  assign n4149 = ~pi222 & ~n4148;
  assign n4150 = pi861 & ~n2442;
  assign n4151 = ~pi224 & ~n4150;
  assign n4152 = n4149 & ~n4151;
  assign n4153 = ~pi935 & n2595;
  assign n4154 = ~pi1141 & ~n2595;
  assign n4155 = pi222 & ~n4154;
  assign n4156 = ~n4153 & n4155;
  assign n4157 = ~n4152 & ~n4156;
  assign n4158 = ~pi223 & ~n4157;
  assign n4159 = ~n4147 & ~n4158;
  assign n4160 = ~pi299 & ~n4159;
  assign n4161 = pi215 & pi1141;
  assign n4162 = pi216 & pi270;
  assign n4163 = ~pi221 & ~n4162;
  assign n4164 = pi105 & ~n4150;
  assign n4165 = ~pi105 & pi171;
  assign n4166 = pi228 & ~n4165;
  assign n4167 = ~n4164 & n4166;
  assign n4168 = ~pi216 & ~n4167;
  assign n4169 = ~pi171 & ~pi228;
  assign n4170 = n4168 & ~n4169;
  assign n4171 = n4163 & ~n4170;
  assign n4172 = ~pi935 & n2452;
  assign n4173 = ~pi1141 & ~n2452;
  assign n4174 = pi221 & ~n4173;
  assign n4175 = ~n4172 & n4174;
  assign n4176 = ~n4171 & ~n4175;
  assign n4177 = ~pi215 & ~n4176;
  assign n4178 = ~n4161 & ~n4177;
  assign n4179 = pi299 & ~n4178;
  assign n4180 = ~n4160 & ~n4179;
  assign n4181 = ~n2534 & n4180;
  assign n4182 = ~n2535 & n4180;
  assign n4183 = ~n2615 & n4180;
  assign n4184 = pi171 & ~n2522;
  assign n4185 = ~pi861 & n2522;
  assign n4186 = ~pi228 & ~n4185;
  assign n4187 = ~n4184 & n4186;
  assign n4188 = n4168 & ~n4187;
  assign n4189 = n4163 & ~n4188;
  assign n4190 = ~n4175 & ~n4189;
  assign n4191 = ~pi215 & ~n4190;
  assign n4192 = ~n4161 & ~n4191;
  assign n4193 = pi299 & ~n4192;
  assign n4194 = ~n4160 & ~n4193;
  assign n4195 = n2615 & n4194;
  assign n4196 = ~n4183 & ~n4195;
  assign n4197 = n2535 & ~n4196;
  assign n4198 = pi92 & ~n4197;
  assign n4199 = ~n4182 & n4198;
  assign n4200 = pi75 & n4180;
  assign n4201 = pi87 & n4196;
  assign n4202 = pi39 & ~n4194;
  assign n4203 = ~pi299 & ~n4147;
  assign n4204 = pi861 & n3087;
  assign n4205 = ~pi224 & ~n4204;
  assign n4206 = n4149 & ~n4205;
  assign n4207 = ~n4156 & ~n4206;
  assign n4208 = ~n3087 & n4149;
  assign n4209 = n4207 & ~n4208;
  assign n4210 = ~pi223 & ~n4209;
  assign n4211 = n4203 & ~n4210;
  assign n4212 = ~pi39 & ~n4211;
  assign n4213 = n4203 & n4207;
  assign n4214 = pi299 & ~n4161;
  assign n4215 = pi861 & n3088;
  assign n4216 = ~pi861 & n3380;
  assign n4217 = ~pi171 & ~n4216;
  assign n4218 = ~n4215 & n4217;
  assign n4219 = pi171 & n3474;
  assign n4220 = pi861 & n4219;
  assign n4221 = ~n4218 & ~n4220;
  assign n4222 = ~pi228 & ~n4221;
  assign n4223 = ~n3464 & n4167;
  assign n4224 = ~pi216 & ~n4223;
  assign n4225 = ~n4222 & n4224;
  assign n4226 = n4163 & ~n4225;
  assign n4227 = ~n4175 & ~n4226;
  assign n4228 = ~pi215 & ~n4227;
  assign n4229 = n4214 & ~n4228;
  assign n4230 = ~n4213 & ~n4229;
  assign n4231 = n4212 & n4230;
  assign n4232 = ~pi38 & ~n4231;
  assign n4233 = ~n4202 & n4232;
  assign n4234 = pi38 & n4180;
  assign n4235 = ~pi100 & ~n4234;
  assign n4236 = ~n4233 & n4235;
  assign n4237 = ~n2532 & n4180;
  assign n4238 = pi100 & ~n4237;
  assign n4239 = ~pi861 & n3400;
  assign n4240 = ~n3401 & ~n4169;
  assign n4241 = ~n4239 & ~n4240;
  assign n4242 = n4168 & ~n4241;
  assign n4243 = n4163 & ~n4242;
  assign n4244 = ~n4175 & ~n4243;
  assign n4245 = ~pi215 & ~n4244;
  assign n4246 = ~n4161 & ~n4245;
  assign n4247 = pi299 & ~n4246;
  assign n4248 = ~n4160 & ~n4247;
  assign n4249 = n2532 & n4248;
  assign n4250 = n4238 & ~n4249;
  assign n4251 = ~n4236 & ~n4250;
  assign n4252 = ~pi87 & ~n4251;
  assign n4253 = ~pi75 & ~n4252;
  assign n4254 = ~n4201 & n4253;
  assign n4255 = ~pi92 & ~n4254;
  assign n4256 = ~n4200 & n4255;
  assign n4257 = n2534 & ~n4256;
  assign n4258 = ~n4199 & n4257;
  assign n4259 = ~pi55 & ~n4258;
  assign n4260 = ~n4181 & n4259;
  assign n4261 = ~n2576 & n4178;
  assign n4262 = pi55 & ~n4261;
  assign n4263 = n2576 & n4192;
  assign n4264 = n4262 & ~n4263;
  assign n4265 = ~pi56 & ~n4264;
  assign n4266 = ~n4260 & n4265;
  assign n4267 = ~n2539 & ~n4178;
  assign n4268 = pi56 & ~n4267;
  assign n4269 = n2539 & ~n4192;
  assign n4270 = n4268 & ~n4269;
  assign n4271 = ~pi62 & ~n4270;
  assign n4272 = ~n4266 & n4271;
  assign n4273 = n3327 & ~n4272;
  assign n4274 = ~n3315 & n4178;
  assign n4275 = n3315 & n4192;
  assign n4276 = ~n4274 & ~n4275;
  assign n4277 = pi62 & n4276;
  assign n4278 = ~pi241 & ~n4277;
  assign n4279 = n4273 & n4278;
  assign n4280 = ~n3432 & n4168;
  assign n4281 = ~n4187 & n4280;
  assign n4282 = n4163 & ~n4281;
  assign n4283 = ~n4175 & ~n4282;
  assign n4284 = ~pi215 & ~n4283;
  assign n4285 = ~n4161 & ~n4284;
  assign n4286 = n3315 & n4285;
  assign n4287 = n3532 & ~n4162;
  assign n4288 = n4178 & ~n4287;
  assign n4289 = ~n3315 & n4288;
  assign n4290 = ~n4286 & ~n4289;
  assign n4291 = pi62 & n4290;
  assign n4292 = pi241 & ~n4291;
  assign n4293 = ~n3446 & ~n4160;
  assign n4294 = pi299 & ~n4288;
  assign n4295 = n4293 & ~n4294;
  assign n4296 = ~n2534 & n4295;
  assign n4297 = ~n2615 & n4295;
  assign n4298 = pi299 & ~n4285;
  assign n4299 = n4293 & ~n4298;
  assign n4300 = n2615 & n4299;
  assign n4301 = ~n4297 & ~n4300;
  assign n4302 = n2535 & ~n4301;
  assign n4303 = pi92 & ~n4302;
  assign n4304 = ~n2535 & n4295;
  assign n4305 = n4303 & ~n4304;
  assign n4306 = pi75 & n4295;
  assign n4307 = pi87 & n4301;
  assign n4308 = pi39 & ~n4299;
  assign n4309 = ~pi861 & n3474;
  assign n4310 = ~pi171 & ~n4309;
  assign n4311 = pi861 & ~n3380;
  assign n4312 = ~pi861 & ~n3088;
  assign n4313 = pi171 & ~n4312;
  assign n4314 = ~n4311 & n4313;
  assign n4315 = ~n4310 & ~n4314;
  assign n4316 = ~pi228 & n4315;
  assign n4317 = ~n3465 & ~n4316;
  assign n4318 = n4168 & ~n4317;
  assign n4319 = n4163 & ~n4318;
  assign n4320 = ~n4175 & ~n4319;
  assign n4321 = ~pi215 & ~n4320;
  assign n4322 = n4214 & ~n4321;
  assign n4323 = n4212 & ~n4322;
  assign n4324 = ~pi38 & ~n4323;
  assign n4325 = ~n4308 & n4324;
  assign n4326 = pi38 & n4295;
  assign n4327 = ~pi100 & ~n4326;
  assign n4328 = ~n4325 & n4327;
  assign n4329 = ~n2532 & n4295;
  assign n4330 = pi100 & ~n4329;
  assign n4331 = ~n4241 & n4280;
  assign n4332 = n4163 & ~n4331;
  assign n4333 = ~n4175 & ~n4332;
  assign n4334 = ~pi215 & ~n4333;
  assign n4335 = ~n4161 & ~n4334;
  assign n4336 = pi299 & ~n4335;
  assign n4337 = n2532 & ~n4336;
  assign n4338 = n4293 & n4337;
  assign n4339 = n4330 & ~n4338;
  assign n4340 = ~n4328 & ~n4339;
  assign n4341 = ~pi87 & ~n4340;
  assign n4342 = ~pi75 & ~n4341;
  assign n4343 = ~n4307 & n4342;
  assign n4344 = ~pi92 & ~n4343;
  assign n4345 = ~n4306 & n4344;
  assign n4346 = n2534 & ~n4345;
  assign n4347 = ~n4305 & n4346;
  assign n4348 = ~pi55 & ~n4347;
  assign n4349 = ~n4296 & n4348;
  assign n4350 = ~n2576 & n4288;
  assign n4351 = n2576 & n4285;
  assign n4352 = pi55 & ~n4351;
  assign n4353 = ~n4350 & n4352;
  assign n4354 = ~pi56 & ~n4353;
  assign n4355 = ~n4349 & n4354;
  assign n4356 = ~n2539 & ~n4288;
  assign n4357 = pi56 & ~n4356;
  assign n4358 = n2539 & ~n4285;
  assign n4359 = n4357 & ~n4358;
  assign n4360 = ~pi62 & ~n4359;
  assign n4361 = ~n4355 & n4360;
  assign n4362 = n4292 & ~n4361;
  assign n4363 = n3327 & n4362;
  assign n4364 = pi241 & n4287;
  assign n4365 = ~n3327 & ~n4364;
  assign n4366 = n4178 & n4365;
  assign n4367 = ~n4363 & ~n4366;
  assign po158 = ~n4279 & n4367;
  assign n4369 = pi223 & pi1140;
  assign n4370 = pi224 & pi282;
  assign n4371 = ~pi222 & ~n4370;
  assign n4372 = pi869 & ~n2442;
  assign n4373 = ~pi224 & ~n4372;
  assign n4374 = n4371 & ~n4373;
  assign n4375 = ~pi921 & n2595;
  assign n4376 = ~pi1140 & ~n2595;
  assign n4377 = pi222 & ~n4376;
  assign n4378 = ~n4375 & n4377;
  assign n4379 = ~n4374 & ~n4378;
  assign n4380 = ~pi223 & ~n4379;
  assign n4381 = ~n4369 & ~n4380;
  assign n4382 = ~pi299 & ~n4381;
  assign n4383 = pi215 & pi1140;
  assign n4384 = pi216 & pi282;
  assign n4385 = ~pi221 & ~n4384;
  assign n4386 = pi105 & ~n4372;
  assign n4387 = ~pi105 & pi170;
  assign n4388 = pi228 & ~n4387;
  assign n4389 = ~n4386 & n4388;
  assign n4390 = ~pi216 & ~n4389;
  assign n4391 = ~pi170 & ~pi228;
  assign n4392 = n4390 & ~n4391;
  assign n4393 = n4385 & ~n4392;
  assign n4394 = ~pi921 & n2452;
  assign n4395 = ~pi1140 & ~n2452;
  assign n4396 = pi221 & ~n4395;
  assign n4397 = ~n4394 & n4396;
  assign n4398 = ~n4393 & ~n4397;
  assign n4399 = ~pi215 & ~n4398;
  assign n4400 = ~n4383 & ~n4399;
  assign n4401 = pi299 & ~n4400;
  assign n4402 = ~n4382 & ~n4401;
  assign n4403 = ~n2534 & n4402;
  assign n4404 = ~n2535 & n4402;
  assign n4405 = ~n2615 & n4402;
  assign n4406 = pi170 & ~n2522;
  assign n4407 = ~pi869 & n2522;
  assign n4408 = ~pi228 & ~n4407;
  assign n4409 = ~n4406 & n4408;
  assign n4410 = n4390 & ~n4409;
  assign n4411 = n4385 & ~n4410;
  assign n4412 = ~n4397 & ~n4411;
  assign n4413 = ~pi215 & ~n4412;
  assign n4414 = ~n4383 & ~n4413;
  assign n4415 = pi299 & ~n4414;
  assign n4416 = ~n4382 & ~n4415;
  assign n4417 = n2615 & n4416;
  assign n4418 = ~n4405 & ~n4417;
  assign n4419 = n2535 & ~n4418;
  assign n4420 = pi92 & ~n4419;
  assign n4421 = ~n4404 & n4420;
  assign n4422 = pi75 & n4402;
  assign n4423 = pi87 & n4418;
  assign n4424 = pi39 & ~n4416;
  assign n4425 = ~pi299 & ~n4369;
  assign n4426 = pi869 & n3087;
  assign n4427 = ~pi224 & ~n4426;
  assign n4428 = n4371 & ~n4427;
  assign n4429 = ~n4378 & ~n4428;
  assign n4430 = ~n3087 & n4371;
  assign n4431 = n4429 & ~n4430;
  assign n4432 = ~pi223 & ~n4431;
  assign n4433 = n4425 & ~n4432;
  assign n4434 = ~pi39 & ~n4433;
  assign n4435 = n4425 & n4429;
  assign n4436 = pi299 & ~n4383;
  assign n4437 = pi869 & n3088;
  assign n4438 = ~pi869 & n3380;
  assign n4439 = ~pi170 & ~n4438;
  assign n4440 = ~n4437 & n4439;
  assign n4441 = pi170 & n3474;
  assign n4442 = pi869 & n4441;
  assign n4443 = ~n4440 & ~n4442;
  assign n4444 = ~pi228 & ~n4443;
  assign n4445 = ~n3464 & n4389;
  assign n4446 = ~pi216 & ~n4445;
  assign n4447 = ~n4444 & n4446;
  assign n4448 = n4385 & ~n4447;
  assign n4449 = ~n4397 & ~n4448;
  assign n4450 = ~pi215 & ~n4449;
  assign n4451 = n4436 & ~n4450;
  assign n4452 = ~n4435 & ~n4451;
  assign n4453 = n4434 & n4452;
  assign n4454 = ~pi38 & ~n4453;
  assign n4455 = ~n4424 & n4454;
  assign n4456 = pi38 & n4402;
  assign n4457 = ~pi100 & ~n4456;
  assign n4458 = ~n4455 & n4457;
  assign n4459 = ~n2532 & n4402;
  assign n4460 = pi100 & ~n4459;
  assign n4461 = ~pi869 & n3400;
  assign n4462 = ~n3401 & ~n4391;
  assign n4463 = ~n4461 & ~n4462;
  assign n4464 = n4390 & ~n4463;
  assign n4465 = n4385 & ~n4464;
  assign n4466 = ~n4397 & ~n4465;
  assign n4467 = ~pi215 & ~n4466;
  assign n4468 = ~n4383 & ~n4467;
  assign n4469 = pi299 & ~n4468;
  assign n4470 = ~n4382 & ~n4469;
  assign n4471 = n2532 & n4470;
  assign n4472 = n4460 & ~n4471;
  assign n4473 = ~n4458 & ~n4472;
  assign n4474 = ~pi87 & ~n4473;
  assign n4475 = ~pi75 & ~n4474;
  assign n4476 = ~n4423 & n4475;
  assign n4477 = ~pi92 & ~n4476;
  assign n4478 = ~n4422 & n4477;
  assign n4479 = n2534 & ~n4478;
  assign n4480 = ~n4421 & n4479;
  assign n4481 = ~pi55 & ~n4480;
  assign n4482 = ~n4403 & n4481;
  assign n4483 = ~n2576 & n4400;
  assign n4484 = pi55 & ~n4483;
  assign n4485 = n2576 & n4414;
  assign n4486 = n4484 & ~n4485;
  assign n4487 = ~pi56 & ~n4486;
  assign n4488 = ~n4482 & n4487;
  assign n4489 = ~n2539 & ~n4400;
  assign n4490 = pi56 & ~n4489;
  assign n4491 = n2539 & ~n4414;
  assign n4492 = n4490 & ~n4491;
  assign n4493 = ~pi62 & ~n4492;
  assign n4494 = ~n4488 & n4493;
  assign n4495 = n3327 & ~n4494;
  assign n4496 = ~n3315 & n4400;
  assign n4497 = n3315 & n4414;
  assign n4498 = ~n4496 & ~n4497;
  assign n4499 = pi62 & n4498;
  assign n4500 = ~pi248 & ~n4499;
  assign n4501 = n4495 & n4500;
  assign n4502 = ~n3432 & n4390;
  assign n4503 = ~n4409 & n4502;
  assign n4504 = n4385 & ~n4503;
  assign n4505 = ~n4397 & ~n4504;
  assign n4506 = ~pi215 & ~n4505;
  assign n4507 = ~n4383 & ~n4506;
  assign n4508 = n3315 & n4507;
  assign n4509 = n3532 & ~n4384;
  assign n4510 = n4400 & ~n4509;
  assign n4511 = ~n3315 & n4510;
  assign n4512 = ~n4508 & ~n4511;
  assign n4513 = pi62 & n4512;
  assign n4514 = pi248 & ~n4513;
  assign n4515 = ~n3446 & ~n4382;
  assign n4516 = pi299 & ~n4510;
  assign n4517 = n4515 & ~n4516;
  assign n4518 = ~n2534 & n4517;
  assign n4519 = ~n2615 & n4517;
  assign n4520 = pi299 & ~n4507;
  assign n4521 = n4515 & ~n4520;
  assign n4522 = n2615 & n4521;
  assign n4523 = ~n4519 & ~n4522;
  assign n4524 = n2535 & ~n4523;
  assign n4525 = pi92 & ~n4524;
  assign n4526 = ~n2535 & n4517;
  assign n4527 = n4525 & ~n4526;
  assign n4528 = pi75 & n4517;
  assign n4529 = pi87 & n4523;
  assign n4530 = pi39 & ~n4521;
  assign n4531 = ~pi869 & n3474;
  assign n4532 = ~pi170 & ~n4531;
  assign n4533 = pi869 & ~n3380;
  assign n4534 = ~pi869 & ~n3088;
  assign n4535 = pi170 & ~n4534;
  assign n4536 = ~n4533 & n4535;
  assign n4537 = ~n4532 & ~n4536;
  assign n4538 = ~pi228 & n4537;
  assign n4539 = ~n3465 & ~n4538;
  assign n4540 = n4390 & ~n4539;
  assign n4541 = n4385 & ~n4540;
  assign n4542 = ~n4397 & ~n4541;
  assign n4543 = ~pi215 & ~n4542;
  assign n4544 = n4436 & ~n4543;
  assign n4545 = n4434 & ~n4544;
  assign n4546 = ~pi38 & ~n4545;
  assign n4547 = ~n4530 & n4546;
  assign n4548 = pi38 & n4517;
  assign n4549 = ~pi100 & ~n4548;
  assign n4550 = ~n4547 & n4549;
  assign n4551 = ~n2532 & n4517;
  assign n4552 = pi100 & ~n4551;
  assign n4553 = ~n4463 & n4502;
  assign n4554 = n4385 & ~n4553;
  assign n4555 = ~n4397 & ~n4554;
  assign n4556 = ~pi215 & ~n4555;
  assign n4557 = ~n4383 & ~n4556;
  assign n4558 = pi299 & ~n4557;
  assign n4559 = n2532 & ~n4558;
  assign n4560 = n4515 & n4559;
  assign n4561 = n4552 & ~n4560;
  assign n4562 = ~n4550 & ~n4561;
  assign n4563 = ~pi87 & ~n4562;
  assign n4564 = ~pi75 & ~n4563;
  assign n4565 = ~n4529 & n4564;
  assign n4566 = ~pi92 & ~n4565;
  assign n4567 = ~n4528 & n4566;
  assign n4568 = n2534 & ~n4567;
  assign n4569 = ~n4527 & n4568;
  assign n4570 = ~pi55 & ~n4569;
  assign n4571 = ~n4518 & n4570;
  assign n4572 = ~n2576 & n4510;
  assign n4573 = n2576 & n4507;
  assign n4574 = pi55 & ~n4573;
  assign n4575 = ~n4572 & n4574;
  assign n4576 = ~pi56 & ~n4575;
  assign n4577 = ~n4571 & n4576;
  assign n4578 = ~n2539 & ~n4510;
  assign n4579 = pi56 & ~n4578;
  assign n4580 = n2539 & ~n4507;
  assign n4581 = n4579 & ~n4580;
  assign n4582 = ~pi62 & ~n4581;
  assign n4583 = ~n4577 & n4582;
  assign n4584 = n4514 & ~n4583;
  assign n4585 = n3327 & n4584;
  assign n4586 = pi248 & n4509;
  assign n4587 = ~n3327 & ~n4586;
  assign n4588 = n4400 & n4587;
  assign n4589 = ~n4585 & ~n4588;
  assign po159 = ~n4501 & n4589;
  assign n4591 = pi215 & pi1139;
  assign n4592 = pi216 & ~pi1139;
  assign n4593 = ~pi833 & pi1139;
  assign n4594 = pi833 & pi920;
  assign n4595 = ~pi216 & ~n4594;
  assign n4596 = ~n4593 & n4595;
  assign n4597 = pi221 & ~n4596;
  assign n4598 = ~n4592 & n4597;
  assign n4599 = pi216 & pi281;
  assign n4600 = ~pi221 & ~n4599;
  assign n4601 = ~pi216 & ~pi862;
  assign n4602 = n3600 & n4601;
  assign n4603 = n4600 & ~n4602;
  assign n4604 = ~n4598 & ~n4603;
  assign n4605 = ~pi216 & ~n4597;
  assign n4606 = pi148 & ~n2441;
  assign n4607 = n4605 & n4606;
  assign n4608 = ~pi215 & ~n4607;
  assign n4609 = ~n4604 & n4608;
  assign n4610 = ~n4591 & ~n4609;
  assign n4611 = ~n3433 & ~n4610;
  assign n4612 = ~n3315 & ~n4611;
  assign n4613 = pi62 & ~n4612;
  assign n4614 = ~pi148 & ~pi215;
  assign n4615 = ~n2441 & ~n3537;
  assign n4616 = pi862 & ~n3432;
  assign n4617 = ~pi216 & ~n4616;
  assign n4618 = ~n4615 & n4617;
  assign n4619 = n4600 & ~n4618;
  assign n4620 = ~n4598 & ~n4619;
  assign n4621 = n4614 & ~n4620;
  assign n4622 = ~n3537 & ~n3600;
  assign n4623 = n4605 & n4622;
  assign n4624 = n4601 & ~n4622;
  assign n4625 = n4600 & ~n4624;
  assign n4626 = ~n4598 & ~n4625;
  assign n4627 = pi148 & ~pi215;
  assign n4628 = ~n4626 & n4627;
  assign n4629 = ~n4623 & n4628;
  assign n4630 = ~n4591 & ~n4629;
  assign n4631 = ~n4621 & n4630;
  assign n4632 = n3315 & n4631;
  assign n4633 = n4613 & ~n4632;
  assign n4634 = pi299 & n4611;
  assign n4635 = ~pi920 & n2595;
  assign n4636 = ~pi1139 & ~n2595;
  assign n4637 = pi222 & ~n4636;
  assign n4638 = ~n4635 & n4637;
  assign n4639 = pi223 & pi1139;
  assign n4640 = ~pi224 & ~n4639;
  assign n4641 = ~n4638 & n4640;
  assign n4642 = ~pi862 & n4641;
  assign n4643 = pi224 & pi281;
  assign n4644 = ~pi222 & ~n4643;
  assign n4645 = ~n4638 & ~n4644;
  assign n4646 = ~pi223 & ~n4645;
  assign n4647 = ~n4639 & ~n4646;
  assign n4648 = ~pi299 & ~n4647;
  assign n4649 = ~n4642 & n4648;
  assign n4650 = ~n3445 & n4649;
  assign n4651 = ~n4634 & ~n4650;
  assign n4652 = ~n2534 & n4651;
  assign n4653 = ~n2535 & n4651;
  assign n4654 = ~n2615 & n4651;
  assign n4655 = pi299 & ~n4631;
  assign n4656 = ~n4650 & ~n4655;
  assign n4657 = n2615 & n4656;
  assign n4658 = ~n4654 & ~n4657;
  assign n4659 = n2535 & ~n4658;
  assign n4660 = pi92 & ~n4659;
  assign n4661 = ~n4653 & n4660;
  assign n4662 = pi75 & n4651;
  assign n4663 = pi87 & n4658;
  assign n4664 = ~n2532 & n4651;
  assign n4665 = pi100 & ~n4664;
  assign n4666 = ~n2441 & ~n3401;
  assign n4667 = n4600 & n4666;
  assign n4668 = n4620 & ~n4667;
  assign n4669 = n4614 & ~n4668;
  assign n4670 = n3601 & n4600;
  assign n4671 = n4626 & ~n4670;
  assign n4672 = n3601 & n4605;
  assign n4673 = ~n4671 & ~n4672;
  assign n4674 = n4627 & n4673;
  assign n4675 = ~n4591 & ~n4674;
  assign n4676 = ~n4669 & n4675;
  assign n4677 = pi299 & ~n4676;
  assign n4678 = ~n4650 & ~n4677;
  assign n4679 = n2532 & n4678;
  assign n4680 = n4665 & ~n4679;
  assign n4681 = pi39 & ~n4656;
  assign n4682 = ~n3087 & n4641;
  assign n4683 = ~n4647 & ~n4682;
  assign n4684 = ~n4642 & n4683;
  assign n4685 = ~pi299 & ~n4684;
  assign n4686 = ~pi228 & n3380;
  assign n4687 = ~n2441 & ~n4686;
  assign n4688 = ~pi862 & n4687;
  assign n4689 = pi862 & ~n3467;
  assign n4690 = ~pi216 & ~n4689;
  assign n4691 = ~n4688 & n4690;
  assign n4692 = n4600 & ~n4691;
  assign n4693 = ~n4598 & ~n4692;
  assign n4694 = n4614 & ~n4693;
  assign n4695 = ~n4591 & ~n4694;
  assign n4696 = ~n3477 & n4601;
  assign n4697 = n4600 & ~n4696;
  assign n4698 = ~n4598 & ~n4697;
  assign n4699 = n3477 & n4605;
  assign n4700 = ~n4698 & ~n4699;
  assign n4701 = n4627 & n4700;
  assign n4702 = pi299 & ~n4701;
  assign n4703 = n4695 & n4702;
  assign n4704 = ~pi39 & ~n4703;
  assign n4705 = ~n4685 & n4704;
  assign n4706 = ~pi38 & ~n4705;
  assign n4707 = ~n4681 & n4706;
  assign n4708 = pi38 & n4651;
  assign n4709 = ~pi100 & ~n4708;
  assign n4710 = ~n4707 & n4709;
  assign n4711 = ~n4680 & ~n4710;
  assign n4712 = ~pi87 & ~n4711;
  assign n4713 = ~pi75 & ~n4712;
  assign n4714 = ~n4663 & n4713;
  assign n4715 = ~pi92 & ~n4714;
  assign n4716 = ~n4662 & n4715;
  assign n4717 = n2534 & ~n4716;
  assign n4718 = ~n4661 & n4717;
  assign n4719 = ~pi55 & ~n4718;
  assign n4720 = ~n4652 & n4719;
  assign n4721 = ~n2576 & ~n4611;
  assign n4722 = pi55 & ~n4721;
  assign n4723 = n2576 & n4631;
  assign n4724 = n4722 & ~n4723;
  assign n4725 = ~pi56 & ~n4724;
  assign n4726 = ~n4720 & n4725;
  assign n4727 = ~n2539 & n4611;
  assign n4728 = n2539 & ~n4631;
  assign n4729 = pi56 & ~n4728;
  assign n4730 = ~n4727 & n4729;
  assign n4731 = ~pi62 & ~n4730;
  assign n4732 = ~n4726 & n4731;
  assign n4733 = n3327 & ~n4732;
  assign n4734 = ~n4633 & n4733;
  assign n4735 = ~n3327 & ~n4611;
  assign n4736 = ~pi247 & ~n4735;
  assign n4737 = ~n4734 & n4736;
  assign n4738 = ~n3315 & n4610;
  assign n4739 = pi62 & ~n4738;
  assign n4740 = n4608 & ~n4626;
  assign n4741 = n4630 & ~n4740;
  assign n4742 = n3315 & n4741;
  assign n4743 = n4739 & ~n4742;
  assign n4744 = ~n3446 & ~n4649;
  assign n4745 = pi299 & ~n4610;
  assign n4746 = n4744 & ~n4745;
  assign n4747 = ~n2534 & n4746;
  assign n4748 = ~n2615 & n4746;
  assign n4749 = pi299 & ~n4741;
  assign n4750 = n4744 & ~n4749;
  assign n4751 = n2615 & n4750;
  assign n4752 = ~n4748 & ~n4751;
  assign n4753 = n2535 & ~n4752;
  assign n4754 = pi92 & ~n4753;
  assign n4755 = ~n2535 & n4746;
  assign n4756 = n4754 & ~n4755;
  assign n4757 = pi75 & n4746;
  assign n4758 = pi87 & n4752;
  assign n4759 = ~n2532 & n4746;
  assign n4760 = pi100 & ~n4759;
  assign n4761 = n4614 & ~n4671;
  assign n4762 = n4605 & n4666;
  assign n4763 = n4628 & ~n4762;
  assign n4764 = ~n4591 & ~n4763;
  assign n4765 = ~n4761 & n4764;
  assign n4766 = pi299 & ~n4765;
  assign n4767 = n2532 & ~n4766;
  assign n4768 = n4744 & n4767;
  assign n4769 = n4760 & ~n4768;
  assign n4770 = pi39 & ~n4750;
  assign n4771 = n3087 & n4642;
  assign n4772 = n4648 & ~n4771;
  assign n4773 = pi862 & ~n4687;
  assign n4774 = ~pi862 & n3467;
  assign n4775 = ~pi216 & ~n4774;
  assign n4776 = ~n4773 & n4775;
  assign n4777 = n4600 & ~n4776;
  assign n4778 = ~n4598 & ~n4777;
  assign n4779 = n4627 & ~n4778;
  assign n4780 = n4614 & ~n4698;
  assign n4781 = ~n4591 & ~n4780;
  assign n4782 = ~n4779 & n4781;
  assign n4783 = pi299 & ~n4782;
  assign n4784 = ~n4772 & ~n4783;
  assign n4785 = ~pi39 & ~n4784;
  assign n4786 = ~pi38 & ~n4785;
  assign n4787 = ~n4770 & n4786;
  assign n4788 = pi38 & n4746;
  assign n4789 = ~pi100 & ~n4788;
  assign n4790 = ~n4787 & n4789;
  assign n4791 = ~n4769 & ~n4790;
  assign n4792 = ~pi87 & ~n4791;
  assign n4793 = ~pi75 & ~n4792;
  assign n4794 = ~n4758 & n4793;
  assign n4795 = ~pi92 & ~n4794;
  assign n4796 = ~n4757 & n4795;
  assign n4797 = n2534 & ~n4796;
  assign n4798 = ~n4756 & n4797;
  assign n4799 = ~pi55 & ~n4798;
  assign n4800 = ~n4747 & n4799;
  assign n4801 = ~n2576 & n4610;
  assign n4802 = pi55 & ~n4801;
  assign n4803 = n2576 & n4741;
  assign n4804 = n4802 & ~n4803;
  assign n4805 = ~pi56 & ~n4804;
  assign n4806 = ~n4800 & n4805;
  assign n4807 = ~n2539 & ~n4610;
  assign n4808 = pi56 & ~n4807;
  assign n4809 = n2539 & ~n4741;
  assign n4810 = n4808 & ~n4809;
  assign n4811 = ~pi62 & ~n4810;
  assign n4812 = ~n4806 & n4811;
  assign n4813 = n3327 & ~n4812;
  assign n4814 = ~n4743 & n4813;
  assign n4815 = ~n3327 & n4610;
  assign n4816 = pi247 & ~n4815;
  assign n4817 = ~n4814 & n4816;
  assign po160 = n4737 | n4817;
  assign n4819 = pi223 & pi1138;
  assign n4820 = pi224 & pi269;
  assign n4821 = ~pi222 & ~n4820;
  assign n4822 = pi877 & ~n2442;
  assign n4823 = ~pi224 & ~n4822;
  assign n4824 = n4821 & ~n4823;
  assign n4825 = ~pi940 & n2595;
  assign n4826 = ~pi1138 & ~n2595;
  assign n4827 = pi222 & ~n4826;
  assign n4828 = ~n4825 & n4827;
  assign n4829 = ~n4824 & ~n4828;
  assign n4830 = ~pi223 & ~n4829;
  assign n4831 = ~n4819 & ~n4830;
  assign n4832 = ~pi299 & ~n4831;
  assign n4833 = pi215 & pi1138;
  assign n4834 = pi216 & pi269;
  assign n4835 = ~pi221 & ~n4834;
  assign n4836 = pi105 & ~n4822;
  assign n4837 = ~pi105 & pi169;
  assign n4838 = pi228 & ~n4837;
  assign n4839 = ~n4836 & n4838;
  assign n4840 = ~pi216 & ~n4839;
  assign n4841 = ~pi169 & ~pi228;
  assign n4842 = n4840 & ~n4841;
  assign n4843 = n4835 & ~n4842;
  assign n4844 = ~pi940 & n2452;
  assign n4845 = ~pi1138 & ~n2452;
  assign n4846 = pi221 & ~n4845;
  assign n4847 = ~n4844 & n4846;
  assign n4848 = ~n4843 & ~n4847;
  assign n4849 = ~pi215 & ~n4848;
  assign n4850 = ~n4833 & ~n4849;
  assign n4851 = pi299 & ~n4850;
  assign n4852 = ~n4832 & ~n4851;
  assign n4853 = ~n2534 & n4852;
  assign n4854 = ~n2535 & n4852;
  assign n4855 = ~n2615 & n4852;
  assign n4856 = pi169 & ~n2522;
  assign n4857 = ~pi877 & n2522;
  assign n4858 = ~pi228 & ~n4857;
  assign n4859 = ~n4856 & n4858;
  assign n4860 = n4840 & ~n4859;
  assign n4861 = n4835 & ~n4860;
  assign n4862 = ~n4847 & ~n4861;
  assign n4863 = ~pi215 & ~n4862;
  assign n4864 = ~n4833 & ~n4863;
  assign n4865 = pi299 & ~n4864;
  assign n4866 = ~n4832 & ~n4865;
  assign n4867 = n2615 & n4866;
  assign n4868 = ~n4855 & ~n4867;
  assign n4869 = n2535 & ~n4868;
  assign n4870 = pi92 & ~n4869;
  assign n4871 = ~n4854 & n4870;
  assign n4872 = pi75 & n4852;
  assign n4873 = pi87 & n4868;
  assign n4874 = pi39 & ~n4866;
  assign n4875 = ~pi299 & ~n4819;
  assign n4876 = pi877 & n3087;
  assign n4877 = ~pi224 & ~n4876;
  assign n4878 = n4821 & ~n4877;
  assign n4879 = ~n4828 & ~n4878;
  assign n4880 = ~n3087 & n4821;
  assign n4881 = n4879 & ~n4880;
  assign n4882 = ~pi223 & ~n4881;
  assign n4883 = n4875 & ~n4882;
  assign n4884 = ~pi39 & ~n4883;
  assign n4885 = n4875 & n4879;
  assign n4886 = pi299 & ~n4833;
  assign n4887 = pi877 & n3088;
  assign n4888 = ~pi877 & n3380;
  assign n4889 = ~pi169 & ~n4888;
  assign n4890 = ~n4887 & n4889;
  assign n4891 = pi169 & n3474;
  assign n4892 = pi877 & n4891;
  assign n4893 = ~n4890 & ~n4892;
  assign n4894 = ~pi228 & ~n4893;
  assign n4895 = ~n3464 & n4839;
  assign n4896 = ~pi216 & ~n4895;
  assign n4897 = ~n4894 & n4896;
  assign n4898 = n4835 & ~n4897;
  assign n4899 = ~n4847 & ~n4898;
  assign n4900 = ~pi215 & ~n4899;
  assign n4901 = n4886 & ~n4900;
  assign n4902 = ~n4885 & ~n4901;
  assign n4903 = n4884 & n4902;
  assign n4904 = ~pi38 & ~n4903;
  assign n4905 = ~n4874 & n4904;
  assign n4906 = pi38 & n4852;
  assign n4907 = ~pi100 & ~n4906;
  assign n4908 = ~n4905 & n4907;
  assign n4909 = ~n2532 & n4852;
  assign n4910 = pi100 & ~n4909;
  assign n4911 = ~pi877 & n3400;
  assign n4912 = ~n3401 & ~n4841;
  assign n4913 = ~n4911 & ~n4912;
  assign n4914 = n4840 & ~n4913;
  assign n4915 = n4835 & ~n4914;
  assign n4916 = ~n4847 & ~n4915;
  assign n4917 = ~pi215 & ~n4916;
  assign n4918 = ~n4833 & ~n4917;
  assign n4919 = pi299 & ~n4918;
  assign n4920 = ~n4832 & ~n4919;
  assign n4921 = n2532 & n4920;
  assign n4922 = n4910 & ~n4921;
  assign n4923 = ~n4908 & ~n4922;
  assign n4924 = ~pi87 & ~n4923;
  assign n4925 = ~pi75 & ~n4924;
  assign n4926 = ~n4873 & n4925;
  assign n4927 = ~pi92 & ~n4926;
  assign n4928 = ~n4872 & n4927;
  assign n4929 = n2534 & ~n4928;
  assign n4930 = ~n4871 & n4929;
  assign n4931 = ~pi55 & ~n4930;
  assign n4932 = ~n4853 & n4931;
  assign n4933 = ~n2576 & n4850;
  assign n4934 = pi55 & ~n4933;
  assign n4935 = n2576 & n4864;
  assign n4936 = n4934 & ~n4935;
  assign n4937 = ~pi56 & ~n4936;
  assign n4938 = ~n4932 & n4937;
  assign n4939 = ~n2539 & ~n4850;
  assign n4940 = pi56 & ~n4939;
  assign n4941 = n2539 & ~n4864;
  assign n4942 = n4940 & ~n4941;
  assign n4943 = ~pi62 & ~n4942;
  assign n4944 = ~n4938 & n4943;
  assign n4945 = n3327 & ~n4944;
  assign n4946 = ~n3315 & n4850;
  assign n4947 = n3315 & n4864;
  assign n4948 = ~n4946 & ~n4947;
  assign n4949 = pi62 & n4948;
  assign n4950 = ~pi246 & ~n4949;
  assign n4951 = n4945 & n4950;
  assign n4952 = ~n3432 & n4840;
  assign n4953 = ~n4859 & n4952;
  assign n4954 = n4835 & ~n4953;
  assign n4955 = ~n4847 & ~n4954;
  assign n4956 = ~pi215 & ~n4955;
  assign n4957 = ~n4833 & ~n4956;
  assign n4958 = n3315 & n4957;
  assign n4959 = n3532 & ~n4834;
  assign n4960 = n4850 & ~n4959;
  assign n4961 = ~n3315 & n4960;
  assign n4962 = ~n4958 & ~n4961;
  assign n4963 = pi62 & n4962;
  assign n4964 = pi246 & ~n4963;
  assign n4965 = ~n3446 & ~n4832;
  assign n4966 = pi299 & ~n4960;
  assign n4967 = n4965 & ~n4966;
  assign n4968 = ~n2534 & n4967;
  assign n4969 = ~n2615 & n4967;
  assign n4970 = pi299 & ~n4957;
  assign n4971 = n4965 & ~n4970;
  assign n4972 = n2615 & n4971;
  assign n4973 = ~n4969 & ~n4972;
  assign n4974 = n2535 & ~n4973;
  assign n4975 = pi92 & ~n4974;
  assign n4976 = ~n2535 & n4967;
  assign n4977 = n4975 & ~n4976;
  assign n4978 = pi75 & n4967;
  assign n4979 = pi87 & n4973;
  assign n4980 = pi39 & ~n4971;
  assign n4981 = ~pi877 & n3474;
  assign n4982 = ~pi169 & ~n4981;
  assign n4983 = pi877 & ~n3380;
  assign n4984 = ~pi877 & ~n3088;
  assign n4985 = pi169 & ~n4984;
  assign n4986 = ~n4983 & n4985;
  assign n4987 = ~n4982 & ~n4986;
  assign n4988 = ~pi228 & n4987;
  assign n4989 = ~n3465 & ~n4988;
  assign n4990 = n4840 & ~n4989;
  assign n4991 = n4835 & ~n4990;
  assign n4992 = ~n4847 & ~n4991;
  assign n4993 = ~pi215 & ~n4992;
  assign n4994 = n4886 & ~n4993;
  assign n4995 = n4884 & ~n4994;
  assign n4996 = ~pi38 & ~n4995;
  assign n4997 = ~n4980 & n4996;
  assign n4998 = pi38 & n4967;
  assign n4999 = ~pi100 & ~n4998;
  assign n5000 = ~n4997 & n4999;
  assign n5001 = ~n2532 & n4967;
  assign n5002 = pi100 & ~n5001;
  assign n5003 = ~n4913 & n4952;
  assign n5004 = n4835 & ~n5003;
  assign n5005 = ~n4847 & ~n5004;
  assign n5006 = ~pi215 & ~n5005;
  assign n5007 = ~n4833 & ~n5006;
  assign n5008 = pi299 & ~n5007;
  assign n5009 = n2532 & ~n5008;
  assign n5010 = n4965 & n5009;
  assign n5011 = n5002 & ~n5010;
  assign n5012 = ~n5000 & ~n5011;
  assign n5013 = ~pi87 & ~n5012;
  assign n5014 = ~pi75 & ~n5013;
  assign n5015 = ~n4979 & n5014;
  assign n5016 = ~pi92 & ~n5015;
  assign n5017 = ~n4978 & n5016;
  assign n5018 = n2534 & ~n5017;
  assign n5019 = ~n4977 & n5018;
  assign n5020 = ~pi55 & ~n5019;
  assign n5021 = ~n4968 & n5020;
  assign n5022 = ~n2576 & n4960;
  assign n5023 = n2576 & n4957;
  assign n5024 = pi55 & ~n5023;
  assign n5025 = ~n5022 & n5024;
  assign n5026 = ~pi56 & ~n5025;
  assign n5027 = ~n5021 & n5026;
  assign n5028 = ~n2539 & ~n4960;
  assign n5029 = pi56 & ~n5028;
  assign n5030 = n2539 & ~n4957;
  assign n5031 = n5029 & ~n5030;
  assign n5032 = ~pi62 & ~n5031;
  assign n5033 = ~n5027 & n5032;
  assign n5034 = n4964 & ~n5033;
  assign n5035 = n3327 & n5034;
  assign n5036 = pi246 & n4959;
  assign n5037 = ~n3327 & ~n5036;
  assign n5038 = n4850 & n5037;
  assign n5039 = ~n5035 & ~n5038;
  assign po161 = ~n4951 & n5039;
  assign n5041 = pi223 & pi1137;
  assign n5042 = pi224 & pi280;
  assign n5043 = ~pi222 & ~n5042;
  assign n5044 = pi878 & ~n2442;
  assign n5045 = ~pi224 & ~n5044;
  assign n5046 = n5043 & ~n5045;
  assign n5047 = ~pi933 & n2595;
  assign n5048 = ~pi1137 & ~n2595;
  assign n5049 = pi222 & ~n5048;
  assign n5050 = ~n5047 & n5049;
  assign n5051 = ~n5046 & ~n5050;
  assign n5052 = ~pi223 & ~n5051;
  assign n5053 = ~n5041 & ~n5052;
  assign n5054 = ~pi299 & ~n5053;
  assign n5055 = pi215 & pi1137;
  assign n5056 = pi216 & pi280;
  assign n5057 = ~pi221 & ~n5056;
  assign n5058 = pi105 & ~n5044;
  assign n5059 = ~pi105 & pi168;
  assign n5060 = pi228 & ~n5059;
  assign n5061 = ~n5058 & n5060;
  assign n5062 = ~pi216 & ~n5061;
  assign n5063 = ~pi168 & ~pi228;
  assign n5064 = n5062 & ~n5063;
  assign n5065 = n5057 & ~n5064;
  assign n5066 = ~pi933 & n2452;
  assign n5067 = ~pi1137 & ~n2452;
  assign n5068 = pi221 & ~n5067;
  assign n5069 = ~n5066 & n5068;
  assign n5070 = ~n5065 & ~n5069;
  assign n5071 = ~pi215 & ~n5070;
  assign n5072 = ~n5055 & ~n5071;
  assign n5073 = pi299 & ~n5072;
  assign n5074 = ~n5054 & ~n5073;
  assign n5075 = ~n2534 & n5074;
  assign n5076 = ~n2535 & n5074;
  assign n5077 = ~n2615 & n5074;
  assign n5078 = ~pi878 & n2522;
  assign n5079 = ~n3537 & ~n5063;
  assign n5080 = ~n5078 & ~n5079;
  assign n5081 = n5062 & ~n5080;
  assign n5082 = n5057 & ~n5081;
  assign n5083 = ~n5069 & ~n5082;
  assign n5084 = ~pi215 & ~n5083;
  assign n5085 = ~n5055 & ~n5084;
  assign n5086 = pi299 & ~n5085;
  assign n5087 = ~n5054 & ~n5086;
  assign n5088 = n2615 & n5087;
  assign n5089 = ~n5077 & ~n5088;
  assign n5090 = n2535 & ~n5089;
  assign n5091 = pi92 & ~n5090;
  assign n5092 = ~n5076 & n5091;
  assign n5093 = pi75 & n5074;
  assign n5094 = pi87 & n5089;
  assign n5095 = pi39 & ~n5087;
  assign n5096 = ~pi299 & ~n5041;
  assign n5097 = pi878 & n3087;
  assign n5098 = ~pi224 & ~n5097;
  assign n5099 = n5043 & ~n5098;
  assign n5100 = ~n5050 & ~n5099;
  assign n5101 = ~n3087 & n5043;
  assign n5102 = n5100 & ~n5101;
  assign n5103 = ~pi223 & ~n5102;
  assign n5104 = n5096 & ~n5103;
  assign n5105 = ~pi39 & ~n5104;
  assign n5106 = n5096 & n5100;
  assign n5107 = pi299 & ~n5055;
  assign n5108 = pi878 & n3088;
  assign n5109 = ~pi878 & n3380;
  assign n5110 = ~pi168 & ~n5109;
  assign n5111 = ~n5108 & n5110;
  assign n5112 = pi168 & n3474;
  assign n5113 = pi878 & n5112;
  assign n5114 = ~n5111 & ~n5113;
  assign n5115 = ~pi228 & ~n5114;
  assign n5116 = ~n3464 & n5061;
  assign n5117 = ~pi216 & ~n5116;
  assign n5118 = ~n5115 & n5117;
  assign n5119 = n5057 & ~n5118;
  assign n5120 = ~n5069 & ~n5119;
  assign n5121 = ~pi215 & ~n5120;
  assign n5122 = n5107 & ~n5121;
  assign n5123 = ~n5106 & ~n5122;
  assign n5124 = n5105 & n5123;
  assign n5125 = ~pi38 & ~n5124;
  assign n5126 = ~n5095 & n5125;
  assign n5127 = pi38 & n5074;
  assign n5128 = ~pi100 & ~n5127;
  assign n5129 = ~n5126 & n5128;
  assign n5130 = ~n2532 & n5074;
  assign n5131 = pi100 & ~n5130;
  assign n5132 = ~pi878 & n3400;
  assign n5133 = ~n3401 & ~n5063;
  assign n5134 = ~n5132 & ~n5133;
  assign n5135 = n5062 & ~n5134;
  assign n5136 = n5057 & ~n5135;
  assign n5137 = ~n5069 & ~n5136;
  assign n5138 = ~pi215 & ~n5137;
  assign n5139 = ~n5055 & ~n5138;
  assign n5140 = pi299 & ~n5139;
  assign n5141 = ~n5054 & ~n5140;
  assign n5142 = n2532 & n5141;
  assign n5143 = n5131 & ~n5142;
  assign n5144 = ~n5129 & ~n5143;
  assign n5145 = ~pi87 & ~n5144;
  assign n5146 = ~pi75 & ~n5145;
  assign n5147 = ~n5094 & n5146;
  assign n5148 = ~pi92 & ~n5147;
  assign n5149 = ~n5093 & n5148;
  assign n5150 = n2534 & ~n5149;
  assign n5151 = ~n5092 & n5150;
  assign n5152 = ~pi55 & ~n5151;
  assign n5153 = ~n5075 & n5152;
  assign n5154 = ~n2576 & n5072;
  assign n5155 = pi55 & ~n5154;
  assign n5156 = n2576 & n5085;
  assign n5157 = n5155 & ~n5156;
  assign n5158 = ~pi56 & ~n5157;
  assign n5159 = ~n5153 & n5158;
  assign n5160 = ~n2539 & ~n5072;
  assign n5161 = pi56 & ~n5160;
  assign n5162 = n2539 & ~n5085;
  assign n5163 = n5161 & ~n5162;
  assign n5164 = ~pi62 & ~n5163;
  assign n5165 = ~n5159 & n5164;
  assign n5166 = n3327 & ~n5165;
  assign n5167 = ~n3315 & n5072;
  assign n5168 = n3315 & n5085;
  assign n5169 = ~n5167 & ~n5168;
  assign n5170 = pi62 & n5169;
  assign n5171 = ~pi240 & ~n5170;
  assign n5172 = n5166 & n5171;
  assign n5173 = ~n3432 & n5062;
  assign n5174 = ~n5080 & n5173;
  assign n5175 = n5057 & ~n5174;
  assign n5176 = ~n5069 & ~n5175;
  assign n5177 = ~pi215 & ~n5176;
  assign n5178 = ~n5055 & ~n5177;
  assign n5179 = n3315 & n5178;
  assign n5180 = n3532 & ~n5056;
  assign n5181 = n5072 & ~n5180;
  assign n5182 = ~n3315 & n5181;
  assign n5183 = ~n5179 & ~n5182;
  assign n5184 = pi62 & n5183;
  assign n5185 = pi240 & ~n5184;
  assign n5186 = ~n3446 & ~n5054;
  assign n5187 = pi299 & ~n5181;
  assign n5188 = n5186 & ~n5187;
  assign n5189 = ~n2534 & n5188;
  assign n5190 = ~n2615 & n5188;
  assign n5191 = pi299 & ~n5178;
  assign n5192 = n5186 & ~n5191;
  assign n5193 = n2615 & n5192;
  assign n5194 = ~n5190 & ~n5193;
  assign n5195 = n2535 & ~n5194;
  assign n5196 = pi92 & ~n5195;
  assign n5197 = ~n2535 & n5188;
  assign n5198 = n5196 & ~n5197;
  assign n5199 = pi75 & n5188;
  assign n5200 = pi87 & n5194;
  assign n5201 = pi39 & ~n5192;
  assign n5202 = ~pi878 & n3474;
  assign n5203 = ~pi168 & ~n5202;
  assign n5204 = pi878 & ~n3380;
  assign n5205 = ~pi878 & ~n3088;
  assign n5206 = pi168 & ~n5205;
  assign n5207 = ~n5204 & n5206;
  assign n5208 = ~n5203 & ~n5207;
  assign n5209 = ~pi228 & n5208;
  assign n5210 = ~n3465 & ~n5209;
  assign n5211 = n5062 & ~n5210;
  assign n5212 = n5057 & ~n5211;
  assign n5213 = ~n5069 & ~n5212;
  assign n5214 = ~pi215 & ~n5213;
  assign n5215 = n5107 & ~n5214;
  assign n5216 = n5105 & ~n5215;
  assign n5217 = ~pi38 & ~n5216;
  assign n5218 = ~n5201 & n5217;
  assign n5219 = pi38 & n5188;
  assign n5220 = ~pi100 & ~n5219;
  assign n5221 = ~n5218 & n5220;
  assign n5222 = ~n2532 & n5188;
  assign n5223 = pi100 & ~n5222;
  assign n5224 = ~n5134 & n5173;
  assign n5225 = n5057 & ~n5224;
  assign n5226 = ~n5069 & ~n5225;
  assign n5227 = ~pi215 & ~n5226;
  assign n5228 = ~n5055 & ~n5227;
  assign n5229 = pi299 & ~n5228;
  assign n5230 = n2532 & ~n5229;
  assign n5231 = n5186 & n5230;
  assign n5232 = n5223 & ~n5231;
  assign n5233 = ~n5221 & ~n5232;
  assign n5234 = ~pi87 & ~n5233;
  assign n5235 = ~pi75 & ~n5234;
  assign n5236 = ~n5200 & n5235;
  assign n5237 = ~pi92 & ~n5236;
  assign n5238 = ~n5199 & n5237;
  assign n5239 = n2534 & ~n5238;
  assign n5240 = ~n5198 & n5239;
  assign n5241 = ~pi55 & ~n5240;
  assign n5242 = ~n5189 & n5241;
  assign n5243 = ~n2576 & n5181;
  assign n5244 = n2576 & n5178;
  assign n5245 = pi55 & ~n5244;
  assign n5246 = ~n5243 & n5245;
  assign n5247 = ~pi56 & ~n5246;
  assign n5248 = ~n5242 & n5247;
  assign n5249 = ~n2539 & ~n5181;
  assign n5250 = pi56 & ~n5249;
  assign n5251 = n2539 & ~n5178;
  assign n5252 = n5250 & ~n5251;
  assign n5253 = ~pi62 & ~n5252;
  assign n5254 = ~n5248 & n5253;
  assign n5255 = n5185 & ~n5254;
  assign n5256 = n3327 & n5255;
  assign n5257 = pi240 & n5180;
  assign n5258 = ~n3327 & ~n5257;
  assign n5259 = n5072 & n5258;
  assign n5260 = ~n5256 & ~n5259;
  assign po162 = ~n5172 & n5260;
  assign n5262 = pi215 & pi1136;
  assign n5263 = pi216 & pi266;
  assign n5264 = pi875 & ~n2442;
  assign n5265 = pi105 & ~n5264;
  assign n5266 = ~pi105 & ~pi166;
  assign n5267 = ~n5265 & ~n5266;
  assign n5268 = pi228 & n5267;
  assign n5269 = pi166 & ~pi228;
  assign n5270 = ~n5268 & ~n5269;
  assign n5271 = ~pi216 & ~n5270;
  assign n5272 = ~n5263 & ~n5271;
  assign n5273 = ~pi221 & ~n5272;
  assign n5274 = ~pi928 & n2452;
  assign n5275 = ~pi1136 & ~n2452;
  assign n5276 = pi221 & ~n5275;
  assign n5277 = ~n5274 & n5276;
  assign n5278 = ~n5273 & ~n5277;
  assign n5279 = ~pi215 & ~n5278;
  assign n5280 = ~n5262 & ~n5279;
  assign n5281 = ~n3433 & n5280;
  assign n5282 = ~n3315 & n5281;
  assign n5283 = ~pi875 & n2522;
  assign n5284 = ~n3537 & ~n5269;
  assign n5285 = ~n5283 & ~n5284;
  assign n5286 = ~n3432 & ~n5268;
  assign n5287 = ~n5285 & n5286;
  assign n5288 = ~pi216 & ~n5287;
  assign n5289 = ~n5263 & ~n5288;
  assign n5290 = ~pi221 & ~n5289;
  assign n5291 = ~n5277 & ~n5290;
  assign n5292 = ~pi215 & ~n5291;
  assign n5293 = ~n5262 & ~n5292;
  assign n5294 = n3315 & n5293;
  assign n5295 = pi62 & ~n5294;
  assign n5296 = ~n5282 & n5295;
  assign n5297 = pi223 & pi1136;
  assign n5298 = pi224 & ~pi266;
  assign n5299 = ~pi222 & ~n5298;
  assign n5300 = ~pi224 & ~pi875;
  assign n5301 = ~n2442 & n5300;
  assign n5302 = n5299 & ~n5301;
  assign n5303 = ~pi928 & n2595;
  assign n5304 = ~pi1136 & ~n2595;
  assign n5305 = pi222 & ~n5304;
  assign n5306 = ~n5303 & n5305;
  assign n5307 = ~n5302 & ~n5306;
  assign n5308 = ~pi223 & ~n5307;
  assign n5309 = ~n5297 & ~n5308;
  assign n5310 = ~pi299 & ~n5309;
  assign n5311 = pi299 & ~n5281;
  assign n5312 = ~n5310 & ~n5311;
  assign n5313 = ~n2534 & n5312;
  assign n5314 = ~n2535 & n5312;
  assign n5315 = ~n2615 & n5312;
  assign n5316 = pi299 & ~n5293;
  assign n5317 = ~n5310 & ~n5316;
  assign n5318 = n2615 & n5317;
  assign n5319 = ~n5315 & ~n5318;
  assign n5320 = n2535 & ~n5319;
  assign n5321 = pi92 & ~n5320;
  assign n5322 = ~n5314 & n5321;
  assign n5323 = pi75 & n5312;
  assign n5324 = pi87 & n5319;
  assign n5325 = pi39 & ~n5317;
  assign n5326 = ~pi299 & ~n5297;
  assign n5327 = n2607 & ~n3087;
  assign n5328 = n5307 & ~n5327;
  assign n5329 = ~pi223 & ~n5328;
  assign n5330 = n5326 & ~n5329;
  assign n5331 = ~pi39 & ~n5330;
  assign n5332 = pi299 & ~n5262;
  assign n5333 = n3465 & ~n5267;
  assign n5334 = ~pi216 & ~n5333;
  assign n5335 = ~pi166 & ~n3380;
  assign n5336 = pi875 & ~n5335;
  assign n5337 = pi166 & n3474;
  assign n5338 = ~pi166 & ~n3088;
  assign n5339 = ~pi875 & ~n5338;
  assign n5340 = ~n5337 & n5339;
  assign n5341 = ~pi228 & ~n5340;
  assign n5342 = ~n5336 & n5341;
  assign n5343 = n5334 & ~n5342;
  assign n5344 = ~n5263 & ~n5343;
  assign n5345 = ~pi221 & ~n5344;
  assign n5346 = ~n5277 & ~n5345;
  assign n5347 = ~pi215 & ~n5346;
  assign n5348 = n5332 & ~n5347;
  assign n5349 = n5331 & ~n5348;
  assign n5350 = ~pi38 & ~n5349;
  assign n5351 = ~n5325 & n5350;
  assign n5352 = pi38 & n5312;
  assign n5353 = ~pi100 & ~n5352;
  assign n5354 = ~n5351 & n5353;
  assign n5355 = ~n2532 & n5312;
  assign n5356 = pi100 & ~n5355;
  assign n5357 = ~pi875 & n3393;
  assign n5358 = pi166 & ~n5357;
  assign n5359 = ~n2626 & ~n3393;
  assign n5360 = n2626 & ~n3391;
  assign n5361 = pi875 & ~n5360;
  assign n5362 = ~n5359 & n5361;
  assign n5363 = ~n5358 & ~n5362;
  assign n5364 = ~pi228 & ~n5363;
  assign n5365 = n5286 & ~n5364;
  assign n5366 = ~pi216 & ~n5365;
  assign n5367 = ~n5263 & ~n5366;
  assign n5368 = ~pi221 & ~n5367;
  assign n5369 = ~n5277 & ~n5368;
  assign n5370 = ~pi215 & ~n5369;
  assign n5371 = ~n5262 & ~n5370;
  assign n5372 = pi299 & ~n5371;
  assign n5373 = ~n5310 & ~n5372;
  assign n5374 = n2532 & n5373;
  assign n5375 = n5356 & ~n5374;
  assign n5376 = ~n5354 & ~n5375;
  assign n5377 = ~pi87 & ~n5376;
  assign n5378 = ~pi75 & ~n5377;
  assign n5379 = ~n5324 & n5378;
  assign n5380 = ~pi92 & ~n5379;
  assign n5381 = ~n5323 & n5380;
  assign n5382 = n2534 & ~n5381;
  assign n5383 = ~n5322 & n5382;
  assign n5384 = ~pi55 & ~n5383;
  assign n5385 = ~n5313 & n5384;
  assign n5386 = ~n2576 & n5281;
  assign n5387 = n2576 & n5293;
  assign n5388 = pi55 & ~n5387;
  assign n5389 = ~n5386 & n5388;
  assign n5390 = ~pi56 & ~n5389;
  assign n5391 = ~n5385 & n5390;
  assign n5392 = ~n2539 & ~n5281;
  assign n5393 = pi56 & ~n5392;
  assign n5394 = n2539 & ~n5293;
  assign n5395 = n5393 & ~n5394;
  assign n5396 = ~pi62 & ~n5395;
  assign n5397 = ~n5391 & n5396;
  assign n5398 = n3327 & ~n5397;
  assign n5399 = ~n5296 & n5398;
  assign n5400 = ~n3327 & n5280;
  assign n5401 = ~n3433 & n5400;
  assign n5402 = pi245 & ~n5401;
  assign n5403 = ~n5399 & n5402;
  assign n5404 = ~n3315 & n5280;
  assign n5405 = pi62 & ~n5404;
  assign n5406 = ~n5268 & ~n5285;
  assign n5407 = ~pi216 & ~n5406;
  assign n5408 = ~n5263 & ~n5407;
  assign n5409 = ~pi221 & ~n5408;
  assign n5410 = ~n5277 & ~n5409;
  assign n5411 = ~pi215 & ~n5410;
  assign n5412 = ~n5262 & ~n5411;
  assign n5413 = n3315 & n5412;
  assign n5414 = n5405 & ~n5413;
  assign n5415 = pi299 & ~n5280;
  assign n5416 = ~n3445 & n5310;
  assign n5417 = ~n5415 & ~n5416;
  assign n5418 = ~n2534 & n5417;
  assign n5419 = ~n2535 & n5417;
  assign n5420 = ~n2615 & n5417;
  assign n5421 = pi299 & ~n5412;
  assign n5422 = ~n5416 & ~n5421;
  assign n5423 = n2615 & n5422;
  assign n5424 = ~n5420 & ~n5423;
  assign n5425 = n2535 & ~n5424;
  assign n5426 = pi92 & ~n5425;
  assign n5427 = ~n5419 & n5426;
  assign n5428 = pi75 & n5417;
  assign n5429 = pi87 & n5424;
  assign n5430 = pi39 & ~n5422;
  assign n5431 = ~pi166 & ~n3474;
  assign n5432 = pi166 & n3088;
  assign n5433 = pi875 & ~n5432;
  assign n5434 = ~n5431 & n5433;
  assign n5435 = ~pi875 & ~n3380;
  assign n5436 = pi166 & n5435;
  assign n5437 = ~pi228 & ~n5436;
  assign n5438 = ~n5434 & n5437;
  assign n5439 = ~n3859 & ~n5438;
  assign n5440 = n5334 & n5439;
  assign n5441 = ~n5263 & ~n5440;
  assign n5442 = ~pi221 & ~n5441;
  assign n5443 = ~n5277 & ~n5442;
  assign n5444 = ~pi215 & ~n5443;
  assign n5445 = n5332 & ~n5444;
  assign n5446 = n5302 & ~n5327;
  assign n5447 = n5326 & ~n5446;
  assign n5448 = ~n5306 & n5447;
  assign n5449 = ~n5445 & ~n5448;
  assign n5450 = n5331 & n5449;
  assign n5451 = ~pi38 & ~n5450;
  assign n5452 = ~n5430 & n5451;
  assign n5453 = pi38 & n5417;
  assign n5454 = ~pi100 & ~n5453;
  assign n5455 = ~n5452 & n5454;
  assign n5456 = ~n2532 & n5417;
  assign n5457 = pi100 & ~n5456;
  assign n5458 = ~n5268 & ~n5364;
  assign n5459 = ~pi216 & ~n5458;
  assign n5460 = ~n5263 & ~n5459;
  assign n5461 = ~pi221 & ~n5460;
  assign n5462 = ~n5277 & ~n5461;
  assign n5463 = ~pi215 & ~n5462;
  assign n5464 = ~n5262 & ~n5463;
  assign n5465 = pi299 & ~n5464;
  assign n5466 = ~n5416 & ~n5465;
  assign n5467 = n2532 & n5466;
  assign n5468 = n5457 & ~n5467;
  assign n5469 = ~n5455 & ~n5468;
  assign n5470 = ~pi87 & ~n5469;
  assign n5471 = ~pi75 & ~n5470;
  assign n5472 = ~n5429 & n5471;
  assign n5473 = ~pi92 & ~n5472;
  assign n5474 = ~n5428 & n5473;
  assign n5475 = n2534 & ~n5474;
  assign n5476 = ~n5427 & n5475;
  assign n5477 = ~pi55 & ~n5476;
  assign n5478 = ~n5418 & n5477;
  assign n5479 = ~n2576 & n5280;
  assign n5480 = pi55 & ~n5479;
  assign n5481 = n2576 & n5412;
  assign n5482 = n5480 & ~n5481;
  assign n5483 = ~pi56 & ~n5482;
  assign n5484 = ~n5478 & n5483;
  assign n5485 = ~n2539 & ~n5280;
  assign n5486 = pi56 & ~n5485;
  assign n5487 = n2539 & ~n5412;
  assign n5488 = n5486 & ~n5487;
  assign n5489 = ~pi62 & ~n5488;
  assign n5490 = ~n5484 & n5489;
  assign n5491 = n3327 & ~n5490;
  assign n5492 = ~n5414 & n5491;
  assign n5493 = ~pi245 & ~n5492;
  assign n5494 = ~n5400 & n5493;
  assign po163 = n5403 | n5494;
  assign n5496 = pi215 & pi1135;
  assign n5497 = pi216 & pi279;
  assign n5498 = pi879 & ~n2442;
  assign n5499 = pi105 & ~n5498;
  assign n5500 = ~pi105 & ~pi161;
  assign n5501 = ~n5499 & ~n5500;
  assign n5502 = pi228 & n5501;
  assign n5503 = pi161 & ~pi228;
  assign n5504 = ~n5502 & ~n5503;
  assign n5505 = ~pi216 & ~n5504;
  assign n5506 = ~n5497 & ~n5505;
  assign n5507 = ~pi221 & ~n5506;
  assign n5508 = ~pi938 & n2452;
  assign n5509 = ~pi1135 & ~n2452;
  assign n5510 = pi221 & ~n5509;
  assign n5511 = ~n5508 & n5510;
  assign n5512 = ~n5507 & ~n5511;
  assign n5513 = ~pi215 & ~n5512;
  assign n5514 = ~n5496 & ~n5513;
  assign n5515 = ~n3433 & n5514;
  assign n5516 = ~n3315 & n5515;
  assign n5517 = ~pi879 & n2522;
  assign n5518 = ~n3537 & ~n5503;
  assign n5519 = ~n5517 & ~n5518;
  assign n5520 = ~n3432 & ~n5502;
  assign n5521 = ~n5519 & n5520;
  assign n5522 = ~pi216 & ~n5521;
  assign n5523 = ~n5497 & ~n5522;
  assign n5524 = ~pi221 & ~n5523;
  assign n5525 = ~n5511 & ~n5524;
  assign n5526 = ~pi215 & ~n5525;
  assign n5527 = ~n5496 & ~n5526;
  assign n5528 = n3315 & n5527;
  assign n5529 = pi62 & ~n5528;
  assign n5530 = ~n5516 & n5529;
  assign n5531 = pi223 & pi1135;
  assign n5532 = ~pi938 & n2595;
  assign n5533 = ~pi1135 & ~n2595;
  assign n5534 = pi222 & ~n5533;
  assign n5535 = ~n5532 & n5534;
  assign n5536 = pi224 & ~pi279;
  assign n5537 = ~pi879 & ~n2442;
  assign n5538 = ~pi224 & n5537;
  assign n5539 = ~pi222 & ~n5538;
  assign n5540 = ~n5536 & n5539;
  assign n5541 = ~n5535 & ~n5540;
  assign n5542 = ~pi223 & ~n5541;
  assign n5543 = ~n5531 & ~n5542;
  assign n5544 = ~pi299 & ~n5543;
  assign n5545 = pi299 & ~n5515;
  assign n5546 = ~n5544 & ~n5545;
  assign n5547 = ~n2534 & n5546;
  assign n5548 = ~n2535 & n5546;
  assign n5549 = ~n2615 & n5546;
  assign n5550 = pi299 & ~n5527;
  assign n5551 = ~n5544 & ~n5550;
  assign n5552 = n2615 & n5551;
  assign n5553 = ~n5549 & ~n5552;
  assign n5554 = n2535 & ~n5553;
  assign n5555 = pi92 & ~n5554;
  assign n5556 = ~n5548 & n5555;
  assign n5557 = pi75 & n5546;
  assign n5558 = pi87 & n5553;
  assign n5559 = pi39 & ~n5551;
  assign n5560 = ~pi299 & ~n5531;
  assign n5561 = ~n5327 & n5541;
  assign n5562 = ~pi223 & ~n5561;
  assign n5563 = n5560 & ~n5562;
  assign n5564 = pi299 & ~n5496;
  assign n5565 = n3465 & ~n5501;
  assign n5566 = ~pi216 & ~n5565;
  assign n5567 = ~pi161 & ~n3380;
  assign n5568 = pi879 & ~n5567;
  assign n5569 = pi161 & n3474;
  assign n5570 = ~pi161 & ~n3088;
  assign n5571 = ~pi879 & ~n5570;
  assign n5572 = ~n5569 & n5571;
  assign n5573 = ~pi228 & ~n5572;
  assign n5574 = ~n5568 & n5573;
  assign n5575 = n5566 & ~n5574;
  assign n5576 = ~n5497 & ~n5575;
  assign n5577 = ~pi221 & ~n5576;
  assign n5578 = ~n5511 & ~n5577;
  assign n5579 = ~pi215 & ~n5578;
  assign n5580 = n5564 & ~n5579;
  assign n5581 = ~pi39 & ~n5580;
  assign n5582 = ~n5563 & n5581;
  assign n5583 = ~pi38 & ~n5582;
  assign n5584 = ~n5559 & n5583;
  assign n5585 = pi38 & n5546;
  assign n5586 = ~pi100 & ~n5585;
  assign n5587 = ~n5584 & n5586;
  assign n5588 = ~n2532 & n5546;
  assign n5589 = pi100 & ~n5588;
  assign n5590 = ~pi879 & n3393;
  assign n5591 = pi161 & ~n5590;
  assign n5592 = ~pi152 & ~pi166;
  assign n5593 = ~n3393 & ~n5592;
  assign n5594 = ~n3391 & n5592;
  assign n5595 = pi879 & ~n5594;
  assign n5596 = ~n5593 & n5595;
  assign n5597 = ~n5591 & ~n5596;
  assign n5598 = ~pi228 & ~n5597;
  assign n5599 = n5520 & ~n5598;
  assign n5600 = ~pi216 & ~n5599;
  assign n5601 = ~n5497 & ~n5600;
  assign n5602 = ~pi221 & ~n5601;
  assign n5603 = ~n5511 & ~n5602;
  assign n5604 = ~pi215 & ~n5603;
  assign n5605 = ~n5496 & ~n5604;
  assign n5606 = pi299 & ~n5605;
  assign n5607 = ~n5544 & ~n5606;
  assign n5608 = n2532 & n5607;
  assign n5609 = n5589 & ~n5608;
  assign n5610 = ~n5587 & ~n5609;
  assign n5611 = ~pi87 & ~n5610;
  assign n5612 = ~pi75 & ~n5611;
  assign n5613 = ~n5558 & n5612;
  assign n5614 = ~pi92 & ~n5613;
  assign n5615 = ~n5557 & n5614;
  assign n5616 = n2534 & ~n5615;
  assign n5617 = ~n5556 & n5616;
  assign n5618 = ~pi55 & ~n5617;
  assign n5619 = ~n5547 & n5618;
  assign n5620 = ~n2576 & n5515;
  assign n5621 = n2576 & n5527;
  assign n5622 = pi55 & ~n5621;
  assign n5623 = ~n5620 & n5622;
  assign n5624 = ~pi56 & ~n5623;
  assign n5625 = ~n5619 & n5624;
  assign n5626 = ~n2539 & ~n5515;
  assign n5627 = pi56 & ~n5626;
  assign n5628 = n2539 & ~n5527;
  assign n5629 = n5627 & ~n5628;
  assign n5630 = ~pi62 & ~n5629;
  assign n5631 = ~n5625 & n5630;
  assign n5632 = n3327 & ~n5631;
  assign n5633 = ~n5530 & n5632;
  assign n5634 = ~n3327 & n5514;
  assign n5635 = ~n3433 & n5634;
  assign n5636 = pi244 & ~n5635;
  assign n5637 = ~n5633 & n5636;
  assign n5638 = ~n3315 & n5514;
  assign n5639 = pi62 & ~n5638;
  assign n5640 = ~n5502 & ~n5519;
  assign n5641 = ~pi216 & ~n5640;
  assign n5642 = ~n5497 & ~n5641;
  assign n5643 = ~pi221 & ~n5642;
  assign n5644 = ~n5511 & ~n5643;
  assign n5645 = ~pi215 & ~n5644;
  assign n5646 = ~n5496 & ~n5645;
  assign n5647 = n3315 & n5646;
  assign n5648 = n5639 & ~n5647;
  assign n5649 = pi299 & ~n5514;
  assign n5650 = ~n3445 & n5544;
  assign n5651 = ~n5649 & ~n5650;
  assign n5652 = ~n2534 & n5651;
  assign n5653 = ~n2535 & n5651;
  assign n5654 = ~n2615 & n5651;
  assign n5655 = pi299 & ~n5646;
  assign n5656 = ~n5650 & ~n5655;
  assign n5657 = n2615 & n5656;
  assign n5658 = ~n5654 & ~n5657;
  assign n5659 = n2535 & ~n5658;
  assign n5660 = pi92 & ~n5659;
  assign n5661 = ~n5653 & n5660;
  assign n5662 = pi75 & n5651;
  assign n5663 = pi87 & n5658;
  assign n5664 = pi39 & ~n5656;
  assign n5665 = n5327 & ~n5535;
  assign n5666 = n5542 & ~n5665;
  assign n5667 = n5560 & ~n5666;
  assign n5668 = ~pi161 & ~n3474;
  assign n5669 = pi161 & n3088;
  assign n5670 = pi879 & ~n5669;
  assign n5671 = ~n5668 & n5670;
  assign n5672 = ~pi879 & ~n3380;
  assign n5673 = pi161 & n5672;
  assign n5674 = ~pi228 & ~n5673;
  assign n5675 = ~n5671 & n5674;
  assign n5676 = ~n3859 & ~n5675;
  assign n5677 = n5566 & n5676;
  assign n5678 = ~n5497 & ~n5677;
  assign n5679 = ~pi221 & ~n5678;
  assign n5680 = ~n5511 & ~n5679;
  assign n5681 = ~pi215 & ~n5680;
  assign n5682 = n5564 & ~n5681;
  assign n5683 = ~pi39 & ~n5682;
  assign n5684 = ~n5667 & n5683;
  assign n5685 = ~pi38 & ~n5684;
  assign n5686 = ~n5664 & n5685;
  assign n5687 = pi38 & n5651;
  assign n5688 = ~pi100 & ~n5687;
  assign n5689 = ~n5686 & n5688;
  assign n5690 = ~n2532 & n5651;
  assign n5691 = pi100 & ~n5690;
  assign n5692 = ~n5502 & ~n5598;
  assign n5693 = ~pi216 & ~n5692;
  assign n5694 = ~n5497 & ~n5693;
  assign n5695 = ~pi221 & ~n5694;
  assign n5696 = ~n5511 & ~n5695;
  assign n5697 = ~pi215 & ~n5696;
  assign n5698 = ~n5496 & ~n5697;
  assign n5699 = pi299 & ~n5698;
  assign n5700 = ~n5650 & ~n5699;
  assign n5701 = n2532 & n5700;
  assign n5702 = n5691 & ~n5701;
  assign n5703 = ~n5689 & ~n5702;
  assign n5704 = ~pi87 & ~n5703;
  assign n5705 = ~pi75 & ~n5704;
  assign n5706 = ~n5663 & n5705;
  assign n5707 = ~pi92 & ~n5706;
  assign n5708 = ~n5662 & n5707;
  assign n5709 = n2534 & ~n5708;
  assign n5710 = ~n5661 & n5709;
  assign n5711 = ~pi55 & ~n5710;
  assign n5712 = ~n5652 & n5711;
  assign n5713 = ~n2576 & n5514;
  assign n5714 = pi55 & ~n5713;
  assign n5715 = n2576 & n5646;
  assign n5716 = n5714 & ~n5715;
  assign n5717 = ~pi56 & ~n5716;
  assign n5718 = ~n5712 & n5717;
  assign n5719 = ~n2539 & ~n5514;
  assign n5720 = pi56 & ~n5719;
  assign n5721 = n2539 & ~n5646;
  assign n5722 = n5720 & ~n5721;
  assign n5723 = ~pi62 & ~n5722;
  assign n5724 = ~n5718 & n5723;
  assign n5725 = n3327 & ~n5724;
  assign n5726 = ~n5648 & n5725;
  assign n5727 = ~pi244 & ~n5726;
  assign n5728 = ~n5634 & n5727;
  assign po164 = n5637 | n5728;
  assign n5730 = pi216 & pi278;
  assign n5731 = ~pi221 & ~n5730;
  assign n5732 = ~pi105 & pi152;
  assign n5733 = pi846 & ~n2442;
  assign n5734 = pi105 & n5733;
  assign n5735 = ~n5732 & ~n5734;
  assign n5736 = pi228 & ~n5735;
  assign n5737 = pi152 & ~pi228;
  assign n5738 = ~n5736 & ~n5737;
  assign n5739 = ~pi216 & ~n5738;
  assign n5740 = n5731 & ~n5739;
  assign n5741 = pi833 & ~pi930;
  assign n5742 = ~pi216 & pi221;
  assign n5743 = n5741 & n5742;
  assign n5744 = ~pi215 & pi221;
  assign n5745 = ~pi216 & n5744;
  assign n5746 = pi833 & n5745;
  assign n5747 = ~n3531 & ~n5746;
  assign n5748 = ~n5743 & ~n5747;
  assign n5749 = ~n5740 & n5748;
  assign n5750 = ~n3433 & ~n5749;
  assign n5751 = ~n3315 & ~n5750;
  assign n5752 = pi62 & ~n5751;
  assign n5753 = ~n3432 & ~n5736;
  assign n5754 = ~pi846 & n2522;
  assign n5755 = ~n3537 & ~n5737;
  assign n5756 = ~n5754 & ~n5755;
  assign n5757 = n5753 & ~n5756;
  assign n5758 = ~pi216 & ~n5757;
  assign n5759 = n5731 & ~n5758;
  assign n5760 = n5748 & ~n5759;
  assign n5761 = n3315 & n5760;
  assign n5762 = n5752 & ~n5761;
  assign n5763 = pi222 & ~pi224;
  assign n5764 = n5741 & n5763;
  assign n5765 = pi224 & pi278;
  assign n5766 = ~pi222 & ~n5765;
  assign n5767 = ~pi224 & n5733;
  assign n5768 = n5766 & ~n5767;
  assign n5769 = ~n5764 & ~n5768;
  assign n5770 = n2597 & n5769;
  assign n5771 = ~pi299 & ~n5770;
  assign n5772 = ~n3445 & n5771;
  assign n5773 = pi299 & n5750;
  assign n5774 = ~n5772 & ~n5773;
  assign n5775 = ~n2534 & n5774;
  assign n5776 = ~n2535 & n5774;
  assign n5777 = ~n2615 & n5774;
  assign n5778 = pi299 & ~n5760;
  assign n5779 = ~n5772 & ~n5778;
  assign n5780 = n2615 & n5779;
  assign n5781 = ~n5777 & ~n5780;
  assign n5782 = n2535 & ~n5781;
  assign n5783 = pi92 & ~n5782;
  assign n5784 = ~n5776 & n5783;
  assign n5785 = pi75 & n5774;
  assign n5786 = pi87 & n5781;
  assign n5787 = pi39 & ~n5779;
  assign n5788 = ~pi846 & n3087;
  assign n5789 = ~pi224 & ~n5788;
  assign n5790 = n5766 & ~n5789;
  assign n5791 = ~n5764 & ~n5790;
  assign n5792 = ~pi223 & ~pi299;
  assign n5793 = ~n2596 & n5792;
  assign n5794 = n5791 & n5793;
  assign n5795 = pi228 & ~n5732;
  assign n5796 = pi105 & ~n5788;
  assign n5797 = n5795 & ~n5796;
  assign n5798 = ~pi216 & ~n5797;
  assign n5799 = pi152 & ~n3474;
  assign n5800 = ~pi152 & n3088;
  assign n5801 = ~pi846 & ~n5800;
  assign n5802 = ~n5799 & n5801;
  assign n5803 = ~pi152 & ~n3380;
  assign n5804 = pi846 & n5803;
  assign n5805 = ~n5802 & ~n5804;
  assign n5806 = ~pi228 & ~n5805;
  assign n5807 = n5798 & ~n5806;
  assign n5808 = n5731 & ~n5807;
  assign n5809 = ~n5743 & ~n5808;
  assign n5810 = pi299 & ~n5747;
  assign n5811 = n5809 & n5810;
  assign n5812 = ~pi39 & ~n5811;
  assign n5813 = ~n5794 & n5812;
  assign n5814 = ~pi38 & ~n5813;
  assign n5815 = ~n5787 & n5814;
  assign n5816 = pi38 & n5774;
  assign n5817 = ~pi100 & ~n5816;
  assign n5818 = ~n5815 & n5817;
  assign n5819 = ~n2532 & n5774;
  assign n5820 = pi100 & ~n5819;
  assign n5821 = pi846 & ~n3399;
  assign n5822 = ~n3394 & ~n5821;
  assign n5823 = ~pi228 & ~n5822;
  assign n5824 = n5753 & ~n5823;
  assign n5825 = ~pi216 & ~n5824;
  assign n5826 = n5731 & ~n5825;
  assign n5827 = n5748 & ~n5826;
  assign n5828 = pi299 & ~n5827;
  assign n5829 = ~n5772 & ~n5828;
  assign n5830 = n2532 & n5829;
  assign n5831 = n5820 & ~n5830;
  assign n5832 = ~n5818 & ~n5831;
  assign n5833 = ~pi87 & ~n5832;
  assign n5834 = ~pi75 & ~n5833;
  assign n5835 = ~n5786 & n5834;
  assign n5836 = ~pi92 & ~n5835;
  assign n5837 = ~n5785 & n5836;
  assign n5838 = n2534 & ~n5837;
  assign n5839 = ~n5784 & n5838;
  assign n5840 = ~pi55 & ~n5839;
  assign n5841 = ~n5775 & n5840;
  assign n5842 = ~n2576 & ~n5750;
  assign n5843 = pi55 & ~n5842;
  assign n5844 = n2576 & n5760;
  assign n5845 = n5843 & ~n5844;
  assign n5846 = ~pi56 & ~n5845;
  assign n5847 = ~n5841 & n5846;
  assign n5848 = ~n2539 & n5750;
  assign n5849 = n2539 & ~n5760;
  assign n5850 = pi56 & ~n5849;
  assign n5851 = ~n5848 & n5850;
  assign n5852 = ~pi62 & ~n5851;
  assign n5853 = ~n5847 & n5852;
  assign n5854 = n3327 & ~n5853;
  assign n5855 = ~n5762 & n5854;
  assign n5856 = ~n3327 & ~n5750;
  assign n5857 = pi242 & ~n5856;
  assign n5858 = ~n5855 & n5857;
  assign n5859 = ~n3315 & n5749;
  assign n5860 = pi62 & ~n5859;
  assign n5861 = ~n5736 & ~n5756;
  assign n5862 = ~pi216 & ~n5861;
  assign n5863 = n5731 & ~n5862;
  assign n5864 = n5748 & ~n5863;
  assign n5865 = n3315 & n5864;
  assign n5866 = n5860 & ~n5865;
  assign n5867 = pi299 & ~n5749;
  assign n5868 = ~n5771 & ~n5867;
  assign n5869 = ~n2534 & n5868;
  assign n5870 = ~n2535 & n5868;
  assign n5871 = ~n2615 & n5868;
  assign n5872 = pi299 & ~n5864;
  assign n5873 = ~n5771 & ~n5872;
  assign n5874 = n2615 & n5873;
  assign n5875 = ~n5871 & ~n5874;
  assign n5876 = n2535 & ~n5875;
  assign n5877 = pi92 & ~n5876;
  assign n5878 = ~n5870 & n5877;
  assign n5879 = pi75 & n5868;
  assign n5880 = pi87 & n5875;
  assign n5881 = pi39 & ~n5873;
  assign n5882 = ~n3087 & n5795;
  assign n5883 = pi152 & n3088;
  assign n5884 = ~pi152 & ~n3474;
  assign n5885 = ~n5883 & ~n5884;
  assign n5886 = pi846 & n5885;
  assign n5887 = pi152 & ~pi846;
  assign n5888 = ~n3380 & n5887;
  assign n5889 = ~pi228 & ~n5888;
  assign n5890 = ~n5886 & n5889;
  assign n5891 = ~n5882 & ~n5890;
  assign n5892 = n5798 & n5891;
  assign n5893 = n5731 & ~n5892;
  assign n5894 = ~n5743 & ~n5893;
  assign n5895 = n5810 & n5894;
  assign n5896 = ~n3086 & n5767;
  assign n5897 = n5766 & ~n5896;
  assign n5898 = ~n5764 & n5793;
  assign n5899 = ~n5897 & n5898;
  assign n5900 = ~pi39 & ~n5899;
  assign n5901 = ~n5895 & n5900;
  assign n5902 = ~pi38 & ~n5901;
  assign n5903 = ~n5881 & n5902;
  assign n5904 = pi38 & n5868;
  assign n5905 = ~pi100 & ~n5904;
  assign n5906 = ~n5903 & n5905;
  assign n5907 = ~n2532 & n5868;
  assign n5908 = pi100 & ~n5907;
  assign n5909 = ~n5736 & ~n5823;
  assign n5910 = ~pi216 & ~n5909;
  assign n5911 = n5731 & ~n5910;
  assign n5912 = n5748 & ~n5911;
  assign n5913 = pi299 & ~n5912;
  assign n5914 = ~n5771 & ~n5913;
  assign n5915 = n2532 & n5914;
  assign n5916 = n5908 & ~n5915;
  assign n5917 = ~n5906 & ~n5916;
  assign n5918 = ~pi87 & ~n5917;
  assign n5919 = ~pi75 & ~n5918;
  assign n5920 = ~n5880 & n5919;
  assign n5921 = ~pi92 & ~n5920;
  assign n5922 = ~n5879 & n5921;
  assign n5923 = n2534 & ~n5922;
  assign n5924 = ~n5878 & n5923;
  assign n5925 = ~pi55 & ~n5924;
  assign n5926 = ~n5869 & n5925;
  assign n5927 = ~n2576 & n5749;
  assign n5928 = pi55 & ~n5927;
  assign n5929 = n2576 & n5864;
  assign n5930 = n5928 & ~n5929;
  assign n5931 = ~pi56 & ~n5930;
  assign n5932 = ~n5926 & n5931;
  assign n5933 = ~n2539 & ~n5749;
  assign n5934 = pi56 & ~n5933;
  assign n5935 = n2539 & ~n5864;
  assign n5936 = n5934 & ~n5935;
  assign n5937 = ~pi62 & ~n5936;
  assign n5938 = ~n5932 & n5937;
  assign n5939 = n3327 & ~n5938;
  assign n5940 = ~n5866 & n5939;
  assign n5941 = ~n3327 & n5749;
  assign n5942 = ~pi242 & ~n5941;
  assign n5943 = ~n5940 & n5942;
  assign n5944 = ~n5858 & ~n5943;
  assign n5945 = ~pi1134 & ~n5944;
  assign n5946 = ~n5747 & ~n5749;
  assign n5947 = ~n3433 & n5946;
  assign n5948 = ~n3315 & n5947;
  assign n5949 = ~n5743 & ~n5759;
  assign n5950 = ~pi215 & ~n5949;
  assign n5951 = n3315 & n5950;
  assign n5952 = pi62 & ~n5951;
  assign n5953 = ~n5948 & n5952;
  assign n5954 = pi299 & ~n5946;
  assign n5955 = n2597 & n5772;
  assign n5956 = ~pi299 & ~n5955;
  assign n5957 = ~n3445 & n5956;
  assign n5958 = ~n5954 & ~n5957;
  assign n5959 = ~n5774 & n5958;
  assign n5960 = ~n2534 & n5959;
  assign n5961 = ~n2535 & n5959;
  assign n5962 = ~n2615 & n5959;
  assign n5963 = pi299 & ~n5950;
  assign n5964 = ~n5956 & ~n5963;
  assign n5965 = n2615 & n5964;
  assign n5966 = ~n5962 & ~n5965;
  assign n5967 = n2535 & ~n5966;
  assign n5968 = pi92 & ~n5967;
  assign n5969 = ~n5961 & n5968;
  assign n5970 = pi75 & n5959;
  assign n5971 = pi87 & n5966;
  assign n5972 = pi39 & ~n5964;
  assign n5973 = ~n5791 & n5792;
  assign n5974 = ~pi39 & ~n5973;
  assign n5975 = ~pi215 & pi299;
  assign n5976 = ~n5809 & n5975;
  assign n5977 = n5974 & ~n5976;
  assign n5978 = ~pi38 & ~n5977;
  assign n5979 = ~n5972 & n5978;
  assign n5980 = pi38 & n5959;
  assign n5981 = ~pi100 & ~n5980;
  assign n5982 = ~n5979 & n5981;
  assign n5983 = ~n2532 & n5959;
  assign n5984 = pi100 & ~n5983;
  assign n5985 = ~n5743 & ~n5826;
  assign n5986 = ~pi215 & ~n5985;
  assign n5987 = pi299 & ~n5986;
  assign n5988 = ~n5956 & ~n5987;
  assign n5989 = n2532 & n5988;
  assign n5990 = n5984 & ~n5989;
  assign n5991 = ~n5982 & ~n5990;
  assign n5992 = ~pi87 & ~n5991;
  assign n5993 = ~pi75 & ~n5992;
  assign n5994 = ~n5971 & n5993;
  assign n5995 = ~pi92 & ~n5994;
  assign n5996 = ~n5970 & n5995;
  assign n5997 = n2534 & ~n5996;
  assign n5998 = ~n5969 & n5997;
  assign n5999 = ~pi55 & ~n5998;
  assign n6000 = ~n5960 & n5999;
  assign n6001 = ~n2576 & n5947;
  assign n6002 = n2576 & n5950;
  assign n6003 = pi55 & ~n6002;
  assign n6004 = ~n6001 & n6003;
  assign n6005 = ~pi56 & ~n6004;
  assign n6006 = ~n6000 & n6005;
  assign n6007 = ~n2539 & ~n5947;
  assign n6008 = pi56 & ~n6007;
  assign n6009 = n2539 & ~n5950;
  assign n6010 = n6008 & ~n6009;
  assign n6011 = ~pi62 & ~n6010;
  assign n6012 = ~n6006 & n6011;
  assign n6013 = n3327 & ~n6012;
  assign n6014 = ~n5953 & n6013;
  assign n6015 = ~n3327 & n5946;
  assign n6016 = ~n3433 & n6015;
  assign n6017 = pi242 & ~n6016;
  assign n6018 = ~n6014 & n6017;
  assign n6019 = ~n3315 & n5946;
  assign n6020 = pi62 & ~n6019;
  assign n6021 = ~n5743 & ~n5863;
  assign n6022 = ~pi215 & ~n6021;
  assign n6023 = n3315 & n6022;
  assign n6024 = n6020 & ~n6023;
  assign n6025 = ~n2534 & n5958;
  assign n6026 = ~n2535 & n5958;
  assign n6027 = ~n2615 & n5958;
  assign n6028 = pi299 & ~n6022;
  assign n6029 = ~n5957 & ~n6028;
  assign n6030 = n2615 & n6029;
  assign n6031 = ~n6027 & ~n6030;
  assign n6032 = n2535 & ~n6031;
  assign n6033 = pi92 & ~n6032;
  assign n6034 = ~n6026 & n6033;
  assign n6035 = pi75 & n5958;
  assign n6036 = pi87 & n6031;
  assign n6037 = pi39 & ~n6029;
  assign n6038 = n5792 & n5897;
  assign n6039 = ~n5894 & n5975;
  assign n6040 = ~n6038 & ~n6039;
  assign n6041 = n5974 & n6040;
  assign n6042 = ~pi38 & ~n6041;
  assign n6043 = ~n6037 & n6042;
  assign n6044 = pi38 & n5958;
  assign n6045 = ~pi100 & ~n6044;
  assign n6046 = ~n6043 & n6045;
  assign n6047 = ~n2532 & n5958;
  assign n6048 = pi100 & ~n6047;
  assign n6049 = ~n5743 & ~n5911;
  assign n6050 = ~pi215 & ~n6049;
  assign n6051 = pi299 & ~n6050;
  assign n6052 = ~n5957 & ~n6051;
  assign n6053 = n2532 & n6052;
  assign n6054 = n6048 & ~n6053;
  assign n6055 = ~n6046 & ~n6054;
  assign n6056 = ~pi87 & ~n6055;
  assign n6057 = ~pi75 & ~n6056;
  assign n6058 = ~n6036 & n6057;
  assign n6059 = ~pi92 & ~n6058;
  assign n6060 = ~n6035 & n6059;
  assign n6061 = n2534 & ~n6060;
  assign n6062 = ~n6034 & n6061;
  assign n6063 = ~pi55 & ~n6062;
  assign n6064 = ~n6025 & n6063;
  assign n6065 = ~n2576 & n5946;
  assign n6066 = pi55 & ~n6065;
  assign n6067 = n2576 & n6022;
  assign n6068 = n6066 & ~n6067;
  assign n6069 = ~pi56 & ~n6068;
  assign n6070 = ~n6064 & n6069;
  assign n6071 = ~n2539 & ~n5946;
  assign n6072 = pi56 & ~n6071;
  assign n6073 = n2539 & ~n6022;
  assign n6074 = n6072 & ~n6073;
  assign n6075 = ~pi62 & ~n6074;
  assign n6076 = ~n6070 & n6075;
  assign n6077 = ~n6024 & ~n6076;
  assign n6078 = n3327 & n6077;
  assign n6079 = ~pi242 & ~n6015;
  assign n6080 = ~n6078 & n6079;
  assign n6081 = pi1134 & ~n6080;
  assign n6082 = ~n6018 & n6081;
  assign po165 = ~n5945 & ~n6082;
  assign n6084 = pi57 & pi59;
  assign n6085 = n2522 & n2540;
  assign n6086 = ~n3327 & ~n6085;
  assign n6087 = ~n6084 & ~n6086;
  assign n6088 = pi57 & ~n6087;
  assign n6089 = n2512 & n2615;
  assign n6090 = ~pi54 & n2536;
  assign n6091 = n6089 & n6090;
  assign n6092 = pi74 & ~n6091;
  assign n6093 = ~pi55 & ~n6092;
  assign n6094 = ~pi54 & ~pi92;
  assign n6095 = pi87 & ~n6089;
  assign n6096 = ~pi75 & ~n6095;
  assign n6097 = ~pi39 & n2522;
  assign n6098 = ~pi38 & pi100;
  assign n6099 = n6097 & n6098;
  assign n6100 = ~pi299 & ~n2658;
  assign n6101 = pi299 & ~n2627;
  assign n6102 = ~n6100 & ~n6101;
  assign n6103 = pi146 & n6101;
  assign n6104 = pi142 & n6100;
  assign n6105 = ~n6103 & ~n6104;
  assign n6106 = ~n6102 & n6105;
  assign n6107 = n3391 & ~n6106;
  assign n6108 = ~pi41 & ~pi99;
  assign n6109 = ~pi101 & n6108;
  assign n6110 = ~pi42 & ~pi43;
  assign n6111 = ~pi52 & n6110;
  assign n6112 = ~pi113 & ~pi116;
  assign n6113 = ~pi114 & ~pi115;
  assign n6114 = n6112 & n6113;
  assign n6115 = n6111 & n6114;
  assign n6116 = n6109 & n6115;
  assign po1057 = pi44 | ~n6116;
  assign n6118 = ~pi683 & po1057;
  assign n6119 = pi129 & pi250;
  assign n6120 = pi950 & pi1092;
  assign n6121 = ~pi824 & ~pi829;
  assign n6122 = n6120 & ~n6121;
  assign po740 = ~pi1093 & n6122;
  assign n6124 = ~pi250 & ~po740;
  assign n6125 = ~n6119 & ~n6124;
  assign n6126 = ~n6118 & ~n6125;
  assign n6127 = n6106 & ~n6126;
  assign n6128 = n6106 & ~po1057;
  assign n6129 = ~n6127 & ~n6128;
  assign n6130 = ~n6107 & n6129;
  assign n6131 = n6099 & ~n6130;
  assign n6132 = ~pi39 & n2512;
  assign n6133 = pi38 & ~n6132;
  assign n6134 = ~pi100 & ~n6133;
  assign n6135 = pi58 & n2503;
  assign n6136 = ~pi90 & ~n6135;
  assign n6137 = n2706 & n2760;
  assign n6138 = n2866 & n6137;
  assign n6139 = n2772 & ~n6138;
  assign n6140 = ~n2769 & ~n6139;
  assign n6141 = ~pi108 & ~n6140;
  assign n6142 = n2768 & ~n6141;
  assign n6143 = ~n2880 & ~n6142;
  assign n6144 = n2691 & n6143;
  assign n6145 = ~n2752 & ~n6144;
  assign n6146 = ~n2759 & n6145;
  assign n6147 = ~pi47 & ~n6146;
  assign n6148 = n2692 & ~n2755;
  assign n6149 = ~n6147 & n6148;
  assign n6150 = n6136 & ~n6149;
  assign n6151 = ~n2888 & ~n6150;
  assign n6152 = ~pi93 & ~n6151;
  assign n6153 = ~pi841 & n2504;
  assign n6154 = pi93 & ~n6153;
  assign n6155 = ~n6152 & ~n6154;
  assign n6156 = ~pi35 & ~n6155;
  assign n6157 = ~pi70 & ~n6156;
  assign n6158 = ~n2717 & n6157;
  assign n6159 = ~pi51 & ~n6158;
  assign n6160 = n2743 & ~n6159;
  assign n6161 = n3065 & ~n6160;
  assign n6162 = n2740 & ~n6161;
  assign n6163 = n2738 & ~n6162;
  assign n6164 = ~pi198 & ~pi299;
  assign n6165 = ~pi210 & pi299;
  assign n6166 = ~n6164 & ~n6165;
  assign n6167 = ~n3376 & n6166;
  assign n6168 = pi32 & ~n2921;
  assign n6169 = ~n6166 & ~n6168;
  assign n6170 = ~n6167 & ~n6169;
  assign n6171 = ~n6163 & ~n6170;
  assign n6172 = ~pi95 & ~n6171;
  assign n6173 = ~n2907 & ~n6172;
  assign n6174 = ~pi39 & ~n6173;
  assign n6175 = pi835 & pi984;
  assign n6176 = ~pi252 & ~pi1001;
  assign n6177 = ~pi979 & ~n6176;
  assign n6178 = ~n6175 & n6177;
  assign n6179 = ~pi287 & n6178;
  assign n6180 = pi835 & pi950;
  assign n6181 = n6179 & n6180;
  assign n6182 = n2978 & n6181;
  assign n6183 = pi603 & ~pi642;
  assign n6184 = ~pi614 & ~pi616;
  assign n6185 = n6183 & n6184;
  assign n6186 = ~pi661 & ~pi681;
  assign n6187 = ~pi662 & n6186;
  assign n6188 = pi680 & n6187;
  assign po1101 = n6185 | n6188;
  assign n6190 = ~pi332 & ~pi468;
  assign n6191 = po1101 & ~n6190;
  assign n6192 = ~pi907 & ~pi947;
  assign n6193 = ~pi960 & ~pi963;
  assign n6194 = ~pi975 & n6193;
  assign n6195 = ~pi978 & n6194;
  assign n6196 = ~pi970 & ~pi972;
  assign n6197 = n6195 & n6196;
  assign n6198 = n6192 & n6197;
  assign n6199 = n6190 & ~n6198;
  assign n6200 = ~n6191 & ~n6199;
  assign n6201 = pi216 & ~n6200;
  assign n6202 = pi221 & n6201;
  assign n6203 = n6182 & n6202;
  assign n6204 = n2522 & ~n6203;
  assign n6205 = ~pi215 & ~n6204;
  assign n6206 = pi1092 & n6181;
  assign n6207 = pi1093 & ~n2914;
  assign n6208 = pi829 & ~n6207;
  assign n6209 = ~pi824 & ~n6208;
  assign n6210 = pi1091 & pi1093;
  assign n6211 = n2913 & n6210;
  assign n6212 = ~n6209 & ~n6211;
  assign n6213 = n6206 & n6212;
  assign n6214 = ~n6185 & ~n6190;
  assign n6215 = ~n6188 & n6214;
  assign n6216 = n6213 & ~n6215;
  assign n6217 = n2522 & ~n6216;
  assign n6218 = ~n6198 & n6217;
  assign n6219 = ~n6190 & ~n6213;
  assign n6220 = po1101 & ~n6219;
  assign n6221 = n2522 & ~n6220;
  assign n6222 = n2512 & n6190;
  assign n6223 = po1101 & n6222;
  assign n6224 = ~n6221 & ~n6223;
  assign n6225 = n6198 & ~n6224;
  assign n6226 = ~n6218 & ~n6225;
  assign n6227 = pi215 & n6226;
  assign n6228 = ~n6205 & ~n6227;
  assign n6229 = pi299 & n6228;
  assign n6230 = ~pi587 & ~pi967;
  assign n6231 = ~pi602 & n6230;
  assign n6232 = ~pi969 & n6231;
  assign n6233 = ~pi971 & ~pi977;
  assign n6234 = ~pi974 & n6233;
  assign n6235 = ~pi961 & n6234;
  assign n6236 = n6232 & n6235;
  assign n6237 = n6190 & ~n6236;
  assign n6238 = ~n6191 & ~n6237;
  assign n6239 = pi222 & ~n6238;
  assign n6240 = pi224 & n6239;
  assign n6241 = n6182 & n6240;
  assign n6242 = n2522 & ~n6241;
  assign n6243 = ~pi223 & ~n6242;
  assign n6244 = ~n6224 & n6236;
  assign n6245 = n6217 & ~n6236;
  assign n6246 = pi223 & ~n6245;
  assign n6247 = ~n6244 & n6246;
  assign n6248 = ~pi299 & ~n6247;
  assign n6249 = ~n6243 & n6248;
  assign n6250 = pi39 & ~n6249;
  assign n6251 = ~n6229 & n6250;
  assign n6252 = ~n6174 & ~n6251;
  assign n6253 = ~pi38 & ~n6252;
  assign n6254 = n6134 & ~n6253;
  assign n6255 = ~pi87 & ~n6254;
  assign n6256 = ~n6131 & n6255;
  assign n6257 = n6096 & ~n6256;
  assign n6258 = n6094 & n6257;
  assign n6259 = ~pi74 & ~n6258;
  assign n6260 = n6093 & ~n6259;
  assign n6261 = ~pi56 & ~n6260;
  assign n6262 = ~pi55 & ~pi74;
  assign n6263 = n6091 & n6262;
  assign n6264 = pi56 & ~n6263;
  assign n6265 = ~n6261 & ~n6264;
  assign n6266 = ~pi62 & ~n6265;
  assign n6267 = n3314 & n6089;
  assign n6268 = pi62 & ~n6267;
  assign n6269 = ~pi59 & ~n6268;
  assign n6270 = ~n6266 & n6269;
  assign n6271 = ~pi57 & ~n6270;
  assign po167 = ~n6088 & ~n6271;
  assign n6273 = ~pi55 & n2531;
  assign n6274 = ~pi59 & n6273;
  assign n6275 = ~pi228 & ~n6274;
  assign n6276 = pi57 & ~n6275;
  assign n6277 = ~n6188 & ~n6190;
  assign n6278 = ~pi907 & n6190;
  assign n6279 = ~n6277 & ~n6278;
  assign n6280 = ~pi228 & ~n2576;
  assign n6281 = pi30 & pi228;
  assign n6282 = ~n3537 & ~n6281;
  assign n6283 = ~n6280 & ~n6282;
  assign n6284 = n6279 & n6283;
  assign n6285 = n6276 & n6284;
  assign n6286 = n6279 & n6281;
  assign n6287 = ~n2531 & n6286;
  assign n6288 = pi55 & ~n6284;
  assign n6289 = pi299 & n6279;
  assign n6290 = ~pi602 & n6190;
  assign n6291 = ~n6277 & ~n6290;
  assign n6292 = ~pi299 & n6291;
  assign n6293 = ~n6289 & ~n6292;
  assign n6294 = n6281 & ~n6293;
  assign n6295 = ~n2573 & ~n6294;
  assign n6296 = ~n3258 & n6294;
  assign n6297 = ~pi39 & ~n6282;
  assign n6298 = ~n6293 & n6297;
  assign n6299 = n2572 & n6298;
  assign n6300 = ~n6296 & ~n6299;
  assign n6301 = n2573 & n6300;
  assign n6302 = ~n6295 & ~n6301;
  assign n6303 = pi54 & ~n6302;
  assign n6304 = pi75 & n6300;
  assign n6305 = pi87 & n6294;
  assign n6306 = n2442 & n2511;
  assign n6307 = ~pi91 & ~pi314;
  assign n6308 = n2758 & ~n2759;
  assign n6309 = pi85 & n2817;
  assign n6310 = n2470 & ~n6309;
  assign n6311 = n2821 & ~n6310;
  assign n6312 = n2471 & ~n6311;
  assign n6313 = ~n2801 & ~n2826;
  assign n6314 = ~n6312 & n6313;
  assign n6315 = n2472 & n6314;
  assign n6316 = ~n2798 & ~n6315;
  assign n6317 = n2795 & ~n6316;
  assign n6318 = pi67 & n2484;
  assign n6319 = ~n6317 & ~n6318;
  assign n6320 = n2788 & n6319;
  assign n6321 = n2787 & ~n6320;
  assign n6322 = ~pi71 & ~n6321;
  assign po1049 = pi64 | ~n2488;
  assign n6324 = n2782 & ~po1049;
  assign n6325 = ~n6322 & n6324;
  assign n6326 = ~pi81 & ~n6325;
  assign n6327 = n2836 & n6324;
  assign n6328 = n6326 & ~n6327;
  assign n6329 = ~pi102 & ~n2777;
  assign n6330 = ~pi77 & n2463;
  assign n6331 = n6329 & n6330;
  assign n6332 = ~n6328 & n6331;
  assign n6333 = n2776 & ~n6332;
  assign n6334 = n2869 & ~n6333;
  assign n6335 = n2705 & ~n6334;
  assign n6336 = ~n2708 & ~n6335;
  assign n6337 = ~pi86 & ~n6336;
  assign n6338 = n2688 & ~n2773;
  assign n6339 = ~n6337 & n6338;
  assign n6340 = n2881 & ~n6339;
  assign n6341 = n6308 & ~n6340;
  assign n6342 = n6307 & ~n6341;
  assign n6343 = ~pi91 & pi314;
  assign n6344 = ~n6326 & n6331;
  assign n6345 = n2776 & ~n6344;
  assign n6346 = n2869 & ~n6345;
  assign n6347 = n2705 & ~n6346;
  assign n6348 = ~n2708 & ~n6347;
  assign n6349 = ~pi86 & ~n6348;
  assign n6350 = n6338 & ~n6349;
  assign n6351 = n2881 & ~n6350;
  assign n6352 = n6308 & ~n6351;
  assign n6353 = n6343 & ~n6352;
  assign n6354 = ~pi58 & n2749;
  assign n6355 = ~n2692 & ~n6354;
  assign n6356 = ~n6353 & ~n6355;
  assign n6357 = ~n6342 & n6356;
  assign n6358 = ~pi90 & ~n6357;
  assign n6359 = ~n2888 & ~n6358;
  assign n6360 = ~pi93 & ~n6359;
  assign n6361 = pi93 & ~n2915;
  assign n6362 = ~pi35 & ~n6361;
  assign n6363 = ~n6360 & n6362;
  assign n6364 = ~pi70 & ~n6363;
  assign n6365 = n3078 & ~n6364;
  assign n6366 = ~pi72 & ~n6365;
  assign n6367 = ~n2739 & n3084;
  assign n6368 = ~n6366 & n6367;
  assign n6369 = ~n6306 & ~n6368;
  assign n6370 = ~pi841 & n2505;
  assign n6371 = n2508 & n6370;
  assign n6372 = n2515 & n6371;
  assign n6373 = pi32 & n6372;
  assign n6374 = ~pi95 & n6373;
  assign n6375 = ~pi198 & n6374;
  assign n6376 = n6369 & ~n6375;
  assign n6377 = ~pi228 & ~n6376;
  assign n6378 = ~n6281 & ~n6377;
  assign n6379 = n6291 & ~n6378;
  assign n6380 = ~pi299 & ~n6379;
  assign n6381 = pi180 & pi182;
  assign n6382 = pi145 & pi181;
  assign n6383 = n6381 & n6382;
  assign n6384 = ~pi299 & n6383;
  assign n6385 = ~n6380 & ~n6384;
  assign n6386 = n6281 & n6291;
  assign n6387 = ~n6190 & ~n6376;
  assign n6388 = ~pi47 & n2691;
  assign n6389 = ~n2880 & ~n6339;
  assign n6390 = n6388 & ~n6389;
  assign n6391 = n6307 & ~n6390;
  assign n6392 = ~n2880 & ~n6350;
  assign n6393 = n6388 & ~n6392;
  assign n6394 = n6343 & ~n6393;
  assign n6395 = ~n6355 & ~n6394;
  assign n6396 = ~n6391 & n6395;
  assign n6397 = ~pi90 & ~n6396;
  assign n6398 = ~n2888 & ~n6397;
  assign n6399 = ~pi93 & ~n6398;
  assign n6400 = n6362 & ~n6399;
  assign n6401 = ~pi70 & ~n6400;
  assign n6402 = n3078 & ~n6401;
  assign n6403 = ~pi72 & ~n6402;
  assign n6404 = n6367 & ~n6403;
  assign n6405 = ~n6306 & ~n6404;
  assign n6406 = ~n6375 & n6405;
  assign n6407 = n6190 & ~n6406;
  assign n6408 = ~n6387 & ~n6407;
  assign n6409 = ~pi228 & n6291;
  assign n6410 = ~n6408 & n6409;
  assign n6411 = ~n6386 & ~n6410;
  assign n6412 = n6383 & ~n6411;
  assign n6413 = ~n6385 & ~n6412;
  assign n6414 = pi299 & ~n6286;
  assign n6415 = pi158 & pi159;
  assign n6416 = pi160 & pi197;
  assign n6417 = n6415 & n6416;
  assign n6418 = ~pi210 & n6374;
  assign n6419 = n6369 & ~n6418;
  assign n6420 = ~n6190 & ~n6419;
  assign n6421 = n6405 & ~n6418;
  assign n6422 = n6190 & ~n6421;
  assign n6423 = ~n6420 & ~n6422;
  assign n6424 = n6279 & ~n6423;
  assign n6425 = n6417 & ~n6424;
  assign n6426 = n6279 & ~n6419;
  assign n6427 = ~n6417 & ~n6426;
  assign n6428 = ~pi228 & ~n6427;
  assign n6429 = ~n6425 & n6428;
  assign n6430 = n6414 & ~n6429;
  assign n6431 = pi232 & ~n6430;
  assign n6432 = ~n6413 & n6431;
  assign n6433 = ~pi228 & n6426;
  assign n6434 = n6414 & ~n6433;
  assign n6435 = ~pi232 & ~n6434;
  assign n6436 = ~n6380 & n6435;
  assign n6437 = ~n6432 & ~n6436;
  assign n6438 = ~pi39 & ~n6437;
  assign n6439 = pi222 & ~pi223;
  assign n6440 = ~pi287 & n2522;
  assign n6441 = pi835 & n6178;
  assign n6442 = n6440 & n6441;
  assign n6443 = pi824 & pi1093;
  assign n6444 = n6120 & n6443;
  assign n6445 = n6442 & n6444;
  assign n6446 = ~pi829 & ~n2913;
  assign n6447 = pi1091 & ~n6446;
  assign n6448 = n6445 & ~n6447;
  assign n6449 = ~pi224 & ~n6448;
  assign n6450 = ~pi1091 & n6445;
  assign n6451 = pi1091 & n2913;
  assign n6452 = n6444 & ~n6451;
  assign n6453 = ~n2978 & ~n6452;
  assign n6454 = pi1091 & ~n6453;
  assign n6455 = n6442 & n6454;
  assign n6456 = ~n6450 & ~n6455;
  assign n6457 = pi224 & n6456;
  assign n6458 = ~n6449 & ~n6457;
  assign n6459 = n6439 & n6458;
  assign n6460 = ~pi228 & n6459;
  assign n6461 = ~n6281 & ~n6460;
  assign n6462 = n6291 & ~n6461;
  assign n6463 = ~pi299 & ~n6462;
  assign n6464 = pi216 & ~n6456;
  assign n6465 = ~pi216 & n6448;
  assign n6466 = ~n6464 & ~n6465;
  assign n6467 = ~pi228 & ~n6466;
  assign n6468 = ~n6281 & ~n6467;
  assign n6469 = n5744 & ~n6468;
  assign n6470 = ~n6281 & ~n6469;
  assign n6471 = n6279 & ~n6470;
  assign n6472 = pi299 & ~n6471;
  assign n6473 = pi39 & ~n6472;
  assign n6474 = ~n6463 & n6473;
  assign n6475 = ~pi38 & ~n6474;
  assign n6476 = ~n6438 & n6475;
  assign n6477 = ~n6294 & ~n6298;
  assign n6478 = pi38 & n6477;
  assign n6479 = ~n6476 & ~n6478;
  assign n6480 = ~pi100 & ~n6479;
  assign n6481 = ~n2532 & n6294;
  assign n6482 = pi100 & ~n6481;
  assign n6483 = pi252 & n6222;
  assign n6484 = ~n6188 & n6483;
  assign n6485 = pi252 & n2522;
  assign n6486 = n6188 & n6485;
  assign n6487 = ~n6484 & ~n6486;
  assign n6488 = ~n2628 & n6487;
  assign n6489 = n2522 & ~n6125;
  assign n6490 = pi683 & n6489;
  assign n6491 = po1057 & n6490;
  assign n6492 = ~n6277 & n6491;
  assign n6493 = n2628 & ~n6492;
  assign n6494 = ~pi228 & ~n6493;
  assign n6495 = ~n6278 & n6494;
  assign n6496 = ~n6488 & n6495;
  assign n6497 = n6414 & ~n6496;
  assign n6498 = ~pi142 & ~n2658;
  assign n6499 = n6492 & n6498;
  assign n6500 = pi252 & ~n6498;
  assign n6501 = ~n6487 & n6500;
  assign n6502 = ~n6499 & ~n6501;
  assign n6503 = ~pi228 & ~n6290;
  assign n6504 = ~n6502 & n6503;
  assign n6505 = ~pi299 & ~n6504;
  assign n6506 = ~n6386 & n6505;
  assign n6507 = ~n6497 & ~n6506;
  assign n6508 = n2532 & n6507;
  assign n6509 = n6482 & ~n6508;
  assign n6510 = ~n6480 & ~n6509;
  assign n6511 = ~pi87 & n6510;
  assign n6512 = ~pi75 & ~n6511;
  assign n6513 = ~n6305 & n6512;
  assign n6514 = ~pi92 & ~n6513;
  assign n6515 = ~n6304 & n6514;
  assign n6516 = pi75 & ~n6294;
  assign n6517 = pi92 & ~n6516;
  assign n6518 = ~pi75 & n6300;
  assign n6519 = n6517 & ~n6518;
  assign n6520 = ~pi54 & ~n6519;
  assign n6521 = ~n6515 & n6520;
  assign n6522 = ~pi74 & ~n6521;
  assign n6523 = ~n6303 & n6522;
  assign n6524 = ~pi54 & n6301;
  assign n6525 = ~pi54 & n2573;
  assign n6526 = ~n6294 & ~n6525;
  assign n6527 = pi74 & ~n6526;
  assign n6528 = ~n6524 & n6527;
  assign n6529 = ~pi55 & ~n6528;
  assign n6530 = ~n6523 & n6529;
  assign n6531 = n2531 & ~n6530;
  assign n6532 = ~n6288 & n6531;
  assign n6533 = ~pi59 & ~n6532;
  assign n6534 = ~n6287 & n6533;
  assign n6535 = ~pi228 & ~n6273;
  assign n6536 = n6284 & ~n6535;
  assign n6537 = pi59 & ~n6536;
  assign n6538 = ~pi57 & ~n6537;
  assign n6539 = ~n6534 & n6538;
  assign po171 = ~n6285 & ~n6539;
  assign n6541 = ~pi947 & n6190;
  assign n6542 = ~n6214 & ~n6541;
  assign n6543 = n6283 & n6542;
  assign n6544 = n6276 & n6543;
  assign n6545 = n6281 & n6542;
  assign n6546 = ~n2531 & n6545;
  assign n6547 = pi55 & ~n6543;
  assign n6548 = pi299 & ~n6542;
  assign n6549 = ~pi587 & n6190;
  assign n6550 = ~n6214 & ~n6549;
  assign n6551 = ~pi299 & ~n6550;
  assign n6552 = ~n6548 & ~n6551;
  assign n6553 = n6281 & n6552;
  assign n6554 = ~n2573 & ~n6553;
  assign n6555 = ~n3258 & n6553;
  assign n6556 = n6297 & n6552;
  assign n6557 = n2572 & n6556;
  assign n6558 = ~n6555 & ~n6557;
  assign n6559 = n2573 & n6558;
  assign n6560 = ~n6554 & ~n6559;
  assign n6561 = pi54 & ~n6560;
  assign n6562 = pi75 & n6558;
  assign n6563 = pi87 & n6553;
  assign n6564 = ~n6378 & n6550;
  assign n6565 = ~n6383 & n6564;
  assign n6566 = n6281 & n6550;
  assign n6567 = ~pi228 & n6550;
  assign n6568 = ~n6408 & n6567;
  assign n6569 = ~n6566 & ~n6568;
  assign n6570 = n6383 & ~n6569;
  assign n6571 = ~pi299 & ~n6570;
  assign n6572 = ~n6565 & n6571;
  assign n6573 = pi299 & ~n6545;
  assign n6574 = ~n6423 & n6542;
  assign n6575 = n6417 & ~n6574;
  assign n6576 = ~n6419 & n6542;
  assign n6577 = ~n6417 & ~n6576;
  assign n6578 = ~pi228 & ~n6577;
  assign n6579 = ~n6575 & n6578;
  assign n6580 = n6573 & ~n6579;
  assign n6581 = pi232 & ~n6580;
  assign n6582 = ~n6572 & n6581;
  assign n6583 = ~pi299 & ~n6564;
  assign n6584 = ~pi228 & n6576;
  assign n6585 = n6573 & ~n6584;
  assign n6586 = ~pi232 & ~n6585;
  assign n6587 = ~n6583 & n6586;
  assign n6588 = ~n6582 & ~n6587;
  assign n6589 = ~pi39 & ~n6588;
  assign n6590 = ~n6461 & n6550;
  assign n6591 = ~pi299 & ~n6590;
  assign n6592 = pi299 & n5744;
  assign n6593 = ~n6573 & ~n6592;
  assign n6594 = n6469 & n6542;
  assign n6595 = ~n6593 & ~n6594;
  assign n6596 = pi39 & ~n6595;
  assign n6597 = ~n6591 & n6596;
  assign n6598 = ~pi38 & ~n6597;
  assign n6599 = ~n6589 & n6598;
  assign n6600 = ~n6553 & ~n6556;
  assign n6601 = pi38 & n6600;
  assign n6602 = ~n6599 & ~n6601;
  assign n6603 = ~pi100 & ~n6602;
  assign n6604 = ~n2532 & n6553;
  assign n6605 = pi100 & ~n6604;
  assign n6606 = ~n6214 & n6491;
  assign n6607 = n2628 & ~n6541;
  assign n6608 = n6606 & n6607;
  assign n6609 = n6185 & ~n6485;
  assign n6610 = ~n6185 & ~n6483;
  assign n6611 = ~n6609 & ~n6610;
  assign n6612 = n6185 & ~n6190;
  assign n6613 = ~pi947 & ~n6612;
  assign n6614 = ~n2628 & ~n6613;
  assign n6615 = n6611 & n6614;
  assign n6616 = ~n6608 & ~n6615;
  assign n6617 = ~pi228 & ~n6616;
  assign n6618 = n6573 & ~n6617;
  assign n6619 = ~pi228 & n2658;
  assign n6620 = ~n6549 & n6611;
  assign n6621 = n6619 & ~n6620;
  assign n6622 = ~pi142 & ~n6606;
  assign n6623 = ~pi587 & ~n6612;
  assign n6624 = pi142 & ~n6611;
  assign n6625 = ~pi228 & ~n6624;
  assign n6626 = ~n6623 & n6625;
  assign n6627 = ~n6622 & n6626;
  assign n6628 = ~n6566 & ~n6619;
  assign n6629 = ~n6627 & n6628;
  assign n6630 = ~n6621 & ~n6629;
  assign n6631 = ~pi299 & ~n6630;
  assign n6632 = ~n6618 & ~n6631;
  assign n6633 = n2532 & n6632;
  assign n6634 = n6605 & ~n6633;
  assign n6635 = ~n6603 & ~n6634;
  assign n6636 = ~pi87 & n6635;
  assign n6637 = ~pi75 & ~n6636;
  assign n6638 = ~n6563 & n6637;
  assign n6639 = ~pi92 & ~n6638;
  assign n6640 = ~n6562 & n6639;
  assign n6641 = pi75 & ~n6553;
  assign n6642 = pi92 & ~n6641;
  assign n6643 = ~pi75 & n6558;
  assign n6644 = n6642 & ~n6643;
  assign n6645 = ~pi54 & ~n6644;
  assign n6646 = ~n6640 & n6645;
  assign n6647 = ~pi74 & ~n6646;
  assign n6648 = ~n6561 & n6647;
  assign n6649 = ~pi54 & n6559;
  assign n6650 = ~n6525 & ~n6553;
  assign n6651 = pi74 & ~n6650;
  assign n6652 = ~n6649 & n6651;
  assign n6653 = ~pi55 & ~n6652;
  assign n6654 = ~n6648 & n6653;
  assign n6655 = n2531 & ~n6654;
  assign n6656 = ~n6547 & n6655;
  assign n6657 = ~pi59 & ~n6656;
  assign n6658 = ~n6546 & n6657;
  assign n6659 = ~n6535 & n6543;
  assign n6660 = pi59 & ~n6659;
  assign n6661 = ~pi57 & ~n6660;
  assign n6662 = ~n6658 & n6661;
  assign po172 = ~n6544 & ~n6662;
  assign n6664 = n6190 & n6281;
  assign n6665 = pi970 & n6664;
  assign n6666 = ~pi228 & pi970;
  assign n6667 = n2576 & n6222;
  assign n6668 = n6666 & n6667;
  assign n6669 = n6274 & n6668;
  assign n6670 = ~n6665 & ~n6669;
  assign n6671 = pi57 & ~n6670;
  assign n6672 = ~n2531 & n6665;
  assign n6673 = pi55 & ~n6665;
  assign n6674 = ~n6668 & n6673;
  assign n6675 = pi299 & pi970;
  assign n6676 = ~pi299 & pi967;
  assign n6677 = ~n6675 & ~n6676;
  assign n6678 = n6664 & ~n6677;
  assign n6679 = ~n2573 & ~n6678;
  assign n6680 = ~n3258 & n6678;
  assign n6681 = ~pi228 & ~n6222;
  assign n6682 = pi228 & ~n6664;
  assign n6683 = ~n6681 & ~n6682;
  assign n6684 = ~pi39 & ~n6677;
  assign n6685 = n6683 & n6684;
  assign n6686 = n2572 & n6685;
  assign n6687 = ~n6680 & ~n6686;
  assign n6688 = n2573 & n6687;
  assign n6689 = ~n6679 & ~n6688;
  assign n6690 = pi54 & ~n6689;
  assign n6691 = pi75 & n6687;
  assign n6692 = pi87 & n6678;
  assign n6693 = pi299 & ~n6665;
  assign n6694 = n6190 & ~n6419;
  assign n6695 = n6666 & n6694;
  assign n6696 = n6693 & ~n6695;
  assign n6697 = pi299 & n6415;
  assign n6698 = ~n6696 & ~n6697;
  assign n6699 = n6416 & ~n6422;
  assign n6700 = ~n6416 & n6419;
  assign n6701 = ~n6699 & ~n6700;
  assign n6702 = n6190 & n6701;
  assign n6703 = n6666 & n6702;
  assign n6704 = ~n6665 & ~n6703;
  assign n6705 = n6415 & ~n6704;
  assign n6706 = ~n6698 & ~n6705;
  assign n6707 = n6190 & ~n6378;
  assign n6708 = ~n6383 & ~n6707;
  assign n6709 = ~n6376 & ~n6383;
  assign n6710 = ~pi228 & n6407;
  assign n6711 = ~n6664 & ~n6710;
  assign n6712 = ~n6709 & n6711;
  assign n6713 = ~n6708 & ~n6712;
  assign n6714 = pi967 & n6713;
  assign n6715 = ~pi299 & ~n6714;
  assign n6716 = pi232 & ~n6715;
  assign n6717 = ~n6706 & n6716;
  assign n6718 = pi967 & n6707;
  assign n6719 = ~pi299 & ~n6718;
  assign n6720 = ~pi232 & ~n6696;
  assign n6721 = ~n6719 & n6720;
  assign n6722 = ~n6717 & ~n6721;
  assign n6723 = ~pi39 & ~n6722;
  assign n6724 = n5744 & ~n6466;
  assign n6725 = n6190 & n6724;
  assign n6726 = ~pi228 & ~n6725;
  assign n6727 = n6675 & ~n6726;
  assign n6728 = n6190 & n6459;
  assign n6729 = ~pi228 & ~n6728;
  assign n6730 = n6676 & ~n6729;
  assign n6731 = ~n6727 & ~n6730;
  assign n6732 = pi39 & ~n6682;
  assign n6733 = ~n6731 & n6732;
  assign n6734 = ~pi38 & ~n6733;
  assign n6735 = ~n6723 & n6734;
  assign n6736 = pi39 & n6678;
  assign n6737 = ~n6685 & ~n6736;
  assign n6738 = pi38 & n6737;
  assign n6739 = ~n6735 & ~n6738;
  assign n6740 = ~pi100 & ~n6739;
  assign n6741 = ~n2532 & n6678;
  assign n6742 = pi100 & ~n6741;
  assign n6743 = n6190 & n6491;
  assign n6744 = n2628 & ~n6743;
  assign n6745 = ~n2628 & ~n6483;
  assign n6746 = ~pi228 & ~n6745;
  assign n6747 = ~n6744 & n6746;
  assign n6748 = pi970 & n6747;
  assign n6749 = n6693 & ~n6748;
  assign n6750 = n6498 & n6743;
  assign n6751 = n6483 & ~n6498;
  assign n6752 = ~pi228 & ~n6751;
  assign n6753 = ~n6750 & n6752;
  assign n6754 = ~n6682 & ~n6753;
  assign n6755 = pi967 & n6754;
  assign n6756 = ~pi299 & ~n6755;
  assign n6757 = ~n6749 & ~n6756;
  assign n6758 = n2532 & n6757;
  assign n6759 = n6742 & ~n6758;
  assign n6760 = ~n6740 & ~n6759;
  assign n6761 = ~pi87 & n6760;
  assign n6762 = ~pi75 & ~n6761;
  assign n6763 = ~n6692 & n6762;
  assign n6764 = ~pi92 & ~n6763;
  assign n6765 = ~n6691 & n6764;
  assign n6766 = pi75 & ~n6678;
  assign n6767 = pi92 & ~n6766;
  assign n6768 = ~pi75 & n6687;
  assign n6769 = n6767 & ~n6768;
  assign n6770 = ~pi54 & ~n6769;
  assign n6771 = ~n6765 & n6770;
  assign n6772 = ~pi74 & ~n6771;
  assign n6773 = ~n6690 & n6772;
  assign n6774 = ~pi54 & n6688;
  assign n6775 = ~n6525 & ~n6678;
  assign n6776 = pi74 & ~n6775;
  assign n6777 = ~n6774 & n6776;
  assign n6778 = ~pi55 & ~n6777;
  assign n6779 = ~n6773 & n6778;
  assign n6780 = n2531 & ~n6779;
  assign n6781 = ~n6674 & n6780;
  assign n6782 = ~pi59 & ~n6781;
  assign n6783 = ~n6672 & n6782;
  assign n6784 = ~pi57 & ~n6783;
  assign n6785 = n6273 & n6668;
  assign n6786 = ~n6665 & ~n6785;
  assign n6787 = pi59 & n6786;
  assign n6788 = n6784 & ~n6787;
  assign po173 = ~n6671 & ~n6788;
  assign n6790 = pi972 & n6664;
  assign n6791 = ~pi228 & pi972;
  assign n6792 = n6667 & n6791;
  assign n6793 = n6274 & n6792;
  assign n6794 = ~n6790 & ~n6793;
  assign n6795 = pi57 & ~n6794;
  assign n6796 = ~n2531 & n6790;
  assign n6797 = pi55 & ~n6790;
  assign n6798 = ~n6792 & n6797;
  assign n6799 = ~pi299 & pi961;
  assign n6800 = pi299 & pi972;
  assign n6801 = ~n6799 & ~n6800;
  assign n6802 = n6664 & ~n6801;
  assign n6803 = ~n2573 & ~n6802;
  assign n6804 = ~n3258 & n6802;
  assign n6805 = ~pi39 & ~n6801;
  assign n6806 = n6683 & n6805;
  assign n6807 = n2572 & n6806;
  assign n6808 = ~n6804 & ~n6807;
  assign n6809 = n2573 & n6808;
  assign n6810 = ~n6803 & ~n6809;
  assign n6811 = pi54 & ~n6810;
  assign n6812 = pi75 & n6808;
  assign n6813 = pi87 & n6802;
  assign n6814 = pi299 & ~n6790;
  assign n6815 = n6694 & n6791;
  assign n6816 = n6814 & ~n6815;
  assign n6817 = ~n6697 & ~n6816;
  assign n6818 = n6702 & n6791;
  assign n6819 = ~n6790 & ~n6818;
  assign n6820 = n6415 & ~n6819;
  assign n6821 = ~n6817 & ~n6820;
  assign n6822 = pi961 & n6713;
  assign n6823 = ~pi299 & ~n6822;
  assign n6824 = pi232 & ~n6823;
  assign n6825 = ~n6821 & n6824;
  assign n6826 = pi961 & n6707;
  assign n6827 = ~pi299 & ~n6826;
  assign n6828 = ~pi232 & ~n6816;
  assign n6829 = ~n6827 & n6828;
  assign n6830 = ~n6825 & ~n6829;
  assign n6831 = ~pi39 & ~n6830;
  assign n6832 = ~n6729 & n6799;
  assign n6833 = ~n6726 & n6800;
  assign n6834 = ~n6832 & ~n6833;
  assign n6835 = n6732 & ~n6834;
  assign n6836 = ~pi38 & ~n6835;
  assign n6837 = ~n6831 & n6836;
  assign n6838 = pi39 & n6802;
  assign n6839 = ~n6806 & ~n6838;
  assign n6840 = pi38 & n6839;
  assign n6841 = ~n6837 & ~n6840;
  assign n6842 = ~pi100 & ~n6841;
  assign n6843 = ~n2532 & n6802;
  assign n6844 = pi100 & ~n6843;
  assign n6845 = pi972 & n6747;
  assign n6846 = n6814 & ~n6845;
  assign n6847 = pi961 & n6754;
  assign n6848 = ~pi299 & ~n6847;
  assign n6849 = ~n6846 & ~n6848;
  assign n6850 = n2532 & n6849;
  assign n6851 = n6844 & ~n6850;
  assign n6852 = ~n6842 & ~n6851;
  assign n6853 = ~pi87 & n6852;
  assign n6854 = ~pi75 & ~n6853;
  assign n6855 = ~n6813 & n6854;
  assign n6856 = ~pi92 & ~n6855;
  assign n6857 = ~n6812 & n6856;
  assign n6858 = pi75 & ~n6802;
  assign n6859 = pi92 & ~n6858;
  assign n6860 = ~pi75 & n6808;
  assign n6861 = n6859 & ~n6860;
  assign n6862 = ~pi54 & ~n6861;
  assign n6863 = ~n6857 & n6862;
  assign n6864 = ~pi74 & ~n6863;
  assign n6865 = ~n6811 & n6864;
  assign n6866 = ~pi54 & n6809;
  assign n6867 = ~n6525 & ~n6802;
  assign n6868 = pi74 & ~n6867;
  assign n6869 = ~n6866 & n6868;
  assign n6870 = ~pi55 & ~n6869;
  assign n6871 = ~n6865 & n6870;
  assign n6872 = n2531 & ~n6871;
  assign n6873 = ~n6798 & n6872;
  assign n6874 = ~pi59 & ~n6873;
  assign n6875 = ~n6796 & n6874;
  assign n6876 = ~pi57 & ~n6875;
  assign n6877 = n6273 & n6792;
  assign n6878 = ~n6790 & ~n6877;
  assign n6879 = pi59 & n6878;
  assign n6880 = n6876 & ~n6879;
  assign po174 = ~n6795 & ~n6880;
  assign n6882 = pi960 & n6664;
  assign n6883 = ~pi228 & pi960;
  assign n6884 = n6667 & n6883;
  assign n6885 = n6274 & n6884;
  assign n6886 = ~n6882 & ~n6885;
  assign n6887 = pi57 & ~n6886;
  assign n6888 = ~n2531 & n6882;
  assign n6889 = pi55 & ~n6882;
  assign n6890 = ~n6884 & n6889;
  assign n6891 = ~pi299 & pi977;
  assign n6892 = pi299 & pi960;
  assign n6893 = ~n6891 & ~n6892;
  assign n6894 = n6664 & ~n6893;
  assign n6895 = ~n2573 & ~n6894;
  assign n6896 = ~n3258 & n6894;
  assign n6897 = ~pi39 & ~n6893;
  assign n6898 = n6683 & n6897;
  assign n6899 = n2572 & n6898;
  assign n6900 = ~n6896 & ~n6899;
  assign n6901 = n2573 & n6900;
  assign n6902 = ~n6895 & ~n6901;
  assign n6903 = pi54 & ~n6902;
  assign n6904 = pi75 & n6900;
  assign n6905 = pi87 & n6894;
  assign n6906 = pi299 & ~n6882;
  assign n6907 = n6694 & n6883;
  assign n6908 = n6906 & ~n6907;
  assign n6909 = ~n6697 & ~n6908;
  assign n6910 = n6702 & n6883;
  assign n6911 = ~n6882 & ~n6910;
  assign n6912 = n6415 & ~n6911;
  assign n6913 = ~n6909 & ~n6912;
  assign n6914 = pi977 & n6713;
  assign n6915 = ~pi299 & ~n6914;
  assign n6916 = pi232 & ~n6915;
  assign n6917 = ~n6913 & n6916;
  assign n6918 = pi977 & n6707;
  assign n6919 = ~pi299 & ~n6918;
  assign n6920 = ~pi232 & ~n6908;
  assign n6921 = ~n6919 & n6920;
  assign n6922 = ~n6917 & ~n6921;
  assign n6923 = ~pi39 & ~n6922;
  assign n6924 = ~n6729 & n6891;
  assign n6925 = ~n6726 & n6892;
  assign n6926 = ~n6924 & ~n6925;
  assign n6927 = n6732 & ~n6926;
  assign n6928 = ~pi38 & ~n6927;
  assign n6929 = ~n6923 & n6928;
  assign n6930 = pi39 & n6894;
  assign n6931 = ~n6898 & ~n6930;
  assign n6932 = pi38 & n6931;
  assign n6933 = ~n6929 & ~n6932;
  assign n6934 = ~pi100 & ~n6933;
  assign n6935 = ~n2532 & n6894;
  assign n6936 = pi100 & ~n6935;
  assign n6937 = pi960 & n6747;
  assign n6938 = n6906 & ~n6937;
  assign n6939 = pi977 & n6754;
  assign n6940 = ~pi299 & ~n6939;
  assign n6941 = ~n6938 & ~n6940;
  assign n6942 = n2532 & n6941;
  assign n6943 = n6936 & ~n6942;
  assign n6944 = ~n6934 & ~n6943;
  assign n6945 = ~pi87 & n6944;
  assign n6946 = ~pi75 & ~n6945;
  assign n6947 = ~n6905 & n6946;
  assign n6948 = ~pi92 & ~n6947;
  assign n6949 = ~n6904 & n6948;
  assign n6950 = pi75 & ~n6894;
  assign n6951 = pi92 & ~n6950;
  assign n6952 = ~pi75 & n6900;
  assign n6953 = n6951 & ~n6952;
  assign n6954 = ~pi54 & ~n6953;
  assign n6955 = ~n6949 & n6954;
  assign n6956 = ~pi74 & ~n6955;
  assign n6957 = ~n6903 & n6956;
  assign n6958 = ~pi54 & n6901;
  assign n6959 = ~n6525 & ~n6894;
  assign n6960 = pi74 & ~n6959;
  assign n6961 = ~n6958 & n6960;
  assign n6962 = ~pi55 & ~n6961;
  assign n6963 = ~n6957 & n6962;
  assign n6964 = n2531 & ~n6963;
  assign n6965 = ~n6890 & n6964;
  assign n6966 = ~pi59 & ~n6965;
  assign n6967 = ~n6888 & n6966;
  assign n6968 = ~pi57 & ~n6967;
  assign n6969 = n6273 & n6884;
  assign n6970 = ~n6882 & ~n6969;
  assign n6971 = pi59 & n6970;
  assign n6972 = n6968 & ~n6971;
  assign po175 = ~n6887 & ~n6972;
  assign n6974 = pi963 & n6664;
  assign n6975 = ~pi228 & pi963;
  assign n6976 = n6667 & n6975;
  assign n6977 = n6274 & n6976;
  assign n6978 = ~n6974 & ~n6977;
  assign n6979 = pi57 & ~n6978;
  assign n6980 = ~n2531 & n6974;
  assign n6981 = pi55 & ~n6974;
  assign n6982 = ~n6976 & n6981;
  assign n6983 = ~pi299 & pi969;
  assign n6984 = pi299 & pi963;
  assign n6985 = ~n6983 & ~n6984;
  assign n6986 = n6664 & ~n6985;
  assign n6987 = ~n2573 & ~n6986;
  assign n6988 = ~n3258 & n6986;
  assign n6989 = ~pi39 & ~n6985;
  assign n6990 = n6683 & n6989;
  assign n6991 = n2572 & n6990;
  assign n6992 = ~n6988 & ~n6991;
  assign n6993 = n2573 & n6992;
  assign n6994 = ~n6987 & ~n6993;
  assign n6995 = pi54 & ~n6994;
  assign n6996 = pi75 & n6992;
  assign n6997 = pi87 & n6986;
  assign n6998 = pi299 & ~n6974;
  assign n6999 = n6694 & n6975;
  assign n7000 = n6998 & ~n6999;
  assign n7001 = ~n6697 & ~n7000;
  assign n7002 = n6702 & n6975;
  assign n7003 = ~n6974 & ~n7002;
  assign n7004 = n6415 & ~n7003;
  assign n7005 = ~n7001 & ~n7004;
  assign n7006 = pi969 & n6713;
  assign n7007 = ~pi299 & ~n7006;
  assign n7008 = pi232 & ~n7007;
  assign n7009 = ~n7005 & n7008;
  assign n7010 = pi969 & n6707;
  assign n7011 = ~pi299 & ~n7010;
  assign n7012 = ~pi232 & ~n7000;
  assign n7013 = ~n7011 & n7012;
  assign n7014 = ~n7009 & ~n7013;
  assign n7015 = ~pi39 & ~n7014;
  assign n7016 = ~n6729 & n6983;
  assign n7017 = ~n6726 & n6984;
  assign n7018 = ~n7016 & ~n7017;
  assign n7019 = n6732 & ~n7018;
  assign n7020 = ~pi38 & ~n7019;
  assign n7021 = ~n7015 & n7020;
  assign n7022 = pi39 & n6986;
  assign n7023 = ~n6990 & ~n7022;
  assign n7024 = pi38 & n7023;
  assign n7025 = ~n7021 & ~n7024;
  assign n7026 = ~pi100 & ~n7025;
  assign n7027 = ~n2532 & n6986;
  assign n7028 = pi100 & ~n7027;
  assign n7029 = pi963 & n6747;
  assign n7030 = n6998 & ~n7029;
  assign n7031 = pi969 & n6754;
  assign n7032 = ~pi299 & ~n7031;
  assign n7033 = ~n7030 & ~n7032;
  assign n7034 = n2532 & n7033;
  assign n7035 = n7028 & ~n7034;
  assign n7036 = ~n7026 & ~n7035;
  assign n7037 = ~pi87 & n7036;
  assign n7038 = ~pi75 & ~n7037;
  assign n7039 = ~n6997 & n7038;
  assign n7040 = ~pi92 & ~n7039;
  assign n7041 = ~n6996 & n7040;
  assign n7042 = pi75 & ~n6986;
  assign n7043 = pi92 & ~n7042;
  assign n7044 = ~pi75 & n6992;
  assign n7045 = n7043 & ~n7044;
  assign n7046 = ~pi54 & ~n7045;
  assign n7047 = ~n7041 & n7046;
  assign n7048 = ~pi74 & ~n7047;
  assign n7049 = ~n6995 & n7048;
  assign n7050 = ~pi54 & n6993;
  assign n7051 = ~n6525 & ~n6986;
  assign n7052 = pi74 & ~n7051;
  assign n7053 = ~n7050 & n7052;
  assign n7054 = ~pi55 & ~n7053;
  assign n7055 = ~n7049 & n7054;
  assign n7056 = n2531 & ~n7055;
  assign n7057 = ~n6982 & n7056;
  assign n7058 = ~pi59 & ~n7057;
  assign n7059 = ~n6980 & n7058;
  assign n7060 = ~pi57 & ~n7059;
  assign n7061 = n6273 & n6976;
  assign n7062 = ~n6974 & ~n7061;
  assign n7063 = pi59 & n7062;
  assign n7064 = n7060 & ~n7063;
  assign po176 = ~n6979 & ~n7064;
  assign n7066 = pi975 & n6664;
  assign n7067 = ~pi228 & pi975;
  assign n7068 = n6667 & n7067;
  assign n7069 = n6274 & n7068;
  assign n7070 = ~n7066 & ~n7069;
  assign n7071 = pi57 & ~n7070;
  assign n7072 = ~n2531 & n7066;
  assign n7073 = pi55 & ~n7066;
  assign n7074 = ~n7068 & n7073;
  assign n7075 = ~pi299 & pi971;
  assign n7076 = pi299 & pi975;
  assign n7077 = ~n7075 & ~n7076;
  assign n7078 = n6664 & ~n7077;
  assign n7079 = ~n2573 & ~n7078;
  assign n7080 = ~n3258 & n7078;
  assign n7081 = ~pi39 & ~n7077;
  assign n7082 = n6683 & n7081;
  assign n7083 = n2572 & n7082;
  assign n7084 = ~n7080 & ~n7083;
  assign n7085 = n2573 & n7084;
  assign n7086 = ~n7079 & ~n7085;
  assign n7087 = pi54 & ~n7086;
  assign n7088 = pi75 & n7084;
  assign n7089 = pi87 & n7078;
  assign n7090 = pi299 & ~n7066;
  assign n7091 = n6694 & n7067;
  assign n7092 = n7090 & ~n7091;
  assign n7093 = ~n6697 & ~n7092;
  assign n7094 = n6702 & n7067;
  assign n7095 = ~n7066 & ~n7094;
  assign n7096 = n6415 & ~n7095;
  assign n7097 = ~n7093 & ~n7096;
  assign n7098 = pi971 & n6713;
  assign n7099 = ~pi299 & ~n7098;
  assign n7100 = pi232 & ~n7099;
  assign n7101 = ~n7097 & n7100;
  assign n7102 = pi971 & n6707;
  assign n7103 = ~pi299 & ~n7102;
  assign n7104 = ~pi232 & ~n7092;
  assign n7105 = ~n7103 & n7104;
  assign n7106 = ~n7101 & ~n7105;
  assign n7107 = ~pi39 & ~n7106;
  assign n7108 = ~n6729 & n7075;
  assign n7109 = ~n6726 & n7076;
  assign n7110 = ~n7108 & ~n7109;
  assign n7111 = n6732 & ~n7110;
  assign n7112 = ~pi38 & ~n7111;
  assign n7113 = ~n7107 & n7112;
  assign n7114 = pi39 & n7078;
  assign n7115 = ~n7082 & ~n7114;
  assign n7116 = pi38 & n7115;
  assign n7117 = ~n7113 & ~n7116;
  assign n7118 = ~pi100 & ~n7117;
  assign n7119 = ~n2532 & n7078;
  assign n7120 = pi100 & ~n7119;
  assign n7121 = pi975 & n6747;
  assign n7122 = n7090 & ~n7121;
  assign n7123 = pi971 & n6754;
  assign n7124 = ~pi299 & ~n7123;
  assign n7125 = ~n7122 & ~n7124;
  assign n7126 = n2532 & n7125;
  assign n7127 = n7120 & ~n7126;
  assign n7128 = ~n7118 & ~n7127;
  assign n7129 = ~pi87 & n7128;
  assign n7130 = ~pi75 & ~n7129;
  assign n7131 = ~n7089 & n7130;
  assign n7132 = ~pi92 & ~n7131;
  assign n7133 = ~n7088 & n7132;
  assign n7134 = pi75 & ~n7078;
  assign n7135 = pi92 & ~n7134;
  assign n7136 = ~pi75 & n7084;
  assign n7137 = n7135 & ~n7136;
  assign n7138 = ~pi54 & ~n7137;
  assign n7139 = ~n7133 & n7138;
  assign n7140 = ~pi74 & ~n7139;
  assign n7141 = ~n7087 & n7140;
  assign n7142 = ~pi54 & n7085;
  assign n7143 = ~n6525 & ~n7078;
  assign n7144 = pi74 & ~n7143;
  assign n7145 = ~n7142 & n7144;
  assign n7146 = ~pi55 & ~n7145;
  assign n7147 = ~n7141 & n7146;
  assign n7148 = n2531 & ~n7147;
  assign n7149 = ~n7074 & n7148;
  assign n7150 = ~pi59 & ~n7149;
  assign n7151 = ~n7072 & n7150;
  assign n7152 = ~pi57 & ~n7151;
  assign n7153 = n6273 & n7068;
  assign n7154 = ~n7066 & ~n7153;
  assign n7155 = pi59 & n7154;
  assign n7156 = n7152 & ~n7155;
  assign po177 = ~n7071 & ~n7156;
  assign n7158 = pi978 & n6664;
  assign n7159 = ~pi228 & pi978;
  assign n7160 = n6667 & n7159;
  assign n7161 = n6274 & n7160;
  assign n7162 = ~n7158 & ~n7161;
  assign n7163 = pi57 & ~n7162;
  assign n7164 = ~n2531 & n7158;
  assign n7165 = pi55 & ~n7158;
  assign n7166 = ~n7160 & n7165;
  assign n7167 = ~pi299 & pi974;
  assign n7168 = pi299 & pi978;
  assign n7169 = ~n7167 & ~n7168;
  assign n7170 = n6664 & ~n7169;
  assign n7171 = ~n2573 & ~n7170;
  assign n7172 = n6683 & ~n7169;
  assign n7173 = ~pi228 & ~n3258;
  assign n7174 = n7172 & ~n7173;
  assign n7175 = n2573 & ~n7174;
  assign n7176 = ~n7171 & ~n7175;
  assign n7177 = pi54 & ~n7176;
  assign n7178 = pi75 & ~n7174;
  assign n7179 = pi87 & n7170;
  assign n7180 = ~pi39 & n7172;
  assign n7181 = pi39 & n7170;
  assign n7182 = pi38 & ~n7181;
  assign n7183 = ~n7180 & n7182;
  assign n7184 = pi299 & ~n7158;
  assign n7185 = n6694 & n7159;
  assign n7186 = n7184 & ~n7185;
  assign n7187 = ~n6697 & ~n7186;
  assign n7188 = n6702 & n7159;
  assign n7189 = ~n7158 & ~n7188;
  assign n7190 = n6415 & ~n7189;
  assign n7191 = ~n7187 & ~n7190;
  assign n7192 = pi974 & n6713;
  assign n7193 = ~pi299 & ~n7192;
  assign n7194 = pi232 & ~n7193;
  assign n7195 = ~n7191 & n7194;
  assign n7196 = pi974 & n6707;
  assign n7197 = ~pi299 & ~n7196;
  assign n7198 = ~pi232 & ~n7186;
  assign n7199 = ~n7197 & n7198;
  assign n7200 = ~n7195 & ~n7199;
  assign n7201 = ~pi39 & ~n7200;
  assign n7202 = ~n6729 & n7167;
  assign n7203 = ~n6726 & n7168;
  assign n7204 = ~n7202 & ~n7203;
  assign n7205 = n6732 & ~n7204;
  assign n7206 = ~pi38 & ~n7205;
  assign n7207 = ~n7201 & n7206;
  assign n7208 = ~n7183 & ~n7207;
  assign n7209 = ~pi100 & ~n7208;
  assign n7210 = ~n2532 & n7170;
  assign n7211 = pi100 & ~n7210;
  assign n7212 = pi978 & n6747;
  assign n7213 = n7184 & ~n7212;
  assign n7214 = pi974 & n6754;
  assign n7215 = ~pi299 & ~n7214;
  assign n7216 = ~n7213 & ~n7215;
  assign n7217 = n2532 & n7216;
  assign n7218 = n7211 & ~n7217;
  assign n7219 = ~n7209 & ~n7218;
  assign n7220 = ~pi87 & n7219;
  assign n7221 = ~pi75 & ~n7220;
  assign n7222 = ~n7179 & n7221;
  assign n7223 = ~pi92 & ~n7222;
  assign n7224 = ~n7178 & n7223;
  assign n7225 = pi75 & ~n7170;
  assign n7226 = ~pi75 & ~n7174;
  assign n7227 = pi92 & ~n7226;
  assign n7228 = ~n7225 & n7227;
  assign n7229 = ~pi54 & ~n7228;
  assign n7230 = ~n7224 & n7229;
  assign n7231 = ~pi74 & ~n7230;
  assign n7232 = ~n7177 & n7231;
  assign n7233 = ~pi54 & n7175;
  assign n7234 = ~n6525 & ~n7170;
  assign n7235 = pi74 & ~n7234;
  assign n7236 = ~n7233 & n7235;
  assign n7237 = ~pi55 & ~n7236;
  assign n7238 = ~n7232 & n7237;
  assign n7239 = n2531 & ~n7238;
  assign n7240 = ~n7166 & n7239;
  assign n7241 = ~pi59 & ~n7240;
  assign n7242 = ~n7164 & n7241;
  assign n7243 = ~pi57 & ~n7242;
  assign n7244 = n6273 & n7160;
  assign n7245 = ~n7158 & ~n7244;
  assign n7246 = pi59 & n7245;
  assign n7247 = n7243 & ~n7246;
  assign po178 = ~n7163 & ~n7247;
  assign n7249 = ~pi74 & n6091;
  assign n7250 = pi55 & ~n7249;
  assign n7251 = ~n6092 & ~n7250;
  assign n7252 = n2572 & n6097;
  assign n7253 = pi75 & ~n7252;
  assign n7254 = ~pi38 & ~pi87;
  assign n7255 = ~pi75 & ~pi100;
  assign n7256 = n6097 & n7255;
  assign n7257 = n7254 & n7256;
  assign n7258 = pi92 & ~n7257;
  assign n7259 = ~n7253 & ~n7258;
  assign n7260 = ~pi38 & n6097;
  assign n7261 = pi100 & ~n7260;
  assign n7262 = ~pi87 & ~n7261;
  assign n7263 = pi299 & ~n6200;
  assign n7264 = n6724 & n7263;
  assign n7265 = n5792 & n6239;
  assign n7266 = n6458 & n7265;
  assign n7267 = pi39 & ~n7266;
  assign n7268 = ~n7264 & n7267;
  assign n7269 = pi299 & n6419;
  assign n7270 = ~n6415 & n7269;
  assign n7271 = pi232 & ~n7270;
  assign n7272 = n6383 & n6407;
  assign n7273 = ~pi299 & ~n7272;
  assign n7274 = ~n6387 & n7273;
  assign n7275 = ~n6709 & n7274;
  assign n7276 = n7271 & ~n7275;
  assign n7277 = ~n6420 & ~n6701;
  assign n7278 = n6697 & n7277;
  assign n7279 = n7276 & ~n7278;
  assign n7280 = ~pi39 & ~n7279;
  assign n7281 = ~pi299 & n6376;
  assign n7282 = ~pi232 & ~n7281;
  assign n7283 = ~n7269 & n7282;
  assign n7284 = n7280 & ~n7283;
  assign n7285 = ~n7268 & ~n7284;
  assign n7286 = ~pi38 & ~n7285;
  assign n7287 = ~n6133 & ~n7286;
  assign n7288 = ~pi100 & ~n7287;
  assign n7289 = ~n6131 & ~n7288;
  assign n7290 = n7262 & n7289;
  assign n7291 = n2573 & ~n7290;
  assign n7292 = n7259 & ~n7291;
  assign n7293 = ~pi54 & ~n7292;
  assign n7294 = ~pi92 & n7257;
  assign n7295 = pi54 & ~n7294;
  assign n7296 = ~n7293 & ~n7295;
  assign n7297 = ~pi74 & ~n7296;
  assign n7298 = ~pi55 & n7297;
  assign n7299 = n7251 & ~n7298;
  assign n7300 = n2531 & n7299;
  assign n7301 = n3327 & ~n7300;
  assign po195 = n6087 & ~n7301;
  assign n7303 = ~pi954 & ~po195;
  assign n7304 = pi24 & pi954;
  assign po182 = ~n7303 & ~n7304;
  assign n7306 = n3315 & n3537;
  assign n7307 = ~n2441 & ~n7306;
  assign n7308 = pi62 & ~n7307;
  assign n7309 = n2534 & n2573;
  assign n7310 = n2532 & n3537;
  assign n7311 = n2571 & n7310;
  assign n7312 = n7309 & n7311;
  assign n7313 = ~n2441 & ~n7312;
  assign n7314 = pi55 & ~n7313;
  assign n7315 = ~n2441 & ~n2534;
  assign n7316 = ~pi75 & n7311;
  assign n7317 = ~n2441 & ~n7316;
  assign n7318 = pi92 & ~n7317;
  assign n7319 = pi75 & ~n2441;
  assign n7320 = n2533 & n3537;
  assign n7321 = ~n2441 & ~n7320;
  assign n7322 = pi87 & ~n7321;
  assign n7323 = ~pi100 & n4686;
  assign n7324 = ~pi39 & ~n7323;
  assign n7325 = n2522 & ~n6500;
  assign n7326 = ~pi299 & ~n7325;
  assign n7327 = pi299 & ~n3400;
  assign n7328 = ~n7326 & ~n7327;
  assign n7329 = pi100 & n7328;
  assign n7330 = n3537 & n7329;
  assign n7331 = n7324 & ~n7330;
  assign n7332 = ~pi100 & n3537;
  assign n7333 = pi39 & ~n7332;
  assign n7334 = ~pi38 & ~n7333;
  assign n7335 = ~n7331 & n7334;
  assign n7336 = ~n2441 & ~n7335;
  assign n7337 = ~pi87 & ~n7336;
  assign n7338 = ~pi75 & ~n7337;
  assign n7339 = ~n7322 & n7338;
  assign n7340 = ~pi92 & ~n7339;
  assign n7341 = ~n7319 & n7340;
  assign n7342 = n2534 & ~n7341;
  assign n7343 = ~n7318 & n7342;
  assign n7344 = ~pi55 & ~n7343;
  assign n7345 = ~n7315 & n7344;
  assign n7346 = ~pi56 & ~n7345;
  assign n7347 = ~n7314 & n7346;
  assign n7348 = n2538 & n7320;
  assign n7349 = pi56 & ~n2441;
  assign n7350 = ~n7348 & n7349;
  assign n7351 = ~pi62 & ~n7350;
  assign n7352 = ~n7347 & n7351;
  assign n7353 = ~n7308 & ~n7352;
  assign n7354 = n3327 & ~n7353;
  assign n7355 = n2441 & ~n3327;
  assign po183 = n7354 | n7355;
  assign n7357 = pi119 & pi1056;
  assign n7358 = ~pi228 & pi252;
  assign n7359 = ~pi119 & ~n7358;
  assign n7360 = ~pi468 & ~n7359;
  assign po184 = n7357 | ~n7360;
  assign n7362 = pi119 & pi1077;
  assign po185 = ~n7360 | n7362;
  assign n7364 = pi119 & pi1073;
  assign po186 = ~n7360 | n7364;
  assign n7366 = pi119 & pi1041;
  assign po187 = ~n7360 | n7366;
  assign n7368 = pi824 & n6120;
  assign n7369 = ~pi122 & pi1093;
  assign n7370 = n7368 & n7369;
  assign n7371 = ~pi1091 & n7370;
  assign n7372 = ~pi98 & n7371;
  assign n7373 = pi567 & n7372;
  assign n7374 = ~pi285 & ~pi286;
  assign n7375 = ~pi289 & n7374;
  assign n7376 = ~pi288 & n7375;
  assign po1038 = pi57 | ~n6274;
  assign n7378 = ~n7376 & po1038;
  assign n7379 = n7373 & n7378;
  assign n7380 = ~pi74 & n6094;
  assign n7381 = n2507 & ~n6154;
  assign n7382 = ~pi841 & n2695;
  assign n7383 = pi90 & n7382;
  assign n7384 = ~pi93 & ~n7383;
  assign n7385 = n7381 & ~n7384;
  assign n7386 = ~pi51 & ~n7385;
  assign n7387 = pi98 & n2761;
  assign n7388 = ~pi88 & n7387;
  assign n7389 = ~pi77 & n2760;
  assign n7390 = n2706 & n7389;
  assign n7391 = n7388 & n7390;
  assign n7392 = ~pi97 & ~n7391;
  assign n7393 = n2712 & ~n7392;
  assign n7394 = ~pi35 & n2696;
  assign n7395 = ~pi70 & n7394;
  assign n7396 = n7393 & n7395;
  assign n7397 = n7386 & ~n7396;
  assign n7398 = n2743 & n3085;
  assign n7399 = ~n7397 & n7398;
  assign n7400 = n6122 & n7399;
  assign n7401 = ~n2742 & ~n7397;
  assign n7402 = ~pi96 & ~n7401;
  assign n7403 = ~pi122 & pi829;
  assign n7404 = n6120 & n7403;
  assign n7405 = ~n7402 & n7404;
  assign n7406 = pi96 & ~n6371;
  assign n7407 = n3085 & ~n7406;
  assign n7408 = n7405 & n7407;
  assign n7409 = ~n7400 & ~n7408;
  assign n7410 = ~pi1093 & ~n7409;
  assign n7411 = ~pi87 & ~n7410;
  assign n7412 = n2522 & n6122;
  assign n7413 = ~pi1093 & n7412;
  assign n7414 = pi87 & ~n7413;
  assign n7415 = ~pi75 & n2533;
  assign n7416 = ~n7414 & n7415;
  assign n7417 = ~n7411 & n7416;
  assign n7418 = ~pi567 & ~n7417;
  assign n7419 = n7380 & ~n7418;
  assign n7420 = pi232 & n6190;
  assign n7421 = n6102 & n7420;
  assign n7422 = n3258 & ~n7421;
  assign n7423 = ~pi24 & n6485;
  assign n7424 = ~n2913 & po1057;
  assign n7425 = pi1091 & n7424;
  assign n7426 = n7404 & n7425;
  assign n7427 = n7423 & n7426;
  assign n7428 = pi1093 & n7427;
  assign n7429 = n7422 & n7428;
  assign n7430 = pi75 & ~n7429;
  assign n7431 = pi1093 & ~n2913;
  assign n7432 = ~n7386 & n7398;
  assign n7433 = n7368 & n7432;
  assign n7434 = ~pi829 & n7433;
  assign n7435 = ~pi24 & n2749;
  assign n7436 = ~pi46 & pi97;
  assign n7437 = ~pi108 & n7436;
  assign n7438 = n6388 & n7437;
  assign n7439 = n2765 & n7438;
  assign n7440 = ~pi91 & n7439;
  assign n7441 = ~n7435 & ~n7440;
  assign n7442 = n2462 & ~n7441;
  assign n7443 = n7381 & n7442;
  assign n7444 = n7386 & ~n7443;
  assign n7445 = ~n2742 & ~n7444;
  assign n7446 = ~pi96 & ~n7445;
  assign n7447 = pi829 & n6120;
  assign n7448 = n7407 & n7447;
  assign n7449 = ~n7446 & n7448;
  assign n7450 = ~n7434 & ~n7449;
  assign n7451 = ~pi122 & ~n7450;
  assign n7452 = pi122 & n6122;
  assign n7453 = n7432 & n7452;
  assign n7454 = ~n7451 & ~n7453;
  assign n7455 = n7431 & ~n7454;
  assign n7456 = pi1091 & ~n7455;
  assign n7457 = ~n7410 & n7456;
  assign n7458 = ~pi1091 & ~n7410;
  assign n7459 = ~n7457 & ~n7458;
  assign n7460 = ~pi39 & ~n7459;
  assign n7461 = n2914 & n7447;
  assign n7462 = n6442 & n7461;
  assign n7463 = pi1093 & n7462;
  assign n7464 = ~n6238 & n7463;
  assign n7465 = ~pi299 & n6439;
  assign n7466 = ~pi224 & n7465;
  assign n7467 = n7464 & n7466;
  assign n7468 = ~n6200 & n7463;
  assign n7469 = ~pi216 & n6592;
  assign n7470 = n7468 & n7469;
  assign n7471 = ~n7467 & ~n7470;
  assign n7472 = pi39 & n7471;
  assign n7473 = ~pi38 & ~n7472;
  assign n7474 = ~n7460 & n7473;
  assign n7475 = ~pi100 & ~n7474;
  assign n7476 = n6444 & n7473;
  assign n7477 = n7432 & n7476;
  assign n7478 = ~n7456 & n7477;
  assign n7479 = n7475 & ~n7478;
  assign n7480 = pi1093 & n7404;
  assign n7481 = n7424 & n7480;
  assign n7482 = n2522 & n7481;
  assign n7483 = pi1091 & n7482;
  assign n7484 = pi228 & ~n7421;
  assign n7485 = n2532 & n7484;
  assign n7486 = n7483 & n7485;
  assign n7487 = pi100 & ~n7486;
  assign n7488 = ~n7479 & ~n7487;
  assign n7489 = ~pi87 & ~n7488;
  assign n7490 = ~pi1091 & pi1093;
  assign n7491 = n2522 & n7368;
  assign n7492 = n7490 & ~n7491;
  assign n7493 = pi1093 & n2913;
  assign n7494 = n7412 & ~n7493;
  assign n7495 = ~n7490 & ~n7494;
  assign n7496 = n2615 & ~n7495;
  assign n7497 = ~n7492 & n7496;
  assign n7498 = pi87 & ~n7497;
  assign n7499 = ~n7489 & ~n7498;
  assign n7500 = ~pi75 & ~n7499;
  assign n7501 = ~n7430 & ~n7500;
  assign n7502 = pi567 & ~n7501;
  assign n7503 = n7419 & ~n7502;
  assign n7504 = n7376 & ~n7503;
  assign n7505 = ~po1038 & ~n7504;
  assign n7506 = n7423 & n7481;
  assign n7507 = pi1091 & ~n7506;
  assign n7508 = n7422 & ~n7507;
  assign n7509 = ~pi98 & n7368;
  assign n7510 = ~pi122 & n7509;
  assign n7511 = pi1093 & n7510;
  assign n7512 = ~pi1091 & ~n7511;
  assign n7513 = n7508 & ~n7512;
  assign n7514 = pi75 & ~n7513;
  assign n7515 = n7372 & ~n7422;
  assign n7516 = n7514 & ~n7515;
  assign n7517 = pi1091 & ~n7482;
  assign n7518 = ~n7512 & ~n7517;
  assign n7519 = n7485 & n7518;
  assign n7520 = n7372 & ~n7485;
  assign n7521 = pi100 & ~n7520;
  assign n7522 = ~n7519 & n7521;
  assign n7523 = ~pi39 & ~n7457;
  assign n7524 = pi122 & n7433;
  assign n7525 = ~n7510 & ~n7524;
  assign n7526 = pi1093 & ~n7525;
  assign n7527 = n7458 & ~n7526;
  assign n7528 = n7523 & ~n7527;
  assign n7529 = ~pi223 & n5763;
  assign n7530 = n7371 & ~n7529;
  assign n7531 = ~pi98 & n7530;
  assign n7532 = ~n6191 & ~n7372;
  assign n7533 = ~n2913 & n2935;
  assign n7534 = n6442 & n7533;
  assign n7535 = n2934 & n7534;
  assign n7536 = pi1091 & ~n7535;
  assign n7537 = ~n7512 & ~n7536;
  assign n7538 = n6191 & ~n7537;
  assign n7539 = ~n7532 & ~n7538;
  assign n7540 = n6236 & ~n7539;
  assign n7541 = ~n6215 & n7537;
  assign n7542 = n6215 & n7372;
  assign n7543 = ~n7541 & ~n7542;
  assign n7544 = ~n6236 & n7543;
  assign n7545 = ~n7540 & ~n7544;
  assign n7546 = n7529 & n7545;
  assign n7547 = ~pi299 & ~n7546;
  assign n7548 = ~n7531 & n7547;
  assign n7549 = n6198 & ~n7539;
  assign n7550 = ~n6198 & n7543;
  assign n7551 = ~n7549 & ~n7550;
  assign n7552 = n5745 & n7551;
  assign n7553 = ~n5745 & n7372;
  assign n7554 = pi299 & ~n7553;
  assign n7555 = ~n7552 & n7554;
  assign n7556 = pi39 & ~n7555;
  assign n7557 = ~n7548 & n7556;
  assign n7558 = ~n7528 & ~n7557;
  assign n7559 = ~pi38 & ~n7558;
  assign n7560 = pi38 & n7371;
  assign n7561 = ~pi98 & n7560;
  assign n7562 = ~pi100 & ~n7561;
  assign n7563 = ~n7559 & n7562;
  assign n7564 = ~n7522 & ~n7563;
  assign n7565 = ~pi87 & n7564;
  assign n7566 = ~pi1091 & ~n7413;
  assign n7567 = pi122 & n7491;
  assign n7568 = ~n7510 & ~n7567;
  assign n7569 = pi1093 & ~n7568;
  assign n7570 = n7566 & ~n7569;
  assign n7571 = pi1091 & ~n7494;
  assign n7572 = n2615 & ~n7571;
  assign n7573 = ~n7570 & n7572;
  assign n7574 = ~n7372 & ~n7573;
  assign n7575 = pi87 & ~n7574;
  assign n7576 = ~pi75 & ~n7575;
  assign n7577 = ~n7565 & n7576;
  assign n7578 = ~n7516 & ~n7577;
  assign n7579 = pi567 & ~n7578;
  assign n7580 = n7419 & ~n7579;
  assign n7581 = n7373 & ~n7380;
  assign n7582 = ~n7580 & ~n7581;
  assign n7583 = ~n7376 & n7582;
  assign n7584 = n7505 & ~n7583;
  assign n7585 = pi217 & ~n7584;
  assign n7586 = ~n7379 & n7585;
  assign n7587 = ~pi1161 & ~pi1162;
  assign n7588 = ~pi1163 & n7587;
  assign n7589 = ~pi351 & pi1199;
  assign n7590 = ~pi327 & ~pi362;
  assign n7591 = pi327 & pi362;
  assign n7592 = ~n7590 & ~n7591;
  assign n7593 = pi343 & ~n7592;
  assign n7594 = ~pi343 & n7592;
  assign n7595 = ~n7593 & ~n7594;
  assign n7596 = pi345 & ~pi346;
  assign n7597 = ~pi345 & pi346;
  assign n7598 = ~n7596 & ~n7597;
  assign n7599 = pi323 & ~n7598;
  assign n7600 = ~pi323 & n7598;
  assign n7601 = ~n7599 & ~n7600;
  assign n7602 = pi358 & ~n7601;
  assign n7603 = ~pi358 & n7601;
  assign n7604 = ~n7602 & ~n7603;
  assign n7605 = pi450 & n7604;
  assign n7606 = ~pi450 & ~n7604;
  assign n7607 = ~n7605 & ~n7606;
  assign n7608 = pi344 & ~n7607;
  assign n7609 = ~pi344 & n7607;
  assign n7610 = ~n7608 & ~n7609;
  assign n7611 = n7595 & ~n7610;
  assign n7612 = ~n7595 & n7610;
  assign n7613 = ~n7611 & ~n7612;
  assign n7614 = pi1197 & n7613;
  assign n7615 = pi452 & ~pi455;
  assign n7616 = ~pi452 & pi455;
  assign n7617 = ~n7615 & ~n7616;
  assign n7618 = pi320 & ~pi460;
  assign n7619 = ~pi320 & pi460;
  assign n7620 = ~n7618 & ~n7619;
  assign n7621 = pi342 & ~n7620;
  assign n7622 = ~pi342 & n7620;
  assign n7623 = ~n7621 & ~n7622;
  assign n7624 = pi361 & ~pi441;
  assign n7625 = ~pi361 & pi441;
  assign n7626 = ~n7624 & ~n7625;
  assign n7627 = n7623 & n7626;
  assign n7628 = ~n7623 & ~n7626;
  assign n7629 = ~n7627 & ~n7628;
  assign n7630 = pi355 & ~n7629;
  assign n7631 = ~pi355 & n7629;
  assign n7632 = ~n7630 & ~n7631;
  assign n7633 = pi458 & n7632;
  assign n7634 = ~pi458 & ~n7632;
  assign n7635 = ~n7633 & ~n7634;
  assign n7636 = n7617 & n7635;
  assign n7637 = ~n7617 & ~n7635;
  assign n7638 = ~n7636 & ~n7637;
  assign n7639 = ~pi592 & ~n7638;
  assign n7640 = n7373 & ~n7639;
  assign n7641 = pi1196 & ~n7640;
  assign n7642 = ~pi1198 & ~n7641;
  assign n7643 = pi1196 & ~n7638;
  assign n7644 = pi315 & ~pi359;
  assign n7645 = ~pi315 & pi359;
  assign n7646 = ~n7644 & ~n7645;
  assign n7647 = pi321 & ~pi347;
  assign n7648 = ~pi321 & pi347;
  assign n7649 = ~n7647 & ~n7648;
  assign n7650 = pi316 & ~pi349;
  assign n7651 = ~pi316 & pi349;
  assign n7652 = ~n7650 & ~n7651;
  assign n7653 = pi322 & ~pi348;
  assign n7654 = ~pi322 & pi348;
  assign n7655 = ~n7653 & ~n7654;
  assign n7656 = n7652 & n7655;
  assign n7657 = ~n7652 & ~n7655;
  assign n7658 = ~n7656 & ~n7657;
  assign n7659 = n7649 & ~n7658;
  assign n7660 = ~n7649 & n7658;
  assign n7661 = ~n7659 & ~n7660;
  assign n7662 = n7646 & n7661;
  assign n7663 = ~n7646 & ~n7661;
  assign n7664 = ~n7662 & ~n7663;
  assign n7665 = ~pi350 & ~n7664;
  assign n7666 = pi350 & n7664;
  assign n7667 = ~n7665 & ~n7666;
  assign n7668 = ~n7643 & n7667;
  assign n7669 = ~pi592 & n7373;
  assign n7670 = pi1198 & n7669;
  assign n7671 = n7668 & n7670;
  assign n7672 = ~n7642 & ~n7671;
  assign n7673 = ~n7614 & ~n7672;
  assign n7674 = ~pi592 & ~n7673;
  assign n7675 = n7373 & ~n7674;
  assign n7676 = ~n7589 & ~n7675;
  assign n7677 = pi592 & n7373;
  assign n7678 = pi1199 & ~n7677;
  assign n7679 = ~pi351 & n7678;
  assign n7680 = ~n7676 & ~n7679;
  assign n7681 = ~pi461 & n7680;
  assign n7682 = pi360 & ~pi462;
  assign n7683 = ~pi360 & pi462;
  assign n7684 = ~n7682 & ~n7683;
  assign n7685 = pi352 & ~pi353;
  assign n7686 = ~pi352 & pi353;
  assign n7687 = ~n7685 & ~n7686;
  assign n7688 = n7684 & n7687;
  assign n7689 = ~n7684 & ~n7687;
  assign n7690 = ~n7688 & ~n7689;
  assign n7691 = pi354 & n7690;
  assign n7692 = ~pi354 & ~n7690;
  assign n7693 = ~n7691 & ~n7692;
  assign n7694 = pi356 & ~pi357;
  assign n7695 = ~pi356 & pi357;
  assign n7696 = ~n7694 & ~n7695;
  assign n7697 = n7693 & n7696;
  assign n7698 = ~n7693 & ~n7696;
  assign n7699 = ~n7697 & ~n7698;
  assign n7700 = pi351 & pi1199;
  assign n7701 = ~n7675 & ~n7700;
  assign n7702 = pi351 & n7678;
  assign n7703 = ~n7701 & ~n7702;
  assign n7704 = pi461 & n7703;
  assign n7705 = ~n7699 & ~n7704;
  assign n7706 = ~n7681 & n7705;
  assign n7707 = ~pi461 & n7703;
  assign n7708 = n7699 & ~n7707;
  assign n7709 = pi461 & n7680;
  assign n7710 = n7708 & ~n7709;
  assign n7711 = ~n7706 & ~n7710;
  assign n7712 = pi590 & n7711;
  assign n7713 = pi380 & ~pi387;
  assign n7714 = ~pi380 & pi387;
  assign n7715 = ~n7713 & ~n7714;
  assign n7716 = ~pi363 & ~pi372;
  assign n7717 = pi363 & pi372;
  assign n7718 = ~n7716 & ~n7717;
  assign n7719 = pi386 & ~n7718;
  assign n7720 = ~pi386 & n7718;
  assign n7721 = ~n7719 & ~n7720;
  assign n7722 = pi338 & ~pi388;
  assign n7723 = ~pi338 & pi388;
  assign n7724 = ~n7722 & ~n7723;
  assign n7725 = pi337 & ~pi339;
  assign n7726 = ~pi337 & pi339;
  assign n7727 = ~n7725 & ~n7726;
  assign n7728 = n7724 & n7727;
  assign n7729 = ~n7724 & ~n7727;
  assign n7730 = ~n7728 & ~n7729;
  assign n7731 = n7721 & ~n7730;
  assign n7732 = ~n7721 & n7730;
  assign n7733 = ~n7731 & ~n7732;
  assign n7734 = n7715 & n7733;
  assign n7735 = ~n7715 & ~n7733;
  assign n7736 = ~n7734 & ~n7735;
  assign n7737 = pi1196 & ~n7736;
  assign n7738 = ~pi368 & ~pi389;
  assign n7739 = pi368 & pi389;
  assign n7740 = ~n7738 & ~n7739;
  assign n7741 = pi336 & ~pi383;
  assign n7742 = ~pi336 & pi383;
  assign n7743 = ~n7741 & ~n7742;
  assign n7744 = n7740 & ~n7743;
  assign n7745 = ~n7740 & n7743;
  assign n7746 = ~n7744 & ~n7745;
  assign n7747 = pi365 & ~pi447;
  assign n7748 = ~pi365 & pi447;
  assign n7749 = ~n7747 & ~n7748;
  assign n7750 = pi367 & ~n7749;
  assign n7751 = ~pi367 & n7749;
  assign n7752 = ~n7750 & ~n7751;
  assign n7753 = pi364 & ~pi366;
  assign n7754 = ~pi364 & pi366;
  assign n7755 = ~n7753 & ~n7754;
  assign n7756 = n7752 & ~n7755;
  assign n7757 = ~n7752 & n7755;
  assign n7758 = ~n7756 & ~n7757;
  assign n7759 = n7746 & n7758;
  assign n7760 = ~n7746 & ~n7758;
  assign n7761 = ~n7759 & ~n7760;
  assign n7762 = pi1197 & n7761;
  assign n7763 = ~n7737 & ~n7762;
  assign n7764 = pi317 & ~pi385;
  assign n7765 = ~pi317 & pi385;
  assign n7766 = ~n7764 & ~n7765;
  assign n7767 = pi379 & ~pi382;
  assign n7768 = ~pi379 & pi382;
  assign n7769 = ~n7767 & ~n7768;
  assign n7770 = pi376 & ~pi439;
  assign n7771 = ~pi376 & pi439;
  assign n7772 = ~n7770 & ~n7771;
  assign n7773 = pi378 & ~pi381;
  assign n7774 = ~pi378 & pi381;
  assign n7775 = ~n7773 & ~n7774;
  assign n7776 = n7772 & n7775;
  assign n7777 = ~n7772 & ~n7775;
  assign n7778 = ~n7776 & ~n7777;
  assign n7779 = n7769 & ~n7778;
  assign n7780 = ~n7769 & n7778;
  assign n7781 = ~n7779 & ~n7780;
  assign n7782 = n7766 & n7781;
  assign n7783 = ~n7766 & ~n7781;
  assign n7784 = ~n7782 & ~n7783;
  assign n7785 = ~pi377 & ~n7784;
  assign n7786 = pi377 & n7784;
  assign n7787 = ~n7785 & ~n7786;
  assign n7788 = n7763 & n7787;
  assign n7789 = pi592 & ~n7788;
  assign n7790 = n7373 & ~n7789;
  assign n7791 = pi1199 & ~n7790;
  assign n7792 = n7763 & ~n7791;
  assign n7793 = ~pi369 & ~pi374;
  assign n7794 = pi369 & pi374;
  assign n7795 = ~n7793 & ~n7794;
  assign n7796 = pi370 & ~pi371;
  assign n7797 = ~pi370 & pi371;
  assign n7798 = ~n7796 & ~n7797;
  assign n7799 = pi384 & ~pi442;
  assign n7800 = ~pi384 & pi442;
  assign n7801 = ~n7799 & ~n7800;
  assign n7802 = pi440 & ~n7801;
  assign n7803 = ~pi440 & n7801;
  assign n7804 = ~n7802 & ~n7803;
  assign n7805 = pi373 & ~n7804;
  assign n7806 = ~pi373 & n7804;
  assign n7807 = ~n7805 & ~n7806;
  assign n7808 = pi375 & n7807;
  assign n7809 = ~pi375 & ~n7807;
  assign n7810 = ~n7808 & ~n7809;
  assign n7811 = n7798 & n7810;
  assign n7812 = ~n7798 & ~n7810;
  assign n7813 = ~n7811 & ~n7812;
  assign n7814 = ~n7795 & ~n7813;
  assign n7815 = n7795 & n7813;
  assign n7816 = pi1198 & ~n7815;
  assign n7817 = ~n7814 & n7816;
  assign n7818 = n7792 & ~n7817;
  assign n7819 = n7677 & ~n7818;
  assign n7820 = n7373 & ~n7819;
  assign n7821 = ~pi590 & n7820;
  assign n7822 = ~pi591 & ~n7821;
  assign n7823 = ~n7712 & n7822;
  assign n7824 = pi1197 & ~n7677;
  assign n7825 = ~pi333 & n7824;
  assign n7826 = pi319 & ~pi324;
  assign n7827 = ~pi319 & pi324;
  assign n7828 = ~n7826 & ~n7827;
  assign n7829 = pi456 & ~n7828;
  assign n7830 = ~pi456 & n7828;
  assign n7831 = ~n7829 & ~n7830;
  assign n7832 = pi397 & ~pi404;
  assign n7833 = ~pi397 & pi404;
  assign n7834 = ~n7832 & ~n7833;
  assign n7835 = pi412 & ~n7834;
  assign n7836 = ~pi412 & n7834;
  assign n7837 = ~n7835 & ~n7836;
  assign n7838 = pi390 & ~pi410;
  assign n7839 = ~pi390 & pi410;
  assign n7840 = ~n7838 & ~n7839;
  assign n7841 = n7837 & ~n7840;
  assign n7842 = ~n7837 & n7840;
  assign n7843 = ~n7841 & ~n7842;
  assign n7844 = n7831 & n7843;
  assign n7845 = ~n7831 & ~n7843;
  assign n7846 = ~n7844 & ~n7845;
  assign n7847 = pi411 & n7846;
  assign n7848 = ~pi411 & ~n7846;
  assign n7849 = ~n7847 & ~n7848;
  assign n7850 = pi1196 & n7849;
  assign n7851 = pi318 & ~pi409;
  assign n7852 = ~pi318 & pi409;
  assign n7853 = ~n7851 & ~n7852;
  assign n7854 = pi325 & ~n7853;
  assign n7855 = ~pi325 & n7853;
  assign n7856 = ~n7854 & ~n7855;
  assign n7857 = ~pi403 & ~pi405;
  assign n7858 = pi403 & pi405;
  assign n7859 = ~n7857 & ~n7858;
  assign n7860 = pi401 & ~pi402;
  assign n7861 = ~pi401 & pi402;
  assign n7862 = ~n7860 & ~n7861;
  assign n7863 = pi326 & ~pi406;
  assign n7864 = ~pi326 & pi406;
  assign n7865 = ~n7863 & ~n7864;
  assign n7866 = n7862 & n7865;
  assign n7867 = ~n7862 & ~n7865;
  assign n7868 = ~n7866 & ~n7867;
  assign n7869 = n7859 & ~n7868;
  assign n7870 = ~n7859 & n7868;
  assign n7871 = ~n7869 & ~n7870;
  assign n7872 = n7856 & n7871;
  assign n7873 = ~n7856 & ~n7871;
  assign n7874 = ~n7872 & ~n7873;
  assign n7875 = n7511 & n7874;
  assign n7876 = ~pi1091 & n7875;
  assign n7877 = pi567 & n7876;
  assign n7878 = ~pi592 & n7877;
  assign n7879 = ~n7850 & n7878;
  assign n7880 = n7678 & ~n7879;
  assign n7881 = ~pi592 & pi1196;
  assign n7882 = n7511 & ~n7849;
  assign n7883 = ~pi1091 & n7882;
  assign n7884 = pi567 & n7883;
  assign n7885 = n7881 & n7884;
  assign n7886 = n7373 & ~n7881;
  assign n7887 = ~pi1199 & ~n7886;
  assign n7888 = ~n7885 & n7887;
  assign n7889 = ~n7880 & ~n7888;
  assign n7890 = pi1198 & ~n7677;
  assign n7891 = n7889 & ~n7890;
  assign n7892 = pi329 & ~pi395;
  assign n7893 = ~pi329 & pi395;
  assign n7894 = ~n7892 & ~n7893;
  assign n7895 = pi396 & ~n7894;
  assign n7896 = ~pi396 & n7894;
  assign n7897 = ~n7895 & ~n7896;
  assign n7898 = pi398 & ~pi399;
  assign n7899 = ~pi398 & pi399;
  assign n7900 = ~n7898 & ~n7899;
  assign n7901 = pi400 & ~n7900;
  assign n7902 = ~pi400 & n7900;
  assign n7903 = ~n7901 & ~n7902;
  assign n7904 = pi328 & ~pi408;
  assign n7905 = ~pi328 & pi408;
  assign n7906 = ~n7904 & ~n7905;
  assign n7907 = pi394 & ~n7906;
  assign n7908 = ~pi394 & n7906;
  assign n7909 = ~n7907 & ~n7908;
  assign n7910 = n7903 & ~n7909;
  assign n7911 = ~n7903 & n7909;
  assign n7912 = ~n7910 & ~n7911;
  assign n7913 = n7897 & n7912;
  assign n7914 = ~n7897 & ~n7912;
  assign n7915 = ~n7913 & ~n7914;
  assign n7916 = ~n7891 & ~n7915;
  assign n7917 = n7889 & ~n7916;
  assign n7918 = ~n7825 & n7917;
  assign n7919 = ~pi391 & n7918;
  assign n7920 = pi407 & ~pi463;
  assign n7921 = ~pi407 & pi463;
  assign n7922 = ~n7920 & ~n7921;
  assign n7923 = pi335 & ~pi413;
  assign n7924 = ~pi335 & pi413;
  assign n7925 = ~n7923 & ~n7924;
  assign n7926 = n7922 & n7925;
  assign n7927 = ~n7922 & ~n7925;
  assign n7928 = ~n7926 & ~n7927;
  assign n7929 = pi334 & n7928;
  assign n7930 = ~pi334 & ~n7928;
  assign n7931 = ~n7929 & ~n7930;
  assign n7932 = pi393 & ~n7931;
  assign n7933 = ~pi393 & n7931;
  assign n7934 = ~n7932 & ~n7933;
  assign n7935 = pi392 & n7934;
  assign n7936 = ~pi392 & ~n7934;
  assign n7937 = ~n7935 & ~n7936;
  assign n7938 = ~pi1197 & ~n7889;
  assign n7939 = ~n7824 & ~n7938;
  assign n7940 = pi333 & ~n7939;
  assign n7941 = ~pi333 & ~n7889;
  assign n7942 = ~n7916 & ~n7941;
  assign n7943 = ~n7940 & n7942;
  assign n7944 = pi391 & n7943;
  assign n7945 = ~n7937 & ~n7944;
  assign n7946 = ~n7919 & n7945;
  assign n7947 = ~pi391 & n7943;
  assign n7948 = n7937 & ~n7947;
  assign n7949 = pi391 & n7918;
  assign n7950 = n7948 & ~n7949;
  assign n7951 = ~pi590 & ~n7950;
  assign n7952 = ~n7946 & n7951;
  assign n7953 = pi590 & n7373;
  assign n7954 = pi591 & ~n7953;
  assign n7955 = ~n7952 & n7954;
  assign n7956 = ~n7823 & ~n7955;
  assign n7957 = ~pi588 & ~n7956;
  assign n7958 = ~pi590 & ~pi591;
  assign n7959 = n7373 & ~n7958;
  assign n7960 = pi588 & ~n7959;
  assign n7961 = pi416 & ~pi438;
  assign n7962 = ~pi416 & pi438;
  assign n7963 = ~n7961 & ~n7962;
  assign n7964 = pi415 & ~pi431;
  assign n7965 = ~pi415 & pi431;
  assign n7966 = ~n7964 & ~n7965;
  assign n7967 = pi437 & ~pi453;
  assign n7968 = ~pi437 & pi453;
  assign n7969 = ~n7967 & ~n7968;
  assign n7970 = ~pi417 & ~pi418;
  assign n7971 = pi417 & pi418;
  assign n7972 = ~n7970 & ~n7971;
  assign n7973 = pi464 & ~n7972;
  assign n7974 = ~pi464 & n7972;
  assign n7975 = ~n7973 & ~n7974;
  assign n7976 = n7969 & n7975;
  assign n7977 = ~n7969 & ~n7975;
  assign n7978 = ~n7976 & ~n7977;
  assign n7979 = n7966 & ~n7978;
  assign n7980 = ~n7966 & n7978;
  assign n7981 = ~n7979 & ~n7980;
  assign n7982 = n7963 & ~n7981;
  assign n7983 = ~n7963 & n7981;
  assign n7984 = ~n7982 & ~n7983;
  assign n7985 = pi1197 & n7984;
  assign n7986 = ~pi419 & ~pi420;
  assign n7987 = pi419 & pi420;
  assign n7988 = ~n7986 & ~n7987;
  assign n7989 = pi459 & ~n7988;
  assign n7990 = ~pi459 & n7988;
  assign n7991 = ~n7989 & ~n7990;
  assign n7992 = pi423 & ~pi424;
  assign n7993 = ~pi423 & pi424;
  assign n7994 = ~n7992 & ~n7993;
  assign n7995 = pi421 & ~pi454;
  assign n7996 = ~pi421 & pi454;
  assign n7997 = ~n7995 & ~n7996;
  assign n7998 = pi432 & ~n7997;
  assign n7999 = ~pi432 & n7997;
  assign n8000 = ~n7998 & ~n7999;
  assign n8001 = n7994 & ~n8000;
  assign n8002 = ~n7994 & n8000;
  assign n8003 = ~n8001 & ~n8002;
  assign n8004 = pi425 & ~n8003;
  assign n8005 = ~pi425 & n8003;
  assign n8006 = ~n8004 & ~n8005;
  assign n8007 = n7991 & n8006;
  assign n8008 = ~n7991 & ~n8006;
  assign n8009 = ~n8007 & ~n8008;
  assign n8010 = pi1198 & n8009;
  assign n8011 = ~n7985 & ~n8010;
  assign n8012 = pi436 & ~pi443;
  assign n8013 = ~pi436 & pi443;
  assign n8014 = ~n8012 & ~n8013;
  assign n8015 = ~pi444 & n8014;
  assign n8016 = pi444 & ~n8014;
  assign n8017 = ~n8015 & ~n8016;
  assign n8018 = pi434 & ~pi446;
  assign n8019 = ~pi434 & pi446;
  assign n8020 = ~n8018 & ~n8019;
  assign n8021 = pi414 & ~pi422;
  assign n8022 = ~pi414 & pi422;
  assign n8023 = ~n8021 & ~n8022;
  assign n8024 = n8020 & n8023;
  assign n8025 = ~n8020 & ~n8023;
  assign n8026 = ~n8024 & ~n8025;
  assign n8027 = pi429 & ~n8026;
  assign n8028 = ~pi429 & n8026;
  assign n8029 = ~n8027 & ~n8028;
  assign n8030 = pi435 & n8029;
  assign n8031 = ~pi435 & ~n8029;
  assign n8032 = ~n8030 & ~n8031;
  assign n8033 = n8017 & ~n8032;
  assign n8034 = ~n8017 & n8032;
  assign n8035 = n7881 & ~n8034;
  assign n8036 = ~n8033 & n8035;
  assign n8037 = n8011 & ~n8036;
  assign n8038 = n7669 & n8037;
  assign n8039 = ~pi1199 & ~n8038;
  assign n8040 = ~n7677 & n8039;
  assign n8041 = pi433 & ~pi451;
  assign n8042 = ~pi433 & pi451;
  assign n8043 = ~n8041 & ~n8042;
  assign n8044 = pi449 & n8043;
  assign n8045 = ~pi449 & ~n8043;
  assign n8046 = ~n8044 & ~n8045;
  assign n8047 = pi426 & ~pi430;
  assign n8048 = ~pi426 & pi430;
  assign n8049 = ~n8047 & ~n8048;
  assign n8050 = ~pi427 & pi428;
  assign n8051 = pi427 & ~pi428;
  assign n8052 = ~n8050 & ~n8051;
  assign n8053 = pi445 & ~n8052;
  assign n8054 = ~pi445 & n8052;
  assign n8055 = ~n8053 & ~n8054;
  assign n8056 = pi448 & ~n8055;
  assign n8057 = ~pi448 & n8055;
  assign n8058 = ~n8056 & ~n8057;
  assign n8059 = n8049 & n8058;
  assign n8060 = ~n8049 & ~n8058;
  assign n8061 = ~n8059 & ~n8060;
  assign n8062 = n8038 & ~n8061;
  assign n8063 = ~n7677 & ~n8062;
  assign n8064 = n8046 & ~n8063;
  assign n8065 = n8038 & n8061;
  assign n8066 = ~n7677 & ~n8065;
  assign n8067 = ~n8046 & ~n8066;
  assign n8068 = ~n8064 & ~n8067;
  assign n8069 = pi1199 & n8068;
  assign n8070 = ~n8040 & ~n8069;
  assign n8071 = n7958 & n8070;
  assign n8072 = n7960 & ~n8071;
  assign n8073 = n7378 & ~n8072;
  assign n8074 = ~n7957 & n8073;
  assign n8075 = ~pi87 & ~n7487;
  assign n8076 = ~n7475 & n8075;
  assign n8077 = ~n7566 & n7572;
  assign n8078 = pi87 & n8077;
  assign n8079 = ~pi75 & ~n8078;
  assign n8080 = ~n8076 & n8079;
  assign n8081 = ~n7430 & ~n8080;
  assign n8082 = pi567 & ~n8081;
  assign n8083 = n7419 & ~n8082;
  assign n8084 = ~pi592 & ~n8083;
  assign n8085 = pi592 & ~n7503;
  assign n8086 = ~n8084 & ~n8085;
  assign n8087 = ~n8011 & n8086;
  assign n8088 = ~pi1196 & ~n7503;
  assign n8089 = ~pi443 & ~pi592;
  assign n8090 = ~n7503 & ~n8089;
  assign n8091 = ~n8083 & n8089;
  assign n8092 = ~n8090 & ~n8091;
  assign n8093 = ~pi444 & ~n8092;
  assign n8094 = pi443 & ~pi592;
  assign n8095 = ~n7503 & ~n8094;
  assign n8096 = ~n8083 & n8094;
  assign n8097 = ~n8095 & ~n8096;
  assign n8098 = pi444 & ~n8097;
  assign n8099 = ~n8093 & ~n8098;
  assign n8100 = pi436 & ~n8099;
  assign n8101 = ~pi444 & ~n8097;
  assign n8102 = pi444 & ~n8092;
  assign n8103 = ~n8101 & ~n8102;
  assign n8104 = ~pi436 & ~n8103;
  assign n8105 = n8032 & ~n8104;
  assign n8106 = ~n8100 & n8105;
  assign n8107 = pi436 & ~n8103;
  assign n8108 = ~pi436 & ~n8099;
  assign n8109 = ~n8032 & ~n8108;
  assign n8110 = ~n8107 & n8109;
  assign n8111 = ~n8106 & ~n8110;
  assign n8112 = pi1196 & n8111;
  assign n8113 = ~n8088 & ~n8112;
  assign n8114 = n8011 & n8113;
  assign n8115 = ~n8087 & ~n8114;
  assign n8116 = ~pi1199 & n8115;
  assign n8117 = pi448 & n8046;
  assign n8118 = ~pi448 & ~n8046;
  assign n8119 = ~n8117 & ~n8118;
  assign n8120 = pi428 & ~n8115;
  assign n8121 = ~pi428 & n8086;
  assign n8122 = ~n8120 & ~n8121;
  assign n8123 = pi427 & ~n8122;
  assign n8124 = ~pi428 & ~n8115;
  assign n8125 = pi428 & n8086;
  assign n8126 = ~n8124 & ~n8125;
  assign n8127 = ~pi427 & ~n8126;
  assign n8128 = ~n8123 & ~n8127;
  assign n8129 = pi430 & ~n8128;
  assign n8130 = ~pi427 & ~n8122;
  assign n8131 = pi427 & ~n8126;
  assign n8132 = ~n8130 & ~n8131;
  assign n8133 = ~pi430 & ~n8132;
  assign n8134 = ~n8129 & ~n8133;
  assign n8135 = pi426 & ~n8134;
  assign n8136 = pi430 & ~n8132;
  assign n8137 = ~pi430 & ~n8128;
  assign n8138 = ~n8136 & ~n8137;
  assign n8139 = ~pi426 & ~n8138;
  assign n8140 = ~n8135 & ~n8139;
  assign n8141 = ~pi445 & n8140;
  assign n8142 = n8119 & ~n8141;
  assign n8143 = pi426 & ~n8138;
  assign n8144 = ~pi426 & ~n8134;
  assign n8145 = ~n8143 & ~n8144;
  assign n8146 = pi445 & n8145;
  assign n8147 = n8142 & ~n8146;
  assign n8148 = pi445 & n8140;
  assign n8149 = ~pi445 & n8145;
  assign n8150 = ~n8119 & ~n8149;
  assign n8151 = ~n8148 & n8150;
  assign n8152 = ~n8147 & ~n8151;
  assign n8153 = pi1199 & n8152;
  assign n8154 = ~n8116 & ~n8153;
  assign n8155 = n7958 & n8154;
  assign n8156 = n7503 & ~n7958;
  assign n8157 = n7376 & ~n8156;
  assign n8158 = ~n8155 & n8157;
  assign n8159 = ~pi1196 & n7582;
  assign n8160 = ~pi436 & pi444;
  assign n8161 = pi436 & ~pi444;
  assign n8162 = ~n8160 & ~n8161;
  assign n8163 = ~n8032 & ~n8162;
  assign n8164 = n8032 & n8162;
  assign n8165 = ~n8163 & ~n8164;
  assign n8166 = n7582 & ~n8094;
  assign n8167 = ~n8096 & ~n8166;
  assign n8168 = ~n8165 & n8167;
  assign n8169 = n7582 & ~n8089;
  assign n8170 = ~n8091 & ~n8169;
  assign n8171 = n8165 & n8170;
  assign n8172 = ~n8168 & ~n8171;
  assign n8173 = pi1196 & n8172;
  assign n8174 = ~n8159 & ~n8173;
  assign n8175 = n8011 & ~n8174;
  assign n8176 = pi592 & n7582;
  assign n8177 = ~n8084 & ~n8176;
  assign n8178 = ~n8011 & ~n8177;
  assign n8179 = ~n8175 & ~n8178;
  assign n8180 = ~pi1199 & ~n8179;
  assign n8181 = pi445 & ~n8119;
  assign n8182 = ~pi445 & n8119;
  assign n8183 = ~n8181 & ~n8182;
  assign n8184 = n8052 & n8177;
  assign n8185 = ~n8052 & n8179;
  assign n8186 = ~n8184 & ~n8185;
  assign n8187 = pi430 & ~n8186;
  assign n8188 = pi428 & n8179;
  assign n8189 = ~pi428 & n8177;
  assign n8190 = pi427 & ~n8189;
  assign n8191 = ~n8188 & n8190;
  assign n8192 = ~pi428 & n8179;
  assign n8193 = pi428 & n8177;
  assign n8194 = ~pi427 & ~n8193;
  assign n8195 = ~n8192 & n8194;
  assign n8196 = ~n8191 & ~n8195;
  assign n8197 = ~pi430 & n8196;
  assign n8198 = ~n8187 & ~n8197;
  assign n8199 = ~pi426 & n8198;
  assign n8200 = ~n8183 & ~n8199;
  assign n8201 = ~pi430 & ~n8186;
  assign n8202 = pi430 & n8196;
  assign n8203 = ~n8201 & ~n8202;
  assign n8204 = pi426 & n8203;
  assign n8205 = n8200 & ~n8204;
  assign n8206 = ~pi426 & n8203;
  assign n8207 = pi426 & n8198;
  assign n8208 = ~n8206 & ~n8207;
  assign n8209 = n8183 & n8208;
  assign n8210 = ~n8205 & ~n8209;
  assign n8211 = pi1199 & n8210;
  assign n8212 = ~n8180 & ~n8211;
  assign n8213 = n7958 & n8212;
  assign n8214 = ~n7582 & ~n7958;
  assign n8215 = ~n7376 & ~n8214;
  assign n8216 = ~n8213 & n8215;
  assign n8217 = ~n8158 & ~n8216;
  assign n8218 = pi588 & ~n8217;
  assign n8219 = pi377 & pi592;
  assign n8220 = ~n7503 & ~n8219;
  assign n8221 = ~n8083 & n8219;
  assign n8222 = n7784 & ~n8221;
  assign n8223 = ~n8220 & n8222;
  assign n8224 = ~pi377 & pi592;
  assign n8225 = ~n7503 & ~n8224;
  assign n8226 = ~n8083 & n8224;
  assign n8227 = ~n7784 & ~n8226;
  assign n8228 = ~n8225 & n8227;
  assign n8229 = ~n8223 & ~n8228;
  assign n8230 = n7763 & ~n8229;
  assign n8231 = pi592 & ~n8083;
  assign n8232 = ~pi592 & ~n7503;
  assign n8233 = ~n8231 & ~n8232;
  assign n8234 = ~n7763 & n8233;
  assign n8235 = ~n8230 & ~n8234;
  assign n8236 = pi1199 & n8235;
  assign n8237 = ~pi1196 & ~n7762;
  assign n8238 = n8233 & ~n8237;
  assign n8239 = n7503 & ~n7762;
  assign n8240 = ~pi1196 & n8239;
  assign n8241 = ~n8238 & ~n8240;
  assign n8242 = ~n7736 & ~n8241;
  assign n8243 = n7762 & n8233;
  assign n8244 = ~n8239 & ~n8243;
  assign n8245 = n7736 & ~n8244;
  assign n8246 = ~pi1199 & ~n8245;
  assign n8247 = ~n8242 & n8246;
  assign n8248 = ~n8236 & ~n8247;
  assign n8249 = ~pi374 & ~n8248;
  assign n8250 = ~pi1198 & ~n8248;
  assign n8251 = pi1198 & ~n8233;
  assign n8252 = ~n8250 & ~n8251;
  assign n8253 = pi374 & ~n8252;
  assign n8254 = ~n8249 & ~n8253;
  assign n8255 = ~pi369 & ~n8254;
  assign n8256 = ~pi374 & ~n8252;
  assign n8257 = pi374 & ~n8248;
  assign n8258 = ~n8256 & ~n8257;
  assign n8259 = pi369 & ~n8258;
  assign n8260 = ~n8255 & ~n8259;
  assign n8261 = n7798 & n8260;
  assign n8262 = pi369 & ~n8254;
  assign n8263 = ~pi369 & ~n8258;
  assign n8264 = ~n8262 & ~n8263;
  assign n8265 = ~n7798 & n8264;
  assign n8266 = ~n8261 & ~n8265;
  assign n8267 = ~pi373 & ~n8266;
  assign n8268 = ~pi370 & n8264;
  assign n8269 = ~pi371 & ~n8268;
  assign n8270 = pi370 & n8260;
  assign n8271 = n8269 & ~n8270;
  assign n8272 = ~pi370 & n8260;
  assign n8273 = pi371 & ~n8272;
  assign n8274 = pi370 & n8264;
  assign n8275 = n8273 & ~n8274;
  assign n8276 = ~n8271 & ~n8275;
  assign n8277 = pi373 & n8276;
  assign n8278 = ~n8267 & ~n8277;
  assign n8279 = ~pi375 & ~n8278;
  assign n8280 = pi373 & ~n8266;
  assign n8281 = ~pi373 & n8276;
  assign n8282 = ~n8280 & ~n8281;
  assign n8283 = pi375 & ~n8282;
  assign n8284 = ~n8279 & ~n8283;
  assign n8285 = ~n7804 & n8284;
  assign n8286 = ~pi375 & ~n8282;
  assign n8287 = pi375 & ~n8278;
  assign n8288 = n7804 & ~n8287;
  assign n8289 = ~n8286 & n8288;
  assign n8290 = ~pi591 & ~n8289;
  assign n8291 = ~n8285 & n8290;
  assign n8292 = pi1197 & ~n8086;
  assign n8293 = pi1198 & ~n7915;
  assign n8294 = n8086 & n8293;
  assign n8295 = ~pi75 & ~pi592;
  assign n8296 = ~n7501 & ~n8295;
  assign n8297 = n7491 & ~n7849;
  assign n8298 = n7490 & ~n8297;
  assign n8299 = pi87 & n2615;
  assign n8300 = ~n7495 & n8299;
  assign n8301 = ~n8298 & n8300;
  assign n8302 = n7478 & ~n7849;
  assign n8303 = n7475 & ~n8302;
  assign n8304 = n8075 & ~n8303;
  assign n8305 = n8295 & ~n8304;
  assign n8306 = ~n8301 & n8305;
  assign n8307 = pi1196 & ~n8306;
  assign n8308 = ~pi1196 & ~n7500;
  assign n8309 = ~pi1199 & ~n8308;
  assign n8310 = ~n8307 & n8309;
  assign n8311 = n7491 & n7874;
  assign n8312 = n7490 & ~n8311;
  assign n8313 = pi1196 & n8298;
  assign n8314 = n8300 & ~n8313;
  assign n8315 = ~n8312 & n8314;
  assign n8316 = pi1199 & ~n8315;
  assign n8317 = ~pi75 & n7850;
  assign n8318 = n7874 & ~n8317;
  assign n8319 = n7478 & n8318;
  assign n8320 = n7475 & ~n8319;
  assign n8321 = n8075 & ~n8320;
  assign n8322 = n8295 & ~n8321;
  assign n8323 = n8316 & n8322;
  assign n8324 = ~n8310 & ~n8323;
  assign n8325 = ~n8296 & n8324;
  assign n8326 = pi567 & ~n8325;
  assign n8327 = ~n8293 & ~n8326;
  assign n8328 = n7419 & n8327;
  assign n8329 = ~n8294 & ~n8328;
  assign n8330 = ~pi1197 & n8329;
  assign n8331 = ~n8292 & ~n8330;
  assign n8332 = pi333 & ~n8331;
  assign n8333 = ~pi333 & n8329;
  assign n8334 = ~n8332 & ~n8333;
  assign n8335 = ~pi391 & ~n8334;
  assign n8336 = ~pi333 & ~n8331;
  assign n8337 = pi333 & n8329;
  assign n8338 = ~n8336 & ~n8337;
  assign n8339 = pi391 & ~n8338;
  assign n8340 = ~n8335 & ~n8339;
  assign n8341 = ~pi392 & ~n8340;
  assign n8342 = pi391 & ~n8334;
  assign n8343 = ~pi391 & ~n8338;
  assign n8344 = ~n8342 & ~n8343;
  assign n8345 = pi392 & ~n8344;
  assign n8346 = ~n8341 & ~n8345;
  assign n8347 = ~pi393 & ~n8346;
  assign n8348 = ~pi392 & ~n8344;
  assign n8349 = pi392 & ~n8340;
  assign n8350 = ~n8348 & ~n8349;
  assign n8351 = pi393 & ~n8350;
  assign n8352 = ~n8347 & ~n8351;
  assign n8353 = ~pi334 & n8352;
  assign n8354 = ~n7928 & ~n8353;
  assign n8355 = ~pi393 & ~n8350;
  assign n8356 = pi393 & ~n8346;
  assign n8357 = ~n8355 & ~n8356;
  assign n8358 = pi334 & n8357;
  assign n8359 = n8354 & ~n8358;
  assign n8360 = ~pi334 & n8357;
  assign n8361 = n7928 & ~n8360;
  assign n8362 = pi334 & n8352;
  assign n8363 = n8361 & ~n8362;
  assign n8364 = pi591 & ~n8363;
  assign n8365 = ~n8359 & n8364;
  assign n8366 = ~pi590 & ~n8365;
  assign n8367 = ~n8291 & n8366;
  assign n8368 = ~pi350 & ~pi592;
  assign n8369 = ~n7503 & ~n8368;
  assign n8370 = ~n8083 & n8368;
  assign n8371 = ~n7664 & ~n8370;
  assign n8372 = ~n8369 & n8371;
  assign n8373 = pi350 & ~pi592;
  assign n8374 = ~n7503 & ~n8373;
  assign n8375 = ~n8083 & n8373;
  assign n8376 = n7664 & ~n8375;
  assign n8377 = ~n8374 & n8376;
  assign n8378 = ~n7643 & ~n8377;
  assign n8379 = ~n8372 & n8378;
  assign n8380 = n7643 & ~n8086;
  assign n8381 = pi1198 & ~n8380;
  assign n8382 = ~n8379 & n8381;
  assign n8383 = ~pi455 & n8086;
  assign n8384 = ~pi452 & ~n8383;
  assign n8385 = pi455 & n7503;
  assign n8386 = n8384 & ~n8385;
  assign n8387 = ~pi455 & n7503;
  assign n8388 = pi452 & ~n8387;
  assign n8389 = pi455 & n8086;
  assign n8390 = n8388 & ~n8389;
  assign n8391 = ~n8386 & ~n8390;
  assign n8392 = ~pi355 & ~n8391;
  assign n8393 = ~n7617 & ~n8086;
  assign n8394 = ~n7503 & n7617;
  assign n8395 = ~n8393 & ~n8394;
  assign n8396 = pi355 & ~n8395;
  assign n8397 = ~n8392 & ~n8396;
  assign n8398 = pi458 & ~n8397;
  assign n8399 = pi355 & ~n8391;
  assign n8400 = ~pi355 & ~n8395;
  assign n8401 = ~n8399 & ~n8400;
  assign n8402 = ~pi458 & ~n8401;
  assign n8403 = n7629 & ~n8402;
  assign n8404 = ~n8398 & n8403;
  assign n8405 = pi458 & ~n8401;
  assign n8406 = ~pi458 & ~n8397;
  assign n8407 = ~n7629 & ~n8406;
  assign n8408 = ~n8405 & n8407;
  assign n8409 = pi1196 & ~n8408;
  assign n8410 = ~n8404 & n8409;
  assign n8411 = ~pi1198 & ~n8088;
  assign n8412 = ~n8410 & n8411;
  assign n8413 = ~n8382 & ~n8412;
  assign n8414 = ~n7614 & ~n8413;
  assign n8415 = n7614 & n8086;
  assign n8416 = ~n8414 & ~n8415;
  assign n8417 = ~n7589 & n8416;
  assign n8418 = pi1199 & ~n8086;
  assign n8419 = ~pi351 & n8418;
  assign n8420 = ~n8417 & ~n8419;
  assign n8421 = ~pi461 & ~n8420;
  assign n8422 = ~n7700 & n8416;
  assign n8423 = pi351 & n8418;
  assign n8424 = ~n8422 & ~n8423;
  assign n8425 = pi461 & ~n8424;
  assign n8426 = ~n8421 & ~n8425;
  assign n8427 = ~pi357 & ~n8426;
  assign n8428 = ~pi461 & ~n8424;
  assign n8429 = pi461 & ~n8420;
  assign n8430 = ~n8428 & ~n8429;
  assign n8431 = pi357 & ~n8430;
  assign n8432 = ~n8427 & ~n8431;
  assign n8433 = ~pi356 & n8432;
  assign n8434 = n7693 & ~n8433;
  assign n8435 = ~pi357 & ~n8430;
  assign n8436 = pi357 & ~n8426;
  assign n8437 = ~n8435 & ~n8436;
  assign n8438 = pi356 & n8437;
  assign n8439 = n8434 & ~n8438;
  assign n8440 = ~pi356 & n8437;
  assign n8441 = pi356 & n8432;
  assign n8442 = ~n8440 & ~n8441;
  assign n8443 = ~n7693 & n8442;
  assign n8444 = ~pi591 & ~n8443;
  assign n8445 = ~n8439 & n8444;
  assign n8446 = pi591 & n7503;
  assign n8447 = pi590 & ~n8446;
  assign n8448 = ~n8445 & n8447;
  assign n8449 = ~n8367 & ~n8448;
  assign n8450 = n7376 & n8449;
  assign n8451 = pi455 & ~n8177;
  assign n8452 = ~pi455 & n7582;
  assign n8453 = ~n8451 & ~n8452;
  assign n8454 = pi452 & ~n8453;
  assign n8455 = ~pi455 & ~n8177;
  assign n8456 = pi455 & n7582;
  assign n8457 = ~n8455 & ~n8456;
  assign n8458 = ~pi452 & ~n8457;
  assign n8459 = n7635 & ~n8458;
  assign n8460 = ~n8454 & n8459;
  assign n8461 = pi452 & ~n8457;
  assign n8462 = ~pi452 & ~n8453;
  assign n8463 = ~n7635 & ~n8462;
  assign n8464 = ~n8461 & n8463;
  assign n8465 = ~n8460 & ~n8464;
  assign n8466 = pi1196 & n8465;
  assign n8467 = ~pi1198 & ~n8466;
  assign n8468 = ~n8159 & n8467;
  assign n8469 = n7643 & ~n8177;
  assign n8470 = pi1198 & ~n8469;
  assign n8471 = n7582 & ~n8373;
  assign n8472 = n8376 & ~n8471;
  assign n8473 = n7582 & ~n8368;
  assign n8474 = n8371 & ~n8473;
  assign n8475 = ~n8472 & ~n8474;
  assign n8476 = ~n7643 & n8475;
  assign n8477 = n8470 & ~n8476;
  assign n8478 = ~n7614 & ~n8477;
  assign n8479 = ~n8468 & n8478;
  assign n8480 = n7614 & ~n8177;
  assign n8481 = ~n8479 & ~n8480;
  assign n8482 = ~n7589 & ~n8481;
  assign n8483 = pi1199 & ~n8177;
  assign n8484 = ~pi351 & n8483;
  assign n8485 = ~n8482 & ~n8484;
  assign n8486 = ~pi461 & ~n8485;
  assign n8487 = ~n7700 & ~n8481;
  assign n8488 = pi351 & n8483;
  assign n8489 = ~n8487 & ~n8488;
  assign n8490 = pi461 & ~n8489;
  assign n8491 = ~n8486 & ~n8490;
  assign n8492 = ~pi357 & ~n8491;
  assign n8493 = ~pi461 & ~n8489;
  assign n8494 = pi461 & ~n8485;
  assign n8495 = ~n8493 & ~n8494;
  assign n8496 = pi357 & ~n8495;
  assign n8497 = ~n8492 & ~n8496;
  assign n8498 = ~pi356 & n8497;
  assign n8499 = n7693 & ~n8498;
  assign n8500 = ~pi357 & ~n8495;
  assign n8501 = pi357 & ~n8491;
  assign n8502 = ~n8500 & ~n8501;
  assign n8503 = pi356 & n8502;
  assign n8504 = n8499 & ~n8503;
  assign n8505 = ~pi356 & n8502;
  assign n8506 = pi356 & n8497;
  assign n8507 = ~n8505 & ~n8506;
  assign n8508 = ~n7693 & n8507;
  assign n8509 = ~pi591 & ~n8508;
  assign n8510 = ~n8504 & n8509;
  assign n8511 = pi591 & ~n7582;
  assign n8512 = pi590 & ~n8511;
  assign n8513 = ~n8510 & n8512;
  assign n8514 = n7582 & ~n8224;
  assign n8515 = n8227 & ~n8514;
  assign n8516 = n7582 & ~n8219;
  assign n8517 = n8222 & ~n8516;
  assign n8518 = ~n8515 & ~n8517;
  assign n8519 = pi1199 & ~n8518;
  assign n8520 = ~pi1199 & ~n7582;
  assign n8521 = ~n8519 & ~n8520;
  assign n8522 = n7763 & ~n8521;
  assign n8523 = ~pi592 & n7582;
  assign n8524 = ~n8231 & ~n8523;
  assign n8525 = ~n7763 & n8524;
  assign n8526 = ~n8522 & ~n8525;
  assign n8527 = pi374 & ~n8526;
  assign n8528 = ~pi1198 & ~n8526;
  assign n8529 = pi1198 & n8524;
  assign n8530 = ~n8528 & ~n8529;
  assign n8531 = ~pi374 & ~n8530;
  assign n8532 = ~n8527 & ~n8531;
  assign n8533 = ~pi369 & ~n8532;
  assign n8534 = pi374 & ~n8530;
  assign n8535 = ~pi374 & ~n8526;
  assign n8536 = ~n8534 & ~n8535;
  assign n8537 = pi369 & ~n8536;
  assign n8538 = ~n8533 & ~n8537;
  assign n8539 = pi370 & ~n8538;
  assign n8540 = pi369 & ~n8532;
  assign n8541 = ~pi369 & ~n8536;
  assign n8542 = ~n8540 & ~n8541;
  assign n8543 = ~pi370 & ~n8542;
  assign n8544 = ~n8539 & ~n8543;
  assign n8545 = ~pi371 & ~n8544;
  assign n8546 = pi370 & ~n8542;
  assign n8547 = ~pi370 & ~n8538;
  assign n8548 = ~n8546 & ~n8547;
  assign n8549 = pi371 & ~n8548;
  assign n8550 = n7810 & ~n8549;
  assign n8551 = ~n8545 & n8550;
  assign n8552 = pi371 & ~n8544;
  assign n8553 = ~pi371 & ~n8548;
  assign n8554 = ~n7810 & ~n8553;
  assign n8555 = ~n8552 & n8554;
  assign n8556 = ~pi591 & ~n8555;
  assign n8557 = ~n8551 & n8556;
  assign n8558 = n8084 & n8293;
  assign n8559 = ~n7380 & n7884;
  assign n8560 = pi38 & n7883;
  assign n8561 = ~pi100 & ~n8560;
  assign n8562 = n7458 & n7849;
  assign n8563 = n7528 & ~n8562;
  assign n8564 = n6215 & ~n6236;
  assign n8565 = ~n6191 & n6236;
  assign n8566 = n7463 & ~n8565;
  assign n8567 = ~n8564 & n8566;
  assign n8568 = n7529 & n8567;
  assign n8569 = ~pi299 & n8568;
  assign n8570 = ~n6198 & n6215;
  assign n8571 = ~n6191 & n6198;
  assign n8572 = n7463 & ~n8571;
  assign n8573 = ~n8570 & n8572;
  assign n8574 = n5745 & n8573;
  assign n8575 = pi299 & n8574;
  assign n8576 = ~n7883 & ~n8575;
  assign n8577 = ~n8569 & n8576;
  assign n8578 = pi39 & ~n8577;
  assign n8579 = ~n8563 & ~n8578;
  assign n8580 = ~pi38 & ~n8579;
  assign n8581 = n8561 & ~n8580;
  assign n8582 = n7487 & ~n7883;
  assign n8583 = ~n8581 & ~n8582;
  assign n8584 = ~pi87 & ~n8583;
  assign n8585 = ~n2615 & n7883;
  assign n8586 = pi87 & ~n8585;
  assign n8587 = n7566 & n7849;
  assign n8588 = n7573 & ~n8587;
  assign n8589 = n8586 & ~n8588;
  assign n8590 = ~n8584 & ~n8589;
  assign n8591 = ~pi75 & ~n8590;
  assign n8592 = ~n7422 & n7883;
  assign n8593 = pi75 & ~n8592;
  assign n8594 = ~pi1091 & ~n7882;
  assign n8595 = n7508 & ~n8594;
  assign n8596 = n8593 & ~n8595;
  assign n8597 = ~n8591 & ~n8596;
  assign n8598 = pi567 & ~n8597;
  assign n8599 = n7419 & ~n8598;
  assign n8600 = ~n8559 & ~n8599;
  assign n8601 = n7881 & n8600;
  assign n8602 = ~pi1199 & ~n8159;
  assign n8603 = ~n8601 & n8602;
  assign n8604 = n7509 & n7874;
  assign n8605 = n8559 & n8604;
  assign n8606 = n7881 & ~n8605;
  assign n8607 = ~n7380 & n7877;
  assign n8608 = ~pi592 & ~pi1196;
  assign n8609 = ~n8607 & n8608;
  assign n8610 = ~n8606 & ~n8609;
  assign n8611 = ~n7419 & ~n8610;
  assign n8612 = n7526 & n7874;
  assign n8613 = n7458 & ~n8612;
  assign n8614 = n8563 & ~n8613;
  assign n8615 = n7874 & n7883;
  assign n8616 = ~n8573 & ~n8615;
  assign n8617 = n5745 & ~n8616;
  assign n8618 = ~n5745 & n7876;
  assign n8619 = n7883 & n8618;
  assign n8620 = ~n8617 & ~n8619;
  assign n8621 = pi299 & n8620;
  assign n8622 = ~n7529 & n7876;
  assign n8623 = n7883 & n8622;
  assign n8624 = ~pi299 & ~n8568;
  assign n8625 = n7529 & n8615;
  assign n8626 = n8624 & ~n8625;
  assign n8627 = ~n8623 & n8626;
  assign n8628 = pi39 & ~n8627;
  assign n8629 = ~n8621 & n8628;
  assign n8630 = ~n8614 & ~n8629;
  assign n8631 = ~pi38 & ~n8630;
  assign n8632 = pi38 & n7876;
  assign n8633 = ~pi100 & ~n8632;
  assign n8634 = ~n8561 & ~n8633;
  assign n8635 = ~n8631 & ~n8634;
  assign n8636 = n6100 & n7483;
  assign n8637 = ~n6101 & n6190;
  assign n8638 = ~n6100 & ~n8637;
  assign n8639 = ~pi1091 & ~n8615;
  assign n8640 = ~n7517 & ~n8639;
  assign n8641 = n8638 & n8640;
  assign n8642 = ~n8636 & ~n8641;
  assign n8643 = pi228 & ~n8642;
  assign n8644 = pi228 & n8638;
  assign n8645 = n8615 & ~n8644;
  assign n8646 = pi232 & ~n8645;
  assign n8647 = ~n8643 & n8646;
  assign n8648 = pi228 & n7483;
  assign n8649 = ~pi232 & ~n8615;
  assign n8650 = ~n8648 & n8649;
  assign n8651 = ~n8647 & ~n8650;
  assign n8652 = n2532 & n8651;
  assign n8653 = ~n2532 & n8615;
  assign n8654 = pi100 & ~n8653;
  assign n8655 = ~n8652 & n8654;
  assign n8656 = ~n8635 & ~n8655;
  assign n8657 = ~pi87 & ~n8656;
  assign n8658 = ~n2615 & n7876;
  assign n8659 = pi87 & ~n8658;
  assign n8660 = ~n8586 & ~n8659;
  assign n8661 = n7566 & ~n7874;
  assign n8662 = n7573 & ~n8661;
  assign n8663 = ~n8587 & n8662;
  assign n8664 = ~n8660 & ~n8663;
  assign n8665 = ~n8657 & ~n8664;
  assign n8666 = ~pi75 & ~n8665;
  assign n8667 = ~n7422 & n7876;
  assign n8668 = pi75 & ~n8667;
  assign n8669 = ~n8593 & ~n8668;
  assign n8670 = n7508 & ~n8639;
  assign n8671 = ~n8669 & ~n8670;
  assign n8672 = ~n8666 & ~n8671;
  assign n8673 = n8606 & ~n8672;
  assign n8674 = n8659 & ~n8662;
  assign n8675 = n7487 & ~n7876;
  assign n8676 = n7523 & ~n8613;
  assign n8677 = ~n7876 & n8624;
  assign n8678 = pi299 & ~n7876;
  assign n8679 = ~n8574 & n8678;
  assign n8680 = pi39 & ~n8679;
  assign n8681 = ~n8677 & n8680;
  assign n8682 = ~n8676 & ~n8681;
  assign n8683 = ~pi38 & ~n8682;
  assign n8684 = n8633 & ~n8683;
  assign n8685 = ~n8675 & ~n8684;
  assign n8686 = ~pi87 & ~n8685;
  assign n8687 = ~n8674 & ~n8686;
  assign n8688 = ~pi75 & ~n8687;
  assign n8689 = ~pi1091 & ~n7875;
  assign n8690 = n7508 & ~n8689;
  assign n8691 = n8668 & ~n8690;
  assign n8692 = ~n8688 & ~n8691;
  assign n8693 = n8609 & ~n8692;
  assign n8694 = ~n8673 & ~n8693;
  assign n8695 = pi567 & ~n8694;
  assign n8696 = ~n8611 & ~n8695;
  assign n8697 = pi1199 & n8696;
  assign n8698 = ~n8293 & ~n8697;
  assign n8699 = ~n8603 & n8698;
  assign n8700 = ~n8558 & ~n8699;
  assign n8701 = ~n8176 & n8700;
  assign n8702 = ~pi1197 & ~n8701;
  assign n8703 = pi1197 & ~n8177;
  assign n8704 = ~n8702 & ~n8703;
  assign n8705 = ~pi333 & ~n8704;
  assign n8706 = pi333 & ~n8701;
  assign n8707 = ~n8705 & ~n8706;
  assign n8708 = ~pi391 & ~n8707;
  assign n8709 = ~pi333 & ~n8701;
  assign n8710 = pi333 & ~n8704;
  assign n8711 = ~n8709 & ~n8710;
  assign n8712 = pi391 & ~n8711;
  assign n8713 = ~n8708 & ~n8712;
  assign n8714 = ~n7937 & ~n8713;
  assign n8715 = ~pi391 & ~n8711;
  assign n8716 = pi391 & ~n8707;
  assign n8717 = ~n8715 & ~n8716;
  assign n8718 = n7937 & ~n8717;
  assign n8719 = ~n8714 & ~n8718;
  assign n8720 = pi591 & n8719;
  assign n8721 = ~pi590 & ~n8720;
  assign n8722 = ~n8557 & n8721;
  assign n8723 = ~n8513 & ~n8722;
  assign n8724 = ~n7376 & n8723;
  assign n8725 = ~pi588 & ~n8724;
  assign n8726 = ~n8450 & n8725;
  assign n8727 = ~n8218 & ~n8726;
  assign n8728 = ~po1038 & n8727;
  assign n8729 = ~pi217 & ~n8728;
  assign n8730 = ~n8074 & n8729;
  assign n8731 = n7588 & ~n8730;
  assign n8732 = ~n7586 & n8731;
  assign n8733 = pi1161 & ~pi1163;
  assign n8734 = pi1162 & n2934;
  assign n8735 = n8733 & n8734;
  assign n8736 = ~pi31 & n8735;
  assign po189 = n8732 | n8736;
  assign n8738 = ~pi74 & ~po1038;
  assign n8739 = n6094 & n8738;
  assign n8740 = pi100 & n2532;
  assign n8741 = n6128 & n6489;
  assign n8742 = ~pi137 & n8741;
  assign n8743 = pi129 & n2522;
  assign n8744 = po1057 & ~n7421;
  assign n8745 = pi252 & ~n8744;
  assign n8746 = ~pi137 & n8745;
  assign n8747 = ~n6106 & n8746;
  assign n8748 = n8743 & n8747;
  assign n8749 = ~n8742 & ~n8748;
  assign n8750 = n8740 & ~n8749;
  assign n8751 = pi829 & ~pi1093;
  assign n8752 = n6120 & n8751;
  assign po840 = n2978 | n8752;
  assign n8754 = ~n7376 & ~po840;
  assign n8755 = ~pi137 & ~n8754;
  assign n8756 = pi50 & n2763;
  assign n8757 = ~pi103 & n2795;
  assign n8758 = n2463 & n2476;
  assign n8759 = n8757 & n8758;
  assign n8760 = n2467 & n2788;
  assign n8761 = ~pi45 & ~pi48;
  assign n8762 = ~pi61 & n8761;
  assign n8763 = ~pi104 & n8762;
  assign n8764 = n8760 & n8763;
  assign n8765 = n8759 & n8764;
  assign n8766 = ~pi68 & ~pi73;
  assign n8767 = ~pi49 & n8766;
  assign n8768 = n8765 & n8767;
  assign n8769 = ~pi111 & n8768;
  assign n8770 = ~pi89 & ~pi102;
  assign n8771 = n2464 & n8770;
  assign n8772 = ~pi64 & ~pi81;
  assign n8773 = n2488 & n8772;
  assign n8774 = n8771 & n8773;
  assign n8775 = ~pi82 & ~pi84;
  assign n8776 = n8774 & n8775;
  assign n8777 = ~pi66 & n8776;
  assign n8778 = pi76 & n8777;
  assign n8779 = n8769 & n8778;
  assign n8780 = ~n8756 & ~n8779;
  assign n8781 = n2689 & n2694;
  assign n8782 = ~n8780 & n8781;
  assign n8783 = ~pi24 & ~n8782;
  assign n8784 = n2688 & n2694;
  assign n8785 = n2494 & n8779;
  assign n8786 = n8784 & n8785;
  assign n8787 = pi24 & ~n8786;
  assign n8788 = n2919 & ~n8787;
  assign n8789 = ~n8783 & n8788;
  assign n8790 = n7394 & n8789;
  assign n8791 = n8755 & ~n8790;
  assign n8792 = ~pi24 & ~pi90;
  assign n8793 = n2920 & n8792;
  assign n8794 = n2494 & n8756;
  assign n8795 = ~pi93 & n8784;
  assign n8796 = n8794 & n8795;
  assign n8797 = n8793 & n8796;
  assign n8798 = ~n8755 & ~n8797;
  assign n8799 = ~pi32 & ~n8798;
  assign n8800 = ~n8791 & n8799;
  assign n8801 = ~pi24 & ~pi841;
  assign n8802 = pi32 & ~n8801;
  assign n8803 = n2700 & n8802;
  assign n8804 = ~n8800 & ~n8803;
  assign n8805 = ~n6166 & n8804;
  assign n8806 = ~pi39 & ~pi95;
  assign n8807 = ~pi32 & ~n8797;
  assign n8808 = ~n6168 & ~n8807;
  assign n8809 = n6166 & ~n8808;
  assign n8810 = n8806 & ~n8809;
  assign n8811 = n2614 & n8810;
  assign n8812 = ~n8805 & n8811;
  assign n8813 = ~n8750 & ~n8812;
  assign n8814 = n2535 & ~n8813;
  assign n8815 = ~pi24 & n2520;
  assign n8816 = n2517 & n2917;
  assign n8817 = n8815 & n8816;
  assign n8818 = ~po840 & n8817;
  assign n8819 = n6106 & po1057;
  assign n8820 = ~pi87 & n2532;
  assign n8821 = pi75 & ~pi100;
  assign n8822 = n8820 & n8821;
  assign n8823 = ~n8745 & n8822;
  assign n8824 = ~n8819 & n8823;
  assign n8825 = ~pi137 & n8824;
  assign n8826 = n8818 & n8825;
  assign n8827 = ~n8814 & ~n8826;
  assign po190 = n8739 & ~n8827;
  assign n8829 = ~pi195 & ~pi196;
  assign n8830 = ~pi138 & n8829;
  assign n8831 = ~pi139 & n8830;
  assign n8832 = ~pi118 & n8831;
  assign n8833 = ~pi79 & n8832;
  assign n8834 = ~pi34 & n8833;
  assign n8835 = ~pi33 & ~n8834;
  assign n8836 = pi149 & pi157;
  assign n8837 = ~pi149 & ~pi157;
  assign n8838 = n6190 & ~n8837;
  assign n8839 = ~n8836 & n8838;
  assign n8840 = pi232 & n8839;
  assign n8841 = pi75 & ~n8840;
  assign n8842 = pi100 & ~n8840;
  assign n8843 = ~n8841 & ~n8842;
  assign n8844 = pi169 & n7420;
  assign n8845 = n7255 & n8844;
  assign n8846 = n8843 & ~n8845;
  assign n8847 = pi74 & ~n8846;
  assign n8848 = pi164 & n7420;
  assign n8849 = n7255 & n8848;
  assign n8850 = n8843 & ~n8849;
  assign n8851 = ~pi74 & ~n8850;
  assign n8852 = ~n3327 & ~n8851;
  assign n8853 = ~n8847 & n8852;
  assign n8854 = pi54 & ~n8850;
  assign n8855 = pi38 & n8849;
  assign n8856 = n8843 & ~n8855;
  assign n8857 = ~n8854 & n8856;
  assign n8858 = ~pi74 & ~n8857;
  assign n8859 = ~n8847 & ~n8858;
  assign n8860 = ~n2531 & ~n8859;
  assign n8861 = n3327 & ~n8860;
  assign n8862 = ~pi40 & n2488;
  assign n8863 = ~pi38 & n8862;
  assign n8864 = n7255 & n8863;
  assign n8865 = n2534 & n8864;
  assign n8866 = ~n2531 & n8865;
  assign n8867 = pi55 & ~n8847;
  assign n8868 = ~pi92 & ~n8841;
  assign n8869 = n2466 & n8772;
  assign n8870 = n2487 & n8869;
  assign n8871 = ~pi60 & n8870;
  assign n8872 = n2498 & n2501;
  assign n8873 = n2706 & n8872;
  assign n8874 = ~pi53 & n8873;
  assign n8875 = n8871 & n8874;
  assign n8876 = ~pi58 & n8875;
  assign n8877 = n7394 & n8876;
  assign n8878 = n2918 & n8877;
  assign n8879 = n2516 & n8878;
  assign n8880 = pi149 & n7420;
  assign n8881 = ~pi39 & ~n8880;
  assign n8882 = n8879 & n8881;
  assign n8883 = n8862 & ~n8882;
  assign n8884 = ~pi38 & ~n8883;
  assign n8885 = pi38 & ~n8848;
  assign n8886 = ~pi100 & ~n8885;
  assign n8887 = ~pi87 & n8886;
  assign n8888 = ~n8884 & n8887;
  assign n8889 = ~pi38 & ~n8862;
  assign n8890 = n8886 & ~n8889;
  assign n8891 = pi87 & n8890;
  assign n8892 = ~n8842 & ~n8891;
  assign n8893 = ~n8888 & n8892;
  assign n8894 = ~pi75 & ~n8893;
  assign n8895 = n8868 & ~n8894;
  assign n8896 = ~pi75 & n8890;
  assign n8897 = pi92 & ~n8896;
  assign n8898 = n8843 & n8897;
  assign n8899 = ~pi54 & ~n8898;
  assign n8900 = ~n8895 & n8899;
  assign n8901 = ~n8854 & ~n8900;
  assign n8902 = ~pi74 & ~n8901;
  assign n8903 = n8867 & ~n8902;
  assign n8904 = pi178 & pi183;
  assign n8905 = ~pi178 & ~pi183;
  assign n8906 = n6190 & ~n8905;
  assign n8907 = ~n8904 & n8906;
  assign n8908 = ~pi299 & ~n8907;
  assign n8909 = pi299 & ~n8839;
  assign n8910 = pi232 & ~n8909;
  assign n8911 = ~n8908 & n8910;
  assign n8912 = pi100 & ~n8911;
  assign n8913 = pi75 & ~n8911;
  assign n8914 = ~n8912 & ~n8913;
  assign n8915 = n7255 & n7420;
  assign n8916 = pi191 & ~pi299;
  assign n8917 = pi169 & pi299;
  assign n8918 = ~n8916 & ~n8917;
  assign n8919 = n8915 & ~n8918;
  assign n8920 = n8914 & ~n8919;
  assign n8921 = pi74 & ~n8920;
  assign n8922 = ~pi55 & ~n8921;
  assign n8923 = ~pi186 & ~pi299;
  assign n8924 = ~pi299 & n7420;
  assign n8925 = ~n8848 & ~n8924;
  assign n8926 = ~n8923 & ~n8925;
  assign n8927 = n7255 & n8926;
  assign n8928 = n8914 & ~n8927;
  assign n8929 = pi54 & ~n8928;
  assign n8930 = ~pi75 & pi92;
  assign n8931 = pi38 & n8926;
  assign n8932 = ~pi100 & n8931;
  assign n8933 = ~n8912 & ~n8932;
  assign n8934 = n3257 & n8879;
  assign n8935 = pi232 & ~n3403;
  assign n8936 = ~pi176 & ~pi299;
  assign n8937 = n6190 & ~n8936;
  assign n8938 = n8935 & n8937;
  assign n8939 = n8934 & ~n8938;
  assign n8940 = n2614 & n8862;
  assign n8941 = ~n8939 & n8940;
  assign n8942 = n8933 & ~n8941;
  assign n8943 = n8930 & ~n8942;
  assign n8944 = pi87 & ~n8940;
  assign n8945 = n8933 & n8944;
  assign n8946 = n2573 & ~n8945;
  assign n8947 = pi299 & n7420;
  assign n8948 = ~n6132 & n8947;
  assign n8949 = ~pi186 & ~n8948;
  assign n8950 = ~n6097 & n7420;
  assign n8951 = pi186 & ~n8950;
  assign n8952 = pi164 & ~n8951;
  assign n8953 = ~n8949 & n8952;
  assign n8954 = ~n6132 & n8924;
  assign n8955 = ~pi164 & pi186;
  assign n8956 = n8954 & n8955;
  assign n8957 = ~n8953 & ~n8956;
  assign n8958 = pi38 & ~n8957;
  assign n8959 = pi216 & n5744;
  assign n8960 = n8862 & ~n8959;
  assign n8961 = pi299 & ~n8960;
  assign n8962 = n6206 & ~n6447;
  assign n8963 = n6443 & n8962;
  assign n8964 = ~n6182 & ~n8963;
  assign n8965 = n8879 & ~n8964;
  assign n8966 = n6191 & n8965;
  assign n8967 = n8862 & ~n8966;
  assign n8968 = n6190 & n8965;
  assign n8969 = n8862 & ~n8968;
  assign n8970 = ~n6198 & ~n8969;
  assign n8971 = n8967 & ~n8970;
  assign n8972 = n8961 & ~n8971;
  assign n8973 = pi224 & n6439;
  assign n8974 = n8862 & ~n8973;
  assign n8975 = ~n8967 & ~n8974;
  assign n8976 = ~n6236 & ~n8969;
  assign n8977 = ~n8974 & n8976;
  assign n8978 = ~n8975 & ~n8977;
  assign n8979 = ~pi299 & ~n8978;
  assign n8980 = ~n8972 & ~n8979;
  assign n8981 = ~pi232 & ~n8980;
  assign n8982 = n8879 & n8963;
  assign n8983 = n8862 & ~n8982;
  assign n8984 = n6199 & ~n8983;
  assign n8985 = pi152 & n8984;
  assign n8986 = n8967 & ~n8985;
  assign n8987 = pi154 & ~n8986;
  assign n8988 = n6182 & n8879;
  assign n8989 = ~n6215 & n8988;
  assign n8990 = n8862 & ~n8989;
  assign n8991 = n6190 & n8990;
  assign n8992 = ~pi152 & n8991;
  assign n8993 = ~pi154 & ~n8992;
  assign n8994 = ~n8971 & n8993;
  assign n8995 = ~n8987 & ~n8994;
  assign n8996 = n8959 & n8995;
  assign n8997 = n8961 & ~n8996;
  assign n8998 = n6190 & n8982;
  assign n8999 = n8862 & ~n8998;
  assign n9000 = ~n6236 & ~n8999;
  assign n9001 = ~n8974 & n9000;
  assign n9002 = ~n8975 & ~n9001;
  assign n9003 = ~pi174 & ~n8975;
  assign n9004 = ~pi299 & ~n9003;
  assign n9005 = ~n9002 & n9004;
  assign n9006 = ~n8997 & ~n9005;
  assign n9007 = n6237 & n8988;
  assign n9008 = n8862 & n8973;
  assign n9009 = ~n9007 & n9008;
  assign n9010 = ~n8974 & ~n9009;
  assign n9011 = n8936 & n9010;
  assign n9012 = n9006 & ~n9011;
  assign n9013 = pi232 & ~n9012;
  assign n9014 = pi39 & ~n9013;
  assign n9015 = ~n8981 & n9014;
  assign n9016 = pi95 & ~n8862;
  assign n9017 = ~n2442 & ~n9016;
  assign n9018 = ~pi40 & ~pi479;
  assign n9019 = ~pi32 & n8878;
  assign n9020 = n2488 & ~n9019;
  assign n9021 = n9018 & n9020;
  assign n9022 = ~n9017 & ~n9021;
  assign n9023 = pi32 & ~n8862;
  assign n9024 = n2488 & ~n2506;
  assign n9025 = n2488 & ~n8877;
  assign n9026 = pi70 & ~n9025;
  assign n9027 = n2488 & ~n2519;
  assign n9028 = ~pi70 & ~n9027;
  assign n9029 = ~pi841 & n8876;
  assign n9030 = n2488 & ~n9029;
  assign n9031 = pi90 & ~n9030;
  assign n9032 = n2519 & ~n9031;
  assign n9033 = n2488 & ~n8875;
  assign n9034 = pi58 & ~n9033;
  assign n9035 = pi53 & ~n8871;
  assign n9036 = ~pi60 & n8756;
  assign n9037 = n2705 & ~n9036;
  assign n9038 = ~n9035 & ~n9037;
  assign n9039 = n8873 & n9038;
  assign n9040 = n2488 & ~n9039;
  assign n9041 = ~pi58 & ~n9040;
  assign n9042 = ~n9034 & ~n9041;
  assign n9043 = ~pi90 & ~n9042;
  assign n9044 = n9032 & ~n9043;
  assign n9045 = ~pi111 & n2468;
  assign n9046 = ~pi68 & n2469;
  assign n9047 = ~pi36 & n9046;
  assign n9048 = n9045 & n9047;
  assign n9049 = pi73 & n9048;
  assign n9050 = ~pi102 & n8772;
  assign n9051 = n2467 & n9050;
  assign n9052 = n2465 & n8775;
  assign n9053 = n9051 & n9052;
  assign n9054 = n2821 & n9053;
  assign n9055 = n9049 & n9054;
  assign n9056 = n2493 & n9055;
  assign n9057 = ~n9038 & ~n9056;
  assign n9058 = n2488 & n9057;
  assign n9059 = n2706 & ~n9058;
  assign n9060 = n8872 & n9059;
  assign n9061 = n2488 & ~n9060;
  assign n9062 = ~pi58 & ~n9061;
  assign n9063 = ~pi90 & n9062;
  assign n9064 = n9044 & ~n9063;
  assign n9065 = n9028 & ~n9064;
  assign n9066 = ~n9026 & ~n9065;
  assign n9067 = ~pi51 & ~n9066;
  assign n9068 = pi51 & ~n2488;
  assign n9069 = n2506 & ~n9068;
  assign n9070 = ~n9067 & n9069;
  assign n9071 = ~n9024 & ~n9070;
  assign n9072 = ~pi40 & ~n9071;
  assign n9073 = ~pi32 & ~n9072;
  assign n9074 = ~n9023 & ~n9073;
  assign n9075 = ~pi95 & ~n9074;
  assign n9076 = ~n9022 & ~n9075;
  assign n9077 = ~pi96 & n7395;
  assign n9078 = n2900 & n9077;
  assign n9079 = n9029 & n9078;
  assign n9080 = n8862 & ~n9079;
  assign n9081 = pi32 & ~n9080;
  assign n9082 = ~n9073 & ~n9081;
  assign n9083 = ~pi95 & ~n9082;
  assign n9084 = ~pi198 & n9083;
  assign n9085 = n9076 & ~n9084;
  assign n9086 = ~n6190 & n9085;
  assign n9087 = n9028 & ~n9044;
  assign n9088 = ~n9026 & ~n9087;
  assign n9089 = ~pi51 & ~n9088;
  assign n9090 = n9069 & ~n9089;
  assign n9091 = ~n9024 & ~n9090;
  assign n9092 = ~pi40 & ~n9091;
  assign n9093 = ~pi32 & ~n9092;
  assign n9094 = ~n9081 & ~n9093;
  assign n9095 = ~pi95 & ~n9094;
  assign n9096 = ~pi198 & n9095;
  assign n9097 = n6190 & ~n9016;
  assign n9098 = ~n9023 & ~n9093;
  assign n9099 = ~pi95 & ~n9098;
  assign n9100 = n9097 & ~n9099;
  assign n9101 = ~n9096 & n9100;
  assign n9102 = ~n9086 & ~n9101;
  assign n9103 = ~pi183 & ~n9102;
  assign n9104 = ~pi40 & ~n9023;
  assign n9105 = n2488 & ~n2509;
  assign n9106 = ~pi32 & ~n9105;
  assign n9107 = pi93 & ~n2488;
  assign n9108 = n2509 & ~n9107;
  assign n9109 = n2488 & ~n9034;
  assign n9110 = ~pi90 & ~n9109;
  assign n9111 = ~n9031 & ~n9110;
  assign n9112 = ~pi93 & ~n9111;
  assign n9113 = n9108 & ~n9112;
  assign n9114 = n9106 & ~n9113;
  assign n9115 = n9104 & ~n9114;
  assign n9116 = ~pi95 & ~n9115;
  assign n9117 = n9097 & ~n9116;
  assign n9118 = ~n9086 & ~n9117;
  assign n9119 = pi183 & ~n9118;
  assign n9120 = ~n9103 & ~n9119;
  assign n9121 = ~pi95 & n9120;
  assign n9122 = ~pi174 & ~n9121;
  assign n9123 = ~n9022 & n9122;
  assign n9124 = n8781 & n9055;
  assign n9125 = ~pi90 & n9124;
  assign n9126 = n9111 & ~n9125;
  assign n9127 = ~pi93 & ~n9126;
  assign n9128 = n9108 & ~n9127;
  assign n9129 = n9106 & ~n9128;
  assign n9130 = n9104 & ~n9129;
  assign n9131 = ~pi95 & ~n9130;
  assign n9132 = ~n9022 & ~n9131;
  assign n9133 = n6190 & ~n9132;
  assign n9134 = pi183 & n9133;
  assign n9135 = pi183 & n6190;
  assign n9136 = ~n9085 & ~n9135;
  assign n9137 = pi174 & ~n9136;
  assign n9138 = ~n9134 & n9137;
  assign n9139 = ~pi180 & ~n9138;
  assign n9140 = ~n9123 & n9139;
  assign n9141 = ~pi40 & n6190;
  assign n9142 = ~n9016 & ~n9075;
  assign n9143 = ~n9084 & n9142;
  assign n9144 = n9141 & n9143;
  assign n9145 = ~n9086 & ~n9144;
  assign n9146 = ~pi183 & n9145;
  assign n9147 = n9097 & ~n9131;
  assign n9148 = ~n9086 & ~n9147;
  assign n9149 = pi183 & n9148;
  assign n9150 = ~n9146 & ~n9149;
  assign n9151 = pi174 & n9150;
  assign n9152 = ~pi174 & ~n9120;
  assign n9153 = pi180 & ~n9152;
  assign n9154 = ~n9151 & n9153;
  assign n9155 = ~n9140 & ~n9154;
  assign n9156 = ~pi193 & ~n9155;
  assign n9157 = n8781 & n9078;
  assign n9158 = ~pi32 & n9157;
  assign n9159 = n9055 & n9158;
  assign n9160 = n8862 & ~n9159;
  assign n9161 = ~pi95 & ~n9160;
  assign n9162 = n9097 & ~n9161;
  assign n9163 = ~n9086 & ~n9162;
  assign n9164 = pi183 & ~n9163;
  assign n9165 = ~pi40 & ~n2488;
  assign n9166 = pi32 & ~n9165;
  assign n9167 = n2462 & n2519;
  assign n9168 = ~n2488 & ~n9167;
  assign n9169 = n7394 & n9062;
  assign n9170 = ~n9168 & ~n9169;
  assign n9171 = ~pi70 & ~n9170;
  assign n9172 = ~n9026 & ~n9171;
  assign n9173 = ~pi51 & ~n9172;
  assign n9174 = n9069 & ~n9173;
  assign n9175 = ~pi40 & ~n9174;
  assign n9176 = ~n9024 & n9175;
  assign n9177 = ~pi32 & ~n9176;
  assign n9178 = ~n9166 & ~n9177;
  assign n9179 = ~n2515 & ~n8862;
  assign n9180 = ~n9178 & ~n9179;
  assign n9181 = ~pi95 & ~n9180;
  assign n9182 = ~n9016 & ~n9181;
  assign n9183 = pi95 & ~n9165;
  assign n9184 = ~pi40 & ~n9080;
  assign n9185 = pi32 & ~n9184;
  assign n9186 = ~n9177 & ~n9185;
  assign n9187 = ~pi95 & ~n9186;
  assign n9188 = ~n9183 & ~n9187;
  assign n9189 = n9182 & ~n9188;
  assign n9190 = ~pi198 & ~n9189;
  assign n9191 = n6190 & ~n9190;
  assign n9192 = n9182 & n9191;
  assign n9193 = ~n9086 & ~n9192;
  assign n9194 = ~pi183 & ~n9193;
  assign n9195 = pi174 & ~n9194;
  assign n9196 = ~n9164 & n9195;
  assign n9197 = n6190 & ~n8862;
  assign n9198 = ~n6190 & ~n9085;
  assign n9199 = ~n9197 & ~n9198;
  assign n9200 = pi183 & n9199;
  assign n9201 = n7394 & n9041;
  assign n9202 = ~n9168 & ~n9201;
  assign n9203 = ~pi70 & ~n9202;
  assign n9204 = ~n9026 & ~n9203;
  assign n9205 = ~pi51 & ~n9204;
  assign n9206 = n9069 & ~n9205;
  assign n9207 = ~n9024 & ~n9206;
  assign n9208 = ~pi40 & n9207;
  assign n9209 = ~pi32 & ~n9208;
  assign n9210 = ~n9166 & ~n9209;
  assign n9211 = ~pi95 & ~n9210;
  assign n9212 = ~n9183 & ~n9211;
  assign n9213 = pi198 & ~n9212;
  assign n9214 = ~n9185 & ~n9209;
  assign n9215 = ~pi95 & ~n9214;
  assign n9216 = ~n9183 & ~n9215;
  assign n9217 = ~pi198 & ~n9216;
  assign n9218 = ~n9213 & ~n9217;
  assign n9219 = n9141 & ~n9218;
  assign n9220 = ~n9086 & ~n9219;
  assign n9221 = ~pi183 & ~n9220;
  assign n9222 = ~pi174 & ~n9221;
  assign n9223 = ~n9200 & n9222;
  assign n9224 = pi180 & ~n9223;
  assign n9225 = ~n9196 & n9224;
  assign n9226 = ~pi40 & ~n9207;
  assign n9227 = ~pi32 & ~n9226;
  assign n9228 = ~n9023 & ~n9227;
  assign n9229 = ~pi95 & ~n9228;
  assign n9230 = ~n9022 & ~n9229;
  assign n9231 = ~n9081 & ~n9227;
  assign n9232 = ~pi95 & ~n9231;
  assign n9233 = ~pi198 & n9232;
  assign n9234 = n9230 & ~n9233;
  assign n9235 = n6190 & ~n9234;
  assign n9236 = ~n9198 & ~n9235;
  assign n9237 = ~pi183 & n9236;
  assign n9238 = ~pi95 & ~n8862;
  assign n9239 = ~n9022 & ~n9238;
  assign n9240 = n6190 & n9239;
  assign n9241 = ~n9086 & ~n9240;
  assign n9242 = pi183 & ~n9241;
  assign n9243 = ~pi174 & ~n9242;
  assign n9244 = ~n9237 & n9243;
  assign n9245 = n6190 & ~n9022;
  assign n9246 = ~n9161 & n9245;
  assign n9247 = ~n9086 & ~n9246;
  assign n9248 = pi183 & ~n9247;
  assign n9249 = ~n9022 & ~n9181;
  assign n9250 = ~n9191 & ~n9197;
  assign n9251 = n9249 & ~n9250;
  assign n9252 = ~n9086 & ~n9251;
  assign n9253 = ~pi183 & ~n9252;
  assign n9254 = ~n9248 & ~n9253;
  assign n9255 = pi174 & n9254;
  assign n9256 = ~pi180 & ~n9255;
  assign n9257 = ~n9244 & n9256;
  assign n9258 = pi193 & ~n9257;
  assign n9259 = ~n9225 & n9258;
  assign n9260 = ~n9156 & ~n9259;
  assign n9261 = ~pi299 & ~n9260;
  assign n9262 = pi158 & pi299;
  assign n9263 = ~pi210 & n9083;
  assign n9264 = n9076 & ~n9263;
  assign n9265 = ~n6190 & ~n9264;
  assign n9266 = n9142 & ~n9263;
  assign n9267 = n6190 & ~n9266;
  assign n9268 = ~n9265 & ~n9267;
  assign n9269 = pi152 & n9268;
  assign n9270 = ~n6190 & n9264;
  assign n9271 = ~pi210 & n9095;
  assign n9272 = n9100 & ~n9271;
  assign n9273 = ~n9270 & ~n9272;
  assign n9274 = ~pi152 & ~n9273;
  assign n9275 = ~pi172 & ~n9274;
  assign n9276 = ~n9269 & n9275;
  assign n9277 = ~pi210 & ~n9189;
  assign n9278 = n6190 & ~n9277;
  assign n9279 = n9182 & n9278;
  assign n9280 = ~n9270 & ~n9279;
  assign n9281 = pi152 & ~n9280;
  assign n9282 = ~pi210 & ~n9216;
  assign n9283 = pi210 & ~n9212;
  assign n9284 = ~n9282 & ~n9283;
  assign n9285 = n9141 & ~n9284;
  assign n9286 = ~n9270 & ~n9285;
  assign n9287 = ~pi152 & ~n9286;
  assign n9288 = pi172 & ~n9287;
  assign n9289 = ~n9281 & n9288;
  assign n9290 = ~n9276 & ~n9289;
  assign n9291 = n9262 & ~n9290;
  assign n9292 = ~pi158 & pi299;
  assign n9293 = ~n9022 & ~n9099;
  assign n9294 = ~n9271 & n9293;
  assign n9295 = n6190 & n9294;
  assign n9296 = ~pi152 & ~n9295;
  assign n9297 = pi152 & ~n9264;
  assign n9298 = ~pi172 & ~n9297;
  assign n9299 = ~n9296 & n9298;
  assign n9300 = n9292 & ~n9299;
  assign n9301 = ~n9197 & ~n9278;
  assign n9302 = n9249 & ~n9301;
  assign n9303 = pi152 & ~n9302;
  assign n9304 = ~n9197 & ~n9285;
  assign n9305 = n9230 & ~n9304;
  assign n9306 = ~pi152 & ~n9305;
  assign n9307 = pi172 & ~n9306;
  assign n9308 = ~n9303 & n9307;
  assign n9309 = ~n9270 & ~n9308;
  assign n9310 = n9300 & n9309;
  assign n9311 = ~pi149 & ~n9310;
  assign n9312 = ~n9291 & n9311;
  assign n9313 = ~n9240 & ~n9270;
  assign n9314 = ~pi152 & ~n9313;
  assign n9315 = ~n9246 & ~n9270;
  assign n9316 = pi152 & ~n9315;
  assign n9317 = pi172 & ~n9316;
  assign n9318 = ~n9314 & n9317;
  assign n9319 = ~n9133 & ~n9265;
  assign n9320 = pi152 & n9319;
  assign n9321 = ~n9022 & ~n9116;
  assign n9322 = n6190 & ~n9321;
  assign n9323 = ~n9265 & ~n9322;
  assign n9324 = ~pi152 & n9323;
  assign n9325 = ~pi172 & ~n9324;
  assign n9326 = ~n9320 & n9325;
  assign n9327 = ~n9318 & ~n9326;
  assign n9328 = n9292 & ~n9327;
  assign n9329 = ~n9117 & ~n9270;
  assign n9330 = ~pi152 & ~n9329;
  assign n9331 = ~n9147 & ~n9270;
  assign n9332 = pi152 & ~n9331;
  assign n9333 = ~pi172 & ~n9332;
  assign n9334 = ~n9330 & n9333;
  assign n9335 = ~n9197 & ~n9265;
  assign n9336 = ~pi152 & n9335;
  assign n9337 = ~n9162 & ~n9270;
  assign n9338 = pi152 & ~n9337;
  assign n9339 = pi172 & ~n9338;
  assign n9340 = ~n9336 & n9339;
  assign n9341 = ~n9334 & ~n9340;
  assign n9342 = n9262 & ~n9341;
  assign n9343 = pi149 & ~n9342;
  assign n9344 = ~n9328 & n9343;
  assign n9345 = ~n9312 & ~n9344;
  assign n9346 = ~n9261 & ~n9345;
  assign n9347 = pi232 & ~n9346;
  assign n9348 = ~n6166 & n9083;
  assign n9349 = n9076 & ~n9348;
  assign n9350 = ~pi232 & ~n9349;
  assign n9351 = ~pi39 & ~n9350;
  assign n9352 = ~n9347 & n9351;
  assign n9353 = ~n9015 & ~n9352;
  assign n9354 = ~pi38 & ~n9353;
  assign n9355 = ~n8958 & ~n9354;
  assign n9356 = ~pi100 & ~n9355;
  assign n9357 = ~pi87 & ~n8912;
  assign n9358 = ~n9356 & n9357;
  assign n9359 = n8946 & ~n9358;
  assign n9360 = ~n8943 & ~n9359;
  assign n9361 = ~n8913 & n9360;
  assign n9362 = ~pi54 & ~n9361;
  assign n9363 = ~n8929 & ~n9362;
  assign n9364 = ~pi74 & ~n9363;
  assign n9365 = n8922 & ~n9364;
  assign n9366 = ~n8903 & ~n9365;
  assign n9367 = n2531 & n9366;
  assign n9368 = ~n8866 & ~n9367;
  assign n9369 = n8861 & n9368;
  assign n9370 = ~n8853 & ~n9369;
  assign n9371 = ~n8835 & ~n9370;
  assign n9372 = pi87 & ~n8931;
  assign n9373 = ~pi176 & pi232;
  assign n9374 = n6237 & n6448;
  assign n9375 = n8973 & n9374;
  assign n9376 = ~pi174 & n9375;
  assign n9377 = ~pi299 & ~n9376;
  assign n9378 = n9373 & ~n9377;
  assign n9379 = pi176 & pi232;
  assign n9380 = n6237 & ~n6456;
  assign n9381 = n8973 & n9380;
  assign n9382 = ~pi174 & n9381;
  assign n9383 = n6190 & n7463;
  assign n9384 = ~n6236 & n8973;
  assign n9385 = n9383 & n9384;
  assign n9386 = pi174 & n9385;
  assign n9387 = ~pi299 & ~n9386;
  assign n9388 = ~n9382 & n9387;
  assign n9389 = n9379 & ~n9388;
  assign n9390 = ~n9378 & ~n9389;
  assign n9391 = n6199 & ~n6456;
  assign n9392 = pi154 & ~n9391;
  assign n9393 = n6199 & n6448;
  assign n9394 = ~pi154 & ~n9393;
  assign n9395 = ~pi152 & ~n9394;
  assign n9396 = ~n9392 & n9395;
  assign n9397 = ~n6198 & n9383;
  assign n9398 = pi152 & pi154;
  assign n9399 = n9397 & n9398;
  assign n9400 = ~n9396 & ~n9399;
  assign n9401 = n8959 & ~n9400;
  assign n9402 = pi299 & ~n9401;
  assign n9403 = pi39 & ~n9402;
  assign n9404 = ~n9390 & n9403;
  assign n9405 = ~pi93 & n2509;
  assign n9406 = ~pi90 & n6135;
  assign n9407 = ~n7383 & ~n9406;
  assign n9408 = n9405 & ~n9407;
  assign n9409 = n2516 & n6190;
  assign n9410 = ~pi40 & n9409;
  assign n9411 = n9408 & n9410;
  assign n9412 = n2488 & n9124;
  assign n9413 = n9078 & n9412;
  assign n9414 = ~n9408 & ~n9413;
  assign n9415 = n9410 & ~n9414;
  assign n9416 = ~pi152 & n9415;
  assign n9417 = ~n9411 & ~n9416;
  assign n9418 = pi172 & ~n9417;
  assign n9419 = n2516 & n9413;
  assign n9420 = n9141 & n9419;
  assign n9421 = ~pi152 & ~pi172;
  assign n9422 = n9420 & n9421;
  assign n9423 = ~n9418 & ~n9422;
  assign n9424 = ~pi149 & ~n9423;
  assign n9425 = n6190 & n6306;
  assign n9426 = pi158 & n9425;
  assign n9427 = n3078 & n3085;
  assign n9428 = n2709 & n2712;
  assign n9429 = n7394 & n9428;
  assign n9430 = n2488 & n9429;
  assign n9431 = n9059 & n9430;
  assign n9432 = ~pi70 & ~n9431;
  assign n9433 = n9427 & ~n9432;
  assign n9434 = ~n6418 & ~n9433;
  assign n9435 = n2519 & ~n9407;
  assign n9436 = n9432 & ~n9435;
  assign n9437 = n9427 & ~n9436;
  assign n9438 = pi172 & n9437;
  assign n9439 = ~pi152 & ~n9438;
  assign n9440 = n9434 & n9439;
  assign n9441 = pi149 & n6190;
  assign n9442 = ~n9037 & n9429;
  assign n9443 = ~pi70 & ~n9442;
  assign n9444 = ~n9435 & n9443;
  assign n9445 = n9427 & ~n9444;
  assign n9446 = pi172 & n9445;
  assign n9447 = n9427 & ~n9443;
  assign n9448 = ~n6418 & ~n9447;
  assign n9449 = pi152 & n9448;
  assign n9450 = ~n9446 & n9449;
  assign n9451 = n9441 & ~n9450;
  assign n9452 = ~n9440 & n9451;
  assign n9453 = pi299 & ~n9452;
  assign n9454 = ~n9426 & n9453;
  assign n9455 = ~n9424 & n9454;
  assign n9456 = ~pi39 & pi232;
  assign n9457 = ~n6374 & ~n9433;
  assign n9458 = ~pi198 & ~n9457;
  assign n9459 = ~n9437 & ~n9458;
  assign n9460 = n9135 & ~n9459;
  assign n9461 = ~pi183 & n9415;
  assign n9462 = ~pi174 & ~n9461;
  assign n9463 = ~n9460 & n9462;
  assign n9464 = ~pi183 & n9411;
  assign n9465 = pi174 & ~n9464;
  assign n9466 = ~n6375 & ~n9445;
  assign n9467 = n6190 & ~n9466;
  assign n9468 = pi183 & n9467;
  assign n9469 = n9465 & ~n9468;
  assign n9470 = ~n9463 & ~n9469;
  assign n9471 = pi193 & ~n9470;
  assign n9472 = ~n6375 & ~n9447;
  assign n9473 = pi174 & n9472;
  assign n9474 = ~n6375 & ~n9433;
  assign n9475 = ~pi174 & n9474;
  assign n9476 = ~n9473 & ~n9475;
  assign n9477 = n9135 & n9476;
  assign n9478 = ~pi174 & n9420;
  assign n9479 = ~pi183 & n9478;
  assign n9480 = ~pi193 & ~n9479;
  assign n9481 = ~n9477 & n9480;
  assign n9482 = ~n9471 & ~n9481;
  assign n9483 = pi180 & n9425;
  assign n9484 = ~pi299 & ~n9483;
  assign n9485 = ~n9482 & n9484;
  assign n9486 = n9456 & ~n9485;
  assign n9487 = ~n9455 & n9486;
  assign n9488 = ~n9404 & ~n9487;
  assign n9489 = ~pi38 & ~n9488;
  assign n9490 = ~pi87 & ~n8958;
  assign n9491 = ~n9489 & n9490;
  assign n9492 = ~pi100 & ~n9491;
  assign n9493 = ~n9372 & n9492;
  assign n9494 = ~n8912 & ~n9493;
  assign n9495 = n2573 & ~n9494;
  assign n9496 = n2572 & n8938;
  assign n9497 = n6132 & n9496;
  assign n9498 = n8933 & ~n9497;
  assign n9499 = n8930 & ~n9498;
  assign n9500 = ~n8913 & ~n9499;
  assign n9501 = ~n9495 & n9500;
  assign n9502 = ~pi54 & ~n9501;
  assign n9503 = ~n8929 & ~n9502;
  assign n9504 = ~pi74 & ~n9503;
  assign n9505 = n8922 & ~n9504;
  assign n9506 = n6132 & n8880;
  assign n9507 = ~pi38 & ~n9506;
  assign n9508 = n8887 & ~n9507;
  assign n9509 = pi38 & pi87;
  assign n9510 = n8886 & n9509;
  assign n9511 = ~n8842 & ~n9510;
  assign n9512 = ~n9508 & n9511;
  assign n9513 = ~pi75 & ~n9512;
  assign n9514 = n8868 & ~n9513;
  assign n9515 = pi92 & n8856;
  assign n9516 = ~pi54 & ~n9515;
  assign n9517 = ~n9514 & n9516;
  assign n9518 = ~n8854 & ~n9517;
  assign n9519 = ~pi74 & ~n9518;
  assign n9520 = n8867 & ~n9519;
  assign n9521 = ~n9505 & ~n9520;
  assign n9522 = n2531 & n9521;
  assign n9523 = n8861 & ~n9522;
  assign n9524 = ~n8853 & ~n9523;
  assign n9525 = n8835 & ~n9524;
  assign n9526 = ~pi954 & ~n9525;
  assign n9527 = ~n9371 & n9526;
  assign n9528 = ~pi33 & ~n9370;
  assign n9529 = pi33 & ~n9524;
  assign n9530 = pi954 & ~n9529;
  assign n9531 = ~n9528 & n9530;
  assign po191 = ~n9527 & ~n9531;
  assign n9533 = ~pi33 & ~pi954;
  assign n9534 = pi197 & n8837;
  assign n9535 = ~pi197 & ~n8837;
  assign n9536 = ~n9534 & ~n9535;
  assign n9537 = pi162 & n6190;
  assign n9538 = n9536 & ~n9537;
  assign n9539 = n9534 & n9537;
  assign n9540 = ~pi162 & ~pi197;
  assign n9541 = n8838 & ~n9540;
  assign n9542 = n6190 & ~n9541;
  assign n9543 = ~n9539 & n9542;
  assign n9544 = ~n9536 & ~n9543;
  assign n9545 = ~n9538 & ~n9544;
  assign n9546 = pi232 & ~n7255;
  assign n9547 = n9545 & n9546;
  assign n9548 = pi167 & n8915;
  assign n9549 = ~n9547 & ~n9548;
  assign n9550 = ~pi74 & n9549;
  assign n9551 = pi74 & ~n9547;
  assign n9552 = pi148 & n8915;
  assign n9553 = n9551 & ~n9552;
  assign n9554 = ~n9550 & ~n9553;
  assign n9555 = ~n3327 & n9554;
  assign n9556 = ~pi54 & ~n9547;
  assign n9557 = pi38 & n9548;
  assign n9558 = n9556 & ~n9557;
  assign n9559 = ~pi74 & n9558;
  assign n9560 = n9554 & ~n9559;
  assign n9561 = ~n2531 & ~n9560;
  assign n9562 = n3327 & ~n9561;
  assign n9563 = ~n2531 & ~n8865;
  assign n9564 = n3327 & ~n9563;
  assign n9565 = ~n9562 & ~n9564;
  assign n9566 = pi299 & ~n9545;
  assign n9567 = pi140 & pi145;
  assign n9568 = n8905 & ~n9567;
  assign n9569 = ~pi140 & ~pi145;
  assign n9570 = n6190 & ~n9569;
  assign n9571 = n9568 & n9570;
  assign n9572 = ~n9567 & ~n9569;
  assign n9573 = n8906 & ~n9572;
  assign n9574 = ~pi299 & ~n9573;
  assign n9575 = ~n9571 & n9574;
  assign n9576 = pi232 & ~n9575;
  assign n9577 = ~n9566 & n9576;
  assign n9578 = pi100 & ~n9577;
  assign n9579 = pi75 & ~n9577;
  assign n9580 = ~n9578 & ~n9579;
  assign n9581 = pi141 & ~pi299;
  assign n9582 = pi148 & pi299;
  assign n9583 = ~n9581 & ~n9582;
  assign n9584 = n7420 & ~n9583;
  assign n9585 = n7255 & ~n9584;
  assign n9586 = n9580 & ~n9585;
  assign n9587 = pi74 & ~n9586;
  assign n9588 = ~pi55 & ~n9587;
  assign n9589 = pi188 & ~pi299;
  assign n9590 = pi167 & pi299;
  assign n9591 = ~n9589 & ~n9590;
  assign n9592 = n7420 & ~n9591;
  assign n9593 = ~pi100 & ~n9592;
  assign n9594 = ~pi75 & n9593;
  assign n9595 = n9580 & ~n9594;
  assign n9596 = pi54 & ~n9595;
  assign n9597 = pi38 & ~n9592;
  assign n9598 = ~n8889 & ~n9597;
  assign n9599 = pi87 & n9598;
  assign n9600 = pi167 & ~n8950;
  assign n9601 = pi188 & n9600;
  assign n9602 = ~pi188 & ~n8948;
  assign n9603 = pi188 & n8954;
  assign n9604 = ~pi167 & ~n9603;
  assign n9605 = ~n9602 & ~n9604;
  assign n9606 = ~n9601 & n9605;
  assign n9607 = pi38 & ~n9606;
  assign n9608 = ~pi142 & ~n9252;
  assign n9609 = pi142 & n9085;
  assign n9610 = ~pi140 & ~n9609;
  assign n9611 = ~n9608 & n9610;
  assign n9612 = ~pi142 & ~n9247;
  assign n9613 = pi140 & ~n9612;
  assign n9614 = ~n9133 & ~n9198;
  assign n9615 = pi142 & n9614;
  assign n9616 = n9613 & ~n9615;
  assign n9617 = ~n9611 & ~n9616;
  assign n9618 = ~pi181 & ~n9617;
  assign n9619 = ~pi142 & ~n9193;
  assign n9620 = pi142 & ~n9145;
  assign n9621 = ~pi140 & ~n9620;
  assign n9622 = ~n9619 & n9621;
  assign n9623 = ~pi142 & ~n9163;
  assign n9624 = pi142 & ~n9148;
  assign n9625 = pi140 & ~n9624;
  assign n9626 = ~n9623 & n9625;
  assign n9627 = ~n9622 & ~n9626;
  assign n9628 = pi181 & ~n9627;
  assign n9629 = pi144 & ~n9628;
  assign n9630 = ~n9618 & n9629;
  assign n9631 = ~pi142 & ~n9220;
  assign n9632 = pi142 & ~n9102;
  assign n9633 = ~pi140 & ~n9632;
  assign n9634 = ~n9631 & n9633;
  assign n9635 = pi142 & ~n9118;
  assign n9636 = ~pi142 & n9199;
  assign n9637 = pi140 & ~n9636;
  assign n9638 = ~n9635 & n9637;
  assign n9639 = ~n9634 & ~n9638;
  assign n9640 = pi181 & ~n9639;
  assign n9641 = ~pi142 & n9236;
  assign n9642 = ~pi140 & ~n9641;
  assign n9643 = ~n9096 & n9293;
  assign n9644 = n6190 & ~n9643;
  assign n9645 = ~n9198 & ~n9644;
  assign n9646 = pi142 & n9645;
  assign n9647 = n9642 & ~n9646;
  assign n9648 = ~pi142 & ~n9241;
  assign n9649 = pi140 & ~n9648;
  assign n9650 = ~n9198 & ~n9322;
  assign n9651 = pi142 & n9650;
  assign n9652 = n9649 & ~n9651;
  assign n9653 = ~n9647 & ~n9652;
  assign n9654 = ~pi181 & ~n9653;
  assign n9655 = ~pi144 & ~n9654;
  assign n9656 = ~n9640 & n9655;
  assign n9657 = ~pi299 & ~n9656;
  assign n9658 = ~n9630 & n9657;
  assign n9659 = ~pi159 & pi299;
  assign n9660 = ~pi146 & ~n9313;
  assign n9661 = pi146 & n9323;
  assign n9662 = ~pi161 & ~n9661;
  assign n9663 = ~n9660 & n9662;
  assign n9664 = ~pi146 & ~n9315;
  assign n9665 = pi146 & n9319;
  assign n9666 = pi161 & ~n9665;
  assign n9667 = ~n9664 & n9666;
  assign n9668 = ~n9663 & ~n9667;
  assign n9669 = pi162 & ~n9668;
  assign n9670 = ~pi161 & ~n9295;
  assign n9671 = pi161 & ~n9264;
  assign n9672 = ~n9670 & ~n9671;
  assign n9673 = pi146 & n9672;
  assign n9674 = ~pi162 & ~n9673;
  assign n9675 = ~pi161 & ~n9305;
  assign n9676 = pi161 & ~n9302;
  assign n9677 = ~pi146 & ~n9676;
  assign n9678 = ~n9675 & n9677;
  assign n9679 = n9674 & ~n9678;
  assign n9680 = ~n9270 & n9679;
  assign n9681 = ~n9669 & ~n9680;
  assign n9682 = n9659 & ~n9681;
  assign n9683 = ~pi146 & ~n9280;
  assign n9684 = pi146 & n9268;
  assign n9685 = ~n9683 & ~n9684;
  assign n9686 = pi161 & n9685;
  assign n9687 = ~pi146 & ~n9286;
  assign n9688 = pi146 & ~n9273;
  assign n9689 = ~pi161 & ~n9688;
  assign n9690 = ~n9687 & n9689;
  assign n9691 = ~pi162 & ~n9690;
  assign n9692 = ~n9686 & n9691;
  assign n9693 = pi159 & pi299;
  assign n9694 = ~pi146 & ~n9337;
  assign n9695 = pi146 & ~n9331;
  assign n9696 = pi161 & ~n9695;
  assign n9697 = ~n9694 & n9696;
  assign n9698 = pi146 & ~n9329;
  assign n9699 = ~pi146 & n9335;
  assign n9700 = ~pi161 & ~n9699;
  assign n9701 = ~n9698 & n9700;
  assign n9702 = pi162 & ~n9701;
  assign n9703 = ~n9697 & n9702;
  assign n9704 = n9693 & ~n9703;
  assign n9705 = ~n9692 & n9704;
  assign n9706 = ~n9682 & ~n9705;
  assign n9707 = ~n9658 & n9706;
  assign n9708 = pi232 & ~n9707;
  assign n9709 = ~n9350 & ~n9708;
  assign n9710 = n2532 & ~n9709;
  assign n9711 = ~pi177 & ~pi299;
  assign n9712 = ~pi144 & ~n8975;
  assign n9713 = ~n9002 & ~n9712;
  assign n9714 = ~n9010 & ~n9713;
  assign n9715 = n9711 & ~n9714;
  assign n9716 = pi177 & ~pi299;
  assign n9717 = n9713 & n9716;
  assign n9718 = ~n9715 & ~n9717;
  assign n9719 = pi232 & ~n9718;
  assign n9720 = ~n8981 & ~n9719;
  assign n9721 = ~pi38 & ~n9720;
  assign n9722 = ~pi161 & n8991;
  assign n9723 = ~n8971 & ~n9722;
  assign n9724 = n8959 & ~n9723;
  assign n9725 = ~pi38 & ~pi155;
  assign n9726 = ~n9724 & n9725;
  assign n9727 = ~pi38 & pi155;
  assign n9728 = pi161 & n8984;
  assign n9729 = n8959 & ~n9728;
  assign n9730 = n8967 & n9729;
  assign n9731 = n9727 & ~n9730;
  assign n9732 = ~n9726 & ~n9731;
  assign n9733 = pi232 & ~n9732;
  assign n9734 = n8961 & n9733;
  assign n9735 = ~n9721 & ~n9734;
  assign n9736 = pi39 & ~n9735;
  assign n9737 = ~pi87 & ~n9736;
  assign n9738 = ~n9710 & n9737;
  assign n9739 = ~n9607 & n9738;
  assign n9740 = ~pi100 & ~n9739;
  assign n9741 = ~n9599 & n9740;
  assign n9742 = ~n9578 & ~n9741;
  assign n9743 = n2573 & ~n9742;
  assign n9744 = pi155 & pi299;
  assign n9745 = ~n9716 & ~n9744;
  assign n9746 = ~pi38 & n9745;
  assign n9747 = n7420 & ~n9746;
  assign n9748 = n8934 & ~n9747;
  assign n9749 = n9598 & ~n9748;
  assign n9750 = ~pi100 & ~n9749;
  assign n9751 = ~n9578 & ~n9750;
  assign n9752 = n8930 & ~n9751;
  assign n9753 = ~n9579 & ~n9752;
  assign n9754 = ~n9743 & n9753;
  assign n9755 = ~pi54 & ~n9754;
  assign n9756 = ~n9596 & ~n9755;
  assign n9757 = ~pi74 & ~n9756;
  assign n9758 = n9588 & ~n9757;
  assign n9759 = pi55 & ~n9553;
  assign n9760 = pi54 & n9549;
  assign n9761 = ~n8864 & n9558;
  assign n9762 = ~n6094 & ~n9761;
  assign n9763 = pi232 & n9545;
  assign n9764 = pi100 & ~n9763;
  assign n9765 = pi167 & n7420;
  assign n9766 = pi38 & n9765;
  assign n9767 = n8934 & ~n9537;
  assign n9768 = n8863 & ~n9767;
  assign n9769 = ~pi100 & ~n9768;
  assign n9770 = ~pi232 & n8934;
  assign n9771 = ~n9769 & ~n9770;
  assign n9772 = ~n9766 & ~n9771;
  assign n9773 = ~n9764 & ~n9772;
  assign n9774 = ~pi75 & ~n9773;
  assign n9775 = pi75 & ~n9763;
  assign n9776 = ~pi92 & ~n9775;
  assign n9777 = ~n9774 & n9776;
  assign n9778 = ~n9762 & ~n9777;
  assign n9779 = ~n9760 & ~n9778;
  assign n9780 = ~pi74 & ~n9779;
  assign n9781 = n9759 & ~n9780;
  assign n9782 = n2531 & ~n9781;
  assign n9783 = ~n9758 & n9782;
  assign n9784 = ~n9565 & ~n9783;
  assign n9785 = ~n9555 & ~n9784;
  assign n9786 = ~pi34 & n9785;
  assign n9787 = ~n9533 & ~n9786;
  assign n9788 = pi161 & ~n9397;
  assign n9789 = ~pi161 & ~n9391;
  assign n9790 = ~n9788 & ~n9789;
  assign n9791 = n8959 & n9790;
  assign n9792 = n9727 & ~n9791;
  assign n9793 = ~pi161 & n8959;
  assign n9794 = n9393 & n9793;
  assign n9795 = n9725 & ~n9794;
  assign n9796 = ~n9792 & ~n9795;
  assign n9797 = pi299 & ~n9796;
  assign n9798 = ~pi144 & n9375;
  assign n9799 = n9711 & ~n9798;
  assign n9800 = ~pi144 & n9381;
  assign n9801 = pi144 & n9385;
  assign n9802 = n9716 & ~n9801;
  assign n9803 = ~n9800 & n9802;
  assign n9804 = ~n9799 & ~n9803;
  assign n9805 = pi232 & n9804;
  assign n9806 = ~pi38 & ~n9805;
  assign n9807 = ~n9797 & ~n9806;
  assign n9808 = pi39 & ~n9807;
  assign n9809 = ~pi142 & n9411;
  assign n9810 = ~pi140 & ~n9809;
  assign n9811 = ~pi142 & n9445;
  assign n9812 = pi140 & ~n9811;
  assign n9813 = n9472 & n9812;
  assign n9814 = ~n9810 & ~n9813;
  assign n9815 = pi144 & ~n9814;
  assign n9816 = pi140 & ~n6190;
  assign n9817 = ~n9420 & n9810;
  assign n9818 = ~pi142 & n9437;
  assign n9819 = pi140 & ~n9818;
  assign n9820 = n9474 & n9819;
  assign n9821 = ~n9817 & ~n9820;
  assign n9822 = ~pi144 & ~n9821;
  assign n9823 = ~n9816 & ~n9822;
  assign n9824 = ~n9815 & n9823;
  assign n9825 = pi181 & n9425;
  assign n9826 = ~pi299 & ~n9825;
  assign n9827 = ~n9824 & n9826;
  assign n9828 = ~pi146 & ~n9415;
  assign n9829 = pi146 & ~n9420;
  assign n9830 = ~pi161 & ~n9829;
  assign n9831 = ~n9828 & n9830;
  assign n9832 = ~pi146 & pi161;
  assign n9833 = n9411 & n9832;
  assign n9834 = ~n9831 & ~n9833;
  assign n9835 = ~pi162 & ~n9834;
  assign n9836 = ~pi146 & n9445;
  assign n9837 = n9448 & ~n9836;
  assign n9838 = pi161 & ~n9837;
  assign n9839 = pi159 & n6306;
  assign n9840 = ~pi146 & n9437;
  assign n9841 = n9434 & ~n9840;
  assign n9842 = ~pi161 & ~n9841;
  assign n9843 = pi299 & ~n9842;
  assign n9844 = ~n9839 & n9843;
  assign n9845 = ~n9838 & n9844;
  assign n9846 = pi159 & n9425;
  assign n9847 = ~n9537 & ~n9846;
  assign n9848 = pi299 & n9847;
  assign n9849 = ~n9845 & ~n9848;
  assign n9850 = ~n9835 & ~n9849;
  assign n9851 = pi232 & ~n9850;
  assign n9852 = ~n9827 & n9851;
  assign n9853 = n2532 & ~n9852;
  assign n9854 = ~n9607 & ~n9853;
  assign n9855 = ~n9808 & n9854;
  assign n9856 = ~pi100 & ~n9855;
  assign n9857 = ~n9578 & ~n9856;
  assign n9858 = ~pi87 & ~n9857;
  assign n9859 = ~n2614 & ~n9593;
  assign n9860 = ~n9578 & n9859;
  assign n9861 = pi87 & ~n9860;
  assign n9862 = ~n9858 & ~n9861;
  assign n9863 = n2573 & ~n9862;
  assign n9864 = pi38 & ~n9591;
  assign n9865 = n2532 & ~n9745;
  assign n9866 = n2512 & n9865;
  assign n9867 = ~n9864 & ~n9866;
  assign n9868 = n7420 & ~n9867;
  assign n9869 = ~pi100 & ~n9868;
  assign n9870 = ~n9578 & ~n9869;
  assign n9871 = ~pi87 & ~n9870;
  assign n9872 = ~n9861 & ~n9871;
  assign n9873 = n8930 & ~n9872;
  assign n9874 = ~n9579 & ~n9873;
  assign n9875 = ~n9863 & n9874;
  assign n9876 = ~pi54 & ~n9875;
  assign n9877 = ~n9596 & ~n9876;
  assign n9878 = ~pi74 & ~n9877;
  assign n9879 = n9588 & ~n9878;
  assign n9880 = ~pi92 & n9456;
  assign n9881 = pi162 & n9880;
  assign n9882 = n7254 & n9881;
  assign n9883 = n6222 & n9882;
  assign n9884 = ~n9766 & ~n9883;
  assign n9885 = n7255 & ~n9884;
  assign n9886 = n9556 & ~n9885;
  assign n9887 = ~n9760 & ~n9886;
  assign n9888 = ~pi74 & ~n9887;
  assign n9889 = n9759 & ~n9888;
  assign n9890 = ~n9879 & ~n9889;
  assign n9891 = n2531 & n9890;
  assign n9892 = n9562 & ~n9891;
  assign n9893 = ~n9555 & ~n9892;
  assign n9894 = pi34 & n9893;
  assign n9895 = n9787 & ~n9894;
  assign n9896 = ~pi34 & ~n8833;
  assign n9897 = n9785 & ~n9896;
  assign n9898 = n9893 & n9896;
  assign n9899 = n9533 & ~n9898;
  assign n9900 = ~n9897 & n9899;
  assign po192 = ~n9895 & ~n9900;
  assign n9902 = pi137 & n8741;
  assign n9903 = ~n6211 & n7368;
  assign n9904 = pi683 & n9903;
  assign n9905 = pi252 & po1057;
  assign n9906 = ~n9904 & n9905;
  assign n9907 = ~n6106 & ~n9906;
  assign n9908 = ~n7421 & ~n9907;
  assign n9909 = ~n8746 & ~n9908;
  assign n9910 = n8743 & n9909;
  assign n9911 = ~n9902 & ~n9910;
  assign n9912 = n8740 & ~n9911;
  assign n9913 = pi38 & ~n8817;
  assign n9914 = pi35 & ~n2916;
  assign n9915 = n2919 & ~n9914;
  assign n9916 = ~pi93 & ~n9406;
  assign n9917 = ~n6154 & ~n9916;
  assign n9918 = ~pi35 & ~n9917;
  assign n9919 = n9915 & ~n9918;
  assign n9920 = ~n2737 & ~n9919;
  assign n9921 = pi1082 & ~n9920;
  assign n9922 = n2516 & n9921;
  assign n9923 = n2696 & n8786;
  assign n9924 = n9918 & ~n9923;
  assign n9925 = n2516 & ~n9924;
  assign n9926 = n6166 & ~n9918;
  assign n9927 = ~pi122 & ~po740;
  assign n9928 = n7376 & ~n9927;
  assign n9929 = n2978 & n7404;
  assign n9930 = ~n7376 & ~n9929;
  assign n9931 = ~pi137 & ~n6166;
  assign n9932 = ~n9930 & ~n9931;
  assign n9933 = ~n9928 & n9932;
  assign n9934 = ~n9926 & ~n9933;
  assign n9935 = n9915 & ~n9934;
  assign n9936 = n9925 & n9935;
  assign n9937 = ~pi38 & ~n9936;
  assign n9938 = ~n9922 & n9937;
  assign n9939 = ~pi32 & n9919;
  assign n9940 = pi32 & ~pi93;
  assign n9941 = n7382 & n9940;
  assign n9942 = n8793 & n9941;
  assign n9943 = ~n9939 & ~n9942;
  assign n9944 = ~pi95 & ~n6166;
  assign n9945 = ~n9943 & n9944;
  assign n9946 = n9938 & ~n9945;
  assign n9947 = n3351 & ~n9946;
  assign n9948 = ~n9913 & n9947;
  assign n9949 = ~n9912 & ~n9948;
  assign n9950 = n2535 & ~n9949;
  assign n9951 = pi137 & ~n8819;
  assign n9952 = ~po840 & n9951;
  assign n9953 = ~n8745 & ~n9952;
  assign n9954 = n8822 & ~n9953;
  assign n9955 = n8817 & n9954;
  assign n9956 = ~n9950 & ~n9955;
  assign n9957 = ~pi92 & ~n9956;
  assign n9958 = ~pi54 & ~n9957;
  assign n9959 = ~pi24 & n7294;
  assign n9960 = pi54 & ~n9959;
  assign n9961 = n2531 & ~n9960;
  assign n9962 = ~n9958 & n9961;
  assign n9963 = n6262 & n9962;
  assign n9964 = ~pi59 & ~n9963;
  assign n9965 = n2531 & n2576;
  assign n9966 = n8817 & n9965;
  assign n9967 = ~pi55 & n9966;
  assign n9968 = pi59 & ~n9967;
  assign n9969 = ~pi57 & ~n9968;
  assign po193 = ~n9964 & n9969;
  assign n9971 = n2712 & n7390;
  assign n9972 = pi36 & ~pi71;
  assign n9973 = n2463 & n2488;
  assign n9974 = n9050 & n9973;
  assign n9975 = ~pi65 & n9974;
  assign n9976 = ~pi69 & n9975;
  assign n9977 = ~pi67 & ~pi103;
  assign n9978 = n9976 & n9977;
  assign n9979 = ~pi83 & n2793;
  assign n9980 = n9978 & n9979;
  assign n9981 = n9972 & n9980;
  assign n9982 = n9971 & n9981;
  assign n9983 = ~pi58 & n7435;
  assign n9984 = ~n9982 & ~n9983;
  assign n9985 = n2533 & n6090;
  assign n9986 = n8738 & n9985;
  assign n9987 = n3084 & n9078;
  assign n9988 = n9986 & n9987;
  assign n9989 = po740 & n9988;
  assign po194 = ~n9984 & n9989;
  assign n9991 = n3084 & n9167;
  assign n9992 = n2502 & n9991;
  assign n9993 = n2918 & n9992;
  assign n9994 = ~pi45 & ~pi49;
  assign n9995 = n2470 & n9994;
  assign n9996 = pi89 & n9995;
  assign n9997 = ~pi48 & ~pi65;
  assign n9998 = n8775 & n9997;
  assign n9999 = n9996 & n9998;
  assign n10000 = ~pi71 & n2488;
  assign n10001 = ~pi104 & n10000;
  assign n10002 = n2477 & n9045;
  assign n10003 = n10001 & n10002;
  assign n10004 = n9999 & n10003;
  assign n10005 = n9047 & n10004;
  assign n10006 = pi332 & n10005;
  assign n10007 = ~pi64 & ~n10006;
  assign n10008 = n2466 & ~n10007;
  assign n10009 = ~pi81 & ~n2780;
  assign n10010 = ~pi841 & n10009;
  assign n10011 = ~pi39 & n10010;
  assign n10012 = n10008 & n10011;
  assign n10013 = n9993 & n10012;
  assign n10014 = ~pi38 & ~n10013;
  assign n10015 = pi24 & n2699;
  assign n10016 = ~pi32 & n8806;
  assign n10017 = n2686 & n10016;
  assign n10018 = n10015 & n10017;
  assign n10019 = pi38 & ~n10018;
  assign n10020 = n2571 & n7309;
  assign n10021 = ~po1038 & n10020;
  assign n10022 = ~n10019 & n10021;
  assign po196 = ~n10014 & n10022;
  assign n10024 = ~pi38 & n10021;
  assign n10025 = pi786 & ~pi1082;
  assign n10026 = ~pi984 & ~n6120;
  assign n10027 = pi835 & ~n10026;
  assign n10028 = n6177 & ~n10027;
  assign n10029 = n6212 & ~n10028;
  assign n10030 = pi1093 & n10029;
  assign n10031 = n6178 & n6440;
  assign n10032 = ~n10030 & n10031;
  assign n10033 = ~pi223 & n10032;
  assign n10034 = ~n6215 & n10029;
  assign n10035 = n10031 & ~n10034;
  assign n10036 = ~n6236 & n10035;
  assign n10037 = n6191 & n10029;
  assign n10038 = n10031 & ~n10037;
  assign n10039 = n6236 & n10038;
  assign n10040 = ~pi299 & ~n10039;
  assign n10041 = ~n10036 & n10040;
  assign n10042 = ~n10033 & n10041;
  assign n10043 = ~pi215 & n10032;
  assign n10044 = ~n6198 & n10035;
  assign n10045 = n6198 & n10038;
  assign n10046 = pi299 & ~n10045;
  assign n10047 = ~n10044 & n10046;
  assign n10048 = ~n10043 & n10047;
  assign n10049 = ~n10042 & ~n10048;
  assign n10050 = ~n10025 & n10049;
  assign n10051 = n5975 & ~n6200;
  assign n10052 = n5792 & ~n6238;
  assign n10053 = ~n10051 & ~n10052;
  assign n10054 = po740 & ~n10053;
  assign n10055 = n10025 & n10054;
  assign n10056 = n6442 & n10055;
  assign n10057 = ~n10050 & ~n10056;
  assign n10058 = pi39 & ~n10057;
  assign n10059 = n6166 & n6373;
  assign n10060 = pi35 & ~n6370;
  assign n10061 = n2918 & ~n10060;
  assign n10062 = ~pi986 & ~po740;
  assign n10063 = pi252 & ~n10062;
  assign n10064 = pi314 & ~n10063;
  assign n10065 = n6148 & n10064;
  assign n10066 = ~pi46 & n2691;
  assign n10067 = pi108 & n10066;
  assign n10068 = n2766 & n10067;
  assign n10069 = ~n2767 & n10066;
  assign n10070 = n8771 & n10003;
  assign n10071 = n2463 & n2795;
  assign n10072 = ~pi66 & ~pi84;
  assign n10073 = n8772 & n10072;
  assign n10074 = ~pi65 & ~pi69;
  assign n10075 = n10073 & n10074;
  assign n10076 = pi48 & n10075;
  assign n10077 = ~pi82 & n10076;
  assign n10078 = ~pi45 & n10077;
  assign n10079 = n10071 & n10078;
  assign n10080 = n8767 & n10079;
  assign n10081 = n10070 & n10080;
  assign n10082 = ~pi841 & n2493;
  assign n10083 = n2706 & n10082;
  assign n10084 = ~pi97 & n10083;
  assign n10085 = n10081 & n10084;
  assign n10086 = n10069 & n10085;
  assign n10087 = ~pi47 & ~n10086;
  assign n10088 = ~n10068 & n10087;
  assign n10089 = n10065 & ~n10088;
  assign n10090 = ~pi47 & ~pi841;
  assign n10091 = n10081 & n10090;
  assign n10092 = ~n2753 & ~n10091;
  assign n10093 = n2500 & ~n10092;
  assign n10094 = ~n10064 & n10093;
  assign n10095 = n2692 & n10094;
  assign n10096 = ~n10089 & ~n10095;
  assign n10097 = n2696 & ~n10096;
  assign n10098 = ~pi35 & ~n10097;
  assign n10099 = n2461 & ~n10098;
  assign n10100 = n10061 & n10099;
  assign n10101 = ~n10059 & ~n10100;
  assign n10102 = n8806 & ~n10101;
  assign n10103 = ~n10058 & ~n10102;
  assign po197 = n10024 & ~n10103;
  assign n10105 = pi102 & n2509;
  assign n10106 = n2941 & n10105;
  assign n10107 = n2491 & n2502;
  assign n10108 = n2465 & n10107;
  assign n10109 = n10106 & n10108;
  assign n10110 = n3084 & n10109;
  assign n10111 = pi1082 & ~n10110;
  assign n10112 = n2516 & ~n3375;
  assign n10113 = ~pi40 & ~n10109;
  assign n10114 = n10112 & ~n10113;
  assign n10115 = ~pi1082 & ~n10114;
  assign n10116 = n9986 & ~n10115;
  assign po198 = ~n10111 & n10116;
  assign n10118 = ~pi166 & n6190;
  assign n10119 = pi161 & n10118;
  assign n10120 = ~pi152 & n10119;
  assign n10121 = ~n6100 & ~n10120;
  assign n10122 = ~pi189 & n6190;
  assign n10123 = pi144 & n10122;
  assign n10124 = ~pi174 & n10123;
  assign n10125 = ~pi299 & ~n10124;
  assign n10126 = pi232 & ~n10125;
  assign n10127 = ~n10121 & n10126;
  assign n10128 = ~pi72 & ~n10127;
  assign n10129 = pi39 & ~n10128;
  assign n10130 = ~pi41 & ~pi72;
  assign n10131 = ~pi39 & ~n10130;
  assign n10132 = ~n10129 & ~n10131;
  assign n10133 = ~n7380 & ~n10132;
  assign n10134 = ~po1038 & ~n10133;
  assign n10135 = ~n7484 & ~n10130;
  assign n10136 = ~n2914 & n10130;
  assign n10137 = n7484 & ~n10136;
  assign n10138 = ~pi44 & n2522;
  assign n10139 = ~pi101 & n10138;
  assign n10140 = n7480 & n10139;
  assign n10141 = pi41 & ~n10140;
  assign n10142 = ~pi41 & pi72;
  assign n10143 = n2914 & ~n10142;
  assign n10144 = ~pi99 & n6115;
  assign n10145 = n2914 & ~n10144;
  assign n10146 = ~n10143 & ~n10145;
  assign n10147 = ~pi72 & pi101;
  assign n10148 = ~pi41 & ~n10147;
  assign n10149 = n2699 & n3084;
  assign n10150 = ~pi44 & n10149;
  assign n10151 = n10148 & n10150;
  assign n10152 = ~n10142 & ~n10151;
  assign n10153 = ~pi72 & ~n7480;
  assign n10154 = ~n10152 & ~n10153;
  assign n10155 = ~n10144 & n10154;
  assign n10156 = ~n10146 & ~n10155;
  assign n10157 = ~n10141 & n10156;
  assign n10158 = n10137 & ~n10157;
  assign n10159 = ~n10135 & ~n10158;
  assign n10160 = ~pi39 & ~n10159;
  assign n10161 = ~n10129 & ~n10160;
  assign n10162 = n6098 & ~n10161;
  assign n10163 = pi38 & ~n10132;
  assign n10164 = pi287 & n2522;
  assign n10165 = n10127 & n10164;
  assign n10166 = ~n10128 & ~n10165;
  assign n10167 = pi39 & ~n10166;
  assign n10168 = pi901 & ~pi959;
  assign n10169 = n2497 & n2771;
  assign n10170 = n2711 & n10169;
  assign n10171 = n2698 & n10170;
  assign n10172 = ~pi480 & pi949;
  assign n10173 = n2698 & n10172;
  assign n10174 = n2693 & n2751;
  assign n10175 = pi110 & n10174;
  assign n10176 = n10173 & n10175;
  assign n10177 = ~n10171 & ~n10176;
  assign n10178 = n10168 & n10177;
  assign n10179 = ~n10168 & ~n10176;
  assign n10180 = ~pi250 & pi252;
  assign n10181 = ~n10179 & n10180;
  assign n10182 = n3084 & n10181;
  assign n10183 = ~n10178 & n10182;
  assign n10184 = ~pi72 & n10183;
  assign n10185 = n9987 & n10175;
  assign n10186 = n10172 & ~n10180;
  assign n10187 = n10185 & n10186;
  assign n10188 = ~n10184 & ~n10187;
  assign n10189 = ~pi44 & ~n10188;
  assign n10190 = ~pi101 & n10189;
  assign n10191 = pi41 & ~n10190;
  assign n10192 = pi44 & ~pi72;
  assign n10193 = ~pi72 & ~n10183;
  assign n10194 = n3084 & ~n10180;
  assign n10195 = n10176 & n10194;
  assign n10196 = n10193 & ~n10195;
  assign n10197 = ~n10192 & ~n10196;
  assign n10198 = ~pi101 & ~n10197;
  assign n10199 = n10148 & ~n10198;
  assign n10200 = ~n10191 & ~n10199;
  assign n10201 = ~pi228 & ~n10200;
  assign n10202 = n7399 & ~n7404;
  assign n10203 = ~pi1093 & ~n7408;
  assign n10204 = ~n10202 & n10203;
  assign n10205 = ~pi1093 & ~n10204;
  assign n10206 = ~n7399 & ~n10205;
  assign n10207 = ~pi44 & ~n10206;
  assign n10208 = ~pi101 & n10207;
  assign n10209 = pi41 & ~n10208;
  assign n10210 = ~pi72 & n10206;
  assign n10211 = ~n10192 & ~n10210;
  assign n10212 = ~pi101 & ~n10211;
  assign n10213 = n10148 & ~n10212;
  assign n10214 = ~n2914 & ~n10213;
  assign n10215 = ~n10209 & n10214;
  assign n10216 = n2940 & ~n7392;
  assign n10217 = n2938 & n10216;
  assign n10218 = ~n7435 & ~n10217;
  assign n10219 = n2462 & ~n10218;
  assign n10220 = n7384 & ~n10219;
  assign n10221 = n7381 & ~n10220;
  assign n10222 = ~pi51 & ~n10221;
  assign n10223 = ~n2742 & ~n10222;
  assign n10224 = ~pi96 & ~n10223;
  assign n10225 = n7448 & ~n10224;
  assign n10226 = ~pi122 & n10225;
  assign n10227 = ~n10202 & ~n10226;
  assign n10228 = pi1093 & n10227;
  assign n10229 = ~n10204 & ~n10228;
  assign n10230 = ~pi44 & n10229;
  assign n10231 = ~pi101 & n10230;
  assign n10232 = pi41 & ~n10231;
  assign n10233 = ~pi72 & ~n10231;
  assign n10234 = ~pi41 & ~n10233;
  assign n10235 = n2914 & ~n10234;
  assign n10236 = ~n10232 & n10235;
  assign n10237 = ~n10215 & ~n10236;
  assign n10238 = pi228 & n10237;
  assign n10239 = ~pi39 & ~n10238;
  assign n10240 = ~n10201 & n10239;
  assign n10241 = ~n10167 & ~n10240;
  assign n10242 = n2614 & n10241;
  assign n10243 = ~pi87 & ~n10242;
  assign n10244 = ~n10163 & n10243;
  assign n10245 = ~n10162 & n10244;
  assign n10246 = ~pi75 & ~n10245;
  assign n10247 = ~pi228 & n10130;
  assign n10248 = pi41 & ~n10139;
  assign n10249 = pi228 & ~n10248;
  assign n10250 = n10152 & n10249;
  assign n10251 = ~n10247 & ~n10250;
  assign n10252 = n2533 & n10251;
  assign n10253 = pi87 & ~n10252;
  assign n10254 = ~n2614 & n10131;
  assign n10255 = ~n10129 & ~n10254;
  assign n10256 = n10253 & n10255;
  assign n10257 = n10246 & ~n10256;
  assign n10258 = ~n2572 & n10132;
  assign n10259 = pi75 & ~n10258;
  assign n10260 = n7423 & n10140;
  assign n10261 = pi41 & ~n10260;
  assign n10262 = pi252 & n3084;
  assign n10263 = ~pi24 & n2699;
  assign n10264 = n7480 & n10263;
  assign n10265 = n10262 & n10264;
  assign n10266 = ~pi44 & n10265;
  assign n10267 = n10148 & n10266;
  assign n10268 = ~n10144 & n10267;
  assign n10269 = ~n10261 & ~n10268;
  assign n10270 = n10143 & n10269;
  assign n10271 = n10137 & ~n10270;
  assign n10272 = ~n10135 & ~n10271;
  assign n10273 = ~pi39 & ~n10272;
  assign n10274 = ~n10129 & ~n10273;
  assign n10275 = n2572 & n10274;
  assign n10276 = n10259 & ~n10275;
  assign n10277 = ~n10257 & ~n10276;
  assign n10278 = n7380 & ~n10277;
  assign n10279 = n10134 & ~n10278;
  assign n10280 = pi39 & pi232;
  assign n10281 = n10120 & n10280;
  assign n10282 = ~n10131 & ~n10281;
  assign n10283 = ~pi72 & n10282;
  assign n10284 = po1038 & n10283;
  assign po199 = ~n10279 & ~n10284;
  assign n10286 = pi42 & ~pi72;
  assign n10287 = ~pi39 & ~n10286;
  assign n10288 = ~pi72 & pi199;
  assign n10289 = ~pi232 & ~n10288;
  assign n10290 = ~pi299 & ~n10289;
  assign n10291 = ~pi72 & ~n10122;
  assign n10292 = pi199 & n10291;
  assign n10293 = pi232 & ~n10292;
  assign n10294 = n10290 & ~n10293;
  assign n10295 = pi232 & n10118;
  assign n10296 = ~pi72 & ~n10295;
  assign n10297 = pi299 & n10296;
  assign n10298 = pi39 & ~n10297;
  assign n10299 = ~n10294 & n10298;
  assign n10300 = ~n10287 & ~n10299;
  assign n10301 = ~n7380 & n10300;
  assign n10302 = pi207 & pi208;
  assign n10303 = ~n2572 & n10286;
  assign n10304 = ~pi39 & ~n10303;
  assign n10305 = ~n7484 & ~n10286;
  assign n10306 = ~pi115 & n2914;
  assign n10307 = n10286 & ~n10306;
  assign n10308 = n7484 & ~n10307;
  assign n10309 = pi114 & ~n10286;
  assign n10310 = n10306 & ~n10309;
  assign n10311 = n6108 & n10139;
  assign n10312 = n6112 & n10311;
  assign n10313 = n7480 & n10312;
  assign n10314 = n7423 & n10313;
  assign n10315 = ~pi114 & ~n6111;
  assign n10316 = n10314 & n10315;
  assign n10317 = ~pi42 & n10316;
  assign n10318 = n6109 & n10266;
  assign n10319 = ~pi113 & n10318;
  assign n10320 = ~pi116 & n10319;
  assign n10321 = n10286 & ~n10320;
  assign n10322 = ~pi114 & ~n10321;
  assign n10323 = ~n10317 & n10322;
  assign n10324 = n10310 & ~n10323;
  assign n10325 = n10308 & ~n10324;
  assign n10326 = ~n10305 & ~n10325;
  assign n10327 = n2572 & n10326;
  assign n10328 = n10304 & ~n10327;
  assign n10329 = ~n10299 & ~n10328;
  assign n10330 = pi75 & ~n10329;
  assign n10331 = pi38 & ~n10300;
  assign n10332 = ~pi87 & ~n10331;
  assign n10333 = n10313 & n10315;
  assign n10334 = ~pi42 & n10333;
  assign n10335 = n6109 & n10150;
  assign n10336 = n6112 & n10335;
  assign n10337 = ~pi72 & ~n10336;
  assign n10338 = ~n10153 & ~n10337;
  assign n10339 = pi42 & ~n10338;
  assign n10340 = ~pi114 & ~n10339;
  assign n10341 = ~n10334 & n10340;
  assign n10342 = n10310 & ~n10341;
  assign n10343 = n10308 & ~n10342;
  assign n10344 = ~n10305 & ~n10343;
  assign n10345 = ~pi39 & ~n10344;
  assign n10346 = ~n10299 & ~n10345;
  assign n10347 = n6098 & ~n10346;
  assign n10348 = pi42 & ~pi114;
  assign n10349 = ~pi113 & n6108;
  assign n10350 = n10231 & n10349;
  assign n10351 = ~pi116 & n10350;
  assign n10352 = ~pi72 & ~n10351;
  assign n10353 = n10348 & ~n10352;
  assign n10354 = ~pi42 & ~n10351;
  assign n10355 = ~n10309 & ~n10354;
  assign n10356 = ~n10353 & n10355;
  assign n10357 = n10306 & ~n10356;
  assign n10358 = pi228 & ~n10357;
  assign n10359 = pi115 & ~n10286;
  assign n10360 = ~pi115 & ~n2914;
  assign n10361 = ~pi72 & pi116;
  assign n10362 = n6108 & n10208;
  assign n10363 = ~pi113 & n10362;
  assign n10364 = ~pi72 & ~n10363;
  assign n10365 = ~n10361 & ~n10364;
  assign n10366 = pi42 & ~n10365;
  assign n10367 = n6112 & n10362;
  assign n10368 = ~pi42 & n10367;
  assign n10369 = ~pi114 & ~n10368;
  assign n10370 = ~n10366 & n10369;
  assign n10371 = ~n10309 & ~n10370;
  assign n10372 = n10360 & ~n10371;
  assign n10373 = ~n10359 & ~n10372;
  assign n10374 = n10358 & n10373;
  assign n10375 = ~pi39 & ~n10374;
  assign n10376 = pi72 & ~n6108;
  assign n10377 = ~pi99 & n10199;
  assign n10378 = ~n10376 & ~n10377;
  assign n10379 = ~pi72 & pi113;
  assign n10380 = ~n10378 & ~n10379;
  assign n10381 = ~n10361 & n10380;
  assign n10382 = n10348 & n10381;
  assign n10383 = n10190 & n10349;
  assign n10384 = ~pi116 & n10383;
  assign n10385 = ~pi42 & ~n10384;
  assign n10386 = ~n10309 & ~n10385;
  assign n10387 = ~n10382 & n10386;
  assign n10388 = ~pi115 & ~n10387;
  assign n10389 = ~pi228 & ~n10388;
  assign n10390 = ~n10359 & n10389;
  assign n10391 = n10375 & ~n10390;
  assign n10392 = pi232 & pi299;
  assign n10393 = ~n10296 & n10392;
  assign n10394 = n10118 & n10164;
  assign n10395 = n10393 & ~n10394;
  assign n10396 = pi72 & ~pi232;
  assign n10397 = pi299 & ~n10396;
  assign n10398 = n10289 & ~n10397;
  assign n10399 = n6190 & n10164;
  assign n10400 = ~pi189 & n10399;
  assign n10401 = ~n10291 & ~n10400;
  assign n10402 = pi199 & ~n10401;
  assign n10403 = pi232 & ~n10402;
  assign n10404 = ~pi299 & n10403;
  assign n10405 = ~n10398 & ~n10404;
  assign n10406 = ~n10395 & n10405;
  assign n10407 = pi39 & ~n10406;
  assign n10408 = ~n10391 & ~n10407;
  assign n10409 = n2614 & ~n10408;
  assign n10410 = ~n10347 & ~n10409;
  assign n10411 = n10332 & n10410;
  assign n10412 = pi228 & n10336;
  assign n10413 = ~pi115 & n10412;
  assign n10414 = ~pi114 & n10413;
  assign n10415 = n10286 & ~n10414;
  assign n10416 = ~pi42 & n6113;
  assign n10417 = pi228 & n10312;
  assign n10418 = n10416 & n10417;
  assign n10419 = ~n10415 & ~n10418;
  assign n10420 = n2533 & n10419;
  assign n10421 = ~n2614 & n10287;
  assign n10422 = pi87 & ~n10421;
  assign n10423 = ~n10420 & n10422;
  assign n10424 = ~n10299 & n10423;
  assign n10425 = ~pi75 & ~n10424;
  assign n10426 = ~n10411 & n10425;
  assign n10427 = ~n10330 & ~n10426;
  assign n10428 = n7380 & n10427;
  assign n10429 = ~n10302 & ~n10428;
  assign n10430 = ~pi72 & pi200;
  assign n10431 = ~pi232 & ~n10430;
  assign n10432 = ~pi299 & ~n10431;
  assign n10433 = pi200 & n10291;
  assign n10434 = pi232 & ~n10433;
  assign n10435 = n10432 & ~n10434;
  assign n10436 = pi39 & ~n10435;
  assign n10437 = ~n10294 & n10436;
  assign n10438 = ~n10287 & ~n10437;
  assign n10439 = ~n7380 & n10438;
  assign n10440 = n10302 & ~n10439;
  assign n10441 = n10299 & n10436;
  assign n10442 = ~n10328 & ~n10441;
  assign n10443 = pi75 & ~n10442;
  assign n10444 = ~n10345 & ~n10441;
  assign n10445 = n6098 & ~n10444;
  assign n10446 = pi38 & ~n10438;
  assign n10447 = ~pi87 & ~n10446;
  assign n10448 = ~n10332 & ~n10447;
  assign n10449 = pi200 & ~n10401;
  assign n10450 = pi232 & ~n10449;
  assign n10451 = ~pi299 & n10450;
  assign n10452 = ~n10402 & n10451;
  assign n10453 = n10398 & ~n10430;
  assign n10454 = ~n10395 & ~n10453;
  assign n10455 = ~n10452 & n10454;
  assign n10456 = pi39 & ~n10455;
  assign n10457 = ~n10391 & ~n10456;
  assign n10458 = n2614 & ~n10457;
  assign n10459 = ~n10448 & ~n10458;
  assign n10460 = ~n10445 & n10459;
  assign n10461 = n10423 & ~n10441;
  assign n10462 = ~pi75 & ~n10461;
  assign n10463 = ~n10460 & n10462;
  assign n10464 = ~n10443 & ~n10463;
  assign n10465 = n7380 & n10464;
  assign n10466 = n10440 & ~n10465;
  assign n10467 = ~n10429 & ~n10466;
  assign n10468 = pi212 & pi214;
  assign n10469 = pi211 & n10468;
  assign n10470 = ~pi219 & ~n10469;
  assign n10471 = ~n10467 & ~n10470;
  assign n10472 = ~n10301 & n10471;
  assign n10473 = pi39 & ~n10294;
  assign n10474 = ~n10287 & ~n10473;
  assign n10475 = ~n7380 & n10474;
  assign n10476 = n10423 & ~n10473;
  assign n10477 = ~n10345 & ~n10473;
  assign n10478 = n6098 & ~n10477;
  assign n10479 = pi38 & ~n10474;
  assign n10480 = n10290 & ~n10403;
  assign n10481 = pi39 & ~n10480;
  assign n10482 = ~n10391 & ~n10481;
  assign n10483 = n2614 & ~n10482;
  assign n10484 = ~pi87 & ~n10483;
  assign n10485 = ~n10479 & n10484;
  assign n10486 = ~n10478 & n10485;
  assign n10487 = ~pi75 & ~n10486;
  assign n10488 = ~n10476 & n10487;
  assign n10489 = ~n10328 & ~n10473;
  assign n10490 = pi75 & ~n10489;
  assign n10491 = n7380 & ~n10490;
  assign n10492 = ~n10488 & n10491;
  assign n10493 = ~n10475 & ~n10492;
  assign n10494 = ~n10302 & n10493;
  assign n10495 = ~n10328 & ~n10437;
  assign n10496 = pi75 & ~n10495;
  assign n10497 = ~n10345 & ~n10437;
  assign n10498 = n6098 & ~n10497;
  assign n10499 = ~n10290 & ~n10432;
  assign n10500 = ~n10402 & n10450;
  assign n10501 = ~n10499 & ~n10500;
  assign n10502 = pi39 & ~n10501;
  assign n10503 = ~n10391 & ~n10502;
  assign n10504 = n2614 & ~n10503;
  assign n10505 = ~n10498 & ~n10504;
  assign n10506 = n10447 & n10505;
  assign n10507 = n10423 & ~n10437;
  assign n10508 = ~pi75 & ~n10507;
  assign n10509 = ~n10506 & n10508;
  assign n10510 = ~n10496 & ~n10509;
  assign n10511 = n7380 & n10510;
  assign n10512 = n10440 & ~n10511;
  assign n10513 = ~n10494 & ~n10512;
  assign n10514 = n10470 & ~n10513;
  assign n10515 = ~po1038 & ~n10514;
  assign n10516 = ~n10472 & n10515;
  assign n10517 = n10296 & ~n10470;
  assign n10518 = pi39 & ~n10517;
  assign n10519 = po1038 & ~n10287;
  assign n10520 = ~n10518 & n10519;
  assign po200 = n10516 | n10520;
  assign n10522 = ~pi211 & pi219;
  assign n10523 = ~pi211 & ~n10468;
  assign n10524 = ~n10469 & ~n10523;
  assign n10525 = ~n10522 & n10524;
  assign n10526 = pi43 & ~pi72;
  assign n10527 = ~pi39 & ~n10526;
  assign n10528 = ~n10436 & ~n10527;
  assign n10529 = ~n7380 & n10528;
  assign n10530 = pi228 & n10416;
  assign n10531 = n10526 & ~n10530;
  assign n10532 = ~pi43 & ~n10312;
  assign n10533 = pi43 & ~n10337;
  assign n10534 = ~n10532 & ~n10533;
  assign n10535 = n10530 & n10534;
  assign n10536 = ~n10531 & ~n10535;
  assign n10537 = n2533 & n10536;
  assign n10538 = ~n2614 & n10527;
  assign n10539 = pi87 & ~n10538;
  assign n10540 = ~n10537 & n10539;
  assign n10541 = ~n10436 & n10540;
  assign n10542 = ~n7484 & ~n10526;
  assign n10543 = n2914 & n10416;
  assign n10544 = n10526 & ~n10543;
  assign n10545 = n7484 & ~n10544;
  assign n10546 = ~pi43 & pi52;
  assign n10547 = n10313 & n10546;
  assign n10548 = pi43 & ~n10338;
  assign n10549 = ~n10547 & ~n10548;
  assign n10550 = n10543 & ~n10549;
  assign n10551 = n10545 & ~n10550;
  assign n10552 = ~n10542 & ~n10551;
  assign n10553 = ~pi39 & ~n10552;
  assign n10554 = ~n10436 & ~n10553;
  assign n10555 = n6098 & ~n10554;
  assign n10556 = pi38 & ~n10528;
  assign n10557 = n6108 & n10190;
  assign n10558 = ~pi228 & ~n10557;
  assign n10559 = ~n2914 & ~n10362;
  assign n10560 = n6108 & n10231;
  assign n10561 = n2914 & ~n10560;
  assign n10562 = ~n10559 & ~n10561;
  assign n10563 = pi228 & ~n10562;
  assign n10564 = n6112 & ~n10563;
  assign n10565 = ~n10558 & n10564;
  assign n10566 = ~pi43 & ~n10565;
  assign n10567 = n10416 & ~n10566;
  assign n10568 = ~n10526 & ~n10567;
  assign n10569 = ~n2914 & n10367;
  assign n10570 = pi116 & n10364;
  assign n10571 = ~n2914 & ~n10570;
  assign n10572 = pi116 & ~n2914;
  assign n10573 = ~n10351 & ~n10572;
  assign n10574 = ~n10350 & n10361;
  assign n10575 = n10573 & ~n10574;
  assign n10576 = ~n10571 & ~n10575;
  assign n10577 = ~n10569 & ~n10576;
  assign n10578 = ~pi116 & ~n10577;
  assign n10579 = ~pi72 & ~n10578;
  assign n10580 = pi228 & ~n10579;
  assign n10581 = ~pi228 & n10381;
  assign n10582 = ~n10580 & ~n10581;
  assign n10583 = n10416 & ~n10582;
  assign n10584 = pi43 & n10583;
  assign n10585 = ~n10568 & ~n10584;
  assign n10586 = ~pi39 & ~n10585;
  assign n10587 = n10432 & ~n10450;
  assign n10588 = pi39 & ~n10587;
  assign n10589 = ~n10586 & ~n10588;
  assign n10590 = n2614 & ~n10589;
  assign n10591 = ~pi87 & ~n10590;
  assign n10592 = ~n10556 & n10591;
  assign n10593 = ~n10555 & n10592;
  assign n10594 = ~pi75 & ~n10593;
  assign n10595 = ~n10541 & n10594;
  assign n10596 = ~n2572 & n10526;
  assign n10597 = ~pi39 & ~n10596;
  assign n10598 = ~pi72 & ~n10320;
  assign n10599 = pi43 & n10598;
  assign n10600 = n10314 & n10546;
  assign n10601 = ~n10599 & ~n10600;
  assign n10602 = n10543 & ~n10601;
  assign n10603 = n10545 & ~n10602;
  assign n10604 = ~n10542 & ~n10603;
  assign n10605 = n2572 & n10604;
  assign n10606 = n10597 & ~n10605;
  assign n10607 = ~n10436 & ~n10606;
  assign n10608 = pi75 & ~n10607;
  assign n10609 = n7380 & ~n10608;
  assign n10610 = ~n10595 & n10609;
  assign n10611 = ~n10529 & ~n10610;
  assign n10612 = ~n10302 & ~n10611;
  assign n10613 = ~n10525 & ~n10612;
  assign n10614 = ~pi199 & ~pi200;
  assign n10615 = ~pi299 & ~n10614;
  assign n10616 = ~pi72 & ~n10615;
  assign n10617 = ~pi232 & ~n10616;
  assign n10618 = ~pi299 & ~n10617;
  assign n10619 = n10291 & n10614;
  assign n10620 = pi232 & ~n10619;
  assign n10621 = n10618 & ~n10620;
  assign n10622 = pi39 & ~n10621;
  assign n10623 = ~n10527 & ~n10622;
  assign n10624 = ~n7380 & n10623;
  assign n10625 = ~n2533 & ~n10623;
  assign n10626 = n10540 & ~n10625;
  assign n10627 = ~n10553 & ~n10622;
  assign n10628 = n6098 & ~n10627;
  assign n10629 = pi38 & ~n10623;
  assign n10630 = ~n10401 & n10614;
  assign n10631 = pi232 & ~n10630;
  assign n10632 = n10618 & ~n10631;
  assign n10633 = pi39 & ~n10632;
  assign n10634 = ~n10586 & ~n10633;
  assign n10635 = n2614 & ~n10634;
  assign n10636 = ~pi87 & ~n10635;
  assign n10637 = ~n10629 & n10636;
  assign n10638 = ~n10628 & n10637;
  assign n10639 = ~pi75 & ~n10638;
  assign n10640 = ~n10626 & n10639;
  assign n10641 = ~n10606 & ~n10622;
  assign n10642 = pi75 & ~n10641;
  assign n10643 = n7380 & ~n10642;
  assign n10644 = ~n10640 & n10643;
  assign n10645 = ~n10624 & ~n10644;
  assign n10646 = n10302 & ~n10645;
  assign n10647 = n10613 & ~n10646;
  assign n10648 = n10298 & ~n10435;
  assign n10649 = ~n10527 & ~n10648;
  assign n10650 = ~n7380 & n10649;
  assign n10651 = n10540 & ~n10648;
  assign n10652 = ~n10553 & ~n10648;
  assign n10653 = n6098 & ~n10652;
  assign n10654 = pi38 & ~n10649;
  assign n10655 = ~n10397 & n10431;
  assign n10656 = ~n10451 & ~n10655;
  assign n10657 = ~n10395 & n10656;
  assign n10658 = pi39 & ~n10657;
  assign n10659 = ~n10586 & ~n10658;
  assign n10660 = n2614 & ~n10659;
  assign n10661 = ~pi87 & ~n10660;
  assign n10662 = ~n10654 & n10661;
  assign n10663 = ~n10653 & n10662;
  assign n10664 = ~pi75 & ~n10663;
  assign n10665 = ~n10651 & n10664;
  assign n10666 = ~n10606 & ~n10648;
  assign n10667 = pi75 & ~n10666;
  assign n10668 = n7380 & ~n10667;
  assign n10669 = ~n10665 & n10668;
  assign n10670 = ~n10650 & ~n10669;
  assign n10671 = ~n10302 & ~n10670;
  assign n10672 = n10525 & ~n10671;
  assign n10673 = ~n10297 & n10622;
  assign n10674 = ~n10527 & ~n10673;
  assign n10675 = ~n7380 & n10674;
  assign n10676 = n10540 & ~n10673;
  assign n10677 = ~n10553 & ~n10673;
  assign n10678 = n6098 & ~n10677;
  assign n10679 = pi38 & ~n10674;
  assign n10680 = pi232 & ~pi299;
  assign n10681 = ~n10630 & n10680;
  assign n10682 = ~n10617 & ~n10681;
  assign n10683 = ~n10395 & n10682;
  assign n10684 = pi39 & ~n10683;
  assign n10685 = ~n10586 & ~n10684;
  assign n10686 = n2614 & ~n10685;
  assign n10687 = ~pi87 & ~n10686;
  assign n10688 = ~n10679 & n10687;
  assign n10689 = ~n10678 & n10688;
  assign n10690 = ~pi75 & ~n10689;
  assign n10691 = ~n10676 & n10690;
  assign n10692 = ~n10606 & ~n10673;
  assign n10693 = pi75 & ~n10692;
  assign n10694 = n7380 & ~n10693;
  assign n10695 = ~n10691 & n10694;
  assign n10696 = ~n10675 & ~n10695;
  assign n10697 = n10302 & ~n10696;
  assign n10698 = n10672 & ~n10697;
  assign n10699 = ~po1038 & ~n10698;
  assign n10700 = ~n10647 & n10699;
  assign n10701 = n10296 & n10525;
  assign n10702 = pi39 & ~n10701;
  assign n10703 = po1038 & ~n10527;
  assign n10704 = ~n10702 & n10703;
  assign po201 = n10700 | n10704;
  assign n10706 = ~pi39 & ~n10192;
  assign n10707 = pi39 & n7421;
  assign n10708 = ~pi72 & n10707;
  assign n10709 = pi39 & ~n10708;
  assign n10710 = ~n10706 & ~n10709;
  assign n10711 = ~n7380 & ~n10710;
  assign n10712 = ~po1038 & ~n10711;
  assign n10713 = ~n7484 & ~n10192;
  assign n10714 = ~pi39 & ~n10713;
  assign n10715 = ~n2914 & n10192;
  assign n10716 = n7484 & ~n10715;
  assign n10717 = pi44 & pi72;
  assign n10718 = n7425 & ~n10717;
  assign n10719 = n7480 & n10138;
  assign n10720 = n7423 & n10719;
  assign n10721 = pi44 & ~n10265;
  assign n10722 = ~n10720 & ~n10721;
  assign n10723 = n10718 & ~n10722;
  assign n10724 = n10716 & ~n10723;
  assign n10725 = n10714 & ~n10724;
  assign n10726 = ~n10708 & ~n10725;
  assign n10727 = n2572 & ~n10726;
  assign n10728 = ~n2572 & n10710;
  assign n10729 = pi75 & ~n10728;
  assign n10730 = ~n10727 & n10729;
  assign n10731 = pi287 & n10149;
  assign n10732 = n10708 & ~n10731;
  assign n10733 = n10192 & ~n10229;
  assign n10734 = n2914 & ~n10230;
  assign n10735 = ~n10733 & n10734;
  assign n10736 = pi44 & n10210;
  assign n10737 = ~n2914 & ~n10207;
  assign n10738 = ~n10736 & n10737;
  assign n10739 = ~n10735 & ~n10738;
  assign n10740 = pi228 & ~n10739;
  assign n10741 = pi44 & n10196;
  assign n10742 = ~pi228 & ~n10741;
  assign n10743 = ~n10189 & n10742;
  assign n10744 = ~pi39 & ~n10743;
  assign n10745 = ~n10740 & n10744;
  assign n10746 = ~n10732 & ~n10745;
  assign n10747 = n2614 & n10746;
  assign n10748 = pi38 & ~n10710;
  assign n10749 = ~pi87 & ~n10748;
  assign n10750 = n7480 & n10149;
  assign n10751 = pi44 & ~n10750;
  assign n10752 = ~n10719 & ~n10751;
  assign n10753 = n10718 & ~n10752;
  assign n10754 = n10716 & ~n10753;
  assign n10755 = n10714 & ~n10754;
  assign n10756 = ~n10708 & ~n10755;
  assign n10757 = n6098 & n10756;
  assign n10758 = n10749 & ~n10757;
  assign n10759 = ~n10747 & n10758;
  assign n10760 = ~pi75 & ~n10759;
  assign n10761 = pi228 & n2614;
  assign n10762 = n10138 & n10761;
  assign n10763 = n10149 & n10761;
  assign n10764 = n10192 & ~n10763;
  assign n10765 = ~pi39 & ~n10764;
  assign n10766 = ~n10762 & n10765;
  assign n10767 = ~n10709 & ~n10766;
  assign n10768 = pi87 & n10767;
  assign n10769 = n10760 & ~n10768;
  assign n10770 = ~n10730 & ~n10769;
  assign n10771 = n7380 & ~n10770;
  assign n10772 = n10712 & ~n10771;
  assign n10773 = n2627 & n7420;
  assign n10774 = ~pi72 & n10773;
  assign n10775 = pi39 & ~n10774;
  assign n10776 = po1038 & ~n10706;
  assign n10777 = ~n10775 & n10776;
  assign po202 = n10772 | n10777;
  assign n10779 = ~pi38 & pi39;
  assign n10780 = n10021 & n10779;
  assign n10781 = pi979 & n10780;
  assign po203 = n6440 & n10781;
  assign n10783 = ~pi76 & n8767;
  assign n10784 = ~pi102 & ~pi104;
  assign n10785 = ~pi111 & n10784;
  assign n10786 = pi61 & ~pi89;
  assign n10787 = n10785 & n10786;
  assign n10788 = n10783 & n10787;
  assign n10789 = ~pi83 & n2464;
  assign n10790 = ~pi82 & n10789;
  assign n10791 = n8759 & n8761;
  assign n10792 = n10790 & n10791;
  assign n10793 = n10075 & n10792;
  assign n10794 = n10000 & n10793;
  assign n10795 = n8781 & n10794;
  assign n10796 = n10788 & n10795;
  assign n10797 = ~pi841 & n10796;
  assign n10798 = n2694 & n2880;
  assign n10799 = pi24 & n10798;
  assign n10800 = ~n10797 & ~n10799;
  assign po204 = n9988 & ~n10800;
  assign n10802 = n2464 & ~n2863;
  assign n10803 = n2488 & n9977;
  assign n10804 = ~pi82 & n2479;
  assign n10805 = ~pi84 & n9995;
  assign n10806 = pi104 & n10805;
  assign n10807 = n2796 & n10806;
  assign n10808 = n10804 & n10807;
  assign n10809 = ~pi36 & ~n10808;
  assign n10810 = n8760 & n9050;
  assign n10811 = ~n10809 & n10810;
  assign n10812 = ~pi98 & n10811;
  assign n10813 = n10803 & n10812;
  assign n10814 = ~n2794 & n10813;
  assign n10815 = ~pi88 & ~n10814;
  assign n10816 = n2725 & ~n10815;
  assign n10817 = n10802 & n10816;
  assign n10818 = n2692 & n10817;
  assign n10819 = ~n9983 & ~n10818;
  assign n10820 = n9987 & ~n10819;
  assign n10821 = n7493 & ~n10820;
  assign n10822 = ~n6120 & n10820;
  assign n10823 = ~pi36 & n10813;
  assign n10824 = ~pi88 & ~n10823;
  assign n10825 = n10802 & ~n10824;
  assign n10826 = n9993 & n10825;
  assign n10827 = ~pi824 & n6120;
  assign n10828 = n10826 & n10827;
  assign n10829 = pi829 & ~n10828;
  assign n10830 = ~n10822 & n10829;
  assign n10831 = ~n2913 & n10830;
  assign n10832 = ~n10821 & ~n10831;
  assign n10833 = pi1091 & ~n10832;
  assign n10834 = ~n7368 & n10820;
  assign n10835 = ~pi829 & ~n10834;
  assign n10836 = ~n10830 & ~n10835;
  assign n10837 = ~pi1093 & ~n10836;
  assign n10838 = ~n6446 & ~n7490;
  assign n10839 = n7368 & n9987;
  assign n10840 = ~n9984 & n10839;
  assign n10841 = ~n10834 & ~n10840;
  assign n10842 = ~n10838 & n10841;
  assign n10843 = ~n10837 & ~n10842;
  assign n10844 = n9986 & n10843;
  assign po205 = ~n10833 & n10844;
  assign n10846 = pi841 & n9986;
  assign n10847 = n10081 & n10846;
  assign po206 = n9993 & n10847;
  assign n10849 = ~pi45 & n10804;
  assign n10850 = pi49 & n10849;
  assign n10851 = n8757 & n10073;
  assign n10852 = n8760 & n8766;
  assign n10853 = n10851 & n10852;
  assign n10854 = n2465 & n2488;
  assign n10855 = n10853 & n10854;
  assign n10856 = n10785 & n10855;
  assign n10857 = n10850 & n10856;
  assign n10858 = ~pi35 & ~pi51;
  assign n10859 = n8781 & n10858;
  assign n10860 = n10857 & n10859;
  assign n10861 = pi841 & n2696;
  assign n10862 = n2518 & n10861;
  assign n10863 = n10860 & n10862;
  assign n10864 = ~pi74 & ~n10863;
  assign n10865 = ~po1038 & ~n10864;
  assign n10866 = pi74 & ~n8817;
  assign n10867 = n10865 & ~n10866;
  assign po207 = n9985 & n10867;
  assign n10869 = ~pi94 & ~n8794;
  assign n10870 = pi24 & n10869;
  assign n10871 = pi24 & n8784;
  assign n10872 = ~n10170 & ~n10871;
  assign n10873 = pi252 & po840;
  assign n10874 = ~pi252 & n8744;
  assign n10875 = ~n10873 & ~n10874;
  assign n10876 = ~n10872 & ~n10875;
  assign n10877 = n9987 & n10876;
  assign n10878 = ~n10870 & n10877;
  assign n10879 = n2508 & n2517;
  assign n10880 = pi24 & ~pi90;
  assign n10881 = n10875 & n10880;
  assign n10882 = n8796 & n10881;
  assign n10883 = n10879 & n10882;
  assign n10884 = ~n10878 & ~n10883;
  assign n10885 = ~pi100 & ~n10884;
  assign n10886 = pi100 & n8819;
  assign n10887 = n6490 & n10886;
  assign n10888 = ~n10885 & ~n10887;
  assign n10889 = n2532 & ~n10888;
  assign n10890 = n2535 & n10889;
  assign n10891 = n8818 & n8819;
  assign n10892 = n8822 & n10891;
  assign n10893 = ~n10890 & ~n10892;
  assign po208 = n8739 & ~n10893;
  assign n10895 = n9051 & n10854;
  assign n10896 = n2468 & n10895;
  assign n10897 = ~pi69 & n10896;
  assign n10898 = n2795 & n10897;
  assign n10899 = n2692 & n9988;
  assign n10900 = n2725 & n10899;
  assign n10901 = n2798 & n10900;
  assign po209 = n10898 & n10901;
  assign n10903 = pi52 & ~pi72;
  assign n10904 = ~pi39 & n10903;
  assign n10905 = ~pi114 & n6110;
  assign n10906 = n7484 & n10306;
  assign n10907 = n10905 & n10906;
  assign n10908 = n2572 & n10907;
  assign n10909 = n10320 & n10908;
  assign n10910 = n10904 & ~n10909;
  assign n10911 = pi75 & n10910;
  assign n10912 = ~pi100 & n10779;
  assign n10913 = pi87 & ~n10912;
  assign n10914 = ~n2614 & ~n10904;
  assign n10915 = n10913 & ~n10914;
  assign n10916 = ~pi43 & n10530;
  assign n10917 = ~pi52 & n10312;
  assign n10918 = pi52 & n10337;
  assign n10919 = ~n10917 & ~n10918;
  assign n10920 = n10916 & ~n10919;
  assign n10921 = n10903 & ~n10916;
  assign n10922 = ~n10920 & ~n10921;
  assign n10923 = n2614 & n10922;
  assign n10924 = n10915 & ~n10923;
  assign n10925 = pi38 & ~n10904;
  assign n10926 = n6110 & n6113;
  assign n10927 = ~n10903 & ~n10926;
  assign n10928 = pi52 & n10352;
  assign n10929 = ~pi52 & n10351;
  assign n10930 = n10306 & ~n10929;
  assign n10931 = ~n10928 & n10930;
  assign n10932 = pi52 & ~n10365;
  assign n10933 = ~pi52 & n10367;
  assign n10934 = n10360 & ~n10933;
  assign n10935 = ~n10932 & n10934;
  assign n10936 = ~n10931 & ~n10935;
  assign n10937 = n10905 & ~n10936;
  assign n10938 = ~n10927 & ~n10937;
  assign n10939 = pi228 & n10938;
  assign n10940 = pi52 & ~n10381;
  assign n10941 = ~pi52 & n10384;
  assign n10942 = ~n10940 & ~n10941;
  assign n10943 = n10926 & n10942;
  assign n10944 = ~pi228 & ~n10927;
  assign n10945 = ~n10943 & n10944;
  assign n10946 = ~pi39 & ~n10945;
  assign n10947 = ~n10939 & n10946;
  assign n10948 = ~pi100 & n10947;
  assign n10949 = n10336 & n10907;
  assign n10950 = n7480 & n10949;
  assign n10951 = n10903 & ~n10950;
  assign n10952 = pi100 & ~n10951;
  assign n10953 = ~pi39 & ~n10952;
  assign n10954 = ~n10948 & n10953;
  assign n10955 = ~pi38 & ~n10954;
  assign n10956 = ~pi87 & ~n10955;
  assign n10957 = ~n10925 & n10956;
  assign n10958 = ~n10924 & ~n10957;
  assign n10959 = ~pi75 & ~n10958;
  assign n10960 = ~n10911 & ~n10959;
  assign n10961 = n7380 & n10960;
  assign n10962 = ~n7380 & ~n10904;
  assign n10963 = n10302 & ~n10962;
  assign n10964 = ~n10961 & n10963;
  assign n10965 = ~pi39 & ~n10903;
  assign n10966 = ~n10622 & ~n10965;
  assign n10967 = ~pi39 & ~n10910;
  assign n10968 = n10966 & ~n10967;
  assign n10969 = pi75 & ~n10968;
  assign n10970 = n7380 & ~n10969;
  assign n10971 = ~pi39 & ~n10951;
  assign n10972 = ~n10622 & ~n10971;
  assign n10973 = n6098 & ~n10972;
  assign n10974 = ~pi87 & ~n10973;
  assign n10975 = pi38 & ~n10966;
  assign n10976 = ~n10633 & ~n10947;
  assign n10977 = n2614 & ~n10976;
  assign n10978 = ~n10975 & ~n10977;
  assign n10979 = n10974 & n10978;
  assign n10980 = ~n2614 & n10966;
  assign n10981 = ~pi39 & n10922;
  assign n10982 = ~n10622 & ~n10981;
  assign n10983 = n2614 & n10982;
  assign n10984 = ~n10980 & ~n10983;
  assign n10985 = pi87 & ~n10984;
  assign n10986 = ~pi75 & ~n10985;
  assign n10987 = ~n10979 & n10986;
  assign n10988 = n10970 & ~n10987;
  assign n10989 = ~n10302 & n10988;
  assign n10990 = ~n10964 & ~n10989;
  assign n10991 = ~pi219 & n10523;
  assign n10992 = ~n10990 & ~n10991;
  assign n10993 = ~n10298 & ~n10965;
  assign n10994 = ~n7380 & ~n10993;
  assign n10995 = ~n10298 & ~n10971;
  assign n10996 = n6098 & ~n10995;
  assign n10997 = pi38 & ~n10993;
  assign n10998 = ~n10395 & n10397;
  assign n10999 = pi39 & ~n10998;
  assign n11000 = ~n10947 & ~n10999;
  assign n11001 = n2614 & ~n11000;
  assign n11002 = ~n10997 & ~n11001;
  assign n11003 = ~n10996 & n11002;
  assign n11004 = ~pi87 & ~n11003;
  assign n11005 = ~n2614 & n10993;
  assign n11006 = pi87 & ~n11005;
  assign n11007 = ~n10298 & ~n10981;
  assign n11008 = n2614 & n11007;
  assign n11009 = n11006 & ~n11008;
  assign n11010 = n10302 & ~n11009;
  assign n11011 = ~n11004 & n11010;
  assign n11012 = ~n10684 & ~n10947;
  assign n11013 = n2614 & ~n11012;
  assign n11014 = ~n10673 & ~n10971;
  assign n11015 = n6098 & ~n11014;
  assign n11016 = ~n11013 & ~n11015;
  assign n11017 = n10975 & ~n10993;
  assign n11018 = n11016 & ~n11017;
  assign n11019 = ~pi87 & ~n11018;
  assign n11020 = ~n10302 & ~n11019;
  assign n11021 = ~n10673 & ~n10981;
  assign n11022 = n2614 & n11021;
  assign n11023 = ~n10980 & ~n11022;
  assign n11024 = n11006 & n11023;
  assign n11025 = n11020 & ~n11024;
  assign n11026 = ~n11011 & ~n11025;
  assign n11027 = ~pi75 & ~n11026;
  assign n11028 = ~n10302 & n10621;
  assign n11029 = n10298 & ~n11028;
  assign n11030 = ~n10967 & ~n11029;
  assign n11031 = pi75 & n11030;
  assign n11032 = ~n11027 & ~n11031;
  assign n11033 = n7380 & n11032;
  assign n11034 = ~n10994 & ~n11033;
  assign n11035 = n10991 & n11034;
  assign n11036 = ~n7380 & n10966;
  assign n11037 = ~n10302 & n11036;
  assign n11038 = ~po1038 & ~n11037;
  assign n11039 = ~n11035 & n11038;
  assign n11040 = ~n10992 & n11039;
  assign n11041 = pi39 & n10991;
  assign n11042 = n10296 & n11041;
  assign n11043 = ~n10904 & ~n11042;
  assign n11044 = po1038 & n11043;
  assign po210 = ~n11040 & ~n11044;
  assign n11046 = pi24 & n9987;
  assign n11047 = pi53 & n2712;
  assign n11048 = n2706 & n11047;
  assign n11049 = n2707 & n11048;
  assign n11050 = n11046 & n11049;
  assign n11051 = ~pi39 & ~n11050;
  assign n11052 = ~pi287 & ~pi979;
  assign n11053 = n6175 & n11052;
  assign n11054 = pi39 & ~n11053;
  assign n11055 = n10024 & ~n11054;
  assign n11056 = ~n3366 & n11055;
  assign po211 = ~n11051 & n11056;
  assign n11058 = n2574 & n10018;
  assign n11059 = pi54 & ~n11058;
  assign n11060 = n8784 & n8874;
  assign n11061 = n8764 & n10851;
  assign n11062 = n8770 & n11061;
  assign n11063 = n10783 & n11062;
  assign n11064 = ~pi85 & pi106;
  assign n11065 = ~pi60 & n11064;
  assign n11066 = n2472 & n11065;
  assign n11067 = n10854 & n11066;
  assign n11068 = n11063 & n11067;
  assign n11069 = n11060 & n11068;
  assign n11070 = ~pi841 & n2696;
  assign n11071 = n2518 & n11070;
  assign n11072 = n3275 & n11071;
  assign n11073 = n10858 & n11072;
  assign n11074 = n11069 & n11073;
  assign n11075 = ~pi54 & ~n11074;
  assign n11076 = n8738 & ~n11075;
  assign po212 = ~n11059 & n11076;
  assign n11078 = n2575 & n10018;
  assign n11079 = pi55 & ~n11078;
  assign n11080 = pi45 & n10853;
  assign n11081 = n2472 & n2488;
  assign n11082 = n2481 & n11081;
  assign n11083 = n11080 & n11082;
  assign n11084 = n3084 & n9157;
  assign n11085 = n2466 & n2576;
  assign n11086 = n11084 & n11085;
  assign n11087 = n11083 & n11086;
  assign n11088 = ~pi55 & ~n11087;
  assign n11089 = n2531 & ~n11088;
  assign n11090 = n3327 & n11089;
  assign po213 = ~n11079 & n11090;
  assign n11092 = pi56 & ~pi62;
  assign n11093 = pi55 & n9966;
  assign n11094 = ~n11092 & ~n11093;
  assign n11095 = n2516 & n2539;
  assign n11096 = n2921 & n11095;
  assign n11097 = pi56 & ~n11096;
  assign n11098 = n3327 & ~n11097;
  assign po214 = ~n11094 & n11098;
  assign n11100 = n6372 & n11095;
  assign n11101 = ~pi56 & pi62;
  assign n11102 = ~pi924 & n11101;
  assign n11103 = ~n11092 & ~n11102;
  assign n11104 = n11100 & ~n11103;
  assign n11105 = ~pi57 & ~n11104;
  assign n11106 = n6273 & n11078;
  assign n11107 = pi57 & ~n11106;
  assign n11108 = ~pi59 & ~n11107;
  assign po215 = ~n11105 & n11108;
  assign n11110 = n9986 & n10879;
  assign n11111 = ~pi93 & n7383;
  assign po216 = n11110 & n11111;
  assign n11113 = pi924 & n11101;
  assign n11114 = n11100 & n11113;
  assign n11115 = ~pi59 & ~n11114;
  assign n11116 = pi59 & ~n11106;
  assign n11117 = ~pi57 & ~n11116;
  assign po217 = ~n11115 & n11117;
  assign n11119 = pi39 & ~n6175;
  assign n11120 = n6176 & n6440;
  assign n11121 = ~pi979 & n11120;
  assign n11122 = n11119 & n11121;
  assign n11123 = ~pi39 & n11060;
  assign n11124 = n2704 & n11123;
  assign n11125 = n11046 & n11124;
  assign n11126 = ~n11122 & ~n11125;
  assign po218 = n10024 & ~n11126;
  assign n11128 = pi841 & n10796;
  assign n11129 = ~pi24 & n11060;
  assign n11130 = n2704 & n11129;
  assign n11131 = ~n11128 & ~n11130;
  assign po219 = n9988 & ~n11131;
  assign n11133 = n11096 & n11101;
  assign n11134 = ~pi57 & ~n11133;
  assign n11135 = pi57 & ~n9967;
  assign n11136 = ~pi59 & ~n11135;
  assign po220 = ~n11134 & n11136;
  assign n11138 = n8781 & n8869;
  assign n11139 = n2854 & n11138;
  assign n11140 = pi999 & n11139;
  assign n11141 = ~pi24 & n10798;
  assign n11142 = ~n11140 & ~n11141;
  assign po221 = n9988 & ~n11142;
  assign n11144 = ~pi64 & ~n2842;
  assign n11145 = n2466 & ~n11144;
  assign n11146 = n10009 & n11145;
  assign n11147 = pi841 & ~n11146;
  assign n11148 = n2841 & n8870;
  assign n11149 = ~pi841 & ~n11148;
  assign n11150 = n10900 & ~n11149;
  assign po222 = ~n11147 & n11150;
  assign n11152 = pi39 & n10025;
  assign n11153 = n10024 & ~n10041;
  assign n11154 = ~n10047 & n11153;
  assign po223 = n11152 & n11154;
  assign n11156 = ~pi199 & ~pi299;
  assign n11157 = pi81 & n2490;
  assign n11158 = pi314 & n11084;
  assign n11159 = n11157 & n11158;
  assign n11160 = n11085 & n11159;
  assign n11161 = ~n11156 & n11160;
  assign n11162 = pi219 & ~n11161;
  assign n11163 = n2614 & n7309;
  assign n11164 = pi199 & ~pi299;
  assign n11165 = n2466 & n11159;
  assign n11166 = n3257 & n11165;
  assign n11167 = n11164 & n11166;
  assign n11168 = n11163 & n11167;
  assign n11169 = ~pi219 & ~n11168;
  assign n11170 = ~po1038 & ~n11169;
  assign po224 = ~n11162 & n11170;
  assign n11172 = pi83 & ~pi103;
  assign n11173 = n10895 & n11172;
  assign n11174 = n2465 & n11158;
  assign n11175 = n9986 & n11174;
  assign n11176 = n2485 & n11175;
  assign po225 = n11173 & n11176;
  assign n11178 = ~n6200 & n6448;
  assign n11179 = n3300 & n5975;
  assign n11180 = n11178 & n11179;
  assign n11181 = ~n6238 & n6448;
  assign n11182 = n3332 & n5792;
  assign n11183 = n11181 & n11182;
  assign n11184 = ~n11180 & ~n11183;
  assign po226 = n10780 & ~n11184;
  assign n11186 = n2782 & n8773;
  assign n11187 = pi69 & n8757;
  assign n11188 = n9979 & n11187;
  assign n11189 = ~pi71 & ~n11188;
  assign n11190 = n11186 & ~n11189;
  assign n11191 = ~pi314 & n2466;
  assign n11192 = n11190 & n11191;
  assign n11193 = pi71 & n2464;
  assign n11194 = pi314 & n11193;
  assign n11195 = n2486 & n11194;
  assign n11196 = n9975 & n11195;
  assign n11197 = ~n11192 & ~n11196;
  assign po227 = n10900 & ~n11197;
  assign n11199 = pi24 & n10016;
  assign n11200 = n2520 & n2744;
  assign n11201 = ~pi96 & n11200;
  assign n11202 = n2686 & n11201;
  assign n11203 = n11199 & n11202;
  assign n11204 = pi198 & pi589;
  assign n11205 = ~pi299 & ~n6238;
  assign n11206 = n2608 & n11205;
  assign n11207 = n11204 & n11206;
  assign n11208 = pi210 & pi589;
  assign n11209 = n2527 & n5975;
  assign n11210 = ~n6200 & n11209;
  assign n11211 = n11208 & n11210;
  assign n11212 = ~n11207 & ~n11211;
  assign n11213 = n6441 & ~n11212;
  assign n11214 = ~n6453 & n11213;
  assign n11215 = ~pi593 & n11214;
  assign n11216 = ~pi287 & ~n11215;
  assign n11217 = pi39 & ~n11216;
  assign n11218 = n2522 & n11217;
  assign n11219 = ~n11203 & ~n11218;
  assign po228 = n10024 & ~n11219;
  assign n11221 = ~pi199 & pi200;
  assign n11222 = ~pi299 & n11221;
  assign n11223 = pi211 & ~pi219;
  assign n11224 = pi299 & n11223;
  assign n11225 = ~n11222 & ~n11224;
  assign n11226 = pi314 & ~n11225;
  assign n11227 = n2470 & n2474;
  assign n11228 = n6309 & n11227;
  assign n11229 = n10803 & n11228;
  assign n11230 = ~pi64 & n8760;
  assign n11231 = n11229 & n11230;
  assign n11232 = ~pi81 & ~n11231;
  assign n11233 = n9987 & ~n11232;
  assign n11234 = ~pi50 & n8781;
  assign n11235 = n6331 & n11234;
  assign n11236 = n11233 & n11235;
  assign n11237 = n11226 & n11236;
  assign n11238 = n10810 & n11174;
  assign n11239 = n11229 & n11238;
  assign n11240 = n11225 & n11239;
  assign n11241 = ~n11237 & ~n11240;
  assign po229 = n9986 & ~n11241;
  assign n11243 = pi72 & n10015;
  assign n11244 = pi88 & n2862;
  assign n11245 = n9971 & n11244;
  assign n11246 = n6452 & n11245;
  assign n11247 = n9078 & n11246;
  assign n11248 = ~n11243 & ~n11247;
  assign n11249 = n3084 & ~n11248;
  assign n11250 = ~pi39 & ~n11249;
  assign n11251 = n7466 & n11181;
  assign n11252 = n7469 & n11178;
  assign n11253 = ~n11251 & ~n11252;
  assign n11254 = pi39 & n11253;
  assign n11255 = n10024 & ~n11254;
  assign po230 = ~n11250 & n11255;
  assign n11257 = n8973 & n11181;
  assign n11258 = ~pi299 & ~n11257;
  assign n11259 = n8959 & n11178;
  assign n11260 = pi299 & ~n11259;
  assign n11261 = ~n11258 & ~n11260;
  assign n11262 = pi39 & ~n11261;
  assign n11263 = ~pi314 & pi1050;
  assign n11264 = n3084 & n9413;
  assign n11265 = n11263 & n11264;
  assign n11266 = ~pi39 & ~n11265;
  assign n11267 = n10024 & ~n11266;
  assign po231 = ~n11262 & n11267;
  assign n11269 = ~pi96 & n7368;
  assign n11270 = ~pi1093 & n11269;
  assign n11271 = n7380 & ~n11270;
  assign n11272 = ~pi96 & ~n6166;
  assign n11273 = pi479 & ~n11272;
  assign n11274 = ~po840 & ~n11273;
  assign n11275 = n2728 & n7439;
  assign n11276 = ~pi96 & ~n11275;
  assign n11277 = n3345 & ~n11276;
  assign n11278 = n11274 & n11277;
  assign n11279 = n7407 & n11278;
  assign n11280 = n11271 & n11279;
  assign n11281 = n2572 & n10018;
  assign n11282 = pi74 & n11281;
  assign n11283 = n6525 & n11282;
  assign n11284 = ~n11280 & ~n11283;
  assign po232 = ~po1038 & ~n11284;
  assign n11286 = pi1093 & n11275;
  assign n11287 = ~pi96 & ~n11286;
  assign n11288 = n3258 & ~n11287;
  assign n11289 = ~n6207 & n11288;
  assign n11290 = n7448 & n11289;
  assign n11291 = ~pi75 & ~n11290;
  assign n11292 = pi75 & ~n11281;
  assign n11293 = n8739 & ~n11292;
  assign po233 = ~n11291 & n11293;
  assign n11295 = ~pi94 & ~n8785;
  assign n11296 = ~n8784 & ~n10170;
  assign n11297 = ~n11295 & ~n11296;
  assign n11298 = n9987 & n11297;
  assign n11299 = ~n7447 & ~n11298;
  assign n11300 = ~pi252 & n11298;
  assign n11301 = n8779 & n9993;
  assign n11302 = pi252 & n11301;
  assign n11303 = n7447 & ~n11302;
  assign n11304 = ~n11300 & n11303;
  assign n11305 = ~n11299 & ~n11304;
  assign n11306 = pi122 & ~n11305;
  assign n11307 = n3085 & n10171;
  assign n11308 = n7447 & ~n11307;
  assign n11309 = pi252 & n7447;
  assign n11310 = ~n11299 & ~n11309;
  assign n11311 = ~n11308 & n11310;
  assign n11312 = n7369 & ~n11311;
  assign n11313 = ~n11306 & ~n11312;
  assign n11314 = n2914 & ~n11313;
  assign n11315 = ~pi1093 & ~n11305;
  assign n11316 = n6207 & ~n11298;
  assign n11317 = ~n11315 & ~n11316;
  assign n11318 = ~n11314 & n11317;
  assign n11319 = ~po1057 & n11318;
  assign n11320 = po1057 & n11301;
  assign n11321 = ~n9929 & n11320;
  assign n11322 = ~n11319 & ~n11321;
  assign n11323 = pi210 & ~n11322;
  assign n11324 = pi1093 & ~n11298;
  assign n11325 = ~pi137 & ~n11311;
  assign n11326 = pi137 & n11315;
  assign n11327 = ~n11325 & ~n11326;
  assign n11328 = ~pi1093 & ~n11327;
  assign n11329 = ~n11324 & ~n11328;
  assign n11330 = ~po1057 & n11329;
  assign n11331 = ~n11320 & ~n11330;
  assign n11332 = ~pi137 & po1057;
  assign n11333 = n8752 & n11332;
  assign n11334 = ~n2914 & ~n11333;
  assign n11335 = ~n11331 & n11334;
  assign n11336 = pi137 & ~n11313;
  assign n11337 = n11327 & ~n11336;
  assign n11338 = ~po1057 & ~n11337;
  assign n11339 = pi137 & ~n7369;
  assign n11340 = n7447 & ~n11339;
  assign n11341 = n11301 & ~n11340;
  assign n11342 = po1057 & ~n11341;
  assign n11343 = n2914 & ~n11342;
  assign n11344 = ~n11338 & n11343;
  assign n11345 = ~n11335 & ~n11344;
  assign n11346 = ~pi210 & ~n11345;
  assign n11347 = ~n11323 & ~n11346;
  assign n11348 = n2626 & n10118;
  assign n11349 = ~n11347 & ~n11348;
  assign n11350 = ~n6207 & ~n11337;
  assign n11351 = ~n11316 & ~n11350;
  assign n11352 = ~pi210 & ~n11351;
  assign n11353 = pi210 & ~n11318;
  assign n11354 = ~n11352 & ~n11353;
  assign n11355 = n11348 & n11354;
  assign n11356 = pi299 & ~n11355;
  assign n11357 = ~n11349 & n11356;
  assign n11358 = pi198 & ~n11322;
  assign n11359 = ~pi198 & ~n11345;
  assign n11360 = ~n11358 & ~n11359;
  assign n11361 = n2658 & n6190;
  assign n11362 = ~n11360 & ~n11361;
  assign n11363 = ~pi198 & ~n11351;
  assign n11364 = pi198 & ~n11318;
  assign n11365 = n11361 & ~n11364;
  assign n11366 = ~n11363 & n11365;
  assign n11367 = ~pi299 & ~n11366;
  assign n11368 = ~n11362 & n11367;
  assign n11369 = ~n11357 & ~n11368;
  assign n11370 = pi232 & ~n11369;
  assign n11371 = ~pi299 & ~n11360;
  assign n11372 = pi299 & ~n11347;
  assign n11373 = ~pi232 & ~n11372;
  assign n11374 = ~n11371 & n11373;
  assign n11375 = ~n11370 & ~n11374;
  assign n11376 = ~n7376 & ~n11375;
  assign n11377 = ~n9927 & n11301;
  assign n11378 = po1057 & ~n11377;
  assign n11379 = n11307 & ~n11309;
  assign n11380 = ~pi137 & n11379;
  assign n11381 = ~pi137 & n2914;
  assign n11382 = n7368 & n11299;
  assign n11383 = ~n6122 & ~n11307;
  assign n11384 = ~n11304 & ~n11383;
  assign n11385 = ~n11382 & n11384;
  assign n11386 = ~pi122 & ~n11385;
  assign n11387 = ~n11306 & ~n11386;
  assign n11388 = ~pi1093 & ~n11387;
  assign n11389 = ~pi122 & ~n11379;
  assign n11390 = ~n11306 & ~n11389;
  assign n11391 = pi1093 & ~n11390;
  assign n11392 = ~n11388 & ~n11391;
  assign n11393 = n2914 & ~n11392;
  assign n11394 = ~n11381 & ~n11393;
  assign n11395 = ~n11380 & ~n11394;
  assign n11396 = ~pi122 & n11307;
  assign n11397 = ~n7369 & ~n11324;
  assign n11398 = ~n11396 & ~n11397;
  assign n11399 = ~n11388 & ~n11398;
  assign n11400 = ~n2914 & ~n11399;
  assign n11401 = ~pi137 & ~n2914;
  assign n11402 = ~n11400 & ~n11401;
  assign n11403 = pi252 & pi1092;
  assign n11404 = ~pi1093 & n11403;
  assign n11405 = n2935 & n11404;
  assign n11406 = ~pi137 & ~n11405;
  assign n11407 = n11307 & n11406;
  assign n11408 = ~n11402 & ~n11407;
  assign n11409 = ~n11395 & ~n11408;
  assign n11410 = ~po1057 & ~n11409;
  assign n11411 = ~n11332 & ~n11410;
  assign n11412 = ~n11378 & n11411;
  assign n11413 = ~pi210 & ~n11412;
  assign n11414 = ~n11393 & ~n11400;
  assign n11415 = ~po1057 & ~n11414;
  assign n11416 = ~n11378 & ~n11415;
  assign n11417 = pi210 & ~n11416;
  assign n11418 = ~n11413 & ~n11417;
  assign n11419 = ~n11348 & ~n11418;
  assign n11420 = ~pi210 & n11409;
  assign n11421 = n11348 & ~n11420;
  assign n11422 = pi210 & n11414;
  assign n11423 = n11421 & ~n11422;
  assign n11424 = pi299 & ~n11423;
  assign n11425 = ~n11419 & n11424;
  assign n11426 = ~pi198 & ~n11412;
  assign n11427 = pi198 & ~n11416;
  assign n11428 = ~n11426 & ~n11427;
  assign n11429 = ~n11361 & ~n11428;
  assign n11430 = ~pi198 & n11409;
  assign n11431 = n11361 & ~n11430;
  assign n11432 = pi198 & n11414;
  assign n11433 = n11431 & ~n11432;
  assign n11434 = ~pi299 & ~n11433;
  assign n11435 = ~n11429 & n11434;
  assign n11436 = ~n11425 & ~n11435;
  assign n11437 = pi232 & ~n11436;
  assign n11438 = ~pi299 & ~n11428;
  assign n11439 = pi299 & ~n11418;
  assign n11440 = ~pi232 & ~n11439;
  assign n11441 = ~n11438 & n11440;
  assign n11442 = n7376 & ~n11441;
  assign n11443 = ~n11437 & n11442;
  assign n11444 = n9986 & ~n11443;
  assign po234 = ~n11376 & n11444;
  assign n11446 = n2760 & n2775;
  assign n11447 = ~pi86 & ~n11446;
  assign n11448 = n6338 & ~n11447;
  assign n11449 = n2694 & n11448;
  assign n11450 = ~pi314 & ~n11449;
  assign n11451 = pi86 & n8784;
  assign n11452 = n2764 & n11451;
  assign n11453 = pi314 & ~n11452;
  assign n11454 = n9988 & ~n11453;
  assign po235 = ~n11450 & n11454;
  assign n11456 = pi119 & pi232;
  assign po236 = ~pi468 & n11456;
  assign n11458 = ~pi34 & n9533;
  assign n11459 = pi163 & ~n9543;
  assign n11460 = ~pi163 & ~n9539;
  assign n11461 = ~n9541 & n11460;
  assign n11462 = ~n11459 & ~n11461;
  assign n11463 = pi232 & n11462;
  assign n11464 = ~n7255 & n11463;
  assign n11465 = pi74 & ~n11464;
  assign n11466 = pi75 & ~n11463;
  assign n11467 = pi100 & ~n11463;
  assign n11468 = ~n11466 & ~n11467;
  assign n11469 = pi147 & n7420;
  assign n11470 = n7255 & n11469;
  assign n11471 = n11468 & ~n11470;
  assign n11472 = ~n11465 & n11471;
  assign n11473 = ~n3327 & n11472;
  assign n11474 = pi54 & ~n11471;
  assign n11475 = ~pi38 & ~pi40;
  assign n11476 = pi38 & ~n11469;
  assign n11477 = ~pi100 & ~n11476;
  assign n11478 = ~n11475 & n11477;
  assign n11479 = ~n11467 & ~n11478;
  assign n11480 = ~pi75 & ~n11479;
  assign n11481 = ~n11466 & ~n11480;
  assign n11482 = ~pi54 & ~n11481;
  assign n11483 = ~n11474 & ~n11482;
  assign n11484 = ~pi74 & ~n11483;
  assign n11485 = ~n11465 & ~n11484;
  assign n11486 = ~n2531 & ~n11485;
  assign n11487 = n3327 & ~n11486;
  assign n11488 = pi55 & ~n11465;
  assign n11489 = pi39 & ~n9165;
  assign n11490 = n7254 & ~n11489;
  assign n11491 = n2488 & ~n8879;
  assign n11492 = ~pi40 & ~n11491;
  assign n11493 = pi163 & pi232;
  assign n11494 = ~n6190 & n8879;
  assign n11495 = n8862 & ~n11494;
  assign n11496 = n11493 & n11495;
  assign n11497 = n11492 & ~n11496;
  assign n11498 = ~pi39 & ~n11497;
  assign n11499 = n11490 & ~n11498;
  assign n11500 = pi87 & ~n2488;
  assign n11501 = n11475 & n11500;
  assign n11502 = ~n11499 & ~n11501;
  assign n11503 = n11477 & n11502;
  assign n11504 = ~n11467 & ~n11503;
  assign n11505 = n2573 & ~n11504;
  assign n11506 = ~n8940 & n11479;
  assign n11507 = n8930 & ~n11506;
  assign n11508 = ~n11466 & ~n11507;
  assign n11509 = ~n11505 & n11508;
  assign n11510 = ~pi54 & ~n11509;
  assign n11511 = ~n11474 & ~n11510;
  assign n11512 = ~pi74 & ~n11511;
  assign n11513 = n11488 & ~n11512;
  assign n11514 = pi299 & ~n11462;
  assign n11515 = ~n9568 & n9570;
  assign n11516 = ~pi184 & n11515;
  assign n11517 = pi184 & n6190;
  assign n11518 = ~n11515 & n11517;
  assign n11519 = ~pi299 & ~n11518;
  assign n11520 = ~n11516 & n11519;
  assign n11521 = pi232 & ~n11520;
  assign n11522 = ~n11514 & n11521;
  assign n11523 = ~n7255 & n11522;
  assign n11524 = pi74 & ~n11523;
  assign n11525 = ~pi55 & ~n11524;
  assign n11526 = ~pi187 & ~pi299;
  assign n11527 = ~n8924 & ~n11469;
  assign n11528 = ~n11526 & ~n11527;
  assign n11529 = n7255 & ~n11528;
  assign n11530 = pi54 & ~n11529;
  assign n11531 = ~n11523 & n11530;
  assign n11532 = pi100 & ~n11522;
  assign n11533 = pi38 & ~n11528;
  assign n11534 = ~pi100 & ~n11533;
  assign n11535 = ~n11501 & n11534;
  assign n11536 = ~pi179 & ~pi299;
  assign n11537 = ~pi156 & pi299;
  assign n11538 = n7420 & ~n11537;
  assign n11539 = ~n11536 & n11538;
  assign n11540 = n2488 & n11539;
  assign n11541 = n11492 & ~n11540;
  assign n11542 = ~pi39 & ~n11541;
  assign n11543 = n11490 & ~n11542;
  assign n11544 = n11535 & ~n11543;
  assign n11545 = ~n11532 & ~n11544;
  assign n11546 = n8930 & ~n11545;
  assign n11547 = pi75 & ~n11522;
  assign n11548 = ~pi187 & ~n8948;
  assign n11549 = pi187 & ~n8950;
  assign n11550 = pi147 & ~n11549;
  assign n11551 = ~n11548 & n11550;
  assign n11552 = ~pi147 & pi187;
  assign n11553 = n8954 & n11552;
  assign n11554 = ~n11551 & ~n11553;
  assign n11555 = pi38 & ~n11554;
  assign n11556 = ~n8973 & ~n9165;
  assign n11557 = ~pi40 & ~n8967;
  assign n11558 = ~pi189 & ~n11557;
  assign n11559 = n2488 & ~n8982;
  assign n11560 = n9141 & ~n11559;
  assign n11561 = n6215 & n9165;
  assign n11562 = n2488 & ~n8965;
  assign n11563 = ~pi40 & ~n11562;
  assign n11564 = n6191 & n11563;
  assign n11565 = ~n11561 & ~n11564;
  assign n11566 = ~n11560 & n11565;
  assign n11567 = pi189 & ~n6236;
  assign n11568 = n11566 & n11567;
  assign n11569 = ~n11558 & ~n11568;
  assign n11570 = pi179 & ~n11569;
  assign n11571 = n6236 & ~n11557;
  assign n11572 = n2488 & ~n8988;
  assign n11573 = n9141 & ~n11572;
  assign n11574 = n11565 & ~n11573;
  assign n11575 = ~pi189 & ~n11574;
  assign n11576 = ~n6215 & n11563;
  assign n11577 = ~n11561 & ~n11576;
  assign n11578 = pi189 & ~n11577;
  assign n11579 = ~n11575 & ~n11578;
  assign n11580 = ~pi179 & n11579;
  assign n11581 = ~n6236 & n11580;
  assign n11582 = ~n11571 & ~n11581;
  assign n11583 = ~n11570 & n11582;
  assign n11584 = n8973 & ~n11583;
  assign n11585 = ~n11556 & ~n11584;
  assign n11586 = ~pi299 & ~n11585;
  assign n11587 = ~n8959 & n9165;
  assign n11588 = pi299 & ~n11587;
  assign n11589 = ~pi166 & ~n6198;
  assign n11590 = n6198 & ~n11557;
  assign n11591 = ~n6198 & n11577;
  assign n11592 = ~n11590 & ~n11591;
  assign n11593 = ~n11589 & ~n11592;
  assign n11594 = n11574 & n11589;
  assign n11595 = ~n11593 & ~n11594;
  assign n11596 = n8959 & n11595;
  assign n11597 = n11588 & ~n11596;
  assign n11598 = ~n11586 & ~n11597;
  assign n11599 = ~pi156 & ~n11598;
  assign n11600 = pi232 & n11599;
  assign n11601 = ~n6236 & n11577;
  assign n11602 = ~n11571 & ~n11601;
  assign n11603 = n8973 & ~n11602;
  assign n11604 = ~pi299 & ~n11556;
  assign n11605 = ~n11603 & n11604;
  assign n11606 = n8961 & n11592;
  assign n11607 = ~pi232 & ~n11606;
  assign n11608 = ~n11605 & n11607;
  assign n11609 = pi39 & ~n11608;
  assign n11610 = ~n11600 & n11609;
  assign n11611 = pi166 & ~n6198;
  assign n11612 = ~n11557 & ~n11611;
  assign n11613 = n11566 & n11611;
  assign n11614 = ~n11612 & ~n11613;
  assign n11615 = n8959 & n11614;
  assign n11616 = n11588 & ~n11615;
  assign n11617 = ~n11586 & ~n11616;
  assign n11618 = pi156 & ~n11617;
  assign n11619 = pi232 & n11618;
  assign n11620 = n11610 & ~n11619;
  assign n11621 = ~n2442 & ~n9183;
  assign n11622 = n9018 & ~n9020;
  assign n11623 = ~n11621 & ~n11622;
  assign n11624 = ~pi40 & ~n9160;
  assign n11625 = ~pi95 & ~n11624;
  assign n11626 = ~pi166 & n11264;
  assign n11627 = ~n11625 & ~n11626;
  assign n11628 = pi153 & ~n11627;
  assign n11629 = ~pi40 & ~n9115;
  assign n11630 = ~pi95 & ~n11629;
  assign n11631 = ~pi40 & ~n9130;
  assign n11632 = pi166 & n11631;
  assign n11633 = n11630 & ~n11632;
  assign n11634 = ~pi153 & n11633;
  assign n11635 = n6190 & ~n11634;
  assign n11636 = ~n11628 & n11635;
  assign n11637 = ~pi160 & n11636;
  assign n11638 = ~n11623 & n11637;
  assign n11639 = pi166 & n6190;
  assign n11640 = ~n9183 & n11639;
  assign n11641 = ~n11625 & n11640;
  assign n11642 = n9165 & n10118;
  assign n11643 = pi153 & ~n11642;
  assign n11644 = ~n11641 & n11643;
  assign n11645 = pi160 & ~n11644;
  assign n11646 = ~n9183 & n11635;
  assign n11647 = ~pi153 & ~n11646;
  assign n11648 = n11645 & ~n11647;
  assign n11649 = pi163 & ~n11648;
  assign n11650 = ~n11638 & n11649;
  assign n11651 = ~n9211 & ~n11623;
  assign n11652 = pi210 & ~n11651;
  assign n11653 = ~n9215 & ~n11623;
  assign n11654 = ~pi210 & ~n11653;
  assign n11655 = n10118 & ~n11654;
  assign n11656 = ~n11652 & n11655;
  assign n11657 = ~pi95 & ~n9178;
  assign n11658 = ~n11623 & ~n11657;
  assign n11659 = pi210 & ~n11658;
  assign n11660 = ~n9187 & ~n11623;
  assign n11661 = ~pi210 & ~n11660;
  assign n11662 = n11639 & ~n11661;
  assign n11663 = ~n11659 & n11662;
  assign n11664 = ~n11656 & ~n11663;
  assign n11665 = pi153 & n11664;
  assign n11666 = ~pi40 & ~n9266;
  assign n11667 = ~pi95 & ~n11666;
  assign n11668 = ~n11623 & ~n11667;
  assign n11669 = pi166 & n11668;
  assign n11670 = ~pi40 & n9091;
  assign n11671 = ~pi32 & ~n11670;
  assign n11672 = ~n9166 & ~n11671;
  assign n11673 = ~pi95 & ~n11672;
  assign n11674 = ~n9183 & ~n11673;
  assign n11675 = pi210 & ~n11674;
  assign n11676 = ~n9185 & ~n11671;
  assign n11677 = ~pi95 & ~n11676;
  assign n11678 = ~n9183 & ~n11677;
  assign n11679 = ~pi210 & ~n11678;
  assign n11680 = ~n11675 & ~n11679;
  assign n11681 = ~pi95 & ~n11680;
  assign n11682 = ~n11623 & ~n11681;
  assign n11683 = n10118 & n11682;
  assign n11684 = ~pi153 & ~n11683;
  assign n11685 = ~n11669 & n11684;
  assign n11686 = ~pi160 & ~n11685;
  assign n11687 = ~n11665 & n11686;
  assign n11688 = n11639 & n11666;
  assign n11689 = n10118 & n11680;
  assign n11690 = ~pi153 & ~n11689;
  assign n11691 = ~n11688 & n11690;
  assign n11692 = n9284 & n10118;
  assign n11693 = ~n9183 & ~n11657;
  assign n11694 = pi210 & ~n11693;
  assign n11695 = ~pi210 & ~n9188;
  assign n11696 = n11639 & ~n11695;
  assign n11697 = ~n11694 & n11696;
  assign n11698 = pi153 & ~n11697;
  assign n11699 = ~n11692 & n11698;
  assign n11700 = ~n11691 & ~n11699;
  assign n11701 = pi160 & n11700;
  assign n11702 = ~pi163 & ~n11701;
  assign n11703 = ~n11687 & n11702;
  assign n11704 = ~n11650 & ~n11703;
  assign n11705 = ~n6190 & n11668;
  assign n11706 = pi299 & ~n11705;
  assign n11707 = ~n11704 & n11706;
  assign n11708 = ~pi40 & ~n9143;
  assign n11709 = ~pi95 & ~n11708;
  assign n11710 = ~n11623 & ~n11709;
  assign n11711 = ~n6190 & n11710;
  assign n11712 = ~pi175 & ~pi299;
  assign n11713 = pi189 & n11631;
  assign n11714 = n11630 & ~n11713;
  assign n11715 = ~pi182 & n11623;
  assign n11716 = pi182 & n9183;
  assign n11717 = n6190 & ~n11716;
  assign n11718 = ~n11715 & n11717;
  assign n11719 = ~n11714 & n11718;
  assign n11720 = pi184 & ~n11719;
  assign n11721 = ~pi198 & ~n11678;
  assign n11722 = pi198 & ~n11674;
  assign n11723 = ~n11721 & ~n11722;
  assign n11724 = n10122 & n11723;
  assign n11725 = pi189 & n6190;
  assign n11726 = n11708 & n11725;
  assign n11727 = ~pi184 & ~n11726;
  assign n11728 = pi182 & n11727;
  assign n11729 = ~n11724 & n11728;
  assign n11730 = ~n11720 & ~n11729;
  assign n11731 = n11712 & ~n11730;
  assign n11732 = ~pi198 & ~n9188;
  assign n11733 = pi198 & ~n11693;
  assign n11734 = ~n11732 & ~n11733;
  assign n11735 = n11725 & n11734;
  assign n11736 = n9218 & n10122;
  assign n11737 = pi182 & ~n11736;
  assign n11738 = ~n11735 & n11737;
  assign n11739 = ~pi95 & ~n11734;
  assign n11740 = ~n11623 & ~n11739;
  assign n11741 = n11725 & n11740;
  assign n11742 = ~pi182 & ~n11741;
  assign n11743 = ~n11738 & ~n11742;
  assign n11744 = pi95 & ~pi182;
  assign n11745 = ~n9218 & ~n11744;
  assign n11746 = ~n11623 & ~n11745;
  assign n11747 = n10122 & n11746;
  assign n11748 = ~n11743 & ~n11747;
  assign n11749 = ~pi184 & ~n11748;
  assign n11750 = pi175 & ~pi299;
  assign n11751 = ~n11749 & n11750;
  assign n11752 = ~pi95 & pi189;
  assign n11753 = n2488 & ~n11752;
  assign n11754 = n11624 & ~n11753;
  assign n11755 = ~n11744 & ~n11754;
  assign n11756 = ~n11715 & ~n11755;
  assign n11757 = n11517 & n11756;
  assign n11758 = n11751 & ~n11757;
  assign n11759 = ~n11731 & ~n11758;
  assign n11760 = ~n11711 & ~n11759;
  assign n11761 = ~n10122 & n11710;
  assign n11762 = ~pi184 & ~pi299;
  assign n11763 = ~pi95 & ~n11723;
  assign n11764 = ~n11623 & ~n11763;
  assign n11765 = n10122 & n11764;
  assign n11766 = n11762 & ~n11765;
  assign n11767 = ~n11761 & n11766;
  assign n11768 = ~pi175 & n11767;
  assign n11769 = ~pi182 & n11768;
  assign n11770 = ~n11760 & ~n11769;
  assign n11771 = ~n11707 & n11770;
  assign n11772 = pi232 & ~n11771;
  assign n11773 = ~pi299 & n11710;
  assign n11774 = pi299 & n11668;
  assign n11775 = ~pi232 & ~n11774;
  assign n11776 = ~n11773 & n11775;
  assign n11777 = ~n11772 & ~n11776;
  assign n11778 = ~pi39 & n11777;
  assign n11779 = ~pi38 & ~n11778;
  assign n11780 = ~n11620 & n11779;
  assign n11781 = ~n11555 & ~n11780;
  assign n11782 = n2571 & ~n11781;
  assign n11783 = pi87 & n11535;
  assign n11784 = ~n11532 & ~n11783;
  assign n11785 = ~n11782 & n11784;
  assign n11786 = n2573 & ~n11785;
  assign n11787 = ~n11547 & ~n11786;
  assign n11788 = ~n11546 & n11787;
  assign n11789 = ~pi54 & ~n11788;
  assign n11790 = ~n11531 & ~n11789;
  assign n11791 = ~pi74 & ~n11790;
  assign n11792 = n11525 & ~n11791;
  assign n11793 = ~n11513 & ~n11792;
  assign n11794 = n2531 & n11793;
  assign n11795 = ~n8866 & ~n11794;
  assign n11796 = n11487 & n11795;
  assign n11797 = ~n11473 & ~n11796;
  assign n11798 = ~pi79 & n11797;
  assign n11799 = ~n11458 & ~n11798;
  assign n11800 = ~pi87 & n11539;
  assign n11801 = n2510 & n11800;
  assign n11802 = n10016 & n11801;
  assign n11803 = n11475 & ~n11802;
  assign n11804 = n11534 & ~n11803;
  assign n11805 = ~n11532 & ~n11804;
  assign n11806 = n8930 & ~n11805;
  assign n11807 = pi184 & n9474;
  assign n11808 = ~pi184 & ~n9419;
  assign n11809 = ~pi189 & ~n11808;
  assign n11810 = ~n11807 & n11809;
  assign n11811 = ~pi32 & pi95;
  assign n11812 = ~pi479 & n2510;
  assign n11813 = n11811 & n11812;
  assign n11814 = pi182 & n11813;
  assign n11815 = pi184 & ~n9472;
  assign n11816 = pi189 & n11815;
  assign n11817 = ~n11814 & ~n11816;
  assign n11818 = ~n11810 & n11817;
  assign n11819 = n6190 & ~n11818;
  assign n11820 = ~pi40 & ~n11819;
  assign n11821 = n11712 & ~n11820;
  assign n11822 = pi189 & ~n9408;
  assign n11823 = ~n9414 & ~n11822;
  assign n11824 = n2516 & n11823;
  assign n11825 = ~n11814 & ~n11824;
  assign n11826 = n6190 & ~n11825;
  assign n11827 = ~pi184 & ~n11826;
  assign n11828 = ~n9466 & n11725;
  assign n11829 = pi184 & ~n11828;
  assign n11830 = ~n9459 & n10122;
  assign n11831 = ~pi182 & ~n11830;
  assign n11832 = n11829 & n11831;
  assign n11833 = ~n11827 & ~n11832;
  assign n11834 = ~pi40 & ~n11833;
  assign n11835 = ~pi40 & ~n11813;
  assign n11836 = ~n9437 & n11835;
  assign n11837 = ~n9458 & n11836;
  assign n11838 = n10122 & ~n11837;
  assign n11839 = pi184 & ~n11838;
  assign n11840 = n9466 & n11835;
  assign n11841 = n11725 & ~n11840;
  assign n11842 = pi182 & ~n11841;
  assign n11843 = pi40 & ~n6190;
  assign n11844 = n11842 & ~n11843;
  assign n11845 = n11839 & n11844;
  assign n11846 = n11750 & ~n11845;
  assign n11847 = ~n11834 & n11846;
  assign n11848 = ~n11821 & ~n11847;
  assign n11849 = n9434 & n11835;
  assign n11850 = n10118 & ~n11849;
  assign n11851 = n9448 & n11835;
  assign n11852 = n11639 & ~n11851;
  assign n11853 = ~pi153 & ~n11852;
  assign n11854 = ~n11850 & n11853;
  assign n11855 = pi153 & n9445;
  assign n11856 = n9448 & ~n11855;
  assign n11857 = n11639 & ~n11856;
  assign n11858 = ~pi210 & ~n9457;
  assign n11859 = n11836 & ~n11858;
  assign n11860 = n10118 & ~n11859;
  assign n11861 = ~n11852 & ~n11860;
  assign n11862 = ~n11853 & n11861;
  assign n11863 = ~n11857 & n11862;
  assign n11864 = ~n11854 & ~n11863;
  assign n11865 = ~n11843 & ~n11864;
  assign n11866 = pi163 & n11865;
  assign n11867 = pi160 & ~n11866;
  assign n11868 = pi153 & n9408;
  assign n11869 = n9409 & n11868;
  assign n11870 = n9419 & n10118;
  assign n11871 = ~pi163 & ~n11870;
  assign n11872 = ~pi40 & n11871;
  assign n11873 = ~n11869 & n11872;
  assign n11874 = pi153 & n9437;
  assign n11875 = n9434 & ~n11874;
  assign n11876 = n10118 & ~n11875;
  assign n11877 = pi163 & ~n11876;
  assign n11878 = ~pi40 & n11877;
  assign n11879 = ~n11857 & n11878;
  assign n11880 = ~pi160 & ~n11879;
  assign n11881 = ~n11873 & n11880;
  assign n11882 = ~n11867 & ~n11881;
  assign n11883 = n6190 & n11813;
  assign n11884 = n11873 & ~n11883;
  assign n11885 = pi299 & ~n11884;
  assign n11886 = ~n11882 & n11885;
  assign n11887 = n11848 & ~n11886;
  assign n11888 = ~pi39 & ~n11887;
  assign n11889 = n2510 & n9409;
  assign n11890 = ~pi189 & n8963;
  assign n11891 = pi179 & n6182;
  assign n11892 = ~n11890 & ~n11891;
  assign n11893 = n9384 & ~n11892;
  assign n11894 = n11889 & n11893;
  assign n11895 = ~pi299 & n11894;
  assign n11896 = ~n6198 & n8959;
  assign n11897 = pi156 & n6182;
  assign n11898 = ~pi166 & n8963;
  assign n11899 = ~n11897 & ~n11898;
  assign n11900 = n11889 & ~n11899;
  assign n11901 = n11896 & n11900;
  assign n11902 = pi299 & n11901;
  assign n11903 = ~pi40 & ~n11902;
  assign n11904 = ~n11895 & n11903;
  assign n11905 = pi39 & ~n11904;
  assign n11906 = pi232 & ~n11905;
  assign n11907 = ~n11888 & n11906;
  assign n11908 = ~pi40 & ~pi232;
  assign n11909 = ~pi38 & ~n11908;
  assign n11910 = ~n11907 & n11909;
  assign n11911 = ~n11555 & ~n11910;
  assign n11912 = n2571 & ~n11911;
  assign n11913 = pi87 & ~n11475;
  assign n11914 = n11534 & n11913;
  assign n11915 = ~n11532 & ~n11914;
  assign n11916 = ~n11912 & n11915;
  assign n11917 = n2573 & ~n11916;
  assign n11918 = ~n11547 & ~n11917;
  assign n11919 = ~n11806 & n11918;
  assign n11920 = ~pi54 & ~n11919;
  assign n11921 = ~n11531 & ~n11920;
  assign n11922 = ~pi74 & ~n11921;
  assign n11923 = n11525 & ~n11922;
  assign n11924 = ~pi92 & n11889;
  assign n11925 = n3257 & n11924;
  assign n11926 = n11493 & n11925;
  assign n11927 = n11475 & ~n11926;
  assign n11928 = ~n11476 & ~n11927;
  assign n11929 = n7255 & n11928;
  assign n11930 = n11468 & ~n11929;
  assign n11931 = ~pi54 & ~n11930;
  assign n11932 = ~n11474 & ~n11931;
  assign n11933 = ~pi74 & ~n11932;
  assign n11934 = n11488 & ~n11933;
  assign n11935 = ~n11923 & ~n11934;
  assign n11936 = n2531 & n11935;
  assign n11937 = n11487 & ~n11936;
  assign n11938 = ~n11473 & ~n11937;
  assign n11939 = pi79 & n11938;
  assign n11940 = n11799 & ~n11939;
  assign n11941 = ~pi79 & ~n8832;
  assign n11942 = n11797 & ~n11941;
  assign n11943 = n11938 & n11941;
  assign n11944 = n11458 & ~n11943;
  assign n11945 = ~n11942 & n11944;
  assign po237 = n11940 | n11945;
  assign n11947 = pi98 & pi1092;
  assign n11948 = pi1093 & n11947;
  assign n11949 = ~pi567 & n2934;
  assign n11950 = ~n11948 & ~n11949;
  assign n11951 = n7376 & n11950;
  assign n11952 = ~n7958 & n11950;
  assign n11953 = pi588 & ~n11952;
  assign n11954 = n7669 & ~n8037;
  assign n11955 = n11950 & ~n11954;
  assign n11956 = ~pi1199 & ~n11955;
  assign n11957 = ~pi428 & n8037;
  assign n11958 = n7669 & ~n11957;
  assign n11959 = ~pi427 & n11958;
  assign n11960 = n11950 & ~n11959;
  assign n11961 = pi428 & n8037;
  assign n11962 = n7669 & ~n11961;
  assign n11963 = pi427 & n11962;
  assign n11964 = n11960 & ~n11963;
  assign n11965 = pi430 & ~n11964;
  assign n11966 = ~n8052 & ~n11955;
  assign n11967 = ~n7669 & n11950;
  assign n11968 = n8052 & ~n11967;
  assign n11969 = ~n11966 & ~n11968;
  assign n11970 = ~pi430 & ~n11969;
  assign n11971 = ~n11965 & ~n11970;
  assign n11972 = ~pi426 & ~n11971;
  assign n11973 = ~pi430 & ~n11964;
  assign n11974 = pi430 & ~n11969;
  assign n11975 = ~n11973 & ~n11974;
  assign n11976 = pi426 & ~n11975;
  assign n11977 = ~n11972 & ~n11976;
  assign n11978 = ~pi445 & ~n11977;
  assign n11979 = ~pi426 & ~n11975;
  assign n11980 = pi426 & ~n11971;
  assign n11981 = ~n11979 & ~n11980;
  assign n11982 = pi445 & ~n11981;
  assign n11983 = ~n11978 & ~n11982;
  assign n11984 = pi448 & ~n11983;
  assign n11985 = ~pi445 & ~n11981;
  assign n11986 = pi445 & ~n11977;
  assign n11987 = ~n11985 & ~n11986;
  assign n11988 = ~pi448 & ~n11987;
  assign n11989 = n8046 & ~n11988;
  assign n11990 = ~n11984 & n11989;
  assign n11991 = ~pi448 & ~n11983;
  assign n11992 = pi448 & ~n11987;
  assign n11993 = ~n8046 & ~n11992;
  assign n11994 = ~n11991 & n11993;
  assign n11995 = ~n11990 & ~n11994;
  assign n11996 = pi1199 & n11995;
  assign n11997 = ~n11956 & ~n11996;
  assign n11998 = n7958 & n11997;
  assign n11999 = n11953 & ~n11998;
  assign n12000 = pi591 & ~n11950;
  assign n12001 = pi590 & ~n12000;
  assign n12002 = ~n7677 & n11950;
  assign n12003 = n7673 & n12002;
  assign n12004 = ~n7589 & n12003;
  assign n12005 = ~n11967 & ~n12004;
  assign n12006 = pi461 & ~n12005;
  assign n12007 = ~n7700 & n12003;
  assign n12008 = ~n11967 & ~n12007;
  assign n12009 = ~pi461 & ~n12008;
  assign n12010 = ~n12006 & ~n12009;
  assign n12011 = n7696 & n12010;
  assign n12012 = pi461 & ~n12008;
  assign n12013 = ~pi461 & ~n12005;
  assign n12014 = ~n12012 & ~n12013;
  assign n12015 = ~n7696 & n12014;
  assign n12016 = ~n12011 & ~n12015;
  assign n12017 = ~pi354 & ~n12016;
  assign n12018 = ~pi357 & n12010;
  assign n12019 = pi356 & ~n12018;
  assign n12020 = pi357 & n12014;
  assign n12021 = n12019 & ~n12020;
  assign n12022 = ~pi357 & n12014;
  assign n12023 = ~pi356 & ~n12022;
  assign n12024 = pi357 & n12010;
  assign n12025 = n12023 & ~n12024;
  assign n12026 = ~n12021 & ~n12025;
  assign n12027 = pi354 & n12026;
  assign n12028 = ~n7690 & ~n12027;
  assign n12029 = ~n12017 & n12028;
  assign n12030 = ~pi354 & n12026;
  assign n12031 = pi354 & ~n12016;
  assign n12032 = n7690 & ~n12031;
  assign n12033 = ~n12030 & n12032;
  assign n12034 = ~pi591 & ~n12033;
  assign n12035 = ~n12029 & n12034;
  assign n12036 = n12001 & ~n12035;
  assign n12037 = ~n7819 & n11950;
  assign n12038 = ~pi591 & ~n12037;
  assign n12039 = ~pi1197 & ~n8293;
  assign n12040 = ~n11967 & ~n12039;
  assign n12041 = pi592 & ~n11950;
  assign n12042 = ~pi1196 & ~n11950;
  assign n12043 = ~n12041 & ~n12042;
  assign n12044 = pi411 & ~n7834;
  assign n12045 = ~pi411 & n7834;
  assign n12046 = ~n12044 & ~n12045;
  assign n12047 = n7840 & n12046;
  assign n12048 = ~n7840 & ~n12046;
  assign n12049 = ~n12047 & ~n12048;
  assign n12050 = n7368 & n12049;
  assign n12051 = ~n11947 & ~n12050;
  assign n12052 = ~pi412 & ~n12051;
  assign n12053 = n7368 & ~n12049;
  assign n12054 = ~n11947 & ~n12053;
  assign n12055 = pi412 & ~n12054;
  assign n12056 = n7831 & ~n12055;
  assign n12057 = ~n12052 & n12056;
  assign n12058 = pi412 & ~n12051;
  assign n12059 = ~pi412 & ~n12054;
  assign n12060 = ~n7831 & ~n12059;
  assign n12061 = ~n12058 & n12060;
  assign n12062 = ~pi122 & ~n12061;
  assign n12063 = ~n12057 & n12062;
  assign n12064 = ~n11947 & ~n12063;
  assign n12065 = n7490 & ~n12064;
  assign n12066 = pi1091 & n11948;
  assign n12067 = ~n12065 & ~n12066;
  assign n12068 = pi567 & ~n12067;
  assign n12069 = ~n11949 & ~n12068;
  assign n12070 = n7881 & ~n12069;
  assign n12071 = n12043 & ~n12070;
  assign n12072 = ~pi1199 & ~n12071;
  assign n12073 = n7368 & ~n7874;
  assign n12074 = ~pi122 & ~n11947;
  assign n12075 = ~n12073 & n12074;
  assign n12076 = ~n7371 & ~n11948;
  assign n12077 = ~n12075 & ~n12076;
  assign n12078 = pi567 & n12077;
  assign n12079 = ~n11949 & ~n12078;
  assign n12080 = ~n12068 & n12079;
  assign n12081 = n7881 & ~n12080;
  assign n12082 = n8608 & ~n12079;
  assign n12083 = ~n12041 & ~n12082;
  assign n12084 = ~n12081 & n12083;
  assign n12085 = pi1199 & ~n12084;
  assign n12086 = ~n12072 & ~n12085;
  assign n12087 = n12039 & ~n12086;
  assign n12088 = ~n12040 & ~n12087;
  assign n12089 = pi333 & ~n12088;
  assign n12090 = n8293 & ~n11967;
  assign n12091 = ~n8293 & ~n12086;
  assign n12092 = ~n12090 & ~n12091;
  assign n12093 = ~pi333 & ~n12092;
  assign n12094 = ~n12089 & ~n12093;
  assign n12095 = ~pi391 & ~n12094;
  assign n12096 = ~pi333 & ~n12088;
  assign n12097 = pi333 & ~n12092;
  assign n12098 = ~n12096 & ~n12097;
  assign n12099 = pi391 & ~n12098;
  assign n12100 = n7937 & ~n12099;
  assign n12101 = ~n12095 & n12100;
  assign n12102 = ~pi391 & ~n12098;
  assign n12103 = pi391 & ~n12094;
  assign n12104 = ~n7937 & ~n12103;
  assign n12105 = ~n12102 & n12104;
  assign n12106 = ~n12101 & ~n12105;
  assign n12107 = pi591 & n12106;
  assign n12108 = ~pi590 & ~n12107;
  assign n12109 = ~n12038 & n12108;
  assign n12110 = ~pi588 & ~n12109;
  assign n12111 = ~n12036 & n12110;
  assign n12112 = ~n7376 & ~n12111;
  assign n12113 = ~n11999 & n12112;
  assign n12114 = ~pi80 & ~n12113;
  assign n12115 = po1038 & n12114;
  assign n12116 = ~n11951 & n12115;
  assign n12117 = ~n7380 & n11950;
  assign n12118 = n7380 & ~n11949;
  assign n12119 = pi75 & n11948;
  assign n12120 = pi824 & pi950;
  assign n12121 = ~pi94 & n2464;
  assign n12122 = n2711 & n12121;
  assign n12123 = ~pi88 & n2494;
  assign n12124 = n2497 & n12123;
  assign n12125 = n2761 & n12124;
  assign n12126 = n12122 & n12125;
  assign n12127 = n7395 & n12126;
  assign n12128 = pi51 & n12127;
  assign n12129 = pi90 & pi93;
  assign n12130 = n2508 & ~n12129;
  assign n12131 = ~n2696 & n12130;
  assign n12132 = ~pi841 & n12131;
  assign n12133 = n12126 & n12132;
  assign n12134 = ~n12128 & ~n12133;
  assign n12135 = n12120 & ~n12134;
  assign n12136 = n2517 & n12135;
  assign n12137 = ~pi98 & ~n12136;
  assign n12138 = pi1092 & ~n12137;
  assign n12139 = ~n7490 & ~n12066;
  assign n12140 = n3258 & ~n12139;
  assign n12141 = n12138 & n12140;
  assign n12142 = ~pi51 & n2517;
  assign n12143 = n12120 & n12127;
  assign n12144 = n12142 & n12143;
  assign n12145 = ~pi98 & ~n12144;
  assign n12146 = pi1092 & ~n12145;
  assign n12147 = n8299 & ~n12139;
  assign n12148 = n12146 & n12147;
  assign n12149 = ~n2615 & n11948;
  assign n12150 = ~n12148 & ~n12149;
  assign n12151 = ~n12141 & n12150;
  assign n12152 = ~pi75 & ~n12151;
  assign n12153 = ~n12119 & ~n12152;
  assign n12154 = pi567 & ~n12153;
  assign n12155 = n12118 & ~n12154;
  assign n12156 = ~n12117 & ~n12155;
  assign n12157 = ~pi592 & n12156;
  assign n12158 = ~n12041 & ~n12157;
  assign n12159 = ~n8011 & n12158;
  assign n12160 = n8011 & ~n12042;
  assign n12161 = pi443 & ~n11950;
  assign n12162 = ~pi443 & ~n12158;
  assign n12163 = ~n12161 & ~n12162;
  assign n12164 = ~n8162 & n12163;
  assign n12165 = ~pi443 & ~n11950;
  assign n12166 = pi443 & ~n12158;
  assign n12167 = ~n12165 & ~n12166;
  assign n12168 = n8162 & n12167;
  assign n12169 = ~n12164 & ~n12168;
  assign n12170 = pi435 & ~n12169;
  assign n12171 = n8162 & n12163;
  assign n12172 = ~n8162 & n12167;
  assign n12173 = ~n12171 & ~n12172;
  assign n12174 = ~pi435 & ~n12173;
  assign n12175 = ~n12170 & ~n12174;
  assign n12176 = ~pi429 & n12175;
  assign n12177 = n8026 & ~n12176;
  assign n12178 = ~pi435 & ~n12169;
  assign n12179 = pi435 & ~n12173;
  assign n12180 = ~n12178 & ~n12179;
  assign n12181 = pi429 & n12180;
  assign n12182 = n12177 & ~n12181;
  assign n12183 = ~pi429 & n12180;
  assign n12184 = ~n8026 & ~n12183;
  assign n12185 = pi429 & n12175;
  assign n12186 = n12184 & ~n12185;
  assign n12187 = pi1196 & ~n12186;
  assign n12188 = ~n12182 & n12187;
  assign n12189 = n12160 & ~n12188;
  assign n12190 = ~n12159 & ~n12189;
  assign n12191 = ~pi1199 & n12190;
  assign n12192 = pi428 & ~n12190;
  assign n12193 = ~pi428 & n12158;
  assign n12194 = ~n12192 & ~n12193;
  assign n12195 = ~pi427 & ~n12194;
  assign n12196 = ~pi428 & ~n12190;
  assign n12197 = pi428 & n12158;
  assign n12198 = ~n12196 & ~n12197;
  assign n12199 = pi427 & ~n12198;
  assign n12200 = ~n12195 & ~n12199;
  assign n12201 = pi430 & ~n12200;
  assign n12202 = pi427 & ~n12194;
  assign n12203 = ~pi427 & ~n12198;
  assign n12204 = ~n12202 & ~n12203;
  assign n12205 = ~pi430 & ~n12204;
  assign n12206 = ~n12201 & ~n12205;
  assign n12207 = pi426 & ~n12206;
  assign n12208 = pi430 & ~n12204;
  assign n12209 = ~pi430 & ~n12200;
  assign n12210 = ~n12208 & ~n12209;
  assign n12211 = ~pi426 & ~n12210;
  assign n12212 = ~n12207 & ~n12211;
  assign n12213 = pi445 & ~n12212;
  assign n12214 = pi426 & ~n12210;
  assign n12215 = ~pi426 & ~n12206;
  assign n12216 = ~n12214 & ~n12215;
  assign n12217 = ~pi445 & ~n12216;
  assign n12218 = ~n12213 & ~n12217;
  assign n12219 = ~pi448 & n12218;
  assign n12220 = n8046 & ~n12219;
  assign n12221 = pi445 & ~n12216;
  assign n12222 = ~pi445 & ~n12212;
  assign n12223 = ~n12221 & ~n12222;
  assign n12224 = pi448 & n12223;
  assign n12225 = n12220 & ~n12224;
  assign n12226 = ~pi448 & n12223;
  assign n12227 = pi448 & n12218;
  assign n12228 = ~n12226 & ~n12227;
  assign n12229 = ~n8046 & n12228;
  assign n12230 = ~n12225 & ~n12229;
  assign n12231 = pi1199 & n12230;
  assign n12232 = ~n12191 & ~n12231;
  assign n12233 = n7958 & n12232;
  assign n12234 = n11953 & ~n12233;
  assign n12235 = ~n12039 & ~n12158;
  assign n12236 = n7881 & ~n12117;
  assign n12237 = ~n7849 & n11947;
  assign n12238 = n7849 & n12146;
  assign n12239 = ~n12237 & ~n12238;
  assign n12240 = n12147 & ~n12239;
  assign n12241 = n7849 & n12138;
  assign n12242 = ~n12237 & ~n12241;
  assign n12243 = ~n12066 & n12242;
  assign n12244 = n12140 & ~n12243;
  assign n12245 = ~n12149 & ~n12244;
  assign n12246 = ~n12240 & n12245;
  assign n12247 = ~pi75 & n12246;
  assign n12248 = n12154 & ~n12247;
  assign n12249 = n12118 & ~n12248;
  assign n12250 = n12236 & ~n12249;
  assign n12251 = ~pi1199 & ~n12250;
  assign n12252 = n12043 & n12251;
  assign n12253 = n7874 & n11947;
  assign n12254 = ~n7874 & n12146;
  assign n12255 = ~n12253 & ~n12254;
  assign n12256 = n12148 & ~n12255;
  assign n12257 = ~n7874 & n12138;
  assign n12258 = ~n12253 & ~n12257;
  assign n12259 = n12141 & ~n12258;
  assign n12260 = ~n12149 & ~n12259;
  assign n12261 = ~n12256 & n12260;
  assign n12262 = n12246 & n12261;
  assign n12263 = n12236 & ~n12262;
  assign n12264 = ~n12117 & ~n12261;
  assign n12265 = n8608 & n12264;
  assign n12266 = ~n12263 & ~n12265;
  assign n12267 = ~pi75 & ~n12266;
  assign n12268 = pi567 & n12267;
  assign n12269 = n8295 & n12118;
  assign n12270 = ~n11950 & ~n12269;
  assign n12271 = pi1199 & ~n12270;
  assign n12272 = ~n12268 & n12271;
  assign n12273 = ~n8293 & ~n12272;
  assign n12274 = ~n12252 & n12273;
  assign n12275 = ~pi1197 & n12274;
  assign n12276 = ~n12235 & ~n12275;
  assign n12277 = ~pi333 & ~n12276;
  assign n12278 = n8293 & ~n12158;
  assign n12279 = ~n12274 & ~n12278;
  assign n12280 = pi333 & ~n12279;
  assign n12281 = ~n12277 & ~n12280;
  assign n12282 = ~pi391 & ~n12281;
  assign n12283 = pi333 & ~n12276;
  assign n12284 = ~pi333 & ~n12279;
  assign n12285 = ~n12283 & ~n12284;
  assign n12286 = pi391 & ~n12285;
  assign n12287 = ~n12282 & ~n12286;
  assign n12288 = ~pi392 & ~n12287;
  assign n12289 = ~pi391 & ~n12285;
  assign n12290 = pi391 & ~n12281;
  assign n12291 = ~n12289 & ~n12290;
  assign n12292 = pi392 & ~n12291;
  assign n12293 = ~n12288 & ~n12292;
  assign n12294 = ~pi393 & ~n12293;
  assign n12295 = ~pi392 & ~n12291;
  assign n12296 = pi392 & ~n12287;
  assign n12297 = ~n12295 & ~n12296;
  assign n12298 = pi393 & ~n12297;
  assign n12299 = n7931 & ~n12298;
  assign n12300 = ~n12294 & n12299;
  assign n12301 = pi393 & ~n12293;
  assign n12302 = ~pi393 & ~n12297;
  assign n12303 = ~n7931 & ~n12302;
  assign n12304 = ~n12301 & n12303;
  assign n12305 = pi591 & ~n12304;
  assign n12306 = ~n12300 & n12305;
  assign n12307 = ~pi1197 & ~n11950;
  assign n12308 = ~n7737 & ~n12307;
  assign n12309 = ~n7761 & n11950;
  assign n12310 = ~pi592 & ~n11950;
  assign n12311 = pi592 & n12156;
  assign n12312 = ~n12310 & ~n12311;
  assign n12313 = n7761 & n12312;
  assign n12314 = ~n12309 & ~n12313;
  assign n12315 = pi1197 & n12314;
  assign n12316 = n12308 & ~n12315;
  assign n12317 = n7737 & n12312;
  assign n12318 = ~pi1199 & ~n12317;
  assign n12319 = ~n12316 & n12318;
  assign n12320 = n7788 & n11950;
  assign n12321 = ~n7788 & n12312;
  assign n12322 = ~n12320 & ~n12321;
  assign n12323 = pi1199 & n12322;
  assign n12324 = ~n12319 & ~n12323;
  assign n12325 = ~pi374 & ~n12324;
  assign n12326 = ~pi1198 & ~n12324;
  assign n12327 = pi1198 & ~n12312;
  assign n12328 = ~n12326 & ~n12327;
  assign n12329 = pi374 & ~n12328;
  assign n12330 = ~n12325 & ~n12329;
  assign n12331 = pi369 & ~n7813;
  assign n12332 = ~pi369 & n7813;
  assign n12333 = ~n12331 & ~n12332;
  assign n12334 = n12330 & n12333;
  assign n12335 = ~pi374 & ~n12328;
  assign n12336 = pi374 & ~n12324;
  assign n12337 = ~n12335 & ~n12336;
  assign n12338 = ~n12333 & n12337;
  assign n12339 = ~pi591 & ~n12338;
  assign n12340 = ~n12334 & n12339;
  assign n12341 = ~n12306 & ~n12340;
  assign n12342 = ~pi590 & n12341;
  assign n12343 = n7668 & n11950;
  assign n12344 = ~n7668 & n12158;
  assign n12345 = ~n12343 & ~n12344;
  assign n12346 = pi1198 & ~n12345;
  assign n12347 = ~pi1198 & ~n12042;
  assign n12348 = n7617 & n11950;
  assign n12349 = ~n7617 & n12158;
  assign n12350 = ~n12348 & ~n12349;
  assign n12351 = pi355 & ~n12350;
  assign n12352 = pi455 & ~n11950;
  assign n12353 = ~pi455 & ~n12158;
  assign n12354 = ~n12352 & ~n12353;
  assign n12355 = ~pi452 & ~n12354;
  assign n12356 = ~pi455 & ~n11950;
  assign n12357 = pi455 & ~n12158;
  assign n12358 = ~n12356 & ~n12357;
  assign n12359 = pi452 & ~n12358;
  assign n12360 = ~n12355 & ~n12359;
  assign n12361 = ~pi355 & n12360;
  assign n12362 = ~n12351 & ~n12361;
  assign n12363 = pi458 & n12362;
  assign n12364 = ~pi355 & ~n12350;
  assign n12365 = pi355 & n12360;
  assign n12366 = ~n12364 & ~n12365;
  assign n12367 = ~pi458 & n12366;
  assign n12368 = n7629 & ~n12367;
  assign n12369 = ~n12363 & n12368;
  assign n12370 = ~pi458 & n12362;
  assign n12371 = pi458 & n12366;
  assign n12372 = ~n12370 & ~n12371;
  assign n12373 = ~n7629 & n12372;
  assign n12374 = ~n12369 & ~n12373;
  assign n12375 = pi1196 & n12374;
  assign n12376 = n12347 & ~n12375;
  assign n12377 = ~n12346 & ~n12376;
  assign n12378 = ~n7614 & ~n12377;
  assign n12379 = n7614 & n12158;
  assign n12380 = ~n12378 & ~n12379;
  assign n12381 = ~n7700 & n12380;
  assign n12382 = pi1199 & ~n12158;
  assign n12383 = pi351 & n12382;
  assign n12384 = ~n12381 & ~n12383;
  assign n12385 = ~pi461 & ~n12384;
  assign n12386 = ~n7589 & n12380;
  assign n12387 = ~pi351 & n12382;
  assign n12388 = ~n12386 & ~n12387;
  assign n12389 = pi461 & ~n12388;
  assign n12390 = ~n12385 & ~n12389;
  assign n12391 = n7696 & n12390;
  assign n12392 = ~pi461 & ~n12388;
  assign n12393 = pi461 & ~n12384;
  assign n12394 = ~n12392 & ~n12393;
  assign n12395 = ~n7696 & n12394;
  assign n12396 = ~n12391 & ~n12395;
  assign n12397 = ~pi354 & n12396;
  assign n12398 = ~n7690 & ~n12397;
  assign n12399 = ~pi357 & n12394;
  assign n12400 = ~pi356 & ~n12399;
  assign n12401 = pi357 & n12390;
  assign n12402 = n12400 & ~n12401;
  assign n12403 = ~pi357 & n12390;
  assign n12404 = pi356 & ~n12403;
  assign n12405 = pi357 & n12394;
  assign n12406 = n12404 & ~n12405;
  assign n12407 = ~n12402 & ~n12406;
  assign n12408 = pi354 & ~n12407;
  assign n12409 = n12398 & ~n12408;
  assign n12410 = ~pi354 & ~n12407;
  assign n12411 = pi354 & n12396;
  assign n12412 = ~n12410 & ~n12411;
  assign n12413 = n7690 & n12412;
  assign n12414 = ~pi591 & ~n12413;
  assign n12415 = ~n12409 & n12414;
  assign n12416 = n12001 & ~n12415;
  assign n12417 = ~pi588 & ~n12416;
  assign n12418 = ~n12342 & n12417;
  assign n12419 = ~n12234 & ~n12418;
  assign n12420 = n7376 & n12419;
  assign n12421 = ~n7380 & ~n12076;
  assign n12422 = ~n7415 & n12076;
  assign n12423 = ~pi122 & n12076;
  assign n12424 = n7490 & ~n12423;
  assign n12425 = n2615 & ~n12066;
  assign n12426 = ~n12424 & n12425;
  assign n12427 = n3258 & ~n12066;
  assign n12428 = ~n12138 & n12427;
  assign n12429 = pi87 & n12425;
  assign n12430 = ~n12146 & n12429;
  assign n12431 = ~n12428 & ~n12430;
  assign n12432 = pi122 & ~n12431;
  assign n12433 = ~n12426 & ~n12432;
  assign n12434 = ~pi75 & ~n12433;
  assign n12435 = pi567 & n7380;
  assign n12436 = ~n12434 & n12435;
  assign n12437 = ~n12422 & n12436;
  assign n12438 = ~n12421 & ~n12437;
  assign n12439 = ~n11949 & n12438;
  assign n12440 = pi592 & ~n12439;
  assign n12441 = ~n12310 & ~n12440;
  assign n12442 = n7761 & n12441;
  assign n12443 = ~n12309 & ~n12442;
  assign n12444 = pi1197 & n12443;
  assign n12445 = n12308 & ~n12444;
  assign n12446 = n7737 & n12441;
  assign n12447 = ~pi1199 & ~n12446;
  assign n12448 = ~n12445 & n12447;
  assign n12449 = ~n7788 & n12441;
  assign n12450 = ~n12320 & ~n12449;
  assign n12451 = pi1199 & n12450;
  assign n12452 = ~n12448 & ~n12451;
  assign n12453 = ~pi374 & ~n12452;
  assign n12454 = ~pi1198 & ~n12452;
  assign n12455 = pi1198 & ~n12441;
  assign n12456 = ~n12454 & ~n12455;
  assign n12457 = pi374 & ~n12456;
  assign n12458 = ~n12453 & ~n12457;
  assign n12459 = pi369 & ~n12458;
  assign n12460 = ~pi374 & ~n12456;
  assign n12461 = pi374 & ~n12452;
  assign n12462 = ~n12460 & ~n12461;
  assign n12463 = ~pi369 & ~n12462;
  assign n12464 = n7813 & ~n12463;
  assign n12465 = ~n12459 & n12464;
  assign n12466 = pi369 & ~n12462;
  assign n12467 = ~pi369 & ~n12458;
  assign n12468 = ~n7813 & ~n12467;
  assign n12469 = ~n12466 & n12468;
  assign n12470 = ~pi591 & ~n12469;
  assign n12471 = ~n12465 & n12470;
  assign n12472 = ~pi592 & ~n12439;
  assign n12473 = ~n12041 & ~n12472;
  assign n12474 = ~n12039 & n12473;
  assign n12475 = ~n12069 & ~n12118;
  assign n12476 = pi122 & ~n12239;
  assign n12477 = ~n12063 & ~n12476;
  assign n12478 = n7490 & ~n12477;
  assign n12479 = n12429 & ~n12478;
  assign n12480 = pi122 & ~n12242;
  assign n12481 = ~n12063 & ~n12480;
  assign n12482 = n7490 & ~n12481;
  assign n12483 = n12427 & ~n12482;
  assign n12484 = ~n2615 & n12067;
  assign n12485 = ~n12483 & ~n12484;
  assign n12486 = ~n12479 & n12485;
  assign n12487 = ~pi75 & ~n12486;
  assign n12488 = pi75 & n12067;
  assign n12489 = n12435 & ~n12488;
  assign n12490 = ~n12487 & n12489;
  assign n12491 = ~n12475 & ~n12490;
  assign n12492 = n7881 & ~n12491;
  assign n12493 = ~n12042 & ~n12492;
  assign n12494 = ~pi1199 & ~n12493;
  assign n12495 = ~n12080 & ~n12118;
  assign n12496 = ~n12075 & ~n12139;
  assign n12497 = n2615 & ~n12496;
  assign n12498 = ~n12065 & n12497;
  assign n12499 = n12258 & n12427;
  assign n12500 = n12242 & n12499;
  assign n12501 = ~n12254 & n12429;
  assign n12502 = n12239 & n12501;
  assign n12503 = ~n12500 & ~n12502;
  assign n12504 = ~n12063 & ~n12503;
  assign n12505 = ~pi122 & n12073;
  assign n12506 = n12504 & ~n12505;
  assign n12507 = ~n12498 & ~n12506;
  assign n12508 = ~pi75 & ~n12507;
  assign n12509 = ~n7415 & ~n12077;
  assign n12510 = ~n12065 & n12509;
  assign n12511 = n12435 & ~n12510;
  assign n12512 = ~n12508 & n12511;
  assign n12513 = ~n12495 & ~n12512;
  assign n12514 = n7881 & ~n12513;
  assign n12515 = ~n12079 & ~n12118;
  assign n12516 = n12255 & n12429;
  assign n12517 = ~n12499 & ~n12516;
  assign n12518 = pi122 & ~n12517;
  assign n12519 = ~n12497 & ~n12518;
  assign n12520 = ~pi75 & ~n12519;
  assign n12521 = ~n12509 & ~n12520;
  assign n12522 = n12435 & n12521;
  assign n12523 = ~n12515 & ~n12522;
  assign n12524 = n8608 & ~n12523;
  assign n12525 = ~n12514 & ~n12524;
  assign n12526 = pi1199 & ~n12525;
  assign n12527 = ~n12041 & ~n12526;
  assign n12528 = ~n12494 & n12527;
  assign n12529 = n12039 & n12528;
  assign n12530 = ~n12474 & ~n12529;
  assign n12531 = pi333 & ~n12530;
  assign n12532 = n8293 & ~n12473;
  assign n12533 = ~n8293 & ~n12528;
  assign n12534 = ~n12532 & ~n12533;
  assign n12535 = ~pi333 & n12534;
  assign n12536 = ~n12531 & ~n12535;
  assign n12537 = pi391 & ~n12536;
  assign n12538 = pi333 & ~n12534;
  assign n12539 = ~pi333 & n12530;
  assign n12540 = ~n12538 & ~n12539;
  assign n12541 = ~pi391 & n12540;
  assign n12542 = ~n12537 & ~n12541;
  assign n12543 = pi392 & ~n12542;
  assign n12544 = pi391 & ~n12540;
  assign n12545 = ~pi391 & n12536;
  assign n12546 = ~n12544 & ~n12545;
  assign n12547 = ~pi392 & n12546;
  assign n12548 = ~n12543 & ~n12547;
  assign n12549 = n7934 & ~n12548;
  assign n12550 = pi392 & ~n12546;
  assign n12551 = ~pi392 & n12542;
  assign n12552 = ~n12550 & ~n12551;
  assign n12553 = ~n7934 & n12552;
  assign n12554 = ~n12549 & ~n12553;
  assign n12555 = pi591 & n12554;
  assign n12556 = ~pi590 & ~n12555;
  assign n12557 = ~n12471 & n12556;
  assign n12558 = ~n7668 & n12473;
  assign n12559 = ~n12343 & ~n12558;
  assign n12560 = pi1198 & ~n12559;
  assign n12561 = ~n7617 & n12473;
  assign n12562 = ~n12348 & ~n12561;
  assign n12563 = ~pi355 & ~n12562;
  assign n12564 = ~pi455 & ~n12473;
  assign n12565 = ~n12352 & ~n12564;
  assign n12566 = ~pi452 & ~n12565;
  assign n12567 = pi455 & ~n12473;
  assign n12568 = ~n12356 & ~n12567;
  assign n12569 = pi452 & ~n12568;
  assign n12570 = ~n12566 & ~n12569;
  assign n12571 = pi355 & n12570;
  assign n12572 = ~n12563 & ~n12571;
  assign n12573 = ~pi458 & n12572;
  assign n12574 = n7629 & ~n12573;
  assign n12575 = pi355 & ~n12562;
  assign n12576 = ~pi355 & n12570;
  assign n12577 = ~n12575 & ~n12576;
  assign n12578 = pi458 & n12577;
  assign n12579 = n12574 & ~n12578;
  assign n12580 = ~pi458 & n12577;
  assign n12581 = ~n7629 & ~n12580;
  assign n12582 = pi458 & n12572;
  assign n12583 = n12581 & ~n12582;
  assign n12584 = pi1196 & ~n12583;
  assign n12585 = ~n12579 & n12584;
  assign n12586 = n12347 & ~n12585;
  assign n12587 = ~n12560 & ~n12586;
  assign n12588 = ~n7614 & ~n12587;
  assign n12589 = n7614 & n12473;
  assign n12590 = ~n12588 & ~n12589;
  assign n12591 = ~n7700 & n12590;
  assign n12592 = pi1199 & ~n12473;
  assign n12593 = pi351 & n12592;
  assign n12594 = ~n12591 & ~n12593;
  assign n12595 = ~pi461 & ~n12594;
  assign n12596 = ~n7589 & n12590;
  assign n12597 = ~pi351 & n12592;
  assign n12598 = ~n12596 & ~n12597;
  assign n12599 = pi461 & ~n12598;
  assign n12600 = ~n12595 & ~n12599;
  assign n12601 = n7696 & n12600;
  assign n12602 = ~pi461 & ~n12598;
  assign n12603 = pi461 & ~n12594;
  assign n12604 = ~n12602 & ~n12603;
  assign n12605 = ~n7696 & n12604;
  assign n12606 = ~n12601 & ~n12605;
  assign n12607 = ~pi354 & n12606;
  assign n12608 = ~n7690 & ~n12607;
  assign n12609 = ~pi357 & n12604;
  assign n12610 = ~pi356 & ~n12609;
  assign n12611 = pi357 & n12600;
  assign n12612 = n12610 & ~n12611;
  assign n12613 = ~pi357 & n12600;
  assign n12614 = pi356 & ~n12613;
  assign n12615 = pi357 & n12604;
  assign n12616 = n12614 & ~n12615;
  assign n12617 = ~n12612 & ~n12616;
  assign n12618 = pi354 & ~n12617;
  assign n12619 = n12608 & ~n12618;
  assign n12620 = ~pi354 & ~n12617;
  assign n12621 = pi354 & n12606;
  assign n12622 = ~n12620 & ~n12621;
  assign n12623 = n7690 & n12622;
  assign n12624 = ~pi591 & ~n12623;
  assign n12625 = ~n12619 & n12624;
  assign n12626 = n12001 & ~n12625;
  assign n12627 = ~pi588 & ~n12626;
  assign n12628 = ~n12557 & n12627;
  assign n12629 = ~n8011 & n12473;
  assign n12630 = ~pi443 & ~n12473;
  assign n12631 = ~n12161 & ~n12630;
  assign n12632 = ~n8162 & n12631;
  assign n12633 = pi443 & ~n12473;
  assign n12634 = ~n12165 & ~n12633;
  assign n12635 = n8162 & n12634;
  assign n12636 = ~n12632 & ~n12635;
  assign n12637 = pi435 & ~n12636;
  assign n12638 = n8162 & n12631;
  assign n12639 = ~n8162 & n12634;
  assign n12640 = ~n12638 & ~n12639;
  assign n12641 = ~pi435 & ~n12640;
  assign n12642 = ~n12637 & ~n12641;
  assign n12643 = ~pi429 & n12642;
  assign n12644 = n8026 & ~n12643;
  assign n12645 = ~pi435 & ~n12636;
  assign n12646 = pi435 & ~n12640;
  assign n12647 = ~n12645 & ~n12646;
  assign n12648 = pi429 & n12647;
  assign n12649 = n12644 & ~n12648;
  assign n12650 = ~pi429 & n12647;
  assign n12651 = ~n8026 & ~n12650;
  assign n12652 = pi429 & n12642;
  assign n12653 = n12651 & ~n12652;
  assign n12654 = pi1196 & ~n12653;
  assign n12655 = ~n12649 & n12654;
  assign n12656 = n12160 & ~n12655;
  assign n12657 = ~n12629 & ~n12656;
  assign n12658 = ~pi1199 & n12657;
  assign n12659 = pi428 & ~n12657;
  assign n12660 = ~pi428 & n12473;
  assign n12661 = ~n12659 & ~n12660;
  assign n12662 = pi427 & ~n12661;
  assign n12663 = ~pi428 & ~n12657;
  assign n12664 = pi428 & n12473;
  assign n12665 = ~n12663 & ~n12664;
  assign n12666 = ~pi427 & ~n12665;
  assign n12667 = ~n12662 & ~n12666;
  assign n12668 = pi430 & ~n12667;
  assign n12669 = ~pi427 & ~n12661;
  assign n12670 = pi427 & ~n12665;
  assign n12671 = ~n12669 & ~n12670;
  assign n12672 = ~pi430 & ~n12671;
  assign n12673 = ~n12668 & ~n12672;
  assign n12674 = pi426 & ~n12673;
  assign n12675 = pi430 & ~n12671;
  assign n12676 = ~pi430 & ~n12667;
  assign n12677 = ~n12675 & ~n12676;
  assign n12678 = ~pi426 & ~n12677;
  assign n12679 = ~n12674 & ~n12678;
  assign n12680 = pi445 & ~n12679;
  assign n12681 = pi426 & ~n12677;
  assign n12682 = ~pi426 & ~n12673;
  assign n12683 = ~n12681 & ~n12682;
  assign n12684 = ~pi445 & ~n12683;
  assign n12685 = ~n12680 & ~n12684;
  assign n12686 = pi448 & n12685;
  assign n12687 = pi445 & ~n12683;
  assign n12688 = ~pi445 & ~n12679;
  assign n12689 = ~n12687 & ~n12688;
  assign n12690 = ~pi448 & n12689;
  assign n12691 = n8046 & ~n12690;
  assign n12692 = ~n12686 & n12691;
  assign n12693 = ~pi448 & n12685;
  assign n12694 = pi448 & n12689;
  assign n12695 = ~n8046 & ~n12694;
  assign n12696 = ~n12693 & n12695;
  assign n12697 = ~n12692 & ~n12696;
  assign n12698 = pi1199 & n12697;
  assign n12699 = ~n12658 & ~n12698;
  assign n12700 = n7958 & n12699;
  assign n12701 = n11953 & ~n12700;
  assign n12702 = ~n7376 & ~n12701;
  assign n12703 = ~n12628 & n12702;
  assign n12704 = ~po1038 & ~n12703;
  assign n12705 = ~pi80 & n12704;
  assign n12706 = ~n12420 & n12705;
  assign n12707 = ~pi217 & ~n12706;
  assign n12708 = ~n12116 & n12707;
  assign n12709 = ~pi80 & ~n11950;
  assign n12710 = pi217 & ~n12709;
  assign n12711 = n7588 & ~n12710;
  assign po238 = ~n12708 & n12711;
  assign n12713 = ~po1038 & n11086;
  assign n12714 = ~pi314 & n11157;
  assign n12715 = pi68 & ~pi81;
  assign n12716 = n2473 & n12715;
  assign n12717 = n2791 & n12716;
  assign n12718 = n10803 & n12717;
  assign n12719 = n11230 & n12718;
  assign n12720 = ~n12714 & ~n12719;
  assign po239 = n12713 & ~n12720;
  assign n12722 = pi69 & pi314;
  assign n12723 = n2783 & n12722;
  assign n12724 = pi66 & ~pi73;
  assign n12725 = n2469 & n12724;
  assign n12726 = n2483 & n12725;
  assign n12727 = ~n12723 & ~n12726;
  assign n12728 = n10896 & n10900;
  assign po240 = ~n12727 & n12728;
  assign n12730 = n8781 & n10895;
  assign n12731 = pi84 & n9046;
  assign n12732 = n2473 & n2790;
  assign n12733 = n2468 & n12732;
  assign n12734 = n12731 & n12733;
  assign n12735 = n2485 & n11172;
  assign n12736 = ~n12734 & ~n12735;
  assign n12737 = n12730 & ~n12736;
  assign n12738 = ~pi314 & ~n12737;
  assign n12739 = n12730 & n12734;
  assign n12740 = pi314 & ~n12739;
  assign n12741 = n9988 & ~n12740;
  assign po241 = ~n12738 & n12741;
  assign n12743 = pi211 & pi299;
  assign n12744 = pi219 & pi299;
  assign n12745 = ~n10615 & ~n12744;
  assign n12746 = ~n12743 & n12745;
  assign n12747 = ~po1038 & n12746;
  assign po242 = n11160 & n12747;
  assign n12749 = n6318 & n10897;
  assign n12750 = ~pi314 & n10898;
  assign n12751 = n11228 & n12750;
  assign n12752 = ~n12749 & ~n12751;
  assign po243 = n10900 & ~n12752;
  assign n12754 = n7468 & n11179;
  assign n12755 = n7464 & n11182;
  assign n12756 = ~n12754 & ~n12755;
  assign po244 = n10780 & ~n12756;
  assign n12758 = n2689 & n10895;
  assign n12759 = n2836 & n12758;
  assign n12760 = pi314 & n9988;
  assign n12761 = n2694 & n12760;
  assign po245 = n12759 & n12761;
  assign n12763 = n7368 & n10826;
  assign n12764 = ~pi1093 & ~n12763;
  assign n12765 = n12121 & n12124;
  assign n12766 = n10823 & n12765;
  assign n12767 = n2711 & n12766;
  assign n12768 = n10839 & n12767;
  assign n12769 = pi1093 & ~n12768;
  assign n12770 = ~n12764 & ~n12769;
  assign n12771 = ~n6211 & n12770;
  assign n12772 = n2576 & n12771;
  assign n12773 = n7376 & ~n12772;
  assign n12774 = n2698 & n7368;
  assign n12775 = n2575 & n10017;
  assign n12776 = ~pi1093 & n12775;
  assign n12777 = n12774 & n12776;
  assign n12778 = n11245 & n12777;
  assign n12779 = ~n7376 & ~n12778;
  assign n12780 = ~po1038 & ~n12779;
  assign po246 = ~n12773 & n12780;
  assign n12782 = pi70 & ~n8815;
  assign n12783 = n10005 & n11138;
  assign n12784 = pi841 & n12783;
  assign n12785 = n7394 & n12784;
  assign n12786 = ~pi70 & ~n12785;
  assign n12787 = n9986 & ~n12786;
  assign n12788 = n12142 & n12787;
  assign po247 = ~n12782 & n12788;
  assign n12790 = ~pi1050 & n9412;
  assign n12791 = ~pi90 & ~n12790;
  assign n12792 = n2889 & ~n12791;
  assign n12793 = ~n7383 & n12792;
  assign po248 = n11110 & n12793;
  assign n12795 = pi24 & ~n2978;
  assign n12796 = n2941 & n12795;
  assign n12797 = n2749 & n12796;
  assign n12798 = n10879 & n12797;
  assign n12799 = ~n6354 & ~n9982;
  assign n12800 = n2978 & ~n12799;
  assign n12801 = n9987 & n12800;
  assign n12802 = ~pi39 & ~n12801;
  assign n12803 = ~n12798 & n12802;
  assign n12804 = n10024 & ~n12803;
  assign po249 = ~n7472 & n12804;
  assign n12806 = n2534 & ~po1038;
  assign n12807 = pi92 & n2522;
  assign n12808 = n3345 & n11263;
  assign n12809 = n12807 & n12808;
  assign n12810 = pi224 & n7465;
  assign n12811 = n7464 & n12810;
  assign n12812 = pi299 & n8959;
  assign n12813 = n7468 & n12812;
  assign n12814 = ~n12811 & ~n12813;
  assign n12815 = n10912 & ~n12814;
  assign n12816 = n2536 & n12815;
  assign n12817 = ~n12809 & ~n12816;
  assign po250 = n12806 & ~n12817;
  assign n12819 = ~pi1050 & n2522;
  assign n12820 = pi92 & ~n12819;
  assign n12821 = n3345 & n12806;
  assign n12822 = pi93 & n10879;
  assign n12823 = n2915 & n12822;
  assign n12824 = ~pi92 & ~n12823;
  assign n12825 = n12821 & ~n12824;
  assign po251 = ~n12820 & n12825;
  assign n12827 = n10083 & n10857;
  assign n12828 = ~n2771 & ~n12827;
  assign n12829 = n2712 & n9987;
  assign n12830 = ~n12828 & n12829;
  assign n12831 = pi252 & n12830;
  assign n12832 = n10860 & n11071;
  assign n12833 = n2914 & n12832;
  assign n12834 = pi1093 & ~n12833;
  assign n12835 = n7447 & ~n12834;
  assign n12836 = ~pi252 & n12832;
  assign n12837 = ~n12835 & ~n12836;
  assign n12838 = ~n12831 & n12837;
  assign n12839 = n8744 & n12838;
  assign n12840 = n8744 & ~po840;
  assign n12841 = ~n12832 & ~n12840;
  assign n12842 = n9986 & ~n12841;
  assign po252 = ~n12839 & n12842;
  assign n12844 = ~pi332 & n9987;
  assign n12845 = n11070 & n12844;
  assign n12846 = n12783 & n12845;
  assign n12847 = n2686 & n11811;
  assign n12848 = n10015 & n12847;
  assign n12849 = ~pi39 & ~n12848;
  assign n12850 = ~n12846 & n12849;
  assign n12851 = n2607 & n5792;
  assign n12852 = n6191 & ~n6456;
  assign n12853 = ~n9380 & ~n12852;
  assign n12854 = ~n11204 & ~n12853;
  assign n12855 = n12851 & n12854;
  assign n12856 = ~n6456 & ~n11208;
  assign n12857 = n11210 & n12856;
  assign n12858 = pi39 & ~n12857;
  assign n12859 = ~n12855 & n12858;
  assign n12860 = n10024 & ~n12859;
  assign po253 = ~n12850 & n12860;
  assign n12862 = n10263 & n12847;
  assign n12863 = ~pi72 & n2899;
  assign n12864 = n2461 & n12863;
  assign n12865 = pi479 & ~po840;
  assign n12866 = n12864 & n12865;
  assign n12867 = pi96 & ~n12865;
  assign n12868 = n2461 & n12867;
  assign n12869 = n2900 & n2916;
  assign n12870 = n2507 & n12869;
  assign n12871 = n12868 & n12870;
  assign n12872 = ~n12866 & ~n12871;
  assign n12873 = ~pi95 & ~n12872;
  assign n12874 = ~n12862 & ~n12873;
  assign po254 = n9986 & ~n12874;
  assign n12876 = pi39 & ~n11212;
  assign n12877 = pi593 & n12876;
  assign n12878 = ~n6456 & n12877;
  assign n12879 = n6166 & n12865;
  assign n12880 = ~po740 & ~n12879;
  assign n12881 = n2515 & n10016;
  assign n12882 = ~n12880 & n12881;
  assign n12883 = n11275 & n12882;
  assign n12884 = ~n12878 & ~n12883;
  assign po255 = n10024 & ~n12884;
  assign n12886 = ~pi92 & n11264;
  assign n12887 = ~n12807 & ~n12886;
  assign n12888 = pi314 & ~n12887;
  assign n12889 = pi1050 & n12888;
  assign po256 = n12821 & n12889;
  assign n12891 = ~pi72 & pi152;
  assign n12892 = n10119 & n12891;
  assign n12893 = pi299 & n12892;
  assign n12894 = ~pi72 & n10123;
  assign n12895 = n10125 & n12894;
  assign n12896 = ~n12893 & ~n12895;
  assign n12897 = pi232 & ~n12896;
  assign n12898 = pi39 & ~n12897;
  assign n12899 = ~pi72 & pi99;
  assign n12900 = ~pi39 & ~n12899;
  assign n12901 = ~n12898 & ~n12900;
  assign n12902 = ~n7380 & ~n12901;
  assign n12903 = ~po1038 & ~n12902;
  assign n12904 = ~n7484 & ~n12899;
  assign n12905 = ~n2914 & n12899;
  assign n12906 = n7484 & ~n12905;
  assign n12907 = ~n10154 & n12899;
  assign n12908 = n6108 & n10140;
  assign n12909 = ~n12907 & ~n12908;
  assign n12910 = n10145 & ~n12909;
  assign n12911 = n12906 & ~n12910;
  assign n12912 = ~n12904 & ~n12911;
  assign n12913 = ~pi39 & ~n12912;
  assign n12914 = ~n12898 & ~n12913;
  assign n12915 = n6098 & ~n12914;
  assign n12916 = pi38 & ~n12901;
  assign n12917 = pi39 & ~n10731;
  assign n12918 = n12897 & n12917;
  assign n12919 = pi41 & pi72;
  assign n12920 = pi99 & ~n12919;
  assign n12921 = ~n10199 & n12920;
  assign n12922 = n10558 & ~n12921;
  assign n12923 = ~n10234 & n12920;
  assign n12924 = n10561 & ~n12923;
  assign n12925 = ~n10213 & n12920;
  assign n12926 = n10559 & ~n12925;
  assign n12927 = ~n12924 & ~n12926;
  assign n12928 = pi228 & ~n12927;
  assign n12929 = ~pi39 & ~n12928;
  assign n12930 = ~n12922 & n12929;
  assign n12931 = ~n12918 & ~n12930;
  assign n12932 = n2614 & n12931;
  assign n12933 = ~pi87 & ~n12932;
  assign n12934 = ~n12916 & n12933;
  assign n12935 = ~n12915 & n12934;
  assign n12936 = ~pi75 & ~n12935;
  assign n12937 = pi228 & n10311;
  assign n12938 = pi228 & n10151;
  assign n12939 = n12899 & ~n12938;
  assign n12940 = ~n12937 & ~n12939;
  assign n12941 = n2615 & n12940;
  assign n12942 = ~n2533 & ~n12901;
  assign n12943 = pi87 & ~n12942;
  assign n12944 = ~n12941 & n12943;
  assign n12945 = n12936 & ~n12944;
  assign n12946 = ~n2572 & n12901;
  assign n12947 = pi75 & ~n12946;
  assign n12948 = ~n10267 & n12899;
  assign n12949 = n6109 & n10720;
  assign n12950 = ~n12948 & ~n12949;
  assign n12951 = n10145 & ~n12950;
  assign n12952 = n12906 & ~n12951;
  assign n12953 = ~n12904 & ~n12952;
  assign n12954 = ~pi39 & ~n12953;
  assign n12955 = ~n12898 & ~n12954;
  assign n12956 = n2572 & n12955;
  assign n12957 = n12947 & ~n12956;
  assign n12958 = ~n12945 & ~n12957;
  assign n12959 = n7380 & ~n12958;
  assign n12960 = n12903 & ~n12959;
  assign n12961 = pi232 & n12892;
  assign n12962 = pi39 & ~n12961;
  assign n12963 = po1038 & ~n12900;
  assign n12964 = ~n12962 & n12963;
  assign po257 = n12960 | n12964;
  assign n12966 = ~pi75 & n3257;
  assign n12967 = pi129 & ~n9906;
  assign n12968 = ~n6105 & ~n12967;
  assign n12969 = ~n7420 & n9906;
  assign n12970 = pi129 & ~n12969;
  assign n12971 = n6102 & ~n12970;
  assign n12972 = ~n6127 & ~n12971;
  assign n12973 = ~n12968 & n12972;
  assign n12974 = n12966 & ~n12973;
  assign n12975 = n6098 & n12974;
  assign n12976 = ~pi24 & n8823;
  assign n12977 = po840 & n12976;
  assign n12978 = ~n12975 & ~n12977;
  assign n12979 = n2522 & ~n12978;
  assign po258 = n8739 & n12979;
  assign n12981 = ~pi39 & ~n10147;
  assign n12982 = n3395 & n6190;
  assign n12983 = n12891 & n12982;
  assign n12984 = pi299 & ~n12983;
  assign n12985 = ~pi144 & pi174;
  assign n12986 = ~pi72 & n12985;
  assign n12987 = n10122 & n12986;
  assign n12988 = ~pi299 & ~n12987;
  assign n12989 = ~n12984 & ~n12988;
  assign n12990 = pi232 & n12989;
  assign n12991 = pi39 & ~n12990;
  assign n12992 = ~n12981 & ~n12991;
  assign n12993 = ~n7380 & ~n12992;
  assign n12994 = ~po1038 & ~n12993;
  assign n12995 = ~n2572 & n12992;
  assign n12996 = pi75 & ~n12995;
  assign n12997 = ~n7484 & ~n10147;
  assign n12998 = ~n2914 & n10147;
  assign n12999 = n7484 & ~n12998;
  assign n13000 = n2914 & ~n6116;
  assign n13001 = n10147 & ~n10266;
  assign n13002 = ~n10260 & ~n13001;
  assign n13003 = n13000 & ~n13002;
  assign n13004 = n12999 & ~n13003;
  assign n13005 = ~n12997 & ~n13004;
  assign n13006 = ~pi39 & ~n13005;
  assign n13007 = ~n12991 & ~n13006;
  assign n13008 = n2572 & n13007;
  assign n13009 = n12996 & ~n13008;
  assign n13010 = n7480 & n10150;
  assign n13011 = n10147 & ~n13010;
  assign n13012 = ~n10140 & ~n13011;
  assign n13013 = n13000 & ~n13012;
  assign n13014 = n12999 & ~n13013;
  assign n13015 = ~n12997 & ~n13014;
  assign n13016 = ~pi39 & ~n13015;
  assign n13017 = ~n12991 & ~n13016;
  assign n13018 = n6098 & ~n13017;
  assign n13019 = pi38 & ~n12992;
  assign n13020 = ~n10731 & n12989;
  assign n13021 = ~pi72 & n10280;
  assign n13022 = n13020 & n13021;
  assign n13023 = n10147 & ~n10230;
  assign n13024 = n2914 & ~n10231;
  assign n13025 = ~n13023 & n13024;
  assign n13026 = pi101 & ~n10211;
  assign n13027 = ~n2914 & ~n10208;
  assign n13028 = ~n13026 & n13027;
  assign n13029 = ~n13025 & ~n13028;
  assign n13030 = pi228 & ~n13029;
  assign n13031 = pi101 & ~n10197;
  assign n13032 = ~pi228 & ~n13031;
  assign n13033 = ~n10190 & n13032;
  assign n13034 = ~pi39 & ~n13033;
  assign n13035 = ~n13030 & n13034;
  assign n13036 = ~n13022 & ~n13035;
  assign n13037 = n2614 & n13036;
  assign n13038 = ~pi87 & ~n13037;
  assign n13039 = ~n13019 & n13038;
  assign n13040 = ~n13018 & n13039;
  assign n13041 = ~pi75 & ~n13040;
  assign n13042 = n10150 & n10761;
  assign n13043 = n10147 & ~n13042;
  assign n13044 = ~pi101 & n10762;
  assign n13045 = ~pi39 & ~n13044;
  assign n13046 = ~n13043 & n13045;
  assign n13047 = ~n12991 & ~n13046;
  assign n13048 = pi87 & n13047;
  assign n13049 = n13041 & ~n13048;
  assign n13050 = ~n13009 & ~n13049;
  assign n13051 = n7380 & ~n13050;
  assign n13052 = n12994 & ~n13051;
  assign n13053 = pi232 & n12983;
  assign n13054 = pi39 & ~n13053;
  assign n13055 = po1038 & ~n12981;
  assign n13056 = ~n13054 & n13055;
  assign po259 = n13052 | n13056;
  assign n13058 = n2846 & n8773;
  assign po260 = n12713 & n13058;
  assign n13060 = ~pi109 & ~n12759;
  assign n13061 = n6308 & ~n13060;
  assign n13062 = ~pi314 & ~n13061;
  assign n13063 = pi109 & n2758;
  assign n13064 = n2690 & n13063;
  assign n13065 = pi314 & ~n13064;
  assign n13066 = n10899 & ~n13065;
  assign po261 = ~n13062 & n13066;
  assign n13068 = n7376 & ~n8744;
  assign n13069 = n9903 & ~n13068;
  assign n13070 = n10185 & ~n13069;
  assign n13071 = n8744 & ~n12768;
  assign n13072 = ~n10175 & ~n12767;
  assign n13073 = n10839 & ~n13072;
  assign n13074 = ~n8744 & ~n13073;
  assign n13075 = ~n7376 & ~n13074;
  assign n13076 = ~n6211 & n13075;
  assign n13077 = ~n13071 & n13076;
  assign n13078 = ~n13070 & ~n13077;
  assign po262 = n9986 & ~n13078;
  assign n13080 = pi24 & n11069;
  assign n13081 = ~pi53 & ~n11068;
  assign n13082 = n2709 & ~n13081;
  assign n13083 = ~pi24 & n2712;
  assign n13084 = n13082 & n13083;
  assign n13085 = ~n13080 & ~n13084;
  assign n13086 = pi841 & ~n13085;
  assign n13087 = n8801 & n11049;
  assign n13088 = ~n13086 & ~n13087;
  assign po264 = n9988 & ~n13088;
  assign n13090 = ~pi999 & n9988;
  assign po265 = n11139 & n13090;
  assign n13092 = ~pi97 & n7391;
  assign n13093 = ~pi108 & ~n13092;
  assign n13094 = n2768 & ~n13093;
  assign n13095 = n2694 & n13094;
  assign n13096 = n7395 & n10063;
  assign n13097 = n13095 & n13096;
  assign n13098 = pi314 & ~n7393;
  assign n13099 = n7395 & ~n13098;
  assign n13100 = ~pi314 & ~n13095;
  assign n13101 = ~n10063 & ~n13100;
  assign n13102 = n13099 & n13101;
  assign n13103 = ~pi51 & ~n13102;
  assign n13104 = ~n13097 & n13103;
  assign n13105 = n2533 & ~n13104;
  assign n13106 = n7398 & n13105;
  assign n13107 = ~pi87 & ~n13106;
  assign n13108 = n6096 & n8739;
  assign po266 = ~n13107 & n13108;
  assign n13110 = n2775 & n11234;
  assign po267 = n12760 & n13110;
  assign n13112 = ~pi82 & n8781;
  assign n13113 = n2792 & n10898;
  assign n13114 = pi111 & n13113;
  assign n13115 = n13112 & n13114;
  assign n13116 = pi314 & n13115;
  assign n13117 = n8744 & n9903;
  assign n13118 = n10175 & n13117;
  assign n13119 = ~n13116 & ~n13118;
  assign po268 = n9988 & ~n13119;
  assign n13121 = pi72 & n10263;
  assign n13122 = ~pi314 & n13115;
  assign n13123 = n9078 & n13122;
  assign n13124 = ~n13121 & ~n13123;
  assign n13125 = n3084 & n9986;
  assign po269 = ~n13124 & n13125;
  assign po270 = ~pi124 | pi468;
  assign n13128 = pi113 & n10378;
  assign n13129 = ~pi228 & ~n10383;
  assign n13130 = ~n13128 & n13129;
  assign n13131 = ~pi113 & n10562;
  assign n13132 = pi228 & ~n13131;
  assign n13133 = n6108 & n10237;
  assign n13134 = ~n10376 & ~n13133;
  assign n13135 = pi113 & n13134;
  assign n13136 = n13132 & ~n13135;
  assign n13137 = ~pi39 & ~n13136;
  assign n13138 = ~n13130 & n13137;
  assign n13139 = n2614 & ~n13138;
  assign n13140 = ~pi39 & n10379;
  assign n13141 = pi38 & ~n13140;
  assign n13142 = n2914 & n7484;
  assign n13143 = n7480 & n10335;
  assign n13144 = ~n6115 & ~n13143;
  assign n13145 = n13142 & ~n13144;
  assign n13146 = n10379 & ~n13145;
  assign n13147 = ~n6115 & n13142;
  assign n13148 = n10140 & n13147;
  assign n13149 = n10349 & n13148;
  assign n13150 = ~n13146 & ~n13149;
  assign n13151 = ~pi39 & ~n13150;
  assign n13152 = n6098 & ~n13151;
  assign n13153 = ~n13141 & ~n13152;
  assign n13154 = ~n13139 & n13153;
  assign n13155 = ~pi87 & ~n13154;
  assign n13156 = pi228 & n10335;
  assign n13157 = n10379 & ~n13156;
  assign n13158 = ~pi113 & n12937;
  assign n13159 = ~n13157 & ~n13158;
  assign n13160 = n2533 & ~n13159;
  assign n13161 = ~n2614 & n13140;
  assign n13162 = pi87 & ~n13161;
  assign n13163 = ~n13160 & n13162;
  assign n13164 = ~n13155 & ~n13163;
  assign n13165 = ~pi75 & ~n13164;
  assign n13166 = n7423 & n13149;
  assign n13167 = ~n6115 & ~n10318;
  assign n13168 = n13142 & ~n13167;
  assign n13169 = n10379 & ~n13168;
  assign n13170 = ~n13166 & ~n13169;
  assign n13171 = n3258 & ~n13170;
  assign n13172 = ~n2572 & n13140;
  assign n13173 = pi75 & ~n13172;
  assign n13174 = ~n13171 & n13173;
  assign n13175 = ~n13165 & ~n13174;
  assign n13176 = n8739 & ~n13175;
  assign n13177 = ~n8739 & ~n13140;
  assign po271 = ~n13176 & ~n13177;
  assign n13179 = ~pi72 & pi114;
  assign n13180 = ~n10906 & ~n13179;
  assign n13181 = pi114 & ~n10338;
  assign n13182 = ~n10333 & ~n13181;
  assign n13183 = n10906 & n13182;
  assign n13184 = ~pi39 & ~n13183;
  assign n13185 = ~n13180 & n13184;
  assign n13186 = n6098 & ~n13185;
  assign n13187 = ~pi39 & n13179;
  assign n13188 = pi38 & ~n13187;
  assign n13189 = pi114 & n10582;
  assign n13190 = ~pi114 & n10565;
  assign n13191 = ~pi115 & ~n13190;
  assign n13192 = ~n13189 & n13191;
  assign n13193 = pi115 & ~n13179;
  assign n13194 = ~pi39 & ~n13193;
  assign n13195 = ~n13192 & n13194;
  assign n13196 = n2614 & ~n13195;
  assign n13197 = ~pi87 & ~n13196;
  assign n13198 = ~n13188 & n13197;
  assign n13199 = ~n13186 & n13198;
  assign n13200 = ~pi75 & ~n13199;
  assign n13201 = ~n2614 & ~n13187;
  assign n13202 = n10913 & ~n13201;
  assign n13203 = ~n10413 & n13179;
  assign n13204 = ~pi115 & n10417;
  assign n13205 = ~pi114 & n13204;
  assign n13206 = ~n13203 & ~n13205;
  assign n13207 = n2614 & n13206;
  assign n13208 = n13202 & ~n13207;
  assign n13209 = n13200 & ~n13208;
  assign n13210 = ~n2572 & n13187;
  assign n13211 = pi75 & ~n13210;
  assign n13212 = pi114 & n10598;
  assign n13213 = ~n10316 & ~n13212;
  assign n13214 = n10906 & n13213;
  assign n13215 = ~n13180 & ~n13214;
  assign n13216 = n3258 & n13215;
  assign n13217 = n13211 & ~n13216;
  assign n13218 = ~n13209 & ~n13217;
  assign n13219 = n8739 & ~n13218;
  assign n13220 = ~n8739 & ~n13187;
  assign po272 = ~n13219 & ~n13220;
  assign n13222 = ~pi72 & pi115;
  assign n13223 = ~n13142 & ~n13222;
  assign n13224 = pi115 & ~n10338;
  assign n13225 = ~pi115 & n10313;
  assign n13226 = ~pi52 & n10905;
  assign n13227 = n13225 & ~n13226;
  assign n13228 = ~n13224 & ~n13227;
  assign n13229 = n13142 & n13228;
  assign n13230 = ~pi39 & ~n13229;
  assign n13231 = ~n13223 & n13230;
  assign n13232 = n6098 & ~n13231;
  assign n13233 = ~pi39 & n13222;
  assign n13234 = pi38 & ~n13233;
  assign n13235 = pi115 & ~n10582;
  assign n13236 = ~pi115 & ~n10565;
  assign n13237 = ~pi39 & ~n13236;
  assign n13238 = ~n13235 & n13237;
  assign n13239 = n2614 & ~n13238;
  assign n13240 = ~pi87 & ~n13239;
  assign n13241 = ~n13234 & n13240;
  assign n13242 = ~n13232 & n13241;
  assign n13243 = ~pi75 & ~n13242;
  assign n13244 = ~n10412 & n13222;
  assign n13245 = ~n13204 & ~n13244;
  assign n13246 = n2614 & n13245;
  assign n13247 = ~n2614 & ~n13233;
  assign n13248 = n10913 & ~n13247;
  assign n13249 = ~n13246 & n13248;
  assign n13250 = n13243 & ~n13249;
  assign n13251 = ~n2572 & n13233;
  assign n13252 = pi75 & ~n13251;
  assign n13253 = n7423 & n13227;
  assign n13254 = pi115 & n10598;
  assign n13255 = ~n13253 & ~n13254;
  assign n13256 = n13142 & n13255;
  assign n13257 = ~n13223 & ~n13256;
  assign n13258 = n3258 & n13257;
  assign n13259 = n13252 & ~n13258;
  assign n13260 = ~n13250 & ~n13259;
  assign n13261 = n8739 & ~n13260;
  assign n13262 = ~n8739 & ~n13233;
  assign po273 = ~n13261 & ~n13262;
  assign n13264 = ~pi39 & n10361;
  assign n13265 = pi38 & ~n13264;
  assign n13266 = pi116 & ~n10380;
  assign n13267 = ~pi228 & ~n13266;
  assign n13268 = ~n10384 & n13267;
  assign n13269 = pi228 & n10577;
  assign n13270 = ~pi39 & ~n13269;
  assign n13271 = ~n13268 & n13270;
  assign n13272 = n2614 & ~n13271;
  assign n13273 = ~pi87 & ~n13272;
  assign n13274 = n10361 & ~n13142;
  assign n13275 = ~pi113 & n13143;
  assign n13276 = n10361 & ~n13275;
  assign n13277 = ~n10313 & ~n13276;
  assign n13278 = n13147 & ~n13277;
  assign n13279 = ~n13274 & ~n13278;
  assign n13280 = ~pi39 & ~n13279;
  assign n13281 = n6098 & ~n13280;
  assign n13282 = n13273 & ~n13281;
  assign n13283 = ~n13265 & n13282;
  assign n13284 = ~pi75 & ~n13283;
  assign n13285 = ~pi113 & n13156;
  assign n13286 = n10361 & ~n13285;
  assign n13287 = ~pi38 & ~n13286;
  assign n13288 = ~n10417 & n13287;
  assign n13289 = ~pi100 & n13288;
  assign n13290 = ~n2614 & ~n13264;
  assign n13291 = n10913 & ~n13290;
  assign n13292 = ~n13289 & n13291;
  assign n13293 = n13284 & ~n13292;
  assign n13294 = ~n10319 & n10361;
  assign n13295 = ~n10314 & ~n13294;
  assign n13296 = n13147 & ~n13295;
  assign n13297 = ~n13274 & ~n13296;
  assign n13298 = n3258 & ~n13297;
  assign n13299 = ~n2572 & n13264;
  assign n13300 = pi75 & ~n13299;
  assign n13301 = ~n13298 & n13300;
  assign n13302 = ~n13293 & ~n13301;
  assign n13303 = n8739 & ~n13302;
  assign n13304 = ~n8739 & ~n13264;
  assign po274 = ~n13303 & ~n13304;
  assign n13306 = n3657 & n7328;
  assign n13307 = ~n3656 & ~n13306;
  assign n13308 = ~pi38 & ~n13307;
  assign n13309 = ~pi87 & ~n13308;
  assign n13310 = n6096 & ~n13309;
  assign n13311 = ~pi92 & ~n13310;
  assign n13312 = ~n7258 & ~n13311;
  assign n13313 = n2534 & n13312;
  assign n13314 = ~pi55 & ~n13313;
  assign n13315 = ~n7250 & ~n13314;
  assign n13316 = ~pi56 & ~n13315;
  assign n13317 = ~n6264 & ~n13316;
  assign n13318 = ~pi62 & ~n13317;
  assign n13319 = ~pi57 & n6269;
  assign po275 = ~n13318 & n13319;
  assign n13321 = ~pi79 & n11458;
  assign n13322 = pi163 & n6190;
  assign n13323 = ~n11462 & ~n13322;
  assign n13324 = ~pi150 & ~n13323;
  assign n13325 = pi150 & n9542;
  assign n13326 = n11460 & n13325;
  assign n13327 = ~n13324 & ~n13326;
  assign n13328 = n9546 & ~n13327;
  assign n13329 = pi74 & ~n13328;
  assign n13330 = pi165 & n7420;
  assign n13331 = n7255 & ~n13330;
  assign n13332 = ~n13328 & ~n13331;
  assign n13333 = ~n3327 & ~n13332;
  assign n13334 = ~n13329 & n13333;
  assign n13335 = ~pi74 & ~n13328;
  assign n13336 = ~pi38 & ~pi54;
  assign n13337 = ~n13330 & ~n13336;
  assign n13338 = n7255 & n13337;
  assign n13339 = n13335 & ~n13338;
  assign n13340 = ~n13329 & ~n13339;
  assign n13341 = ~n2531 & ~n13340;
  assign n13342 = n3327 & ~n13341;
  assign n13343 = pi299 & n13327;
  assign n13344 = ~pi184 & ~n11515;
  assign n13345 = ~pi185 & n13344;
  assign n13346 = pi185 & ~n13344;
  assign n13347 = n6190 & ~n13346;
  assign n13348 = ~n13345 & n13347;
  assign n13349 = ~pi299 & ~n13348;
  assign n13350 = pi232 & ~n13349;
  assign n13351 = ~n13343 & n13350;
  assign n13352 = ~n7255 & n13351;
  assign n13353 = pi74 & ~n13352;
  assign n13354 = ~pi55 & ~n13353;
  assign n13355 = ~pi143 & ~pi299;
  assign n13356 = ~n8924 & ~n13330;
  assign n13357 = ~n13355 & ~n13356;
  assign n13358 = n7255 & ~n13357;
  assign n13359 = pi54 & ~n13358;
  assign n13360 = ~n13352 & n13359;
  assign n13361 = pi100 & ~n13351;
  assign n13362 = pi38 & ~n13357;
  assign n13363 = ~pi100 & ~n13362;
  assign n13364 = ~pi178 & ~pi299;
  assign n13365 = ~pi157 & pi299;
  assign n13366 = n7420 & ~n13365;
  assign n13367 = ~n13364 & n13366;
  assign n13368 = n2522 & ~n13367;
  assign n13369 = n8820 & n13368;
  assign n13370 = n13363 & ~n13369;
  assign n13371 = ~n13361 & ~n13370;
  assign n13372 = n8930 & ~n13371;
  assign n13373 = pi75 & ~n13351;
  assign n13374 = ~pi157 & ~pi168;
  assign n13375 = ~n9391 & n13374;
  assign n13376 = pi157 & ~n9393;
  assign n13377 = ~pi157 & n9397;
  assign n13378 = pi168 & ~n13377;
  assign n13379 = ~n13376 & ~n13378;
  assign n13380 = ~n13375 & n13379;
  assign n13381 = ~n12852 & ~n13380;
  assign n13382 = n12812 & ~n13381;
  assign n13383 = ~pi178 & ~n6236;
  assign n13384 = n9383 & n13383;
  assign n13385 = ~n12852 & ~n13384;
  assign n13386 = pi190 & ~n13385;
  assign n13387 = ~pi178 & n12853;
  assign n13388 = ~pi190 & ~n13387;
  assign n13389 = ~n9374 & ~n12852;
  assign n13390 = pi178 & n13389;
  assign n13391 = n13388 & ~n13390;
  assign n13392 = ~n13386 & ~n13391;
  assign n13393 = n12810 & ~n13392;
  assign n13394 = pi232 & ~n13393;
  assign n13395 = ~n13382 & n13394;
  assign n13396 = n12810 & ~n12853;
  assign n13397 = n5744 & n6464;
  assign n13398 = n7263 & n13397;
  assign n13399 = ~pi232 & ~n13398;
  assign n13400 = ~n13396 & n13399;
  assign n13401 = pi39 & ~n13400;
  assign n13402 = ~n13395 & n13401;
  assign n13403 = ~pi151 & n9408;
  assign n13404 = ~pi168 & n9413;
  assign n13405 = ~n13403 & ~n13404;
  assign n13406 = n9410 & ~n13405;
  assign n13407 = pi150 & ~n13406;
  assign n13408 = ~pi151 & n9437;
  assign n13409 = n9434 & ~n13408;
  assign n13410 = ~pi168 & ~n13409;
  assign n13411 = pi168 & n6190;
  assign n13412 = ~pi151 & n9445;
  assign n13413 = n9448 & ~n13412;
  assign n13414 = n13411 & ~n13413;
  assign n13415 = ~pi150 & ~n13414;
  assign n13416 = ~n13410 & n13415;
  assign n13417 = ~n13407 & ~n13416;
  assign n13418 = ~n9437 & ~n11858;
  assign n13419 = ~n6190 & ~n13418;
  assign n13420 = pi299 & ~n13419;
  assign n13421 = ~n13417 & n13420;
  assign n13422 = ~pi173 & n9408;
  assign n13423 = ~n9413 & ~n13422;
  assign n13424 = n6190 & ~n13423;
  assign n13425 = ~pi190 & n13424;
  assign n13426 = n3084 & n13425;
  assign n13427 = ~pi173 & pi190;
  assign n13428 = n9411 & n13427;
  assign n13429 = pi185 & ~n13428;
  assign n13430 = ~n13426 & n13429;
  assign n13431 = ~pi173 & n9437;
  assign n13432 = n9474 & ~n13431;
  assign n13433 = ~pi190 & ~n13432;
  assign n13434 = ~pi185 & ~n13433;
  assign n13435 = pi173 & n9472;
  assign n13436 = pi190 & ~n13435;
  assign n13437 = n9467 & n13436;
  assign n13438 = n13434 & ~n13437;
  assign n13439 = ~n13430 & ~n13438;
  assign n13440 = ~n6190 & ~n9459;
  assign n13441 = ~pi299 & ~n13440;
  assign n13442 = ~n13439 & n13441;
  assign n13443 = ~n13421 & ~n13442;
  assign n13444 = pi232 & ~n13443;
  assign n13445 = ~pi39 & ~n13444;
  assign n13446 = ~n6166 & ~n9457;
  assign n13447 = ~pi232 & ~n13446;
  assign n13448 = ~n9437 & n13447;
  assign n13449 = n13445 & ~n13448;
  assign n13450 = ~n13402 & ~n13449;
  assign n13451 = ~pi38 & ~n13450;
  assign n13452 = ~pi143 & ~n8948;
  assign n13453 = pi143 & ~n8950;
  assign n13454 = pi165 & ~n13453;
  assign n13455 = ~n13452 & n13454;
  assign n13456 = ~pi165 & n8954;
  assign n13457 = pi143 & n13456;
  assign n13458 = ~n13455 & ~n13457;
  assign n13459 = pi38 & n13458;
  assign n13460 = n2571 & ~n13459;
  assign n13461 = ~n13451 & n13460;
  assign n13462 = pi87 & n13363;
  assign n13463 = ~n13361 & ~n13462;
  assign n13464 = ~n13461 & n13463;
  assign n13465 = n2573 & ~n13464;
  assign n13466 = ~n13373 & ~n13465;
  assign n13467 = ~n13372 & n13466;
  assign n13468 = ~pi54 & ~n13467;
  assign n13469 = ~n13360 & ~n13468;
  assign n13470 = ~pi74 & ~n13469;
  assign n13471 = n13354 & ~n13470;
  assign n13472 = pi55 & ~n13329;
  assign n13473 = pi54 & n13330;
  assign n13474 = ~pi92 & ~n13473;
  assign n13475 = pi150 & n7420;
  assign n13476 = n2522 & ~n13475;
  assign n13477 = n3345 & n13476;
  assign n13478 = n13474 & n13477;
  assign n13479 = n13339 & ~n13478;
  assign n13480 = n13472 & ~n13479;
  assign n13481 = ~n13471 & ~n13480;
  assign n13482 = n2531 & n13481;
  assign n13483 = n13342 & ~n13482;
  assign n13484 = ~n13334 & ~n13483;
  assign n13485 = ~pi118 & n13484;
  assign n13486 = ~n9564 & ~n13342;
  assign n13487 = n8934 & n13367;
  assign n13488 = n8863 & ~n13487;
  assign n13489 = n13363 & ~n13488;
  assign n13490 = ~n13361 & ~n13489;
  assign n13491 = n8930 & ~n13490;
  assign n13492 = ~n6190 & n9239;
  assign n13493 = ~n9251 & ~n13492;
  assign n13494 = ~pi173 & ~n13493;
  assign n13495 = pi185 & ~n13494;
  assign n13496 = ~n6190 & ~n9239;
  assign n13497 = n6190 & ~n9085;
  assign n13498 = ~n13496 & ~n13497;
  assign n13499 = pi173 & n13498;
  assign n13500 = n13495 & ~n13499;
  assign n13501 = ~n9133 & ~n13496;
  assign n13502 = pi173 & n13501;
  assign n13503 = ~n9246 & ~n13492;
  assign n13504 = ~pi173 & ~n13503;
  assign n13505 = ~pi185 & ~n13504;
  assign n13506 = ~n13502 & n13505;
  assign n13507 = pi190 & ~n13506;
  assign n13508 = ~n13500 & n13507;
  assign n13509 = ~n9322 & ~n13496;
  assign n13510 = pi173 & n13509;
  assign n13511 = ~pi173 & n9239;
  assign n13512 = ~pi185 & ~n13511;
  assign n13513 = ~n13510 & n13512;
  assign n13514 = ~pi190 & ~n13513;
  assign n13515 = ~pi173 & ~n9234;
  assign n13516 = pi173 & ~n9643;
  assign n13517 = ~n13515 & ~n13516;
  assign n13518 = n6190 & n13517;
  assign n13519 = ~n13492 & ~n13518;
  assign n13520 = pi185 & n13519;
  assign n13521 = n13514 & ~n13520;
  assign n13522 = ~n13508 & ~n13521;
  assign n13523 = ~pi299 & n13522;
  assign n13524 = ~pi168 & n9305;
  assign n13525 = ~pi151 & ~n13524;
  assign n13526 = ~n9302 & n13525;
  assign n13527 = pi168 & ~n13526;
  assign n13528 = pi151 & ~n9295;
  assign n13529 = ~n13525 & ~n13528;
  assign n13530 = ~n13492 & ~n13529;
  assign n13531 = ~n13527 & n13530;
  assign n13532 = pi150 & ~n13531;
  assign n13533 = n6190 & ~n9264;
  assign n13534 = ~n13496 & ~n13533;
  assign n13535 = pi151 & ~n13534;
  assign n13536 = pi168 & n13535;
  assign n13537 = n13532 & ~n13536;
  assign n13538 = n9239 & ~n13411;
  assign n13539 = pi168 & n9246;
  assign n13540 = ~pi151 & ~n13539;
  assign n13541 = ~n13538 & n13540;
  assign n13542 = ~pi168 & n13509;
  assign n13543 = pi168 & n13501;
  assign n13544 = ~n13542 & ~n13543;
  assign n13545 = pi151 & n13544;
  assign n13546 = ~pi150 & ~n13545;
  assign n13547 = ~n13541 & n13546;
  assign n13548 = ~n13537 & ~n13547;
  assign n13549 = pi299 & n13548;
  assign n13550 = ~n13523 & ~n13549;
  assign n13551 = pi232 & n13550;
  assign n13552 = ~pi232 & n9239;
  assign n13553 = ~pi39 & ~n13552;
  assign n13554 = ~n13551 & n13553;
  assign n13555 = pi168 & n8982;
  assign n13556 = pi157 & n8988;
  assign n13557 = ~n13555 & ~n13556;
  assign n13558 = n6199 & ~n13557;
  assign n13559 = n8959 & n13558;
  assign n13560 = pi299 & ~n13559;
  assign n13561 = ~n13364 & ~n13560;
  assign n13562 = n8862 & ~n13561;
  assign n13563 = pi178 & ~n9010;
  assign n13564 = ~pi190 & ~n13563;
  assign n13565 = ~pi299 & ~n13564;
  assign n13566 = ~n13562 & ~n13565;
  assign n13567 = pi232 & ~n13566;
  assign n13568 = ~n9008 & ~n9384;
  assign n13569 = ~pi178 & ~n9000;
  assign n13570 = ~n13568 & n13569;
  assign n13571 = pi190 & ~n13570;
  assign n13572 = ~pi299 & ~n8974;
  assign n13573 = pi178 & ~n13568;
  assign n13574 = ~n8976 & n13573;
  assign n13575 = n13572 & ~n13574;
  assign n13576 = n13571 & n13575;
  assign n13577 = n13567 & ~n13576;
  assign n13578 = ~pi232 & n8862;
  assign n13579 = ~n13577 & ~n13578;
  assign n13580 = pi39 & n13579;
  assign n13581 = ~pi38 & ~n13580;
  assign n13582 = ~n13554 & n13581;
  assign n13583 = n13460 & ~n13582;
  assign n13584 = ~n8863 & n13462;
  assign n13585 = ~n13361 & ~n13584;
  assign n13586 = ~n13583 & n13585;
  assign n13587 = n2573 & ~n13586;
  assign n13588 = ~n13373 & ~n13587;
  assign n13589 = ~n13491 & n13588;
  assign n13590 = ~pi54 & ~n13589;
  assign n13591 = ~n13360 & ~n13590;
  assign n13592 = ~pi74 & ~n13591;
  assign n13593 = n13354 & ~n13592;
  assign n13594 = ~pi92 & n8934;
  assign n13595 = n13475 & n13594;
  assign n13596 = n13336 & ~n13595;
  assign n13597 = n8862 & n13596;
  assign n13598 = ~n13337 & ~n13597;
  assign n13599 = n7255 & ~n13598;
  assign n13600 = n13335 & ~n13599;
  assign n13601 = n13472 & ~n13600;
  assign n13602 = n2531 & ~n13601;
  assign n13603 = ~n13593 & n13602;
  assign n13604 = ~n13486 & ~n13603;
  assign n13605 = ~n13334 & ~n13604;
  assign n13606 = pi118 & n13605;
  assign n13607 = ~n13485 & ~n13606;
  assign n13608 = ~n13321 & n13607;
  assign n13609 = ~pi118 & ~n8831;
  assign n13610 = n13605 & n13609;
  assign n13611 = n13484 & ~n13609;
  assign n13612 = n13321 & ~n13611;
  assign n13613 = ~n13610 & n13612;
  assign po276 = n13608 | n13613;
  assign n13615 = pi128 & pi228;
  assign n13616 = ~n12806 & n13615;
  assign n13617 = pi87 & ~n13615;
  assign n13618 = ~n7310 & ~n13615;
  assign n13619 = pi100 & ~n13618;
  assign n13620 = ~n2607 & n5792;
  assign n13621 = n7464 & n13620;
  assign n13622 = ~n2527 & n5975;
  assign n13623 = n7468 & n13622;
  assign n13624 = ~n13621 & ~n13623;
  assign n13625 = pi39 & ~n13624;
  assign n13626 = pi299 & n6417;
  assign n13627 = ~n6384 & ~n13626;
  assign n13628 = n7420 & ~n13627;
  assign n13629 = pi109 & ~n13628;
  assign n13630 = ~n2978 & n11448;
  assign n13631 = ~n13629 & ~n13630;
  assign n13632 = n7389 & n9981;
  assign n13633 = n11447 & ~n13632;
  assign n13634 = n2774 & ~n13633;
  assign n13635 = ~pi97 & ~n13634;
  assign n13636 = n2939 & ~n13635;
  assign n13637 = ~pi46 & n13636;
  assign n13638 = n2978 & n13637;
  assign n13639 = n13631 & ~n13638;
  assign n13640 = ~n6308 & ~n13628;
  assign n13641 = ~n6388 & n13628;
  assign n13642 = ~n13640 & ~n13641;
  assign n13643 = ~n13639 & n13642;
  assign n13644 = ~pi91 & ~n13643;
  assign n13645 = ~n6355 & ~n13644;
  assign n13646 = n2696 & n13645;
  assign n13647 = ~n2747 & ~n13646;
  assign n13648 = n2508 & ~n13647;
  assign n13649 = n12881 & n13648;
  assign n13650 = ~n13625 & ~n13649;
  assign n13651 = ~pi38 & ~n13650;
  assign n13652 = ~pi228 & n13651;
  assign n13653 = ~n13615 & ~n13652;
  assign n13654 = ~pi100 & ~n13653;
  assign n13655 = ~pi87 & ~n13654;
  assign n13656 = ~n13619 & n13655;
  assign n13657 = ~pi75 & ~n13656;
  assign n13658 = ~n13617 & n13657;
  assign n13659 = ~n7311 & ~n13615;
  assign n13660 = pi75 & ~n13659;
  assign n13661 = ~pi92 & ~n13660;
  assign n13662 = ~n13658 & n13661;
  assign n13663 = ~n7316 & ~n13615;
  assign n13664 = pi92 & n13663;
  assign n13665 = ~n13662 & ~n13664;
  assign n13666 = n12806 & n13665;
  assign po277 = n13616 | n13666;
  assign n13668 = ~pi31 & ~pi80;
  assign n13669 = pi818 & n13668;
  assign n13670 = n7371 & ~n7380;
  assign n13671 = ~n7376 & ~n13670;
  assign n13672 = ~pi120 & ~n7380;
  assign n13673 = ~pi1093 & n13672;
  assign n13674 = n13671 & ~n13673;
  assign n13675 = n2522 & n7426;
  assign n13676 = pi120 & ~n7371;
  assign n13677 = ~n7483 & n13676;
  assign n13678 = n13675 & ~n13677;
  assign n13679 = ~pi120 & pi1093;
  assign n13680 = n7483 & ~n13679;
  assign n13681 = ~n13678 & ~n13680;
  assign n13682 = n7485 & ~n13681;
  assign n13683 = ~pi120 & ~pi1093;
  assign n13684 = pi100 & ~n13683;
  assign n13685 = ~n7371 & n13684;
  assign n13686 = ~n13682 & n13685;
  assign n13687 = ~pi1093 & n7409;
  assign n13688 = pi120 & n13687;
  assign n13689 = ~pi39 & ~n13688;
  assign n13690 = pi122 & ~n7400;
  assign n13691 = n7368 & n7399;
  assign n13692 = ~pi829 & n13691;
  assign n13693 = ~pi122 & ~n13692;
  assign n13694 = ~n10225 & n13693;
  assign n13695 = ~n2913 & ~n13694;
  assign n13696 = ~n13690 & n13695;
  assign n13697 = n6210 & ~n13696;
  assign n13698 = ~pi122 & n7368;
  assign n13699 = n7490 & ~n13691;
  assign n13700 = ~n13698 & n13699;
  assign n13701 = ~n13697 & ~n13700;
  assign n13702 = n13689 & n13701;
  assign n13703 = ~n7371 & n13679;
  assign n13704 = ~n13676 & ~n13703;
  assign n13705 = ~n5745 & n13704;
  assign n13706 = pi299 & ~n13705;
  assign n13707 = ~n8573 & ~n13704;
  assign n13708 = n5745 & ~n13707;
  assign n13709 = n13706 & ~n13708;
  assign n13710 = pi39 & ~n13709;
  assign n13711 = n8624 & ~n13704;
  assign n13712 = n13710 & ~n13711;
  assign n13713 = ~n13702 & ~n13712;
  assign n13714 = ~pi38 & ~n13713;
  assign n13715 = pi38 & n13683;
  assign n13716 = ~pi100 & ~n13715;
  assign n13717 = ~n7560 & n13716;
  assign n13718 = ~n13714 & n13717;
  assign n13719 = ~n13686 & ~n13718;
  assign n13720 = ~pi87 & ~n13719;
  assign n13721 = n7498 & ~n13683;
  assign n13722 = n7490 & ~n13698;
  assign n13723 = ~n7567 & n13722;
  assign n13724 = n7496 & ~n13723;
  assign n13725 = ~n2615 & n7371;
  assign n13726 = pi87 & ~n13725;
  assign n13727 = ~n13724 & n13726;
  assign n13728 = n13721 & n13727;
  assign n13729 = ~n13720 & ~n13728;
  assign n13730 = ~pi75 & ~n13729;
  assign n13731 = ~n7427 & n13703;
  assign n13732 = ~pi1091 & ~n7370;
  assign n13733 = ~n7507 & ~n13732;
  assign n13734 = pi120 & ~n13733;
  assign n13735 = ~n7421 & ~n13734;
  assign n13736 = ~n13731 & n13735;
  assign n13737 = n3258 & n13736;
  assign n13738 = ~n7422 & n13704;
  assign n13739 = pi75 & ~n13738;
  assign n13740 = ~n13737 & n13739;
  assign n13741 = ~n13730 & ~n13740;
  assign n13742 = n7380 & n13741;
  assign n13743 = n13674 & ~n13742;
  assign n13744 = n7430 & ~n13683;
  assign n13745 = ~n13697 & ~n13699;
  assign n13746 = n13689 & n13745;
  assign n13747 = n8624 & ~n13683;
  assign n13748 = pi39 & ~n13747;
  assign n13749 = ~n8574 & ~n13683;
  assign n13750 = pi299 & n13749;
  assign n13751 = n13748 & ~n13750;
  assign n13752 = ~n13746 & ~n13751;
  assign n13753 = ~pi38 & ~n13752;
  assign n13754 = n13716 & ~n13753;
  assign n13755 = pi120 & n7483;
  assign n13756 = ~pi120 & n13675;
  assign n13757 = ~n13755 & ~n13756;
  assign n13758 = n7485 & ~n13757;
  assign n13759 = n13684 & ~n13758;
  assign n13760 = ~n13754 & ~n13759;
  assign n13761 = ~pi87 & ~n13760;
  assign n13762 = ~n13721 & ~n13761;
  assign n13763 = ~pi75 & ~n13762;
  assign n13764 = ~n13744 & ~n13763;
  assign n13765 = n7380 & n13764;
  assign n13766 = ~n13673 & ~n13765;
  assign n13767 = n7376 & n13766;
  assign n13768 = ~n13743 & ~n13767;
  assign n13769 = n13669 & ~n13768;
  assign n13770 = ~po1038 & ~n13769;
  assign n13771 = ~n7376 & n13704;
  assign n13772 = pi120 & ~n13771;
  assign n13773 = ~n13683 & ~n13771;
  assign n13774 = n13669 & n13773;
  assign n13775 = po1038 & ~n13774;
  assign n13776 = ~n13772 & n13775;
  assign n13777 = ~n7588 & ~n13776;
  assign n13778 = pi951 & pi982;
  assign n13779 = pi1092 & n13778;
  assign n13780 = pi1093 & n13779;
  assign n13781 = ~pi120 & ~n13780;
  assign n13782 = ~n13771 & ~n13781;
  assign n13783 = n13775 & ~n13782;
  assign n13784 = n7588 & ~n13783;
  assign n13785 = ~n13777 & ~n13784;
  assign n13786 = ~n13770 & ~n13785;
  assign n13787 = pi120 & n7428;
  assign n13788 = ~pi1091 & n13780;
  assign n13789 = ~pi120 & ~n13788;
  assign n13790 = n6210 & n13779;
  assign n13791 = ~pi122 & n9405;
  assign n13792 = n2935 & n10262;
  assign n13793 = n7424 & n13792;
  assign n13794 = n8792 & n13793;
  assign n13795 = n13791 & n13794;
  assign n13796 = n2695 & n13795;
  assign n13797 = n13790 & ~n13796;
  assign n13798 = n13789 & ~n13797;
  assign n13799 = ~n13787 & ~n13798;
  assign n13800 = ~n7421 & ~n13799;
  assign n13801 = n7421 & n13781;
  assign n13802 = ~n13800 & ~n13801;
  assign n13803 = n3258 & n13802;
  assign n13804 = ~n3258 & ~n13781;
  assign n13805 = pi75 & ~n13804;
  assign n13806 = ~n13803 & n13805;
  assign n13807 = pi950 & n2522;
  assign n13808 = n7403 & n7424;
  assign n13809 = n13807 & n13808;
  assign n13810 = n13790 & ~n13809;
  assign n13811 = n13789 & ~n13810;
  assign n13812 = ~n13755 & ~n13811;
  assign n13813 = ~pi39 & n7484;
  assign n13814 = ~n13812 & n13813;
  assign n13815 = pi100 & ~n13814;
  assign n13816 = ~pi38 & ~n13815;
  assign n13817 = ~n7485 & n13781;
  assign n13818 = ~n13816 & ~n13817;
  assign n13819 = ~n13687 & n13745;
  assign n13820 = pi120 & n13819;
  assign n13821 = ~pi39 & ~n13820;
  assign n13822 = pi829 & pi1092;
  assign n13823 = n2713 & n7391;
  assign n13824 = n7381 & n13823;
  assign n13825 = n7386 & ~n13824;
  assign n13826 = pi950 & n7398;
  assign n13827 = ~n13825 & n13826;
  assign n13828 = pi122 & ~n13827;
  assign n13829 = n13778 & n13828;
  assign n13830 = n13822 & n13829;
  assign n13831 = pi824 & n13827;
  assign n13832 = n13779 & ~n13831;
  assign n13833 = ~pi829 & n13832;
  assign n13834 = n7403 & n13779;
  assign n13835 = n7407 & ~n10224;
  assign n13836 = pi950 & n13835;
  assign n13837 = n13834 & ~n13836;
  assign n13838 = ~n13833 & ~n13837;
  assign n13839 = ~n13830 & n13838;
  assign n13840 = n7431 & ~n13839;
  assign n13841 = n7493 & n13779;
  assign n13842 = ~n13840 & ~n13841;
  assign n13843 = pi1091 & ~n13842;
  assign n13844 = n7490 & n13832;
  assign n13845 = ~pi120 & ~n13844;
  assign n13846 = ~n13843 & n13845;
  assign n13847 = n13821 & ~n13846;
  assign n13848 = ~n8569 & ~n13781;
  assign n13849 = ~n8575 & n13848;
  assign n13850 = pi39 & n13849;
  assign n13851 = ~n13847 & ~n13850;
  assign n13852 = n2614 & ~n13851;
  assign n13853 = ~n13818 & ~n13852;
  assign n13854 = ~pi87 & ~n13853;
  assign n13855 = ~n2615 & n13781;
  assign n13856 = pi87 & ~n13855;
  assign n13857 = ~n2913 & ~n6121;
  assign n13858 = n13807 & n13857;
  assign n13859 = n13790 & ~n13858;
  assign n13860 = pi824 & n13807;
  assign n13861 = n13788 & ~n13860;
  assign n13862 = ~n13859 & ~n13861;
  assign n13863 = ~pi120 & ~n13862;
  assign n13864 = ~n7492 & ~n7495;
  assign n13865 = pi120 & ~n13864;
  assign n13866 = n2615 & ~n13865;
  assign n13867 = ~n13863 & n13866;
  assign n13868 = n13856 & ~n13867;
  assign n13869 = ~pi75 & ~n13868;
  assign n13870 = ~n13854 & n13869;
  assign n13871 = ~n13806 & ~n13870;
  assign n13872 = n7380 & ~n13871;
  assign n13873 = n7376 & ~n13872;
  assign n13874 = ~n13704 & ~n13781;
  assign n13875 = ~n7484 & n13874;
  assign n13876 = ~n13698 & n13788;
  assign n13877 = ~n13810 & ~n13876;
  assign n13878 = ~pi120 & ~n13877;
  assign n13879 = ~n13677 & ~n13878;
  assign n13880 = n7484 & ~n13879;
  assign n13881 = ~n13875 & ~n13880;
  assign n13882 = n2532 & n13881;
  assign n13883 = ~n2532 & ~n13874;
  assign n13884 = pi100 & ~n13883;
  assign n13885 = ~n13882 & n13884;
  assign n13886 = ~n13687 & n13701;
  assign n13887 = pi120 & n13886;
  assign n13888 = n13722 & n13832;
  assign n13889 = ~pi120 & ~n13888;
  assign n13890 = ~n13843 & n13889;
  assign n13891 = ~n13887 & ~n13890;
  assign n13892 = ~pi39 & ~n13891;
  assign n13893 = ~n5745 & n7371;
  assign n13894 = pi299 & ~n13893;
  assign n13895 = ~n5745 & n13781;
  assign n13896 = ~n6191 & ~n13874;
  assign n13897 = ~n7463 & n13676;
  assign n13898 = ~n7534 & n13790;
  assign n13899 = ~n13876 & ~n13898;
  assign n13900 = ~pi120 & ~n13899;
  assign n13901 = ~n13897 & ~n13900;
  assign n13902 = n6191 & n13901;
  assign n13903 = ~n13896 & ~n13902;
  assign n13904 = n6198 & n13903;
  assign n13905 = ~n6215 & ~n13901;
  assign n13906 = n6215 & n13874;
  assign n13907 = ~n13905 & ~n13906;
  assign n13908 = ~n6198 & ~n13907;
  assign n13909 = ~n13904 & ~n13908;
  assign n13910 = n5745 & n13909;
  assign n13911 = ~n13895 & ~n13910;
  assign n13912 = n13894 & n13911;
  assign n13913 = n6236 & n13903;
  assign n13914 = ~n6236 & ~n13907;
  assign n13915 = ~n13913 & ~n13914;
  assign n13916 = n7529 & n13915;
  assign n13917 = ~n7529 & ~n13874;
  assign n13918 = ~pi299 & ~n13917;
  assign n13919 = ~n13916 & n13918;
  assign n13920 = pi39 & ~n13919;
  assign n13921 = ~n13912 & n13920;
  assign n13922 = ~n13892 & ~n13921;
  assign n13923 = ~pi38 & ~n13922;
  assign n13924 = pi38 & ~n13874;
  assign n13925 = ~pi100 & ~n13924;
  assign n13926 = ~n13923 & n13925;
  assign n13927 = ~n13885 & ~n13926;
  assign n13928 = ~pi87 & ~n13927;
  assign n13929 = ~n13724 & ~n13866;
  assign n13930 = ~n13859 & ~n13876;
  assign n13931 = n13863 & ~n13930;
  assign n13932 = ~n13929 & ~n13931;
  assign n13933 = ~n13725 & ~n13932;
  assign n13934 = n13856 & n13933;
  assign n13935 = ~n13928 & ~n13934;
  assign n13936 = ~pi75 & ~n13935;
  assign n13937 = ~n13797 & ~n13876;
  assign n13938 = ~pi120 & ~n13937;
  assign n13939 = n13735 & ~n13938;
  assign n13940 = n3258 & n13939;
  assign n13941 = ~n7422 & ~n13874;
  assign n13942 = pi75 & ~n13941;
  assign n13943 = ~n13940 & n13942;
  assign n13944 = ~n13936 & ~n13943;
  assign n13945 = n7380 & n13944;
  assign n13946 = n13674 & ~n13945;
  assign n13947 = ~n13873 & ~n13946;
  assign n13948 = n13784 & ~n13947;
  assign n13949 = n13672 & ~n13780;
  assign n13950 = n13948 & ~n13949;
  assign n13951 = ~n7371 & n7487;
  assign n13952 = ~pi39 & ~n13886;
  assign n13953 = ~pi38 & ~n13952;
  assign n13954 = ~n7371 & ~n8569;
  assign n13955 = ~n8575 & n13954;
  assign n13956 = pi39 & n13955;
  assign n13957 = n13953 & ~n13956;
  assign n13958 = ~pi100 & ~n7560;
  assign n13959 = ~n13957 & n13958;
  assign n13960 = ~n13951 & ~n13959;
  assign n13961 = ~pi87 & ~n13960;
  assign n13962 = ~n13727 & ~n13961;
  assign n13963 = ~pi75 & ~n13962;
  assign n13964 = n7371 & ~n7422;
  assign n13965 = pi75 & ~n13964;
  assign n13966 = n7422 & n13733;
  assign n13967 = n13965 & ~n13966;
  assign n13968 = ~n13963 & ~n13967;
  assign n13969 = n13671 & ~n13968;
  assign n13970 = ~n7380 & ~n13771;
  assign n13971 = ~n13969 & ~n13970;
  assign n13972 = ~pi39 & ~n13819;
  assign n13973 = n7473 & ~n13972;
  assign n13974 = ~pi100 & ~n13973;
  assign n13975 = ~n7487 & ~n13974;
  assign n13976 = ~pi87 & ~n13975;
  assign n13977 = ~n7498 & ~n13976;
  assign n13978 = ~pi75 & ~n13977;
  assign n13979 = ~n7430 & ~n13978;
  assign n13980 = ~n13672 & ~n13979;
  assign n13981 = n7376 & n13980;
  assign n13982 = n13971 & ~n13981;
  assign n13983 = pi120 & ~n13982;
  assign n13984 = n13777 & n13983;
  assign n13985 = ~n13950 & ~n13984;
  assign n13986 = ~n13669 & ~n13985;
  assign po278 = n13786 | n13986;
  assign n13988 = pi51 & pi146;
  assign n13989 = pi51 & n6190;
  assign n13990 = ~pi146 & n13989;
  assign n13991 = pi161 & ~n13990;
  assign n13992 = ~pi67 & ~pi71;
  assign n13993 = n2471 & n13992;
  assign n13994 = ~pi51 & n13993;
  assign n13995 = n6190 & ~n13994;
  assign n13996 = ~n13991 & n13995;
  assign n13997 = ~n13988 & n13996;
  assign n13998 = ~pi87 & ~n13997;
  assign n13999 = pi87 & ~n13322;
  assign n14000 = pi232 & ~n13999;
  assign n14001 = ~n13998 & n14000;
  assign n14002 = ~pi134 & ~pi135;
  assign n14003 = ~pi136 & n14002;
  assign n14004 = ~pi130 & n14003;
  assign n14005 = ~pi132 & n14004;
  assign n14006 = ~pi126 & n14005;
  assign n14007 = ~pi121 & n14006;
  assign n14008 = ~pi125 & ~pi133;
  assign n14009 = pi121 & ~n14008;
  assign n14010 = ~pi121 & n14008;
  assign n14011 = ~n14009 & ~n14010;
  assign n14012 = ~n14007 & ~n14011;
  assign n14013 = ~pi87 & n13994;
  assign n14014 = ~n14012 & n14013;
  assign n14015 = po1038 & ~n14014;
  assign n14016 = ~n14001 & n14015;
  assign n14017 = ~pi163 & pi299;
  assign n14018 = ~n11762 & ~n14017;
  assign n14019 = n7420 & n14018;
  assign n14020 = pi87 & ~n14019;
  assign n14021 = ~pi87 & ~n7309;
  assign n14022 = pi299 & ~n13997;
  assign n14023 = ~pi142 & n13989;
  assign n14024 = pi144 & ~n14023;
  assign n14025 = pi51 & pi142;
  assign n14026 = n13995 & ~n14025;
  assign n14027 = ~n14024 & n14026;
  assign n14028 = ~pi299 & ~n14027;
  assign n14029 = pi232 & ~n14028;
  assign n14030 = ~n14022 & n14029;
  assign n14031 = n14021 & ~n14030;
  assign n14032 = ~n13994 & n14031;
  assign n14033 = pi100 & n14030;
  assign n14034 = n2537 & ~n14033;
  assign n14035 = pi38 & ~n14030;
  assign n14036 = ~pi100 & ~n14035;
  assign n14037 = pi38 & ~n13994;
  assign n14038 = ~pi100 & ~n14037;
  assign n14039 = ~n14036 & ~n14038;
  assign n14040 = n2760 & n9976;
  assign n14041 = n12733 & n14040;
  assign n14042 = pi77 & n14041;
  assign n14043 = ~pi86 & n14042;
  assign n14044 = ~pi24 & pi314;
  assign n14045 = n9077 & n14044;
  assign n14046 = n8784 & n14045;
  assign n14047 = n14043 & n14046;
  assign n14048 = n3085 & n14047;
  assign n14049 = ~pi51 & ~n13993;
  assign n14050 = ~n2698 & ~n14049;
  assign n14051 = ~pi77 & n14041;
  assign n14052 = pi86 & n14051;
  assign n14053 = ~n14043 & ~n14052;
  assign n14054 = n10871 & ~n14053;
  assign n14055 = n13993 & ~n14054;
  assign n14056 = ~pi24 & n11451;
  assign n14057 = n14051 & n14056;
  assign n14058 = n14055 & ~n14057;
  assign n14059 = ~n14050 & ~n14058;
  assign n14060 = n3085 & n14059;
  assign n14061 = n13994 & ~n14060;
  assign n14062 = ~pi58 & n14051;
  assign n14063 = n8873 & n14062;
  assign n14064 = n9077 & n14063;
  assign n14065 = pi72 & n3084;
  assign n14066 = n14064 & n14065;
  assign n14067 = n14061 & ~n14066;
  assign n14068 = ~n14048 & n14067;
  assign n14069 = ~n6190 & ~n14068;
  assign n14070 = ~pi51 & n6190;
  assign n14071 = ~n14067 & n14070;
  assign n14072 = ~n14069 & ~n14071;
  assign n14073 = n6190 & ~n14061;
  assign n14074 = ~pi142 & ~n14073;
  assign n14075 = n6190 & n14049;
  assign n14076 = n2686 & n9409;
  assign n14077 = ~n14075 & ~n14076;
  assign n14078 = n3085 & ~n14059;
  assign n14079 = ~n14077 & ~n14078;
  assign n14080 = pi142 & ~n14079;
  assign n14081 = ~n14074 & ~n14080;
  assign n14082 = n13994 & ~n14048;
  assign n14083 = ~n14060 & n14082;
  assign n14084 = ~n6190 & ~n14083;
  assign n14085 = ~n13995 & ~n14084;
  assign n14086 = ~n14081 & ~n14085;
  assign n14087 = n14072 & ~n14086;
  assign n14088 = pi144 & ~n14087;
  assign n14089 = ~n6190 & n14068;
  assign n14090 = ~n10871 & ~n11451;
  assign n14091 = n11448 & ~n14090;
  assign n14092 = n2698 & n14091;
  assign n14093 = ~pi72 & ~n14092;
  assign n14094 = n6367 & ~n14093;
  assign n14095 = n6190 & ~n14094;
  assign n14096 = ~n14089 & ~n14095;
  assign n14097 = ~pi142 & ~n14096;
  assign n14098 = n14076 & n14092;
  assign n14099 = n2699 & n14065;
  assign n14100 = ~n13989 & ~n14099;
  assign n14101 = n6190 & ~n14100;
  assign n14102 = ~n14069 & ~n14101;
  assign n14103 = ~n14098 & n14102;
  assign n14104 = pi142 & n14103;
  assign n14105 = ~pi144 & ~n14104;
  assign n14106 = ~n14097 & n14105;
  assign n14107 = pi180 & ~n14106;
  assign n14108 = ~n14088 & n14107;
  assign n14109 = n14024 & ~n14068;
  assign n14110 = ~pi314 & ~n14091;
  assign n14111 = pi314 & ~n11449;
  assign n14112 = ~n14110 & ~n14111;
  assign n14113 = n2518 & n14112;
  assign n14114 = n7394 & n14113;
  assign n14115 = ~pi51 & ~n14114;
  assign n14116 = ~n14099 & n14115;
  assign n14117 = n6190 & ~n14116;
  assign n14118 = ~n14069 & ~n14117;
  assign n14119 = pi142 & n14118;
  assign n14120 = n2698 & n14112;
  assign n14121 = ~pi72 & ~n14120;
  assign n14122 = n6367 & ~n14121;
  assign n14123 = n6190 & ~n14122;
  assign n14124 = ~n14089 & ~n14123;
  assign n14125 = ~pi142 & ~n14124;
  assign n14126 = ~pi144 & ~n14125;
  assign n14127 = ~n14119 & n14126;
  assign n14128 = ~pi180 & ~n14127;
  assign n14129 = ~n14109 & n14128;
  assign n14130 = ~pi179 & ~n14129;
  assign n14131 = ~n14108 & n14130;
  assign n14132 = ~n14066 & n14085;
  assign n14133 = ~n14048 & n14132;
  assign n14134 = n14024 & ~n14133;
  assign n14135 = n13110 & n14045;
  assign n14136 = ~pi51 & n14135;
  assign n14137 = ~pi72 & ~n14136;
  assign n14138 = n6367 & ~n14137;
  assign n14139 = n6190 & ~n14138;
  assign n14140 = ~n14089 & ~n14139;
  assign n14141 = ~pi142 & ~n14140;
  assign n14142 = n14076 & n14136;
  assign n14143 = n14102 & ~n14142;
  assign n14144 = pi142 & n14143;
  assign n14145 = ~pi144 & ~n14144;
  assign n14146 = ~n14141 & n14145;
  assign n14147 = ~pi180 & ~n14146;
  assign n14148 = ~n14134 & n14147;
  assign n14149 = ~pi144 & n14102;
  assign n14150 = pi144 & n14132;
  assign n14151 = ~n14023 & ~n14150;
  assign n14152 = ~n14149 & n14151;
  assign n14153 = pi180 & ~n14152;
  assign n14154 = pi179 & ~n14153;
  assign n14155 = ~n14148 & n14154;
  assign n14156 = ~n14131 & ~n14155;
  assign n14157 = ~pi299 & ~n14156;
  assign n14158 = ~pi161 & ~n13990;
  assign n14159 = ~n14102 & n14158;
  assign n14160 = n13991 & ~n14132;
  assign n14161 = ~n14159 & ~n14160;
  assign n14162 = n9262 & ~n14161;
  assign n14163 = pi146 & n14143;
  assign n14164 = ~pi146 & ~n14140;
  assign n14165 = ~pi161 & ~n14164;
  assign n14166 = ~n14163 & n14165;
  assign n14167 = n13991 & ~n14133;
  assign n14168 = ~n14166 & ~n14167;
  assign n14169 = n9292 & ~n14168;
  assign n14170 = ~n14162 & ~n14169;
  assign n14171 = pi156 & ~n14170;
  assign n14172 = ~n13990 & ~n14068;
  assign n14173 = n9292 & n14172;
  assign n14174 = ~pi146 & ~n14073;
  assign n14175 = pi146 & ~n14079;
  assign n14176 = ~n14174 & ~n14175;
  assign n14177 = ~n14085 & ~n14176;
  assign n14178 = n14072 & ~n14177;
  assign n14179 = n9262 & ~n14178;
  assign n14180 = pi161 & ~n14179;
  assign n14181 = ~n14173 & n14180;
  assign n14182 = ~pi146 & ~n14096;
  assign n14183 = n9262 & ~n14182;
  assign n14184 = pi146 & n14103;
  assign n14185 = n14183 & ~n14184;
  assign n14186 = ~pi146 & ~n14124;
  assign n14187 = pi146 & n14118;
  assign n14188 = ~n14186 & ~n14187;
  assign n14189 = n9292 & n14188;
  assign n14190 = ~pi161 & ~n14189;
  assign n14191 = ~n14185 & n14190;
  assign n14192 = ~pi156 & ~n14191;
  assign n14193 = ~n14181 & n14192;
  assign n14194 = ~n14171 & ~n14193;
  assign n14195 = ~n14157 & n14194;
  assign n14196 = n9456 & ~n14195;
  assign n14197 = n3085 & n14064;
  assign n14198 = n13994 & ~n14197;
  assign n14199 = ~n6190 & ~n14198;
  assign n14200 = ~pi51 & ~n2521;
  assign n14201 = n6190 & ~n14200;
  assign n14202 = ~n14199 & ~n14201;
  assign n14203 = pi142 & ~n14202;
  assign n14204 = ~n6222 & ~n14199;
  assign n14205 = ~pi142 & ~n14204;
  assign n14206 = n6439 & ~n14205;
  assign n14207 = ~n14203 & n14206;
  assign n14208 = ~n8973 & ~n14207;
  assign n14209 = ~pi287 & n6190;
  assign n14210 = ~pi51 & n14209;
  assign n14211 = ~n14202 & ~n14210;
  assign n14212 = pi224 & ~n14023;
  assign n14213 = n14211 & n14212;
  assign n14214 = ~n14208 & ~n14213;
  assign n14215 = ~n13994 & ~n14023;
  assign n14216 = ~n6439 & ~n14215;
  assign n14217 = ~n6439 & n14075;
  assign n14218 = ~pi144 & ~n14217;
  assign n14219 = ~n14216 & n14218;
  assign n14220 = ~n14214 & n14219;
  assign n14221 = ~pi51 & ~n14198;
  assign n14222 = ~pi287 & ~n14221;
  assign n14223 = ~n14075 & ~n14209;
  assign n14224 = ~n14222 & ~n14223;
  assign n14225 = ~n14026 & ~n14224;
  assign n14226 = n8973 & ~n14225;
  assign n14227 = n13993 & n14226;
  assign n14228 = pi144 & ~n14216;
  assign n14229 = pi51 & ~n6190;
  assign n14230 = ~n14221 & ~n14229;
  assign n14231 = n6439 & ~n14025;
  assign n14232 = n14230 & n14231;
  assign n14233 = n14228 & ~n14232;
  assign n14234 = ~n14227 & n14233;
  assign n14235 = pi181 & ~n14234;
  assign n14236 = ~n14220 & n14235;
  assign n14237 = ~n14207 & n14219;
  assign n14238 = ~pi181 & ~n14233;
  assign n14239 = ~n14237 & n14238;
  assign n14240 = ~n14236 & ~n14239;
  assign n14241 = ~pi299 & n14240;
  assign n14242 = ~n13994 & ~n13997;
  assign n14243 = ~n5744 & ~n14242;
  assign n14244 = ~n13990 & ~n14198;
  assign n14245 = pi161 & ~n14244;
  assign n14246 = pi146 & ~n14202;
  assign n14247 = ~pi146 & ~n14204;
  assign n14248 = ~pi161 & ~n14247;
  assign n14249 = ~n14246 & n14248;
  assign n14250 = ~n14245 & ~n14249;
  assign n14251 = n5744 & ~n14250;
  assign n14252 = n9659 & ~n14251;
  assign n14253 = ~n14243 & n14252;
  assign n14254 = pi232 & ~n14253;
  assign n14255 = ~n14241 & n14254;
  assign n14256 = ~n8959 & ~n14251;
  assign n14257 = n14158 & n14211;
  assign n14258 = n14197 & ~n14209;
  assign n14259 = n13994 & ~n14258;
  assign n14260 = n13991 & ~n14259;
  assign n14261 = ~n14257 & ~n14260;
  assign n14262 = pi216 & ~n14261;
  assign n14263 = ~n14256 & ~n14262;
  assign n14264 = ~n14243 & ~n14263;
  assign n14265 = n9693 & n14264;
  assign n14266 = n14255 & ~n14265;
  assign n14267 = pi39 & ~n14266;
  assign n14268 = ~n6592 & ~n7465;
  assign n14269 = n14197 & ~n14268;
  assign n14270 = ~pi232 & ~n14269;
  assign n14271 = n13994 & n14270;
  assign n14272 = n14267 & ~n14271;
  assign n14273 = ~pi39 & ~pi232;
  assign n14274 = ~n14068 & n14273;
  assign n14275 = ~n14272 & ~n14274;
  assign n14276 = ~n14196 & n14275;
  assign n14277 = ~pi38 & ~n14276;
  assign n14278 = ~n14039 & ~n14277;
  assign n14279 = pi100 & n13994;
  assign n14280 = ~n14278 & ~n14279;
  assign n14281 = n14034 & n14280;
  assign n14282 = ~n14012 & ~n14281;
  assign n14283 = ~n14032 & n14282;
  assign n14284 = ~n14020 & n14283;
  assign n14285 = ~n8959 & n13997;
  assign n14286 = n14158 & ~n14224;
  assign n14287 = n6190 & n6440;
  assign n14288 = n13991 & ~n14287;
  assign n14289 = ~n14286 & ~n14288;
  assign n14290 = n8959 & n14289;
  assign n14291 = ~n14285 & ~n14290;
  assign n14292 = n9693 & n14291;
  assign n14293 = n9659 & ~n13997;
  assign n14294 = n8973 & n14209;
  assign n14295 = n2521 & ~n14025;
  assign n14296 = n14294 & n14295;
  assign n14297 = n14024 & ~n14296;
  assign n14298 = ~pi144 & ~n14026;
  assign n14299 = ~n14226 & n14298;
  assign n14300 = ~n14297 & ~n14299;
  assign n14301 = pi181 & n14300;
  assign n14302 = ~pi181 & n14027;
  assign n14303 = ~pi299 & ~n14302;
  assign n14304 = ~n14301 & n14303;
  assign n14305 = n10280 & ~n14304;
  assign n14306 = ~n14293 & n14305;
  assign n14307 = ~n14292 & n14306;
  assign n14308 = ~pi38 & ~n14307;
  assign n14309 = n6190 & ~n14115;
  assign n14310 = ~n14025 & n14309;
  assign n14311 = pi144 & ~n14310;
  assign n14312 = n6190 & ~n14083;
  assign n14313 = ~pi142 & n14312;
  assign n14314 = n13993 & ~n14047;
  assign n14315 = n9077 & n14058;
  assign n14316 = n14314 & n14315;
  assign n14317 = ~n14050 & ~n14316;
  assign n14318 = n3085 & ~n14317;
  assign n14319 = ~n14077 & ~n14318;
  assign n14320 = pi142 & n14319;
  assign n14321 = ~pi144 & ~n14320;
  assign n14322 = ~n14313 & n14321;
  assign n14323 = pi180 & ~n14322;
  assign n14324 = ~n14311 & n14323;
  assign n14325 = n14024 & ~n14098;
  assign n14326 = ~pi144 & ~n14081;
  assign n14327 = ~pi180 & ~n14326;
  assign n14328 = ~n14325 & n14327;
  assign n14329 = pi179 & ~n14328;
  assign n14330 = ~n14324 & n14329;
  assign n14331 = n14024 & ~n14142;
  assign n14332 = n6190 & ~n14082;
  assign n14333 = ~pi142 & n14332;
  assign n14334 = ~pi51 & ~n14314;
  assign n14335 = n3085 & ~n14334;
  assign n14336 = ~n14077 & ~n14335;
  assign n14337 = pi142 & n14336;
  assign n14338 = ~pi144 & ~n14337;
  assign n14339 = ~n14333 & n14338;
  assign n14340 = ~n14331 & ~n14339;
  assign n14341 = pi180 & n14340;
  assign n14342 = ~pi180 & n14027;
  assign n14343 = ~pi179 & ~n14342;
  assign n14344 = ~n14341 & n14343;
  assign n14345 = ~n14330 & ~n14344;
  assign n14346 = ~pi299 & ~n14345;
  assign n14347 = ~n13988 & n14309;
  assign n14348 = pi161 & ~n14347;
  assign n14349 = pi146 & n14319;
  assign n14350 = ~pi146 & n14312;
  assign n14351 = ~pi161 & ~n14350;
  assign n14352 = ~n14349 & n14351;
  assign n14353 = ~n14348 & ~n14352;
  assign n14354 = n9262 & ~n14353;
  assign n14355 = n13991 & ~n14098;
  assign n14356 = ~pi161 & ~n14176;
  assign n14357 = ~n14355 & ~n14356;
  assign n14358 = n9292 & ~n14357;
  assign n14359 = ~n14354 & ~n14358;
  assign n14360 = pi232 & n14359;
  assign n14361 = pi156 & ~n14360;
  assign n14362 = ~pi39 & ~n14361;
  assign n14363 = ~n14346 & n14362;
  assign n14364 = n14308 & ~n14363;
  assign n14365 = n13991 & ~n14142;
  assign n14366 = pi146 & n14336;
  assign n14367 = ~pi146 & n14332;
  assign n14368 = ~pi161 & ~n14367;
  assign n14369 = ~n14366 & n14368;
  assign n14370 = ~n14365 & ~n14369;
  assign n14371 = n9262 & ~n14370;
  assign n14372 = ~pi158 & n14022;
  assign n14373 = ~n14371 & ~n14372;
  assign n14374 = pi232 & n14373;
  assign n14375 = ~pi156 & ~n14374;
  assign n14376 = n2532 & n14375;
  assign n14377 = ~n14364 & ~n14376;
  assign n14378 = n14036 & n14377;
  assign n14379 = n14034 & ~n14378;
  assign n14380 = n14012 & ~n14379;
  assign n14381 = ~n14020 & ~n14031;
  assign n14382 = n14380 & n14381;
  assign n14383 = ~po1038 & ~n14382;
  assign n14384 = ~n14284 & n14383;
  assign po279 = n14016 | n14384;
  assign n14386 = n7371 & n7378;
  assign n14387 = n7380 & n13968;
  assign n14388 = n13671 & ~n14387;
  assign n14389 = n7380 & n13979;
  assign n14390 = n7376 & ~n14389;
  assign n14391 = ~po1038 & ~n14390;
  assign n14392 = ~n14388 & n14391;
  assign po280 = n14386 | n14392;
  assign n14394 = ~pi110 & n8963;
  assign n14395 = ~n6200 & n14394;
  assign n14396 = n5744 & n14395;
  assign n14397 = pi39 & ~n14396;
  assign n14398 = pi110 & ~n10773;
  assign n14399 = po1057 & n14398;
  assign n14400 = n9903 & n14399;
  assign n14401 = ~pi39 & ~n14400;
  assign n14402 = ~n14397 & ~n14401;
  assign n14403 = po1038 & n14402;
  assign n14404 = pi90 & ~n10174;
  assign n14405 = ~pi111 & ~n6314;
  assign n14406 = ~pi36 & n2800;
  assign n14407 = ~n14405 & n14406;
  assign n14408 = n2469 & ~n14407;
  assign n14409 = ~n2784 & ~n14408;
  assign n14410 = ~n2789 & n14409;
  assign n14411 = ~pi83 & ~n14410;
  assign n14412 = n2786 & ~n14411;
  assign n14413 = ~pi71 & ~n14412;
  assign n14414 = n6324 & ~n14413;
  assign n14415 = ~pi81 & ~n14414;
  assign n14416 = n11235 & ~n14415;
  assign n14417 = ~pi90 & ~n14416;
  assign n14418 = n2697 & ~n14417;
  assign n14419 = ~n14404 & n14418;
  assign n14420 = ~pi72 & ~pi93;
  assign n14421 = n14419 & n14420;
  assign n14422 = pi72 & n2698;
  assign n14423 = n10174 & n14422;
  assign n14424 = ~n14421 & ~n14423;
  assign n14425 = n3084 & ~n14424;
  assign n14426 = ~pi110 & ~n14425;
  assign n14427 = n13117 & ~n14426;
  assign n14428 = n2889 & n14418;
  assign n14429 = ~pi72 & ~n14428;
  assign n14430 = n6367 & ~n14429;
  assign n14431 = ~n13117 & n14430;
  assign n14432 = ~pi39 & ~n14431;
  assign n14433 = ~n14427 & n14432;
  assign n14434 = n2575 & n14433;
  assign n14435 = n6592 & n14395;
  assign n14436 = n7265 & n14394;
  assign n14437 = pi39 & ~n14436;
  assign n14438 = ~n14435 & n14437;
  assign n14439 = pi110 & n13117;
  assign n14440 = ~pi39 & ~n14439;
  assign n14441 = ~n2575 & n14440;
  assign n14442 = ~n14438 & ~n14441;
  assign n14443 = ~po1038 & n14442;
  assign n14444 = ~n14434 & n14443;
  assign po281 = ~n14403 & ~n14444;
  assign n14446 = pi87 & n7420;
  assign n14447 = pi162 & n14446;
  assign n14448 = ~pi125 & n14007;
  assign n14449 = pi125 & pi133;
  assign n14450 = ~n14008 & ~n14449;
  assign n14451 = ~n14448 & ~n14450;
  assign n14452 = n13994 & ~n14451;
  assign n14453 = pi172 & n13989;
  assign n14454 = ~pi152 & n14075;
  assign n14455 = ~n14453 & ~n14454;
  assign n14456 = pi232 & ~n14455;
  assign n14457 = ~n14452 & ~n14456;
  assign n14458 = ~pi87 & ~n14457;
  assign n14459 = po1038 & ~n14458;
  assign n14460 = ~n14447 & n14459;
  assign n14461 = pi299 & n14455;
  assign n14462 = pi232 & ~n14461;
  assign n14463 = pi193 & n13989;
  assign n14464 = ~pi174 & n14075;
  assign n14465 = ~pi299 & ~n14464;
  assign n14466 = ~n14463 & n14465;
  assign n14467 = n14462 & ~n14466;
  assign n14468 = n14021 & ~n14467;
  assign n14469 = ~n13994 & n14468;
  assign n14470 = pi140 & ~pi299;
  assign n14471 = pi162 & pi299;
  assign n14472 = ~n14470 & ~n14471;
  assign n14473 = n7420 & ~n14472;
  assign n14474 = pi87 & ~n14473;
  assign n14475 = n2537 & ~n14279;
  assign n14476 = pi100 & n14467;
  assign n14477 = ~n13994 & n14455;
  assign n14478 = ~n8959 & ~n14477;
  assign n14479 = ~pi152 & n6190;
  assign n14480 = ~n14198 & ~n14479;
  assign n14481 = ~pi152 & n14201;
  assign n14482 = ~n14480 & ~n14481;
  assign n14483 = ~pi172 & ~n14482;
  assign n14484 = ~pi152 & n14204;
  assign n14485 = pi152 & n14230;
  assign n14486 = pi172 & ~n14485;
  assign n14487 = ~n14484 & n14486;
  assign n14488 = ~n14483 & ~n14487;
  assign n14489 = n8959 & n14488;
  assign n14490 = n9292 & ~n14489;
  assign n14491 = ~pi152 & ~n14453;
  assign n14492 = n14211 & n14491;
  assign n14493 = ~n14259 & ~n14453;
  assign n14494 = pi152 & n14493;
  assign n14495 = ~n14492 & ~n14494;
  assign n14496 = n8959 & n14495;
  assign n14497 = n9262 & ~n14496;
  assign n14498 = ~n14490 & ~n14497;
  assign n14499 = ~n14478 & ~n14498;
  assign n14500 = n8973 & n14197;
  assign n14501 = n13994 & ~n14500;
  assign n14502 = ~pi51 & ~n14259;
  assign n14503 = n6190 & ~n14502;
  assign n14504 = ~n14501 & ~n14503;
  assign n14505 = pi174 & ~n14504;
  assign n14506 = ~n6190 & ~n13993;
  assign n14507 = ~n8973 & ~n14506;
  assign n14508 = ~n14229 & n14507;
  assign n14509 = ~n10399 & ~n14199;
  assign n14510 = n8973 & n14509;
  assign n14511 = ~n14508 & ~n14510;
  assign n14512 = ~pi174 & ~n14511;
  assign n14513 = pi180 & ~n14512;
  assign n14514 = ~n14505 & n14513;
  assign n14515 = ~n13989 & ~n14501;
  assign n14516 = pi174 & ~n14515;
  assign n14517 = n8973 & n14204;
  assign n14518 = ~n14508 & ~n14517;
  assign n14519 = ~pi174 & ~n14518;
  assign n14520 = ~pi180 & ~n14519;
  assign n14521 = ~n14516 & n14520;
  assign n14522 = pi193 & ~n14521;
  assign n14523 = ~n14514 & n14522;
  assign n14524 = pi180 & n14210;
  assign n14525 = ~pi51 & ~n14202;
  assign n14526 = n14507 & n14525;
  assign n14527 = ~n14202 & ~n14526;
  assign n14528 = ~n14524 & n14527;
  assign n14529 = ~pi174 & n14528;
  assign n14530 = pi180 & n14259;
  assign n14531 = ~n14501 & ~n14530;
  assign n14532 = pi174 & n14531;
  assign n14533 = ~pi193 & ~n14532;
  assign n14534 = ~n14529 & n14533;
  assign n14535 = ~pi299 & ~n14534;
  assign n14536 = ~n14523 & n14535;
  assign n14537 = ~n14499 & ~n14536;
  assign n14538 = pi232 & ~n14537;
  assign n14539 = ~pi299 & ~n14501;
  assign n14540 = n8959 & n14197;
  assign n14541 = n13994 & ~n14540;
  assign n14542 = pi299 & ~n14541;
  assign n14543 = ~n14539 & ~n14542;
  assign n14544 = ~pi232 & ~n14543;
  assign n14545 = pi39 & ~n14544;
  assign n14546 = ~n14538 & n14545;
  assign n14547 = ~pi232 & ~n14083;
  assign n14548 = ~pi39 & ~n14547;
  assign n14549 = ~pi38 & ~n14548;
  assign n14550 = ~n14546 & n14549;
  assign n14551 = pi38 & ~n14467;
  assign n14552 = ~pi100 & ~n14551;
  assign n14553 = ~n14038 & ~n14552;
  assign n14554 = ~pi145 & ~n14082;
  assign n14555 = ~n6190 & ~n14082;
  assign n14556 = ~n13995 & ~n14555;
  assign n14557 = ~n14060 & n14556;
  assign n14558 = ~n14554 & n14557;
  assign n14559 = n3085 & n14558;
  assign n14560 = ~n14084 & ~n14319;
  assign n14561 = ~n14559 & ~n14560;
  assign n14562 = pi174 & n14561;
  assign n14563 = ~n14084 & ~n14098;
  assign n14564 = pi145 & n14563;
  assign n14565 = ~pi174 & ~n14564;
  assign n14566 = n14076 & n14120;
  assign n14567 = ~n14084 & ~n14566;
  assign n14568 = ~pi145 & n14567;
  assign n14569 = n14565 & ~n14568;
  assign n14570 = pi193 & ~n14569;
  assign n14571 = ~n14562 & n14570;
  assign n14572 = pi174 & ~n14558;
  assign n14573 = ~pi51 & n14564;
  assign n14574 = ~pi145 & ~n14084;
  assign n14575 = ~n14309 & n14574;
  assign n14576 = ~pi174 & ~n14575;
  assign n14577 = ~n14573 & n14576;
  assign n14578 = ~pi193 & ~n14577;
  assign n14579 = ~n14572 & n14578;
  assign n14580 = ~n14571 & ~n14579;
  assign n14581 = n9711 & n14580;
  assign n14582 = ~n13989 & ~n14084;
  assign n14583 = ~pi145 & n14142;
  assign n14584 = ~pi174 & ~n14583;
  assign n14585 = pi145 & n13993;
  assign n14586 = ~n14584 & ~n14585;
  assign n14587 = n14582 & ~n14586;
  assign n14588 = ~n14084 & ~n14332;
  assign n14589 = pi174 & n14588;
  assign n14590 = ~n14587 & ~n14589;
  assign n14591 = ~pi193 & ~n14590;
  assign n14592 = n9716 & ~n14591;
  assign n14593 = pi145 & ~n14075;
  assign n14594 = ~pi145 & ~n14336;
  assign n14595 = pi174 & n14594;
  assign n14596 = ~n14584 & ~n14595;
  assign n14597 = ~n14593 & n14596;
  assign n14598 = ~n14084 & ~n14597;
  assign n14599 = pi193 & n14598;
  assign n14600 = n14592 & ~n14599;
  assign n14601 = ~n14581 & ~n14600;
  assign n14602 = ~pi38 & ~n14601;
  assign n14603 = ~pi152 & ~n14567;
  assign n14604 = pi152 & ~n14560;
  assign n14605 = pi172 & ~n14604;
  assign n14606 = ~n14603 & n14605;
  assign n14607 = ~n14083 & ~n14479;
  assign n14608 = ~pi172 & ~n14607;
  assign n14609 = ~pi152 & n14309;
  assign n14610 = n14608 & ~n14609;
  assign n14611 = ~n14606 & ~n14610;
  assign n14612 = ~pi197 & ~n14611;
  assign n14613 = ~pi172 & n14557;
  assign n14614 = ~n14079 & ~n14084;
  assign n14615 = pi172 & n14614;
  assign n14616 = ~n14613 & ~n14615;
  assign n14617 = pi152 & n14616;
  assign n14618 = pi51 & ~pi172;
  assign n14619 = n6190 & n14618;
  assign n14620 = ~pi152 & ~n14563;
  assign n14621 = pi197 & ~n14620;
  assign n14622 = ~n14619 & n14621;
  assign n14623 = ~n14617 & n14622;
  assign n14624 = pi299 & ~n14623;
  assign n14625 = n9725 & n14624;
  assign n14626 = ~n14612 & n14625;
  assign n14627 = pi152 & n14075;
  assign n14628 = ~n14084 & ~n14627;
  assign n14629 = pi172 & ~n14628;
  assign n14630 = ~pi172 & ~n14454;
  assign n14631 = ~n14085 & n14630;
  assign n14632 = ~n14629 & ~n14631;
  assign n14633 = pi197 & n14632;
  assign n14634 = pi299 & ~n14633;
  assign n14635 = ~n14084 & ~n14336;
  assign n14636 = pi152 & ~n14635;
  assign n14637 = ~n14084 & ~n14142;
  assign n14638 = ~pi152 & ~n14637;
  assign n14639 = ~n14636 & ~n14638;
  assign n14640 = ~pi197 & ~n14618;
  assign n14641 = n14639 & n14640;
  assign n14642 = n14634 & ~n14641;
  assign n14643 = n9727 & n14642;
  assign n14644 = ~n14626 & ~n14643;
  assign n14645 = ~n14602 & n14644;
  assign n14646 = n9456 & ~n14645;
  assign n14647 = ~n14553 & ~n14646;
  assign n14648 = ~n14550 & n14647;
  assign n14649 = ~n14476 & ~n14648;
  assign n14650 = n14475 & n14649;
  assign n14651 = ~n14474 & ~n14650;
  assign n14652 = ~n14469 & n14651;
  assign n14653 = ~n14451 & n14652;
  assign n14654 = ~po1038 & ~n14653;
  assign n14655 = n14099 & ~n14479;
  assign n14656 = n13993 & ~n14066;
  assign n14657 = n14070 & ~n14656;
  assign n14658 = ~pi152 & n14657;
  assign n14659 = ~pi197 & ~n14658;
  assign n14660 = ~n14655 & n14659;
  assign n14661 = ~n6190 & n14099;
  assign n14662 = ~n14657 & ~n14661;
  assign n14663 = ~pi51 & n14332;
  assign n14664 = n14662 & ~n14663;
  assign n14665 = ~pi152 & n14664;
  assign n14666 = pi197 & n14665;
  assign n14667 = ~n14660 & ~n14666;
  assign n14668 = ~n14453 & ~n14667;
  assign n14669 = ~n6190 & ~n14099;
  assign n14670 = ~n14139 & ~n14669;
  assign n14671 = ~pi172 & n14670;
  assign n14672 = n14100 & ~n14142;
  assign n14673 = pi172 & ~n14672;
  assign n14674 = pi152 & ~n14673;
  assign n14675 = pi197 & n14674;
  assign n14676 = ~n14671 & n14675;
  assign n14677 = ~n14668 & ~n14676;
  assign n14678 = n9725 & ~n14677;
  assign n14679 = ~n14098 & n14100;
  assign n14680 = pi152 & ~n14679;
  assign n14681 = n14070 & n14656;
  assign n14682 = n14061 & n14681;
  assign n14683 = ~n14669 & ~n14682;
  assign n14684 = ~pi152 & n14683;
  assign n14685 = ~n14680 & ~n14684;
  assign n14686 = pi172 & n14685;
  assign n14687 = ~n14095 & ~n14669;
  assign n14688 = pi152 & n14687;
  assign n14689 = ~n14071 & ~n14661;
  assign n14690 = ~pi152 & ~n14689;
  assign n14691 = ~pi172 & ~n14690;
  assign n14692 = ~n14688 & n14691;
  assign n14693 = ~pi197 & ~n14692;
  assign n14694 = ~n14686 & n14693;
  assign n14695 = ~n14116 & ~n14669;
  assign n14696 = pi172 & n14695;
  assign n14697 = ~n14123 & ~n14669;
  assign n14698 = ~pi172 & n14697;
  assign n14699 = ~n14696 & ~n14698;
  assign n14700 = pi152 & n14699;
  assign n14701 = ~n14071 & n14664;
  assign n14702 = n14491 & n14701;
  assign n14703 = pi197 & ~n14702;
  assign n14704 = ~n14700 & n14703;
  assign n14705 = n9727 & ~n14704;
  assign n14706 = ~n14694 & n14705;
  assign n14707 = ~n14678 & ~n14706;
  assign n14708 = pi299 & ~n14707;
  assign n14709 = ~n13989 & ~n14048;
  assign n14710 = pi145 & ~n14709;
  assign n14711 = n14681 & ~n14710;
  assign n14712 = ~pi174 & ~n14669;
  assign n14713 = ~n14711 & n14712;
  assign n14714 = ~n14583 & ~n14672;
  assign n14715 = ~n14584 & n14714;
  assign n14716 = ~n14713 & ~n14715;
  assign n14717 = pi193 & ~n14716;
  assign n14718 = n9711 & ~n14717;
  assign n14719 = ~n13989 & n14713;
  assign n14720 = ~pi174 & ~n14719;
  assign n14721 = pi145 & n14670;
  assign n14722 = ~pi145 & n14099;
  assign n14723 = pi174 & ~n14722;
  assign n14724 = ~n14721 & n14723;
  assign n14725 = ~n14720 & ~n14724;
  assign n14726 = ~pi193 & n14725;
  assign n14727 = n14718 & ~n14726;
  assign n14728 = ~n14463 & n14701;
  assign n14729 = pi145 & n14728;
  assign n14730 = ~pi174 & ~n14729;
  assign n14731 = ~pi145 & ~n14463;
  assign n14732 = n14689 & n14731;
  assign n14733 = n14730 & ~n14732;
  assign n14734 = ~pi145 & ~n14679;
  assign n14735 = pi193 & ~n14734;
  assign n14736 = pi145 & n14695;
  assign n14737 = n14735 & ~n14736;
  assign n14738 = ~pi145 & n14687;
  assign n14739 = pi145 & n14697;
  assign n14740 = ~pi193 & ~n14739;
  assign n14741 = ~n14738 & n14740;
  assign n14742 = pi174 & ~n14741;
  assign n14743 = ~n14737 & n14742;
  assign n14744 = n9716 & ~n14743;
  assign n14745 = ~n14733 & n14744;
  assign n14746 = ~n14727 & ~n14745;
  assign n14747 = ~pi38 & ~n14746;
  assign n14748 = ~n14708 & ~n14747;
  assign n14749 = n9456 & ~n14748;
  assign n14750 = ~n7466 & ~n7469;
  assign n14751 = n2522 & ~n14750;
  assign n14752 = ~pi232 & ~n14751;
  assign n14753 = pi39 & ~n14752;
  assign n14754 = ~n5745 & n14455;
  assign n14755 = n2522 & ~n6190;
  assign n14756 = n6190 & ~n14198;
  assign n14757 = ~n14755 & ~n14756;
  assign n14758 = ~pi152 & n14757;
  assign n14759 = ~n14200 & ~n14229;
  assign n14760 = pi152 & ~n14759;
  assign n14761 = ~n14758 & ~n14760;
  assign n14762 = ~n14618 & n14761;
  assign n14763 = ~pi216 & ~n14762;
  assign n14764 = n5744 & n14763;
  assign n14765 = ~n14754 & ~n14764;
  assign n14766 = n9292 & ~n14765;
  assign n14767 = ~n5744 & ~n14455;
  assign n14768 = n9262 & ~n14767;
  assign n14769 = n14197 & n14209;
  assign n14770 = ~n13995 & ~n14769;
  assign n14771 = ~pi152 & n14770;
  assign n14772 = pi172 & ~n14771;
  assign n14773 = n2521 & n14209;
  assign n14774 = ~n13989 & ~n14773;
  assign n14775 = pi152 & n14774;
  assign n14776 = n14772 & ~n14775;
  assign n14777 = pi152 & ~n14287;
  assign n14778 = ~pi152 & ~n14224;
  assign n14779 = ~pi172 & ~n14778;
  assign n14780 = ~n14777 & n14779;
  assign n14781 = pi216 & ~n14780;
  assign n14782 = ~n14776 & n14781;
  assign n14783 = ~n14763 & ~n14782;
  assign n14784 = n5744 & n14783;
  assign n14785 = n14768 & ~n14784;
  assign n14786 = ~n14766 & ~n14785;
  assign n14787 = pi224 & n14774;
  assign n14788 = n6439 & ~n14787;
  assign n14789 = n7529 & ~n14759;
  assign n14790 = n14788 & ~n14789;
  assign n14791 = ~n13989 & ~n14790;
  assign n14792 = pi174 & ~n14791;
  assign n14793 = n7529 & n14757;
  assign n14794 = pi224 & ~n14769;
  assign n14795 = n6439 & ~n14794;
  assign n14796 = ~n13995 & ~n14795;
  assign n14797 = ~n14793 & ~n14796;
  assign n14798 = ~pi174 & n14797;
  assign n14799 = pi193 & ~n14798;
  assign n14800 = ~n14792 & n14799;
  assign n14801 = n6190 & n14221;
  assign n14802 = ~n14755 & ~n14801;
  assign n14803 = ~n14796 & ~n14802;
  assign n14804 = ~pi174 & n14803;
  assign n14805 = ~n7529 & ~n14294;
  assign n14806 = n2522 & ~n14805;
  assign n14807 = pi174 & n14806;
  assign n14808 = ~pi193 & ~n14807;
  assign n14809 = ~n14804 & n14808;
  assign n14810 = ~n14800 & ~n14809;
  assign n14811 = pi180 & n14810;
  assign n14812 = ~n7529 & ~n13995;
  assign n14813 = ~n14802 & ~n14812;
  assign n14814 = ~pi174 & n14813;
  assign n14815 = n2522 & n7529;
  assign n14816 = pi174 & n14815;
  assign n14817 = ~n14463 & ~n14816;
  assign n14818 = ~n14814 & n14817;
  assign n14819 = ~pi180 & ~n14818;
  assign n14820 = ~pi299 & ~n14819;
  assign n14821 = ~n14811 & n14820;
  assign n14822 = n14786 & ~n14821;
  assign n14823 = pi232 & ~n14822;
  assign n14824 = n14753 & ~n14823;
  assign n14825 = ~pi232 & ~n14099;
  assign n14826 = ~pi39 & ~n14825;
  assign n14827 = ~pi38 & ~n14826;
  assign n14828 = ~n14824 & n14827;
  assign n14829 = ~n14749 & ~n14828;
  assign n14830 = n14552 & n14829;
  assign n14831 = ~n14476 & ~n14830;
  assign n14832 = n2537 & n14831;
  assign n14833 = n14451 & ~n14832;
  assign n14834 = ~n14474 & n14833;
  assign n14835 = ~n14468 & n14834;
  assign n14836 = n14654 & ~n14835;
  assign po282 = n14460 | n14836;
  assign n14838 = pi182 & n14259;
  assign n14839 = pi189 & ~n14501;
  assign n14840 = ~n14838 & n14839;
  assign n14841 = pi182 & n14210;
  assign n14842 = ~pi189 & ~n14841;
  assign n14843 = n14527 & n14842;
  assign n14844 = ~n14840 & ~n14843;
  assign n14845 = n11712 & ~n14844;
  assign n14846 = ~pi189 & ~n14518;
  assign n14847 = pi189 & ~n14515;
  assign n14848 = ~pi182 & ~n14847;
  assign n14849 = ~n14846 & n14848;
  assign n14850 = ~pi189 & ~n14511;
  assign n14851 = pi189 & ~n14504;
  assign n14852 = pi182 & ~n14851;
  assign n14853 = ~n14850 & n14852;
  assign n14854 = ~n14849 & ~n14853;
  assign n14855 = n11750 & ~n14854;
  assign n14856 = ~n14845 & ~n14855;
  assign n14857 = ~n10118 & ~n14198;
  assign n14858 = ~pi166 & n14201;
  assign n14859 = ~n14857 & ~n14858;
  assign n14860 = ~pi153 & ~n14859;
  assign n14861 = ~pi166 & n14204;
  assign n14862 = pi166 & n14230;
  assign n14863 = pi153 & ~n14862;
  assign n14864 = ~n14861 & n14863;
  assign n14865 = ~n14860 & ~n14864;
  assign n14866 = ~pi160 & ~n14865;
  assign n14867 = ~pi166 & ~n14211;
  assign n14868 = pi160 & ~n14867;
  assign n14869 = pi153 & n13989;
  assign n14870 = pi166 & n14259;
  assign n14871 = ~n14869 & ~n14870;
  assign n14872 = n14868 & n14871;
  assign n14873 = ~n14866 & ~n14872;
  assign n14874 = n8959 & n14873;
  assign n14875 = ~n10118 & ~n13993;
  assign n14876 = ~pi51 & ~n14875;
  assign n14877 = ~n14869 & ~n14876;
  assign n14878 = ~n8959 & ~n14877;
  assign n14879 = pi299 & ~n14878;
  assign n14880 = ~n14874 & n14879;
  assign n14881 = n14856 & ~n14880;
  assign n14882 = pi232 & ~n14881;
  assign n14883 = n14545 & ~n14882;
  assign n14884 = ~pi126 & n14010;
  assign n14885 = pi126 & ~n14010;
  assign n14886 = ~n14884 & ~n14885;
  assign n14887 = ~n14006 & ~n14886;
  assign n14888 = ~pi189 & n14637;
  assign n14889 = pi189 & n14635;
  assign n14890 = pi178 & ~n14889;
  assign n14891 = ~n14888 & n14890;
  assign n14892 = pi189 & n14560;
  assign n14893 = ~pi189 & n14567;
  assign n14894 = ~pi178 & ~n14893;
  assign n14895 = ~n14892 & n14894;
  assign n14896 = ~pi181 & ~n14895;
  assign n14897 = ~n14891 & n14896;
  assign n14898 = pi178 & n11725;
  assign n14899 = n14049 & n14898;
  assign n14900 = pi181 & ~n14899;
  assign n14901 = ~pi189 & ~n14098;
  assign n14902 = pi189 & ~n14079;
  assign n14903 = ~pi178 & ~n14902;
  assign n14904 = ~n14901 & n14903;
  assign n14905 = ~n14084 & ~n14904;
  assign n14906 = n14900 & n14905;
  assign n14907 = n11750 & ~n14906;
  assign n14908 = ~n14897 & n14907;
  assign n14909 = ~pi51 & ~n14075;
  assign n14910 = ~n14877 & ~n14909;
  assign n14911 = ~pi153 & ~n14910;
  assign n14912 = ~n14085 & n14911;
  assign n14913 = n11639 & n14049;
  assign n14914 = ~n14084 & ~n14913;
  assign n14915 = pi153 & ~n14914;
  assign n14916 = pi157 & ~n14915;
  assign n14917 = ~n14912 & n14916;
  assign n14918 = pi166 & ~n14557;
  assign n14919 = pi51 & n10118;
  assign n14920 = ~n14918 & ~n14919;
  assign n14921 = ~pi153 & ~n14920;
  assign n14922 = pi153 & pi166;
  assign n14923 = ~n14614 & n14922;
  assign n14924 = ~pi166 & ~n14563;
  assign n14925 = ~pi157 & ~n14924;
  assign n14926 = ~n14923 & n14925;
  assign n14927 = ~n14921 & n14926;
  assign n14928 = ~n14917 & ~n14927;
  assign n14929 = n9693 & n14928;
  assign n14930 = ~n14908 & ~n14929;
  assign n14931 = pi189 & n14557;
  assign n14932 = ~pi189 & n14582;
  assign n14933 = ~n14098 & n14932;
  assign n14934 = ~pi178 & ~n14933;
  assign n14935 = ~n14931 & n14934;
  assign n14936 = pi178 & ~n14085;
  assign n14937 = ~n14932 & n14936;
  assign n14938 = pi181 & ~n14937;
  assign n14939 = ~n14935 & n14938;
  assign n14940 = ~n10122 & ~n14083;
  assign n14941 = ~pi189 & n14309;
  assign n14942 = ~n14940 & ~n14941;
  assign n14943 = ~pi178 & ~n14942;
  assign n14944 = ~pi181 & ~n14943;
  assign n14945 = ~n14891 & ~n14937;
  assign n14946 = n14944 & n14945;
  assign n14947 = ~n14939 & ~n14946;
  assign n14948 = n11712 & n14947;
  assign n14949 = n14930 & ~n14948;
  assign n14950 = ~pi166 & ~n14567;
  assign n14951 = pi166 & ~n14560;
  assign n14952 = pi153 & ~n14951;
  assign n14953 = ~n14950 & n14952;
  assign n14954 = ~n10118 & ~n14083;
  assign n14955 = ~pi153 & ~n14954;
  assign n14956 = ~pi166 & n14309;
  assign n14957 = n14955 & ~n14956;
  assign n14958 = ~n14953 & ~n14957;
  assign n14959 = ~pi157 & ~n14958;
  assign n14960 = ~pi166 & ~n14637;
  assign n14961 = ~n14635 & n14922;
  assign n14962 = pi166 & ~n14588;
  assign n14963 = ~n14919 & ~n14962;
  assign n14964 = ~pi153 & ~n14963;
  assign n14965 = pi157 & ~n14964;
  assign n14966 = ~n14961 & n14965;
  assign n14967 = ~n14960 & n14966;
  assign n14968 = n9659 & ~n14967;
  assign n14969 = ~n14959 & n14968;
  assign n14970 = n14949 & ~n14969;
  assign n14971 = pi232 & ~n14970;
  assign n14972 = n14548 & ~n14971;
  assign n14973 = ~n14887 & ~n14972;
  assign n14974 = ~n14883 & n14973;
  assign n14975 = ~pi153 & n14697;
  assign n14976 = pi153 & n14695;
  assign n14977 = pi157 & ~n14976;
  assign n14978 = ~n14975 & n14977;
  assign n14979 = ~pi153 & n14670;
  assign n14980 = pi153 & ~n14672;
  assign n14981 = ~pi157 & ~n14980;
  assign n14982 = ~n14979 & n14981;
  assign n14983 = ~n14978 & ~n14982;
  assign n14984 = pi166 & ~n14983;
  assign n14985 = pi157 & n14071;
  assign n14986 = ~pi166 & n14664;
  assign n14987 = ~n14869 & n14986;
  assign n14988 = ~n14985 & n14987;
  assign n14989 = ~n14984 & ~n14988;
  assign n14990 = n9693 & ~n14989;
  assign n14991 = pi166 & ~n14679;
  assign n14992 = ~pi166 & n14683;
  assign n14993 = pi153 & ~n14992;
  assign n14994 = ~n14991 & n14993;
  assign n14995 = pi166 & n14687;
  assign n14996 = ~pi166 & ~n14689;
  assign n14997 = ~pi153 & ~n14996;
  assign n14998 = ~n14995 & n14997;
  assign n14999 = ~n14994 & ~n14998;
  assign n15000 = pi157 & ~n14999;
  assign n15001 = ~pi166 & ~n14662;
  assign n15002 = pi166 & n14099;
  assign n15003 = ~pi157 & ~n15002;
  assign n15004 = ~n14869 & n15003;
  assign n15005 = ~n15001 & n15004;
  assign n15006 = ~n15000 & ~n15005;
  assign n15007 = n9659 & ~n15006;
  assign n15008 = pi189 & n14672;
  assign n15009 = ~pi189 & n14664;
  assign n15010 = ~n13989 & n15009;
  assign n15011 = ~n15008 & ~n15010;
  assign n15012 = ~pi178 & ~n15011;
  assign n15013 = ~pi189 & ~n14701;
  assign n15014 = n14695 & ~n14932;
  assign n15015 = ~n15013 & ~n15014;
  assign n15016 = pi178 & n15015;
  assign n15017 = ~n15012 & ~n15016;
  assign n15018 = pi181 & n15017;
  assign n15019 = ~pi189 & ~n14662;
  assign n15020 = pi189 & n14099;
  assign n15021 = ~pi178 & ~n15020;
  assign n15022 = ~n15019 & n15021;
  assign n15023 = ~n13989 & n15022;
  assign n15024 = ~pi181 & ~n15023;
  assign n15025 = pi189 & ~n14679;
  assign n15026 = ~pi189 & n14683;
  assign n15027 = ~n15025 & ~n15026;
  assign n15028 = pi178 & n15027;
  assign n15029 = n15024 & ~n15028;
  assign n15030 = n11750 & ~n15029;
  assign n15031 = ~n15018 & n15030;
  assign n15032 = ~n15007 & ~n15031;
  assign n15033 = ~n14990 & n15032;
  assign n15034 = pi189 & n14697;
  assign n15035 = ~n15013 & ~n15034;
  assign n15036 = pi178 & ~n15035;
  assign n15037 = pi189 & ~n14670;
  assign n15038 = ~pi178 & ~n15009;
  assign n15039 = ~n15037 & n15038;
  assign n15040 = ~n15036 & ~n15039;
  assign n15041 = pi181 & ~n15040;
  assign n15042 = n14662 & n15021;
  assign n15043 = pi189 & n14687;
  assign n15044 = ~pi189 & ~n14689;
  assign n15045 = pi178 & ~n15044;
  assign n15046 = ~n15043 & n15045;
  assign n15047 = n15024 & ~n15046;
  assign n15048 = ~n15042 & n15047;
  assign n15049 = n11712 & ~n15048;
  assign n15050 = ~n15041 & n15049;
  assign n15051 = n15033 & ~n15050;
  assign n15052 = pi232 & ~n15051;
  assign n15053 = n14826 & ~n15052;
  assign n15054 = ~pi189 & n14813;
  assign n15055 = pi189 & n14815;
  assign n15056 = ~pi182 & ~n15055;
  assign n15057 = ~n15054 & n15056;
  assign n15058 = ~n13989 & n15057;
  assign n15059 = pi189 & ~n14791;
  assign n15060 = ~pi189 & n14797;
  assign n15061 = pi182 & ~n15060;
  assign n15062 = ~n15059 & n15061;
  assign n15063 = ~n15058 & ~n15062;
  assign n15064 = n11750 & ~n15063;
  assign n15065 = ~pi189 & n14803;
  assign n15066 = pi189 & n14806;
  assign n15067 = ~n15065 & ~n15066;
  assign n15068 = pi182 & n15067;
  assign n15069 = ~n15057 & ~n15068;
  assign n15070 = n11712 & ~n15069;
  assign n15071 = ~n15064 & ~n15070;
  assign n15072 = pi166 & ~n14759;
  assign n15073 = ~pi166 & n14757;
  assign n15074 = pi51 & ~pi153;
  assign n15075 = ~n15073 & ~n15074;
  assign n15076 = ~n15072 & n15075;
  assign n15077 = ~pi216 & ~n15076;
  assign n15078 = ~pi166 & n14224;
  assign n15079 = ~pi153 & ~n15078;
  assign n15080 = n6440 & n11639;
  assign n15081 = n15079 & ~n15080;
  assign n15082 = pi166 & ~n14774;
  assign n15083 = ~pi166 & ~n14770;
  assign n15084 = pi153 & ~n15083;
  assign n15085 = ~n15082 & n15084;
  assign n15086 = pi160 & ~n15085;
  assign n15087 = ~n15081 & n15086;
  assign n15088 = pi216 & ~n15087;
  assign n15089 = ~n15077 & ~n15088;
  assign n15090 = n5744 & n15089;
  assign n15091 = ~pi160 & pi216;
  assign n15092 = n5744 & ~n15091;
  assign n15093 = n14910 & ~n15092;
  assign n15094 = pi299 & ~n15093;
  assign n15095 = ~n15090 & n15094;
  assign n15096 = n15071 & ~n15095;
  assign n15097 = pi232 & ~n15096;
  assign n15098 = n14753 & ~n15097;
  assign n15099 = n14887 & ~n15098;
  assign n15100 = ~n15053 & n15099;
  assign n15101 = n2614 & ~n15100;
  assign n15102 = ~n14974 & n15101;
  assign n15103 = pi299 & ~n14910;
  assign n15104 = n10122 & n14049;
  assign n15105 = pi175 & n13989;
  assign n15106 = ~pi299 & ~n15105;
  assign n15107 = ~n15104 & n15106;
  assign n15108 = pi232 & ~n15107;
  assign n15109 = ~n15103 & n15108;
  assign n15110 = n13994 & ~n14887;
  assign n15111 = ~n15109 & ~n15110;
  assign n15112 = ~n2614 & ~n15111;
  assign n15113 = ~n15102 & ~n15112;
  assign n15114 = n2537 & n15113;
  assign n15115 = n14021 & ~n15109;
  assign n15116 = ~pi150 & pi299;
  assign n15117 = ~pi185 & ~pi299;
  assign n15118 = ~n15116 & ~n15117;
  assign n15119 = n7420 & n15118;
  assign n15120 = pi87 & ~n15119;
  assign n15121 = ~n15115 & ~n15120;
  assign n15122 = n14013 & ~n14887;
  assign n15123 = ~n15121 & ~n15122;
  assign n15124 = ~po1038 & ~n15123;
  assign n15125 = ~n15114 & n15124;
  assign n15126 = pi232 & n14910;
  assign n15127 = ~n15110 & ~n15126;
  assign n15128 = ~pi87 & n15127;
  assign n15129 = pi87 & ~n13475;
  assign n15130 = po1038 & ~n15129;
  assign n15131 = ~n15128 & n15130;
  assign po283 = ~n15125 & ~n15131;
  assign n15133 = n2539 & n8743;
  assign n15134 = ~n2531 & ~n15133;
  assign n15135 = pi54 & n3275;
  assign n15136 = n8743 & n15135;
  assign n15137 = pi92 & ~pi129;
  assign n15138 = ~pi54 & ~n7258;
  assign n15139 = pi129 & n7252;
  assign n15140 = pi75 & n15139;
  assign n15141 = ~n2615 & ~n8820;
  assign n15142 = n8743 & ~n15141;
  assign n15143 = ~n2571 & ~n15142;
  assign n15144 = pi129 & n6132;
  assign n15145 = pi38 & ~n15144;
  assign n15146 = pi39 & n8743;
  assign n15147 = ~pi38 & ~n15146;
  assign n15148 = ~n2717 & ~n3043;
  assign n15149 = n2779 & ~n2852;
  assign n15150 = n2463 & ~n15149;
  assign n15151 = n2865 & ~n15150;
  assign n15152 = n2776 & ~n15151;
  assign n15153 = n2869 & ~n15152;
  assign n15154 = n2705 & ~n15153;
  assign n15155 = ~n2708 & ~n15154;
  assign n15156 = ~pi86 & ~n15155;
  assign n15157 = n2774 & ~n15156;
  assign n15158 = n2772 & ~n15157;
  assign n15159 = ~n2769 & ~n15158;
  assign n15160 = ~pi108 & ~n15159;
  assign n15161 = n2768 & ~n15160;
  assign n15162 = n2881 & ~n15161;
  assign n15163 = ~n2759 & ~n15162;
  assign n15164 = n2758 & ~n15163;
  assign n15165 = n2757 & ~n15164;
  assign n15166 = ~po740 & n15165;
  assign n15167 = ~pi97 & ~n15157;
  assign n15168 = ~n2769 & ~n15167;
  assign n15169 = ~pi108 & ~n15168;
  assign n15170 = n2768 & ~n15169;
  assign n15171 = n2881 & ~n15170;
  assign n15172 = ~n2759 & ~n15171;
  assign n15173 = n2758 & ~n15172;
  assign n15174 = n2757 & ~n15173;
  assign n15175 = po740 & n15174;
  assign n15176 = pi250 & ~n7421;
  assign n15177 = n9905 & n15176;
  assign n15178 = ~n15175 & n15177;
  assign n15179 = ~n15166 & n15178;
  assign n15180 = pi127 & n15165;
  assign n15181 = ~pi127 & n15174;
  assign n15182 = ~n15177 & ~n15181;
  assign n15183 = ~n15180 & n15182;
  assign n15184 = ~n15179 & ~n15183;
  assign n15185 = n2750 & ~n15184;
  assign n15186 = n3045 & ~n15185;
  assign n15187 = n2519 & ~n15186;
  assign n15188 = n15148 & ~n15187;
  assign n15189 = ~pi70 & ~n15188;
  assign n15190 = ~n3062 & ~n15189;
  assign n15191 = ~pi51 & ~n15190;
  assign n15192 = n2743 & ~n15191;
  assign n15193 = n3065 & ~n15192;
  assign n15194 = ~n2739 & ~n15193;
  assign n15195 = n2461 & ~n15194;
  assign n15196 = n3377 & ~n15195;
  assign n15197 = ~pi95 & ~n15196;
  assign n15198 = pi129 & ~n15197;
  assign n15199 = ~pi39 & n15198;
  assign n15200 = ~n2907 & n15199;
  assign n15201 = n15147 & ~n15200;
  assign n15202 = ~n15145 & ~n15201;
  assign n15203 = n2571 & ~n15202;
  assign n15204 = ~pi75 & ~n15203;
  assign n15205 = ~n15143 & n15204;
  assign n15206 = ~pi92 & ~n15205;
  assign n15207 = ~n15140 & n15206;
  assign n15208 = n15138 & ~n15207;
  assign n15209 = ~n15137 & n15208;
  assign n15210 = ~pi74 & ~n15209;
  assign n15211 = ~n15136 & n15210;
  assign n15212 = n6525 & n15139;
  assign n15213 = pi74 & ~n15212;
  assign n15214 = ~pi55 & ~n15213;
  assign n15215 = ~n15211 & n15214;
  assign n15216 = pi55 & n7309;
  assign n15217 = n15139 & n15216;
  assign n15218 = ~n15215 & ~n15217;
  assign n15219 = ~pi56 & ~n15218;
  assign n15220 = ~n11092 & ~n11101;
  assign n15221 = ~n15219 & n15220;
  assign n15222 = ~n15134 & ~n15221;
  assign n15223 = n3327 & ~n15222;
  assign n15224 = ~pi129 & ~n3327;
  assign n15225 = n6087 & ~n15224;
  assign po284 = ~n15223 & n15225;
  assign n15227 = ~pi38 & ~n3382;
  assign n15228 = n6134 & ~n15227;
  assign n15229 = n6489 & n8740;
  assign n15230 = ~pi87 & ~n15229;
  assign n15231 = ~n15228 & n15230;
  assign n15232 = n6096 & ~n15231;
  assign n15233 = n8744 & n10180;
  assign n15234 = ~pi129 & ~n15233;
  assign n15235 = n8822 & ~n15234;
  assign n15236 = po740 & n15233;
  assign n15237 = n2522 & ~n15236;
  assign n15238 = n15235 & n15237;
  assign n15239 = n6094 & ~n15238;
  assign n15240 = ~n15232 & n15239;
  assign n15241 = ~n7295 & ~n15240;
  assign n15242 = ~n7258 & n15241;
  assign n15243 = n6262 & ~n15242;
  assign n15244 = n7251 & ~n15243;
  assign n15245 = ~pi56 & ~n15244;
  assign n15246 = ~n6264 & ~n15245;
  assign n15247 = ~pi62 & ~n15246;
  assign n15248 = ~n6268 & ~n15247;
  assign n15249 = n3327 & ~n15248;
  assign po286 = n6087 & ~n15249;
  assign n15251 = pi87 & ~n9592;
  assign n15252 = n7420 & ~n8918;
  assign n15253 = n14049 & ~n15252;
  assign n15254 = ~n14909 & ~n15253;
  assign n15255 = n14021 & ~n15254;
  assign n15256 = ~n15251 & ~n15255;
  assign n15257 = ~n14013 & ~n15256;
  assign n15258 = ~pi132 & n14884;
  assign n15259 = pi130 & ~n15258;
  assign n15260 = ~pi130 & n15258;
  assign n15261 = ~n15259 & ~n15260;
  assign n15262 = ~n14004 & ~n15261;
  assign n15263 = ~n15257 & ~n15262;
  assign n15264 = pi100 & n15254;
  assign n15265 = ~n10779 & n15253;
  assign n15266 = ~pi51 & ~n14543;
  assign n15267 = ~pi232 & ~n15266;
  assign n15268 = n10779 & ~n15267;
  assign n15269 = ~pi191 & ~pi299;
  assign n15270 = ~pi51 & ~n14501;
  assign n15271 = pi140 & n14503;
  assign n15272 = n15270 & ~n15271;
  assign n15273 = n15269 & ~n15272;
  assign n15274 = ~pi51 & n14527;
  assign n15275 = pi140 & n14209;
  assign n15276 = n15274 & ~n15275;
  assign n15277 = n8916 & ~n15276;
  assign n15278 = ~n15273 & ~n15277;
  assign n15279 = ~pi169 & ~n14502;
  assign n15280 = ~n14209 & n14525;
  assign n15281 = pi169 & ~n15280;
  assign n15282 = pi162 & n8959;
  assign n15283 = ~n15281 & n15282;
  assign n15284 = ~n15279 & n15283;
  assign n15285 = pi169 & n6190;
  assign n15286 = ~n8959 & n14049;
  assign n15287 = ~n15285 & n15286;
  assign n15288 = ~n14221 & ~n15285;
  assign n15289 = ~pi162 & ~n15288;
  assign n15290 = n4856 & n6190;
  assign n15291 = n8959 & ~n15290;
  assign n15292 = n15289 & n15291;
  assign n15293 = pi299 & ~n15292;
  assign n15294 = ~n15287 & n15293;
  assign n15295 = ~n15284 & n15294;
  assign n15296 = n15278 & ~n15295;
  assign n15297 = pi232 & ~n15296;
  assign n15298 = n15268 & ~n15297;
  assign n15299 = ~pi100 & ~n15298;
  assign n15300 = ~n15265 & n15299;
  assign n15301 = ~n15264 & ~n15300;
  assign n15302 = n14475 & n15301;
  assign n15303 = n15263 & ~n15302;
  assign n15304 = ~n2614 & n15254;
  assign n15305 = ~n14200 & ~n15285;
  assign n15306 = pi169 & n14756;
  assign n15307 = ~n15305 & ~n15306;
  assign n15308 = ~pi216 & ~n15307;
  assign n15309 = pi162 & pi216;
  assign n15310 = ~pi51 & ~n14773;
  assign n15311 = ~pi169 & n15310;
  assign n15312 = n15309 & ~n15311;
  assign n15313 = ~n14229 & n14770;
  assign n15314 = pi169 & n15313;
  assign n15315 = n15312 & ~n15314;
  assign n15316 = ~n15308 & ~n15315;
  assign n15317 = n5744 & ~n15316;
  assign n15318 = pi169 & n14075;
  assign n15319 = ~pi51 & ~n15318;
  assign n15320 = ~n5745 & ~n15282;
  assign n15321 = ~n15319 & n15320;
  assign n15322 = ~n15317 & ~n15321;
  assign n15323 = pi299 & ~n15322;
  assign n15324 = n2521 & n14788;
  assign n15325 = ~pi51 & ~n15324;
  assign n15326 = pi140 & n15325;
  assign n15327 = ~pi51 & ~n14815;
  assign n15328 = ~pi140 & n15327;
  assign n15329 = n15269 & ~n15328;
  assign n15330 = ~n15326 & n15329;
  assign n15331 = ~n15323 & ~n15330;
  assign n15332 = ~pi51 & ~n14803;
  assign n15333 = pi140 & n15332;
  assign n15334 = ~pi51 & ~n14813;
  assign n15335 = ~pi140 & n15334;
  assign n15336 = n8916 & ~n15335;
  assign n15337 = ~n15333 & n15336;
  assign n15338 = n15331 & ~n15337;
  assign n15339 = pi232 & ~n15338;
  assign n15340 = ~pi51 & ~n14751;
  assign n15341 = ~pi232 & ~n15340;
  assign n15342 = pi39 & ~n15341;
  assign n15343 = ~n15339 & n15342;
  assign n15344 = ~pi232 & ~n14116;
  assign n15345 = ~pi39 & ~n15344;
  assign n15346 = n6190 & n14068;
  assign n15347 = ~n6190 & n14116;
  assign n15348 = ~n15346 & ~n15347;
  assign n15349 = ~n8918 & ~n15348;
  assign n15350 = n8918 & n14116;
  assign n15351 = ~n15349 & ~n15350;
  assign n15352 = pi232 & n15351;
  assign n15353 = n15345 & ~n15352;
  assign n15354 = ~n15343 & ~n15353;
  assign n15355 = n2614 & n15354;
  assign n15356 = ~n15304 & ~n15355;
  assign n15357 = n2537 & n15356;
  assign n15358 = n15256 & ~n15357;
  assign n15359 = n15262 & n15358;
  assign n15360 = ~n15303 & ~n15359;
  assign n15361 = ~po1038 & ~n15360;
  assign n15362 = pi87 & ~n9765;
  assign n15363 = po1038 & ~n15362;
  assign n15364 = ~pi51 & ~pi87;
  assign n15365 = ~n8844 & ~n13993;
  assign n15366 = n15364 & n15365;
  assign n15367 = n15363 & ~n15366;
  assign n15368 = ~n15318 & n15364;
  assign n15369 = n15262 & n15368;
  assign n15370 = n15367 & ~n15369;
  assign po287 = ~n15361 & ~n15370;
  assign n15372 = ~pi100 & ~n13651;
  assign n15373 = n7262 & ~n15372;
  assign n15374 = ~pi75 & ~n15373;
  assign n15375 = ~n7253 & ~n15374;
  assign n15376 = ~pi92 & ~n15375;
  assign n15377 = n8738 & n15138;
  assign po288 = ~n15376 & n15377;
  assign n15379 = pi51 & ~pi151;
  assign n15380 = ~n13411 & ~n13989;
  assign n15381 = ~n15379 & ~n15380;
  assign n15382 = n13995 & n15381;
  assign n15383 = pi232 & n15382;
  assign n15384 = pi132 & ~n14884;
  assign n15385 = ~n15258 & ~n15384;
  assign n15386 = ~n14005 & ~n15385;
  assign n15387 = n13994 & ~n15386;
  assign n15388 = ~n15383 & ~n15387;
  assign n15389 = ~pi87 & ~n15388;
  assign n15390 = po1038 & ~n15389;
  assign n15391 = pi164 & n14446;
  assign n15392 = n15390 & ~n15391;
  assign n15393 = pi299 & ~n15382;
  assign n15394 = pi190 & n14075;
  assign n15395 = pi173 & n13989;
  assign n15396 = ~pi299 & ~n15395;
  assign n15397 = ~n15394 & n15396;
  assign n15398 = pi232 & ~n15397;
  assign n15399 = ~n15393 & n15398;
  assign n15400 = n14021 & ~n15399;
  assign n15401 = ~n13994 & n15400;
  assign n15402 = pi87 & ~n8926;
  assign n15403 = ~n2614 & n15399;
  assign n15404 = n2537 & ~n15403;
  assign n15405 = ~n2614 & n13994;
  assign n15406 = pi190 & ~pi299;
  assign n15407 = ~pi183 & ~n14518;
  assign n15408 = pi183 & ~n14511;
  assign n15409 = pi173 & ~n15408;
  assign n15410 = ~n15407 & n15409;
  assign n15411 = pi183 & n14210;
  assign n15412 = ~pi173 & ~n15411;
  assign n15413 = n14527 & n15412;
  assign n15414 = ~n15410 & ~n15413;
  assign n15415 = n15406 & ~n15414;
  assign n15416 = ~n13994 & n15393;
  assign n15417 = ~n12812 & ~n15416;
  assign n15418 = ~pi168 & ~n14230;
  assign n15419 = pi168 & ~n14204;
  assign n15420 = ~n15418 & ~n15419;
  assign n15421 = pi151 & n15420;
  assign n15422 = pi168 & n14201;
  assign n15423 = ~n13411 & ~n14198;
  assign n15424 = ~pi151 & ~n15423;
  assign n15425 = ~n15422 & n15424;
  assign n15426 = ~pi149 & ~n15425;
  assign n15427 = ~n15421 & n15426;
  assign n15428 = n6190 & n15379;
  assign n15429 = pi168 & ~n15428;
  assign n15430 = n14509 & n15429;
  assign n15431 = ~n14259 & ~n15381;
  assign n15432 = ~pi168 & ~n15431;
  assign n15433 = pi149 & ~n15432;
  assign n15434 = ~n15430 & n15433;
  assign n15435 = n8959 & ~n15434;
  assign n15436 = ~n15427 & n15435;
  assign n15437 = ~n15417 & ~n15436;
  assign n15438 = pi183 & n14259;
  assign n15439 = ~pi190 & ~pi299;
  assign n15440 = ~n15395 & n15439;
  assign n15441 = ~n14501 & n15440;
  assign n15442 = ~n15438 & n15441;
  assign n15443 = ~n15437 & ~n15442;
  assign n15444 = ~n15415 & n15443;
  assign n15445 = pi232 & ~n15444;
  assign n15446 = ~n14544 & ~n15445;
  assign n15447 = pi39 & ~n15446;
  assign n15448 = ~pi232 & n14082;
  assign n15449 = pi151 & n14336;
  assign n15450 = ~pi151 & ~n14082;
  assign n15451 = ~pi168 & ~n15450;
  assign n15452 = ~n15449 & n15451;
  assign n15453 = ~n14142 & n15429;
  assign n15454 = ~n15452 & ~n15453;
  assign n15455 = ~pi160 & ~n15454;
  assign n15456 = ~n14555 & n15455;
  assign n15457 = ~pi151 & ~n15382;
  assign n15458 = ~n14556 & n15457;
  assign n15459 = ~pi168 & n14075;
  assign n15460 = ~n14555 & ~n15459;
  assign n15461 = pi151 & ~n15460;
  assign n15462 = pi160 & ~n15461;
  assign n15463 = ~n15458 & n15462;
  assign n15464 = pi299 & ~n15463;
  assign n15465 = ~n15456 & n15464;
  assign n15466 = ~pi182 & n14142;
  assign n15467 = pi51 & ~pi173;
  assign n15468 = ~n14555 & ~n15467;
  assign n15469 = ~n15466 & n15468;
  assign n15470 = n15406 & ~n15469;
  assign n15471 = pi232 & ~n15470;
  assign n15472 = pi182 & n14556;
  assign n15473 = ~n14082 & n15440;
  assign n15474 = ~n15472 & n15473;
  assign n15475 = n15471 & ~n15474;
  assign n15476 = ~n15465 & n15475;
  assign n15477 = ~pi39 & ~n15476;
  assign n15478 = ~n15448 & n15477;
  assign n15479 = ~n15447 & ~n15478;
  assign n15480 = n2614 & n15479;
  assign n15481 = ~n15405 & ~n15480;
  assign n15482 = n15404 & n15481;
  assign n15483 = ~n15386 & ~n15482;
  assign n15484 = ~n15402 & n15483;
  assign n15485 = ~n15401 & n15484;
  assign n15486 = ~po1038 & ~n15485;
  assign n15487 = ~pi182 & n14094;
  assign n15488 = ~pi173 & ~n15487;
  assign n15489 = ~n6190 & ~n14094;
  assign n15490 = ~n14123 & ~n15489;
  assign n15491 = pi182 & n15490;
  assign n15492 = n15488 & ~n15491;
  assign n15493 = ~n6190 & n14094;
  assign n15494 = ~n14117 & ~n15493;
  assign n15495 = pi182 & ~n15494;
  assign n15496 = n14679 & ~n15493;
  assign n15497 = ~pi182 & ~n15496;
  assign n15498 = pi173 & ~n15497;
  assign n15499 = ~n15495 & n15498;
  assign n15500 = ~n15492 & ~n15499;
  assign n15501 = n15439 & ~n15500;
  assign n15502 = ~pi168 & ~n15496;
  assign n15503 = ~n14682 & ~n15489;
  assign n15504 = pi168 & n15503;
  assign n15505 = ~n15502 & ~n15504;
  assign n15506 = pi151 & n15505;
  assign n15507 = pi168 & n14071;
  assign n15508 = ~n13411 & n14094;
  assign n15509 = ~pi151 & ~n15508;
  assign n15510 = ~n15507 & n15509;
  assign n15511 = ~pi160 & ~n15510;
  assign n15512 = ~n15506 & n15511;
  assign n15513 = pi168 & ~n15379;
  assign n15514 = ~n14068 & n15513;
  assign n15515 = pi151 & n14116;
  assign n15516 = ~pi151 & ~n14122;
  assign n15517 = ~pi168 & ~n15516;
  assign n15518 = ~n15515 & n15517;
  assign n15519 = n6190 & ~n15518;
  assign n15520 = ~n15514 & n15519;
  assign n15521 = ~n15489 & ~n15520;
  assign n15522 = pi160 & n15521;
  assign n15523 = ~n15512 & ~n15522;
  assign n15524 = pi299 & n15523;
  assign n15525 = pi182 & n14048;
  assign n15526 = n14067 & ~n15525;
  assign n15527 = ~n15467 & ~n15526;
  assign n15528 = n6190 & n15527;
  assign n15529 = n15406 & ~n15493;
  assign n15530 = ~n15528 & n15529;
  assign n15531 = pi232 & ~n15530;
  assign n15532 = ~n15524 & n15531;
  assign n15533 = ~n15501 & n15532;
  assign n15534 = ~pi232 & n14094;
  assign n15535 = ~n15533 & ~n15534;
  assign n15536 = ~pi39 & ~n15535;
  assign n15537 = pi183 & n14796;
  assign n15538 = ~n14793 & ~n15537;
  assign n15539 = pi173 & ~n15538;
  assign n15540 = ~n14802 & ~n15537;
  assign n15541 = ~pi173 & ~n15540;
  assign n15542 = ~n15539 & ~n15541;
  assign n15543 = ~pi183 & ~n7529;
  assign n15544 = ~n13995 & n15543;
  assign n15545 = n15542 & ~n15544;
  assign n15546 = n15406 & ~n15545;
  assign n15547 = ~n14229 & ~n15327;
  assign n15548 = ~pi183 & ~n15547;
  assign n15549 = pi183 & n14791;
  assign n15550 = ~n15548 & ~n15549;
  assign n15551 = pi173 & n15550;
  assign n15552 = ~pi173 & n14806;
  assign n15553 = ~n15543 & n15552;
  assign n15554 = n15439 & ~n15553;
  assign n15555 = ~n15551 & n15554;
  assign n15556 = ~n15546 & ~n15555;
  assign n15557 = pi168 & n14224;
  assign n15558 = ~pi168 & n14287;
  assign n15559 = ~pi151 & ~n15558;
  assign n15560 = ~n15557 & n15559;
  assign n15561 = ~pi168 & ~n14774;
  assign n15562 = pi168 & ~n14770;
  assign n15563 = pi151 & ~n15562;
  assign n15564 = ~n15561 & n15563;
  assign n15565 = pi149 & ~n15564;
  assign n15566 = ~n15560 & n15565;
  assign n15567 = pi216 & ~n15566;
  assign n15568 = ~pi168 & ~n14759;
  assign n15569 = pi168 & n14757;
  assign n15570 = ~n15379 & ~n15569;
  assign n15571 = ~n15568 & n15570;
  assign n15572 = ~pi216 & ~n15571;
  assign n15573 = ~n15567 & ~n15572;
  assign n15574 = n5744 & n15573;
  assign n15575 = ~pi149 & pi216;
  assign n15576 = n5744 & ~n15575;
  assign n15577 = n15382 & ~n15576;
  assign n15578 = pi299 & ~n15577;
  assign n15579 = ~n15574 & n15578;
  assign n15580 = n15556 & ~n15579;
  assign n15581 = pi232 & ~n15580;
  assign n15582 = n14753 & ~n15581;
  assign n15583 = ~n15536 & ~n15582;
  assign n15584 = n2614 & ~n15583;
  assign n15585 = n15404 & ~n15584;
  assign n15586 = ~n15402 & ~n15585;
  assign n15587 = ~n15400 & n15586;
  assign n15588 = n15386 & n15587;
  assign n15589 = n15486 & ~n15588;
  assign po289 = n15392 | n15589;
  assign n15591 = ~pi133 & ~n14448;
  assign n15592 = ~n13994 & n14021;
  assign n15593 = pi145 & n14259;
  assign n15594 = n14539 & ~n15593;
  assign n15595 = pi197 & n14209;
  assign n15596 = n14540 & ~n15595;
  assign n15597 = n13994 & ~n15596;
  assign n15598 = pi299 & ~n15597;
  assign n15599 = ~n15594 & ~n15598;
  assign n15600 = pi232 & ~n15599;
  assign n15601 = n14545 & ~n15600;
  assign n15602 = ~n8938 & n14060;
  assign n15603 = ~pi39 & ~n15602;
  assign n15604 = n13994 & n15603;
  assign n15605 = ~pi38 & ~n15604;
  assign n15606 = ~n15601 & n15605;
  assign n15607 = n14038 & ~n15606;
  assign n15608 = n14475 & ~n15607;
  assign n15609 = ~n15592 & ~n15608;
  assign n15610 = ~n15591 & ~n15609;
  assign n15611 = ~pi183 & ~pi299;
  assign n15612 = ~pi149 & pi299;
  assign n15613 = ~n15611 & ~n15612;
  assign n15614 = n7420 & n15613;
  assign n15615 = pi87 & ~n15614;
  assign n15616 = ~n15610 & ~n15615;
  assign n15617 = ~n6190 & ~n14138;
  assign n15618 = n8935 & ~n15617;
  assign n15619 = ~n14123 & n15618;
  assign n15620 = pi299 & n15619;
  assign n15621 = pi299 & n8935;
  assign n15622 = n14138 & ~n15621;
  assign n15623 = ~pi39 & ~n15622;
  assign n15624 = ~pi176 & n15623;
  assign n15625 = ~n15620 & n15624;
  assign n15626 = ~n5742 & ~n15595;
  assign n15627 = n6592 & ~n15626;
  assign n15628 = ~pi145 & ~n7529;
  assign n15629 = ~pi299 & ~n15628;
  assign n15630 = ~n14805 & n15629;
  assign n15631 = ~n15627 & ~n15630;
  assign n15632 = n2522 & ~n15631;
  assign n15633 = pi232 & ~n15632;
  assign n15634 = ~n14752 & ~n15633;
  assign n15635 = pi39 & ~n15634;
  assign n15636 = n11163 & ~n15635;
  assign n15637 = ~n8935 & n14138;
  assign n15638 = ~pi39 & ~n15637;
  assign n15639 = ~n15619 & n15638;
  assign n15640 = pi176 & n15639;
  assign n15641 = n15636 & ~n15640;
  assign n15642 = ~n15625 & n15641;
  assign n15643 = ~pi87 & n15591;
  assign n15644 = ~n15642 & n15643;
  assign n15645 = n15616 & ~n15644;
  assign n15646 = ~po1038 & ~n15645;
  assign n15647 = n14013 & ~n15591;
  assign n15648 = po1038 & ~n15647;
  assign n15649 = pi87 & n8880;
  assign n15650 = n15648 & ~n15649;
  assign po290 = n15646 | n15650;
  assign n15652 = po1038 & n15364;
  assign n15653 = pi171 & n6190;
  assign n15654 = ~n13993 & n15653;
  assign n15655 = pi232 & n15654;
  assign n15656 = ~pi136 & n15260;
  assign n15657 = ~pi135 & n15656;
  assign n15658 = pi134 & ~n15657;
  assign n15659 = n13993 & ~n15658;
  assign n15660 = ~n15655 & ~n15659;
  assign n15661 = n15652 & n15660;
  assign n15662 = pi192 & ~pi299;
  assign n15663 = pi171 & pi299;
  assign n15664 = ~n15662 & ~n15663;
  assign n15665 = n7420 & ~n15664;
  assign n15666 = n14049 & ~n15665;
  assign n15667 = ~n14909 & ~n15666;
  assign n15668 = ~n2614 & n15667;
  assign n15669 = n2537 & ~n15668;
  assign n15670 = ~pi51 & ~n15654;
  assign n15671 = ~pi164 & pi216;
  assign n15672 = n5744 & ~n15671;
  assign n15673 = ~n15670 & ~n15672;
  assign n15674 = ~n14200 & ~n15653;
  assign n15675 = pi171 & n14756;
  assign n15676 = ~n15674 & ~n15675;
  assign n15677 = ~pi216 & ~n15676;
  assign n15678 = ~pi171 & n15310;
  assign n15679 = pi171 & n15313;
  assign n15680 = pi164 & ~n15679;
  assign n15681 = pi216 & n15680;
  assign n15682 = ~n15678 & n15681;
  assign n15683 = ~n15677 & ~n15682;
  assign n15684 = n5744 & ~n15683;
  assign n15685 = ~n15673 & ~n15684;
  assign n15686 = pi299 & ~n15685;
  assign n15687 = ~n15334 & n15662;
  assign n15688 = ~pi192 & ~pi299;
  assign n15689 = ~n15327 & n15688;
  assign n15690 = pi39 & pi186;
  assign n15691 = ~n15689 & ~n15690;
  assign n15692 = ~n15687 & n15691;
  assign n15693 = ~n15332 & n15662;
  assign n15694 = ~n15325 & n15688;
  assign n15695 = pi186 & ~n15694;
  assign n15696 = ~n15693 & n15695;
  assign n15697 = ~n15692 & ~n15696;
  assign n15698 = ~n15686 & ~n15697;
  assign n15699 = pi232 & ~n15698;
  assign n15700 = n15342 & ~n15699;
  assign n15701 = pi232 & ~n15664;
  assign n15702 = n15348 & n15701;
  assign n15703 = ~n14116 & ~n15701;
  assign n15704 = ~pi39 & ~n15703;
  assign n15705 = ~n15702 & n15704;
  assign n15706 = ~n15700 & ~n15705;
  assign n15707 = n2614 & n15706;
  assign n15708 = n15669 & ~n15707;
  assign n15709 = n14021 & ~n15667;
  assign n15710 = n15658 & ~n15709;
  assign n15711 = ~n15708 & n15710;
  assign n15712 = n14021 & n15666;
  assign n15713 = pi39 & ~pi186;
  assign n15714 = ~n15274 & n15662;
  assign n15715 = ~n15270 & n15688;
  assign n15716 = ~n15714 & ~n15715;
  assign n15717 = n15286 & ~n15653;
  assign n15718 = pi299 & ~n15717;
  assign n15719 = ~n14221 & ~n15653;
  assign n15720 = n4184 & n6190;
  assign n15721 = ~n15719 & ~n15720;
  assign n15722 = n8959 & n15721;
  assign n15723 = n15718 & ~n15722;
  assign n15724 = n15716 & ~n15723;
  assign n15725 = pi232 & ~n15724;
  assign n15726 = ~n15267 & ~n15725;
  assign n15727 = n15713 & ~n15726;
  assign n15728 = ~pi164 & ~n15727;
  assign n15729 = ~pi39 & ~n15666;
  assign n15730 = ~n14209 & n15274;
  assign n15731 = n15662 & ~n15730;
  assign n15732 = ~n14503 & n15270;
  assign n15733 = n15688 & ~n15732;
  assign n15734 = ~n15731 & ~n15733;
  assign n15735 = ~n15723 & n15734;
  assign n15736 = pi232 & ~n15735;
  assign n15737 = ~n15267 & ~n15736;
  assign n15738 = n15690 & ~n15737;
  assign n15739 = ~n15729 & ~n15738;
  assign n15740 = n15728 & n15739;
  assign n15741 = pi171 & ~n15280;
  assign n15742 = ~pi171 & ~n14502;
  assign n15743 = ~n15741 & ~n15742;
  assign n15744 = n8959 & n15743;
  assign n15745 = n15718 & ~n15744;
  assign n15746 = n15734 & ~n15745;
  assign n15747 = pi232 & ~n15746;
  assign n15748 = ~n15267 & ~n15747;
  assign n15749 = n15690 & ~n15748;
  assign n15750 = n15716 & ~n15745;
  assign n15751 = pi232 & ~n15750;
  assign n15752 = ~n15267 & ~n15751;
  assign n15753 = n15713 & ~n15752;
  assign n15754 = pi164 & ~n15753;
  assign n15755 = ~n15749 & n15754;
  assign n15756 = ~n15729 & n15755;
  assign n15757 = ~n15740 & ~n15756;
  assign n15758 = n2614 & n15757;
  assign n15759 = ~n15405 & ~n15758;
  assign n15760 = n15669 & n15759;
  assign n15761 = ~n15658 & ~n15760;
  assign n15762 = ~n15712 & n15761;
  assign n15763 = ~n15711 & ~n15762;
  assign n15764 = ~po1038 & n15763;
  assign po291 = n15661 | n15764;
  assign n15766 = pi170 & n6190;
  assign n15767 = n10392 & n15766;
  assign n15768 = n14049 & ~n15767;
  assign n15769 = pi194 & n8924;
  assign n15770 = n15768 & ~n15769;
  assign n15771 = ~n14909 & ~n15770;
  assign n15772 = pi100 & n15771;
  assign n15773 = pi185 & n14503;
  assign n15774 = n15270 & ~n15773;
  assign n15775 = ~n10779 & n15768;
  assign n15776 = ~pi194 & ~n15775;
  assign n15777 = ~n15774 & n15776;
  assign n15778 = ~pi185 & n15274;
  assign n15779 = pi170 & n7420;
  assign n15780 = ~n8924 & ~n15779;
  assign n15781 = n14049 & n15780;
  assign n15782 = ~n10779 & n15781;
  assign n15783 = pi194 & ~n15782;
  assign n15784 = ~n15730 & n15783;
  assign n15785 = ~n15778 & n15784;
  assign n15786 = ~n15777 & ~n15785;
  assign n15787 = ~pi299 & ~n15786;
  assign n15788 = n15286 & ~n15766;
  assign n15789 = ~n15776 & ~n15783;
  assign n15790 = pi150 & pi299;
  assign n15791 = pi170 & ~n15280;
  assign n15792 = ~pi170 & ~n14502;
  assign n15793 = ~n15791 & ~n15792;
  assign n15794 = n8959 & n15793;
  assign n15795 = n15790 & ~n15794;
  assign n15796 = ~n14221 & ~n15766;
  assign n15797 = n4406 & n6190;
  assign n15798 = ~n15796 & ~n15797;
  assign n15799 = n8959 & n15798;
  assign n15800 = n15116 & ~n15799;
  assign n15801 = ~n15795 & ~n15800;
  assign n15802 = ~n15789 & ~n15801;
  assign n15803 = ~n15788 & n15802;
  assign n15804 = ~n15787 & ~n15803;
  assign n15805 = pi232 & ~n15804;
  assign n15806 = ~n15268 & ~n15789;
  assign n15807 = ~n15805 & ~n15806;
  assign n15808 = ~pi100 & ~n15807;
  assign n15809 = ~n15772 & ~n15808;
  assign n15810 = n14475 & n15809;
  assign n15811 = pi135 & ~n15656;
  assign n15812 = pi134 & n15657;
  assign n15813 = ~n15811 & ~n15812;
  assign n15814 = n14021 & n15770;
  assign n15815 = n15813 & ~n15814;
  assign n15816 = ~n15810 & n15815;
  assign n15817 = n14021 & ~n15771;
  assign n15818 = ~n13993 & n15766;
  assign n15819 = ~pi51 & ~n15818;
  assign n15820 = ~n5744 & n15819;
  assign n15821 = ~n14200 & ~n15766;
  assign n15822 = n5745 & ~n15821;
  assign n15823 = pi170 & n14756;
  assign n15824 = n15822 & ~n15823;
  assign n15825 = ~n8959 & ~n15824;
  assign n15826 = ~pi170 & n15310;
  assign n15827 = pi170 & n15313;
  assign n15828 = pi216 & ~n15827;
  assign n15829 = ~n15826 & n15828;
  assign n15830 = ~n15825 & ~n15829;
  assign n15831 = ~n15820 & ~n15830;
  assign n15832 = n15790 & n15831;
  assign n15833 = ~n5745 & n15819;
  assign n15834 = ~n15824 & ~n15833;
  assign n15835 = n15116 & n15834;
  assign n15836 = ~n15832 & ~n15835;
  assign n15837 = pi185 & n15325;
  assign n15838 = ~pi185 & n15327;
  assign n15839 = ~pi299 & ~n15838;
  assign n15840 = ~n15837 & n15839;
  assign n15841 = n15836 & ~n15840;
  assign n15842 = pi232 & ~n15841;
  assign n15843 = n15342 & ~n15842;
  assign n15844 = ~pi299 & ~n14116;
  assign n15845 = pi170 & ~n15348;
  assign n15846 = ~pi170 & n14116;
  assign n15847 = ~n15845 & ~n15846;
  assign n15848 = n10392 & n15847;
  assign n15849 = n15345 & ~n15848;
  assign n15850 = ~n15844 & n15849;
  assign n15851 = ~n15843 & ~n15850;
  assign n15852 = ~pi38 & ~n15851;
  assign n15853 = ~n14909 & ~n15768;
  assign n15854 = pi38 & ~n15853;
  assign n15855 = ~pi194 & ~n15854;
  assign n15856 = ~n15852 & n15855;
  assign n15857 = pi185 & n15332;
  assign n15858 = ~pi185 & n15334;
  assign n15859 = ~pi299 & ~n15858;
  assign n15860 = ~n15857 & n15859;
  assign n15861 = n15836 & ~n15860;
  assign n15862 = pi232 & ~n15861;
  assign n15863 = n15342 & ~n15862;
  assign n15864 = n10680 & n15348;
  assign n15865 = n15849 & ~n15864;
  assign n15866 = ~n15863 & ~n15865;
  assign n15867 = ~pi38 & ~n15866;
  assign n15868 = ~n14909 & ~n15781;
  assign n15869 = pi38 & ~n15868;
  assign n15870 = pi194 & ~n15869;
  assign n15871 = ~n15867 & n15870;
  assign n15872 = ~n15856 & ~n15871;
  assign n15873 = ~pi100 & ~n15872;
  assign n15874 = ~n15772 & ~n15873;
  assign n15875 = n2537 & n15874;
  assign n15876 = ~n15813 & ~n15875;
  assign n15877 = ~n15817 & n15876;
  assign n15878 = ~n15816 & ~n15877;
  assign n15879 = ~po1038 & n15878;
  assign n15880 = n13993 & n15813;
  assign n15881 = pi232 & n15818;
  assign n15882 = n15652 & ~n15881;
  assign n15883 = ~n15880 & n15882;
  assign po292 = n15879 | n15883;
  assign n15885 = pi136 & ~n15260;
  assign n15886 = ~n15656 & ~n15885;
  assign n15887 = ~n14003 & ~n15886;
  assign n15888 = ~n14049 & n15887;
  assign n15889 = pi148 & n7420;
  assign n15890 = ~n13993 & ~n15889;
  assign n15891 = ~n15888 & ~n15890;
  assign n15892 = n15652 & ~n15891;
  assign n15893 = n9584 & ~n13993;
  assign n15894 = ~pi51 & ~n15893;
  assign n15895 = n14021 & n15894;
  assign n15896 = ~n2614 & ~n15894;
  assign n15897 = ~pi141 & ~pi299;
  assign n15898 = ~pi184 & n15327;
  assign n15899 = pi184 & n15325;
  assign n15900 = ~n15898 & ~n15899;
  assign n15901 = n15897 & n15900;
  assign n15902 = pi163 & n5744;
  assign n15903 = ~n14909 & ~n15902;
  assign n15904 = ~n5745 & n15903;
  assign n15905 = ~n15313 & n15902;
  assign n15906 = ~pi51 & n14757;
  assign n15907 = n5745 & ~n15906;
  assign n15908 = pi148 & ~n15907;
  assign n15909 = ~n15905 & n15908;
  assign n15910 = ~n15904 & n15909;
  assign n15911 = pi299 & ~n15910;
  assign n15912 = ~pi287 & n13322;
  assign n15913 = pi216 & ~n15912;
  assign n15914 = n2521 & ~n15913;
  assign n15915 = n5744 & n15914;
  assign n15916 = ~pi51 & ~n15915;
  assign n15917 = ~pi148 & n15916;
  assign n15918 = n15911 & ~n15917;
  assign n15919 = ~n15901 & ~n15918;
  assign n15920 = pi184 & n15332;
  assign n15921 = ~pi184 & n15334;
  assign n15922 = n9581 & ~n15921;
  assign n15923 = ~n15920 & n15922;
  assign n15924 = n15919 & ~n15923;
  assign n15925 = pi232 & ~n15924;
  assign n15926 = n15342 & ~n15925;
  assign n15927 = ~n9583 & ~n15348;
  assign n15928 = n9583 & n14116;
  assign n15929 = ~n15927 & ~n15928;
  assign n15930 = pi232 & n15929;
  assign n15931 = n15345 & ~n15930;
  assign n15932 = ~n15926 & ~n15931;
  assign n15933 = n2614 & n15932;
  assign n15934 = ~n15896 & ~n15933;
  assign n15935 = n2537 & n15934;
  assign n15936 = ~n15895 & ~n15935;
  assign n15937 = n15887 & n15936;
  assign n15938 = ~n13993 & n15895;
  assign n15939 = ~n13993 & n15894;
  assign n15940 = ~n10912 & ~n15939;
  assign n15941 = n2537 & ~n15940;
  assign n15942 = ~pi51 & n14540;
  assign n15943 = ~pi148 & ~n15942;
  assign n15944 = ~n15912 & ~n15943;
  assign n15945 = ~pi148 & n14049;
  assign n15946 = ~n15944 & ~n15945;
  assign n15947 = n8959 & n14525;
  assign n15948 = ~n6190 & n15286;
  assign n15949 = pi148 & ~n15948;
  assign n15950 = ~n15947 & n15949;
  assign n15951 = ~n15946 & ~n15950;
  assign n15952 = pi299 & ~n15951;
  assign n15953 = pi184 & n14503;
  assign n15954 = n15270 & ~n15953;
  assign n15955 = n15897 & ~n15954;
  assign n15956 = pi184 & n14209;
  assign n15957 = n15274 & ~n15956;
  assign n15958 = n9581 & ~n15957;
  assign n15959 = ~n15955 & ~n15958;
  assign n15960 = ~n15952 & n15959;
  assign n15961 = pi232 & ~n15960;
  assign n15962 = ~n15267 & ~n15961;
  assign n15963 = n10912 & ~n15962;
  assign n15964 = n15941 & ~n15963;
  assign n15965 = ~n15887 & ~n15964;
  assign n15966 = ~n15938 & n15965;
  assign n15967 = ~po1038 & ~n15966;
  assign n15968 = ~n15937 & n15967;
  assign po293 = n15892 | n15968;
  assign n15970 = ~pi39 & pi137;
  assign n15971 = n2575 & n10164;
  assign n15972 = n6165 & n11348;
  assign n15973 = ~pi299 & ~po1038;
  assign n15974 = ~pi198 & n11361;
  assign n15975 = n15973 & n15974;
  assign n15976 = ~n15972 & ~n15975;
  assign n15977 = ~n15971 & ~n15976;
  assign n15978 = ~pi210 & po1038;
  assign n15979 = n11348 & n15978;
  assign n15980 = ~n15977 & ~n15979;
  assign n15981 = n10280 & ~n15980;
  assign po294 = n15970 | n15981;
  assign n15983 = ~pi118 & n13321;
  assign n15984 = ~pi139 & n15983;
  assign n15985 = ~pi232 & ~n11261;
  assign n15986 = ~n6191 & n9582;
  assign n15987 = ~n9581 & ~n11261;
  assign n15988 = ~n15986 & ~n15987;
  assign n15989 = n6191 & n6448;
  assign n15990 = n8973 & n15989;
  assign n15991 = n9581 & ~n15990;
  assign n15992 = n15988 & ~n15991;
  assign n15993 = pi232 & ~n15992;
  assign n15994 = ~n15985 & ~n15993;
  assign n15995 = pi39 & ~n15994;
  assign n15996 = ~n9584 & n11264;
  assign n15997 = ~pi39 & ~n15996;
  assign n15998 = n10024 & ~n15997;
  assign n15999 = ~n15995 & n15998;
  assign n16000 = ~pi138 & n15999;
  assign n16001 = ~n15984 & ~n16000;
  assign n16002 = n8864 & ~n8934;
  assign n16003 = pi92 & ~n16002;
  assign n16004 = n2534 & ~n16003;
  assign n16005 = ~pi75 & ~n8944;
  assign n16006 = ~pi299 & ~n9643;
  assign n16007 = pi299 & ~n9294;
  assign n16008 = ~pi232 & ~n16007;
  assign n16009 = ~n16006 & n16008;
  assign n16010 = ~pi39 & ~n16009;
  assign n16011 = ~n6190 & ~n9643;
  assign n16012 = ~n13497 & ~n16011;
  assign n16013 = n9581 & ~n16012;
  assign n16014 = ~n9643 & n15897;
  assign n16015 = pi148 & n6190;
  assign n16016 = ~n9294 & ~n16015;
  assign n16017 = pi148 & n13533;
  assign n16018 = ~n16016 & ~n16017;
  assign n16019 = pi299 & ~n16018;
  assign n16020 = pi232 & ~n16019;
  assign n16021 = ~n16014 & n16020;
  assign n16022 = ~n16013 & n16021;
  assign n16023 = n16010 & ~n16022;
  assign n16024 = ~n8990 & ~n11495;
  assign n16025 = n9009 & ~n16024;
  assign n16026 = n13572 & ~n16025;
  assign n16027 = n6198 & n11495;
  assign n16028 = ~n8990 & ~n16027;
  assign n16029 = n8959 & ~n16028;
  assign n16030 = n8961 & ~n16029;
  assign n16031 = ~n16026 & ~n16030;
  assign n16032 = ~pi232 & ~n16031;
  assign n16033 = ~pi141 & n16026;
  assign n16034 = ~n8970 & ~n16024;
  assign n16035 = ~n8960 & ~n16034;
  assign n16036 = pi148 & ~n16035;
  assign n16037 = ~n9582 & ~n16030;
  assign n16038 = ~n16036 & ~n16037;
  assign n16039 = ~n8976 & n16025;
  assign n16040 = n13572 & ~n16039;
  assign n16041 = pi141 & n16040;
  assign n16042 = ~n16038 & ~n16041;
  assign n16043 = ~n16033 & n16042;
  assign n16044 = pi232 & ~n16043;
  assign n16045 = ~n16032 & ~n16044;
  assign n16046 = pi39 & ~n16045;
  assign n16047 = ~n16023 & ~n16046;
  assign n16048 = n2614 & n16047;
  assign n16049 = ~pi87 & ~n16048;
  assign n16050 = n16005 & ~n16049;
  assign n16051 = ~pi92 & ~n16050;
  assign n16052 = n16004 & ~n16051;
  assign n16053 = ~pi55 & ~n16052;
  assign n16054 = n8865 & ~n13594;
  assign n16055 = pi55 & ~n16054;
  assign n16056 = ~n16053 & ~n16055;
  assign n16057 = n2531 & ~n16056;
  assign n16058 = n9564 & ~n16057;
  assign n16059 = pi138 & n16058;
  assign n16060 = n16001 & ~n16059;
  assign n16061 = ~pi138 & ~n8829;
  assign n16062 = n16058 & n16061;
  assign n16063 = n15999 & ~n16061;
  assign n16064 = n15984 & ~n16063;
  assign n16065 = ~n16062 & n16064;
  assign po295 = ~n16060 & ~n16065;
  assign n16067 = n8916 & ~n16012;
  assign n16068 = ~n9643 & n15269;
  assign n16069 = ~n9294 & ~n15285;
  assign n16070 = pi169 & n13533;
  assign n16071 = ~n16069 & ~n16070;
  assign n16072 = pi299 & ~n16071;
  assign n16073 = pi232 & ~n16072;
  assign n16074 = ~n16068 & n16073;
  assign n16075 = ~n16067 & n16074;
  assign n16076 = n16010 & ~n16075;
  assign n16077 = pi191 & n16040;
  assign n16078 = ~pi191 & n16026;
  assign n16079 = ~pi169 & n8990;
  assign n16080 = ~n16034 & ~n16079;
  assign n16081 = n8959 & ~n16080;
  assign n16082 = n8961 & ~n16081;
  assign n16083 = ~n16078 & ~n16082;
  assign n16084 = ~n16077 & n16083;
  assign n16085 = pi232 & ~n16084;
  assign n16086 = ~n16032 & ~n16085;
  assign n16087 = pi39 & ~n16086;
  assign n16088 = ~n16076 & ~n16087;
  assign n16089 = n2614 & n16088;
  assign n16090 = ~pi87 & ~n16089;
  assign n16091 = n16005 & ~n16090;
  assign n16092 = ~pi92 & ~n16091;
  assign n16093 = n16004 & ~n16092;
  assign n16094 = ~pi55 & ~n16093;
  assign n16095 = ~n16055 & ~n16094;
  assign n16096 = n2531 & ~n16095;
  assign n16097 = n9564 & ~n16096;
  assign n16098 = pi139 & n16097;
  assign n16099 = ~n6191 & n8917;
  assign n16100 = ~pi191 & n11258;
  assign n16101 = n8916 & ~n15990;
  assign n16102 = ~n11260 & ~n16101;
  assign n16103 = ~n16100 & n16102;
  assign n16104 = ~n16099 & n16103;
  assign n16105 = pi232 & ~n16104;
  assign n16106 = ~n15985 & ~n16105;
  assign n16107 = pi39 & ~n16106;
  assign n16108 = n11264 & ~n15252;
  assign n16109 = ~pi39 & ~n16108;
  assign n16110 = n10024 & ~n16109;
  assign n16111 = ~n16107 & n16110;
  assign n16112 = ~pi139 & n16111;
  assign n16113 = ~n15983 & ~n16112;
  assign n16114 = ~n16098 & n16113;
  assign n16115 = ~pi139 & ~n8830;
  assign n16116 = n16097 & n16115;
  assign n16117 = n16111 & ~n16115;
  assign n16118 = n15983 & ~n16117;
  assign n16119 = ~n16116 & n16118;
  assign po296 = ~n16114 & ~n16119;
  assign n16121 = ~pi629 & pi1156;
  assign n16122 = pi629 & ~pi1156;
  assign n16123 = ~n16121 & ~n16122;
  assign n16124 = pi792 & ~n16123;
  assign n16125 = pi140 & ~n10020;
  assign n16126 = ~pi102 & ~n11083;
  assign n16127 = ~pi98 & ~n2778;
  assign n16128 = ~n16126 & n16127;
  assign n16129 = n2464 & n12123;
  assign n16130 = n16128 & n16129;
  assign n16131 = n8784 & n9078;
  assign n16132 = n16130 & n16131;
  assign n16133 = ~pi40 & ~n16132;
  assign n16134 = n10112 & ~n16133;
  assign n16135 = ~pi252 & ~n16134;
  assign n16136 = n2727 & ~n2755;
  assign n16137 = n2499 & n16130;
  assign n16138 = ~pi47 & ~n16137;
  assign n16139 = pi314 & n10068;
  assign n16140 = n16138 & ~n16139;
  assign n16141 = n16136 & ~n16140;
  assign n16142 = ~pi35 & ~n16141;
  assign n16143 = ~pi40 & n10061;
  assign n16144 = ~n16142 & n16143;
  assign n16145 = ~n2737 & ~n16144;
  assign n16146 = pi252 & n16145;
  assign n16147 = ~n16135 & ~n16146;
  assign n16148 = n2516 & n16147;
  assign n16149 = pi1092 & ~n12120;
  assign n16150 = n16148 & n16149;
  assign n16151 = ~pi88 & ~n16128;
  assign n16152 = n10802 & ~n16151;
  assign n16153 = n2500 & n16152;
  assign n16154 = ~pi47 & ~n16139;
  assign n16155 = ~n16153 & n16154;
  assign n16156 = n16136 & ~n16155;
  assign n16157 = ~pi35 & ~n16156;
  assign n16158 = pi252 & ~n16157;
  assign n16159 = n10061 & n16158;
  assign n16160 = ~pi252 & n16152;
  assign n16161 = n9157 & n16160;
  assign n16162 = ~pi40 & ~n16161;
  assign n16163 = ~n16159 & n16162;
  assign n16164 = n7368 & n10112;
  assign n16165 = ~n16163 & n16164;
  assign n16166 = ~n16150 & ~n16165;
  assign n16167 = pi1093 & ~n16166;
  assign n16168 = ~n2913 & ~n16167;
  assign n16169 = pi1092 & n6210;
  assign po1106 = n2913 & n16169;
  assign n16171 = n16148 & po1106;
  assign n16172 = ~n2914 & ~n16171;
  assign n16173 = ~n16168 & ~n16172;
  assign n16174 = ~pi1091 & n16167;
  assign n16175 = ~n16173 & ~n16174;
  assign n16176 = ~pi210 & n16175;
  assign n16177 = ~n3375 & ~n16163;
  assign n16178 = ~pi32 & ~n16177;
  assign n16179 = ~n2516 & ~n6374;
  assign n16180 = n6120 & ~n16179;
  assign n16181 = ~n16178 & n16180;
  assign n16182 = pi824 & n16181;
  assign n16183 = ~n16150 & ~n16182;
  assign n16184 = n7490 & ~n16183;
  assign n16185 = ~pi32 & ~n16147;
  assign n16186 = n16180 & ~n16185;
  assign n16187 = ~pi824 & pi829;
  assign n16188 = n16186 & n16187;
  assign n16189 = n16183 & ~n16188;
  assign n16190 = pi1093 & ~n16189;
  assign n16191 = ~n2913 & ~n16190;
  assign n16192 = ~n16172 & ~n16191;
  assign n16193 = ~n16184 & ~n16192;
  assign n16194 = pi210 & n16193;
  assign n16195 = ~n16176 & ~n16194;
  assign n16196 = pi299 & ~n16195;
  assign n16197 = ~pi198 & n16175;
  assign n16198 = pi198 & n16193;
  assign n16199 = ~n16197 & ~n16198;
  assign n16200 = ~pi299 & ~n16199;
  assign n16201 = ~n16196 & ~n16200;
  assign n16202 = ~pi39 & ~n16201;
  assign n16203 = ~n6178 & n6440;
  assign n16204 = ~pi120 & ~n16203;
  assign n16205 = pi120 & ~n2522;
  assign n16206 = ~n16204 & ~n16205;
  assign n16207 = n2934 & n16206;
  assign n16208 = pi616 & ~n16207;
  assign n16209 = ~n6183 & ~n16207;
  assign n16210 = n2934 & n16203;
  assign n16211 = ~pi120 & ~n16210;
  assign n16212 = n2522 & n2934;
  assign n16213 = n6181 & n13857;
  assign n16214 = n16212 & ~n16213;
  assign n16215 = pi120 & ~n16214;
  assign n16216 = pi1091 & ~n16215;
  assign n16217 = ~n16211 & n16216;
  assign n16218 = pi120 & ~n16212;
  assign n16219 = ~pi1091 & ~n16218;
  assign n16220 = pi120 & pi824;
  assign n16221 = n6181 & n16220;
  assign n16222 = ~n16211 & ~n16221;
  assign n16223 = n16219 & n16222;
  assign n16224 = ~n16217 & ~n16223;
  assign n16225 = ~n6190 & n16224;
  assign n16226 = n6190 & ~n16207;
  assign n16227 = ~n16225 & ~n16226;
  assign n16228 = n6183 & ~n16227;
  assign n16229 = ~n16209 & ~n16228;
  assign n16230 = ~pi614 & ~n16229;
  assign n16231 = pi614 & ~n16207;
  assign n16232 = ~n16230 & ~n16231;
  assign n16233 = ~pi616 & ~n16232;
  assign n16234 = ~n16208 & ~n16233;
  assign n16235 = pi681 & ~n16234;
  assign n16236 = pi680 & ~n16227;
  assign n16237 = ~pi680 & ~n16207;
  assign n16238 = pi616 & n6187;
  assign n16239 = ~n16237 & n16238;
  assign n16240 = ~n16236 & n16239;
  assign n16241 = pi616 & ~n6187;
  assign n16242 = n16207 & n16241;
  assign n16243 = ~n16240 & ~n16242;
  assign n16244 = ~pi681 & n16243;
  assign n16245 = ~n6188 & ~n16234;
  assign n16246 = n6188 & ~n16227;
  assign n16247 = ~pi616 & ~n16246;
  assign n16248 = ~n16245 & n16247;
  assign n16249 = n16244 & ~n16248;
  assign n16250 = ~n16235 & ~n16249;
  assign n16251 = n6236 & ~n16250;
  assign n16252 = n6190 & ~n16224;
  assign n16253 = ~pi662 & pi680;
  assign n16254 = ~n16234 & ~n16253;
  assign n16255 = n16224 & n16253;
  assign n16256 = ~n6190 & ~n16255;
  assign n16257 = ~n16254 & n16256;
  assign n16258 = ~n16252 & ~n16257;
  assign n16259 = ~pi661 & ~n16258;
  assign n16260 = ~n6190 & n16207;
  assign n16261 = ~n16252 & ~n16260;
  assign n16262 = ~n6185 & ~n16261;
  assign n16263 = n16224 & ~n16262;
  assign n16264 = pi661 & ~n16263;
  assign n16265 = ~pi681 & ~n16264;
  assign n16266 = ~n16259 & n16265;
  assign n16267 = ~n16263 & ~n16266;
  assign n16268 = ~n6236 & ~n16267;
  assign n16269 = ~n16251 & ~n16268;
  assign n16270 = pi223 & ~n16269;
  assign n16271 = n2607 & n16207;
  assign n16272 = ~pi824 & ~n16203;
  assign n16273 = n6440 & ~n10028;
  assign n16274 = pi1092 & n16273;
  assign n16275 = ~n10827 & ~n16274;
  assign n16276 = ~n16272 & ~n16275;
  assign n16277 = pi1093 & n16276;
  assign n16278 = ~pi120 & ~n16277;
  assign n16279 = n16219 & ~n16278;
  assign n16280 = n2913 & n16210;
  assign n16281 = ~pi829 & ~n16276;
  assign n16282 = pi829 & ~n16274;
  assign n16283 = n7431 & ~n16282;
  assign n16284 = ~n16281 & n16283;
  assign n16285 = ~n16280 & ~n16284;
  assign n16286 = pi1091 & ~n16285;
  assign n16287 = ~pi120 & ~n16286;
  assign n16288 = ~n16218 & ~n16287;
  assign n16289 = ~n16279 & ~n16288;
  assign n16290 = n6185 & ~n16289;
  assign n16291 = n6190 & ~n16289;
  assign n16292 = ~n16260 & ~n16291;
  assign n16293 = ~n6185 & ~n16292;
  assign n16294 = ~n16290 & ~n16293;
  assign n16295 = ~n6188 & n16294;
  assign n16296 = n6188 & n16289;
  assign n16297 = ~n16295 & ~n16296;
  assign n16298 = ~n6236 & n16297;
  assign n16299 = ~pi603 & ~n16207;
  assign n16300 = ~n6190 & n16289;
  assign n16301 = ~n16226 & ~n16300;
  assign n16302 = pi603 & ~n16301;
  assign n16303 = ~n16299 & ~n16302;
  assign n16304 = ~pi642 & ~n16303;
  assign n16305 = ~n16209 & ~n16304;
  assign n16306 = ~pi614 & ~n16305;
  assign n16307 = ~n16231 & ~n16306;
  assign n16308 = ~pi616 & ~n16307;
  assign n16309 = ~n16208 & ~n16308;
  assign n16310 = pi681 & ~n16309;
  assign n16311 = pi614 & ~n6187;
  assign n16312 = n16207 & n16311;
  assign n16313 = pi680 & ~n16301;
  assign n16314 = pi614 & n6187;
  assign n16315 = ~n16237 & n16314;
  assign n16316 = ~n16313 & n16315;
  assign n16317 = ~pi616 & ~n16305;
  assign n16318 = ~pi614 & ~n6188;
  assign n16319 = ~n16208 & n16318;
  assign n16320 = ~n16317 & n16319;
  assign n16321 = ~pi614 & n6188;
  assign n16322 = n16301 & n16321;
  assign n16323 = ~n16320 & ~n16322;
  assign n16324 = ~n16316 & n16323;
  assign n16325 = ~pi681 & n16324;
  assign n16326 = ~n16312 & n16325;
  assign n16327 = ~n16310 & ~n16326;
  assign n16328 = n6236 & n16327;
  assign n16329 = ~n16298 & ~n16328;
  assign n16330 = ~pi223 & n16329;
  assign n16331 = ~n2608 & ~n16330;
  assign n16332 = ~n16271 & ~n16331;
  assign n16333 = ~n16270 & ~n16332;
  assign n16334 = ~pi299 & ~n16333;
  assign n16335 = n6197 & ~n16327;
  assign n16336 = ~n6197 & ~n16297;
  assign n16337 = n6192 & ~n16336;
  assign n16338 = ~n16335 & n16337;
  assign n16339 = ~n2527 & n16338;
  assign n16340 = ~n6192 & n16297;
  assign n16341 = ~n2527 & n16340;
  assign n16342 = n2527 & n16207;
  assign n16343 = ~pi215 & ~n16342;
  assign n16344 = ~n16341 & n16343;
  assign n16345 = ~n16339 & n16344;
  assign n16346 = ~n6192 & n16267;
  assign n16347 = ~n6197 & ~n16267;
  assign n16348 = n6197 & ~n16250;
  assign n16349 = n6192 & ~n16348;
  assign n16350 = ~n16347 & n16349;
  assign n16351 = ~n16346 & ~n16350;
  assign n16352 = pi215 & n16351;
  assign n16353 = ~n16345 & ~n16352;
  assign n16354 = pi299 & ~n16353;
  assign n16355 = ~n16334 & ~n16354;
  assign n16356 = pi39 & ~n16355;
  assign n16357 = ~n16202 & ~n16356;
  assign n16358 = pi761 & n16357;
  assign n16359 = pi621 & n16173;
  assign n16360 = ~pi210 & ~n16359;
  assign n16361 = pi621 & n16192;
  assign n16362 = pi210 & ~n16361;
  assign n16363 = ~n16360 & ~n16362;
  assign n16364 = pi603 & ~n16363;
  assign n16365 = n16195 & ~n16364;
  assign n16366 = pi299 & ~n16365;
  assign n16367 = ~pi198 & ~n16359;
  assign n16368 = pi198 & ~n16361;
  assign n16369 = ~n16367 & ~n16368;
  assign n16370 = pi621 & ~n16174;
  assign n16371 = ~n16175 & ~n16370;
  assign n16372 = ~pi198 & n16371;
  assign n16373 = pi621 & ~n16184;
  assign n16374 = ~n16193 & ~n16373;
  assign n16375 = pi198 & n16374;
  assign n16376 = ~n16372 & ~n16375;
  assign n16377 = ~pi603 & ~n16376;
  assign n16378 = ~n16369 & ~n16377;
  assign n16379 = ~pi299 & n16378;
  assign n16380 = ~n16366 & ~n16379;
  assign n16381 = ~pi39 & ~n16380;
  assign n16382 = pi621 & pi1091;
  assign n16383 = n16207 & n16382;
  assign n16384 = n6190 & ~n16383;
  assign n16385 = n16288 & n16382;
  assign n16386 = ~n6190 & ~n16385;
  assign n16387 = ~n16384 & ~n16386;
  assign n16388 = pi603 & ~n16387;
  assign n16389 = n16301 & ~n16388;
  assign n16390 = n6188 & ~n16389;
  assign n16391 = ~pi614 & ~pi642;
  assign n16392 = ~pi616 & n16391;
  assign n16393 = pi603 & ~n16382;
  assign n16394 = n16207 & ~n16393;
  assign n16395 = ~n16392 & n16394;
  assign n16396 = ~n16299 & n16392;
  assign n16397 = ~n16388 & n16396;
  assign n16398 = ~n16395 & ~n16397;
  assign n16399 = ~n6188 & n16398;
  assign n16400 = ~n16390 & ~n16399;
  assign n16401 = n6198 & ~n16400;
  assign n16402 = n16297 & ~n16393;
  assign n16403 = ~n6198 & ~n16402;
  assign n16404 = ~n2527 & ~n16403;
  assign n16405 = ~n16401 & n16404;
  assign n16406 = n2527 & n16394;
  assign n16407 = ~n16405 & ~n16406;
  assign n16408 = ~pi215 & ~n16407;
  assign n16409 = pi621 & n16217;
  assign n16410 = ~n6190 & ~n16409;
  assign n16411 = ~n16384 & ~n16410;
  assign n16412 = pi603 & ~n16411;
  assign n16413 = n16396 & ~n16412;
  assign n16414 = ~n16395 & ~n16413;
  assign n16415 = ~n6188 & ~n16414;
  assign n16416 = n6188 & n16227;
  assign n16417 = ~n16412 & n16416;
  assign n16418 = ~n16415 & ~n16417;
  assign n16419 = n6198 & n16418;
  assign n16420 = n2934 & ~n16393;
  assign n16421 = ~n16261 & n16420;
  assign n16422 = n6185 & ~n16217;
  assign n16423 = n16421 & ~n16422;
  assign n16424 = ~n6188 & ~n16423;
  assign n16425 = ~n16224 & n16420;
  assign n16426 = pi680 & ~n16425;
  assign n16427 = n6187 & n16426;
  assign n16428 = ~n16424 & ~n16427;
  assign n16429 = ~n6198 & ~n16428;
  assign n16430 = pi215 & ~n16429;
  assign n16431 = ~n16419 & n16430;
  assign n16432 = ~n16408 & ~n16431;
  assign n16433 = pi299 & ~n16432;
  assign n16434 = n6236 & ~n16400;
  assign n16435 = ~n6236 & ~n16402;
  assign n16436 = ~n2607 & ~n16435;
  assign n16437 = ~n16434 & n16436;
  assign n16438 = n2607 & n16394;
  assign n16439 = ~n16437 & ~n16438;
  assign n16440 = ~pi223 & ~n16439;
  assign n16441 = n6236 & n16418;
  assign n16442 = ~n6236 & ~n16428;
  assign n16443 = pi223 & ~n16442;
  assign n16444 = ~n16441 & n16443;
  assign n16445 = ~n16440 & ~n16444;
  assign n16446 = ~pi299 & ~n16445;
  assign n16447 = ~n16433 & ~n16446;
  assign n16448 = pi39 & n16447;
  assign n16449 = ~n16381 & ~n16448;
  assign n16450 = ~pi761 & n16449;
  assign n16451 = ~pi140 & ~n16450;
  assign n16452 = ~n16358 & n16451;
  assign n16453 = pi603 & ~n16376;
  assign n16454 = ~pi299 & ~n16453;
  assign n16455 = ~pi210 & ~n16371;
  assign n16456 = pi210 & ~n16374;
  assign n16457 = ~n16455 & ~n16456;
  assign n16458 = pi603 & n16457;
  assign n16459 = pi299 & ~n16458;
  assign n16460 = ~n16454 & ~n16459;
  assign n16461 = ~pi39 & ~n16460;
  assign n16462 = n16342 & n16393;
  assign n16463 = n16301 & n16393;
  assign n16464 = n6188 & n16463;
  assign n16465 = n16207 & n16393;
  assign n16466 = ~n16392 & n16465;
  assign n16467 = n16392 & n16463;
  assign n16468 = ~n16466 & ~n16467;
  assign n16469 = ~n6188 & ~n16468;
  assign n16470 = ~n16464 & ~n16469;
  assign n16471 = n6198 & n16470;
  assign n16472 = n16297 & n16393;
  assign n16473 = ~n6198 & ~n16472;
  assign n16474 = ~n2527 & ~n16473;
  assign n16475 = ~n16471 & n16474;
  assign n16476 = ~pi215 & ~n16475;
  assign n16477 = ~n16462 & n16476;
  assign n16478 = ~n6198 & n16261;
  assign n16479 = ~n16225 & n16465;
  assign n16480 = ~n16261 & n16465;
  assign n16481 = n16225 & n16392;
  assign n16482 = n16480 & ~n16481;
  assign n16483 = ~n6188 & n16482;
  assign n16484 = ~n16479 & ~n16483;
  assign n16485 = ~n16478 & ~n16484;
  assign n16486 = pi215 & ~n16485;
  assign n16487 = pi299 & ~n16486;
  assign n16488 = ~n16477 & n16487;
  assign n16489 = ~n6236 & n16261;
  assign n16490 = ~n16484 & ~n16489;
  assign n16491 = pi223 & ~n16490;
  assign n16492 = ~pi299 & ~n16491;
  assign n16493 = ~n6236 & ~n16472;
  assign n16494 = n6236 & n16470;
  assign n16495 = ~n2607 & ~n16494;
  assign n16496 = ~n16493 & n16495;
  assign n16497 = n16271 & n16393;
  assign n16498 = ~pi223 & ~n16497;
  assign n16499 = ~n16496 & n16498;
  assign n16500 = n16492 & ~n16499;
  assign n16501 = ~n16488 & ~n16500;
  assign n16502 = pi39 & n16501;
  assign n16503 = ~n16461 & ~n16502;
  assign n16504 = pi140 & ~pi761;
  assign n16505 = n16503 & n16504;
  assign n16506 = ~n16452 & ~n16505;
  assign n16507 = ~pi38 & ~n16506;
  assign n16508 = n2934 & n6097;
  assign n16509 = ~pi140 & ~n16508;
  assign n16510 = n2934 & n16393;
  assign n16511 = n6097 & n16510;
  assign n16512 = ~pi761 & n16511;
  assign n16513 = ~n16509 & ~n16512;
  assign n16514 = pi38 & ~n16513;
  assign n16515 = ~n16507 & ~n16514;
  assign n16516 = n10020 & n16515;
  assign n16517 = ~n16125 & ~n16516;
  assign n16518 = ~pi608 & pi1153;
  assign n16519 = pi608 & ~pi1153;
  assign n16520 = ~n16518 & ~n16519;
  assign n16521 = pi778 & ~n16520;
  assign n16522 = ~n16517 & ~n16521;
  assign n16523 = ~pi38 & ~n16357;
  assign n16524 = n2934 & n6132;
  assign n16525 = pi38 & ~n16524;
  assign n16526 = ~n16523 & ~n16525;
  assign n16527 = n10020 & n16526;
  assign n16528 = ~pi140 & ~n16527;
  assign n16529 = n16521 & ~n16528;
  assign n16530 = ~n16522 & ~n16529;
  assign n16531 = ~pi785 & ~n16530;
  assign n16532 = pi609 & ~n16521;
  assign n16533 = ~n16528 & ~n16532;
  assign n16534 = pi609 & n16522;
  assign n16535 = ~n16533 & ~n16534;
  assign n16536 = pi1155 & ~n16535;
  assign n16537 = ~pi609 & ~n16521;
  assign n16538 = ~n16528 & ~n16537;
  assign n16539 = ~pi609 & n16522;
  assign n16540 = ~n16538 & ~n16539;
  assign n16541 = ~pi1155 & ~n16540;
  assign n16542 = ~n16536 & ~n16541;
  assign n16543 = pi785 & ~n16542;
  assign n16544 = ~n16531 & ~n16543;
  assign n16545 = ~pi781 & ~n16544;
  assign n16546 = pi618 & n16544;
  assign n16547 = ~pi618 & n16528;
  assign n16548 = pi1154 & ~n16547;
  assign n16549 = ~n16546 & n16548;
  assign n16550 = ~pi618 & n16544;
  assign n16551 = pi618 & n16528;
  assign n16552 = ~pi1154 & ~n16551;
  assign n16553 = ~n16550 & n16552;
  assign n16554 = ~n16549 & ~n16553;
  assign n16555 = pi781 & ~n16554;
  assign n16556 = ~n16545 & ~n16555;
  assign n16557 = ~pi789 & ~n16556;
  assign n16558 = pi619 & n16556;
  assign n16559 = ~pi619 & n16528;
  assign n16560 = pi1159 & ~n16559;
  assign n16561 = ~n16558 & n16560;
  assign n16562 = ~pi619 & n16556;
  assign n16563 = pi619 & n16528;
  assign n16564 = ~pi1159 & ~n16563;
  assign n16565 = ~n16562 & n16564;
  assign n16566 = ~n16561 & ~n16565;
  assign n16567 = pi789 & ~n16566;
  assign n16568 = ~n16557 & ~n16567;
  assign n16569 = ~pi626 & n16568;
  assign n16570 = pi626 & n16528;
  assign n16571 = ~pi1158 & ~n16570;
  assign n16572 = ~n16569 & n16571;
  assign n16573 = pi626 & n16568;
  assign n16574 = ~pi626 & n16528;
  assign n16575 = pi1158 & ~n16574;
  assign n16576 = ~n16573 & n16575;
  assign n16577 = ~n16572 & ~n16576;
  assign n16578 = pi788 & ~n16577;
  assign n16579 = ~pi788 & ~n16568;
  assign n16580 = ~n16578 & ~n16579;
  assign n16581 = ~n16124 & n16580;
  assign n16582 = n16124 & n16528;
  assign n16583 = ~n16581 & ~n16582;
  assign n16584 = pi647 & ~n16583;
  assign n16585 = pi628 & n16580;
  assign n16586 = ~pi627 & ~pi1154;
  assign n16587 = pi627 & pi1154;
  assign n16588 = pi781 & ~n16587;
  assign n16589 = ~n16586 & n16588;
  assign n16590 = ~pi660 & ~pi1155;
  assign n16591 = pi660 & pi1155;
  assign n16592 = pi785 & ~n16591;
  assign n16593 = ~n16590 & n16592;
  assign n16594 = ~n16528 & n16593;
  assign n16595 = pi665 & pi1091;
  assign n16596 = pi680 & ~n16595;
  assign n16597 = n16271 & n16596;
  assign n16598 = n16297 & n16596;
  assign n16599 = ~n6236 & ~n16598;
  assign n16600 = n16207 & ~n16595;
  assign n16601 = ~n6185 & n16600;
  assign n16602 = ~pi665 & n16288;
  assign n16603 = ~n16279 & ~n16602;
  assign n16604 = ~n16600 & n16603;
  assign n16605 = n16301 & ~n16604;
  assign n16606 = n6185 & n16605;
  assign n16607 = ~n16601 & ~n16606;
  assign n16608 = ~n6187 & n16607;
  assign n16609 = n6187 & ~n16605;
  assign n16610 = pi680 & ~n16609;
  assign n16611 = ~n16608 & n16610;
  assign n16612 = n6236 & ~n16611;
  assign n16613 = ~n2607 & ~n16612;
  assign n16614 = ~n16599 & n16613;
  assign n16615 = ~n16597 & ~n16614;
  assign n16616 = ~pi223 & ~n16615;
  assign n16617 = ~n16225 & n16600;
  assign n16618 = ~n16601 & ~n16617;
  assign n16619 = pi680 & ~n16618;
  assign n16620 = ~n16489 & n16619;
  assign n16621 = n6187 & ~n16617;
  assign n16622 = pi223 & ~n16621;
  assign n16623 = n16620 & n16622;
  assign n16624 = ~n16616 & ~n16623;
  assign n16625 = ~pi299 & ~n16624;
  assign n16626 = ~n6198 & n16598;
  assign n16627 = n6198 & n16611;
  assign n16628 = ~n2527 & ~n16627;
  assign n16629 = ~n16626 & n16628;
  assign n16630 = pi680 & n16600;
  assign n16631 = n2527 & ~n16630;
  assign n16632 = ~pi215 & ~n16631;
  assign n16633 = ~n16629 & n16632;
  assign n16634 = ~n16478 & n16619;
  assign n16635 = pi215 & ~n16621;
  assign n16636 = n16634 & n16635;
  assign n16637 = ~n16633 & ~n16636;
  assign n16638 = pi299 & ~n16637;
  assign n16639 = ~n16625 & ~n16638;
  assign n16640 = pi140 & ~n16639;
  assign n16641 = pi39 & pi140;
  assign n16642 = n16297 & ~n16598;
  assign n16643 = ~n6236 & ~n16642;
  assign n16644 = n16288 & n16595;
  assign n16645 = ~n6214 & n16644;
  assign n16646 = n16260 & n16595;
  assign n16647 = ~n6185 & n16646;
  assign n16648 = ~n16645 & ~n16647;
  assign n16649 = ~pi680 & ~n16309;
  assign n16650 = n16207 & n16595;
  assign n16651 = n6190 & ~n16650;
  assign n16652 = ~n6190 & ~n16644;
  assign n16653 = ~n16651 & ~n16652;
  assign n16654 = pi680 & ~n16653;
  assign n16655 = ~n16649 & ~n16654;
  assign n16656 = n16648 & ~n16655;
  assign n16657 = n16309 & ~n16656;
  assign n16658 = ~n6187 & n16657;
  assign n16659 = n6187 & n16655;
  assign n16660 = ~n16658 & ~n16659;
  assign n16661 = n6236 & n16660;
  assign n16662 = ~n2607 & ~n16661;
  assign n16663 = ~n16643 & n16662;
  assign n16664 = n2607 & n16206;
  assign n16665 = n2934 & ~n16596;
  assign n16666 = n16664 & n16665;
  assign n16667 = ~pi223 & ~n16666;
  assign n16668 = ~n16663 & n16667;
  assign n16669 = pi665 & n16217;
  assign n16670 = ~n6190 & ~n16669;
  assign n16671 = ~n16651 & ~n16670;
  assign n16672 = n6188 & ~n16671;
  assign n16673 = pi680 & ~n16669;
  assign n16674 = ~n16647 & n16673;
  assign n16675 = pi680 & ~n16671;
  assign n16676 = n16674 & n16675;
  assign n16677 = ~n16672 & ~n16676;
  assign n16678 = ~pi680 & n16263;
  assign n16679 = ~n16674 & ~n16678;
  assign n16680 = n16677 & n16679;
  assign n16681 = ~n6236 & n16680;
  assign n16682 = ~pi680 & ~n16234;
  assign n16683 = n16677 & ~n16682;
  assign n16684 = n6236 & n16683;
  assign n16685 = pi223 & ~n16684;
  assign n16686 = ~n16681 & n16685;
  assign n16687 = ~n16668 & ~n16686;
  assign n16688 = ~pi299 & ~n16687;
  assign n16689 = ~n6198 & ~n16642;
  assign n16690 = n6198 & n16660;
  assign n16691 = ~n2527 & ~n16690;
  assign n16692 = ~n16689 & n16691;
  assign n16693 = n16342 & ~n16596;
  assign n16694 = ~pi215 & ~n16693;
  assign n16695 = ~n16692 & n16694;
  assign n16696 = ~n6198 & n16680;
  assign n16697 = n6198 & n16683;
  assign n16698 = pi215 & ~n16697;
  assign n16699 = ~n16696 & n16698;
  assign n16700 = ~n16695 & ~n16699;
  assign n16701 = pi299 & ~n16700;
  assign n16702 = ~n16688 & ~n16701;
  assign n16703 = pi39 & n16702;
  assign n16704 = ~n16641 & ~n16703;
  assign n16705 = ~n16640 & ~n16704;
  assign n16706 = pi665 & n16192;
  assign n16707 = pi198 & ~n16706;
  assign n16708 = pi665 & n16173;
  assign n16709 = ~pi198 & ~n16708;
  assign n16710 = ~n16707 & ~n16709;
  assign n16711 = pi680 & ~n16710;
  assign n16712 = n16199 & ~n16711;
  assign n16713 = ~pi299 & ~n16712;
  assign n16714 = ~pi210 & ~n16708;
  assign n16715 = pi210 & ~n16706;
  assign n16716 = ~n16714 & ~n16715;
  assign n16717 = pi680 & ~n16716;
  assign n16718 = n16195 & ~n16717;
  assign n16719 = pi299 & ~n16718;
  assign n16720 = ~n16713 & ~n16719;
  assign n16721 = ~pi140 & ~n16720;
  assign n16722 = pi665 & ~n16174;
  assign n16723 = ~n16175 & ~n16722;
  assign n16724 = ~pi198 & ~n16723;
  assign n16725 = pi665 & ~n16184;
  assign n16726 = ~n16193 & ~n16725;
  assign n16727 = pi198 & ~n16726;
  assign n16728 = ~n16724 & ~n16727;
  assign n16729 = pi680 & n16728;
  assign n16730 = ~pi299 & ~n16729;
  assign n16731 = pi210 & ~n16726;
  assign n16732 = ~pi210 & ~n16723;
  assign n16733 = ~n16731 & ~n16732;
  assign n16734 = pi680 & n16733;
  assign n16735 = pi299 & ~n16734;
  assign n16736 = ~n16730 & ~n16735;
  assign n16737 = pi140 & n16736;
  assign n16738 = ~pi39 & ~n16737;
  assign n16739 = ~n16721 & n16738;
  assign n16740 = ~n16705 & ~n16739;
  assign n16741 = ~pi38 & ~n16740;
  assign n16742 = n2934 & n16596;
  assign n16743 = n6097 & n16742;
  assign n16744 = pi38 & ~n16743;
  assign n16745 = ~n16509 & n16744;
  assign n16746 = ~pi738 & ~n16745;
  assign n16747 = ~n16741 & n16746;
  assign n16748 = ~pi140 & ~n16526;
  assign n16749 = pi738 & n16748;
  assign n16750 = ~n16747 & ~n16749;
  assign n16751 = n10020 & n16750;
  assign n16752 = ~n16125 & ~n16751;
  assign n16753 = ~pi778 & ~n16752;
  assign n16754 = pi625 & n16752;
  assign n16755 = pi1153 & ~n16754;
  assign n16756 = ~pi625 & n16528;
  assign n16757 = n16755 & ~n16756;
  assign n16758 = ~pi625 & n16752;
  assign n16759 = ~pi1153 & ~n16758;
  assign n16760 = pi625 & n16528;
  assign n16761 = n16759 & ~n16760;
  assign n16762 = ~n16757 & ~n16761;
  assign n16763 = pi778 & ~n16762;
  assign n16764 = ~n16753 & ~n16763;
  assign n16765 = ~n16593 & ~n16764;
  assign n16766 = ~n16594 & ~n16765;
  assign n16767 = ~n16589 & n16766;
  assign n16768 = n16528 & n16589;
  assign n16769 = ~n16767 & ~n16768;
  assign n16770 = pi619 & ~n16769;
  assign n16771 = pi618 & n16766;
  assign n16772 = pi609 & n16764;
  assign n16773 = pi625 & n16517;
  assign n16774 = pi680 & ~n6187;
  assign n16775 = ~n16393 & ~n16595;
  assign n16776 = n16207 & ~n16775;
  assign n16777 = pi616 & ~n16776;
  assign n16778 = pi614 & ~n16776;
  assign n16779 = pi642 & ~n16776;
  assign n16780 = ~n16224 & n16465;
  assign n16781 = ~n16669 & ~n16780;
  assign n16782 = ~pi603 & n16646;
  assign n16783 = n16781 & ~n16782;
  assign n16784 = ~pi642 & ~n16479;
  assign n16785 = ~n16671 & n16784;
  assign n16786 = n16783 & n16785;
  assign n16787 = ~n16779 & ~n16786;
  assign n16788 = ~pi614 & ~n16787;
  assign n16789 = ~n16778 & ~n16788;
  assign n16790 = ~pi616 & ~n16789;
  assign n16791 = ~n16777 & ~n16790;
  assign n16792 = n16774 & ~n16791;
  assign n16793 = ~n16479 & n16672;
  assign n16794 = ~n16682 & ~n16793;
  assign n16795 = ~n16792 & n16794;
  assign n16796 = n6236 & ~n16795;
  assign n16797 = n6188 & n16781;
  assign n16798 = ~n16646 & ~n16669;
  assign n16799 = ~n16480 & n16798;
  assign n16800 = n16392 & n16783;
  assign n16801 = ~n16799 & ~n16800;
  assign n16802 = n16774 & ~n16801;
  assign n16803 = ~n16678 & ~n16802;
  assign n16804 = ~n16797 & n16803;
  assign n16805 = ~n6236 & ~n16804;
  assign n16806 = pi223 & ~n16805;
  assign n16807 = ~n16796 & n16806;
  assign n16808 = ~n16289 & ~n16385;
  assign n16809 = pi603 & n16808;
  assign n16810 = pi603 & ~pi621;
  assign n16811 = n16644 & ~n16810;
  assign n16812 = n6188 & ~n16811;
  assign n16813 = ~n16809 & n16812;
  assign n16814 = pi680 & n16775;
  assign n16815 = ~n16294 & ~n16814;
  assign n16816 = ~n6188 & ~n16815;
  assign n16817 = ~n16813 & ~n16816;
  assign n16818 = ~n6236 & n16817;
  assign n16819 = n16303 & ~n16775;
  assign n16820 = ~pi642 & ~n16819;
  assign n16821 = ~n16779 & ~n16820;
  assign n16822 = ~pi614 & ~n16821;
  assign n16823 = ~n16778 & ~n16822;
  assign n16824 = ~pi616 & ~n16823;
  assign n16825 = ~n16777 & ~n16824;
  assign n16826 = n16774 & ~n16825;
  assign n16827 = ~n16463 & ~n16653;
  assign n16828 = n6188 & n16827;
  assign n16829 = ~n16649 & ~n16828;
  assign n16830 = ~n16826 & n16829;
  assign n16831 = n6236 & n16830;
  assign n16832 = ~n2607 & ~n16831;
  assign n16833 = ~n16818 & n16832;
  assign n16834 = n16207 & ~n16814;
  assign n16835 = n2607 & ~n16834;
  assign n16836 = ~pi223 & ~n16835;
  assign n16837 = ~n16833 & n16836;
  assign n16838 = ~n16807 & ~n16837;
  assign n16839 = ~pi299 & ~n16838;
  assign n16840 = n2527 & ~n16834;
  assign n16841 = ~pi215 & ~n16840;
  assign n16842 = ~n6198 & n16817;
  assign n16843 = n6198 & n16830;
  assign n16844 = ~n2527 & ~n16843;
  assign n16845 = ~n16842 & n16844;
  assign n16846 = n16841 & ~n16845;
  assign n16847 = n6198 & ~n16795;
  assign n16848 = ~n6198 & ~n16804;
  assign n16849 = pi215 & ~n16848;
  assign n16850 = ~n16847 & n16849;
  assign n16851 = ~n16846 & ~n16850;
  assign n16852 = pi299 & ~n16851;
  assign n16853 = ~n16839 & ~n16852;
  assign n16854 = ~pi140 & n16853;
  assign n16855 = ~n16343 & ~n16841;
  assign n16856 = n6188 & ~n16603;
  assign n16857 = ~n16774 & ~n16856;
  assign n16858 = n16382 & n16602;
  assign n16859 = pi603 & ~n16858;
  assign n16860 = ~n16774 & n16859;
  assign n16861 = ~n16292 & ~n16393;
  assign n16862 = ~n16604 & n16861;
  assign n16863 = pi616 & ~n16862;
  assign n16864 = ~n16292 & ~n16604;
  assign n16865 = ~pi603 & ~n16864;
  assign n16866 = ~n16859 & ~n16865;
  assign n16867 = n16392 & ~n16866;
  assign n16868 = n16862 & ~n16867;
  assign n16869 = n16391 & n16866;
  assign n16870 = ~pi616 & ~n16869;
  assign n16871 = ~n16868 & n16870;
  assign n16872 = ~n16863 & ~n16871;
  assign n16873 = ~n6187 & ~n16872;
  assign n16874 = ~n16860 & ~n16873;
  assign n16875 = ~n16857 & n16874;
  assign n16876 = ~n6198 & ~n16875;
  assign n16877 = ~n16393 & n16600;
  assign n16878 = pi616 & ~n16877;
  assign n16879 = n16774 & ~n16878;
  assign n16880 = pi603 & pi665;
  assign n16881 = ~pi603 & ~n16600;
  assign n16882 = ~n16880 & ~n16881;
  assign n16883 = ~n16388 & n16882;
  assign n16884 = n16391 & n16883;
  assign n16885 = ~n16391 & n16877;
  assign n16886 = ~pi616 & ~n16885;
  assign n16887 = ~n16884 & n16886;
  assign n16888 = n16879 & ~n16887;
  assign n16889 = n16301 & n16828;
  assign n16890 = ~n16888 & ~n16889;
  assign n16891 = n6198 & n16890;
  assign n16892 = ~n2527 & ~n16891;
  assign n16893 = ~n16876 & n16892;
  assign n16894 = ~n16855 & ~n16893;
  assign n16895 = n16421 & n16882;
  assign n16896 = ~n16412 & n16882;
  assign n16897 = ~pi642 & ~n16896;
  assign n16898 = n16895 & ~n16897;
  assign n16899 = n6184 & ~n16898;
  assign n16900 = n16895 & ~n16899;
  assign n16901 = ~n6187 & ~n16900;
  assign n16902 = ~n16224 & n16814;
  assign n16903 = ~n16774 & ~n16902;
  assign n16904 = ~n16901 & ~n16903;
  assign n16905 = ~n6198 & n16904;
  assign n16906 = ~n16414 & ~n16595;
  assign n16907 = ~pi616 & ~n16906;
  assign n16908 = n16879 & ~n16907;
  assign n16909 = n16417 & n16882;
  assign n16910 = ~n16908 & ~n16909;
  assign n16911 = n6198 & ~n16910;
  assign n16912 = pi215 & ~n16911;
  assign n16913 = ~n16905 & n16912;
  assign n16914 = ~n16894 & ~n16913;
  assign n16915 = pi299 & ~n16914;
  assign n16916 = ~n16393 & ~n16596;
  assign n16917 = n16212 & n16916;
  assign n16918 = ~n16204 & n16917;
  assign n16919 = n2607 & n16918;
  assign n16920 = n2607 & ~n16207;
  assign n16921 = ~pi223 & ~n16920;
  assign n16922 = ~n16919 & n16921;
  assign n16923 = n6236 & ~n16890;
  assign n16924 = ~n6236 & n16875;
  assign n16925 = ~n2607 & ~n16924;
  assign n16926 = ~n16923 & n16925;
  assign n16927 = ~n16497 & ~n16926;
  assign n16928 = n16922 & n16927;
  assign n16929 = ~n6236 & ~n16904;
  assign n16930 = pi223 & ~n16929;
  assign n16931 = n6236 & n16910;
  assign n16932 = n16930 & ~n16931;
  assign n16933 = ~pi299 & ~n16932;
  assign n16934 = ~n16928 & n16933;
  assign n16935 = ~n16915 & ~n16934;
  assign n16936 = pi140 & n16935;
  assign n16937 = pi761 & ~n16936;
  assign n16938 = ~n16854 & n16937;
  assign n16939 = ~n16472 & n16857;
  assign n16940 = ~n16809 & ~n16866;
  assign n16941 = n16392 & ~n16940;
  assign n16942 = ~n16292 & n16393;
  assign n16943 = ~n16864 & ~n16942;
  assign n16944 = ~n16392 & ~n16943;
  assign n16945 = n16774 & ~n16944;
  assign n16946 = ~n16941 & n16945;
  assign n16947 = ~n16939 & ~n16946;
  assign n16948 = ~n6198 & ~n16947;
  assign n16949 = pi680 & ~n16463;
  assign n16950 = n16609 & n16949;
  assign n16951 = ~pi680 & n16468;
  assign n16952 = n16595 & ~n16810;
  assign n16953 = n16207 & ~n16952;
  assign n16954 = ~n16392 & n16953;
  assign n16955 = n16774 & ~n16954;
  assign n16956 = n16397 & n16595;
  assign n16957 = n16303 & n16392;
  assign n16958 = ~n16956 & n16957;
  assign n16959 = n16955 & ~n16958;
  assign n16960 = ~n16951 & ~n16959;
  assign n16961 = ~n16950 & n16960;
  assign n16962 = n6198 & ~n16961;
  assign n16963 = ~n2527 & ~n16962;
  assign n16964 = ~n16948 & n16963;
  assign n16965 = n2527 & n16206;
  assign n16966 = n2934 & ~n16916;
  assign n16967 = n16965 & n16966;
  assign n16968 = ~pi215 & ~n16967;
  assign n16969 = ~n16964 & n16968;
  assign n16970 = ~n16479 & n16618;
  assign n16971 = n16392 & ~n16970;
  assign n16972 = n16955 & ~n16971;
  assign n16973 = pi680 & ~n16621;
  assign n16974 = n16484 & ~n16973;
  assign n16975 = ~n16972 & ~n16974;
  assign n16976 = n6198 & n16975;
  assign n16977 = ~n16483 & ~n16780;
  assign n16978 = ~n16261 & n16600;
  assign n16979 = ~n16618 & n16973;
  assign n16980 = n16978 & n16979;
  assign n16981 = n16977 & ~n16980;
  assign n16982 = ~n6198 & ~n16981;
  assign n16983 = pi215 & ~n16982;
  assign n16984 = ~n16976 & n16983;
  assign n16985 = ~n16969 & ~n16984;
  assign n16986 = pi299 & ~n16985;
  assign n16987 = ~n6236 & n16947;
  assign n16988 = n6236 & n16961;
  assign n16989 = ~n2607 & ~n16988;
  assign n16990 = ~n16987 & n16989;
  assign n16991 = n16922 & ~n16990;
  assign n16992 = n6236 & ~n16975;
  assign n16993 = pi223 & ~n16992;
  assign n16994 = ~n6236 & n16981;
  assign n16995 = n16993 & ~n16994;
  assign n16996 = ~pi299 & ~n16995;
  assign n16997 = ~n16991 & n16996;
  assign n16998 = ~n16986 & ~n16997;
  assign n16999 = pi140 & n16998;
  assign n17000 = ~n16673 & ~n16810;
  assign n17001 = n6188 & ~n17000;
  assign n17002 = ~pi680 & ~n16423;
  assign n17003 = ~n16414 & ~n16798;
  assign n17004 = n16774 & ~n17003;
  assign n17005 = ~n17002 & ~n17004;
  assign n17006 = ~n17001 & n17005;
  assign n17007 = ~n6236 & n17006;
  assign n17008 = n16415 & ~n16596;
  assign n17009 = n6188 & ~n16810;
  assign n17010 = n16671 & n17009;
  assign n17011 = ~n17008 & ~n17010;
  assign n17012 = n6236 & ~n17011;
  assign n17013 = pi223 & ~n17012;
  assign n17014 = ~n17007 & n17013;
  assign n17015 = ~n16294 & ~n16393;
  assign n17016 = ~pi680 & ~n17015;
  assign n17017 = ~n16648 & n16952;
  assign n17018 = n16774 & ~n17017;
  assign n17019 = ~n16812 & ~n17018;
  assign n17020 = ~n17016 & n17019;
  assign n17021 = ~n6236 & ~n17020;
  assign n17022 = n16650 & ~n16810;
  assign n17023 = ~n16392 & n17022;
  assign n17024 = n16774 & ~n17023;
  assign n17025 = ~n16956 & n17024;
  assign n17026 = ~pi680 & n16398;
  assign n17027 = n16653 & n16952;
  assign n17028 = n6188 & ~n17027;
  assign n17029 = ~n17026 & ~n17028;
  assign n17030 = ~n17025 & n17029;
  assign n17031 = n6236 & ~n17030;
  assign n17032 = ~n2607 & ~n17031;
  assign n17033 = ~n17021 & n17032;
  assign n17034 = ~pi223 & ~n17033;
  assign n17035 = ~n16919 & n17034;
  assign n17036 = ~n17014 & ~n17035;
  assign n17037 = ~pi299 & ~n17036;
  assign n17038 = ~n6198 & ~n17020;
  assign n17039 = n6198 & ~n17030;
  assign n17040 = ~n2527 & ~n17039;
  assign n17041 = ~n17038 & n17040;
  assign n17042 = n2527 & n16918;
  assign n17043 = ~pi215 & ~n17042;
  assign n17044 = ~n17041 & n17043;
  assign n17045 = ~n6198 & n17006;
  assign n17046 = n6198 & ~n17011;
  assign n17047 = pi215 & ~n17046;
  assign n17048 = ~n17045 & n17047;
  assign n17049 = ~n17044 & ~n17048;
  assign n17050 = pi299 & ~n17049;
  assign n17051 = ~n17037 & ~n17050;
  assign n17052 = ~pi140 & ~n17051;
  assign n17053 = ~pi761 & ~n17052;
  assign n17054 = ~n16999 & n17053;
  assign n17055 = ~n16938 & ~n17054;
  assign n17056 = pi39 & ~n17055;
  assign n17057 = n16736 & ~n16880;
  assign n17058 = n16380 & n17057;
  assign n17059 = pi140 & ~n17058;
  assign n17060 = pi680 & n16460;
  assign n17061 = ~n16720 & ~n17060;
  assign n17062 = ~pi140 & ~n17061;
  assign n17063 = pi761 & ~n17062;
  assign n17064 = ~n17059 & n17063;
  assign n17065 = ~n16460 & ~n16736;
  assign n17066 = pi140 & n17065;
  assign n17067 = n16380 & n16720;
  assign n17068 = ~pi140 & n17067;
  assign n17069 = ~pi761 & ~n17068;
  assign n17070 = ~n17066 & n17069;
  assign n17071 = ~n17064 & ~n17070;
  assign n17072 = ~pi39 & n17071;
  assign n17073 = ~pi38 & ~n17072;
  assign n17074 = ~n17056 & n17073;
  assign n17075 = ~pi140 & ~n16212;
  assign n17076 = n16212 & ~n16916;
  assign n17077 = ~pi761 & n17076;
  assign n17078 = ~n17075 & ~n17077;
  assign n17079 = ~n16393 & n16742;
  assign n17080 = n2522 & n17079;
  assign n17081 = pi761 & n17080;
  assign n17082 = ~pi39 & ~n17081;
  assign n17083 = n17078 & n17082;
  assign n17084 = ~n16641 & ~n17083;
  assign n17085 = pi38 & n17084;
  assign n17086 = ~n17074 & ~n17085;
  assign n17087 = ~pi738 & ~n17086;
  assign n17088 = pi738 & ~n16515;
  assign n17089 = ~n17087 & ~n17088;
  assign n17090 = n10020 & n17089;
  assign n17091 = ~n16125 & ~n17090;
  assign n17092 = ~pi625 & n17091;
  assign n17093 = ~pi1153 & ~n17092;
  assign n17094 = ~n16773 & n17093;
  assign n17095 = ~pi608 & ~n16757;
  assign n17096 = ~n17094 & n17095;
  assign n17097 = ~pi625 & n16517;
  assign n17098 = pi625 & n17091;
  assign n17099 = ~n17097 & ~n17098;
  assign n17100 = pi1153 & n17099;
  assign n17101 = ~n16761 & ~n17100;
  assign n17102 = pi608 & n17101;
  assign n17103 = ~n17096 & ~n17102;
  assign n17104 = pi778 & ~n17103;
  assign n17105 = ~pi778 & n17091;
  assign n17106 = ~n17104 & ~n17105;
  assign n17107 = ~pi609 & ~n17106;
  assign n17108 = ~pi1155 & ~n17107;
  assign n17109 = ~n16772 & n17108;
  assign n17110 = ~pi660 & ~n16536;
  assign n17111 = ~n17109 & n17110;
  assign n17112 = ~pi609 & n16764;
  assign n17113 = pi609 & ~n17106;
  assign n17114 = ~n17112 & ~n17113;
  assign n17115 = pi1155 & n17114;
  assign n17116 = ~n16541 & ~n17115;
  assign n17117 = pi660 & n17116;
  assign n17118 = ~n17111 & ~n17117;
  assign n17119 = pi785 & ~n17118;
  assign n17120 = ~pi785 & ~n17106;
  assign n17121 = ~n17119 & ~n17120;
  assign n17122 = ~pi618 & ~n17121;
  assign n17123 = ~pi1154 & ~n17122;
  assign n17124 = ~n16771 & n17123;
  assign n17125 = ~pi627 & ~n16549;
  assign n17126 = ~n17124 & n17125;
  assign n17127 = ~pi618 & n16766;
  assign n17128 = pi618 & ~n17121;
  assign n17129 = ~n17127 & ~n17128;
  assign n17130 = pi1154 & n17129;
  assign n17131 = ~n16553 & ~n17130;
  assign n17132 = pi627 & n17131;
  assign n17133 = ~n17126 & ~n17132;
  assign n17134 = pi781 & ~n17133;
  assign n17135 = ~pi781 & ~n17121;
  assign n17136 = ~n17134 & ~n17135;
  assign n17137 = ~pi619 & ~n17136;
  assign n17138 = ~pi1159 & ~n17137;
  assign n17139 = ~n16770 & n17138;
  assign n17140 = ~pi648 & ~n16561;
  assign n17141 = ~n17139 & n17140;
  assign n17142 = ~pi619 & ~n16769;
  assign n17143 = pi619 & ~n17136;
  assign n17144 = ~n17142 & ~n17143;
  assign n17145 = pi1159 & n17144;
  assign n17146 = ~n16565 & ~n17145;
  assign n17147 = pi648 & n17146;
  assign n17148 = ~n17141 & ~n17147;
  assign n17149 = pi789 & ~n17148;
  assign n17150 = ~pi789 & ~n17136;
  assign n17151 = ~n17149 & ~n17150;
  assign n17152 = ~pi788 & n17151;
  assign n17153 = ~pi641 & ~pi1158;
  assign n17154 = ~n16572 & ~n17153;
  assign n17155 = ~pi626 & n17151;
  assign n17156 = ~pi648 & pi1159;
  assign n17157 = pi648 & ~pi1159;
  assign n17158 = ~n17156 & ~n17157;
  assign n17159 = pi789 & ~n17158;
  assign n17160 = ~n16528 & n17159;
  assign n17161 = n16769 & ~n17159;
  assign n17162 = ~n17160 & ~n17161;
  assign n17163 = pi626 & ~n17162;
  assign n17164 = ~pi641 & ~n17163;
  assign n17165 = ~n17155 & n17164;
  assign n17166 = ~n17154 & ~n17165;
  assign n17167 = pi641 & pi1158;
  assign n17168 = ~n16576 & ~n17167;
  assign n17169 = pi626 & n17151;
  assign n17170 = ~pi626 & ~n17162;
  assign n17171 = pi641 & ~n17170;
  assign n17172 = ~n17169 & n17171;
  assign n17173 = ~n17168 & ~n17172;
  assign n17174 = ~n17166 & ~n17173;
  assign n17175 = pi788 & ~n17174;
  assign n17176 = ~n17152 & ~n17175;
  assign n17177 = ~pi628 & n17176;
  assign n17178 = ~pi1156 & ~n17177;
  assign n17179 = ~n16585 & n17178;
  assign n17180 = ~pi641 & pi1158;
  assign n17181 = pi641 & ~pi1158;
  assign n17182 = ~n17180 & ~n17181;
  assign n17183 = pi788 & ~n17182;
  assign n17184 = n17162 & ~n17183;
  assign n17185 = n16528 & n17183;
  assign n17186 = ~n17184 & ~n17185;
  assign n17187 = pi628 & ~n17186;
  assign n17188 = pi1156 & ~n17187;
  assign n17189 = ~pi628 & n16528;
  assign n17190 = n17188 & ~n17189;
  assign n17191 = ~pi629 & ~n17190;
  assign n17192 = ~n17179 & n17191;
  assign n17193 = ~pi628 & ~n17186;
  assign n17194 = pi628 & n16528;
  assign n17195 = ~pi1156 & ~n17194;
  assign n17196 = ~n17193 & n17195;
  assign n17197 = ~pi628 & n16580;
  assign n17198 = pi628 & n17176;
  assign n17199 = ~n17197 & ~n17198;
  assign n17200 = pi1156 & n17199;
  assign n17201 = ~n17196 & ~n17200;
  assign n17202 = pi629 & n17201;
  assign n17203 = ~n17192 & ~n17202;
  assign n17204 = pi792 & ~n17203;
  assign n17205 = ~pi792 & n17176;
  assign n17206 = ~n17204 & ~n17205;
  assign n17207 = ~pi647 & ~n17206;
  assign n17208 = ~pi1157 & ~n17207;
  assign n17209 = ~n16584 & n17208;
  assign n17210 = ~pi792 & n17186;
  assign n17211 = ~n17190 & ~n17196;
  assign n17212 = pi792 & ~n17211;
  assign n17213 = ~n17210 & ~n17212;
  assign n17214 = pi647 & n17213;
  assign n17215 = pi1157 & ~n17214;
  assign n17216 = ~pi647 & n16528;
  assign n17217 = n17215 & ~n17216;
  assign n17218 = ~pi630 & ~n17217;
  assign n17219 = ~n17209 & n17218;
  assign n17220 = ~pi647 & n17213;
  assign n17221 = pi647 & n16528;
  assign n17222 = ~pi1157 & ~n17221;
  assign n17223 = ~n17220 & n17222;
  assign n17224 = ~pi647 & ~n16583;
  assign n17225 = pi647 & ~n17206;
  assign n17226 = ~n17224 & ~n17225;
  assign n17227 = pi1157 & n17226;
  assign n17228 = ~n17223 & ~n17227;
  assign n17229 = pi630 & n17228;
  assign n17230 = ~n17219 & ~n17229;
  assign n17231 = pi787 & ~n17230;
  assign n17232 = ~pi787 & ~n17206;
  assign n17233 = ~n17231 & ~n17232;
  assign n17234 = ~pi790 & n17233;
  assign n17235 = pi644 & ~n17233;
  assign n17236 = ~pi787 & ~n17213;
  assign n17237 = ~n17217 & ~n17223;
  assign n17238 = pi787 & ~n17237;
  assign n17239 = ~n17236 & ~n17238;
  assign n17240 = ~pi644 & n17239;
  assign n17241 = pi715 & ~n17240;
  assign n17242 = ~n17235 & n17241;
  assign n17243 = ~pi644 & n16528;
  assign n17244 = ~pi630 & pi1157;
  assign n17245 = pi630 & ~pi1157;
  assign n17246 = ~n17244 & ~n17245;
  assign n17247 = pi787 & ~n17246;
  assign n17248 = ~n16528 & n17247;
  assign n17249 = n16583 & ~n17247;
  assign n17250 = ~n17248 & ~n17249;
  assign n17251 = pi644 & n17250;
  assign n17252 = ~pi715 & ~n17251;
  assign n17253 = ~n17243 & n17252;
  assign n17254 = ~n17242 & ~n17253;
  assign n17255 = pi1160 & n17254;
  assign n17256 = ~pi644 & n17250;
  assign n17257 = pi715 & ~n17256;
  assign n17258 = pi644 & n16528;
  assign n17259 = n17257 & ~n17258;
  assign n17260 = pi644 & n17239;
  assign n17261 = ~pi644 & ~n17233;
  assign n17262 = ~pi715 & ~n17261;
  assign n17263 = ~n17260 & n17262;
  assign n17264 = ~n17259 & ~n17263;
  assign n17265 = ~pi1160 & n17264;
  assign n17266 = ~n17255 & ~n17265;
  assign n17267 = pi790 & n17266;
  assign n17268 = ~n17234 & ~n17267;
  assign n17269 = ~po1038 & n17268;
  assign n17270 = ~pi140 & po1038;
  assign n17271 = ~pi832 & ~n17270;
  assign n17272 = ~n17269 & n17271;
  assign n17273 = n2934 & n16521;
  assign n17274 = ~pi140 & ~n2934;
  assign n17275 = ~pi761 & n16510;
  assign n17276 = ~n17274 & ~n17275;
  assign n17277 = ~n17273 & ~n17276;
  assign n17278 = ~pi785 & ~n17277;
  assign n17279 = n2934 & ~n16532;
  assign n17280 = ~n17276 & ~n17279;
  assign n17281 = pi1155 & ~n17280;
  assign n17282 = pi609 & n2934;
  assign n17283 = n17277 & ~n17282;
  assign n17284 = ~pi1155 & ~n17283;
  assign n17285 = ~n17281 & ~n17284;
  assign n17286 = pi785 & ~n17285;
  assign n17287 = ~n17278 & ~n17286;
  assign n17288 = ~pi781 & ~n17287;
  assign n17289 = ~pi618 & n2934;
  assign n17290 = n17287 & ~n17289;
  assign n17291 = pi1154 & ~n17290;
  assign n17292 = pi618 & n2934;
  assign n17293 = n17287 & ~n17292;
  assign n17294 = ~pi1154 & ~n17293;
  assign n17295 = ~n17291 & ~n17294;
  assign n17296 = pi781 & ~n17295;
  assign n17297 = ~n17288 & ~n17296;
  assign n17298 = ~pi789 & ~n17297;
  assign n17299 = pi619 & n17297;
  assign n17300 = ~pi619 & n17274;
  assign n17301 = pi1159 & ~n17300;
  assign n17302 = ~n17299 & n17301;
  assign n17303 = ~pi619 & n17297;
  assign n17304 = pi619 & n17274;
  assign n17305 = ~pi1159 & ~n17304;
  assign n17306 = ~n17303 & n17305;
  assign n17307 = ~n17302 & ~n17306;
  assign n17308 = pi789 & ~n17307;
  assign n17309 = ~n17298 & ~n17308;
  assign n17310 = ~pi788 & ~n17309;
  assign n17311 = pi626 & n17309;
  assign n17312 = ~pi626 & n17274;
  assign n17313 = pi1158 & ~n17312;
  assign n17314 = ~n17311 & n17313;
  assign n17315 = ~pi626 & n17309;
  assign n17316 = pi626 & n17274;
  assign n17317 = ~pi1158 & ~n17316;
  assign n17318 = ~n17315 & n17317;
  assign n17319 = ~n17314 & ~n17318;
  assign n17320 = pi788 & ~n17319;
  assign n17321 = ~n17310 & ~n17320;
  assign n17322 = ~n16124 & n17321;
  assign n17323 = n16124 & n17274;
  assign n17324 = ~n17322 & ~n17323;
  assign n17325 = pi647 & ~n17324;
  assign n17326 = pi628 & n17321;
  assign n17327 = ~pi738 & n16742;
  assign n17328 = ~n17274 & ~n17327;
  assign n17329 = ~pi778 & n17328;
  assign n17330 = ~pi625 & n17327;
  assign n17331 = ~n17328 & ~n17330;
  assign n17332 = pi1153 & ~n17331;
  assign n17333 = ~pi1153 & ~n17274;
  assign n17334 = ~n17330 & n17333;
  assign n17335 = ~n17332 & ~n17334;
  assign n17336 = pi778 & ~n17335;
  assign n17337 = ~n17329 & ~n17336;
  assign n17338 = n2934 & n16593;
  assign n17339 = n17337 & ~n17338;
  assign n17340 = n2934 & n16589;
  assign n17341 = n17339 & ~n17340;
  assign n17342 = n2934 & n17159;
  assign n17343 = n17341 & ~n17342;
  assign n17344 = ~pi626 & pi1158;
  assign n17345 = pi626 & ~pi1158;
  assign n17346 = ~n17344 & ~n17345;
  assign n17347 = ~pi626 & pi641;
  assign n17348 = pi626 & ~pi641;
  assign n17349 = ~n17347 & ~n17348;
  assign n17350 = ~n17346 & ~n17349;
  assign n17351 = n17343 & n17350;
  assign n17352 = ~n17182 & n17319;
  assign n17353 = ~n17351 & ~n17352;
  assign n17354 = pi788 & ~n17353;
  assign n17355 = pi788 & ~n17346;
  assign n17356 = ~n17183 & ~n17355;
  assign n17357 = pi618 & n17339;
  assign n17358 = pi609 & n17337;
  assign n17359 = ~n16393 & ~n17328;
  assign n17360 = pi625 & n17359;
  assign n17361 = n17276 & ~n17359;
  assign n17362 = ~n17360 & ~n17361;
  assign n17363 = n17333 & ~n17362;
  assign n17364 = ~pi608 & ~n17332;
  assign n17365 = ~n17363 & n17364;
  assign n17366 = pi1153 & ~n17360;
  assign n17367 = n17276 & n17366;
  assign n17368 = ~n17334 & ~n17367;
  assign n17369 = pi608 & n17368;
  assign n17370 = ~n17365 & ~n17369;
  assign n17371 = pi778 & ~n17370;
  assign n17372 = ~pi778 & ~n17361;
  assign n17373 = ~n17371 & ~n17372;
  assign n17374 = ~pi609 & ~n17373;
  assign n17375 = ~pi1155 & ~n17374;
  assign n17376 = ~n17358 & n17375;
  assign n17377 = ~pi660 & ~n17281;
  assign n17378 = ~n17376 & n17377;
  assign n17379 = ~pi609 & n17337;
  assign n17380 = pi609 & ~n17373;
  assign n17381 = ~n17379 & ~n17380;
  assign n17382 = pi1155 & n17381;
  assign n17383 = ~n17284 & ~n17382;
  assign n17384 = pi660 & n17383;
  assign n17385 = ~n17378 & ~n17384;
  assign n17386 = pi785 & ~n17385;
  assign n17387 = ~pi785 & ~n17373;
  assign n17388 = ~n17386 & ~n17387;
  assign n17389 = ~pi618 & ~n17388;
  assign n17390 = ~pi1154 & ~n17389;
  assign n17391 = ~n17357 & n17390;
  assign n17392 = ~pi627 & ~n17291;
  assign n17393 = ~n17391 & n17392;
  assign n17394 = ~pi618 & n17339;
  assign n17395 = pi618 & ~n17388;
  assign n17396 = ~n17394 & ~n17395;
  assign n17397 = pi1154 & n17396;
  assign n17398 = ~n17294 & ~n17397;
  assign n17399 = pi627 & n17398;
  assign n17400 = ~n17393 & ~n17399;
  assign n17401 = pi781 & ~n17400;
  assign n17402 = ~pi781 & ~n17388;
  assign n17403 = ~n17401 & ~n17402;
  assign n17404 = ~pi789 & n17403;
  assign n17405 = n17356 & ~n17404;
  assign n17406 = ~pi619 & ~n17403;
  assign n17407 = pi619 & n17341;
  assign n17408 = ~pi1159 & ~n17407;
  assign n17409 = ~n17406 & n17408;
  assign n17410 = ~pi648 & ~n17409;
  assign n17411 = ~n17302 & n17410;
  assign n17412 = ~pi619 & n17341;
  assign n17413 = pi619 & ~n17403;
  assign n17414 = ~n17412 & ~n17413;
  assign n17415 = pi1159 & n17414;
  assign n17416 = ~n17306 & ~n17415;
  assign n17417 = pi648 & n17416;
  assign n17418 = ~n17411 & ~n17417;
  assign n17419 = pi789 & n17418;
  assign n17420 = n17405 & ~n17419;
  assign n17421 = ~n17354 & ~n17420;
  assign n17422 = ~pi628 & ~n17421;
  assign n17423 = ~pi1156 & ~n17422;
  assign n17424 = ~n17326 & n17423;
  assign n17425 = n2934 & n17183;
  assign n17426 = n17343 & ~n17425;
  assign n17427 = ~pi628 & n2934;
  assign n17428 = n17426 & ~n17427;
  assign n17429 = pi1156 & ~n17428;
  assign n17430 = ~pi629 & ~n17429;
  assign n17431 = ~n17424 & n17430;
  assign n17432 = ~pi628 & n17321;
  assign n17433 = pi628 & ~n17421;
  assign n17434 = ~n17432 & ~n17433;
  assign n17435 = pi1156 & n17434;
  assign n17436 = pi628 & n2934;
  assign n17437 = n17426 & ~n17436;
  assign n17438 = ~pi1156 & ~n17437;
  assign n17439 = pi629 & ~n17438;
  assign n17440 = ~n17435 & n17439;
  assign n17441 = ~n17431 & ~n17440;
  assign n17442 = pi792 & ~n17441;
  assign n17443 = ~pi792 & ~n17421;
  assign n17444 = ~n17442 & ~n17443;
  assign n17445 = ~pi647 & ~n17444;
  assign n17446 = ~pi1157 & ~n17445;
  assign n17447 = ~n17325 & n17446;
  assign n17448 = ~pi628 & pi1156;
  assign n17449 = pi628 & ~pi1156;
  assign n17450 = ~n17448 & ~n17449;
  assign n17451 = pi792 & ~n17450;
  assign n17452 = n2934 & n17451;
  assign n17453 = n17426 & ~n17452;
  assign n17454 = pi647 & n17453;
  assign n17455 = ~pi647 & n17274;
  assign n17456 = pi1157 & ~n17455;
  assign n17457 = ~n17454 & n17456;
  assign n17458 = ~pi630 & ~n17457;
  assign n17459 = ~n17447 & n17458;
  assign n17460 = ~pi647 & n17453;
  assign n17461 = pi647 & n17274;
  assign n17462 = ~pi1157 & ~n17461;
  assign n17463 = ~n17460 & n17462;
  assign n17464 = ~pi647 & ~n17324;
  assign n17465 = pi647 & ~n17444;
  assign n17466 = ~n17464 & ~n17465;
  assign n17467 = pi1157 & n17466;
  assign n17468 = ~n17463 & ~n17467;
  assign n17469 = pi630 & n17468;
  assign n17470 = ~n17459 & ~n17469;
  assign n17471 = pi787 & ~n17470;
  assign n17472 = ~pi787 & ~n17444;
  assign n17473 = ~n17471 & ~n17472;
  assign n17474 = pi644 & ~n17473;
  assign n17475 = ~pi787 & ~n17453;
  assign n17476 = ~n17457 & ~n17463;
  assign n17477 = pi787 & ~n17476;
  assign n17478 = ~n17475 & ~n17477;
  assign n17479 = ~pi644 & n17478;
  assign n17480 = pi715 & ~n17479;
  assign n17481 = ~n17474 & n17480;
  assign n17482 = n17247 & ~n17274;
  assign n17483 = ~n17247 & n17324;
  assign n17484 = ~n17482 & ~n17483;
  assign n17485 = pi644 & n17484;
  assign n17486 = ~pi644 & n17274;
  assign n17487 = ~pi715 & ~n17486;
  assign n17488 = ~n17485 & n17487;
  assign n17489 = pi1160 & ~n17488;
  assign n17490 = ~n17481 & n17489;
  assign n17491 = ~pi644 & n17484;
  assign n17492 = pi715 & ~n17491;
  assign n17493 = pi644 & n17274;
  assign n17494 = n17492 & ~n17493;
  assign n17495 = pi644 & n17478;
  assign n17496 = ~pi644 & ~n17473;
  assign n17497 = ~pi715 & ~n17496;
  assign n17498 = ~n17495 & n17497;
  assign n17499 = ~pi1160 & ~n17498;
  assign n17500 = ~n17494 & n17499;
  assign n17501 = ~n17490 & ~n17500;
  assign n17502 = pi790 & ~n17501;
  assign n17503 = ~pi790 & ~n17473;
  assign n17504 = pi832 & ~n17503;
  assign n17505 = ~n17502 & n17504;
  assign po297 = ~n17272 & ~n17505;
  assign n17507 = pi141 & ~n10020;
  assign n17508 = ~pi141 & ~n16508;
  assign n17509 = pi749 & n16511;
  assign n17510 = ~n17508 & ~n17509;
  assign n17511 = pi38 & ~n17510;
  assign n17512 = ~pi749 & n16355;
  assign n17513 = pi141 & n16501;
  assign n17514 = ~n17512 & ~n17513;
  assign n17515 = pi39 & ~n17514;
  assign n17516 = ~pi141 & n16449;
  assign n17517 = pi141 & n16461;
  assign n17518 = pi749 & ~n17517;
  assign n17519 = ~n17516 & n17518;
  assign n17520 = ~pi39 & n16201;
  assign n17521 = ~pi141 & ~pi749;
  assign n17522 = ~n17520 & n17521;
  assign n17523 = ~n17519 & ~n17522;
  assign n17524 = ~n17515 & ~n17523;
  assign n17525 = ~pi38 & n17524;
  assign n17526 = ~n17511 & ~n17525;
  assign n17527 = n10020 & n17526;
  assign n17528 = ~n17507 & ~n17527;
  assign n17529 = ~n16521 & ~n17528;
  assign n17530 = ~pi141 & ~n16527;
  assign n17531 = n16521 & ~n17530;
  assign n17532 = ~n17529 & ~n17531;
  assign n17533 = ~pi785 & ~n17532;
  assign n17534 = ~n16532 & ~n17530;
  assign n17535 = pi609 & n17529;
  assign n17536 = ~n17534 & ~n17535;
  assign n17537 = pi1155 & ~n17536;
  assign n17538 = ~n16537 & ~n17530;
  assign n17539 = ~pi609 & n17529;
  assign n17540 = ~n17538 & ~n17539;
  assign n17541 = ~pi1155 & ~n17540;
  assign n17542 = ~n17537 & ~n17541;
  assign n17543 = pi785 & ~n17542;
  assign n17544 = ~n17533 & ~n17543;
  assign n17545 = ~pi781 & ~n17544;
  assign n17546 = pi618 & n17544;
  assign n17547 = ~pi618 & n17530;
  assign n17548 = pi1154 & ~n17547;
  assign n17549 = ~n17546 & n17548;
  assign n17550 = ~pi618 & n17544;
  assign n17551 = pi618 & n17530;
  assign n17552 = ~pi1154 & ~n17551;
  assign n17553 = ~n17550 & n17552;
  assign n17554 = ~n17549 & ~n17553;
  assign n17555 = pi781 & ~n17554;
  assign n17556 = ~n17545 & ~n17555;
  assign n17557 = ~pi789 & ~n17556;
  assign n17558 = pi619 & n17556;
  assign n17559 = ~pi619 & n17530;
  assign n17560 = pi1159 & ~n17559;
  assign n17561 = ~n17558 & n17560;
  assign n17562 = ~pi619 & n17556;
  assign n17563 = pi619 & n17530;
  assign n17564 = ~pi1159 & ~n17563;
  assign n17565 = ~n17562 & n17564;
  assign n17566 = ~n17561 & ~n17565;
  assign n17567 = pi789 & ~n17566;
  assign n17568 = ~n17557 & ~n17567;
  assign n17569 = ~pi626 & n17568;
  assign n17570 = pi626 & n17530;
  assign n17571 = ~pi1158 & ~n17570;
  assign n17572 = ~n17569 & n17571;
  assign n17573 = pi626 & n17568;
  assign n17574 = ~pi626 & n17530;
  assign n17575 = pi1158 & ~n17574;
  assign n17576 = ~n17573 & n17575;
  assign n17577 = ~n17572 & ~n17576;
  assign n17578 = pi788 & ~n17577;
  assign n17579 = ~pi788 & ~n17568;
  assign n17580 = ~n17578 & ~n17579;
  assign n17581 = ~n16124 & n17580;
  assign n17582 = n16124 & n17530;
  assign n17583 = ~n17581 & ~n17582;
  assign n17584 = pi647 & ~n17583;
  assign n17585 = pi628 & n17580;
  assign n17586 = n16593 & ~n17530;
  assign n17587 = ~pi39 & ~n16736;
  assign n17588 = pi39 & n16639;
  assign n17589 = ~n17587 & ~n17588;
  assign n17590 = pi141 & n17589;
  assign n17591 = ~pi39 & n16720;
  assign n17592 = ~n16703 & ~n17591;
  assign n17593 = ~pi141 & n17592;
  assign n17594 = ~pi38 & ~n17593;
  assign n17595 = ~n17590 & n17594;
  assign n17596 = n16744 & ~n17508;
  assign n17597 = pi706 & ~n17596;
  assign n17598 = ~n17595 & n17597;
  assign n17599 = ~pi141 & ~pi706;
  assign n17600 = ~n16526 & n17599;
  assign n17601 = ~n17598 & ~n17600;
  assign n17602 = n10020 & n17601;
  assign n17603 = ~n17507 & ~n17602;
  assign n17604 = ~pi778 & ~n17603;
  assign n17605 = pi625 & n17603;
  assign n17606 = pi1153 & ~n17605;
  assign n17607 = ~pi625 & n17530;
  assign n17608 = n17606 & ~n17607;
  assign n17609 = ~pi625 & n17603;
  assign n17610 = ~pi1153 & ~n17609;
  assign n17611 = pi625 & n17530;
  assign n17612 = n17610 & ~n17611;
  assign n17613 = ~n17608 & ~n17612;
  assign n17614 = pi778 & ~n17613;
  assign n17615 = ~n17604 & ~n17614;
  assign n17616 = ~n16593 & ~n17615;
  assign n17617 = ~n17586 & ~n17616;
  assign n17618 = ~n16589 & n17617;
  assign n17619 = n16589 & n17530;
  assign n17620 = ~n17618 & ~n17619;
  assign n17621 = pi619 & ~n17620;
  assign n17622 = pi618 & n17617;
  assign n17623 = pi609 & n17615;
  assign n17624 = pi625 & n17528;
  assign n17625 = ~pi706 & ~n17526;
  assign n17626 = ~n16393 & n16743;
  assign n17627 = pi38 & ~n17626;
  assign n17628 = n17510 & n17627;
  assign n17629 = pi141 & n17058;
  assign n17630 = ~pi141 & n17061;
  assign n17631 = ~pi749 & ~n17630;
  assign n17632 = ~n17629 & n17631;
  assign n17633 = ~pi141 & ~n17067;
  assign n17634 = pi141 & ~n17065;
  assign n17635 = ~n17633 & ~n17634;
  assign n17636 = pi749 & n17635;
  assign n17637 = ~pi39 & ~n17636;
  assign n17638 = ~n17632 & n17637;
  assign n17639 = ~pi141 & ~n17051;
  assign n17640 = pi749 & ~n17639;
  assign n17641 = pi141 & n16998;
  assign n17642 = n17640 & ~n17641;
  assign n17643 = pi141 & n16935;
  assign n17644 = ~pi141 & n16853;
  assign n17645 = ~pi749 & ~n17644;
  assign n17646 = ~n17643 & n17645;
  assign n17647 = pi39 & ~n17646;
  assign n17648 = ~n17642 & n17647;
  assign n17649 = ~pi38 & ~n17648;
  assign n17650 = ~n17638 & n17649;
  assign n17651 = ~n17628 & ~n17650;
  assign n17652 = pi706 & n17651;
  assign n17653 = ~n17625 & ~n17652;
  assign n17654 = n10020 & n17653;
  assign n17655 = ~n17507 & ~n17654;
  assign n17656 = ~pi625 & n17655;
  assign n17657 = ~pi1153 & ~n17656;
  assign n17658 = ~n17624 & n17657;
  assign n17659 = ~pi608 & ~n17608;
  assign n17660 = ~n17658 & n17659;
  assign n17661 = ~pi625 & n17528;
  assign n17662 = pi625 & n17655;
  assign n17663 = ~n17661 & ~n17662;
  assign n17664 = pi1153 & n17663;
  assign n17665 = ~n17612 & ~n17664;
  assign n17666 = pi608 & n17665;
  assign n17667 = ~n17660 & ~n17666;
  assign n17668 = pi778 & ~n17667;
  assign n17669 = ~pi778 & n17655;
  assign n17670 = ~n17668 & ~n17669;
  assign n17671 = ~pi609 & ~n17670;
  assign n17672 = ~pi1155 & ~n17671;
  assign n17673 = ~n17623 & n17672;
  assign n17674 = ~pi660 & ~n17537;
  assign n17675 = ~n17673 & n17674;
  assign n17676 = ~pi609 & n17615;
  assign n17677 = pi609 & ~n17670;
  assign n17678 = ~n17676 & ~n17677;
  assign n17679 = pi1155 & n17678;
  assign n17680 = ~n17541 & ~n17679;
  assign n17681 = pi660 & n17680;
  assign n17682 = ~n17675 & ~n17681;
  assign n17683 = pi785 & ~n17682;
  assign n17684 = ~pi785 & ~n17670;
  assign n17685 = ~n17683 & ~n17684;
  assign n17686 = ~pi618 & ~n17685;
  assign n17687 = ~pi1154 & ~n17686;
  assign n17688 = ~n17622 & n17687;
  assign n17689 = ~pi627 & ~n17549;
  assign n17690 = ~n17688 & n17689;
  assign n17691 = ~pi618 & n17617;
  assign n17692 = pi618 & ~n17685;
  assign n17693 = ~n17691 & ~n17692;
  assign n17694 = pi1154 & n17693;
  assign n17695 = ~n17553 & ~n17694;
  assign n17696 = pi627 & n17695;
  assign n17697 = ~n17690 & ~n17696;
  assign n17698 = pi781 & ~n17697;
  assign n17699 = ~pi781 & ~n17685;
  assign n17700 = ~n17698 & ~n17699;
  assign n17701 = ~pi619 & ~n17700;
  assign n17702 = ~pi1159 & ~n17701;
  assign n17703 = ~n17621 & n17702;
  assign n17704 = ~pi648 & ~n17561;
  assign n17705 = ~n17703 & n17704;
  assign n17706 = ~pi619 & ~n17620;
  assign n17707 = pi619 & ~n17700;
  assign n17708 = ~n17706 & ~n17707;
  assign n17709 = pi1159 & n17708;
  assign n17710 = ~n17565 & ~n17709;
  assign n17711 = pi648 & n17710;
  assign n17712 = ~n17705 & ~n17711;
  assign n17713 = pi789 & ~n17712;
  assign n17714 = ~pi789 & ~n17700;
  assign n17715 = ~n17713 & ~n17714;
  assign n17716 = ~pi788 & n17715;
  assign n17717 = ~n17153 & ~n17572;
  assign n17718 = ~pi626 & n17715;
  assign n17719 = n17159 & ~n17530;
  assign n17720 = ~n17159 & n17620;
  assign n17721 = ~n17719 & ~n17720;
  assign n17722 = pi626 & ~n17721;
  assign n17723 = ~pi641 & ~n17722;
  assign n17724 = ~n17718 & n17723;
  assign n17725 = ~n17717 & ~n17724;
  assign n17726 = ~n17167 & ~n17576;
  assign n17727 = pi626 & n17715;
  assign n17728 = ~pi626 & ~n17721;
  assign n17729 = pi641 & ~n17728;
  assign n17730 = ~n17727 & n17729;
  assign n17731 = ~n17726 & ~n17730;
  assign n17732 = ~n17725 & ~n17731;
  assign n17733 = pi788 & ~n17732;
  assign n17734 = ~n17716 & ~n17733;
  assign n17735 = ~pi628 & n17734;
  assign n17736 = ~pi1156 & ~n17735;
  assign n17737 = ~n17585 & n17736;
  assign n17738 = ~n17183 & n17721;
  assign n17739 = n17183 & n17530;
  assign n17740 = ~n17738 & ~n17739;
  assign n17741 = pi628 & ~n17740;
  assign n17742 = pi1156 & ~n17741;
  assign n17743 = ~pi628 & n17530;
  assign n17744 = n17742 & ~n17743;
  assign n17745 = ~pi629 & ~n17744;
  assign n17746 = ~n17737 & n17745;
  assign n17747 = ~pi628 & ~n17740;
  assign n17748 = pi628 & n17530;
  assign n17749 = ~pi1156 & ~n17748;
  assign n17750 = ~n17747 & n17749;
  assign n17751 = ~pi628 & n17580;
  assign n17752 = pi628 & n17734;
  assign n17753 = ~n17751 & ~n17752;
  assign n17754 = pi1156 & n17753;
  assign n17755 = ~n17750 & ~n17754;
  assign n17756 = pi629 & n17755;
  assign n17757 = ~n17746 & ~n17756;
  assign n17758 = pi792 & ~n17757;
  assign n17759 = ~pi792 & n17734;
  assign n17760 = ~n17758 & ~n17759;
  assign n17761 = ~pi647 & ~n17760;
  assign n17762 = ~pi1157 & ~n17761;
  assign n17763 = ~n17584 & n17762;
  assign n17764 = ~pi792 & n17740;
  assign n17765 = ~n17744 & ~n17750;
  assign n17766 = pi792 & ~n17765;
  assign n17767 = ~n17764 & ~n17766;
  assign n17768 = pi647 & n17767;
  assign n17769 = pi1157 & ~n17768;
  assign n17770 = ~pi647 & n17530;
  assign n17771 = n17769 & ~n17770;
  assign n17772 = ~pi630 & ~n17771;
  assign n17773 = ~n17763 & n17772;
  assign n17774 = ~pi647 & n17767;
  assign n17775 = pi647 & n17530;
  assign n17776 = ~pi1157 & ~n17775;
  assign n17777 = ~n17774 & n17776;
  assign n17778 = ~pi647 & ~n17583;
  assign n17779 = pi647 & ~n17760;
  assign n17780 = ~n17778 & ~n17779;
  assign n17781 = pi1157 & n17780;
  assign n17782 = ~n17777 & ~n17781;
  assign n17783 = pi630 & n17782;
  assign n17784 = ~n17773 & ~n17783;
  assign n17785 = pi787 & ~n17784;
  assign n17786 = ~pi787 & ~n17760;
  assign n17787 = ~n17785 & ~n17786;
  assign n17788 = ~pi790 & n17787;
  assign n17789 = pi644 & ~n17787;
  assign n17790 = ~pi787 & ~n17767;
  assign n17791 = ~n17771 & ~n17777;
  assign n17792 = pi787 & ~n17791;
  assign n17793 = ~n17790 & ~n17792;
  assign n17794 = ~pi644 & n17793;
  assign n17795 = pi715 & ~n17794;
  assign n17796 = ~n17789 & n17795;
  assign n17797 = ~pi644 & n17530;
  assign n17798 = n17247 & ~n17530;
  assign n17799 = ~n17247 & n17583;
  assign n17800 = ~n17798 & ~n17799;
  assign n17801 = pi644 & n17800;
  assign n17802 = ~pi715 & ~n17801;
  assign n17803 = ~n17797 & n17802;
  assign n17804 = ~n17796 & ~n17803;
  assign n17805 = pi1160 & n17804;
  assign n17806 = ~pi644 & n17800;
  assign n17807 = pi715 & ~n17806;
  assign n17808 = pi644 & n17530;
  assign n17809 = n17807 & ~n17808;
  assign n17810 = pi644 & n17793;
  assign n17811 = ~pi644 & ~n17787;
  assign n17812 = ~pi715 & ~n17811;
  assign n17813 = ~n17810 & n17812;
  assign n17814 = ~n17809 & ~n17813;
  assign n17815 = ~pi1160 & n17814;
  assign n17816 = ~n17805 & ~n17815;
  assign n17817 = pi790 & n17816;
  assign n17818 = ~n17788 & ~n17817;
  assign n17819 = ~po1038 & n17818;
  assign n17820 = ~pi141 & po1038;
  assign n17821 = ~pi832 & ~n17820;
  assign n17822 = ~n17819 & n17821;
  assign n17823 = ~pi141 & ~n2934;
  assign n17824 = pi749 & n16510;
  assign n17825 = ~n17823 & ~n17824;
  assign n17826 = ~n17273 & ~n17825;
  assign n17827 = ~pi785 & ~n17826;
  assign n17828 = ~n17279 & ~n17825;
  assign n17829 = pi1155 & ~n17828;
  assign n17830 = ~n17282 & n17826;
  assign n17831 = ~pi1155 & ~n17830;
  assign n17832 = ~n17829 & ~n17831;
  assign n17833 = pi785 & ~n17832;
  assign n17834 = ~n17827 & ~n17833;
  assign n17835 = ~pi781 & ~n17834;
  assign n17836 = ~n17289 & n17834;
  assign n17837 = pi1154 & ~n17836;
  assign n17838 = ~n17292 & n17834;
  assign n17839 = ~pi1154 & ~n17838;
  assign n17840 = ~n17837 & ~n17839;
  assign n17841 = pi781 & ~n17840;
  assign n17842 = ~n17835 & ~n17841;
  assign n17843 = ~pi789 & ~n17842;
  assign n17844 = pi619 & n17842;
  assign n17845 = ~pi619 & n17823;
  assign n17846 = pi1159 & ~n17845;
  assign n17847 = ~n17844 & n17846;
  assign n17848 = ~pi619 & n17842;
  assign n17849 = pi619 & n17823;
  assign n17850 = ~pi1159 & ~n17849;
  assign n17851 = ~n17848 & n17850;
  assign n17852 = ~n17847 & ~n17851;
  assign n17853 = pi789 & ~n17852;
  assign n17854 = ~n17843 & ~n17853;
  assign n17855 = ~pi788 & ~n17854;
  assign n17856 = pi626 & n17854;
  assign n17857 = ~pi626 & n17823;
  assign n17858 = pi1158 & ~n17857;
  assign n17859 = ~n17856 & n17858;
  assign n17860 = ~pi626 & n17854;
  assign n17861 = pi626 & n17823;
  assign n17862 = ~pi1158 & ~n17861;
  assign n17863 = ~n17860 & n17862;
  assign n17864 = ~n17859 & ~n17863;
  assign n17865 = pi788 & ~n17864;
  assign n17866 = ~n17855 & ~n17865;
  assign n17867 = ~n16124 & n17866;
  assign n17868 = n16124 & n17823;
  assign n17869 = ~n17867 & ~n17868;
  assign n17870 = pi647 & ~n17869;
  assign n17871 = pi628 & n17866;
  assign n17872 = pi706 & n16742;
  assign n17873 = ~n17823 & ~n17872;
  assign n17874 = ~pi778 & n17873;
  assign n17875 = ~pi625 & n17872;
  assign n17876 = ~n17873 & ~n17875;
  assign n17877 = pi1153 & ~n17876;
  assign n17878 = ~pi1153 & ~n17823;
  assign n17879 = ~n17875 & n17878;
  assign n17880 = ~n17877 & ~n17879;
  assign n17881 = pi778 & ~n17880;
  assign n17882 = ~n17874 & ~n17881;
  assign n17883 = ~n17338 & n17882;
  assign n17884 = ~n17340 & n17883;
  assign n17885 = ~n17342 & n17884;
  assign n17886 = n17350 & n17885;
  assign n17887 = ~n17182 & n17864;
  assign n17888 = ~n17886 & ~n17887;
  assign n17889 = pi788 & ~n17888;
  assign n17890 = pi618 & n17883;
  assign n17891 = pi609 & n17882;
  assign n17892 = ~n16393 & ~n17873;
  assign n17893 = pi625 & n17892;
  assign n17894 = n17825 & ~n17892;
  assign n17895 = ~n17893 & ~n17894;
  assign n17896 = n17878 & ~n17895;
  assign n17897 = ~pi608 & ~n17877;
  assign n17898 = ~n17896 & n17897;
  assign n17899 = pi1153 & ~n17893;
  assign n17900 = n17825 & n17899;
  assign n17901 = ~n17879 & ~n17900;
  assign n17902 = pi608 & n17901;
  assign n17903 = ~n17898 & ~n17902;
  assign n17904 = pi778 & ~n17903;
  assign n17905 = ~pi778 & ~n17894;
  assign n17906 = ~n17904 & ~n17905;
  assign n17907 = ~pi609 & ~n17906;
  assign n17908 = ~pi1155 & ~n17907;
  assign n17909 = ~n17891 & n17908;
  assign n17910 = ~pi660 & ~n17829;
  assign n17911 = ~n17909 & n17910;
  assign n17912 = ~pi609 & n17882;
  assign n17913 = pi609 & ~n17906;
  assign n17914 = ~n17912 & ~n17913;
  assign n17915 = pi1155 & n17914;
  assign n17916 = ~n17831 & ~n17915;
  assign n17917 = pi660 & n17916;
  assign n17918 = ~n17911 & ~n17917;
  assign n17919 = pi785 & ~n17918;
  assign n17920 = ~pi785 & ~n17906;
  assign n17921 = ~n17919 & ~n17920;
  assign n17922 = ~pi618 & ~n17921;
  assign n17923 = ~pi1154 & ~n17922;
  assign n17924 = ~n17890 & n17923;
  assign n17925 = ~pi627 & ~n17837;
  assign n17926 = ~n17924 & n17925;
  assign n17927 = ~pi618 & n17883;
  assign n17928 = pi618 & ~n17921;
  assign n17929 = ~n17927 & ~n17928;
  assign n17930 = pi1154 & n17929;
  assign n17931 = ~n17839 & ~n17930;
  assign n17932 = pi627 & n17931;
  assign n17933 = ~n17926 & ~n17932;
  assign n17934 = pi781 & ~n17933;
  assign n17935 = ~pi781 & ~n17921;
  assign n17936 = ~n17934 & ~n17935;
  assign n17937 = ~pi619 & ~n17936;
  assign n17938 = pi619 & n17884;
  assign n17939 = ~pi1159 & ~n17938;
  assign n17940 = ~n17937 & n17939;
  assign n17941 = ~pi648 & ~n17940;
  assign n17942 = ~n17847 & n17941;
  assign n17943 = ~pi619 & n17884;
  assign n17944 = pi619 & ~n17936;
  assign n17945 = ~n17943 & ~n17944;
  assign n17946 = pi1159 & n17945;
  assign n17947 = ~n17851 & ~n17946;
  assign n17948 = pi648 & n17947;
  assign n17949 = ~n17942 & ~n17948;
  assign n17950 = pi789 & n17949;
  assign n17951 = ~pi789 & n17936;
  assign n17952 = n17356 & ~n17951;
  assign n17953 = ~n17950 & n17952;
  assign n17954 = ~n17889 & ~n17953;
  assign n17955 = ~pi628 & ~n17954;
  assign n17956 = ~pi1156 & ~n17955;
  assign n17957 = ~n17871 & n17956;
  assign n17958 = ~n17425 & n17885;
  assign n17959 = ~n17427 & n17958;
  assign n17960 = pi1156 & ~n17959;
  assign n17961 = ~pi629 & ~n17960;
  assign n17962 = ~n17957 & n17961;
  assign n17963 = ~pi628 & n17866;
  assign n17964 = pi628 & ~n17954;
  assign n17965 = ~n17963 & ~n17964;
  assign n17966 = pi1156 & n17965;
  assign n17967 = ~n17436 & n17958;
  assign n17968 = ~pi1156 & ~n17967;
  assign n17969 = pi629 & ~n17968;
  assign n17970 = ~n17966 & n17969;
  assign n17971 = ~n17962 & ~n17970;
  assign n17972 = pi792 & ~n17971;
  assign n17973 = ~pi792 & ~n17954;
  assign n17974 = ~n17972 & ~n17973;
  assign n17975 = ~pi647 & ~n17974;
  assign n17976 = ~pi1157 & ~n17975;
  assign n17977 = ~n17870 & n17976;
  assign n17978 = ~n17452 & n17958;
  assign n17979 = pi647 & n17978;
  assign n17980 = ~pi647 & n17823;
  assign n17981 = pi1157 & ~n17980;
  assign n17982 = ~n17979 & n17981;
  assign n17983 = ~pi630 & ~n17982;
  assign n17984 = ~n17977 & n17983;
  assign n17985 = ~pi647 & n17978;
  assign n17986 = pi647 & n17823;
  assign n17987 = ~pi1157 & ~n17986;
  assign n17988 = ~n17985 & n17987;
  assign n17989 = ~pi647 & ~n17869;
  assign n17990 = pi647 & ~n17974;
  assign n17991 = ~n17989 & ~n17990;
  assign n17992 = pi1157 & n17991;
  assign n17993 = ~n17988 & ~n17992;
  assign n17994 = pi630 & n17993;
  assign n17995 = ~n17984 & ~n17994;
  assign n17996 = pi787 & ~n17995;
  assign n17997 = ~pi787 & ~n17974;
  assign n17998 = ~n17996 & ~n17997;
  assign n17999 = pi644 & ~n17998;
  assign n18000 = ~pi787 & ~n17978;
  assign n18001 = ~n17982 & ~n17988;
  assign n18002 = pi787 & ~n18001;
  assign n18003 = ~n18000 & ~n18002;
  assign n18004 = ~pi644 & n18003;
  assign n18005 = pi715 & ~n18004;
  assign n18006 = ~n17999 & n18005;
  assign n18007 = n17247 & ~n17823;
  assign n18008 = ~n17247 & n17869;
  assign n18009 = ~n18007 & ~n18008;
  assign n18010 = pi644 & n18009;
  assign n18011 = ~pi644 & n17823;
  assign n18012 = ~pi715 & ~n18011;
  assign n18013 = ~n18010 & n18012;
  assign n18014 = pi1160 & ~n18013;
  assign n18015 = ~n18006 & n18014;
  assign n18016 = ~pi644 & n18009;
  assign n18017 = pi715 & ~n18016;
  assign n18018 = pi644 & n17823;
  assign n18019 = n18017 & ~n18018;
  assign n18020 = pi644 & n18003;
  assign n18021 = ~pi644 & ~n17998;
  assign n18022 = ~pi715 & ~n18021;
  assign n18023 = ~n18020 & n18022;
  assign n18024 = ~pi1160 & ~n18023;
  assign n18025 = ~n18019 & n18024;
  assign n18026 = ~n18015 & ~n18025;
  assign n18027 = pi790 & ~n18026;
  assign n18028 = ~pi790 & ~n17998;
  assign n18029 = pi832 & ~n18028;
  assign n18030 = ~n18027 & n18029;
  assign po298 = ~n17822 & ~n18030;
  assign n18032 = ~pi142 & ~n6274;
  assign n18033 = pi142 & ~n10020;
  assign n18034 = pi39 & pi142;
  assign n18035 = pi38 & ~n18034;
  assign n18036 = pi142 & ~n16212;
  assign n18037 = pi743 & n16510;
  assign n18038 = n2522 & n18037;
  assign n18039 = ~n18036 & ~n18038;
  assign n18040 = ~pi39 & ~n18039;
  assign n18041 = n18035 & ~n18040;
  assign n18042 = pi142 & n16365;
  assign n18043 = pi142 & ~n16195;
  assign n18044 = ~pi142 & ~n16458;
  assign n18045 = pi743 & ~n18044;
  assign n18046 = ~n18043 & ~n18045;
  assign n18047 = ~n18042 & ~n18046;
  assign n18048 = pi299 & ~n18047;
  assign n18049 = ~pi142 & ~n16453;
  assign n18050 = pi142 & ~n16378;
  assign n18051 = ~n18049 & ~n18050;
  assign n18052 = pi743 & n18051;
  assign n18053 = pi142 & ~pi743;
  assign n18054 = ~n16199 & n18053;
  assign n18055 = ~pi299 & ~n18054;
  assign n18056 = ~n18052 & n18055;
  assign n18057 = ~n18048 & ~n18056;
  assign n18058 = ~pi39 & n18057;
  assign n18059 = ~pi142 & n16470;
  assign n18060 = pi743 & ~n18059;
  assign n18061 = pi142 & n16400;
  assign n18062 = n18060 & ~n18061;
  assign n18063 = pi142 & ~n16327;
  assign n18064 = ~pi743 & n18063;
  assign n18065 = ~n18062 & ~n18064;
  assign n18066 = n6198 & n18065;
  assign n18067 = pi142 & ~n16297;
  assign n18068 = pi743 & n16472;
  assign n18069 = ~n18067 & ~n18068;
  assign n18070 = ~n6198 & n18069;
  assign n18071 = ~n2527 & ~n18070;
  assign n18072 = ~n18066 & n18071;
  assign n18073 = pi142 & ~n16207;
  assign n18074 = n16206 & n18037;
  assign n18075 = ~n18073 & ~n18074;
  assign n18076 = n2527 & ~n18075;
  assign n18077 = ~pi215 & ~n18076;
  assign n18078 = ~n18072 & n18077;
  assign n18079 = pi142 & ~n16267;
  assign n18080 = ~pi743 & ~n18079;
  assign n18081 = pi142 & ~n16428;
  assign n18082 = pi743 & ~n18081;
  assign n18083 = n16977 & n18082;
  assign n18084 = ~n18080 & ~n18083;
  assign n18085 = ~n6198 & n18084;
  assign n18086 = pi142 & ~n16250;
  assign n18087 = ~pi743 & ~n18086;
  assign n18088 = pi142 & n16418;
  assign n18089 = pi743 & ~n18088;
  assign n18090 = n16484 & n18089;
  assign n18091 = ~n18087 & ~n18090;
  assign n18092 = n6198 & n18091;
  assign n18093 = pi215 & ~n18092;
  assign n18094 = ~n18085 & n18093;
  assign n18095 = ~n18078 & ~n18094;
  assign n18096 = pi299 & ~n18095;
  assign n18097 = ~n6236 & ~n18084;
  assign n18098 = n6236 & ~n18091;
  assign n18099 = ~n18097 & ~n18098;
  assign n18100 = pi223 & n18099;
  assign n18101 = ~n6236 & ~n18069;
  assign n18102 = n6236 & ~n18065;
  assign n18103 = ~n2607 & ~n18102;
  assign n18104 = ~n18101 & n18103;
  assign n18105 = n2607 & ~n18073;
  assign n18106 = ~n18074 & n18105;
  assign n18107 = ~pi223 & ~n18106;
  assign n18108 = ~n18104 & n18107;
  assign n18109 = ~pi299 & ~n18108;
  assign n18110 = ~n18100 & n18109;
  assign n18111 = ~n18096 & ~n18110;
  assign n18112 = pi39 & n18111;
  assign n18113 = ~pi38 & ~n18112;
  assign n18114 = ~n18058 & n18113;
  assign n18115 = ~n18041 & ~n18114;
  assign n18116 = n10020 & n18115;
  assign n18117 = ~n18033 & ~n18116;
  assign n18118 = ~n16521 & ~n18117;
  assign n18119 = n10020 & ~n16525;
  assign n18120 = pi142 & ~n18119;
  assign n18121 = pi39 & ~n16334;
  assign n18122 = pi142 & ~n17520;
  assign n18123 = ~n18121 & n18122;
  assign n18124 = ~n6198 & ~n18079;
  assign n18125 = n6198 & ~n18086;
  assign n18126 = pi215 & ~n18125;
  assign n18127 = ~n18124 & n18126;
  assign n18128 = n6198 & n18063;
  assign n18129 = ~n6198 & n18067;
  assign n18130 = ~n2527 & ~n18129;
  assign n18131 = ~n18128 & n18130;
  assign n18132 = n2527 & ~n18073;
  assign n18133 = ~pi215 & ~n18132;
  assign n18134 = ~n18131 & n18133;
  assign n18135 = ~n18127 & ~n18134;
  assign n18136 = pi39 & ~n18135;
  assign n18137 = pi299 & n18136;
  assign n18138 = ~n18123 & ~n18137;
  assign n18139 = n2575 & ~n18138;
  assign n18140 = ~n18120 & ~n18139;
  assign n18141 = n16521 & ~n18140;
  assign n18142 = ~n18118 & ~n18141;
  assign n18143 = ~pi785 & ~n18142;
  assign n18144 = ~n16532 & ~n18140;
  assign n18145 = pi609 & n18118;
  assign n18146 = ~n18144 & ~n18145;
  assign n18147 = pi1155 & ~n18146;
  assign n18148 = ~n16537 & ~n18140;
  assign n18149 = ~pi609 & n18118;
  assign n18150 = ~n18148 & ~n18149;
  assign n18151 = ~pi1155 & ~n18150;
  assign n18152 = ~n18147 & ~n18151;
  assign n18153 = pi785 & ~n18152;
  assign n18154 = ~n18143 & ~n18153;
  assign n18155 = ~pi781 & ~n18154;
  assign n18156 = pi618 & n18154;
  assign n18157 = ~pi618 & n18140;
  assign n18158 = pi1154 & ~n18157;
  assign n18159 = ~n18156 & n18158;
  assign n18160 = ~pi618 & n18154;
  assign n18161 = pi618 & n18140;
  assign n18162 = ~pi1154 & ~n18161;
  assign n18163 = ~n18160 & n18162;
  assign n18164 = ~n18159 & ~n18163;
  assign n18165 = pi781 & ~n18164;
  assign n18166 = ~n18155 & ~n18165;
  assign n18167 = ~pi789 & ~n18166;
  assign n18168 = pi619 & n18166;
  assign n18169 = ~pi619 & n18140;
  assign n18170 = pi1159 & ~n18169;
  assign n18171 = ~n18168 & n18170;
  assign n18172 = ~pi619 & n18166;
  assign n18173 = pi619 & n18140;
  assign n18174 = ~pi1159 & ~n18173;
  assign n18175 = ~n18172 & n18174;
  assign n18176 = ~n18171 & ~n18175;
  assign n18177 = pi789 & ~n18176;
  assign n18178 = ~n18167 & ~n18177;
  assign n18179 = ~pi626 & n18178;
  assign n18180 = pi626 & n18140;
  assign n18181 = ~pi1158 & ~n18180;
  assign n18182 = ~n18179 & n18181;
  assign n18183 = pi626 & n18178;
  assign n18184 = ~pi626 & n18140;
  assign n18185 = pi1158 & ~n18184;
  assign n18186 = ~n18183 & n18185;
  assign n18187 = ~n18182 & ~n18186;
  assign n18188 = pi788 & ~n18187;
  assign n18189 = ~pi788 & ~n18178;
  assign n18190 = ~n18188 & ~n18189;
  assign n18191 = ~n16124 & n18190;
  assign n18192 = n16124 & n18140;
  assign n18193 = ~n18191 & ~n18192;
  assign n18194 = pi647 & ~n18193;
  assign n18195 = pi628 & n18190;
  assign n18196 = n16589 & ~n18140;
  assign n18197 = pi735 & n16742;
  assign n18198 = n2522 & n18197;
  assign n18199 = ~n18036 & ~n18198;
  assign n18200 = ~pi39 & ~n18199;
  assign n18201 = n18035 & ~n18200;
  assign n18202 = pi735 & n16598;
  assign n18203 = ~n18067 & ~n18202;
  assign n18204 = ~n6198 & ~n18203;
  assign n18205 = pi142 & ~n16660;
  assign n18206 = ~pi142 & ~n16611;
  assign n18207 = ~n18205 & ~n18206;
  assign n18208 = pi735 & ~n18207;
  assign n18209 = ~pi735 & ~n18063;
  assign n18210 = ~n18208 & ~n18209;
  assign n18211 = n6198 & n18210;
  assign n18212 = ~n2527 & ~n18211;
  assign n18213 = ~n18204 & n18212;
  assign n18214 = n16206 & n18197;
  assign n18215 = n18132 & ~n18214;
  assign n18216 = ~pi215 & ~n18215;
  assign n18217 = ~n18213 & n18216;
  assign n18218 = ~pi735 & ~n18079;
  assign n18219 = pi142 & ~n16680;
  assign n18220 = ~pi142 & n16979;
  assign n18221 = n16978 & n18220;
  assign n18222 = ~n18219 & ~n18221;
  assign n18223 = pi735 & n18222;
  assign n18224 = ~n18218 & ~n18223;
  assign n18225 = ~n6198 & ~n18224;
  assign n18226 = pi215 & ~n18225;
  assign n18227 = ~pi735 & ~n18086;
  assign n18228 = pi142 & ~n16683;
  assign n18229 = ~n18220 & ~n18228;
  assign n18230 = pi735 & n18229;
  assign n18231 = ~n18227 & ~n18230;
  assign n18232 = n6198 & ~n18231;
  assign n18233 = n18226 & ~n18232;
  assign n18234 = ~n18217 & ~n18233;
  assign n18235 = pi299 & n18234;
  assign n18236 = ~n6236 & ~n18224;
  assign n18237 = pi223 & ~n18236;
  assign n18238 = n6236 & ~n18231;
  assign n18239 = n18237 & ~n18238;
  assign n18240 = n18105 & ~n18214;
  assign n18241 = ~n6236 & ~n18203;
  assign n18242 = n6236 & n18210;
  assign n18243 = ~n2607 & ~n18242;
  assign n18244 = ~n18241 & n18243;
  assign n18245 = ~pi223 & ~n18244;
  assign n18246 = ~n18240 & n18245;
  assign n18247 = ~n18239 & ~n18246;
  assign n18248 = ~pi299 & n18247;
  assign n18249 = ~n18235 & ~n18248;
  assign n18250 = pi39 & n18249;
  assign n18251 = pi142 & n16720;
  assign n18252 = ~pi142 & ~n16736;
  assign n18253 = pi735 & ~n18252;
  assign n18254 = ~n18251 & n18253;
  assign n18255 = ~pi735 & ~n16201;
  assign n18256 = pi142 & n18255;
  assign n18257 = ~n18254 & ~n18256;
  assign n18258 = ~pi39 & ~n18257;
  assign n18259 = ~pi38 & ~n18258;
  assign n18260 = ~n18250 & n18259;
  assign n18261 = ~n18201 & ~n18260;
  assign n18262 = n10020 & n18261;
  assign n18263 = ~n18033 & ~n18262;
  assign n18264 = ~pi778 & ~n18263;
  assign n18265 = ~pi625 & n18263;
  assign n18266 = pi625 & n18140;
  assign n18267 = ~pi1153 & ~n18266;
  assign n18268 = ~n18265 & n18267;
  assign n18269 = pi625 & n18263;
  assign n18270 = ~pi625 & n18140;
  assign n18271 = pi1153 & ~n18270;
  assign n18272 = ~n18269 & n18271;
  assign n18273 = ~n18268 & ~n18272;
  assign n18274 = pi778 & ~n18273;
  assign n18275 = ~n18264 & ~n18274;
  assign n18276 = ~n16593 & n18275;
  assign n18277 = n16593 & n18140;
  assign n18278 = ~n18276 & ~n18277;
  assign n18279 = ~n16589 & n18278;
  assign n18280 = ~n18196 & ~n18279;
  assign n18281 = pi619 & n18280;
  assign n18282 = pi618 & ~n18278;
  assign n18283 = pi609 & n18275;
  assign n18284 = ~pi625 & n18117;
  assign n18285 = n16712 & n18050;
  assign n18286 = ~n16729 & n18049;
  assign n18287 = ~n18285 & ~n18286;
  assign n18288 = pi743 & ~n18287;
  assign n18289 = ~n16453 & ~n16712;
  assign n18290 = pi142 & n18289;
  assign n18291 = n16728 & ~n16880;
  assign n18292 = ~n16378 & n18291;
  assign n18293 = pi680 & n18292;
  assign n18294 = ~pi142 & n18293;
  assign n18295 = ~pi743 & ~n18294;
  assign n18296 = ~n18290 & n18295;
  assign n18297 = ~pi299 & ~n18296;
  assign n18298 = ~n18288 & n18297;
  assign n18299 = n16733 & ~n16880;
  assign n18300 = n16365 & n18299;
  assign n18301 = pi680 & n18300;
  assign n18302 = ~pi142 & n18301;
  assign n18303 = ~n16458 & ~n16718;
  assign n18304 = pi142 & n18303;
  assign n18305 = ~pi743 & ~n18304;
  assign n18306 = ~n18302 & n18305;
  assign n18307 = ~n16734 & n18044;
  assign n18308 = ~n16717 & n18042;
  assign n18309 = ~n18307 & ~n18308;
  assign n18310 = pi743 & ~n18309;
  assign n18311 = pi299 & ~n18310;
  assign n18312 = ~n18306 & n18311;
  assign n18313 = ~n18298 & ~n18312;
  assign n18314 = pi735 & ~n18313;
  assign n18315 = ~pi735 & n18057;
  assign n18316 = ~pi39 & ~n18315;
  assign n18317 = ~n18314 & n18316;
  assign n18318 = pi142 & n17006;
  assign n18319 = ~pi142 & n16981;
  assign n18320 = pi743 & ~n18319;
  assign n18321 = ~n18318 & n18320;
  assign n18322 = ~pi142 & ~n16904;
  assign n18323 = pi142 & n16804;
  assign n18324 = ~pi743 & ~n18323;
  assign n18325 = ~n18322 & n18324;
  assign n18326 = ~n18321 & ~n18325;
  assign n18327 = pi735 & ~n18326;
  assign n18328 = ~pi735 & n18084;
  assign n18329 = ~n18327 & ~n18328;
  assign n18330 = ~n6198 & n18329;
  assign n18331 = pi142 & ~n17011;
  assign n18332 = ~pi142 & ~n16975;
  assign n18333 = pi743 & ~n18332;
  assign n18334 = ~n18331 & n18333;
  assign n18335 = pi142 & n16795;
  assign n18336 = ~pi142 & n16910;
  assign n18337 = ~pi743 & ~n18336;
  assign n18338 = ~n18335 & n18337;
  assign n18339 = ~n18334 & ~n18338;
  assign n18340 = pi735 & ~n18339;
  assign n18341 = ~pi735 & n18091;
  assign n18342 = ~n18340 & ~n18341;
  assign n18343 = n6198 & n18342;
  assign n18344 = pi215 & ~n18343;
  assign n18345 = ~n18330 & n18344;
  assign n18346 = ~pi142 & ~n16947;
  assign n18347 = pi142 & n17020;
  assign n18348 = pi743 & ~n18347;
  assign n18349 = ~n18346 & n18348;
  assign n18350 = ~pi142 & ~n16875;
  assign n18351 = pi142 & n16817;
  assign n18352 = ~pi743 & ~n18351;
  assign n18353 = ~n18350 & n18352;
  assign n18354 = ~n18349 & ~n18353;
  assign n18355 = pi735 & ~n18354;
  assign n18356 = ~pi735 & ~n18069;
  assign n18357 = ~n18355 & ~n18356;
  assign n18358 = ~n6198 & ~n18357;
  assign n18359 = ~pi142 & ~n16961;
  assign n18360 = pi142 & n17030;
  assign n18361 = pi743 & ~n18360;
  assign n18362 = ~n18359 & n18361;
  assign n18363 = pi142 & n16830;
  assign n18364 = ~pi142 & n16890;
  assign n18365 = ~pi743 & ~n18364;
  assign n18366 = ~n18363 & n18365;
  assign n18367 = ~n18362 & ~n18366;
  assign n18368 = pi735 & ~n18367;
  assign n18369 = ~pi735 & ~n18065;
  assign n18370 = ~n18368 & ~n18369;
  assign n18371 = n6198 & ~n18370;
  assign n18372 = ~n2527 & ~n18371;
  assign n18373 = ~n18358 & n18372;
  assign n18374 = pi735 & n17079;
  assign n18375 = pi142 & ~n2934;
  assign n18376 = ~n18037 & ~n18375;
  assign n18377 = ~n18374 & n18376;
  assign n18378 = n16206 & ~n18377;
  assign n18379 = ~n18073 & ~n18378;
  assign n18380 = n2527 & n18379;
  assign n18381 = ~pi215 & ~n18380;
  assign n18382 = ~n18373 & n18381;
  assign n18383 = ~n18345 & ~n18382;
  assign n18384 = pi299 & ~n18383;
  assign n18385 = ~n6236 & n18329;
  assign n18386 = n6236 & n18342;
  assign n18387 = pi223 & ~n18386;
  assign n18388 = ~n18385 & n18387;
  assign n18389 = ~n6236 & ~n18357;
  assign n18390 = n6236 & ~n18370;
  assign n18391 = ~n2607 & ~n18390;
  assign n18392 = ~n18389 & n18391;
  assign n18393 = n2607 & n18379;
  assign n18394 = ~pi223 & ~n18393;
  assign n18395 = ~n18392 & n18394;
  assign n18396 = ~n18388 & ~n18395;
  assign n18397 = ~pi299 & ~n18396;
  assign n18398 = pi39 & ~n18397;
  assign n18399 = ~n18384 & n18398;
  assign n18400 = ~n18317 & ~n18399;
  assign n18401 = ~pi38 & ~n18400;
  assign n18402 = n6097 & n18374;
  assign n18403 = n18041 & ~n18402;
  assign n18404 = ~n18401 & ~n18403;
  assign n18405 = n10020 & n18404;
  assign n18406 = ~n18033 & ~n18405;
  assign n18407 = pi625 & n18406;
  assign n18408 = ~n18284 & ~n18407;
  assign n18409 = pi1153 & n18408;
  assign n18410 = pi608 & ~n18268;
  assign n18411 = ~n18409 & n18410;
  assign n18412 = ~pi625 & n18406;
  assign n18413 = pi625 & n18117;
  assign n18414 = ~pi1153 & ~n18413;
  assign n18415 = ~n18412 & n18414;
  assign n18416 = ~pi608 & ~n18272;
  assign n18417 = ~n18415 & n18416;
  assign n18418 = ~n18411 & ~n18417;
  assign n18419 = pi778 & ~n18418;
  assign n18420 = ~pi778 & n18406;
  assign n18421 = ~n18419 & ~n18420;
  assign n18422 = ~pi609 & ~n18421;
  assign n18423 = ~pi1155 & ~n18422;
  assign n18424 = ~n18283 & n18423;
  assign n18425 = ~pi660 & ~n18147;
  assign n18426 = ~n18424 & n18425;
  assign n18427 = ~pi609 & n18275;
  assign n18428 = pi609 & ~n18421;
  assign n18429 = ~n18427 & ~n18428;
  assign n18430 = pi1155 & n18429;
  assign n18431 = ~n18151 & ~n18430;
  assign n18432 = pi660 & n18431;
  assign n18433 = ~n18426 & ~n18432;
  assign n18434 = pi785 & ~n18433;
  assign n18435 = ~pi785 & ~n18421;
  assign n18436 = ~n18434 & ~n18435;
  assign n18437 = ~pi618 & ~n18436;
  assign n18438 = ~pi1154 & ~n18437;
  assign n18439 = ~n18282 & n18438;
  assign n18440 = ~pi627 & ~n18159;
  assign n18441 = ~n18439 & n18440;
  assign n18442 = ~pi618 & ~n18278;
  assign n18443 = pi618 & ~n18436;
  assign n18444 = ~n18442 & ~n18443;
  assign n18445 = pi1154 & n18444;
  assign n18446 = ~n18163 & ~n18445;
  assign n18447 = pi627 & n18446;
  assign n18448 = ~n18441 & ~n18447;
  assign n18449 = pi781 & ~n18448;
  assign n18450 = ~pi781 & ~n18436;
  assign n18451 = ~n18449 & ~n18450;
  assign n18452 = ~pi619 & ~n18451;
  assign n18453 = ~pi1159 & ~n18452;
  assign n18454 = ~n18281 & n18453;
  assign n18455 = ~pi648 & ~n18171;
  assign n18456 = ~n18454 & n18455;
  assign n18457 = ~pi619 & n18280;
  assign n18458 = pi619 & ~n18451;
  assign n18459 = ~n18457 & ~n18458;
  assign n18460 = pi1159 & n18459;
  assign n18461 = ~n18175 & ~n18460;
  assign n18462 = pi648 & n18461;
  assign n18463 = ~n18456 & ~n18462;
  assign n18464 = pi789 & ~n18463;
  assign n18465 = ~pi789 & ~n18451;
  assign n18466 = ~n18464 & ~n18465;
  assign n18467 = ~pi788 & n18466;
  assign n18468 = ~n17153 & ~n18182;
  assign n18469 = ~pi626 & n18466;
  assign n18470 = ~n17159 & n18280;
  assign n18471 = n17159 & n18140;
  assign n18472 = ~n18470 & ~n18471;
  assign n18473 = pi626 & n18472;
  assign n18474 = ~pi641 & ~n18473;
  assign n18475 = ~n18469 & n18474;
  assign n18476 = ~n18468 & ~n18475;
  assign n18477 = ~n17167 & ~n18186;
  assign n18478 = pi626 & n18466;
  assign n18479 = ~pi626 & n18472;
  assign n18480 = pi641 & ~n18479;
  assign n18481 = ~n18478 & n18480;
  assign n18482 = ~n18477 & ~n18481;
  assign n18483 = ~n18476 & ~n18482;
  assign n18484 = pi788 & ~n18483;
  assign n18485 = ~n18467 & ~n18484;
  assign n18486 = ~pi628 & n18485;
  assign n18487 = ~pi1156 & ~n18486;
  assign n18488 = ~n18195 & n18487;
  assign n18489 = ~n17183 & ~n18472;
  assign n18490 = n17183 & n18140;
  assign n18491 = ~n18489 & ~n18490;
  assign n18492 = pi628 & ~n18491;
  assign n18493 = ~pi628 & n18140;
  assign n18494 = pi1156 & ~n18493;
  assign n18495 = ~n18492 & n18494;
  assign n18496 = ~pi629 & ~n18495;
  assign n18497 = ~n18488 & n18496;
  assign n18498 = ~pi628 & ~n18491;
  assign n18499 = pi628 & n18140;
  assign n18500 = ~pi1156 & ~n18499;
  assign n18501 = ~n18498 & n18500;
  assign n18502 = ~pi628 & n18190;
  assign n18503 = pi628 & n18485;
  assign n18504 = ~n18502 & ~n18503;
  assign n18505 = pi1156 & n18504;
  assign n18506 = ~n18501 & ~n18505;
  assign n18507 = pi629 & n18506;
  assign n18508 = ~n18497 & ~n18507;
  assign n18509 = pi792 & ~n18508;
  assign n18510 = ~pi792 & n18485;
  assign n18511 = ~n18509 & ~n18510;
  assign n18512 = ~pi647 & ~n18511;
  assign n18513 = ~pi1157 & ~n18512;
  assign n18514 = ~n18194 & n18513;
  assign n18515 = ~pi792 & n18491;
  assign n18516 = ~n18495 & ~n18501;
  assign n18517 = pi792 & ~n18516;
  assign n18518 = ~n18515 & ~n18517;
  assign n18519 = pi647 & n18518;
  assign n18520 = ~pi647 & n18140;
  assign n18521 = pi1157 & ~n18520;
  assign n18522 = ~n18519 & n18521;
  assign n18523 = ~pi630 & ~n18522;
  assign n18524 = ~n18514 & n18523;
  assign n18525 = ~pi647 & n18518;
  assign n18526 = pi647 & n18140;
  assign n18527 = ~pi1157 & ~n18526;
  assign n18528 = ~n18525 & n18527;
  assign n18529 = ~pi647 & ~n18193;
  assign n18530 = pi647 & ~n18511;
  assign n18531 = ~n18529 & ~n18530;
  assign n18532 = pi1157 & n18531;
  assign n18533 = ~n18528 & ~n18532;
  assign n18534 = pi630 & n18533;
  assign n18535 = ~n18524 & ~n18534;
  assign n18536 = pi787 & ~n18535;
  assign n18537 = ~pi787 & ~n18511;
  assign n18538 = ~n18536 & ~n18537;
  assign n18539 = ~pi790 & n18538;
  assign n18540 = pi644 & ~n18538;
  assign n18541 = ~pi787 & ~n18518;
  assign n18542 = ~n18522 & ~n18528;
  assign n18543 = pi787 & ~n18542;
  assign n18544 = ~n18541 & ~n18543;
  assign n18545 = ~pi644 & n18544;
  assign n18546 = pi715 & ~n18545;
  assign n18547 = ~n18540 & n18546;
  assign n18548 = ~pi644 & n18140;
  assign n18549 = n17247 & ~n18140;
  assign n18550 = ~n17247 & n18193;
  assign n18551 = ~n18549 & ~n18550;
  assign n18552 = pi644 & n18551;
  assign n18553 = ~pi715 & ~n18552;
  assign n18554 = ~n18548 & n18553;
  assign n18555 = ~n18547 & ~n18554;
  assign n18556 = pi1160 & n18555;
  assign n18557 = ~pi644 & n18551;
  assign n18558 = pi715 & ~n18557;
  assign n18559 = pi644 & n18140;
  assign n18560 = n18558 & ~n18559;
  assign n18561 = pi644 & n18544;
  assign n18562 = ~pi644 & ~n18538;
  assign n18563 = ~pi715 & ~n18562;
  assign n18564 = ~n18561 & n18563;
  assign n18565 = ~n18560 & ~n18564;
  assign n18566 = ~pi1160 & n18565;
  assign n18567 = ~n18556 & ~n18566;
  assign n18568 = pi790 & n18567;
  assign n18569 = ~n18539 & ~n18568;
  assign n18570 = n6274 & n18569;
  assign n18571 = ~pi57 & ~n18570;
  assign n18572 = ~n18032 & n18571;
  assign n18573 = pi57 & pi142;
  assign n18574 = ~pi832 & ~n18573;
  assign n18575 = ~n18572 & n18574;
  assign n18576 = pi1155 & ~n18375;
  assign n18577 = ~n16521 & n18037;
  assign n18578 = pi609 & n18577;
  assign n18579 = n18576 & ~n18578;
  assign n18580 = ~pi1155 & ~n18375;
  assign n18581 = ~pi609 & n18577;
  assign n18582 = n18580 & ~n18581;
  assign n18583 = ~n18579 & ~n18582;
  assign n18584 = pi785 & ~n18583;
  assign n18585 = ~pi785 & ~n18375;
  assign n18586 = ~n18577 & n18585;
  assign n18587 = ~n18584 & ~n18586;
  assign n18588 = ~pi781 & ~n18587;
  assign n18589 = pi618 & n18587;
  assign n18590 = ~pi618 & n18375;
  assign n18591 = pi1154 & ~n18590;
  assign n18592 = ~n18589 & n18591;
  assign n18593 = ~pi618 & n18587;
  assign n18594 = pi618 & n18375;
  assign n18595 = ~pi1154 & ~n18594;
  assign n18596 = ~n18593 & n18595;
  assign n18597 = ~n18592 & ~n18596;
  assign n18598 = pi781 & ~n18597;
  assign n18599 = ~n18588 & ~n18598;
  assign n18600 = ~pi789 & ~n18599;
  assign n18601 = pi619 & n18599;
  assign n18602 = ~pi619 & n18375;
  assign n18603 = pi1159 & ~n18602;
  assign n18604 = ~n18601 & n18603;
  assign n18605 = ~pi619 & n18599;
  assign n18606 = pi619 & n18375;
  assign n18607 = ~pi1159 & ~n18606;
  assign n18608 = ~n18605 & n18607;
  assign n18609 = ~n18604 & ~n18608;
  assign n18610 = pi789 & ~n18609;
  assign n18611 = ~n18600 & ~n18610;
  assign n18612 = ~pi788 & ~n18611;
  assign n18613 = pi626 & n18611;
  assign n18614 = ~pi626 & n18375;
  assign n18615 = pi1158 & ~n18614;
  assign n18616 = ~n18613 & n18615;
  assign n18617 = ~pi626 & n18611;
  assign n18618 = pi626 & n18375;
  assign n18619 = ~pi1158 & ~n18618;
  assign n18620 = ~n18617 & n18619;
  assign n18621 = ~n18616 & ~n18620;
  assign n18622 = pi788 & ~n18621;
  assign n18623 = ~n18612 & ~n18622;
  assign n18624 = ~n16124 & n18623;
  assign n18625 = n16124 & n18375;
  assign n18626 = ~n18624 & ~n18625;
  assign n18627 = pi647 & ~n18626;
  assign n18628 = pi628 & ~n18623;
  assign n18629 = ~n17182 & n18621;
  assign n18630 = ~pi625 & pi1153;
  assign n18631 = pi625 & ~pi1153;
  assign n18632 = ~n18630 & ~n18631;
  assign n18633 = pi778 & ~n18632;
  assign n18634 = n18197 & ~n18633;
  assign n18635 = ~n18375 & ~n18634;
  assign n18636 = ~n16593 & ~n18635;
  assign n18637 = ~n18375 & ~n18636;
  assign n18638 = ~n17340 & ~n18637;
  assign n18639 = ~n17342 & n18638;
  assign n18640 = n17350 & n18639;
  assign n18641 = ~n18629 & ~n18640;
  assign n18642 = pi788 & ~n18641;
  assign n18643 = pi618 & ~n18637;
  assign n18644 = pi609 & ~n18635;
  assign n18645 = pi625 & n18374;
  assign n18646 = ~n18377 & ~n18645;
  assign n18647 = ~pi1153 & ~n18646;
  assign n18648 = ~pi608 & ~n18647;
  assign n18649 = pi625 & n18197;
  assign n18650 = ~n18375 & ~n18649;
  assign n18651 = pi1153 & n18650;
  assign n18652 = n18648 & ~n18651;
  assign n18653 = ~n18037 & ~n18645;
  assign n18654 = pi1153 & ~n18653;
  assign n18655 = ~pi625 & ~pi1153;
  assign n18656 = n18197 & n18655;
  assign n18657 = ~n18375 & ~n18656;
  assign n18658 = ~n18654 & n18657;
  assign n18659 = pi608 & ~n18658;
  assign n18660 = ~n18652 & ~n18659;
  assign n18661 = pi778 & ~n18660;
  assign n18662 = ~pi778 & ~n18377;
  assign n18663 = ~n18661 & ~n18662;
  assign n18664 = ~pi609 & ~n18663;
  assign n18665 = ~pi1155 & ~n18664;
  assign n18666 = ~n18644 & n18665;
  assign n18667 = ~pi660 & ~n18579;
  assign n18668 = ~n18666 & n18667;
  assign n18669 = ~pi609 & ~n18635;
  assign n18670 = pi609 & ~n18663;
  assign n18671 = ~n18669 & ~n18670;
  assign n18672 = pi1155 & n18671;
  assign n18673 = ~n18582 & ~n18672;
  assign n18674 = pi660 & n18673;
  assign n18675 = ~n18668 & ~n18674;
  assign n18676 = pi785 & ~n18675;
  assign n18677 = ~pi785 & ~n18663;
  assign n18678 = ~n18676 & ~n18677;
  assign n18679 = ~pi618 & ~n18678;
  assign n18680 = ~pi1154 & ~n18679;
  assign n18681 = ~n18643 & n18680;
  assign n18682 = ~pi627 & ~n18592;
  assign n18683 = ~n18681 & n18682;
  assign n18684 = ~pi618 & ~n18637;
  assign n18685 = pi618 & ~n18678;
  assign n18686 = ~n18684 & ~n18685;
  assign n18687 = pi1154 & n18686;
  assign n18688 = ~n18596 & ~n18687;
  assign n18689 = pi627 & n18688;
  assign n18690 = ~n18683 & ~n18689;
  assign n18691 = pi781 & ~n18690;
  assign n18692 = ~pi781 & ~n18678;
  assign n18693 = ~n18691 & ~n18692;
  assign n18694 = ~pi619 & ~n18693;
  assign n18695 = pi619 & n18638;
  assign n18696 = ~pi1159 & ~n18695;
  assign n18697 = ~n18694 & n18696;
  assign n18698 = ~pi648 & ~n18697;
  assign n18699 = ~n18604 & n18698;
  assign n18700 = ~pi619 & n18638;
  assign n18701 = pi619 & ~n18693;
  assign n18702 = ~n18700 & ~n18701;
  assign n18703 = pi1159 & n18702;
  assign n18704 = ~n18608 & ~n18703;
  assign n18705 = pi648 & n18704;
  assign n18706 = ~n18699 & ~n18705;
  assign n18707 = pi789 & n18706;
  assign n18708 = ~pi789 & n18693;
  assign n18709 = n17356 & ~n18708;
  assign n18710 = ~n18707 & n18709;
  assign n18711 = ~n18642 & ~n18710;
  assign n18712 = ~pi628 & n18711;
  assign n18713 = ~pi1156 & ~n18712;
  assign n18714 = ~n18628 & n18713;
  assign n18715 = ~n16589 & ~n16593;
  assign n18716 = ~n17159 & n18715;
  assign n18717 = ~n17183 & n18716;
  assign n18718 = ~n18635 & n18717;
  assign n18719 = pi628 & n18718;
  assign n18720 = ~n18375 & ~n18719;
  assign n18721 = pi1156 & ~n18720;
  assign n18722 = ~pi629 & ~n18721;
  assign n18723 = ~n18714 & n18722;
  assign n18724 = ~pi628 & ~n18623;
  assign n18725 = pi628 & n18711;
  assign n18726 = ~n18724 & ~n18725;
  assign n18727 = pi1156 & n18726;
  assign n18728 = ~pi628 & n18718;
  assign n18729 = ~n18375 & ~n18728;
  assign n18730 = ~pi1156 & ~n18729;
  assign n18731 = pi629 & ~n18730;
  assign n18732 = ~n18727 & n18731;
  assign n18733 = ~n18723 & ~n18732;
  assign n18734 = pi792 & ~n18733;
  assign n18735 = ~pi792 & n18711;
  assign n18736 = ~n18734 & ~n18735;
  assign n18737 = ~pi647 & n18736;
  assign n18738 = ~pi1157 & ~n18737;
  assign n18739 = ~n18627 & n18738;
  assign n18740 = ~pi630 & ~n18739;
  assign n18741 = ~pi628 & ~pi1156;
  assign n18742 = pi628 & pi1156;
  assign n18743 = pi792 & ~n18742;
  assign n18744 = ~n18741 & n18743;
  assign n18745 = n18718 & ~n18744;
  assign n18746 = pi647 & n18745;
  assign n18747 = ~n18375 & ~n18746;
  assign n18748 = pi1157 & n18747;
  assign n18749 = n18740 & ~n18748;
  assign n18750 = ~pi647 & ~n18626;
  assign n18751 = pi647 & n18736;
  assign n18752 = ~n18750 & ~n18751;
  assign n18753 = pi1157 & n18752;
  assign n18754 = ~pi647 & n18745;
  assign n18755 = ~pi1157 & ~n18375;
  assign n18756 = ~n18754 & n18755;
  assign n18757 = pi630 & ~n18756;
  assign n18758 = ~n18753 & n18757;
  assign n18759 = ~n18749 & ~n18758;
  assign n18760 = pi787 & ~n18759;
  assign n18761 = ~pi787 & n18736;
  assign n18762 = ~n18760 & ~n18761;
  assign n18763 = pi644 & ~n18762;
  assign n18764 = ~pi647 & pi1157;
  assign n18765 = pi647 & ~pi1157;
  assign n18766 = ~n18764 & ~n18765;
  assign n18767 = pi787 & ~n18766;
  assign n18768 = n18745 & ~n18767;
  assign n18769 = ~n18375 & ~n18768;
  assign n18770 = ~pi644 & ~n18769;
  assign n18771 = pi715 & ~n18770;
  assign n18772 = ~n18763 & n18771;
  assign n18773 = n17247 & ~n18375;
  assign n18774 = ~n17247 & n18626;
  assign n18775 = ~n18773 & ~n18774;
  assign n18776 = pi644 & n18775;
  assign n18777 = ~pi644 & n18375;
  assign n18778 = ~pi715 & ~n18777;
  assign n18779 = ~n18776 & n18778;
  assign n18780 = pi1160 & ~n18779;
  assign n18781 = ~n18772 & n18780;
  assign n18782 = ~pi644 & n18775;
  assign n18783 = pi715 & ~n18782;
  assign n18784 = pi644 & n18375;
  assign n18785 = n18783 & ~n18784;
  assign n18786 = pi644 & ~n18769;
  assign n18787 = ~pi644 & ~n18762;
  assign n18788 = ~pi715 & ~n18787;
  assign n18789 = ~n18786 & n18788;
  assign n18790 = ~pi1160 & ~n18789;
  assign n18791 = ~n18785 & n18790;
  assign n18792 = ~n18781 & ~n18791;
  assign n18793 = pi790 & ~n18792;
  assign n18794 = ~pi790 & ~n18762;
  assign n18795 = pi832 & ~n18794;
  assign n18796 = ~n18793 & n18795;
  assign po299 = ~n18575 & ~n18796;
  assign n18798 = pi143 & ~n10020;
  assign n18799 = ~pi143 & ~n16526;
  assign n18800 = pi774 & ~n18799;
  assign n18801 = pi38 & n16524;
  assign n18802 = n16393 & n18801;
  assign n18803 = ~pi38 & n16503;
  assign n18804 = pi143 & ~n18803;
  assign n18805 = ~pi38 & ~n16449;
  assign n18806 = ~n16393 & n16508;
  assign n18807 = pi38 & ~n18806;
  assign n18808 = ~n18805 & ~n18807;
  assign n18809 = ~pi143 & ~pi774;
  assign n18810 = n18808 & n18809;
  assign n18811 = ~n18804 & ~n18810;
  assign n18812 = ~n18802 & ~n18811;
  assign n18813 = ~n18800 & ~n18812;
  assign n18814 = n10020 & ~n18813;
  assign n18815 = ~n18798 & ~n18814;
  assign n18816 = ~n16521 & ~n18815;
  assign n18817 = ~pi143 & ~n16527;
  assign n18818 = n16521 & ~n18817;
  assign n18819 = ~n18816 & ~n18818;
  assign n18820 = ~pi785 & ~n18819;
  assign n18821 = ~n16532 & ~n18817;
  assign n18822 = pi609 & n18816;
  assign n18823 = ~n18821 & ~n18822;
  assign n18824 = pi1155 & ~n18823;
  assign n18825 = ~n16537 & ~n18817;
  assign n18826 = ~pi609 & n18816;
  assign n18827 = ~n18825 & ~n18826;
  assign n18828 = ~pi1155 & ~n18827;
  assign n18829 = ~n18824 & ~n18828;
  assign n18830 = pi785 & ~n18829;
  assign n18831 = ~n18820 & ~n18830;
  assign n18832 = ~pi781 & ~n18831;
  assign n18833 = pi618 & n18831;
  assign n18834 = ~pi618 & n18817;
  assign n18835 = pi1154 & ~n18834;
  assign n18836 = ~n18833 & n18835;
  assign n18837 = ~pi618 & n18831;
  assign n18838 = pi618 & n18817;
  assign n18839 = ~pi1154 & ~n18838;
  assign n18840 = ~n18837 & n18839;
  assign n18841 = ~n18836 & ~n18840;
  assign n18842 = pi781 & ~n18841;
  assign n18843 = ~n18832 & ~n18842;
  assign n18844 = ~pi789 & ~n18843;
  assign n18845 = pi619 & n18843;
  assign n18846 = ~pi619 & n18817;
  assign n18847 = pi1159 & ~n18846;
  assign n18848 = ~n18845 & n18847;
  assign n18849 = ~pi619 & n18843;
  assign n18850 = pi619 & n18817;
  assign n18851 = ~pi1159 & ~n18850;
  assign n18852 = ~n18849 & n18851;
  assign n18853 = ~n18848 & ~n18852;
  assign n18854 = pi789 & ~n18853;
  assign n18855 = ~n18844 & ~n18854;
  assign n18856 = ~pi626 & n18855;
  assign n18857 = pi626 & n18817;
  assign n18858 = ~pi1158 & ~n18857;
  assign n18859 = ~n18856 & n18858;
  assign n18860 = pi626 & n18855;
  assign n18861 = ~pi626 & n18817;
  assign n18862 = pi1158 & ~n18861;
  assign n18863 = ~n18860 & n18862;
  assign n18864 = ~n18859 & ~n18863;
  assign n18865 = pi788 & ~n18864;
  assign n18866 = ~pi788 & ~n18855;
  assign n18867 = ~n18865 & ~n18866;
  assign n18868 = ~n16124 & n18867;
  assign n18869 = n16124 & n18817;
  assign n18870 = ~n18868 & ~n18869;
  assign n18871 = pi647 & ~n18870;
  assign n18872 = pi628 & n18867;
  assign n18873 = n16593 & ~n18817;
  assign n18874 = ~pi687 & n18799;
  assign n18875 = ~pi143 & ~n16508;
  assign n18876 = n16744 & ~n18875;
  assign n18877 = pi143 & n17589;
  assign n18878 = ~pi143 & n17592;
  assign n18879 = ~pi38 & ~n18878;
  assign n18880 = ~n18877 & n18879;
  assign n18881 = ~n18876 & ~n18880;
  assign n18882 = pi687 & n18881;
  assign n18883 = ~n18874 & ~n18882;
  assign n18884 = n10020 & n18883;
  assign n18885 = ~n18798 & ~n18884;
  assign n18886 = ~pi778 & ~n18885;
  assign n18887 = pi625 & n18885;
  assign n18888 = pi1153 & ~n18887;
  assign n18889 = ~pi625 & n18817;
  assign n18890 = n18888 & ~n18889;
  assign n18891 = ~pi625 & n18885;
  assign n18892 = ~pi1153 & ~n18891;
  assign n18893 = pi625 & n18817;
  assign n18894 = n18892 & ~n18893;
  assign n18895 = ~n18890 & ~n18894;
  assign n18896 = pi778 & ~n18895;
  assign n18897 = ~n18886 & ~n18896;
  assign n18898 = ~n16593 & ~n18897;
  assign n18899 = ~n18873 & ~n18898;
  assign n18900 = ~n16589 & n18899;
  assign n18901 = n16589 & n18817;
  assign n18902 = ~n18900 & ~n18901;
  assign n18903 = pi619 & ~n18902;
  assign n18904 = pi618 & n18899;
  assign n18905 = pi609 & n18897;
  assign n18906 = pi625 & n18815;
  assign n18907 = ~pi687 & n18813;
  assign n18908 = pi39 & ~n17051;
  assign n18909 = ~pi39 & n16917;
  assign n18910 = pi38 & ~n18909;
  assign n18911 = ~n18908 & ~n18910;
  assign n18912 = ~pi39 & ~n17067;
  assign n18913 = ~pi38 & n18912;
  assign n18914 = n18911 & ~n18913;
  assign n18915 = ~pi143 & ~n18914;
  assign n18916 = pi39 & ~n16998;
  assign n18917 = ~n16460 & n17587;
  assign n18918 = ~n18916 & ~n18917;
  assign n18919 = ~pi38 & ~n18918;
  assign n18920 = n16508 & ~n16916;
  assign n18921 = pi38 & ~n18920;
  assign n18922 = ~n18919 & ~n18921;
  assign n18923 = pi143 & n18922;
  assign n18924 = ~pi774 & ~n18923;
  assign n18925 = ~n18915 & n18924;
  assign n18926 = ~pi39 & ~n17058;
  assign n18927 = pi39 & ~n16935;
  assign n18928 = ~n18926 & ~n18927;
  assign n18929 = ~pi38 & n18928;
  assign n18930 = pi143 & n18929;
  assign n18931 = pi38 & ~pi39;
  assign n18932 = n17080 & n18931;
  assign n18933 = n16508 & ~n16814;
  assign n18934 = pi38 & n18933;
  assign n18935 = pi39 & ~n16853;
  assign n18936 = ~pi39 & ~n17061;
  assign n18937 = ~n18935 & ~n18936;
  assign n18938 = ~pi38 & ~n18937;
  assign n18939 = ~n18934 & ~n18938;
  assign n18940 = ~pi143 & n18939;
  assign n18941 = ~n18932 & ~n18940;
  assign n18942 = pi774 & n18941;
  assign n18943 = ~n18930 & n18942;
  assign n18944 = ~n18925 & ~n18943;
  assign n18945 = pi687 & n18944;
  assign n18946 = ~n18907 & ~n18945;
  assign n18947 = n10020 & n18946;
  assign n18948 = ~n18798 & ~n18947;
  assign n18949 = ~pi625 & n18948;
  assign n18950 = ~pi1153 & ~n18949;
  assign n18951 = ~n18906 & n18950;
  assign n18952 = ~pi608 & ~n18890;
  assign n18953 = ~n18951 & n18952;
  assign n18954 = ~pi625 & n18815;
  assign n18955 = pi625 & n18948;
  assign n18956 = ~n18954 & ~n18955;
  assign n18957 = pi1153 & n18956;
  assign n18958 = ~n18894 & ~n18957;
  assign n18959 = pi608 & n18958;
  assign n18960 = ~n18953 & ~n18959;
  assign n18961 = pi778 & ~n18960;
  assign n18962 = ~pi778 & n18948;
  assign n18963 = ~n18961 & ~n18962;
  assign n18964 = ~pi609 & ~n18963;
  assign n18965 = ~pi1155 & ~n18964;
  assign n18966 = ~n18905 & n18965;
  assign n18967 = ~pi660 & ~n18824;
  assign n18968 = ~n18966 & n18967;
  assign n18969 = ~pi609 & n18897;
  assign n18970 = pi609 & ~n18963;
  assign n18971 = ~n18969 & ~n18970;
  assign n18972 = pi1155 & n18971;
  assign n18973 = ~n18828 & ~n18972;
  assign n18974 = pi660 & n18973;
  assign n18975 = ~n18968 & ~n18974;
  assign n18976 = pi785 & ~n18975;
  assign n18977 = ~pi785 & ~n18963;
  assign n18978 = ~n18976 & ~n18977;
  assign n18979 = ~pi618 & ~n18978;
  assign n18980 = ~pi1154 & ~n18979;
  assign n18981 = ~n18904 & n18980;
  assign n18982 = ~pi627 & ~n18836;
  assign n18983 = ~n18981 & n18982;
  assign n18984 = ~pi618 & n18899;
  assign n18985 = pi618 & ~n18978;
  assign n18986 = ~n18984 & ~n18985;
  assign n18987 = pi1154 & n18986;
  assign n18988 = ~n18840 & ~n18987;
  assign n18989 = pi627 & n18988;
  assign n18990 = ~n18983 & ~n18989;
  assign n18991 = pi781 & ~n18990;
  assign n18992 = ~pi781 & ~n18978;
  assign n18993 = ~n18991 & ~n18992;
  assign n18994 = ~pi619 & ~n18993;
  assign n18995 = ~pi1159 & ~n18994;
  assign n18996 = ~n18903 & n18995;
  assign n18997 = ~pi648 & ~n18848;
  assign n18998 = ~n18996 & n18997;
  assign n18999 = ~pi619 & ~n18902;
  assign n19000 = pi619 & ~n18993;
  assign n19001 = ~n18999 & ~n19000;
  assign n19002 = pi1159 & n19001;
  assign n19003 = ~n18852 & ~n19002;
  assign n19004 = pi648 & n19003;
  assign n19005 = ~n18998 & ~n19004;
  assign n19006 = pi789 & ~n19005;
  assign n19007 = ~pi789 & ~n18993;
  assign n19008 = ~n19006 & ~n19007;
  assign n19009 = ~pi788 & n19008;
  assign n19010 = ~n17153 & ~n18859;
  assign n19011 = ~pi626 & n19008;
  assign n19012 = n17159 & ~n18817;
  assign n19013 = ~n17159 & n18902;
  assign n19014 = ~n19012 & ~n19013;
  assign n19015 = pi626 & ~n19014;
  assign n19016 = ~pi641 & ~n19015;
  assign n19017 = ~n19011 & n19016;
  assign n19018 = ~n19010 & ~n19017;
  assign n19019 = ~n17167 & ~n18863;
  assign n19020 = pi626 & n19008;
  assign n19021 = ~pi626 & ~n19014;
  assign n19022 = pi641 & ~n19021;
  assign n19023 = ~n19020 & n19022;
  assign n19024 = ~n19019 & ~n19023;
  assign n19025 = ~n19018 & ~n19024;
  assign n19026 = pi788 & ~n19025;
  assign n19027 = ~n19009 & ~n19026;
  assign n19028 = ~pi628 & n19027;
  assign n19029 = ~pi1156 & ~n19028;
  assign n19030 = ~n18872 & n19029;
  assign n19031 = ~n17183 & n19014;
  assign n19032 = n17183 & n18817;
  assign n19033 = ~n19031 & ~n19032;
  assign n19034 = pi628 & ~n19033;
  assign n19035 = pi1156 & ~n19034;
  assign n19036 = ~pi628 & n18817;
  assign n19037 = n19035 & ~n19036;
  assign n19038 = ~pi629 & ~n19037;
  assign n19039 = ~n19030 & n19038;
  assign n19040 = ~pi628 & ~n19033;
  assign n19041 = pi628 & n18817;
  assign n19042 = ~pi1156 & ~n19041;
  assign n19043 = ~n19040 & n19042;
  assign n19044 = ~pi628 & n18867;
  assign n19045 = pi628 & n19027;
  assign n19046 = ~n19044 & ~n19045;
  assign n19047 = pi1156 & n19046;
  assign n19048 = ~n19043 & ~n19047;
  assign n19049 = pi629 & n19048;
  assign n19050 = ~n19039 & ~n19049;
  assign n19051 = pi792 & ~n19050;
  assign n19052 = ~pi792 & n19027;
  assign n19053 = ~n19051 & ~n19052;
  assign n19054 = ~pi647 & ~n19053;
  assign n19055 = ~pi1157 & ~n19054;
  assign n19056 = ~n18871 & n19055;
  assign n19057 = ~pi792 & n19033;
  assign n19058 = ~n19037 & ~n19043;
  assign n19059 = pi792 & ~n19058;
  assign n19060 = ~n19057 & ~n19059;
  assign n19061 = pi647 & n19060;
  assign n19062 = pi1157 & ~n19061;
  assign n19063 = ~pi647 & n18817;
  assign n19064 = n19062 & ~n19063;
  assign n19065 = ~pi630 & ~n19064;
  assign n19066 = ~n19056 & n19065;
  assign n19067 = ~pi647 & n19060;
  assign n19068 = pi647 & n18817;
  assign n19069 = ~pi1157 & ~n19068;
  assign n19070 = ~n19067 & n19069;
  assign n19071 = ~pi647 & ~n18870;
  assign n19072 = pi647 & ~n19053;
  assign n19073 = ~n19071 & ~n19072;
  assign n19074 = pi1157 & n19073;
  assign n19075 = ~n19070 & ~n19074;
  assign n19076 = pi630 & n19075;
  assign n19077 = ~n19066 & ~n19076;
  assign n19078 = pi787 & ~n19077;
  assign n19079 = ~pi787 & ~n19053;
  assign n19080 = ~n19078 & ~n19079;
  assign n19081 = ~pi790 & n19080;
  assign n19082 = pi644 & ~n19080;
  assign n19083 = ~pi787 & ~n19060;
  assign n19084 = ~n19064 & ~n19070;
  assign n19085 = pi787 & ~n19084;
  assign n19086 = ~n19083 & ~n19085;
  assign n19087 = ~pi644 & n19086;
  assign n19088 = pi715 & ~n19087;
  assign n19089 = ~n19082 & n19088;
  assign n19090 = ~pi644 & n18817;
  assign n19091 = n17247 & ~n18817;
  assign n19092 = ~n17247 & n18870;
  assign n19093 = ~n19091 & ~n19092;
  assign n19094 = pi644 & n19093;
  assign n19095 = ~pi715 & ~n19094;
  assign n19096 = ~n19090 & n19095;
  assign n19097 = ~n19089 & ~n19096;
  assign n19098 = pi1160 & n19097;
  assign n19099 = ~pi644 & n19093;
  assign n19100 = pi715 & ~n19099;
  assign n19101 = pi644 & n18817;
  assign n19102 = n19100 & ~n19101;
  assign n19103 = pi644 & n19086;
  assign n19104 = ~pi644 & ~n19080;
  assign n19105 = ~pi715 & ~n19104;
  assign n19106 = ~n19103 & n19105;
  assign n19107 = ~n19102 & ~n19106;
  assign n19108 = ~pi1160 & n19107;
  assign n19109 = ~n19098 & ~n19108;
  assign n19110 = pi790 & n19109;
  assign n19111 = ~n19081 & ~n19110;
  assign n19112 = ~po1038 & n19111;
  assign n19113 = ~pi143 & po1038;
  assign n19114 = ~pi832 & ~n19113;
  assign n19115 = ~n19112 & n19114;
  assign n19116 = ~pi143 & ~n2934;
  assign n19117 = ~pi774 & n16510;
  assign n19118 = ~n19116 & ~n19117;
  assign n19119 = ~n17273 & ~n19118;
  assign n19120 = ~pi785 & ~n19119;
  assign n19121 = ~n17279 & ~n19118;
  assign n19122 = pi1155 & ~n19121;
  assign n19123 = ~n17282 & n19119;
  assign n19124 = ~pi1155 & ~n19123;
  assign n19125 = ~n19122 & ~n19124;
  assign n19126 = pi785 & ~n19125;
  assign n19127 = ~n19120 & ~n19126;
  assign n19128 = ~pi781 & ~n19127;
  assign n19129 = ~n17289 & n19127;
  assign n19130 = pi1154 & ~n19129;
  assign n19131 = ~n17292 & n19127;
  assign n19132 = ~pi1154 & ~n19131;
  assign n19133 = ~n19130 & ~n19132;
  assign n19134 = pi781 & ~n19133;
  assign n19135 = ~n19128 & ~n19134;
  assign n19136 = ~pi789 & ~n19135;
  assign n19137 = pi619 & n19135;
  assign n19138 = ~pi619 & n19116;
  assign n19139 = pi1159 & ~n19138;
  assign n19140 = ~n19137 & n19139;
  assign n19141 = ~pi619 & n19135;
  assign n19142 = pi619 & n19116;
  assign n19143 = ~pi1159 & ~n19142;
  assign n19144 = ~n19141 & n19143;
  assign n19145 = ~n19140 & ~n19144;
  assign n19146 = pi789 & ~n19145;
  assign n19147 = ~n19136 & ~n19146;
  assign n19148 = ~pi788 & ~n19147;
  assign n19149 = pi626 & n19147;
  assign n19150 = ~pi626 & n19116;
  assign n19151 = pi1158 & ~n19150;
  assign n19152 = ~n19149 & n19151;
  assign n19153 = ~pi626 & n19147;
  assign n19154 = pi626 & n19116;
  assign n19155 = ~pi1158 & ~n19154;
  assign n19156 = ~n19153 & n19155;
  assign n19157 = ~n19152 & ~n19156;
  assign n19158 = pi788 & ~n19157;
  assign n19159 = ~n19148 & ~n19158;
  assign n19160 = ~n16124 & n19159;
  assign n19161 = n16124 & n19116;
  assign n19162 = ~n19160 & ~n19161;
  assign n19163 = pi647 & ~n19162;
  assign n19164 = pi628 & n19159;
  assign n19165 = pi687 & n16742;
  assign n19166 = ~n19116 & ~n19165;
  assign n19167 = ~pi778 & n19166;
  assign n19168 = ~pi625 & n19165;
  assign n19169 = ~n19166 & ~n19168;
  assign n19170 = pi1153 & ~n19169;
  assign n19171 = ~pi1153 & ~n19116;
  assign n19172 = ~n19168 & n19171;
  assign n19173 = ~n19170 & ~n19172;
  assign n19174 = pi778 & ~n19173;
  assign n19175 = ~n19167 & ~n19174;
  assign n19176 = ~n17338 & n19175;
  assign n19177 = ~n17340 & n19176;
  assign n19178 = ~n17342 & n19177;
  assign n19179 = n17350 & n19178;
  assign n19180 = ~n17182 & n19157;
  assign n19181 = ~n19179 & ~n19180;
  assign n19182 = pi788 & ~n19181;
  assign n19183 = pi618 & n19176;
  assign n19184 = pi609 & n19175;
  assign n19185 = ~n16393 & ~n19166;
  assign n19186 = pi625 & n19185;
  assign n19187 = n19118 & ~n19185;
  assign n19188 = ~n19186 & ~n19187;
  assign n19189 = n19171 & ~n19188;
  assign n19190 = ~pi608 & ~n19170;
  assign n19191 = ~n19189 & n19190;
  assign n19192 = pi1153 & ~n19186;
  assign n19193 = n19118 & n19192;
  assign n19194 = ~n19172 & ~n19193;
  assign n19195 = pi608 & n19194;
  assign n19196 = ~n19191 & ~n19195;
  assign n19197 = pi778 & ~n19196;
  assign n19198 = ~pi778 & ~n19187;
  assign n19199 = ~n19197 & ~n19198;
  assign n19200 = ~pi609 & ~n19199;
  assign n19201 = ~pi1155 & ~n19200;
  assign n19202 = ~n19184 & n19201;
  assign n19203 = ~pi660 & ~n19122;
  assign n19204 = ~n19202 & n19203;
  assign n19205 = ~pi609 & n19175;
  assign n19206 = pi609 & ~n19199;
  assign n19207 = ~n19205 & ~n19206;
  assign n19208 = pi1155 & n19207;
  assign n19209 = ~n19124 & ~n19208;
  assign n19210 = pi660 & n19209;
  assign n19211 = ~n19204 & ~n19210;
  assign n19212 = pi785 & ~n19211;
  assign n19213 = ~pi785 & ~n19199;
  assign n19214 = ~n19212 & ~n19213;
  assign n19215 = ~pi618 & ~n19214;
  assign n19216 = ~pi1154 & ~n19215;
  assign n19217 = ~n19183 & n19216;
  assign n19218 = ~pi627 & ~n19130;
  assign n19219 = ~n19217 & n19218;
  assign n19220 = ~pi618 & n19176;
  assign n19221 = pi618 & ~n19214;
  assign n19222 = ~n19220 & ~n19221;
  assign n19223 = pi1154 & n19222;
  assign n19224 = ~n19132 & ~n19223;
  assign n19225 = pi627 & n19224;
  assign n19226 = ~n19219 & ~n19225;
  assign n19227 = pi781 & ~n19226;
  assign n19228 = ~pi781 & ~n19214;
  assign n19229 = ~n19227 & ~n19228;
  assign n19230 = ~pi619 & ~n19229;
  assign n19231 = pi619 & n19177;
  assign n19232 = ~pi1159 & ~n19231;
  assign n19233 = ~n19230 & n19232;
  assign n19234 = ~pi648 & ~n19233;
  assign n19235 = ~n19140 & n19234;
  assign n19236 = ~pi619 & n19177;
  assign n19237 = pi619 & ~n19229;
  assign n19238 = ~n19236 & ~n19237;
  assign n19239 = pi1159 & n19238;
  assign n19240 = ~n19144 & ~n19239;
  assign n19241 = pi648 & n19240;
  assign n19242 = ~n19235 & ~n19241;
  assign n19243 = pi789 & n19242;
  assign n19244 = ~pi789 & n19229;
  assign n19245 = n17356 & ~n19244;
  assign n19246 = ~n19243 & n19245;
  assign n19247 = ~n19182 & ~n19246;
  assign n19248 = ~pi628 & ~n19247;
  assign n19249 = ~pi1156 & ~n19248;
  assign n19250 = ~n19164 & n19249;
  assign n19251 = ~n17425 & n19178;
  assign n19252 = ~n17427 & n19251;
  assign n19253 = pi1156 & ~n19252;
  assign n19254 = ~pi629 & ~n19253;
  assign n19255 = ~n19250 & n19254;
  assign n19256 = ~pi628 & n19159;
  assign n19257 = pi628 & ~n19247;
  assign n19258 = ~n19256 & ~n19257;
  assign n19259 = pi1156 & n19258;
  assign n19260 = ~n17436 & n19251;
  assign n19261 = ~pi1156 & ~n19260;
  assign n19262 = pi629 & ~n19261;
  assign n19263 = ~n19259 & n19262;
  assign n19264 = ~n19255 & ~n19263;
  assign n19265 = pi792 & ~n19264;
  assign n19266 = ~pi792 & ~n19247;
  assign n19267 = ~n19265 & ~n19266;
  assign n19268 = ~pi647 & ~n19267;
  assign n19269 = ~pi1157 & ~n19268;
  assign n19270 = ~n19163 & n19269;
  assign n19271 = ~n17452 & n19251;
  assign n19272 = pi647 & n19271;
  assign n19273 = ~pi647 & n19116;
  assign n19274 = pi1157 & ~n19273;
  assign n19275 = ~n19272 & n19274;
  assign n19276 = ~pi630 & ~n19275;
  assign n19277 = ~n19270 & n19276;
  assign n19278 = ~pi647 & n19271;
  assign n19279 = pi647 & n19116;
  assign n19280 = ~pi1157 & ~n19279;
  assign n19281 = ~n19278 & n19280;
  assign n19282 = ~pi647 & ~n19162;
  assign n19283 = pi647 & ~n19267;
  assign n19284 = ~n19282 & ~n19283;
  assign n19285 = pi1157 & n19284;
  assign n19286 = ~n19281 & ~n19285;
  assign n19287 = pi630 & n19286;
  assign n19288 = ~n19277 & ~n19287;
  assign n19289 = pi787 & ~n19288;
  assign n19290 = ~pi787 & ~n19267;
  assign n19291 = ~n19289 & ~n19290;
  assign n19292 = pi644 & ~n19291;
  assign n19293 = ~pi787 & ~n19271;
  assign n19294 = ~n19275 & ~n19281;
  assign n19295 = pi787 & ~n19294;
  assign n19296 = ~n19293 & ~n19295;
  assign n19297 = ~pi644 & n19296;
  assign n19298 = pi715 & ~n19297;
  assign n19299 = ~n19292 & n19298;
  assign n19300 = n17247 & ~n19116;
  assign n19301 = ~n17247 & n19162;
  assign n19302 = ~n19300 & ~n19301;
  assign n19303 = pi644 & n19302;
  assign n19304 = ~pi644 & n19116;
  assign n19305 = ~pi715 & ~n19304;
  assign n19306 = ~n19303 & n19305;
  assign n19307 = pi1160 & ~n19306;
  assign n19308 = ~n19299 & n19307;
  assign n19309 = ~pi644 & n19302;
  assign n19310 = pi715 & ~n19309;
  assign n19311 = pi644 & n19116;
  assign n19312 = n19310 & ~n19311;
  assign n19313 = pi644 & n19296;
  assign n19314 = ~pi644 & ~n19291;
  assign n19315 = ~pi715 & ~n19314;
  assign n19316 = ~n19313 & n19315;
  assign n19317 = ~pi1160 & ~n19316;
  assign n19318 = ~n19312 & n19317;
  assign n19319 = ~n19308 & ~n19318;
  assign n19320 = pi790 & ~n19319;
  assign n19321 = ~pi790 & ~n19291;
  assign n19322 = pi832 & ~n19321;
  assign n19323 = ~n19320 & n19322;
  assign po300 = ~n19115 & ~n19323;
  assign n19325 = ~pi144 & ~n6274;
  assign n19326 = pi144 & ~n10020;
  assign n19327 = ~pi758 & ~n16355;
  assign n19328 = pi758 & n16447;
  assign n19329 = ~n19327 & ~n19328;
  assign n19330 = pi39 & ~n19329;
  assign n19331 = pi758 & n16380;
  assign n19332 = ~pi758 & n16201;
  assign n19333 = ~pi39 & ~n19332;
  assign n19334 = ~n19331 & n19333;
  assign n19335 = ~n19330 & ~n19334;
  assign n19336 = pi144 & ~n19335;
  assign n19337 = ~pi144 & pi758;
  assign n19338 = n16503 & n19337;
  assign n19339 = ~n19336 & ~n19338;
  assign n19340 = ~pi38 & ~n19339;
  assign n19341 = pi758 & n16393;
  assign n19342 = n16508 & ~n19341;
  assign n19343 = ~pi144 & ~n16508;
  assign n19344 = pi38 & ~n19343;
  assign n19345 = ~n19342 & n19344;
  assign n19346 = ~n19340 & ~n19345;
  assign n19347 = n10020 & ~n19346;
  assign n19348 = ~n19326 & ~n19347;
  assign n19349 = ~n16521 & ~n19348;
  assign n19350 = pi144 & ~n16527;
  assign n19351 = n16521 & n19350;
  assign n19352 = ~n19349 & ~n19351;
  assign n19353 = ~pi785 & ~n19352;
  assign n19354 = pi609 & n19352;
  assign n19355 = ~pi609 & ~n19350;
  assign n19356 = pi1155 & ~n19355;
  assign n19357 = ~n19354 & n19356;
  assign n19358 = ~pi609 & n19352;
  assign n19359 = pi609 & ~n19350;
  assign n19360 = ~pi1155 & ~n19359;
  assign n19361 = ~n19358 & n19360;
  assign n19362 = ~n19357 & ~n19361;
  assign n19363 = pi785 & ~n19362;
  assign n19364 = ~n19353 & ~n19363;
  assign n19365 = ~pi781 & ~n19364;
  assign n19366 = pi618 & n19364;
  assign n19367 = ~pi618 & ~n19350;
  assign n19368 = pi1154 & ~n19367;
  assign n19369 = ~n19366 & n19368;
  assign n19370 = ~pi618 & n19364;
  assign n19371 = pi618 & ~n19350;
  assign n19372 = ~pi1154 & ~n19371;
  assign n19373 = ~n19370 & n19372;
  assign n19374 = ~n19369 & ~n19373;
  assign n19375 = pi781 & ~n19374;
  assign n19376 = ~n19365 & ~n19375;
  assign n19377 = ~pi789 & ~n19376;
  assign n19378 = pi619 & n19376;
  assign n19379 = ~pi619 & ~n19350;
  assign n19380 = pi1159 & ~n19379;
  assign n19381 = ~n19378 & n19380;
  assign n19382 = ~pi619 & n19376;
  assign n19383 = pi619 & ~n19350;
  assign n19384 = ~pi1159 & ~n19383;
  assign n19385 = ~n19382 & n19384;
  assign n19386 = ~n19381 & ~n19385;
  assign n19387 = pi789 & ~n19386;
  assign n19388 = ~n19377 & ~n19387;
  assign n19389 = ~pi626 & n19388;
  assign n19390 = pi626 & ~n19350;
  assign n19391 = ~pi1158 & ~n19390;
  assign n19392 = ~n19389 & n19391;
  assign n19393 = pi626 & n19388;
  assign n19394 = ~pi626 & ~n19350;
  assign n19395 = pi1158 & ~n19394;
  assign n19396 = ~n19393 & n19395;
  assign n19397 = ~n19392 & ~n19396;
  assign n19398 = pi788 & ~n19397;
  assign n19399 = ~pi788 & ~n19388;
  assign n19400 = ~n19398 & ~n19399;
  assign n19401 = ~n16124 & ~n19400;
  assign n19402 = n16124 & n19350;
  assign n19403 = ~n19401 & ~n19402;
  assign n19404 = pi647 & n19403;
  assign n19405 = pi628 & n19400;
  assign n19406 = n16593 & ~n19350;
  assign n19407 = pi736 & n10020;
  assign n19408 = ~n19350 & ~n19407;
  assign n19409 = n6097 & n16665;
  assign n19410 = pi38 & ~n19409;
  assign n19411 = ~n19343 & n19410;
  assign n19412 = pi144 & ~n17592;
  assign n19413 = ~pi144 & ~n17589;
  assign n19414 = ~pi38 & ~n19413;
  assign n19415 = ~n19412 & n19414;
  assign n19416 = ~n19411 & ~n19415;
  assign n19417 = n19407 & n19416;
  assign n19418 = ~n19408 & ~n19417;
  assign n19419 = ~pi778 & n19418;
  assign n19420 = pi625 & ~n19418;
  assign n19421 = ~pi625 & ~n19350;
  assign n19422 = pi1153 & ~n19421;
  assign n19423 = ~n19420 & n19422;
  assign n19424 = ~pi625 & ~n19418;
  assign n19425 = pi625 & ~n19350;
  assign n19426 = ~pi1153 & ~n19425;
  assign n19427 = ~n19424 & n19426;
  assign n19428 = ~n19423 & ~n19427;
  assign n19429 = pi778 & ~n19428;
  assign n19430 = ~n19419 & ~n19429;
  assign n19431 = ~n16593 & n19430;
  assign n19432 = ~n19406 & ~n19431;
  assign n19433 = ~n16589 & n19432;
  assign n19434 = n16589 & n19350;
  assign n19435 = ~n19433 & ~n19434;
  assign n19436 = pi619 & n19435;
  assign n19437 = pi618 & ~n19432;
  assign n19438 = pi609 & n19430;
  assign n19439 = pi625 & n19348;
  assign n19440 = ~n19347 & ~n19407;
  assign n19441 = pi144 & ~n17061;
  assign n19442 = ~pi144 & ~n17058;
  assign n19443 = ~pi758 & ~n19442;
  assign n19444 = ~n19441 & n19443;
  assign n19445 = ~pi144 & n17065;
  assign n19446 = pi144 & n17067;
  assign n19447 = ~n19445 & ~n19446;
  assign n19448 = pi758 & n19447;
  assign n19449 = ~pi39 & ~n19448;
  assign n19450 = ~n19444 & n19449;
  assign n19451 = ~pi144 & ~n16998;
  assign n19452 = pi758 & ~n19451;
  assign n19453 = pi144 & n17051;
  assign n19454 = n19452 & ~n19453;
  assign n19455 = ~pi144 & ~n16935;
  assign n19456 = pi144 & ~n16853;
  assign n19457 = ~pi758 & ~n19456;
  assign n19458 = ~n19455 & n19457;
  assign n19459 = pi39 & ~n19458;
  assign n19460 = ~n19454 & n19459;
  assign n19461 = ~pi38 & ~n19460;
  assign n19462 = ~n19450 & n19461;
  assign n19463 = pi736 & ~n19462;
  assign n19464 = ~n18932 & n19463;
  assign n19465 = ~n19345 & n19464;
  assign n19466 = ~n19440 & ~n19465;
  assign n19467 = ~n19326 & ~n19466;
  assign n19468 = ~pi625 & n19467;
  assign n19469 = ~pi1153 & ~n19468;
  assign n19470 = ~n19439 & n19469;
  assign n19471 = ~pi608 & ~n19423;
  assign n19472 = ~n19470 & n19471;
  assign n19473 = ~pi625 & n19348;
  assign n19474 = pi625 & n19467;
  assign n19475 = ~n19473 & ~n19474;
  assign n19476 = pi1153 & n19475;
  assign n19477 = ~n19427 & ~n19476;
  assign n19478 = pi608 & n19477;
  assign n19479 = ~n19472 & ~n19478;
  assign n19480 = pi778 & ~n19479;
  assign n19481 = ~pi778 & n19467;
  assign n19482 = ~n19480 & ~n19481;
  assign n19483 = ~pi609 & ~n19482;
  assign n19484 = ~pi1155 & ~n19483;
  assign n19485 = ~n19438 & n19484;
  assign n19486 = ~pi660 & ~n19357;
  assign n19487 = ~n19485 & n19486;
  assign n19488 = ~pi609 & n19430;
  assign n19489 = pi609 & ~n19482;
  assign n19490 = ~n19488 & ~n19489;
  assign n19491 = pi1155 & n19490;
  assign n19492 = ~n19361 & ~n19491;
  assign n19493 = pi660 & n19492;
  assign n19494 = ~n19487 & ~n19493;
  assign n19495 = pi785 & ~n19494;
  assign n19496 = ~pi785 & ~n19482;
  assign n19497 = ~n19495 & ~n19496;
  assign n19498 = ~pi618 & ~n19497;
  assign n19499 = ~pi1154 & ~n19498;
  assign n19500 = ~n19437 & n19499;
  assign n19501 = ~pi627 & ~n19369;
  assign n19502 = ~n19500 & n19501;
  assign n19503 = ~pi618 & ~n19432;
  assign n19504 = pi618 & ~n19497;
  assign n19505 = ~n19503 & ~n19504;
  assign n19506 = pi1154 & n19505;
  assign n19507 = ~n19373 & ~n19506;
  assign n19508 = pi627 & n19507;
  assign n19509 = ~n19502 & ~n19508;
  assign n19510 = pi781 & ~n19509;
  assign n19511 = ~pi781 & ~n19497;
  assign n19512 = ~n19510 & ~n19511;
  assign n19513 = ~pi619 & ~n19512;
  assign n19514 = ~pi1159 & ~n19513;
  assign n19515 = ~n19436 & n19514;
  assign n19516 = ~pi648 & ~n19381;
  assign n19517 = ~n19515 & n19516;
  assign n19518 = ~pi619 & n19435;
  assign n19519 = pi619 & ~n19512;
  assign n19520 = ~n19518 & ~n19519;
  assign n19521 = pi1159 & n19520;
  assign n19522 = ~n19385 & ~n19521;
  assign n19523 = pi648 & n19522;
  assign n19524 = ~n19517 & ~n19523;
  assign n19525 = pi789 & ~n19524;
  assign n19526 = ~pi789 & ~n19512;
  assign n19527 = ~n19525 & ~n19526;
  assign n19528 = ~pi788 & n19527;
  assign n19529 = ~n17153 & ~n19392;
  assign n19530 = ~pi626 & n19527;
  assign n19531 = n17159 & ~n19350;
  assign n19532 = ~n17159 & n19435;
  assign n19533 = ~n19531 & ~n19532;
  assign n19534 = pi626 & n19533;
  assign n19535 = ~pi641 & ~n19534;
  assign n19536 = ~n19530 & n19535;
  assign n19537 = ~n19529 & ~n19536;
  assign n19538 = ~n17167 & ~n19396;
  assign n19539 = pi626 & n19527;
  assign n19540 = ~pi626 & n19533;
  assign n19541 = pi641 & ~n19540;
  assign n19542 = ~n19539 & n19541;
  assign n19543 = ~n19538 & ~n19542;
  assign n19544 = ~n19537 & ~n19543;
  assign n19545 = pi788 & ~n19544;
  assign n19546 = ~n19528 & ~n19545;
  assign n19547 = ~pi628 & n19546;
  assign n19548 = ~pi1156 & ~n19547;
  assign n19549 = ~n19405 & n19548;
  assign n19550 = ~n17183 & n19533;
  assign n19551 = n17183 & n19350;
  assign n19552 = ~n19550 & ~n19551;
  assign n19553 = pi628 & n19552;
  assign n19554 = ~pi628 & ~n19350;
  assign n19555 = pi1156 & ~n19554;
  assign n19556 = ~n19553 & n19555;
  assign n19557 = ~pi629 & ~n19556;
  assign n19558 = ~n19549 & n19557;
  assign n19559 = ~pi628 & n19552;
  assign n19560 = pi628 & ~n19350;
  assign n19561 = ~pi1156 & ~n19560;
  assign n19562 = ~n19559 & n19561;
  assign n19563 = ~pi628 & n19400;
  assign n19564 = pi628 & n19546;
  assign n19565 = ~n19563 & ~n19564;
  assign n19566 = pi1156 & n19565;
  assign n19567 = ~n19562 & ~n19566;
  assign n19568 = pi629 & n19567;
  assign n19569 = ~n19558 & ~n19568;
  assign n19570 = pi792 & ~n19569;
  assign n19571 = ~pi792 & n19546;
  assign n19572 = ~n19570 & ~n19571;
  assign n19573 = ~pi647 & ~n19572;
  assign n19574 = ~pi1157 & ~n19573;
  assign n19575 = ~n19404 & n19574;
  assign n19576 = ~pi792 & ~n19552;
  assign n19577 = ~n19556 & ~n19562;
  assign n19578 = pi792 & ~n19577;
  assign n19579 = ~n19576 & ~n19578;
  assign n19580 = pi647 & n19579;
  assign n19581 = ~pi647 & ~n19350;
  assign n19582 = pi1157 & ~n19581;
  assign n19583 = ~n19580 & n19582;
  assign n19584 = ~pi630 & ~n19583;
  assign n19585 = ~n19575 & n19584;
  assign n19586 = ~pi647 & n19579;
  assign n19587 = pi647 & ~n19350;
  assign n19588 = ~pi1157 & ~n19587;
  assign n19589 = ~n19586 & n19588;
  assign n19590 = ~pi647 & n19403;
  assign n19591 = pi647 & ~n19572;
  assign n19592 = ~n19590 & ~n19591;
  assign n19593 = pi1157 & n19592;
  assign n19594 = ~n19589 & ~n19593;
  assign n19595 = pi630 & n19594;
  assign n19596 = ~n19585 & ~n19595;
  assign n19597 = pi787 & ~n19596;
  assign n19598 = ~pi787 & ~n19572;
  assign n19599 = ~n19597 & ~n19598;
  assign n19600 = ~pi790 & n19599;
  assign n19601 = pi644 & ~n19599;
  assign n19602 = ~pi787 & ~n19579;
  assign n19603 = ~n19583 & ~n19589;
  assign n19604 = pi787 & ~n19603;
  assign n19605 = ~n19602 & ~n19604;
  assign n19606 = ~pi644 & n19605;
  assign n19607 = pi715 & ~n19606;
  assign n19608 = ~n19601 & n19607;
  assign n19609 = ~pi644 & ~n19350;
  assign n19610 = n17247 & ~n19350;
  assign n19611 = ~n17247 & n19403;
  assign n19612 = ~n19610 & ~n19611;
  assign n19613 = pi644 & ~n19612;
  assign n19614 = ~pi715 & ~n19613;
  assign n19615 = ~n19609 & n19614;
  assign n19616 = ~n19608 & ~n19615;
  assign n19617 = pi1160 & n19616;
  assign n19618 = pi644 & ~n19350;
  assign n19619 = ~pi644 & ~n19612;
  assign n19620 = pi715 & ~n19619;
  assign n19621 = ~n19618 & n19620;
  assign n19622 = pi644 & n19605;
  assign n19623 = ~pi644 & ~n19599;
  assign n19624 = ~pi715 & ~n19623;
  assign n19625 = ~n19622 & n19624;
  assign n19626 = ~n19621 & ~n19625;
  assign n19627 = ~pi1160 & n19626;
  assign n19628 = ~n19617 & ~n19627;
  assign n19629 = pi790 & n19628;
  assign n19630 = ~n19600 & ~n19629;
  assign n19631 = n6274 & n19630;
  assign n19632 = ~pi57 & ~n19631;
  assign n19633 = ~n19325 & n19632;
  assign n19634 = pi57 & pi144;
  assign n19635 = ~pi832 & ~n19634;
  assign n19636 = ~n19633 & n19635;
  assign n19637 = ~n17247 & ~n18767;
  assign n19638 = pi144 & ~n2934;
  assign n19639 = pi736 & n16742;
  assign n19640 = ~n19638 & ~n19639;
  assign n19641 = ~pi778 & n19640;
  assign n19642 = pi625 & n19639;
  assign n19643 = ~n19640 & ~n19642;
  assign n19644 = ~pi1153 & ~n19643;
  assign n19645 = pi1153 & ~n19638;
  assign n19646 = ~n19642 & n19645;
  assign n19647 = ~n19644 & ~n19646;
  assign n19648 = pi778 & ~n19647;
  assign n19649 = ~n19641 & ~n19648;
  assign n19650 = n18717 & n19649;
  assign n19651 = ~pi628 & n19650;
  assign n19652 = pi629 & ~n19651;
  assign n19653 = pi609 & pi1155;
  assign n19654 = ~pi609 & ~pi1155;
  assign n19655 = pi785 & ~n19654;
  assign n19656 = ~n19653 & n19655;
  assign n19657 = pi758 & n16510;
  assign n19658 = ~n19656 & n19657;
  assign n19659 = pi618 & pi1154;
  assign n19660 = ~pi618 & ~pi1154;
  assign n19661 = pi781 & ~n19660;
  assign n19662 = ~n19659 & n19661;
  assign n19663 = n19658 & ~n19662;
  assign n19664 = ~pi619 & pi1159;
  assign n19665 = pi619 & ~pi1159;
  assign n19666 = ~n19664 & ~n19665;
  assign n19667 = pi789 & ~n19666;
  assign n19668 = ~n16521 & ~n19667;
  assign n19669 = n19663 & n19668;
  assign n19670 = ~n17355 & n19669;
  assign n19671 = pi628 & ~n19670;
  assign n19672 = ~n19652 & ~n19671;
  assign n19673 = ~pi1156 & ~n19672;
  assign n19674 = pi628 & n19650;
  assign n19675 = ~pi628 & ~n19670;
  assign n19676 = pi629 & ~n19675;
  assign n19677 = pi1156 & ~n19676;
  assign n19678 = ~n19674 & n19677;
  assign n19679 = ~n19673 & ~n19678;
  assign n19680 = ~n19638 & ~n19679;
  assign n19681 = pi792 & n19680;
  assign n19682 = ~pi626 & n19669;
  assign n19683 = ~n19638 & ~n19682;
  assign n19684 = ~pi1158 & ~n19683;
  assign n19685 = n18715 & n19649;
  assign n19686 = ~n19638 & ~n19685;
  assign n19687 = n17159 & ~n19638;
  assign n19688 = ~n19686 & ~n19687;
  assign n19689 = n17344 & n19688;
  assign n19690 = pi641 & ~n19689;
  assign n19691 = ~n19684 & n19690;
  assign n19692 = pi626 & n19669;
  assign n19693 = ~n19638 & ~n19692;
  assign n19694 = pi1158 & ~n19693;
  assign n19695 = n17345 & n19688;
  assign n19696 = ~pi641 & ~n19695;
  assign n19697 = ~n19694 & n19696;
  assign n19698 = pi788 & ~n19697;
  assign n19699 = ~n19691 & n19698;
  assign n19700 = ~pi619 & ~n19686;
  assign n19701 = ~n17338 & n19649;
  assign n19702 = pi618 & n19701;
  assign n19703 = pi609 & n19649;
  assign n19704 = ~n19638 & ~n19657;
  assign n19705 = ~n16393 & n19639;
  assign n19706 = n19704 & ~n19705;
  assign n19707 = pi625 & n19705;
  assign n19708 = ~n19706 & ~n19707;
  assign n19709 = ~pi1153 & ~n19708;
  assign n19710 = ~pi608 & ~n19646;
  assign n19711 = ~n19709 & n19710;
  assign n19712 = pi1153 & ~n19707;
  assign n19713 = n19704 & n19712;
  assign n19714 = ~n19644 & ~n19713;
  assign n19715 = pi608 & n19714;
  assign n19716 = ~n19711 & ~n19715;
  assign n19717 = pi778 & ~n19716;
  assign n19718 = ~pi778 & ~n19706;
  assign n19719 = ~n19717 & ~n19718;
  assign n19720 = ~pi609 & ~n19719;
  assign n19721 = ~pi1155 & ~n19720;
  assign n19722 = ~n19703 & n19721;
  assign n19723 = ~n17279 & ~n19704;
  assign n19724 = pi1155 & ~n19723;
  assign n19725 = ~pi660 & ~n19724;
  assign n19726 = ~n19722 & n19725;
  assign n19727 = ~pi609 & n19649;
  assign n19728 = pi609 & ~n19719;
  assign n19729 = ~n19727 & ~n19728;
  assign n19730 = pi1155 & n19729;
  assign n19731 = ~pi1155 & ~n19638;
  assign n19732 = n16537 & n19657;
  assign n19733 = n19731 & ~n19732;
  assign n19734 = pi660 & ~n19733;
  assign n19735 = ~n19730 & n19734;
  assign n19736 = ~n19726 & ~n19735;
  assign n19737 = pi785 & ~n19736;
  assign n19738 = ~pi785 & ~n19719;
  assign n19739 = ~n19737 & ~n19738;
  assign n19740 = ~pi618 & ~n19739;
  assign n19741 = ~pi1154 & ~n19740;
  assign n19742 = ~n19702 & n19741;
  assign n19743 = ~pi627 & ~n19742;
  assign n19744 = pi618 & ~n16521;
  assign n19745 = n19658 & n19744;
  assign n19746 = ~n19638 & ~n19745;
  assign n19747 = pi1154 & n19746;
  assign n19748 = n19743 & ~n19747;
  assign n19749 = ~pi618 & n19701;
  assign n19750 = pi618 & ~n19739;
  assign n19751 = ~n19749 & ~n19750;
  assign n19752 = pi1154 & n19751;
  assign n19753 = ~pi618 & ~n16521;
  assign n19754 = n19658 & n19753;
  assign n19755 = ~pi1154 & ~n19638;
  assign n19756 = ~n19754 & n19755;
  assign n19757 = pi627 & ~n19756;
  assign n19758 = ~n19752 & n19757;
  assign n19759 = ~n19748 & ~n19758;
  assign n19760 = pi781 & ~n19759;
  assign n19761 = ~pi781 & ~n19739;
  assign n19762 = ~n19760 & ~n19761;
  assign n19763 = pi619 & ~n19762;
  assign n19764 = ~n19700 & ~n19763;
  assign n19765 = pi1159 & n19764;
  assign n19766 = ~pi619 & ~n16521;
  assign n19767 = n19663 & n19766;
  assign n19768 = ~pi1159 & ~n19638;
  assign n19769 = ~n19767 & n19768;
  assign n19770 = pi648 & ~n19769;
  assign n19771 = ~n19765 & n19770;
  assign n19772 = ~pi619 & ~n19762;
  assign n19773 = pi619 & ~n19686;
  assign n19774 = ~pi1159 & ~n19773;
  assign n19775 = ~n19772 & n19774;
  assign n19776 = pi619 & ~n16521;
  assign n19777 = n19663 & n19776;
  assign n19778 = ~n19638 & ~n19777;
  assign n19779 = pi1159 & n19778;
  assign n19780 = ~pi648 & ~n19779;
  assign n19781 = ~n19775 & n19780;
  assign n19782 = ~n19771 & ~n19781;
  assign n19783 = pi789 & n19782;
  assign n19784 = ~pi789 & n19762;
  assign n19785 = n17356 & ~n19784;
  assign n19786 = ~n19783 & n19785;
  assign n19787 = ~n19699 & ~n19786;
  assign n19788 = ~n16124 & ~n17451;
  assign n19789 = ~n19680 & ~n19788;
  assign n19790 = n19787 & ~n19789;
  assign n19791 = ~n19681 & ~n19790;
  assign n19792 = n19637 & ~n19791;
  assign n19793 = ~n16124 & n19670;
  assign n19794 = ~pi630 & n19793;
  assign n19795 = pi647 & ~n19794;
  assign n19796 = ~n18744 & n19650;
  assign n19797 = pi630 & ~n19796;
  assign n19798 = ~n19795 & ~n19797;
  assign n19799 = ~pi1157 & ~n19798;
  assign n19800 = ~pi630 & ~n19796;
  assign n19801 = pi647 & ~n19800;
  assign n19802 = pi630 & n19793;
  assign n19803 = pi1157 & ~n19802;
  assign n19804 = ~n19801 & n19803;
  assign n19805 = ~n19799 & ~n19804;
  assign n19806 = ~n19638 & ~n19805;
  assign n19807 = pi787 & n19806;
  assign n19808 = ~n19792 & ~n19807;
  assign n19809 = pi644 & n19808;
  assign n19810 = ~n18767 & n19796;
  assign n19811 = ~n19638 & ~n19810;
  assign n19812 = ~pi644 & ~n19811;
  assign n19813 = pi715 & ~n19812;
  assign n19814 = ~n19809 & n19813;
  assign n19815 = ~n17247 & n19793;
  assign n19816 = pi644 & n19815;
  assign n19817 = ~pi715 & ~n19638;
  assign n19818 = ~n19816 & n19817;
  assign n19819 = pi1160 & ~n19818;
  assign n19820 = ~n19814 & n19819;
  assign n19821 = pi644 & ~n19811;
  assign n19822 = ~pi644 & n19808;
  assign n19823 = ~pi715 & ~n19822;
  assign n19824 = ~n19821 & n19823;
  assign n19825 = ~pi1160 & ~n19824;
  assign n19826 = ~pi644 & n19815;
  assign n19827 = ~n19638 & ~n19826;
  assign n19828 = pi715 & n19827;
  assign n19829 = n19825 & ~n19828;
  assign n19830 = ~n19820 & ~n19829;
  assign n19831 = pi790 & ~n19830;
  assign n19832 = ~pi790 & n19808;
  assign n19833 = pi832 & ~n19832;
  assign n19834 = ~n19831 & n19833;
  assign po301 = ~n19636 & ~n19834;
  assign n19836 = ~pi145 & ~n16527;
  assign n19837 = n17159 & ~n19836;
  assign n19838 = n16593 & ~n19836;
  assign n19839 = ~pi698 & n10020;
  assign n19840 = n19836 & ~n19839;
  assign n19841 = ~pi145 & n17592;
  assign n19842 = ~pi38 & ~n17589;
  assign n19843 = n10020 & ~n19842;
  assign n19844 = ~pi38 & ~pi145;
  assign n19845 = n19843 & ~n19844;
  assign n19846 = ~n19841 & ~n19845;
  assign n19847 = ~pi145 & ~n16508;
  assign n19848 = n16744 & ~n19847;
  assign n19849 = ~pi698 & ~n19848;
  assign n19850 = ~n19846 & n19849;
  assign n19851 = ~n19840 & ~n19850;
  assign n19852 = ~pi778 & n19851;
  assign n19853 = pi625 & ~n19851;
  assign n19854 = pi1153 & ~n19853;
  assign n19855 = ~pi625 & n19836;
  assign n19856 = n19854 & ~n19855;
  assign n19857 = ~pi625 & ~n19851;
  assign n19858 = ~pi1153 & ~n19857;
  assign n19859 = pi625 & n19836;
  assign n19860 = n19858 & ~n19859;
  assign n19861 = ~n19856 & ~n19860;
  assign n19862 = pi778 & ~n19861;
  assign n19863 = ~n19852 & ~n19862;
  assign n19864 = ~n16593 & ~n19863;
  assign n19865 = ~n19838 & ~n19864;
  assign n19866 = ~n16589 & n19865;
  assign n19867 = n16589 & n19836;
  assign n19868 = ~n19866 & ~n19867;
  assign n19869 = ~n17159 & n19868;
  assign n19870 = ~n19837 & ~n19869;
  assign n19871 = ~n17183 & n19870;
  assign n19872 = n17183 & n19836;
  assign n19873 = ~n19871 & ~n19872;
  assign n19874 = ~pi792 & n19873;
  assign n19875 = pi628 & ~n19873;
  assign n19876 = pi1156 & ~n19875;
  assign n19877 = ~pi628 & n19836;
  assign n19878 = n19876 & ~n19877;
  assign n19879 = ~pi628 & ~n19873;
  assign n19880 = pi628 & n19836;
  assign n19881 = ~pi1156 & ~n19880;
  assign n19882 = ~n19879 & n19881;
  assign n19883 = ~n19878 & ~n19882;
  assign n19884 = pi792 & ~n19883;
  assign n19885 = ~n19874 & ~n19884;
  assign n19886 = pi647 & ~n19885;
  assign n19887 = ~pi647 & ~n19836;
  assign n19888 = ~n19886 & ~n19887;
  assign n19889 = pi1157 & ~n19888;
  assign n19890 = ~pi647 & n19885;
  assign n19891 = ~pi1157 & ~n19890;
  assign n19892 = pi647 & n19836;
  assign n19893 = n19891 & ~n19892;
  assign n19894 = ~n19889 & ~n19893;
  assign n19895 = pi787 & ~n19894;
  assign n19896 = ~pi787 & ~n19885;
  assign n19897 = ~n19895 & ~n19896;
  assign n19898 = ~pi644 & n19897;
  assign n19899 = pi715 & ~n19898;
  assign n19900 = n17247 & ~n19836;
  assign n19901 = pi145 & ~n10020;
  assign n19902 = ~pi767 & n16511;
  assign n19903 = ~n19847 & ~n19902;
  assign n19904 = pi38 & ~n19903;
  assign n19905 = n10020 & ~n19904;
  assign n19906 = ~pi145 & ~pi767;
  assign n19907 = n16449 & n19906;
  assign n19908 = pi145 & ~n16503;
  assign n19909 = ~pi145 & ~n16357;
  assign n19910 = pi767 & ~n19909;
  assign n19911 = ~n19908 & ~n19910;
  assign n19912 = ~n19907 & n19911;
  assign n19913 = ~pi38 & n19912;
  assign n19914 = n19905 & ~n19913;
  assign n19915 = ~n19901 & ~n19914;
  assign n19916 = ~n16521 & ~n19915;
  assign n19917 = n16521 & ~n19836;
  assign n19918 = ~n19916 & ~n19917;
  assign n19919 = ~pi785 & ~n19918;
  assign n19920 = ~n16532 & ~n19836;
  assign n19921 = pi609 & n19916;
  assign n19922 = ~n19920 & ~n19921;
  assign n19923 = pi1155 & ~n19922;
  assign n19924 = ~n16537 & ~n19836;
  assign n19925 = ~pi609 & n19916;
  assign n19926 = ~n19924 & ~n19925;
  assign n19927 = ~pi1155 & ~n19926;
  assign n19928 = ~n19923 & ~n19927;
  assign n19929 = pi785 & ~n19928;
  assign n19930 = ~n19919 & ~n19929;
  assign n19931 = ~pi781 & ~n19930;
  assign n19932 = pi618 & n19930;
  assign n19933 = ~pi618 & n19836;
  assign n19934 = pi1154 & ~n19933;
  assign n19935 = ~n19932 & n19934;
  assign n19936 = ~pi618 & n19930;
  assign n19937 = pi618 & n19836;
  assign n19938 = ~pi1154 & ~n19937;
  assign n19939 = ~n19936 & n19938;
  assign n19940 = ~n19935 & ~n19939;
  assign n19941 = pi781 & ~n19940;
  assign n19942 = ~n19931 & ~n19941;
  assign n19943 = ~pi789 & ~n19942;
  assign n19944 = pi619 & n19942;
  assign n19945 = ~pi619 & n19836;
  assign n19946 = pi1159 & ~n19945;
  assign n19947 = ~n19944 & n19946;
  assign n19948 = ~pi619 & n19942;
  assign n19949 = pi619 & n19836;
  assign n19950 = ~pi1159 & ~n19949;
  assign n19951 = ~n19948 & n19950;
  assign n19952 = ~n19947 & ~n19951;
  assign n19953 = pi789 & ~n19952;
  assign n19954 = ~n19943 & ~n19953;
  assign n19955 = ~pi788 & ~n19954;
  assign n19956 = pi626 & n19954;
  assign n19957 = ~pi626 & n19836;
  assign n19958 = pi1158 & ~n19957;
  assign n19959 = ~n19956 & n19958;
  assign n19960 = ~pi626 & n19954;
  assign n19961 = pi626 & n19836;
  assign n19962 = ~pi1158 & ~n19961;
  assign n19963 = ~n19960 & n19962;
  assign n19964 = ~n19959 & ~n19963;
  assign n19965 = pi788 & ~n19964;
  assign n19966 = ~n19955 & ~n19965;
  assign n19967 = ~n16124 & n19966;
  assign n19968 = n16124 & n19836;
  assign n19969 = ~n19967 & ~n19968;
  assign n19970 = ~n17247 & n19969;
  assign n19971 = ~n19900 & ~n19970;
  assign n19972 = pi644 & n19971;
  assign n19973 = ~pi644 & n19836;
  assign n19974 = ~pi715 & ~n19973;
  assign n19975 = ~n19972 & n19974;
  assign n19976 = pi1160 & ~n19975;
  assign n19977 = ~n19899 & n19976;
  assign n19978 = ~pi644 & n19971;
  assign n19979 = pi715 & ~n19978;
  assign n19980 = pi644 & n19836;
  assign n19981 = n19979 & ~n19980;
  assign n19982 = pi644 & n19897;
  assign n19983 = pi630 & ~pi647;
  assign n19984 = pi1157 & n19983;
  assign n19985 = ~pi630 & pi647;
  assign n19986 = ~pi1157 & n19985;
  assign n19987 = ~n19984 & ~n19986;
  assign n19988 = n19969 & ~n19987;
  assign n19989 = pi630 & n19893;
  assign n19990 = ~n19988 & ~n19989;
  assign n19991 = n17244 & ~n19888;
  assign n19992 = n19990 & ~n19991;
  assign n19993 = pi787 & ~n19992;
  assign n19994 = ~pi629 & n19878;
  assign n19995 = ~pi628 & pi629;
  assign n19996 = pi1156 & n19995;
  assign n19997 = pi628 & ~pi629;
  assign n19998 = ~pi1156 & n19997;
  assign n19999 = ~n19996 & ~n19998;
  assign n20000 = ~n19966 & ~n19999;
  assign n20001 = pi629 & n19882;
  assign n20002 = ~n20000 & ~n20001;
  assign n20003 = ~n19994 & n20002;
  assign n20004 = pi792 & ~n20003;
  assign n20005 = pi618 & n19865;
  assign n20006 = pi609 & n19863;
  assign n20007 = pi625 & n19915;
  assign n20008 = ~n19839 & ~n19914;
  assign n20009 = ~pi767 & ~n16917;
  assign n20010 = n18933 & ~n20009;
  assign n20011 = ~pi145 & ~n20010;
  assign n20012 = ~pi767 & n16510;
  assign n20013 = ~n17079 & ~n20012;
  assign n20014 = pi145 & ~n20013;
  assign n20015 = n6097 & n20014;
  assign n20016 = ~n20011 & ~n20015;
  assign n20017 = pi38 & n20016;
  assign n20018 = ~pi145 & n16853;
  assign n20019 = pi145 & n16935;
  assign n20020 = pi767 & ~n20019;
  assign n20021 = ~n20018 & n20020;
  assign n20022 = pi145 & n16998;
  assign n20023 = ~pi145 & ~n17051;
  assign n20024 = ~pi767 & ~n20023;
  assign n20025 = ~n20022 & n20024;
  assign n20026 = ~n20021 & ~n20025;
  assign n20027 = pi39 & n20026;
  assign n20028 = ~pi145 & ~n17061;
  assign n20029 = pi145 & ~n17058;
  assign n20030 = pi767 & ~n20029;
  assign n20031 = ~n20028 & n20030;
  assign n20032 = ~pi145 & n17067;
  assign n20033 = pi145 & n17065;
  assign n20034 = ~pi767 & ~n20033;
  assign n20035 = ~n20032 & n20034;
  assign n20036 = ~n20031 & ~n20035;
  assign n20037 = ~pi39 & ~n20036;
  assign n20038 = ~pi38 & ~n20037;
  assign n20039 = ~n20027 & n20038;
  assign n20040 = ~pi698 & ~n20039;
  assign n20041 = ~n20017 & n20040;
  assign n20042 = ~n20008 & ~n20041;
  assign n20043 = ~n19901 & ~n20042;
  assign n20044 = ~pi625 & n20043;
  assign n20045 = ~pi1153 & ~n20044;
  assign n20046 = ~n20007 & n20045;
  assign n20047 = ~pi608 & ~n19856;
  assign n20048 = ~n20046 & n20047;
  assign n20049 = ~pi625 & n19915;
  assign n20050 = pi625 & n20043;
  assign n20051 = ~n20049 & ~n20050;
  assign n20052 = pi1153 & n20051;
  assign n20053 = ~n19860 & ~n20052;
  assign n20054 = pi608 & n20053;
  assign n20055 = ~n20048 & ~n20054;
  assign n20056 = pi778 & ~n20055;
  assign n20057 = ~pi778 & n20043;
  assign n20058 = ~n20056 & ~n20057;
  assign n20059 = ~pi609 & ~n20058;
  assign n20060 = ~pi1155 & ~n20059;
  assign n20061 = ~n20006 & n20060;
  assign n20062 = ~pi660 & ~n19923;
  assign n20063 = ~n20061 & n20062;
  assign n20064 = ~pi609 & n19863;
  assign n20065 = pi609 & ~n20058;
  assign n20066 = ~n20064 & ~n20065;
  assign n20067 = pi1155 & n20066;
  assign n20068 = ~n19927 & ~n20067;
  assign n20069 = pi660 & n20068;
  assign n20070 = ~n20063 & ~n20069;
  assign n20071 = pi785 & ~n20070;
  assign n20072 = ~pi785 & ~n20058;
  assign n20073 = ~n20071 & ~n20072;
  assign n20074 = ~pi618 & ~n20073;
  assign n20075 = ~pi1154 & ~n20074;
  assign n20076 = ~n20005 & n20075;
  assign n20077 = ~pi627 & ~n19935;
  assign n20078 = ~n20076 & n20077;
  assign n20079 = ~pi618 & n19865;
  assign n20080 = pi618 & ~n20073;
  assign n20081 = ~n20079 & ~n20080;
  assign n20082 = pi1154 & n20081;
  assign n20083 = ~n19939 & ~n20082;
  assign n20084 = pi627 & n20083;
  assign n20085 = ~n20078 & ~n20084;
  assign n20086 = pi781 & ~n20085;
  assign n20087 = ~pi781 & ~n20073;
  assign n20088 = ~n20086 & ~n20087;
  assign n20089 = ~pi789 & n20088;
  assign n20090 = ~pi619 & ~n20088;
  assign n20091 = pi619 & ~n19868;
  assign n20092 = ~pi1159 & ~n20091;
  assign n20093 = ~n20090 & n20092;
  assign n20094 = ~pi648 & ~n20093;
  assign n20095 = ~n19947 & n20094;
  assign n20096 = ~pi619 & ~n19868;
  assign n20097 = pi619 & ~n20088;
  assign n20098 = ~n20096 & ~n20097;
  assign n20099 = pi1159 & n20098;
  assign n20100 = ~n19951 & ~n20099;
  assign n20101 = pi648 & n20100;
  assign n20102 = ~n20095 & ~n20101;
  assign n20103 = pi789 & n20102;
  assign n20104 = ~n20089 & ~n20103;
  assign n20105 = n17356 & n20104;
  assign n20106 = n17350 & n19870;
  assign n20107 = ~n17182 & n19964;
  assign n20108 = ~n20106 & ~n20107;
  assign n20109 = pi788 & ~n20108;
  assign n20110 = n19788 & ~n20109;
  assign n20111 = ~n20105 & n20110;
  assign n20112 = ~n20004 & ~n20111;
  assign n20113 = n19637 & ~n20112;
  assign n20114 = ~n19993 & ~n20113;
  assign n20115 = ~pi644 & n20114;
  assign n20116 = ~pi715 & ~n20115;
  assign n20117 = ~n19982 & n20116;
  assign n20118 = ~pi1160 & ~n20117;
  assign n20119 = ~n19981 & n20118;
  assign n20120 = ~n19977 & ~n20119;
  assign n20121 = pi790 & ~n20120;
  assign n20122 = pi644 & n19976;
  assign n20123 = pi790 & ~n20122;
  assign n20124 = n20114 & ~n20123;
  assign n20125 = ~n20121 & ~n20124;
  assign n20126 = ~po1038 & ~n20125;
  assign n20127 = ~pi145 & po1038;
  assign n20128 = ~pi832 & ~n20127;
  assign n20129 = ~n20126 & n20128;
  assign n20130 = ~pi145 & ~n2934;
  assign n20131 = ~n20012 & ~n20130;
  assign n20132 = ~n17273 & ~n20131;
  assign n20133 = ~pi785 & ~n20132;
  assign n20134 = ~n17279 & ~n20131;
  assign n20135 = pi1155 & ~n20134;
  assign n20136 = ~n17282 & n20132;
  assign n20137 = ~pi1155 & ~n20136;
  assign n20138 = ~n20135 & ~n20137;
  assign n20139 = pi785 & ~n20138;
  assign n20140 = ~n20133 & ~n20139;
  assign n20141 = ~pi781 & ~n20140;
  assign n20142 = ~n17289 & n20140;
  assign n20143 = pi1154 & ~n20142;
  assign n20144 = ~n17292 & n20140;
  assign n20145 = ~pi1154 & ~n20144;
  assign n20146 = ~n20143 & ~n20145;
  assign n20147 = pi781 & ~n20146;
  assign n20148 = ~n20141 & ~n20147;
  assign n20149 = ~pi789 & ~n20148;
  assign n20150 = pi619 & n20148;
  assign n20151 = ~pi619 & n20130;
  assign n20152 = pi1159 & ~n20151;
  assign n20153 = ~n20150 & n20152;
  assign n20154 = ~pi619 & n20148;
  assign n20155 = pi619 & n20130;
  assign n20156 = ~pi1159 & ~n20155;
  assign n20157 = ~n20154 & n20156;
  assign n20158 = ~n20153 & ~n20157;
  assign n20159 = pi789 & ~n20158;
  assign n20160 = ~n20149 & ~n20159;
  assign n20161 = ~pi788 & ~n20160;
  assign n20162 = pi626 & n20160;
  assign n20163 = ~pi626 & n20130;
  assign n20164 = pi1158 & ~n20163;
  assign n20165 = ~n20162 & n20164;
  assign n20166 = ~pi626 & n20160;
  assign n20167 = pi626 & n20130;
  assign n20168 = ~pi1158 & ~n20167;
  assign n20169 = ~n20166 & n20168;
  assign n20170 = ~n20165 & ~n20169;
  assign n20171 = pi788 & ~n20170;
  assign n20172 = ~n20161 & ~n20171;
  assign n20173 = ~n16124 & n20172;
  assign n20174 = n16124 & n20130;
  assign n20175 = ~n20173 & ~n20174;
  assign n20176 = ~n19987 & n20175;
  assign n20177 = ~pi698 & n16742;
  assign n20178 = ~n20130 & ~n20177;
  assign n20179 = ~pi778 & n20178;
  assign n20180 = ~pi625 & n20177;
  assign n20181 = ~n20178 & ~n20180;
  assign n20182 = pi1153 & ~n20181;
  assign n20183 = ~pi1153 & ~n20130;
  assign n20184 = ~n20180 & n20183;
  assign n20185 = ~n20182 & ~n20184;
  assign n20186 = pi778 & ~n20185;
  assign n20187 = ~n20179 & ~n20186;
  assign n20188 = ~n17338 & n20187;
  assign n20189 = ~n17340 & n20188;
  assign n20190 = ~n17342 & n20189;
  assign n20191 = ~n17425 & n20190;
  assign n20192 = ~n17452 & n20191;
  assign n20193 = ~pi647 & n20192;
  assign n20194 = pi647 & n20130;
  assign n20195 = ~pi1157 & ~n20194;
  assign n20196 = ~n20193 & n20195;
  assign n20197 = ~pi647 & n20130;
  assign n20198 = pi647 & n20192;
  assign n20199 = pi1157 & ~n20198;
  assign n20200 = ~n20197 & n20199;
  assign n20201 = ~n20196 & ~n20200;
  assign n20202 = ~n17246 & ~n20201;
  assign n20203 = ~n20176 & ~n20202;
  assign n20204 = pi787 & ~n20203;
  assign n20205 = n17350 & n20190;
  assign n20206 = ~n17182 & n20170;
  assign n20207 = ~n20205 & ~n20206;
  assign n20208 = pi788 & ~n20207;
  assign n20209 = pi618 & n20188;
  assign n20210 = pi609 & n20187;
  assign n20211 = ~n16393 & ~n20178;
  assign n20212 = pi625 & n20211;
  assign n20213 = n20131 & ~n20211;
  assign n20214 = ~n20212 & ~n20213;
  assign n20215 = n20183 & ~n20214;
  assign n20216 = ~pi608 & ~n20182;
  assign n20217 = ~n20215 & n20216;
  assign n20218 = pi1153 & ~n20212;
  assign n20219 = n20131 & n20218;
  assign n20220 = ~n20184 & ~n20219;
  assign n20221 = pi608 & n20220;
  assign n20222 = ~n20217 & ~n20221;
  assign n20223 = pi778 & ~n20222;
  assign n20224 = ~pi778 & ~n20213;
  assign n20225 = ~n20223 & ~n20224;
  assign n20226 = ~pi609 & ~n20225;
  assign n20227 = ~pi1155 & ~n20226;
  assign n20228 = ~n20210 & n20227;
  assign n20229 = ~pi660 & ~n20135;
  assign n20230 = ~n20228 & n20229;
  assign n20231 = ~pi609 & n20187;
  assign n20232 = pi609 & ~n20225;
  assign n20233 = ~n20231 & ~n20232;
  assign n20234 = pi1155 & n20233;
  assign n20235 = ~n20137 & ~n20234;
  assign n20236 = pi660 & n20235;
  assign n20237 = ~n20230 & ~n20236;
  assign n20238 = pi785 & ~n20237;
  assign n20239 = ~pi785 & ~n20225;
  assign n20240 = ~n20238 & ~n20239;
  assign n20241 = ~pi618 & ~n20240;
  assign n20242 = ~pi1154 & ~n20241;
  assign n20243 = ~n20209 & n20242;
  assign n20244 = ~pi627 & ~n20143;
  assign n20245 = ~n20243 & n20244;
  assign n20246 = ~pi618 & n20188;
  assign n20247 = pi618 & ~n20240;
  assign n20248 = ~n20246 & ~n20247;
  assign n20249 = pi1154 & n20248;
  assign n20250 = ~n20145 & ~n20249;
  assign n20251 = pi627 & n20250;
  assign n20252 = ~n20245 & ~n20251;
  assign n20253 = pi781 & ~n20252;
  assign n20254 = ~pi781 & ~n20240;
  assign n20255 = ~n20253 & ~n20254;
  assign n20256 = ~pi619 & ~n20255;
  assign n20257 = pi619 & n20189;
  assign n20258 = ~pi1159 & ~n20257;
  assign n20259 = ~n20256 & n20258;
  assign n20260 = ~pi648 & ~n20259;
  assign n20261 = ~n20153 & n20260;
  assign n20262 = ~pi619 & n20189;
  assign n20263 = pi619 & ~n20255;
  assign n20264 = ~n20262 & ~n20263;
  assign n20265 = pi1159 & n20264;
  assign n20266 = ~n20157 & ~n20265;
  assign n20267 = pi648 & n20266;
  assign n20268 = ~n20261 & ~n20267;
  assign n20269 = pi789 & n20268;
  assign n20270 = ~pi789 & n20255;
  assign n20271 = n17356 & ~n20270;
  assign n20272 = ~n20269 & n20271;
  assign n20273 = ~n20208 & ~n20272;
  assign n20274 = n19788 & ~n20273;
  assign n20275 = pi1156 & ~n17427;
  assign n20276 = n20191 & n20275;
  assign n20277 = n17449 & n20172;
  assign n20278 = ~pi629 & ~n20277;
  assign n20279 = ~n20276 & n20278;
  assign n20280 = n17448 & n20172;
  assign n20281 = ~pi1156 & ~n17436;
  assign n20282 = n20191 & n20281;
  assign n20283 = pi629 & ~n20282;
  assign n20284 = ~n20280 & n20283;
  assign n20285 = ~n20279 & ~n20284;
  assign n20286 = pi792 & n20285;
  assign n20287 = n19637 & ~n20286;
  assign n20288 = ~n20274 & n20287;
  assign n20289 = ~n20204 & ~n20288;
  assign n20290 = pi644 & n20289;
  assign n20291 = ~pi787 & ~n20192;
  assign n20292 = pi787 & ~n20201;
  assign n20293 = ~n20291 & ~n20292;
  assign n20294 = ~pi644 & n20293;
  assign n20295 = pi715 & ~n20294;
  assign n20296 = ~n20290 & n20295;
  assign n20297 = ~n17247 & ~n20175;
  assign n20298 = n17247 & n20130;
  assign n20299 = ~n20297 & ~n20298;
  assign n20300 = pi644 & ~n20299;
  assign n20301 = ~pi644 & n20130;
  assign n20302 = ~pi715 & ~n20301;
  assign n20303 = ~n20300 & n20302;
  assign n20304 = pi1160 & ~n20303;
  assign n20305 = ~n20296 & n20304;
  assign n20306 = ~pi644 & ~n20299;
  assign n20307 = pi715 & ~n20306;
  assign n20308 = pi644 & n20130;
  assign n20309 = n20307 & ~n20308;
  assign n20310 = pi644 & n20293;
  assign n20311 = ~pi644 & n20289;
  assign n20312 = ~pi715 & ~n20311;
  assign n20313 = ~n20310 & n20312;
  assign n20314 = ~pi1160 & ~n20313;
  assign n20315 = ~n20309 & n20314;
  assign n20316 = ~n20305 & ~n20315;
  assign n20317 = pi790 & ~n20316;
  assign n20318 = ~pi790 & n20289;
  assign n20319 = pi832 & ~n20318;
  assign n20320 = ~n20317 & n20319;
  assign po302 = ~n20129 & ~n20320;
  assign n20322 = pi743 & pi947;
  assign n20323 = pi907 & ~pi947;
  assign n20324 = pi735 & n20323;
  assign n20325 = ~n20322 & ~n20324;
  assign n20326 = n16508 & n20325;
  assign n20327 = ~pi146 & ~n16508;
  assign n20328 = pi38 & ~n20327;
  assign n20329 = ~n20326 & n20328;
  assign n20330 = ~pi146 & ~n16195;
  assign n20331 = n16195 & n20325;
  assign n20332 = ~n20330 & ~n20331;
  assign n20333 = pi299 & n20332;
  assign n20334 = n16199 & n20325;
  assign n20335 = ~pi146 & ~n16199;
  assign n20336 = ~pi299 & ~n20335;
  assign n20337 = ~n20334 & n20336;
  assign n20338 = ~pi39 & ~n20337;
  assign n20339 = ~n20333 & n20338;
  assign n20340 = ~pi907 & n6197;
  assign n20341 = pi146 & ~n16297;
  assign n20342 = ~n20340 & n20341;
  assign n20343 = pi146 & ~n16327;
  assign n20344 = n20340 & n20343;
  assign n20345 = ~pi947 & ~n20344;
  assign n20346 = pi735 & pi907;
  assign n20347 = n16297 & n20346;
  assign n20348 = n20345 & ~n20347;
  assign n20349 = pi743 & n16297;
  assign n20350 = ~n20341 & ~n20349;
  assign n20351 = pi947 & n20350;
  assign n20352 = ~n20348 & ~n20351;
  assign n20353 = ~n20342 & ~n20352;
  assign n20354 = ~n2527 & ~n20353;
  assign n20355 = n16207 & ~n20325;
  assign n20356 = pi146 & ~n16207;
  assign n20357 = ~n20355 & ~n20356;
  assign n20358 = n2527 & ~n20357;
  assign n20359 = ~pi215 & ~n20358;
  assign n20360 = ~n20354 & n20359;
  assign n20361 = pi146 & n16351;
  assign n20362 = n16267 & ~n20325;
  assign n20363 = ~n20361 & ~n20362;
  assign n20364 = pi215 & n20363;
  assign n20365 = ~n20360 & ~n20364;
  assign n20366 = pi299 & ~n20365;
  assign n20367 = n2607 & n20357;
  assign n20368 = n16297 & ~n20325;
  assign n20369 = ~n6236 & ~n20341;
  assign n20370 = ~n20368 & n20369;
  assign n20371 = n16327 & ~n20325;
  assign n20372 = ~n20343 & ~n20371;
  assign n20373 = n6236 & n20372;
  assign n20374 = ~n20370 & ~n20373;
  assign n20375 = ~n2607 & ~n20374;
  assign n20376 = ~pi223 & ~n20375;
  assign n20377 = ~n20367 & n20376;
  assign n20378 = pi146 & ~n16267;
  assign n20379 = ~n20362 & ~n20378;
  assign n20380 = ~n6236 & ~n20379;
  assign n20381 = n16250 & n20325;
  assign n20382 = ~pi146 & ~n16250;
  assign n20383 = n6236 & ~n20382;
  assign n20384 = ~n20381 & n20383;
  assign n20385 = ~n20380 & ~n20384;
  assign n20386 = pi223 & ~n20385;
  assign n20387 = ~pi299 & ~n20386;
  assign n20388 = ~n20377 & n20387;
  assign n20389 = ~n20366 & ~n20388;
  assign n20390 = pi39 & ~n20389;
  assign n20391 = ~pi38 & ~n20390;
  assign n20392 = ~n20339 & n20391;
  assign n20393 = n10021 & ~n20392;
  assign n20394 = ~n20329 & n20393;
  assign n20395 = ~pi146 & ~n10021;
  assign n20396 = ~pi832 & ~n20395;
  assign n20397 = ~n20394 & n20396;
  assign n20398 = n2934 & n20325;
  assign n20399 = ~pi146 & ~n2934;
  assign n20400 = pi832 & ~n20399;
  assign n20401 = ~n20398 & n20400;
  assign po303 = n20397 | n20401;
  assign n20403 = ~pi770 & pi947;
  assign n20404 = pi726 & n20323;
  assign n20405 = ~n20403 & ~n20404;
  assign n20406 = n2934 & ~n20405;
  assign n20407 = ~pi147 & ~n2934;
  assign n20408 = pi832 & ~n20407;
  assign n20409 = ~n20406 & n20408;
  assign n20410 = n16267 & n20323;
  assign n20411 = pi215 & ~n20410;
  assign n20412 = n16297 & n20323;
  assign n20413 = ~n2527 & ~n20412;
  assign n20414 = pi907 & n16207;
  assign n20415 = ~pi947 & n20414;
  assign n20416 = n2527 & ~n20415;
  assign n20417 = ~n20413 & ~n20416;
  assign n20418 = ~pi215 & ~n20417;
  assign n20419 = ~n20411 & ~n20418;
  assign n20420 = pi299 & ~n20419;
  assign n20421 = n16333 & n20323;
  assign n20422 = ~pi299 & ~n20421;
  assign n20423 = ~n20420 & ~n20422;
  assign n20424 = pi39 & ~n20423;
  assign n20425 = n16201 & n20323;
  assign n20426 = ~pi39 & ~n20425;
  assign n20427 = ~n20424 & ~n20426;
  assign n20428 = pi147 & n20427;
  assign n20429 = pi215 & ~n16350;
  assign n20430 = n16342 & ~n20323;
  assign n20431 = pi947 & n16297;
  assign n20432 = ~n16338 & ~n20431;
  assign n20433 = ~n2527 & ~n20432;
  assign n20434 = ~pi215 & ~n20433;
  assign n20435 = ~n20430 & n20434;
  assign n20436 = ~n20429 & ~n20435;
  assign n20437 = pi215 & pi947;
  assign n20438 = n16267 & n20437;
  assign n20439 = ~n20436 & ~n20438;
  assign n20440 = pi299 & ~n20439;
  assign n20441 = ~pi299 & n16333;
  assign n20442 = ~n20323 & n20441;
  assign n20443 = ~n20440 & ~n20442;
  assign n20444 = pi39 & ~n20443;
  assign n20445 = n16201 & ~n20323;
  assign n20446 = ~pi39 & n20445;
  assign n20447 = ~n20444 & ~n20446;
  assign n20448 = ~pi147 & n20447;
  assign n20449 = ~pi38 & ~n20448;
  assign n20450 = ~n20428 & n20449;
  assign n20451 = ~pi147 & ~n16508;
  assign n20452 = n16508 & n20323;
  assign n20453 = pi38 & ~n20452;
  assign n20454 = ~n20451 & n20453;
  assign n20455 = pi770 & ~n20454;
  assign n20456 = ~n20450 & n20455;
  assign n20457 = n6192 & n16524;
  assign n20458 = ~pi147 & ~n20457;
  assign n20459 = ~n6192 & n16508;
  assign n20460 = pi38 & ~n20459;
  assign n20461 = ~n20458 & n20460;
  assign n20462 = pi299 & pi947;
  assign n20463 = pi299 & ~n20436;
  assign n20464 = ~n20462 & ~n20463;
  assign n20465 = ~n6192 & n20441;
  assign n20466 = ~n16334 & ~n20465;
  assign n20467 = n20464 & n20466;
  assign n20468 = pi39 & n20467;
  assign n20469 = ~n6192 & n16201;
  assign n20470 = ~pi39 & ~n20469;
  assign n20471 = n16201 & n20470;
  assign n20472 = ~n20468 & ~n20471;
  assign n20473 = ~pi147 & n20472;
  assign n20474 = pi215 & ~n16346;
  assign n20475 = ~n6192 & ~n16344;
  assign n20476 = ~n20474 & n20475;
  assign n20477 = pi299 & n20476;
  assign n20478 = ~n20465 & ~n20477;
  assign n20479 = pi39 & n20478;
  assign n20480 = ~n20470 & ~n20479;
  assign n20481 = pi147 & n20480;
  assign n20482 = ~pi38 & ~n20481;
  assign n20483 = ~n20473 & n20482;
  assign n20484 = ~pi770 & ~n20483;
  assign n20485 = ~n20461 & n20484;
  assign n20486 = ~n20456 & ~n20485;
  assign n20487 = pi726 & n20486;
  assign n20488 = ~pi947 & n18801;
  assign n20489 = ~pi947 & n16201;
  assign n20490 = ~pi39 & ~n20489;
  assign n20491 = ~pi947 & n16342;
  assign n20492 = ~n16338 & ~n20412;
  assign n20493 = ~n2527 & ~n20492;
  assign n20494 = ~pi215 & ~n20493;
  assign n20495 = ~n20491 & n20494;
  assign n20496 = ~n20410 & n20429;
  assign n20497 = ~n20495 & ~n20496;
  assign n20498 = pi299 & ~n20497;
  assign n20499 = ~n16334 & ~n20498;
  assign n20500 = pi947 & n20441;
  assign n20501 = n20499 & ~n20500;
  assign n20502 = pi39 & ~n20501;
  assign n20503 = ~n20490 & ~n20502;
  assign n20504 = ~pi38 & n20503;
  assign n20505 = ~n20488 & ~n20504;
  assign n20506 = ~pi770 & n20505;
  assign n20507 = pi770 & ~n16526;
  assign n20508 = ~n20506 & ~n20507;
  assign n20509 = ~pi147 & ~n20508;
  assign n20510 = ~n16525 & ~n20488;
  assign n20511 = pi947 & n16201;
  assign n20512 = ~pi39 & ~n20511;
  assign n20513 = pi947 & n16333;
  assign n20514 = ~pi299 & ~n20513;
  assign n20515 = pi299 & ~n20438;
  assign n20516 = ~n2527 & ~n20431;
  assign n20517 = pi947 & n16207;
  assign n20518 = n2527 & ~n20517;
  assign n20519 = ~pi215 & ~n20518;
  assign n20520 = ~n20516 & n20519;
  assign n20521 = n20515 & ~n20520;
  assign n20522 = ~n20514 & ~n20521;
  assign n20523 = pi39 & ~n20522;
  assign n20524 = ~n20512 & ~n20523;
  assign n20525 = ~pi38 & ~n20524;
  assign n20526 = n20510 & ~n20525;
  assign n20527 = pi147 & ~pi770;
  assign n20528 = n20526 & n20527;
  assign n20529 = ~pi726 & ~n20528;
  assign n20530 = ~n20509 & n20529;
  assign n20531 = n10021 & ~n20530;
  assign n20532 = ~n20487 & n20531;
  assign n20533 = ~pi147 & ~n10021;
  assign n20534 = ~pi832 & ~n20533;
  assign n20535 = ~n20532 & n20534;
  assign po304 = ~n20409 & ~n20535;
  assign n20537 = n6274 & n10020;
  assign n20538 = ~pi148 & ~n20537;
  assign n20539 = ~pi148 & ~n16201;
  assign n20540 = ~pi39 & ~n20539;
  assign n20541 = ~pi749 & pi947;
  assign n20542 = n20469 & ~n20541;
  assign n20543 = n20540 & ~n20542;
  assign n20544 = ~pi148 & n20467;
  assign n20545 = pi148 & n20478;
  assign n20546 = pi749 & ~n20545;
  assign n20547 = ~n20544 & n20546;
  assign n20548 = ~n9582 & ~n20443;
  assign n20549 = ~n16334 & ~n20420;
  assign n20550 = pi148 & ~n20549;
  assign n20551 = ~pi749 & ~n20550;
  assign n20552 = ~n20548 & n20551;
  assign n20553 = ~n20547 & ~n20552;
  assign n20554 = pi39 & n20553;
  assign n20555 = ~pi38 & ~n20554;
  assign n20556 = ~n20543 & n20555;
  assign n20557 = n20459 & ~n20541;
  assign n20558 = ~pi148 & ~n16508;
  assign n20559 = ~n20557 & ~n20558;
  assign n20560 = pi38 & ~n20559;
  assign n20561 = pi706 & ~n20560;
  assign n20562 = ~n20556 & n20561;
  assign n20563 = pi148 & ~n16524;
  assign n20564 = pi749 & pi947;
  assign n20565 = n2934 & ~n20564;
  assign n20566 = n6097 & n20565;
  assign n20567 = ~n20563 & ~n20566;
  assign n20568 = pi38 & n20567;
  assign n20569 = ~pi148 & ~pi749;
  assign n20570 = ~n16355 & n20569;
  assign n20571 = ~pi148 & ~n16333;
  assign n20572 = n20514 & ~n20571;
  assign n20573 = ~n20438 & ~n20520;
  assign n20574 = pi148 & ~n20573;
  assign n20575 = ~pi148 & ~n20497;
  assign n20576 = ~n20574 & ~n20575;
  assign n20577 = pi299 & n20576;
  assign n20578 = ~n20572 & ~n20577;
  assign n20579 = pi749 & n20578;
  assign n20580 = ~n20570 & ~n20579;
  assign n20581 = pi39 & n20580;
  assign n20582 = n16201 & n20564;
  assign n20583 = n20540 & ~n20582;
  assign n20584 = ~pi38 & ~n20583;
  assign n20585 = ~n20581 & n20584;
  assign n20586 = ~pi706 & ~n20585;
  assign n20587 = ~n20568 & n20586;
  assign n20588 = ~n20562 & ~n20587;
  assign n20589 = n20537 & n20588;
  assign n20590 = ~pi57 & ~n20589;
  assign n20591 = ~n20538 & n20590;
  assign n20592 = pi57 & pi148;
  assign n20593 = ~pi832 & ~n20592;
  assign n20594 = ~n20591 & n20593;
  assign n20595 = pi706 & n20323;
  assign n20596 = n20565 & ~n20595;
  assign n20597 = pi148 & ~n2934;
  assign n20598 = pi832 & ~n20597;
  assign n20599 = ~n20596 & n20598;
  assign po305 = n20594 | n20599;
  assign n20601 = ~pi755 & pi947;
  assign n20602 = ~pi725 & n20323;
  assign n20603 = ~n20601 & ~n20602;
  assign n20604 = n2934 & ~n20603;
  assign n20605 = ~pi149 & ~n2934;
  assign n20606 = pi832 & ~n20605;
  assign n20607 = ~n20604 & n20606;
  assign n20608 = pi149 & ~n16524;
  assign n20609 = n16508 & ~n20601;
  assign n20610 = pi38 & ~n20609;
  assign n20611 = ~n20608 & n20610;
  assign n20612 = ~pi149 & ~n16333;
  assign n20613 = n20514 & ~n20612;
  assign n20614 = ~pi149 & ~n20497;
  assign n20615 = ~n15612 & ~n20521;
  assign n20616 = ~n20614 & ~n20615;
  assign n20617 = ~pi755 & ~n20616;
  assign n20618 = ~n20613 & n20617;
  assign n20619 = ~pi149 & pi755;
  assign n20620 = ~n16355 & n20619;
  assign n20621 = pi39 & ~n20620;
  assign n20622 = ~n20618 & n20621;
  assign n20623 = ~pi149 & ~n16201;
  assign n20624 = ~pi39 & ~n20623;
  assign n20625 = n16201 & n20601;
  assign n20626 = n20624 & ~n20625;
  assign n20627 = ~pi38 & ~n20626;
  assign n20628 = ~n20622 & n20627;
  assign n20629 = ~n20611 & ~n20628;
  assign n20630 = pi725 & ~n20629;
  assign n20631 = ~n20425 & n20626;
  assign n20632 = ~pi149 & n20467;
  assign n20633 = pi149 & n20478;
  assign n20634 = ~pi755 & ~n20633;
  assign n20635 = ~n20632 & n20634;
  assign n20636 = pi149 & ~n20549;
  assign n20637 = n15612 & ~n20439;
  assign n20638 = pi755 & ~n20637;
  assign n20639 = ~n20442 & n20638;
  assign n20640 = ~n20636 & n20639;
  assign n20641 = pi39 & ~n20640;
  assign n20642 = ~n20635 & n20641;
  assign n20643 = ~n20631 & ~n20642;
  assign n20644 = ~pi38 & ~n20643;
  assign n20645 = pi149 & ~n16508;
  assign n20646 = ~n20609 & ~n20645;
  assign n20647 = n20453 & ~n20646;
  assign n20648 = ~pi725 & ~n20647;
  assign n20649 = ~n20644 & n20648;
  assign n20650 = ~n20630 & ~n20649;
  assign n20651 = n10021 & ~n20650;
  assign n20652 = ~pi149 & ~n10021;
  assign n20653 = ~pi832 & ~n20652;
  assign n20654 = ~n20651 & n20653;
  assign po306 = ~n20607 & ~n20654;
  assign n20656 = ~pi150 & n20501;
  assign n20657 = pi150 & ~n20522;
  assign n20658 = ~pi751 & ~n20657;
  assign n20659 = ~n20656 & n20658;
  assign n20660 = ~pi150 & ~n16355;
  assign n20661 = pi751 & n20660;
  assign n20662 = ~n20659 & ~n20661;
  assign n20663 = pi39 & ~n20662;
  assign n20664 = pi150 & ~n16201;
  assign n20665 = pi751 & n16201;
  assign n20666 = ~n20664 & ~n20665;
  assign n20667 = n20490 & n20666;
  assign n20668 = ~pi38 & ~n20667;
  assign n20669 = ~n20663 & n20668;
  assign n20670 = pi150 & ~n16524;
  assign n20671 = ~pi751 & pi947;
  assign n20672 = n16508 & ~n20671;
  assign n20673 = ~n20670 & ~n20672;
  assign n20674 = pi38 & ~n20673;
  assign n20675 = pi701 & ~n20674;
  assign n20676 = ~n20669 & n20675;
  assign n20677 = ~pi150 & ~n20443;
  assign n20678 = pi150 & ~n20423;
  assign n20679 = pi751 & ~n20678;
  assign n20680 = ~n20677 & n20679;
  assign n20681 = ~pi150 & n20467;
  assign n20682 = pi150 & n20478;
  assign n20683 = ~pi751 & ~n20682;
  assign n20684 = ~n20681 & n20683;
  assign n20685 = ~n20680 & ~n20684;
  assign n20686 = pi39 & ~n20685;
  assign n20687 = n20445 & ~n20671;
  assign n20688 = ~pi39 & ~n20687;
  assign n20689 = ~n20664 & n20688;
  assign n20690 = ~pi38 & ~n20689;
  assign n20691 = ~n20686 & n20690;
  assign n20692 = pi150 & ~n16508;
  assign n20693 = ~n20672 & ~n20692;
  assign n20694 = n20453 & ~n20693;
  assign n20695 = ~pi701 & ~n20694;
  assign n20696 = ~n20691 & n20695;
  assign n20697 = ~n20676 & ~n20696;
  assign n20698 = n10021 & ~n20697;
  assign n20699 = ~pi150 & ~n10021;
  assign n20700 = ~pi832 & ~n20699;
  assign n20701 = ~n20698 & n20700;
  assign n20702 = ~pi701 & n20323;
  assign n20703 = ~n20671 & ~n20702;
  assign n20704 = n2934 & ~n20703;
  assign n20705 = ~pi150 & ~n2934;
  assign n20706 = pi832 & ~n20705;
  assign n20707 = ~n20704 & n20706;
  assign po307 = ~n20701 & ~n20707;
  assign n20709 = ~pi745 & pi947;
  assign n20710 = ~pi723 & n20323;
  assign n20711 = ~n20709 & ~n20710;
  assign n20712 = n2934 & ~n20711;
  assign n20713 = ~pi151 & ~n2934;
  assign n20714 = pi832 & ~n20713;
  assign n20715 = ~n20712 & n20714;
  assign n20716 = ~pi151 & ~n16201;
  assign n20717 = ~pi745 & n20511;
  assign n20718 = ~n20716 & ~n20717;
  assign n20719 = n20426 & n20718;
  assign n20720 = ~n16350 & ~n20410;
  assign n20721 = ~pi151 & n20720;
  assign n20722 = ~n16346 & ~n20721;
  assign n20723 = pi215 & ~n20722;
  assign n20724 = ~n2527 & ~n16340;
  assign n20725 = pi151 & n20724;
  assign n20726 = ~n16339 & ~n20725;
  assign n20727 = ~pi151 & ~n16207;
  assign n20728 = n20416 & ~n20727;
  assign n20729 = ~n6192 & n16207;
  assign n20730 = n20728 & ~n20729;
  assign n20731 = ~pi215 & ~n20730;
  assign n20732 = n20726 & n20731;
  assign n20733 = ~n20723 & ~n20732;
  assign n20734 = pi299 & ~n20733;
  assign n20735 = ~n6192 & n16333;
  assign n20736 = pi151 & ~n20735;
  assign n20737 = ~n20466 & ~n20736;
  assign n20738 = ~n20734 & ~n20737;
  assign n20739 = ~pi745 & ~n20738;
  assign n20740 = ~pi151 & ~n16333;
  assign n20741 = n20422 & ~n20740;
  assign n20742 = n20726 & ~n20728;
  assign n20743 = n20434 & n20742;
  assign n20744 = ~n20723 & ~n20743;
  assign n20745 = ~n20438 & ~n20744;
  assign n20746 = pi299 & ~n20745;
  assign n20747 = pi745 & ~n20746;
  assign n20748 = ~n20741 & n20747;
  assign n20749 = pi39 & ~n20748;
  assign n20750 = ~n20739 & n20749;
  assign n20751 = ~n20719 & ~n20750;
  assign n20752 = ~pi38 & ~n20751;
  assign n20753 = n16508 & ~n20709;
  assign n20754 = pi151 & ~n16508;
  assign n20755 = ~n20753 & ~n20754;
  assign n20756 = n20453 & ~n20755;
  assign n20757 = ~pi723 & ~n20756;
  assign n20758 = ~n20752 & n20757;
  assign n20759 = ~pi39 & ~n20718;
  assign n20760 = ~pi745 & ~n16334;
  assign n20761 = ~pi151 & ~n16355;
  assign n20762 = ~n20760 & n20761;
  assign n20763 = n20518 & ~n20727;
  assign n20764 = n20494 & ~n20763;
  assign n20765 = n20726 & n20764;
  assign n20766 = ~n20410 & n20723;
  assign n20767 = pi299 & ~n20766;
  assign n20768 = ~n20765 & n20767;
  assign n20769 = ~pi745 & ~n20514;
  assign n20770 = ~n20768 & n20769;
  assign n20771 = ~n20762 & ~n20770;
  assign n20772 = pi39 & ~n20771;
  assign n20773 = ~pi38 & ~n20772;
  assign n20774 = ~n20759 & n20773;
  assign n20775 = pi151 & ~n16524;
  assign n20776 = ~n20753 & ~n20775;
  assign n20777 = pi38 & ~n20776;
  assign n20778 = pi723 & ~n20777;
  assign n20779 = ~n20774 & n20778;
  assign n20780 = ~n20758 & ~n20779;
  assign n20781 = n10021 & ~n20780;
  assign n20782 = ~pi151 & ~n10021;
  assign n20783 = ~pi832 & ~n20782;
  assign n20784 = ~n20781 & n20783;
  assign po308 = ~n20715 & ~n20784;
  assign n20786 = pi759 & pi947;
  assign n20787 = n16508 & ~n20786;
  assign n20788 = ~n20323 & n20787;
  assign n20789 = ~pi152 & ~n16508;
  assign n20790 = pi38 & ~n20789;
  assign n20791 = ~n20788 & n20790;
  assign n20792 = pi759 & n20511;
  assign n20793 = pi152 & ~n16201;
  assign n20794 = ~pi39 & ~n20793;
  assign n20795 = ~n20792 & n20794;
  assign n20796 = ~n20425 & n20795;
  assign n20797 = ~pi947 & n16269;
  assign n20798 = pi223 & ~n20797;
  assign n20799 = ~pi152 & ~n16269;
  assign n20800 = n20798 & ~n20799;
  assign n20801 = ~pi299 & ~n20800;
  assign n20802 = n16269 & ~n20323;
  assign n20803 = pi223 & ~n20802;
  assign n20804 = ~n20799 & n20803;
  assign n20805 = pi152 & ~n16207;
  assign n20806 = ~n20729 & ~n20805;
  assign n20807 = n2607 & n20806;
  assign n20808 = ~pi152 & n16329;
  assign n20809 = ~pi947 & ~n16329;
  assign n20810 = ~n2607 & ~n20809;
  assign n20811 = ~n20808 & n20810;
  assign n20812 = ~n6192 & ~n16329;
  assign n20813 = ~n2607 & ~n20812;
  assign n20814 = ~n20811 & n20813;
  assign n20815 = ~pi223 & ~n20814;
  assign n20816 = ~n20807 & n20815;
  assign n20817 = ~n20804 & ~n20816;
  assign n20818 = n20801 & n20817;
  assign n20819 = ~pi152 & ~n16346;
  assign n20820 = n20429 & ~n20819;
  assign n20821 = n2527 & n20806;
  assign n20822 = ~pi215 & ~n20821;
  assign n20823 = pi152 & n20432;
  assign n20824 = n20413 & ~n20823;
  assign n20825 = ~n16340 & n20824;
  assign n20826 = n20822 & ~n20825;
  assign n20827 = pi299 & ~n20826;
  assign n20828 = ~n20820 & n20827;
  assign n20829 = pi759 & ~n20828;
  assign n20830 = ~n20818 & n20829;
  assign n20831 = ~n20415 & ~n20805;
  assign n20832 = n2607 & ~n20831;
  assign n20833 = ~n16329 & ~n20323;
  assign n20834 = ~n2607 & ~n20833;
  assign n20835 = ~n20808 & n20834;
  assign n20836 = ~n20832 & ~n20835;
  assign n20837 = ~pi223 & ~n20836;
  assign n20838 = ~pi299 & ~n20804;
  assign n20839 = ~n20837 & n20838;
  assign n20840 = ~n20323 & ~n20474;
  assign n20841 = n20820 & ~n20840;
  assign n20842 = ~n20430 & n20822;
  assign n20843 = ~n20824 & n20842;
  assign n20844 = ~n20841 & ~n20843;
  assign n20845 = pi299 & n20844;
  assign n20846 = ~pi759 & ~n20845;
  assign n20847 = ~n20839 & n20846;
  assign n20848 = ~n20830 & ~n20847;
  assign n20849 = pi39 & n20848;
  assign n20850 = ~pi38 & ~n20849;
  assign n20851 = ~n20796 & n20850;
  assign n20852 = pi696 & ~n20851;
  assign n20853 = ~n20791 & n20852;
  assign n20854 = ~pi759 & ~n16355;
  assign n20855 = pi152 & n20854;
  assign n20856 = ~n20517 & ~n20805;
  assign n20857 = n2607 & ~n20856;
  assign n20858 = ~n20811 & ~n20857;
  assign n20859 = ~pi223 & ~n20858;
  assign n20860 = n20801 & ~n20859;
  assign n20861 = pi152 & n20496;
  assign n20862 = n2527 & n20856;
  assign n20863 = ~n20825 & ~n20862;
  assign n20864 = n20494 & n20863;
  assign n20865 = ~n20861 & ~n20864;
  assign n20866 = n20515 & n20865;
  assign n20867 = ~n20860 & ~n20866;
  assign n20868 = pi759 & n20867;
  assign n20869 = ~n20855 & ~n20868;
  assign n20870 = pi39 & n20869;
  assign n20871 = ~pi38 & ~n20870;
  assign n20872 = ~n20795 & n20871;
  assign n20873 = ~pi152 & ~n16524;
  assign n20874 = pi38 & ~n20873;
  assign n20875 = ~n20787 & n20874;
  assign n20876 = ~pi696 & ~n20875;
  assign n20877 = ~n20872 & n20876;
  assign n20878 = ~n20853 & ~n20877;
  assign n20879 = n10021 & ~n20878;
  assign n20880 = ~pi152 & ~n10021;
  assign n20881 = ~pi832 & ~n20880;
  assign n20882 = ~n20879 & n20881;
  assign n20883 = pi696 & n20323;
  assign n20884 = ~n20786 & ~n20883;
  assign n20885 = n2934 & n20884;
  assign n20886 = ~pi152 & ~n2934;
  assign n20887 = pi832 & ~n20886;
  assign n20888 = ~n20885 & n20887;
  assign po309 = n20882 | n20888;
  assign n20890 = pi766 & pi947;
  assign n20891 = pi700 & n20323;
  assign n20892 = ~n20890 & ~n20891;
  assign n20893 = n2934 & n20892;
  assign n20894 = pi153 & ~n2934;
  assign n20895 = pi832 & ~n20894;
  assign n20896 = ~n20893 & n20895;
  assign n20897 = ~pi153 & ~n20537;
  assign n20898 = ~pi153 & ~n16201;
  assign n20899 = ~pi766 & n17520;
  assign n20900 = ~n20512 & ~n20899;
  assign n20901 = ~n20898 & ~n20900;
  assign n20902 = ~n20425 & n20901;
  assign n20903 = pi153 & ~n16346;
  assign n20904 = n20429 & ~n20903;
  assign n20905 = pi153 & n20724;
  assign n20906 = ~n16339 & ~n20905;
  assign n20907 = ~pi153 & ~n16207;
  assign n20908 = n20518 & ~n20907;
  assign n20909 = ~n20414 & n20908;
  assign n20910 = ~pi215 & ~n20909;
  assign n20911 = n20906 & n20910;
  assign n20912 = ~n20904 & ~n20911;
  assign n20913 = pi299 & ~n20912;
  assign n20914 = pi153 & ~n20735;
  assign n20915 = ~n20466 & ~n20914;
  assign n20916 = ~n20913 & ~n20915;
  assign n20917 = pi766 & ~n20916;
  assign n20918 = n20474 & ~n20904;
  assign n20919 = n20416 & ~n20907;
  assign n20920 = ~n20433 & ~n20919;
  assign n20921 = n20906 & n20920;
  assign n20922 = ~pi215 & ~n20921;
  assign n20923 = ~n20918 & ~n20922;
  assign n20924 = ~n20438 & n20923;
  assign n20925 = pi299 & ~n20924;
  assign n20926 = ~pi153 & ~n16333;
  assign n20927 = n20422 & ~n20926;
  assign n20928 = ~pi766 & ~n20927;
  assign n20929 = ~n20925 & n20928;
  assign n20930 = pi39 & ~n20929;
  assign n20931 = ~n20917 & n20930;
  assign n20932 = ~n20902 & ~n20931;
  assign n20933 = ~pi38 & ~n20932;
  assign n20934 = ~n20323 & ~n20890;
  assign n20935 = n16508 & ~n20934;
  assign n20936 = ~pi153 & ~n16508;
  assign n20937 = pi38 & ~n20936;
  assign n20938 = ~n20935 & n20937;
  assign n20939 = ~n20933 & ~n20938;
  assign n20940 = pi700 & ~n20939;
  assign n20941 = pi153 & ~n16524;
  assign n20942 = n16508 & ~n20890;
  assign n20943 = ~n20941 & ~n20942;
  assign n20944 = pi38 & n20943;
  assign n20945 = ~pi153 & ~pi766;
  assign n20946 = ~n16355 & n20945;
  assign n20947 = n20514 & ~n20926;
  assign n20948 = n20494 & ~n20908;
  assign n20949 = n20906 & n20948;
  assign n20950 = n20496 & ~n20903;
  assign n20951 = pi299 & ~n20950;
  assign n20952 = ~n20949 & n20951;
  assign n20953 = ~n20947 & ~n20952;
  assign n20954 = pi766 & n20953;
  assign n20955 = ~n20946 & ~n20954;
  assign n20956 = pi39 & n20955;
  assign n20957 = ~pi38 & ~n20901;
  assign n20958 = ~n20956 & n20957;
  assign n20959 = ~pi700 & ~n20958;
  assign n20960 = ~n20944 & n20959;
  assign n20961 = ~n20940 & ~n20960;
  assign n20962 = n20537 & n20961;
  assign n20963 = ~pi57 & ~n20962;
  assign n20964 = ~n20897 & n20963;
  assign n20965 = pi57 & pi153;
  assign n20966 = ~pi832 & ~n20965;
  assign n20967 = ~n20964 & n20966;
  assign po310 = n20896 | n20967;
  assign n20969 = ~pi742 & pi947;
  assign n20970 = ~pi704 & n20323;
  assign n20971 = ~n20969 & ~n20970;
  assign n20972 = n2934 & ~n20971;
  assign n20973 = ~pi154 & ~n2934;
  assign n20974 = pi832 & ~n20973;
  assign n20975 = ~n20972 & n20974;
  assign n20976 = ~pi154 & ~n16526;
  assign n20977 = pi742 & n20976;
  assign n20978 = ~pi154 & ~n16201;
  assign n20979 = n20512 & ~n20978;
  assign n20980 = ~pi154 & ~n20501;
  assign n20981 = pi154 & n20522;
  assign n20982 = pi39 & ~n20981;
  assign n20983 = ~n20980 & n20982;
  assign n20984 = ~n20979 & ~n20983;
  assign n20985 = ~pi38 & ~n20984;
  assign n20986 = ~pi154 & ~n16524;
  assign n20987 = ~n20510 & ~n20986;
  assign n20988 = ~pi742 & ~n20987;
  assign n20989 = ~n20985 & n20988;
  assign n20990 = pi704 & ~n20989;
  assign n20991 = ~n20977 & n20990;
  assign n20992 = ~pi154 & ~n16508;
  assign n20993 = n20460 & ~n20992;
  assign n20994 = n20426 & ~n20978;
  assign n20995 = ~n20469 & n20994;
  assign n20996 = ~pi154 & ~n20467;
  assign n20997 = pi154 & ~n20478;
  assign n20998 = pi39 & ~n20997;
  assign n20999 = ~n20996 & n20998;
  assign n21000 = ~n20995 & ~n20999;
  assign n21001 = ~pi38 & ~n21000;
  assign n21002 = ~pi742 & ~n21001;
  assign n21003 = ~n20993 & n21002;
  assign n21004 = n20453 & ~n20992;
  assign n21005 = ~pi154 & n20443;
  assign n21006 = pi154 & n20423;
  assign n21007 = ~n21005 & ~n21006;
  assign n21008 = pi39 & n21007;
  assign n21009 = ~n20994 & ~n21008;
  assign n21010 = ~pi38 & ~n21009;
  assign n21011 = pi742 & ~n21010;
  assign n21012 = ~n21004 & n21011;
  assign n21013 = ~pi704 & ~n21012;
  assign n21014 = ~n21003 & n21013;
  assign n21015 = n10021 & ~n21014;
  assign n21016 = ~n20991 & n21015;
  assign n21017 = ~pi154 & ~n10021;
  assign n21018 = ~pi832 & ~n21017;
  assign n21019 = ~n21016 & n21018;
  assign po311 = ~n20975 & ~n21019;
  assign n21021 = ~pi757 & n20526;
  assign n21022 = pi686 & ~n21021;
  assign n21023 = ~pi38 & ~n20480;
  assign n21024 = ~n20460 & ~n21023;
  assign n21025 = ~pi757 & n21024;
  assign n21026 = ~pi38 & ~n20427;
  assign n21027 = ~n20453 & ~n21026;
  assign n21028 = pi757 & n21027;
  assign n21029 = ~pi686 & ~n21028;
  assign n21030 = ~n21025 & n21029;
  assign n21031 = n10021 & ~n21030;
  assign n21032 = ~n21022 & n21031;
  assign n21033 = pi155 & ~n21032;
  assign n21034 = ~pi38 & ~n20447;
  assign n21035 = n16212 & ~n20323;
  assign n21036 = n18931 & n21035;
  assign n21037 = ~n21034 & ~n21036;
  assign n21038 = pi757 & n21037;
  assign n21039 = ~pi38 & ~n20472;
  assign n21040 = pi38 & n20457;
  assign n21041 = ~n21039 & ~n21040;
  assign n21042 = ~pi757 & n21041;
  assign n21043 = ~pi686 & ~n21042;
  assign n21044 = ~n21038 & n21043;
  assign n21045 = ~pi757 & n20505;
  assign n21046 = pi757 & ~n16526;
  assign n21047 = ~n21045 & ~n21046;
  assign n21048 = pi686 & n21047;
  assign n21049 = ~n21044 & ~n21048;
  assign n21050 = ~pi155 & ~n21049;
  assign n21051 = n10021 & n21050;
  assign n21052 = ~n21033 & ~n21051;
  assign n21053 = ~pi832 & ~n21052;
  assign n21054 = ~pi757 & pi947;
  assign n21055 = ~pi686 & n20323;
  assign n21056 = ~n21054 & ~n21055;
  assign n21057 = n2934 & ~n21056;
  assign n21058 = ~pi155 & ~n2934;
  assign n21059 = pi832 & ~n21058;
  assign n21060 = ~n21057 & n21059;
  assign po312 = ~n21053 & ~n21060;
  assign n21062 = ~pi741 & pi947;
  assign n21063 = ~pi724 & n20323;
  assign n21064 = ~n21062 & ~n21063;
  assign n21065 = n2934 & ~n21064;
  assign n21066 = ~pi156 & ~n2934;
  assign n21067 = pi832 & ~n21066;
  assign n21068 = ~n21065 & n21067;
  assign n21069 = pi741 & ~n21037;
  assign n21070 = ~pi741 & ~n21041;
  assign n21071 = ~pi724 & ~n21070;
  assign n21072 = ~n21069 & n21071;
  assign n21073 = ~pi741 & ~n20505;
  assign n21074 = pi741 & n16526;
  assign n21075 = ~n21073 & ~n21074;
  assign n21076 = pi724 & n21075;
  assign n21077 = ~n21072 & ~n21076;
  assign n21078 = n10021 & n21077;
  assign n21079 = ~pi156 & ~n21078;
  assign n21080 = ~pi832 & ~n21079;
  assign n21081 = pi741 & ~n21027;
  assign n21082 = ~pi741 & ~n21024;
  assign n21083 = ~pi724 & ~n21082;
  assign n21084 = ~n21081 & n21083;
  assign n21085 = pi724 & ~pi741;
  assign n21086 = n20526 & n21085;
  assign n21087 = ~n21084 & ~n21086;
  assign n21088 = pi156 & ~n21087;
  assign n21089 = n10021 & n21088;
  assign n21090 = n21080 & ~n21089;
  assign po313 = ~n21068 & ~n21090;
  assign n21092 = ~pi760 & pi947;
  assign n21093 = ~pi688 & n20323;
  assign n21094 = ~n21092 & ~n21093;
  assign n21095 = n2934 & ~n21094;
  assign n21096 = ~pi157 & ~n2934;
  assign n21097 = pi832 & ~n21096;
  assign n21098 = ~n21095 & n21097;
  assign n21099 = pi157 & ~n16524;
  assign n21100 = n16508 & ~n21092;
  assign n21101 = pi38 & ~n21100;
  assign n21102 = ~n21099 & n21101;
  assign n21103 = ~pi157 & ~n16333;
  assign n21104 = n20514 & ~n21103;
  assign n21105 = ~pi157 & ~n20497;
  assign n21106 = ~n13365 & ~n20521;
  assign n21107 = ~n21105 & ~n21106;
  assign n21108 = ~pi760 & ~n21107;
  assign n21109 = ~n21104 & n21108;
  assign n21110 = ~pi157 & pi760;
  assign n21111 = ~n16355 & n21110;
  assign n21112 = pi39 & ~n21111;
  assign n21113 = ~n21109 & n21112;
  assign n21114 = ~pi157 & ~n16201;
  assign n21115 = ~pi39 & ~n21114;
  assign n21116 = n16201 & n21092;
  assign n21117 = n21115 & ~n21116;
  assign n21118 = ~pi38 & ~n21117;
  assign n21119 = ~n21113 & n21118;
  assign n21120 = ~n21102 & ~n21119;
  assign n21121 = pi688 & ~n21120;
  assign n21122 = ~n20425 & n21117;
  assign n21123 = pi760 & ~n20423;
  assign n21124 = pi157 & ~n21123;
  assign n21125 = ~pi760 & n20478;
  assign n21126 = n21124 & ~n21125;
  assign n21127 = pi760 & ~n20443;
  assign n21128 = ~pi760 & n20467;
  assign n21129 = ~pi157 & ~n21128;
  assign n21130 = ~n21127 & n21129;
  assign n21131 = pi39 & ~n21130;
  assign n21132 = ~n21126 & n21131;
  assign n21133 = ~n21122 & ~n21132;
  assign n21134 = ~pi38 & ~n21133;
  assign n21135 = pi157 & ~n16508;
  assign n21136 = ~n21100 & ~n21135;
  assign n21137 = n20453 & ~n21136;
  assign n21138 = ~pi688 & ~n21137;
  assign n21139 = ~n21134 & n21138;
  assign n21140 = ~n21121 & ~n21139;
  assign n21141 = n10021 & ~n21140;
  assign n21142 = ~pi157 & ~n10021;
  assign n21143 = ~pi832 & ~n21142;
  assign n21144 = ~n21141 & n21143;
  assign po314 = ~n21098 & ~n21144;
  assign n21146 = ~pi158 & n20501;
  assign n21147 = pi158 & ~n20522;
  assign n21148 = ~pi753 & ~n21147;
  assign n21149 = ~n21146 & n21148;
  assign n21150 = ~pi158 & ~n16355;
  assign n21151 = pi753 & n21150;
  assign n21152 = ~n21149 & ~n21151;
  assign n21153 = pi39 & ~n21152;
  assign n21154 = pi158 & ~n16201;
  assign n21155 = pi753 & n16201;
  assign n21156 = ~n21154 & ~n21155;
  assign n21157 = n20490 & n21156;
  assign n21158 = ~pi38 & ~n21157;
  assign n21159 = ~n21153 & n21158;
  assign n21160 = pi158 & ~n16524;
  assign n21161 = ~pi753 & pi947;
  assign n21162 = n16508 & ~n21161;
  assign n21163 = ~n21160 & ~n21162;
  assign n21164 = pi38 & ~n21163;
  assign n21165 = pi702 & ~n21164;
  assign n21166 = ~n21159 & n21165;
  assign n21167 = ~pi158 & ~n20443;
  assign n21168 = pi158 & ~n20423;
  assign n21169 = pi753 & ~n21168;
  assign n21170 = ~n21167 & n21169;
  assign n21171 = ~pi158 & n20467;
  assign n21172 = pi158 & n20478;
  assign n21173 = ~pi753 & ~n21172;
  assign n21174 = ~n21171 & n21173;
  assign n21175 = ~n21170 & ~n21174;
  assign n21176 = pi39 & ~n21175;
  assign n21177 = n20445 & ~n21161;
  assign n21178 = ~pi39 & ~n21177;
  assign n21179 = ~n21154 & n21178;
  assign n21180 = ~pi38 & ~n21179;
  assign n21181 = ~n21176 & n21180;
  assign n21182 = pi158 & ~n16508;
  assign n21183 = ~n21162 & ~n21182;
  assign n21184 = n20453 & ~n21183;
  assign n21185 = ~pi702 & ~n21184;
  assign n21186 = ~n21181 & n21185;
  assign n21187 = ~n21166 & ~n21186;
  assign n21188 = n10021 & ~n21187;
  assign n21189 = ~pi158 & ~n10021;
  assign n21190 = ~pi832 & ~n21189;
  assign n21191 = ~n21188 & n21190;
  assign n21192 = ~pi702 & n20323;
  assign n21193 = ~n21161 & ~n21192;
  assign n21194 = n2934 & ~n21193;
  assign n21195 = ~pi158 & ~n2934;
  assign n21196 = pi832 & ~n21195;
  assign n21197 = ~n21194 & n21196;
  assign po315 = ~n21191 & ~n21197;
  assign n21199 = ~pi159 & n20501;
  assign n21200 = pi159 & ~n20522;
  assign n21201 = ~pi754 & ~n21200;
  assign n21202 = ~n21199 & n21201;
  assign n21203 = ~pi159 & ~n16355;
  assign n21204 = pi754 & n21203;
  assign n21205 = ~n21202 & ~n21204;
  assign n21206 = pi39 & ~n21205;
  assign n21207 = pi159 & ~n16201;
  assign n21208 = pi754 & n16201;
  assign n21209 = ~n21207 & ~n21208;
  assign n21210 = n20490 & n21209;
  assign n21211 = ~pi38 & ~n21210;
  assign n21212 = ~n21206 & n21211;
  assign n21213 = pi159 & ~n16524;
  assign n21214 = ~pi754 & pi947;
  assign n21215 = n16508 & ~n21214;
  assign n21216 = ~n21213 & ~n21215;
  assign n21217 = pi38 & ~n21216;
  assign n21218 = pi709 & ~n21217;
  assign n21219 = ~n21212 & n21218;
  assign n21220 = ~pi159 & ~n20443;
  assign n21221 = pi159 & ~n20423;
  assign n21222 = pi754 & ~n21221;
  assign n21223 = ~n21220 & n21222;
  assign n21224 = ~pi159 & n20467;
  assign n21225 = pi159 & n20478;
  assign n21226 = ~pi754 & ~n21225;
  assign n21227 = ~n21224 & n21226;
  assign n21228 = ~n21223 & ~n21227;
  assign n21229 = pi39 & ~n21228;
  assign n21230 = n20445 & ~n21214;
  assign n21231 = ~pi39 & ~n21230;
  assign n21232 = ~n21207 & n21231;
  assign n21233 = ~pi38 & ~n21232;
  assign n21234 = ~n21229 & n21233;
  assign n21235 = pi159 & ~n16508;
  assign n21236 = ~n21215 & ~n21235;
  assign n21237 = n20453 & ~n21236;
  assign n21238 = ~pi709 & ~n21237;
  assign n21239 = ~n21234 & n21238;
  assign n21240 = ~n21219 & ~n21239;
  assign n21241 = n10021 & ~n21240;
  assign n21242 = ~pi159 & ~n10021;
  assign n21243 = ~pi832 & ~n21242;
  assign n21244 = ~n21241 & n21243;
  assign n21245 = ~pi709 & n20323;
  assign n21246 = ~n21214 & ~n21245;
  assign n21247 = n2934 & ~n21246;
  assign n21248 = ~pi159 & ~n2934;
  assign n21249 = pi832 & ~n21248;
  assign n21250 = ~n21247 & n21249;
  assign po316 = ~n21244 & ~n21250;
  assign n21252 = ~pi756 & pi947;
  assign n21253 = ~pi734 & n20323;
  assign n21254 = ~n21252 & ~n21253;
  assign n21255 = n2934 & ~n21254;
  assign n21256 = ~pi160 & ~n2934;
  assign n21257 = pi832 & ~n21256;
  assign n21258 = ~n21255 & n21257;
  assign n21259 = pi160 & ~n16524;
  assign n21260 = n16508 & ~n21252;
  assign n21261 = pi38 & ~n21260;
  assign n21262 = ~n21259 & n21261;
  assign n21263 = ~pi160 & ~n16333;
  assign n21264 = n20514 & ~n21263;
  assign n21265 = pi160 & ~n20573;
  assign n21266 = ~pi160 & ~n20497;
  assign n21267 = ~n21265 & ~n21266;
  assign n21268 = pi299 & n21267;
  assign n21269 = ~pi756 & ~n21268;
  assign n21270 = ~n21264 & n21269;
  assign n21271 = ~pi160 & pi756;
  assign n21272 = ~n16355 & n21271;
  assign n21273 = pi39 & ~n21272;
  assign n21274 = ~n21270 & n21273;
  assign n21275 = ~pi160 & ~n16201;
  assign n21276 = ~pi39 & ~n21275;
  assign n21277 = n16201 & n21252;
  assign n21278 = n21276 & ~n21277;
  assign n21279 = ~pi38 & ~n21278;
  assign n21280 = ~n21274 & n21279;
  assign n21281 = ~n21262 & ~n21280;
  assign n21282 = pi734 & ~n21281;
  assign n21283 = ~n20425 & n21278;
  assign n21284 = ~pi160 & n20440;
  assign n21285 = pi160 & ~n20549;
  assign n21286 = ~n20442 & ~n21285;
  assign n21287 = pi756 & n21286;
  assign n21288 = ~n21284 & n21287;
  assign n21289 = pi160 & n20478;
  assign n21290 = ~pi160 & n20467;
  assign n21291 = ~pi756 & ~n21290;
  assign n21292 = ~n21289 & n21291;
  assign n21293 = pi39 & ~n21292;
  assign n21294 = ~n21288 & n21293;
  assign n21295 = ~n21283 & ~n21294;
  assign n21296 = ~pi38 & ~n21295;
  assign n21297 = pi160 & ~n16508;
  assign n21298 = ~n21260 & ~n21297;
  assign n21299 = n20453 & ~n21298;
  assign n21300 = ~pi734 & ~n21299;
  assign n21301 = ~n21296 & n21300;
  assign n21302 = ~n21282 & ~n21301;
  assign n21303 = n10021 & ~n21302;
  assign n21304 = ~pi160 & ~n10021;
  assign n21305 = ~pi832 & ~n21304;
  assign n21306 = ~n21303 & n21305;
  assign po317 = ~n21258 & ~n21306;
  assign n21308 = pi758 & pi947;
  assign n21309 = n16508 & ~n21308;
  assign n21310 = ~n20323 & n21309;
  assign n21311 = ~pi161 & ~n16508;
  assign n21312 = pi38 & ~n21311;
  assign n21313 = ~n21310 & n21312;
  assign n21314 = pi758 & n20511;
  assign n21315 = pi161 & ~n16201;
  assign n21316 = ~pi39 & ~n21315;
  assign n21317 = ~n21314 & n21316;
  assign n21318 = ~n20425 & n21317;
  assign n21319 = ~pi161 & ~n16269;
  assign n21320 = n20798 & ~n21319;
  assign n21321 = ~pi299 & ~n21320;
  assign n21322 = n20803 & ~n21319;
  assign n21323 = pi161 & ~n16207;
  assign n21324 = ~n20729 & ~n21323;
  assign n21325 = n2607 & n21324;
  assign n21326 = ~pi161 & n16329;
  assign n21327 = n20810 & ~n21326;
  assign n21328 = n20813 & ~n21327;
  assign n21329 = ~pi223 & ~n21328;
  assign n21330 = ~n21325 & n21329;
  assign n21331 = ~n21322 & ~n21330;
  assign n21332 = n21321 & n21331;
  assign n21333 = ~pi161 & ~n16346;
  assign n21334 = n20429 & ~n21333;
  assign n21335 = n2527 & n21324;
  assign n21336 = ~pi215 & ~n21335;
  assign n21337 = pi161 & n20432;
  assign n21338 = n20413 & ~n21337;
  assign n21339 = ~n16340 & n21338;
  assign n21340 = n21336 & ~n21339;
  assign n21341 = pi299 & ~n21340;
  assign n21342 = ~n21334 & n21341;
  assign n21343 = pi758 & ~n21342;
  assign n21344 = ~n21332 & n21343;
  assign n21345 = ~n20415 & ~n21323;
  assign n21346 = n2607 & ~n21345;
  assign n21347 = n20834 & ~n21326;
  assign n21348 = ~n21346 & ~n21347;
  assign n21349 = ~pi223 & ~n21348;
  assign n21350 = ~pi299 & ~n21322;
  assign n21351 = ~n21349 & n21350;
  assign n21352 = ~n20840 & n21334;
  assign n21353 = ~n20430 & n21336;
  assign n21354 = ~n21338 & n21353;
  assign n21355 = ~n21352 & ~n21354;
  assign n21356 = pi299 & n21355;
  assign n21357 = ~pi758 & ~n21356;
  assign n21358 = ~n21351 & n21357;
  assign n21359 = ~n21344 & ~n21358;
  assign n21360 = pi39 & n21359;
  assign n21361 = ~pi38 & ~n21360;
  assign n21362 = ~n21318 & n21361;
  assign n21363 = pi736 & ~n21362;
  assign n21364 = ~n21313 & n21363;
  assign n21365 = pi161 & n19327;
  assign n21366 = ~n20517 & ~n21323;
  assign n21367 = n2607 & ~n21366;
  assign n21368 = ~n21327 & ~n21367;
  assign n21369 = ~pi223 & ~n21368;
  assign n21370 = n21321 & ~n21369;
  assign n21371 = pi161 & n20496;
  assign n21372 = n2527 & n21366;
  assign n21373 = ~n21339 & ~n21372;
  assign n21374 = n20494 & n21373;
  assign n21375 = ~n21371 & ~n21374;
  assign n21376 = n20515 & n21375;
  assign n21377 = ~n21370 & ~n21376;
  assign n21378 = pi758 & n21377;
  assign n21379 = ~n21365 & ~n21378;
  assign n21380 = pi39 & n21379;
  assign n21381 = ~pi38 & ~n21380;
  assign n21382 = ~n21317 & n21381;
  assign n21383 = ~pi161 & ~n16524;
  assign n21384 = pi38 & ~n21383;
  assign n21385 = ~n21309 & n21384;
  assign n21386 = ~pi736 & ~n21385;
  assign n21387 = ~n21382 & n21386;
  assign n21388 = ~n21364 & ~n21387;
  assign n21389 = n10021 & ~n21388;
  assign n21390 = ~pi161 & ~n10021;
  assign n21391 = ~pi832 & ~n21390;
  assign n21392 = ~n21389 & n21391;
  assign n21393 = pi736 & n20323;
  assign n21394 = ~n21308 & ~n21393;
  assign n21395 = n2934 & n21394;
  assign n21396 = ~pi161 & ~n2934;
  assign n21397 = pi832 & ~n21396;
  assign n21398 = ~n21395 & n21397;
  assign po318 = n21392 | n21398;
  assign n21400 = pi162 & ~n16524;
  assign n21401 = ~pi761 & pi947;
  assign n21402 = n16508 & ~n21401;
  assign n21403 = pi38 & ~n21402;
  assign n21404 = ~n21400 & n21403;
  assign n21405 = pi761 & n16355;
  assign n21406 = ~pi761 & n20499;
  assign n21407 = ~pi162 & ~n21406;
  assign n21408 = ~n21405 & n21407;
  assign n21409 = n14471 & ~n20573;
  assign n21410 = ~n20500 & ~n21409;
  assign n21411 = ~pi761 & ~n21410;
  assign n21412 = pi39 & ~n21411;
  assign n21413 = ~n21408 & n21412;
  assign n21414 = ~pi162 & ~n16201;
  assign n21415 = ~pi39 & ~n21414;
  assign n21416 = n16201 & n21401;
  assign n21417 = n21415 & ~n21416;
  assign n21418 = ~pi38 & ~n21417;
  assign n21419 = ~n21413 & n21418;
  assign n21420 = ~n21404 & ~n21419;
  assign n21421 = pi738 & ~n21420;
  assign n21422 = ~n20425 & n21417;
  assign n21423 = pi162 & ~n20549;
  assign n21424 = ~n14471 & ~n20443;
  assign n21425 = pi761 & ~n21424;
  assign n21426 = ~n21423 & n21425;
  assign n21427 = pi162 & n20478;
  assign n21428 = ~pi162 & n20467;
  assign n21429 = ~pi761 & ~n21428;
  assign n21430 = ~n21427 & n21429;
  assign n21431 = pi39 & ~n21430;
  assign n21432 = ~n21426 & n21431;
  assign n21433 = ~n21422 & ~n21432;
  assign n21434 = ~pi38 & ~n21433;
  assign n21435 = pi162 & ~n16508;
  assign n21436 = ~n21402 & ~n21435;
  assign n21437 = n20453 & ~n21436;
  assign n21438 = ~pi738 & ~n21437;
  assign n21439 = ~n21434 & n21438;
  assign n21440 = ~n21421 & ~n21439;
  assign n21441 = n10021 & ~n21440;
  assign n21442 = ~pi162 & ~n10021;
  assign n21443 = ~pi832 & ~n21442;
  assign n21444 = ~n21441 & n21443;
  assign n21445 = ~pi738 & n20323;
  assign n21446 = ~n21401 & ~n21445;
  assign n21447 = n2934 & ~n21446;
  assign n21448 = ~pi162 & ~n2934;
  assign n21449 = pi832 & ~n21448;
  assign n21450 = ~n21447 & n21449;
  assign po319 = ~n21444 & ~n21450;
  assign n21452 = ~pi777 & pi947;
  assign n21453 = ~pi737 & n20323;
  assign n21454 = ~n21452 & ~n21453;
  assign n21455 = n2934 & ~n21454;
  assign n21456 = ~pi163 & ~n2934;
  assign n21457 = pi832 & ~n21456;
  assign n21458 = ~n21455 & n21457;
  assign n21459 = pi163 & ~n16524;
  assign n21460 = n16508 & ~n21452;
  assign n21461 = pi38 & ~n21460;
  assign n21462 = ~n21459 & n21461;
  assign n21463 = ~pi163 & ~n16333;
  assign n21464 = n20514 & ~n21463;
  assign n21465 = ~pi163 & ~n20497;
  assign n21466 = ~n14017 & ~n20521;
  assign n21467 = ~n21465 & ~n21466;
  assign n21468 = ~pi777 & ~n21467;
  assign n21469 = ~n21464 & n21468;
  assign n21470 = ~pi163 & pi777;
  assign n21471 = ~n16355 & n21470;
  assign n21472 = pi39 & ~n21471;
  assign n21473 = ~n21469 & n21472;
  assign n21474 = ~pi163 & ~n16201;
  assign n21475 = ~pi39 & ~n21474;
  assign n21476 = n16201 & n21452;
  assign n21477 = n21475 & ~n21476;
  assign n21478 = ~pi38 & ~n21477;
  assign n21479 = ~n21473 & n21478;
  assign n21480 = ~n21462 & ~n21479;
  assign n21481 = pi737 & ~n21480;
  assign n21482 = ~n20425 & n21477;
  assign n21483 = ~pi163 & n20467;
  assign n21484 = pi163 & n20478;
  assign n21485 = ~pi777 & ~n21484;
  assign n21486 = ~n21483 & n21485;
  assign n21487 = pi163 & ~n20549;
  assign n21488 = n14017 & ~n20439;
  assign n21489 = pi777 & ~n21488;
  assign n21490 = ~n20442 & n21489;
  assign n21491 = ~n21487 & n21490;
  assign n21492 = pi39 & ~n21491;
  assign n21493 = ~n21486 & n21492;
  assign n21494 = ~n21482 & ~n21493;
  assign n21495 = ~pi38 & ~n21494;
  assign n21496 = pi163 & ~n16508;
  assign n21497 = ~n21460 & ~n21496;
  assign n21498 = n20453 & ~n21497;
  assign n21499 = ~pi737 & ~n21498;
  assign n21500 = ~n21495 & n21499;
  assign n21501 = ~n21481 & ~n21500;
  assign n21502 = n10021 & ~n21501;
  assign n21503 = ~pi163 & ~n10021;
  assign n21504 = ~pi832 & ~n21503;
  assign n21505 = ~n21502 & n21504;
  assign po320 = ~n21458 & ~n21505;
  assign n21507 = ~pi752 & pi947;
  assign n21508 = pi703 & n20323;
  assign n21509 = ~n21507 & ~n21508;
  assign n21510 = n2934 & ~n21509;
  assign n21511 = ~pi164 & ~n2934;
  assign n21512 = pi832 & ~n21511;
  assign n21513 = ~n21510 & n21512;
  assign n21514 = pi164 & n20480;
  assign n21515 = ~pi164 & n20472;
  assign n21516 = ~pi38 & ~n21515;
  assign n21517 = ~n21514 & n21516;
  assign n21518 = ~pi164 & ~n20457;
  assign n21519 = n20460 & ~n21518;
  assign n21520 = ~pi752 & ~n21519;
  assign n21521 = ~n21517 & n21520;
  assign n21522 = pi164 & n20427;
  assign n21523 = ~pi164 & n20447;
  assign n21524 = ~pi38 & ~n21523;
  assign n21525 = ~n21522 & n21524;
  assign n21526 = ~pi164 & ~n16508;
  assign n21527 = n20453 & ~n21526;
  assign n21528 = pi752 & ~n21527;
  assign n21529 = ~n21525 & n21528;
  assign n21530 = ~n21521 & ~n21529;
  assign n21531 = pi703 & ~n21530;
  assign n21532 = pi164 & ~n20488;
  assign n21533 = ~pi752 & ~n20505;
  assign n21534 = ~n21532 & n21533;
  assign n21535 = pi752 & n16526;
  assign n21536 = ~pi752 & n20526;
  assign n21537 = pi164 & ~n21536;
  assign n21538 = ~pi703 & ~n21537;
  assign n21539 = ~n21535 & n21538;
  assign n21540 = ~n21534 & n21539;
  assign n21541 = ~n21531 & ~n21540;
  assign n21542 = n10021 & ~n21541;
  assign n21543 = ~pi164 & ~n10021;
  assign n21544 = ~pi832 & ~n21543;
  assign n21545 = ~n21542 & n21544;
  assign po321 = ~n21513 & ~n21545;
  assign n21547 = ~pi774 & pi947;
  assign n21548 = pi687 & n20323;
  assign n21549 = ~n21547 & ~n21548;
  assign n21550 = n2934 & ~n21549;
  assign n21551 = ~pi165 & ~n2934;
  assign n21552 = pi832 & ~n21551;
  assign n21553 = ~n21550 & n21552;
  assign n21554 = pi165 & n20480;
  assign n21555 = ~pi165 & n20472;
  assign n21556 = ~pi38 & ~n21555;
  assign n21557 = ~n21554 & n21556;
  assign n21558 = ~pi165 & ~n20457;
  assign n21559 = n20460 & ~n21558;
  assign n21560 = ~pi774 & ~n21559;
  assign n21561 = ~n21557 & n21560;
  assign n21562 = pi165 & n20427;
  assign n21563 = ~pi165 & n20447;
  assign n21564 = ~pi38 & ~n21563;
  assign n21565 = ~n21562 & n21564;
  assign n21566 = ~pi165 & ~n16508;
  assign n21567 = n20453 & ~n21566;
  assign n21568 = pi774 & ~n21567;
  assign n21569 = ~n21565 & n21568;
  assign n21570 = ~n21561 & ~n21569;
  assign n21571 = pi687 & ~n21570;
  assign n21572 = pi165 & ~n20488;
  assign n21573 = ~pi774 & ~n20505;
  assign n21574 = ~n21572 & n21573;
  assign n21575 = pi774 & n16526;
  assign n21576 = ~pi774 & n20526;
  assign n21577 = pi165 & ~n21576;
  assign n21578 = ~pi687 & ~n21577;
  assign n21579 = ~n21575 & n21578;
  assign n21580 = ~n21574 & n21579;
  assign n21581 = ~n21571 & ~n21580;
  assign n21582 = n10021 & ~n21581;
  assign n21583 = ~pi165 & ~n10021;
  assign n21584 = ~pi832 & ~n21583;
  assign n21585 = ~n21582 & n21584;
  assign po322 = ~n21553 & ~n21585;
  assign n21587 = pi772 & pi947;
  assign n21588 = ~pi39 & ~n21587;
  assign n21589 = n21035 & n21588;
  assign n21590 = ~pi166 & ~n16508;
  assign n21591 = pi38 & ~n21590;
  assign n21592 = ~n21589 & n21591;
  assign n21593 = pi166 & ~n16201;
  assign n21594 = ~n16202 & ~n21588;
  assign n21595 = ~n21593 & ~n21594;
  assign n21596 = ~n20425 & n21595;
  assign n21597 = ~n6192 & n16269;
  assign n21598 = ~pi166 & ~n21597;
  assign n21599 = n20803 & ~n21598;
  assign n21600 = ~pi299 & ~n21599;
  assign n21601 = ~pi166 & ~n16269;
  assign n21602 = n20798 & ~n21601;
  assign n21603 = pi166 & ~n16207;
  assign n21604 = ~n20729 & ~n21603;
  assign n21605 = n2607 & n21604;
  assign n21606 = ~pi223 & ~n21605;
  assign n21607 = ~pi166 & n16329;
  assign n21608 = ~n20833 & ~n21607;
  assign n21609 = n20813 & ~n21608;
  assign n21610 = n21606 & ~n21609;
  assign n21611 = ~n21602 & ~n21610;
  assign n21612 = n21600 & n21611;
  assign n21613 = pi166 & n20432;
  assign n21614 = n20413 & ~n21613;
  assign n21615 = ~n16340 & n21614;
  assign n21616 = n2527 & n21604;
  assign n21617 = ~pi215 & ~n21616;
  assign n21618 = ~n21615 & n21617;
  assign n21619 = ~pi166 & ~n16346;
  assign n21620 = n20429 & ~n21619;
  assign n21621 = pi299 & ~n21620;
  assign n21622 = ~n21618 & n21621;
  assign n21623 = pi772 & ~n21622;
  assign n21624 = ~n21612 & n21623;
  assign n21625 = ~n20840 & n21620;
  assign n21626 = pi299 & ~n21625;
  assign n21627 = ~n20430 & n21617;
  assign n21628 = ~n21614 & n21627;
  assign n21629 = n21626 & ~n21628;
  assign n21630 = ~n2607 & ~n21608;
  assign n21631 = pi947 & n16271;
  assign n21632 = ~n21630 & ~n21631;
  assign n21633 = n21606 & n21632;
  assign n21634 = n21600 & ~n21633;
  assign n21635 = ~pi772 & ~n21634;
  assign n21636 = ~n21629 & n21635;
  assign n21637 = ~n21624 & ~n21636;
  assign n21638 = pi39 & n21637;
  assign n21639 = ~pi38 & ~n21638;
  assign n21640 = ~n21596 & n21639;
  assign n21641 = pi727 & ~n21640;
  assign n21642 = ~n21592 & n21641;
  assign n21643 = ~pi772 & ~n16355;
  assign n21644 = pi166 & n21643;
  assign n21645 = ~n20517 & ~n21603;
  assign n21646 = n2607 & ~n21645;
  assign n21647 = n20810 & ~n21607;
  assign n21648 = ~n21646 & ~n21647;
  assign n21649 = ~pi223 & ~n21648;
  assign n21650 = ~pi299 & ~n21649;
  assign n21651 = ~n21602 & n21650;
  assign n21652 = pi166 & n20496;
  assign n21653 = n2527 & n21645;
  assign n21654 = ~n21615 & ~n21653;
  assign n21655 = n20494 & n21654;
  assign n21656 = ~n21652 & ~n21655;
  assign n21657 = n20515 & n21656;
  assign n21658 = ~n21651 & ~n21657;
  assign n21659 = pi772 & n21658;
  assign n21660 = ~n21644 & ~n21659;
  assign n21661 = pi39 & n21660;
  assign n21662 = ~pi38 & ~n21661;
  assign n21663 = ~n21595 & n21662;
  assign n21664 = n2934 & ~n21587;
  assign n21665 = n6097 & n21664;
  assign n21666 = ~pi166 & ~n16524;
  assign n21667 = pi38 & ~n21666;
  assign n21668 = ~n21665 & n21667;
  assign n21669 = ~pi727 & ~n21668;
  assign n21670 = ~n21663 & n21669;
  assign n21671 = ~n21642 & ~n21670;
  assign n21672 = n10021 & ~n21671;
  assign n21673 = ~pi166 & ~n10021;
  assign n21674 = ~pi832 & ~n21673;
  assign n21675 = ~n21672 & n21674;
  assign n21676 = pi727 & n20323;
  assign n21677 = n21664 & ~n21676;
  assign n21678 = ~pi166 & ~n2934;
  assign n21679 = pi832 & ~n21678;
  assign n21680 = ~n21677 & n21679;
  assign po323 = n21675 | n21680;
  assign n21682 = ~pi768 & pi947;
  assign n21683 = pi705 & n20323;
  assign n21684 = ~n21682 & ~n21683;
  assign n21685 = n2934 & ~n21684;
  assign n21686 = ~pi167 & ~n2934;
  assign n21687 = pi832 & ~n21686;
  assign n21688 = ~n21685 & n21687;
  assign n21689 = ~pi167 & ~n16508;
  assign n21690 = n20453 & ~n21689;
  assign n21691 = ~pi167 & n20447;
  assign n21692 = pi167 & n20427;
  assign n21693 = ~pi38 & ~n21692;
  assign n21694 = ~n21691 & n21693;
  assign n21695 = pi768 & ~n21694;
  assign n21696 = ~n21690 & n21695;
  assign n21697 = ~pi167 & ~n20457;
  assign n21698 = n20460 & ~n21697;
  assign n21699 = pi167 & n20480;
  assign n21700 = ~pi167 & n20472;
  assign n21701 = ~pi38 & ~n21700;
  assign n21702 = ~n21699 & n21701;
  assign n21703 = ~pi768 & ~n21702;
  assign n21704 = ~n21698 & n21703;
  assign n21705 = pi705 & ~n21704;
  assign n21706 = ~n21696 & n21705;
  assign n21707 = pi768 & ~n16526;
  assign n21708 = ~pi167 & n21707;
  assign n21709 = pi167 & n20524;
  assign n21710 = ~pi167 & ~n20503;
  assign n21711 = ~pi38 & ~n21710;
  assign n21712 = ~n21709 & n21711;
  assign n21713 = ~pi167 & ~n16524;
  assign n21714 = ~n20510 & ~n21713;
  assign n21715 = ~pi768 & ~n21714;
  assign n21716 = ~n21712 & n21715;
  assign n21717 = ~pi705 & ~n21716;
  assign n21718 = ~n21708 & n21717;
  assign n21719 = ~n21706 & ~n21718;
  assign n21720 = n10021 & n21719;
  assign n21721 = ~pi167 & ~n10021;
  assign n21722 = ~pi832 & ~n21721;
  assign n21723 = ~n21720 & n21722;
  assign po324 = ~n21688 & ~n21723;
  assign n21725 = pi763 & pi947;
  assign n21726 = pi699 & n20323;
  assign n21727 = ~n21725 & ~n21726;
  assign n21728 = n2934 & n21727;
  assign n21729 = pi168 & ~n2934;
  assign n21730 = pi832 & ~n21729;
  assign n21731 = ~n21728 & n21730;
  assign n21732 = ~pi168 & ~n20537;
  assign n21733 = ~pi168 & ~n16201;
  assign n21734 = ~pi763 & n17520;
  assign n21735 = ~n20512 & ~n21734;
  assign n21736 = ~n21733 & ~n21735;
  assign n21737 = ~n20425 & n21736;
  assign n21738 = pi168 & ~n16346;
  assign n21739 = n20429 & ~n21738;
  assign n21740 = pi168 & n20724;
  assign n21741 = ~n16339 & ~n21740;
  assign n21742 = ~pi168 & ~n16207;
  assign n21743 = n20518 & ~n21742;
  assign n21744 = ~n20414 & n21743;
  assign n21745 = ~pi215 & ~n21744;
  assign n21746 = n21741 & n21745;
  assign n21747 = ~n21739 & ~n21746;
  assign n21748 = pi299 & ~n21747;
  assign n21749 = pi168 & ~n20735;
  assign n21750 = ~n20466 & ~n21749;
  assign n21751 = ~n21748 & ~n21750;
  assign n21752 = pi763 & ~n21751;
  assign n21753 = n20474 & ~n21739;
  assign n21754 = n20416 & ~n21742;
  assign n21755 = ~n20433 & ~n21754;
  assign n21756 = n21741 & n21755;
  assign n21757 = ~pi215 & ~n21756;
  assign n21758 = ~n21753 & ~n21757;
  assign n21759 = ~n20438 & n21758;
  assign n21760 = pi299 & ~n21759;
  assign n21761 = ~pi168 & ~n16333;
  assign n21762 = n20422 & ~n21761;
  assign n21763 = ~pi763 & ~n21762;
  assign n21764 = ~n21760 & n21763;
  assign n21765 = pi39 & ~n21764;
  assign n21766 = ~n21752 & n21765;
  assign n21767 = ~n21737 & ~n21766;
  assign n21768 = ~pi38 & ~n21767;
  assign n21769 = ~n20323 & ~n21725;
  assign n21770 = n16508 & ~n21769;
  assign n21771 = ~pi168 & ~n16508;
  assign n21772 = pi38 & ~n21771;
  assign n21773 = ~n21770 & n21772;
  assign n21774 = ~n21768 & ~n21773;
  assign n21775 = pi699 & ~n21774;
  assign n21776 = pi168 & ~n16524;
  assign n21777 = n16508 & ~n21725;
  assign n21778 = ~n21776 & ~n21777;
  assign n21779 = pi38 & n21778;
  assign n21780 = ~pi168 & ~pi763;
  assign n21781 = ~n16355 & n21780;
  assign n21782 = n20514 & ~n21761;
  assign n21783 = n20494 & ~n21743;
  assign n21784 = n21741 & n21783;
  assign n21785 = n20496 & ~n21738;
  assign n21786 = pi299 & ~n21785;
  assign n21787 = ~n21784 & n21786;
  assign n21788 = ~n21782 & ~n21787;
  assign n21789 = pi763 & n21788;
  assign n21790 = ~n21781 & ~n21789;
  assign n21791 = pi39 & n21790;
  assign n21792 = ~pi38 & ~n21736;
  assign n21793 = ~n21791 & n21792;
  assign n21794 = ~pi699 & ~n21793;
  assign n21795 = ~n21779 & n21794;
  assign n21796 = ~n21775 & ~n21795;
  assign n21797 = n20537 & n21796;
  assign n21798 = ~pi57 & ~n21797;
  assign n21799 = ~n21732 & n21798;
  assign n21800 = pi57 & pi168;
  assign n21801 = ~pi832 & ~n21800;
  assign n21802 = ~n21799 & n21801;
  assign po325 = n21731 | n21802;
  assign n21804 = pi746 & pi947;
  assign n21805 = pi729 & n20323;
  assign n21806 = ~n21804 & ~n21805;
  assign n21807 = n2934 & n21806;
  assign n21808 = pi169 & ~n2934;
  assign n21809 = pi832 & ~n21808;
  assign n21810 = ~n21807 & n21809;
  assign n21811 = ~pi169 & ~n20537;
  assign n21812 = ~pi169 & ~n16201;
  assign n21813 = ~pi746 & n17520;
  assign n21814 = ~n20512 & ~n21813;
  assign n21815 = ~n21812 & ~n21814;
  assign n21816 = ~n20425 & n21815;
  assign n21817 = pi169 & ~n16346;
  assign n21818 = n20429 & ~n21817;
  assign n21819 = pi169 & n20724;
  assign n21820 = ~n16339 & ~n21819;
  assign n21821 = ~pi169 & ~n16207;
  assign n21822 = n20518 & ~n21821;
  assign n21823 = ~n20414 & n21822;
  assign n21824 = ~pi215 & ~n21823;
  assign n21825 = n21820 & n21824;
  assign n21826 = ~n21818 & ~n21825;
  assign n21827 = pi299 & ~n21826;
  assign n21828 = pi169 & ~n20735;
  assign n21829 = ~n20466 & ~n21828;
  assign n21830 = ~n21827 & ~n21829;
  assign n21831 = pi746 & ~n21830;
  assign n21832 = n20474 & ~n21818;
  assign n21833 = n20416 & ~n21821;
  assign n21834 = ~n20433 & ~n21833;
  assign n21835 = n21820 & n21834;
  assign n21836 = ~pi215 & ~n21835;
  assign n21837 = ~n21832 & ~n21836;
  assign n21838 = ~n20438 & n21837;
  assign n21839 = pi299 & ~n21838;
  assign n21840 = ~pi169 & ~n16333;
  assign n21841 = n20422 & ~n21840;
  assign n21842 = ~pi746 & ~n21841;
  assign n21843 = ~n21839 & n21842;
  assign n21844 = pi39 & ~n21843;
  assign n21845 = ~n21831 & n21844;
  assign n21846 = ~n21816 & ~n21845;
  assign n21847 = ~pi38 & ~n21846;
  assign n21848 = ~n20323 & ~n21804;
  assign n21849 = n16508 & ~n21848;
  assign n21850 = ~pi169 & ~n16508;
  assign n21851 = pi38 & ~n21850;
  assign n21852 = ~n21849 & n21851;
  assign n21853 = ~n21847 & ~n21852;
  assign n21854 = pi729 & ~n21853;
  assign n21855 = pi169 & ~n16524;
  assign n21856 = n16508 & ~n21804;
  assign n21857 = ~n21855 & ~n21856;
  assign n21858 = pi38 & n21857;
  assign n21859 = ~pi169 & ~pi746;
  assign n21860 = ~n16355 & n21859;
  assign n21861 = n20514 & ~n21840;
  assign n21862 = n20494 & ~n21822;
  assign n21863 = n21820 & n21862;
  assign n21864 = n20496 & ~n21817;
  assign n21865 = pi299 & ~n21864;
  assign n21866 = ~n21863 & n21865;
  assign n21867 = ~n21861 & ~n21866;
  assign n21868 = pi746 & n21867;
  assign n21869 = ~n21860 & ~n21868;
  assign n21870 = pi39 & n21869;
  assign n21871 = ~pi38 & ~n21815;
  assign n21872 = ~n21870 & n21871;
  assign n21873 = ~pi729 & ~n21872;
  assign n21874 = ~n21858 & n21873;
  assign n21875 = ~n21854 & ~n21874;
  assign n21876 = n20537 & n21875;
  assign n21877 = ~pi57 & ~n21876;
  assign n21878 = ~n21811 & n21877;
  assign n21879 = pi57 & pi169;
  assign n21880 = ~pi832 & ~n21879;
  assign n21881 = ~n21878 & n21880;
  assign po326 = n21810 | n21881;
  assign n21883 = pi748 & pi947;
  assign n21884 = pi730 & n20323;
  assign n21885 = ~n21883 & ~n21884;
  assign n21886 = n2934 & n21885;
  assign n21887 = pi170 & ~n2934;
  assign n21888 = pi832 & ~n21887;
  assign n21889 = ~n21886 & n21888;
  assign n21890 = ~pi170 & ~n20537;
  assign n21891 = ~pi170 & ~n16508;
  assign n21892 = n20460 & ~n21891;
  assign n21893 = ~pi170 & ~n16201;
  assign n21894 = n20470 & ~n21893;
  assign n21895 = pi170 & ~n20735;
  assign n21896 = ~n20466 & ~n21895;
  assign n21897 = pi170 & ~n16346;
  assign n21898 = n20429 & ~n21897;
  assign n21899 = pi170 & n20724;
  assign n21900 = ~n16339 & ~n21899;
  assign n21901 = ~pi170 & ~n16207;
  assign n21902 = n20518 & ~n21901;
  assign n21903 = ~n20414 & n21902;
  assign n21904 = ~pi215 & ~n21903;
  assign n21905 = n21900 & n21904;
  assign n21906 = ~n21898 & ~n21905;
  assign n21907 = pi299 & ~n21906;
  assign n21908 = pi39 & ~n21907;
  assign n21909 = ~n21896 & n21908;
  assign n21910 = ~n21894 & ~n21909;
  assign n21911 = ~pi38 & ~n21910;
  assign n21912 = pi748 & ~n21911;
  assign n21913 = ~n21892 & n21912;
  assign n21914 = n20453 & ~n21891;
  assign n21915 = n20474 & ~n21898;
  assign n21916 = n20416 & ~n21901;
  assign n21917 = ~n20433 & ~n21916;
  assign n21918 = n21900 & n21917;
  assign n21919 = ~pi215 & ~n21918;
  assign n21920 = ~n21915 & ~n21919;
  assign n21921 = ~n20438 & n21920;
  assign n21922 = pi299 & ~n21921;
  assign n21923 = ~pi170 & ~n16333;
  assign n21924 = ~pi299 & ~n21923;
  assign n21925 = ~n20421 & n21924;
  assign n21926 = ~n21922 & ~n21925;
  assign n21927 = pi39 & ~n21926;
  assign n21928 = n20426 & ~n21893;
  assign n21929 = ~n21927 & ~n21928;
  assign n21930 = ~pi38 & ~n21929;
  assign n21931 = ~pi748 & ~n21930;
  assign n21932 = ~n21914 & n21931;
  assign n21933 = pi730 & ~n21932;
  assign n21934 = ~n21913 & n21933;
  assign n21935 = ~pi170 & ~pi748;
  assign n21936 = ~n16526 & n21935;
  assign n21937 = n20512 & ~n21893;
  assign n21938 = ~n20410 & n21898;
  assign n21939 = pi299 & ~n21938;
  assign n21940 = n20494 & ~n21902;
  assign n21941 = n21900 & n21940;
  assign n21942 = n21939 & ~n21941;
  assign n21943 = ~n20513 & n21924;
  assign n21944 = ~n21942 & ~n21943;
  assign n21945 = pi39 & ~n21944;
  assign n21946 = ~n21937 & ~n21945;
  assign n21947 = ~pi38 & ~n21946;
  assign n21948 = ~pi170 & ~n16524;
  assign n21949 = ~n20510 & ~n21948;
  assign n21950 = pi748 & ~n21949;
  assign n21951 = ~n21947 & n21950;
  assign n21952 = ~pi730 & ~n21951;
  assign n21953 = ~n21936 & n21952;
  assign n21954 = ~n21934 & ~n21953;
  assign n21955 = n20537 & n21954;
  assign n21956 = ~pi57 & ~n21955;
  assign n21957 = ~n21890 & n21956;
  assign n21958 = pi57 & pi170;
  assign n21959 = ~pi832 & ~n21958;
  assign n21960 = ~n21957 & n21959;
  assign po327 = n21889 | n21960;
  assign n21962 = pi764 & pi947;
  assign n21963 = pi691 & n20323;
  assign n21964 = ~n21962 & ~n21963;
  assign n21965 = n2934 & n21964;
  assign n21966 = pi171 & ~n2934;
  assign n21967 = pi832 & ~n21966;
  assign n21968 = ~n21965 & n21967;
  assign n21969 = ~pi171 & ~n20537;
  assign n21970 = ~pi171 & ~n16201;
  assign n21971 = ~pi764 & n17520;
  assign n21972 = ~n20512 & ~n21971;
  assign n21973 = ~n21970 & ~n21972;
  assign n21974 = ~n20425 & n21973;
  assign n21975 = pi171 & ~n16346;
  assign n21976 = n20429 & ~n21975;
  assign n21977 = pi171 & n20724;
  assign n21978 = ~n16339 & ~n21977;
  assign n21979 = ~pi171 & ~n16207;
  assign n21980 = n20518 & ~n21979;
  assign n21981 = ~n20414 & n21980;
  assign n21982 = ~pi215 & ~n21981;
  assign n21983 = n21978 & n21982;
  assign n21984 = ~n21976 & ~n21983;
  assign n21985 = pi299 & ~n21984;
  assign n21986 = pi171 & ~n20735;
  assign n21987 = ~n20466 & ~n21986;
  assign n21988 = ~n21985 & ~n21987;
  assign n21989 = pi764 & ~n21988;
  assign n21990 = n20474 & ~n21976;
  assign n21991 = n20416 & ~n21979;
  assign n21992 = ~n20433 & ~n21991;
  assign n21993 = n21978 & n21992;
  assign n21994 = ~pi215 & ~n21993;
  assign n21995 = ~n21990 & ~n21994;
  assign n21996 = ~n20438 & n21995;
  assign n21997 = pi299 & ~n21996;
  assign n21998 = ~pi171 & ~n16333;
  assign n21999 = n20422 & ~n21998;
  assign n22000 = ~pi764 & ~n21999;
  assign n22001 = ~n21997 & n22000;
  assign n22002 = pi39 & ~n22001;
  assign n22003 = ~n21989 & n22002;
  assign n22004 = ~n21974 & ~n22003;
  assign n22005 = ~pi38 & ~n22004;
  assign n22006 = ~n20323 & ~n21962;
  assign n22007 = n16508 & ~n22006;
  assign n22008 = ~pi171 & ~n16508;
  assign n22009 = pi38 & ~n22008;
  assign n22010 = ~n22007 & n22009;
  assign n22011 = ~n22005 & ~n22010;
  assign n22012 = pi691 & ~n22011;
  assign n22013 = pi171 & ~n16524;
  assign n22014 = n16508 & ~n21962;
  assign n22015 = ~n22013 & ~n22014;
  assign n22016 = pi38 & n22015;
  assign n22017 = ~pi171 & ~pi764;
  assign n22018 = ~n16355 & n22017;
  assign n22019 = n20514 & ~n21998;
  assign n22020 = n20494 & ~n21980;
  assign n22021 = n21978 & n22020;
  assign n22022 = n20496 & ~n21975;
  assign n22023 = pi299 & ~n22022;
  assign n22024 = ~n22021 & n22023;
  assign n22025 = ~n22019 & ~n22024;
  assign n22026 = pi764 & n22025;
  assign n22027 = ~n22018 & ~n22026;
  assign n22028 = pi39 & n22027;
  assign n22029 = ~pi38 & ~n21973;
  assign n22030 = ~n22028 & n22029;
  assign n22031 = ~pi691 & ~n22030;
  assign n22032 = ~n22016 & n22031;
  assign n22033 = ~n22012 & ~n22032;
  assign n22034 = n20537 & n22033;
  assign n22035 = ~pi57 & ~n22034;
  assign n22036 = ~n21969 & n22035;
  assign n22037 = pi57 & pi171;
  assign n22038 = ~pi832 & ~n22037;
  assign n22039 = ~n22036 & n22038;
  assign po328 = n21968 | n22039;
  assign n22041 = pi739 & pi947;
  assign n22042 = pi690 & n20323;
  assign n22043 = ~n22041 & ~n22042;
  assign n22044 = n2934 & n22043;
  assign n22045 = pi172 & ~n2934;
  assign n22046 = pi832 & ~n22045;
  assign n22047 = ~n22044 & n22046;
  assign n22048 = ~pi172 & ~n20537;
  assign n22049 = ~pi172 & ~n16201;
  assign n22050 = ~pi39 & ~n22049;
  assign n22051 = n16201 & n22041;
  assign n22052 = n22050 & ~n22051;
  assign n22053 = ~n20425 & n22052;
  assign n22054 = pi172 & ~n16346;
  assign n22055 = n20429 & ~n22054;
  assign n22056 = pi172 & n20724;
  assign n22057 = ~n16339 & ~n22056;
  assign n22058 = ~pi172 & ~n16207;
  assign n22059 = n20518 & ~n22058;
  assign n22060 = ~n20414 & n22059;
  assign n22061 = ~pi215 & ~n22060;
  assign n22062 = n22057 & n22061;
  assign n22063 = ~n22055 & ~n22062;
  assign n22064 = pi299 & ~n22063;
  assign n22065 = pi172 & ~n20735;
  assign n22066 = ~n20466 & ~n22065;
  assign n22067 = ~n22064 & ~n22066;
  assign n22068 = pi739 & ~n22067;
  assign n22069 = n20474 & ~n22055;
  assign n22070 = n20416 & ~n22058;
  assign n22071 = ~n20433 & ~n22070;
  assign n22072 = n22057 & n22071;
  assign n22073 = ~pi215 & ~n22072;
  assign n22074 = ~n22069 & ~n22073;
  assign n22075 = ~n20438 & n22074;
  assign n22076 = pi299 & ~n22075;
  assign n22077 = ~pi172 & ~n16333;
  assign n22078 = n20422 & ~n22077;
  assign n22079 = ~pi739 & ~n22078;
  assign n22080 = ~n22076 & n22079;
  assign n22081 = pi39 & ~n22080;
  assign n22082 = ~n22068 & n22081;
  assign n22083 = ~n22053 & ~n22082;
  assign n22084 = ~pi38 & ~n22083;
  assign n22085 = ~n20323 & ~n22041;
  assign n22086 = n16508 & ~n22085;
  assign n22087 = ~pi172 & ~n16508;
  assign n22088 = pi38 & ~n22087;
  assign n22089 = ~n22086 & n22088;
  assign n22090 = ~n22084 & ~n22089;
  assign n22091 = pi690 & ~n22090;
  assign n22092 = pi172 & ~n16524;
  assign n22093 = n16508 & ~n22041;
  assign n22094 = ~n22092 & ~n22093;
  assign n22095 = pi38 & n22094;
  assign n22096 = ~pi172 & ~pi739;
  assign n22097 = ~n16355 & n22096;
  assign n22098 = n20514 & ~n22077;
  assign n22099 = n20494 & ~n22059;
  assign n22100 = n22057 & n22099;
  assign n22101 = n20496 & ~n22054;
  assign n22102 = pi299 & ~n22101;
  assign n22103 = ~n22100 & n22102;
  assign n22104 = ~n22098 & ~n22103;
  assign n22105 = pi739 & n22104;
  assign n22106 = ~n22097 & ~n22105;
  assign n22107 = pi39 & n22106;
  assign n22108 = ~pi38 & ~n22052;
  assign n22109 = ~n22107 & n22108;
  assign n22110 = ~pi690 & ~n22109;
  assign n22111 = ~n22095 & n22110;
  assign n22112 = ~n22091 & ~n22111;
  assign n22113 = n20537 & n22112;
  assign n22114 = ~pi57 & ~n22113;
  assign n22115 = ~n22048 & n22114;
  assign n22116 = pi57 & pi172;
  assign n22117 = ~pi832 & ~n22116;
  assign n22118 = ~n22115 & n22117;
  assign po329 = n22047 | n22118;
  assign n22120 = ~pi173 & ~n16527;
  assign n22121 = n17159 & ~n22120;
  assign n22122 = n16593 & ~n22120;
  assign n22123 = ~pi723 & n10020;
  assign n22124 = n22120 & ~n22123;
  assign n22125 = ~pi173 & n17592;
  assign n22126 = ~pi38 & ~pi173;
  assign n22127 = n19843 & ~n22126;
  assign n22128 = ~n22125 & ~n22127;
  assign n22129 = ~pi173 & ~n16508;
  assign n22130 = n16744 & ~n22129;
  assign n22131 = ~pi723 & ~n22130;
  assign n22132 = ~n22128 & n22131;
  assign n22133 = ~n22124 & ~n22132;
  assign n22134 = ~pi778 & n22133;
  assign n22135 = pi625 & ~n22133;
  assign n22136 = pi1153 & ~n22135;
  assign n22137 = ~pi625 & n22120;
  assign n22138 = n22136 & ~n22137;
  assign n22139 = ~pi625 & ~n22133;
  assign n22140 = ~pi1153 & ~n22139;
  assign n22141 = pi625 & n22120;
  assign n22142 = n22140 & ~n22141;
  assign n22143 = ~n22138 & ~n22142;
  assign n22144 = pi778 & ~n22143;
  assign n22145 = ~n22134 & ~n22144;
  assign n22146 = ~n16593 & ~n22145;
  assign n22147 = ~n22122 & ~n22146;
  assign n22148 = ~n16589 & n22147;
  assign n22149 = n16589 & n22120;
  assign n22150 = ~n22148 & ~n22149;
  assign n22151 = ~n17159 & n22150;
  assign n22152 = ~n22121 & ~n22151;
  assign n22153 = ~n17183 & n22152;
  assign n22154 = n17183 & n22120;
  assign n22155 = ~n22153 & ~n22154;
  assign n22156 = ~pi792 & n22155;
  assign n22157 = pi628 & ~n22155;
  assign n22158 = pi1156 & ~n22157;
  assign n22159 = ~pi628 & n22120;
  assign n22160 = n22158 & ~n22159;
  assign n22161 = ~pi628 & ~n22155;
  assign n22162 = pi628 & n22120;
  assign n22163 = ~pi1156 & ~n22162;
  assign n22164 = ~n22161 & n22163;
  assign n22165 = ~n22160 & ~n22164;
  assign n22166 = pi792 & ~n22165;
  assign n22167 = ~n22156 & ~n22166;
  assign n22168 = pi647 & ~n22167;
  assign n22169 = ~pi647 & ~n22120;
  assign n22170 = ~n22168 & ~n22169;
  assign n22171 = pi1157 & ~n22170;
  assign n22172 = ~pi647 & n22167;
  assign n22173 = ~pi1157 & ~n22172;
  assign n22174 = pi647 & n22120;
  assign n22175 = n22173 & ~n22174;
  assign n22176 = ~n22171 & ~n22175;
  assign n22177 = pi787 & ~n22176;
  assign n22178 = ~pi787 & ~n22167;
  assign n22179 = ~n22177 & ~n22178;
  assign n22180 = ~pi644 & n22179;
  assign n22181 = pi715 & ~n22180;
  assign n22182 = n17247 & ~n22120;
  assign n22183 = pi173 & ~n10020;
  assign n22184 = ~pi745 & n16511;
  assign n22185 = ~n22129 & ~n22184;
  assign n22186 = pi38 & ~n22185;
  assign n22187 = n10020 & ~n22186;
  assign n22188 = ~pi173 & ~pi745;
  assign n22189 = n16449 & n22188;
  assign n22190 = pi173 & ~n16503;
  assign n22191 = ~pi173 & ~n16357;
  assign n22192 = pi745 & ~n22191;
  assign n22193 = ~n22190 & ~n22192;
  assign n22194 = ~n22189 & n22193;
  assign n22195 = ~pi38 & n22194;
  assign n22196 = n22187 & ~n22195;
  assign n22197 = ~n22183 & ~n22196;
  assign n22198 = ~n16521 & ~n22197;
  assign n22199 = n16521 & ~n22120;
  assign n22200 = ~n22198 & ~n22199;
  assign n22201 = ~pi785 & ~n22200;
  assign n22202 = ~n16532 & ~n22120;
  assign n22203 = pi609 & n22198;
  assign n22204 = ~n22202 & ~n22203;
  assign n22205 = pi1155 & ~n22204;
  assign n22206 = ~n16537 & ~n22120;
  assign n22207 = ~pi609 & n22198;
  assign n22208 = ~n22206 & ~n22207;
  assign n22209 = ~pi1155 & ~n22208;
  assign n22210 = ~n22205 & ~n22209;
  assign n22211 = pi785 & ~n22210;
  assign n22212 = ~n22201 & ~n22211;
  assign n22213 = ~pi781 & ~n22212;
  assign n22214 = pi618 & n22212;
  assign n22215 = ~pi618 & n22120;
  assign n22216 = pi1154 & ~n22215;
  assign n22217 = ~n22214 & n22216;
  assign n22218 = ~pi618 & n22212;
  assign n22219 = pi618 & n22120;
  assign n22220 = ~pi1154 & ~n22219;
  assign n22221 = ~n22218 & n22220;
  assign n22222 = ~n22217 & ~n22221;
  assign n22223 = pi781 & ~n22222;
  assign n22224 = ~n22213 & ~n22223;
  assign n22225 = ~pi789 & ~n22224;
  assign n22226 = pi619 & n22224;
  assign n22227 = ~pi619 & n22120;
  assign n22228 = pi1159 & ~n22227;
  assign n22229 = ~n22226 & n22228;
  assign n22230 = ~pi619 & n22224;
  assign n22231 = pi619 & n22120;
  assign n22232 = ~pi1159 & ~n22231;
  assign n22233 = ~n22230 & n22232;
  assign n22234 = ~n22229 & ~n22233;
  assign n22235 = pi789 & ~n22234;
  assign n22236 = ~n22225 & ~n22235;
  assign n22237 = ~pi788 & ~n22236;
  assign n22238 = pi626 & n22236;
  assign n22239 = ~pi626 & n22120;
  assign n22240 = pi1158 & ~n22239;
  assign n22241 = ~n22238 & n22240;
  assign n22242 = ~pi626 & n22236;
  assign n22243 = pi626 & n22120;
  assign n22244 = ~pi1158 & ~n22243;
  assign n22245 = ~n22242 & n22244;
  assign n22246 = ~n22241 & ~n22245;
  assign n22247 = pi788 & ~n22246;
  assign n22248 = ~n22237 & ~n22247;
  assign n22249 = ~n16124 & n22248;
  assign n22250 = n16124 & n22120;
  assign n22251 = ~n22249 & ~n22250;
  assign n22252 = ~n17247 & n22251;
  assign n22253 = ~n22182 & ~n22252;
  assign n22254 = pi644 & n22253;
  assign n22255 = ~pi644 & n22120;
  assign n22256 = ~pi715 & ~n22255;
  assign n22257 = ~n22254 & n22256;
  assign n22258 = pi1160 & ~n22257;
  assign n22259 = ~n22181 & n22258;
  assign n22260 = ~pi644 & n22253;
  assign n22261 = pi715 & ~n22260;
  assign n22262 = pi644 & n22120;
  assign n22263 = n22261 & ~n22262;
  assign n22264 = pi644 & n22179;
  assign n22265 = ~n19987 & n22251;
  assign n22266 = pi630 & n22175;
  assign n22267 = ~n22265 & ~n22266;
  assign n22268 = n17244 & ~n22170;
  assign n22269 = n22267 & ~n22268;
  assign n22270 = pi787 & ~n22269;
  assign n22271 = ~pi629 & n22160;
  assign n22272 = ~n19999 & ~n22248;
  assign n22273 = pi629 & n22164;
  assign n22274 = ~n22272 & ~n22273;
  assign n22275 = ~n22271 & n22274;
  assign n22276 = pi792 & ~n22275;
  assign n22277 = pi618 & n22147;
  assign n22278 = pi609 & n22145;
  assign n22279 = pi625 & n22197;
  assign n22280 = ~n22123 & ~n22196;
  assign n22281 = ~pi745 & ~n16917;
  assign n22282 = n18933 & ~n22281;
  assign n22283 = ~pi173 & ~n22282;
  assign n22284 = ~pi745 & n16510;
  assign n22285 = ~n17079 & ~n22284;
  assign n22286 = pi173 & ~n22285;
  assign n22287 = n6097 & n22286;
  assign n22288 = ~n22283 & ~n22287;
  assign n22289 = pi38 & n22288;
  assign n22290 = ~pi173 & n16853;
  assign n22291 = pi173 & n16935;
  assign n22292 = pi745 & ~n22291;
  assign n22293 = ~n22290 & n22292;
  assign n22294 = pi173 & n16998;
  assign n22295 = ~pi173 & ~n17051;
  assign n22296 = ~pi745 & ~n22295;
  assign n22297 = ~n22294 & n22296;
  assign n22298 = ~n22293 & ~n22297;
  assign n22299 = pi39 & n22298;
  assign n22300 = ~pi173 & ~n17061;
  assign n22301 = pi173 & ~n17058;
  assign n22302 = pi745 & ~n22301;
  assign n22303 = ~n22300 & n22302;
  assign n22304 = ~pi173 & n17067;
  assign n22305 = pi173 & n17065;
  assign n22306 = ~pi745 & ~n22305;
  assign n22307 = ~n22304 & n22306;
  assign n22308 = ~n22303 & ~n22307;
  assign n22309 = ~pi39 & ~n22308;
  assign n22310 = ~pi38 & ~n22309;
  assign n22311 = ~n22299 & n22310;
  assign n22312 = ~pi723 & ~n22311;
  assign n22313 = ~n22289 & n22312;
  assign n22314 = ~n22280 & ~n22313;
  assign n22315 = ~n22183 & ~n22314;
  assign n22316 = ~pi625 & n22315;
  assign n22317 = ~pi1153 & ~n22316;
  assign n22318 = ~n22279 & n22317;
  assign n22319 = ~pi608 & ~n22138;
  assign n22320 = ~n22318 & n22319;
  assign n22321 = ~pi625 & n22197;
  assign n22322 = pi625 & n22315;
  assign n22323 = ~n22321 & ~n22322;
  assign n22324 = pi1153 & n22323;
  assign n22325 = ~n22142 & ~n22324;
  assign n22326 = pi608 & n22325;
  assign n22327 = ~n22320 & ~n22326;
  assign n22328 = pi778 & ~n22327;
  assign n22329 = ~pi778 & n22315;
  assign n22330 = ~n22328 & ~n22329;
  assign n22331 = ~pi609 & ~n22330;
  assign n22332 = ~pi1155 & ~n22331;
  assign n22333 = ~n22278 & n22332;
  assign n22334 = ~pi660 & ~n22205;
  assign n22335 = ~n22333 & n22334;
  assign n22336 = ~pi609 & n22145;
  assign n22337 = pi609 & ~n22330;
  assign n22338 = ~n22336 & ~n22337;
  assign n22339 = pi1155 & n22338;
  assign n22340 = ~n22209 & ~n22339;
  assign n22341 = pi660 & n22340;
  assign n22342 = ~n22335 & ~n22341;
  assign n22343 = pi785 & ~n22342;
  assign n22344 = ~pi785 & ~n22330;
  assign n22345 = ~n22343 & ~n22344;
  assign n22346 = ~pi618 & ~n22345;
  assign n22347 = ~pi1154 & ~n22346;
  assign n22348 = ~n22277 & n22347;
  assign n22349 = ~pi627 & ~n22217;
  assign n22350 = ~n22348 & n22349;
  assign n22351 = ~pi618 & n22147;
  assign n22352 = pi618 & ~n22345;
  assign n22353 = ~n22351 & ~n22352;
  assign n22354 = pi1154 & n22353;
  assign n22355 = ~n22221 & ~n22354;
  assign n22356 = pi627 & n22355;
  assign n22357 = ~n22350 & ~n22356;
  assign n22358 = pi781 & ~n22357;
  assign n22359 = ~pi781 & ~n22345;
  assign n22360 = ~n22358 & ~n22359;
  assign n22361 = ~pi789 & n22360;
  assign n22362 = ~pi619 & ~n22360;
  assign n22363 = pi619 & ~n22150;
  assign n22364 = ~pi1159 & ~n22363;
  assign n22365 = ~n22362 & n22364;
  assign n22366 = ~pi648 & ~n22365;
  assign n22367 = ~n22229 & n22366;
  assign n22368 = ~pi619 & ~n22150;
  assign n22369 = pi619 & ~n22360;
  assign n22370 = ~n22368 & ~n22369;
  assign n22371 = pi1159 & n22370;
  assign n22372 = ~n22233 & ~n22371;
  assign n22373 = pi648 & n22372;
  assign n22374 = ~n22367 & ~n22373;
  assign n22375 = pi789 & n22374;
  assign n22376 = ~n22361 & ~n22375;
  assign n22377 = n17356 & n22376;
  assign n22378 = n17350 & n22152;
  assign n22379 = ~n17182 & n22246;
  assign n22380 = ~n22378 & ~n22379;
  assign n22381 = pi788 & ~n22380;
  assign n22382 = n19788 & ~n22381;
  assign n22383 = ~n22377 & n22382;
  assign n22384 = ~n22276 & ~n22383;
  assign n22385 = n19637 & ~n22384;
  assign n22386 = ~n22270 & ~n22385;
  assign n22387 = ~pi644 & n22386;
  assign n22388 = ~pi715 & ~n22387;
  assign n22389 = ~n22264 & n22388;
  assign n22390 = ~pi1160 & ~n22389;
  assign n22391 = ~n22263 & n22390;
  assign n22392 = ~n22259 & ~n22391;
  assign n22393 = pi790 & ~n22392;
  assign n22394 = pi644 & n22258;
  assign n22395 = pi790 & ~n22394;
  assign n22396 = n22386 & ~n22395;
  assign n22397 = ~n22393 & ~n22396;
  assign n22398 = ~po1038 & ~n22397;
  assign n22399 = ~pi173 & po1038;
  assign n22400 = ~pi832 & ~n22399;
  assign n22401 = ~n22398 & n22400;
  assign n22402 = ~pi173 & ~n2934;
  assign n22403 = ~n22284 & ~n22402;
  assign n22404 = ~n17273 & ~n22403;
  assign n22405 = ~pi785 & ~n22404;
  assign n22406 = n16537 & n22284;
  assign n22407 = n22404 & ~n22406;
  assign n22408 = pi1155 & ~n22407;
  assign n22409 = ~pi1155 & ~n22402;
  assign n22410 = ~n22406 & n22409;
  assign n22411 = ~n22408 & ~n22410;
  assign n22412 = pi785 & ~n22411;
  assign n22413 = ~n22405 & ~n22412;
  assign n22414 = ~pi781 & ~n22413;
  assign n22415 = ~n17289 & n22413;
  assign n22416 = pi1154 & ~n22415;
  assign n22417 = ~n17292 & n22413;
  assign n22418 = ~pi1154 & ~n22417;
  assign n22419 = ~n22416 & ~n22418;
  assign n22420 = pi781 & ~n22419;
  assign n22421 = ~n22414 & ~n22420;
  assign n22422 = ~pi789 & ~n22421;
  assign n22423 = ~pi619 & n2934;
  assign n22424 = n22421 & ~n22423;
  assign n22425 = pi1159 & ~n22424;
  assign n22426 = pi619 & n2934;
  assign n22427 = n22421 & ~n22426;
  assign n22428 = ~pi1159 & ~n22427;
  assign n22429 = ~n22425 & ~n22428;
  assign n22430 = pi789 & ~n22429;
  assign n22431 = ~n22422 & ~n22430;
  assign n22432 = ~pi788 & ~n22431;
  assign n22433 = pi626 & n22431;
  assign n22434 = ~pi626 & n22402;
  assign n22435 = pi1158 & ~n22434;
  assign n22436 = ~n22433 & n22435;
  assign n22437 = ~pi626 & n22431;
  assign n22438 = pi626 & n22402;
  assign n22439 = ~pi1158 & ~n22438;
  assign n22440 = ~n22437 & n22439;
  assign n22441 = ~n22436 & ~n22440;
  assign n22442 = pi788 & ~n22441;
  assign n22443 = ~n22432 & ~n22442;
  assign n22444 = ~n16124 & n22443;
  assign n22445 = n16124 & n22402;
  assign n22446 = ~n22444 & ~n22445;
  assign n22447 = ~n19987 & n22446;
  assign n22448 = ~pi723 & n16742;
  assign n22449 = ~n22402 & ~n22448;
  assign n22450 = ~pi778 & ~n22449;
  assign n22451 = ~pi625 & n22448;
  assign n22452 = ~n22449 & ~n22451;
  assign n22453 = pi1153 & ~n22452;
  assign n22454 = ~pi1153 & ~n22402;
  assign n22455 = ~n22451 & n22454;
  assign n22456 = ~n22453 & ~n22455;
  assign n22457 = pi778 & n22456;
  assign n22458 = ~n22450 & ~n22457;
  assign n22459 = ~n17338 & ~n22458;
  assign n22460 = ~n17340 & n22459;
  assign n22461 = ~n17342 & n22460;
  assign n22462 = ~n17425 & n22461;
  assign n22463 = ~n17452 & n22462;
  assign n22464 = ~pi647 & n22463;
  assign n22465 = pi647 & n22402;
  assign n22466 = ~pi1157 & ~n22465;
  assign n22467 = ~n22464 & n22466;
  assign n22468 = ~pi647 & n22402;
  assign n22469 = pi647 & n22463;
  assign n22470 = pi1157 & ~n22469;
  assign n22471 = ~n22468 & n22470;
  assign n22472 = ~n22467 & ~n22471;
  assign n22473 = ~n17246 & ~n22472;
  assign n22474 = ~n22447 & ~n22473;
  assign n22475 = pi787 & ~n22474;
  assign n22476 = n17350 & n22461;
  assign n22477 = ~n17182 & n22441;
  assign n22478 = ~n22476 & ~n22477;
  assign n22479 = pi788 & ~n22478;
  assign n22480 = pi618 & n22459;
  assign n22481 = pi609 & ~n22458;
  assign n22482 = ~n16393 & ~n22449;
  assign n22483 = pi625 & n22482;
  assign n22484 = n22403 & ~n22482;
  assign n22485 = ~n22483 & ~n22484;
  assign n22486 = n22454 & ~n22485;
  assign n22487 = ~pi608 & ~n22453;
  assign n22488 = ~n22486 & n22487;
  assign n22489 = pi1153 & ~n22483;
  assign n22490 = n22403 & n22489;
  assign n22491 = ~n22455 & ~n22490;
  assign n22492 = pi608 & n22491;
  assign n22493 = ~n22488 & ~n22492;
  assign n22494 = pi778 & ~n22493;
  assign n22495 = ~pi778 & ~n22484;
  assign n22496 = ~n22494 & ~n22495;
  assign n22497 = ~pi609 & ~n22496;
  assign n22498 = ~pi1155 & ~n22497;
  assign n22499 = ~n22481 & n22498;
  assign n22500 = ~pi660 & ~n22408;
  assign n22501 = ~n22499 & n22500;
  assign n22502 = ~pi609 & ~n22458;
  assign n22503 = pi609 & ~n22496;
  assign n22504 = ~n22502 & ~n22503;
  assign n22505 = pi1155 & n22504;
  assign n22506 = ~n22410 & ~n22505;
  assign n22507 = pi660 & n22506;
  assign n22508 = ~n22501 & ~n22507;
  assign n22509 = pi785 & ~n22508;
  assign n22510 = ~pi785 & ~n22496;
  assign n22511 = ~n22509 & ~n22510;
  assign n22512 = ~pi618 & ~n22511;
  assign n22513 = ~pi1154 & ~n22512;
  assign n22514 = ~n22480 & n22513;
  assign n22515 = ~pi627 & ~n22416;
  assign n22516 = ~n22514 & n22515;
  assign n22517 = ~pi618 & n22459;
  assign n22518 = pi618 & ~n22511;
  assign n22519 = ~n22517 & ~n22518;
  assign n22520 = pi1154 & n22519;
  assign n22521 = ~n22418 & ~n22520;
  assign n22522 = pi627 & n22521;
  assign n22523 = ~n22516 & ~n22522;
  assign n22524 = pi781 & ~n22523;
  assign n22525 = ~pi781 & ~n22511;
  assign n22526 = ~n22524 & ~n22525;
  assign n22527 = ~pi619 & ~n22526;
  assign n22528 = pi619 & n22460;
  assign n22529 = ~pi1159 & ~n22528;
  assign n22530 = ~n22527 & n22529;
  assign n22531 = ~pi648 & ~n22530;
  assign n22532 = ~n22425 & n22531;
  assign n22533 = ~pi619 & n22460;
  assign n22534 = pi619 & ~n22526;
  assign n22535 = ~n22533 & ~n22534;
  assign n22536 = pi1159 & n22535;
  assign n22537 = ~n22428 & ~n22536;
  assign n22538 = pi648 & n22537;
  assign n22539 = ~n22532 & ~n22538;
  assign n22540 = pi789 & n22539;
  assign n22541 = ~pi789 & n22526;
  assign n22542 = n17356 & ~n22541;
  assign n22543 = ~n22540 & n22542;
  assign n22544 = ~n22479 & ~n22543;
  assign n22545 = n19788 & ~n22544;
  assign n22546 = n20275 & n22462;
  assign n22547 = n17449 & n22443;
  assign n22548 = ~pi629 & ~n22547;
  assign n22549 = ~n22546 & n22548;
  assign n22550 = n17448 & n22443;
  assign n22551 = n20281 & n22462;
  assign n22552 = pi629 & ~n22551;
  assign n22553 = ~n22550 & n22552;
  assign n22554 = ~n22549 & ~n22553;
  assign n22555 = pi792 & n22554;
  assign n22556 = n19637 & ~n22555;
  assign n22557 = ~n22545 & n22556;
  assign n22558 = ~n22475 & ~n22557;
  assign n22559 = pi644 & n22558;
  assign n22560 = ~pi787 & ~n22463;
  assign n22561 = pi787 & ~n22472;
  assign n22562 = ~n22560 & ~n22561;
  assign n22563 = ~pi644 & n22562;
  assign n22564 = pi715 & ~n22563;
  assign n22565 = ~n22559 & n22564;
  assign n22566 = ~n17247 & ~n22446;
  assign n22567 = n17247 & n22402;
  assign n22568 = ~n22566 & ~n22567;
  assign n22569 = pi644 & ~n22568;
  assign n22570 = ~pi644 & n22402;
  assign n22571 = ~pi715 & ~n22570;
  assign n22572 = ~n22569 & n22571;
  assign n22573 = pi1160 & ~n22572;
  assign n22574 = ~n22565 & n22573;
  assign n22575 = ~pi644 & ~n22568;
  assign n22576 = pi715 & ~n22575;
  assign n22577 = pi644 & n22402;
  assign n22578 = n22576 & ~n22577;
  assign n22579 = pi644 & n22562;
  assign n22580 = ~pi644 & n22558;
  assign n22581 = ~pi715 & ~n22580;
  assign n22582 = ~n22579 & n22581;
  assign n22583 = ~pi1160 & ~n22582;
  assign n22584 = ~n22578 & n22583;
  assign n22585 = ~n22574 & ~n22584;
  assign n22586 = pi790 & ~n22585;
  assign n22587 = ~pi790 & n22558;
  assign n22588 = pi832 & ~n22587;
  assign n22589 = ~n22586 & n22588;
  assign po330 = ~n22401 & ~n22589;
  assign n22591 = ~pi174 & ~n6274;
  assign n22592 = pi174 & ~n10020;
  assign n22593 = pi759 & n16447;
  assign n22594 = ~n20854 & ~n22593;
  assign n22595 = pi39 & ~n22594;
  assign n22596 = pi759 & n16380;
  assign n22597 = ~pi759 & n16201;
  assign n22598 = ~pi39 & ~n22597;
  assign n22599 = ~n22596 & n22598;
  assign n22600 = ~n22595 & ~n22599;
  assign n22601 = pi174 & ~n22600;
  assign n22602 = ~pi174 & pi759;
  assign n22603 = n16503 & n22602;
  assign n22604 = ~n22601 & ~n22603;
  assign n22605 = ~pi38 & ~n22604;
  assign n22606 = pi759 & n16393;
  assign n22607 = n16508 & ~n22606;
  assign n22608 = ~pi174 & ~n16508;
  assign n22609 = pi38 & ~n22608;
  assign n22610 = ~n22607 & n22609;
  assign n22611 = ~n22605 & ~n22610;
  assign n22612 = n10020 & ~n22611;
  assign n22613 = ~n22592 & ~n22612;
  assign n22614 = ~n16521 & ~n22613;
  assign n22615 = pi174 & ~n16527;
  assign n22616 = n16521 & n22615;
  assign n22617 = ~n22614 & ~n22616;
  assign n22618 = ~pi785 & ~n22617;
  assign n22619 = pi609 & n22617;
  assign n22620 = ~pi609 & ~n22615;
  assign n22621 = pi1155 & ~n22620;
  assign n22622 = ~n22619 & n22621;
  assign n22623 = ~pi609 & n22617;
  assign n22624 = pi609 & ~n22615;
  assign n22625 = ~pi1155 & ~n22624;
  assign n22626 = ~n22623 & n22625;
  assign n22627 = ~n22622 & ~n22626;
  assign n22628 = pi785 & ~n22627;
  assign n22629 = ~n22618 & ~n22628;
  assign n22630 = ~pi781 & ~n22629;
  assign n22631 = pi618 & n22629;
  assign n22632 = ~pi618 & ~n22615;
  assign n22633 = pi1154 & ~n22632;
  assign n22634 = ~n22631 & n22633;
  assign n22635 = ~pi618 & n22629;
  assign n22636 = pi618 & ~n22615;
  assign n22637 = ~pi1154 & ~n22636;
  assign n22638 = ~n22635 & n22637;
  assign n22639 = ~n22634 & ~n22638;
  assign n22640 = pi781 & ~n22639;
  assign n22641 = ~n22630 & ~n22640;
  assign n22642 = ~pi789 & ~n22641;
  assign n22643 = pi619 & n22641;
  assign n22644 = ~pi619 & ~n22615;
  assign n22645 = pi1159 & ~n22644;
  assign n22646 = ~n22643 & n22645;
  assign n22647 = ~pi619 & n22641;
  assign n22648 = pi619 & ~n22615;
  assign n22649 = ~pi1159 & ~n22648;
  assign n22650 = ~n22647 & n22649;
  assign n22651 = ~n22646 & ~n22650;
  assign n22652 = pi789 & ~n22651;
  assign n22653 = ~n22642 & ~n22652;
  assign n22654 = ~n17355 & ~n22653;
  assign n22655 = n17355 & n22615;
  assign n22656 = ~n22654 & ~n22655;
  assign n22657 = ~n16124 & ~n22656;
  assign n22658 = n16124 & n22615;
  assign n22659 = ~n22657 & ~n22658;
  assign n22660 = pi647 & n22659;
  assign n22661 = pi628 & n22656;
  assign n22662 = n16593 & ~n22615;
  assign n22663 = pi696 & n10020;
  assign n22664 = ~n22615 & ~n22663;
  assign n22665 = n19410 & ~n22608;
  assign n22666 = pi174 & ~n17592;
  assign n22667 = ~pi174 & ~n17589;
  assign n22668 = ~pi38 & ~n22667;
  assign n22669 = ~n22666 & n22668;
  assign n22670 = ~n22665 & ~n22669;
  assign n22671 = n22663 & n22670;
  assign n22672 = ~n22664 & ~n22671;
  assign n22673 = ~pi778 & n22672;
  assign n22674 = pi625 & ~n22672;
  assign n22675 = ~pi625 & ~n22615;
  assign n22676 = pi1153 & ~n22675;
  assign n22677 = ~n22674 & n22676;
  assign n22678 = ~pi625 & ~n22672;
  assign n22679 = pi625 & ~n22615;
  assign n22680 = ~pi1153 & ~n22679;
  assign n22681 = ~n22678 & n22680;
  assign n22682 = ~n22677 & ~n22681;
  assign n22683 = pi778 & ~n22682;
  assign n22684 = ~n22673 & ~n22683;
  assign n22685 = ~n16593 & n22684;
  assign n22686 = ~n22662 & ~n22685;
  assign n22687 = ~n16589 & n22686;
  assign n22688 = n16589 & n22615;
  assign n22689 = ~n22687 & ~n22688;
  assign n22690 = pi619 & n22689;
  assign n22691 = pi618 & ~n22686;
  assign n22692 = pi609 & n22684;
  assign n22693 = pi625 & n22613;
  assign n22694 = ~n22612 & ~n22663;
  assign n22695 = pi174 & ~n17061;
  assign n22696 = ~pi174 & ~n17058;
  assign n22697 = ~pi759 & ~n22696;
  assign n22698 = ~n22695 & n22697;
  assign n22699 = ~pi174 & n17065;
  assign n22700 = pi174 & n17067;
  assign n22701 = ~n22699 & ~n22700;
  assign n22702 = pi759 & n22701;
  assign n22703 = ~pi39 & ~n22702;
  assign n22704 = ~n22698 & n22703;
  assign n22705 = ~pi174 & ~n16998;
  assign n22706 = pi759 & ~n22705;
  assign n22707 = pi174 & n17051;
  assign n22708 = n22706 & ~n22707;
  assign n22709 = ~pi174 & ~n16935;
  assign n22710 = pi174 & ~n16853;
  assign n22711 = ~pi759 & ~n22710;
  assign n22712 = ~n22709 & n22711;
  assign n22713 = pi39 & ~n22712;
  assign n22714 = ~n22708 & n22713;
  assign n22715 = ~pi38 & ~n22714;
  assign n22716 = ~n22704 & n22715;
  assign n22717 = pi696 & ~n22716;
  assign n22718 = ~n18932 & n22717;
  assign n22719 = ~n22610 & n22718;
  assign n22720 = ~n22694 & ~n22719;
  assign n22721 = ~n22592 & ~n22720;
  assign n22722 = ~pi625 & n22721;
  assign n22723 = ~pi1153 & ~n22722;
  assign n22724 = ~n22693 & n22723;
  assign n22725 = ~pi608 & ~n22677;
  assign n22726 = ~n22724 & n22725;
  assign n22727 = ~pi625 & n22613;
  assign n22728 = pi625 & n22721;
  assign n22729 = ~n22727 & ~n22728;
  assign n22730 = pi1153 & n22729;
  assign n22731 = ~n22681 & ~n22730;
  assign n22732 = pi608 & n22731;
  assign n22733 = ~n22726 & ~n22732;
  assign n22734 = pi778 & ~n22733;
  assign n22735 = ~pi778 & n22721;
  assign n22736 = ~n22734 & ~n22735;
  assign n22737 = ~pi609 & ~n22736;
  assign n22738 = ~pi1155 & ~n22737;
  assign n22739 = ~n22692 & n22738;
  assign n22740 = ~pi660 & ~n22622;
  assign n22741 = ~n22739 & n22740;
  assign n22742 = ~pi609 & n22684;
  assign n22743 = pi609 & ~n22736;
  assign n22744 = ~n22742 & ~n22743;
  assign n22745 = pi1155 & n22744;
  assign n22746 = ~n22626 & ~n22745;
  assign n22747 = pi660 & n22746;
  assign n22748 = ~n22741 & ~n22747;
  assign n22749 = pi785 & ~n22748;
  assign n22750 = ~pi785 & ~n22736;
  assign n22751 = ~n22749 & ~n22750;
  assign n22752 = ~pi618 & ~n22751;
  assign n22753 = ~pi1154 & ~n22752;
  assign n22754 = ~n22691 & n22753;
  assign n22755 = ~pi627 & ~n22634;
  assign n22756 = ~n22754 & n22755;
  assign n22757 = ~pi618 & ~n22686;
  assign n22758 = pi618 & ~n22751;
  assign n22759 = ~n22757 & ~n22758;
  assign n22760 = pi1154 & n22759;
  assign n22761 = ~n22638 & ~n22760;
  assign n22762 = pi627 & n22761;
  assign n22763 = ~n22756 & ~n22762;
  assign n22764 = pi781 & ~n22763;
  assign n22765 = ~pi781 & ~n22751;
  assign n22766 = ~n22764 & ~n22765;
  assign n22767 = ~pi619 & ~n22766;
  assign n22768 = ~pi1159 & ~n22767;
  assign n22769 = ~n22690 & n22768;
  assign n22770 = ~pi648 & ~n22646;
  assign n22771 = ~n22769 & n22770;
  assign n22772 = ~pi619 & n22689;
  assign n22773 = pi619 & ~n22766;
  assign n22774 = ~n22772 & ~n22773;
  assign n22775 = pi1159 & n22774;
  assign n22776 = ~n22650 & ~n22775;
  assign n22777 = pi648 & n22776;
  assign n22778 = ~n22771 & ~n22777;
  assign n22779 = pi789 & ~n22778;
  assign n22780 = ~pi789 & ~n22766;
  assign n22781 = ~n22779 & ~n22780;
  assign n22782 = ~pi788 & n22781;
  assign n22783 = pi626 & n22781;
  assign n22784 = n17159 & ~n22615;
  assign n22785 = ~n17159 & n22689;
  assign n22786 = ~n22784 & ~n22785;
  assign n22787 = ~pi626 & n22786;
  assign n22788 = pi641 & ~n22787;
  assign n22789 = ~n22783 & n22788;
  assign n22790 = pi626 & ~n22653;
  assign n22791 = ~pi626 & n22615;
  assign n22792 = ~pi641 & ~n22791;
  assign n22793 = ~n22790 & n22792;
  assign n22794 = pi1158 & ~n22793;
  assign n22795 = ~n22789 & n22794;
  assign n22796 = ~pi626 & ~n22653;
  assign n22797 = pi641 & ~n22796;
  assign n22798 = pi626 & n22615;
  assign n22799 = n22797 & ~n22798;
  assign n22800 = pi626 & n22786;
  assign n22801 = ~pi626 & n22781;
  assign n22802 = ~pi641 & ~n22801;
  assign n22803 = ~n22800 & n22802;
  assign n22804 = ~pi1158 & ~n22803;
  assign n22805 = ~n22799 & n22804;
  assign n22806 = ~n22795 & ~n22805;
  assign n22807 = pi788 & ~n22806;
  assign n22808 = ~n22782 & ~n22807;
  assign n22809 = ~pi628 & n22808;
  assign n22810 = ~pi1156 & ~n22809;
  assign n22811 = ~n22661 & n22810;
  assign n22812 = ~n17183 & n22786;
  assign n22813 = n17183 & n22615;
  assign n22814 = ~n22812 & ~n22813;
  assign n22815 = pi628 & n22814;
  assign n22816 = ~pi628 & ~n22615;
  assign n22817 = pi1156 & ~n22816;
  assign n22818 = ~n22815 & n22817;
  assign n22819 = ~pi629 & ~n22818;
  assign n22820 = ~n22811 & n22819;
  assign n22821 = ~pi628 & n22814;
  assign n22822 = pi628 & ~n22615;
  assign n22823 = ~pi1156 & ~n22822;
  assign n22824 = ~n22821 & n22823;
  assign n22825 = ~pi628 & n22656;
  assign n22826 = pi628 & n22808;
  assign n22827 = ~n22825 & ~n22826;
  assign n22828 = pi1156 & n22827;
  assign n22829 = ~n22824 & ~n22828;
  assign n22830 = pi629 & n22829;
  assign n22831 = ~n22820 & ~n22830;
  assign n22832 = pi792 & ~n22831;
  assign n22833 = ~pi792 & n22808;
  assign n22834 = ~n22832 & ~n22833;
  assign n22835 = ~pi647 & ~n22834;
  assign n22836 = ~pi1157 & ~n22835;
  assign n22837 = ~n22660 & n22836;
  assign n22838 = ~pi792 & ~n22814;
  assign n22839 = ~n22818 & ~n22824;
  assign n22840 = pi792 & ~n22839;
  assign n22841 = ~n22838 & ~n22840;
  assign n22842 = pi647 & n22841;
  assign n22843 = ~pi647 & ~n22615;
  assign n22844 = pi1157 & ~n22843;
  assign n22845 = ~n22842 & n22844;
  assign n22846 = ~pi630 & ~n22845;
  assign n22847 = ~n22837 & n22846;
  assign n22848 = ~pi647 & n22841;
  assign n22849 = pi647 & ~n22615;
  assign n22850 = ~pi1157 & ~n22849;
  assign n22851 = ~n22848 & n22850;
  assign n22852 = ~pi647 & n22659;
  assign n22853 = pi647 & ~n22834;
  assign n22854 = ~n22852 & ~n22853;
  assign n22855 = pi1157 & n22854;
  assign n22856 = ~n22851 & ~n22855;
  assign n22857 = pi630 & n22856;
  assign n22858 = ~n22847 & ~n22857;
  assign n22859 = pi787 & ~n22858;
  assign n22860 = ~pi787 & ~n22834;
  assign n22861 = ~n22859 & ~n22860;
  assign n22862 = ~pi790 & n22861;
  assign n22863 = pi644 & ~n22861;
  assign n22864 = ~pi787 & ~n22841;
  assign n22865 = ~n22845 & ~n22851;
  assign n22866 = pi787 & ~n22865;
  assign n22867 = ~n22864 & ~n22866;
  assign n22868 = ~pi644 & n22867;
  assign n22869 = pi715 & ~n22868;
  assign n22870 = ~n22863 & n22869;
  assign n22871 = ~pi644 & ~n22615;
  assign n22872 = n17247 & ~n22615;
  assign n22873 = ~n17247 & n22659;
  assign n22874 = ~n22872 & ~n22873;
  assign n22875 = pi644 & ~n22874;
  assign n22876 = ~pi715 & ~n22875;
  assign n22877 = ~n22871 & n22876;
  assign n22878 = ~n22870 & ~n22877;
  assign n22879 = pi1160 & n22878;
  assign n22880 = pi644 & ~n22615;
  assign n22881 = ~pi644 & ~n22874;
  assign n22882 = pi715 & ~n22881;
  assign n22883 = ~n22880 & n22882;
  assign n22884 = pi644 & n22867;
  assign n22885 = ~pi644 & ~n22861;
  assign n22886 = ~pi715 & ~n22885;
  assign n22887 = ~n22884 & n22886;
  assign n22888 = ~n22883 & ~n22887;
  assign n22889 = ~pi1160 & n22888;
  assign n22890 = ~n22879 & ~n22889;
  assign n22891 = pi790 & n22890;
  assign n22892 = ~n22862 & ~n22891;
  assign n22893 = n6274 & n22892;
  assign n22894 = ~pi57 & ~n22893;
  assign n22895 = ~n22591 & n22894;
  assign n22896 = pi57 & pi174;
  assign n22897 = ~pi832 & ~n22896;
  assign n22898 = ~n22895 & n22897;
  assign n22899 = pi174 & ~n2934;
  assign n22900 = pi696 & n16742;
  assign n22901 = ~n22899 & ~n22900;
  assign n22902 = ~pi778 & n22901;
  assign n22903 = pi625 & n22900;
  assign n22904 = ~n22901 & ~n22903;
  assign n22905 = ~pi1153 & ~n22904;
  assign n22906 = pi1153 & ~n22899;
  assign n22907 = ~n22903 & n22906;
  assign n22908 = ~n22905 & ~n22907;
  assign n22909 = pi778 & ~n22908;
  assign n22910 = ~n22902 & ~n22909;
  assign n22911 = n18715 & n22910;
  assign n22912 = ~n17159 & n22911;
  assign n22913 = ~n22899 & ~n22912;
  assign n22914 = n17345 & ~n22913;
  assign n22915 = pi759 & n16510;
  assign n22916 = ~n19656 & n22915;
  assign n22917 = ~n19662 & n22916;
  assign n22918 = n19668 & n22917;
  assign n22919 = pi626 & n22918;
  assign n22920 = ~n22899 & ~n22919;
  assign n22921 = pi1158 & ~n22920;
  assign n22922 = ~pi641 & ~n22921;
  assign n22923 = ~n22914 & n22922;
  assign n22924 = ~pi626 & n22918;
  assign n22925 = ~n22899 & ~n22924;
  assign n22926 = ~pi1158 & ~n22925;
  assign n22927 = n17344 & ~n22913;
  assign n22928 = pi641 & ~n22927;
  assign n22929 = ~n22926 & n22928;
  assign n22930 = ~n22923 & ~n22929;
  assign n22931 = pi788 & n22930;
  assign n22932 = ~n17338 & n22910;
  assign n22933 = pi618 & n22932;
  assign n22934 = pi609 & n22910;
  assign n22935 = ~n22899 & ~n22915;
  assign n22936 = ~n16393 & n22900;
  assign n22937 = n22935 & ~n22936;
  assign n22938 = pi625 & n22936;
  assign n22939 = ~n22937 & ~n22938;
  assign n22940 = ~pi1153 & ~n22939;
  assign n22941 = ~pi608 & ~n22907;
  assign n22942 = ~n22940 & n22941;
  assign n22943 = pi1153 & ~n22938;
  assign n22944 = n22935 & n22943;
  assign n22945 = ~n22905 & ~n22944;
  assign n22946 = pi608 & n22945;
  assign n22947 = ~n22942 & ~n22946;
  assign n22948 = pi778 & ~n22947;
  assign n22949 = ~pi778 & ~n22937;
  assign n22950 = ~n22948 & ~n22949;
  assign n22951 = ~pi609 & ~n22950;
  assign n22952 = ~pi1155 & ~n22951;
  assign n22953 = ~n22934 & n22952;
  assign n22954 = ~n17279 & ~n22935;
  assign n22955 = pi1155 & ~n22954;
  assign n22956 = ~pi660 & ~n22955;
  assign n22957 = ~n22953 & n22956;
  assign n22958 = ~pi609 & n22910;
  assign n22959 = pi609 & ~n22950;
  assign n22960 = ~n22958 & ~n22959;
  assign n22961 = pi1155 & n22960;
  assign n22962 = ~pi1155 & ~n22899;
  assign n22963 = n16537 & n22915;
  assign n22964 = n22962 & ~n22963;
  assign n22965 = pi660 & ~n22964;
  assign n22966 = ~n22961 & n22965;
  assign n22967 = ~n22957 & ~n22966;
  assign n22968 = pi785 & ~n22967;
  assign n22969 = ~pi785 & ~n22950;
  assign n22970 = ~n22968 & ~n22969;
  assign n22971 = ~pi618 & ~n22970;
  assign n22972 = ~pi1154 & ~n22971;
  assign n22973 = ~n22933 & n22972;
  assign n22974 = ~pi627 & ~n22973;
  assign n22975 = n19744 & n22916;
  assign n22976 = ~n22899 & ~n22975;
  assign n22977 = pi1154 & n22976;
  assign n22978 = n22974 & ~n22977;
  assign n22979 = ~pi618 & n22932;
  assign n22980 = pi618 & ~n22970;
  assign n22981 = ~n22979 & ~n22980;
  assign n22982 = pi1154 & n22981;
  assign n22983 = n19753 & n22916;
  assign n22984 = ~pi1154 & ~n22899;
  assign n22985 = ~n22983 & n22984;
  assign n22986 = pi627 & ~n22985;
  assign n22987 = ~n22982 & n22986;
  assign n22988 = ~n22978 & ~n22987;
  assign n22989 = pi781 & ~n22988;
  assign n22990 = ~pi781 & ~n22970;
  assign n22991 = ~n17159 & ~n19667;
  assign n22992 = ~n22990 & n22991;
  assign n22993 = ~n22989 & n22992;
  assign n22994 = pi648 & n19664;
  assign n22995 = ~pi648 & n19665;
  assign n22996 = ~n22994 & ~n22995;
  assign n22997 = ~n22911 & ~n22996;
  assign n22998 = n19776 & n22917;
  assign n22999 = n17156 & ~n22998;
  assign n23000 = n19766 & n22917;
  assign n23001 = n17157 & ~n23000;
  assign n23002 = ~n22999 & ~n23001;
  assign n23003 = ~n22997 & n23002;
  assign n23004 = pi789 & ~n22899;
  assign n23005 = ~n23003 & n23004;
  assign n23006 = n17356 & ~n23005;
  assign n23007 = ~n22993 & n23006;
  assign n23008 = ~n22931 & ~n23007;
  assign n23009 = n19788 & n23008;
  assign n23010 = ~n17355 & n22918;
  assign n23011 = ~pi629 & n23010;
  assign n23012 = pi628 & ~n23011;
  assign n23013 = n18717 & n22910;
  assign n23014 = pi629 & ~n23013;
  assign n23015 = ~n23012 & ~n23014;
  assign n23016 = ~pi1156 & ~n23015;
  assign n23017 = pi628 & n23013;
  assign n23018 = ~pi628 & ~n23010;
  assign n23019 = pi629 & ~n23018;
  assign n23020 = pi1156 & ~n23019;
  assign n23021 = ~n23017 & n23020;
  assign n23022 = ~n23016 & ~n23021;
  assign n23023 = ~n22899 & ~n23022;
  assign n23024 = pi792 & n23023;
  assign n23025 = ~n23009 & ~n23024;
  assign n23026 = n19637 & ~n23025;
  assign n23027 = ~n16124 & n23010;
  assign n23028 = ~pi630 & n23027;
  assign n23029 = pi647 & ~n23028;
  assign n23030 = ~n18744 & n23013;
  assign n23031 = pi630 & ~n23030;
  assign n23032 = ~n23029 & ~n23031;
  assign n23033 = ~pi1157 & ~n23032;
  assign n23034 = ~pi630 & ~n23030;
  assign n23035 = pi647 & ~n23034;
  assign n23036 = pi630 & n23027;
  assign n23037 = pi1157 & ~n23036;
  assign n23038 = ~n23035 & n23037;
  assign n23039 = ~n23033 & ~n23038;
  assign n23040 = ~n22899 & ~n23039;
  assign n23041 = pi787 & n23040;
  assign n23042 = ~n23026 & ~n23041;
  assign n23043 = pi644 & n23042;
  assign n23044 = ~n18767 & n23030;
  assign n23045 = ~n22899 & ~n23044;
  assign n23046 = ~pi644 & ~n23045;
  assign n23047 = pi715 & ~n23046;
  assign n23048 = ~n23043 & n23047;
  assign n23049 = ~n16124 & ~n17247;
  assign n23050 = n23010 & n23049;
  assign n23051 = pi644 & n23050;
  assign n23052 = ~pi715 & ~n22899;
  assign n23053 = ~n23051 & n23052;
  assign n23054 = pi1160 & ~n23053;
  assign n23055 = ~n23048 & n23054;
  assign n23056 = pi644 & ~n23045;
  assign n23057 = ~pi644 & n23042;
  assign n23058 = ~pi715 & ~n23057;
  assign n23059 = ~n23056 & n23058;
  assign n23060 = ~pi1160 & ~n23059;
  assign n23061 = ~pi644 & n23050;
  assign n23062 = ~n22899 & ~n23061;
  assign n23063 = pi715 & n23062;
  assign n23064 = n23060 & ~n23063;
  assign n23065 = ~n23055 & ~n23064;
  assign n23066 = pi790 & ~n23065;
  assign n23067 = ~pi790 & n23042;
  assign n23068 = pi832 & ~n23067;
  assign n23069 = ~n23066 & n23068;
  assign po331 = ~n22898 & ~n23069;
  assign n23071 = ~pi175 & ~n2934;
  assign n23072 = pi766 & n16510;
  assign n23073 = ~n23071 & ~n23072;
  assign n23074 = ~n17273 & ~n23073;
  assign n23075 = ~pi785 & ~n23074;
  assign n23076 = n16537 & n23072;
  assign n23077 = n23074 & ~n23076;
  assign n23078 = pi1155 & ~n23077;
  assign n23079 = ~pi1155 & ~n23071;
  assign n23080 = ~n23076 & n23079;
  assign n23081 = ~n23078 & ~n23080;
  assign n23082 = pi785 & ~n23081;
  assign n23083 = ~n23075 & ~n23082;
  assign n23084 = ~pi781 & ~n23083;
  assign n23085 = ~n17289 & n23083;
  assign n23086 = pi1154 & ~n23085;
  assign n23087 = ~n17292 & n23083;
  assign n23088 = ~pi1154 & ~n23087;
  assign n23089 = ~n23086 & ~n23088;
  assign n23090 = pi781 & ~n23089;
  assign n23091 = ~n23084 & ~n23090;
  assign n23092 = ~pi789 & ~n23091;
  assign n23093 = ~n22423 & n23091;
  assign n23094 = pi1159 & ~n23093;
  assign n23095 = ~n22426 & n23091;
  assign n23096 = ~pi1159 & ~n23095;
  assign n23097 = ~n23094 & ~n23096;
  assign n23098 = pi789 & ~n23097;
  assign n23099 = ~n23092 & ~n23098;
  assign n23100 = ~n17355 & n23099;
  assign n23101 = n17355 & n23071;
  assign n23102 = ~n23100 & ~n23101;
  assign n23103 = ~n16124 & ~n23102;
  assign n23104 = n16124 & n23071;
  assign n23105 = ~n23103 & ~n23104;
  assign n23106 = ~n19987 & n23105;
  assign n23107 = pi700 & n16742;
  assign n23108 = ~n23071 & ~n23107;
  assign n23109 = ~pi778 & ~n23108;
  assign n23110 = ~pi625 & n23107;
  assign n23111 = ~n23108 & ~n23110;
  assign n23112 = pi1153 & ~n23111;
  assign n23113 = ~pi1153 & ~n23071;
  assign n23114 = ~n23110 & n23113;
  assign n23115 = ~n23112 & ~n23114;
  assign n23116 = pi778 & n23115;
  assign n23117 = ~n23109 & ~n23116;
  assign n23118 = ~n17338 & ~n23117;
  assign n23119 = ~n17340 & n23118;
  assign n23120 = ~n17342 & n23119;
  assign n23121 = ~n17425 & n23120;
  assign n23122 = ~n17452 & n23121;
  assign n23123 = ~pi647 & n23122;
  assign n23124 = pi647 & n23071;
  assign n23125 = ~pi1157 & ~n23124;
  assign n23126 = ~n23123 & n23125;
  assign n23127 = ~pi647 & n23071;
  assign n23128 = pi647 & n23122;
  assign n23129 = pi1157 & ~n23128;
  assign n23130 = ~n23127 & n23129;
  assign n23131 = ~n23126 & ~n23130;
  assign n23132 = ~n17246 & ~n23131;
  assign n23133 = ~n23106 & ~n23132;
  assign n23134 = pi787 & ~n23133;
  assign n23135 = ~pi626 & ~n23099;
  assign n23136 = pi626 & ~n23071;
  assign n23137 = n17181 & ~n23136;
  assign n23138 = ~n23135 & n23137;
  assign n23139 = n17350 & n23120;
  assign n23140 = pi626 & ~n23099;
  assign n23141 = ~pi626 & ~n23071;
  assign n23142 = n17180 & ~n23141;
  assign n23143 = ~n23140 & n23142;
  assign n23144 = ~n23139 & ~n23143;
  assign n23145 = ~n23138 & n23144;
  assign n23146 = pi788 & ~n23145;
  assign n23147 = pi618 & n23118;
  assign n23148 = pi609 & ~n23117;
  assign n23149 = ~n16393 & ~n23108;
  assign n23150 = pi625 & n23149;
  assign n23151 = n23073 & ~n23149;
  assign n23152 = ~n23150 & ~n23151;
  assign n23153 = n23113 & ~n23152;
  assign n23154 = ~pi608 & ~n23112;
  assign n23155 = ~n23153 & n23154;
  assign n23156 = pi1153 & ~n23150;
  assign n23157 = n23073 & n23156;
  assign n23158 = ~n23114 & ~n23157;
  assign n23159 = pi608 & n23158;
  assign n23160 = ~n23155 & ~n23159;
  assign n23161 = pi778 & ~n23160;
  assign n23162 = ~pi778 & ~n23151;
  assign n23163 = ~n23161 & ~n23162;
  assign n23164 = ~pi609 & ~n23163;
  assign n23165 = ~pi1155 & ~n23164;
  assign n23166 = ~n23148 & n23165;
  assign n23167 = ~pi660 & ~n23078;
  assign n23168 = ~n23166 & n23167;
  assign n23169 = ~pi609 & ~n23117;
  assign n23170 = pi609 & ~n23163;
  assign n23171 = ~n23169 & ~n23170;
  assign n23172 = pi1155 & n23171;
  assign n23173 = ~n23080 & ~n23172;
  assign n23174 = pi660 & n23173;
  assign n23175 = ~n23168 & ~n23174;
  assign n23176 = pi785 & ~n23175;
  assign n23177 = ~pi785 & ~n23163;
  assign n23178 = ~n23176 & ~n23177;
  assign n23179 = ~pi618 & ~n23178;
  assign n23180 = ~pi1154 & ~n23179;
  assign n23181 = ~n23147 & n23180;
  assign n23182 = ~pi627 & ~n23086;
  assign n23183 = ~n23181 & n23182;
  assign n23184 = ~pi618 & n23118;
  assign n23185 = pi618 & ~n23178;
  assign n23186 = ~n23184 & ~n23185;
  assign n23187 = pi1154 & n23186;
  assign n23188 = ~n23088 & ~n23187;
  assign n23189 = pi627 & n23188;
  assign n23190 = ~n23183 & ~n23189;
  assign n23191 = pi781 & ~n23190;
  assign n23192 = ~pi781 & ~n23178;
  assign n23193 = ~n23191 & ~n23192;
  assign n23194 = ~pi619 & ~n23193;
  assign n23195 = pi619 & n23119;
  assign n23196 = ~pi1159 & ~n23195;
  assign n23197 = ~n23194 & n23196;
  assign n23198 = ~pi648 & ~n23197;
  assign n23199 = ~n23094 & n23198;
  assign n23200 = ~pi619 & n23119;
  assign n23201 = pi619 & ~n23193;
  assign n23202 = ~n23200 & ~n23201;
  assign n23203 = pi1159 & n23202;
  assign n23204 = ~n23096 & ~n23203;
  assign n23205 = pi648 & n23204;
  assign n23206 = ~n23199 & ~n23205;
  assign n23207 = pi789 & n23206;
  assign n23208 = ~pi789 & n23193;
  assign n23209 = n17356 & ~n23208;
  assign n23210 = ~n23207 & n23209;
  assign n23211 = ~n23146 & ~n23210;
  assign n23212 = n19788 & ~n23211;
  assign n23213 = n20275 & n23121;
  assign n23214 = n17449 & ~n23102;
  assign n23215 = ~pi629 & ~n23214;
  assign n23216 = ~n23213 & n23215;
  assign n23217 = n17448 & ~n23102;
  assign n23218 = n20281 & n23121;
  assign n23219 = pi629 & ~n23218;
  assign n23220 = ~n23217 & n23219;
  assign n23221 = ~n23216 & ~n23220;
  assign n23222 = pi792 & n23221;
  assign n23223 = n19637 & ~n23222;
  assign n23224 = ~n23212 & n23223;
  assign n23225 = ~n23134 & ~n23224;
  assign n23226 = pi644 & n23225;
  assign n23227 = ~pi787 & ~n23122;
  assign n23228 = pi787 & ~n23131;
  assign n23229 = ~n23227 & ~n23228;
  assign n23230 = ~pi644 & n23229;
  assign n23231 = pi715 & ~n23230;
  assign n23232 = ~n23226 & n23231;
  assign n23233 = ~n17247 & ~n23105;
  assign n23234 = n17247 & n23071;
  assign n23235 = ~n23233 & ~n23234;
  assign n23236 = pi644 & ~n23235;
  assign n23237 = ~pi644 & n23071;
  assign n23238 = ~pi715 & ~n23237;
  assign n23239 = ~n23236 & n23238;
  assign n23240 = pi1160 & ~n23239;
  assign n23241 = ~n23232 & n23240;
  assign n23242 = ~pi644 & ~n23235;
  assign n23243 = pi715 & ~n23242;
  assign n23244 = pi644 & n23071;
  assign n23245 = n23243 & ~n23244;
  assign n23246 = pi644 & n23229;
  assign n23247 = ~pi644 & n23225;
  assign n23248 = ~pi715 & ~n23247;
  assign n23249 = ~n23246 & n23248;
  assign n23250 = ~pi1160 & ~n23249;
  assign n23251 = ~n23245 & n23250;
  assign n23252 = ~n23241 & ~n23251;
  assign n23253 = pi790 & ~n23252;
  assign n23254 = ~pi790 & n23225;
  assign n23255 = pi832 & ~n23254;
  assign n23256 = ~n23253 & n23255;
  assign n23257 = ~pi175 & ~n16527;
  assign n23258 = n17451 & ~n23257;
  assign n23259 = n17159 & ~n23257;
  assign n23260 = n16593 & ~n23257;
  assign n23261 = pi175 & ~n10020;
  assign n23262 = pi175 & n17589;
  assign n23263 = ~pi175 & n17592;
  assign n23264 = ~pi38 & ~n23263;
  assign n23265 = ~n23262 & n23264;
  assign n23266 = ~pi175 & ~n16508;
  assign n23267 = n16744 & ~n23266;
  assign n23268 = pi700 & ~n23267;
  assign n23269 = ~n23265 & n23268;
  assign n23270 = ~pi175 & ~pi700;
  assign n23271 = ~n16526 & n23270;
  assign n23272 = ~n23269 & ~n23271;
  assign n23273 = n10020 & n23272;
  assign n23274 = ~n23261 & ~n23273;
  assign n23275 = ~pi778 & ~n23274;
  assign n23276 = pi625 & n23274;
  assign n23277 = pi1153 & ~n23276;
  assign n23278 = ~pi625 & n23257;
  assign n23279 = n23277 & ~n23278;
  assign n23280 = ~pi625 & n23274;
  assign n23281 = ~pi1153 & ~n23280;
  assign n23282 = pi625 & n23257;
  assign n23283 = n23281 & ~n23282;
  assign n23284 = ~n23279 & ~n23283;
  assign n23285 = pi778 & ~n23284;
  assign n23286 = ~n23275 & ~n23285;
  assign n23287 = ~n16593 & ~n23286;
  assign n23288 = ~n23260 & ~n23287;
  assign n23289 = ~n16589 & n23288;
  assign n23290 = n16589 & n23257;
  assign n23291 = ~n23289 & ~n23290;
  assign n23292 = ~n17159 & n23291;
  assign n23293 = ~n23259 & ~n23292;
  assign n23294 = ~n17183 & n23293;
  assign n23295 = n17183 & n23257;
  assign n23296 = ~n23294 & ~n23295;
  assign n23297 = ~n17451 & n23296;
  assign n23298 = ~n23258 & ~n23297;
  assign n23299 = ~n18767 & n23298;
  assign n23300 = n18767 & n23257;
  assign n23301 = ~n23299 & ~n23300;
  assign n23302 = ~pi644 & ~n23301;
  assign n23303 = pi715 & ~n23302;
  assign n23304 = n17247 & ~n23257;
  assign n23305 = ~pi766 & n16355;
  assign n23306 = pi175 & n16501;
  assign n23307 = ~n23305 & ~n23306;
  assign n23308 = pi39 & ~n23307;
  assign n23309 = pi766 & ~n16461;
  assign n23310 = pi175 & ~n23309;
  assign n23311 = ~n20899 & ~n23310;
  assign n23312 = ~pi175 & n16449;
  assign n23313 = pi766 & n23312;
  assign n23314 = n23311 & ~n23313;
  assign n23315 = ~n23308 & n23314;
  assign n23316 = ~pi38 & ~n23315;
  assign n23317 = pi766 & n16511;
  assign n23318 = ~n23266 & ~n23317;
  assign n23319 = pi38 & n23318;
  assign n23320 = ~n23316 & ~n23319;
  assign n23321 = n10020 & ~n23320;
  assign n23322 = ~n23261 & ~n23321;
  assign n23323 = ~n16521 & ~n23322;
  assign n23324 = n16521 & ~n23257;
  assign n23325 = ~n23323 & ~n23324;
  assign n23326 = ~pi785 & ~n23325;
  assign n23327 = ~n16532 & ~n23257;
  assign n23328 = pi609 & n23323;
  assign n23329 = ~n23327 & ~n23328;
  assign n23330 = pi1155 & ~n23329;
  assign n23331 = ~n16537 & ~n23257;
  assign n23332 = ~pi609 & n23323;
  assign n23333 = ~n23331 & ~n23332;
  assign n23334 = ~pi1155 & ~n23333;
  assign n23335 = ~n23330 & ~n23334;
  assign n23336 = pi785 & ~n23335;
  assign n23337 = ~n23326 & ~n23336;
  assign n23338 = ~pi781 & ~n23337;
  assign n23339 = pi618 & n23337;
  assign n23340 = ~pi618 & n23257;
  assign n23341 = pi1154 & ~n23340;
  assign n23342 = ~n23339 & n23341;
  assign n23343 = ~pi618 & n23337;
  assign n23344 = pi618 & n23257;
  assign n23345 = ~pi1154 & ~n23344;
  assign n23346 = ~n23343 & n23345;
  assign n23347 = ~n23342 & ~n23346;
  assign n23348 = pi781 & ~n23347;
  assign n23349 = ~n23338 & ~n23348;
  assign n23350 = ~pi789 & ~n23349;
  assign n23351 = pi619 & n23349;
  assign n23352 = ~pi619 & n23257;
  assign n23353 = pi1159 & ~n23352;
  assign n23354 = ~n23351 & n23353;
  assign n23355 = ~pi619 & n23349;
  assign n23356 = pi619 & n23257;
  assign n23357 = ~pi1159 & ~n23356;
  assign n23358 = ~n23355 & n23357;
  assign n23359 = ~n23354 & ~n23358;
  assign n23360 = pi789 & ~n23359;
  assign n23361 = ~n23350 & ~n23360;
  assign n23362 = ~n17355 & n23361;
  assign n23363 = n17355 & n23257;
  assign n23364 = ~n23362 & ~n23363;
  assign n23365 = ~n16124 & ~n23364;
  assign n23366 = n16124 & n23257;
  assign n23367 = ~n23365 & ~n23366;
  assign n23368 = ~n17247 & n23367;
  assign n23369 = ~n23304 & ~n23368;
  assign n23370 = pi644 & n23369;
  assign n23371 = ~pi644 & n23257;
  assign n23372 = ~pi715 & ~n23371;
  assign n23373 = ~n23370 & n23372;
  assign n23374 = pi1160 & ~n23373;
  assign n23375 = ~n23303 & n23374;
  assign n23376 = pi644 & ~n23301;
  assign n23377 = ~pi715 & ~n23376;
  assign n23378 = ~pi644 & n23369;
  assign n23379 = pi644 & n23257;
  assign n23380 = ~n23378 & ~n23379;
  assign n23381 = pi715 & n23380;
  assign n23382 = ~pi1160 & ~n23381;
  assign n23383 = ~n23377 & n23382;
  assign n23384 = ~n23375 & ~n23383;
  assign n23385 = pi790 & ~n23384;
  assign n23386 = ~n19999 & n23364;
  assign n23387 = pi628 & ~n23296;
  assign n23388 = n16121 & ~n23387;
  assign n23389 = ~pi628 & n23257;
  assign n23390 = n23388 & ~n23389;
  assign n23391 = ~pi628 & ~n23296;
  assign n23392 = pi628 & n23257;
  assign n23393 = n16122 & ~n23392;
  assign n23394 = ~n23391 & n23393;
  assign n23395 = ~n23390 & ~n23394;
  assign n23396 = ~n23386 & n23395;
  assign n23397 = pi792 & ~n23396;
  assign n23398 = pi618 & n23288;
  assign n23399 = pi609 & n23286;
  assign n23400 = pi625 & n23322;
  assign n23401 = ~pi700 & n23320;
  assign n23402 = ~pi175 & ~n17051;
  assign n23403 = pi766 & ~n23402;
  assign n23404 = pi175 & n16998;
  assign n23405 = n23403 & ~n23404;
  assign n23406 = pi175 & n16935;
  assign n23407 = ~pi175 & n16853;
  assign n23408 = ~pi766 & ~n23407;
  assign n23409 = ~n23406 & n23408;
  assign n23410 = pi39 & ~n23409;
  assign n23411 = ~n23405 & n23410;
  assign n23412 = pi175 & n17058;
  assign n23413 = ~pi175 & n17061;
  assign n23414 = ~pi766 & ~n23413;
  assign n23415 = ~n23412 & n23414;
  assign n23416 = ~pi175 & ~n17067;
  assign n23417 = pi175 & ~n17065;
  assign n23418 = ~n23416 & ~n23417;
  assign n23419 = pi766 & n23418;
  assign n23420 = ~pi39 & ~n23419;
  assign n23421 = ~n23415 & n23420;
  assign n23422 = ~pi38 & ~n23421;
  assign n23423 = ~n23411 & n23422;
  assign n23424 = ~n17079 & ~n23072;
  assign n23425 = pi175 & ~n23424;
  assign n23426 = n6097 & n23425;
  assign n23427 = n16212 & ~n16775;
  assign n23428 = ~pi766 & n23427;
  assign n23429 = ~n16917 & ~n23428;
  assign n23430 = ~pi39 & ~n23429;
  assign n23431 = ~pi175 & ~n23430;
  assign n23432 = pi38 & ~n23431;
  assign n23433 = ~n23426 & n23432;
  assign n23434 = ~n23423 & ~n23433;
  assign n23435 = pi700 & n23434;
  assign n23436 = ~n23401 & ~n23435;
  assign n23437 = n10020 & n23436;
  assign n23438 = ~n23261 & ~n23437;
  assign n23439 = ~pi625 & n23438;
  assign n23440 = ~pi1153 & ~n23439;
  assign n23441 = ~n23400 & n23440;
  assign n23442 = ~pi608 & ~n23279;
  assign n23443 = ~n23441 & n23442;
  assign n23444 = ~pi625 & n23322;
  assign n23445 = pi625 & n23438;
  assign n23446 = ~n23444 & ~n23445;
  assign n23447 = pi1153 & n23446;
  assign n23448 = ~n23283 & ~n23447;
  assign n23449 = pi608 & n23448;
  assign n23450 = ~n23443 & ~n23449;
  assign n23451 = pi778 & ~n23450;
  assign n23452 = ~pi778 & n23438;
  assign n23453 = ~n23451 & ~n23452;
  assign n23454 = ~pi609 & ~n23453;
  assign n23455 = ~pi1155 & ~n23454;
  assign n23456 = ~n23399 & n23455;
  assign n23457 = ~pi660 & ~n23330;
  assign n23458 = ~n23456 & n23457;
  assign n23459 = ~pi609 & n23286;
  assign n23460 = pi609 & ~n23453;
  assign n23461 = ~n23459 & ~n23460;
  assign n23462 = pi1155 & n23461;
  assign n23463 = ~n23334 & ~n23462;
  assign n23464 = pi660 & n23463;
  assign n23465 = ~n23458 & ~n23464;
  assign n23466 = pi785 & ~n23465;
  assign n23467 = ~pi785 & ~n23453;
  assign n23468 = ~n23466 & ~n23467;
  assign n23469 = ~pi618 & ~n23468;
  assign n23470 = ~pi1154 & ~n23469;
  assign n23471 = ~n23398 & n23470;
  assign n23472 = ~pi627 & ~n23342;
  assign n23473 = ~n23471 & n23472;
  assign n23474 = ~pi618 & n23288;
  assign n23475 = pi618 & ~n23468;
  assign n23476 = ~n23474 & ~n23475;
  assign n23477 = pi1154 & n23476;
  assign n23478 = ~n23346 & ~n23477;
  assign n23479 = pi627 & n23478;
  assign n23480 = ~n23473 & ~n23479;
  assign n23481 = pi781 & ~n23480;
  assign n23482 = ~pi781 & ~n23468;
  assign n23483 = ~n23481 & ~n23482;
  assign n23484 = ~pi789 & n23483;
  assign n23485 = ~pi619 & ~n23483;
  assign n23486 = pi619 & ~n23291;
  assign n23487 = ~pi1159 & ~n23486;
  assign n23488 = ~n23485 & n23487;
  assign n23489 = ~pi648 & ~n23488;
  assign n23490 = ~n23354 & n23489;
  assign n23491 = ~pi619 & ~n23291;
  assign n23492 = pi619 & ~n23483;
  assign n23493 = ~n23491 & ~n23492;
  assign n23494 = pi1159 & n23493;
  assign n23495 = ~n23358 & ~n23494;
  assign n23496 = pi648 & n23495;
  assign n23497 = ~n23490 & ~n23496;
  assign n23498 = pi789 & n23497;
  assign n23499 = ~n23484 & ~n23498;
  assign n23500 = n17356 & n23499;
  assign n23501 = ~pi626 & ~n23361;
  assign n23502 = pi626 & ~n23257;
  assign n23503 = n17181 & ~n23502;
  assign n23504 = ~n23501 & n23503;
  assign n23505 = n17350 & n23293;
  assign n23506 = pi626 & ~n23361;
  assign n23507 = ~pi626 & ~n23257;
  assign n23508 = n17180 & ~n23507;
  assign n23509 = ~n23506 & n23508;
  assign n23510 = ~n23505 & ~n23509;
  assign n23511 = ~n23504 & n23510;
  assign n23512 = pi788 & ~n23511;
  assign n23513 = n19788 & ~n23512;
  assign n23514 = ~n23500 & n23513;
  assign n23515 = ~n23397 & ~n23514;
  assign n23516 = n19637 & ~n23515;
  assign n23517 = ~pi647 & n23298;
  assign n23518 = pi647 & n23257;
  assign n23519 = n17245 & ~n23518;
  assign n23520 = ~n23517 & n23519;
  assign n23521 = ~n19987 & n23367;
  assign n23522 = pi647 & n23298;
  assign n23523 = n17244 & ~n23522;
  assign n23524 = ~pi647 & n23257;
  assign n23525 = n23523 & ~n23524;
  assign n23526 = ~n23521 & ~n23525;
  assign n23527 = ~n23520 & n23526;
  assign n23528 = pi787 & ~n23527;
  assign n23529 = ~n23516 & ~n23528;
  assign n23530 = pi644 & n23374;
  assign n23531 = ~pi644 & n23382;
  assign n23532 = pi790 & ~n23531;
  assign n23533 = ~n23530 & n23532;
  assign n23534 = n23529 & ~n23533;
  assign n23535 = ~n23385 & ~n23534;
  assign n23536 = ~po1038 & ~n23535;
  assign n23537 = ~pi175 & po1038;
  assign n23538 = ~pi832 & ~n23537;
  assign n23539 = ~n23536 & n23538;
  assign po332 = ~n23256 & ~n23539;
  assign n23541 = ~pi176 & ~n2934;
  assign n23542 = ~pi742 & n16510;
  assign n23543 = ~n23541 & ~n23542;
  assign n23544 = ~n17273 & ~n23543;
  assign n23545 = ~pi785 & ~n23544;
  assign n23546 = ~n17279 & ~n23543;
  assign n23547 = pi1155 & ~n23546;
  assign n23548 = ~n17282 & n23544;
  assign n23549 = ~pi1155 & ~n23548;
  assign n23550 = ~n23547 & ~n23549;
  assign n23551 = pi785 & ~n23550;
  assign n23552 = ~n23545 & ~n23551;
  assign n23553 = ~pi781 & ~n23552;
  assign n23554 = ~n17289 & n23552;
  assign n23555 = pi1154 & ~n23554;
  assign n23556 = ~n17292 & n23552;
  assign n23557 = ~pi1154 & ~n23556;
  assign n23558 = ~n23555 & ~n23557;
  assign n23559 = pi781 & ~n23558;
  assign n23560 = ~n23553 & ~n23559;
  assign n23561 = ~pi789 & ~n23560;
  assign n23562 = pi619 & n23560;
  assign n23563 = ~pi619 & n23541;
  assign n23564 = pi1159 & ~n23563;
  assign n23565 = ~n23562 & n23564;
  assign n23566 = ~pi619 & n23560;
  assign n23567 = pi619 & n23541;
  assign n23568 = ~pi1159 & ~n23567;
  assign n23569 = ~n23566 & n23568;
  assign n23570 = ~n23565 & ~n23569;
  assign n23571 = pi789 & ~n23570;
  assign n23572 = ~n23561 & ~n23571;
  assign n23573 = ~n17355 & n23572;
  assign n23574 = n17355 & n23541;
  assign n23575 = ~n23573 & ~n23574;
  assign n23576 = ~n16124 & ~n23575;
  assign n23577 = n16124 & n23541;
  assign n23578 = ~n23576 & ~n23577;
  assign n23579 = ~n19987 & n23578;
  assign n23580 = ~pi704 & n16742;
  assign n23581 = ~n23541 & ~n23580;
  assign n23582 = ~pi778 & n23581;
  assign n23583 = ~pi625 & n23580;
  assign n23584 = ~n23581 & ~n23583;
  assign n23585 = pi1153 & ~n23584;
  assign n23586 = ~pi1153 & ~n23541;
  assign n23587 = ~n23583 & n23586;
  assign n23588 = ~n23585 & ~n23587;
  assign n23589 = pi778 & ~n23588;
  assign n23590 = ~n23582 & ~n23589;
  assign n23591 = ~n17338 & n23590;
  assign n23592 = ~n17340 & n23591;
  assign n23593 = ~n17342 & n23592;
  assign n23594 = ~n17425 & n23593;
  assign n23595 = ~n17452 & n23594;
  assign n23596 = ~pi647 & n23595;
  assign n23597 = pi647 & n23541;
  assign n23598 = ~pi1157 & ~n23597;
  assign n23599 = ~n23596 & n23598;
  assign n23600 = ~pi647 & n23541;
  assign n23601 = pi647 & n23595;
  assign n23602 = pi1157 & ~n23601;
  assign n23603 = ~n23600 & n23602;
  assign n23604 = ~n23599 & ~n23603;
  assign n23605 = ~n17246 & ~n23604;
  assign n23606 = ~n23579 & ~n23605;
  assign n23607 = pi787 & ~n23606;
  assign n23608 = ~pi626 & ~n23572;
  assign n23609 = pi626 & ~n23541;
  assign n23610 = n17181 & ~n23609;
  assign n23611 = ~n23608 & n23610;
  assign n23612 = n17350 & n23593;
  assign n23613 = pi626 & ~n23572;
  assign n23614 = ~pi626 & ~n23541;
  assign n23615 = n17180 & ~n23614;
  assign n23616 = ~n23613 & n23615;
  assign n23617 = ~n23612 & ~n23616;
  assign n23618 = ~n23611 & n23617;
  assign n23619 = pi788 & ~n23618;
  assign n23620 = pi618 & n23591;
  assign n23621 = pi609 & n23590;
  assign n23622 = ~n16393 & ~n23581;
  assign n23623 = pi625 & n23622;
  assign n23624 = n23543 & ~n23622;
  assign n23625 = ~n23623 & ~n23624;
  assign n23626 = n23586 & ~n23625;
  assign n23627 = ~pi608 & ~n23585;
  assign n23628 = ~n23626 & n23627;
  assign n23629 = pi1153 & ~n23623;
  assign n23630 = n23543 & n23629;
  assign n23631 = ~n23587 & ~n23630;
  assign n23632 = pi608 & n23631;
  assign n23633 = ~n23628 & ~n23632;
  assign n23634 = pi778 & ~n23633;
  assign n23635 = ~pi778 & ~n23624;
  assign n23636 = ~n23634 & ~n23635;
  assign n23637 = ~pi609 & ~n23636;
  assign n23638 = ~pi1155 & ~n23637;
  assign n23639 = ~n23621 & n23638;
  assign n23640 = ~pi660 & ~n23547;
  assign n23641 = ~n23639 & n23640;
  assign n23642 = ~pi609 & n23590;
  assign n23643 = pi609 & ~n23636;
  assign n23644 = ~n23642 & ~n23643;
  assign n23645 = pi1155 & n23644;
  assign n23646 = ~n23549 & ~n23645;
  assign n23647 = pi660 & n23646;
  assign n23648 = ~n23641 & ~n23647;
  assign n23649 = pi785 & ~n23648;
  assign n23650 = ~pi785 & ~n23636;
  assign n23651 = ~n23649 & ~n23650;
  assign n23652 = ~pi618 & ~n23651;
  assign n23653 = ~pi1154 & ~n23652;
  assign n23654 = ~n23620 & n23653;
  assign n23655 = ~pi627 & ~n23555;
  assign n23656 = ~n23654 & n23655;
  assign n23657 = ~pi618 & n23591;
  assign n23658 = pi618 & ~n23651;
  assign n23659 = ~n23657 & ~n23658;
  assign n23660 = pi1154 & n23659;
  assign n23661 = ~n23557 & ~n23660;
  assign n23662 = pi627 & n23661;
  assign n23663 = ~n23656 & ~n23662;
  assign n23664 = pi781 & ~n23663;
  assign n23665 = ~pi781 & ~n23651;
  assign n23666 = ~n23664 & ~n23665;
  assign n23667 = ~pi619 & ~n23666;
  assign n23668 = pi619 & n23592;
  assign n23669 = ~pi1159 & ~n23668;
  assign n23670 = ~n23667 & n23669;
  assign n23671 = ~pi648 & ~n23670;
  assign n23672 = ~n23565 & n23671;
  assign n23673 = ~pi619 & n23592;
  assign n23674 = pi619 & ~n23666;
  assign n23675 = ~n23673 & ~n23674;
  assign n23676 = pi1159 & n23675;
  assign n23677 = ~n23569 & ~n23676;
  assign n23678 = pi648 & n23677;
  assign n23679 = ~n23672 & ~n23678;
  assign n23680 = pi789 & n23679;
  assign n23681 = ~pi789 & n23666;
  assign n23682 = n17356 & ~n23681;
  assign n23683 = ~n23680 & n23682;
  assign n23684 = ~n23619 & ~n23683;
  assign n23685 = n19788 & ~n23684;
  assign n23686 = n20275 & n23594;
  assign n23687 = n17449 & ~n23575;
  assign n23688 = ~pi629 & ~n23687;
  assign n23689 = ~n23686 & n23688;
  assign n23690 = n17448 & ~n23575;
  assign n23691 = n20281 & n23594;
  assign n23692 = pi629 & ~n23691;
  assign n23693 = ~n23690 & n23692;
  assign n23694 = ~n23689 & ~n23693;
  assign n23695 = pi792 & n23694;
  assign n23696 = n19637 & ~n23695;
  assign n23697 = ~n23685 & n23696;
  assign n23698 = ~n23607 & ~n23697;
  assign n23699 = pi644 & n23698;
  assign n23700 = ~pi787 & ~n23595;
  assign n23701 = pi787 & ~n23604;
  assign n23702 = ~n23700 & ~n23701;
  assign n23703 = ~pi644 & n23702;
  assign n23704 = pi715 & ~n23703;
  assign n23705 = ~n23699 & n23704;
  assign n23706 = ~n17247 & ~n23578;
  assign n23707 = n17247 & n23541;
  assign n23708 = ~n23706 & ~n23707;
  assign n23709 = pi644 & ~n23708;
  assign n23710 = ~pi644 & n23541;
  assign n23711 = ~pi715 & ~n23710;
  assign n23712 = ~n23709 & n23711;
  assign n23713 = pi1160 & ~n23712;
  assign n23714 = ~n23705 & n23713;
  assign n23715 = ~pi644 & ~n23708;
  assign n23716 = pi715 & ~n23715;
  assign n23717 = pi644 & n23541;
  assign n23718 = n23716 & ~n23717;
  assign n23719 = pi644 & n23702;
  assign n23720 = ~pi644 & n23698;
  assign n23721 = ~pi715 & ~n23720;
  assign n23722 = ~n23719 & n23721;
  assign n23723 = ~pi1160 & ~n23722;
  assign n23724 = ~n23718 & n23723;
  assign n23725 = ~n23714 & ~n23724;
  assign n23726 = pi790 & ~n23725;
  assign n23727 = ~pi790 & n23698;
  assign n23728 = pi832 & ~n23727;
  assign n23729 = ~n23726 & n23728;
  assign n23730 = ~pi176 & ~n16527;
  assign n23731 = n17451 & ~n23730;
  assign n23732 = n17159 & ~n23730;
  assign n23733 = n16593 & ~n23730;
  assign n23734 = ~n16744 & n19843;
  assign n23735 = pi176 & ~n23734;
  assign n23736 = ~pi38 & n17592;
  assign n23737 = ~n19410 & ~n23736;
  assign n23738 = ~pi176 & n23737;
  assign n23739 = ~pi704 & ~n23738;
  assign n23740 = ~pi176 & ~n16526;
  assign n23741 = pi704 & n23740;
  assign n23742 = n10020 & ~n23741;
  assign n23743 = ~n23739 & n23742;
  assign n23744 = ~n23735 & ~n23743;
  assign n23745 = ~pi778 & ~n23744;
  assign n23746 = pi625 & n23744;
  assign n23747 = pi1153 & ~n23746;
  assign n23748 = ~pi625 & n23730;
  assign n23749 = n23747 & ~n23748;
  assign n23750 = ~pi625 & n23744;
  assign n23751 = ~pi1153 & ~n23750;
  assign n23752 = pi625 & n23730;
  assign n23753 = n23751 & ~n23752;
  assign n23754 = ~n23749 & ~n23753;
  assign n23755 = pi778 & ~n23754;
  assign n23756 = ~n23745 & ~n23755;
  assign n23757 = ~n16593 & ~n23756;
  assign n23758 = ~n23733 & ~n23757;
  assign n23759 = ~n16589 & n23758;
  assign n23760 = n16589 & n23730;
  assign n23761 = ~n23759 & ~n23760;
  assign n23762 = ~n17159 & n23761;
  assign n23763 = ~n23732 & ~n23762;
  assign n23764 = ~n17183 & n23763;
  assign n23765 = n17183 & n23730;
  assign n23766 = ~n23764 & ~n23765;
  assign n23767 = ~n17451 & n23766;
  assign n23768 = ~n23731 & ~n23767;
  assign n23769 = ~n18767 & n23768;
  assign n23770 = n18767 & n23730;
  assign n23771 = ~n23769 & ~n23770;
  assign n23772 = ~pi644 & ~n23771;
  assign n23773 = pi715 & ~n23772;
  assign n23774 = n17247 & ~n23730;
  assign n23775 = pi176 & ~n10020;
  assign n23776 = ~pi176 & n18808;
  assign n23777 = ~n18802 & ~n18803;
  assign n23778 = pi176 & n23777;
  assign n23779 = ~n23776 & ~n23778;
  assign n23780 = ~pi742 & ~n23779;
  assign n23781 = pi742 & ~n23740;
  assign n23782 = ~n23780 & ~n23781;
  assign n23783 = n10020 & ~n23782;
  assign n23784 = ~n23775 & ~n23783;
  assign n23785 = ~n16521 & ~n23784;
  assign n23786 = n16521 & ~n23730;
  assign n23787 = ~n23785 & ~n23786;
  assign n23788 = ~pi785 & ~n23787;
  assign n23789 = ~n16532 & ~n23730;
  assign n23790 = pi609 & n23785;
  assign n23791 = ~n23789 & ~n23790;
  assign n23792 = pi1155 & ~n23791;
  assign n23793 = ~n16537 & ~n23730;
  assign n23794 = ~pi609 & n23785;
  assign n23795 = ~n23793 & ~n23794;
  assign n23796 = ~pi1155 & ~n23795;
  assign n23797 = ~n23792 & ~n23796;
  assign n23798 = pi785 & ~n23797;
  assign n23799 = ~n23788 & ~n23798;
  assign n23800 = ~pi781 & ~n23799;
  assign n23801 = pi618 & n23799;
  assign n23802 = ~pi618 & n23730;
  assign n23803 = pi1154 & ~n23802;
  assign n23804 = ~n23801 & n23803;
  assign n23805 = ~pi618 & n23799;
  assign n23806 = pi618 & n23730;
  assign n23807 = ~pi1154 & ~n23806;
  assign n23808 = ~n23805 & n23807;
  assign n23809 = ~n23804 & ~n23808;
  assign n23810 = pi781 & ~n23809;
  assign n23811 = ~n23800 & ~n23810;
  assign n23812 = ~pi789 & ~n23811;
  assign n23813 = pi619 & n23811;
  assign n23814 = ~pi619 & n23730;
  assign n23815 = pi1159 & ~n23814;
  assign n23816 = ~n23813 & n23815;
  assign n23817 = ~pi619 & n23811;
  assign n23818 = pi619 & n23730;
  assign n23819 = ~pi1159 & ~n23818;
  assign n23820 = ~n23817 & n23819;
  assign n23821 = ~n23816 & ~n23820;
  assign n23822 = pi789 & ~n23821;
  assign n23823 = ~n23812 & ~n23822;
  assign n23824 = ~n17355 & n23823;
  assign n23825 = n17355 & n23730;
  assign n23826 = ~n23824 & ~n23825;
  assign n23827 = ~n16124 & ~n23826;
  assign n23828 = n16124 & n23730;
  assign n23829 = ~n23827 & ~n23828;
  assign n23830 = ~n17247 & n23829;
  assign n23831 = ~n23774 & ~n23830;
  assign n23832 = pi644 & n23831;
  assign n23833 = ~pi644 & n23730;
  assign n23834 = ~pi715 & ~n23833;
  assign n23835 = ~n23832 & n23834;
  assign n23836 = pi1160 & ~n23835;
  assign n23837 = ~n23773 & n23836;
  assign n23838 = pi644 & ~n23771;
  assign n23839 = ~pi715 & ~n23838;
  assign n23840 = ~pi644 & n23831;
  assign n23841 = pi644 & n23730;
  assign n23842 = ~n23840 & ~n23841;
  assign n23843 = pi715 & n23842;
  assign n23844 = ~pi1160 & ~n23843;
  assign n23845 = ~n23839 & n23844;
  assign n23846 = ~n23837 & ~n23845;
  assign n23847 = pi790 & ~n23846;
  assign n23848 = ~pi647 & n23768;
  assign n23849 = pi647 & n23730;
  assign n23850 = n17245 & ~n23849;
  assign n23851 = ~n23848 & n23850;
  assign n23852 = ~n19987 & n23829;
  assign n23853 = pi647 & n23768;
  assign n23854 = n17244 & ~n23853;
  assign n23855 = ~pi647 & n23730;
  assign n23856 = n23854 & ~n23855;
  assign n23857 = ~n23852 & ~n23856;
  assign n23858 = ~n23851 & n23857;
  assign n23859 = pi787 & ~n23858;
  assign n23860 = ~n19999 & n23826;
  assign n23861 = pi628 & ~n23766;
  assign n23862 = n16121 & ~n23861;
  assign n23863 = ~pi628 & n23730;
  assign n23864 = n23862 & ~n23863;
  assign n23865 = ~pi628 & ~n23766;
  assign n23866 = pi628 & n23730;
  assign n23867 = n16122 & ~n23866;
  assign n23868 = ~n23865 & n23867;
  assign n23869 = ~n23864 & ~n23868;
  assign n23870 = ~n23860 & n23869;
  assign n23871 = ~n19788 & n23870;
  assign n23872 = pi792 & ~n23870;
  assign n23873 = ~pi626 & ~n23823;
  assign n23874 = pi626 & ~n23730;
  assign n23875 = n17181 & ~n23874;
  assign n23876 = ~n23873 & n23875;
  assign n23877 = n17350 & n23763;
  assign n23878 = pi626 & ~n23823;
  assign n23879 = ~pi626 & ~n23730;
  assign n23880 = n17180 & ~n23879;
  assign n23881 = ~n23878 & n23880;
  assign n23882 = ~n23877 & ~n23881;
  assign n23883 = ~n23876 & n23882;
  assign n23884 = pi788 & ~n23883;
  assign n23885 = pi618 & n23758;
  assign n23886 = pi609 & n23756;
  assign n23887 = pi625 & n23784;
  assign n23888 = pi704 & n23782;
  assign n23889 = ~n18929 & ~n18932;
  assign n23890 = pi176 & ~n23889;
  assign n23891 = ~pi176 & n18939;
  assign n23892 = ~n23890 & ~n23891;
  assign n23893 = pi742 & n23892;
  assign n23894 = ~pi176 & ~n18914;
  assign n23895 = pi176 & n18922;
  assign n23896 = ~pi742 & ~n23895;
  assign n23897 = ~n23894 & n23896;
  assign n23898 = ~pi704 & ~n23897;
  assign n23899 = ~n23893 & n23898;
  assign n23900 = ~n23888 & ~n23899;
  assign n23901 = n10020 & n23900;
  assign n23902 = ~n23775 & ~n23901;
  assign n23903 = ~pi625 & n23902;
  assign n23904 = ~pi1153 & ~n23903;
  assign n23905 = ~n23887 & n23904;
  assign n23906 = ~pi608 & ~n23749;
  assign n23907 = ~n23905 & n23906;
  assign n23908 = ~pi625 & n23784;
  assign n23909 = pi625 & n23902;
  assign n23910 = ~n23908 & ~n23909;
  assign n23911 = pi1153 & n23910;
  assign n23912 = ~n23753 & ~n23911;
  assign n23913 = pi608 & n23912;
  assign n23914 = ~n23907 & ~n23913;
  assign n23915 = pi778 & ~n23914;
  assign n23916 = ~pi778 & n23902;
  assign n23917 = ~n23915 & ~n23916;
  assign n23918 = ~pi609 & ~n23917;
  assign n23919 = ~pi1155 & ~n23918;
  assign n23920 = ~n23886 & n23919;
  assign n23921 = ~pi660 & ~n23792;
  assign n23922 = ~n23920 & n23921;
  assign n23923 = ~pi609 & n23756;
  assign n23924 = pi609 & ~n23917;
  assign n23925 = ~n23923 & ~n23924;
  assign n23926 = pi1155 & n23925;
  assign n23927 = ~n23796 & ~n23926;
  assign n23928 = pi660 & n23927;
  assign n23929 = ~n23922 & ~n23928;
  assign n23930 = pi785 & ~n23929;
  assign n23931 = ~pi785 & ~n23917;
  assign n23932 = ~n23930 & ~n23931;
  assign n23933 = ~pi618 & ~n23932;
  assign n23934 = ~pi1154 & ~n23933;
  assign n23935 = ~n23885 & n23934;
  assign n23936 = ~pi627 & ~n23804;
  assign n23937 = ~n23935 & n23936;
  assign n23938 = ~pi618 & n23758;
  assign n23939 = pi618 & ~n23932;
  assign n23940 = ~n23938 & ~n23939;
  assign n23941 = pi1154 & n23940;
  assign n23942 = ~n23808 & ~n23941;
  assign n23943 = pi627 & n23942;
  assign n23944 = ~n23937 & ~n23943;
  assign n23945 = pi781 & ~n23944;
  assign n23946 = ~pi781 & ~n23932;
  assign n23947 = ~n23945 & ~n23946;
  assign n23948 = ~pi619 & ~n23947;
  assign n23949 = pi619 & ~n23761;
  assign n23950 = ~pi1159 & ~n23949;
  assign n23951 = ~n23948 & n23950;
  assign n23952 = ~pi648 & ~n23951;
  assign n23953 = ~n23816 & n23952;
  assign n23954 = ~pi619 & ~n23761;
  assign n23955 = pi619 & ~n23947;
  assign n23956 = ~n23954 & ~n23955;
  assign n23957 = pi1159 & n23956;
  assign n23958 = ~n23820 & ~n23957;
  assign n23959 = pi648 & n23958;
  assign n23960 = ~n23953 & ~n23959;
  assign n23961 = pi789 & n23960;
  assign n23962 = ~pi789 & n23947;
  assign n23963 = n17356 & ~n23962;
  assign n23964 = ~n23961 & n23963;
  assign n23965 = ~n23884 & ~n23964;
  assign n23966 = ~n23872 & ~n23965;
  assign n23967 = ~n23871 & ~n23966;
  assign n23968 = n19637 & n23967;
  assign n23969 = ~n23859 & ~n23968;
  assign n23970 = pi644 & n23836;
  assign n23971 = ~pi644 & n23844;
  assign n23972 = pi790 & ~n23971;
  assign n23973 = ~n23970 & n23972;
  assign n23974 = n23969 & ~n23973;
  assign n23975 = ~n23847 & ~n23974;
  assign n23976 = ~po1038 & ~n23975;
  assign n23977 = ~pi176 & po1038;
  assign n23978 = ~pi832 & ~n23977;
  assign n23979 = ~n23976 & n23978;
  assign po333 = ~n23729 & ~n23979;
  assign n23981 = pi177 & ~n10020;
  assign n23982 = ~pi757 & ~n18808;
  assign n23983 = ~n21046 & ~n23982;
  assign n23984 = ~pi177 & ~n23983;
  assign n23985 = ~pi177 & ~n18802;
  assign n23986 = ~pi757 & ~n23985;
  assign n23987 = ~n23777 & n23986;
  assign n23988 = ~n23984 & ~n23987;
  assign n23989 = n10020 & n23988;
  assign n23990 = ~n23981 & ~n23989;
  assign n23991 = ~n16521 & ~n23990;
  assign n23992 = ~pi177 & ~n16527;
  assign n23993 = n16521 & ~n23992;
  assign n23994 = ~n23991 & ~n23993;
  assign n23995 = ~pi785 & ~n23994;
  assign n23996 = ~n16532 & ~n23992;
  assign n23997 = pi609 & n23991;
  assign n23998 = ~n23996 & ~n23997;
  assign n23999 = pi1155 & ~n23998;
  assign n24000 = ~n16537 & ~n23992;
  assign n24001 = ~pi609 & n23991;
  assign n24002 = ~n24000 & ~n24001;
  assign n24003 = ~pi1155 & ~n24002;
  assign n24004 = ~n23999 & ~n24003;
  assign n24005 = pi785 & ~n24004;
  assign n24006 = ~n23995 & ~n24005;
  assign n24007 = ~pi781 & ~n24006;
  assign n24008 = pi618 & n24006;
  assign n24009 = ~pi618 & n23992;
  assign n24010 = pi1154 & ~n24009;
  assign n24011 = ~n24008 & n24010;
  assign n24012 = ~pi618 & n24006;
  assign n24013 = pi618 & n23992;
  assign n24014 = ~pi1154 & ~n24013;
  assign n24015 = ~n24012 & n24014;
  assign n24016 = ~n24011 & ~n24015;
  assign n24017 = pi781 & ~n24016;
  assign n24018 = ~n24007 & ~n24017;
  assign n24019 = ~pi789 & ~n24018;
  assign n24020 = pi619 & n24018;
  assign n24021 = ~pi619 & n23992;
  assign n24022 = pi1159 & ~n24021;
  assign n24023 = ~n24020 & n24022;
  assign n24024 = ~pi619 & n24018;
  assign n24025 = pi619 & n23992;
  assign n24026 = ~pi1159 & ~n24025;
  assign n24027 = ~n24024 & n24026;
  assign n24028 = ~n24023 & ~n24027;
  assign n24029 = pi789 & ~n24028;
  assign n24030 = ~n24019 & ~n24029;
  assign n24031 = ~n17355 & n24030;
  assign n24032 = n17355 & n23992;
  assign n24033 = ~n24031 & ~n24032;
  assign n24034 = ~n16124 & ~n24033;
  assign n24035 = n16124 & n23992;
  assign n24036 = ~n24034 & ~n24035;
  assign n24037 = pi647 & ~n24036;
  assign n24038 = pi628 & ~n24033;
  assign n24039 = n16593 & ~n23992;
  assign n24040 = pi177 & n17589;
  assign n24041 = ~pi177 & n17592;
  assign n24042 = ~pi38 & ~n24041;
  assign n24043 = ~n24040 & n24042;
  assign n24044 = ~pi177 & ~n16508;
  assign n24045 = n16744 & ~n24044;
  assign n24046 = ~pi686 & ~n24045;
  assign n24047 = ~n24043 & n24046;
  assign n24048 = ~pi177 & ~n16526;
  assign n24049 = pi686 & n24048;
  assign n24050 = ~n24047 & ~n24049;
  assign n24051 = n10020 & n24050;
  assign n24052 = ~n23981 & ~n24051;
  assign n24053 = ~pi778 & ~n24052;
  assign n24054 = pi625 & n24052;
  assign n24055 = pi1153 & ~n24054;
  assign n24056 = ~pi625 & n23992;
  assign n24057 = n24055 & ~n24056;
  assign n24058 = ~pi625 & n24052;
  assign n24059 = ~pi1153 & ~n24058;
  assign n24060 = pi625 & n23992;
  assign n24061 = n24059 & ~n24060;
  assign n24062 = ~n24057 & ~n24061;
  assign n24063 = pi778 & ~n24062;
  assign n24064 = ~n24053 & ~n24063;
  assign n24065 = ~n16593 & ~n24064;
  assign n24066 = ~n24039 & ~n24065;
  assign n24067 = ~n16589 & n24066;
  assign n24068 = n16589 & n23992;
  assign n24069 = ~n24067 & ~n24068;
  assign n24070 = pi619 & ~n24069;
  assign n24071 = pi618 & n24066;
  assign n24072 = pi609 & n24064;
  assign n24073 = pi625 & n23990;
  assign n24074 = pi686 & ~n23988;
  assign n24075 = pi177 & n18928;
  assign n24076 = ~pi177 & n18937;
  assign n24077 = ~pi38 & ~n24076;
  assign n24078 = ~n24075 & n24077;
  assign n24079 = n17627 & ~n24044;
  assign n24080 = pi757 & ~n24079;
  assign n24081 = ~n24078 & n24080;
  assign n24082 = ~n18908 & ~n18912;
  assign n24083 = ~pi177 & ~n24082;
  assign n24084 = pi177 & n18918;
  assign n24085 = ~pi38 & ~n24084;
  assign n24086 = ~n24083 & n24085;
  assign n24087 = n18921 & ~n24044;
  assign n24088 = ~pi757 & ~n24087;
  assign n24089 = ~n24086 & n24088;
  assign n24090 = ~n24081 & ~n24089;
  assign n24091 = ~pi686 & ~n24090;
  assign n24092 = ~n24074 & ~n24091;
  assign n24093 = n10020 & n24092;
  assign n24094 = ~n23981 & ~n24093;
  assign n24095 = ~pi625 & n24094;
  assign n24096 = ~pi1153 & ~n24095;
  assign n24097 = ~n24073 & n24096;
  assign n24098 = ~pi608 & ~n24057;
  assign n24099 = ~n24097 & n24098;
  assign n24100 = ~pi625 & n23990;
  assign n24101 = pi625 & n24094;
  assign n24102 = ~n24100 & ~n24101;
  assign n24103 = pi1153 & n24102;
  assign n24104 = ~n24061 & ~n24103;
  assign n24105 = pi608 & n24104;
  assign n24106 = ~n24099 & ~n24105;
  assign n24107 = pi778 & ~n24106;
  assign n24108 = ~pi778 & n24094;
  assign n24109 = ~n24107 & ~n24108;
  assign n24110 = ~pi609 & ~n24109;
  assign n24111 = ~pi1155 & ~n24110;
  assign n24112 = ~n24072 & n24111;
  assign n24113 = ~pi660 & ~n23999;
  assign n24114 = ~n24112 & n24113;
  assign n24115 = ~pi609 & n24064;
  assign n24116 = pi609 & ~n24109;
  assign n24117 = ~n24115 & ~n24116;
  assign n24118 = pi1155 & n24117;
  assign n24119 = ~n24003 & ~n24118;
  assign n24120 = pi660 & n24119;
  assign n24121 = ~n24114 & ~n24120;
  assign n24122 = pi785 & ~n24121;
  assign n24123 = ~pi785 & ~n24109;
  assign n24124 = ~n24122 & ~n24123;
  assign n24125 = ~pi618 & ~n24124;
  assign n24126 = ~pi1154 & ~n24125;
  assign n24127 = ~n24071 & n24126;
  assign n24128 = ~pi627 & ~n24011;
  assign n24129 = ~n24127 & n24128;
  assign n24130 = ~pi618 & n24066;
  assign n24131 = pi618 & ~n24124;
  assign n24132 = ~n24130 & ~n24131;
  assign n24133 = pi1154 & n24132;
  assign n24134 = ~n24015 & ~n24133;
  assign n24135 = pi627 & n24134;
  assign n24136 = ~n24129 & ~n24135;
  assign n24137 = pi781 & ~n24136;
  assign n24138 = ~pi781 & ~n24124;
  assign n24139 = ~n24137 & ~n24138;
  assign n24140 = ~pi619 & ~n24139;
  assign n24141 = ~pi1159 & ~n24140;
  assign n24142 = ~n24070 & n24141;
  assign n24143 = ~pi648 & ~n24023;
  assign n24144 = ~n24142 & n24143;
  assign n24145 = ~pi619 & ~n24069;
  assign n24146 = pi619 & ~n24139;
  assign n24147 = ~n24145 & ~n24146;
  assign n24148 = pi1159 & n24147;
  assign n24149 = ~n24027 & ~n24148;
  assign n24150 = pi648 & n24149;
  assign n24151 = ~n24144 & ~n24150;
  assign n24152 = pi789 & ~n24151;
  assign n24153 = ~pi789 & ~n24139;
  assign n24154 = ~n24152 & ~n24153;
  assign n24155 = ~pi788 & n24154;
  assign n24156 = pi626 & n24154;
  assign n24157 = n17159 & ~n23992;
  assign n24158 = ~n17159 & n24069;
  assign n24159 = ~n24157 & ~n24158;
  assign n24160 = ~pi626 & ~n24159;
  assign n24161 = pi641 & ~n24160;
  assign n24162 = ~n24156 & n24161;
  assign n24163 = pi626 & ~n24030;
  assign n24164 = ~pi626 & ~n23992;
  assign n24165 = ~pi641 & ~n24164;
  assign n24166 = ~n24163 & n24165;
  assign n24167 = pi1158 & ~n24166;
  assign n24168 = ~n24162 & n24167;
  assign n24169 = pi626 & ~n23992;
  assign n24170 = ~pi626 & ~n24030;
  assign n24171 = pi641 & ~n24170;
  assign n24172 = ~n24169 & n24171;
  assign n24173 = pi626 & ~n24159;
  assign n24174 = ~pi626 & n24154;
  assign n24175 = ~pi641 & ~n24174;
  assign n24176 = ~n24173 & n24175;
  assign n24177 = ~pi1158 & ~n24176;
  assign n24178 = ~n24172 & n24177;
  assign n24179 = ~n24168 & ~n24178;
  assign n24180 = pi788 & ~n24179;
  assign n24181 = ~n24155 & ~n24180;
  assign n24182 = ~pi628 & n24181;
  assign n24183 = ~pi1156 & ~n24182;
  assign n24184 = ~n24038 & n24183;
  assign n24185 = ~n17183 & n24159;
  assign n24186 = n17183 & n23992;
  assign n24187 = ~n24185 & ~n24186;
  assign n24188 = pi628 & ~n24187;
  assign n24189 = pi1156 & ~n24188;
  assign n24190 = ~pi628 & n23992;
  assign n24191 = n24189 & ~n24190;
  assign n24192 = ~pi629 & ~n24191;
  assign n24193 = ~n24184 & n24192;
  assign n24194 = ~pi628 & ~n24187;
  assign n24195 = pi628 & n23992;
  assign n24196 = ~pi1156 & ~n24195;
  assign n24197 = ~n24194 & n24196;
  assign n24198 = ~pi628 & ~n24033;
  assign n24199 = pi628 & n24181;
  assign n24200 = ~n24198 & ~n24199;
  assign n24201 = pi1156 & n24200;
  assign n24202 = ~n24197 & ~n24201;
  assign n24203 = pi629 & n24202;
  assign n24204 = ~n24193 & ~n24203;
  assign n24205 = pi792 & ~n24204;
  assign n24206 = ~pi792 & n24181;
  assign n24207 = ~n24205 & ~n24206;
  assign n24208 = ~pi647 & ~n24207;
  assign n24209 = ~pi1157 & ~n24208;
  assign n24210 = ~n24037 & n24209;
  assign n24211 = ~pi792 & n24187;
  assign n24212 = ~n24191 & ~n24197;
  assign n24213 = pi792 & ~n24212;
  assign n24214 = ~n24211 & ~n24213;
  assign n24215 = pi647 & n24214;
  assign n24216 = pi1157 & ~n24215;
  assign n24217 = ~pi647 & n23992;
  assign n24218 = n24216 & ~n24217;
  assign n24219 = ~pi630 & ~n24218;
  assign n24220 = ~n24210 & n24219;
  assign n24221 = ~pi647 & n24214;
  assign n24222 = pi647 & n23992;
  assign n24223 = ~pi1157 & ~n24222;
  assign n24224 = ~n24221 & n24223;
  assign n24225 = ~pi647 & ~n24036;
  assign n24226 = pi647 & ~n24207;
  assign n24227 = ~n24225 & ~n24226;
  assign n24228 = pi1157 & n24227;
  assign n24229 = ~n24224 & ~n24228;
  assign n24230 = pi630 & n24229;
  assign n24231 = ~n24220 & ~n24230;
  assign n24232 = pi787 & ~n24231;
  assign n24233 = ~pi787 & ~n24207;
  assign n24234 = ~n24232 & ~n24233;
  assign n24235 = ~pi790 & n24234;
  assign n24236 = pi644 & ~n24234;
  assign n24237 = ~pi787 & ~n24214;
  assign n24238 = ~n24218 & ~n24224;
  assign n24239 = pi787 & ~n24238;
  assign n24240 = ~n24237 & ~n24239;
  assign n24241 = ~pi644 & n24240;
  assign n24242 = pi715 & ~n24241;
  assign n24243 = ~n24236 & n24242;
  assign n24244 = ~pi644 & n23992;
  assign n24245 = n17247 & ~n23992;
  assign n24246 = ~n17247 & n24036;
  assign n24247 = ~n24245 & ~n24246;
  assign n24248 = pi644 & n24247;
  assign n24249 = ~pi715 & ~n24248;
  assign n24250 = ~n24244 & n24249;
  assign n24251 = ~n24243 & ~n24250;
  assign n24252 = pi1160 & n24251;
  assign n24253 = ~pi644 & n24247;
  assign n24254 = pi715 & ~n24253;
  assign n24255 = pi644 & n23992;
  assign n24256 = n24254 & ~n24255;
  assign n24257 = pi644 & n24240;
  assign n24258 = ~pi644 & ~n24234;
  assign n24259 = ~pi715 & ~n24258;
  assign n24260 = ~n24257 & n24259;
  assign n24261 = ~n24256 & ~n24260;
  assign n24262 = ~pi1160 & n24261;
  assign n24263 = ~n24252 & ~n24262;
  assign n24264 = pi790 & n24263;
  assign n24265 = ~n24235 & ~n24264;
  assign n24266 = ~po1038 & n24265;
  assign n24267 = ~pi177 & po1038;
  assign n24268 = ~pi832 & ~n24267;
  assign n24269 = ~n24266 & n24268;
  assign n24270 = ~pi177 & ~n2934;
  assign n24271 = ~pi757 & n16510;
  assign n24272 = ~n24270 & ~n24271;
  assign n24273 = ~n17273 & ~n24272;
  assign n24274 = ~pi785 & ~n24273;
  assign n24275 = ~n17279 & ~n24272;
  assign n24276 = pi1155 & ~n24275;
  assign n24277 = ~n17282 & n24273;
  assign n24278 = ~pi1155 & ~n24277;
  assign n24279 = ~n24276 & ~n24278;
  assign n24280 = pi785 & ~n24279;
  assign n24281 = ~n24274 & ~n24280;
  assign n24282 = ~pi781 & ~n24281;
  assign n24283 = ~n17289 & n24281;
  assign n24284 = pi1154 & ~n24283;
  assign n24285 = ~n17292 & n24281;
  assign n24286 = ~pi1154 & ~n24285;
  assign n24287 = ~n24284 & ~n24286;
  assign n24288 = pi781 & ~n24287;
  assign n24289 = ~n24282 & ~n24288;
  assign n24290 = ~pi789 & ~n24289;
  assign n24291 = pi619 & n24289;
  assign n24292 = ~pi619 & n24270;
  assign n24293 = pi1159 & ~n24292;
  assign n24294 = ~n24291 & n24293;
  assign n24295 = ~pi619 & n24289;
  assign n24296 = pi619 & n24270;
  assign n24297 = ~pi1159 & ~n24296;
  assign n24298 = ~n24295 & n24297;
  assign n24299 = ~n24294 & ~n24298;
  assign n24300 = pi789 & ~n24299;
  assign n24301 = ~n24290 & ~n24300;
  assign n24302 = ~n17355 & n24301;
  assign n24303 = n17355 & n24270;
  assign n24304 = ~n24302 & ~n24303;
  assign n24305 = ~n16124 & ~n24304;
  assign n24306 = n16124 & n24270;
  assign n24307 = ~n24305 & ~n24306;
  assign n24308 = ~n19987 & n24307;
  assign n24309 = ~pi686 & n16742;
  assign n24310 = ~n24270 & ~n24309;
  assign n24311 = ~pi778 & n24310;
  assign n24312 = ~pi625 & n24309;
  assign n24313 = ~n24310 & ~n24312;
  assign n24314 = pi1153 & ~n24313;
  assign n24315 = ~pi1153 & ~n24270;
  assign n24316 = ~n24312 & n24315;
  assign n24317 = ~n24314 & ~n24316;
  assign n24318 = pi778 & ~n24317;
  assign n24319 = ~n24311 & ~n24318;
  assign n24320 = ~n17338 & n24319;
  assign n24321 = ~n17340 & n24320;
  assign n24322 = ~n17342 & n24321;
  assign n24323 = ~n17425 & n24322;
  assign n24324 = ~n17452 & n24323;
  assign n24325 = ~pi647 & n24324;
  assign n24326 = pi647 & n24270;
  assign n24327 = ~pi1157 & ~n24326;
  assign n24328 = ~n24325 & n24327;
  assign n24329 = ~pi647 & n24270;
  assign n24330 = pi647 & n24324;
  assign n24331 = pi1157 & ~n24330;
  assign n24332 = ~n24329 & n24331;
  assign n24333 = ~n24328 & ~n24332;
  assign n24334 = ~n17246 & ~n24333;
  assign n24335 = ~n24308 & ~n24334;
  assign n24336 = pi787 & ~n24335;
  assign n24337 = ~pi626 & ~n24301;
  assign n24338 = pi626 & ~n24270;
  assign n24339 = n17181 & ~n24338;
  assign n24340 = ~n24337 & n24339;
  assign n24341 = n17350 & n24322;
  assign n24342 = pi626 & ~n24301;
  assign n24343 = ~pi626 & ~n24270;
  assign n24344 = n17180 & ~n24343;
  assign n24345 = ~n24342 & n24344;
  assign n24346 = ~n24341 & ~n24345;
  assign n24347 = ~n24340 & n24346;
  assign n24348 = pi788 & ~n24347;
  assign n24349 = pi618 & n24320;
  assign n24350 = pi609 & n24319;
  assign n24351 = ~n16393 & ~n24310;
  assign n24352 = pi625 & n24351;
  assign n24353 = n24272 & ~n24351;
  assign n24354 = ~n24352 & ~n24353;
  assign n24355 = n24315 & ~n24354;
  assign n24356 = ~pi608 & ~n24314;
  assign n24357 = ~n24355 & n24356;
  assign n24358 = pi1153 & ~n24352;
  assign n24359 = n24272 & n24358;
  assign n24360 = ~n24316 & ~n24359;
  assign n24361 = pi608 & n24360;
  assign n24362 = ~n24357 & ~n24361;
  assign n24363 = pi778 & ~n24362;
  assign n24364 = ~pi778 & ~n24353;
  assign n24365 = ~n24363 & ~n24364;
  assign n24366 = ~pi609 & ~n24365;
  assign n24367 = ~pi1155 & ~n24366;
  assign n24368 = ~n24350 & n24367;
  assign n24369 = ~pi660 & ~n24276;
  assign n24370 = ~n24368 & n24369;
  assign n24371 = ~pi609 & n24319;
  assign n24372 = pi609 & ~n24365;
  assign n24373 = ~n24371 & ~n24372;
  assign n24374 = pi1155 & n24373;
  assign n24375 = ~n24278 & ~n24374;
  assign n24376 = pi660 & n24375;
  assign n24377 = ~n24370 & ~n24376;
  assign n24378 = pi785 & ~n24377;
  assign n24379 = ~pi785 & ~n24365;
  assign n24380 = ~n24378 & ~n24379;
  assign n24381 = ~pi618 & ~n24380;
  assign n24382 = ~pi1154 & ~n24381;
  assign n24383 = ~n24349 & n24382;
  assign n24384 = ~pi627 & ~n24284;
  assign n24385 = ~n24383 & n24384;
  assign n24386 = ~pi618 & n24320;
  assign n24387 = pi618 & ~n24380;
  assign n24388 = ~n24386 & ~n24387;
  assign n24389 = pi1154 & n24388;
  assign n24390 = ~n24286 & ~n24389;
  assign n24391 = pi627 & n24390;
  assign n24392 = ~n24385 & ~n24391;
  assign n24393 = pi781 & ~n24392;
  assign n24394 = ~pi781 & ~n24380;
  assign n24395 = ~n24393 & ~n24394;
  assign n24396 = ~pi619 & ~n24395;
  assign n24397 = pi619 & n24321;
  assign n24398 = ~pi1159 & ~n24397;
  assign n24399 = ~n24396 & n24398;
  assign n24400 = ~pi648 & ~n24399;
  assign n24401 = ~n24294 & n24400;
  assign n24402 = ~pi619 & n24321;
  assign n24403 = pi619 & ~n24395;
  assign n24404 = ~n24402 & ~n24403;
  assign n24405 = pi1159 & n24404;
  assign n24406 = ~n24298 & ~n24405;
  assign n24407 = pi648 & n24406;
  assign n24408 = ~n24401 & ~n24407;
  assign n24409 = pi789 & n24408;
  assign n24410 = ~pi789 & n24395;
  assign n24411 = n17356 & ~n24410;
  assign n24412 = ~n24409 & n24411;
  assign n24413 = ~n24348 & ~n24412;
  assign n24414 = n19788 & ~n24413;
  assign n24415 = n20275 & n24323;
  assign n24416 = n17449 & ~n24304;
  assign n24417 = ~pi629 & ~n24416;
  assign n24418 = ~n24415 & n24417;
  assign n24419 = n17448 & ~n24304;
  assign n24420 = n20281 & n24323;
  assign n24421 = pi629 & ~n24420;
  assign n24422 = ~n24419 & n24421;
  assign n24423 = ~n24418 & ~n24422;
  assign n24424 = pi792 & n24423;
  assign n24425 = n19637 & ~n24424;
  assign n24426 = ~n24414 & n24425;
  assign n24427 = ~n24336 & ~n24426;
  assign n24428 = pi644 & n24427;
  assign n24429 = ~pi787 & ~n24324;
  assign n24430 = pi787 & ~n24333;
  assign n24431 = ~n24429 & ~n24430;
  assign n24432 = ~pi644 & n24431;
  assign n24433 = pi715 & ~n24432;
  assign n24434 = ~n24428 & n24433;
  assign n24435 = ~n17247 & ~n24307;
  assign n24436 = n17247 & n24270;
  assign n24437 = ~n24435 & ~n24436;
  assign n24438 = pi644 & ~n24437;
  assign n24439 = ~pi644 & n24270;
  assign n24440 = ~pi715 & ~n24439;
  assign n24441 = ~n24438 & n24440;
  assign n24442 = pi1160 & ~n24441;
  assign n24443 = ~n24434 & n24442;
  assign n24444 = ~pi644 & ~n24437;
  assign n24445 = pi715 & ~n24444;
  assign n24446 = pi644 & n24270;
  assign n24447 = n24445 & ~n24446;
  assign n24448 = pi644 & n24431;
  assign n24449 = ~pi644 & n24427;
  assign n24450 = ~pi715 & ~n24449;
  assign n24451 = ~n24448 & n24450;
  assign n24452 = ~pi1160 & ~n24451;
  assign n24453 = ~n24447 & n24452;
  assign n24454 = ~n24443 & ~n24453;
  assign n24455 = pi790 & ~n24454;
  assign n24456 = ~pi790 & n24427;
  assign n24457 = pi832 & ~n24456;
  assign n24458 = ~n24455 & n24457;
  assign po334 = ~n24269 & ~n24458;
  assign n24460 = ~pi178 & ~n2934;
  assign n24461 = ~pi760 & n16510;
  assign n24462 = ~n24460 & ~n24461;
  assign n24463 = ~n17273 & ~n24462;
  assign n24464 = ~pi785 & ~n24463;
  assign n24465 = n16537 & n24461;
  assign n24466 = n24463 & ~n24465;
  assign n24467 = pi1155 & ~n24466;
  assign n24468 = ~pi1155 & ~n24460;
  assign n24469 = ~n24465 & n24468;
  assign n24470 = ~n24467 & ~n24469;
  assign n24471 = pi785 & ~n24470;
  assign n24472 = ~n24464 & ~n24471;
  assign n24473 = ~pi781 & ~n24472;
  assign n24474 = ~n17289 & n24472;
  assign n24475 = pi1154 & ~n24474;
  assign n24476 = ~n17292 & n24472;
  assign n24477 = ~pi1154 & ~n24476;
  assign n24478 = ~n24475 & ~n24477;
  assign n24479 = pi781 & ~n24478;
  assign n24480 = ~n24473 & ~n24479;
  assign n24481 = ~pi789 & ~n24480;
  assign n24482 = ~n22423 & n24480;
  assign n24483 = pi1159 & ~n24482;
  assign n24484 = ~n22426 & n24480;
  assign n24485 = ~pi1159 & ~n24484;
  assign n24486 = ~n24483 & ~n24485;
  assign n24487 = pi789 & ~n24486;
  assign n24488 = ~n24481 & ~n24487;
  assign n24489 = ~n17355 & n24488;
  assign n24490 = n17355 & n24460;
  assign n24491 = ~n24489 & ~n24490;
  assign n24492 = ~n16124 & ~n24491;
  assign n24493 = n16124 & n24460;
  assign n24494 = ~n24492 & ~n24493;
  assign n24495 = ~n19987 & n24494;
  assign n24496 = ~pi688 & n16742;
  assign n24497 = ~n24460 & ~n24496;
  assign n24498 = ~pi778 & ~n24497;
  assign n24499 = ~pi625 & n24496;
  assign n24500 = ~n24497 & ~n24499;
  assign n24501 = pi1153 & ~n24500;
  assign n24502 = ~pi1153 & ~n24460;
  assign n24503 = ~n24499 & n24502;
  assign n24504 = ~n24501 & ~n24503;
  assign n24505 = pi778 & n24504;
  assign n24506 = ~n24498 & ~n24505;
  assign n24507 = ~n17338 & ~n24506;
  assign n24508 = ~n17340 & n24507;
  assign n24509 = ~n17342 & n24508;
  assign n24510 = ~n17425 & n24509;
  assign n24511 = ~n17452 & n24510;
  assign n24512 = ~pi647 & n24511;
  assign n24513 = pi647 & n24460;
  assign n24514 = ~pi1157 & ~n24513;
  assign n24515 = ~n24512 & n24514;
  assign n24516 = ~pi647 & n24460;
  assign n24517 = pi647 & n24511;
  assign n24518 = pi1157 & ~n24517;
  assign n24519 = ~n24516 & n24518;
  assign n24520 = ~n24515 & ~n24519;
  assign n24521 = ~n17246 & ~n24520;
  assign n24522 = ~n24495 & ~n24521;
  assign n24523 = pi787 & ~n24522;
  assign n24524 = ~pi626 & ~n24488;
  assign n24525 = pi626 & ~n24460;
  assign n24526 = n17181 & ~n24525;
  assign n24527 = ~n24524 & n24526;
  assign n24528 = n17350 & n24509;
  assign n24529 = pi626 & ~n24488;
  assign n24530 = ~pi626 & ~n24460;
  assign n24531 = n17180 & ~n24530;
  assign n24532 = ~n24529 & n24531;
  assign n24533 = ~n24528 & ~n24532;
  assign n24534 = ~n24527 & n24533;
  assign n24535 = pi788 & ~n24534;
  assign n24536 = pi618 & n24507;
  assign n24537 = pi609 & ~n24506;
  assign n24538 = ~n16393 & ~n24497;
  assign n24539 = pi625 & n24538;
  assign n24540 = n24462 & ~n24538;
  assign n24541 = ~n24539 & ~n24540;
  assign n24542 = n24502 & ~n24541;
  assign n24543 = ~pi608 & ~n24501;
  assign n24544 = ~n24542 & n24543;
  assign n24545 = pi1153 & ~n24539;
  assign n24546 = n24462 & n24545;
  assign n24547 = ~n24503 & ~n24546;
  assign n24548 = pi608 & n24547;
  assign n24549 = ~n24544 & ~n24548;
  assign n24550 = pi778 & ~n24549;
  assign n24551 = ~pi778 & ~n24540;
  assign n24552 = ~n24550 & ~n24551;
  assign n24553 = ~pi609 & ~n24552;
  assign n24554 = ~pi1155 & ~n24553;
  assign n24555 = ~n24537 & n24554;
  assign n24556 = ~pi660 & ~n24467;
  assign n24557 = ~n24555 & n24556;
  assign n24558 = ~pi609 & ~n24506;
  assign n24559 = pi609 & ~n24552;
  assign n24560 = ~n24558 & ~n24559;
  assign n24561 = pi1155 & n24560;
  assign n24562 = ~n24469 & ~n24561;
  assign n24563 = pi660 & n24562;
  assign n24564 = ~n24557 & ~n24563;
  assign n24565 = pi785 & ~n24564;
  assign n24566 = ~pi785 & ~n24552;
  assign n24567 = ~n24565 & ~n24566;
  assign n24568 = ~pi618 & ~n24567;
  assign n24569 = ~pi1154 & ~n24568;
  assign n24570 = ~n24536 & n24569;
  assign n24571 = ~pi627 & ~n24475;
  assign n24572 = ~n24570 & n24571;
  assign n24573 = ~pi618 & n24507;
  assign n24574 = pi618 & ~n24567;
  assign n24575 = ~n24573 & ~n24574;
  assign n24576 = pi1154 & n24575;
  assign n24577 = ~n24477 & ~n24576;
  assign n24578 = pi627 & n24577;
  assign n24579 = ~n24572 & ~n24578;
  assign n24580 = pi781 & ~n24579;
  assign n24581 = ~pi781 & ~n24567;
  assign n24582 = ~n24580 & ~n24581;
  assign n24583 = ~pi619 & ~n24582;
  assign n24584 = pi619 & n24508;
  assign n24585 = ~pi1159 & ~n24584;
  assign n24586 = ~n24583 & n24585;
  assign n24587 = ~pi648 & ~n24586;
  assign n24588 = ~n24483 & n24587;
  assign n24589 = ~pi619 & n24508;
  assign n24590 = pi619 & ~n24582;
  assign n24591 = ~n24589 & ~n24590;
  assign n24592 = pi1159 & n24591;
  assign n24593 = ~n24485 & ~n24592;
  assign n24594 = pi648 & n24593;
  assign n24595 = ~n24588 & ~n24594;
  assign n24596 = pi789 & n24595;
  assign n24597 = ~pi789 & n24582;
  assign n24598 = n17356 & ~n24597;
  assign n24599 = ~n24596 & n24598;
  assign n24600 = ~n24535 & ~n24599;
  assign n24601 = n19788 & ~n24600;
  assign n24602 = n20275 & n24510;
  assign n24603 = n17449 & ~n24491;
  assign n24604 = ~pi629 & ~n24603;
  assign n24605 = ~n24602 & n24604;
  assign n24606 = n17448 & ~n24491;
  assign n24607 = n20281 & n24510;
  assign n24608 = pi629 & ~n24607;
  assign n24609 = ~n24606 & n24608;
  assign n24610 = ~n24605 & ~n24609;
  assign n24611 = pi792 & n24610;
  assign n24612 = n19637 & ~n24611;
  assign n24613 = ~n24601 & n24612;
  assign n24614 = ~n24523 & ~n24613;
  assign n24615 = pi644 & n24614;
  assign n24616 = ~pi787 & ~n24511;
  assign n24617 = pi787 & ~n24520;
  assign n24618 = ~n24616 & ~n24617;
  assign n24619 = ~pi644 & n24618;
  assign n24620 = pi715 & ~n24619;
  assign n24621 = ~n24615 & n24620;
  assign n24622 = ~n17247 & ~n24494;
  assign n24623 = n17247 & n24460;
  assign n24624 = ~n24622 & ~n24623;
  assign n24625 = pi644 & ~n24624;
  assign n24626 = ~pi644 & n24460;
  assign n24627 = ~pi715 & ~n24626;
  assign n24628 = ~n24625 & n24627;
  assign n24629 = pi1160 & ~n24628;
  assign n24630 = ~n24621 & n24629;
  assign n24631 = ~pi644 & ~n24624;
  assign n24632 = pi715 & ~n24631;
  assign n24633 = pi644 & n24460;
  assign n24634 = n24632 & ~n24633;
  assign n24635 = pi644 & n24618;
  assign n24636 = ~pi644 & n24614;
  assign n24637 = ~pi715 & ~n24636;
  assign n24638 = ~n24635 & n24637;
  assign n24639 = ~pi1160 & ~n24638;
  assign n24640 = ~n24634 & n24639;
  assign n24641 = ~n24630 & ~n24640;
  assign n24642 = pi790 & ~n24641;
  assign n24643 = ~pi790 & n24614;
  assign n24644 = pi832 & ~n24643;
  assign n24645 = ~n24642 & n24644;
  assign n24646 = ~pi178 & ~n16527;
  assign n24647 = n17159 & ~n24646;
  assign n24648 = n16593 & ~n24646;
  assign n24649 = ~pi688 & n10020;
  assign n24650 = n24646 & ~n24649;
  assign n24651 = ~pi178 & n17592;
  assign n24652 = ~pi38 & ~pi178;
  assign n24653 = n19843 & ~n24652;
  assign n24654 = ~n24651 & ~n24653;
  assign n24655 = ~pi178 & ~n16508;
  assign n24656 = n16744 & ~n24655;
  assign n24657 = ~pi688 & ~n24656;
  assign n24658 = ~n24654 & n24657;
  assign n24659 = ~n24650 & ~n24658;
  assign n24660 = ~pi778 & n24659;
  assign n24661 = pi625 & ~n24659;
  assign n24662 = pi1153 & ~n24661;
  assign n24663 = ~pi625 & n24646;
  assign n24664 = n24662 & ~n24663;
  assign n24665 = ~pi625 & ~n24659;
  assign n24666 = ~pi1153 & ~n24665;
  assign n24667 = pi625 & n24646;
  assign n24668 = n24666 & ~n24667;
  assign n24669 = ~n24664 & ~n24668;
  assign n24670 = pi778 & ~n24669;
  assign n24671 = ~n24660 & ~n24670;
  assign n24672 = ~n16593 & ~n24671;
  assign n24673 = ~n24648 & ~n24672;
  assign n24674 = ~n16589 & n24673;
  assign n24675 = n16589 & n24646;
  assign n24676 = ~n24674 & ~n24675;
  assign n24677 = ~n17159 & n24676;
  assign n24678 = ~n24647 & ~n24677;
  assign n24679 = ~n17183 & n24678;
  assign n24680 = n17183 & n24646;
  assign n24681 = ~n24679 & ~n24680;
  assign n24682 = ~pi792 & n24681;
  assign n24683 = pi628 & ~n24681;
  assign n24684 = pi1156 & ~n24683;
  assign n24685 = ~pi628 & n24646;
  assign n24686 = n24684 & ~n24685;
  assign n24687 = ~pi628 & ~n24681;
  assign n24688 = pi628 & n24646;
  assign n24689 = ~pi1156 & ~n24688;
  assign n24690 = ~n24687 & n24689;
  assign n24691 = ~n24686 & ~n24690;
  assign n24692 = pi792 & ~n24691;
  assign n24693 = ~n24682 & ~n24692;
  assign n24694 = pi647 & ~n24693;
  assign n24695 = ~pi647 & ~n24646;
  assign n24696 = ~n24694 & ~n24695;
  assign n24697 = pi1157 & ~n24696;
  assign n24698 = ~pi647 & n24693;
  assign n24699 = ~pi1157 & ~n24698;
  assign n24700 = pi647 & n24646;
  assign n24701 = n24699 & ~n24700;
  assign n24702 = ~n24697 & ~n24701;
  assign n24703 = pi787 & ~n24702;
  assign n24704 = ~pi787 & ~n24693;
  assign n24705 = ~n24703 & ~n24704;
  assign n24706 = ~pi644 & n24705;
  assign n24707 = pi715 & ~n24706;
  assign n24708 = n17247 & ~n24646;
  assign n24709 = pi178 & ~n10020;
  assign n24710 = ~pi178 & n16449;
  assign n24711 = pi178 & ~n16503;
  assign n24712 = ~pi760 & ~n24711;
  assign n24713 = ~n24710 & n24712;
  assign n24714 = ~pi178 & ~n16357;
  assign n24715 = pi760 & n24714;
  assign n24716 = ~n24713 & ~n24715;
  assign n24717 = ~pi38 & ~n24716;
  assign n24718 = ~pi760 & n16511;
  assign n24719 = ~n24655 & ~n24718;
  assign n24720 = pi38 & ~n24719;
  assign n24721 = n10020 & ~n24720;
  assign n24722 = ~n24717 & n24721;
  assign n24723 = ~n24709 & ~n24722;
  assign n24724 = ~n16521 & ~n24723;
  assign n24725 = n16521 & ~n24646;
  assign n24726 = ~n24724 & ~n24725;
  assign n24727 = ~pi785 & ~n24726;
  assign n24728 = ~n16532 & ~n24646;
  assign n24729 = pi609 & n24724;
  assign n24730 = ~n24728 & ~n24729;
  assign n24731 = pi1155 & ~n24730;
  assign n24732 = ~n16537 & ~n24646;
  assign n24733 = ~pi609 & n24724;
  assign n24734 = ~n24732 & ~n24733;
  assign n24735 = ~pi1155 & ~n24734;
  assign n24736 = ~n24731 & ~n24735;
  assign n24737 = pi785 & ~n24736;
  assign n24738 = ~n24727 & ~n24737;
  assign n24739 = ~pi781 & ~n24738;
  assign n24740 = pi618 & n24738;
  assign n24741 = ~pi618 & n24646;
  assign n24742 = pi1154 & ~n24741;
  assign n24743 = ~n24740 & n24742;
  assign n24744 = ~pi618 & n24738;
  assign n24745 = pi618 & n24646;
  assign n24746 = ~pi1154 & ~n24745;
  assign n24747 = ~n24744 & n24746;
  assign n24748 = ~n24743 & ~n24747;
  assign n24749 = pi781 & ~n24748;
  assign n24750 = ~n24739 & ~n24749;
  assign n24751 = ~pi789 & ~n24750;
  assign n24752 = pi619 & n24750;
  assign n24753 = ~pi619 & n24646;
  assign n24754 = pi1159 & ~n24753;
  assign n24755 = ~n24752 & n24754;
  assign n24756 = ~pi619 & n24750;
  assign n24757 = pi619 & n24646;
  assign n24758 = ~pi1159 & ~n24757;
  assign n24759 = ~n24756 & n24758;
  assign n24760 = ~n24755 & ~n24759;
  assign n24761 = pi789 & ~n24760;
  assign n24762 = ~n24751 & ~n24761;
  assign n24763 = ~n17355 & n24762;
  assign n24764 = n17355 & n24646;
  assign n24765 = ~n24763 & ~n24764;
  assign n24766 = ~n16124 & ~n24765;
  assign n24767 = n16124 & n24646;
  assign n24768 = ~n24766 & ~n24767;
  assign n24769 = ~n17247 & n24768;
  assign n24770 = ~n24708 & ~n24769;
  assign n24771 = pi644 & n24770;
  assign n24772 = ~pi644 & n24646;
  assign n24773 = ~pi715 & ~n24772;
  assign n24774 = ~n24771 & n24773;
  assign n24775 = pi1160 & ~n24774;
  assign n24776 = ~n24707 & n24775;
  assign n24777 = pi644 & n24705;
  assign n24778 = ~pi715 & ~n24777;
  assign n24779 = ~pi644 & n24770;
  assign n24780 = pi644 & n24646;
  assign n24781 = ~n24779 & ~n24780;
  assign n24782 = pi715 & n24781;
  assign n24783 = ~pi1160 & ~n24782;
  assign n24784 = ~n24778 & n24783;
  assign n24785 = ~n24776 & ~n24784;
  assign n24786 = pi790 & ~n24785;
  assign n24787 = ~pi629 & n24686;
  assign n24788 = ~n19999 & n24765;
  assign n24789 = pi629 & n24690;
  assign n24790 = ~n24788 & ~n24789;
  assign n24791 = ~n24787 & n24790;
  assign n24792 = pi792 & ~n24791;
  assign n24793 = pi618 & n24673;
  assign n24794 = pi609 & n24671;
  assign n24795 = pi625 & n24723;
  assign n24796 = ~n24649 & ~n24722;
  assign n24797 = ~pi760 & ~n16917;
  assign n24798 = n18933 & ~n24797;
  assign n24799 = ~pi178 & ~n24798;
  assign n24800 = ~n17079 & ~n24461;
  assign n24801 = pi178 & ~n24800;
  assign n24802 = n6097 & n24801;
  assign n24803 = ~n24799 & ~n24802;
  assign n24804 = pi38 & n24803;
  assign n24805 = ~pi178 & n16853;
  assign n24806 = pi178 & n16935;
  assign n24807 = pi760 & ~n24806;
  assign n24808 = ~n24805 & n24807;
  assign n24809 = pi178 & n16998;
  assign n24810 = ~pi178 & ~n17051;
  assign n24811 = ~pi760 & ~n24810;
  assign n24812 = ~n24809 & n24811;
  assign n24813 = ~n24808 & ~n24812;
  assign n24814 = pi39 & n24813;
  assign n24815 = ~pi178 & ~n17061;
  assign n24816 = pi178 & ~n17058;
  assign n24817 = pi760 & ~n24816;
  assign n24818 = ~n24815 & n24817;
  assign n24819 = ~pi178 & n17067;
  assign n24820 = pi178 & n17065;
  assign n24821 = ~pi760 & ~n24820;
  assign n24822 = ~n24819 & n24821;
  assign n24823 = ~n24818 & ~n24822;
  assign n24824 = ~pi39 & ~n24823;
  assign n24825 = ~pi38 & ~n24824;
  assign n24826 = ~n24814 & n24825;
  assign n24827 = ~pi688 & ~n24826;
  assign n24828 = ~n24804 & n24827;
  assign n24829 = ~n24796 & ~n24828;
  assign n24830 = ~n24709 & ~n24829;
  assign n24831 = ~pi625 & n24830;
  assign n24832 = ~pi1153 & ~n24831;
  assign n24833 = ~n24795 & n24832;
  assign n24834 = ~pi608 & ~n24664;
  assign n24835 = ~n24833 & n24834;
  assign n24836 = ~pi625 & n24723;
  assign n24837 = pi625 & n24830;
  assign n24838 = ~n24836 & ~n24837;
  assign n24839 = pi1153 & n24838;
  assign n24840 = ~n24668 & ~n24839;
  assign n24841 = pi608 & n24840;
  assign n24842 = ~n24835 & ~n24841;
  assign n24843 = pi778 & ~n24842;
  assign n24844 = ~pi778 & n24830;
  assign n24845 = ~n24843 & ~n24844;
  assign n24846 = ~pi609 & ~n24845;
  assign n24847 = ~pi1155 & ~n24846;
  assign n24848 = ~n24794 & n24847;
  assign n24849 = ~pi660 & ~n24731;
  assign n24850 = ~n24848 & n24849;
  assign n24851 = ~pi609 & n24671;
  assign n24852 = pi609 & ~n24845;
  assign n24853 = ~n24851 & ~n24852;
  assign n24854 = pi1155 & n24853;
  assign n24855 = ~n24735 & ~n24854;
  assign n24856 = pi660 & n24855;
  assign n24857 = ~n24850 & ~n24856;
  assign n24858 = pi785 & ~n24857;
  assign n24859 = ~pi785 & ~n24845;
  assign n24860 = ~n24858 & ~n24859;
  assign n24861 = ~pi618 & ~n24860;
  assign n24862 = ~pi1154 & ~n24861;
  assign n24863 = ~n24793 & n24862;
  assign n24864 = ~pi627 & ~n24743;
  assign n24865 = ~n24863 & n24864;
  assign n24866 = ~pi618 & n24673;
  assign n24867 = pi618 & ~n24860;
  assign n24868 = ~n24866 & ~n24867;
  assign n24869 = pi1154 & n24868;
  assign n24870 = ~n24747 & ~n24869;
  assign n24871 = pi627 & n24870;
  assign n24872 = ~n24865 & ~n24871;
  assign n24873 = pi781 & ~n24872;
  assign n24874 = ~pi781 & ~n24860;
  assign n24875 = ~n24873 & ~n24874;
  assign n24876 = ~pi789 & n24875;
  assign n24877 = ~pi619 & ~n24875;
  assign n24878 = pi619 & ~n24676;
  assign n24879 = ~pi1159 & ~n24878;
  assign n24880 = ~n24877 & n24879;
  assign n24881 = ~pi648 & ~n24880;
  assign n24882 = ~n24755 & n24881;
  assign n24883 = ~pi619 & ~n24676;
  assign n24884 = pi619 & ~n24875;
  assign n24885 = ~n24883 & ~n24884;
  assign n24886 = pi1159 & n24885;
  assign n24887 = ~n24759 & ~n24886;
  assign n24888 = pi648 & n24887;
  assign n24889 = ~n24882 & ~n24888;
  assign n24890 = pi789 & n24889;
  assign n24891 = ~n24876 & ~n24890;
  assign n24892 = n17356 & n24891;
  assign n24893 = ~pi626 & ~n24762;
  assign n24894 = pi626 & ~n24646;
  assign n24895 = n17181 & ~n24894;
  assign n24896 = ~n24893 & n24895;
  assign n24897 = n17350 & n24678;
  assign n24898 = pi626 & ~n24762;
  assign n24899 = ~pi626 & ~n24646;
  assign n24900 = n17180 & ~n24899;
  assign n24901 = ~n24898 & n24900;
  assign n24902 = ~n24897 & ~n24901;
  assign n24903 = ~n24896 & n24902;
  assign n24904 = pi788 & ~n24903;
  assign n24905 = n19788 & ~n24904;
  assign n24906 = ~n24892 & n24905;
  assign n24907 = ~n24792 & ~n24906;
  assign n24908 = n19637 & ~n24907;
  assign n24909 = ~n19987 & n24768;
  assign n24910 = pi630 & n24701;
  assign n24911 = ~n24909 & ~n24910;
  assign n24912 = n17244 & ~n24696;
  assign n24913 = n24911 & ~n24912;
  assign n24914 = pi787 & ~n24913;
  assign n24915 = ~n24908 & ~n24914;
  assign n24916 = pi644 & n24775;
  assign n24917 = ~pi644 & n24783;
  assign n24918 = pi790 & ~n24917;
  assign n24919 = ~n24916 & n24918;
  assign n24920 = n24915 & ~n24919;
  assign n24921 = ~n24786 & ~n24920;
  assign n24922 = ~po1038 & ~n24921;
  assign n24923 = ~pi178 & po1038;
  assign n24924 = ~pi832 & ~n24923;
  assign n24925 = ~n24922 & n24924;
  assign po335 = ~n24645 & ~n24925;
  assign n24927 = pi179 & ~n10020;
  assign n24928 = ~pi741 & ~n23777;
  assign n24929 = pi179 & ~n24928;
  assign n24930 = ~n18802 & n18808;
  assign n24931 = ~pi179 & n24930;
  assign n24932 = ~pi741 & n24931;
  assign n24933 = ~n21074 & ~n24932;
  assign n24934 = ~n24929 & n24933;
  assign n24935 = n10020 & ~n24934;
  assign n24936 = ~n24927 & ~n24935;
  assign n24937 = ~n16521 & ~n24936;
  assign n24938 = ~pi179 & ~n16527;
  assign n24939 = n16521 & ~n24938;
  assign n24940 = ~n24937 & ~n24939;
  assign n24941 = ~pi785 & ~n24940;
  assign n24942 = ~n16532 & ~n24938;
  assign n24943 = pi609 & n24937;
  assign n24944 = ~n24942 & ~n24943;
  assign n24945 = pi1155 & ~n24944;
  assign n24946 = ~n16537 & ~n24938;
  assign n24947 = ~pi609 & n24937;
  assign n24948 = ~n24946 & ~n24947;
  assign n24949 = ~pi1155 & ~n24948;
  assign n24950 = ~n24945 & ~n24949;
  assign n24951 = pi785 & ~n24950;
  assign n24952 = ~n24941 & ~n24951;
  assign n24953 = ~pi781 & ~n24952;
  assign n24954 = pi618 & n24952;
  assign n24955 = ~pi618 & n24938;
  assign n24956 = pi1154 & ~n24955;
  assign n24957 = ~n24954 & n24956;
  assign n24958 = ~pi618 & n24952;
  assign n24959 = pi618 & n24938;
  assign n24960 = ~pi1154 & ~n24959;
  assign n24961 = ~n24958 & n24960;
  assign n24962 = ~n24957 & ~n24961;
  assign n24963 = pi781 & ~n24962;
  assign n24964 = ~n24953 & ~n24963;
  assign n24965 = ~pi789 & ~n24964;
  assign n24966 = pi619 & n24964;
  assign n24967 = ~pi619 & n24938;
  assign n24968 = pi1159 & ~n24967;
  assign n24969 = ~n24966 & n24968;
  assign n24970 = ~pi619 & n24964;
  assign n24971 = pi619 & n24938;
  assign n24972 = ~pi1159 & ~n24971;
  assign n24973 = ~n24970 & n24972;
  assign n24974 = ~n24969 & ~n24973;
  assign n24975 = pi789 & ~n24974;
  assign n24976 = ~n24965 & ~n24975;
  assign n24977 = ~n17355 & n24976;
  assign n24978 = n17355 & n24938;
  assign n24979 = ~n24977 & ~n24978;
  assign n24980 = ~n16124 & ~n24979;
  assign n24981 = n16124 & n24938;
  assign n24982 = ~n24980 & ~n24981;
  assign n24983 = pi647 & ~n24982;
  assign n24984 = pi628 & ~n24979;
  assign n24985 = n16593 & ~n24938;
  assign n24986 = ~pi724 & n10020;
  assign n24987 = n24938 & ~n24986;
  assign n24988 = ~pi179 & n17592;
  assign n24989 = ~pi38 & ~pi179;
  assign n24990 = n19843 & ~n24989;
  assign n24991 = ~n24988 & ~n24990;
  assign n24992 = ~pi179 & ~n16508;
  assign n24993 = n16744 & ~n24992;
  assign n24994 = ~pi724 & ~n24993;
  assign n24995 = ~n24991 & n24994;
  assign n24996 = ~n24987 & ~n24995;
  assign n24997 = ~pi778 & n24996;
  assign n24998 = pi625 & ~n24996;
  assign n24999 = pi1153 & ~n24998;
  assign n25000 = ~pi625 & n24938;
  assign n25001 = n24999 & ~n25000;
  assign n25002 = ~pi625 & ~n24996;
  assign n25003 = ~pi1153 & ~n25002;
  assign n25004 = pi625 & n24938;
  assign n25005 = n25003 & ~n25004;
  assign n25006 = ~n25001 & ~n25005;
  assign n25007 = pi778 & ~n25006;
  assign n25008 = ~n24997 & ~n25007;
  assign n25009 = ~n16593 & ~n25008;
  assign n25010 = ~n24985 & ~n25009;
  assign n25011 = ~n16589 & n25010;
  assign n25012 = n16589 & n24938;
  assign n25013 = ~n25011 & ~n25012;
  assign n25014 = pi619 & ~n25013;
  assign n25015 = pi618 & n25010;
  assign n25016 = pi609 & n25008;
  assign n25017 = pi625 & n24936;
  assign n25018 = ~n24935 & ~n24986;
  assign n25019 = n17627 & ~n24992;
  assign n25020 = ~pi179 & n16853;
  assign n25021 = pi179 & n16935;
  assign n25022 = pi39 & ~n25021;
  assign n25023 = ~n25020 & n25022;
  assign n25024 = pi179 & n17058;
  assign n25025 = ~pi179 & n17061;
  assign n25026 = ~pi39 & ~n25025;
  assign n25027 = ~n25024 & n25026;
  assign n25028 = ~n25023 & ~n25027;
  assign n25029 = ~pi38 & ~n25028;
  assign n25030 = ~n25019 & ~n25029;
  assign n25031 = pi741 & ~n25030;
  assign n25032 = ~pi179 & ~n18914;
  assign n25033 = pi179 & n18922;
  assign n25034 = ~pi741 & ~n25033;
  assign n25035 = ~n25032 & n25034;
  assign n25036 = ~pi724 & ~n25035;
  assign n25037 = ~n25031 & n25036;
  assign n25038 = ~n25018 & ~n25037;
  assign n25039 = ~n24927 & ~n25038;
  assign n25040 = ~pi625 & n25039;
  assign n25041 = ~pi1153 & ~n25040;
  assign n25042 = ~n25017 & n25041;
  assign n25043 = ~pi608 & ~n25001;
  assign n25044 = ~n25042 & n25043;
  assign n25045 = ~pi625 & n24936;
  assign n25046 = pi625 & n25039;
  assign n25047 = ~n25045 & ~n25046;
  assign n25048 = pi1153 & n25047;
  assign n25049 = ~n25005 & ~n25048;
  assign n25050 = pi608 & n25049;
  assign n25051 = ~n25044 & ~n25050;
  assign n25052 = pi778 & ~n25051;
  assign n25053 = ~pi778 & n25039;
  assign n25054 = ~n25052 & ~n25053;
  assign n25055 = ~pi609 & ~n25054;
  assign n25056 = ~pi1155 & ~n25055;
  assign n25057 = ~n25016 & n25056;
  assign n25058 = ~pi660 & ~n24945;
  assign n25059 = ~n25057 & n25058;
  assign n25060 = ~pi609 & n25008;
  assign n25061 = pi609 & ~n25054;
  assign n25062 = ~n25060 & ~n25061;
  assign n25063 = pi1155 & n25062;
  assign n25064 = ~n24949 & ~n25063;
  assign n25065 = pi660 & n25064;
  assign n25066 = ~n25059 & ~n25065;
  assign n25067 = pi785 & ~n25066;
  assign n25068 = ~pi785 & ~n25054;
  assign n25069 = ~n25067 & ~n25068;
  assign n25070 = ~pi618 & ~n25069;
  assign n25071 = ~pi1154 & ~n25070;
  assign n25072 = ~n25015 & n25071;
  assign n25073 = ~pi627 & ~n24957;
  assign n25074 = ~n25072 & n25073;
  assign n25075 = ~pi618 & n25010;
  assign n25076 = pi618 & ~n25069;
  assign n25077 = ~n25075 & ~n25076;
  assign n25078 = pi1154 & n25077;
  assign n25079 = ~n24961 & ~n25078;
  assign n25080 = pi627 & n25079;
  assign n25081 = ~n25074 & ~n25080;
  assign n25082 = pi781 & ~n25081;
  assign n25083 = ~pi781 & ~n25069;
  assign n25084 = ~n25082 & ~n25083;
  assign n25085 = ~pi619 & ~n25084;
  assign n25086 = ~pi1159 & ~n25085;
  assign n25087 = ~n25014 & n25086;
  assign n25088 = ~pi648 & ~n24969;
  assign n25089 = ~n25087 & n25088;
  assign n25090 = ~pi619 & ~n25013;
  assign n25091 = pi619 & ~n25084;
  assign n25092 = ~n25090 & ~n25091;
  assign n25093 = pi1159 & n25092;
  assign n25094 = ~n24973 & ~n25093;
  assign n25095 = pi648 & n25094;
  assign n25096 = ~n25089 & ~n25095;
  assign n25097 = pi789 & ~n25096;
  assign n25098 = ~pi789 & ~n25084;
  assign n25099 = ~n25097 & ~n25098;
  assign n25100 = ~pi788 & n25099;
  assign n25101 = pi626 & n25099;
  assign n25102 = n17159 & ~n24938;
  assign n25103 = ~n17159 & n25013;
  assign n25104 = ~n25102 & ~n25103;
  assign n25105 = ~pi626 & ~n25104;
  assign n25106 = pi641 & ~n25105;
  assign n25107 = ~n25101 & n25106;
  assign n25108 = pi626 & ~n24976;
  assign n25109 = ~pi626 & ~n24938;
  assign n25110 = ~pi641 & ~n25109;
  assign n25111 = ~n25108 & n25110;
  assign n25112 = pi1158 & ~n25111;
  assign n25113 = ~n25107 & n25112;
  assign n25114 = pi626 & ~n24938;
  assign n25115 = ~pi626 & ~n24976;
  assign n25116 = pi641 & ~n25115;
  assign n25117 = ~n25114 & n25116;
  assign n25118 = pi626 & ~n25104;
  assign n25119 = ~pi626 & n25099;
  assign n25120 = ~pi641 & ~n25119;
  assign n25121 = ~n25118 & n25120;
  assign n25122 = ~pi1158 & ~n25121;
  assign n25123 = ~n25117 & n25122;
  assign n25124 = ~n25113 & ~n25123;
  assign n25125 = pi788 & ~n25124;
  assign n25126 = ~n25100 & ~n25125;
  assign n25127 = ~pi628 & n25126;
  assign n25128 = ~pi1156 & ~n25127;
  assign n25129 = ~n24984 & n25128;
  assign n25130 = ~n17183 & n25104;
  assign n25131 = n17183 & n24938;
  assign n25132 = ~n25130 & ~n25131;
  assign n25133 = pi628 & ~n25132;
  assign n25134 = pi1156 & ~n25133;
  assign n25135 = ~pi628 & n24938;
  assign n25136 = n25134 & ~n25135;
  assign n25137 = ~pi629 & ~n25136;
  assign n25138 = ~n25129 & n25137;
  assign n25139 = ~pi628 & ~n25132;
  assign n25140 = pi628 & n24938;
  assign n25141 = ~pi1156 & ~n25140;
  assign n25142 = ~n25139 & n25141;
  assign n25143 = ~pi628 & ~n24979;
  assign n25144 = pi628 & n25126;
  assign n25145 = ~n25143 & ~n25144;
  assign n25146 = pi1156 & n25145;
  assign n25147 = ~n25142 & ~n25146;
  assign n25148 = pi629 & n25147;
  assign n25149 = ~n25138 & ~n25148;
  assign n25150 = pi792 & ~n25149;
  assign n25151 = ~pi792 & n25126;
  assign n25152 = ~n25150 & ~n25151;
  assign n25153 = ~pi647 & ~n25152;
  assign n25154 = ~pi1157 & ~n25153;
  assign n25155 = ~n24983 & n25154;
  assign n25156 = ~pi792 & n25132;
  assign n25157 = ~n25136 & ~n25142;
  assign n25158 = pi792 & ~n25157;
  assign n25159 = ~n25156 & ~n25158;
  assign n25160 = pi647 & n25159;
  assign n25161 = pi1157 & ~n25160;
  assign n25162 = ~pi647 & n24938;
  assign n25163 = n25161 & ~n25162;
  assign n25164 = ~pi630 & ~n25163;
  assign n25165 = ~n25155 & n25164;
  assign n25166 = ~pi647 & n25159;
  assign n25167 = pi647 & n24938;
  assign n25168 = ~pi1157 & ~n25167;
  assign n25169 = ~n25166 & n25168;
  assign n25170 = ~pi647 & ~n24982;
  assign n25171 = pi647 & ~n25152;
  assign n25172 = ~n25170 & ~n25171;
  assign n25173 = pi1157 & n25172;
  assign n25174 = ~n25169 & ~n25173;
  assign n25175 = pi630 & n25174;
  assign n25176 = ~n25165 & ~n25175;
  assign n25177 = pi787 & ~n25176;
  assign n25178 = ~pi787 & ~n25152;
  assign n25179 = ~n25177 & ~n25178;
  assign n25180 = ~pi790 & n25179;
  assign n25181 = pi644 & ~n25179;
  assign n25182 = ~pi787 & ~n25159;
  assign n25183 = ~n25163 & ~n25169;
  assign n25184 = pi787 & ~n25183;
  assign n25185 = ~n25182 & ~n25184;
  assign n25186 = ~pi644 & n25185;
  assign n25187 = pi715 & ~n25186;
  assign n25188 = ~n25181 & n25187;
  assign n25189 = ~pi644 & n24938;
  assign n25190 = n17247 & ~n24938;
  assign n25191 = ~n17247 & n24982;
  assign n25192 = ~n25190 & ~n25191;
  assign n25193 = pi644 & n25192;
  assign n25194 = ~pi715 & ~n25193;
  assign n25195 = ~n25189 & n25194;
  assign n25196 = ~n25188 & ~n25195;
  assign n25197 = pi1160 & n25196;
  assign n25198 = ~pi644 & n25192;
  assign n25199 = pi715 & ~n25198;
  assign n25200 = pi644 & n24938;
  assign n25201 = n25199 & ~n25200;
  assign n25202 = pi644 & n25185;
  assign n25203 = ~pi644 & ~n25179;
  assign n25204 = ~pi715 & ~n25203;
  assign n25205 = ~n25202 & n25204;
  assign n25206 = ~n25201 & ~n25205;
  assign n25207 = ~pi1160 & n25206;
  assign n25208 = ~n25197 & ~n25207;
  assign n25209 = pi790 & n25208;
  assign n25210 = ~n25180 & ~n25209;
  assign n25211 = ~po1038 & n25210;
  assign n25212 = ~pi179 & po1038;
  assign n25213 = ~pi832 & ~n25212;
  assign n25214 = ~n25211 & n25213;
  assign n25215 = ~pi179 & ~n2934;
  assign n25216 = ~pi741 & n16510;
  assign n25217 = ~n25215 & ~n25216;
  assign n25218 = ~n17273 & ~n25217;
  assign n25219 = ~pi785 & ~n25218;
  assign n25220 = ~n17279 & ~n25217;
  assign n25221 = pi1155 & ~n25220;
  assign n25222 = ~n17282 & n25218;
  assign n25223 = ~pi1155 & ~n25222;
  assign n25224 = ~n25221 & ~n25223;
  assign n25225 = pi785 & ~n25224;
  assign n25226 = ~n25219 & ~n25225;
  assign n25227 = ~pi781 & ~n25226;
  assign n25228 = ~n17289 & n25226;
  assign n25229 = pi1154 & ~n25228;
  assign n25230 = ~n17292 & n25226;
  assign n25231 = ~pi1154 & ~n25230;
  assign n25232 = ~n25229 & ~n25231;
  assign n25233 = pi781 & ~n25232;
  assign n25234 = ~n25227 & ~n25233;
  assign n25235 = ~pi789 & ~n25234;
  assign n25236 = pi619 & n25234;
  assign n25237 = ~pi619 & n25215;
  assign n25238 = pi1159 & ~n25237;
  assign n25239 = ~n25236 & n25238;
  assign n25240 = ~pi619 & n25234;
  assign n25241 = pi619 & n25215;
  assign n25242 = ~pi1159 & ~n25241;
  assign n25243 = ~n25240 & n25242;
  assign n25244 = ~n25239 & ~n25243;
  assign n25245 = pi789 & ~n25244;
  assign n25246 = ~n25235 & ~n25245;
  assign n25247 = ~n17355 & n25246;
  assign n25248 = n17355 & n25215;
  assign n25249 = ~n25247 & ~n25248;
  assign n25250 = ~n16124 & ~n25249;
  assign n25251 = n16124 & n25215;
  assign n25252 = ~n25250 & ~n25251;
  assign n25253 = ~n19987 & n25252;
  assign n25254 = ~pi724 & n16742;
  assign n25255 = ~n25215 & ~n25254;
  assign n25256 = ~pi778 & n25255;
  assign n25257 = ~pi625 & n25254;
  assign n25258 = ~n25255 & ~n25257;
  assign n25259 = pi1153 & ~n25258;
  assign n25260 = ~pi1153 & ~n25215;
  assign n25261 = ~n25257 & n25260;
  assign n25262 = ~n25259 & ~n25261;
  assign n25263 = pi778 & ~n25262;
  assign n25264 = ~n25256 & ~n25263;
  assign n25265 = ~n17338 & n25264;
  assign n25266 = ~n17340 & n25265;
  assign n25267 = ~n17342 & n25266;
  assign n25268 = ~n17425 & n25267;
  assign n25269 = ~n17452 & n25268;
  assign n25270 = ~pi647 & n25269;
  assign n25271 = pi647 & n25215;
  assign n25272 = ~pi1157 & ~n25271;
  assign n25273 = ~n25270 & n25272;
  assign n25274 = ~pi647 & n25215;
  assign n25275 = pi647 & n25269;
  assign n25276 = pi1157 & ~n25275;
  assign n25277 = ~n25274 & n25276;
  assign n25278 = ~n25273 & ~n25277;
  assign n25279 = ~n17246 & ~n25278;
  assign n25280 = ~n25253 & ~n25279;
  assign n25281 = pi787 & ~n25280;
  assign n25282 = ~pi626 & ~n25246;
  assign n25283 = pi626 & ~n25215;
  assign n25284 = n17181 & ~n25283;
  assign n25285 = ~n25282 & n25284;
  assign n25286 = n17350 & n25267;
  assign n25287 = pi626 & ~n25246;
  assign n25288 = ~pi626 & ~n25215;
  assign n25289 = n17180 & ~n25288;
  assign n25290 = ~n25287 & n25289;
  assign n25291 = ~n25286 & ~n25290;
  assign n25292 = ~n25285 & n25291;
  assign n25293 = pi788 & ~n25292;
  assign n25294 = pi618 & n25265;
  assign n25295 = pi609 & n25264;
  assign n25296 = ~n16393 & ~n25255;
  assign n25297 = pi625 & n25296;
  assign n25298 = n25217 & ~n25296;
  assign n25299 = ~n25297 & ~n25298;
  assign n25300 = n25260 & ~n25299;
  assign n25301 = ~pi608 & ~n25259;
  assign n25302 = ~n25300 & n25301;
  assign n25303 = pi1153 & ~n25297;
  assign n25304 = n25217 & n25303;
  assign n25305 = ~n25261 & ~n25304;
  assign n25306 = pi608 & n25305;
  assign n25307 = ~n25302 & ~n25306;
  assign n25308 = pi778 & ~n25307;
  assign n25309 = ~pi778 & ~n25298;
  assign n25310 = ~n25308 & ~n25309;
  assign n25311 = ~pi609 & ~n25310;
  assign n25312 = ~pi1155 & ~n25311;
  assign n25313 = ~n25295 & n25312;
  assign n25314 = ~pi660 & ~n25221;
  assign n25315 = ~n25313 & n25314;
  assign n25316 = ~pi609 & n25264;
  assign n25317 = pi609 & ~n25310;
  assign n25318 = ~n25316 & ~n25317;
  assign n25319 = pi1155 & n25318;
  assign n25320 = ~n25223 & ~n25319;
  assign n25321 = pi660 & n25320;
  assign n25322 = ~n25315 & ~n25321;
  assign n25323 = pi785 & ~n25322;
  assign n25324 = ~pi785 & ~n25310;
  assign n25325 = ~n25323 & ~n25324;
  assign n25326 = ~pi618 & ~n25325;
  assign n25327 = ~pi1154 & ~n25326;
  assign n25328 = ~n25294 & n25327;
  assign n25329 = ~pi627 & ~n25229;
  assign n25330 = ~n25328 & n25329;
  assign n25331 = ~pi618 & n25265;
  assign n25332 = pi618 & ~n25325;
  assign n25333 = ~n25331 & ~n25332;
  assign n25334 = pi1154 & n25333;
  assign n25335 = ~n25231 & ~n25334;
  assign n25336 = pi627 & n25335;
  assign n25337 = ~n25330 & ~n25336;
  assign n25338 = pi781 & ~n25337;
  assign n25339 = ~pi781 & ~n25325;
  assign n25340 = ~n25338 & ~n25339;
  assign n25341 = ~pi619 & ~n25340;
  assign n25342 = pi619 & n25266;
  assign n25343 = ~pi1159 & ~n25342;
  assign n25344 = ~n25341 & n25343;
  assign n25345 = ~pi648 & ~n25344;
  assign n25346 = ~n25239 & n25345;
  assign n25347 = ~pi619 & n25266;
  assign n25348 = pi619 & ~n25340;
  assign n25349 = ~n25347 & ~n25348;
  assign n25350 = pi1159 & n25349;
  assign n25351 = ~n25243 & ~n25350;
  assign n25352 = pi648 & n25351;
  assign n25353 = ~n25346 & ~n25352;
  assign n25354 = pi789 & n25353;
  assign n25355 = ~pi789 & n25340;
  assign n25356 = n17356 & ~n25355;
  assign n25357 = ~n25354 & n25356;
  assign n25358 = ~n25293 & ~n25357;
  assign n25359 = n19788 & ~n25358;
  assign n25360 = n20275 & n25268;
  assign n25361 = n17449 & ~n25249;
  assign n25362 = ~pi629 & ~n25361;
  assign n25363 = ~n25360 & n25362;
  assign n25364 = n17448 & ~n25249;
  assign n25365 = n20281 & n25268;
  assign n25366 = pi629 & ~n25365;
  assign n25367 = ~n25364 & n25366;
  assign n25368 = ~n25363 & ~n25367;
  assign n25369 = pi792 & n25368;
  assign n25370 = n19637 & ~n25369;
  assign n25371 = ~n25359 & n25370;
  assign n25372 = ~n25281 & ~n25371;
  assign n25373 = pi644 & n25372;
  assign n25374 = ~pi787 & ~n25269;
  assign n25375 = pi787 & ~n25278;
  assign n25376 = ~n25374 & ~n25375;
  assign n25377 = ~pi644 & n25376;
  assign n25378 = pi715 & ~n25377;
  assign n25379 = ~n25373 & n25378;
  assign n25380 = ~n17247 & ~n25252;
  assign n25381 = n17247 & n25215;
  assign n25382 = ~n25380 & ~n25381;
  assign n25383 = pi644 & ~n25382;
  assign n25384 = ~pi644 & n25215;
  assign n25385 = ~pi715 & ~n25384;
  assign n25386 = ~n25383 & n25385;
  assign n25387 = pi1160 & ~n25386;
  assign n25388 = ~n25379 & n25387;
  assign n25389 = ~pi644 & ~n25382;
  assign n25390 = pi715 & ~n25389;
  assign n25391 = pi644 & n25215;
  assign n25392 = n25390 & ~n25391;
  assign n25393 = pi644 & n25376;
  assign n25394 = ~pi644 & n25372;
  assign n25395 = ~pi715 & ~n25394;
  assign n25396 = ~n25393 & n25395;
  assign n25397 = ~pi1160 & ~n25396;
  assign n25398 = ~n25392 & n25397;
  assign n25399 = ~n25388 & ~n25398;
  assign n25400 = pi790 & ~n25399;
  assign n25401 = ~pi790 & n25372;
  assign n25402 = pi832 & ~n25401;
  assign n25403 = ~n25400 & n25402;
  assign po336 = ~n25214 & ~n25403;
  assign n25405 = ~pi180 & ~n2934;
  assign n25406 = ~pi753 & n16510;
  assign n25407 = ~n25405 & ~n25406;
  assign n25408 = ~n17273 & ~n25407;
  assign n25409 = ~pi785 & ~n25408;
  assign n25410 = n16537 & n25406;
  assign n25411 = n25408 & ~n25410;
  assign n25412 = pi1155 & ~n25411;
  assign n25413 = ~pi1155 & ~n25405;
  assign n25414 = ~n25410 & n25413;
  assign n25415 = ~n25412 & ~n25414;
  assign n25416 = pi785 & ~n25415;
  assign n25417 = ~n25409 & ~n25416;
  assign n25418 = ~pi781 & ~n25417;
  assign n25419 = ~n17289 & n25417;
  assign n25420 = pi1154 & ~n25419;
  assign n25421 = ~n17292 & n25417;
  assign n25422 = ~pi1154 & ~n25421;
  assign n25423 = ~n25420 & ~n25422;
  assign n25424 = pi781 & ~n25423;
  assign n25425 = ~n25418 & ~n25424;
  assign n25426 = ~pi789 & ~n25425;
  assign n25427 = ~n22423 & n25425;
  assign n25428 = pi1159 & ~n25427;
  assign n25429 = ~n22426 & n25425;
  assign n25430 = ~pi1159 & ~n25429;
  assign n25431 = ~n25428 & ~n25430;
  assign n25432 = pi789 & ~n25431;
  assign n25433 = ~n25426 & ~n25432;
  assign n25434 = ~n17355 & n25433;
  assign n25435 = n17355 & n25405;
  assign n25436 = ~n25434 & ~n25435;
  assign n25437 = ~n16124 & ~n25436;
  assign n25438 = n16124 & n25405;
  assign n25439 = ~n25437 & ~n25438;
  assign n25440 = ~n19987 & n25439;
  assign n25441 = ~pi702 & n16742;
  assign n25442 = ~n25405 & ~n25441;
  assign n25443 = ~pi778 & ~n25442;
  assign n25444 = ~pi625 & n25441;
  assign n25445 = ~n25442 & ~n25444;
  assign n25446 = pi1153 & ~n25445;
  assign n25447 = ~pi1153 & ~n25405;
  assign n25448 = ~n25444 & n25447;
  assign n25449 = ~n25446 & ~n25448;
  assign n25450 = pi778 & n25449;
  assign n25451 = ~n25443 & ~n25450;
  assign n25452 = ~n17338 & ~n25451;
  assign n25453 = ~n17340 & n25452;
  assign n25454 = ~n17342 & n25453;
  assign n25455 = ~n17425 & n25454;
  assign n25456 = ~n17452 & n25455;
  assign n25457 = ~pi647 & n25456;
  assign n25458 = pi647 & n25405;
  assign n25459 = ~pi1157 & ~n25458;
  assign n25460 = ~n25457 & n25459;
  assign n25461 = ~pi647 & n25405;
  assign n25462 = pi647 & n25456;
  assign n25463 = pi1157 & ~n25462;
  assign n25464 = ~n25461 & n25463;
  assign n25465 = ~n25460 & ~n25464;
  assign n25466 = ~n17246 & ~n25465;
  assign n25467 = ~n25440 & ~n25466;
  assign n25468 = pi787 & ~n25467;
  assign n25469 = ~pi626 & ~n25433;
  assign n25470 = pi626 & ~n25405;
  assign n25471 = n17181 & ~n25470;
  assign n25472 = ~n25469 & n25471;
  assign n25473 = n17350 & n25454;
  assign n25474 = pi626 & ~n25433;
  assign n25475 = ~pi626 & ~n25405;
  assign n25476 = n17180 & ~n25475;
  assign n25477 = ~n25474 & n25476;
  assign n25478 = ~n25473 & ~n25477;
  assign n25479 = ~n25472 & n25478;
  assign n25480 = pi788 & ~n25479;
  assign n25481 = pi618 & n25452;
  assign n25482 = pi609 & ~n25451;
  assign n25483 = ~n16393 & ~n25442;
  assign n25484 = pi625 & n25483;
  assign n25485 = n25407 & ~n25483;
  assign n25486 = ~n25484 & ~n25485;
  assign n25487 = n25447 & ~n25486;
  assign n25488 = ~pi608 & ~n25446;
  assign n25489 = ~n25487 & n25488;
  assign n25490 = pi1153 & ~n25484;
  assign n25491 = n25407 & n25490;
  assign n25492 = ~n25448 & ~n25491;
  assign n25493 = pi608 & n25492;
  assign n25494 = ~n25489 & ~n25493;
  assign n25495 = pi778 & ~n25494;
  assign n25496 = ~pi778 & ~n25485;
  assign n25497 = ~n25495 & ~n25496;
  assign n25498 = ~pi609 & ~n25497;
  assign n25499 = ~pi1155 & ~n25498;
  assign n25500 = ~n25482 & n25499;
  assign n25501 = ~pi660 & ~n25412;
  assign n25502 = ~n25500 & n25501;
  assign n25503 = ~pi609 & ~n25451;
  assign n25504 = pi609 & ~n25497;
  assign n25505 = ~n25503 & ~n25504;
  assign n25506 = pi1155 & n25505;
  assign n25507 = ~n25414 & ~n25506;
  assign n25508 = pi660 & n25507;
  assign n25509 = ~n25502 & ~n25508;
  assign n25510 = pi785 & ~n25509;
  assign n25511 = ~pi785 & ~n25497;
  assign n25512 = ~n25510 & ~n25511;
  assign n25513 = ~pi618 & ~n25512;
  assign n25514 = ~pi1154 & ~n25513;
  assign n25515 = ~n25481 & n25514;
  assign n25516 = ~pi627 & ~n25420;
  assign n25517 = ~n25515 & n25516;
  assign n25518 = ~pi618 & n25452;
  assign n25519 = pi618 & ~n25512;
  assign n25520 = ~n25518 & ~n25519;
  assign n25521 = pi1154 & n25520;
  assign n25522 = ~n25422 & ~n25521;
  assign n25523 = pi627 & n25522;
  assign n25524 = ~n25517 & ~n25523;
  assign n25525 = pi781 & ~n25524;
  assign n25526 = ~pi781 & ~n25512;
  assign n25527 = ~n25525 & ~n25526;
  assign n25528 = ~pi619 & ~n25527;
  assign n25529 = pi619 & n25453;
  assign n25530 = ~pi1159 & ~n25529;
  assign n25531 = ~n25528 & n25530;
  assign n25532 = ~pi648 & ~n25531;
  assign n25533 = ~n25428 & n25532;
  assign n25534 = ~pi619 & n25453;
  assign n25535 = pi619 & ~n25527;
  assign n25536 = ~n25534 & ~n25535;
  assign n25537 = pi1159 & n25536;
  assign n25538 = ~n25430 & ~n25537;
  assign n25539 = pi648 & n25538;
  assign n25540 = ~n25533 & ~n25539;
  assign n25541 = pi789 & n25540;
  assign n25542 = ~pi789 & n25527;
  assign n25543 = n17356 & ~n25542;
  assign n25544 = ~n25541 & n25543;
  assign n25545 = ~n25480 & ~n25544;
  assign n25546 = n19788 & ~n25545;
  assign n25547 = n20275 & n25455;
  assign n25548 = n17449 & ~n25436;
  assign n25549 = ~pi629 & ~n25548;
  assign n25550 = ~n25547 & n25549;
  assign n25551 = n17448 & ~n25436;
  assign n25552 = n20281 & n25455;
  assign n25553 = pi629 & ~n25552;
  assign n25554 = ~n25551 & n25553;
  assign n25555 = ~n25550 & ~n25554;
  assign n25556 = pi792 & n25555;
  assign n25557 = n19637 & ~n25556;
  assign n25558 = ~n25546 & n25557;
  assign n25559 = ~n25468 & ~n25558;
  assign n25560 = pi644 & n25559;
  assign n25561 = ~pi787 & ~n25456;
  assign n25562 = pi787 & ~n25465;
  assign n25563 = ~n25561 & ~n25562;
  assign n25564 = ~pi644 & n25563;
  assign n25565 = pi715 & ~n25564;
  assign n25566 = ~n25560 & n25565;
  assign n25567 = ~n17247 & ~n25439;
  assign n25568 = n17247 & n25405;
  assign n25569 = ~n25567 & ~n25568;
  assign n25570 = pi644 & ~n25569;
  assign n25571 = ~pi644 & n25405;
  assign n25572 = ~pi715 & ~n25571;
  assign n25573 = ~n25570 & n25572;
  assign n25574 = pi1160 & ~n25573;
  assign n25575 = ~n25566 & n25574;
  assign n25576 = ~pi644 & ~n25569;
  assign n25577 = pi715 & ~n25576;
  assign n25578 = pi644 & n25405;
  assign n25579 = n25577 & ~n25578;
  assign n25580 = pi644 & n25563;
  assign n25581 = ~pi644 & n25559;
  assign n25582 = ~pi715 & ~n25581;
  assign n25583 = ~n25580 & n25582;
  assign n25584 = ~pi1160 & ~n25583;
  assign n25585 = ~n25579 & n25584;
  assign n25586 = ~n25575 & ~n25585;
  assign n25587 = pi790 & ~n25586;
  assign n25588 = ~pi790 & n25559;
  assign n25589 = pi832 & ~n25588;
  assign n25590 = ~n25587 & n25589;
  assign n25591 = ~pi180 & ~n16527;
  assign n25592 = n17159 & ~n25591;
  assign n25593 = n16593 & ~n25591;
  assign n25594 = ~pi702 & n10020;
  assign n25595 = n25591 & ~n25594;
  assign n25596 = ~pi180 & n17592;
  assign n25597 = ~pi38 & ~pi180;
  assign n25598 = n19843 & ~n25597;
  assign n25599 = ~n25596 & ~n25598;
  assign n25600 = ~pi180 & ~n16508;
  assign n25601 = n16744 & ~n25600;
  assign n25602 = ~pi702 & ~n25601;
  assign n25603 = ~n25599 & n25602;
  assign n25604 = ~n25595 & ~n25603;
  assign n25605 = ~pi778 & n25604;
  assign n25606 = pi625 & ~n25604;
  assign n25607 = pi1153 & ~n25606;
  assign n25608 = ~pi625 & n25591;
  assign n25609 = n25607 & ~n25608;
  assign n25610 = ~pi625 & ~n25604;
  assign n25611 = ~pi1153 & ~n25610;
  assign n25612 = pi625 & n25591;
  assign n25613 = n25611 & ~n25612;
  assign n25614 = ~n25609 & ~n25613;
  assign n25615 = pi778 & ~n25614;
  assign n25616 = ~n25605 & ~n25615;
  assign n25617 = ~n16593 & ~n25616;
  assign n25618 = ~n25593 & ~n25617;
  assign n25619 = ~n16589 & n25618;
  assign n25620 = n16589 & n25591;
  assign n25621 = ~n25619 & ~n25620;
  assign n25622 = ~n17159 & n25621;
  assign n25623 = ~n25592 & ~n25622;
  assign n25624 = ~n17183 & n25623;
  assign n25625 = n17183 & n25591;
  assign n25626 = ~n25624 & ~n25625;
  assign n25627 = ~pi792 & n25626;
  assign n25628 = pi628 & ~n25626;
  assign n25629 = pi1156 & ~n25628;
  assign n25630 = ~pi628 & n25591;
  assign n25631 = n25629 & ~n25630;
  assign n25632 = ~pi628 & ~n25626;
  assign n25633 = pi628 & n25591;
  assign n25634 = ~pi1156 & ~n25633;
  assign n25635 = ~n25632 & n25634;
  assign n25636 = ~n25631 & ~n25635;
  assign n25637 = pi792 & ~n25636;
  assign n25638 = ~n25627 & ~n25637;
  assign n25639 = pi647 & ~n25638;
  assign n25640 = ~pi647 & ~n25591;
  assign n25641 = ~n25639 & ~n25640;
  assign n25642 = pi1157 & ~n25641;
  assign n25643 = ~pi647 & n25638;
  assign n25644 = ~pi1157 & ~n25643;
  assign n25645 = pi647 & n25591;
  assign n25646 = n25644 & ~n25645;
  assign n25647 = ~n25642 & ~n25646;
  assign n25648 = pi787 & ~n25647;
  assign n25649 = ~pi787 & ~n25638;
  assign n25650 = ~n25648 & ~n25649;
  assign n25651 = ~pi644 & n25650;
  assign n25652 = pi715 & ~n25651;
  assign n25653 = n17247 & ~n25591;
  assign n25654 = pi180 & ~n10020;
  assign n25655 = ~pi753 & n16511;
  assign n25656 = ~n25600 & ~n25655;
  assign n25657 = pi38 & ~n25656;
  assign n25658 = n10020 & ~n25657;
  assign n25659 = pi753 & n16355;
  assign n25660 = pi180 & n16501;
  assign n25661 = ~n25659 & ~n25660;
  assign n25662 = pi39 & ~n25661;
  assign n25663 = pi180 & pi753;
  assign n25664 = pi180 & ~n16460;
  assign n25665 = ~n21155 & ~n25664;
  assign n25666 = ~pi39 & ~n25665;
  assign n25667 = ~n25663 & ~n25666;
  assign n25668 = ~pi180 & ~pi753;
  assign n25669 = n16449 & n25668;
  assign n25670 = n25667 & ~n25669;
  assign n25671 = ~n25662 & n25670;
  assign n25672 = ~pi38 & n25671;
  assign n25673 = n25658 & ~n25672;
  assign n25674 = ~n25654 & ~n25673;
  assign n25675 = ~n16521 & ~n25674;
  assign n25676 = n16521 & ~n25591;
  assign n25677 = ~n25675 & ~n25676;
  assign n25678 = ~pi785 & ~n25677;
  assign n25679 = ~n16532 & ~n25591;
  assign n25680 = pi609 & n25675;
  assign n25681 = ~n25679 & ~n25680;
  assign n25682 = pi1155 & ~n25681;
  assign n25683 = ~n16537 & ~n25591;
  assign n25684 = ~pi609 & n25675;
  assign n25685 = ~n25683 & ~n25684;
  assign n25686 = ~pi1155 & ~n25685;
  assign n25687 = ~n25682 & ~n25686;
  assign n25688 = pi785 & ~n25687;
  assign n25689 = ~n25678 & ~n25688;
  assign n25690 = ~pi781 & ~n25689;
  assign n25691 = pi618 & n25689;
  assign n25692 = ~pi618 & n25591;
  assign n25693 = pi1154 & ~n25692;
  assign n25694 = ~n25691 & n25693;
  assign n25695 = ~pi618 & n25689;
  assign n25696 = pi618 & n25591;
  assign n25697 = ~pi1154 & ~n25696;
  assign n25698 = ~n25695 & n25697;
  assign n25699 = ~n25694 & ~n25698;
  assign n25700 = pi781 & ~n25699;
  assign n25701 = ~n25690 & ~n25700;
  assign n25702 = ~pi789 & ~n25701;
  assign n25703 = pi619 & n25701;
  assign n25704 = ~pi619 & n25591;
  assign n25705 = pi1159 & ~n25704;
  assign n25706 = ~n25703 & n25705;
  assign n25707 = ~pi619 & n25701;
  assign n25708 = pi619 & n25591;
  assign n25709 = ~pi1159 & ~n25708;
  assign n25710 = ~n25707 & n25709;
  assign n25711 = ~n25706 & ~n25710;
  assign n25712 = pi789 & ~n25711;
  assign n25713 = ~n25702 & ~n25712;
  assign n25714 = ~n17355 & n25713;
  assign n25715 = n17355 & n25591;
  assign n25716 = ~n25714 & ~n25715;
  assign n25717 = ~n16124 & ~n25716;
  assign n25718 = n16124 & n25591;
  assign n25719 = ~n25717 & ~n25718;
  assign n25720 = ~n17247 & n25719;
  assign n25721 = ~n25653 & ~n25720;
  assign n25722 = pi644 & n25721;
  assign n25723 = ~pi644 & n25591;
  assign n25724 = ~pi715 & ~n25723;
  assign n25725 = ~n25722 & n25724;
  assign n25726 = pi1160 & ~n25725;
  assign n25727 = ~n25652 & n25726;
  assign n25728 = pi644 & n25650;
  assign n25729 = ~pi715 & ~n25728;
  assign n25730 = ~pi644 & n25721;
  assign n25731 = pi644 & n25591;
  assign n25732 = ~n25730 & ~n25731;
  assign n25733 = pi715 & n25732;
  assign n25734 = ~pi1160 & ~n25733;
  assign n25735 = ~n25729 & n25734;
  assign n25736 = ~n25727 & ~n25735;
  assign n25737 = pi790 & ~n25736;
  assign n25738 = ~pi629 & n25631;
  assign n25739 = ~n19999 & n25716;
  assign n25740 = pi629 & n25635;
  assign n25741 = ~n25739 & ~n25740;
  assign n25742 = ~n25738 & n25741;
  assign n25743 = pi792 & ~n25742;
  assign n25744 = pi618 & n25618;
  assign n25745 = pi609 & n25616;
  assign n25746 = pi625 & n25674;
  assign n25747 = ~n25594 & ~n25673;
  assign n25748 = ~pi753 & ~n16917;
  assign n25749 = n18933 & ~n25748;
  assign n25750 = ~pi180 & ~n25749;
  assign n25751 = ~n17079 & ~n25406;
  assign n25752 = pi180 & ~n25751;
  assign n25753 = n6097 & n25752;
  assign n25754 = ~n25750 & ~n25753;
  assign n25755 = pi38 & n25754;
  assign n25756 = ~pi180 & n16853;
  assign n25757 = pi180 & n16935;
  assign n25758 = pi753 & ~n25757;
  assign n25759 = ~n25756 & n25758;
  assign n25760 = pi180 & n16998;
  assign n25761 = ~pi180 & ~n17051;
  assign n25762 = ~pi753 & ~n25761;
  assign n25763 = ~n25760 & n25762;
  assign n25764 = ~n25759 & ~n25763;
  assign n25765 = pi39 & n25764;
  assign n25766 = ~pi180 & ~n17061;
  assign n25767 = pi180 & ~n17058;
  assign n25768 = pi753 & ~n25767;
  assign n25769 = ~n25766 & n25768;
  assign n25770 = ~pi180 & n17067;
  assign n25771 = ~pi753 & ~n25770;
  assign n25772 = pi180 & n17065;
  assign n25773 = n25771 & ~n25772;
  assign n25774 = ~n25769 & ~n25773;
  assign n25775 = ~pi39 & ~n25774;
  assign n25776 = ~pi38 & ~n25775;
  assign n25777 = ~n25765 & n25776;
  assign n25778 = ~pi702 & ~n25777;
  assign n25779 = ~n25755 & n25778;
  assign n25780 = ~n25747 & ~n25779;
  assign n25781 = ~n25654 & ~n25780;
  assign n25782 = ~pi625 & n25781;
  assign n25783 = ~pi1153 & ~n25782;
  assign n25784 = ~n25746 & n25783;
  assign n25785 = ~pi608 & ~n25609;
  assign n25786 = ~n25784 & n25785;
  assign n25787 = ~pi625 & n25674;
  assign n25788 = pi625 & n25781;
  assign n25789 = ~n25787 & ~n25788;
  assign n25790 = pi1153 & n25789;
  assign n25791 = ~n25613 & ~n25790;
  assign n25792 = pi608 & n25791;
  assign n25793 = ~n25786 & ~n25792;
  assign n25794 = pi778 & ~n25793;
  assign n25795 = ~pi778 & n25781;
  assign n25796 = ~n25794 & ~n25795;
  assign n25797 = ~pi609 & ~n25796;
  assign n25798 = ~pi1155 & ~n25797;
  assign n25799 = ~n25745 & n25798;
  assign n25800 = ~pi660 & ~n25682;
  assign n25801 = ~n25799 & n25800;
  assign n25802 = ~pi609 & n25616;
  assign n25803 = pi609 & ~n25796;
  assign n25804 = ~n25802 & ~n25803;
  assign n25805 = pi1155 & n25804;
  assign n25806 = ~n25686 & ~n25805;
  assign n25807 = pi660 & n25806;
  assign n25808 = ~n25801 & ~n25807;
  assign n25809 = pi785 & ~n25808;
  assign n25810 = ~pi785 & ~n25796;
  assign n25811 = ~n25809 & ~n25810;
  assign n25812 = ~pi618 & ~n25811;
  assign n25813 = ~pi1154 & ~n25812;
  assign n25814 = ~n25744 & n25813;
  assign n25815 = ~pi627 & ~n25694;
  assign n25816 = ~n25814 & n25815;
  assign n25817 = ~pi618 & n25618;
  assign n25818 = pi618 & ~n25811;
  assign n25819 = ~n25817 & ~n25818;
  assign n25820 = pi1154 & n25819;
  assign n25821 = ~n25698 & ~n25820;
  assign n25822 = pi627 & n25821;
  assign n25823 = ~n25816 & ~n25822;
  assign n25824 = pi781 & ~n25823;
  assign n25825 = ~pi781 & ~n25811;
  assign n25826 = ~n25824 & ~n25825;
  assign n25827 = ~pi789 & n25826;
  assign n25828 = ~pi619 & ~n25826;
  assign n25829 = pi619 & ~n25621;
  assign n25830 = ~pi1159 & ~n25829;
  assign n25831 = ~n25828 & n25830;
  assign n25832 = ~pi648 & ~n25831;
  assign n25833 = ~n25706 & n25832;
  assign n25834 = ~pi619 & ~n25621;
  assign n25835 = pi619 & ~n25826;
  assign n25836 = ~n25834 & ~n25835;
  assign n25837 = pi1159 & n25836;
  assign n25838 = ~n25710 & ~n25837;
  assign n25839 = pi648 & n25838;
  assign n25840 = ~n25833 & ~n25839;
  assign n25841 = pi789 & n25840;
  assign n25842 = ~n25827 & ~n25841;
  assign n25843 = n17356 & n25842;
  assign n25844 = ~pi626 & ~n25713;
  assign n25845 = pi626 & ~n25591;
  assign n25846 = n17181 & ~n25845;
  assign n25847 = ~n25844 & n25846;
  assign n25848 = n17350 & n25623;
  assign n25849 = pi626 & ~n25713;
  assign n25850 = ~pi626 & ~n25591;
  assign n25851 = n17180 & ~n25850;
  assign n25852 = ~n25849 & n25851;
  assign n25853 = ~n25848 & ~n25852;
  assign n25854 = ~n25847 & n25853;
  assign n25855 = pi788 & ~n25854;
  assign n25856 = n19788 & ~n25855;
  assign n25857 = ~n25843 & n25856;
  assign n25858 = ~n25743 & ~n25857;
  assign n25859 = n19637 & ~n25858;
  assign n25860 = ~n19987 & n25719;
  assign n25861 = pi630 & n25646;
  assign n25862 = ~n25860 & ~n25861;
  assign n25863 = n17244 & ~n25641;
  assign n25864 = n25862 & ~n25863;
  assign n25865 = pi787 & ~n25864;
  assign n25866 = ~n25859 & ~n25865;
  assign n25867 = pi644 & n25726;
  assign n25868 = ~pi644 & n25734;
  assign n25869 = pi790 & ~n25868;
  assign n25870 = ~n25867 & n25869;
  assign n25871 = n25866 & ~n25870;
  assign n25872 = ~n25737 & ~n25871;
  assign n25873 = ~po1038 & ~n25872;
  assign n25874 = ~pi180 & po1038;
  assign n25875 = ~pi832 & ~n25874;
  assign n25876 = ~n25873 & n25875;
  assign po337 = ~n25590 & ~n25876;
  assign n25878 = ~pi181 & ~n2934;
  assign n25879 = ~pi754 & n16510;
  assign n25880 = ~n25878 & ~n25879;
  assign n25881 = ~n17273 & ~n25880;
  assign n25882 = ~pi785 & ~n25881;
  assign n25883 = n16537 & n25879;
  assign n25884 = n25881 & ~n25883;
  assign n25885 = pi1155 & ~n25884;
  assign n25886 = ~pi1155 & ~n25878;
  assign n25887 = ~n25883 & n25886;
  assign n25888 = ~n25885 & ~n25887;
  assign n25889 = pi785 & ~n25888;
  assign n25890 = ~n25882 & ~n25889;
  assign n25891 = ~pi781 & ~n25890;
  assign n25892 = ~n17289 & n25890;
  assign n25893 = pi1154 & ~n25892;
  assign n25894 = ~n17292 & n25890;
  assign n25895 = ~pi1154 & ~n25894;
  assign n25896 = ~n25893 & ~n25895;
  assign n25897 = pi781 & ~n25896;
  assign n25898 = ~n25891 & ~n25897;
  assign n25899 = ~pi789 & ~n25898;
  assign n25900 = ~n22423 & n25898;
  assign n25901 = pi1159 & ~n25900;
  assign n25902 = ~n22426 & n25898;
  assign n25903 = ~pi1159 & ~n25902;
  assign n25904 = ~n25901 & ~n25903;
  assign n25905 = pi789 & ~n25904;
  assign n25906 = ~n25899 & ~n25905;
  assign n25907 = ~n17355 & n25906;
  assign n25908 = n17355 & n25878;
  assign n25909 = ~n25907 & ~n25908;
  assign n25910 = ~n16124 & ~n25909;
  assign n25911 = n16124 & n25878;
  assign n25912 = ~n25910 & ~n25911;
  assign n25913 = ~n19987 & n25912;
  assign n25914 = ~pi709 & n16742;
  assign n25915 = ~n25878 & ~n25914;
  assign n25916 = ~pi778 & ~n25915;
  assign n25917 = ~pi625 & n25914;
  assign n25918 = ~n25915 & ~n25917;
  assign n25919 = pi1153 & ~n25918;
  assign n25920 = ~pi1153 & ~n25878;
  assign n25921 = ~n25917 & n25920;
  assign n25922 = ~n25919 & ~n25921;
  assign n25923 = pi778 & n25922;
  assign n25924 = ~n25916 & ~n25923;
  assign n25925 = ~n17338 & ~n25924;
  assign n25926 = ~n17340 & n25925;
  assign n25927 = ~n17342 & n25926;
  assign n25928 = ~n17425 & n25927;
  assign n25929 = ~n17452 & n25928;
  assign n25930 = ~pi647 & n25929;
  assign n25931 = pi647 & n25878;
  assign n25932 = ~pi1157 & ~n25931;
  assign n25933 = ~n25930 & n25932;
  assign n25934 = ~pi647 & n25878;
  assign n25935 = pi647 & n25929;
  assign n25936 = pi1157 & ~n25935;
  assign n25937 = ~n25934 & n25936;
  assign n25938 = ~n25933 & ~n25937;
  assign n25939 = ~n17246 & ~n25938;
  assign n25940 = ~n25913 & ~n25939;
  assign n25941 = pi787 & ~n25940;
  assign n25942 = ~pi626 & ~n25906;
  assign n25943 = pi626 & ~n25878;
  assign n25944 = n17181 & ~n25943;
  assign n25945 = ~n25942 & n25944;
  assign n25946 = n17350 & n25927;
  assign n25947 = pi626 & ~n25906;
  assign n25948 = ~pi626 & ~n25878;
  assign n25949 = n17180 & ~n25948;
  assign n25950 = ~n25947 & n25949;
  assign n25951 = ~n25946 & ~n25950;
  assign n25952 = ~n25945 & n25951;
  assign n25953 = pi788 & ~n25952;
  assign n25954 = pi618 & n25925;
  assign n25955 = pi609 & ~n25924;
  assign n25956 = ~n16393 & ~n25915;
  assign n25957 = pi625 & n25956;
  assign n25958 = n25880 & ~n25956;
  assign n25959 = ~n25957 & ~n25958;
  assign n25960 = n25920 & ~n25959;
  assign n25961 = ~pi608 & ~n25919;
  assign n25962 = ~n25960 & n25961;
  assign n25963 = pi1153 & ~n25957;
  assign n25964 = n25880 & n25963;
  assign n25965 = ~n25921 & ~n25964;
  assign n25966 = pi608 & n25965;
  assign n25967 = ~n25962 & ~n25966;
  assign n25968 = pi778 & ~n25967;
  assign n25969 = ~pi778 & ~n25958;
  assign n25970 = ~n25968 & ~n25969;
  assign n25971 = ~pi609 & ~n25970;
  assign n25972 = ~pi1155 & ~n25971;
  assign n25973 = ~n25955 & n25972;
  assign n25974 = ~pi660 & ~n25885;
  assign n25975 = ~n25973 & n25974;
  assign n25976 = ~pi609 & ~n25924;
  assign n25977 = pi609 & ~n25970;
  assign n25978 = ~n25976 & ~n25977;
  assign n25979 = pi1155 & n25978;
  assign n25980 = ~n25887 & ~n25979;
  assign n25981 = pi660 & n25980;
  assign n25982 = ~n25975 & ~n25981;
  assign n25983 = pi785 & ~n25982;
  assign n25984 = ~pi785 & ~n25970;
  assign n25985 = ~n25983 & ~n25984;
  assign n25986 = ~pi618 & ~n25985;
  assign n25987 = ~pi1154 & ~n25986;
  assign n25988 = ~n25954 & n25987;
  assign n25989 = ~pi627 & ~n25893;
  assign n25990 = ~n25988 & n25989;
  assign n25991 = ~pi618 & n25925;
  assign n25992 = pi618 & ~n25985;
  assign n25993 = ~n25991 & ~n25992;
  assign n25994 = pi1154 & n25993;
  assign n25995 = ~n25895 & ~n25994;
  assign n25996 = pi627 & n25995;
  assign n25997 = ~n25990 & ~n25996;
  assign n25998 = pi781 & ~n25997;
  assign n25999 = ~pi781 & ~n25985;
  assign n26000 = ~n25998 & ~n25999;
  assign n26001 = ~pi619 & ~n26000;
  assign n26002 = pi619 & n25926;
  assign n26003 = ~pi1159 & ~n26002;
  assign n26004 = ~n26001 & n26003;
  assign n26005 = ~pi648 & ~n26004;
  assign n26006 = ~n25901 & n26005;
  assign n26007 = ~pi619 & n25926;
  assign n26008 = pi619 & ~n26000;
  assign n26009 = ~n26007 & ~n26008;
  assign n26010 = pi1159 & n26009;
  assign n26011 = ~n25903 & ~n26010;
  assign n26012 = pi648 & n26011;
  assign n26013 = ~n26006 & ~n26012;
  assign n26014 = pi789 & n26013;
  assign n26015 = ~pi789 & n26000;
  assign n26016 = n17356 & ~n26015;
  assign n26017 = ~n26014 & n26016;
  assign n26018 = ~n25953 & ~n26017;
  assign n26019 = n19788 & ~n26018;
  assign n26020 = n20275 & n25928;
  assign n26021 = n17449 & ~n25909;
  assign n26022 = ~pi629 & ~n26021;
  assign n26023 = ~n26020 & n26022;
  assign n26024 = n17448 & ~n25909;
  assign n26025 = n20281 & n25928;
  assign n26026 = pi629 & ~n26025;
  assign n26027 = ~n26024 & n26026;
  assign n26028 = ~n26023 & ~n26027;
  assign n26029 = pi792 & n26028;
  assign n26030 = n19637 & ~n26029;
  assign n26031 = ~n26019 & n26030;
  assign n26032 = ~n25941 & ~n26031;
  assign n26033 = pi644 & n26032;
  assign n26034 = ~pi787 & ~n25929;
  assign n26035 = pi787 & ~n25938;
  assign n26036 = ~n26034 & ~n26035;
  assign n26037 = ~pi644 & n26036;
  assign n26038 = pi715 & ~n26037;
  assign n26039 = ~n26033 & n26038;
  assign n26040 = ~n17247 & ~n25912;
  assign n26041 = n17247 & n25878;
  assign n26042 = ~n26040 & ~n26041;
  assign n26043 = pi644 & ~n26042;
  assign n26044 = ~pi644 & n25878;
  assign n26045 = ~pi715 & ~n26044;
  assign n26046 = ~n26043 & n26045;
  assign n26047 = pi1160 & ~n26046;
  assign n26048 = ~n26039 & n26047;
  assign n26049 = ~pi644 & ~n26042;
  assign n26050 = pi715 & ~n26049;
  assign n26051 = pi644 & n25878;
  assign n26052 = n26050 & ~n26051;
  assign n26053 = pi644 & n26036;
  assign n26054 = ~pi644 & n26032;
  assign n26055 = ~pi715 & ~n26054;
  assign n26056 = ~n26053 & n26055;
  assign n26057 = ~pi1160 & ~n26056;
  assign n26058 = ~n26052 & n26057;
  assign n26059 = ~n26048 & ~n26058;
  assign n26060 = pi790 & ~n26059;
  assign n26061 = ~pi790 & n26032;
  assign n26062 = pi832 & ~n26061;
  assign n26063 = ~n26060 & n26062;
  assign n26064 = ~pi181 & ~n16527;
  assign n26065 = n17159 & ~n26064;
  assign n26066 = n16593 & ~n26064;
  assign n26067 = ~pi709 & n10020;
  assign n26068 = n26064 & ~n26067;
  assign n26069 = ~pi181 & n17592;
  assign n26070 = ~pi38 & ~pi181;
  assign n26071 = n19843 & ~n26070;
  assign n26072 = ~n26069 & ~n26071;
  assign n26073 = ~pi181 & ~n16508;
  assign n26074 = n16744 & ~n26073;
  assign n26075 = ~pi709 & ~n26074;
  assign n26076 = ~n26072 & n26075;
  assign n26077 = ~n26068 & ~n26076;
  assign n26078 = ~pi778 & n26077;
  assign n26079 = pi625 & ~n26077;
  assign n26080 = pi1153 & ~n26079;
  assign n26081 = ~pi625 & n26064;
  assign n26082 = n26080 & ~n26081;
  assign n26083 = ~pi625 & ~n26077;
  assign n26084 = ~pi1153 & ~n26083;
  assign n26085 = pi625 & n26064;
  assign n26086 = n26084 & ~n26085;
  assign n26087 = ~n26082 & ~n26086;
  assign n26088 = pi778 & ~n26087;
  assign n26089 = ~n26078 & ~n26088;
  assign n26090 = ~n16593 & ~n26089;
  assign n26091 = ~n26066 & ~n26090;
  assign n26092 = ~n16589 & n26091;
  assign n26093 = n16589 & n26064;
  assign n26094 = ~n26092 & ~n26093;
  assign n26095 = ~n17159 & n26094;
  assign n26096 = ~n26065 & ~n26095;
  assign n26097 = ~n17183 & n26096;
  assign n26098 = n17183 & n26064;
  assign n26099 = ~n26097 & ~n26098;
  assign n26100 = ~pi792 & n26099;
  assign n26101 = pi628 & ~n26099;
  assign n26102 = pi1156 & ~n26101;
  assign n26103 = ~pi628 & n26064;
  assign n26104 = n26102 & ~n26103;
  assign n26105 = ~pi628 & ~n26099;
  assign n26106 = pi628 & n26064;
  assign n26107 = ~pi1156 & ~n26106;
  assign n26108 = ~n26105 & n26107;
  assign n26109 = ~n26104 & ~n26108;
  assign n26110 = pi792 & ~n26109;
  assign n26111 = ~n26100 & ~n26110;
  assign n26112 = pi647 & ~n26111;
  assign n26113 = ~pi647 & ~n26064;
  assign n26114 = ~n26112 & ~n26113;
  assign n26115 = pi1157 & ~n26114;
  assign n26116 = ~pi647 & n26111;
  assign n26117 = ~pi1157 & ~n26116;
  assign n26118 = pi647 & n26064;
  assign n26119 = n26117 & ~n26118;
  assign n26120 = ~n26115 & ~n26119;
  assign n26121 = pi787 & ~n26120;
  assign n26122 = ~pi787 & ~n26111;
  assign n26123 = ~n26121 & ~n26122;
  assign n26124 = ~pi644 & n26123;
  assign n26125 = pi715 & ~n26124;
  assign n26126 = n17247 & ~n26064;
  assign n26127 = pi181 & ~n10020;
  assign n26128 = ~pi754 & n16511;
  assign n26129 = ~n26073 & ~n26128;
  assign n26130 = pi38 & ~n26129;
  assign n26131 = n10020 & ~n26130;
  assign n26132 = pi754 & n16355;
  assign n26133 = pi181 & n16501;
  assign n26134 = ~n26132 & ~n26133;
  assign n26135 = pi39 & ~n26134;
  assign n26136 = pi181 & pi754;
  assign n26137 = pi181 & ~n16460;
  assign n26138 = ~n21208 & ~n26137;
  assign n26139 = ~pi39 & ~n26138;
  assign n26140 = ~n26136 & ~n26139;
  assign n26141 = ~pi181 & ~pi754;
  assign n26142 = n16449 & n26141;
  assign n26143 = n26140 & ~n26142;
  assign n26144 = ~n26135 & n26143;
  assign n26145 = ~pi38 & n26144;
  assign n26146 = n26131 & ~n26145;
  assign n26147 = ~n26127 & ~n26146;
  assign n26148 = ~n16521 & ~n26147;
  assign n26149 = n16521 & ~n26064;
  assign n26150 = ~n26148 & ~n26149;
  assign n26151 = ~pi785 & ~n26150;
  assign n26152 = ~n16532 & ~n26064;
  assign n26153 = pi609 & n26148;
  assign n26154 = ~n26152 & ~n26153;
  assign n26155 = pi1155 & ~n26154;
  assign n26156 = ~n16537 & ~n26064;
  assign n26157 = ~pi609 & n26148;
  assign n26158 = ~n26156 & ~n26157;
  assign n26159 = ~pi1155 & ~n26158;
  assign n26160 = ~n26155 & ~n26159;
  assign n26161 = pi785 & ~n26160;
  assign n26162 = ~n26151 & ~n26161;
  assign n26163 = ~pi781 & ~n26162;
  assign n26164 = pi618 & n26162;
  assign n26165 = ~pi618 & n26064;
  assign n26166 = pi1154 & ~n26165;
  assign n26167 = ~n26164 & n26166;
  assign n26168 = ~pi618 & n26162;
  assign n26169 = pi618 & n26064;
  assign n26170 = ~pi1154 & ~n26169;
  assign n26171 = ~n26168 & n26170;
  assign n26172 = ~n26167 & ~n26171;
  assign n26173 = pi781 & ~n26172;
  assign n26174 = ~n26163 & ~n26173;
  assign n26175 = ~pi789 & ~n26174;
  assign n26176 = pi619 & n26174;
  assign n26177 = ~pi619 & n26064;
  assign n26178 = pi1159 & ~n26177;
  assign n26179 = ~n26176 & n26178;
  assign n26180 = ~pi619 & n26174;
  assign n26181 = pi619 & n26064;
  assign n26182 = ~pi1159 & ~n26181;
  assign n26183 = ~n26180 & n26182;
  assign n26184 = ~n26179 & ~n26183;
  assign n26185 = pi789 & ~n26184;
  assign n26186 = ~n26175 & ~n26185;
  assign n26187 = ~n17355 & n26186;
  assign n26188 = n17355 & n26064;
  assign n26189 = ~n26187 & ~n26188;
  assign n26190 = ~n16124 & ~n26189;
  assign n26191 = n16124 & n26064;
  assign n26192 = ~n26190 & ~n26191;
  assign n26193 = ~n17247 & n26192;
  assign n26194 = ~n26126 & ~n26193;
  assign n26195 = pi644 & n26194;
  assign n26196 = ~pi644 & n26064;
  assign n26197 = ~pi715 & ~n26196;
  assign n26198 = ~n26195 & n26197;
  assign n26199 = pi1160 & ~n26198;
  assign n26200 = ~n26125 & n26199;
  assign n26201 = pi644 & n26123;
  assign n26202 = ~pi715 & ~n26201;
  assign n26203 = ~pi644 & n26194;
  assign n26204 = pi644 & n26064;
  assign n26205 = ~n26203 & ~n26204;
  assign n26206 = pi715 & n26205;
  assign n26207 = ~pi1160 & ~n26206;
  assign n26208 = ~n26202 & n26207;
  assign n26209 = ~n26200 & ~n26208;
  assign n26210 = pi790 & ~n26209;
  assign n26211 = ~pi629 & n26104;
  assign n26212 = ~n19999 & n26189;
  assign n26213 = pi629 & n26108;
  assign n26214 = ~n26212 & ~n26213;
  assign n26215 = ~n26211 & n26214;
  assign n26216 = pi792 & ~n26215;
  assign n26217 = pi618 & n26091;
  assign n26218 = pi609 & n26089;
  assign n26219 = pi625 & n26147;
  assign n26220 = ~n26067 & ~n26146;
  assign n26221 = ~pi754 & ~n16917;
  assign n26222 = n18933 & ~n26221;
  assign n26223 = ~pi181 & ~n26222;
  assign n26224 = ~n17079 & ~n25879;
  assign n26225 = pi181 & ~n26224;
  assign n26226 = n6097 & n26225;
  assign n26227 = ~n26223 & ~n26226;
  assign n26228 = pi38 & n26227;
  assign n26229 = ~pi181 & n16853;
  assign n26230 = pi181 & n16935;
  assign n26231 = pi754 & ~n26230;
  assign n26232 = ~n26229 & n26231;
  assign n26233 = pi181 & n16998;
  assign n26234 = ~pi181 & ~n17051;
  assign n26235 = ~pi754 & ~n26234;
  assign n26236 = ~n26233 & n26235;
  assign n26237 = ~n26232 & ~n26236;
  assign n26238 = pi39 & n26237;
  assign n26239 = ~pi181 & ~n17061;
  assign n26240 = pi181 & ~n17058;
  assign n26241 = pi754 & ~n26240;
  assign n26242 = ~n26239 & n26241;
  assign n26243 = ~pi181 & n17067;
  assign n26244 = ~pi754 & ~n26243;
  assign n26245 = pi181 & n17065;
  assign n26246 = n26244 & ~n26245;
  assign n26247 = ~n26242 & ~n26246;
  assign n26248 = ~pi39 & ~n26247;
  assign n26249 = ~pi38 & ~n26248;
  assign n26250 = ~n26238 & n26249;
  assign n26251 = ~pi709 & ~n26250;
  assign n26252 = ~n26228 & n26251;
  assign n26253 = ~n26220 & ~n26252;
  assign n26254 = ~n26127 & ~n26253;
  assign n26255 = ~pi625 & n26254;
  assign n26256 = ~pi1153 & ~n26255;
  assign n26257 = ~n26219 & n26256;
  assign n26258 = ~pi608 & ~n26082;
  assign n26259 = ~n26257 & n26258;
  assign n26260 = ~pi625 & n26147;
  assign n26261 = pi625 & n26254;
  assign n26262 = ~n26260 & ~n26261;
  assign n26263 = pi1153 & n26262;
  assign n26264 = ~n26086 & ~n26263;
  assign n26265 = pi608 & n26264;
  assign n26266 = ~n26259 & ~n26265;
  assign n26267 = pi778 & ~n26266;
  assign n26268 = ~pi778 & n26254;
  assign n26269 = ~n26267 & ~n26268;
  assign n26270 = ~pi609 & ~n26269;
  assign n26271 = ~pi1155 & ~n26270;
  assign n26272 = ~n26218 & n26271;
  assign n26273 = ~pi660 & ~n26155;
  assign n26274 = ~n26272 & n26273;
  assign n26275 = ~pi609 & n26089;
  assign n26276 = pi609 & ~n26269;
  assign n26277 = ~n26275 & ~n26276;
  assign n26278 = pi1155 & n26277;
  assign n26279 = ~n26159 & ~n26278;
  assign n26280 = pi660 & n26279;
  assign n26281 = ~n26274 & ~n26280;
  assign n26282 = pi785 & ~n26281;
  assign n26283 = ~pi785 & ~n26269;
  assign n26284 = ~n26282 & ~n26283;
  assign n26285 = ~pi618 & ~n26284;
  assign n26286 = ~pi1154 & ~n26285;
  assign n26287 = ~n26217 & n26286;
  assign n26288 = ~pi627 & ~n26167;
  assign n26289 = ~n26287 & n26288;
  assign n26290 = ~pi618 & n26091;
  assign n26291 = pi618 & ~n26284;
  assign n26292 = ~n26290 & ~n26291;
  assign n26293 = pi1154 & n26292;
  assign n26294 = ~n26171 & ~n26293;
  assign n26295 = pi627 & n26294;
  assign n26296 = ~n26289 & ~n26295;
  assign n26297 = pi781 & ~n26296;
  assign n26298 = ~pi781 & ~n26284;
  assign n26299 = ~n26297 & ~n26298;
  assign n26300 = ~pi789 & n26299;
  assign n26301 = ~pi619 & ~n26299;
  assign n26302 = pi619 & ~n26094;
  assign n26303 = ~pi1159 & ~n26302;
  assign n26304 = ~n26301 & n26303;
  assign n26305 = ~pi648 & ~n26304;
  assign n26306 = ~n26179 & n26305;
  assign n26307 = ~pi619 & ~n26094;
  assign n26308 = pi619 & ~n26299;
  assign n26309 = ~n26307 & ~n26308;
  assign n26310 = pi1159 & n26309;
  assign n26311 = ~n26183 & ~n26310;
  assign n26312 = pi648 & n26311;
  assign n26313 = ~n26306 & ~n26312;
  assign n26314 = pi789 & n26313;
  assign n26315 = ~n26300 & ~n26314;
  assign n26316 = n17356 & n26315;
  assign n26317 = ~pi626 & ~n26186;
  assign n26318 = pi626 & ~n26064;
  assign n26319 = n17181 & ~n26318;
  assign n26320 = ~n26317 & n26319;
  assign n26321 = n17350 & n26096;
  assign n26322 = pi626 & ~n26186;
  assign n26323 = ~pi626 & ~n26064;
  assign n26324 = n17180 & ~n26323;
  assign n26325 = ~n26322 & n26324;
  assign n26326 = ~n26321 & ~n26325;
  assign n26327 = ~n26320 & n26326;
  assign n26328 = pi788 & ~n26327;
  assign n26329 = n19788 & ~n26328;
  assign n26330 = ~n26316 & n26329;
  assign n26331 = ~n26216 & ~n26330;
  assign n26332 = n19637 & ~n26331;
  assign n26333 = ~n19987 & n26192;
  assign n26334 = pi630 & n26119;
  assign n26335 = ~n26333 & ~n26334;
  assign n26336 = n17244 & ~n26114;
  assign n26337 = n26335 & ~n26336;
  assign n26338 = pi787 & ~n26337;
  assign n26339 = ~n26332 & ~n26338;
  assign n26340 = pi644 & n26199;
  assign n26341 = ~pi644 & n26207;
  assign n26342 = pi790 & ~n26341;
  assign n26343 = ~n26340 & n26342;
  assign n26344 = n26339 & ~n26343;
  assign n26345 = ~n26210 & ~n26344;
  assign n26346 = ~po1038 & ~n26345;
  assign n26347 = ~pi181 & po1038;
  assign n26348 = ~pi832 & ~n26347;
  assign n26349 = ~n26346 & n26348;
  assign po338 = ~n26063 & ~n26349;
  assign n26351 = ~pi182 & ~n2934;
  assign n26352 = ~pi756 & n16510;
  assign n26353 = ~n26351 & ~n26352;
  assign n26354 = ~n17273 & ~n26353;
  assign n26355 = ~pi785 & ~n26354;
  assign n26356 = n16537 & n26352;
  assign n26357 = n26354 & ~n26356;
  assign n26358 = pi1155 & ~n26357;
  assign n26359 = ~pi1155 & ~n26351;
  assign n26360 = ~n26356 & n26359;
  assign n26361 = ~n26358 & ~n26360;
  assign n26362 = pi785 & ~n26361;
  assign n26363 = ~n26355 & ~n26362;
  assign n26364 = ~pi781 & ~n26363;
  assign n26365 = ~n17289 & n26363;
  assign n26366 = pi1154 & ~n26365;
  assign n26367 = ~n17292 & n26363;
  assign n26368 = ~pi1154 & ~n26367;
  assign n26369 = ~n26366 & ~n26368;
  assign n26370 = pi781 & ~n26369;
  assign n26371 = ~n26364 & ~n26370;
  assign n26372 = ~pi789 & ~n26371;
  assign n26373 = ~n22423 & n26371;
  assign n26374 = pi1159 & ~n26373;
  assign n26375 = ~n22426 & n26371;
  assign n26376 = ~pi1159 & ~n26375;
  assign n26377 = ~n26374 & ~n26376;
  assign n26378 = pi789 & ~n26377;
  assign n26379 = ~n26372 & ~n26378;
  assign n26380 = ~n17355 & n26379;
  assign n26381 = n17355 & n26351;
  assign n26382 = ~n26380 & ~n26381;
  assign n26383 = ~n16124 & ~n26382;
  assign n26384 = n16124 & n26351;
  assign n26385 = ~n26383 & ~n26384;
  assign n26386 = ~n19987 & n26385;
  assign n26387 = ~pi734 & n16742;
  assign n26388 = ~n26351 & ~n26387;
  assign n26389 = ~pi778 & ~n26388;
  assign n26390 = ~pi625 & n26387;
  assign n26391 = ~n26388 & ~n26390;
  assign n26392 = pi1153 & ~n26391;
  assign n26393 = ~pi1153 & ~n26351;
  assign n26394 = ~n26390 & n26393;
  assign n26395 = ~n26392 & ~n26394;
  assign n26396 = pi778 & n26395;
  assign n26397 = ~n26389 & ~n26396;
  assign n26398 = ~n17338 & ~n26397;
  assign n26399 = ~n17340 & n26398;
  assign n26400 = ~n17342 & n26399;
  assign n26401 = ~n17425 & n26400;
  assign n26402 = ~n17452 & n26401;
  assign n26403 = ~pi647 & n26402;
  assign n26404 = pi647 & n26351;
  assign n26405 = ~pi1157 & ~n26404;
  assign n26406 = ~n26403 & n26405;
  assign n26407 = ~pi647 & n26351;
  assign n26408 = pi647 & n26402;
  assign n26409 = pi1157 & ~n26408;
  assign n26410 = ~n26407 & n26409;
  assign n26411 = ~n26406 & ~n26410;
  assign n26412 = ~n17246 & ~n26411;
  assign n26413 = ~n26386 & ~n26412;
  assign n26414 = pi787 & ~n26413;
  assign n26415 = ~pi626 & ~n26379;
  assign n26416 = pi626 & ~n26351;
  assign n26417 = n17181 & ~n26416;
  assign n26418 = ~n26415 & n26417;
  assign n26419 = n17350 & n26400;
  assign n26420 = pi626 & ~n26379;
  assign n26421 = ~pi626 & ~n26351;
  assign n26422 = n17180 & ~n26421;
  assign n26423 = ~n26420 & n26422;
  assign n26424 = ~n26419 & ~n26423;
  assign n26425 = ~n26418 & n26424;
  assign n26426 = pi788 & ~n26425;
  assign n26427 = pi618 & n26398;
  assign n26428 = pi609 & ~n26397;
  assign n26429 = ~n16393 & ~n26388;
  assign n26430 = pi625 & n26429;
  assign n26431 = n26353 & ~n26429;
  assign n26432 = ~n26430 & ~n26431;
  assign n26433 = n26393 & ~n26432;
  assign n26434 = ~pi608 & ~n26392;
  assign n26435 = ~n26433 & n26434;
  assign n26436 = pi1153 & ~n26430;
  assign n26437 = n26353 & n26436;
  assign n26438 = ~n26394 & ~n26437;
  assign n26439 = pi608 & n26438;
  assign n26440 = ~n26435 & ~n26439;
  assign n26441 = pi778 & ~n26440;
  assign n26442 = ~pi778 & ~n26431;
  assign n26443 = ~n26441 & ~n26442;
  assign n26444 = ~pi609 & ~n26443;
  assign n26445 = ~pi1155 & ~n26444;
  assign n26446 = ~n26428 & n26445;
  assign n26447 = ~pi660 & ~n26358;
  assign n26448 = ~n26446 & n26447;
  assign n26449 = ~pi609 & ~n26397;
  assign n26450 = pi609 & ~n26443;
  assign n26451 = ~n26449 & ~n26450;
  assign n26452 = pi1155 & n26451;
  assign n26453 = ~n26360 & ~n26452;
  assign n26454 = pi660 & n26453;
  assign n26455 = ~n26448 & ~n26454;
  assign n26456 = pi785 & ~n26455;
  assign n26457 = ~pi785 & ~n26443;
  assign n26458 = ~n26456 & ~n26457;
  assign n26459 = ~pi618 & ~n26458;
  assign n26460 = ~pi1154 & ~n26459;
  assign n26461 = ~n26427 & n26460;
  assign n26462 = ~pi627 & ~n26366;
  assign n26463 = ~n26461 & n26462;
  assign n26464 = ~pi618 & n26398;
  assign n26465 = pi618 & ~n26458;
  assign n26466 = ~n26464 & ~n26465;
  assign n26467 = pi1154 & n26466;
  assign n26468 = ~n26368 & ~n26467;
  assign n26469 = pi627 & n26468;
  assign n26470 = ~n26463 & ~n26469;
  assign n26471 = pi781 & ~n26470;
  assign n26472 = ~pi781 & ~n26458;
  assign n26473 = ~n26471 & ~n26472;
  assign n26474 = ~pi619 & ~n26473;
  assign n26475 = pi619 & n26399;
  assign n26476 = ~pi1159 & ~n26475;
  assign n26477 = ~n26474 & n26476;
  assign n26478 = ~pi648 & ~n26477;
  assign n26479 = ~n26374 & n26478;
  assign n26480 = ~pi619 & n26399;
  assign n26481 = pi619 & ~n26473;
  assign n26482 = ~n26480 & ~n26481;
  assign n26483 = pi1159 & n26482;
  assign n26484 = ~n26376 & ~n26483;
  assign n26485 = pi648 & n26484;
  assign n26486 = ~n26479 & ~n26485;
  assign n26487 = pi789 & n26486;
  assign n26488 = ~pi789 & n26473;
  assign n26489 = n17356 & ~n26488;
  assign n26490 = ~n26487 & n26489;
  assign n26491 = ~n26426 & ~n26490;
  assign n26492 = n19788 & ~n26491;
  assign n26493 = n20275 & n26401;
  assign n26494 = n17449 & ~n26382;
  assign n26495 = ~pi629 & ~n26494;
  assign n26496 = ~n26493 & n26495;
  assign n26497 = n17448 & ~n26382;
  assign n26498 = n20281 & n26401;
  assign n26499 = pi629 & ~n26498;
  assign n26500 = ~n26497 & n26499;
  assign n26501 = ~n26496 & ~n26500;
  assign n26502 = pi792 & n26501;
  assign n26503 = n19637 & ~n26502;
  assign n26504 = ~n26492 & n26503;
  assign n26505 = ~n26414 & ~n26504;
  assign n26506 = pi644 & n26505;
  assign n26507 = ~pi787 & ~n26402;
  assign n26508 = pi787 & ~n26411;
  assign n26509 = ~n26507 & ~n26508;
  assign n26510 = ~pi644 & n26509;
  assign n26511 = pi715 & ~n26510;
  assign n26512 = ~n26506 & n26511;
  assign n26513 = ~n17247 & ~n26385;
  assign n26514 = n17247 & n26351;
  assign n26515 = ~n26513 & ~n26514;
  assign n26516 = pi644 & ~n26515;
  assign n26517 = ~pi644 & n26351;
  assign n26518 = ~pi715 & ~n26517;
  assign n26519 = ~n26516 & n26518;
  assign n26520 = pi1160 & ~n26519;
  assign n26521 = ~n26512 & n26520;
  assign n26522 = ~pi644 & ~n26515;
  assign n26523 = pi715 & ~n26522;
  assign n26524 = pi644 & n26351;
  assign n26525 = n26523 & ~n26524;
  assign n26526 = pi644 & n26509;
  assign n26527 = ~pi644 & n26505;
  assign n26528 = ~pi715 & ~n26527;
  assign n26529 = ~n26526 & n26528;
  assign n26530 = ~pi1160 & ~n26529;
  assign n26531 = ~n26525 & n26530;
  assign n26532 = ~n26521 & ~n26531;
  assign n26533 = pi790 & ~n26532;
  assign n26534 = ~pi790 & n26505;
  assign n26535 = pi832 & ~n26534;
  assign n26536 = ~n26533 & n26535;
  assign n26537 = ~pi182 & ~n16527;
  assign n26538 = n17159 & ~n26537;
  assign n26539 = n16593 & ~n26537;
  assign n26540 = ~pi734 & n10020;
  assign n26541 = n26537 & ~n26540;
  assign n26542 = ~pi182 & n17592;
  assign n26543 = ~pi38 & ~pi182;
  assign n26544 = n19843 & ~n26543;
  assign n26545 = ~n26542 & ~n26544;
  assign n26546 = ~pi182 & ~n16508;
  assign n26547 = n16744 & ~n26546;
  assign n26548 = ~pi734 & ~n26547;
  assign n26549 = ~n26545 & n26548;
  assign n26550 = ~n26541 & ~n26549;
  assign n26551 = ~pi778 & n26550;
  assign n26552 = pi625 & ~n26550;
  assign n26553 = pi1153 & ~n26552;
  assign n26554 = ~pi625 & n26537;
  assign n26555 = n26553 & ~n26554;
  assign n26556 = ~pi625 & ~n26550;
  assign n26557 = ~pi1153 & ~n26556;
  assign n26558 = pi625 & n26537;
  assign n26559 = n26557 & ~n26558;
  assign n26560 = ~n26555 & ~n26559;
  assign n26561 = pi778 & ~n26560;
  assign n26562 = ~n26551 & ~n26561;
  assign n26563 = ~n16593 & ~n26562;
  assign n26564 = ~n26539 & ~n26563;
  assign n26565 = ~n16589 & n26564;
  assign n26566 = n16589 & n26537;
  assign n26567 = ~n26565 & ~n26566;
  assign n26568 = ~n17159 & n26567;
  assign n26569 = ~n26538 & ~n26568;
  assign n26570 = ~n17183 & n26569;
  assign n26571 = n17183 & n26537;
  assign n26572 = ~n26570 & ~n26571;
  assign n26573 = ~pi792 & n26572;
  assign n26574 = pi628 & ~n26572;
  assign n26575 = pi1156 & ~n26574;
  assign n26576 = ~pi628 & n26537;
  assign n26577 = n26575 & ~n26576;
  assign n26578 = ~pi628 & ~n26572;
  assign n26579 = pi628 & n26537;
  assign n26580 = ~pi1156 & ~n26579;
  assign n26581 = ~n26578 & n26580;
  assign n26582 = ~n26577 & ~n26581;
  assign n26583 = pi792 & ~n26582;
  assign n26584 = ~n26573 & ~n26583;
  assign n26585 = pi647 & ~n26584;
  assign n26586 = ~pi647 & ~n26537;
  assign n26587 = ~n26585 & ~n26586;
  assign n26588 = pi1157 & ~n26587;
  assign n26589 = ~pi647 & n26584;
  assign n26590 = ~pi1157 & ~n26589;
  assign n26591 = pi647 & n26537;
  assign n26592 = n26590 & ~n26591;
  assign n26593 = ~n26588 & ~n26592;
  assign n26594 = pi787 & ~n26593;
  assign n26595 = ~pi787 & ~n26584;
  assign n26596 = ~n26594 & ~n26595;
  assign n26597 = ~pi644 & n26596;
  assign n26598 = pi715 & ~n26597;
  assign n26599 = n17247 & ~n26537;
  assign n26600 = pi182 & ~n10020;
  assign n26601 = ~pi182 & n16449;
  assign n26602 = pi182 & ~n16503;
  assign n26603 = ~pi756 & ~n26602;
  assign n26604 = ~n26601 & n26603;
  assign n26605 = ~pi182 & ~n16357;
  assign n26606 = pi756 & n26605;
  assign n26607 = ~n26604 & ~n26606;
  assign n26608 = ~pi38 & ~n26607;
  assign n26609 = ~pi756 & n16511;
  assign n26610 = ~n26546 & ~n26609;
  assign n26611 = pi38 & ~n26610;
  assign n26612 = n10020 & ~n26611;
  assign n26613 = ~n26608 & n26612;
  assign n26614 = ~n26600 & ~n26613;
  assign n26615 = ~n16521 & ~n26614;
  assign n26616 = n16521 & ~n26537;
  assign n26617 = ~n26615 & ~n26616;
  assign n26618 = ~pi785 & ~n26617;
  assign n26619 = ~n16532 & ~n26537;
  assign n26620 = pi609 & n26615;
  assign n26621 = ~n26619 & ~n26620;
  assign n26622 = pi1155 & ~n26621;
  assign n26623 = ~n16537 & ~n26537;
  assign n26624 = ~pi609 & n26615;
  assign n26625 = ~n26623 & ~n26624;
  assign n26626 = ~pi1155 & ~n26625;
  assign n26627 = ~n26622 & ~n26626;
  assign n26628 = pi785 & ~n26627;
  assign n26629 = ~n26618 & ~n26628;
  assign n26630 = ~pi781 & ~n26629;
  assign n26631 = pi618 & n26629;
  assign n26632 = ~pi618 & n26537;
  assign n26633 = pi1154 & ~n26632;
  assign n26634 = ~n26631 & n26633;
  assign n26635 = ~pi618 & n26629;
  assign n26636 = pi618 & n26537;
  assign n26637 = ~pi1154 & ~n26636;
  assign n26638 = ~n26635 & n26637;
  assign n26639 = ~n26634 & ~n26638;
  assign n26640 = pi781 & ~n26639;
  assign n26641 = ~n26630 & ~n26640;
  assign n26642 = ~pi789 & ~n26641;
  assign n26643 = pi619 & n26641;
  assign n26644 = ~pi619 & n26537;
  assign n26645 = pi1159 & ~n26644;
  assign n26646 = ~n26643 & n26645;
  assign n26647 = ~pi619 & n26641;
  assign n26648 = pi619 & n26537;
  assign n26649 = ~pi1159 & ~n26648;
  assign n26650 = ~n26647 & n26649;
  assign n26651 = ~n26646 & ~n26650;
  assign n26652 = pi789 & ~n26651;
  assign n26653 = ~n26642 & ~n26652;
  assign n26654 = ~n17355 & n26653;
  assign n26655 = n17355 & n26537;
  assign n26656 = ~n26654 & ~n26655;
  assign n26657 = ~n16124 & ~n26656;
  assign n26658 = n16124 & n26537;
  assign n26659 = ~n26657 & ~n26658;
  assign n26660 = ~n17247 & n26659;
  assign n26661 = ~n26599 & ~n26660;
  assign n26662 = pi644 & n26661;
  assign n26663 = ~pi644 & n26537;
  assign n26664 = ~pi715 & ~n26663;
  assign n26665 = ~n26662 & n26664;
  assign n26666 = pi1160 & ~n26665;
  assign n26667 = ~n26598 & n26666;
  assign n26668 = pi644 & n26596;
  assign n26669 = ~pi715 & ~n26668;
  assign n26670 = ~pi644 & n26661;
  assign n26671 = pi644 & n26537;
  assign n26672 = ~n26670 & ~n26671;
  assign n26673 = pi715 & n26672;
  assign n26674 = ~pi1160 & ~n26673;
  assign n26675 = ~n26669 & n26674;
  assign n26676 = ~n26667 & ~n26675;
  assign n26677 = pi790 & ~n26676;
  assign n26678 = ~pi629 & n26577;
  assign n26679 = ~n19999 & n26656;
  assign n26680 = pi629 & n26581;
  assign n26681 = ~n26679 & ~n26680;
  assign n26682 = ~n26678 & n26681;
  assign n26683 = pi792 & ~n26682;
  assign n26684 = pi618 & n26564;
  assign n26685 = pi609 & n26562;
  assign n26686 = pi625 & n26614;
  assign n26687 = ~n26540 & ~n26613;
  assign n26688 = ~pi756 & ~n16917;
  assign n26689 = n18933 & ~n26688;
  assign n26690 = ~pi182 & ~n26689;
  assign n26691 = ~n17079 & ~n26352;
  assign n26692 = pi182 & ~n26691;
  assign n26693 = n6097 & n26692;
  assign n26694 = ~n26690 & ~n26693;
  assign n26695 = pi38 & n26694;
  assign n26696 = ~pi182 & n16853;
  assign n26697 = pi182 & n16935;
  assign n26698 = pi756 & ~n26697;
  assign n26699 = ~n26696 & n26698;
  assign n26700 = pi182 & n16998;
  assign n26701 = ~pi182 & ~n17051;
  assign n26702 = ~pi756 & ~n26701;
  assign n26703 = ~n26700 & n26702;
  assign n26704 = ~n26699 & ~n26703;
  assign n26705 = pi39 & n26704;
  assign n26706 = ~pi182 & ~n17061;
  assign n26707 = pi182 & ~n17058;
  assign n26708 = pi756 & ~n26707;
  assign n26709 = ~n26706 & n26708;
  assign n26710 = ~pi182 & n17067;
  assign n26711 = pi182 & n17065;
  assign n26712 = ~pi756 & ~n26711;
  assign n26713 = ~n26710 & n26712;
  assign n26714 = ~n26709 & ~n26713;
  assign n26715 = ~pi39 & ~n26714;
  assign n26716 = ~pi38 & ~n26715;
  assign n26717 = ~n26705 & n26716;
  assign n26718 = ~pi734 & ~n26717;
  assign n26719 = ~n26695 & n26718;
  assign n26720 = ~n26687 & ~n26719;
  assign n26721 = ~n26600 & ~n26720;
  assign n26722 = ~pi625 & n26721;
  assign n26723 = ~pi1153 & ~n26722;
  assign n26724 = ~n26686 & n26723;
  assign n26725 = ~pi608 & ~n26555;
  assign n26726 = ~n26724 & n26725;
  assign n26727 = ~pi625 & n26614;
  assign n26728 = pi625 & n26721;
  assign n26729 = ~n26727 & ~n26728;
  assign n26730 = pi1153 & n26729;
  assign n26731 = ~n26559 & ~n26730;
  assign n26732 = pi608 & n26731;
  assign n26733 = ~n26726 & ~n26732;
  assign n26734 = pi778 & ~n26733;
  assign n26735 = ~pi778 & n26721;
  assign n26736 = ~n26734 & ~n26735;
  assign n26737 = ~pi609 & ~n26736;
  assign n26738 = ~pi1155 & ~n26737;
  assign n26739 = ~n26685 & n26738;
  assign n26740 = ~pi660 & ~n26622;
  assign n26741 = ~n26739 & n26740;
  assign n26742 = ~pi609 & n26562;
  assign n26743 = pi609 & ~n26736;
  assign n26744 = ~n26742 & ~n26743;
  assign n26745 = pi1155 & n26744;
  assign n26746 = ~n26626 & ~n26745;
  assign n26747 = pi660 & n26746;
  assign n26748 = ~n26741 & ~n26747;
  assign n26749 = pi785 & ~n26748;
  assign n26750 = ~pi785 & ~n26736;
  assign n26751 = ~n26749 & ~n26750;
  assign n26752 = ~pi618 & ~n26751;
  assign n26753 = ~pi1154 & ~n26752;
  assign n26754 = ~n26684 & n26753;
  assign n26755 = ~pi627 & ~n26634;
  assign n26756 = ~n26754 & n26755;
  assign n26757 = ~pi618 & n26564;
  assign n26758 = pi618 & ~n26751;
  assign n26759 = ~n26757 & ~n26758;
  assign n26760 = pi1154 & n26759;
  assign n26761 = ~n26638 & ~n26760;
  assign n26762 = pi627 & n26761;
  assign n26763 = ~n26756 & ~n26762;
  assign n26764 = pi781 & ~n26763;
  assign n26765 = ~pi781 & ~n26751;
  assign n26766 = ~n26764 & ~n26765;
  assign n26767 = ~pi789 & n26766;
  assign n26768 = ~pi619 & ~n26766;
  assign n26769 = pi619 & ~n26567;
  assign n26770 = ~pi1159 & ~n26769;
  assign n26771 = ~n26768 & n26770;
  assign n26772 = ~pi648 & ~n26771;
  assign n26773 = ~n26646 & n26772;
  assign n26774 = ~pi619 & ~n26567;
  assign n26775 = pi619 & ~n26766;
  assign n26776 = ~n26774 & ~n26775;
  assign n26777 = pi1159 & n26776;
  assign n26778 = ~n26650 & ~n26777;
  assign n26779 = pi648 & n26778;
  assign n26780 = ~n26773 & ~n26779;
  assign n26781 = pi789 & n26780;
  assign n26782 = ~n26767 & ~n26781;
  assign n26783 = n17356 & n26782;
  assign n26784 = ~pi626 & ~n26653;
  assign n26785 = pi626 & ~n26537;
  assign n26786 = n17181 & ~n26785;
  assign n26787 = ~n26784 & n26786;
  assign n26788 = n17350 & n26569;
  assign n26789 = pi626 & ~n26653;
  assign n26790 = ~pi626 & ~n26537;
  assign n26791 = n17180 & ~n26790;
  assign n26792 = ~n26789 & n26791;
  assign n26793 = ~n26788 & ~n26792;
  assign n26794 = ~n26787 & n26793;
  assign n26795 = pi788 & ~n26794;
  assign n26796 = n19788 & ~n26795;
  assign n26797 = ~n26783 & n26796;
  assign n26798 = ~n26683 & ~n26797;
  assign n26799 = n19637 & ~n26798;
  assign n26800 = ~n19987 & n26659;
  assign n26801 = pi630 & n26592;
  assign n26802 = ~n26800 & ~n26801;
  assign n26803 = n17244 & ~n26587;
  assign n26804 = n26802 & ~n26803;
  assign n26805 = pi787 & ~n26804;
  assign n26806 = ~n26799 & ~n26805;
  assign n26807 = pi644 & n26666;
  assign n26808 = ~pi644 & n26674;
  assign n26809 = pi790 & ~n26808;
  assign n26810 = ~n26807 & n26809;
  assign n26811 = n26806 & ~n26810;
  assign n26812 = ~n26677 & ~n26811;
  assign n26813 = ~po1038 & ~n26812;
  assign n26814 = ~pi182 & po1038;
  assign n26815 = ~pi832 & ~n26814;
  assign n26816 = ~n26813 & n26815;
  assign po339 = ~n26536 & ~n26816;
  assign n26818 = ~pi183 & ~n2934;
  assign n26819 = ~pi755 & n16510;
  assign n26820 = ~n26818 & ~n26819;
  assign n26821 = ~n17273 & ~n26820;
  assign n26822 = ~pi785 & ~n26821;
  assign n26823 = n16537 & n26819;
  assign n26824 = n26821 & ~n26823;
  assign n26825 = pi1155 & ~n26824;
  assign n26826 = ~pi1155 & ~n26818;
  assign n26827 = ~n26823 & n26826;
  assign n26828 = ~n26825 & ~n26827;
  assign n26829 = pi785 & ~n26828;
  assign n26830 = ~n26822 & ~n26829;
  assign n26831 = ~pi781 & ~n26830;
  assign n26832 = ~n17289 & n26830;
  assign n26833 = pi1154 & ~n26832;
  assign n26834 = ~n17292 & n26830;
  assign n26835 = ~pi1154 & ~n26834;
  assign n26836 = ~n26833 & ~n26835;
  assign n26837 = pi781 & ~n26836;
  assign n26838 = ~n26831 & ~n26837;
  assign n26839 = ~pi789 & ~n26838;
  assign n26840 = ~n22423 & n26838;
  assign n26841 = pi1159 & ~n26840;
  assign n26842 = ~n22426 & n26838;
  assign n26843 = ~pi1159 & ~n26842;
  assign n26844 = ~n26841 & ~n26843;
  assign n26845 = pi789 & ~n26844;
  assign n26846 = ~n26839 & ~n26845;
  assign n26847 = ~n17355 & n26846;
  assign n26848 = n17355 & n26818;
  assign n26849 = ~n26847 & ~n26848;
  assign n26850 = ~n16124 & ~n26849;
  assign n26851 = n16124 & n26818;
  assign n26852 = ~n26850 & ~n26851;
  assign n26853 = ~n19987 & n26852;
  assign n26854 = ~pi725 & n16742;
  assign n26855 = ~n26818 & ~n26854;
  assign n26856 = ~pi778 & ~n26855;
  assign n26857 = ~pi625 & n26854;
  assign n26858 = ~n26855 & ~n26857;
  assign n26859 = pi1153 & ~n26858;
  assign n26860 = ~pi1153 & ~n26818;
  assign n26861 = ~n26857 & n26860;
  assign n26862 = ~n26859 & ~n26861;
  assign n26863 = pi778 & n26862;
  assign n26864 = ~n26856 & ~n26863;
  assign n26865 = ~n17338 & ~n26864;
  assign n26866 = ~n17340 & n26865;
  assign n26867 = ~n17342 & n26866;
  assign n26868 = ~n17425 & n26867;
  assign n26869 = ~n17452 & n26868;
  assign n26870 = ~pi647 & n26869;
  assign n26871 = pi647 & n26818;
  assign n26872 = ~pi1157 & ~n26871;
  assign n26873 = ~n26870 & n26872;
  assign n26874 = ~pi647 & n26818;
  assign n26875 = pi647 & n26869;
  assign n26876 = pi1157 & ~n26875;
  assign n26877 = ~n26874 & n26876;
  assign n26878 = ~n26873 & ~n26877;
  assign n26879 = ~n17246 & ~n26878;
  assign n26880 = ~n26853 & ~n26879;
  assign n26881 = pi787 & ~n26880;
  assign n26882 = ~pi626 & ~n26846;
  assign n26883 = pi626 & ~n26818;
  assign n26884 = n17181 & ~n26883;
  assign n26885 = ~n26882 & n26884;
  assign n26886 = n17350 & n26867;
  assign n26887 = pi626 & ~n26846;
  assign n26888 = ~pi626 & ~n26818;
  assign n26889 = n17180 & ~n26888;
  assign n26890 = ~n26887 & n26889;
  assign n26891 = ~n26886 & ~n26890;
  assign n26892 = ~n26885 & n26891;
  assign n26893 = pi788 & ~n26892;
  assign n26894 = pi618 & n26865;
  assign n26895 = pi609 & ~n26864;
  assign n26896 = ~n16393 & ~n26855;
  assign n26897 = pi625 & n26896;
  assign n26898 = n26820 & ~n26896;
  assign n26899 = ~n26897 & ~n26898;
  assign n26900 = n26860 & ~n26899;
  assign n26901 = ~pi608 & ~n26859;
  assign n26902 = ~n26900 & n26901;
  assign n26903 = pi1153 & ~n26897;
  assign n26904 = n26820 & n26903;
  assign n26905 = ~n26861 & ~n26904;
  assign n26906 = pi608 & n26905;
  assign n26907 = ~n26902 & ~n26906;
  assign n26908 = pi778 & ~n26907;
  assign n26909 = ~pi778 & ~n26898;
  assign n26910 = ~n26908 & ~n26909;
  assign n26911 = ~pi609 & ~n26910;
  assign n26912 = ~pi1155 & ~n26911;
  assign n26913 = ~n26895 & n26912;
  assign n26914 = ~pi660 & ~n26825;
  assign n26915 = ~n26913 & n26914;
  assign n26916 = ~pi609 & ~n26864;
  assign n26917 = pi609 & ~n26910;
  assign n26918 = ~n26916 & ~n26917;
  assign n26919 = pi1155 & n26918;
  assign n26920 = ~n26827 & ~n26919;
  assign n26921 = pi660 & n26920;
  assign n26922 = ~n26915 & ~n26921;
  assign n26923 = pi785 & ~n26922;
  assign n26924 = ~pi785 & ~n26910;
  assign n26925 = ~n26923 & ~n26924;
  assign n26926 = ~pi618 & ~n26925;
  assign n26927 = ~pi1154 & ~n26926;
  assign n26928 = ~n26894 & n26927;
  assign n26929 = ~pi627 & ~n26833;
  assign n26930 = ~n26928 & n26929;
  assign n26931 = ~pi618 & n26865;
  assign n26932 = pi618 & ~n26925;
  assign n26933 = ~n26931 & ~n26932;
  assign n26934 = pi1154 & n26933;
  assign n26935 = ~n26835 & ~n26934;
  assign n26936 = pi627 & n26935;
  assign n26937 = ~n26930 & ~n26936;
  assign n26938 = pi781 & ~n26937;
  assign n26939 = ~pi781 & ~n26925;
  assign n26940 = ~n26938 & ~n26939;
  assign n26941 = ~pi619 & ~n26940;
  assign n26942 = pi619 & n26866;
  assign n26943 = ~pi1159 & ~n26942;
  assign n26944 = ~n26941 & n26943;
  assign n26945 = ~pi648 & ~n26944;
  assign n26946 = ~n26841 & n26945;
  assign n26947 = ~pi619 & n26866;
  assign n26948 = pi619 & ~n26940;
  assign n26949 = ~n26947 & ~n26948;
  assign n26950 = pi1159 & n26949;
  assign n26951 = ~n26843 & ~n26950;
  assign n26952 = pi648 & n26951;
  assign n26953 = ~n26946 & ~n26952;
  assign n26954 = pi789 & n26953;
  assign n26955 = ~pi789 & n26940;
  assign n26956 = n17356 & ~n26955;
  assign n26957 = ~n26954 & n26956;
  assign n26958 = ~n26893 & ~n26957;
  assign n26959 = n19788 & ~n26958;
  assign n26960 = n20275 & n26868;
  assign n26961 = n17449 & ~n26849;
  assign n26962 = ~pi629 & ~n26961;
  assign n26963 = ~n26960 & n26962;
  assign n26964 = n17448 & ~n26849;
  assign n26965 = n20281 & n26868;
  assign n26966 = pi629 & ~n26965;
  assign n26967 = ~n26964 & n26966;
  assign n26968 = ~n26963 & ~n26967;
  assign n26969 = pi792 & n26968;
  assign n26970 = n19637 & ~n26969;
  assign n26971 = ~n26959 & n26970;
  assign n26972 = ~n26881 & ~n26971;
  assign n26973 = pi644 & n26972;
  assign n26974 = ~pi787 & ~n26869;
  assign n26975 = pi787 & ~n26878;
  assign n26976 = ~n26974 & ~n26975;
  assign n26977 = ~pi644 & n26976;
  assign n26978 = pi715 & ~n26977;
  assign n26979 = ~n26973 & n26978;
  assign n26980 = ~n17247 & ~n26852;
  assign n26981 = n17247 & n26818;
  assign n26982 = ~n26980 & ~n26981;
  assign n26983 = pi644 & ~n26982;
  assign n26984 = ~pi644 & n26818;
  assign n26985 = ~pi715 & ~n26984;
  assign n26986 = ~n26983 & n26985;
  assign n26987 = pi1160 & ~n26986;
  assign n26988 = ~n26979 & n26987;
  assign n26989 = ~pi644 & ~n26982;
  assign n26990 = pi715 & ~n26989;
  assign n26991 = pi644 & n26818;
  assign n26992 = n26990 & ~n26991;
  assign n26993 = pi644 & n26976;
  assign n26994 = ~pi644 & n26972;
  assign n26995 = ~pi715 & ~n26994;
  assign n26996 = ~n26993 & n26995;
  assign n26997 = ~pi1160 & ~n26996;
  assign n26998 = ~n26992 & n26997;
  assign n26999 = ~n26988 & ~n26998;
  assign n27000 = pi790 & ~n26999;
  assign n27001 = ~pi790 & n26972;
  assign n27002 = pi832 & ~n27001;
  assign n27003 = ~n27000 & n27002;
  assign n27004 = ~pi183 & ~n16527;
  assign n27005 = n17159 & ~n27004;
  assign n27006 = n16593 & ~n27004;
  assign n27007 = ~pi725 & n10020;
  assign n27008 = n27004 & ~n27007;
  assign n27009 = ~pi183 & n17592;
  assign n27010 = ~pi38 & ~pi183;
  assign n27011 = n19843 & ~n27010;
  assign n27012 = ~n27009 & ~n27011;
  assign n27013 = ~pi183 & ~n16508;
  assign n27014 = n16744 & ~n27013;
  assign n27015 = ~pi725 & ~n27014;
  assign n27016 = ~n27012 & n27015;
  assign n27017 = ~n27008 & ~n27016;
  assign n27018 = ~pi778 & n27017;
  assign n27019 = pi625 & ~n27017;
  assign n27020 = pi1153 & ~n27019;
  assign n27021 = ~pi625 & n27004;
  assign n27022 = n27020 & ~n27021;
  assign n27023 = ~pi625 & ~n27017;
  assign n27024 = ~pi1153 & ~n27023;
  assign n27025 = pi625 & n27004;
  assign n27026 = n27024 & ~n27025;
  assign n27027 = ~n27022 & ~n27026;
  assign n27028 = pi778 & ~n27027;
  assign n27029 = ~n27018 & ~n27028;
  assign n27030 = ~n16593 & ~n27029;
  assign n27031 = ~n27006 & ~n27030;
  assign n27032 = ~n16589 & n27031;
  assign n27033 = n16589 & n27004;
  assign n27034 = ~n27032 & ~n27033;
  assign n27035 = ~n17159 & n27034;
  assign n27036 = ~n27005 & ~n27035;
  assign n27037 = ~n17183 & n27036;
  assign n27038 = n17183 & n27004;
  assign n27039 = ~n27037 & ~n27038;
  assign n27040 = ~pi792 & n27039;
  assign n27041 = pi628 & ~n27039;
  assign n27042 = pi1156 & ~n27041;
  assign n27043 = ~pi628 & n27004;
  assign n27044 = n27042 & ~n27043;
  assign n27045 = ~pi628 & ~n27039;
  assign n27046 = pi628 & n27004;
  assign n27047 = ~pi1156 & ~n27046;
  assign n27048 = ~n27045 & n27047;
  assign n27049 = ~n27044 & ~n27048;
  assign n27050 = pi792 & ~n27049;
  assign n27051 = ~n27040 & ~n27050;
  assign n27052 = pi647 & ~n27051;
  assign n27053 = ~pi647 & ~n27004;
  assign n27054 = ~n27052 & ~n27053;
  assign n27055 = pi1157 & ~n27054;
  assign n27056 = ~pi647 & n27051;
  assign n27057 = ~pi1157 & ~n27056;
  assign n27058 = pi647 & n27004;
  assign n27059 = n27057 & ~n27058;
  assign n27060 = ~n27055 & ~n27059;
  assign n27061 = pi787 & ~n27060;
  assign n27062 = ~pi787 & ~n27051;
  assign n27063 = ~n27061 & ~n27062;
  assign n27064 = ~pi644 & n27063;
  assign n27065 = pi715 & ~n27064;
  assign n27066 = n17247 & ~n27004;
  assign n27067 = pi183 & ~n10020;
  assign n27068 = ~pi183 & n16449;
  assign n27069 = pi183 & ~n16503;
  assign n27070 = ~pi755 & ~n27069;
  assign n27071 = ~n27068 & n27070;
  assign n27072 = ~pi183 & ~n16357;
  assign n27073 = pi755 & n27072;
  assign n27074 = ~n27071 & ~n27073;
  assign n27075 = ~pi38 & ~n27074;
  assign n27076 = ~pi755 & n16511;
  assign n27077 = ~n27013 & ~n27076;
  assign n27078 = pi38 & ~n27077;
  assign n27079 = n10020 & ~n27078;
  assign n27080 = ~n27075 & n27079;
  assign n27081 = ~n27067 & ~n27080;
  assign n27082 = ~n16521 & ~n27081;
  assign n27083 = n16521 & ~n27004;
  assign n27084 = ~n27082 & ~n27083;
  assign n27085 = ~pi785 & ~n27084;
  assign n27086 = ~n16532 & ~n27004;
  assign n27087 = pi609 & n27082;
  assign n27088 = ~n27086 & ~n27087;
  assign n27089 = pi1155 & ~n27088;
  assign n27090 = ~n16537 & ~n27004;
  assign n27091 = ~pi609 & n27082;
  assign n27092 = ~n27090 & ~n27091;
  assign n27093 = ~pi1155 & ~n27092;
  assign n27094 = ~n27089 & ~n27093;
  assign n27095 = pi785 & ~n27094;
  assign n27096 = ~n27085 & ~n27095;
  assign n27097 = ~pi781 & ~n27096;
  assign n27098 = pi618 & n27096;
  assign n27099 = ~pi618 & n27004;
  assign n27100 = pi1154 & ~n27099;
  assign n27101 = ~n27098 & n27100;
  assign n27102 = ~pi618 & n27096;
  assign n27103 = pi618 & n27004;
  assign n27104 = ~pi1154 & ~n27103;
  assign n27105 = ~n27102 & n27104;
  assign n27106 = ~n27101 & ~n27105;
  assign n27107 = pi781 & ~n27106;
  assign n27108 = ~n27097 & ~n27107;
  assign n27109 = ~pi789 & ~n27108;
  assign n27110 = pi619 & n27108;
  assign n27111 = ~pi619 & n27004;
  assign n27112 = pi1159 & ~n27111;
  assign n27113 = ~n27110 & n27112;
  assign n27114 = ~pi619 & n27108;
  assign n27115 = pi619 & n27004;
  assign n27116 = ~pi1159 & ~n27115;
  assign n27117 = ~n27114 & n27116;
  assign n27118 = ~n27113 & ~n27117;
  assign n27119 = pi789 & ~n27118;
  assign n27120 = ~n27109 & ~n27119;
  assign n27121 = ~n17355 & n27120;
  assign n27122 = n17355 & n27004;
  assign n27123 = ~n27121 & ~n27122;
  assign n27124 = ~n16124 & ~n27123;
  assign n27125 = n16124 & n27004;
  assign n27126 = ~n27124 & ~n27125;
  assign n27127 = ~n17247 & n27126;
  assign n27128 = ~n27066 & ~n27127;
  assign n27129 = pi644 & n27128;
  assign n27130 = ~pi644 & n27004;
  assign n27131 = ~pi715 & ~n27130;
  assign n27132 = ~n27129 & n27131;
  assign n27133 = pi1160 & ~n27132;
  assign n27134 = ~n27065 & n27133;
  assign n27135 = pi644 & n27063;
  assign n27136 = ~pi715 & ~n27135;
  assign n27137 = ~pi644 & n27128;
  assign n27138 = pi644 & n27004;
  assign n27139 = ~n27137 & ~n27138;
  assign n27140 = pi715 & n27139;
  assign n27141 = ~pi1160 & ~n27140;
  assign n27142 = ~n27136 & n27141;
  assign n27143 = ~n27134 & ~n27142;
  assign n27144 = pi790 & ~n27143;
  assign n27145 = ~pi629 & n27044;
  assign n27146 = ~n19999 & n27123;
  assign n27147 = pi629 & n27048;
  assign n27148 = ~n27146 & ~n27147;
  assign n27149 = ~n27145 & n27148;
  assign n27150 = pi792 & ~n27149;
  assign n27151 = pi618 & n27031;
  assign n27152 = pi609 & n27029;
  assign n27153 = pi625 & n27081;
  assign n27154 = ~n27007 & ~n27080;
  assign n27155 = ~pi755 & ~n16917;
  assign n27156 = n18933 & ~n27155;
  assign n27157 = ~pi183 & ~n27156;
  assign n27158 = ~n17079 & ~n26819;
  assign n27159 = pi183 & ~n27158;
  assign n27160 = n6097 & n27159;
  assign n27161 = ~n27157 & ~n27160;
  assign n27162 = pi38 & n27161;
  assign n27163 = ~pi183 & n16853;
  assign n27164 = pi183 & n16935;
  assign n27165 = pi755 & ~n27164;
  assign n27166 = ~n27163 & n27165;
  assign n27167 = pi183 & n16998;
  assign n27168 = ~pi183 & ~n17051;
  assign n27169 = ~pi755 & ~n27168;
  assign n27170 = ~n27167 & n27169;
  assign n27171 = ~n27166 & ~n27170;
  assign n27172 = pi39 & n27171;
  assign n27173 = ~pi183 & ~n17061;
  assign n27174 = pi183 & ~n17058;
  assign n27175 = pi755 & ~n27174;
  assign n27176 = ~n27173 & n27175;
  assign n27177 = ~pi183 & n17067;
  assign n27178 = pi183 & n17065;
  assign n27179 = ~pi755 & ~n27178;
  assign n27180 = ~n27177 & n27179;
  assign n27181 = ~n27176 & ~n27180;
  assign n27182 = ~pi39 & ~n27181;
  assign n27183 = ~pi38 & ~n27182;
  assign n27184 = ~n27172 & n27183;
  assign n27185 = ~pi725 & ~n27184;
  assign n27186 = ~n27162 & n27185;
  assign n27187 = ~n27154 & ~n27186;
  assign n27188 = ~n27067 & ~n27187;
  assign n27189 = ~pi625 & n27188;
  assign n27190 = ~pi1153 & ~n27189;
  assign n27191 = ~n27153 & n27190;
  assign n27192 = ~pi608 & ~n27022;
  assign n27193 = ~n27191 & n27192;
  assign n27194 = ~pi625 & n27081;
  assign n27195 = pi625 & n27188;
  assign n27196 = ~n27194 & ~n27195;
  assign n27197 = pi1153 & n27196;
  assign n27198 = ~n27026 & ~n27197;
  assign n27199 = pi608 & n27198;
  assign n27200 = ~n27193 & ~n27199;
  assign n27201 = pi778 & ~n27200;
  assign n27202 = ~pi778 & n27188;
  assign n27203 = ~n27201 & ~n27202;
  assign n27204 = ~pi609 & ~n27203;
  assign n27205 = ~pi1155 & ~n27204;
  assign n27206 = ~n27152 & n27205;
  assign n27207 = ~pi660 & ~n27089;
  assign n27208 = ~n27206 & n27207;
  assign n27209 = ~pi609 & n27029;
  assign n27210 = pi609 & ~n27203;
  assign n27211 = ~n27209 & ~n27210;
  assign n27212 = pi1155 & n27211;
  assign n27213 = ~n27093 & ~n27212;
  assign n27214 = pi660 & n27213;
  assign n27215 = ~n27208 & ~n27214;
  assign n27216 = pi785 & ~n27215;
  assign n27217 = ~pi785 & ~n27203;
  assign n27218 = ~n27216 & ~n27217;
  assign n27219 = ~pi618 & ~n27218;
  assign n27220 = ~pi1154 & ~n27219;
  assign n27221 = ~n27151 & n27220;
  assign n27222 = ~pi627 & ~n27101;
  assign n27223 = ~n27221 & n27222;
  assign n27224 = ~pi618 & n27031;
  assign n27225 = pi618 & ~n27218;
  assign n27226 = ~n27224 & ~n27225;
  assign n27227 = pi1154 & n27226;
  assign n27228 = ~n27105 & ~n27227;
  assign n27229 = pi627 & n27228;
  assign n27230 = ~n27223 & ~n27229;
  assign n27231 = pi781 & ~n27230;
  assign n27232 = ~pi781 & ~n27218;
  assign n27233 = ~n27231 & ~n27232;
  assign n27234 = ~pi789 & n27233;
  assign n27235 = ~pi619 & ~n27233;
  assign n27236 = pi619 & ~n27034;
  assign n27237 = ~pi1159 & ~n27236;
  assign n27238 = ~n27235 & n27237;
  assign n27239 = ~pi648 & ~n27238;
  assign n27240 = ~n27113 & n27239;
  assign n27241 = ~pi619 & ~n27034;
  assign n27242 = pi619 & ~n27233;
  assign n27243 = ~n27241 & ~n27242;
  assign n27244 = pi1159 & n27243;
  assign n27245 = ~n27117 & ~n27244;
  assign n27246 = pi648 & n27245;
  assign n27247 = ~n27240 & ~n27246;
  assign n27248 = pi789 & n27247;
  assign n27249 = ~n27234 & ~n27248;
  assign n27250 = n17356 & n27249;
  assign n27251 = ~pi626 & ~n27120;
  assign n27252 = pi626 & ~n27004;
  assign n27253 = n17181 & ~n27252;
  assign n27254 = ~n27251 & n27253;
  assign n27255 = n17350 & n27036;
  assign n27256 = pi626 & ~n27120;
  assign n27257 = ~pi626 & ~n27004;
  assign n27258 = n17180 & ~n27257;
  assign n27259 = ~n27256 & n27258;
  assign n27260 = ~n27255 & ~n27259;
  assign n27261 = ~n27254 & n27260;
  assign n27262 = pi788 & ~n27261;
  assign n27263 = n19788 & ~n27262;
  assign n27264 = ~n27250 & n27263;
  assign n27265 = ~n27150 & ~n27264;
  assign n27266 = n19637 & ~n27265;
  assign n27267 = ~n19987 & n27126;
  assign n27268 = pi630 & n27059;
  assign n27269 = ~n27267 & ~n27268;
  assign n27270 = n17244 & ~n27054;
  assign n27271 = n27269 & ~n27270;
  assign n27272 = pi787 & ~n27271;
  assign n27273 = ~n27266 & ~n27272;
  assign n27274 = pi644 & n27133;
  assign n27275 = ~pi644 & n27141;
  assign n27276 = pi790 & ~n27275;
  assign n27277 = ~n27274 & n27276;
  assign n27278 = n27273 & ~n27277;
  assign n27279 = ~n27144 & ~n27278;
  assign n27280 = ~po1038 & ~n27279;
  assign n27281 = ~pi183 & po1038;
  assign n27282 = ~pi832 & ~n27281;
  assign n27283 = ~n27280 & n27282;
  assign po340 = ~n27003 & ~n27283;
  assign n27285 = ~pi184 & ~n2934;
  assign n27286 = ~pi777 & n16510;
  assign n27287 = ~n27285 & ~n27286;
  assign n27288 = ~n17273 & ~n27287;
  assign n27289 = ~pi785 & ~n27288;
  assign n27290 = n16537 & n27286;
  assign n27291 = n27288 & ~n27290;
  assign n27292 = pi1155 & ~n27291;
  assign n27293 = ~pi1155 & ~n27285;
  assign n27294 = ~n27290 & n27293;
  assign n27295 = ~n27292 & ~n27294;
  assign n27296 = pi785 & ~n27295;
  assign n27297 = ~n27289 & ~n27296;
  assign n27298 = ~pi781 & ~n27297;
  assign n27299 = ~n17289 & n27297;
  assign n27300 = pi1154 & ~n27299;
  assign n27301 = ~n17292 & n27297;
  assign n27302 = ~pi1154 & ~n27301;
  assign n27303 = ~n27300 & ~n27302;
  assign n27304 = pi781 & ~n27303;
  assign n27305 = ~n27298 & ~n27304;
  assign n27306 = ~pi789 & ~n27305;
  assign n27307 = ~n22423 & n27305;
  assign n27308 = pi1159 & ~n27307;
  assign n27309 = ~n22426 & n27305;
  assign n27310 = ~pi1159 & ~n27309;
  assign n27311 = ~n27308 & ~n27310;
  assign n27312 = pi789 & ~n27311;
  assign n27313 = ~n27306 & ~n27312;
  assign n27314 = ~n17355 & n27313;
  assign n27315 = n17355 & n27285;
  assign n27316 = ~n27314 & ~n27315;
  assign n27317 = ~n16124 & ~n27316;
  assign n27318 = n16124 & n27285;
  assign n27319 = ~n27317 & ~n27318;
  assign n27320 = ~n19987 & n27319;
  assign n27321 = ~pi737 & n16742;
  assign n27322 = ~n27285 & ~n27321;
  assign n27323 = ~pi778 & ~n27322;
  assign n27324 = ~pi625 & n27321;
  assign n27325 = ~n27322 & ~n27324;
  assign n27326 = pi1153 & ~n27325;
  assign n27327 = ~pi1153 & ~n27285;
  assign n27328 = ~n27324 & n27327;
  assign n27329 = ~n27326 & ~n27328;
  assign n27330 = pi778 & n27329;
  assign n27331 = ~n27323 & ~n27330;
  assign n27332 = ~n17338 & ~n27331;
  assign n27333 = ~n17340 & n27332;
  assign n27334 = ~n17342 & n27333;
  assign n27335 = ~n17425 & n27334;
  assign n27336 = ~n17452 & n27335;
  assign n27337 = ~pi647 & n27336;
  assign n27338 = pi647 & n27285;
  assign n27339 = ~pi1157 & ~n27338;
  assign n27340 = ~n27337 & n27339;
  assign n27341 = ~pi647 & n27285;
  assign n27342 = pi647 & n27336;
  assign n27343 = pi1157 & ~n27342;
  assign n27344 = ~n27341 & n27343;
  assign n27345 = ~n27340 & ~n27344;
  assign n27346 = ~n17246 & ~n27345;
  assign n27347 = ~n27320 & ~n27346;
  assign n27348 = pi787 & ~n27347;
  assign n27349 = ~pi626 & ~n27313;
  assign n27350 = pi626 & ~n27285;
  assign n27351 = n17181 & ~n27350;
  assign n27352 = ~n27349 & n27351;
  assign n27353 = n17350 & n27334;
  assign n27354 = pi626 & ~n27313;
  assign n27355 = ~pi626 & ~n27285;
  assign n27356 = n17180 & ~n27355;
  assign n27357 = ~n27354 & n27356;
  assign n27358 = ~n27353 & ~n27357;
  assign n27359 = ~n27352 & n27358;
  assign n27360 = pi788 & ~n27359;
  assign n27361 = pi618 & n27332;
  assign n27362 = pi609 & ~n27331;
  assign n27363 = ~n16393 & ~n27322;
  assign n27364 = pi625 & n27363;
  assign n27365 = n27287 & ~n27363;
  assign n27366 = ~n27364 & ~n27365;
  assign n27367 = n27327 & ~n27366;
  assign n27368 = ~pi608 & ~n27326;
  assign n27369 = ~n27367 & n27368;
  assign n27370 = pi1153 & ~n27364;
  assign n27371 = n27287 & n27370;
  assign n27372 = ~n27328 & ~n27371;
  assign n27373 = pi608 & n27372;
  assign n27374 = ~n27369 & ~n27373;
  assign n27375 = pi778 & ~n27374;
  assign n27376 = ~pi778 & ~n27365;
  assign n27377 = ~n27375 & ~n27376;
  assign n27378 = ~pi609 & ~n27377;
  assign n27379 = ~pi1155 & ~n27378;
  assign n27380 = ~n27362 & n27379;
  assign n27381 = ~pi660 & ~n27292;
  assign n27382 = ~n27380 & n27381;
  assign n27383 = ~pi609 & ~n27331;
  assign n27384 = pi609 & ~n27377;
  assign n27385 = ~n27383 & ~n27384;
  assign n27386 = pi1155 & n27385;
  assign n27387 = ~n27294 & ~n27386;
  assign n27388 = pi660 & n27387;
  assign n27389 = ~n27382 & ~n27388;
  assign n27390 = pi785 & ~n27389;
  assign n27391 = ~pi785 & ~n27377;
  assign n27392 = ~n27390 & ~n27391;
  assign n27393 = ~pi618 & ~n27392;
  assign n27394 = ~pi1154 & ~n27393;
  assign n27395 = ~n27361 & n27394;
  assign n27396 = ~pi627 & ~n27300;
  assign n27397 = ~n27395 & n27396;
  assign n27398 = ~pi618 & n27332;
  assign n27399 = pi618 & ~n27392;
  assign n27400 = ~n27398 & ~n27399;
  assign n27401 = pi1154 & n27400;
  assign n27402 = ~n27302 & ~n27401;
  assign n27403 = pi627 & n27402;
  assign n27404 = ~n27397 & ~n27403;
  assign n27405 = pi781 & ~n27404;
  assign n27406 = ~pi781 & ~n27392;
  assign n27407 = ~n27405 & ~n27406;
  assign n27408 = ~pi619 & ~n27407;
  assign n27409 = pi619 & n27333;
  assign n27410 = ~pi1159 & ~n27409;
  assign n27411 = ~n27408 & n27410;
  assign n27412 = ~pi648 & ~n27411;
  assign n27413 = ~n27308 & n27412;
  assign n27414 = ~pi619 & n27333;
  assign n27415 = pi619 & ~n27407;
  assign n27416 = ~n27414 & ~n27415;
  assign n27417 = pi1159 & n27416;
  assign n27418 = ~n27310 & ~n27417;
  assign n27419 = pi648 & n27418;
  assign n27420 = ~n27413 & ~n27419;
  assign n27421 = pi789 & n27420;
  assign n27422 = ~pi789 & n27407;
  assign n27423 = n17356 & ~n27422;
  assign n27424 = ~n27421 & n27423;
  assign n27425 = ~n27360 & ~n27424;
  assign n27426 = n19788 & ~n27425;
  assign n27427 = n20275 & n27335;
  assign n27428 = n17449 & ~n27316;
  assign n27429 = ~pi629 & ~n27428;
  assign n27430 = ~n27427 & n27429;
  assign n27431 = n17448 & ~n27316;
  assign n27432 = n20281 & n27335;
  assign n27433 = pi629 & ~n27432;
  assign n27434 = ~n27431 & n27433;
  assign n27435 = ~n27430 & ~n27434;
  assign n27436 = pi792 & n27435;
  assign n27437 = n19637 & ~n27436;
  assign n27438 = ~n27426 & n27437;
  assign n27439 = ~n27348 & ~n27438;
  assign n27440 = pi644 & n27439;
  assign n27441 = ~pi787 & ~n27336;
  assign n27442 = pi787 & ~n27345;
  assign n27443 = ~n27441 & ~n27442;
  assign n27444 = ~pi644 & n27443;
  assign n27445 = pi715 & ~n27444;
  assign n27446 = ~n27440 & n27445;
  assign n27447 = ~n17247 & ~n27319;
  assign n27448 = n17247 & n27285;
  assign n27449 = ~n27447 & ~n27448;
  assign n27450 = pi644 & ~n27449;
  assign n27451 = ~pi644 & n27285;
  assign n27452 = ~pi715 & ~n27451;
  assign n27453 = ~n27450 & n27452;
  assign n27454 = pi1160 & ~n27453;
  assign n27455 = ~n27446 & n27454;
  assign n27456 = ~pi644 & ~n27449;
  assign n27457 = pi715 & ~n27456;
  assign n27458 = pi644 & n27285;
  assign n27459 = n27457 & ~n27458;
  assign n27460 = pi644 & n27443;
  assign n27461 = ~pi644 & n27439;
  assign n27462 = ~pi715 & ~n27461;
  assign n27463 = ~n27460 & n27462;
  assign n27464 = ~pi1160 & ~n27463;
  assign n27465 = ~n27459 & n27464;
  assign n27466 = ~n27455 & ~n27465;
  assign n27467 = pi790 & ~n27466;
  assign n27468 = ~pi790 & n27439;
  assign n27469 = pi832 & ~n27468;
  assign n27470 = ~n27467 & n27469;
  assign n27471 = ~pi184 & ~n16527;
  assign n27472 = n17159 & ~n27471;
  assign n27473 = n16593 & ~n27471;
  assign n27474 = ~pi737 & n10020;
  assign n27475 = n27471 & ~n27474;
  assign n27476 = ~pi184 & n17592;
  assign n27477 = ~pi38 & ~pi184;
  assign n27478 = n19843 & ~n27477;
  assign n27479 = ~n27476 & ~n27478;
  assign n27480 = ~pi184 & ~n16508;
  assign n27481 = n16744 & ~n27480;
  assign n27482 = ~pi737 & ~n27481;
  assign n27483 = ~n27479 & n27482;
  assign n27484 = ~n27475 & ~n27483;
  assign n27485 = ~pi778 & n27484;
  assign n27486 = pi625 & ~n27484;
  assign n27487 = pi1153 & ~n27486;
  assign n27488 = ~pi625 & n27471;
  assign n27489 = n27487 & ~n27488;
  assign n27490 = ~pi625 & ~n27484;
  assign n27491 = ~pi1153 & ~n27490;
  assign n27492 = pi625 & n27471;
  assign n27493 = n27491 & ~n27492;
  assign n27494 = ~n27489 & ~n27493;
  assign n27495 = pi778 & ~n27494;
  assign n27496 = ~n27485 & ~n27495;
  assign n27497 = ~n16593 & ~n27496;
  assign n27498 = ~n27473 & ~n27497;
  assign n27499 = ~n16589 & n27498;
  assign n27500 = n16589 & n27471;
  assign n27501 = ~n27499 & ~n27500;
  assign n27502 = ~n17159 & n27501;
  assign n27503 = ~n27472 & ~n27502;
  assign n27504 = ~n17183 & n27503;
  assign n27505 = n17183 & n27471;
  assign n27506 = ~n27504 & ~n27505;
  assign n27507 = ~pi792 & n27506;
  assign n27508 = pi628 & ~n27506;
  assign n27509 = pi1156 & ~n27508;
  assign n27510 = ~pi628 & n27471;
  assign n27511 = n27509 & ~n27510;
  assign n27512 = ~pi628 & ~n27506;
  assign n27513 = pi628 & n27471;
  assign n27514 = ~pi1156 & ~n27513;
  assign n27515 = ~n27512 & n27514;
  assign n27516 = ~n27511 & ~n27515;
  assign n27517 = pi792 & ~n27516;
  assign n27518 = ~n27507 & ~n27517;
  assign n27519 = pi647 & ~n27518;
  assign n27520 = ~pi647 & ~n27471;
  assign n27521 = ~n27519 & ~n27520;
  assign n27522 = pi1157 & ~n27521;
  assign n27523 = ~pi647 & n27518;
  assign n27524 = ~pi1157 & ~n27523;
  assign n27525 = pi647 & n27471;
  assign n27526 = n27524 & ~n27525;
  assign n27527 = ~n27522 & ~n27526;
  assign n27528 = pi787 & ~n27527;
  assign n27529 = ~pi787 & ~n27518;
  assign n27530 = ~n27528 & ~n27529;
  assign n27531 = ~pi644 & n27530;
  assign n27532 = pi715 & ~n27531;
  assign n27533 = n17247 & ~n27471;
  assign n27534 = pi184 & ~n10020;
  assign n27535 = ~pi184 & n16449;
  assign n27536 = pi184 & ~n16503;
  assign n27537 = ~pi777 & ~n27536;
  assign n27538 = ~n27535 & n27537;
  assign n27539 = ~pi184 & ~n16357;
  assign n27540 = pi777 & n27539;
  assign n27541 = ~n27538 & ~n27540;
  assign n27542 = ~pi38 & ~n27541;
  assign n27543 = ~pi777 & n16511;
  assign n27544 = ~n27480 & ~n27543;
  assign n27545 = pi38 & ~n27544;
  assign n27546 = n10020 & ~n27545;
  assign n27547 = ~n27542 & n27546;
  assign n27548 = ~n27534 & ~n27547;
  assign n27549 = ~n16521 & ~n27548;
  assign n27550 = n16521 & ~n27471;
  assign n27551 = ~n27549 & ~n27550;
  assign n27552 = ~pi785 & ~n27551;
  assign n27553 = ~n16532 & ~n27471;
  assign n27554 = pi609 & n27549;
  assign n27555 = ~n27553 & ~n27554;
  assign n27556 = pi1155 & ~n27555;
  assign n27557 = ~n16537 & ~n27471;
  assign n27558 = ~pi609 & n27549;
  assign n27559 = ~n27557 & ~n27558;
  assign n27560 = ~pi1155 & ~n27559;
  assign n27561 = ~n27556 & ~n27560;
  assign n27562 = pi785 & ~n27561;
  assign n27563 = ~n27552 & ~n27562;
  assign n27564 = ~pi781 & ~n27563;
  assign n27565 = pi618 & n27563;
  assign n27566 = ~pi618 & n27471;
  assign n27567 = pi1154 & ~n27566;
  assign n27568 = ~n27565 & n27567;
  assign n27569 = ~pi618 & n27563;
  assign n27570 = pi618 & n27471;
  assign n27571 = ~pi1154 & ~n27570;
  assign n27572 = ~n27569 & n27571;
  assign n27573 = ~n27568 & ~n27572;
  assign n27574 = pi781 & ~n27573;
  assign n27575 = ~n27564 & ~n27574;
  assign n27576 = ~pi789 & ~n27575;
  assign n27577 = pi619 & n27575;
  assign n27578 = ~pi619 & n27471;
  assign n27579 = pi1159 & ~n27578;
  assign n27580 = ~n27577 & n27579;
  assign n27581 = ~pi619 & n27575;
  assign n27582 = pi619 & n27471;
  assign n27583 = ~pi1159 & ~n27582;
  assign n27584 = ~n27581 & n27583;
  assign n27585 = ~n27580 & ~n27584;
  assign n27586 = pi789 & ~n27585;
  assign n27587 = ~n27576 & ~n27586;
  assign n27588 = ~n17355 & n27587;
  assign n27589 = n17355 & n27471;
  assign n27590 = ~n27588 & ~n27589;
  assign n27591 = ~n16124 & ~n27590;
  assign n27592 = n16124 & n27471;
  assign n27593 = ~n27591 & ~n27592;
  assign n27594 = ~n17247 & n27593;
  assign n27595 = ~n27533 & ~n27594;
  assign n27596 = pi644 & n27595;
  assign n27597 = ~pi644 & n27471;
  assign n27598 = ~pi715 & ~n27597;
  assign n27599 = ~n27596 & n27598;
  assign n27600 = pi1160 & ~n27599;
  assign n27601 = ~n27532 & n27600;
  assign n27602 = pi644 & n27530;
  assign n27603 = ~pi715 & ~n27602;
  assign n27604 = ~pi644 & n27595;
  assign n27605 = pi644 & n27471;
  assign n27606 = ~n27604 & ~n27605;
  assign n27607 = pi715 & n27606;
  assign n27608 = ~pi1160 & ~n27607;
  assign n27609 = ~n27603 & n27608;
  assign n27610 = ~n27601 & ~n27609;
  assign n27611 = pi790 & ~n27610;
  assign n27612 = ~pi629 & n27511;
  assign n27613 = ~n19999 & n27590;
  assign n27614 = pi629 & n27515;
  assign n27615 = ~n27613 & ~n27614;
  assign n27616 = ~n27612 & n27615;
  assign n27617 = pi792 & ~n27616;
  assign n27618 = pi618 & n27498;
  assign n27619 = pi609 & n27496;
  assign n27620 = pi625 & n27548;
  assign n27621 = ~n27474 & ~n27547;
  assign n27622 = ~pi777 & ~n16917;
  assign n27623 = n18933 & ~n27622;
  assign n27624 = ~pi184 & ~n27623;
  assign n27625 = ~n17079 & ~n27286;
  assign n27626 = pi184 & ~n27625;
  assign n27627 = n6097 & n27626;
  assign n27628 = ~n27624 & ~n27627;
  assign n27629 = pi38 & n27628;
  assign n27630 = ~pi184 & n16853;
  assign n27631 = pi184 & n16935;
  assign n27632 = pi777 & ~n27631;
  assign n27633 = ~n27630 & n27632;
  assign n27634 = pi184 & n16998;
  assign n27635 = ~pi184 & ~n17051;
  assign n27636 = ~pi777 & ~n27635;
  assign n27637 = ~n27634 & n27636;
  assign n27638 = ~n27633 & ~n27637;
  assign n27639 = pi39 & n27638;
  assign n27640 = ~pi184 & ~n17061;
  assign n27641 = pi184 & ~n17058;
  assign n27642 = pi777 & ~n27641;
  assign n27643 = ~n27640 & n27642;
  assign n27644 = ~pi184 & n17067;
  assign n27645 = pi184 & n17065;
  assign n27646 = ~pi777 & ~n27645;
  assign n27647 = ~n27644 & n27646;
  assign n27648 = ~n27643 & ~n27647;
  assign n27649 = ~pi39 & ~n27648;
  assign n27650 = ~pi38 & ~n27649;
  assign n27651 = ~n27639 & n27650;
  assign n27652 = ~pi737 & ~n27651;
  assign n27653 = ~n27629 & n27652;
  assign n27654 = ~n27621 & ~n27653;
  assign n27655 = ~n27534 & ~n27654;
  assign n27656 = ~pi625 & n27655;
  assign n27657 = ~pi1153 & ~n27656;
  assign n27658 = ~n27620 & n27657;
  assign n27659 = ~pi608 & ~n27489;
  assign n27660 = ~n27658 & n27659;
  assign n27661 = ~pi625 & n27548;
  assign n27662 = pi625 & n27655;
  assign n27663 = ~n27661 & ~n27662;
  assign n27664 = pi1153 & n27663;
  assign n27665 = ~n27493 & ~n27664;
  assign n27666 = pi608 & n27665;
  assign n27667 = ~n27660 & ~n27666;
  assign n27668 = pi778 & ~n27667;
  assign n27669 = ~pi778 & n27655;
  assign n27670 = ~n27668 & ~n27669;
  assign n27671 = ~pi609 & ~n27670;
  assign n27672 = ~pi1155 & ~n27671;
  assign n27673 = ~n27619 & n27672;
  assign n27674 = ~pi660 & ~n27556;
  assign n27675 = ~n27673 & n27674;
  assign n27676 = ~pi609 & n27496;
  assign n27677 = pi609 & ~n27670;
  assign n27678 = ~n27676 & ~n27677;
  assign n27679 = pi1155 & n27678;
  assign n27680 = ~n27560 & ~n27679;
  assign n27681 = pi660 & n27680;
  assign n27682 = ~n27675 & ~n27681;
  assign n27683 = pi785 & ~n27682;
  assign n27684 = ~pi785 & ~n27670;
  assign n27685 = ~n27683 & ~n27684;
  assign n27686 = ~pi618 & ~n27685;
  assign n27687 = ~pi1154 & ~n27686;
  assign n27688 = ~n27618 & n27687;
  assign n27689 = ~pi627 & ~n27568;
  assign n27690 = ~n27688 & n27689;
  assign n27691 = ~pi618 & n27498;
  assign n27692 = pi618 & ~n27685;
  assign n27693 = ~n27691 & ~n27692;
  assign n27694 = pi1154 & n27693;
  assign n27695 = ~n27572 & ~n27694;
  assign n27696 = pi627 & n27695;
  assign n27697 = ~n27690 & ~n27696;
  assign n27698 = pi781 & ~n27697;
  assign n27699 = ~pi781 & ~n27685;
  assign n27700 = ~n27698 & ~n27699;
  assign n27701 = ~pi789 & n27700;
  assign n27702 = ~pi619 & ~n27700;
  assign n27703 = pi619 & ~n27501;
  assign n27704 = ~pi1159 & ~n27703;
  assign n27705 = ~n27702 & n27704;
  assign n27706 = ~pi648 & ~n27705;
  assign n27707 = ~n27580 & n27706;
  assign n27708 = ~pi619 & ~n27501;
  assign n27709 = pi619 & ~n27700;
  assign n27710 = ~n27708 & ~n27709;
  assign n27711 = pi1159 & n27710;
  assign n27712 = ~n27584 & ~n27711;
  assign n27713 = pi648 & n27712;
  assign n27714 = ~n27707 & ~n27713;
  assign n27715 = pi789 & n27714;
  assign n27716 = ~n27701 & ~n27715;
  assign n27717 = n17356 & n27716;
  assign n27718 = ~pi626 & ~n27587;
  assign n27719 = pi626 & ~n27471;
  assign n27720 = n17181 & ~n27719;
  assign n27721 = ~n27718 & n27720;
  assign n27722 = n17350 & n27503;
  assign n27723 = pi626 & ~n27587;
  assign n27724 = ~pi626 & ~n27471;
  assign n27725 = n17180 & ~n27724;
  assign n27726 = ~n27723 & n27725;
  assign n27727 = ~n27722 & ~n27726;
  assign n27728 = ~n27721 & n27727;
  assign n27729 = pi788 & ~n27728;
  assign n27730 = n19788 & ~n27729;
  assign n27731 = ~n27717 & n27730;
  assign n27732 = ~n27617 & ~n27731;
  assign n27733 = n19637 & ~n27732;
  assign n27734 = ~n19987 & n27593;
  assign n27735 = pi630 & n27526;
  assign n27736 = ~n27734 & ~n27735;
  assign n27737 = n17244 & ~n27521;
  assign n27738 = n27736 & ~n27737;
  assign n27739 = pi787 & ~n27738;
  assign n27740 = ~n27733 & ~n27739;
  assign n27741 = pi644 & n27600;
  assign n27742 = ~pi644 & n27608;
  assign n27743 = pi790 & ~n27742;
  assign n27744 = ~n27741 & n27743;
  assign n27745 = n27740 & ~n27744;
  assign n27746 = ~n27611 & ~n27745;
  assign n27747 = ~po1038 & ~n27746;
  assign n27748 = ~pi184 & po1038;
  assign n27749 = ~pi832 & ~n27748;
  assign n27750 = ~n27747 & n27749;
  assign po341 = ~n27470 & ~n27750;
  assign n27752 = ~pi185 & ~n2934;
  assign n27753 = ~pi751 & n16510;
  assign n27754 = ~n27752 & ~n27753;
  assign n27755 = ~n17273 & ~n27754;
  assign n27756 = ~pi785 & ~n27755;
  assign n27757 = n16537 & n27753;
  assign n27758 = n27755 & ~n27757;
  assign n27759 = pi1155 & ~n27758;
  assign n27760 = ~pi1155 & ~n27752;
  assign n27761 = ~n27757 & n27760;
  assign n27762 = ~n27759 & ~n27761;
  assign n27763 = pi785 & ~n27762;
  assign n27764 = ~n27756 & ~n27763;
  assign n27765 = ~pi781 & ~n27764;
  assign n27766 = ~n17289 & n27764;
  assign n27767 = pi1154 & ~n27766;
  assign n27768 = ~n17292 & n27764;
  assign n27769 = ~pi1154 & ~n27768;
  assign n27770 = ~n27767 & ~n27769;
  assign n27771 = pi781 & ~n27770;
  assign n27772 = ~n27765 & ~n27771;
  assign n27773 = ~pi789 & ~n27772;
  assign n27774 = ~n22423 & n27772;
  assign n27775 = pi1159 & ~n27774;
  assign n27776 = ~n22426 & n27772;
  assign n27777 = ~pi1159 & ~n27776;
  assign n27778 = ~n27775 & ~n27777;
  assign n27779 = pi789 & ~n27778;
  assign n27780 = ~n27773 & ~n27779;
  assign n27781 = ~n17355 & n27780;
  assign n27782 = n17355 & n27752;
  assign n27783 = ~n27781 & ~n27782;
  assign n27784 = ~n16124 & ~n27783;
  assign n27785 = n16124 & n27752;
  assign n27786 = ~n27784 & ~n27785;
  assign n27787 = ~n19987 & n27786;
  assign n27788 = ~pi701 & n16742;
  assign n27789 = ~n27752 & ~n27788;
  assign n27790 = ~pi778 & ~n27789;
  assign n27791 = ~pi625 & n27788;
  assign n27792 = ~n27789 & ~n27791;
  assign n27793 = pi1153 & ~n27792;
  assign n27794 = ~pi1153 & ~n27752;
  assign n27795 = ~n27791 & n27794;
  assign n27796 = ~n27793 & ~n27795;
  assign n27797 = pi778 & n27796;
  assign n27798 = ~n27790 & ~n27797;
  assign n27799 = ~n17338 & ~n27798;
  assign n27800 = ~n17340 & n27799;
  assign n27801 = ~n17342 & n27800;
  assign n27802 = ~n17425 & n27801;
  assign n27803 = ~n17452 & n27802;
  assign n27804 = ~pi647 & n27803;
  assign n27805 = pi647 & n27752;
  assign n27806 = ~pi1157 & ~n27805;
  assign n27807 = ~n27804 & n27806;
  assign n27808 = ~pi647 & n27752;
  assign n27809 = pi647 & n27803;
  assign n27810 = pi1157 & ~n27809;
  assign n27811 = ~n27808 & n27810;
  assign n27812 = ~n27807 & ~n27811;
  assign n27813 = ~n17246 & ~n27812;
  assign n27814 = ~n27787 & ~n27813;
  assign n27815 = pi787 & ~n27814;
  assign n27816 = ~pi626 & ~n27780;
  assign n27817 = pi626 & ~n27752;
  assign n27818 = n17181 & ~n27817;
  assign n27819 = ~n27816 & n27818;
  assign n27820 = n17350 & n27801;
  assign n27821 = pi626 & ~n27780;
  assign n27822 = ~pi626 & ~n27752;
  assign n27823 = n17180 & ~n27822;
  assign n27824 = ~n27821 & n27823;
  assign n27825 = ~n27820 & ~n27824;
  assign n27826 = ~n27819 & n27825;
  assign n27827 = pi788 & ~n27826;
  assign n27828 = pi618 & n27799;
  assign n27829 = pi609 & ~n27798;
  assign n27830 = ~n16393 & ~n27789;
  assign n27831 = pi625 & n27830;
  assign n27832 = n27754 & ~n27830;
  assign n27833 = ~n27831 & ~n27832;
  assign n27834 = n27794 & ~n27833;
  assign n27835 = ~pi608 & ~n27793;
  assign n27836 = ~n27834 & n27835;
  assign n27837 = pi1153 & ~n27831;
  assign n27838 = n27754 & n27837;
  assign n27839 = ~n27795 & ~n27838;
  assign n27840 = pi608 & n27839;
  assign n27841 = ~n27836 & ~n27840;
  assign n27842 = pi778 & ~n27841;
  assign n27843 = ~pi778 & ~n27832;
  assign n27844 = ~n27842 & ~n27843;
  assign n27845 = ~pi609 & ~n27844;
  assign n27846 = ~pi1155 & ~n27845;
  assign n27847 = ~n27829 & n27846;
  assign n27848 = ~pi660 & ~n27759;
  assign n27849 = ~n27847 & n27848;
  assign n27850 = ~pi609 & ~n27798;
  assign n27851 = pi609 & ~n27844;
  assign n27852 = ~n27850 & ~n27851;
  assign n27853 = pi1155 & n27852;
  assign n27854 = ~n27761 & ~n27853;
  assign n27855 = pi660 & n27854;
  assign n27856 = ~n27849 & ~n27855;
  assign n27857 = pi785 & ~n27856;
  assign n27858 = ~pi785 & ~n27844;
  assign n27859 = ~n27857 & ~n27858;
  assign n27860 = ~pi618 & ~n27859;
  assign n27861 = ~pi1154 & ~n27860;
  assign n27862 = ~n27828 & n27861;
  assign n27863 = ~pi627 & ~n27767;
  assign n27864 = ~n27862 & n27863;
  assign n27865 = ~pi618 & n27799;
  assign n27866 = pi618 & ~n27859;
  assign n27867 = ~n27865 & ~n27866;
  assign n27868 = pi1154 & n27867;
  assign n27869 = ~n27769 & ~n27868;
  assign n27870 = pi627 & n27869;
  assign n27871 = ~n27864 & ~n27870;
  assign n27872 = pi781 & ~n27871;
  assign n27873 = ~pi781 & ~n27859;
  assign n27874 = ~n27872 & ~n27873;
  assign n27875 = ~pi619 & ~n27874;
  assign n27876 = pi619 & n27800;
  assign n27877 = ~pi1159 & ~n27876;
  assign n27878 = ~n27875 & n27877;
  assign n27879 = ~pi648 & ~n27878;
  assign n27880 = ~n27775 & n27879;
  assign n27881 = ~pi619 & n27800;
  assign n27882 = pi619 & ~n27874;
  assign n27883 = ~n27881 & ~n27882;
  assign n27884 = pi1159 & n27883;
  assign n27885 = ~n27777 & ~n27884;
  assign n27886 = pi648 & n27885;
  assign n27887 = ~n27880 & ~n27886;
  assign n27888 = pi789 & n27887;
  assign n27889 = ~pi789 & n27874;
  assign n27890 = n17356 & ~n27889;
  assign n27891 = ~n27888 & n27890;
  assign n27892 = ~n27827 & ~n27891;
  assign n27893 = n19788 & ~n27892;
  assign n27894 = n20275 & n27802;
  assign n27895 = n17449 & ~n27783;
  assign n27896 = ~pi629 & ~n27895;
  assign n27897 = ~n27894 & n27896;
  assign n27898 = n17448 & ~n27783;
  assign n27899 = n20281 & n27802;
  assign n27900 = pi629 & ~n27899;
  assign n27901 = ~n27898 & n27900;
  assign n27902 = ~n27897 & ~n27901;
  assign n27903 = pi792 & n27902;
  assign n27904 = n19637 & ~n27903;
  assign n27905 = ~n27893 & n27904;
  assign n27906 = ~n27815 & ~n27905;
  assign n27907 = pi644 & n27906;
  assign n27908 = ~pi787 & ~n27803;
  assign n27909 = pi787 & ~n27812;
  assign n27910 = ~n27908 & ~n27909;
  assign n27911 = ~pi644 & n27910;
  assign n27912 = pi715 & ~n27911;
  assign n27913 = ~n27907 & n27912;
  assign n27914 = ~n17247 & ~n27786;
  assign n27915 = n17247 & n27752;
  assign n27916 = ~n27914 & ~n27915;
  assign n27917 = pi644 & ~n27916;
  assign n27918 = ~pi644 & n27752;
  assign n27919 = ~pi715 & ~n27918;
  assign n27920 = ~n27917 & n27919;
  assign n27921 = pi1160 & ~n27920;
  assign n27922 = ~n27913 & n27921;
  assign n27923 = ~pi644 & ~n27916;
  assign n27924 = pi715 & ~n27923;
  assign n27925 = pi644 & n27752;
  assign n27926 = n27924 & ~n27925;
  assign n27927 = pi644 & n27910;
  assign n27928 = ~pi644 & n27906;
  assign n27929 = ~pi715 & ~n27928;
  assign n27930 = ~n27927 & n27929;
  assign n27931 = ~pi1160 & ~n27930;
  assign n27932 = ~n27926 & n27931;
  assign n27933 = ~n27922 & ~n27932;
  assign n27934 = pi790 & ~n27933;
  assign n27935 = ~pi790 & n27906;
  assign n27936 = pi832 & ~n27935;
  assign n27937 = ~n27934 & n27936;
  assign n27938 = ~pi185 & ~n16527;
  assign n27939 = n17159 & ~n27938;
  assign n27940 = n16593 & ~n27938;
  assign n27941 = ~pi701 & n10020;
  assign n27942 = n27938 & ~n27941;
  assign n27943 = ~pi185 & n17592;
  assign n27944 = ~pi38 & ~pi185;
  assign n27945 = n19843 & ~n27944;
  assign n27946 = ~n27943 & ~n27945;
  assign n27947 = ~pi185 & ~n16508;
  assign n27948 = n16744 & ~n27947;
  assign n27949 = ~pi701 & ~n27948;
  assign n27950 = ~n27946 & n27949;
  assign n27951 = ~n27942 & ~n27950;
  assign n27952 = ~pi778 & n27951;
  assign n27953 = pi625 & ~n27951;
  assign n27954 = pi1153 & ~n27953;
  assign n27955 = ~pi625 & n27938;
  assign n27956 = n27954 & ~n27955;
  assign n27957 = ~pi625 & ~n27951;
  assign n27958 = ~pi1153 & ~n27957;
  assign n27959 = pi625 & n27938;
  assign n27960 = n27958 & ~n27959;
  assign n27961 = ~n27956 & ~n27960;
  assign n27962 = pi778 & ~n27961;
  assign n27963 = ~n27952 & ~n27962;
  assign n27964 = ~n16593 & ~n27963;
  assign n27965 = ~n27940 & ~n27964;
  assign n27966 = ~n16589 & n27965;
  assign n27967 = n16589 & n27938;
  assign n27968 = ~n27966 & ~n27967;
  assign n27969 = ~n17159 & n27968;
  assign n27970 = ~n27939 & ~n27969;
  assign n27971 = ~n17183 & n27970;
  assign n27972 = n17183 & n27938;
  assign n27973 = ~n27971 & ~n27972;
  assign n27974 = ~pi792 & n27973;
  assign n27975 = pi628 & ~n27973;
  assign n27976 = pi1156 & ~n27975;
  assign n27977 = ~pi628 & n27938;
  assign n27978 = n27976 & ~n27977;
  assign n27979 = ~pi628 & ~n27973;
  assign n27980 = pi628 & n27938;
  assign n27981 = ~pi1156 & ~n27980;
  assign n27982 = ~n27979 & n27981;
  assign n27983 = ~n27978 & ~n27982;
  assign n27984 = pi792 & ~n27983;
  assign n27985 = ~n27974 & ~n27984;
  assign n27986 = pi647 & ~n27985;
  assign n27987 = ~pi647 & ~n27938;
  assign n27988 = ~n27986 & ~n27987;
  assign n27989 = pi1157 & ~n27988;
  assign n27990 = ~pi647 & n27985;
  assign n27991 = ~pi1157 & ~n27990;
  assign n27992 = pi647 & n27938;
  assign n27993 = n27991 & ~n27992;
  assign n27994 = ~n27989 & ~n27993;
  assign n27995 = pi787 & ~n27994;
  assign n27996 = ~pi787 & ~n27985;
  assign n27997 = ~n27995 & ~n27996;
  assign n27998 = ~pi644 & n27997;
  assign n27999 = pi715 & ~n27998;
  assign n28000 = n17247 & ~n27938;
  assign n28001 = pi185 & ~n10020;
  assign n28002 = ~pi751 & n16511;
  assign n28003 = ~n27947 & ~n28002;
  assign n28004 = pi38 & ~n28003;
  assign n28005 = n10020 & ~n28004;
  assign n28006 = pi751 & n16355;
  assign n28007 = pi185 & n16501;
  assign n28008 = ~n28006 & ~n28007;
  assign n28009 = pi39 & ~n28008;
  assign n28010 = pi185 & pi751;
  assign n28011 = pi185 & ~n16460;
  assign n28012 = ~n20665 & ~n28011;
  assign n28013 = ~pi39 & ~n28012;
  assign n28014 = ~n28010 & ~n28013;
  assign n28015 = ~pi185 & ~pi751;
  assign n28016 = n16449 & n28015;
  assign n28017 = n28014 & ~n28016;
  assign n28018 = ~n28009 & n28017;
  assign n28019 = ~pi38 & n28018;
  assign n28020 = n28005 & ~n28019;
  assign n28021 = ~n28001 & ~n28020;
  assign n28022 = ~n16521 & ~n28021;
  assign n28023 = n16521 & ~n27938;
  assign n28024 = ~n28022 & ~n28023;
  assign n28025 = ~pi785 & ~n28024;
  assign n28026 = ~n16532 & ~n27938;
  assign n28027 = pi609 & n28022;
  assign n28028 = ~n28026 & ~n28027;
  assign n28029 = pi1155 & ~n28028;
  assign n28030 = ~n16537 & ~n27938;
  assign n28031 = ~pi609 & n28022;
  assign n28032 = ~n28030 & ~n28031;
  assign n28033 = ~pi1155 & ~n28032;
  assign n28034 = ~n28029 & ~n28033;
  assign n28035 = pi785 & ~n28034;
  assign n28036 = ~n28025 & ~n28035;
  assign n28037 = ~pi781 & ~n28036;
  assign n28038 = pi618 & n28036;
  assign n28039 = ~pi618 & n27938;
  assign n28040 = pi1154 & ~n28039;
  assign n28041 = ~n28038 & n28040;
  assign n28042 = ~pi618 & n28036;
  assign n28043 = pi618 & n27938;
  assign n28044 = ~pi1154 & ~n28043;
  assign n28045 = ~n28042 & n28044;
  assign n28046 = ~n28041 & ~n28045;
  assign n28047 = pi781 & ~n28046;
  assign n28048 = ~n28037 & ~n28047;
  assign n28049 = ~pi789 & ~n28048;
  assign n28050 = pi619 & n28048;
  assign n28051 = ~pi619 & n27938;
  assign n28052 = pi1159 & ~n28051;
  assign n28053 = ~n28050 & n28052;
  assign n28054 = ~pi619 & n28048;
  assign n28055 = pi619 & n27938;
  assign n28056 = ~pi1159 & ~n28055;
  assign n28057 = ~n28054 & n28056;
  assign n28058 = ~n28053 & ~n28057;
  assign n28059 = pi789 & ~n28058;
  assign n28060 = ~n28049 & ~n28059;
  assign n28061 = ~n17355 & n28060;
  assign n28062 = n17355 & n27938;
  assign n28063 = ~n28061 & ~n28062;
  assign n28064 = ~n16124 & ~n28063;
  assign n28065 = n16124 & n27938;
  assign n28066 = ~n28064 & ~n28065;
  assign n28067 = ~n17247 & n28066;
  assign n28068 = ~n28000 & ~n28067;
  assign n28069 = pi644 & n28068;
  assign n28070 = ~pi644 & n27938;
  assign n28071 = ~pi715 & ~n28070;
  assign n28072 = ~n28069 & n28071;
  assign n28073 = pi1160 & ~n28072;
  assign n28074 = ~n27999 & n28073;
  assign n28075 = pi644 & n27997;
  assign n28076 = ~pi715 & ~n28075;
  assign n28077 = ~pi644 & n28068;
  assign n28078 = pi644 & n27938;
  assign n28079 = ~n28077 & ~n28078;
  assign n28080 = pi715 & n28079;
  assign n28081 = ~pi1160 & ~n28080;
  assign n28082 = ~n28076 & n28081;
  assign n28083 = ~n28074 & ~n28082;
  assign n28084 = pi790 & ~n28083;
  assign n28085 = ~pi629 & n27978;
  assign n28086 = ~n19999 & n28063;
  assign n28087 = pi629 & n27982;
  assign n28088 = ~n28086 & ~n28087;
  assign n28089 = ~n28085 & n28088;
  assign n28090 = pi792 & ~n28089;
  assign n28091 = pi618 & n27965;
  assign n28092 = pi609 & n27963;
  assign n28093 = pi625 & n28021;
  assign n28094 = ~n27941 & ~n28020;
  assign n28095 = ~pi751 & ~n16917;
  assign n28096 = n18933 & ~n28095;
  assign n28097 = ~pi185 & ~n28096;
  assign n28098 = ~n17079 & ~n27753;
  assign n28099 = pi185 & ~n28098;
  assign n28100 = n6097 & n28099;
  assign n28101 = ~n28097 & ~n28100;
  assign n28102 = pi38 & n28101;
  assign n28103 = ~pi185 & n16853;
  assign n28104 = pi185 & n16935;
  assign n28105 = pi751 & ~n28104;
  assign n28106 = ~n28103 & n28105;
  assign n28107 = pi185 & n16998;
  assign n28108 = ~pi185 & ~n17051;
  assign n28109 = ~pi751 & ~n28108;
  assign n28110 = ~n28107 & n28109;
  assign n28111 = ~n28106 & ~n28110;
  assign n28112 = pi39 & n28111;
  assign n28113 = ~pi185 & ~n17061;
  assign n28114 = pi185 & ~n17058;
  assign n28115 = pi751 & ~n28114;
  assign n28116 = ~n28113 & n28115;
  assign n28117 = ~pi185 & n17067;
  assign n28118 = ~pi751 & ~n28117;
  assign n28119 = pi185 & n17065;
  assign n28120 = n28118 & ~n28119;
  assign n28121 = ~n28116 & ~n28120;
  assign n28122 = ~pi39 & ~n28121;
  assign n28123 = ~pi38 & ~n28122;
  assign n28124 = ~n28112 & n28123;
  assign n28125 = ~pi701 & ~n28124;
  assign n28126 = ~n28102 & n28125;
  assign n28127 = ~n28094 & ~n28126;
  assign n28128 = ~n28001 & ~n28127;
  assign n28129 = ~pi625 & n28128;
  assign n28130 = ~pi1153 & ~n28129;
  assign n28131 = ~n28093 & n28130;
  assign n28132 = ~pi608 & ~n27956;
  assign n28133 = ~n28131 & n28132;
  assign n28134 = ~pi625 & n28021;
  assign n28135 = pi625 & n28128;
  assign n28136 = ~n28134 & ~n28135;
  assign n28137 = pi1153 & n28136;
  assign n28138 = ~n27960 & ~n28137;
  assign n28139 = pi608 & n28138;
  assign n28140 = ~n28133 & ~n28139;
  assign n28141 = pi778 & ~n28140;
  assign n28142 = ~pi778 & n28128;
  assign n28143 = ~n28141 & ~n28142;
  assign n28144 = ~pi609 & ~n28143;
  assign n28145 = ~pi1155 & ~n28144;
  assign n28146 = ~n28092 & n28145;
  assign n28147 = ~pi660 & ~n28029;
  assign n28148 = ~n28146 & n28147;
  assign n28149 = ~pi609 & n27963;
  assign n28150 = pi609 & ~n28143;
  assign n28151 = ~n28149 & ~n28150;
  assign n28152 = pi1155 & n28151;
  assign n28153 = ~n28033 & ~n28152;
  assign n28154 = pi660 & n28153;
  assign n28155 = ~n28148 & ~n28154;
  assign n28156 = pi785 & ~n28155;
  assign n28157 = ~pi785 & ~n28143;
  assign n28158 = ~n28156 & ~n28157;
  assign n28159 = ~pi618 & ~n28158;
  assign n28160 = ~pi1154 & ~n28159;
  assign n28161 = ~n28091 & n28160;
  assign n28162 = ~pi627 & ~n28041;
  assign n28163 = ~n28161 & n28162;
  assign n28164 = ~pi618 & n27965;
  assign n28165 = pi618 & ~n28158;
  assign n28166 = ~n28164 & ~n28165;
  assign n28167 = pi1154 & n28166;
  assign n28168 = ~n28045 & ~n28167;
  assign n28169 = pi627 & n28168;
  assign n28170 = ~n28163 & ~n28169;
  assign n28171 = pi781 & ~n28170;
  assign n28172 = ~pi781 & ~n28158;
  assign n28173 = ~n28171 & ~n28172;
  assign n28174 = ~pi789 & n28173;
  assign n28175 = ~pi619 & ~n28173;
  assign n28176 = pi619 & ~n27968;
  assign n28177 = ~pi1159 & ~n28176;
  assign n28178 = ~n28175 & n28177;
  assign n28179 = ~pi648 & ~n28178;
  assign n28180 = ~n28053 & n28179;
  assign n28181 = ~pi619 & ~n27968;
  assign n28182 = pi619 & ~n28173;
  assign n28183 = ~n28181 & ~n28182;
  assign n28184 = pi1159 & n28183;
  assign n28185 = ~n28057 & ~n28184;
  assign n28186 = pi648 & n28185;
  assign n28187 = ~n28180 & ~n28186;
  assign n28188 = pi789 & n28187;
  assign n28189 = ~n28174 & ~n28188;
  assign n28190 = n17356 & n28189;
  assign n28191 = ~pi626 & ~n28060;
  assign n28192 = pi626 & ~n27938;
  assign n28193 = n17181 & ~n28192;
  assign n28194 = ~n28191 & n28193;
  assign n28195 = n17350 & n27970;
  assign n28196 = pi626 & ~n28060;
  assign n28197 = ~pi626 & ~n27938;
  assign n28198 = n17180 & ~n28197;
  assign n28199 = ~n28196 & n28198;
  assign n28200 = ~n28195 & ~n28199;
  assign n28201 = ~n28194 & n28200;
  assign n28202 = pi788 & ~n28201;
  assign n28203 = n19788 & ~n28202;
  assign n28204 = ~n28190 & n28203;
  assign n28205 = ~n28090 & ~n28204;
  assign n28206 = n19637 & ~n28205;
  assign n28207 = ~n19987 & n28066;
  assign n28208 = pi630 & n27993;
  assign n28209 = ~n28207 & ~n28208;
  assign n28210 = n17244 & ~n27988;
  assign n28211 = n28209 & ~n28210;
  assign n28212 = pi787 & ~n28211;
  assign n28213 = ~n28206 & ~n28212;
  assign n28214 = pi644 & n28073;
  assign n28215 = ~pi644 & n28081;
  assign n28216 = pi790 & ~n28215;
  assign n28217 = ~n28214 & n28216;
  assign n28218 = n28213 & ~n28217;
  assign n28219 = ~n28084 & ~n28218;
  assign n28220 = ~po1038 & ~n28219;
  assign n28221 = ~pi185 & po1038;
  assign n28222 = ~pi832 & ~n28221;
  assign n28223 = ~n28220 & n28222;
  assign po342 = ~n27937 & ~n28223;
  assign n28225 = pi186 & ~n10020;
  assign n28226 = ~pi186 & ~n16526;
  assign n28227 = pi752 & ~n28226;
  assign n28228 = pi186 & ~n18803;
  assign n28229 = ~pi186 & ~pi752;
  assign n28230 = n18808 & n28229;
  assign n28231 = ~n28228 & ~n28230;
  assign n28232 = ~n18802 & ~n28231;
  assign n28233 = ~n28227 & ~n28232;
  assign n28234 = n10020 & ~n28233;
  assign n28235 = ~n28225 & ~n28234;
  assign n28236 = ~n16521 & ~n28235;
  assign n28237 = ~pi186 & ~n16527;
  assign n28238 = n16521 & ~n28237;
  assign n28239 = ~n28236 & ~n28238;
  assign n28240 = ~pi785 & ~n28239;
  assign n28241 = ~n16532 & ~n28237;
  assign n28242 = pi609 & n28236;
  assign n28243 = ~n28241 & ~n28242;
  assign n28244 = pi1155 & ~n28243;
  assign n28245 = ~n16537 & ~n28237;
  assign n28246 = ~pi609 & n28236;
  assign n28247 = ~n28245 & ~n28246;
  assign n28248 = ~pi1155 & ~n28247;
  assign n28249 = ~n28244 & ~n28248;
  assign n28250 = pi785 & ~n28249;
  assign n28251 = ~n28240 & ~n28250;
  assign n28252 = ~pi781 & ~n28251;
  assign n28253 = pi618 & n28251;
  assign n28254 = ~pi618 & n28237;
  assign n28255 = pi1154 & ~n28254;
  assign n28256 = ~n28253 & n28255;
  assign n28257 = ~pi618 & n28251;
  assign n28258 = pi618 & n28237;
  assign n28259 = ~pi1154 & ~n28258;
  assign n28260 = ~n28257 & n28259;
  assign n28261 = ~n28256 & ~n28260;
  assign n28262 = pi781 & ~n28261;
  assign n28263 = ~n28252 & ~n28262;
  assign n28264 = ~pi789 & ~n28263;
  assign n28265 = pi619 & n28263;
  assign n28266 = ~pi619 & n28237;
  assign n28267 = pi1159 & ~n28266;
  assign n28268 = ~n28265 & n28267;
  assign n28269 = ~pi619 & n28263;
  assign n28270 = pi619 & n28237;
  assign n28271 = ~pi1159 & ~n28270;
  assign n28272 = ~n28269 & n28271;
  assign n28273 = ~n28268 & ~n28272;
  assign n28274 = pi789 & ~n28273;
  assign n28275 = ~n28264 & ~n28274;
  assign n28276 = ~n17355 & n28275;
  assign n28277 = n17355 & n28237;
  assign n28278 = ~n28276 & ~n28277;
  assign n28279 = ~n16124 & ~n28278;
  assign n28280 = n16124 & n28237;
  assign n28281 = ~n28279 & ~n28280;
  assign n28282 = pi647 & ~n28281;
  assign n28283 = pi628 & ~n28278;
  assign n28284 = n16593 & ~n28237;
  assign n28285 = ~pi703 & n28226;
  assign n28286 = ~pi186 & ~n16508;
  assign n28287 = n16744 & ~n28286;
  assign n28288 = pi186 & n17589;
  assign n28289 = ~pi186 & n17592;
  assign n28290 = ~pi38 & ~n28289;
  assign n28291 = ~n28288 & n28290;
  assign n28292 = ~n28287 & ~n28291;
  assign n28293 = pi703 & n28292;
  assign n28294 = ~n28285 & ~n28293;
  assign n28295 = n10020 & n28294;
  assign n28296 = ~n28225 & ~n28295;
  assign n28297 = ~pi778 & ~n28296;
  assign n28298 = pi625 & n28296;
  assign n28299 = pi1153 & ~n28298;
  assign n28300 = ~pi625 & n28237;
  assign n28301 = n28299 & ~n28300;
  assign n28302 = ~pi625 & n28296;
  assign n28303 = ~pi1153 & ~n28302;
  assign n28304 = pi625 & n28237;
  assign n28305 = n28303 & ~n28304;
  assign n28306 = ~n28301 & ~n28305;
  assign n28307 = pi778 & ~n28306;
  assign n28308 = ~n28297 & ~n28307;
  assign n28309 = ~n16593 & ~n28308;
  assign n28310 = ~n28284 & ~n28309;
  assign n28311 = ~n16589 & n28310;
  assign n28312 = n16589 & n28237;
  assign n28313 = ~n28311 & ~n28312;
  assign n28314 = pi619 & ~n28313;
  assign n28315 = pi618 & n28310;
  assign n28316 = pi609 & n28308;
  assign n28317 = pi625 & n28235;
  assign n28318 = ~pi703 & n28233;
  assign n28319 = ~pi186 & ~n18914;
  assign n28320 = pi186 & n18922;
  assign n28321 = ~pi752 & ~n28320;
  assign n28322 = ~n28319 & n28321;
  assign n28323 = pi186 & n18929;
  assign n28324 = ~pi186 & n18939;
  assign n28325 = ~n18932 & ~n28324;
  assign n28326 = pi752 & n28325;
  assign n28327 = ~n28323 & n28326;
  assign n28328 = ~n28322 & ~n28327;
  assign n28329 = pi703 & n28328;
  assign n28330 = ~n28318 & ~n28329;
  assign n28331 = n10020 & n28330;
  assign n28332 = ~n28225 & ~n28331;
  assign n28333 = ~pi625 & n28332;
  assign n28334 = ~pi1153 & ~n28333;
  assign n28335 = ~n28317 & n28334;
  assign n28336 = ~pi608 & ~n28301;
  assign n28337 = ~n28335 & n28336;
  assign n28338 = ~pi625 & n28235;
  assign n28339 = pi625 & n28332;
  assign n28340 = ~n28338 & ~n28339;
  assign n28341 = pi1153 & n28340;
  assign n28342 = ~n28305 & ~n28341;
  assign n28343 = pi608 & n28342;
  assign n28344 = ~n28337 & ~n28343;
  assign n28345 = pi778 & ~n28344;
  assign n28346 = ~pi778 & n28332;
  assign n28347 = ~n28345 & ~n28346;
  assign n28348 = ~pi609 & ~n28347;
  assign n28349 = ~pi1155 & ~n28348;
  assign n28350 = ~n28316 & n28349;
  assign n28351 = ~pi660 & ~n28244;
  assign n28352 = ~n28350 & n28351;
  assign n28353 = ~pi609 & n28308;
  assign n28354 = pi609 & ~n28347;
  assign n28355 = ~n28353 & ~n28354;
  assign n28356 = pi1155 & n28355;
  assign n28357 = ~n28248 & ~n28356;
  assign n28358 = pi660 & n28357;
  assign n28359 = ~n28352 & ~n28358;
  assign n28360 = pi785 & ~n28359;
  assign n28361 = ~pi785 & ~n28347;
  assign n28362 = ~n28360 & ~n28361;
  assign n28363 = ~pi618 & ~n28362;
  assign n28364 = ~pi1154 & ~n28363;
  assign n28365 = ~n28315 & n28364;
  assign n28366 = ~pi627 & ~n28256;
  assign n28367 = ~n28365 & n28366;
  assign n28368 = ~pi618 & n28310;
  assign n28369 = pi618 & ~n28362;
  assign n28370 = ~n28368 & ~n28369;
  assign n28371 = pi1154 & n28370;
  assign n28372 = ~n28260 & ~n28371;
  assign n28373 = pi627 & n28372;
  assign n28374 = ~n28367 & ~n28373;
  assign n28375 = pi781 & ~n28374;
  assign n28376 = ~pi781 & ~n28362;
  assign n28377 = ~n28375 & ~n28376;
  assign n28378 = ~pi619 & ~n28377;
  assign n28379 = ~pi1159 & ~n28378;
  assign n28380 = ~n28314 & n28379;
  assign n28381 = ~pi648 & ~n28268;
  assign n28382 = ~n28380 & n28381;
  assign n28383 = ~pi619 & ~n28313;
  assign n28384 = pi619 & ~n28377;
  assign n28385 = ~n28383 & ~n28384;
  assign n28386 = pi1159 & n28385;
  assign n28387 = ~n28272 & ~n28386;
  assign n28388 = pi648 & n28387;
  assign n28389 = ~n28382 & ~n28388;
  assign n28390 = pi789 & ~n28389;
  assign n28391 = ~pi789 & ~n28377;
  assign n28392 = ~n28390 & ~n28391;
  assign n28393 = ~pi788 & n28392;
  assign n28394 = pi626 & n28392;
  assign n28395 = n17159 & ~n28237;
  assign n28396 = ~n17159 & n28313;
  assign n28397 = ~n28395 & ~n28396;
  assign n28398 = ~pi626 & ~n28397;
  assign n28399 = pi641 & ~n28398;
  assign n28400 = ~n28394 & n28399;
  assign n28401 = pi626 & ~n28275;
  assign n28402 = ~pi626 & ~n28237;
  assign n28403 = ~pi641 & ~n28402;
  assign n28404 = ~n28401 & n28403;
  assign n28405 = pi1158 & ~n28404;
  assign n28406 = ~n28400 & n28405;
  assign n28407 = pi626 & ~n28237;
  assign n28408 = ~pi626 & ~n28275;
  assign n28409 = pi641 & ~n28408;
  assign n28410 = ~n28407 & n28409;
  assign n28411 = pi626 & ~n28397;
  assign n28412 = ~pi626 & n28392;
  assign n28413 = ~pi641 & ~n28412;
  assign n28414 = ~n28411 & n28413;
  assign n28415 = ~pi1158 & ~n28414;
  assign n28416 = ~n28410 & n28415;
  assign n28417 = ~n28406 & ~n28416;
  assign n28418 = pi788 & ~n28417;
  assign n28419 = ~n28393 & ~n28418;
  assign n28420 = ~pi628 & n28419;
  assign n28421 = ~pi1156 & ~n28420;
  assign n28422 = ~n28283 & n28421;
  assign n28423 = ~n17183 & n28397;
  assign n28424 = n17183 & n28237;
  assign n28425 = ~n28423 & ~n28424;
  assign n28426 = pi628 & ~n28425;
  assign n28427 = pi1156 & ~n28426;
  assign n28428 = ~pi628 & n28237;
  assign n28429 = n28427 & ~n28428;
  assign n28430 = ~pi629 & ~n28429;
  assign n28431 = ~n28422 & n28430;
  assign n28432 = ~pi628 & ~n28425;
  assign n28433 = pi628 & n28237;
  assign n28434 = ~pi1156 & ~n28433;
  assign n28435 = ~n28432 & n28434;
  assign n28436 = ~pi628 & ~n28278;
  assign n28437 = pi628 & n28419;
  assign n28438 = ~n28436 & ~n28437;
  assign n28439 = pi1156 & n28438;
  assign n28440 = ~n28435 & ~n28439;
  assign n28441 = pi629 & n28440;
  assign n28442 = ~n28431 & ~n28441;
  assign n28443 = pi792 & ~n28442;
  assign n28444 = ~pi792 & n28419;
  assign n28445 = ~n28443 & ~n28444;
  assign n28446 = ~pi647 & ~n28445;
  assign n28447 = ~pi1157 & ~n28446;
  assign n28448 = ~n28282 & n28447;
  assign n28449 = ~pi792 & n28425;
  assign n28450 = ~n28429 & ~n28435;
  assign n28451 = pi792 & ~n28450;
  assign n28452 = ~n28449 & ~n28451;
  assign n28453 = pi647 & n28452;
  assign n28454 = pi1157 & ~n28453;
  assign n28455 = ~pi647 & n28237;
  assign n28456 = n28454 & ~n28455;
  assign n28457 = ~pi630 & ~n28456;
  assign n28458 = ~n28448 & n28457;
  assign n28459 = ~pi647 & n28452;
  assign n28460 = pi647 & n28237;
  assign n28461 = ~pi1157 & ~n28460;
  assign n28462 = ~n28459 & n28461;
  assign n28463 = ~pi647 & ~n28281;
  assign n28464 = pi647 & ~n28445;
  assign n28465 = ~n28463 & ~n28464;
  assign n28466 = pi1157 & n28465;
  assign n28467 = ~n28462 & ~n28466;
  assign n28468 = pi630 & n28467;
  assign n28469 = ~n28458 & ~n28468;
  assign n28470 = pi787 & ~n28469;
  assign n28471 = ~pi787 & ~n28445;
  assign n28472 = ~n28470 & ~n28471;
  assign n28473 = ~pi790 & n28472;
  assign n28474 = pi644 & ~n28472;
  assign n28475 = ~pi787 & ~n28452;
  assign n28476 = ~n28456 & ~n28462;
  assign n28477 = pi787 & ~n28476;
  assign n28478 = ~n28475 & ~n28477;
  assign n28479 = ~pi644 & n28478;
  assign n28480 = pi715 & ~n28479;
  assign n28481 = ~n28474 & n28480;
  assign n28482 = ~pi644 & n28237;
  assign n28483 = n17247 & ~n28237;
  assign n28484 = ~n17247 & n28281;
  assign n28485 = ~n28483 & ~n28484;
  assign n28486 = pi644 & n28485;
  assign n28487 = ~pi715 & ~n28486;
  assign n28488 = ~n28482 & n28487;
  assign n28489 = ~n28481 & ~n28488;
  assign n28490 = pi1160 & n28489;
  assign n28491 = ~pi644 & n28485;
  assign n28492 = pi715 & ~n28491;
  assign n28493 = pi644 & n28237;
  assign n28494 = n28492 & ~n28493;
  assign n28495 = pi644 & n28478;
  assign n28496 = ~pi644 & ~n28472;
  assign n28497 = ~pi715 & ~n28496;
  assign n28498 = ~n28495 & n28497;
  assign n28499 = ~n28494 & ~n28498;
  assign n28500 = ~pi1160 & n28499;
  assign n28501 = ~n28490 & ~n28500;
  assign n28502 = pi790 & n28501;
  assign n28503 = ~n28473 & ~n28502;
  assign n28504 = ~po1038 & n28503;
  assign n28505 = ~pi186 & po1038;
  assign n28506 = ~pi832 & ~n28505;
  assign n28507 = ~n28504 & n28506;
  assign n28508 = ~pi186 & ~n2934;
  assign n28509 = ~pi752 & n16510;
  assign n28510 = ~n28508 & ~n28509;
  assign n28511 = ~n17273 & ~n28510;
  assign n28512 = ~pi785 & ~n28511;
  assign n28513 = ~n17279 & ~n28510;
  assign n28514 = pi1155 & ~n28513;
  assign n28515 = ~n17282 & n28511;
  assign n28516 = ~pi1155 & ~n28515;
  assign n28517 = ~n28514 & ~n28516;
  assign n28518 = pi785 & ~n28517;
  assign n28519 = ~n28512 & ~n28518;
  assign n28520 = ~pi781 & ~n28519;
  assign n28521 = ~n17289 & n28519;
  assign n28522 = pi1154 & ~n28521;
  assign n28523 = ~n17292 & n28519;
  assign n28524 = ~pi1154 & ~n28523;
  assign n28525 = ~n28522 & ~n28524;
  assign n28526 = pi781 & ~n28525;
  assign n28527 = ~n28520 & ~n28526;
  assign n28528 = ~pi789 & ~n28527;
  assign n28529 = pi619 & n28527;
  assign n28530 = ~pi619 & n28508;
  assign n28531 = pi1159 & ~n28530;
  assign n28532 = ~n28529 & n28531;
  assign n28533 = ~pi619 & n28527;
  assign n28534 = pi619 & n28508;
  assign n28535 = ~pi1159 & ~n28534;
  assign n28536 = ~n28533 & n28535;
  assign n28537 = ~n28532 & ~n28536;
  assign n28538 = pi789 & ~n28537;
  assign n28539 = ~n28528 & ~n28538;
  assign n28540 = ~n17355 & n28539;
  assign n28541 = n17355 & n28508;
  assign n28542 = ~n28540 & ~n28541;
  assign n28543 = ~n16124 & ~n28542;
  assign n28544 = n16124 & n28508;
  assign n28545 = ~n28543 & ~n28544;
  assign n28546 = ~n19987 & n28545;
  assign n28547 = pi703 & n16742;
  assign n28548 = ~n28508 & ~n28547;
  assign n28549 = ~pi778 & n28548;
  assign n28550 = ~pi625 & n28547;
  assign n28551 = ~n28548 & ~n28550;
  assign n28552 = pi1153 & ~n28551;
  assign n28553 = ~pi1153 & ~n28508;
  assign n28554 = ~n28550 & n28553;
  assign n28555 = ~n28552 & ~n28554;
  assign n28556 = pi778 & ~n28555;
  assign n28557 = ~n28549 & ~n28556;
  assign n28558 = ~n17338 & n28557;
  assign n28559 = ~n17340 & n28558;
  assign n28560 = ~n17342 & n28559;
  assign n28561 = ~n17425 & n28560;
  assign n28562 = ~n17452 & n28561;
  assign n28563 = ~pi647 & n28562;
  assign n28564 = pi647 & n28508;
  assign n28565 = ~pi1157 & ~n28564;
  assign n28566 = ~n28563 & n28565;
  assign n28567 = ~pi647 & n28508;
  assign n28568 = pi647 & n28562;
  assign n28569 = pi1157 & ~n28568;
  assign n28570 = ~n28567 & n28569;
  assign n28571 = ~n28566 & ~n28570;
  assign n28572 = ~n17246 & ~n28571;
  assign n28573 = ~n28546 & ~n28572;
  assign n28574 = pi787 & ~n28573;
  assign n28575 = ~pi626 & ~n28539;
  assign n28576 = pi626 & ~n28508;
  assign n28577 = n17181 & ~n28576;
  assign n28578 = ~n28575 & n28577;
  assign n28579 = n17350 & n28560;
  assign n28580 = pi626 & ~n28539;
  assign n28581 = ~pi626 & ~n28508;
  assign n28582 = n17180 & ~n28581;
  assign n28583 = ~n28580 & n28582;
  assign n28584 = ~n28579 & ~n28583;
  assign n28585 = ~n28578 & n28584;
  assign n28586 = pi788 & ~n28585;
  assign n28587 = pi618 & n28558;
  assign n28588 = pi609 & n28557;
  assign n28589 = ~n16393 & ~n28548;
  assign n28590 = pi625 & n28589;
  assign n28591 = n28510 & ~n28589;
  assign n28592 = ~n28590 & ~n28591;
  assign n28593 = n28553 & ~n28592;
  assign n28594 = ~pi608 & ~n28552;
  assign n28595 = ~n28593 & n28594;
  assign n28596 = pi1153 & ~n28590;
  assign n28597 = n28510 & n28596;
  assign n28598 = ~n28554 & ~n28597;
  assign n28599 = pi608 & n28598;
  assign n28600 = ~n28595 & ~n28599;
  assign n28601 = pi778 & ~n28600;
  assign n28602 = ~pi778 & ~n28591;
  assign n28603 = ~n28601 & ~n28602;
  assign n28604 = ~pi609 & ~n28603;
  assign n28605 = ~pi1155 & ~n28604;
  assign n28606 = ~n28588 & n28605;
  assign n28607 = ~pi660 & ~n28514;
  assign n28608 = ~n28606 & n28607;
  assign n28609 = ~pi609 & n28557;
  assign n28610 = pi609 & ~n28603;
  assign n28611 = ~n28609 & ~n28610;
  assign n28612 = pi1155 & n28611;
  assign n28613 = ~n28516 & ~n28612;
  assign n28614 = pi660 & n28613;
  assign n28615 = ~n28608 & ~n28614;
  assign n28616 = pi785 & ~n28615;
  assign n28617 = ~pi785 & ~n28603;
  assign n28618 = ~n28616 & ~n28617;
  assign n28619 = ~pi618 & ~n28618;
  assign n28620 = ~pi1154 & ~n28619;
  assign n28621 = ~n28587 & n28620;
  assign n28622 = ~pi627 & ~n28522;
  assign n28623 = ~n28621 & n28622;
  assign n28624 = ~pi618 & n28558;
  assign n28625 = pi618 & ~n28618;
  assign n28626 = ~n28624 & ~n28625;
  assign n28627 = pi1154 & n28626;
  assign n28628 = ~n28524 & ~n28627;
  assign n28629 = pi627 & n28628;
  assign n28630 = ~n28623 & ~n28629;
  assign n28631 = pi781 & ~n28630;
  assign n28632 = ~pi781 & ~n28618;
  assign n28633 = ~n28631 & ~n28632;
  assign n28634 = ~pi619 & ~n28633;
  assign n28635 = pi619 & n28559;
  assign n28636 = ~pi1159 & ~n28635;
  assign n28637 = ~n28634 & n28636;
  assign n28638 = ~pi648 & ~n28637;
  assign n28639 = ~n28532 & n28638;
  assign n28640 = ~pi619 & n28559;
  assign n28641 = pi619 & ~n28633;
  assign n28642 = ~n28640 & ~n28641;
  assign n28643 = pi1159 & n28642;
  assign n28644 = ~n28536 & ~n28643;
  assign n28645 = pi648 & n28644;
  assign n28646 = ~n28639 & ~n28645;
  assign n28647 = pi789 & n28646;
  assign n28648 = ~pi789 & n28633;
  assign n28649 = n17356 & ~n28648;
  assign n28650 = ~n28647 & n28649;
  assign n28651 = ~n28586 & ~n28650;
  assign n28652 = n19788 & ~n28651;
  assign n28653 = n20275 & n28561;
  assign n28654 = n17449 & ~n28542;
  assign n28655 = ~pi629 & ~n28654;
  assign n28656 = ~n28653 & n28655;
  assign n28657 = n17448 & ~n28542;
  assign n28658 = n20281 & n28561;
  assign n28659 = pi629 & ~n28658;
  assign n28660 = ~n28657 & n28659;
  assign n28661 = ~n28656 & ~n28660;
  assign n28662 = pi792 & n28661;
  assign n28663 = n19637 & ~n28662;
  assign n28664 = ~n28652 & n28663;
  assign n28665 = ~n28574 & ~n28664;
  assign n28666 = pi644 & n28665;
  assign n28667 = ~pi787 & ~n28562;
  assign n28668 = pi787 & ~n28571;
  assign n28669 = ~n28667 & ~n28668;
  assign n28670 = ~pi644 & n28669;
  assign n28671 = pi715 & ~n28670;
  assign n28672 = ~n28666 & n28671;
  assign n28673 = ~n17247 & ~n28545;
  assign n28674 = n17247 & n28508;
  assign n28675 = ~n28673 & ~n28674;
  assign n28676 = pi644 & ~n28675;
  assign n28677 = ~pi644 & n28508;
  assign n28678 = ~pi715 & ~n28677;
  assign n28679 = ~n28676 & n28678;
  assign n28680 = pi1160 & ~n28679;
  assign n28681 = ~n28672 & n28680;
  assign n28682 = ~pi644 & ~n28675;
  assign n28683 = pi715 & ~n28682;
  assign n28684 = pi644 & n28508;
  assign n28685 = n28683 & ~n28684;
  assign n28686 = pi644 & n28669;
  assign n28687 = ~pi644 & n28665;
  assign n28688 = ~pi715 & ~n28687;
  assign n28689 = ~n28686 & n28688;
  assign n28690 = ~pi1160 & ~n28689;
  assign n28691 = ~n28685 & n28690;
  assign n28692 = ~n28681 & ~n28691;
  assign n28693 = pi790 & ~n28692;
  assign n28694 = ~pi790 & n28665;
  assign n28695 = pi832 & ~n28694;
  assign n28696 = ~n28693 & n28695;
  assign po343 = ~n28507 & ~n28696;
  assign n28698 = pi187 & ~n10020;
  assign n28699 = ~pi770 & ~n18808;
  assign n28700 = ~n20507 & ~n28699;
  assign n28701 = ~pi187 & ~n28700;
  assign n28702 = ~pi187 & ~n18802;
  assign n28703 = ~pi770 & ~n28702;
  assign n28704 = ~n23777 & n28703;
  assign n28705 = ~n28701 & ~n28704;
  assign n28706 = n10020 & n28705;
  assign n28707 = ~n28698 & ~n28706;
  assign n28708 = ~n16521 & ~n28707;
  assign n28709 = ~pi187 & ~n16527;
  assign n28710 = n16521 & ~n28709;
  assign n28711 = ~n28708 & ~n28710;
  assign n28712 = ~pi785 & ~n28711;
  assign n28713 = ~n16532 & ~n28709;
  assign n28714 = pi609 & n28708;
  assign n28715 = ~n28713 & ~n28714;
  assign n28716 = pi1155 & ~n28715;
  assign n28717 = ~n16537 & ~n28709;
  assign n28718 = ~pi609 & n28708;
  assign n28719 = ~n28717 & ~n28718;
  assign n28720 = ~pi1155 & ~n28719;
  assign n28721 = ~n28716 & ~n28720;
  assign n28722 = pi785 & ~n28721;
  assign n28723 = ~n28712 & ~n28722;
  assign n28724 = ~pi781 & ~n28723;
  assign n28725 = pi618 & n28723;
  assign n28726 = ~pi618 & n28709;
  assign n28727 = pi1154 & ~n28726;
  assign n28728 = ~n28725 & n28727;
  assign n28729 = ~pi618 & n28723;
  assign n28730 = pi618 & n28709;
  assign n28731 = ~pi1154 & ~n28730;
  assign n28732 = ~n28729 & n28731;
  assign n28733 = ~n28728 & ~n28732;
  assign n28734 = pi781 & ~n28733;
  assign n28735 = ~n28724 & ~n28734;
  assign n28736 = ~pi789 & ~n28735;
  assign n28737 = pi619 & n28735;
  assign n28738 = ~pi619 & n28709;
  assign n28739 = pi1159 & ~n28738;
  assign n28740 = ~n28737 & n28739;
  assign n28741 = ~pi619 & n28735;
  assign n28742 = pi619 & n28709;
  assign n28743 = ~pi1159 & ~n28742;
  assign n28744 = ~n28741 & n28743;
  assign n28745 = ~n28740 & ~n28744;
  assign n28746 = pi789 & ~n28745;
  assign n28747 = ~n28736 & ~n28746;
  assign n28748 = ~n17355 & n28747;
  assign n28749 = n17355 & n28709;
  assign n28750 = ~n28748 & ~n28749;
  assign n28751 = ~n16124 & ~n28750;
  assign n28752 = n16124 & n28709;
  assign n28753 = ~n28751 & ~n28752;
  assign n28754 = pi647 & ~n28753;
  assign n28755 = pi628 & ~n28750;
  assign n28756 = n16593 & ~n28709;
  assign n28757 = pi187 & n17589;
  assign n28758 = ~pi187 & n17592;
  assign n28759 = ~pi38 & ~n28758;
  assign n28760 = ~n28757 & n28759;
  assign n28761 = ~pi187 & ~n16508;
  assign n28762 = n16744 & ~n28761;
  assign n28763 = pi726 & ~n28762;
  assign n28764 = ~n28760 & n28763;
  assign n28765 = ~pi187 & ~pi726;
  assign n28766 = ~n16526 & n28765;
  assign n28767 = ~n28764 & ~n28766;
  assign n28768 = n10020 & n28767;
  assign n28769 = ~n28698 & ~n28768;
  assign n28770 = ~pi778 & ~n28769;
  assign n28771 = pi625 & n28769;
  assign n28772 = pi1153 & ~n28771;
  assign n28773 = ~pi625 & n28709;
  assign n28774 = n28772 & ~n28773;
  assign n28775 = ~pi625 & n28769;
  assign n28776 = ~pi1153 & ~n28775;
  assign n28777 = pi625 & n28709;
  assign n28778 = n28776 & ~n28777;
  assign n28779 = ~n28774 & ~n28778;
  assign n28780 = pi778 & ~n28779;
  assign n28781 = ~n28770 & ~n28780;
  assign n28782 = ~n16593 & ~n28781;
  assign n28783 = ~n28756 & ~n28782;
  assign n28784 = ~n16589 & n28783;
  assign n28785 = n16589 & n28709;
  assign n28786 = ~n28784 & ~n28785;
  assign n28787 = pi619 & ~n28786;
  assign n28788 = pi618 & n28783;
  assign n28789 = pi609 & n28781;
  assign n28790 = pi625 & n28707;
  assign n28791 = ~pi726 & ~n28705;
  assign n28792 = ~pi187 & ~n18914;
  assign n28793 = pi187 & n18922;
  assign n28794 = ~pi770 & ~n28793;
  assign n28795 = ~n28792 & n28794;
  assign n28796 = pi187 & n18929;
  assign n28797 = ~pi187 & n18939;
  assign n28798 = ~n18932 & ~n28797;
  assign n28799 = pi770 & n28798;
  assign n28800 = ~n28796 & n28799;
  assign n28801 = ~n28795 & ~n28800;
  assign n28802 = pi726 & n28801;
  assign n28803 = ~n28791 & ~n28802;
  assign n28804 = n10020 & n28803;
  assign n28805 = ~n28698 & ~n28804;
  assign n28806 = ~pi625 & n28805;
  assign n28807 = ~pi1153 & ~n28806;
  assign n28808 = ~n28790 & n28807;
  assign n28809 = ~pi608 & ~n28774;
  assign n28810 = ~n28808 & n28809;
  assign n28811 = ~pi625 & n28707;
  assign n28812 = pi625 & n28805;
  assign n28813 = ~n28811 & ~n28812;
  assign n28814 = pi1153 & n28813;
  assign n28815 = ~n28778 & ~n28814;
  assign n28816 = pi608 & n28815;
  assign n28817 = ~n28810 & ~n28816;
  assign n28818 = pi778 & ~n28817;
  assign n28819 = ~pi778 & n28805;
  assign n28820 = ~n28818 & ~n28819;
  assign n28821 = ~pi609 & ~n28820;
  assign n28822 = ~pi1155 & ~n28821;
  assign n28823 = ~n28789 & n28822;
  assign n28824 = ~pi660 & ~n28716;
  assign n28825 = ~n28823 & n28824;
  assign n28826 = ~pi609 & n28781;
  assign n28827 = pi609 & ~n28820;
  assign n28828 = ~n28826 & ~n28827;
  assign n28829 = pi1155 & n28828;
  assign n28830 = ~n28720 & ~n28829;
  assign n28831 = pi660 & n28830;
  assign n28832 = ~n28825 & ~n28831;
  assign n28833 = pi785 & ~n28832;
  assign n28834 = ~pi785 & ~n28820;
  assign n28835 = ~n28833 & ~n28834;
  assign n28836 = ~pi618 & ~n28835;
  assign n28837 = ~pi1154 & ~n28836;
  assign n28838 = ~n28788 & n28837;
  assign n28839 = ~pi627 & ~n28728;
  assign n28840 = ~n28838 & n28839;
  assign n28841 = ~pi618 & n28783;
  assign n28842 = pi618 & ~n28835;
  assign n28843 = ~n28841 & ~n28842;
  assign n28844 = pi1154 & n28843;
  assign n28845 = ~n28732 & ~n28844;
  assign n28846 = pi627 & n28845;
  assign n28847 = ~n28840 & ~n28846;
  assign n28848 = pi781 & ~n28847;
  assign n28849 = ~pi781 & ~n28835;
  assign n28850 = ~n28848 & ~n28849;
  assign n28851 = ~pi619 & ~n28850;
  assign n28852 = ~pi1159 & ~n28851;
  assign n28853 = ~n28787 & n28852;
  assign n28854 = ~pi648 & ~n28740;
  assign n28855 = ~n28853 & n28854;
  assign n28856 = ~pi619 & ~n28786;
  assign n28857 = pi619 & ~n28850;
  assign n28858 = ~n28856 & ~n28857;
  assign n28859 = pi1159 & n28858;
  assign n28860 = ~n28744 & ~n28859;
  assign n28861 = pi648 & n28860;
  assign n28862 = ~n28855 & ~n28861;
  assign n28863 = pi789 & ~n28862;
  assign n28864 = ~pi789 & ~n28850;
  assign n28865 = ~n28863 & ~n28864;
  assign n28866 = ~pi788 & n28865;
  assign n28867 = pi626 & n28865;
  assign n28868 = n17159 & ~n28709;
  assign n28869 = ~n17159 & n28786;
  assign n28870 = ~n28868 & ~n28869;
  assign n28871 = ~pi626 & ~n28870;
  assign n28872 = pi641 & ~n28871;
  assign n28873 = ~n28867 & n28872;
  assign n28874 = pi626 & ~n28747;
  assign n28875 = ~pi626 & ~n28709;
  assign n28876 = ~pi641 & ~n28875;
  assign n28877 = ~n28874 & n28876;
  assign n28878 = pi1158 & ~n28877;
  assign n28879 = ~n28873 & n28878;
  assign n28880 = pi626 & ~n28709;
  assign n28881 = ~pi626 & ~n28747;
  assign n28882 = pi641 & ~n28881;
  assign n28883 = ~n28880 & n28882;
  assign n28884 = pi626 & ~n28870;
  assign n28885 = ~pi626 & n28865;
  assign n28886 = ~pi641 & ~n28885;
  assign n28887 = ~n28884 & n28886;
  assign n28888 = ~pi1158 & ~n28887;
  assign n28889 = ~n28883 & n28888;
  assign n28890 = ~n28879 & ~n28889;
  assign n28891 = pi788 & ~n28890;
  assign n28892 = ~n28866 & ~n28891;
  assign n28893 = ~pi628 & n28892;
  assign n28894 = ~pi1156 & ~n28893;
  assign n28895 = ~n28755 & n28894;
  assign n28896 = ~n17183 & n28870;
  assign n28897 = n17183 & n28709;
  assign n28898 = ~n28896 & ~n28897;
  assign n28899 = pi628 & ~n28898;
  assign n28900 = pi1156 & ~n28899;
  assign n28901 = ~pi628 & n28709;
  assign n28902 = n28900 & ~n28901;
  assign n28903 = ~pi629 & ~n28902;
  assign n28904 = ~n28895 & n28903;
  assign n28905 = ~pi628 & ~n28898;
  assign n28906 = pi628 & n28709;
  assign n28907 = ~pi1156 & ~n28906;
  assign n28908 = ~n28905 & n28907;
  assign n28909 = ~pi628 & ~n28750;
  assign n28910 = pi628 & n28892;
  assign n28911 = ~n28909 & ~n28910;
  assign n28912 = pi1156 & n28911;
  assign n28913 = ~n28908 & ~n28912;
  assign n28914 = pi629 & n28913;
  assign n28915 = ~n28904 & ~n28914;
  assign n28916 = pi792 & ~n28915;
  assign n28917 = ~pi792 & n28892;
  assign n28918 = ~n28916 & ~n28917;
  assign n28919 = ~pi647 & ~n28918;
  assign n28920 = ~pi1157 & ~n28919;
  assign n28921 = ~n28754 & n28920;
  assign n28922 = ~pi792 & n28898;
  assign n28923 = ~n28902 & ~n28908;
  assign n28924 = pi792 & ~n28923;
  assign n28925 = ~n28922 & ~n28924;
  assign n28926 = pi647 & n28925;
  assign n28927 = pi1157 & ~n28926;
  assign n28928 = ~pi647 & n28709;
  assign n28929 = n28927 & ~n28928;
  assign n28930 = ~pi630 & ~n28929;
  assign n28931 = ~n28921 & n28930;
  assign n28932 = ~pi647 & n28925;
  assign n28933 = pi647 & n28709;
  assign n28934 = ~pi1157 & ~n28933;
  assign n28935 = ~n28932 & n28934;
  assign n28936 = ~pi647 & ~n28753;
  assign n28937 = pi647 & ~n28918;
  assign n28938 = ~n28936 & ~n28937;
  assign n28939 = pi1157 & n28938;
  assign n28940 = ~n28935 & ~n28939;
  assign n28941 = pi630 & n28940;
  assign n28942 = ~n28931 & ~n28941;
  assign n28943 = pi787 & ~n28942;
  assign n28944 = ~pi787 & ~n28918;
  assign n28945 = ~n28943 & ~n28944;
  assign n28946 = ~pi790 & n28945;
  assign n28947 = pi644 & ~n28945;
  assign n28948 = ~pi787 & ~n28925;
  assign n28949 = ~n28929 & ~n28935;
  assign n28950 = pi787 & ~n28949;
  assign n28951 = ~n28948 & ~n28950;
  assign n28952 = ~pi644 & n28951;
  assign n28953 = pi715 & ~n28952;
  assign n28954 = ~n28947 & n28953;
  assign n28955 = ~pi644 & n28709;
  assign n28956 = n17247 & ~n28709;
  assign n28957 = ~n17247 & n28753;
  assign n28958 = ~n28956 & ~n28957;
  assign n28959 = pi644 & n28958;
  assign n28960 = ~pi715 & ~n28959;
  assign n28961 = ~n28955 & n28960;
  assign n28962 = ~n28954 & ~n28961;
  assign n28963 = pi1160 & n28962;
  assign n28964 = ~pi644 & n28958;
  assign n28965 = pi715 & ~n28964;
  assign n28966 = pi644 & n28709;
  assign n28967 = n28965 & ~n28966;
  assign n28968 = pi644 & n28951;
  assign n28969 = ~pi644 & ~n28945;
  assign n28970 = ~pi715 & ~n28969;
  assign n28971 = ~n28968 & n28970;
  assign n28972 = ~n28967 & ~n28971;
  assign n28973 = ~pi1160 & n28972;
  assign n28974 = ~n28963 & ~n28973;
  assign n28975 = pi790 & n28974;
  assign n28976 = ~n28946 & ~n28975;
  assign n28977 = ~po1038 & n28976;
  assign n28978 = ~pi187 & po1038;
  assign n28979 = ~pi832 & ~n28978;
  assign n28980 = ~n28977 & n28979;
  assign n28981 = ~pi187 & ~n2934;
  assign n28982 = ~pi770 & n16510;
  assign n28983 = ~n28981 & ~n28982;
  assign n28984 = ~n17273 & ~n28983;
  assign n28985 = ~pi785 & ~n28984;
  assign n28986 = ~n17279 & ~n28983;
  assign n28987 = pi1155 & ~n28986;
  assign n28988 = ~n17282 & n28984;
  assign n28989 = ~pi1155 & ~n28988;
  assign n28990 = ~n28987 & ~n28989;
  assign n28991 = pi785 & ~n28990;
  assign n28992 = ~n28985 & ~n28991;
  assign n28993 = ~pi781 & ~n28992;
  assign n28994 = ~n17289 & n28992;
  assign n28995 = pi1154 & ~n28994;
  assign n28996 = ~n17292 & n28992;
  assign n28997 = ~pi1154 & ~n28996;
  assign n28998 = ~n28995 & ~n28997;
  assign n28999 = pi781 & ~n28998;
  assign n29000 = ~n28993 & ~n28999;
  assign n29001 = ~pi789 & ~n29000;
  assign n29002 = pi619 & n29000;
  assign n29003 = ~pi619 & n28981;
  assign n29004 = pi1159 & ~n29003;
  assign n29005 = ~n29002 & n29004;
  assign n29006 = ~pi619 & n29000;
  assign n29007 = pi619 & n28981;
  assign n29008 = ~pi1159 & ~n29007;
  assign n29009 = ~n29006 & n29008;
  assign n29010 = ~n29005 & ~n29009;
  assign n29011 = pi789 & ~n29010;
  assign n29012 = ~n29001 & ~n29011;
  assign n29013 = ~n17355 & n29012;
  assign n29014 = n17355 & n28981;
  assign n29015 = ~n29013 & ~n29014;
  assign n29016 = ~n16124 & ~n29015;
  assign n29017 = n16124 & n28981;
  assign n29018 = ~n29016 & ~n29017;
  assign n29019 = ~n19987 & n29018;
  assign n29020 = pi726 & n16742;
  assign n29021 = ~n28981 & ~n29020;
  assign n29022 = ~pi778 & n29021;
  assign n29023 = ~pi625 & n29020;
  assign n29024 = ~n29021 & ~n29023;
  assign n29025 = pi1153 & ~n29024;
  assign n29026 = ~pi1153 & ~n28981;
  assign n29027 = ~n29023 & n29026;
  assign n29028 = ~n29025 & ~n29027;
  assign n29029 = pi778 & ~n29028;
  assign n29030 = ~n29022 & ~n29029;
  assign n29031 = ~n17338 & n29030;
  assign n29032 = ~n17340 & n29031;
  assign n29033 = ~n17342 & n29032;
  assign n29034 = ~n17425 & n29033;
  assign n29035 = ~n17452 & n29034;
  assign n29036 = ~pi647 & n29035;
  assign n29037 = pi647 & n28981;
  assign n29038 = ~pi1157 & ~n29037;
  assign n29039 = ~n29036 & n29038;
  assign n29040 = ~pi647 & n28981;
  assign n29041 = pi647 & n29035;
  assign n29042 = pi1157 & ~n29041;
  assign n29043 = ~n29040 & n29042;
  assign n29044 = ~n29039 & ~n29043;
  assign n29045 = ~n17246 & ~n29044;
  assign n29046 = ~n29019 & ~n29045;
  assign n29047 = pi787 & ~n29046;
  assign n29048 = ~pi626 & ~n29012;
  assign n29049 = pi626 & ~n28981;
  assign n29050 = n17181 & ~n29049;
  assign n29051 = ~n29048 & n29050;
  assign n29052 = n17350 & n29033;
  assign n29053 = pi626 & ~n29012;
  assign n29054 = ~pi626 & ~n28981;
  assign n29055 = n17180 & ~n29054;
  assign n29056 = ~n29053 & n29055;
  assign n29057 = ~n29052 & ~n29056;
  assign n29058 = ~n29051 & n29057;
  assign n29059 = pi788 & ~n29058;
  assign n29060 = pi618 & n29031;
  assign n29061 = pi609 & n29030;
  assign n29062 = ~n16393 & ~n29021;
  assign n29063 = pi625 & n29062;
  assign n29064 = n28983 & ~n29062;
  assign n29065 = ~n29063 & ~n29064;
  assign n29066 = n29026 & ~n29065;
  assign n29067 = ~pi608 & ~n29025;
  assign n29068 = ~n29066 & n29067;
  assign n29069 = pi1153 & ~n29063;
  assign n29070 = n28983 & n29069;
  assign n29071 = ~n29027 & ~n29070;
  assign n29072 = pi608 & n29071;
  assign n29073 = ~n29068 & ~n29072;
  assign n29074 = pi778 & ~n29073;
  assign n29075 = ~pi778 & ~n29064;
  assign n29076 = ~n29074 & ~n29075;
  assign n29077 = ~pi609 & ~n29076;
  assign n29078 = ~pi1155 & ~n29077;
  assign n29079 = ~n29061 & n29078;
  assign n29080 = ~pi660 & ~n28987;
  assign n29081 = ~n29079 & n29080;
  assign n29082 = ~pi609 & n29030;
  assign n29083 = pi609 & ~n29076;
  assign n29084 = ~n29082 & ~n29083;
  assign n29085 = pi1155 & n29084;
  assign n29086 = ~n28989 & ~n29085;
  assign n29087 = pi660 & n29086;
  assign n29088 = ~n29081 & ~n29087;
  assign n29089 = pi785 & ~n29088;
  assign n29090 = ~pi785 & ~n29076;
  assign n29091 = ~n29089 & ~n29090;
  assign n29092 = ~pi618 & ~n29091;
  assign n29093 = ~pi1154 & ~n29092;
  assign n29094 = ~n29060 & n29093;
  assign n29095 = ~pi627 & ~n28995;
  assign n29096 = ~n29094 & n29095;
  assign n29097 = ~pi618 & n29031;
  assign n29098 = pi618 & ~n29091;
  assign n29099 = ~n29097 & ~n29098;
  assign n29100 = pi1154 & n29099;
  assign n29101 = ~n28997 & ~n29100;
  assign n29102 = pi627 & n29101;
  assign n29103 = ~n29096 & ~n29102;
  assign n29104 = pi781 & ~n29103;
  assign n29105 = ~pi781 & ~n29091;
  assign n29106 = ~n29104 & ~n29105;
  assign n29107 = ~pi619 & ~n29106;
  assign n29108 = pi619 & n29032;
  assign n29109 = ~pi1159 & ~n29108;
  assign n29110 = ~n29107 & n29109;
  assign n29111 = ~pi648 & ~n29110;
  assign n29112 = ~n29005 & n29111;
  assign n29113 = ~pi619 & n29032;
  assign n29114 = pi619 & ~n29106;
  assign n29115 = ~n29113 & ~n29114;
  assign n29116 = pi1159 & n29115;
  assign n29117 = ~n29009 & ~n29116;
  assign n29118 = pi648 & n29117;
  assign n29119 = ~n29112 & ~n29118;
  assign n29120 = pi789 & n29119;
  assign n29121 = ~pi789 & n29106;
  assign n29122 = n17356 & ~n29121;
  assign n29123 = ~n29120 & n29122;
  assign n29124 = ~n29059 & ~n29123;
  assign n29125 = n19788 & ~n29124;
  assign n29126 = n20275 & n29034;
  assign n29127 = n17449 & ~n29015;
  assign n29128 = ~pi629 & ~n29127;
  assign n29129 = ~n29126 & n29128;
  assign n29130 = n17448 & ~n29015;
  assign n29131 = n20281 & n29034;
  assign n29132 = pi629 & ~n29131;
  assign n29133 = ~n29130 & n29132;
  assign n29134 = ~n29129 & ~n29133;
  assign n29135 = pi792 & n29134;
  assign n29136 = n19637 & ~n29135;
  assign n29137 = ~n29125 & n29136;
  assign n29138 = ~n29047 & ~n29137;
  assign n29139 = pi644 & n29138;
  assign n29140 = ~pi787 & ~n29035;
  assign n29141 = pi787 & ~n29044;
  assign n29142 = ~n29140 & ~n29141;
  assign n29143 = ~pi644 & n29142;
  assign n29144 = pi715 & ~n29143;
  assign n29145 = ~n29139 & n29144;
  assign n29146 = ~n17247 & ~n29018;
  assign n29147 = n17247 & n28981;
  assign n29148 = ~n29146 & ~n29147;
  assign n29149 = pi644 & ~n29148;
  assign n29150 = ~pi644 & n28981;
  assign n29151 = ~pi715 & ~n29150;
  assign n29152 = ~n29149 & n29151;
  assign n29153 = pi1160 & ~n29152;
  assign n29154 = ~n29145 & n29153;
  assign n29155 = ~pi644 & ~n29148;
  assign n29156 = pi715 & ~n29155;
  assign n29157 = pi644 & n28981;
  assign n29158 = n29156 & ~n29157;
  assign n29159 = pi644 & n29142;
  assign n29160 = ~pi644 & n29138;
  assign n29161 = ~pi715 & ~n29160;
  assign n29162 = ~n29159 & n29161;
  assign n29163 = ~pi1160 & ~n29162;
  assign n29164 = ~n29158 & n29163;
  assign n29165 = ~n29154 & ~n29164;
  assign n29166 = pi790 & ~n29165;
  assign n29167 = ~pi790 & n29138;
  assign n29168 = pi832 & ~n29167;
  assign n29169 = ~n29166 & n29168;
  assign po344 = ~n28980 & ~n29169;
  assign n29171 = pi188 & ~n10020;
  assign n29172 = ~pi768 & ~n18808;
  assign n29173 = ~n21707 & ~n29172;
  assign n29174 = ~pi188 & ~n29173;
  assign n29175 = ~pi188 & ~n18802;
  assign n29176 = ~pi768 & ~n29175;
  assign n29177 = ~n23777 & n29176;
  assign n29178 = ~n29174 & ~n29177;
  assign n29179 = n10020 & n29178;
  assign n29180 = ~n29171 & ~n29179;
  assign n29181 = ~n16521 & ~n29180;
  assign n29182 = ~pi188 & ~n16527;
  assign n29183 = n16521 & ~n29182;
  assign n29184 = ~n29181 & ~n29183;
  assign n29185 = ~pi785 & ~n29184;
  assign n29186 = ~n16532 & ~n29182;
  assign n29187 = pi609 & n29181;
  assign n29188 = ~n29186 & ~n29187;
  assign n29189 = pi1155 & ~n29188;
  assign n29190 = ~n16537 & ~n29182;
  assign n29191 = ~pi609 & n29181;
  assign n29192 = ~n29190 & ~n29191;
  assign n29193 = ~pi1155 & ~n29192;
  assign n29194 = ~n29189 & ~n29193;
  assign n29195 = pi785 & ~n29194;
  assign n29196 = ~n29185 & ~n29195;
  assign n29197 = ~pi781 & ~n29196;
  assign n29198 = pi618 & n29196;
  assign n29199 = ~pi618 & n29182;
  assign n29200 = pi1154 & ~n29199;
  assign n29201 = ~n29198 & n29200;
  assign n29202 = ~pi618 & n29196;
  assign n29203 = pi618 & n29182;
  assign n29204 = ~pi1154 & ~n29203;
  assign n29205 = ~n29202 & n29204;
  assign n29206 = ~n29201 & ~n29205;
  assign n29207 = pi781 & ~n29206;
  assign n29208 = ~n29197 & ~n29207;
  assign n29209 = ~pi789 & ~n29208;
  assign n29210 = pi619 & n29208;
  assign n29211 = ~pi619 & n29182;
  assign n29212 = pi1159 & ~n29211;
  assign n29213 = ~n29210 & n29212;
  assign n29214 = ~pi619 & n29208;
  assign n29215 = pi619 & n29182;
  assign n29216 = ~pi1159 & ~n29215;
  assign n29217 = ~n29214 & n29216;
  assign n29218 = ~n29213 & ~n29217;
  assign n29219 = pi789 & ~n29218;
  assign n29220 = ~n29209 & ~n29219;
  assign n29221 = ~n17355 & n29220;
  assign n29222 = n17355 & n29182;
  assign n29223 = ~n29221 & ~n29222;
  assign n29224 = ~n16124 & ~n29223;
  assign n29225 = n16124 & n29182;
  assign n29226 = ~n29224 & ~n29225;
  assign n29227 = pi647 & ~n29226;
  assign n29228 = pi628 & ~n29223;
  assign n29229 = n16593 & ~n29182;
  assign n29230 = pi188 & n17589;
  assign n29231 = ~pi188 & n17592;
  assign n29232 = ~pi38 & ~n29231;
  assign n29233 = ~n29230 & n29232;
  assign n29234 = ~pi188 & ~n16508;
  assign n29235 = n16744 & ~n29234;
  assign n29236 = pi705 & ~n29235;
  assign n29237 = ~n29233 & n29236;
  assign n29238 = ~pi188 & ~pi705;
  assign n29239 = ~n16526 & n29238;
  assign n29240 = ~n29237 & ~n29239;
  assign n29241 = n10020 & n29240;
  assign n29242 = ~n29171 & ~n29241;
  assign n29243 = ~pi778 & ~n29242;
  assign n29244 = pi625 & n29242;
  assign n29245 = pi1153 & ~n29244;
  assign n29246 = ~pi625 & n29182;
  assign n29247 = n29245 & ~n29246;
  assign n29248 = ~pi625 & n29242;
  assign n29249 = ~pi1153 & ~n29248;
  assign n29250 = pi625 & n29182;
  assign n29251 = n29249 & ~n29250;
  assign n29252 = ~n29247 & ~n29251;
  assign n29253 = pi778 & ~n29252;
  assign n29254 = ~n29243 & ~n29253;
  assign n29255 = ~n16593 & ~n29254;
  assign n29256 = ~n29229 & ~n29255;
  assign n29257 = ~n16589 & n29256;
  assign n29258 = n16589 & n29182;
  assign n29259 = ~n29257 & ~n29258;
  assign n29260 = pi619 & ~n29259;
  assign n29261 = pi618 & n29256;
  assign n29262 = pi609 & n29254;
  assign n29263 = pi625 & n29180;
  assign n29264 = ~pi705 & ~n29178;
  assign n29265 = ~pi188 & ~n18914;
  assign n29266 = pi188 & n18922;
  assign n29267 = ~pi768 & ~n29266;
  assign n29268 = ~n29265 & n29267;
  assign n29269 = pi188 & n18929;
  assign n29270 = ~pi188 & n18939;
  assign n29271 = ~n18932 & ~n29270;
  assign n29272 = pi768 & n29271;
  assign n29273 = ~n29269 & n29272;
  assign n29274 = ~n29268 & ~n29273;
  assign n29275 = pi705 & n29274;
  assign n29276 = ~n29264 & ~n29275;
  assign n29277 = n10020 & n29276;
  assign n29278 = ~n29171 & ~n29277;
  assign n29279 = ~pi625 & n29278;
  assign n29280 = ~pi1153 & ~n29279;
  assign n29281 = ~n29263 & n29280;
  assign n29282 = ~pi608 & ~n29247;
  assign n29283 = ~n29281 & n29282;
  assign n29284 = ~pi625 & n29180;
  assign n29285 = pi625 & n29278;
  assign n29286 = ~n29284 & ~n29285;
  assign n29287 = pi1153 & n29286;
  assign n29288 = ~n29251 & ~n29287;
  assign n29289 = pi608 & n29288;
  assign n29290 = ~n29283 & ~n29289;
  assign n29291 = pi778 & ~n29290;
  assign n29292 = ~pi778 & n29278;
  assign n29293 = ~n29291 & ~n29292;
  assign n29294 = ~pi609 & ~n29293;
  assign n29295 = ~pi1155 & ~n29294;
  assign n29296 = ~n29262 & n29295;
  assign n29297 = ~pi660 & ~n29189;
  assign n29298 = ~n29296 & n29297;
  assign n29299 = ~pi609 & n29254;
  assign n29300 = pi609 & ~n29293;
  assign n29301 = ~n29299 & ~n29300;
  assign n29302 = pi1155 & n29301;
  assign n29303 = ~n29193 & ~n29302;
  assign n29304 = pi660 & n29303;
  assign n29305 = ~n29298 & ~n29304;
  assign n29306 = pi785 & ~n29305;
  assign n29307 = ~pi785 & ~n29293;
  assign n29308 = ~n29306 & ~n29307;
  assign n29309 = ~pi618 & ~n29308;
  assign n29310 = ~pi1154 & ~n29309;
  assign n29311 = ~n29261 & n29310;
  assign n29312 = ~pi627 & ~n29201;
  assign n29313 = ~n29311 & n29312;
  assign n29314 = ~pi618 & n29256;
  assign n29315 = pi618 & ~n29308;
  assign n29316 = ~n29314 & ~n29315;
  assign n29317 = pi1154 & n29316;
  assign n29318 = ~n29205 & ~n29317;
  assign n29319 = pi627 & n29318;
  assign n29320 = ~n29313 & ~n29319;
  assign n29321 = pi781 & ~n29320;
  assign n29322 = ~pi781 & ~n29308;
  assign n29323 = ~n29321 & ~n29322;
  assign n29324 = ~pi619 & ~n29323;
  assign n29325 = ~pi1159 & ~n29324;
  assign n29326 = ~n29260 & n29325;
  assign n29327 = ~pi648 & ~n29213;
  assign n29328 = ~n29326 & n29327;
  assign n29329 = ~pi619 & ~n29259;
  assign n29330 = pi619 & ~n29323;
  assign n29331 = ~n29329 & ~n29330;
  assign n29332 = pi1159 & n29331;
  assign n29333 = ~n29217 & ~n29332;
  assign n29334 = pi648 & n29333;
  assign n29335 = ~n29328 & ~n29334;
  assign n29336 = pi789 & ~n29335;
  assign n29337 = ~pi789 & ~n29323;
  assign n29338 = ~n29336 & ~n29337;
  assign n29339 = ~pi788 & n29338;
  assign n29340 = pi626 & n29338;
  assign n29341 = n17159 & ~n29182;
  assign n29342 = ~n17159 & n29259;
  assign n29343 = ~n29341 & ~n29342;
  assign n29344 = ~pi626 & ~n29343;
  assign n29345 = pi641 & ~n29344;
  assign n29346 = ~n29340 & n29345;
  assign n29347 = pi626 & ~n29220;
  assign n29348 = ~pi626 & ~n29182;
  assign n29349 = ~pi641 & ~n29348;
  assign n29350 = ~n29347 & n29349;
  assign n29351 = pi1158 & ~n29350;
  assign n29352 = ~n29346 & n29351;
  assign n29353 = pi626 & ~n29182;
  assign n29354 = ~pi626 & ~n29220;
  assign n29355 = pi641 & ~n29354;
  assign n29356 = ~n29353 & n29355;
  assign n29357 = pi626 & ~n29343;
  assign n29358 = ~pi626 & n29338;
  assign n29359 = ~pi641 & ~n29358;
  assign n29360 = ~n29357 & n29359;
  assign n29361 = ~pi1158 & ~n29360;
  assign n29362 = ~n29356 & n29361;
  assign n29363 = ~n29352 & ~n29362;
  assign n29364 = pi788 & ~n29363;
  assign n29365 = ~n29339 & ~n29364;
  assign n29366 = ~pi628 & n29365;
  assign n29367 = ~pi1156 & ~n29366;
  assign n29368 = ~n29228 & n29367;
  assign n29369 = ~n17183 & n29343;
  assign n29370 = n17183 & n29182;
  assign n29371 = ~n29369 & ~n29370;
  assign n29372 = pi628 & ~n29371;
  assign n29373 = pi1156 & ~n29372;
  assign n29374 = ~pi628 & n29182;
  assign n29375 = n29373 & ~n29374;
  assign n29376 = ~pi629 & ~n29375;
  assign n29377 = ~n29368 & n29376;
  assign n29378 = ~pi628 & ~n29371;
  assign n29379 = pi628 & n29182;
  assign n29380 = ~pi1156 & ~n29379;
  assign n29381 = ~n29378 & n29380;
  assign n29382 = ~pi628 & ~n29223;
  assign n29383 = pi628 & n29365;
  assign n29384 = ~n29382 & ~n29383;
  assign n29385 = pi1156 & n29384;
  assign n29386 = ~n29381 & ~n29385;
  assign n29387 = pi629 & n29386;
  assign n29388 = ~n29377 & ~n29387;
  assign n29389 = pi792 & ~n29388;
  assign n29390 = ~pi792 & n29365;
  assign n29391 = ~n29389 & ~n29390;
  assign n29392 = ~pi647 & ~n29391;
  assign n29393 = ~pi1157 & ~n29392;
  assign n29394 = ~n29227 & n29393;
  assign n29395 = ~pi792 & n29371;
  assign n29396 = ~n29375 & ~n29381;
  assign n29397 = pi792 & ~n29396;
  assign n29398 = ~n29395 & ~n29397;
  assign n29399 = pi647 & n29398;
  assign n29400 = pi1157 & ~n29399;
  assign n29401 = ~pi647 & n29182;
  assign n29402 = n29400 & ~n29401;
  assign n29403 = ~pi630 & ~n29402;
  assign n29404 = ~n29394 & n29403;
  assign n29405 = ~pi647 & n29398;
  assign n29406 = pi647 & n29182;
  assign n29407 = ~pi1157 & ~n29406;
  assign n29408 = ~n29405 & n29407;
  assign n29409 = ~pi647 & ~n29226;
  assign n29410 = pi647 & ~n29391;
  assign n29411 = ~n29409 & ~n29410;
  assign n29412 = pi1157 & n29411;
  assign n29413 = ~n29408 & ~n29412;
  assign n29414 = pi630 & n29413;
  assign n29415 = ~n29404 & ~n29414;
  assign n29416 = pi787 & ~n29415;
  assign n29417 = ~pi787 & ~n29391;
  assign n29418 = ~n29416 & ~n29417;
  assign n29419 = ~pi790 & n29418;
  assign n29420 = pi644 & ~n29418;
  assign n29421 = ~pi787 & ~n29398;
  assign n29422 = ~n29402 & ~n29408;
  assign n29423 = pi787 & ~n29422;
  assign n29424 = ~n29421 & ~n29423;
  assign n29425 = ~pi644 & n29424;
  assign n29426 = pi715 & ~n29425;
  assign n29427 = ~n29420 & n29426;
  assign n29428 = ~pi644 & n29182;
  assign n29429 = n17247 & ~n29182;
  assign n29430 = ~n17247 & n29226;
  assign n29431 = ~n29429 & ~n29430;
  assign n29432 = pi644 & n29431;
  assign n29433 = ~pi715 & ~n29432;
  assign n29434 = ~n29428 & n29433;
  assign n29435 = ~n29427 & ~n29434;
  assign n29436 = pi1160 & n29435;
  assign n29437 = ~pi644 & n29431;
  assign n29438 = pi715 & ~n29437;
  assign n29439 = pi644 & n29182;
  assign n29440 = n29438 & ~n29439;
  assign n29441 = pi644 & n29424;
  assign n29442 = ~pi644 & ~n29418;
  assign n29443 = ~pi715 & ~n29442;
  assign n29444 = ~n29441 & n29443;
  assign n29445 = ~n29440 & ~n29444;
  assign n29446 = ~pi1160 & n29445;
  assign n29447 = ~n29436 & ~n29446;
  assign n29448 = pi790 & n29447;
  assign n29449 = ~n29419 & ~n29448;
  assign n29450 = ~po1038 & n29449;
  assign n29451 = ~pi188 & po1038;
  assign n29452 = ~pi832 & ~n29451;
  assign n29453 = ~n29450 & n29452;
  assign n29454 = ~pi188 & ~n2934;
  assign n29455 = ~pi768 & n16510;
  assign n29456 = ~n29454 & ~n29455;
  assign n29457 = ~n17273 & ~n29456;
  assign n29458 = ~pi785 & ~n29457;
  assign n29459 = ~n17279 & ~n29456;
  assign n29460 = pi1155 & ~n29459;
  assign n29461 = ~n17282 & n29457;
  assign n29462 = ~pi1155 & ~n29461;
  assign n29463 = ~n29460 & ~n29462;
  assign n29464 = pi785 & ~n29463;
  assign n29465 = ~n29458 & ~n29464;
  assign n29466 = ~pi781 & ~n29465;
  assign n29467 = ~n17289 & n29465;
  assign n29468 = pi1154 & ~n29467;
  assign n29469 = ~n17292 & n29465;
  assign n29470 = ~pi1154 & ~n29469;
  assign n29471 = ~n29468 & ~n29470;
  assign n29472 = pi781 & ~n29471;
  assign n29473 = ~n29466 & ~n29472;
  assign n29474 = ~pi789 & ~n29473;
  assign n29475 = pi619 & n29473;
  assign n29476 = ~pi619 & n29454;
  assign n29477 = pi1159 & ~n29476;
  assign n29478 = ~n29475 & n29477;
  assign n29479 = ~pi619 & n29473;
  assign n29480 = pi619 & n29454;
  assign n29481 = ~pi1159 & ~n29480;
  assign n29482 = ~n29479 & n29481;
  assign n29483 = ~n29478 & ~n29482;
  assign n29484 = pi789 & ~n29483;
  assign n29485 = ~n29474 & ~n29484;
  assign n29486 = ~n17355 & n29485;
  assign n29487 = n17355 & n29454;
  assign n29488 = ~n29486 & ~n29487;
  assign n29489 = ~n16124 & ~n29488;
  assign n29490 = n16124 & n29454;
  assign n29491 = ~n29489 & ~n29490;
  assign n29492 = ~n19987 & n29491;
  assign n29493 = pi705 & n16742;
  assign n29494 = ~n29454 & ~n29493;
  assign n29495 = ~pi778 & n29494;
  assign n29496 = ~pi625 & n29493;
  assign n29497 = ~n29494 & ~n29496;
  assign n29498 = pi1153 & ~n29497;
  assign n29499 = ~pi1153 & ~n29454;
  assign n29500 = ~n29496 & n29499;
  assign n29501 = ~n29498 & ~n29500;
  assign n29502 = pi778 & ~n29501;
  assign n29503 = ~n29495 & ~n29502;
  assign n29504 = ~n17338 & n29503;
  assign n29505 = ~n17340 & n29504;
  assign n29506 = ~n17342 & n29505;
  assign n29507 = ~n17425 & n29506;
  assign n29508 = ~n17452 & n29507;
  assign n29509 = ~pi647 & n29508;
  assign n29510 = pi647 & n29454;
  assign n29511 = ~pi1157 & ~n29510;
  assign n29512 = ~n29509 & n29511;
  assign n29513 = ~pi647 & n29454;
  assign n29514 = pi647 & n29508;
  assign n29515 = pi1157 & ~n29514;
  assign n29516 = ~n29513 & n29515;
  assign n29517 = ~n29512 & ~n29516;
  assign n29518 = ~n17246 & ~n29517;
  assign n29519 = ~n29492 & ~n29518;
  assign n29520 = pi787 & ~n29519;
  assign n29521 = ~pi626 & ~n29485;
  assign n29522 = pi626 & ~n29454;
  assign n29523 = n17181 & ~n29522;
  assign n29524 = ~n29521 & n29523;
  assign n29525 = n17350 & n29506;
  assign n29526 = pi626 & ~n29485;
  assign n29527 = ~pi626 & ~n29454;
  assign n29528 = n17180 & ~n29527;
  assign n29529 = ~n29526 & n29528;
  assign n29530 = ~n29525 & ~n29529;
  assign n29531 = ~n29524 & n29530;
  assign n29532 = pi788 & ~n29531;
  assign n29533 = pi618 & n29504;
  assign n29534 = pi609 & n29503;
  assign n29535 = ~n16393 & ~n29494;
  assign n29536 = pi625 & n29535;
  assign n29537 = n29456 & ~n29535;
  assign n29538 = ~n29536 & ~n29537;
  assign n29539 = n29499 & ~n29538;
  assign n29540 = ~pi608 & ~n29498;
  assign n29541 = ~n29539 & n29540;
  assign n29542 = pi1153 & ~n29536;
  assign n29543 = n29456 & n29542;
  assign n29544 = ~n29500 & ~n29543;
  assign n29545 = pi608 & n29544;
  assign n29546 = ~n29541 & ~n29545;
  assign n29547 = pi778 & ~n29546;
  assign n29548 = ~pi778 & ~n29537;
  assign n29549 = ~n29547 & ~n29548;
  assign n29550 = ~pi609 & ~n29549;
  assign n29551 = ~pi1155 & ~n29550;
  assign n29552 = ~n29534 & n29551;
  assign n29553 = ~pi660 & ~n29460;
  assign n29554 = ~n29552 & n29553;
  assign n29555 = ~pi609 & n29503;
  assign n29556 = pi609 & ~n29549;
  assign n29557 = ~n29555 & ~n29556;
  assign n29558 = pi1155 & n29557;
  assign n29559 = ~n29462 & ~n29558;
  assign n29560 = pi660 & n29559;
  assign n29561 = ~n29554 & ~n29560;
  assign n29562 = pi785 & ~n29561;
  assign n29563 = ~pi785 & ~n29549;
  assign n29564 = ~n29562 & ~n29563;
  assign n29565 = ~pi618 & ~n29564;
  assign n29566 = ~pi1154 & ~n29565;
  assign n29567 = ~n29533 & n29566;
  assign n29568 = ~pi627 & ~n29468;
  assign n29569 = ~n29567 & n29568;
  assign n29570 = ~pi618 & n29504;
  assign n29571 = pi618 & ~n29564;
  assign n29572 = ~n29570 & ~n29571;
  assign n29573 = pi1154 & n29572;
  assign n29574 = ~n29470 & ~n29573;
  assign n29575 = pi627 & n29574;
  assign n29576 = ~n29569 & ~n29575;
  assign n29577 = pi781 & ~n29576;
  assign n29578 = ~pi781 & ~n29564;
  assign n29579 = ~n29577 & ~n29578;
  assign n29580 = ~pi619 & ~n29579;
  assign n29581 = pi619 & n29505;
  assign n29582 = ~pi1159 & ~n29581;
  assign n29583 = ~n29580 & n29582;
  assign n29584 = ~pi648 & ~n29583;
  assign n29585 = ~n29478 & n29584;
  assign n29586 = ~pi619 & n29505;
  assign n29587 = pi619 & ~n29579;
  assign n29588 = ~n29586 & ~n29587;
  assign n29589 = pi1159 & n29588;
  assign n29590 = ~n29482 & ~n29589;
  assign n29591 = pi648 & n29590;
  assign n29592 = ~n29585 & ~n29591;
  assign n29593 = pi789 & n29592;
  assign n29594 = ~pi789 & n29579;
  assign n29595 = n17356 & ~n29594;
  assign n29596 = ~n29593 & n29595;
  assign n29597 = ~n29532 & ~n29596;
  assign n29598 = n19788 & ~n29597;
  assign n29599 = n20275 & n29507;
  assign n29600 = n17449 & ~n29488;
  assign n29601 = ~pi629 & ~n29600;
  assign n29602 = ~n29599 & n29601;
  assign n29603 = n17448 & ~n29488;
  assign n29604 = n20281 & n29507;
  assign n29605 = pi629 & ~n29604;
  assign n29606 = ~n29603 & n29605;
  assign n29607 = ~n29602 & ~n29606;
  assign n29608 = pi792 & n29607;
  assign n29609 = n19637 & ~n29608;
  assign n29610 = ~n29598 & n29609;
  assign n29611 = ~n29520 & ~n29610;
  assign n29612 = pi644 & n29611;
  assign n29613 = ~pi787 & ~n29508;
  assign n29614 = pi787 & ~n29517;
  assign n29615 = ~n29613 & ~n29614;
  assign n29616 = ~pi644 & n29615;
  assign n29617 = pi715 & ~n29616;
  assign n29618 = ~n29612 & n29617;
  assign n29619 = ~n17247 & ~n29491;
  assign n29620 = n17247 & n29454;
  assign n29621 = ~n29619 & ~n29620;
  assign n29622 = pi644 & ~n29621;
  assign n29623 = ~pi644 & n29454;
  assign n29624 = ~pi715 & ~n29623;
  assign n29625 = ~n29622 & n29624;
  assign n29626 = pi1160 & ~n29625;
  assign n29627 = ~n29618 & n29626;
  assign n29628 = ~pi644 & ~n29621;
  assign n29629 = pi715 & ~n29628;
  assign n29630 = pi644 & n29454;
  assign n29631 = n29629 & ~n29630;
  assign n29632 = pi644 & n29615;
  assign n29633 = ~pi644 & n29611;
  assign n29634 = ~pi715 & ~n29633;
  assign n29635 = ~n29632 & n29634;
  assign n29636 = ~pi1160 & ~n29635;
  assign n29637 = ~n29631 & n29636;
  assign n29638 = ~n29627 & ~n29637;
  assign n29639 = pi790 & ~n29638;
  assign n29640 = ~pi790 & n29611;
  assign n29641 = pi832 & ~n29640;
  assign n29642 = ~n29639 & n29641;
  assign po345 = ~n29453 & ~n29642;
  assign n29644 = ~pi189 & ~n6274;
  assign n29645 = pi189 & ~n10020;
  assign n29646 = pi772 & n16447;
  assign n29647 = ~n21643 & ~n29646;
  assign n29648 = pi39 & ~n29647;
  assign n29649 = pi772 & n16380;
  assign n29650 = ~pi772 & n16201;
  assign n29651 = ~pi39 & ~n29650;
  assign n29652 = ~n29649 & n29651;
  assign n29653 = ~n29648 & ~n29652;
  assign n29654 = pi189 & ~n29653;
  assign n29655 = ~pi189 & pi772;
  assign n29656 = n16503 & n29655;
  assign n29657 = ~n29654 & ~n29656;
  assign n29658 = ~pi38 & ~n29657;
  assign n29659 = pi772 & n16393;
  assign n29660 = n16508 & ~n29659;
  assign n29661 = ~pi189 & ~n16508;
  assign n29662 = pi38 & ~n29661;
  assign n29663 = ~n29660 & n29662;
  assign n29664 = ~n29658 & ~n29663;
  assign n29665 = n10020 & ~n29664;
  assign n29666 = ~n29645 & ~n29665;
  assign n29667 = ~n16521 & ~n29666;
  assign n29668 = pi189 & ~n16527;
  assign n29669 = n16521 & n29668;
  assign n29670 = ~n29667 & ~n29669;
  assign n29671 = ~pi785 & ~n29670;
  assign n29672 = pi609 & n29670;
  assign n29673 = ~pi609 & ~n29668;
  assign n29674 = pi1155 & ~n29673;
  assign n29675 = ~n29672 & n29674;
  assign n29676 = ~pi609 & n29670;
  assign n29677 = pi609 & ~n29668;
  assign n29678 = ~pi1155 & ~n29677;
  assign n29679 = ~n29676 & n29678;
  assign n29680 = ~n29675 & ~n29679;
  assign n29681 = pi785 & ~n29680;
  assign n29682 = ~n29671 & ~n29681;
  assign n29683 = ~pi781 & ~n29682;
  assign n29684 = pi618 & n29682;
  assign n29685 = ~pi618 & ~n29668;
  assign n29686 = pi1154 & ~n29685;
  assign n29687 = ~n29684 & n29686;
  assign n29688 = ~pi618 & n29682;
  assign n29689 = pi618 & ~n29668;
  assign n29690 = ~pi1154 & ~n29689;
  assign n29691 = ~n29688 & n29690;
  assign n29692 = ~n29687 & ~n29691;
  assign n29693 = pi781 & ~n29692;
  assign n29694 = ~n29683 & ~n29693;
  assign n29695 = ~pi789 & ~n29694;
  assign n29696 = pi619 & n29694;
  assign n29697 = ~pi619 & ~n29668;
  assign n29698 = pi1159 & ~n29697;
  assign n29699 = ~n29696 & n29698;
  assign n29700 = ~pi619 & n29694;
  assign n29701 = pi619 & ~n29668;
  assign n29702 = ~pi1159 & ~n29701;
  assign n29703 = ~n29700 & n29702;
  assign n29704 = ~n29699 & ~n29703;
  assign n29705 = pi789 & ~n29704;
  assign n29706 = ~n29695 & ~n29705;
  assign n29707 = ~n17355 & ~n29706;
  assign n29708 = n17355 & n29668;
  assign n29709 = ~n29707 & ~n29708;
  assign n29710 = ~n16124 & ~n29709;
  assign n29711 = n16124 & n29668;
  assign n29712 = ~n29710 & ~n29711;
  assign n29713 = pi647 & n29712;
  assign n29714 = pi628 & n29709;
  assign n29715 = n16593 & ~n29668;
  assign n29716 = pi727 & n10020;
  assign n29717 = ~n29668 & ~n29716;
  assign n29718 = n19410 & ~n29661;
  assign n29719 = pi189 & ~n17592;
  assign n29720 = ~pi189 & ~n17589;
  assign n29721 = ~pi38 & ~n29720;
  assign n29722 = ~n29719 & n29721;
  assign n29723 = ~n29718 & ~n29722;
  assign n29724 = n29716 & n29723;
  assign n29725 = ~n29717 & ~n29724;
  assign n29726 = ~pi778 & n29725;
  assign n29727 = pi625 & ~n29725;
  assign n29728 = ~pi625 & ~n29668;
  assign n29729 = pi1153 & ~n29728;
  assign n29730 = ~n29727 & n29729;
  assign n29731 = ~pi625 & ~n29725;
  assign n29732 = pi625 & ~n29668;
  assign n29733 = ~pi1153 & ~n29732;
  assign n29734 = ~n29731 & n29733;
  assign n29735 = ~n29730 & ~n29734;
  assign n29736 = pi778 & ~n29735;
  assign n29737 = ~n29726 & ~n29736;
  assign n29738 = ~n16593 & n29737;
  assign n29739 = ~n29715 & ~n29738;
  assign n29740 = ~n16589 & n29739;
  assign n29741 = n16589 & n29668;
  assign n29742 = ~n29740 & ~n29741;
  assign n29743 = pi619 & n29742;
  assign n29744 = pi618 & ~n29739;
  assign n29745 = pi609 & n29737;
  assign n29746 = pi625 & n29666;
  assign n29747 = ~n29665 & ~n29716;
  assign n29748 = pi189 & ~n17061;
  assign n29749 = ~pi189 & ~n17058;
  assign n29750 = ~pi772 & ~n29749;
  assign n29751 = ~n29748 & n29750;
  assign n29752 = ~pi189 & n17065;
  assign n29753 = pi189 & n17067;
  assign n29754 = ~n29752 & ~n29753;
  assign n29755 = pi772 & n29754;
  assign n29756 = ~pi39 & ~n29755;
  assign n29757 = ~n29751 & n29756;
  assign n29758 = ~pi189 & ~n16998;
  assign n29759 = pi772 & ~n29758;
  assign n29760 = pi189 & n17051;
  assign n29761 = n29759 & ~n29760;
  assign n29762 = ~pi189 & ~n16935;
  assign n29763 = pi189 & ~n16853;
  assign n29764 = ~pi772 & ~n29763;
  assign n29765 = ~n29762 & n29764;
  assign n29766 = pi39 & ~n29765;
  assign n29767 = ~n29761 & n29766;
  assign n29768 = ~pi38 & ~n29767;
  assign n29769 = ~n29757 & n29768;
  assign n29770 = pi727 & ~n29769;
  assign n29771 = ~n18932 & n29770;
  assign n29772 = ~n29663 & n29771;
  assign n29773 = ~n29747 & ~n29772;
  assign n29774 = ~n29645 & ~n29773;
  assign n29775 = ~pi625 & n29774;
  assign n29776 = ~pi1153 & ~n29775;
  assign n29777 = ~n29746 & n29776;
  assign n29778 = ~pi608 & ~n29730;
  assign n29779 = ~n29777 & n29778;
  assign n29780 = ~pi625 & n29666;
  assign n29781 = pi625 & n29774;
  assign n29782 = ~n29780 & ~n29781;
  assign n29783 = pi1153 & n29782;
  assign n29784 = ~n29734 & ~n29783;
  assign n29785 = pi608 & n29784;
  assign n29786 = ~n29779 & ~n29785;
  assign n29787 = pi778 & ~n29786;
  assign n29788 = ~pi778 & n29774;
  assign n29789 = ~n29787 & ~n29788;
  assign n29790 = ~pi609 & ~n29789;
  assign n29791 = ~pi1155 & ~n29790;
  assign n29792 = ~n29745 & n29791;
  assign n29793 = ~pi660 & ~n29675;
  assign n29794 = ~n29792 & n29793;
  assign n29795 = ~pi609 & n29737;
  assign n29796 = pi609 & ~n29789;
  assign n29797 = ~n29795 & ~n29796;
  assign n29798 = pi1155 & n29797;
  assign n29799 = ~n29679 & ~n29798;
  assign n29800 = pi660 & n29799;
  assign n29801 = ~n29794 & ~n29800;
  assign n29802 = pi785 & ~n29801;
  assign n29803 = ~pi785 & ~n29789;
  assign n29804 = ~n29802 & ~n29803;
  assign n29805 = ~pi618 & ~n29804;
  assign n29806 = ~pi1154 & ~n29805;
  assign n29807 = ~n29744 & n29806;
  assign n29808 = ~pi627 & ~n29687;
  assign n29809 = ~n29807 & n29808;
  assign n29810 = ~pi618 & ~n29739;
  assign n29811 = pi618 & ~n29804;
  assign n29812 = ~n29810 & ~n29811;
  assign n29813 = pi1154 & n29812;
  assign n29814 = ~n29691 & ~n29813;
  assign n29815 = pi627 & n29814;
  assign n29816 = ~n29809 & ~n29815;
  assign n29817 = pi781 & ~n29816;
  assign n29818 = ~pi781 & ~n29804;
  assign n29819 = ~n29817 & ~n29818;
  assign n29820 = ~pi619 & ~n29819;
  assign n29821 = ~pi1159 & ~n29820;
  assign n29822 = ~n29743 & n29821;
  assign n29823 = ~pi648 & ~n29699;
  assign n29824 = ~n29822 & n29823;
  assign n29825 = ~pi619 & n29742;
  assign n29826 = pi619 & ~n29819;
  assign n29827 = ~n29825 & ~n29826;
  assign n29828 = pi1159 & n29827;
  assign n29829 = ~n29703 & ~n29828;
  assign n29830 = pi648 & n29829;
  assign n29831 = ~n29824 & ~n29830;
  assign n29832 = pi789 & ~n29831;
  assign n29833 = ~pi789 & ~n29819;
  assign n29834 = ~n29832 & ~n29833;
  assign n29835 = ~pi788 & n29834;
  assign n29836 = pi626 & n29834;
  assign n29837 = n17159 & ~n29668;
  assign n29838 = ~n17159 & n29742;
  assign n29839 = ~n29837 & ~n29838;
  assign n29840 = ~pi626 & n29839;
  assign n29841 = pi641 & ~n29840;
  assign n29842 = ~n29836 & n29841;
  assign n29843 = pi626 & ~n29706;
  assign n29844 = ~pi626 & n29668;
  assign n29845 = ~pi641 & ~n29844;
  assign n29846 = ~n29843 & n29845;
  assign n29847 = pi1158 & ~n29846;
  assign n29848 = ~n29842 & n29847;
  assign n29849 = ~pi626 & ~n29706;
  assign n29850 = pi641 & ~n29849;
  assign n29851 = pi626 & n29668;
  assign n29852 = n29850 & ~n29851;
  assign n29853 = pi626 & n29839;
  assign n29854 = ~pi626 & n29834;
  assign n29855 = ~pi641 & ~n29854;
  assign n29856 = ~n29853 & n29855;
  assign n29857 = ~pi1158 & ~n29856;
  assign n29858 = ~n29852 & n29857;
  assign n29859 = ~n29848 & ~n29858;
  assign n29860 = pi788 & ~n29859;
  assign n29861 = ~n29835 & ~n29860;
  assign n29862 = ~pi628 & n29861;
  assign n29863 = ~pi1156 & ~n29862;
  assign n29864 = ~n29714 & n29863;
  assign n29865 = ~n17183 & n29839;
  assign n29866 = n17183 & n29668;
  assign n29867 = ~n29865 & ~n29866;
  assign n29868 = pi628 & n29867;
  assign n29869 = ~pi628 & ~n29668;
  assign n29870 = pi1156 & ~n29869;
  assign n29871 = ~n29868 & n29870;
  assign n29872 = ~pi629 & ~n29871;
  assign n29873 = ~n29864 & n29872;
  assign n29874 = ~pi628 & n29867;
  assign n29875 = pi628 & ~n29668;
  assign n29876 = ~pi1156 & ~n29875;
  assign n29877 = ~n29874 & n29876;
  assign n29878 = ~pi628 & n29709;
  assign n29879 = pi628 & n29861;
  assign n29880 = ~n29878 & ~n29879;
  assign n29881 = pi1156 & n29880;
  assign n29882 = ~n29877 & ~n29881;
  assign n29883 = pi629 & n29882;
  assign n29884 = ~n29873 & ~n29883;
  assign n29885 = pi792 & ~n29884;
  assign n29886 = ~pi792 & n29861;
  assign n29887 = ~n29885 & ~n29886;
  assign n29888 = ~pi647 & ~n29887;
  assign n29889 = ~pi1157 & ~n29888;
  assign n29890 = ~n29713 & n29889;
  assign n29891 = ~pi792 & ~n29867;
  assign n29892 = ~n29871 & ~n29877;
  assign n29893 = pi792 & ~n29892;
  assign n29894 = ~n29891 & ~n29893;
  assign n29895 = pi647 & n29894;
  assign n29896 = ~pi647 & ~n29668;
  assign n29897 = pi1157 & ~n29896;
  assign n29898 = ~n29895 & n29897;
  assign n29899 = ~pi630 & ~n29898;
  assign n29900 = ~n29890 & n29899;
  assign n29901 = ~pi647 & n29894;
  assign n29902 = pi647 & ~n29668;
  assign n29903 = ~pi1157 & ~n29902;
  assign n29904 = ~n29901 & n29903;
  assign n29905 = ~pi647 & n29712;
  assign n29906 = pi647 & ~n29887;
  assign n29907 = ~n29905 & ~n29906;
  assign n29908 = pi1157 & n29907;
  assign n29909 = ~n29904 & ~n29908;
  assign n29910 = pi630 & n29909;
  assign n29911 = ~n29900 & ~n29910;
  assign n29912 = pi787 & ~n29911;
  assign n29913 = ~pi787 & ~n29887;
  assign n29914 = ~n29912 & ~n29913;
  assign n29915 = ~pi790 & n29914;
  assign n29916 = pi644 & ~n29914;
  assign n29917 = ~pi787 & ~n29894;
  assign n29918 = ~n29898 & ~n29904;
  assign n29919 = pi787 & ~n29918;
  assign n29920 = ~n29917 & ~n29919;
  assign n29921 = ~pi644 & n29920;
  assign n29922 = pi715 & ~n29921;
  assign n29923 = ~n29916 & n29922;
  assign n29924 = ~pi644 & ~n29668;
  assign n29925 = n17247 & ~n29668;
  assign n29926 = ~n17247 & n29712;
  assign n29927 = ~n29925 & ~n29926;
  assign n29928 = pi644 & ~n29927;
  assign n29929 = ~pi715 & ~n29928;
  assign n29930 = ~n29924 & n29929;
  assign n29931 = ~n29923 & ~n29930;
  assign n29932 = pi1160 & n29931;
  assign n29933 = pi644 & ~n29668;
  assign n29934 = ~pi644 & ~n29927;
  assign n29935 = pi715 & ~n29934;
  assign n29936 = ~n29933 & n29935;
  assign n29937 = pi644 & n29920;
  assign n29938 = ~pi644 & ~n29914;
  assign n29939 = ~pi715 & ~n29938;
  assign n29940 = ~n29937 & n29939;
  assign n29941 = ~n29936 & ~n29940;
  assign n29942 = ~pi1160 & n29941;
  assign n29943 = ~n29932 & ~n29942;
  assign n29944 = pi790 & n29943;
  assign n29945 = ~n29915 & ~n29944;
  assign n29946 = n6274 & n29945;
  assign n29947 = ~pi57 & ~n29946;
  assign n29948 = ~n29644 & n29947;
  assign n29949 = pi57 & pi189;
  assign n29950 = ~pi832 & ~n29949;
  assign n29951 = ~n29948 & n29950;
  assign n29952 = pi189 & ~n2934;
  assign n29953 = pi727 & n16742;
  assign n29954 = ~n29952 & ~n29953;
  assign n29955 = ~pi778 & n29954;
  assign n29956 = pi625 & n29953;
  assign n29957 = ~n29954 & ~n29956;
  assign n29958 = ~pi1153 & ~n29957;
  assign n29959 = pi1153 & ~n29952;
  assign n29960 = ~n29956 & n29959;
  assign n29961 = ~n29958 & ~n29960;
  assign n29962 = pi778 & ~n29961;
  assign n29963 = ~n29955 & ~n29962;
  assign n29964 = n18715 & n29963;
  assign n29965 = ~n17159 & n29964;
  assign n29966 = ~n29952 & ~n29965;
  assign n29967 = n17345 & ~n29966;
  assign n29968 = pi772 & n16510;
  assign n29969 = ~n19656 & n29968;
  assign n29970 = ~n19662 & n29969;
  assign n29971 = n19668 & n29970;
  assign n29972 = pi626 & n29971;
  assign n29973 = ~n29952 & ~n29972;
  assign n29974 = pi1158 & ~n29973;
  assign n29975 = ~pi641 & ~n29974;
  assign n29976 = ~n29967 & n29975;
  assign n29977 = ~pi626 & n29971;
  assign n29978 = ~n29952 & ~n29977;
  assign n29979 = ~pi1158 & ~n29978;
  assign n29980 = n17344 & ~n29966;
  assign n29981 = pi641 & ~n29980;
  assign n29982 = ~n29979 & n29981;
  assign n29983 = ~n29976 & ~n29982;
  assign n29984 = pi788 & n29983;
  assign n29985 = pi609 & n29963;
  assign n29986 = ~n29952 & ~n29968;
  assign n29987 = ~n16393 & n29953;
  assign n29988 = n29986 & ~n29987;
  assign n29989 = pi625 & n29987;
  assign n29990 = ~n29988 & ~n29989;
  assign n29991 = ~pi1153 & ~n29990;
  assign n29992 = ~pi608 & ~n29960;
  assign n29993 = ~n29991 & n29992;
  assign n29994 = pi1153 & ~n29989;
  assign n29995 = n29986 & n29994;
  assign n29996 = ~n29958 & ~n29995;
  assign n29997 = pi608 & n29996;
  assign n29998 = ~n29993 & ~n29997;
  assign n29999 = pi778 & ~n29998;
  assign n30000 = ~pi778 & ~n29988;
  assign n30001 = ~n29999 & ~n30000;
  assign n30002 = ~pi609 & ~n30001;
  assign n30003 = ~pi1155 & ~n30002;
  assign n30004 = ~n29985 & n30003;
  assign n30005 = ~n17279 & ~n29986;
  assign n30006 = pi1155 & ~n30005;
  assign n30007 = ~pi660 & ~n30006;
  assign n30008 = ~n30004 & n30007;
  assign n30009 = ~pi609 & n29963;
  assign n30010 = pi609 & ~n30001;
  assign n30011 = ~n30009 & ~n30010;
  assign n30012 = pi1155 & n30011;
  assign n30013 = ~pi1155 & ~n29952;
  assign n30014 = n16537 & n29968;
  assign n30015 = n30013 & ~n30014;
  assign n30016 = pi660 & ~n30015;
  assign n30017 = ~n30012 & n30016;
  assign n30018 = ~n30008 & ~n30017;
  assign n30019 = pi785 & ~n30018;
  assign n30020 = ~pi785 & ~n30001;
  assign n30021 = ~n30019 & ~n30020;
  assign n30022 = ~pi781 & ~n30021;
  assign n30023 = ~n17338 & n29963;
  assign n30024 = ~pi618 & n30023;
  assign n30025 = pi618 & ~n30021;
  assign n30026 = ~n30024 & ~n30025;
  assign n30027 = pi1154 & n30026;
  assign n30028 = n19753 & n29969;
  assign n30029 = ~pi1154 & ~n29952;
  assign n30030 = ~n30028 & n30029;
  assign n30031 = pi627 & ~n30030;
  assign n30032 = ~n30027 & n30031;
  assign n30033 = pi618 & n30023;
  assign n30034 = ~pi618 & ~n30021;
  assign n30035 = ~pi1154 & ~n30034;
  assign n30036 = ~n30033 & n30035;
  assign n30037 = ~pi627 & ~n30036;
  assign n30038 = n19744 & n29969;
  assign n30039 = ~n29952 & ~n30038;
  assign n30040 = pi1154 & n30039;
  assign n30041 = n30037 & ~n30040;
  assign n30042 = ~n30032 & ~n30041;
  assign n30043 = pi781 & ~n30042;
  assign n30044 = n22991 & ~n30043;
  assign n30045 = ~n30022 & n30044;
  assign n30046 = ~n22996 & ~n29964;
  assign n30047 = n19776 & n29970;
  assign n30048 = n17156 & ~n30047;
  assign n30049 = n19766 & n29970;
  assign n30050 = n17157 & ~n30049;
  assign n30051 = ~n30048 & ~n30050;
  assign n30052 = ~n30046 & n30051;
  assign n30053 = pi789 & ~n29952;
  assign n30054 = ~n30052 & n30053;
  assign n30055 = n17356 & ~n30054;
  assign n30056 = ~n30045 & n30055;
  assign n30057 = ~n29984 & ~n30056;
  assign n30058 = n19788 & n30057;
  assign n30059 = ~n17355 & n29971;
  assign n30060 = ~pi629 & n30059;
  assign n30061 = pi628 & ~n30060;
  assign n30062 = n18717 & n29963;
  assign n30063 = pi629 & ~n30062;
  assign n30064 = ~n30061 & ~n30063;
  assign n30065 = ~pi1156 & ~n30064;
  assign n30066 = pi628 & n30062;
  assign n30067 = ~pi628 & ~n30059;
  assign n30068 = pi629 & ~n30067;
  assign n30069 = pi1156 & ~n30068;
  assign n30070 = ~n30066 & n30069;
  assign n30071 = ~n30065 & ~n30070;
  assign n30072 = ~n29952 & ~n30071;
  assign n30073 = pi792 & n30072;
  assign n30074 = ~n30058 & ~n30073;
  assign n30075 = n19637 & ~n30074;
  assign n30076 = ~n16124 & n30059;
  assign n30077 = ~pi630 & n30076;
  assign n30078 = pi647 & ~n30077;
  assign n30079 = ~n18744 & n30062;
  assign n30080 = pi630 & ~n30079;
  assign n30081 = ~n30078 & ~n30080;
  assign n30082 = ~pi1157 & ~n30081;
  assign n30083 = ~pi630 & ~n30079;
  assign n30084 = pi647 & ~n30083;
  assign n30085 = pi630 & n30076;
  assign n30086 = pi1157 & ~n30085;
  assign n30087 = ~n30084 & n30086;
  assign n30088 = ~n30082 & ~n30087;
  assign n30089 = ~n29952 & ~n30088;
  assign n30090 = pi787 & n30089;
  assign n30091 = ~n30075 & ~n30090;
  assign n30092 = pi644 & n30091;
  assign n30093 = ~n18767 & n30079;
  assign n30094 = ~n29952 & ~n30093;
  assign n30095 = ~pi644 & ~n30094;
  assign n30096 = pi715 & ~n30095;
  assign n30097 = ~n30092 & n30096;
  assign n30098 = ~n17355 & n23049;
  assign n30099 = n29971 & n30098;
  assign n30100 = pi644 & n30099;
  assign n30101 = ~pi715 & ~n29952;
  assign n30102 = ~n30100 & n30101;
  assign n30103 = pi1160 & ~n30102;
  assign n30104 = ~n30097 & n30103;
  assign n30105 = pi644 & ~n30094;
  assign n30106 = ~pi644 & n30091;
  assign n30107 = ~pi715 & ~n30106;
  assign n30108 = ~n30105 & n30107;
  assign n30109 = ~pi1160 & ~n30108;
  assign n30110 = ~pi644 & n30099;
  assign n30111 = ~n29952 & ~n30110;
  assign n30112 = pi715 & n30111;
  assign n30113 = n30109 & ~n30112;
  assign n30114 = ~n30104 & ~n30113;
  assign n30115 = pi790 & ~n30114;
  assign n30116 = ~pi790 & n30091;
  assign n30117 = pi832 & ~n30116;
  assign n30118 = ~n30115 & n30117;
  assign po346 = ~n29951 & ~n30118;
  assign n30120 = ~pi190 & ~n2934;
  assign n30121 = pi763 & n16510;
  assign n30122 = ~n30120 & ~n30121;
  assign n30123 = ~n17273 & ~n30122;
  assign n30124 = ~pi785 & ~n30123;
  assign n30125 = n16537 & n30121;
  assign n30126 = n30123 & ~n30125;
  assign n30127 = pi1155 & ~n30126;
  assign n30128 = ~pi1155 & ~n30120;
  assign n30129 = ~n30125 & n30128;
  assign n30130 = ~n30127 & ~n30129;
  assign n30131 = pi785 & ~n30130;
  assign n30132 = ~n30124 & ~n30131;
  assign n30133 = ~pi781 & ~n30132;
  assign n30134 = ~n17289 & n30132;
  assign n30135 = pi1154 & ~n30134;
  assign n30136 = ~n17292 & n30132;
  assign n30137 = ~pi1154 & ~n30136;
  assign n30138 = ~n30135 & ~n30137;
  assign n30139 = pi781 & ~n30138;
  assign n30140 = ~n30133 & ~n30139;
  assign n30141 = ~pi789 & ~n30140;
  assign n30142 = ~n22423 & n30140;
  assign n30143 = pi1159 & ~n30142;
  assign n30144 = ~n22426 & n30140;
  assign n30145 = ~pi1159 & ~n30144;
  assign n30146 = ~n30143 & ~n30145;
  assign n30147 = pi789 & ~n30146;
  assign n30148 = ~n30141 & ~n30147;
  assign n30149 = ~n17355 & n30148;
  assign n30150 = n17355 & n30120;
  assign n30151 = ~n30149 & ~n30150;
  assign n30152 = ~n16124 & ~n30151;
  assign n30153 = n16124 & n30120;
  assign n30154 = ~n30152 & ~n30153;
  assign n30155 = ~n19987 & n30154;
  assign n30156 = pi699 & n16742;
  assign n30157 = ~n30120 & ~n30156;
  assign n30158 = ~pi778 & ~n30157;
  assign n30159 = ~pi625 & n30156;
  assign n30160 = ~n30157 & ~n30159;
  assign n30161 = pi1153 & ~n30160;
  assign n30162 = ~pi1153 & ~n30120;
  assign n30163 = ~n30159 & n30162;
  assign n30164 = ~n30161 & ~n30163;
  assign n30165 = pi778 & n30164;
  assign n30166 = ~n30158 & ~n30165;
  assign n30167 = ~n17338 & ~n30166;
  assign n30168 = ~n17340 & n30167;
  assign n30169 = ~n17342 & n30168;
  assign n30170 = ~n17425 & n30169;
  assign n30171 = ~n17452 & n30170;
  assign n30172 = ~pi647 & n30171;
  assign n30173 = pi647 & n30120;
  assign n30174 = ~pi1157 & ~n30173;
  assign n30175 = ~n30172 & n30174;
  assign n30176 = ~pi647 & n30120;
  assign n30177 = pi647 & n30171;
  assign n30178 = pi1157 & ~n30177;
  assign n30179 = ~n30176 & n30178;
  assign n30180 = ~n30175 & ~n30179;
  assign n30181 = ~n17246 & ~n30180;
  assign n30182 = ~n30155 & ~n30181;
  assign n30183 = pi787 & ~n30182;
  assign n30184 = ~pi626 & ~n30148;
  assign n30185 = pi626 & ~n30120;
  assign n30186 = n17181 & ~n30185;
  assign n30187 = ~n30184 & n30186;
  assign n30188 = n17350 & n30169;
  assign n30189 = pi626 & ~n30148;
  assign n30190 = ~pi626 & ~n30120;
  assign n30191 = n17180 & ~n30190;
  assign n30192 = ~n30189 & n30191;
  assign n30193 = ~n30188 & ~n30192;
  assign n30194 = ~n30187 & n30193;
  assign n30195 = pi788 & ~n30194;
  assign n30196 = pi618 & n30167;
  assign n30197 = pi609 & ~n30166;
  assign n30198 = ~n16393 & ~n30157;
  assign n30199 = pi625 & n30198;
  assign n30200 = n30122 & ~n30198;
  assign n30201 = ~n30199 & ~n30200;
  assign n30202 = n30162 & ~n30201;
  assign n30203 = ~pi608 & ~n30161;
  assign n30204 = ~n30202 & n30203;
  assign n30205 = pi1153 & ~n30199;
  assign n30206 = n30122 & n30205;
  assign n30207 = ~n30163 & ~n30206;
  assign n30208 = pi608 & n30207;
  assign n30209 = ~n30204 & ~n30208;
  assign n30210 = pi778 & ~n30209;
  assign n30211 = ~pi778 & ~n30200;
  assign n30212 = ~n30210 & ~n30211;
  assign n30213 = ~pi609 & ~n30212;
  assign n30214 = ~pi1155 & ~n30213;
  assign n30215 = ~n30197 & n30214;
  assign n30216 = ~pi660 & ~n30127;
  assign n30217 = ~n30215 & n30216;
  assign n30218 = ~pi609 & ~n30166;
  assign n30219 = pi609 & ~n30212;
  assign n30220 = ~n30218 & ~n30219;
  assign n30221 = pi1155 & n30220;
  assign n30222 = ~n30129 & ~n30221;
  assign n30223 = pi660 & n30222;
  assign n30224 = ~n30217 & ~n30223;
  assign n30225 = pi785 & ~n30224;
  assign n30226 = ~pi785 & ~n30212;
  assign n30227 = ~n30225 & ~n30226;
  assign n30228 = ~pi618 & ~n30227;
  assign n30229 = ~pi1154 & ~n30228;
  assign n30230 = ~n30196 & n30229;
  assign n30231 = ~pi627 & ~n30135;
  assign n30232 = ~n30230 & n30231;
  assign n30233 = ~pi618 & n30167;
  assign n30234 = pi618 & ~n30227;
  assign n30235 = ~n30233 & ~n30234;
  assign n30236 = pi1154 & n30235;
  assign n30237 = ~n30137 & ~n30236;
  assign n30238 = pi627 & n30237;
  assign n30239 = ~n30232 & ~n30238;
  assign n30240 = pi781 & ~n30239;
  assign n30241 = ~pi781 & ~n30227;
  assign n30242 = ~n30240 & ~n30241;
  assign n30243 = ~pi619 & ~n30242;
  assign n30244 = pi619 & n30168;
  assign n30245 = ~pi1159 & ~n30244;
  assign n30246 = ~n30243 & n30245;
  assign n30247 = ~pi648 & ~n30246;
  assign n30248 = ~n30143 & n30247;
  assign n30249 = ~pi619 & n30168;
  assign n30250 = pi619 & ~n30242;
  assign n30251 = ~n30249 & ~n30250;
  assign n30252 = pi1159 & n30251;
  assign n30253 = ~n30145 & ~n30252;
  assign n30254 = pi648 & n30253;
  assign n30255 = ~n30248 & ~n30254;
  assign n30256 = pi789 & n30255;
  assign n30257 = ~pi789 & n30242;
  assign n30258 = n17356 & ~n30257;
  assign n30259 = ~n30256 & n30258;
  assign n30260 = ~n30195 & ~n30259;
  assign n30261 = n19788 & ~n30260;
  assign n30262 = n20275 & n30170;
  assign n30263 = n17449 & ~n30151;
  assign n30264 = ~pi629 & ~n30263;
  assign n30265 = ~n30262 & n30264;
  assign n30266 = n17448 & ~n30151;
  assign n30267 = n20281 & n30170;
  assign n30268 = pi629 & ~n30267;
  assign n30269 = ~n30266 & n30268;
  assign n30270 = ~n30265 & ~n30269;
  assign n30271 = pi792 & n30270;
  assign n30272 = n19637 & ~n30271;
  assign n30273 = ~n30261 & n30272;
  assign n30274 = ~n30183 & ~n30273;
  assign n30275 = pi644 & n30274;
  assign n30276 = ~pi787 & ~n30171;
  assign n30277 = pi787 & ~n30180;
  assign n30278 = ~n30276 & ~n30277;
  assign n30279 = ~pi644 & n30278;
  assign n30280 = pi715 & ~n30279;
  assign n30281 = ~n30275 & n30280;
  assign n30282 = ~n17247 & ~n30154;
  assign n30283 = n17247 & n30120;
  assign n30284 = ~n30282 & ~n30283;
  assign n30285 = pi644 & ~n30284;
  assign n30286 = ~pi644 & n30120;
  assign n30287 = ~pi715 & ~n30286;
  assign n30288 = ~n30285 & n30287;
  assign n30289 = pi1160 & ~n30288;
  assign n30290 = ~n30281 & n30289;
  assign n30291 = ~pi644 & ~n30284;
  assign n30292 = pi715 & ~n30291;
  assign n30293 = pi644 & n30120;
  assign n30294 = n30292 & ~n30293;
  assign n30295 = pi644 & n30278;
  assign n30296 = ~pi644 & n30274;
  assign n30297 = ~pi715 & ~n30296;
  assign n30298 = ~n30295 & n30297;
  assign n30299 = ~pi1160 & ~n30298;
  assign n30300 = ~n30294 & n30299;
  assign n30301 = ~n30290 & ~n30300;
  assign n30302 = pi790 & ~n30301;
  assign n30303 = ~pi790 & n30274;
  assign n30304 = pi832 & ~n30303;
  assign n30305 = ~n30302 & n30304;
  assign n30306 = ~pi190 & ~n16527;
  assign n30307 = n17451 & ~n30306;
  assign n30308 = n17159 & ~n30306;
  assign n30309 = n16593 & ~n30306;
  assign n30310 = pi190 & ~n10020;
  assign n30311 = pi190 & n17589;
  assign n30312 = ~pi190 & n17592;
  assign n30313 = ~pi38 & ~n30312;
  assign n30314 = ~n30311 & n30313;
  assign n30315 = ~pi190 & ~n16508;
  assign n30316 = n16744 & ~n30315;
  assign n30317 = pi699 & ~n30316;
  assign n30318 = ~n30314 & n30317;
  assign n30319 = ~pi190 & ~pi699;
  assign n30320 = ~n16526 & n30319;
  assign n30321 = ~n30318 & ~n30320;
  assign n30322 = n10020 & n30321;
  assign n30323 = ~n30310 & ~n30322;
  assign n30324 = ~pi778 & ~n30323;
  assign n30325 = pi625 & n30323;
  assign n30326 = pi1153 & ~n30325;
  assign n30327 = ~pi625 & n30306;
  assign n30328 = n30326 & ~n30327;
  assign n30329 = ~pi625 & n30323;
  assign n30330 = ~pi1153 & ~n30329;
  assign n30331 = pi625 & n30306;
  assign n30332 = n30330 & ~n30331;
  assign n30333 = ~n30328 & ~n30332;
  assign n30334 = pi778 & ~n30333;
  assign n30335 = ~n30324 & ~n30334;
  assign n30336 = ~n16593 & ~n30335;
  assign n30337 = ~n30309 & ~n30336;
  assign n30338 = ~n16589 & n30337;
  assign n30339 = n16589 & n30306;
  assign n30340 = ~n30338 & ~n30339;
  assign n30341 = ~n17159 & n30340;
  assign n30342 = ~n30308 & ~n30341;
  assign n30343 = ~n17183 & n30342;
  assign n30344 = n17183 & n30306;
  assign n30345 = ~n30343 & ~n30344;
  assign n30346 = ~n17451 & n30345;
  assign n30347 = ~n30307 & ~n30346;
  assign n30348 = ~n18767 & n30347;
  assign n30349 = n18767 & n30306;
  assign n30350 = ~n30348 & ~n30349;
  assign n30351 = ~pi644 & ~n30350;
  assign n30352 = pi715 & ~n30351;
  assign n30353 = n17247 & ~n30306;
  assign n30354 = ~pi763 & n16355;
  assign n30355 = pi190 & n16501;
  assign n30356 = ~n30354 & ~n30355;
  assign n30357 = pi39 & ~n30356;
  assign n30358 = pi763 & ~n16461;
  assign n30359 = pi190 & ~n30358;
  assign n30360 = ~n21734 & ~n30359;
  assign n30361 = ~pi190 & n16449;
  assign n30362 = pi763 & n30361;
  assign n30363 = n30360 & ~n30362;
  assign n30364 = ~n30357 & n30363;
  assign n30365 = ~pi38 & ~n30364;
  assign n30366 = pi763 & n16511;
  assign n30367 = ~n30315 & ~n30366;
  assign n30368 = pi38 & n30367;
  assign n30369 = ~n30365 & ~n30368;
  assign n30370 = n10020 & ~n30369;
  assign n30371 = ~n30310 & ~n30370;
  assign n30372 = ~n16521 & ~n30371;
  assign n30373 = n16521 & ~n30306;
  assign n30374 = ~n30372 & ~n30373;
  assign n30375 = ~pi785 & ~n30374;
  assign n30376 = ~n16532 & ~n30306;
  assign n30377 = pi609 & n30372;
  assign n30378 = ~n30376 & ~n30377;
  assign n30379 = pi1155 & ~n30378;
  assign n30380 = ~n16537 & ~n30306;
  assign n30381 = ~pi609 & n30372;
  assign n30382 = ~n30380 & ~n30381;
  assign n30383 = ~pi1155 & ~n30382;
  assign n30384 = ~n30379 & ~n30383;
  assign n30385 = pi785 & ~n30384;
  assign n30386 = ~n30375 & ~n30385;
  assign n30387 = ~pi781 & ~n30386;
  assign n30388 = pi618 & n30386;
  assign n30389 = ~pi618 & n30306;
  assign n30390 = pi1154 & ~n30389;
  assign n30391 = ~n30388 & n30390;
  assign n30392 = ~pi618 & n30386;
  assign n30393 = pi618 & n30306;
  assign n30394 = ~pi1154 & ~n30393;
  assign n30395 = ~n30392 & n30394;
  assign n30396 = ~n30391 & ~n30395;
  assign n30397 = pi781 & ~n30396;
  assign n30398 = ~n30387 & ~n30397;
  assign n30399 = ~pi789 & ~n30398;
  assign n30400 = pi619 & n30398;
  assign n30401 = ~pi619 & n30306;
  assign n30402 = pi1159 & ~n30401;
  assign n30403 = ~n30400 & n30402;
  assign n30404 = ~pi619 & n30398;
  assign n30405 = pi619 & n30306;
  assign n30406 = ~pi1159 & ~n30405;
  assign n30407 = ~n30404 & n30406;
  assign n30408 = ~n30403 & ~n30407;
  assign n30409 = pi789 & ~n30408;
  assign n30410 = ~n30399 & ~n30409;
  assign n30411 = ~n17355 & n30410;
  assign n30412 = n17355 & n30306;
  assign n30413 = ~n30411 & ~n30412;
  assign n30414 = ~n16124 & ~n30413;
  assign n30415 = n16124 & n30306;
  assign n30416 = ~n30414 & ~n30415;
  assign n30417 = ~n17247 & n30416;
  assign n30418 = ~n30353 & ~n30417;
  assign n30419 = pi644 & n30418;
  assign n30420 = ~pi644 & n30306;
  assign n30421 = ~pi715 & ~n30420;
  assign n30422 = ~n30419 & n30421;
  assign n30423 = pi1160 & ~n30422;
  assign n30424 = ~n30352 & n30423;
  assign n30425 = pi644 & ~n30350;
  assign n30426 = ~pi715 & ~n30425;
  assign n30427 = ~pi644 & n30418;
  assign n30428 = pi644 & n30306;
  assign n30429 = ~n30427 & ~n30428;
  assign n30430 = pi715 & n30429;
  assign n30431 = ~pi1160 & ~n30430;
  assign n30432 = ~n30426 & n30431;
  assign n30433 = ~n30424 & ~n30432;
  assign n30434 = pi790 & ~n30433;
  assign n30435 = ~n19999 & n30413;
  assign n30436 = pi628 & ~n30345;
  assign n30437 = n16121 & ~n30436;
  assign n30438 = ~pi628 & n30306;
  assign n30439 = n30437 & ~n30438;
  assign n30440 = ~pi628 & ~n30345;
  assign n30441 = pi628 & n30306;
  assign n30442 = n16122 & ~n30441;
  assign n30443 = ~n30440 & n30442;
  assign n30444 = ~n30439 & ~n30443;
  assign n30445 = ~n30435 & n30444;
  assign n30446 = pi792 & ~n30445;
  assign n30447 = pi618 & n30337;
  assign n30448 = pi609 & n30335;
  assign n30449 = pi625 & n30371;
  assign n30450 = ~pi699 & n30369;
  assign n30451 = ~pi190 & ~n17051;
  assign n30452 = pi763 & ~n30451;
  assign n30453 = pi190 & n16998;
  assign n30454 = n30452 & ~n30453;
  assign n30455 = pi190 & n16935;
  assign n30456 = ~pi190 & n16853;
  assign n30457 = ~pi763 & ~n30456;
  assign n30458 = ~n30455 & n30457;
  assign n30459 = pi39 & ~n30458;
  assign n30460 = ~n30454 & n30459;
  assign n30461 = pi190 & n17058;
  assign n30462 = ~pi190 & n17061;
  assign n30463 = ~pi763 & ~n30462;
  assign n30464 = ~n30461 & n30463;
  assign n30465 = ~pi190 & ~n17067;
  assign n30466 = pi190 & ~n17065;
  assign n30467 = ~n30465 & ~n30466;
  assign n30468 = pi763 & n30467;
  assign n30469 = ~pi39 & ~n30468;
  assign n30470 = ~n30464 & n30469;
  assign n30471 = ~pi38 & ~n30470;
  assign n30472 = ~n30460 & n30471;
  assign n30473 = ~n17079 & ~n30121;
  assign n30474 = pi190 & ~n30473;
  assign n30475 = n6097 & n30474;
  assign n30476 = ~pi763 & n23427;
  assign n30477 = ~n16917 & ~n30476;
  assign n30478 = ~pi39 & ~n30477;
  assign n30479 = ~pi190 & ~n30478;
  assign n30480 = pi38 & ~n30479;
  assign n30481 = ~n30475 & n30480;
  assign n30482 = ~n30472 & ~n30481;
  assign n30483 = pi699 & n30482;
  assign n30484 = ~n30450 & ~n30483;
  assign n30485 = n10020 & n30484;
  assign n30486 = ~n30310 & ~n30485;
  assign n30487 = ~pi625 & n30486;
  assign n30488 = ~pi1153 & ~n30487;
  assign n30489 = ~n30449 & n30488;
  assign n30490 = ~pi608 & ~n30328;
  assign n30491 = ~n30489 & n30490;
  assign n30492 = ~pi625 & n30371;
  assign n30493 = pi625 & n30486;
  assign n30494 = ~n30492 & ~n30493;
  assign n30495 = pi1153 & n30494;
  assign n30496 = ~n30332 & ~n30495;
  assign n30497 = pi608 & n30496;
  assign n30498 = ~n30491 & ~n30497;
  assign n30499 = pi778 & ~n30498;
  assign n30500 = ~pi778 & n30486;
  assign n30501 = ~n30499 & ~n30500;
  assign n30502 = ~pi609 & ~n30501;
  assign n30503 = ~pi1155 & ~n30502;
  assign n30504 = ~n30448 & n30503;
  assign n30505 = ~pi660 & ~n30379;
  assign n30506 = ~n30504 & n30505;
  assign n30507 = ~pi609 & n30335;
  assign n30508 = pi609 & ~n30501;
  assign n30509 = ~n30507 & ~n30508;
  assign n30510 = pi1155 & n30509;
  assign n30511 = ~n30383 & ~n30510;
  assign n30512 = pi660 & n30511;
  assign n30513 = ~n30506 & ~n30512;
  assign n30514 = pi785 & ~n30513;
  assign n30515 = ~pi785 & ~n30501;
  assign n30516 = ~n30514 & ~n30515;
  assign n30517 = ~pi618 & ~n30516;
  assign n30518 = ~pi1154 & ~n30517;
  assign n30519 = ~n30447 & n30518;
  assign n30520 = ~pi627 & ~n30391;
  assign n30521 = ~n30519 & n30520;
  assign n30522 = ~pi618 & n30337;
  assign n30523 = pi618 & ~n30516;
  assign n30524 = ~n30522 & ~n30523;
  assign n30525 = pi1154 & n30524;
  assign n30526 = ~n30395 & ~n30525;
  assign n30527 = pi627 & n30526;
  assign n30528 = ~n30521 & ~n30527;
  assign n30529 = pi781 & ~n30528;
  assign n30530 = ~pi781 & ~n30516;
  assign n30531 = ~n30529 & ~n30530;
  assign n30532 = ~pi789 & n30531;
  assign n30533 = ~pi619 & ~n30531;
  assign n30534 = pi619 & ~n30340;
  assign n30535 = ~pi1159 & ~n30534;
  assign n30536 = ~n30533 & n30535;
  assign n30537 = ~pi648 & ~n30536;
  assign n30538 = ~n30403 & n30537;
  assign n30539 = ~pi619 & ~n30340;
  assign n30540 = pi619 & ~n30531;
  assign n30541 = ~n30539 & ~n30540;
  assign n30542 = pi1159 & n30541;
  assign n30543 = ~n30407 & ~n30542;
  assign n30544 = pi648 & n30543;
  assign n30545 = ~n30538 & ~n30544;
  assign n30546 = pi789 & n30545;
  assign n30547 = ~n30532 & ~n30546;
  assign n30548 = n17356 & n30547;
  assign n30549 = ~pi626 & ~n30410;
  assign n30550 = pi626 & ~n30306;
  assign n30551 = n17181 & ~n30550;
  assign n30552 = ~n30549 & n30551;
  assign n30553 = n17350 & n30342;
  assign n30554 = pi626 & ~n30410;
  assign n30555 = ~pi626 & ~n30306;
  assign n30556 = n17180 & ~n30555;
  assign n30557 = ~n30554 & n30556;
  assign n30558 = ~n30553 & ~n30557;
  assign n30559 = ~n30552 & n30558;
  assign n30560 = pi788 & ~n30559;
  assign n30561 = n19788 & ~n30560;
  assign n30562 = ~n30548 & n30561;
  assign n30563 = ~n30446 & ~n30562;
  assign n30564 = n19637 & ~n30563;
  assign n30565 = ~pi647 & n30347;
  assign n30566 = pi647 & n30306;
  assign n30567 = n17245 & ~n30566;
  assign n30568 = ~n30565 & n30567;
  assign n30569 = ~n19987 & n30416;
  assign n30570 = pi647 & n30347;
  assign n30571 = n17244 & ~n30570;
  assign n30572 = ~pi647 & n30306;
  assign n30573 = n30571 & ~n30572;
  assign n30574 = ~n30569 & ~n30573;
  assign n30575 = ~n30568 & n30574;
  assign n30576 = pi787 & ~n30575;
  assign n30577 = ~n30564 & ~n30576;
  assign n30578 = pi644 & n30423;
  assign n30579 = ~pi644 & n30431;
  assign n30580 = pi790 & ~n30579;
  assign n30581 = ~n30578 & n30580;
  assign n30582 = n30577 & ~n30581;
  assign n30583 = ~n30434 & ~n30582;
  assign n30584 = ~po1038 & ~n30583;
  assign n30585 = ~pi190 & po1038;
  assign n30586 = ~pi832 & ~n30585;
  assign n30587 = ~n30584 & n30586;
  assign po347 = ~n30305 & ~n30587;
  assign n30589 = ~pi191 & ~n2934;
  assign n30590 = pi746 & n16510;
  assign n30591 = ~n30589 & ~n30590;
  assign n30592 = ~n17273 & ~n30591;
  assign n30593 = ~pi785 & ~n30592;
  assign n30594 = n16537 & n30590;
  assign n30595 = n30592 & ~n30594;
  assign n30596 = pi1155 & ~n30595;
  assign n30597 = ~pi1155 & ~n30589;
  assign n30598 = ~n30594 & n30597;
  assign n30599 = ~n30596 & ~n30598;
  assign n30600 = pi785 & ~n30599;
  assign n30601 = ~n30593 & ~n30600;
  assign n30602 = ~pi781 & ~n30601;
  assign n30603 = ~n17289 & n30601;
  assign n30604 = pi1154 & ~n30603;
  assign n30605 = ~n17292 & n30601;
  assign n30606 = ~pi1154 & ~n30605;
  assign n30607 = ~n30604 & ~n30606;
  assign n30608 = pi781 & ~n30607;
  assign n30609 = ~n30602 & ~n30608;
  assign n30610 = ~pi789 & ~n30609;
  assign n30611 = ~n22423 & n30609;
  assign n30612 = pi1159 & ~n30611;
  assign n30613 = ~n22426 & n30609;
  assign n30614 = ~pi1159 & ~n30613;
  assign n30615 = ~n30612 & ~n30614;
  assign n30616 = pi789 & ~n30615;
  assign n30617 = ~n30610 & ~n30616;
  assign n30618 = ~n17355 & n30617;
  assign n30619 = n17355 & n30589;
  assign n30620 = ~n30618 & ~n30619;
  assign n30621 = ~n16124 & ~n30620;
  assign n30622 = n16124 & n30589;
  assign n30623 = ~n30621 & ~n30622;
  assign n30624 = ~n19987 & n30623;
  assign n30625 = pi729 & n16742;
  assign n30626 = ~n30589 & ~n30625;
  assign n30627 = ~pi778 & ~n30626;
  assign n30628 = ~pi625 & n30625;
  assign n30629 = ~n30626 & ~n30628;
  assign n30630 = pi1153 & ~n30629;
  assign n30631 = ~pi1153 & ~n30589;
  assign n30632 = ~n30628 & n30631;
  assign n30633 = ~n30630 & ~n30632;
  assign n30634 = pi778 & n30633;
  assign n30635 = ~n30627 & ~n30634;
  assign n30636 = ~n17338 & ~n30635;
  assign n30637 = ~n17340 & n30636;
  assign n30638 = ~n17342 & n30637;
  assign n30639 = ~n17425 & n30638;
  assign n30640 = ~n17452 & n30639;
  assign n30641 = ~pi647 & n30640;
  assign n30642 = pi647 & n30589;
  assign n30643 = ~pi1157 & ~n30642;
  assign n30644 = ~n30641 & n30643;
  assign n30645 = ~pi647 & n30589;
  assign n30646 = pi647 & n30640;
  assign n30647 = pi1157 & ~n30646;
  assign n30648 = ~n30645 & n30647;
  assign n30649 = ~n30644 & ~n30648;
  assign n30650 = ~n17246 & ~n30649;
  assign n30651 = ~n30624 & ~n30650;
  assign n30652 = pi787 & ~n30651;
  assign n30653 = ~pi626 & ~n30617;
  assign n30654 = pi626 & ~n30589;
  assign n30655 = n17181 & ~n30654;
  assign n30656 = ~n30653 & n30655;
  assign n30657 = n17350 & n30638;
  assign n30658 = pi626 & ~n30617;
  assign n30659 = ~pi626 & ~n30589;
  assign n30660 = n17180 & ~n30659;
  assign n30661 = ~n30658 & n30660;
  assign n30662 = ~n30657 & ~n30661;
  assign n30663 = ~n30656 & n30662;
  assign n30664 = pi788 & ~n30663;
  assign n30665 = pi618 & n30636;
  assign n30666 = pi609 & ~n30635;
  assign n30667 = ~n16393 & ~n30626;
  assign n30668 = pi625 & n30667;
  assign n30669 = n30591 & ~n30667;
  assign n30670 = ~n30668 & ~n30669;
  assign n30671 = n30631 & ~n30670;
  assign n30672 = ~pi608 & ~n30630;
  assign n30673 = ~n30671 & n30672;
  assign n30674 = pi1153 & ~n30668;
  assign n30675 = n30591 & n30674;
  assign n30676 = ~n30632 & ~n30675;
  assign n30677 = pi608 & n30676;
  assign n30678 = ~n30673 & ~n30677;
  assign n30679 = pi778 & ~n30678;
  assign n30680 = ~pi778 & ~n30669;
  assign n30681 = ~n30679 & ~n30680;
  assign n30682 = ~pi609 & ~n30681;
  assign n30683 = ~pi1155 & ~n30682;
  assign n30684 = ~n30666 & n30683;
  assign n30685 = ~pi660 & ~n30596;
  assign n30686 = ~n30684 & n30685;
  assign n30687 = ~pi609 & ~n30635;
  assign n30688 = pi609 & ~n30681;
  assign n30689 = ~n30687 & ~n30688;
  assign n30690 = pi1155 & n30689;
  assign n30691 = ~n30598 & ~n30690;
  assign n30692 = pi660 & n30691;
  assign n30693 = ~n30686 & ~n30692;
  assign n30694 = pi785 & ~n30693;
  assign n30695 = ~pi785 & ~n30681;
  assign n30696 = ~n30694 & ~n30695;
  assign n30697 = ~pi618 & ~n30696;
  assign n30698 = ~pi1154 & ~n30697;
  assign n30699 = ~n30665 & n30698;
  assign n30700 = ~pi627 & ~n30604;
  assign n30701 = ~n30699 & n30700;
  assign n30702 = ~pi618 & n30636;
  assign n30703 = pi618 & ~n30696;
  assign n30704 = ~n30702 & ~n30703;
  assign n30705 = pi1154 & n30704;
  assign n30706 = ~n30606 & ~n30705;
  assign n30707 = pi627 & n30706;
  assign n30708 = ~n30701 & ~n30707;
  assign n30709 = pi781 & ~n30708;
  assign n30710 = ~pi781 & ~n30696;
  assign n30711 = ~n30709 & ~n30710;
  assign n30712 = ~pi619 & ~n30711;
  assign n30713 = pi619 & n30637;
  assign n30714 = ~pi1159 & ~n30713;
  assign n30715 = ~n30712 & n30714;
  assign n30716 = ~pi648 & ~n30715;
  assign n30717 = ~n30612 & n30716;
  assign n30718 = ~pi619 & n30637;
  assign n30719 = pi619 & ~n30711;
  assign n30720 = ~n30718 & ~n30719;
  assign n30721 = pi1159 & n30720;
  assign n30722 = ~n30614 & ~n30721;
  assign n30723 = pi648 & n30722;
  assign n30724 = ~n30717 & ~n30723;
  assign n30725 = pi789 & n30724;
  assign n30726 = ~pi789 & n30711;
  assign n30727 = n17356 & ~n30726;
  assign n30728 = ~n30725 & n30727;
  assign n30729 = ~n30664 & ~n30728;
  assign n30730 = n19788 & ~n30729;
  assign n30731 = n20275 & n30639;
  assign n30732 = n17449 & ~n30620;
  assign n30733 = ~pi629 & ~n30732;
  assign n30734 = ~n30731 & n30733;
  assign n30735 = n17448 & ~n30620;
  assign n30736 = n20281 & n30639;
  assign n30737 = pi629 & ~n30736;
  assign n30738 = ~n30735 & n30737;
  assign n30739 = ~n30734 & ~n30738;
  assign n30740 = pi792 & n30739;
  assign n30741 = n19637 & ~n30740;
  assign n30742 = ~n30730 & n30741;
  assign n30743 = ~n30652 & ~n30742;
  assign n30744 = pi644 & n30743;
  assign n30745 = ~pi787 & ~n30640;
  assign n30746 = pi787 & ~n30649;
  assign n30747 = ~n30745 & ~n30746;
  assign n30748 = ~pi644 & n30747;
  assign n30749 = pi715 & ~n30748;
  assign n30750 = ~n30744 & n30749;
  assign n30751 = ~n17247 & ~n30623;
  assign n30752 = n17247 & n30589;
  assign n30753 = ~n30751 & ~n30752;
  assign n30754 = pi644 & ~n30753;
  assign n30755 = ~pi644 & n30589;
  assign n30756 = ~pi715 & ~n30755;
  assign n30757 = ~n30754 & n30756;
  assign n30758 = pi1160 & ~n30757;
  assign n30759 = ~n30750 & n30758;
  assign n30760 = ~pi644 & ~n30753;
  assign n30761 = pi715 & ~n30760;
  assign n30762 = pi644 & n30589;
  assign n30763 = n30761 & ~n30762;
  assign n30764 = pi644 & n30747;
  assign n30765 = ~pi644 & n30743;
  assign n30766 = ~pi715 & ~n30765;
  assign n30767 = ~n30764 & n30766;
  assign n30768 = ~pi1160 & ~n30767;
  assign n30769 = ~n30763 & n30768;
  assign n30770 = ~n30759 & ~n30769;
  assign n30771 = pi790 & ~n30770;
  assign n30772 = ~pi790 & n30743;
  assign n30773 = pi832 & ~n30772;
  assign n30774 = ~n30771 & n30773;
  assign n30775 = ~pi191 & ~n16527;
  assign n30776 = n17451 & ~n30775;
  assign n30777 = n17159 & ~n30775;
  assign n30778 = n16593 & ~n30775;
  assign n30779 = pi191 & ~n10020;
  assign n30780 = pi191 & n17589;
  assign n30781 = ~pi191 & n17592;
  assign n30782 = ~pi38 & ~n30781;
  assign n30783 = ~n30780 & n30782;
  assign n30784 = ~pi191 & ~n16508;
  assign n30785 = n16744 & ~n30784;
  assign n30786 = pi729 & ~n30785;
  assign n30787 = ~n30783 & n30786;
  assign n30788 = ~pi191 & ~pi729;
  assign n30789 = ~n16526 & n30788;
  assign n30790 = ~n30787 & ~n30789;
  assign n30791 = n10020 & n30790;
  assign n30792 = ~n30779 & ~n30791;
  assign n30793 = ~pi778 & ~n30792;
  assign n30794 = pi625 & n30792;
  assign n30795 = pi1153 & ~n30794;
  assign n30796 = ~pi625 & n30775;
  assign n30797 = n30795 & ~n30796;
  assign n30798 = ~pi625 & n30792;
  assign n30799 = ~pi1153 & ~n30798;
  assign n30800 = pi625 & n30775;
  assign n30801 = n30799 & ~n30800;
  assign n30802 = ~n30797 & ~n30801;
  assign n30803 = pi778 & ~n30802;
  assign n30804 = ~n30793 & ~n30803;
  assign n30805 = ~n16593 & ~n30804;
  assign n30806 = ~n30778 & ~n30805;
  assign n30807 = ~n16589 & n30806;
  assign n30808 = n16589 & n30775;
  assign n30809 = ~n30807 & ~n30808;
  assign n30810 = ~n17159 & n30809;
  assign n30811 = ~n30777 & ~n30810;
  assign n30812 = ~n17183 & n30811;
  assign n30813 = n17183 & n30775;
  assign n30814 = ~n30812 & ~n30813;
  assign n30815 = ~n17451 & n30814;
  assign n30816 = ~n30776 & ~n30815;
  assign n30817 = ~n18767 & n30816;
  assign n30818 = n18767 & n30775;
  assign n30819 = ~n30817 & ~n30818;
  assign n30820 = ~pi644 & ~n30819;
  assign n30821 = pi715 & ~n30820;
  assign n30822 = n17247 & ~n30775;
  assign n30823 = ~pi746 & n16355;
  assign n30824 = pi191 & n16501;
  assign n30825 = ~n30823 & ~n30824;
  assign n30826 = pi39 & ~n30825;
  assign n30827 = pi746 & ~n16461;
  assign n30828 = pi191 & ~n30827;
  assign n30829 = ~n21813 & ~n30828;
  assign n30830 = ~pi191 & n16449;
  assign n30831 = pi746 & n30830;
  assign n30832 = n30829 & ~n30831;
  assign n30833 = ~n30826 & n30832;
  assign n30834 = ~pi38 & ~n30833;
  assign n30835 = pi746 & n16511;
  assign n30836 = ~n30784 & ~n30835;
  assign n30837 = pi38 & n30836;
  assign n30838 = ~n30834 & ~n30837;
  assign n30839 = n10020 & ~n30838;
  assign n30840 = ~n30779 & ~n30839;
  assign n30841 = ~n16521 & ~n30840;
  assign n30842 = n16521 & ~n30775;
  assign n30843 = ~n30841 & ~n30842;
  assign n30844 = ~pi785 & ~n30843;
  assign n30845 = ~n16532 & ~n30775;
  assign n30846 = pi609 & n30841;
  assign n30847 = ~n30845 & ~n30846;
  assign n30848 = pi1155 & ~n30847;
  assign n30849 = ~n16537 & ~n30775;
  assign n30850 = ~pi609 & n30841;
  assign n30851 = ~n30849 & ~n30850;
  assign n30852 = ~pi1155 & ~n30851;
  assign n30853 = ~n30848 & ~n30852;
  assign n30854 = pi785 & ~n30853;
  assign n30855 = ~n30844 & ~n30854;
  assign n30856 = ~pi781 & ~n30855;
  assign n30857 = pi618 & n30855;
  assign n30858 = ~pi618 & n30775;
  assign n30859 = pi1154 & ~n30858;
  assign n30860 = ~n30857 & n30859;
  assign n30861 = ~pi618 & n30855;
  assign n30862 = pi618 & n30775;
  assign n30863 = ~pi1154 & ~n30862;
  assign n30864 = ~n30861 & n30863;
  assign n30865 = ~n30860 & ~n30864;
  assign n30866 = pi781 & ~n30865;
  assign n30867 = ~n30856 & ~n30866;
  assign n30868 = ~pi789 & ~n30867;
  assign n30869 = pi619 & n30867;
  assign n30870 = ~pi619 & n30775;
  assign n30871 = pi1159 & ~n30870;
  assign n30872 = ~n30869 & n30871;
  assign n30873 = ~pi619 & n30867;
  assign n30874 = pi619 & n30775;
  assign n30875 = ~pi1159 & ~n30874;
  assign n30876 = ~n30873 & n30875;
  assign n30877 = ~n30872 & ~n30876;
  assign n30878 = pi789 & ~n30877;
  assign n30879 = ~n30868 & ~n30878;
  assign n30880 = ~n17355 & n30879;
  assign n30881 = n17355 & n30775;
  assign n30882 = ~n30880 & ~n30881;
  assign n30883 = ~n16124 & ~n30882;
  assign n30884 = n16124 & n30775;
  assign n30885 = ~n30883 & ~n30884;
  assign n30886 = ~n17247 & n30885;
  assign n30887 = ~n30822 & ~n30886;
  assign n30888 = pi644 & n30887;
  assign n30889 = ~pi644 & n30775;
  assign n30890 = ~pi715 & ~n30889;
  assign n30891 = ~n30888 & n30890;
  assign n30892 = pi1160 & ~n30891;
  assign n30893 = ~n30821 & n30892;
  assign n30894 = pi644 & ~n30819;
  assign n30895 = ~pi715 & ~n30894;
  assign n30896 = ~pi644 & n30887;
  assign n30897 = pi644 & n30775;
  assign n30898 = ~n30896 & ~n30897;
  assign n30899 = pi715 & n30898;
  assign n30900 = ~pi1160 & ~n30899;
  assign n30901 = ~n30895 & n30900;
  assign n30902 = ~n30893 & ~n30901;
  assign n30903 = pi790 & ~n30902;
  assign n30904 = ~n19999 & n30882;
  assign n30905 = pi628 & ~n30814;
  assign n30906 = n16121 & ~n30905;
  assign n30907 = ~pi628 & n30775;
  assign n30908 = n30906 & ~n30907;
  assign n30909 = ~pi628 & ~n30814;
  assign n30910 = pi628 & n30775;
  assign n30911 = n16122 & ~n30910;
  assign n30912 = ~n30909 & n30911;
  assign n30913 = ~n30908 & ~n30912;
  assign n30914 = ~n30904 & n30913;
  assign n30915 = pi792 & ~n30914;
  assign n30916 = pi618 & n30806;
  assign n30917 = pi609 & n30804;
  assign n30918 = pi625 & n30840;
  assign n30919 = ~pi729 & n30838;
  assign n30920 = ~pi191 & ~n17051;
  assign n30921 = pi746 & ~n30920;
  assign n30922 = pi191 & n16998;
  assign n30923 = n30921 & ~n30922;
  assign n30924 = pi191 & n16935;
  assign n30925 = ~pi191 & n16853;
  assign n30926 = ~pi746 & ~n30925;
  assign n30927 = ~n30924 & n30926;
  assign n30928 = pi39 & ~n30927;
  assign n30929 = ~n30923 & n30928;
  assign n30930 = pi191 & n17058;
  assign n30931 = ~pi191 & n17061;
  assign n30932 = ~pi746 & ~n30931;
  assign n30933 = ~n30930 & n30932;
  assign n30934 = ~pi191 & ~n17067;
  assign n30935 = pi191 & ~n17065;
  assign n30936 = ~n30934 & ~n30935;
  assign n30937 = pi746 & n30936;
  assign n30938 = ~pi39 & ~n30937;
  assign n30939 = ~n30933 & n30938;
  assign n30940 = ~pi38 & ~n30939;
  assign n30941 = ~n30929 & n30940;
  assign n30942 = ~n17079 & ~n30590;
  assign n30943 = pi191 & ~n30942;
  assign n30944 = n6097 & n30943;
  assign n30945 = ~pi746 & n23427;
  assign n30946 = ~n16917 & ~n30945;
  assign n30947 = ~pi39 & ~n30946;
  assign n30948 = ~pi191 & ~n30947;
  assign n30949 = pi38 & ~n30948;
  assign n30950 = ~n30944 & n30949;
  assign n30951 = ~n30941 & ~n30950;
  assign n30952 = pi729 & n30951;
  assign n30953 = ~n30919 & ~n30952;
  assign n30954 = n10020 & n30953;
  assign n30955 = ~n30779 & ~n30954;
  assign n30956 = ~pi625 & n30955;
  assign n30957 = ~pi1153 & ~n30956;
  assign n30958 = ~n30918 & n30957;
  assign n30959 = ~pi608 & ~n30797;
  assign n30960 = ~n30958 & n30959;
  assign n30961 = ~pi625 & n30840;
  assign n30962 = pi625 & n30955;
  assign n30963 = ~n30961 & ~n30962;
  assign n30964 = pi1153 & n30963;
  assign n30965 = ~n30801 & ~n30964;
  assign n30966 = pi608 & n30965;
  assign n30967 = ~n30960 & ~n30966;
  assign n30968 = pi778 & ~n30967;
  assign n30969 = ~pi778 & n30955;
  assign n30970 = ~n30968 & ~n30969;
  assign n30971 = ~pi609 & ~n30970;
  assign n30972 = ~pi1155 & ~n30971;
  assign n30973 = ~n30917 & n30972;
  assign n30974 = ~pi660 & ~n30848;
  assign n30975 = ~n30973 & n30974;
  assign n30976 = ~pi609 & n30804;
  assign n30977 = pi609 & ~n30970;
  assign n30978 = ~n30976 & ~n30977;
  assign n30979 = pi1155 & n30978;
  assign n30980 = ~n30852 & ~n30979;
  assign n30981 = pi660 & n30980;
  assign n30982 = ~n30975 & ~n30981;
  assign n30983 = pi785 & ~n30982;
  assign n30984 = ~pi785 & ~n30970;
  assign n30985 = ~n30983 & ~n30984;
  assign n30986 = ~pi618 & ~n30985;
  assign n30987 = ~pi1154 & ~n30986;
  assign n30988 = ~n30916 & n30987;
  assign n30989 = ~pi627 & ~n30860;
  assign n30990 = ~n30988 & n30989;
  assign n30991 = ~pi618 & n30806;
  assign n30992 = pi618 & ~n30985;
  assign n30993 = ~n30991 & ~n30992;
  assign n30994 = pi1154 & n30993;
  assign n30995 = ~n30864 & ~n30994;
  assign n30996 = pi627 & n30995;
  assign n30997 = ~n30990 & ~n30996;
  assign n30998 = pi781 & ~n30997;
  assign n30999 = ~pi781 & ~n30985;
  assign n31000 = ~n30998 & ~n30999;
  assign n31001 = ~pi789 & n31000;
  assign n31002 = ~pi619 & ~n31000;
  assign n31003 = pi619 & ~n30809;
  assign n31004 = ~pi1159 & ~n31003;
  assign n31005 = ~n31002 & n31004;
  assign n31006 = ~pi648 & ~n31005;
  assign n31007 = ~n30872 & n31006;
  assign n31008 = ~pi619 & ~n30809;
  assign n31009 = pi619 & ~n31000;
  assign n31010 = ~n31008 & ~n31009;
  assign n31011 = pi1159 & n31010;
  assign n31012 = ~n30876 & ~n31011;
  assign n31013 = pi648 & n31012;
  assign n31014 = ~n31007 & ~n31013;
  assign n31015 = pi789 & n31014;
  assign n31016 = ~n31001 & ~n31015;
  assign n31017 = n17356 & n31016;
  assign n31018 = ~pi626 & ~n30879;
  assign n31019 = pi626 & ~n30775;
  assign n31020 = n17181 & ~n31019;
  assign n31021 = ~n31018 & n31020;
  assign n31022 = n17350 & n30811;
  assign n31023 = pi626 & ~n30879;
  assign n31024 = ~pi626 & ~n30775;
  assign n31025 = n17180 & ~n31024;
  assign n31026 = ~n31023 & n31025;
  assign n31027 = ~n31022 & ~n31026;
  assign n31028 = ~n31021 & n31027;
  assign n31029 = pi788 & ~n31028;
  assign n31030 = n19788 & ~n31029;
  assign n31031 = ~n31017 & n31030;
  assign n31032 = ~n30915 & ~n31031;
  assign n31033 = n19637 & ~n31032;
  assign n31034 = ~pi647 & n30816;
  assign n31035 = pi647 & n30775;
  assign n31036 = n17245 & ~n31035;
  assign n31037 = ~n31034 & n31036;
  assign n31038 = ~n19987 & n30885;
  assign n31039 = pi647 & n30816;
  assign n31040 = n17244 & ~n31039;
  assign n31041 = ~pi647 & n30775;
  assign n31042 = n31040 & ~n31041;
  assign n31043 = ~n31038 & ~n31042;
  assign n31044 = ~n31037 & n31043;
  assign n31045 = pi787 & ~n31044;
  assign n31046 = ~n31033 & ~n31045;
  assign n31047 = pi644 & n30892;
  assign n31048 = ~pi644 & n30900;
  assign n31049 = pi790 & ~n31048;
  assign n31050 = ~n31047 & n31049;
  assign n31051 = n31046 & ~n31050;
  assign n31052 = ~n30903 & ~n31051;
  assign n31053 = ~po1038 & ~n31052;
  assign n31054 = ~pi191 & po1038;
  assign n31055 = ~pi832 & ~n31054;
  assign n31056 = ~n31053 & n31055;
  assign po348 = ~n30774 & ~n31056;
  assign n31058 = ~pi192 & ~n2934;
  assign n31059 = pi764 & n16510;
  assign n31060 = ~n31058 & ~n31059;
  assign n31061 = ~n17273 & ~n31060;
  assign n31062 = ~pi785 & ~n31061;
  assign n31063 = n16537 & n31059;
  assign n31064 = n31061 & ~n31063;
  assign n31065 = pi1155 & ~n31064;
  assign n31066 = ~pi1155 & ~n31058;
  assign n31067 = ~n31063 & n31066;
  assign n31068 = ~n31065 & ~n31067;
  assign n31069 = pi785 & ~n31068;
  assign n31070 = ~n31062 & ~n31069;
  assign n31071 = ~pi781 & ~n31070;
  assign n31072 = ~n17289 & n31070;
  assign n31073 = pi1154 & ~n31072;
  assign n31074 = ~n17292 & n31070;
  assign n31075 = ~pi1154 & ~n31074;
  assign n31076 = ~n31073 & ~n31075;
  assign n31077 = pi781 & ~n31076;
  assign n31078 = ~n31071 & ~n31077;
  assign n31079 = ~pi789 & ~n31078;
  assign n31080 = ~n22423 & n31078;
  assign n31081 = pi1159 & ~n31080;
  assign n31082 = ~n22426 & n31078;
  assign n31083 = ~pi1159 & ~n31082;
  assign n31084 = ~n31081 & ~n31083;
  assign n31085 = pi789 & ~n31084;
  assign n31086 = ~n31079 & ~n31085;
  assign n31087 = ~n17355 & n31086;
  assign n31088 = n17355 & n31058;
  assign n31089 = ~n31087 & ~n31088;
  assign n31090 = ~n16124 & ~n31089;
  assign n31091 = n16124 & n31058;
  assign n31092 = ~n31090 & ~n31091;
  assign n31093 = ~n19987 & n31092;
  assign n31094 = pi691 & n16742;
  assign n31095 = ~n31058 & ~n31094;
  assign n31096 = ~pi778 & ~n31095;
  assign n31097 = ~pi625 & n31094;
  assign n31098 = ~n31095 & ~n31097;
  assign n31099 = pi1153 & ~n31098;
  assign n31100 = ~pi1153 & ~n31058;
  assign n31101 = ~n31097 & n31100;
  assign n31102 = ~n31099 & ~n31101;
  assign n31103 = pi778 & n31102;
  assign n31104 = ~n31096 & ~n31103;
  assign n31105 = ~n17338 & ~n31104;
  assign n31106 = ~n17340 & n31105;
  assign n31107 = ~n17342 & n31106;
  assign n31108 = ~n17425 & n31107;
  assign n31109 = ~n17452 & n31108;
  assign n31110 = ~pi647 & n31109;
  assign n31111 = pi647 & n31058;
  assign n31112 = ~pi1157 & ~n31111;
  assign n31113 = ~n31110 & n31112;
  assign n31114 = ~pi647 & n31058;
  assign n31115 = pi647 & n31109;
  assign n31116 = pi1157 & ~n31115;
  assign n31117 = ~n31114 & n31116;
  assign n31118 = ~n31113 & ~n31117;
  assign n31119 = ~n17246 & ~n31118;
  assign n31120 = ~n31093 & ~n31119;
  assign n31121 = pi787 & ~n31120;
  assign n31122 = ~pi626 & ~n31086;
  assign n31123 = pi626 & ~n31058;
  assign n31124 = n17181 & ~n31123;
  assign n31125 = ~n31122 & n31124;
  assign n31126 = n17350 & n31107;
  assign n31127 = pi626 & ~n31086;
  assign n31128 = ~pi626 & ~n31058;
  assign n31129 = n17180 & ~n31128;
  assign n31130 = ~n31127 & n31129;
  assign n31131 = ~n31126 & ~n31130;
  assign n31132 = ~n31125 & n31131;
  assign n31133 = pi788 & ~n31132;
  assign n31134 = pi618 & n31105;
  assign n31135 = pi609 & ~n31104;
  assign n31136 = ~n16393 & ~n31095;
  assign n31137 = pi625 & n31136;
  assign n31138 = n31060 & ~n31136;
  assign n31139 = ~n31137 & ~n31138;
  assign n31140 = n31100 & ~n31139;
  assign n31141 = ~pi608 & ~n31099;
  assign n31142 = ~n31140 & n31141;
  assign n31143 = pi1153 & ~n31137;
  assign n31144 = n31060 & n31143;
  assign n31145 = ~n31101 & ~n31144;
  assign n31146 = pi608 & n31145;
  assign n31147 = ~n31142 & ~n31146;
  assign n31148 = pi778 & ~n31147;
  assign n31149 = ~pi778 & ~n31138;
  assign n31150 = ~n31148 & ~n31149;
  assign n31151 = ~pi609 & ~n31150;
  assign n31152 = ~pi1155 & ~n31151;
  assign n31153 = ~n31135 & n31152;
  assign n31154 = ~pi660 & ~n31065;
  assign n31155 = ~n31153 & n31154;
  assign n31156 = ~pi609 & ~n31104;
  assign n31157 = pi609 & ~n31150;
  assign n31158 = ~n31156 & ~n31157;
  assign n31159 = pi1155 & n31158;
  assign n31160 = ~n31067 & ~n31159;
  assign n31161 = pi660 & n31160;
  assign n31162 = ~n31155 & ~n31161;
  assign n31163 = pi785 & ~n31162;
  assign n31164 = ~pi785 & ~n31150;
  assign n31165 = ~n31163 & ~n31164;
  assign n31166 = ~pi618 & ~n31165;
  assign n31167 = ~pi1154 & ~n31166;
  assign n31168 = ~n31134 & n31167;
  assign n31169 = ~pi627 & ~n31073;
  assign n31170 = ~n31168 & n31169;
  assign n31171 = ~pi618 & n31105;
  assign n31172 = pi618 & ~n31165;
  assign n31173 = ~n31171 & ~n31172;
  assign n31174 = pi1154 & n31173;
  assign n31175 = ~n31075 & ~n31174;
  assign n31176 = pi627 & n31175;
  assign n31177 = ~n31170 & ~n31176;
  assign n31178 = pi781 & ~n31177;
  assign n31179 = ~pi781 & ~n31165;
  assign n31180 = ~n31178 & ~n31179;
  assign n31181 = ~pi619 & ~n31180;
  assign n31182 = pi619 & n31106;
  assign n31183 = ~pi1159 & ~n31182;
  assign n31184 = ~n31181 & n31183;
  assign n31185 = ~pi648 & ~n31184;
  assign n31186 = ~n31081 & n31185;
  assign n31187 = ~pi619 & n31106;
  assign n31188 = pi619 & ~n31180;
  assign n31189 = ~n31187 & ~n31188;
  assign n31190 = pi1159 & n31189;
  assign n31191 = ~n31083 & ~n31190;
  assign n31192 = pi648 & n31191;
  assign n31193 = ~n31186 & ~n31192;
  assign n31194 = pi789 & n31193;
  assign n31195 = ~pi789 & n31180;
  assign n31196 = n17356 & ~n31195;
  assign n31197 = ~n31194 & n31196;
  assign n31198 = ~n31133 & ~n31197;
  assign n31199 = n19788 & ~n31198;
  assign n31200 = n20275 & n31108;
  assign n31201 = n17449 & ~n31089;
  assign n31202 = ~pi629 & ~n31201;
  assign n31203 = ~n31200 & n31202;
  assign n31204 = n17448 & ~n31089;
  assign n31205 = n20281 & n31108;
  assign n31206 = pi629 & ~n31205;
  assign n31207 = ~n31204 & n31206;
  assign n31208 = ~n31203 & ~n31207;
  assign n31209 = pi792 & n31208;
  assign n31210 = n19637 & ~n31209;
  assign n31211 = ~n31199 & n31210;
  assign n31212 = ~n31121 & ~n31211;
  assign n31213 = pi644 & n31212;
  assign n31214 = ~pi787 & ~n31109;
  assign n31215 = pi787 & ~n31118;
  assign n31216 = ~n31214 & ~n31215;
  assign n31217 = ~pi644 & n31216;
  assign n31218 = pi715 & ~n31217;
  assign n31219 = ~n31213 & n31218;
  assign n31220 = ~n17247 & ~n31092;
  assign n31221 = n17247 & n31058;
  assign n31222 = ~n31220 & ~n31221;
  assign n31223 = pi644 & ~n31222;
  assign n31224 = ~pi644 & n31058;
  assign n31225 = ~pi715 & ~n31224;
  assign n31226 = ~n31223 & n31225;
  assign n31227 = pi1160 & ~n31226;
  assign n31228 = ~n31219 & n31227;
  assign n31229 = ~pi644 & ~n31222;
  assign n31230 = pi715 & ~n31229;
  assign n31231 = pi644 & n31058;
  assign n31232 = n31230 & ~n31231;
  assign n31233 = pi644 & n31216;
  assign n31234 = ~pi644 & n31212;
  assign n31235 = ~pi715 & ~n31234;
  assign n31236 = ~n31233 & n31235;
  assign n31237 = ~pi1160 & ~n31236;
  assign n31238 = ~n31232 & n31237;
  assign n31239 = ~n31228 & ~n31238;
  assign n31240 = pi790 & ~n31239;
  assign n31241 = ~pi790 & n31212;
  assign n31242 = pi832 & ~n31241;
  assign n31243 = ~n31240 & n31242;
  assign n31244 = ~pi192 & ~n16527;
  assign n31245 = n17451 & ~n31244;
  assign n31246 = n17159 & ~n31244;
  assign n31247 = n16593 & ~n31244;
  assign n31248 = pi192 & ~n10020;
  assign n31249 = pi192 & n17589;
  assign n31250 = ~pi192 & n17592;
  assign n31251 = ~pi38 & ~n31250;
  assign n31252 = ~n31249 & n31251;
  assign n31253 = ~pi192 & ~n16508;
  assign n31254 = n16744 & ~n31253;
  assign n31255 = pi691 & ~n31254;
  assign n31256 = ~n31252 & n31255;
  assign n31257 = ~pi192 & ~pi691;
  assign n31258 = ~n16526 & n31257;
  assign n31259 = ~n31256 & ~n31258;
  assign n31260 = n10020 & n31259;
  assign n31261 = ~n31248 & ~n31260;
  assign n31262 = ~pi778 & ~n31261;
  assign n31263 = pi625 & n31261;
  assign n31264 = pi1153 & ~n31263;
  assign n31265 = ~pi625 & n31244;
  assign n31266 = n31264 & ~n31265;
  assign n31267 = ~pi625 & n31261;
  assign n31268 = ~pi1153 & ~n31267;
  assign n31269 = pi625 & n31244;
  assign n31270 = n31268 & ~n31269;
  assign n31271 = ~n31266 & ~n31270;
  assign n31272 = pi778 & ~n31271;
  assign n31273 = ~n31262 & ~n31272;
  assign n31274 = ~n16593 & ~n31273;
  assign n31275 = ~n31247 & ~n31274;
  assign n31276 = ~n16589 & n31275;
  assign n31277 = n16589 & n31244;
  assign n31278 = ~n31276 & ~n31277;
  assign n31279 = ~n17159 & n31278;
  assign n31280 = ~n31246 & ~n31279;
  assign n31281 = ~n17183 & n31280;
  assign n31282 = n17183 & n31244;
  assign n31283 = ~n31281 & ~n31282;
  assign n31284 = ~n17451 & n31283;
  assign n31285 = ~n31245 & ~n31284;
  assign n31286 = ~n18767 & n31285;
  assign n31287 = n18767 & n31244;
  assign n31288 = ~n31286 & ~n31287;
  assign n31289 = ~pi644 & ~n31288;
  assign n31290 = pi715 & ~n31289;
  assign n31291 = n17247 & ~n31244;
  assign n31292 = ~pi764 & n16355;
  assign n31293 = pi192 & n16501;
  assign n31294 = ~n31292 & ~n31293;
  assign n31295 = pi39 & ~n31294;
  assign n31296 = pi764 & ~n16461;
  assign n31297 = pi192 & ~n31296;
  assign n31298 = ~n21971 & ~n31297;
  assign n31299 = ~pi192 & n16449;
  assign n31300 = pi764 & n31299;
  assign n31301 = n31298 & ~n31300;
  assign n31302 = ~n31295 & n31301;
  assign n31303 = ~pi38 & ~n31302;
  assign n31304 = pi764 & n16511;
  assign n31305 = ~n31253 & ~n31304;
  assign n31306 = pi38 & n31305;
  assign n31307 = ~n31303 & ~n31306;
  assign n31308 = n10020 & ~n31307;
  assign n31309 = ~n31248 & ~n31308;
  assign n31310 = ~n16521 & ~n31309;
  assign n31311 = n16521 & ~n31244;
  assign n31312 = ~n31310 & ~n31311;
  assign n31313 = ~pi785 & ~n31312;
  assign n31314 = ~n16532 & ~n31244;
  assign n31315 = pi609 & n31310;
  assign n31316 = ~n31314 & ~n31315;
  assign n31317 = pi1155 & ~n31316;
  assign n31318 = ~n16537 & ~n31244;
  assign n31319 = ~pi609 & n31310;
  assign n31320 = ~n31318 & ~n31319;
  assign n31321 = ~pi1155 & ~n31320;
  assign n31322 = ~n31317 & ~n31321;
  assign n31323 = pi785 & ~n31322;
  assign n31324 = ~n31313 & ~n31323;
  assign n31325 = ~pi781 & ~n31324;
  assign n31326 = pi618 & n31324;
  assign n31327 = ~pi618 & n31244;
  assign n31328 = pi1154 & ~n31327;
  assign n31329 = ~n31326 & n31328;
  assign n31330 = ~pi618 & n31324;
  assign n31331 = pi618 & n31244;
  assign n31332 = ~pi1154 & ~n31331;
  assign n31333 = ~n31330 & n31332;
  assign n31334 = ~n31329 & ~n31333;
  assign n31335 = pi781 & ~n31334;
  assign n31336 = ~n31325 & ~n31335;
  assign n31337 = ~pi789 & ~n31336;
  assign n31338 = pi619 & n31336;
  assign n31339 = ~pi619 & n31244;
  assign n31340 = pi1159 & ~n31339;
  assign n31341 = ~n31338 & n31340;
  assign n31342 = ~pi619 & n31336;
  assign n31343 = pi619 & n31244;
  assign n31344 = ~pi1159 & ~n31343;
  assign n31345 = ~n31342 & n31344;
  assign n31346 = ~n31341 & ~n31345;
  assign n31347 = pi789 & ~n31346;
  assign n31348 = ~n31337 & ~n31347;
  assign n31349 = ~n17355 & n31348;
  assign n31350 = n17355 & n31244;
  assign n31351 = ~n31349 & ~n31350;
  assign n31352 = ~n16124 & ~n31351;
  assign n31353 = n16124 & n31244;
  assign n31354 = ~n31352 & ~n31353;
  assign n31355 = ~n17247 & n31354;
  assign n31356 = ~n31291 & ~n31355;
  assign n31357 = pi644 & n31356;
  assign n31358 = ~pi644 & n31244;
  assign n31359 = ~pi715 & ~n31358;
  assign n31360 = ~n31357 & n31359;
  assign n31361 = pi1160 & ~n31360;
  assign n31362 = ~n31290 & n31361;
  assign n31363 = pi644 & ~n31288;
  assign n31364 = ~pi715 & ~n31363;
  assign n31365 = ~pi644 & n31356;
  assign n31366 = pi644 & n31244;
  assign n31367 = ~n31365 & ~n31366;
  assign n31368 = pi715 & n31367;
  assign n31369 = ~pi1160 & ~n31368;
  assign n31370 = ~n31364 & n31369;
  assign n31371 = ~n31362 & ~n31370;
  assign n31372 = pi790 & ~n31371;
  assign n31373 = ~n19999 & n31351;
  assign n31374 = pi628 & ~n31283;
  assign n31375 = n16121 & ~n31374;
  assign n31376 = ~pi628 & n31244;
  assign n31377 = n31375 & ~n31376;
  assign n31378 = ~pi628 & ~n31283;
  assign n31379 = pi628 & n31244;
  assign n31380 = n16122 & ~n31379;
  assign n31381 = ~n31378 & n31380;
  assign n31382 = ~n31377 & ~n31381;
  assign n31383 = ~n31373 & n31382;
  assign n31384 = pi792 & ~n31383;
  assign n31385 = pi618 & n31275;
  assign n31386 = pi609 & n31273;
  assign n31387 = pi625 & n31309;
  assign n31388 = ~pi691 & n31307;
  assign n31389 = ~pi192 & ~n17051;
  assign n31390 = pi764 & ~n31389;
  assign n31391 = pi192 & n16998;
  assign n31392 = n31390 & ~n31391;
  assign n31393 = pi192 & n16935;
  assign n31394 = ~pi192 & n16853;
  assign n31395 = ~pi764 & ~n31394;
  assign n31396 = ~n31393 & n31395;
  assign n31397 = pi39 & ~n31396;
  assign n31398 = ~n31392 & n31397;
  assign n31399 = pi192 & n17058;
  assign n31400 = ~pi192 & n17061;
  assign n31401 = ~pi764 & ~n31400;
  assign n31402 = ~n31399 & n31401;
  assign n31403 = ~pi192 & ~n17067;
  assign n31404 = pi192 & ~n17065;
  assign n31405 = ~n31403 & ~n31404;
  assign n31406 = pi764 & n31405;
  assign n31407 = ~pi39 & ~n31406;
  assign n31408 = ~n31402 & n31407;
  assign n31409 = ~pi38 & ~n31408;
  assign n31410 = ~n31398 & n31409;
  assign n31411 = ~n17079 & ~n31059;
  assign n31412 = pi192 & ~n31411;
  assign n31413 = n6097 & n31412;
  assign n31414 = ~pi764 & n23427;
  assign n31415 = ~n16917 & ~n31414;
  assign n31416 = ~pi39 & ~n31415;
  assign n31417 = ~pi192 & ~n31416;
  assign n31418 = pi38 & ~n31417;
  assign n31419 = ~n31413 & n31418;
  assign n31420 = ~n31410 & ~n31419;
  assign n31421 = pi691 & n31420;
  assign n31422 = ~n31388 & ~n31421;
  assign n31423 = n10020 & n31422;
  assign n31424 = ~n31248 & ~n31423;
  assign n31425 = ~pi625 & n31424;
  assign n31426 = ~pi1153 & ~n31425;
  assign n31427 = ~n31387 & n31426;
  assign n31428 = ~pi608 & ~n31266;
  assign n31429 = ~n31427 & n31428;
  assign n31430 = ~pi625 & n31309;
  assign n31431 = pi625 & n31424;
  assign n31432 = ~n31430 & ~n31431;
  assign n31433 = pi1153 & n31432;
  assign n31434 = ~n31270 & ~n31433;
  assign n31435 = pi608 & n31434;
  assign n31436 = ~n31429 & ~n31435;
  assign n31437 = pi778 & ~n31436;
  assign n31438 = ~pi778 & n31424;
  assign n31439 = ~n31437 & ~n31438;
  assign n31440 = ~pi609 & ~n31439;
  assign n31441 = ~pi1155 & ~n31440;
  assign n31442 = ~n31386 & n31441;
  assign n31443 = ~pi660 & ~n31317;
  assign n31444 = ~n31442 & n31443;
  assign n31445 = ~pi609 & n31273;
  assign n31446 = pi609 & ~n31439;
  assign n31447 = ~n31445 & ~n31446;
  assign n31448 = pi1155 & n31447;
  assign n31449 = ~n31321 & ~n31448;
  assign n31450 = pi660 & n31449;
  assign n31451 = ~n31444 & ~n31450;
  assign n31452 = pi785 & ~n31451;
  assign n31453 = ~pi785 & ~n31439;
  assign n31454 = ~n31452 & ~n31453;
  assign n31455 = ~pi618 & ~n31454;
  assign n31456 = ~pi1154 & ~n31455;
  assign n31457 = ~n31385 & n31456;
  assign n31458 = ~pi627 & ~n31329;
  assign n31459 = ~n31457 & n31458;
  assign n31460 = ~pi618 & n31275;
  assign n31461 = pi618 & ~n31454;
  assign n31462 = ~n31460 & ~n31461;
  assign n31463 = pi1154 & n31462;
  assign n31464 = ~n31333 & ~n31463;
  assign n31465 = pi627 & n31464;
  assign n31466 = ~n31459 & ~n31465;
  assign n31467 = pi781 & ~n31466;
  assign n31468 = ~pi781 & ~n31454;
  assign n31469 = ~n31467 & ~n31468;
  assign n31470 = ~pi789 & n31469;
  assign n31471 = ~pi619 & ~n31469;
  assign n31472 = pi619 & ~n31278;
  assign n31473 = ~pi1159 & ~n31472;
  assign n31474 = ~n31471 & n31473;
  assign n31475 = ~pi648 & ~n31474;
  assign n31476 = ~n31341 & n31475;
  assign n31477 = ~pi619 & ~n31278;
  assign n31478 = pi619 & ~n31469;
  assign n31479 = ~n31477 & ~n31478;
  assign n31480 = pi1159 & n31479;
  assign n31481 = ~n31345 & ~n31480;
  assign n31482 = pi648 & n31481;
  assign n31483 = ~n31476 & ~n31482;
  assign n31484 = pi789 & n31483;
  assign n31485 = ~n31470 & ~n31484;
  assign n31486 = n17356 & n31485;
  assign n31487 = ~pi626 & ~n31348;
  assign n31488 = pi626 & ~n31244;
  assign n31489 = n17181 & ~n31488;
  assign n31490 = ~n31487 & n31489;
  assign n31491 = n17350 & n31280;
  assign n31492 = pi626 & ~n31348;
  assign n31493 = ~pi626 & ~n31244;
  assign n31494 = n17180 & ~n31493;
  assign n31495 = ~n31492 & n31494;
  assign n31496 = ~n31491 & ~n31495;
  assign n31497 = ~n31490 & n31496;
  assign n31498 = pi788 & ~n31497;
  assign n31499 = n19788 & ~n31498;
  assign n31500 = ~n31486 & n31499;
  assign n31501 = ~n31384 & ~n31500;
  assign n31502 = n19637 & ~n31501;
  assign n31503 = ~pi647 & n31285;
  assign n31504 = pi647 & n31244;
  assign n31505 = n17245 & ~n31504;
  assign n31506 = ~n31503 & n31505;
  assign n31507 = ~n19987 & n31354;
  assign n31508 = pi647 & n31285;
  assign n31509 = n17244 & ~n31508;
  assign n31510 = ~pi647 & n31244;
  assign n31511 = n31509 & ~n31510;
  assign n31512 = ~n31507 & ~n31511;
  assign n31513 = ~n31506 & n31512;
  assign n31514 = pi787 & ~n31513;
  assign n31515 = ~n31502 & ~n31514;
  assign n31516 = pi644 & n31361;
  assign n31517 = ~pi644 & n31369;
  assign n31518 = pi790 & ~n31517;
  assign n31519 = ~n31516 & n31518;
  assign n31520 = n31515 & ~n31519;
  assign n31521 = ~n31372 & ~n31520;
  assign n31522 = ~po1038 & ~n31521;
  assign n31523 = ~pi192 & po1038;
  assign n31524 = ~pi832 & ~n31523;
  assign n31525 = ~n31522 & n31524;
  assign po349 = ~n31243 & ~n31525;
  assign n31527 = ~pi193 & ~n2934;
  assign n31528 = pi739 & n16510;
  assign n31529 = ~n31527 & ~n31528;
  assign n31530 = ~n17273 & ~n31529;
  assign n31531 = ~pi785 & ~n31530;
  assign n31532 = n16537 & n31528;
  assign n31533 = n31530 & ~n31532;
  assign n31534 = pi1155 & ~n31533;
  assign n31535 = ~pi1155 & ~n31527;
  assign n31536 = ~n31532 & n31535;
  assign n31537 = ~n31534 & ~n31536;
  assign n31538 = pi785 & ~n31537;
  assign n31539 = ~n31531 & ~n31538;
  assign n31540 = ~pi781 & ~n31539;
  assign n31541 = ~n17289 & n31539;
  assign n31542 = pi1154 & ~n31541;
  assign n31543 = ~n17292 & n31539;
  assign n31544 = ~pi1154 & ~n31543;
  assign n31545 = ~n31542 & ~n31544;
  assign n31546 = pi781 & ~n31545;
  assign n31547 = ~n31540 & ~n31546;
  assign n31548 = ~pi789 & ~n31547;
  assign n31549 = ~n22423 & n31547;
  assign n31550 = pi1159 & ~n31549;
  assign n31551 = ~n22426 & n31547;
  assign n31552 = ~pi1159 & ~n31551;
  assign n31553 = ~n31550 & ~n31552;
  assign n31554 = pi789 & ~n31553;
  assign n31555 = ~n31548 & ~n31554;
  assign n31556 = ~n17355 & n31555;
  assign n31557 = n17355 & n31527;
  assign n31558 = ~n31556 & ~n31557;
  assign n31559 = ~n16124 & ~n31558;
  assign n31560 = n16124 & n31527;
  assign n31561 = ~n31559 & ~n31560;
  assign n31562 = ~n19987 & n31561;
  assign n31563 = pi690 & n16742;
  assign n31564 = ~n31527 & ~n31563;
  assign n31565 = ~pi778 & ~n31564;
  assign n31566 = ~pi625 & n31563;
  assign n31567 = ~n31564 & ~n31566;
  assign n31568 = pi1153 & ~n31567;
  assign n31569 = ~pi1153 & ~n31527;
  assign n31570 = ~n31566 & n31569;
  assign n31571 = ~n31568 & ~n31570;
  assign n31572 = pi778 & n31571;
  assign n31573 = ~n31565 & ~n31572;
  assign n31574 = ~n17338 & ~n31573;
  assign n31575 = ~n17340 & n31574;
  assign n31576 = ~n17342 & n31575;
  assign n31577 = ~n17425 & n31576;
  assign n31578 = ~n17452 & n31577;
  assign n31579 = ~pi647 & n31578;
  assign n31580 = pi647 & n31527;
  assign n31581 = ~pi1157 & ~n31580;
  assign n31582 = ~n31579 & n31581;
  assign n31583 = ~pi647 & n31527;
  assign n31584 = pi647 & n31578;
  assign n31585 = pi1157 & ~n31584;
  assign n31586 = ~n31583 & n31585;
  assign n31587 = ~n31582 & ~n31586;
  assign n31588 = ~n17246 & ~n31587;
  assign n31589 = ~n31562 & ~n31588;
  assign n31590 = pi787 & ~n31589;
  assign n31591 = ~pi626 & ~n31555;
  assign n31592 = pi626 & ~n31527;
  assign n31593 = n17181 & ~n31592;
  assign n31594 = ~n31591 & n31593;
  assign n31595 = n17350 & n31576;
  assign n31596 = pi626 & ~n31555;
  assign n31597 = ~pi626 & ~n31527;
  assign n31598 = n17180 & ~n31597;
  assign n31599 = ~n31596 & n31598;
  assign n31600 = ~n31595 & ~n31599;
  assign n31601 = ~n31594 & n31600;
  assign n31602 = pi788 & ~n31601;
  assign n31603 = pi618 & n31574;
  assign n31604 = pi609 & ~n31573;
  assign n31605 = ~n16393 & ~n31564;
  assign n31606 = pi625 & n31605;
  assign n31607 = n31529 & ~n31605;
  assign n31608 = ~n31606 & ~n31607;
  assign n31609 = n31569 & ~n31608;
  assign n31610 = ~pi608 & ~n31568;
  assign n31611 = ~n31609 & n31610;
  assign n31612 = pi1153 & ~n31606;
  assign n31613 = n31529 & n31612;
  assign n31614 = ~n31570 & ~n31613;
  assign n31615 = pi608 & n31614;
  assign n31616 = ~n31611 & ~n31615;
  assign n31617 = pi778 & ~n31616;
  assign n31618 = ~pi778 & ~n31607;
  assign n31619 = ~n31617 & ~n31618;
  assign n31620 = ~pi609 & ~n31619;
  assign n31621 = ~pi1155 & ~n31620;
  assign n31622 = ~n31604 & n31621;
  assign n31623 = ~pi660 & ~n31534;
  assign n31624 = ~n31622 & n31623;
  assign n31625 = ~pi609 & ~n31573;
  assign n31626 = pi609 & ~n31619;
  assign n31627 = ~n31625 & ~n31626;
  assign n31628 = pi1155 & n31627;
  assign n31629 = ~n31536 & ~n31628;
  assign n31630 = pi660 & n31629;
  assign n31631 = ~n31624 & ~n31630;
  assign n31632 = pi785 & ~n31631;
  assign n31633 = ~pi785 & ~n31619;
  assign n31634 = ~n31632 & ~n31633;
  assign n31635 = ~pi618 & ~n31634;
  assign n31636 = ~pi1154 & ~n31635;
  assign n31637 = ~n31603 & n31636;
  assign n31638 = ~pi627 & ~n31542;
  assign n31639 = ~n31637 & n31638;
  assign n31640 = ~pi618 & n31574;
  assign n31641 = pi618 & ~n31634;
  assign n31642 = ~n31640 & ~n31641;
  assign n31643 = pi1154 & n31642;
  assign n31644 = ~n31544 & ~n31643;
  assign n31645 = pi627 & n31644;
  assign n31646 = ~n31639 & ~n31645;
  assign n31647 = pi781 & ~n31646;
  assign n31648 = ~pi781 & ~n31634;
  assign n31649 = ~n31647 & ~n31648;
  assign n31650 = ~pi619 & ~n31649;
  assign n31651 = pi619 & n31575;
  assign n31652 = ~pi1159 & ~n31651;
  assign n31653 = ~n31650 & n31652;
  assign n31654 = ~pi648 & ~n31653;
  assign n31655 = ~n31550 & n31654;
  assign n31656 = ~pi619 & n31575;
  assign n31657 = pi619 & ~n31649;
  assign n31658 = ~n31656 & ~n31657;
  assign n31659 = pi1159 & n31658;
  assign n31660 = ~n31552 & ~n31659;
  assign n31661 = pi648 & n31660;
  assign n31662 = ~n31655 & ~n31661;
  assign n31663 = pi789 & n31662;
  assign n31664 = ~pi789 & n31649;
  assign n31665 = n17356 & ~n31664;
  assign n31666 = ~n31663 & n31665;
  assign n31667 = ~n31602 & ~n31666;
  assign n31668 = n19788 & ~n31667;
  assign n31669 = n20275 & n31577;
  assign n31670 = n17449 & ~n31558;
  assign n31671 = ~pi629 & ~n31670;
  assign n31672 = ~n31669 & n31671;
  assign n31673 = n17448 & ~n31558;
  assign n31674 = n20281 & n31577;
  assign n31675 = pi629 & ~n31674;
  assign n31676 = ~n31673 & n31675;
  assign n31677 = ~n31672 & ~n31676;
  assign n31678 = pi792 & n31677;
  assign n31679 = n19637 & ~n31678;
  assign n31680 = ~n31668 & n31679;
  assign n31681 = ~n31590 & ~n31680;
  assign n31682 = pi644 & n31681;
  assign n31683 = ~pi787 & ~n31578;
  assign n31684 = pi787 & ~n31587;
  assign n31685 = ~n31683 & ~n31684;
  assign n31686 = ~pi644 & n31685;
  assign n31687 = pi715 & ~n31686;
  assign n31688 = ~n31682 & n31687;
  assign n31689 = ~n17247 & ~n31561;
  assign n31690 = n17247 & n31527;
  assign n31691 = ~n31689 & ~n31690;
  assign n31692 = pi644 & ~n31691;
  assign n31693 = ~pi644 & n31527;
  assign n31694 = ~pi715 & ~n31693;
  assign n31695 = ~n31692 & n31694;
  assign n31696 = pi1160 & ~n31695;
  assign n31697 = ~n31688 & n31696;
  assign n31698 = ~pi644 & ~n31691;
  assign n31699 = pi715 & ~n31698;
  assign n31700 = pi644 & n31527;
  assign n31701 = n31699 & ~n31700;
  assign n31702 = pi644 & n31685;
  assign n31703 = ~pi644 & n31681;
  assign n31704 = ~pi715 & ~n31703;
  assign n31705 = ~n31702 & n31704;
  assign n31706 = ~pi1160 & ~n31705;
  assign n31707 = ~n31701 & n31706;
  assign n31708 = ~n31697 & ~n31707;
  assign n31709 = pi790 & ~n31708;
  assign n31710 = ~pi790 & n31681;
  assign n31711 = pi832 & ~n31710;
  assign n31712 = ~n31709 & n31711;
  assign n31713 = ~pi193 & ~n16527;
  assign n31714 = n17159 & ~n31713;
  assign n31715 = n16593 & ~n31713;
  assign n31716 = pi690 & n10020;
  assign n31717 = n31713 & ~n31716;
  assign n31718 = ~pi193 & n17592;
  assign n31719 = ~pi38 & ~pi193;
  assign n31720 = n19843 & ~n31719;
  assign n31721 = ~n31718 & ~n31720;
  assign n31722 = ~pi193 & ~n16508;
  assign n31723 = n16744 & ~n31722;
  assign n31724 = pi690 & ~n31723;
  assign n31725 = ~n31721 & n31724;
  assign n31726 = ~n31717 & ~n31725;
  assign n31727 = ~pi778 & n31726;
  assign n31728 = pi625 & ~n31726;
  assign n31729 = pi1153 & ~n31728;
  assign n31730 = ~pi625 & n31713;
  assign n31731 = n31729 & ~n31730;
  assign n31732 = ~pi625 & ~n31726;
  assign n31733 = ~pi1153 & ~n31732;
  assign n31734 = pi625 & n31713;
  assign n31735 = n31733 & ~n31734;
  assign n31736 = ~n31731 & ~n31735;
  assign n31737 = pi778 & ~n31736;
  assign n31738 = ~n31727 & ~n31737;
  assign n31739 = ~n16593 & ~n31738;
  assign n31740 = ~n31715 & ~n31739;
  assign n31741 = ~n16589 & n31740;
  assign n31742 = n16589 & n31713;
  assign n31743 = ~n31741 & ~n31742;
  assign n31744 = ~n17159 & n31743;
  assign n31745 = ~n31714 & ~n31744;
  assign n31746 = ~n17183 & n31745;
  assign n31747 = n17183 & n31713;
  assign n31748 = ~n31746 & ~n31747;
  assign n31749 = ~pi792 & n31748;
  assign n31750 = pi628 & ~n31748;
  assign n31751 = pi1156 & ~n31750;
  assign n31752 = ~pi628 & n31713;
  assign n31753 = n31751 & ~n31752;
  assign n31754 = ~pi628 & ~n31748;
  assign n31755 = pi628 & n31713;
  assign n31756 = ~pi1156 & ~n31755;
  assign n31757 = ~n31754 & n31756;
  assign n31758 = ~n31753 & ~n31757;
  assign n31759 = pi792 & ~n31758;
  assign n31760 = ~n31749 & ~n31759;
  assign n31761 = pi647 & ~n31760;
  assign n31762 = ~pi647 & ~n31713;
  assign n31763 = ~n31761 & ~n31762;
  assign n31764 = pi1157 & ~n31763;
  assign n31765 = ~pi647 & n31760;
  assign n31766 = ~pi1157 & ~n31765;
  assign n31767 = pi647 & n31713;
  assign n31768 = n31766 & ~n31767;
  assign n31769 = ~n31764 & ~n31768;
  assign n31770 = pi787 & ~n31769;
  assign n31771 = ~pi787 & ~n31760;
  assign n31772 = ~n31770 & ~n31771;
  assign n31773 = ~pi644 & n31772;
  assign n31774 = pi715 & ~n31773;
  assign n31775 = n17247 & ~n31713;
  assign n31776 = pi193 & ~n10020;
  assign n31777 = pi739 & n16511;
  assign n31778 = ~n31722 & ~n31777;
  assign n31779 = pi38 & ~n31778;
  assign n31780 = ~pi193 & n16449;
  assign n31781 = pi193 & ~n16503;
  assign n31782 = pi739 & ~n31781;
  assign n31783 = ~n31780 & n31782;
  assign n31784 = ~pi193 & ~pi739;
  assign n31785 = ~n16357 & n31784;
  assign n31786 = ~n31783 & ~n31785;
  assign n31787 = ~pi38 & ~n31786;
  assign n31788 = ~n31779 & ~n31787;
  assign n31789 = n10020 & n31788;
  assign n31790 = ~n31776 & ~n31789;
  assign n31791 = ~n16521 & ~n31790;
  assign n31792 = n16521 & ~n31713;
  assign n31793 = ~n31791 & ~n31792;
  assign n31794 = ~pi785 & ~n31793;
  assign n31795 = ~n16532 & ~n31713;
  assign n31796 = pi609 & n31791;
  assign n31797 = ~n31795 & ~n31796;
  assign n31798 = pi1155 & ~n31797;
  assign n31799 = ~n16537 & ~n31713;
  assign n31800 = ~pi609 & n31791;
  assign n31801 = ~n31799 & ~n31800;
  assign n31802 = ~pi1155 & ~n31801;
  assign n31803 = ~n31798 & ~n31802;
  assign n31804 = pi785 & ~n31803;
  assign n31805 = ~n31794 & ~n31804;
  assign n31806 = ~pi781 & ~n31805;
  assign n31807 = pi618 & n31805;
  assign n31808 = ~pi618 & n31713;
  assign n31809 = pi1154 & ~n31808;
  assign n31810 = ~n31807 & n31809;
  assign n31811 = ~pi618 & n31805;
  assign n31812 = pi618 & n31713;
  assign n31813 = ~pi1154 & ~n31812;
  assign n31814 = ~n31811 & n31813;
  assign n31815 = ~n31810 & ~n31814;
  assign n31816 = pi781 & ~n31815;
  assign n31817 = ~n31806 & ~n31816;
  assign n31818 = ~pi789 & ~n31817;
  assign n31819 = pi619 & n31817;
  assign n31820 = ~pi619 & n31713;
  assign n31821 = pi1159 & ~n31820;
  assign n31822 = ~n31819 & n31821;
  assign n31823 = ~pi619 & n31817;
  assign n31824 = pi619 & n31713;
  assign n31825 = ~pi1159 & ~n31824;
  assign n31826 = ~n31823 & n31825;
  assign n31827 = ~n31822 & ~n31826;
  assign n31828 = pi789 & ~n31827;
  assign n31829 = ~n31818 & ~n31828;
  assign n31830 = ~n17355 & n31829;
  assign n31831 = n17355 & n31713;
  assign n31832 = ~n31830 & ~n31831;
  assign n31833 = ~n16124 & ~n31832;
  assign n31834 = n16124 & n31713;
  assign n31835 = ~n31833 & ~n31834;
  assign n31836 = ~n17247 & n31835;
  assign n31837 = ~n31775 & ~n31836;
  assign n31838 = pi644 & n31837;
  assign n31839 = ~pi644 & n31713;
  assign n31840 = ~pi715 & ~n31839;
  assign n31841 = ~n31838 & n31840;
  assign n31842 = pi1160 & ~n31841;
  assign n31843 = ~n31774 & n31842;
  assign n31844 = pi644 & n31772;
  assign n31845 = ~pi715 & ~n31844;
  assign n31846 = ~pi644 & n31837;
  assign n31847 = pi644 & n31713;
  assign n31848 = ~n31846 & ~n31847;
  assign n31849 = pi715 & n31848;
  assign n31850 = ~pi1160 & ~n31849;
  assign n31851 = ~n31845 & n31850;
  assign n31852 = ~n31843 & ~n31851;
  assign n31853 = pi790 & ~n31852;
  assign n31854 = ~pi629 & n31753;
  assign n31855 = ~n19999 & n31832;
  assign n31856 = pi629 & n31757;
  assign n31857 = ~n31855 & ~n31856;
  assign n31858 = ~n31854 & n31857;
  assign n31859 = pi792 & ~n31858;
  assign n31860 = pi618 & n31740;
  assign n31861 = pi609 & n31738;
  assign n31862 = pi625 & n31790;
  assign n31863 = ~pi690 & ~n31788;
  assign n31864 = ~pi193 & ~n17051;
  assign n31865 = pi739 & ~n31864;
  assign n31866 = pi193 & n16998;
  assign n31867 = n31865 & ~n31866;
  assign n31868 = pi193 & n16935;
  assign n31869 = ~pi193 & n16853;
  assign n31870 = ~pi739 & ~n31869;
  assign n31871 = ~n31868 & n31870;
  assign n31872 = ~n31867 & ~n31871;
  assign n31873 = pi39 & n31872;
  assign n31874 = ~pi193 & n17067;
  assign n31875 = pi193 & n17065;
  assign n31876 = pi739 & ~n31875;
  assign n31877 = ~n31874 & n31876;
  assign n31878 = ~pi193 & ~n17061;
  assign n31879 = pi193 & ~n17058;
  assign n31880 = ~pi739 & ~n31879;
  assign n31881 = ~n31878 & n31880;
  assign n31882 = ~n31877 & ~n31881;
  assign n31883 = ~pi39 & ~n31882;
  assign n31884 = ~pi38 & ~n31883;
  assign n31885 = ~n31873 & n31884;
  assign n31886 = ~n17079 & ~n31528;
  assign n31887 = pi193 & ~n31886;
  assign n31888 = n6097 & n31887;
  assign n31889 = ~pi739 & n23427;
  assign n31890 = ~n16917 & ~n31889;
  assign n31891 = ~pi39 & ~n31890;
  assign n31892 = ~pi193 & ~n31891;
  assign n31893 = pi38 & ~n31892;
  assign n31894 = ~n31888 & n31893;
  assign n31895 = ~n31885 & ~n31894;
  assign n31896 = pi690 & n31895;
  assign n31897 = ~n31863 & ~n31896;
  assign n31898 = n10020 & n31897;
  assign n31899 = ~n31776 & ~n31898;
  assign n31900 = ~pi625 & n31899;
  assign n31901 = ~pi1153 & ~n31900;
  assign n31902 = ~n31862 & n31901;
  assign n31903 = ~pi608 & ~n31731;
  assign n31904 = ~n31902 & n31903;
  assign n31905 = ~pi625 & n31790;
  assign n31906 = pi625 & n31899;
  assign n31907 = ~n31905 & ~n31906;
  assign n31908 = pi1153 & n31907;
  assign n31909 = ~n31735 & ~n31908;
  assign n31910 = pi608 & n31909;
  assign n31911 = ~n31904 & ~n31910;
  assign n31912 = pi778 & ~n31911;
  assign n31913 = ~pi778 & n31899;
  assign n31914 = ~n31912 & ~n31913;
  assign n31915 = ~pi609 & ~n31914;
  assign n31916 = ~pi1155 & ~n31915;
  assign n31917 = ~n31861 & n31916;
  assign n31918 = ~pi660 & ~n31798;
  assign n31919 = ~n31917 & n31918;
  assign n31920 = ~pi609 & n31738;
  assign n31921 = pi609 & ~n31914;
  assign n31922 = ~n31920 & ~n31921;
  assign n31923 = pi1155 & n31922;
  assign n31924 = ~n31802 & ~n31923;
  assign n31925 = pi660 & n31924;
  assign n31926 = ~n31919 & ~n31925;
  assign n31927 = pi785 & ~n31926;
  assign n31928 = ~pi785 & ~n31914;
  assign n31929 = ~n31927 & ~n31928;
  assign n31930 = ~pi618 & ~n31929;
  assign n31931 = ~pi1154 & ~n31930;
  assign n31932 = ~n31860 & n31931;
  assign n31933 = ~pi627 & ~n31810;
  assign n31934 = ~n31932 & n31933;
  assign n31935 = ~pi618 & n31740;
  assign n31936 = pi618 & ~n31929;
  assign n31937 = ~n31935 & ~n31936;
  assign n31938 = pi1154 & n31937;
  assign n31939 = ~n31814 & ~n31938;
  assign n31940 = pi627 & n31939;
  assign n31941 = ~n31934 & ~n31940;
  assign n31942 = pi781 & ~n31941;
  assign n31943 = ~pi781 & ~n31929;
  assign n31944 = ~n31942 & ~n31943;
  assign n31945 = ~pi789 & n31944;
  assign n31946 = ~pi619 & ~n31944;
  assign n31947 = pi619 & ~n31743;
  assign n31948 = ~pi1159 & ~n31947;
  assign n31949 = ~n31946 & n31948;
  assign n31950 = ~pi648 & ~n31949;
  assign n31951 = ~n31822 & n31950;
  assign n31952 = ~pi619 & ~n31743;
  assign n31953 = pi619 & ~n31944;
  assign n31954 = ~n31952 & ~n31953;
  assign n31955 = pi1159 & n31954;
  assign n31956 = ~n31826 & ~n31955;
  assign n31957 = pi648 & n31956;
  assign n31958 = ~n31951 & ~n31957;
  assign n31959 = pi789 & n31958;
  assign n31960 = ~n31945 & ~n31959;
  assign n31961 = n17356 & n31960;
  assign n31962 = ~pi626 & ~n31829;
  assign n31963 = pi626 & ~n31713;
  assign n31964 = n17181 & ~n31963;
  assign n31965 = ~n31962 & n31964;
  assign n31966 = n17350 & n31745;
  assign n31967 = pi626 & ~n31829;
  assign n31968 = ~pi626 & ~n31713;
  assign n31969 = n17180 & ~n31968;
  assign n31970 = ~n31967 & n31969;
  assign n31971 = ~n31966 & ~n31970;
  assign n31972 = ~n31965 & n31971;
  assign n31973 = pi788 & ~n31972;
  assign n31974 = n19788 & ~n31973;
  assign n31975 = ~n31961 & n31974;
  assign n31976 = ~n31859 & ~n31975;
  assign n31977 = n19637 & ~n31976;
  assign n31978 = ~n19987 & n31835;
  assign n31979 = pi630 & n31768;
  assign n31980 = ~n31978 & ~n31979;
  assign n31981 = n17244 & ~n31763;
  assign n31982 = n31980 & ~n31981;
  assign n31983 = pi787 & ~n31982;
  assign n31984 = ~n31977 & ~n31983;
  assign n31985 = pi644 & n31842;
  assign n31986 = ~pi644 & n31850;
  assign n31987 = pi790 & ~n31986;
  assign n31988 = ~n31985 & n31987;
  assign n31989 = n31984 & ~n31988;
  assign n31990 = ~n31853 & ~n31989;
  assign n31991 = ~po1038 & ~n31990;
  assign n31992 = ~pi193 & po1038;
  assign n31993 = ~pi832 & ~n31992;
  assign n31994 = ~n31991 & n31993;
  assign po350 = ~n31712 & ~n31994;
  assign n31996 = pi194 & ~n10020;
  assign n31997 = ~pi194 & n18808;
  assign n31998 = pi194 & n23777;
  assign n31999 = ~n31997 & ~n31998;
  assign n32000 = pi748 & ~n31999;
  assign n32001 = ~pi194 & ~n16526;
  assign n32002 = ~pi748 & ~n32001;
  assign n32003 = ~n32000 & ~n32002;
  assign n32004 = n10020 & ~n32003;
  assign n32005 = ~n31996 & ~n32004;
  assign n32006 = ~n16521 & ~n32005;
  assign n32007 = ~pi194 & ~n16527;
  assign n32008 = n16521 & ~n32007;
  assign n32009 = ~n32006 & ~n32008;
  assign n32010 = ~pi785 & ~n32009;
  assign n32011 = ~n16532 & ~n32007;
  assign n32012 = pi609 & n32006;
  assign n32013 = ~n32011 & ~n32012;
  assign n32014 = pi1155 & ~n32013;
  assign n32015 = ~n16537 & ~n32007;
  assign n32016 = ~pi609 & n32006;
  assign n32017 = ~n32015 & ~n32016;
  assign n32018 = ~pi1155 & ~n32017;
  assign n32019 = ~n32014 & ~n32018;
  assign n32020 = pi785 & ~n32019;
  assign n32021 = ~n32010 & ~n32020;
  assign n32022 = ~pi781 & ~n32021;
  assign n32023 = pi618 & n32021;
  assign n32024 = ~pi618 & n32007;
  assign n32025 = pi1154 & ~n32024;
  assign n32026 = ~n32023 & n32025;
  assign n32027 = ~pi618 & n32021;
  assign n32028 = pi618 & n32007;
  assign n32029 = ~pi1154 & ~n32028;
  assign n32030 = ~n32027 & n32029;
  assign n32031 = ~n32026 & ~n32030;
  assign n32032 = pi781 & ~n32031;
  assign n32033 = ~n32022 & ~n32032;
  assign n32034 = ~pi789 & ~n32033;
  assign n32035 = pi619 & n32033;
  assign n32036 = ~pi619 & n32007;
  assign n32037 = pi1159 & ~n32036;
  assign n32038 = ~n32035 & n32037;
  assign n32039 = ~pi619 & n32033;
  assign n32040 = pi619 & n32007;
  assign n32041 = ~pi1159 & ~n32040;
  assign n32042 = ~n32039 & n32041;
  assign n32043 = ~n32038 & ~n32042;
  assign n32044 = pi789 & ~n32043;
  assign n32045 = ~n32034 & ~n32044;
  assign n32046 = ~n17355 & n32045;
  assign n32047 = n17355 & n32007;
  assign n32048 = ~n32046 & ~n32047;
  assign n32049 = ~n16124 & ~n32048;
  assign n32050 = n16124 & n32007;
  assign n32051 = ~n32049 & ~n32050;
  assign n32052 = pi647 & ~n32051;
  assign n32053 = pi628 & ~n32048;
  assign n32054 = n16593 & ~n32007;
  assign n32055 = pi194 & ~n23734;
  assign n32056 = ~pi194 & n23737;
  assign n32057 = pi730 & ~n32056;
  assign n32058 = ~pi730 & n32001;
  assign n32059 = n10020 & ~n32058;
  assign n32060 = ~n32057 & n32059;
  assign n32061 = ~n32055 & ~n32060;
  assign n32062 = ~pi778 & ~n32061;
  assign n32063 = pi625 & n32061;
  assign n32064 = pi1153 & ~n32063;
  assign n32065 = ~pi625 & n32007;
  assign n32066 = n32064 & ~n32065;
  assign n32067 = ~pi625 & n32061;
  assign n32068 = ~pi1153 & ~n32067;
  assign n32069 = pi625 & n32007;
  assign n32070 = n32068 & ~n32069;
  assign n32071 = ~n32066 & ~n32070;
  assign n32072 = pi778 & ~n32071;
  assign n32073 = ~n32062 & ~n32072;
  assign n32074 = ~n16593 & ~n32073;
  assign n32075 = ~n32054 & ~n32074;
  assign n32076 = ~n16589 & n32075;
  assign n32077 = n16589 & n32007;
  assign n32078 = ~n32076 & ~n32077;
  assign n32079 = pi619 & ~n32078;
  assign n32080 = pi618 & n32075;
  assign n32081 = pi609 & n32073;
  assign n32082 = pi625 & n32005;
  assign n32083 = ~pi730 & n32003;
  assign n32084 = ~pi194 & ~n18914;
  assign n32085 = pi748 & ~n32084;
  assign n32086 = pi194 & n18922;
  assign n32087 = n32085 & ~n32086;
  assign n32088 = pi194 & ~n23889;
  assign n32089 = ~pi194 & n18939;
  assign n32090 = ~pi748 & ~n32089;
  assign n32091 = ~n32088 & n32090;
  assign n32092 = ~n32087 & ~n32091;
  assign n32093 = pi730 & n32092;
  assign n32094 = ~n32083 & ~n32093;
  assign n32095 = n10020 & n32094;
  assign n32096 = ~n31996 & ~n32095;
  assign n32097 = ~pi625 & n32096;
  assign n32098 = ~pi1153 & ~n32097;
  assign n32099 = ~n32082 & n32098;
  assign n32100 = ~pi608 & ~n32066;
  assign n32101 = ~n32099 & n32100;
  assign n32102 = ~pi625 & n32005;
  assign n32103 = pi625 & n32096;
  assign n32104 = ~n32102 & ~n32103;
  assign n32105 = pi1153 & n32104;
  assign n32106 = ~n32070 & ~n32105;
  assign n32107 = pi608 & n32106;
  assign n32108 = ~n32101 & ~n32107;
  assign n32109 = pi778 & ~n32108;
  assign n32110 = ~pi778 & n32096;
  assign n32111 = ~n32109 & ~n32110;
  assign n32112 = ~pi609 & ~n32111;
  assign n32113 = ~pi1155 & ~n32112;
  assign n32114 = ~n32081 & n32113;
  assign n32115 = ~pi660 & ~n32014;
  assign n32116 = ~n32114 & n32115;
  assign n32117 = ~pi609 & n32073;
  assign n32118 = pi609 & ~n32111;
  assign n32119 = ~n32117 & ~n32118;
  assign n32120 = pi1155 & n32119;
  assign n32121 = ~n32018 & ~n32120;
  assign n32122 = pi660 & n32121;
  assign n32123 = ~n32116 & ~n32122;
  assign n32124 = pi785 & ~n32123;
  assign n32125 = ~pi785 & ~n32111;
  assign n32126 = ~n32124 & ~n32125;
  assign n32127 = ~pi618 & ~n32126;
  assign n32128 = ~pi1154 & ~n32127;
  assign n32129 = ~n32080 & n32128;
  assign n32130 = ~pi627 & ~n32026;
  assign n32131 = ~n32129 & n32130;
  assign n32132 = ~pi618 & n32075;
  assign n32133 = pi618 & ~n32126;
  assign n32134 = ~n32132 & ~n32133;
  assign n32135 = pi1154 & n32134;
  assign n32136 = ~n32030 & ~n32135;
  assign n32137 = pi627 & n32136;
  assign n32138 = ~n32131 & ~n32137;
  assign n32139 = pi781 & ~n32138;
  assign n32140 = ~pi781 & ~n32126;
  assign n32141 = ~n32139 & ~n32140;
  assign n32142 = ~pi619 & ~n32141;
  assign n32143 = ~pi1159 & ~n32142;
  assign n32144 = ~n32079 & n32143;
  assign n32145 = ~pi648 & ~n32038;
  assign n32146 = ~n32144 & n32145;
  assign n32147 = ~pi619 & ~n32078;
  assign n32148 = pi619 & ~n32141;
  assign n32149 = ~n32147 & ~n32148;
  assign n32150 = pi1159 & n32149;
  assign n32151 = ~n32042 & ~n32150;
  assign n32152 = pi648 & n32151;
  assign n32153 = ~n32146 & ~n32152;
  assign n32154 = pi789 & ~n32153;
  assign n32155 = ~pi789 & ~n32141;
  assign n32156 = ~n32154 & ~n32155;
  assign n32157 = ~pi788 & n32156;
  assign n32158 = pi626 & n32156;
  assign n32159 = n17159 & ~n32007;
  assign n32160 = ~n17159 & n32078;
  assign n32161 = ~n32159 & ~n32160;
  assign n32162 = ~pi626 & ~n32161;
  assign n32163 = pi641 & ~n32162;
  assign n32164 = ~n32158 & n32163;
  assign n32165 = pi626 & ~n32045;
  assign n32166 = ~pi626 & ~n32007;
  assign n32167 = ~pi641 & ~n32166;
  assign n32168 = ~n32165 & n32167;
  assign n32169 = pi1158 & ~n32168;
  assign n32170 = ~n32164 & n32169;
  assign n32171 = pi626 & ~n32007;
  assign n32172 = ~pi626 & ~n32045;
  assign n32173 = pi641 & ~n32172;
  assign n32174 = ~n32171 & n32173;
  assign n32175 = pi626 & ~n32161;
  assign n32176 = ~pi626 & n32156;
  assign n32177 = ~pi641 & ~n32176;
  assign n32178 = ~n32175 & n32177;
  assign n32179 = ~pi1158 & ~n32178;
  assign n32180 = ~n32174 & n32179;
  assign n32181 = ~n32170 & ~n32180;
  assign n32182 = pi788 & ~n32181;
  assign n32183 = ~n32157 & ~n32182;
  assign n32184 = ~pi628 & n32183;
  assign n32185 = ~pi1156 & ~n32184;
  assign n32186 = ~n32053 & n32185;
  assign n32187 = ~n17183 & n32161;
  assign n32188 = n17183 & n32007;
  assign n32189 = ~n32187 & ~n32188;
  assign n32190 = pi628 & ~n32189;
  assign n32191 = pi1156 & ~n32190;
  assign n32192 = ~pi628 & n32007;
  assign n32193 = n32191 & ~n32192;
  assign n32194 = ~pi629 & ~n32193;
  assign n32195 = ~n32186 & n32194;
  assign n32196 = ~pi628 & ~n32189;
  assign n32197 = pi628 & n32007;
  assign n32198 = ~pi1156 & ~n32197;
  assign n32199 = ~n32196 & n32198;
  assign n32200 = ~pi628 & ~n32048;
  assign n32201 = pi628 & n32183;
  assign n32202 = ~n32200 & ~n32201;
  assign n32203 = pi1156 & n32202;
  assign n32204 = ~n32199 & ~n32203;
  assign n32205 = pi629 & n32204;
  assign n32206 = ~n32195 & ~n32205;
  assign n32207 = pi792 & ~n32206;
  assign n32208 = ~pi792 & n32183;
  assign n32209 = ~n32207 & ~n32208;
  assign n32210 = ~pi647 & ~n32209;
  assign n32211 = ~pi1157 & ~n32210;
  assign n32212 = ~n32052 & n32211;
  assign n32213 = ~pi792 & n32189;
  assign n32214 = ~n32193 & ~n32199;
  assign n32215 = pi792 & ~n32214;
  assign n32216 = ~n32213 & ~n32215;
  assign n32217 = pi647 & n32216;
  assign n32218 = pi1157 & ~n32217;
  assign n32219 = ~pi647 & n32007;
  assign n32220 = n32218 & ~n32219;
  assign n32221 = ~pi630 & ~n32220;
  assign n32222 = ~n32212 & n32221;
  assign n32223 = ~pi647 & n32216;
  assign n32224 = pi647 & n32007;
  assign n32225 = ~pi1157 & ~n32224;
  assign n32226 = ~n32223 & n32225;
  assign n32227 = ~pi647 & ~n32051;
  assign n32228 = pi647 & ~n32209;
  assign n32229 = ~n32227 & ~n32228;
  assign n32230 = pi1157 & n32229;
  assign n32231 = ~n32226 & ~n32230;
  assign n32232 = pi630 & n32231;
  assign n32233 = ~n32222 & ~n32232;
  assign n32234 = pi787 & ~n32233;
  assign n32235 = ~pi787 & ~n32209;
  assign n32236 = ~n32234 & ~n32235;
  assign n32237 = ~pi790 & n32236;
  assign n32238 = pi644 & ~n32236;
  assign n32239 = ~pi787 & ~n32216;
  assign n32240 = ~n32220 & ~n32226;
  assign n32241 = pi787 & ~n32240;
  assign n32242 = ~n32239 & ~n32241;
  assign n32243 = ~pi644 & n32242;
  assign n32244 = pi715 & ~n32243;
  assign n32245 = ~n32238 & n32244;
  assign n32246 = ~pi644 & n32007;
  assign n32247 = n17247 & ~n32007;
  assign n32248 = ~n17247 & n32051;
  assign n32249 = ~n32247 & ~n32248;
  assign n32250 = pi644 & n32249;
  assign n32251 = ~pi715 & ~n32250;
  assign n32252 = ~n32246 & n32251;
  assign n32253 = ~n32245 & ~n32252;
  assign n32254 = pi1160 & n32253;
  assign n32255 = ~pi644 & n32249;
  assign n32256 = pi715 & ~n32255;
  assign n32257 = pi644 & n32007;
  assign n32258 = n32256 & ~n32257;
  assign n32259 = pi644 & n32242;
  assign n32260 = ~pi644 & ~n32236;
  assign n32261 = ~pi715 & ~n32260;
  assign n32262 = ~n32259 & n32261;
  assign n32263 = ~n32258 & ~n32262;
  assign n32264 = ~pi1160 & n32263;
  assign n32265 = ~n32254 & ~n32264;
  assign n32266 = pi790 & n32265;
  assign n32267 = ~n32237 & ~n32266;
  assign n32268 = ~po1038 & n32267;
  assign n32269 = ~pi194 & po1038;
  assign n32270 = ~pi832 & ~n32269;
  assign n32271 = ~n32268 & n32270;
  assign n32272 = ~pi194 & ~n2934;
  assign n32273 = pi748 & n16510;
  assign n32274 = ~n32272 & ~n32273;
  assign n32275 = ~n17273 & ~n32274;
  assign n32276 = ~pi785 & ~n32275;
  assign n32277 = ~n17279 & ~n32274;
  assign n32278 = pi1155 & ~n32277;
  assign n32279 = ~n17282 & n32275;
  assign n32280 = ~pi1155 & ~n32279;
  assign n32281 = ~n32278 & ~n32280;
  assign n32282 = pi785 & ~n32281;
  assign n32283 = ~n32276 & ~n32282;
  assign n32284 = ~pi781 & ~n32283;
  assign n32285 = ~n17289 & n32283;
  assign n32286 = pi1154 & ~n32285;
  assign n32287 = ~n17292 & n32283;
  assign n32288 = ~pi1154 & ~n32287;
  assign n32289 = ~n32286 & ~n32288;
  assign n32290 = pi781 & ~n32289;
  assign n32291 = ~n32284 & ~n32290;
  assign n32292 = ~pi789 & ~n32291;
  assign n32293 = pi619 & n32291;
  assign n32294 = ~pi619 & n32272;
  assign n32295 = pi1159 & ~n32294;
  assign n32296 = ~n32293 & n32295;
  assign n32297 = ~pi619 & n32291;
  assign n32298 = pi619 & n32272;
  assign n32299 = ~pi1159 & ~n32298;
  assign n32300 = ~n32297 & n32299;
  assign n32301 = ~n32296 & ~n32300;
  assign n32302 = pi789 & ~n32301;
  assign n32303 = ~n32292 & ~n32302;
  assign n32304 = ~n17355 & n32303;
  assign n32305 = n17355 & n32272;
  assign n32306 = ~n32304 & ~n32305;
  assign n32307 = ~n16124 & ~n32306;
  assign n32308 = n16124 & n32272;
  assign n32309 = ~n32307 & ~n32308;
  assign n32310 = ~n19987 & n32309;
  assign n32311 = pi730 & n16742;
  assign n32312 = ~n32272 & ~n32311;
  assign n32313 = ~pi778 & n32312;
  assign n32314 = ~pi625 & n32311;
  assign n32315 = ~n32312 & ~n32314;
  assign n32316 = pi1153 & ~n32315;
  assign n32317 = ~pi1153 & ~n32272;
  assign n32318 = ~n32314 & n32317;
  assign n32319 = ~n32316 & ~n32318;
  assign n32320 = pi778 & ~n32319;
  assign n32321 = ~n32313 & ~n32320;
  assign n32322 = ~n17338 & n32321;
  assign n32323 = ~n17340 & n32322;
  assign n32324 = ~n17342 & n32323;
  assign n32325 = ~n17425 & n32324;
  assign n32326 = ~n17452 & n32325;
  assign n32327 = ~pi647 & n32326;
  assign n32328 = pi647 & n32272;
  assign n32329 = ~pi1157 & ~n32328;
  assign n32330 = ~n32327 & n32329;
  assign n32331 = ~pi647 & n32272;
  assign n32332 = pi647 & n32326;
  assign n32333 = pi1157 & ~n32332;
  assign n32334 = ~n32331 & n32333;
  assign n32335 = ~n32330 & ~n32334;
  assign n32336 = ~n17246 & ~n32335;
  assign n32337 = ~n32310 & ~n32336;
  assign n32338 = pi787 & ~n32337;
  assign n32339 = ~pi626 & ~n32303;
  assign n32340 = pi626 & ~n32272;
  assign n32341 = n17181 & ~n32340;
  assign n32342 = ~n32339 & n32341;
  assign n32343 = n17350 & n32324;
  assign n32344 = pi626 & ~n32303;
  assign n32345 = ~pi626 & ~n32272;
  assign n32346 = n17180 & ~n32345;
  assign n32347 = ~n32344 & n32346;
  assign n32348 = ~n32343 & ~n32347;
  assign n32349 = ~n32342 & n32348;
  assign n32350 = pi788 & ~n32349;
  assign n32351 = pi618 & n32322;
  assign n32352 = pi609 & n32321;
  assign n32353 = ~n16393 & ~n32312;
  assign n32354 = pi625 & n32353;
  assign n32355 = n32274 & ~n32353;
  assign n32356 = ~n32354 & ~n32355;
  assign n32357 = n32317 & ~n32356;
  assign n32358 = ~pi608 & ~n32316;
  assign n32359 = ~n32357 & n32358;
  assign n32360 = pi1153 & ~n32354;
  assign n32361 = n32274 & n32360;
  assign n32362 = ~n32318 & ~n32361;
  assign n32363 = pi608 & n32362;
  assign n32364 = ~n32359 & ~n32363;
  assign n32365 = pi778 & ~n32364;
  assign n32366 = ~pi778 & ~n32355;
  assign n32367 = ~n32365 & ~n32366;
  assign n32368 = ~pi609 & ~n32367;
  assign n32369 = ~pi1155 & ~n32368;
  assign n32370 = ~n32352 & n32369;
  assign n32371 = ~pi660 & ~n32278;
  assign n32372 = ~n32370 & n32371;
  assign n32373 = ~pi609 & n32321;
  assign n32374 = pi609 & ~n32367;
  assign n32375 = ~n32373 & ~n32374;
  assign n32376 = pi1155 & n32375;
  assign n32377 = ~n32280 & ~n32376;
  assign n32378 = pi660 & n32377;
  assign n32379 = ~n32372 & ~n32378;
  assign n32380 = pi785 & ~n32379;
  assign n32381 = ~pi785 & ~n32367;
  assign n32382 = ~n32380 & ~n32381;
  assign n32383 = ~pi618 & ~n32382;
  assign n32384 = ~pi1154 & ~n32383;
  assign n32385 = ~n32351 & n32384;
  assign n32386 = ~pi627 & ~n32286;
  assign n32387 = ~n32385 & n32386;
  assign n32388 = ~pi618 & n32322;
  assign n32389 = pi618 & ~n32382;
  assign n32390 = ~n32388 & ~n32389;
  assign n32391 = pi1154 & n32390;
  assign n32392 = ~n32288 & ~n32391;
  assign n32393 = pi627 & n32392;
  assign n32394 = ~n32387 & ~n32393;
  assign n32395 = pi781 & ~n32394;
  assign n32396 = ~pi781 & ~n32382;
  assign n32397 = ~n32395 & ~n32396;
  assign n32398 = ~pi619 & ~n32397;
  assign n32399 = pi619 & n32323;
  assign n32400 = ~pi1159 & ~n32399;
  assign n32401 = ~n32398 & n32400;
  assign n32402 = ~pi648 & ~n32401;
  assign n32403 = ~n32296 & n32402;
  assign n32404 = ~pi619 & n32323;
  assign n32405 = pi619 & ~n32397;
  assign n32406 = ~n32404 & ~n32405;
  assign n32407 = pi1159 & n32406;
  assign n32408 = ~n32300 & ~n32407;
  assign n32409 = pi648 & n32408;
  assign n32410 = ~n32403 & ~n32409;
  assign n32411 = pi789 & n32410;
  assign n32412 = ~pi789 & n32397;
  assign n32413 = n17356 & ~n32412;
  assign n32414 = ~n32411 & n32413;
  assign n32415 = ~n32350 & ~n32414;
  assign n32416 = n19788 & ~n32415;
  assign n32417 = n20275 & n32325;
  assign n32418 = n17449 & ~n32306;
  assign n32419 = ~pi629 & ~n32418;
  assign n32420 = ~n32417 & n32419;
  assign n32421 = n17448 & ~n32306;
  assign n32422 = n20281 & n32325;
  assign n32423 = pi629 & ~n32422;
  assign n32424 = ~n32421 & n32423;
  assign n32425 = ~n32420 & ~n32424;
  assign n32426 = pi792 & n32425;
  assign n32427 = n19637 & ~n32426;
  assign n32428 = ~n32416 & n32427;
  assign n32429 = ~n32338 & ~n32428;
  assign n32430 = pi644 & n32429;
  assign n32431 = ~pi787 & ~n32326;
  assign n32432 = pi787 & ~n32335;
  assign n32433 = ~n32431 & ~n32432;
  assign n32434 = ~pi644 & n32433;
  assign n32435 = pi715 & ~n32434;
  assign n32436 = ~n32430 & n32435;
  assign n32437 = ~n17247 & ~n32309;
  assign n32438 = n17247 & n32272;
  assign n32439 = ~n32437 & ~n32438;
  assign n32440 = pi644 & ~n32439;
  assign n32441 = ~pi644 & n32272;
  assign n32442 = ~pi715 & ~n32441;
  assign n32443 = ~n32440 & n32442;
  assign n32444 = pi1160 & ~n32443;
  assign n32445 = ~n32436 & n32444;
  assign n32446 = ~pi644 & ~n32439;
  assign n32447 = pi715 & ~n32446;
  assign n32448 = pi644 & n32272;
  assign n32449 = n32447 & ~n32448;
  assign n32450 = pi644 & n32433;
  assign n32451 = ~pi644 & n32429;
  assign n32452 = ~pi715 & ~n32451;
  assign n32453 = ~n32450 & n32452;
  assign n32454 = ~pi1160 & ~n32453;
  assign n32455 = ~n32449 & n32454;
  assign n32456 = ~n32445 & ~n32455;
  assign n32457 = pi790 & ~n32456;
  assign n32458 = ~pi790 & n32429;
  assign n32459 = pi832 & ~n32458;
  assign n32460 = ~n32457 & n32459;
  assign po351 = ~n32271 & ~n32460;
  assign n32462 = n11264 & ~n15665;
  assign n32463 = ~pi39 & ~n32462;
  assign n32464 = n10024 & ~n32463;
  assign n32465 = ~pi138 & n15984;
  assign n32466 = ~pi196 & n32465;
  assign n32467 = pi195 & ~n32466;
  assign n32468 = ~n6191 & n15663;
  assign n32469 = ~pi192 & n11258;
  assign n32470 = n15662 & ~n15990;
  assign n32471 = ~n11260 & ~n32470;
  assign n32472 = ~n32469 & n32471;
  assign n32473 = ~n32468 & n32472;
  assign n32474 = pi232 & ~n32473;
  assign n32475 = ~n15985 & ~n32474;
  assign n32476 = pi39 & ~n32475;
  assign n32477 = ~n32467 & ~n32476;
  assign n32478 = n32464 & n32477;
  assign n32479 = n15662 & ~n16012;
  assign n32480 = ~n9643 & n15688;
  assign n32481 = ~n9294 & ~n15653;
  assign n32482 = pi171 & n13533;
  assign n32483 = ~n32481 & ~n32482;
  assign n32484 = pi299 & ~n32483;
  assign n32485 = pi232 & ~n32484;
  assign n32486 = ~n32480 & n32485;
  assign n32487 = ~n32479 & n32486;
  assign n32488 = n16010 & ~n32487;
  assign n32489 = pi192 & n16040;
  assign n32490 = ~pi192 & n16026;
  assign n32491 = ~pi171 & n8990;
  assign n32492 = ~n16034 & ~n32491;
  assign n32493 = n8959 & ~n32492;
  assign n32494 = n8961 & ~n32493;
  assign n32495 = ~n32490 & ~n32494;
  assign n32496 = ~n32489 & n32495;
  assign n32497 = pi232 & ~n32496;
  assign n32498 = ~n16032 & ~n32497;
  assign n32499 = pi39 & ~n32498;
  assign n32500 = ~n32488 & ~n32499;
  assign n32501 = n2614 & n32500;
  assign n32502 = ~pi87 & ~n32501;
  assign n32503 = n16005 & ~n32502;
  assign n32504 = ~pi92 & ~n32503;
  assign n32505 = n16004 & ~n32504;
  assign n32506 = ~pi55 & ~n32505;
  assign n32507 = ~n16055 & ~n32506;
  assign n32508 = n2531 & ~n32507;
  assign n32509 = n9564 & ~n32508;
  assign n32510 = n32467 & n32509;
  assign po352 = n32478 | n32510;
  assign n32512 = ~pi170 & n8990;
  assign n32513 = ~n16034 & ~n32512;
  assign n32514 = n8959 & ~n32513;
  assign n32515 = n8961 & ~n32514;
  assign n32516 = ~n16026 & ~n32515;
  assign n32517 = pi232 & ~n32516;
  assign n32518 = ~n16032 & ~n32517;
  assign n32519 = pi232 & n16040;
  assign n32520 = n32518 & ~n32519;
  assign n32521 = pi39 & ~n32520;
  assign n32522 = ~pi38 & pi194;
  assign n32523 = ~n32521 & n32522;
  assign n32524 = pi39 & ~n32518;
  assign n32525 = ~pi38 & ~pi194;
  assign n32526 = ~n32524 & n32525;
  assign n32527 = ~n32523 & ~n32526;
  assign n32528 = ~n16010 & ~n32527;
  assign n32529 = ~pi299 & ~n16012;
  assign n32530 = n32523 & ~n32529;
  assign n32531 = ~n16006 & n32526;
  assign n32532 = ~n32530 & ~n32531;
  assign n32533 = ~n9294 & ~n15766;
  assign n32534 = pi170 & n13533;
  assign n32535 = ~n32533 & ~n32534;
  assign n32536 = pi299 & ~n32535;
  assign n32537 = pi232 & ~n32536;
  assign n32538 = ~n32532 & n32537;
  assign n32539 = ~n32528 & ~n32538;
  assign n32540 = ~pi100 & ~n32539;
  assign n32541 = ~pi87 & ~n32540;
  assign n32542 = n16005 & ~n32541;
  assign n32543 = ~pi92 & ~n32542;
  assign n32544 = n16004 & ~n32543;
  assign n32545 = ~pi55 & ~n32544;
  assign n32546 = ~n16055 & ~n32545;
  assign n32547 = n2531 & ~n32546;
  assign n32548 = n9564 & ~n32547;
  assign n32549 = pi196 & ~n32548;
  assign n32550 = ~pi170 & n9393;
  assign n32551 = ~n15989 & ~n32550;
  assign n32552 = n12812 & ~n32551;
  assign n32553 = ~pi299 & n15990;
  assign n32554 = ~n32552 & ~n32553;
  assign n32555 = pi232 & n32554;
  assign n32556 = ~n15985 & ~n32555;
  assign n32557 = pi299 & ~n32556;
  assign n32558 = ~n11258 & ~n32557;
  assign n32559 = pi39 & ~n32558;
  assign n32560 = n11264 & ~n15767;
  assign n32561 = ~pi39 & ~n32560;
  assign n32562 = ~pi38 & ~n32561;
  assign n32563 = ~n32559 & n32562;
  assign n32564 = ~pi194 & ~n32563;
  assign n32565 = pi39 & ~n32556;
  assign n32566 = n11264 & n15780;
  assign n32567 = ~pi39 & ~n32566;
  assign n32568 = ~pi38 & ~n32567;
  assign n32569 = ~n32565 & n32568;
  assign n32570 = pi194 & ~n32569;
  assign n32571 = n10021 & ~n32570;
  assign n32572 = ~n32564 & n32571;
  assign n32573 = ~pi196 & ~n32572;
  assign n32574 = ~n32465 & ~n32573;
  assign n32575 = ~n32549 & n32574;
  assign n32576 = pi195 & ~pi196;
  assign n32577 = ~n32548 & n32576;
  assign n32578 = ~n32572 & ~n32576;
  assign n32579 = n32465 & ~n32578;
  assign n32580 = ~n32577 & n32579;
  assign po353 = n32575 | n32580;
  assign n32582 = ~pi767 & pi947;
  assign n32583 = ~pi698 & n20323;
  assign n32584 = ~n32582 & ~n32583;
  assign n32585 = n2934 & ~n32584;
  assign n32586 = ~pi197 & ~n2934;
  assign n32587 = pi832 & ~n32586;
  assign n32588 = ~n32585 & n32587;
  assign n32589 = pi197 & ~n16524;
  assign n32590 = n16508 & ~n32582;
  assign n32591 = pi38 & ~n32590;
  assign n32592 = ~n32589 & n32591;
  assign n32593 = ~pi197 & ~n16333;
  assign n32594 = n20514 & ~n32593;
  assign n32595 = pi197 & ~n20573;
  assign n32596 = ~pi197 & ~n20497;
  assign n32597 = ~n32595 & ~n32596;
  assign n32598 = pi299 & n32597;
  assign n32599 = ~pi767 & ~n32598;
  assign n32600 = ~n32594 & n32599;
  assign n32601 = ~pi197 & pi767;
  assign n32602 = ~n16355 & n32601;
  assign n32603 = pi39 & ~n32602;
  assign n32604 = ~n32600 & n32603;
  assign n32605 = ~pi197 & ~n16201;
  assign n32606 = ~pi39 & ~n32605;
  assign n32607 = n16201 & n32582;
  assign n32608 = n32606 & ~n32607;
  assign n32609 = ~pi38 & ~n32608;
  assign n32610 = ~n32604 & n32609;
  assign n32611 = ~n32592 & ~n32610;
  assign n32612 = pi698 & ~n32611;
  assign n32613 = ~n20425 & n32608;
  assign n32614 = n20422 & ~n32593;
  assign n32615 = ~pi197 & n20439;
  assign n32616 = pi197 & n20419;
  assign n32617 = pi299 & ~n32616;
  assign n32618 = ~n32615 & n32617;
  assign n32619 = pi767 & ~n32618;
  assign n32620 = ~n32614 & n32619;
  assign n32621 = pi197 & n20478;
  assign n32622 = ~pi197 & n20467;
  assign n32623 = ~pi767 & ~n32622;
  assign n32624 = ~n32621 & n32623;
  assign n32625 = pi39 & ~n32624;
  assign n32626 = ~n32620 & n32625;
  assign n32627 = ~n32613 & ~n32626;
  assign n32628 = ~pi38 & ~n32627;
  assign n32629 = pi197 & ~n16508;
  assign n32630 = ~n32590 & ~n32629;
  assign n32631 = n20453 & ~n32630;
  assign n32632 = ~pi698 & ~n32631;
  assign n32633 = ~n32628 & n32632;
  assign n32634 = ~n32612 & ~n32633;
  assign n32635 = n10021 & ~n32634;
  assign n32636 = ~pi197 & ~n10021;
  assign n32637 = ~pi832 & ~n32636;
  assign n32638 = ~n32635 & n32637;
  assign po354 = ~n32588 & ~n32638;
  assign n32640 = n2532 & ~n16201;
  assign n32641 = n18119 & ~n32640;
  assign n32642 = pi198 & ~n32641;
  assign n32643 = pi198 & ~n16227;
  assign n32644 = pi198 & ~n16207;
  assign n32645 = ~po1101 & ~n32644;
  assign n32646 = n32643 & ~n32645;
  assign n32647 = pi198 & n16263;
  assign n32648 = ~n6198 & n32647;
  assign n32649 = ~n32646 & ~n32648;
  assign n32650 = pi215 & ~n32649;
  assign n32651 = n2527 & ~n32644;
  assign n32652 = pi198 & ~n16301;
  assign n32653 = po1101 & ~n32652;
  assign n32654 = ~n32645 & ~n32653;
  assign n32655 = n6198 & n32654;
  assign n32656 = pi198 & ~n16297;
  assign n32657 = ~n6198 & n32656;
  assign n32658 = ~n2527 & ~n32657;
  assign n32659 = ~n32655 & n32658;
  assign n32660 = ~pi215 & ~n32659;
  assign n32661 = ~n32651 & n32660;
  assign n32662 = ~n32650 & ~n32661;
  assign n32663 = pi299 & n32662;
  assign n32664 = pi39 & ~n32663;
  assign n32665 = ~n6236 & n32647;
  assign n32666 = ~n32646 & ~n32665;
  assign n32667 = pi223 & ~n32666;
  assign n32668 = n2607 & ~n32644;
  assign n32669 = n6236 & n32654;
  assign n32670 = ~n6236 & n32656;
  assign n32671 = ~n2607 & ~n32670;
  assign n32672 = ~n32669 & n32671;
  assign n32673 = ~pi223 & ~n32672;
  assign n32674 = ~n32668 & n32673;
  assign n32675 = ~pi299 & ~n32674;
  assign n32676 = ~n32667 & n32675;
  assign n32677 = n32664 & ~n32676;
  assign n32678 = n2575 & n32677;
  assign n32679 = ~n32642 & ~n32678;
  assign n32680 = n16124 & ~n32679;
  assign n32681 = pi198 & ~n10020;
  assign n32682 = pi603 & pi633;
  assign n32683 = pi198 & ~n16195;
  assign n32684 = ~n32682 & ~n32683;
  assign n32685 = ~pi198 & ~n16457;
  assign n32686 = pi198 & n16363;
  assign n32687 = ~n32685 & ~n32686;
  assign n32688 = n32682 & ~n32687;
  assign n32689 = ~n32684 & ~n32688;
  assign n32690 = pi299 & n32689;
  assign n32691 = ~n16368 & ~n16372;
  assign n32692 = pi633 & ~n32691;
  assign n32693 = ~n16198 & ~n32692;
  assign n32694 = ~n16377 & ~n32693;
  assign n32695 = ~pi299 & n32694;
  assign n32696 = ~pi39 & ~n32695;
  assign n32697 = ~n32690 & n32696;
  assign n32698 = pi633 & n16207;
  assign n32699 = ~n16382 & n32698;
  assign n32700 = ~n32644 & ~n32699;
  assign n32701 = pi603 & ~n32700;
  assign n32702 = ~pi603 & n32644;
  assign n32703 = ~n32701 & ~n32702;
  assign n32704 = ~n16392 & n32703;
  assign n32705 = ~n16224 & n32699;
  assign n32706 = n6190 & ~n32700;
  assign n32707 = ~n32705 & ~n32706;
  assign n32708 = ~n32643 & n32707;
  assign n32709 = pi603 & ~n32708;
  assign n32710 = ~n32702 & ~n32709;
  assign n32711 = n16392 & n32710;
  assign n32712 = ~n32704 & ~n32711;
  assign n32713 = ~n6188 & n32712;
  assign n32714 = ~n32643 & ~n32709;
  assign n32715 = n6188 & ~n32714;
  assign n32716 = ~n32713 & ~n32715;
  assign n32717 = n6198 & n32716;
  assign n32718 = pi633 & n16482;
  assign n32719 = ~n32647 & ~n32718;
  assign n32720 = ~n6188 & ~n32719;
  assign n32721 = pi198 & n16224;
  assign n32722 = ~n32705 & ~n32721;
  assign n32723 = n16427 & ~n32722;
  assign n32724 = ~n32720 & ~n32723;
  assign n32725 = ~n6198 & n32724;
  assign n32726 = pi215 & ~n32725;
  assign n32727 = ~n32717 & n32726;
  assign n32728 = ~pi603 & n16292;
  assign n32729 = pi198 & n32728;
  assign n32730 = pi198 & n16289;
  assign n32731 = pi633 & n16808;
  assign n32732 = ~n32730 & ~n32731;
  assign n32733 = pi603 & ~n32732;
  assign n32734 = n16392 & n32733;
  assign n32735 = n6190 & n32732;
  assign n32736 = ~n6190 & n32700;
  assign n32737 = pi603 & ~n32736;
  assign n32738 = ~n16392 & n32737;
  assign n32739 = ~n32735 & n32738;
  assign n32740 = ~n32734 & ~n32739;
  assign n32741 = ~n32729 & n32740;
  assign n32742 = ~n6188 & n32741;
  assign n32743 = n6188 & ~n32730;
  assign n32744 = ~n32733 & n32743;
  assign n32745 = ~n32742 & ~n32744;
  assign n32746 = ~n6198 & n32745;
  assign n32747 = pi642 & ~n32701;
  assign n32748 = ~n6190 & ~n32732;
  assign n32749 = ~n32706 & ~n32748;
  assign n32750 = pi603 & ~n32749;
  assign n32751 = ~pi642 & ~n32750;
  assign n32752 = ~n32747 & ~n32751;
  assign n32753 = n6184 & n32752;
  assign n32754 = ~n6184 & n32701;
  assign n32755 = ~n32702 & ~n32754;
  assign n32756 = ~n32753 & n32755;
  assign n32757 = ~n6188 & n32756;
  assign n32758 = ~pi603 & n32652;
  assign n32759 = n6188 & ~n32750;
  assign n32760 = ~n32758 & n32759;
  assign n32761 = ~n32757 & ~n32760;
  assign n32762 = n6198 & n32761;
  assign n32763 = ~n2527 & ~n32762;
  assign n32764 = ~n32746 & n32763;
  assign n32765 = n2527 & n32703;
  assign n32766 = ~pi215 & ~n32765;
  assign n32767 = ~n32764 & n32766;
  assign n32768 = ~n32727 & ~n32767;
  assign n32769 = pi299 & ~n32768;
  assign n32770 = n6236 & n32716;
  assign n32771 = ~n6236 & n32724;
  assign n32772 = pi223 & ~n32771;
  assign n32773 = ~n32770 & n32772;
  assign n32774 = ~n6236 & n32745;
  assign n32775 = n6236 & n32761;
  assign n32776 = ~n2607 & ~n32775;
  assign n32777 = ~n32774 & n32776;
  assign n32778 = n2607 & n32703;
  assign n32779 = ~pi223 & ~n32778;
  assign n32780 = ~n32777 & n32779;
  assign n32781 = ~n32773 & ~n32780;
  assign n32782 = ~pi299 & ~n32781;
  assign n32783 = pi39 & ~n32782;
  assign n32784 = ~n32769 & n32783;
  assign n32785 = ~n32697 & ~n32784;
  assign n32786 = ~pi38 & ~n32785;
  assign n32787 = pi39 & pi198;
  assign n32788 = pi38 & ~n32787;
  assign n32789 = pi198 & ~n16212;
  assign n32790 = pi633 & n16393;
  assign n32791 = n16212 & n32790;
  assign n32792 = ~n32789 & ~n32791;
  assign n32793 = ~pi39 & ~n32792;
  assign n32794 = n32788 & ~n32793;
  assign n32795 = ~n32786 & ~n32794;
  assign n32796 = n10020 & n32795;
  assign n32797 = ~n32681 & ~n32796;
  assign n32798 = ~n16521 & ~n32797;
  assign n32799 = n16521 & ~n32679;
  assign n32800 = ~n32798 & ~n32799;
  assign n32801 = ~pi785 & ~n32800;
  assign n32802 = ~n16532 & ~n32679;
  assign n32803 = pi609 & n32798;
  assign n32804 = ~n32802 & ~n32803;
  assign n32805 = pi1155 & ~n32804;
  assign n32806 = ~n16537 & ~n32679;
  assign n32807 = ~pi609 & n32798;
  assign n32808 = ~n32806 & ~n32807;
  assign n32809 = ~pi1155 & ~n32808;
  assign n32810 = ~n32805 & ~n32809;
  assign n32811 = pi785 & ~n32810;
  assign n32812 = ~n32801 & ~n32811;
  assign n32813 = ~pi781 & ~n32812;
  assign n32814 = pi618 & n32812;
  assign n32815 = ~pi618 & n32679;
  assign n32816 = pi1154 & ~n32815;
  assign n32817 = ~n32814 & n32816;
  assign n32818 = ~pi618 & n32812;
  assign n32819 = pi618 & n32679;
  assign n32820 = ~pi1154 & ~n32819;
  assign n32821 = ~n32818 & n32820;
  assign n32822 = ~n32817 & ~n32821;
  assign n32823 = pi781 & ~n32822;
  assign n32824 = ~n32813 & ~n32823;
  assign n32825 = ~pi789 & ~n32824;
  assign n32826 = pi619 & n32824;
  assign n32827 = ~pi619 & n32679;
  assign n32828 = pi1159 & ~n32827;
  assign n32829 = ~n32826 & n32828;
  assign n32830 = ~pi619 & n32824;
  assign n32831 = pi619 & n32679;
  assign n32832 = ~pi1159 & ~n32831;
  assign n32833 = ~n32830 & n32832;
  assign n32834 = ~n32829 & ~n32833;
  assign n32835 = pi789 & ~n32834;
  assign n32836 = ~n32825 & ~n32835;
  assign n32837 = ~n17355 & n32836;
  assign n32838 = n17355 & n32679;
  assign n32839 = ~n32837 & ~n32838;
  assign n32840 = ~n16124 & n32839;
  assign n32841 = ~n32680 & ~n32840;
  assign n32842 = ~n19987 & ~n32841;
  assign n32843 = ~n17159 & ~n17183;
  assign n32844 = n32679 & ~n32843;
  assign n32845 = n16589 & ~n32679;
  assign n32846 = ~n16600 & ~n32644;
  assign n32847 = pi634 & ~n32846;
  assign n32848 = ~n32644 & ~n32847;
  assign n32849 = ~n6190 & n32848;
  assign n32850 = pi634 & ~n16224;
  assign n32851 = n16600 & n32850;
  assign n32852 = ~n32721 & ~n32851;
  assign n32853 = n6190 & n32852;
  assign n32854 = ~n32849 & ~n32853;
  assign n32855 = n6190 & ~n32848;
  assign n32856 = ~n6190 & ~n32852;
  assign n32857 = ~n32855 & ~n32856;
  assign n32858 = n6185 & n32857;
  assign n32859 = n32854 & ~n32858;
  assign n32860 = ~n32647 & ~n32859;
  assign n32861 = n16774 & ~n32860;
  assign n32862 = ~pi680 & n32647;
  assign n32863 = n6188 & ~n32852;
  assign n32864 = ~n32862 & ~n32863;
  assign n32865 = ~n32861 & n32864;
  assign n32866 = ~n6236 & n32865;
  assign n32867 = pi223 & ~n32866;
  assign n32868 = n32643 & n32862;
  assign n32869 = n6188 & ~n32857;
  assign n32870 = ~n6185 & n32848;
  assign n32871 = n16774 & ~n32870;
  assign n32872 = ~n32858 & n32871;
  assign n32873 = ~n32869 & ~n32872;
  assign n32874 = ~n32868 & n32873;
  assign n32875 = n6236 & n32874;
  assign n32876 = n32867 & ~n32875;
  assign n32877 = pi634 & pi680;
  assign n32878 = ~n32846 & n32877;
  assign n32879 = n32668 & ~n32878;
  assign n32880 = ~n6185 & ~n32644;
  assign n32881 = n6185 & ~n32652;
  assign n32882 = ~pi680 & ~n32881;
  assign n32883 = ~n32880 & n32882;
  assign n32884 = pi634 & ~n16603;
  assign n32885 = ~n32730 & ~n32884;
  assign n32886 = ~n6190 & ~n32885;
  assign n32887 = ~n32855 & ~n32886;
  assign n32888 = n6188 & ~n32887;
  assign n32889 = n6185 & n32887;
  assign n32890 = n32871 & ~n32889;
  assign n32891 = ~n32888 & ~n32890;
  assign n32892 = ~n32883 & n32891;
  assign n32893 = n6236 & ~n32892;
  assign n32894 = ~pi680 & n16294;
  assign n32895 = pi198 & n32894;
  assign n32896 = n6188 & ~n32885;
  assign n32897 = n6190 & n32885;
  assign n32898 = ~n32849 & ~n32897;
  assign n32899 = ~n6185 & ~n32898;
  assign n32900 = n6185 & n32885;
  assign n32901 = n16774 & ~n32900;
  assign n32902 = ~n32899 & n32901;
  assign n32903 = ~n32896 & ~n32902;
  assign n32904 = ~n32895 & n32903;
  assign n32905 = ~n6236 & ~n32904;
  assign n32906 = ~n2607 & ~n32905;
  assign n32907 = ~n32893 & n32906;
  assign n32908 = ~pi223 & ~n32907;
  assign n32909 = ~n32879 & n32908;
  assign n32910 = ~pi299 & ~n32909;
  assign n32911 = ~n32876 & n32910;
  assign n32912 = ~n6198 & n32865;
  assign n32913 = pi215 & ~n32912;
  assign n32914 = n6198 & n32874;
  assign n32915 = n32913 & ~n32914;
  assign n32916 = n32651 & ~n32878;
  assign n32917 = ~n6198 & ~n32904;
  assign n32918 = n6198 & ~n32892;
  assign n32919 = ~n2527 & ~n32918;
  assign n32920 = ~n32917 & n32919;
  assign n32921 = ~pi215 & ~n32920;
  assign n32922 = ~n32916 & n32921;
  assign n32923 = pi299 & ~n32922;
  assign n32924 = ~n32915 & n32923;
  assign n32925 = ~n32911 & ~n32924;
  assign n32926 = pi39 & ~n32925;
  assign n32927 = ~pi198 & n16733;
  assign n32928 = pi198 & ~n16716;
  assign n32929 = ~n32927 & ~n32928;
  assign n32930 = n32877 & n32929;
  assign n32931 = ~n32683 & ~n32877;
  assign n32932 = ~n32930 & ~n32931;
  assign n32933 = pi299 & n32932;
  assign n32934 = pi198 & n16706;
  assign n32935 = n32877 & ~n32934;
  assign n32936 = ~n16724 & n32935;
  assign n32937 = ~n16198 & ~n32936;
  assign n32938 = ~pi299 & ~n32937;
  assign n32939 = ~pi39 & ~n32938;
  assign n32940 = ~n32933 & n32939;
  assign n32941 = ~n32926 & ~n32940;
  assign n32942 = ~pi38 & ~n32941;
  assign n32943 = pi634 & n16596;
  assign n32944 = n16212 & n32943;
  assign n32945 = ~n32789 & ~n32944;
  assign n32946 = ~pi39 & ~n32945;
  assign n32947 = n32788 & ~n32946;
  assign n32948 = ~n32942 & ~n32947;
  assign n32949 = n10020 & n32948;
  assign n32950 = ~n32681 & ~n32949;
  assign n32951 = ~pi778 & ~n32950;
  assign n32952 = pi625 & n32950;
  assign n32953 = ~pi625 & n32679;
  assign n32954 = pi1153 & ~n32953;
  assign n32955 = ~n32952 & n32954;
  assign n32956 = ~pi625 & n32950;
  assign n32957 = pi625 & n32679;
  assign n32958 = ~pi1153 & ~n32957;
  assign n32959 = ~n32956 & n32958;
  assign n32960 = ~n32955 & ~n32959;
  assign n32961 = pi778 & ~n32960;
  assign n32962 = ~n32951 & ~n32961;
  assign n32963 = ~n16593 & n32962;
  assign n32964 = n16593 & n32679;
  assign n32965 = ~n32963 & ~n32964;
  assign n32966 = ~n16589 & n32965;
  assign n32967 = ~n32845 & ~n32966;
  assign n32968 = ~n17159 & n32967;
  assign n32969 = ~n17183 & n32968;
  assign n32970 = ~n32844 & ~n32969;
  assign n32971 = ~pi792 & n32970;
  assign n32972 = pi628 & ~n32970;
  assign n32973 = ~pi628 & n32679;
  assign n32974 = ~n32972 & ~n32973;
  assign n32975 = pi1156 & n32974;
  assign n32976 = ~pi628 & ~n32970;
  assign n32977 = pi628 & n32679;
  assign n32978 = ~pi1156 & ~n32977;
  assign n32979 = ~n32976 & n32978;
  assign n32980 = ~n32975 & ~n32979;
  assign n32981 = pi792 & ~n32980;
  assign n32982 = ~n32971 & ~n32981;
  assign n32983 = ~pi647 & n32982;
  assign n32984 = pi647 & n32679;
  assign n32985 = ~pi1157 & ~n32984;
  assign n32986 = ~n32983 & n32985;
  assign n32987 = ~pi647 & n32679;
  assign n32988 = pi647 & n32982;
  assign n32989 = pi1157 & ~n32988;
  assign n32990 = ~n32987 & n32989;
  assign n32991 = ~n32986 & ~n32990;
  assign n32992 = ~n17246 & ~n32991;
  assign n32993 = ~n32842 & ~n32992;
  assign n32994 = pi787 & ~n32993;
  assign n32995 = ~n19999 & n32839;
  assign n32996 = pi629 & n32979;
  assign n32997 = ~n32995 & ~n32996;
  assign n32998 = n16121 & n32974;
  assign n32999 = n32997 & ~n32998;
  assign n33000 = ~n19788 & n32999;
  assign n33001 = pi792 & ~n32999;
  assign n33002 = n17159 & n32679;
  assign n33003 = ~n32968 & ~n33002;
  assign n33004 = n17350 & ~n33003;
  assign n33005 = ~pi626 & ~n32836;
  assign n33006 = pi626 & ~n32679;
  assign n33007 = n17181 & ~n33006;
  assign n33008 = ~n33005 & n33007;
  assign n33009 = ~n33004 & ~n33008;
  assign n33010 = pi626 & ~n32836;
  assign n33011 = ~pi626 & ~n32679;
  assign n33012 = n17180 & ~n33011;
  assign n33013 = ~n33010 & n33012;
  assign n33014 = n33009 & ~n33013;
  assign n33015 = pi788 & ~n33014;
  assign n33016 = pi618 & ~n32965;
  assign n33017 = pi609 & n32962;
  assign n33018 = pi625 & n32797;
  assign n33019 = ~pi603 & n32929;
  assign n33020 = ~pi198 & ~pi665;
  assign n33021 = n16363 & n33020;
  assign n33022 = ~n16457 & n32928;
  assign n33023 = ~pi633 & ~n33022;
  assign n33024 = ~n33021 & n33023;
  assign n33025 = ~n32687 & n32929;
  assign n33026 = ~n33024 & n33025;
  assign n33027 = ~n33024 & ~n33026;
  assign n33028 = pi603 & ~n33027;
  assign n33029 = ~n33019 & ~n33028;
  assign n33030 = n32877 & n33029;
  assign n33031 = n32689 & ~n32877;
  assign n33032 = pi299 & ~n33031;
  assign n33033 = ~n33030 & n33032;
  assign n33034 = ~pi603 & n32937;
  assign n33035 = pi198 & ~pi633;
  assign n33036 = pi634 & ~pi665;
  assign n33037 = ~n33035 & n33036;
  assign n33038 = ~n16367 & n33037;
  assign n33039 = ~pi634 & ~n16198;
  assign n33040 = ~n16374 & n16707;
  assign n33041 = pi634 & ~n33040;
  assign n33042 = ~pi633 & ~n33041;
  assign n33043 = ~n33039 & n33042;
  assign n33044 = pi603 & ~n33043;
  assign n33045 = ~n33038 & n33044;
  assign n33046 = ~n32692 & n33045;
  assign n33047 = ~n33034 & ~n33046;
  assign n33048 = pi680 & n33047;
  assign n33049 = ~pi680 & n32694;
  assign n33050 = ~pi299 & ~n33049;
  assign n33051 = ~n33048 & n33050;
  assign n33052 = ~n33033 & ~n33051;
  assign n33053 = ~pi39 & ~n33052;
  assign n33054 = ~n16393 & ~n32885;
  assign n33055 = ~n32733 & ~n33054;
  assign n33056 = n6188 & ~n33055;
  assign n33057 = ~pi680 & ~n32741;
  assign n33058 = ~pi603 & n32898;
  assign n33059 = n16383 & n33036;
  assign n33060 = n32700 & ~n33059;
  assign n33061 = pi603 & ~n33060;
  assign n33062 = ~n16392 & n33061;
  assign n33063 = ~n32738 & ~n33062;
  assign n33064 = ~n6185 & n33063;
  assign n33065 = pi634 & n16858;
  assign n33066 = n32732 & ~n33065;
  assign n33067 = ~n6190 & ~n33063;
  assign n33068 = n33066 & ~n33067;
  assign n33069 = ~n33064 & ~n33068;
  assign n33070 = ~n33058 & ~n33069;
  assign n33071 = n16774 & ~n33070;
  assign n33072 = ~n33057 & ~n33071;
  assign n33073 = ~n33056 & n33072;
  assign n33074 = ~n6198 & ~n33073;
  assign n33075 = ~pi680 & n32756;
  assign n33076 = n6190 & ~n33060;
  assign n33077 = ~n6190 & ~n33066;
  assign n33078 = ~n33076 & ~n33077;
  assign n33079 = pi603 & ~n33078;
  assign n33080 = ~pi642 & n33079;
  assign n33081 = ~pi603 & ~n32848;
  assign n33082 = pi642 & n33061;
  assign n33083 = ~n33081 & ~n33082;
  assign n33084 = ~n33080 & n33083;
  assign n33085 = n6184 & ~n33084;
  assign n33086 = ~n33061 & ~n33081;
  assign n33087 = ~n6184 & ~n33086;
  assign n33088 = ~n6187 & ~n33087;
  assign n33089 = ~n33085 & n33088;
  assign n33090 = ~pi603 & ~n32887;
  assign n33091 = ~n33079 & ~n33090;
  assign n33092 = n6187 & n33091;
  assign n33093 = ~n33089 & ~n33092;
  assign n33094 = pi680 & ~n33093;
  assign n33095 = ~n33075 & ~n33094;
  assign n33096 = n6198 & n33095;
  assign n33097 = ~n2527 & ~n33096;
  assign n33098 = ~n33074 & n33097;
  assign n33099 = n16814 & n32847;
  assign n33100 = n32765 & ~n33099;
  assign n33101 = ~pi215 & ~n33100;
  assign n33102 = ~n33098 & n33101;
  assign n33103 = ~n16392 & n33086;
  assign n33104 = n16774 & ~n33103;
  assign n33105 = n16409 & n33036;
  assign n33106 = n32722 & ~n33105;
  assign n33107 = ~n6190 & ~n33106;
  assign n33108 = ~n33076 & ~n33107;
  assign n33109 = pi603 & ~n33108;
  assign n33110 = ~n33081 & ~n33109;
  assign n33111 = n16392 & n33110;
  assign n33112 = n33104 & ~n33111;
  assign n33113 = ~pi680 & n32712;
  assign n33114 = pi634 & n16909;
  assign n33115 = ~n32715 & ~n33114;
  assign n33116 = ~n33113 & n33115;
  assign n33117 = ~n33112 & n33116;
  assign n33118 = n6198 & n33117;
  assign n33119 = ~pi603 & n32852;
  assign n33120 = pi603 & n33106;
  assign n33121 = n6188 & ~n33120;
  assign n33122 = ~n33119 & n33121;
  assign n33123 = ~pi680 & ~n32719;
  assign n33124 = ~pi603 & n32854;
  assign n33125 = ~n33064 & ~n33106;
  assign n33126 = ~n33067 & ~n33125;
  assign n33127 = ~n33124 & n33126;
  assign n33128 = n16774 & ~n33127;
  assign n33129 = ~n33123 & ~n33128;
  assign n33130 = ~n33122 & n33129;
  assign n33131 = ~n6198 & n33130;
  assign n33132 = pi215 & ~n33131;
  assign n33133 = ~n33118 & n33132;
  assign n33134 = ~n33102 & ~n33133;
  assign n33135 = pi299 & ~n33134;
  assign n33136 = ~n6236 & ~n33073;
  assign n33137 = n6236 & n33095;
  assign n33138 = ~n2607 & ~n33137;
  assign n33139 = ~n33136 & n33138;
  assign n33140 = n32778 & ~n33099;
  assign n33141 = ~pi223 & ~n33140;
  assign n33142 = ~n33139 & n33141;
  assign n33143 = n6236 & n33117;
  assign n33144 = ~n6236 & n33130;
  assign n33145 = pi223 & ~n33144;
  assign n33146 = ~n33143 & n33145;
  assign n33147 = ~n33142 & ~n33146;
  assign n33148 = ~pi299 & ~n33147;
  assign n33149 = pi39 & ~n33148;
  assign n33150 = ~n33135 & n33149;
  assign n33151 = ~n33053 & ~n33150;
  assign n33152 = ~pi38 & ~n33151;
  assign n33153 = pi634 & n17626;
  assign n33154 = n32794 & ~n33153;
  assign n33155 = ~n33152 & ~n33154;
  assign n33156 = n10020 & n33155;
  assign n33157 = ~n32681 & ~n33156;
  assign n33158 = ~pi625 & n33157;
  assign n33159 = ~pi1153 & ~n33158;
  assign n33160 = ~n33018 & n33159;
  assign n33161 = ~pi608 & ~n32955;
  assign n33162 = ~n33160 & n33161;
  assign n33163 = ~pi625 & n32797;
  assign n33164 = pi625 & n33157;
  assign n33165 = ~n33163 & ~n33164;
  assign n33166 = pi1153 & n33165;
  assign n33167 = ~n32959 & ~n33166;
  assign n33168 = pi608 & n33167;
  assign n33169 = ~n33162 & ~n33168;
  assign n33170 = pi778 & ~n33169;
  assign n33171 = ~pi778 & n33157;
  assign n33172 = ~n33170 & ~n33171;
  assign n33173 = ~pi609 & ~n33172;
  assign n33174 = ~pi1155 & ~n33173;
  assign n33175 = ~n33017 & n33174;
  assign n33176 = ~pi660 & ~n32805;
  assign n33177 = ~n33175 & n33176;
  assign n33178 = ~pi609 & n32962;
  assign n33179 = pi609 & ~n33172;
  assign n33180 = ~n33178 & ~n33179;
  assign n33181 = pi1155 & n33180;
  assign n33182 = ~n32809 & ~n33181;
  assign n33183 = pi660 & n33182;
  assign n33184 = ~n33177 & ~n33183;
  assign n33185 = pi785 & ~n33184;
  assign n33186 = ~pi785 & ~n33172;
  assign n33187 = ~n33185 & ~n33186;
  assign n33188 = ~pi618 & ~n33187;
  assign n33189 = ~pi1154 & ~n33188;
  assign n33190 = ~n33016 & n33189;
  assign n33191 = ~pi627 & ~n32817;
  assign n33192 = ~n33190 & n33191;
  assign n33193 = ~pi618 & ~n32965;
  assign n33194 = pi618 & ~n33187;
  assign n33195 = ~n33193 & ~n33194;
  assign n33196 = pi1154 & n33195;
  assign n33197 = ~n32821 & ~n33196;
  assign n33198 = pi627 & n33197;
  assign n33199 = ~n33192 & ~n33198;
  assign n33200 = pi781 & ~n33199;
  assign n33201 = ~pi781 & ~n33187;
  assign n33202 = ~n33200 & ~n33201;
  assign n33203 = ~pi619 & ~n33202;
  assign n33204 = pi619 & n32967;
  assign n33205 = ~pi1159 & ~n33204;
  assign n33206 = ~n33203 & n33205;
  assign n33207 = ~pi648 & ~n33206;
  assign n33208 = ~n32829 & n33207;
  assign n33209 = ~pi619 & n32967;
  assign n33210 = pi619 & ~n33202;
  assign n33211 = ~n33209 & ~n33210;
  assign n33212 = pi1159 & n33211;
  assign n33213 = ~n32833 & ~n33212;
  assign n33214 = pi648 & n33213;
  assign n33215 = ~n33208 & ~n33214;
  assign n33216 = pi789 & n33215;
  assign n33217 = ~pi789 & n33202;
  assign n33218 = n17356 & ~n33217;
  assign n33219 = ~n33216 & n33218;
  assign n33220 = ~n33015 & ~n33219;
  assign n33221 = ~n33001 & ~n33220;
  assign n33222 = ~n33000 & ~n33221;
  assign n33223 = n19637 & n33222;
  assign n33224 = ~n32994 & ~n33223;
  assign n33225 = ~pi790 & ~n33224;
  assign n33226 = ~n17247 & n32841;
  assign n33227 = n17247 & n32679;
  assign n33228 = ~n33226 & ~n33227;
  assign n33229 = ~pi644 & ~n33228;
  assign n33230 = pi715 & ~n33229;
  assign n33231 = pi644 & n32679;
  assign n33232 = n33230 & ~n33231;
  assign n33233 = ~pi787 & ~n32982;
  assign n33234 = pi787 & ~n32991;
  assign n33235 = ~n33233 & ~n33234;
  assign n33236 = pi644 & n33235;
  assign n33237 = ~pi644 & n33224;
  assign n33238 = ~pi715 & ~n33237;
  assign n33239 = ~n33236 & n33238;
  assign n33240 = ~pi1160 & ~n33239;
  assign n33241 = ~n33232 & n33240;
  assign n33242 = pi644 & n33224;
  assign n33243 = ~pi644 & n33235;
  assign n33244 = pi715 & ~n33243;
  assign n33245 = ~n33242 & n33244;
  assign n33246 = ~pi644 & n32679;
  assign n33247 = pi644 & ~n33228;
  assign n33248 = ~pi715 & ~n33247;
  assign n33249 = ~n33246 & n33248;
  assign n33250 = ~n33245 & ~n33249;
  assign n33251 = pi1160 & n33250;
  assign n33252 = ~n33241 & ~n33251;
  assign n33253 = pi790 & n33252;
  assign n33254 = ~n33225 & ~n33253;
  assign n33255 = ~po1038 & ~n33254;
  assign n33256 = pi198 & po1038;
  assign po355 = n33255 | n33256;
  assign n33258 = pi199 & ~n16527;
  assign n33259 = ~pi617 & ~n33258;
  assign n33260 = n6132 & n16510;
  assign n33261 = ~pi199 & ~n33260;
  assign n33262 = n18807 & ~n33261;
  assign n33263 = pi199 & n16449;
  assign n33264 = ~pi199 & ~n16503;
  assign n33265 = ~pi38 & ~n33264;
  assign n33266 = ~n33263 & n33265;
  assign n33267 = ~n33262 & ~n33266;
  assign n33268 = n10020 & ~n33267;
  assign n33269 = pi199 & ~n10020;
  assign n33270 = ~n33268 & ~n33269;
  assign n33271 = pi617 & n33270;
  assign n33272 = ~n33259 & ~n33271;
  assign n33273 = ~n16521 & n33272;
  assign n33274 = n16521 & n33258;
  assign n33275 = ~n33273 & ~n33274;
  assign n33276 = ~pi785 & ~n33275;
  assign n33277 = pi609 & n33275;
  assign n33278 = ~pi609 & ~n33258;
  assign n33279 = pi1155 & ~n33278;
  assign n33280 = ~n33277 & n33279;
  assign n33281 = ~pi609 & n33275;
  assign n33282 = pi609 & ~n33258;
  assign n33283 = ~pi1155 & ~n33282;
  assign n33284 = ~n33281 & n33283;
  assign n33285 = ~n33280 & ~n33284;
  assign n33286 = pi785 & ~n33285;
  assign n33287 = ~n33276 & ~n33286;
  assign n33288 = ~pi781 & ~n33287;
  assign n33289 = pi618 & n33287;
  assign n33290 = ~pi618 & ~n33258;
  assign n33291 = pi1154 & ~n33290;
  assign n33292 = ~n33289 & n33291;
  assign n33293 = ~pi618 & n33287;
  assign n33294 = pi618 & ~n33258;
  assign n33295 = ~pi1154 & ~n33294;
  assign n33296 = ~n33293 & n33295;
  assign n33297 = ~n33292 & ~n33296;
  assign n33298 = pi781 & ~n33297;
  assign n33299 = ~n33288 & ~n33298;
  assign n33300 = ~pi789 & ~n33299;
  assign n33301 = pi619 & n33299;
  assign n33302 = ~pi619 & ~n33258;
  assign n33303 = pi1159 & ~n33302;
  assign n33304 = ~n33301 & n33303;
  assign n33305 = ~pi619 & n33299;
  assign n33306 = pi619 & ~n33258;
  assign n33307 = ~pi1159 & ~n33306;
  assign n33308 = ~n33305 & n33307;
  assign n33309 = ~n33304 & ~n33308;
  assign n33310 = pi789 & ~n33309;
  assign n33311 = ~n33300 & ~n33310;
  assign n33312 = ~n17355 & ~n33311;
  assign n33313 = n17355 & n33258;
  assign n33314 = ~n33312 & ~n33313;
  assign n33315 = ~n16124 & ~n33314;
  assign n33316 = n16124 & n33258;
  assign n33317 = ~n33315 & ~n33316;
  assign n33318 = pi647 & n33317;
  assign n33319 = pi628 & n33314;
  assign n33320 = n16593 & ~n33258;
  assign n33321 = ~pi637 & ~n33258;
  assign n33322 = ~pi199 & ~n16508;
  assign n33323 = n19410 & ~n33322;
  assign n33324 = pi199 & ~n16702;
  assign n33325 = ~pi199 & ~n16639;
  assign n33326 = pi39 & ~n33325;
  assign n33327 = ~n33324 & n33326;
  assign n33328 = ~pi199 & n16736;
  assign n33329 = pi199 & ~n16720;
  assign n33330 = ~pi39 & ~n33329;
  assign n33331 = ~n33328 & n33330;
  assign n33332 = ~pi38 & ~n33331;
  assign n33333 = ~n33327 & n33332;
  assign n33334 = ~n33323 & ~n33333;
  assign n33335 = n10020 & ~n33334;
  assign n33336 = ~n33269 & ~n33335;
  assign n33337 = pi637 & n33336;
  assign n33338 = ~n33321 & ~n33337;
  assign n33339 = ~pi778 & n33338;
  assign n33340 = pi625 & ~n33338;
  assign n33341 = ~pi625 & ~n33258;
  assign n33342 = pi1153 & ~n33341;
  assign n33343 = ~n33340 & n33342;
  assign n33344 = ~pi625 & ~n33338;
  assign n33345 = pi625 & ~n33258;
  assign n33346 = ~pi1153 & ~n33345;
  assign n33347 = ~n33344 & n33346;
  assign n33348 = ~n33343 & ~n33347;
  assign n33349 = pi778 & ~n33348;
  assign n33350 = ~n33339 & ~n33349;
  assign n33351 = ~n16593 & n33350;
  assign n33352 = ~n33320 & ~n33351;
  assign n33353 = ~n16589 & n33352;
  assign n33354 = n16589 & n33258;
  assign n33355 = ~n33353 & ~n33354;
  assign n33356 = pi619 & n33355;
  assign n33357 = pi618 & ~n33352;
  assign n33358 = pi609 & n33350;
  assign n33359 = pi625 & ~n33272;
  assign n33360 = ~pi637 & n33272;
  assign n33361 = n10020 & ~n23889;
  assign n33362 = ~pi199 & ~n33361;
  assign n33363 = ~pi617 & ~n33362;
  assign n33364 = ~n18934 & n33363;
  assign n33365 = pi199 & n18938;
  assign n33366 = n33364 & ~n33365;
  assign n33367 = n10020 & n18922;
  assign n33368 = ~pi199 & ~n33367;
  assign n33369 = pi199 & n18914;
  assign n33370 = ~n33368 & ~n33369;
  assign n33371 = pi617 & n33370;
  assign n33372 = ~n33269 & ~n33371;
  assign n33373 = ~n33366 & n33372;
  assign n33374 = pi637 & ~n33373;
  assign n33375 = ~n33360 & ~n33374;
  assign n33376 = ~pi625 & n33375;
  assign n33377 = ~pi1153 & ~n33376;
  assign n33378 = ~n33359 & n33377;
  assign n33379 = ~pi608 & ~n33343;
  assign n33380 = ~n33378 & n33379;
  assign n33381 = ~pi625 & ~n33272;
  assign n33382 = pi625 & n33375;
  assign n33383 = ~n33381 & ~n33382;
  assign n33384 = pi1153 & n33383;
  assign n33385 = ~n33347 & ~n33384;
  assign n33386 = pi608 & n33385;
  assign n33387 = ~n33380 & ~n33386;
  assign n33388 = pi778 & ~n33387;
  assign n33389 = ~pi778 & n33375;
  assign n33390 = ~n33388 & ~n33389;
  assign n33391 = ~pi609 & ~n33390;
  assign n33392 = ~pi1155 & ~n33391;
  assign n33393 = ~n33358 & n33392;
  assign n33394 = ~pi660 & ~n33280;
  assign n33395 = ~n33393 & n33394;
  assign n33396 = ~pi609 & n33350;
  assign n33397 = pi609 & ~n33390;
  assign n33398 = ~n33396 & ~n33397;
  assign n33399 = pi1155 & n33398;
  assign n33400 = ~n33284 & ~n33399;
  assign n33401 = pi660 & n33400;
  assign n33402 = ~n33395 & ~n33401;
  assign n33403 = pi785 & ~n33402;
  assign n33404 = ~pi785 & ~n33390;
  assign n33405 = ~n33403 & ~n33404;
  assign n33406 = ~pi618 & ~n33405;
  assign n33407 = ~pi1154 & ~n33406;
  assign n33408 = ~n33357 & n33407;
  assign n33409 = ~pi627 & ~n33292;
  assign n33410 = ~n33408 & n33409;
  assign n33411 = ~pi618 & ~n33352;
  assign n33412 = pi618 & ~n33405;
  assign n33413 = ~n33411 & ~n33412;
  assign n33414 = pi1154 & n33413;
  assign n33415 = ~n33296 & ~n33414;
  assign n33416 = pi627 & n33415;
  assign n33417 = ~n33410 & ~n33416;
  assign n33418 = pi781 & ~n33417;
  assign n33419 = ~pi781 & ~n33405;
  assign n33420 = ~n33418 & ~n33419;
  assign n33421 = ~pi619 & ~n33420;
  assign n33422 = ~pi1159 & ~n33421;
  assign n33423 = ~n33356 & n33422;
  assign n33424 = ~pi648 & ~n33304;
  assign n33425 = ~n33423 & n33424;
  assign n33426 = ~pi619 & n33355;
  assign n33427 = pi619 & ~n33420;
  assign n33428 = ~n33426 & ~n33427;
  assign n33429 = pi1159 & n33428;
  assign n33430 = ~n33308 & ~n33429;
  assign n33431 = pi648 & n33430;
  assign n33432 = ~n33425 & ~n33431;
  assign n33433 = pi789 & ~n33432;
  assign n33434 = ~pi789 & ~n33420;
  assign n33435 = ~n33433 & ~n33434;
  assign n33436 = ~pi788 & n33435;
  assign n33437 = pi626 & n33435;
  assign n33438 = n17159 & ~n33258;
  assign n33439 = ~n17159 & n33355;
  assign n33440 = ~n33438 & ~n33439;
  assign n33441 = ~pi626 & n33440;
  assign n33442 = pi641 & ~n33441;
  assign n33443 = ~n33437 & n33442;
  assign n33444 = pi626 & ~n33311;
  assign n33445 = ~pi626 & n33258;
  assign n33446 = ~pi641 & ~n33445;
  assign n33447 = ~n33444 & n33446;
  assign n33448 = pi1158 & ~n33447;
  assign n33449 = ~n33443 & n33448;
  assign n33450 = ~pi626 & ~n33311;
  assign n33451 = pi641 & ~n33450;
  assign n33452 = pi626 & n33258;
  assign n33453 = n33451 & ~n33452;
  assign n33454 = pi626 & n33440;
  assign n33455 = ~pi626 & n33435;
  assign n33456 = ~pi641 & ~n33455;
  assign n33457 = ~n33454 & n33456;
  assign n33458 = ~pi1158 & ~n33457;
  assign n33459 = ~n33453 & n33458;
  assign n33460 = ~n33449 & ~n33459;
  assign n33461 = pi788 & ~n33460;
  assign n33462 = ~n33436 & ~n33461;
  assign n33463 = ~pi628 & n33462;
  assign n33464 = ~pi1156 & ~n33463;
  assign n33465 = ~n33319 & n33464;
  assign n33466 = ~n17183 & n33440;
  assign n33467 = n17183 & n33258;
  assign n33468 = ~n33466 & ~n33467;
  assign n33469 = pi628 & n33468;
  assign n33470 = ~pi628 & ~n33258;
  assign n33471 = pi1156 & ~n33470;
  assign n33472 = ~n33469 & n33471;
  assign n33473 = ~pi629 & ~n33472;
  assign n33474 = ~n33465 & n33473;
  assign n33475 = ~pi628 & n33468;
  assign n33476 = pi628 & ~n33258;
  assign n33477 = ~pi1156 & ~n33476;
  assign n33478 = ~n33475 & n33477;
  assign n33479 = ~pi628 & n33314;
  assign n33480 = pi628 & n33462;
  assign n33481 = ~n33479 & ~n33480;
  assign n33482 = pi1156 & n33481;
  assign n33483 = ~n33478 & ~n33482;
  assign n33484 = pi629 & n33483;
  assign n33485 = ~n33474 & ~n33484;
  assign n33486 = pi792 & ~n33485;
  assign n33487 = ~pi792 & n33462;
  assign n33488 = ~n33486 & ~n33487;
  assign n33489 = ~pi647 & ~n33488;
  assign n33490 = ~pi1157 & ~n33489;
  assign n33491 = ~n33318 & n33490;
  assign n33492 = ~pi792 & ~n33468;
  assign n33493 = ~n33472 & ~n33478;
  assign n33494 = pi792 & ~n33493;
  assign n33495 = ~n33492 & ~n33494;
  assign n33496 = pi647 & n33495;
  assign n33497 = ~pi647 & ~n33258;
  assign n33498 = pi1157 & ~n33497;
  assign n33499 = ~n33496 & n33498;
  assign n33500 = ~pi630 & ~n33499;
  assign n33501 = ~n33491 & n33500;
  assign n33502 = ~pi647 & n33495;
  assign n33503 = pi647 & ~n33258;
  assign n33504 = ~pi1157 & ~n33503;
  assign n33505 = ~n33502 & n33504;
  assign n33506 = ~pi647 & n33317;
  assign n33507 = pi647 & ~n33488;
  assign n33508 = ~n33506 & ~n33507;
  assign n33509 = pi1157 & n33508;
  assign n33510 = ~n33505 & ~n33509;
  assign n33511 = pi630 & n33510;
  assign n33512 = ~n33501 & ~n33511;
  assign n33513 = pi787 & ~n33512;
  assign n33514 = ~pi787 & ~n33488;
  assign n33515 = ~n33513 & ~n33514;
  assign n33516 = ~pi790 & n33515;
  assign n33517 = pi644 & ~n33258;
  assign n33518 = n17247 & ~n33258;
  assign n33519 = ~n17247 & n33317;
  assign n33520 = ~n33518 & ~n33519;
  assign n33521 = ~pi644 & ~n33520;
  assign n33522 = pi715 & ~n33521;
  assign n33523 = ~n33517 & n33522;
  assign n33524 = ~pi787 & ~n33495;
  assign n33525 = ~n33499 & ~n33505;
  assign n33526 = pi787 & ~n33525;
  assign n33527 = ~n33524 & ~n33526;
  assign n33528 = pi644 & n33527;
  assign n33529 = ~pi644 & ~n33515;
  assign n33530 = ~pi715 & ~n33529;
  assign n33531 = ~n33528 & n33530;
  assign n33532 = ~pi1160 & ~n33531;
  assign n33533 = ~n33523 & n33532;
  assign n33534 = pi644 & ~n33515;
  assign n33535 = ~pi644 & n33527;
  assign n33536 = pi715 & ~n33535;
  assign n33537 = ~n33534 & n33536;
  assign n33538 = ~pi644 & ~n33258;
  assign n33539 = pi644 & ~n33520;
  assign n33540 = ~pi715 & ~n33539;
  assign n33541 = ~n33538 & n33540;
  assign n33542 = ~n33537 & ~n33541;
  assign n33543 = pi1160 & n33542;
  assign n33544 = ~n33533 & ~n33543;
  assign n33545 = pi790 & n33544;
  assign n33546 = ~n33516 & ~n33545;
  assign n33547 = ~po1038 & ~n33546;
  assign n33548 = pi199 & po1038;
  assign po356 = n33547 | n33548;
  assign n33550 = pi200 & ~n16527;
  assign n33551 = n17159 & ~n33550;
  assign n33552 = n16593 & ~n33550;
  assign n33553 = ~pi643 & ~n33550;
  assign n33554 = pi200 & ~n10020;
  assign n33555 = ~pi200 & ~n16508;
  assign n33556 = n19410 & ~n33555;
  assign n33557 = pi200 & n16687;
  assign n33558 = ~pi200 & n16624;
  assign n33559 = ~pi299 & ~n33558;
  assign n33560 = ~n33557 & n33559;
  assign n33561 = pi200 & n16700;
  assign n33562 = ~pi200 & n16637;
  assign n33563 = pi299 & ~n33562;
  assign n33564 = ~n33561 & n33563;
  assign n33565 = ~n33560 & ~n33564;
  assign n33566 = pi39 & ~n33565;
  assign n33567 = pi200 & n16720;
  assign n33568 = ~pi200 & ~n16736;
  assign n33569 = ~pi39 & ~n33568;
  assign n33570 = ~n33567 & n33569;
  assign n33571 = ~n33566 & ~n33570;
  assign n33572 = ~pi38 & ~n33571;
  assign n33573 = ~n33556 & ~n33572;
  assign n33574 = n10020 & ~n33573;
  assign n33575 = ~n33554 & ~n33574;
  assign n33576 = pi643 & n33575;
  assign n33577 = ~n33553 & ~n33576;
  assign n33578 = ~pi778 & n33577;
  assign n33579 = pi625 & ~n33577;
  assign n33580 = ~pi625 & ~n33550;
  assign n33581 = pi1153 & ~n33580;
  assign n33582 = ~n33579 & n33581;
  assign n33583 = ~pi625 & ~n33577;
  assign n33584 = pi625 & ~n33550;
  assign n33585 = ~pi1153 & ~n33584;
  assign n33586 = ~n33583 & n33585;
  assign n33587 = ~n33582 & ~n33586;
  assign n33588 = pi778 & ~n33587;
  assign n33589 = ~n33578 & ~n33588;
  assign n33590 = ~n16593 & n33589;
  assign n33591 = ~n33552 & ~n33590;
  assign n33592 = ~n16589 & n33591;
  assign n33593 = n16589 & n33550;
  assign n33594 = ~n33592 & ~n33593;
  assign n33595 = ~n17159 & n33594;
  assign n33596 = ~n33551 & ~n33595;
  assign n33597 = ~n17183 & n33596;
  assign n33598 = n17183 & n33550;
  assign n33599 = ~n33597 & ~n33598;
  assign n33600 = pi628 & n33599;
  assign n33601 = ~pi628 & ~n33550;
  assign n33602 = pi1156 & ~n33601;
  assign n33603 = ~n33600 & n33602;
  assign n33604 = ~pi629 & n33603;
  assign n33605 = ~pi606 & ~n33550;
  assign n33606 = ~pi200 & ~n33260;
  assign n33607 = n18807 & ~n33606;
  assign n33608 = pi200 & n16449;
  assign n33609 = ~pi200 & ~n16503;
  assign n33610 = ~pi38 & ~n33609;
  assign n33611 = ~n33608 & n33610;
  assign n33612 = ~n33607 & ~n33611;
  assign n33613 = n10020 & ~n33612;
  assign n33614 = ~n33554 & ~n33613;
  assign n33615 = pi606 & n33614;
  assign n33616 = ~n33605 & ~n33615;
  assign n33617 = ~n16521 & n33616;
  assign n33618 = n16521 & n33550;
  assign n33619 = ~n33617 & ~n33618;
  assign n33620 = ~pi785 & ~n33619;
  assign n33621 = pi609 & n33619;
  assign n33622 = ~pi609 & ~n33550;
  assign n33623 = pi1155 & ~n33622;
  assign n33624 = ~n33621 & n33623;
  assign n33625 = ~pi609 & n33619;
  assign n33626 = pi609 & ~n33550;
  assign n33627 = ~pi1155 & ~n33626;
  assign n33628 = ~n33625 & n33627;
  assign n33629 = ~n33624 & ~n33628;
  assign n33630 = pi785 & ~n33629;
  assign n33631 = ~n33620 & ~n33630;
  assign n33632 = ~pi781 & ~n33631;
  assign n33633 = pi618 & n33631;
  assign n33634 = ~pi618 & ~n33550;
  assign n33635 = pi1154 & ~n33634;
  assign n33636 = ~n33633 & n33635;
  assign n33637 = ~pi618 & n33631;
  assign n33638 = pi618 & ~n33550;
  assign n33639 = ~pi1154 & ~n33638;
  assign n33640 = ~n33637 & n33639;
  assign n33641 = ~n33636 & ~n33640;
  assign n33642 = pi781 & ~n33641;
  assign n33643 = ~n33632 & ~n33642;
  assign n33644 = ~pi789 & ~n33643;
  assign n33645 = pi619 & n33643;
  assign n33646 = ~pi619 & ~n33550;
  assign n33647 = pi1159 & ~n33646;
  assign n33648 = ~n33645 & n33647;
  assign n33649 = ~pi619 & n33643;
  assign n33650 = pi619 & ~n33550;
  assign n33651 = ~pi1159 & ~n33650;
  assign n33652 = ~n33649 & n33651;
  assign n33653 = ~n33648 & ~n33652;
  assign n33654 = pi789 & ~n33653;
  assign n33655 = ~n33644 & ~n33654;
  assign n33656 = ~n17355 & ~n33655;
  assign n33657 = n17355 & n33550;
  assign n33658 = ~n33656 & ~n33657;
  assign n33659 = ~n19999 & ~n33658;
  assign n33660 = ~pi628 & n33599;
  assign n33661 = pi628 & ~n33550;
  assign n33662 = ~pi1156 & ~n33661;
  assign n33663 = ~n33660 & n33662;
  assign n33664 = pi629 & n33663;
  assign n33665 = ~n33659 & ~n33664;
  assign n33666 = ~n33604 & n33665;
  assign n33667 = pi792 & ~n33666;
  assign n33668 = pi618 & ~n33591;
  assign n33669 = pi609 & n33589;
  assign n33670 = pi625 & ~n33616;
  assign n33671 = ~pi643 & n33616;
  assign n33672 = pi200 & ~n24082;
  assign n33673 = ~pi200 & ~n18917;
  assign n33674 = ~pi38 & ~n33673;
  assign n33675 = ~n33672 & n33674;
  assign n33676 = pi200 & n18931;
  assign n33677 = n16917 & n33676;
  assign n33678 = ~n18916 & ~n18921;
  assign n33679 = ~pi200 & ~n33678;
  assign n33680 = n10020 & ~n33679;
  assign n33681 = pi606 & n33680;
  assign n33682 = ~n33677 & n33681;
  assign n33683 = ~n33675 & n33682;
  assign n33684 = ~n16511 & n33556;
  assign n33685 = pi200 & ~n18937;
  assign n33686 = ~pi200 & ~n18928;
  assign n33687 = ~pi38 & ~n33686;
  assign n33688 = ~n33685 & n33687;
  assign n33689 = ~n33684 & ~n33688;
  assign n33690 = ~pi606 & n10020;
  assign n33691 = ~n33689 & n33690;
  assign n33692 = ~n33554 & ~n33691;
  assign n33693 = ~n33683 & n33692;
  assign n33694 = pi643 & ~n33693;
  assign n33695 = ~n33671 & ~n33694;
  assign n33696 = ~pi625 & n33695;
  assign n33697 = ~pi1153 & ~n33696;
  assign n33698 = ~n33670 & n33697;
  assign n33699 = ~pi608 & ~n33582;
  assign n33700 = ~n33698 & n33699;
  assign n33701 = ~pi625 & ~n33616;
  assign n33702 = pi625 & n33695;
  assign n33703 = ~n33701 & ~n33702;
  assign n33704 = pi1153 & n33703;
  assign n33705 = ~n33586 & ~n33704;
  assign n33706 = pi608 & n33705;
  assign n33707 = ~n33700 & ~n33706;
  assign n33708 = pi778 & ~n33707;
  assign n33709 = ~pi778 & n33695;
  assign n33710 = ~n33708 & ~n33709;
  assign n33711 = ~pi609 & ~n33710;
  assign n33712 = ~pi1155 & ~n33711;
  assign n33713 = ~n33669 & n33712;
  assign n33714 = ~pi660 & ~n33624;
  assign n33715 = ~n33713 & n33714;
  assign n33716 = ~pi609 & n33589;
  assign n33717 = pi609 & ~n33710;
  assign n33718 = ~n33716 & ~n33717;
  assign n33719 = pi1155 & n33718;
  assign n33720 = ~n33628 & ~n33719;
  assign n33721 = pi660 & n33720;
  assign n33722 = ~n33715 & ~n33721;
  assign n33723 = pi785 & ~n33722;
  assign n33724 = ~pi785 & ~n33710;
  assign n33725 = ~n33723 & ~n33724;
  assign n33726 = ~pi618 & ~n33725;
  assign n33727 = ~pi1154 & ~n33726;
  assign n33728 = ~n33668 & n33727;
  assign n33729 = ~pi627 & ~n33636;
  assign n33730 = ~n33728 & n33729;
  assign n33731 = ~pi618 & ~n33591;
  assign n33732 = pi618 & ~n33725;
  assign n33733 = ~n33731 & ~n33732;
  assign n33734 = pi1154 & n33733;
  assign n33735 = ~n33640 & ~n33734;
  assign n33736 = pi627 & n33735;
  assign n33737 = ~n33730 & ~n33736;
  assign n33738 = pi781 & ~n33737;
  assign n33739 = ~pi781 & ~n33725;
  assign n33740 = ~n33738 & ~n33739;
  assign n33741 = ~pi789 & n33740;
  assign n33742 = ~pi619 & ~n33740;
  assign n33743 = pi619 & n33594;
  assign n33744 = ~pi1159 & ~n33743;
  assign n33745 = ~n33742 & n33744;
  assign n33746 = ~pi648 & ~n33745;
  assign n33747 = ~n33648 & n33746;
  assign n33748 = ~pi619 & n33594;
  assign n33749 = pi619 & ~n33740;
  assign n33750 = ~n33748 & ~n33749;
  assign n33751 = pi1159 & n33750;
  assign n33752 = ~n33652 & ~n33751;
  assign n33753 = pi648 & n33752;
  assign n33754 = ~n33747 & ~n33753;
  assign n33755 = pi789 & n33754;
  assign n33756 = ~n33741 & ~n33755;
  assign n33757 = n17356 & n33756;
  assign n33758 = ~pi626 & ~n33655;
  assign n33759 = pi626 & n33550;
  assign n33760 = n17181 & ~n33759;
  assign n33761 = ~n33758 & n33760;
  assign n33762 = n17350 & ~n33596;
  assign n33763 = pi626 & ~n33655;
  assign n33764 = ~pi626 & n33550;
  assign n33765 = n17180 & ~n33764;
  assign n33766 = ~n33763 & n33765;
  assign n33767 = ~n33762 & ~n33766;
  assign n33768 = ~n33761 & n33767;
  assign n33769 = pi788 & ~n33768;
  assign n33770 = n19788 & ~n33769;
  assign n33771 = ~n33757 & n33770;
  assign n33772 = ~n33667 & ~n33771;
  assign n33773 = n19637 & ~n33772;
  assign n33774 = ~pi792 & ~n33599;
  assign n33775 = ~n33603 & ~n33663;
  assign n33776 = pi792 & ~n33775;
  assign n33777 = ~n33774 & ~n33776;
  assign n33778 = ~pi647 & n33777;
  assign n33779 = pi647 & ~n33550;
  assign n33780 = ~pi1157 & ~n33779;
  assign n33781 = ~n33778 & n33780;
  assign n33782 = pi630 & n33781;
  assign n33783 = ~n16124 & ~n33658;
  assign n33784 = n16124 & n33550;
  assign n33785 = ~n33783 & ~n33784;
  assign n33786 = ~n19987 & ~n33785;
  assign n33787 = ~n33782 & ~n33786;
  assign n33788 = pi647 & ~n33777;
  assign n33789 = ~pi647 & n33550;
  assign n33790 = ~n33788 & ~n33789;
  assign n33791 = n17244 & ~n33790;
  assign n33792 = n33787 & ~n33791;
  assign n33793 = pi787 & ~n33792;
  assign n33794 = ~n33773 & ~n33793;
  assign n33795 = pi644 & n33794;
  assign n33796 = ~pi787 & ~n33777;
  assign n33797 = pi1157 & ~n33790;
  assign n33798 = ~n33781 & ~n33797;
  assign n33799 = pi787 & ~n33798;
  assign n33800 = ~n33796 & ~n33799;
  assign n33801 = ~pi644 & n33800;
  assign n33802 = pi715 & ~n33801;
  assign n33803 = ~n33795 & n33802;
  assign n33804 = n17247 & ~n33550;
  assign n33805 = ~n17247 & n33785;
  assign n33806 = ~n33804 & ~n33805;
  assign n33807 = pi644 & ~n33806;
  assign n33808 = ~pi644 & ~n33550;
  assign n33809 = ~pi715 & ~n33808;
  assign n33810 = ~n33807 & n33809;
  assign n33811 = pi1160 & ~n33810;
  assign n33812 = ~n33803 & n33811;
  assign n33813 = pi644 & ~n33550;
  assign n33814 = ~pi644 & ~n33806;
  assign n33815 = pi715 & ~n33814;
  assign n33816 = ~n33813 & n33815;
  assign n33817 = pi644 & n33800;
  assign n33818 = ~pi644 & n33794;
  assign n33819 = ~pi715 & ~n33818;
  assign n33820 = ~n33817 & n33819;
  assign n33821 = ~pi1160 & ~n33820;
  assign n33822 = ~n33816 & n33821;
  assign n33823 = ~n33812 & ~n33822;
  assign n33824 = pi790 & ~n33823;
  assign n33825 = ~pi790 & n33794;
  assign n33826 = ~n33824 & ~n33825;
  assign n33827 = ~po1038 & ~n33826;
  assign n33828 = ~pi200 & po1038;
  assign po357 = ~n33827 & ~n33828;
  assign n33830 = pi233 & pi237;
  assign n33831 = ~pi332 & ~n6185;
  assign n33832 = ~pi947 & ~n33831;
  assign n33833 = pi96 & pi210;
  assign n33834 = pi332 & n33833;
  assign n33835 = ~pi70 & ~pi841;
  assign n33836 = pi32 & ~n33835;
  assign n33837 = ~pi32 & ~pi70;
  assign n33838 = ~n33836 & ~n33837;
  assign n33839 = ~pi210 & n33838;
  assign n33840 = ~pi32 & ~pi96;
  assign n33841 = pi70 & n33840;
  assign n33842 = ~pi332 & ~n33841;
  assign n33843 = ~n33839 & n33842;
  assign n33844 = ~n33834 & ~n33843;
  assign n33845 = ~n6190 & n33844;
  assign n33846 = n6185 & ~n33845;
  assign n33847 = n33832 & ~n33846;
  assign n33848 = n6185 & ~n33844;
  assign n33849 = pi947 & ~n33848;
  assign n33850 = pi332 & pi468;
  assign n33851 = ~pi468 & ~n33843;
  assign n33852 = ~n33850 & ~n33851;
  assign n33853 = ~n6185 & n33852;
  assign n33854 = n33849 & ~n33853;
  assign n33855 = ~n33847 & ~n33854;
  assign n33856 = pi57 & ~n33855;
  assign n33857 = ~n2576 & n33855;
  assign n33858 = ~pi95 & n2902;
  assign n33859 = ~pi70 & ~n33858;
  assign n33860 = n33840 & ~n33859;
  assign n33861 = pi210 & n33860;
  assign n33862 = ~pi95 & n2686;
  assign n33863 = ~pi96 & n33862;
  assign n33864 = ~n33836 & n33863;
  assign n33865 = n10858 & n33864;
  assign n33866 = n2505 & n33865;
  assign n33867 = ~n33838 & ~n33866;
  assign n33868 = ~pi210 & ~n33867;
  assign n33869 = ~pi332 & ~n33868;
  assign n33870 = ~n33861 & n33869;
  assign n33871 = ~n33834 & ~n33870;
  assign n33872 = ~n6190 & n33871;
  assign n33873 = n6185 & ~n33872;
  assign n33874 = n33832 & ~n33873;
  assign n33875 = n6185 & ~n33871;
  assign n33876 = pi947 & ~n33875;
  assign n33877 = ~pi468 & ~n33870;
  assign n33878 = ~n33850 & ~n33877;
  assign n33879 = ~n6185 & n33878;
  assign n33880 = n33876 & ~n33879;
  assign n33881 = ~n33874 & ~n33880;
  assign n33882 = n2576 & n33881;
  assign n33883 = ~n33857 & ~n33882;
  assign n33884 = n6273 & ~n33883;
  assign n33885 = ~n6273 & n33855;
  assign n33886 = pi59 & ~n33885;
  assign n33887 = ~n33884 & n33886;
  assign n33888 = pi55 & n33883;
  assign n33889 = ~pi74 & n3275;
  assign n33890 = pi299 & ~n33855;
  assign n33891 = ~pi198 & n33838;
  assign n33892 = n33842 & ~n33891;
  assign n33893 = n6550 & ~n33892;
  assign n33894 = n33831 & ~n33893;
  assign n33895 = pi96 & pi198;
  assign n33896 = pi332 & n33895;
  assign n33897 = ~n33892 & ~n33896;
  assign n33898 = n6185 & ~n33897;
  assign n33899 = ~pi299 & ~n33898;
  assign n33900 = ~n6549 & n33899;
  assign n33901 = ~n33894 & n33900;
  assign n33902 = ~n33890 & ~n33901;
  assign n33903 = ~n33889 & n33902;
  assign n33904 = n2508 & n2715;
  assign n33905 = n33862 & n33904;
  assign n33906 = ~pi70 & ~n33905;
  assign n33907 = n33840 & ~n33906;
  assign n33908 = pi210 & n33907;
  assign n33909 = n33864 & n33904;
  assign n33910 = ~n33838 & ~n33909;
  assign n33911 = ~pi210 & ~n33910;
  assign n33912 = ~pi332 & ~n33911;
  assign n33913 = ~n33908 & n33912;
  assign n33914 = ~n33834 & ~n33913;
  assign n33915 = n6185 & ~n33914;
  assign n33916 = ~pi468 & ~n33913;
  assign n33917 = ~n33850 & ~n33916;
  assign n33918 = ~n6185 & n33917;
  assign n33919 = ~n33915 & ~n33918;
  assign n33920 = pi947 & n33919;
  assign n33921 = ~n6190 & n33914;
  assign n33922 = n6185 & ~n33921;
  assign n33923 = n33832 & ~n33922;
  assign n33924 = pi299 & ~n33923;
  assign n33925 = ~n33920 & n33924;
  assign n33926 = pi198 & n33907;
  assign n33927 = ~pi198 & ~n33910;
  assign n33928 = ~pi332 & ~n33927;
  assign n33929 = ~n33926 & n33928;
  assign n33930 = ~n33896 & ~n33929;
  assign n33931 = n6185 & ~n33930;
  assign n33932 = ~pi468 & ~n33929;
  assign n33933 = ~n6185 & ~n33850;
  assign n33934 = ~n33932 & n33933;
  assign n33935 = ~n33931 & ~n33934;
  assign n33936 = pi587 & n33935;
  assign n33937 = ~pi587 & ~n33831;
  assign n33938 = ~n6190 & n33930;
  assign n33939 = n6185 & ~n33938;
  assign n33940 = n33937 & ~n33939;
  assign n33941 = ~pi299 & ~n33940;
  assign n33942 = ~n33936 & n33941;
  assign n33943 = ~n33925 & ~n33942;
  assign n33944 = n9985 & ~n33943;
  assign n33945 = pi198 & n33860;
  assign n33946 = ~pi198 & ~n33867;
  assign n33947 = ~pi332 & ~n33946;
  assign n33948 = ~n33945 & n33947;
  assign n33949 = ~n33896 & ~n33948;
  assign n33950 = ~n6190 & n33949;
  assign n33951 = n6185 & ~n33950;
  assign n33952 = n33937 & ~n33951;
  assign n33953 = ~pi468 & ~n33948;
  assign n33954 = n33933 & ~n33953;
  assign n33955 = n6185 & ~n33949;
  assign n33956 = pi587 & ~n33955;
  assign n33957 = ~n33954 & n33956;
  assign n33958 = ~n33952 & ~n33957;
  assign n33959 = ~pi299 & ~n33958;
  assign n33960 = pi299 & ~n33881;
  assign n33961 = n15135 & ~n33960;
  assign n33962 = ~n33959 & n33961;
  assign n33963 = ~n33944 & ~n33962;
  assign n33964 = ~pi74 & ~n33963;
  assign n33965 = ~pi55 & ~n33964;
  assign n33966 = ~n33903 & n33965;
  assign n33967 = n2531 & ~n33966;
  assign n33968 = ~n33888 & n33967;
  assign n33969 = ~n2531 & n33855;
  assign n33970 = ~pi59 & ~n33969;
  assign n33971 = ~n33968 & n33970;
  assign n33972 = ~n33887 & ~n33971;
  assign n33973 = ~pi57 & ~n33972;
  assign n33974 = ~n33856 & ~n33973;
  assign n33975 = n33830 & ~n33974;
  assign n33976 = pi57 & pi332;
  assign n33977 = pi332 & ~n2531;
  assign n33978 = ~pi59 & ~n33977;
  assign n33979 = pi74 & pi332;
  assign n33980 = ~pi55 & ~n33979;
  assign n33981 = n2715 & n10879;
  assign n33982 = pi468 & ~n6185;
  assign n33983 = ~pi299 & pi587;
  assign n33984 = ~pi468 & ~n33983;
  assign n33985 = ~n20462 & n33984;
  assign n33986 = ~n33982 & ~n33985;
  assign n33987 = n33981 & n33986;
  assign n33988 = ~pi332 & ~n33987;
  assign n33989 = n9985 & ~n33988;
  assign n33990 = n2522 & n6552;
  assign n33991 = ~pi332 & ~n33990;
  assign n33992 = n15135 & ~n33991;
  assign n33993 = pi332 & ~n3275;
  assign n33994 = ~n33992 & ~n33993;
  assign n33995 = ~n33989 & n33994;
  assign n33996 = ~pi74 & ~n33995;
  assign n33997 = n33980 & ~n33996;
  assign n33998 = n2522 & n6542;
  assign n33999 = n2576 & n33998;
  assign n34000 = ~pi332 & ~n33999;
  assign n34001 = pi55 & n34000;
  assign n34002 = ~n33997 & ~n34001;
  assign n34003 = n2531 & n34002;
  assign n34004 = n33978 & ~n34003;
  assign n34005 = n6273 & ~n34000;
  assign n34006 = pi332 & ~n6273;
  assign n34007 = pi59 & ~n34006;
  assign n34008 = ~n34005 & n34007;
  assign n34009 = ~pi57 & ~n34008;
  assign n34010 = ~n34004 & n34009;
  assign n34011 = ~n33976 & ~n34010;
  assign n34012 = ~n33830 & ~n34011;
  assign n34013 = ~n33975 & ~n34012;
  assign n34014 = ~pi201 & ~n34013;
  assign n34015 = ~n6542 & ~n15973;
  assign n34016 = n6551 & ~po1038;
  assign n34017 = ~n34015 & ~n34016;
  assign n34018 = n15973 & ~n33895;
  assign n34019 = ~n15973 & ~n33833;
  assign n34020 = ~n34018 & ~n34019;
  assign n34021 = n34017 & n34020;
  assign n34022 = n33830 & n34021;
  assign n34023 = pi201 & ~n34022;
  assign po358 = ~n34014 & ~n34023;
  assign n34025 = ~pi233 & pi237;
  assign n34026 = ~n33974 & n34025;
  assign n34027 = ~n34011 & ~n34025;
  assign n34028 = ~n34026 & ~n34027;
  assign n34029 = ~pi202 & ~n34028;
  assign n34030 = n34021 & n34025;
  assign n34031 = pi202 & ~n34030;
  assign po359 = ~n34029 & ~n34031;
  assign n34033 = ~pi233 & ~pi237;
  assign n34034 = ~n33974 & n34033;
  assign n34035 = ~n34011 & ~n34033;
  assign n34036 = ~n34034 & ~n34035;
  assign n34037 = ~pi203 & ~n34036;
  assign n34038 = n34021 & n34033;
  assign n34039 = pi203 & ~n34038;
  assign po360 = ~n34037 & ~n34039;
  assign n34041 = ~pi332 & ~n6188;
  assign n34042 = ~pi907 & ~n34041;
  assign n34043 = n6188 & ~n33845;
  assign n34044 = n34042 & ~n34043;
  assign n34045 = ~n6188 & n33852;
  assign n34046 = n6188 & ~n33844;
  assign n34047 = pi907 & ~n34046;
  assign n34048 = ~n34045 & n34047;
  assign n34049 = ~n34044 & ~n34048;
  assign n34050 = pi57 & ~n34049;
  assign n34051 = ~n2576 & n34049;
  assign n34052 = ~n6188 & n33878;
  assign n34053 = n6188 & ~n33871;
  assign n34054 = pi907 & ~n34053;
  assign n34055 = ~n34052 & n34054;
  assign n34056 = pi332 & ~n6187;
  assign n34057 = ~n33872 & ~n34056;
  assign n34058 = pi680 & n34057;
  assign n34059 = n34042 & ~n34058;
  assign n34060 = ~n34055 & ~n34059;
  assign n34061 = n2576 & n34060;
  assign n34062 = ~n34051 & ~n34061;
  assign n34063 = n6273 & ~n34062;
  assign n34064 = ~n6273 & n34049;
  assign n34065 = pi59 & ~n34064;
  assign n34066 = ~n34063 & n34065;
  assign n34067 = pi55 & n34062;
  assign n34068 = n6188 & n33895;
  assign n34069 = pi332 & ~n34068;
  assign n34070 = ~pi468 & pi602;
  assign n34071 = pi468 & n6188;
  assign n34072 = ~n34070 & ~n34071;
  assign n34073 = n33897 & ~n34072;
  assign n34074 = ~n34069 & ~n34073;
  assign n34075 = ~pi299 & ~n34074;
  assign n34076 = pi299 & ~n34049;
  assign n34077 = ~n33889 & ~n34076;
  assign n34078 = ~n34075 & n34077;
  assign n34079 = pi299 & n34060;
  assign n34080 = ~pi299 & ~n34069;
  assign n34081 = n6291 & n33949;
  assign n34082 = n34080 & ~n34081;
  assign n34083 = ~n34079 & ~n34082;
  assign n34084 = n15135 & ~n34083;
  assign n34085 = n6291 & n33930;
  assign n34086 = n34080 & ~n34085;
  assign n34087 = n6188 & ~n33914;
  assign n34088 = ~n6188 & n33917;
  assign n34089 = ~n34087 & ~n34088;
  assign n34090 = pi907 & n34089;
  assign n34091 = n6188 & ~n33921;
  assign n34092 = n34042 & ~n34091;
  assign n34093 = pi299 & ~n34092;
  assign n34094 = ~n34090 & n34093;
  assign n34095 = ~n34086 & ~n34094;
  assign n34096 = n9985 & ~n34095;
  assign n34097 = ~n34084 & ~n34096;
  assign n34098 = ~pi74 & ~n34097;
  assign n34099 = ~pi55 & ~n34098;
  assign n34100 = ~n34078 & n34099;
  assign n34101 = n2531 & ~n34100;
  assign n34102 = ~n34067 & n34101;
  assign n34103 = ~n2531 & n34049;
  assign n34104 = ~pi59 & ~n34103;
  assign n34105 = ~n34102 & n34104;
  assign n34106 = ~n34066 & ~n34105;
  assign n34107 = ~pi57 & ~n34106;
  assign n34108 = ~n34050 & ~n34107;
  assign n34109 = n33830 & ~n34108;
  assign n34110 = n2522 & n6279;
  assign n34111 = n2576 & n34110;
  assign n34112 = ~pi332 & ~n34111;
  assign n34113 = pi55 & n34112;
  assign n34114 = ~pi299 & ~n34072;
  assign n34115 = ~n6289 & ~n34114;
  assign n34116 = n2522 & ~n34115;
  assign n34117 = ~pi332 & ~n34116;
  assign n34118 = n15135 & ~n34117;
  assign n34119 = pi299 & ~pi907;
  assign n34120 = ~pi299 & ~pi602;
  assign n34121 = ~pi468 & ~n34120;
  assign n34122 = ~n34119 & n34121;
  assign n34123 = ~n34071 & ~n34122;
  assign n34124 = n33981 & ~n34123;
  assign n34125 = ~pi332 & ~n34124;
  assign n34126 = n9985 & ~n34125;
  assign n34127 = ~n34118 & ~n34126;
  assign n34128 = ~pi74 & ~n34127;
  assign n34129 = ~n33993 & ~n34128;
  assign n34130 = n33980 & n34129;
  assign n34131 = ~n34113 & ~n34130;
  assign n34132 = n2531 & n34131;
  assign n34133 = n33978 & ~n34132;
  assign n34134 = n6273 & ~n34112;
  assign n34135 = n34007 & ~n34134;
  assign n34136 = ~pi57 & ~n34135;
  assign n34137 = ~n34133 & n34136;
  assign n34138 = ~n33976 & ~n34137;
  assign n34139 = ~n33830 & ~n34138;
  assign n34140 = ~n34109 & ~n34139;
  assign n34141 = ~pi204 & ~n34140;
  assign n34142 = n6279 & ~n15973;
  assign n34143 = n6291 & n15973;
  assign n34144 = ~n34142 & ~n34143;
  assign n34145 = n34020 & ~n34144;
  assign n34146 = n33830 & n34145;
  assign n34147 = pi204 & ~n34146;
  assign po361 = ~n34141 & ~n34147;
  assign n34149 = n34025 & ~n34108;
  assign n34150 = ~n34025 & ~n34138;
  assign n34151 = ~n34149 & ~n34150;
  assign n34152 = ~pi205 & ~n34151;
  assign n34153 = n34025 & n34145;
  assign n34154 = pi205 & ~n34153;
  assign po362 = ~n34152 & ~n34154;
  assign n34156 = pi233 & ~pi237;
  assign n34157 = ~n34108 & n34156;
  assign n34158 = ~n34138 & ~n34156;
  assign n34159 = ~n34157 & ~n34158;
  assign n34160 = ~pi206 & ~n34159;
  assign n34161 = n34145 & n34156;
  assign n34162 = pi206 & ~n34161;
  assign po363 = ~n34160 & ~n34162;
  assign n34164 = n16521 & ~n16527;
  assign n34165 = n10020 & n18808;
  assign n34166 = ~n16521 & ~n34165;
  assign n34167 = ~n34164 & ~n34166;
  assign n34168 = ~pi785 & ~n34167;
  assign n34169 = ~n16527 & ~n16537;
  assign n34170 = ~pi609 & n34166;
  assign n34171 = ~n34169 & ~n34170;
  assign n34172 = ~pi1155 & ~n34171;
  assign n34173 = ~n16527 & ~n16532;
  assign n34174 = pi609 & n34166;
  assign n34175 = ~n34173 & ~n34174;
  assign n34176 = pi1155 & ~n34175;
  assign n34177 = ~n34172 & ~n34176;
  assign n34178 = pi785 & ~n34177;
  assign n34179 = ~n34168 & ~n34178;
  assign n34180 = ~pi781 & ~n34179;
  assign n34181 = ~pi618 & n34179;
  assign n34182 = pi618 & n16527;
  assign n34183 = ~pi1154 & ~n34182;
  assign n34184 = ~n34181 & n34183;
  assign n34185 = pi618 & n34179;
  assign n34186 = ~pi618 & n16527;
  assign n34187 = pi1154 & ~n34186;
  assign n34188 = ~n34185 & n34187;
  assign n34189 = ~n34184 & ~n34188;
  assign n34190 = pi781 & ~n34189;
  assign n34191 = ~n34180 & ~n34190;
  assign n34192 = ~pi789 & ~n34191;
  assign n34193 = ~pi619 & n34191;
  assign n34194 = pi619 & n16527;
  assign n34195 = ~pi1159 & ~n34194;
  assign n34196 = ~n34193 & n34195;
  assign n34197 = pi619 & n34191;
  assign n34198 = ~pi619 & n16527;
  assign n34199 = pi1159 & ~n34198;
  assign n34200 = ~n34197 & n34199;
  assign n34201 = ~n34196 & ~n34200;
  assign n34202 = pi789 & ~n34201;
  assign n34203 = ~n34192 & ~n34202;
  assign n34204 = ~n17355 & n34203;
  assign n34205 = n16527 & n17355;
  assign n34206 = ~n34204 & ~n34205;
  assign n34207 = ~n16124 & ~n34206;
  assign n34208 = n16124 & n16527;
  assign n34209 = ~n34207 & ~n34208;
  assign n34210 = ~pi207 & n34209;
  assign n34211 = n10020 & ~n23777;
  assign n34212 = ~n16521 & n34211;
  assign n34213 = ~n19656 & n34212;
  assign n34214 = ~n19662 & n34213;
  assign n34215 = ~n19667 & n34214;
  assign n34216 = ~n17355 & n34215;
  assign n34217 = ~n16124 & n34216;
  assign n34218 = pi207 & n34217;
  assign n34219 = ~n34210 & ~n34218;
  assign n34220 = pi623 & ~n34219;
  assign n34221 = ~pi207 & ~n16527;
  assign n34222 = ~pi623 & n34221;
  assign n34223 = ~n34220 & ~n34222;
  assign n34224 = ~n19987 & n34223;
  assign n34225 = ~n18633 & n23734;
  assign n34226 = n18717 & n34225;
  assign n34227 = ~n18744 & n34226;
  assign n34228 = pi207 & ~n34227;
  assign n34229 = ~n16527 & n17159;
  assign n34230 = ~n16527 & n16593;
  assign n34231 = n10020 & n23737;
  assign n34232 = ~pi778 & ~n34231;
  assign n34233 = ~pi625 & ~n16527;
  assign n34234 = pi625 & ~n34231;
  assign n34235 = ~n34233 & ~n34234;
  assign n34236 = pi1153 & ~n34235;
  assign n34237 = pi625 & ~n16527;
  assign n34238 = ~pi625 & ~n34231;
  assign n34239 = ~n34237 & ~n34238;
  assign n34240 = ~pi1153 & ~n34239;
  assign n34241 = ~n34236 & ~n34240;
  assign n34242 = pi778 & ~n34241;
  assign n34243 = ~n34232 & ~n34242;
  assign n34244 = ~n16593 & ~n34243;
  assign n34245 = ~n34230 & ~n34244;
  assign n34246 = ~n16589 & n34245;
  assign n34247 = n16527 & n16589;
  assign n34248 = ~n34246 & ~n34247;
  assign n34249 = ~n17159 & n34248;
  assign n34250 = ~n34229 & ~n34249;
  assign n34251 = ~n17183 & n34250;
  assign n34252 = n16527 & n17183;
  assign n34253 = ~n34251 & ~n34252;
  assign n34254 = ~n18744 & ~n34253;
  assign n34255 = n16527 & n17451;
  assign n34256 = ~n34254 & ~n34255;
  assign n34257 = ~pi207 & ~n34256;
  assign n34258 = ~n34228 & ~n34257;
  assign n34259 = pi710 & ~n34258;
  assign n34260 = ~pi710 & ~n34221;
  assign n34261 = ~n34259 & ~n34260;
  assign n34262 = ~pi647 & n34261;
  assign n34263 = pi647 & n34221;
  assign n34264 = ~pi1157 & ~n34263;
  assign n34265 = ~n34262 & n34264;
  assign n34266 = pi647 & n34261;
  assign n34267 = pi1157 & ~n34266;
  assign n34268 = ~pi647 & n34221;
  assign n34269 = n34267 & ~n34268;
  assign n34270 = ~n34265 & ~n34269;
  assign n34271 = ~n17246 & ~n34270;
  assign n34272 = ~n34224 & ~n34271;
  assign n34273 = pi787 & ~n34272;
  assign n34274 = pi1156 & ~n34216;
  assign n34275 = ~pi1156 & ~n34226;
  assign n34276 = n19995 & ~n34275;
  assign n34277 = ~n34274 & n34276;
  assign n34278 = ~pi1156 & ~n34216;
  assign n34279 = pi1156 & ~n34226;
  assign n34280 = n19997 & ~n34279;
  assign n34281 = ~n34278 & n34280;
  assign n34282 = ~n34277 & ~n34281;
  assign n34283 = pi792 & ~n34282;
  assign n34284 = n17347 & n34215;
  assign n34285 = ~pi1158 & ~n34284;
  assign n34286 = n18715 & n34225;
  assign n34287 = ~pi1159 & ~n34286;
  assign n34288 = pi1159 & ~n34214;
  assign n34289 = pi619 & ~n34288;
  assign n34290 = ~pi648 & n34289;
  assign n34291 = ~n34287 & n34290;
  assign n34292 = pi1159 & ~n34286;
  assign n34293 = ~pi1159 & ~n34214;
  assign n34294 = pi648 & ~n34293;
  assign n34295 = ~pi619 & n34294;
  assign n34296 = ~n34292 & n34295;
  assign n34297 = ~n34291 & ~n34296;
  assign n34298 = pi789 & ~n34297;
  assign n34299 = ~pi778 & ~n33367;
  assign n34300 = ~pi625 & n23734;
  assign n34301 = ~pi1153 & ~n34300;
  assign n34302 = pi608 & ~n34301;
  assign n34303 = ~pi625 & n34211;
  assign n34304 = pi625 & n33367;
  assign n34305 = ~n34303 & ~n34304;
  assign n34306 = pi1153 & n34305;
  assign n34307 = n34302 & ~n34306;
  assign n34308 = pi625 & n23734;
  assign n34309 = pi1153 & ~n34308;
  assign n34310 = ~pi608 & ~n34309;
  assign n34311 = ~pi625 & n33367;
  assign n34312 = pi625 & n34211;
  assign n34313 = ~pi1153 & ~n34312;
  assign n34314 = ~n34311 & n34313;
  assign n34315 = n34310 & ~n34314;
  assign n34316 = ~n34307 & ~n34315;
  assign n34317 = pi778 & n34316;
  assign n34318 = ~n34299 & ~n34317;
  assign n34319 = ~pi785 & ~n34318;
  assign n34320 = ~pi609 & ~n34318;
  assign n34321 = pi609 & ~n34225;
  assign n34322 = ~pi1155 & ~n34321;
  assign n34323 = ~n34320 & n34322;
  assign n34324 = n19653 & n34212;
  assign n34325 = ~pi660 & ~n34324;
  assign n34326 = ~n34323 & n34325;
  assign n34327 = pi609 & ~n34318;
  assign n34328 = ~pi609 & ~n34225;
  assign n34329 = pi1155 & ~n34328;
  assign n34330 = ~n34327 & n34329;
  assign n34331 = n19654 & n34212;
  assign n34332 = pi660 & ~n34331;
  assign n34333 = ~n34330 & n34332;
  assign n34334 = ~n34326 & ~n34333;
  assign n34335 = pi785 & ~n34334;
  assign n34336 = ~n34319 & ~n34335;
  assign n34337 = pi618 & ~n34336;
  assign n34338 = ~n16593 & n34225;
  assign n34339 = ~pi618 & ~n34338;
  assign n34340 = pi1154 & ~n34339;
  assign n34341 = ~n34337 & n34340;
  assign n34342 = n19660 & n34213;
  assign n34343 = pi627 & ~n34342;
  assign n34344 = ~n34341 & n34343;
  assign n34345 = pi618 & ~n34338;
  assign n34346 = ~pi1154 & ~n34345;
  assign n34347 = n19659 & n34213;
  assign n34348 = ~pi627 & ~n34347;
  assign n34349 = ~n34346 & n34348;
  assign n34350 = ~n34344 & ~n34349;
  assign n34351 = pi781 & ~n34350;
  assign n34352 = ~pi618 & ~pi627;
  assign n34353 = pi781 & ~n34352;
  assign n34354 = ~n34336 & ~n34353;
  assign n34355 = ~n34351 & ~n34354;
  assign n34356 = n22991 & n34355;
  assign n34357 = ~n34298 & ~n34356;
  assign n34358 = ~pi626 & n34357;
  assign n34359 = ~n17159 & n34286;
  assign n34360 = pi626 & ~n34359;
  assign n34361 = ~pi641 & ~n34360;
  assign n34362 = ~n34358 & n34361;
  assign n34363 = n34285 & ~n34362;
  assign n34364 = n17348 & n34215;
  assign n34365 = pi1158 & ~n34364;
  assign n34366 = ~pi626 & ~n34359;
  assign n34367 = pi626 & n34357;
  assign n34368 = ~n34366 & ~n34367;
  assign n34369 = pi641 & n34368;
  assign n34370 = n34365 & ~n34369;
  assign n34371 = ~n34363 & ~n34370;
  assign n34372 = pi788 & ~n34371;
  assign n34373 = ~pi788 & n34357;
  assign n34374 = n19788 & ~n34373;
  assign n34375 = ~n34372 & n34374;
  assign n34376 = ~n34283 & ~n34375;
  assign n34377 = pi207 & ~n34376;
  assign n34378 = ~n19999 & n34206;
  assign n34379 = ~pi628 & ~n34253;
  assign n34380 = n16122 & ~n34379;
  assign n34381 = pi628 & n16527;
  assign n34382 = n34380 & ~n34381;
  assign n34383 = ~n34378 & ~n34382;
  assign n34384 = ~pi628 & ~n16527;
  assign n34385 = pi628 & n34253;
  assign n34386 = ~n34384 & ~n34385;
  assign n34387 = ~pi629 & ~n34386;
  assign n34388 = pi1156 & n34387;
  assign n34389 = n34383 & ~n34388;
  assign n34390 = pi792 & ~n34389;
  assign n34391 = pi618 & ~n34245;
  assign n34392 = pi609 & ~n34243;
  assign n34393 = n10020 & n18914;
  assign n34394 = ~pi778 & ~n34393;
  assign n34395 = ~pi608 & ~n34236;
  assign n34396 = pi625 & n34165;
  assign n34397 = ~pi625 & n34393;
  assign n34398 = ~pi1153 & ~n34397;
  assign n34399 = ~n34396 & n34398;
  assign n34400 = n34395 & ~n34399;
  assign n34401 = pi608 & ~n34240;
  assign n34402 = ~pi625 & n34165;
  assign n34403 = pi625 & n34393;
  assign n34404 = ~n34402 & ~n34403;
  assign n34405 = pi1153 & n34404;
  assign n34406 = n34401 & ~n34405;
  assign n34407 = ~n34400 & ~n34406;
  assign n34408 = pi778 & n34407;
  assign n34409 = ~n34394 & ~n34408;
  assign n34410 = ~pi609 & ~n34409;
  assign n34411 = ~n34392 & ~n34410;
  assign n34412 = ~pi1155 & ~n34411;
  assign n34413 = ~pi660 & ~n34176;
  assign n34414 = ~n34412 & n34413;
  assign n34415 = ~pi609 & ~n34243;
  assign n34416 = pi609 & ~n34409;
  assign n34417 = ~n34415 & ~n34416;
  assign n34418 = pi1155 & ~n34417;
  assign n34419 = ~n34172 & ~n34418;
  assign n34420 = pi660 & n34419;
  assign n34421 = ~n34414 & ~n34420;
  assign n34422 = pi785 & ~n34421;
  assign n34423 = ~pi785 & n34409;
  assign n34424 = ~n34422 & ~n34423;
  assign n34425 = ~pi618 & n34424;
  assign n34426 = ~n34391 & ~n34425;
  assign n34427 = ~pi1154 & ~n34426;
  assign n34428 = ~pi627 & ~n34188;
  assign n34429 = ~n34427 & n34428;
  assign n34430 = ~pi618 & ~n34245;
  assign n34431 = pi618 & n34424;
  assign n34432 = ~n34430 & ~n34431;
  assign n34433 = pi1154 & ~n34432;
  assign n34434 = ~n34184 & ~n34433;
  assign n34435 = pi627 & n34434;
  assign n34436 = ~n34429 & ~n34435;
  assign n34437 = pi781 & ~n34436;
  assign n34438 = ~pi781 & ~n34424;
  assign n34439 = ~n34437 & ~n34438;
  assign n34440 = ~pi789 & n34439;
  assign n34441 = pi619 & n34248;
  assign n34442 = ~pi619 & n34439;
  assign n34443 = ~n34441 & ~n34442;
  assign n34444 = ~pi1159 & ~n34443;
  assign n34445 = ~pi648 & ~n34444;
  assign n34446 = ~n34200 & n34445;
  assign n34447 = ~pi619 & n34248;
  assign n34448 = pi619 & n34439;
  assign n34449 = ~n34447 & ~n34448;
  assign n34450 = pi1159 & ~n34449;
  assign n34451 = ~n34196 & ~n34450;
  assign n34452 = pi648 & n34451;
  assign n34453 = ~n34446 & ~n34452;
  assign n34454 = pi789 & n34453;
  assign n34455 = ~n34440 & ~n34454;
  assign n34456 = n17356 & n34455;
  assign n34457 = ~n17182 & ~n17349;
  assign n34458 = n34203 & n34457;
  assign n34459 = ~pi641 & ~n34250;
  assign n34460 = pi641 & ~n16527;
  assign n34461 = n17345 & ~n34460;
  assign n34462 = ~n34459 & n34461;
  assign n34463 = ~pi641 & ~n16527;
  assign n34464 = pi641 & ~n34250;
  assign n34465 = ~n34463 & ~n34464;
  assign n34466 = n17344 & n34465;
  assign n34467 = ~n34462 & ~n34466;
  assign n34468 = ~n34458 & n34467;
  assign n34469 = pi788 & ~n34468;
  assign n34470 = n19788 & ~n34469;
  assign n34471 = ~n34456 & n34470;
  assign n34472 = ~n34390 & ~n34471;
  assign n34473 = ~pi207 & ~n34472;
  assign n34474 = pi623 & ~n34473;
  assign n34475 = ~n34377 & n34474;
  assign n34476 = ~pi778 & ~n33361;
  assign n34477 = pi625 & n33361;
  assign n34478 = pi1153 & ~n34477;
  assign n34479 = n34302 & ~n34478;
  assign n34480 = ~pi625 & n33361;
  assign n34481 = ~pi1153 & ~n34480;
  assign n34482 = n34310 & ~n34481;
  assign n34483 = ~n34479 & ~n34482;
  assign n34484 = pi778 & n34483;
  assign n34485 = ~n34476 & ~n34484;
  assign n34486 = ~pi609 & ~n34485;
  assign n34487 = ~pi660 & n34322;
  assign n34488 = ~n34486 & n34487;
  assign n34489 = pi609 & ~n34485;
  assign n34490 = pi660 & ~n34489;
  assign n34491 = n34329 & n34490;
  assign n34492 = ~n34488 & ~n34491;
  assign n34493 = pi785 & ~n34492;
  assign n34494 = ~pi785 & n34485;
  assign n34495 = ~n34493 & ~n34494;
  assign n34496 = ~pi618 & n34495;
  assign n34497 = n16586 & ~n34496;
  assign n34498 = ~n34345 & n34497;
  assign n34499 = pi618 & n34495;
  assign n34500 = pi627 & ~n34499;
  assign n34501 = n34340 & n34500;
  assign n34502 = ~n34498 & ~n34501;
  assign n34503 = pi781 & n34502;
  assign n34504 = ~pi781 & n34495;
  assign n34505 = n22991 & ~n34504;
  assign n34506 = ~n34503 & n34505;
  assign n34507 = n17158 & n19667;
  assign n34508 = n34286 & n34507;
  assign n34509 = ~n34506 & ~n34508;
  assign n34510 = ~pi626 & n34509;
  assign n34511 = n17153 & ~n34360;
  assign n34512 = ~n34510 & n34511;
  assign n34513 = pi626 & n34509;
  assign n34514 = ~n34366 & ~n34513;
  assign n34515 = n17167 & n34514;
  assign n34516 = ~n34512 & ~n34515;
  assign n34517 = pi788 & n34516;
  assign n34518 = ~pi788 & n34509;
  assign n34519 = n19788 & ~n34518;
  assign n34520 = ~n34517 & n34519;
  assign n34521 = n16124 & n17450;
  assign n34522 = n34226 & n34521;
  assign n34523 = ~n34520 & ~n34522;
  assign n34524 = pi207 & ~n34523;
  assign n34525 = ~n34384 & ~n34387;
  assign n34526 = pi1156 & ~n34525;
  assign n34527 = n17449 & ~n34381;
  assign n34528 = ~n34382 & ~n34527;
  assign n34529 = ~n34526 & n34528;
  assign n34530 = pi792 & ~n34529;
  assign n34531 = pi626 & n34250;
  assign n34532 = n10020 & ~n18939;
  assign n34533 = ~pi778 & ~n34532;
  assign n34534 = pi625 & ~n34532;
  assign n34535 = ~n34233 & ~n34534;
  assign n34536 = pi1153 & ~n34535;
  assign n34537 = n34401 & ~n34536;
  assign n34538 = ~pi625 & ~n34532;
  assign n34539 = ~n34237 & ~n34538;
  assign n34540 = ~pi1153 & ~n34539;
  assign n34541 = n34395 & ~n34540;
  assign n34542 = ~n34537 & ~n34541;
  assign n34543 = pi778 & n34542;
  assign n34544 = ~n34533 & ~n34543;
  assign n34545 = ~pi609 & ~n34544;
  assign n34546 = ~n34392 & ~n34545;
  assign n34547 = ~pi1155 & ~n34546;
  assign n34548 = pi1155 & ~n16527;
  assign n34549 = ~pi660 & ~n34548;
  assign n34550 = ~n34547 & n34549;
  assign n34551 = pi609 & ~n34544;
  assign n34552 = ~n34415 & ~n34551;
  assign n34553 = pi1155 & ~n34552;
  assign n34554 = ~pi1155 & ~n16527;
  assign n34555 = pi660 & ~n34554;
  assign n34556 = ~n34553 & n34555;
  assign n34557 = ~n34550 & ~n34556;
  assign n34558 = pi785 & ~n34557;
  assign n34559 = ~pi785 & n34544;
  assign n34560 = ~n34558 & ~n34559;
  assign n34561 = ~pi618 & n34560;
  assign n34562 = ~n34391 & ~n34561;
  assign n34563 = ~pi1154 & ~n34562;
  assign n34564 = pi1154 & ~n16527;
  assign n34565 = ~pi627 & ~n34564;
  assign n34566 = ~n34563 & n34565;
  assign n34567 = pi618 & n34560;
  assign n34568 = ~n34430 & ~n34567;
  assign n34569 = pi1154 & ~n34568;
  assign n34570 = ~pi1154 & ~n16527;
  assign n34571 = pi627 & ~n34570;
  assign n34572 = ~n34569 & n34571;
  assign n34573 = ~n34566 & ~n34572;
  assign n34574 = pi781 & ~n34573;
  assign n34575 = ~pi781 & ~n34560;
  assign n34576 = ~n34574 & ~n34575;
  assign n34577 = ~pi619 & n34576;
  assign n34578 = ~n34441 & ~n34577;
  assign n34579 = ~pi1159 & ~n34578;
  assign n34580 = pi1159 & ~n16527;
  assign n34581 = ~pi648 & ~n34580;
  assign n34582 = ~n34579 & n34581;
  assign n34583 = pi619 & n34576;
  assign n34584 = ~n34447 & ~n34583;
  assign n34585 = pi1159 & ~n34584;
  assign n34586 = ~pi1159 & ~n16527;
  assign n34587 = pi648 & ~n34586;
  assign n34588 = ~n34585 & n34587;
  assign n34589 = ~n34582 & ~n34588;
  assign n34590 = pi789 & ~n34589;
  assign n34591 = ~pi789 & ~n34576;
  assign n34592 = ~n34590 & ~n34591;
  assign n34593 = ~pi626 & ~n34592;
  assign n34594 = ~pi641 & ~n34593;
  assign n34595 = ~n34531 & n34594;
  assign n34596 = ~pi1158 & ~n34460;
  assign n34597 = ~n34595 & n34596;
  assign n34598 = ~pi626 & n34250;
  assign n34599 = pi626 & ~n34592;
  assign n34600 = ~n34598 & ~n34599;
  assign n34601 = pi641 & n34600;
  assign n34602 = ~n34463 & ~n34601;
  assign n34603 = pi1158 & n34602;
  assign n34604 = ~n34597 & ~n34603;
  assign n34605 = pi788 & ~n34604;
  assign n34606 = ~pi788 & ~n34592;
  assign n34607 = n19788 & ~n34606;
  assign n34608 = ~n34605 & n34607;
  assign n34609 = ~n34530 & ~n34608;
  assign n34610 = ~pi207 & ~n34609;
  assign n34611 = ~pi623 & ~n34610;
  assign n34612 = ~n34524 & n34611;
  assign n34613 = ~n34475 & ~n34612;
  assign n34614 = pi710 & n34613;
  assign n34615 = ~pi710 & ~n34223;
  assign n34616 = n19637 & ~n34615;
  assign n34617 = ~n34614 & n34616;
  assign n34618 = ~n34273 & ~n34617;
  assign n34619 = pi644 & n34618;
  assign n34620 = ~pi787 & ~n34261;
  assign n34621 = pi787 & ~n34270;
  assign n34622 = ~n34620 & ~n34621;
  assign n34623 = ~pi644 & n34622;
  assign n34624 = pi715 & ~n34623;
  assign n34625 = ~n34619 & n34624;
  assign n34626 = n17247 & ~n34221;
  assign n34627 = ~n17247 & n34223;
  assign n34628 = ~n34626 & ~n34627;
  assign n34629 = pi644 & n34628;
  assign n34630 = ~pi644 & n34221;
  assign n34631 = ~pi715 & ~n34630;
  assign n34632 = ~n34629 & n34631;
  assign n34633 = pi1160 & ~n34632;
  assign n34634 = ~n34625 & n34633;
  assign n34635 = ~pi644 & n34628;
  assign n34636 = pi715 & ~n34635;
  assign n34637 = pi644 & n34221;
  assign n34638 = n34636 & ~n34637;
  assign n34639 = pi644 & n34622;
  assign n34640 = ~pi644 & n34618;
  assign n34641 = ~pi715 & ~n34640;
  assign n34642 = ~n34639 & n34641;
  assign n34643 = ~pi1160 & ~n34642;
  assign n34644 = ~n34638 & n34643;
  assign n34645 = ~n34634 & ~n34644;
  assign n34646 = pi790 & ~n34645;
  assign n34647 = ~pi790 & n34618;
  assign n34648 = ~n34646 & ~n34647;
  assign n34649 = ~po1038 & ~n34648;
  assign n34650 = ~pi207 & po1038;
  assign po364 = n34649 | n34650;
  assign n34652 = ~pi208 & n34209;
  assign n34653 = pi208 & n34217;
  assign n34654 = ~n34652 & ~n34653;
  assign n34655 = pi607 & ~n34654;
  assign n34656 = ~pi208 & ~n16527;
  assign n34657 = ~pi607 & n34656;
  assign n34658 = ~n34655 & ~n34657;
  assign n34659 = ~n19987 & n34658;
  assign n34660 = pi208 & ~n34227;
  assign n34661 = ~pi208 & ~n34256;
  assign n34662 = ~n34660 & ~n34661;
  assign n34663 = pi638 & ~n34662;
  assign n34664 = ~pi638 & ~n34656;
  assign n34665 = ~n34663 & ~n34664;
  assign n34666 = ~pi647 & n34665;
  assign n34667 = pi647 & n34656;
  assign n34668 = ~pi1157 & ~n34667;
  assign n34669 = ~n34666 & n34668;
  assign n34670 = pi647 & n34665;
  assign n34671 = pi1157 & ~n34670;
  assign n34672 = ~pi647 & n34656;
  assign n34673 = n34671 & ~n34672;
  assign n34674 = ~n34669 & ~n34673;
  assign n34675 = ~n17246 & ~n34674;
  assign n34676 = ~n34659 & ~n34675;
  assign n34677 = pi787 & ~n34676;
  assign n34678 = pi208 & ~n34376;
  assign n34679 = ~pi208 & ~n34472;
  assign n34680 = pi607 & ~n34679;
  assign n34681 = ~n34678 & n34680;
  assign n34682 = pi208 & ~n34523;
  assign n34683 = ~pi208 & ~n34609;
  assign n34684 = ~pi607 & ~n34683;
  assign n34685 = ~n34682 & n34684;
  assign n34686 = ~n34681 & ~n34685;
  assign n34687 = pi638 & n34686;
  assign n34688 = ~pi638 & ~n34658;
  assign n34689 = n19637 & ~n34688;
  assign n34690 = ~n34687 & n34689;
  assign n34691 = ~n34677 & ~n34690;
  assign n34692 = pi644 & n34691;
  assign n34693 = ~pi787 & ~n34665;
  assign n34694 = pi787 & ~n34674;
  assign n34695 = ~n34693 & ~n34694;
  assign n34696 = ~pi644 & n34695;
  assign n34697 = pi715 & ~n34696;
  assign n34698 = ~n34692 & n34697;
  assign n34699 = n17247 & ~n34656;
  assign n34700 = ~n17247 & n34658;
  assign n34701 = ~n34699 & ~n34700;
  assign n34702 = pi644 & n34701;
  assign n34703 = ~pi644 & n34656;
  assign n34704 = ~pi715 & ~n34703;
  assign n34705 = ~n34702 & n34704;
  assign n34706 = pi1160 & ~n34705;
  assign n34707 = ~n34698 & n34706;
  assign n34708 = ~pi644 & n34701;
  assign n34709 = pi715 & ~n34708;
  assign n34710 = pi644 & n34656;
  assign n34711 = n34709 & ~n34710;
  assign n34712 = pi644 & n34695;
  assign n34713 = ~pi644 & n34691;
  assign n34714 = ~pi715 & ~n34713;
  assign n34715 = ~n34712 & n34714;
  assign n34716 = ~pi1160 & ~n34715;
  assign n34717 = ~n34711 & n34716;
  assign n34718 = ~n34707 & ~n34717;
  assign n34719 = pi790 & ~n34718;
  assign n34720 = ~pi790 & n34691;
  assign n34721 = ~n34719 & ~n34720;
  assign n34722 = ~po1038 & ~n34721;
  assign n34723 = ~pi208 & po1038;
  assign po365 = n34722 | n34723;
  assign n34725 = n19637 & ~n34609;
  assign n34726 = ~pi647 & ~n16527;
  assign n34727 = pi647 & n34256;
  assign n34728 = ~n34726 & ~n34727;
  assign n34729 = ~pi630 & ~n34728;
  assign n34730 = ~n34726 & ~n34729;
  assign n34731 = pi1157 & ~n34730;
  assign n34732 = pi647 & n16527;
  assign n34733 = n18765 & ~n34732;
  assign n34734 = ~n34731 & ~n34733;
  assign n34735 = ~pi647 & ~n34256;
  assign n34736 = n17245 & ~n34732;
  assign n34737 = ~n34735 & n34736;
  assign n34738 = n34734 & ~n34737;
  assign n34739 = pi787 & ~n34738;
  assign n34740 = ~n34725 & ~n34739;
  assign n34741 = ~pi790 & ~n34740;
  assign n34742 = ~pi644 & ~n34740;
  assign n34743 = ~n18767 & n34256;
  assign n34744 = ~n16527 & n18767;
  assign n34745 = ~n34743 & ~n34744;
  assign n34746 = pi644 & ~n34745;
  assign n34747 = ~pi715 & ~n34746;
  assign n34748 = ~n34742 & n34747;
  assign n34749 = pi715 & n16527;
  assign n34750 = ~pi1160 & ~n34749;
  assign n34751 = ~n34748 & n34750;
  assign n34752 = pi644 & ~n34740;
  assign n34753 = ~pi644 & ~n34745;
  assign n34754 = pi715 & ~n34753;
  assign n34755 = ~n34752 & n34754;
  assign n34756 = ~pi715 & n16527;
  assign n34757 = pi1160 & ~n34756;
  assign n34758 = ~n34755 & n34757;
  assign n34759 = ~n34751 & ~n34758;
  assign n34760 = pi790 & ~n34759;
  assign n34761 = ~po1038 & ~n34760;
  assign n34762 = ~n34741 & n34761;
  assign n34763 = pi639 & n34762;
  assign n34764 = ~pi622 & ~n34763;
  assign n34765 = ~po1038 & n16527;
  assign n34766 = ~pi639 & n34765;
  assign n34767 = n34764 & ~n34766;
  assign n34768 = n19637 & ~n34472;
  assign n34769 = ~n19987 & n34209;
  assign n34770 = pi1157 & n34729;
  assign n34771 = ~n34769 & ~n34770;
  assign n34772 = ~n34737 & n34771;
  assign n34773 = pi787 & ~n34772;
  assign n34774 = ~n34768 & ~n34773;
  assign n34775 = ~pi790 & ~n34774;
  assign n34776 = ~pi644 & ~n34774;
  assign n34777 = n34747 & ~n34776;
  assign n34778 = pi644 & ~n16527;
  assign n34779 = ~n16527 & n17247;
  assign n34780 = ~n17247 & n34209;
  assign n34781 = ~n34779 & ~n34780;
  assign n34782 = ~pi644 & ~n34781;
  assign n34783 = ~n34778 & ~n34782;
  assign n34784 = pi715 & n34783;
  assign n34785 = ~pi1160 & ~n34784;
  assign n34786 = ~n34777 & n34785;
  assign n34787 = pi644 & ~n34774;
  assign n34788 = n34754 & ~n34787;
  assign n34789 = ~pi644 & ~n16527;
  assign n34790 = pi644 & ~n34781;
  assign n34791 = ~n34789 & ~n34790;
  assign n34792 = ~pi715 & n34791;
  assign n34793 = pi1160 & ~n34792;
  assign n34794 = ~n34788 & n34793;
  assign n34795 = ~n34786 & ~n34794;
  assign n34796 = pi790 & ~n34795;
  assign n34797 = ~po1038 & ~n34796;
  assign n34798 = ~n34775 & n34797;
  assign n34799 = pi639 & n34798;
  assign n34800 = ~pi790 & ~n34781;
  assign n34801 = ~po1038 & ~n34800;
  assign n34802 = pi1160 & n34791;
  assign n34803 = ~pi1160 & n34783;
  assign n34804 = ~n34802 & ~n34803;
  assign n34805 = pi790 & n34804;
  assign n34806 = n34801 & ~n34805;
  assign n34807 = ~pi639 & n34806;
  assign n34808 = pi622 & ~n34807;
  assign n34809 = ~n34799 & n34808;
  assign n34810 = ~n34767 & ~n34809;
  assign n34811 = ~pi209 & ~n34810;
  assign n34812 = n19637 & ~n34523;
  assign n34813 = n17247 & n18766;
  assign n34814 = n34227 & n34813;
  assign n34815 = ~n34812 & ~n34814;
  assign n34816 = ~pi790 & n34815;
  assign n34817 = ~po1038 & ~n34816;
  assign n34818 = pi644 & n34815;
  assign n34819 = ~n18767 & n34227;
  assign n34820 = ~pi644 & ~n34819;
  assign n34821 = pi715 & ~n34820;
  assign n34822 = pi1160 & n34821;
  assign n34823 = ~n34818 & n34822;
  assign n34824 = pi644 & ~n34819;
  assign n34825 = ~pi715 & ~n34824;
  assign n34826 = ~pi644 & n34815;
  assign n34827 = ~pi1160 & ~n34826;
  assign n34828 = n34825 & n34827;
  assign n34829 = ~n34823 & ~n34828;
  assign n34830 = pi790 & n34829;
  assign n34831 = n34817 & ~n34830;
  assign n34832 = ~pi622 & ~n34831;
  assign n34833 = n23049 & n34216;
  assign n34834 = ~pi644 & pi1160;
  assign n34835 = pi644 & ~pi1160;
  assign n34836 = ~n34834 & ~n34835;
  assign n34837 = pi790 & ~n34836;
  assign n34838 = ~po1038 & ~n34837;
  assign n34839 = n34833 & n34838;
  assign n34840 = pi622 & n34839;
  assign n34841 = ~pi639 & ~n34840;
  assign n34842 = pi209 & ~n34841;
  assign n34843 = ~n34832 & n34842;
  assign n34844 = pi647 & n34217;
  assign n34845 = ~pi647 & ~n34376;
  assign n34846 = ~pi1157 & ~n34845;
  assign n34847 = ~n34844 & n34846;
  assign n34848 = pi647 & n34227;
  assign n34849 = pi1157 & ~n34848;
  assign n34850 = ~pi630 & ~n34849;
  assign n34851 = ~n34847 & n34850;
  assign n34852 = ~pi647 & n34217;
  assign n34853 = pi647 & ~n34376;
  assign n34854 = ~n34852 & ~n34853;
  assign n34855 = pi1157 & n34854;
  assign n34856 = ~pi647 & n34227;
  assign n34857 = ~pi1157 & ~n34856;
  assign n34858 = pi630 & ~n34857;
  assign n34859 = ~n34855 & n34858;
  assign n34860 = ~n34851 & ~n34859;
  assign n34861 = pi787 & ~n34860;
  assign n34862 = ~pi787 & ~n34376;
  assign n34863 = ~n34861 & ~n34862;
  assign n34864 = ~pi790 & n34863;
  assign n34865 = ~pi644 & n34863;
  assign n34866 = n34825 & ~n34865;
  assign n34867 = ~pi1160 & ~n34866;
  assign n34868 = ~pi644 & pi715;
  assign n34869 = n34833 & n34868;
  assign n34870 = n34867 & ~n34869;
  assign n34871 = pi644 & n34863;
  assign n34872 = n34821 & ~n34871;
  assign n34873 = pi1160 & ~n34872;
  assign n34874 = pi644 & ~pi715;
  assign n34875 = n34833 & n34874;
  assign n34876 = n34873 & ~n34875;
  assign n34877 = ~n34870 & ~n34876;
  assign n34878 = pi790 & ~n34877;
  assign n34879 = ~po1038 & ~n34878;
  assign n34880 = ~n34864 & n34879;
  assign n34881 = pi622 & ~n34880;
  assign n34882 = pi639 & n34881;
  assign n34883 = n34843 & ~n34882;
  assign po366 = n34811 | n34883;
  assign n34885 = pi210 & ~n16207;
  assign n34886 = ~n32698 & ~n34885;
  assign n34887 = n6215 & n34886;
  assign n34888 = pi947 & ~n34887;
  assign n34889 = pi210 & n16224;
  assign n34890 = pi633 & ~n16224;
  assign n34891 = ~n34889 & ~n34890;
  assign n34892 = ~n6215 & n34891;
  assign n34893 = n34888 & ~n34892;
  assign n34894 = pi634 & n16207;
  assign n34895 = ~n34885 & ~n34894;
  assign n34896 = n6215 & n34895;
  assign n34897 = pi907 & ~n34896;
  assign n34898 = ~n32850 & ~n34889;
  assign n34899 = ~n6215 & n34898;
  assign n34900 = n34897 & ~n34899;
  assign n34901 = n6215 & n16206;
  assign n34902 = n2934 & n34901;
  assign n34903 = n34889 & ~n34902;
  assign n34904 = ~n34900 & ~n34903;
  assign n34905 = ~pi947 & ~n34904;
  assign n34906 = ~n34893 & ~n34905;
  assign n34907 = ~n6236 & n34906;
  assign n34908 = ~n6191 & ~n34895;
  assign n34909 = pi907 & ~n34908;
  assign n34910 = n6191 & ~n34898;
  assign n34911 = n34909 & ~n34910;
  assign n34912 = ~po1101 & n34885;
  assign n34913 = pi210 & po1101;
  assign n34914 = ~n16227 & n34913;
  assign n34915 = ~n34912 & ~n34914;
  assign n34916 = ~pi907 & n34915;
  assign n34917 = ~pi947 & ~n34916;
  assign n34918 = ~n34911 & n34917;
  assign n34919 = ~po1101 & n34886;
  assign n34920 = pi947 & ~n34919;
  assign n34921 = ~n6190 & ~n34891;
  assign n34922 = po1101 & n34886;
  assign n34923 = ~n6191 & ~n34922;
  assign n34924 = ~n34921 & ~n34923;
  assign n34925 = n34920 & ~n34924;
  assign n34926 = n6236 & ~n34925;
  assign n34927 = ~n34918 & n34926;
  assign n34928 = pi223 & ~n34927;
  assign n34929 = ~n34907 & n34928;
  assign n34930 = pi634 & n20323;
  assign n34931 = pi633 & pi947;
  assign n34932 = ~n34930 & ~n34931;
  assign n34933 = n16207 & ~n34932;
  assign n34934 = ~n34885 & ~n34933;
  assign n34935 = n2607 & n34934;
  assign n34936 = pi210 & n16289;
  assign n34937 = pi634 & ~n16289;
  assign n34938 = ~n34936 & ~n34937;
  assign n34939 = n6191 & ~n34938;
  assign n34940 = n34909 & ~n34939;
  assign n34941 = ~n16301 & n34913;
  assign n34942 = ~n34912 & ~n34941;
  assign n34943 = ~pi907 & n34942;
  assign n34944 = ~pi947 & ~n34943;
  assign n34945 = ~n34940 & n34944;
  assign n34946 = pi633 & ~n16289;
  assign n34947 = ~n34936 & ~n34946;
  assign n34948 = ~n6190 & ~n34947;
  assign n34949 = ~n34923 & ~n34948;
  assign n34950 = n34920 & ~n34949;
  assign n34951 = n6236 & ~n34950;
  assign n34952 = ~n34945 & n34951;
  assign n34953 = ~n6215 & n34947;
  assign n34954 = n34888 & ~n34953;
  assign n34955 = ~n6215 & n34938;
  assign n34956 = n34897 & ~n34955;
  assign n34957 = pi210 & ~n16297;
  assign n34958 = ~pi907 & n34957;
  assign n34959 = ~n34956 & ~n34958;
  assign n34960 = ~pi947 & ~n34959;
  assign n34961 = ~n34954 & ~n34960;
  assign n34962 = ~n6236 & n34961;
  assign n34963 = ~n34952 & ~n34962;
  assign n34964 = ~n2607 & ~n34963;
  assign n34965 = ~pi223 & ~n34964;
  assign n34966 = ~n34935 & n34965;
  assign n34967 = ~n34929 & ~n34966;
  assign n34968 = ~pi299 & n34967;
  assign n34969 = n6197 & n34915;
  assign n34970 = ~n6197 & ~n34903;
  assign n34971 = ~pi907 & ~n34970;
  assign n34972 = ~n34969 & n34971;
  assign n34973 = ~n34900 & ~n34972;
  assign n34974 = ~pi947 & ~n34973;
  assign n34975 = ~n34893 & ~n34974;
  assign n34976 = pi215 & ~n34975;
  assign n34977 = n2527 & n34934;
  assign n34978 = ~pi215 & ~n34977;
  assign n34979 = ~n6197 & ~n34957;
  assign n34980 = n6197 & n34942;
  assign n34981 = ~pi907 & ~n34980;
  assign n34982 = ~n34979 & n34981;
  assign n34983 = ~n34956 & ~n34982;
  assign n34984 = ~pi947 & ~n34983;
  assign n34985 = ~n2527 & ~n34954;
  assign n34986 = ~n34984 & n34985;
  assign n34987 = n34978 & ~n34986;
  assign n34988 = pi299 & ~n34987;
  assign n34989 = ~n34976 & n34988;
  assign n34990 = pi39 & ~n34989;
  assign n34991 = ~n34968 & n34990;
  assign n34992 = n16199 & ~n34932;
  assign n34993 = pi210 & ~n16199;
  assign n34994 = ~pi299 & ~n34993;
  assign n34995 = ~n34992 & n34994;
  assign n34996 = ~n16176 & ~n34932;
  assign n34997 = ~n16194 & ~n34996;
  assign n34998 = pi299 & n34997;
  assign n34999 = ~pi39 & ~n34998;
  assign n35000 = ~n34995 & n34999;
  assign n35001 = ~pi38 & ~n35000;
  assign n35002 = ~n34991 & n35001;
  assign n35003 = n16508 & ~n34932;
  assign n35004 = pi210 & ~n16508;
  assign n35005 = pi38 & ~n35004;
  assign n35006 = ~n35003 & n35005;
  assign n35007 = ~n35002 & ~n35006;
  assign n35008 = n10021 & ~n35007;
  assign n35009 = ~pi210 & ~n10021;
  assign po367 = ~n35008 & ~n35009;
  assign n35011 = n10020 & ~n21041;
  assign n35012 = pi606 & n35011;
  assign n35013 = pi643 & ~n35012;
  assign n35014 = n10020 & ~n21037;
  assign n35015 = ~pi606 & n35014;
  assign n35016 = n35013 & ~n35015;
  assign n35017 = n10020 & ~n20505;
  assign n35018 = pi606 & n35017;
  assign n35019 = n16526 & n33690;
  assign n35020 = ~pi643 & ~n35019;
  assign n35021 = ~n35018 & n35020;
  assign n35022 = ~po1038 & ~n35021;
  assign n35023 = ~n35016 & n35022;
  assign n35024 = pi211 & ~n35023;
  assign n35025 = n10020 & n21024;
  assign n35026 = pi606 & ~n35025;
  assign n35027 = n10020 & n21027;
  assign n35028 = ~pi606 & ~n35027;
  assign n35029 = pi643 & ~n35028;
  assign n35030 = ~n35026 & n35029;
  assign n35031 = n10020 & n20526;
  assign n35032 = pi606 & ~pi643;
  assign n35033 = n35031 & n35032;
  assign n35034 = ~n35030 & ~n35033;
  assign n35035 = ~pi211 & ~n35034;
  assign n35036 = ~po1038 & n35035;
  assign po368 = n35024 | n35036;
  assign n35038 = pi607 & n35011;
  assign n35039 = ~pi607 & n35014;
  assign n35040 = pi638 & ~n35039;
  assign n35041 = ~n35038 & n35040;
  assign n35042 = pi607 & n35017;
  assign n35043 = ~pi607 & n16527;
  assign n35044 = ~pi638 & ~n35043;
  assign n35045 = ~n35042 & n35044;
  assign n35046 = ~po1038 & ~n35045;
  assign n35047 = ~n35041 & n35046;
  assign n35048 = ~pi212 & ~n35047;
  assign n35049 = ~pi607 & ~n35027;
  assign n35050 = pi607 & ~n35025;
  assign n35051 = pi638 & ~n35050;
  assign n35052 = ~n35049 & n35051;
  assign n35053 = pi607 & ~pi638;
  assign n35054 = n35031 & n35053;
  assign n35055 = ~n35052 & ~n35054;
  assign n35056 = pi212 & ~n35055;
  assign n35057 = ~po1038 & n35056;
  assign po369 = n35048 | n35057;
  assign n35059 = pi213 & ~po1038;
  assign n35060 = ~pi622 & ~n35027;
  assign n35061 = pi622 & ~n35025;
  assign n35062 = pi639 & ~n35061;
  assign n35063 = ~n35060 & n35062;
  assign n35064 = pi622 & ~pi639;
  assign n35065 = n35031 & n35064;
  assign n35066 = ~n35063 & ~n35065;
  assign n35067 = n35059 & ~n35066;
  assign n35068 = pi639 & n35011;
  assign n35069 = ~pi639 & n35017;
  assign n35070 = pi622 & ~n35069;
  assign n35071 = ~n35068 & n35070;
  assign n35072 = pi639 & n35014;
  assign n35073 = ~pi639 & n16527;
  assign n35074 = ~pi622 & ~n35073;
  assign n35075 = ~n35072 & n35074;
  assign n35076 = ~po1038 & ~n35075;
  assign n35077 = ~n35071 & n35076;
  assign n35078 = ~pi213 & ~n35077;
  assign po370 = n35067 | n35078;
  assign n35080 = pi623 & n35011;
  assign n35081 = ~pi623 & n35014;
  assign n35082 = pi710 & ~n35081;
  assign n35083 = ~n35080 & n35082;
  assign n35084 = pi623 & n35017;
  assign n35085 = ~pi623 & n16527;
  assign n35086 = ~pi710 & ~n35085;
  assign n35087 = ~n35084 & n35086;
  assign n35088 = ~po1038 & ~n35087;
  assign n35089 = ~n35083 & n35088;
  assign n35090 = ~pi214 & ~n35089;
  assign n35091 = ~pi623 & ~n35027;
  assign n35092 = pi623 & ~n35025;
  assign n35093 = pi710 & ~n35092;
  assign n35094 = ~n35091 & n35093;
  assign n35095 = pi623 & ~pi710;
  assign n35096 = n35031 & n35095;
  assign n35097 = ~n35094 & ~n35096;
  assign n35098 = pi214 & ~n35097;
  assign n35099 = ~po1038 & n35098;
  assign po371 = n35090 | n35099;
  assign n35101 = pi215 & ~n10021;
  assign n35102 = ~pi947 & n20720;
  assign n35103 = pi681 & pi907;
  assign n35104 = ~pi947 & n35103;
  assign n35105 = ~n6188 & n16263;
  assign n35106 = n6186 & n16255;
  assign n35107 = ~pi642 & ~n35106;
  assign n35108 = ~n35105 & n35107;
  assign n35109 = pi947 & ~n35108;
  assign n35110 = ~n35104 & ~n35109;
  assign n35111 = ~n35102 & n35110;
  assign n35112 = pi299 & ~n35111;
  assign n35113 = pi642 & pi947;
  assign n35114 = ~n35104 & ~n35113;
  assign n35115 = n16271 & ~n35114;
  assign n35116 = ~pi642 & n16297;
  assign n35117 = ~n6236 & ~n35116;
  assign n35118 = pi947 & ~n35117;
  assign n35119 = ~pi642 & n16301;
  assign n35120 = n6188 & n35119;
  assign n35121 = ~n6184 & n16207;
  assign n35122 = ~pi642 & n35121;
  assign n35123 = ~n16957 & ~n35122;
  assign n35124 = ~n6188 & ~n35123;
  assign n35125 = ~n35120 & ~n35124;
  assign n35126 = n6236 & n35125;
  assign n35127 = n35118 & ~n35126;
  assign n35128 = n20809 & ~n35103;
  assign n35129 = ~n2607 & ~n35128;
  assign n35130 = ~n35127 & n35129;
  assign n35131 = n16921 & ~n35130;
  assign n35132 = ~n35115 & n35131;
  assign n35133 = ~n6236 & ~n35108;
  assign n35134 = ~pi642 & ~n16246;
  assign n35135 = ~n16245 & n35134;
  assign n35136 = n6236 & ~n35135;
  assign n35137 = ~n35133 & ~n35136;
  assign n35138 = pi947 & n35137;
  assign n35139 = n20797 & ~n35104;
  assign n35140 = ~n35138 & ~n35139;
  assign n35141 = pi223 & ~n35140;
  assign n35142 = ~pi299 & ~n35141;
  assign n35143 = ~n35132 & n35142;
  assign n35144 = ~n35112 & ~n35143;
  assign n35145 = pi215 & ~n35144;
  assign n35146 = n6236 & ~n16234;
  assign n35147 = n35103 & ~n35146;
  assign n35148 = ~pi947 & ~n35147;
  assign n35149 = pi947 & ~n16261;
  assign n35150 = n16263 & ~n35149;
  assign n35151 = ~n6236 & n35150;
  assign n35152 = pi642 & ~n6187;
  assign n35153 = n16207 & n35152;
  assign n35154 = pi642 & n6187;
  assign n35155 = ~n16237 & n35154;
  assign n35156 = ~n16236 & n35155;
  assign n35157 = ~n35153 & ~n35156;
  assign n35158 = pi947 & n35157;
  assign n35159 = ~n35151 & ~n35158;
  assign n35160 = ~n35148 & n35159;
  assign n35161 = pi223 & ~n35160;
  assign n35162 = ~n16294 & n35103;
  assign n35163 = ~pi947 & ~n35162;
  assign n35164 = ~n6188 & n16292;
  assign n35165 = ~n16296 & ~n35164;
  assign n35166 = n35154 & n35165;
  assign n35167 = ~n16292 & n35152;
  assign n35168 = ~n35166 & ~n35167;
  assign n35169 = pi947 & n35168;
  assign n35170 = ~n35163 & ~n35169;
  assign n35171 = ~n6236 & ~n35170;
  assign n35172 = ~n16313 & n35155;
  assign n35173 = ~n35153 & ~n35172;
  assign n35174 = pi947 & ~n35173;
  assign n35175 = n16309 & n35104;
  assign n35176 = ~n35174 & ~n35175;
  assign n35177 = n6236 & n35176;
  assign n35178 = ~n2607 & ~n35177;
  assign n35179 = ~n35171 & n35178;
  assign n35180 = ~pi223 & ~n35179;
  assign n35181 = ~n35115 & n35180;
  assign n35182 = ~n35161 & ~n35181;
  assign n35183 = ~pi299 & ~n35182;
  assign n35184 = n16342 & ~n35114;
  assign n35185 = ~n2527 & n35170;
  assign n35186 = pi299 & ~n35185;
  assign n35187 = ~n35184 & n35186;
  assign n35188 = ~pi215 & ~n35187;
  assign n35189 = ~n35183 & n35188;
  assign n35190 = ~n35145 & ~n35189;
  assign n35191 = pi39 & ~n35190;
  assign n35192 = n16195 & ~n35114;
  assign n35193 = pi215 & ~n16195;
  assign n35194 = ~n35192 & ~n35193;
  assign n35195 = pi299 & n35194;
  assign n35196 = pi215 & ~n16199;
  assign n35197 = n16199 & ~n35114;
  assign n35198 = ~pi299 & ~n35197;
  assign n35199 = ~n35196 & n35198;
  assign n35200 = ~pi39 & ~n35199;
  assign n35201 = ~n35195 & n35200;
  assign n35202 = ~pi38 & ~n35201;
  assign n35203 = ~n35191 & n35202;
  assign n35204 = n16508 & ~n35114;
  assign n35205 = pi215 & ~n16508;
  assign n35206 = pi38 & ~n35205;
  assign n35207 = ~n35204 & n35206;
  assign n35208 = ~n35203 & ~n35207;
  assign n35209 = n10021 & n35208;
  assign po372 = n35101 | n35209;
  assign n35211 = pi614 & pi947;
  assign n35212 = n35165 & n35211;
  assign n35213 = pi662 & pi907;
  assign n35214 = ~pi947 & n35213;
  assign n35215 = ~n16294 & n35214;
  assign n35216 = ~n35212 & ~n35215;
  assign n35217 = n5742 & ~n35216;
  assign n35218 = ~n35211 & ~n35214;
  assign n35219 = n16342 & ~n35218;
  assign n35220 = ~pi947 & n20492;
  assign n35221 = pi947 & ~n16297;
  assign n35222 = ~n35220 & ~n35221;
  assign n35223 = n35218 & n35222;
  assign n35224 = pi216 & ~n35223;
  assign n35225 = ~n35219 & ~n35224;
  assign n35226 = ~n35217 & n35225;
  assign n35227 = ~pi215 & ~n35226;
  assign n35228 = ~pi614 & ~n16224;
  assign n35229 = n16262 & n16318;
  assign n35230 = ~n35228 & ~n35229;
  assign n35231 = pi947 & n35230;
  assign n35232 = pi216 & ~n35231;
  assign n35233 = ~n35102 & n35232;
  assign n35234 = ~n35214 & n35233;
  assign n35235 = ~n16236 & n16315;
  assign n35236 = pi947 & ~n16312;
  assign n35237 = ~n35235 & n35236;
  assign n35238 = ~n16263 & n35214;
  assign n35239 = ~n35149 & ~n35238;
  assign n35240 = ~n35237 & ~n35239;
  assign n35241 = ~pi216 & ~n35240;
  assign n35242 = pi215 & ~n35241;
  assign n35243 = ~n35234 & n35242;
  assign n35244 = ~n35227 & ~n35243;
  assign n35245 = pi299 & n35244;
  assign n35246 = n16271 & ~n35218;
  assign n35247 = n16298 & n35218;
  assign n35248 = pi947 & ~n16323;
  assign n35249 = ~pi947 & n16327;
  assign n35250 = ~n35213 & n35249;
  assign n35251 = ~n35248 & ~n35250;
  assign n35252 = n6236 & ~n35251;
  assign n35253 = ~n2607 & ~n35252;
  assign n35254 = ~n35247 & n35253;
  assign n35255 = n16921 & ~n35254;
  assign n35256 = ~n35246 & n35255;
  assign n35257 = ~n6236 & n35230;
  assign n35258 = ~pi614 & ~n16246;
  assign n35259 = ~n16245 & n35258;
  assign n35260 = n6236 & ~n35259;
  assign n35261 = ~n35257 & ~n35260;
  assign n35262 = pi947 & n35261;
  assign n35263 = n20797 & ~n35214;
  assign n35264 = ~n35262 & ~n35263;
  assign n35265 = pi223 & ~n35264;
  assign n35266 = pi216 & ~n35265;
  assign n35267 = ~n35256 & n35266;
  assign n35268 = ~n35146 & n35213;
  assign n35269 = ~pi947 & ~n35268;
  assign n35270 = ~n35151 & ~n35237;
  assign n35271 = ~n35269 & n35270;
  assign n35272 = pi223 & ~n35271;
  assign n35273 = ~pi216 & ~n35272;
  assign n35274 = ~n6236 & n35216;
  assign n35275 = ~n16312 & ~n16316;
  assign n35276 = pi947 & ~n35275;
  assign n35277 = n16309 & n35214;
  assign n35278 = ~n35276 & ~n35277;
  assign n35279 = n6236 & n35278;
  assign n35280 = ~n2607 & ~n35279;
  assign n35281 = ~n35274 & n35280;
  assign n35282 = ~pi223 & ~n35281;
  assign n35283 = ~n35246 & n35282;
  assign n35284 = n35273 & ~n35283;
  assign n35285 = ~n35267 & ~n35284;
  assign n35286 = ~pi299 & n35285;
  assign n35287 = pi39 & ~n35286;
  assign n35288 = ~n35245 & n35287;
  assign n35289 = pi216 & ~n16199;
  assign n35290 = n16199 & ~n35218;
  assign n35291 = ~pi299 & ~n35290;
  assign n35292 = ~n35289 & n35291;
  assign n35293 = n16195 & ~n35218;
  assign n35294 = pi216 & ~n16195;
  assign n35295 = ~n35293 & ~n35294;
  assign n35296 = pi299 & n35295;
  assign n35297 = ~pi39 & ~n35296;
  assign n35298 = ~n35292 & n35297;
  assign n35299 = ~pi38 & ~n35298;
  assign n35300 = ~n35288 & n35299;
  assign n35301 = pi216 & ~n16508;
  assign n35302 = n16508 & ~n35218;
  assign n35303 = pi38 & ~n35302;
  assign n35304 = ~n35301 & n35303;
  assign n35305 = ~n35300 & ~n35304;
  assign n35306 = n10021 & ~n35305;
  assign n35307 = ~pi216 & ~n10021;
  assign po373 = ~n35306 & ~n35307;
  assign n35309 = ~pi695 & n34880;
  assign n35310 = pi217 & ~n35309;
  assign n35311 = pi695 & n34839;
  assign n35312 = n35310 & ~n35311;
  assign n35313 = pi695 & ~n34806;
  assign n35314 = ~pi695 & ~n34798;
  assign n35315 = ~pi217 & ~n35314;
  assign n35316 = ~n35313 & n35315;
  assign n35317 = pi612 & ~n35316;
  assign n35318 = ~n35312 & n35317;
  assign n35319 = pi695 & ~n34765;
  assign n35320 = ~pi695 & ~n34762;
  assign n35321 = ~pi217 & ~n35320;
  assign n35322 = ~n35319 & n35321;
  assign n35323 = ~pi695 & n34831;
  assign n35324 = pi217 & ~n35323;
  assign n35325 = ~pi612 & ~n35324;
  assign n35326 = ~n35322 & n35325;
  assign po374 = n35318 | n35326;
  assign n35328 = n34033 & ~n34108;
  assign n35329 = ~n34033 & ~n34138;
  assign n35330 = ~n35328 & ~n35329;
  assign n35331 = ~pi218 & ~n35330;
  assign n35332 = n34033 & n34145;
  assign n35333 = pi218 & ~n35332;
  assign po375 = ~n35331 & ~n35333;
  assign n35335 = ~pi219 & ~po1038;
  assign n35336 = ~pi617 & ~n35027;
  assign n35337 = pi617 & ~n35025;
  assign n35338 = pi637 & ~n35337;
  assign n35339 = ~n35336 & n35338;
  assign n35340 = pi617 & ~pi637;
  assign n35341 = n35031 & n35340;
  assign n35342 = ~n35339 & ~n35341;
  assign n35343 = n35335 & ~n35342;
  assign n35344 = pi617 & n35011;
  assign n35345 = ~pi617 & n35014;
  assign n35346 = pi637 & ~n35345;
  assign n35347 = ~n35344 & n35346;
  assign n35348 = pi617 & n35017;
  assign n35349 = ~pi617 & n16527;
  assign n35350 = ~pi637 & ~n35349;
  assign n35351 = ~n35348 & n35350;
  assign n35352 = ~po1038 & ~n35351;
  assign n35353 = ~n35347 & n35352;
  assign n35354 = pi219 & ~n35353;
  assign po376 = n35343 | n35354;
  assign n35356 = ~n33974 & n34156;
  assign n35357 = ~n34011 & ~n34156;
  assign n35358 = ~n35356 & ~n35357;
  assign n35359 = ~pi220 & ~n35358;
  assign n35360 = n34021 & n34156;
  assign n35361 = pi220 & ~n35360;
  assign po377 = ~n35359 & ~n35361;
  assign n35363 = pi661 & n20323;
  assign n35364 = pi221 & ~n35363;
  assign n35365 = ~pi616 & ~n35106;
  assign n35366 = ~n35105 & n35365;
  assign n35367 = pi947 & ~n35366;
  assign n35368 = ~n35102 & ~n35367;
  assign n35369 = n35364 & n35368;
  assign n35370 = pi947 & ~n16243;
  assign n35371 = ~n35363 & ~n35370;
  assign n35372 = ~n35150 & ~n35371;
  assign n35373 = ~pi221 & ~n35372;
  assign n35374 = pi215 & ~n35373;
  assign n35375 = ~n35369 & n35374;
  assign n35376 = pi616 & pi947;
  assign n35377 = n35165 & n35376;
  assign n35378 = ~n16294 & n35363;
  assign n35379 = ~n35377 & ~n35378;
  assign n35380 = pi216 & ~n35379;
  assign n35381 = ~n35363 & ~n35376;
  assign n35382 = n16342 & ~n35381;
  assign n35383 = ~pi221 & ~n35382;
  assign n35384 = ~n35380 & n35383;
  assign n35385 = ~pi616 & ~n6187;
  assign n35386 = ~n6190 & n16307;
  assign n35387 = ~n16291 & ~n35386;
  assign n35388 = n35385 & ~n35387;
  assign n35389 = ~pi616 & n6187;
  assign n35390 = ~n35116 & ~n35166;
  assign n35391 = n35389 & ~n35390;
  assign n35392 = pi947 & ~n35391;
  assign n35393 = ~n35388 & n35392;
  assign n35394 = ~n35220 & ~n35393;
  assign n35395 = n35364 & n35394;
  assign n35396 = ~pi215 & ~n35395;
  assign n35397 = ~n35384 & n35396;
  assign n35398 = ~n35375 & ~n35397;
  assign n35399 = pi299 & n35398;
  assign n35400 = n16271 & ~n35381;
  assign n35401 = ~pi223 & ~n35400;
  assign n35402 = ~pi947 & ~n16297;
  assign n35403 = ~n35393 & ~n35402;
  assign n35404 = ~n6236 & ~n35403;
  assign n35405 = n16307 & n35385;
  assign n35406 = ~n16324 & n35389;
  assign n35407 = ~n35405 & ~n35406;
  assign n35408 = pi947 & ~n35407;
  assign n35409 = ~n35249 & ~n35408;
  assign n35410 = n6236 & n35409;
  assign n35411 = ~n35363 & ~n35410;
  assign n35412 = ~n35404 & n35411;
  assign n35413 = ~n2607 & ~n35412;
  assign n35414 = ~n16920 & ~n35413;
  assign n35415 = n35401 & n35414;
  assign n35416 = pi947 & n16248;
  assign n35417 = ~pi947 & n16250;
  assign n35418 = ~n35416 & ~n35417;
  assign n35419 = n6236 & n35418;
  assign n35420 = pi223 & ~n35419;
  assign n35421 = ~pi947 & ~n16267;
  assign n35422 = ~n35367 & ~n35421;
  assign n35423 = ~n6236 & ~n35422;
  assign n35424 = ~n35363 & ~n35423;
  assign n35425 = n35420 & n35424;
  assign n35426 = pi221 & ~n35425;
  assign n35427 = ~n35415 & n35426;
  assign n35428 = ~n35146 & n35363;
  assign n35429 = ~n35370 & ~n35428;
  assign n35430 = ~n35151 & ~n35429;
  assign n35431 = pi223 & ~n35430;
  assign n35432 = n16309 & n35363;
  assign n35433 = n16239 & ~n16313;
  assign n35434 = ~n16242 & ~n35433;
  assign n35435 = pi947 & ~n35434;
  assign n35436 = n6236 & ~n35435;
  assign n35437 = ~n35432 & n35436;
  assign n35438 = ~n6236 & n35379;
  assign n35439 = ~n2607 & ~n35438;
  assign n35440 = ~n35437 & n35439;
  assign n35441 = n35401 & ~n35440;
  assign n35442 = ~pi221 & ~n35441;
  assign n35443 = ~n35431 & n35442;
  assign n35444 = ~n35427 & ~n35443;
  assign n35445 = ~pi299 & n35444;
  assign n35446 = pi39 & ~n35445;
  assign n35447 = ~n35399 & n35446;
  assign n35448 = pi221 & ~n16199;
  assign n35449 = n16199 & ~n35381;
  assign n35450 = ~pi299 & ~n35449;
  assign n35451 = ~n35448 & n35450;
  assign n35452 = n16195 & ~n35381;
  assign n35453 = pi221 & ~n16195;
  assign n35454 = ~n35452 & ~n35453;
  assign n35455 = pi299 & n35454;
  assign n35456 = ~pi39 & ~n35455;
  assign n35457 = ~n35451 & n35456;
  assign n35458 = ~pi38 & ~n35457;
  assign n35459 = ~n35447 & n35458;
  assign n35460 = pi221 & ~n16508;
  assign n35461 = n16508 & ~n35381;
  assign n35462 = pi38 & ~n35461;
  assign n35463 = ~n35460 & n35462;
  assign n35464 = ~n35459 & ~n35463;
  assign n35465 = n10021 & ~n35464;
  assign n35466 = ~pi221 & ~n10021;
  assign po378 = ~n35465 & ~n35466;
  assign n35468 = ~n16270 & ~n16330;
  assign n35469 = ~pi299 & ~n35468;
  assign n35470 = ~n16354 & ~n35469;
  assign n35471 = pi39 & n35470;
  assign n35472 = ~pi38 & ~n35471;
  assign n35473 = ~n17520 & n35472;
  assign n35474 = n18119 & ~n35473;
  assign n35475 = pi222 & ~n35474;
  assign n35476 = n17355 & ~n35475;
  assign n35477 = pi222 & ~n10020;
  assign n35478 = ~pi222 & ~n16460;
  assign n35479 = ~pi616 & n16460;
  assign n35480 = pi222 & n16380;
  assign n35481 = ~pi39 & ~n35480;
  assign n35482 = ~n35479 & n35481;
  assign n35483 = ~n35478 & n35482;
  assign n35484 = ~pi38 & ~n35483;
  assign n35485 = pi616 & n16393;
  assign n35486 = ~n32728 & ~n35485;
  assign n35487 = ~n16294 & n35486;
  assign n35488 = ~n6186 & ~n35487;
  assign n35489 = ~n16253 & n35487;
  assign n35490 = ~n16289 & ~n35485;
  assign n35491 = ~n16385 & ~n35490;
  assign n35492 = n16253 & ~n35491;
  assign n35493 = n6186 & ~n35492;
  assign n35494 = ~n35489 & n35493;
  assign n35495 = ~n35488 & ~n35494;
  assign n35496 = ~n6236 & n35495;
  assign n35497 = pi616 & ~n16394;
  assign n35498 = ~n16308 & ~n35497;
  assign n35499 = ~n6186 & ~n35498;
  assign n35500 = ~n16253 & n35498;
  assign n35501 = n16253 & ~n35485;
  assign n35502 = n16301 & n35501;
  assign n35503 = n6186 & ~n35502;
  assign n35504 = ~n35500 & n35503;
  assign n35505 = ~n35499 & ~n35504;
  assign n35506 = n6236 & n35505;
  assign n35507 = pi222 & ~n35506;
  assign n35508 = ~n35496 & n35507;
  assign n35509 = ~n16292 & n35485;
  assign n35510 = ~n6186 & ~n35509;
  assign n35511 = ~n16253 & n35509;
  assign n35512 = pi616 & n16253;
  assign n35513 = n16809 & n35512;
  assign n35514 = n6186 & ~n35513;
  assign n35515 = ~n35511 & n35514;
  assign n35516 = ~n35510 & ~n35515;
  assign n35517 = ~n6236 & n35516;
  assign n35518 = ~n6188 & n16465;
  assign n35519 = ~n16464 & ~n35518;
  assign n35520 = pi616 & ~n35519;
  assign n35521 = n6236 & n35520;
  assign n35522 = pi224 & ~n35521;
  assign n35523 = ~n35517 & n35522;
  assign n35524 = pi616 & n16465;
  assign n35525 = ~pi224 & ~n35524;
  assign n35526 = ~pi222 & ~n35525;
  assign n35527 = ~n35523 & n35526;
  assign n35528 = ~pi223 & ~n35527;
  assign n35529 = ~n35508 & n35528;
  assign n35530 = pi616 & ~n16420;
  assign n35531 = ~n16263 & ~n35530;
  assign n35532 = ~n16255 & ~n35530;
  assign n35533 = ~n16263 & n35532;
  assign n35534 = n6186 & ~n35533;
  assign n35535 = n35531 & ~n35534;
  assign n35536 = ~n6236 & n35535;
  assign n35537 = ~n16233 & ~n35497;
  assign n35538 = ~n6186 & ~n35537;
  assign n35539 = ~n16253 & n35537;
  assign n35540 = n16227 & n35501;
  assign n35541 = n6186 & ~n35540;
  assign n35542 = ~n35539 & n35541;
  assign n35543 = ~n35538 & ~n35542;
  assign n35544 = n6236 & n35543;
  assign n35545 = ~n35536 & ~n35544;
  assign n35546 = pi222 & n35545;
  assign n35547 = ~n16479 & ~n35518;
  assign n35548 = pi616 & ~n35547;
  assign n35549 = ~pi222 & n35548;
  assign n35550 = ~n16489 & n35549;
  assign n35551 = pi223 & ~n35550;
  assign n35552 = ~n35546 & n35551;
  assign n35553 = ~n35529 & ~n35552;
  assign n35554 = ~pi299 & ~n35553;
  assign n35555 = ~n16478 & n35549;
  assign n35556 = n6198 & n35543;
  assign n35557 = ~n6198 & n35535;
  assign n35558 = pi222 & ~n35557;
  assign n35559 = ~n35556 & n35558;
  assign n35560 = ~n35555 & ~n35559;
  assign n35561 = pi215 & ~n35560;
  assign n35562 = ~n6198 & n35495;
  assign n35563 = n6198 & n35505;
  assign n35564 = pi222 & ~n35563;
  assign n35565 = ~n35562 & n35564;
  assign n35566 = n6198 & ~n35520;
  assign n35567 = ~n6198 & ~n35516;
  assign n35568 = ~pi222 & ~n35567;
  assign n35569 = ~n35566 & n35568;
  assign n35570 = ~n2527 & ~n35569;
  assign n35571 = ~n35565 & n35570;
  assign n35572 = pi222 & ~n16207;
  assign n35573 = n2527 & ~n35572;
  assign n35574 = ~n35524 & n35573;
  assign n35575 = ~pi215 & ~n35574;
  assign n35576 = ~n35571 & n35575;
  assign n35577 = pi299 & ~n35576;
  assign n35578 = ~n35561 & n35577;
  assign n35579 = pi39 & ~n35578;
  assign n35580 = ~n35554 & n35579;
  assign n35581 = n35484 & ~n35580;
  assign n35582 = pi222 & ~n16508;
  assign n35583 = pi38 & ~n35582;
  assign n35584 = n16508 & n35485;
  assign n35585 = n35583 & ~n35584;
  assign n35586 = ~n35581 & ~n35585;
  assign n35587 = n10020 & n35586;
  assign n35588 = ~n35477 & ~n35587;
  assign n35589 = ~n16521 & ~n35588;
  assign n35590 = n16521 & n35475;
  assign n35591 = ~n35589 & ~n35590;
  assign n35592 = ~pi785 & ~n35591;
  assign n35593 = pi609 & n35591;
  assign n35594 = ~pi609 & ~n35475;
  assign n35595 = pi1155 & ~n35594;
  assign n35596 = ~n35593 & n35595;
  assign n35597 = ~pi609 & n35591;
  assign n35598 = pi609 & ~n35475;
  assign n35599 = ~pi1155 & ~n35598;
  assign n35600 = ~n35597 & n35599;
  assign n35601 = ~n35596 & ~n35600;
  assign n35602 = pi785 & ~n35601;
  assign n35603 = ~n35592 & ~n35602;
  assign n35604 = ~pi781 & ~n35603;
  assign n35605 = pi618 & n35603;
  assign n35606 = ~pi618 & ~n35475;
  assign n35607 = pi1154 & ~n35606;
  assign n35608 = ~n35605 & n35607;
  assign n35609 = ~pi618 & n35603;
  assign n35610 = pi618 & ~n35475;
  assign n35611 = ~pi1154 & ~n35610;
  assign n35612 = ~n35609 & n35611;
  assign n35613 = ~n35608 & ~n35612;
  assign n35614 = pi781 & ~n35613;
  assign n35615 = ~n35604 & ~n35614;
  assign n35616 = ~pi789 & ~n35615;
  assign n35617 = pi619 & n35615;
  assign n35618 = ~pi619 & ~n35475;
  assign n35619 = pi1159 & ~n35618;
  assign n35620 = ~n35617 & n35619;
  assign n35621 = ~pi619 & n35615;
  assign n35622 = pi619 & ~n35475;
  assign n35623 = ~pi1159 & ~n35622;
  assign n35624 = ~n35621 & n35623;
  assign n35625 = ~n35620 & ~n35624;
  assign n35626 = pi789 & ~n35625;
  assign n35627 = ~n35616 & ~n35626;
  assign n35628 = ~n17355 & n35627;
  assign n35629 = ~n35476 & ~n35628;
  assign n35630 = ~n19999 & n35629;
  assign n35631 = ~n32843 & ~n35475;
  assign n35632 = pi661 & pi680;
  assign n35633 = n16728 & ~n35632;
  assign n35634 = pi222 & n16710;
  assign n35635 = ~pi222 & ~n16728;
  assign n35636 = ~pi299 & ~n35635;
  assign n35637 = ~n35634 & n35636;
  assign n35638 = ~n35633 & n35637;
  assign n35639 = ~pi39 & ~n35638;
  assign n35640 = n16733 & ~n35632;
  assign n35641 = pi222 & n16716;
  assign n35642 = ~pi222 & ~n16733;
  assign n35643 = pi299 & ~n35642;
  assign n35644 = ~n35641 & n35643;
  assign n35645 = ~n35640 & n35644;
  assign n35646 = n35639 & ~n35645;
  assign n35647 = pi661 & ~n16657;
  assign n35648 = n6186 & ~n16312;
  assign n35649 = n16324 & n35648;
  assign n35650 = ~n35647 & ~n35649;
  assign n35651 = ~pi661 & n16310;
  assign n35652 = n35650 & ~n35651;
  assign n35653 = n6236 & n35652;
  assign n35654 = ~pi661 & ~n16297;
  assign n35655 = ~n16294 & ~n16596;
  assign n35656 = pi661 & ~n35655;
  assign n35657 = ~n35654 & ~n35656;
  assign n35658 = ~n6236 & n35657;
  assign n35659 = pi222 & ~n35658;
  assign n35660 = ~n35653 & n35659;
  assign n35661 = ~n16294 & n16596;
  assign n35662 = pi661 & n35661;
  assign n35663 = ~n6236 & n35662;
  assign n35664 = ~n16607 & n35632;
  assign n35665 = n6236 & n35664;
  assign n35666 = pi224 & ~n35665;
  assign n35667 = ~n35663 & n35666;
  assign n35668 = pi661 & n16630;
  assign n35669 = ~pi224 & ~n35668;
  assign n35670 = ~pi222 & ~n35669;
  assign n35671 = ~n35667 & n35670;
  assign n35672 = ~pi223 & ~n35671;
  assign n35673 = ~n35660 & n35672;
  assign n35674 = ~pi661 & pi681;
  assign n35675 = n16263 & n35674;
  assign n35676 = pi661 & n16679;
  assign n35677 = ~n16259 & ~n35676;
  assign n35678 = ~n35674 & n35677;
  assign n35679 = ~n35675 & ~n35678;
  assign n35680 = ~n6236 & n35679;
  assign n35681 = ~pi661 & ~n16250;
  assign n35682 = ~n16676 & ~n16682;
  assign n35683 = pi661 & ~n35682;
  assign n35684 = ~n35681 & ~n35683;
  assign n35685 = n6236 & n35684;
  assign n35686 = ~n35680 & ~n35685;
  assign n35687 = pi222 & n35686;
  assign n35688 = ~pi222 & pi661;
  assign n35689 = n16620 & n35688;
  assign n35690 = pi223 & ~n35689;
  assign n35691 = ~n35687 & n35690;
  assign n35692 = ~n35673 & ~n35691;
  assign n35693 = ~pi299 & ~n35692;
  assign n35694 = n35573 & ~n35668;
  assign n35695 = n6198 & n35652;
  assign n35696 = ~n6198 & n35657;
  assign n35697 = pi222 & ~n35696;
  assign n35698 = ~n35695 & n35697;
  assign n35699 = ~n6198 & ~n35662;
  assign n35700 = n6198 & ~n35664;
  assign n35701 = ~pi222 & ~n35700;
  assign n35702 = ~n35699 & n35701;
  assign n35703 = ~n2527 & ~n35702;
  assign n35704 = ~n35698 & n35703;
  assign n35705 = ~pi215 & ~n35704;
  assign n35706 = ~n35694 & n35705;
  assign n35707 = n16634 & n35688;
  assign n35708 = n6198 & n35684;
  assign n35709 = ~n6198 & n35679;
  assign n35710 = pi222 & ~n35709;
  assign n35711 = ~n35708 & n35710;
  assign n35712 = ~n35707 & ~n35711;
  assign n35713 = pi215 & ~n35712;
  assign n35714 = pi299 & ~n35713;
  assign n35715 = ~n35706 & n35714;
  assign n35716 = ~n35693 & ~n35715;
  assign n35717 = pi39 & ~n35716;
  assign n35718 = ~n35646 & ~n35717;
  assign n35719 = ~pi38 & ~n35718;
  assign n35720 = pi661 & n16743;
  assign n35721 = n35583 & ~n35720;
  assign n35722 = ~n35719 & ~n35721;
  assign n35723 = n10020 & n35722;
  assign n35724 = ~n35477 & ~n35723;
  assign n35725 = ~pi778 & ~n35724;
  assign n35726 = pi625 & n35724;
  assign n35727 = ~pi625 & ~n35475;
  assign n35728 = pi1153 & ~n35727;
  assign n35729 = ~n35726 & n35728;
  assign n35730 = ~pi625 & n35724;
  assign n35731 = pi625 & ~n35475;
  assign n35732 = ~pi1153 & ~n35731;
  assign n35733 = ~n35730 & n35732;
  assign n35734 = ~n35729 & ~n35733;
  assign n35735 = pi778 & ~n35734;
  assign n35736 = ~n35725 & ~n35735;
  assign n35737 = ~n16593 & ~n35736;
  assign n35738 = n16593 & n35475;
  assign n35739 = ~n35737 & ~n35738;
  assign n35740 = ~n16589 & ~n35739;
  assign n35741 = n16589 & n35475;
  assign n35742 = ~n35740 & ~n35741;
  assign n35743 = ~n17159 & n35742;
  assign n35744 = ~n17183 & n35743;
  assign n35745 = ~n35631 & ~n35744;
  assign n35746 = pi628 & ~n35745;
  assign n35747 = ~pi628 & ~n35475;
  assign n35748 = n16121 & ~n35747;
  assign n35749 = ~n35746 & n35748;
  assign n35750 = ~pi628 & ~n35745;
  assign n35751 = pi628 & ~n35475;
  assign n35752 = n16122 & ~n35751;
  assign n35753 = ~n35750 & n35752;
  assign n35754 = ~n35749 & ~n35753;
  assign n35755 = ~n35630 & n35754;
  assign n35756 = pi792 & ~n35755;
  assign n35757 = pi626 & n35627;
  assign n35758 = ~pi626 & ~n35475;
  assign n35759 = n17180 & ~n35758;
  assign n35760 = ~n35757 & n35759;
  assign n35761 = ~pi626 & n35627;
  assign n35762 = pi626 & ~n35475;
  assign n35763 = n17181 & ~n35762;
  assign n35764 = ~n35761 & n35763;
  assign n35765 = n17159 & ~n35475;
  assign n35766 = ~n35743 & ~n35765;
  assign n35767 = n17350 & n35766;
  assign n35768 = ~n35764 & ~n35767;
  assign n35769 = ~n35760 & n35768;
  assign n35770 = ~n17356 & n35769;
  assign n35771 = pi788 & ~n35769;
  assign n35772 = pi618 & n35739;
  assign n35773 = pi609 & n35736;
  assign n35774 = pi625 & n35588;
  assign n35775 = ~n35485 & ~n35632;
  assign n35776 = pi616 & ~n16953;
  assign n35777 = ~pi616 & ~n16877;
  assign n35778 = ~n35776 & ~n35777;
  assign n35779 = ~n35775 & n35778;
  assign n35780 = n35573 & ~n35779;
  assign n35781 = ~pi680 & n35487;
  assign n35782 = pi614 & n16393;
  assign n35783 = ~n16292 & n35782;
  assign n35784 = n6190 & n16644;
  assign n35785 = ~n16646 & ~n35784;
  assign n35786 = n16952 & ~n35785;
  assign n35787 = pi614 & ~n35786;
  assign n35788 = ~n16942 & n35785;
  assign n35789 = pi642 & ~n35788;
  assign n35790 = ~pi603 & n35785;
  assign n35791 = pi603 & n16289;
  assign n35792 = pi603 & n16775;
  assign n35793 = ~n35791 & ~n35792;
  assign n35794 = ~n35790 & n35793;
  assign n35795 = ~pi642 & n35794;
  assign n35796 = n6184 & ~n35795;
  assign n35797 = ~n35789 & n35796;
  assign n35798 = ~pi614 & pi616;
  assign n35799 = n35788 & n35798;
  assign n35800 = ~n35797 & ~n35799;
  assign n35801 = ~n35787 & n35800;
  assign n35802 = ~n35783 & ~n35801;
  assign n35803 = ~n35485 & ~n35802;
  assign n35804 = pi680 & n35803;
  assign n35805 = ~n35781 & ~n35804;
  assign n35806 = pi661 & n35805;
  assign n35807 = ~n35487 & n35674;
  assign n35808 = ~n35494 & ~n35807;
  assign n35809 = ~n35806 & n35808;
  assign n35810 = ~n6198 & ~n35809;
  assign n35811 = ~pi680 & n35498;
  assign n35812 = pi616 & ~n17022;
  assign n35813 = pi680 & ~n35812;
  assign n35814 = ~n16824 & n35813;
  assign n35815 = ~n35811 & ~n35814;
  assign n35816 = pi661 & n35815;
  assign n35817 = ~n35498 & n35674;
  assign n35818 = ~n35504 & ~n35817;
  assign n35819 = ~n35816 & n35818;
  assign n35820 = n6198 & ~n35819;
  assign n35821 = pi222 & ~n35820;
  assign n35822 = ~n35810 & n35821;
  assign n35823 = pi680 & n16872;
  assign n35824 = ~n35509 & ~n35823;
  assign n35825 = pi661 & n35824;
  assign n35826 = ~n35509 & n35674;
  assign n35827 = ~n35515 & ~n35826;
  assign n35828 = ~n35825 & n35827;
  assign n35829 = ~n6198 & n35828;
  assign n35830 = n16463 & n35512;
  assign n35831 = ~pi681 & n35830;
  assign n35832 = ~pi661 & ~n35831;
  assign n35833 = ~n35524 & n35832;
  assign n35834 = n6188 & ~n35830;
  assign n35835 = pi680 & ~n16887;
  assign n35836 = ~n35776 & n35835;
  assign n35837 = ~pi680 & n35524;
  assign n35838 = pi661 & ~n35837;
  assign n35839 = ~n35836 & n35838;
  assign n35840 = ~n35834 & ~n35839;
  assign n35841 = ~n35833 & n35840;
  assign n35842 = n6198 & n35841;
  assign n35843 = ~pi222 & ~n35842;
  assign n35844 = ~n35829 & n35843;
  assign n35845 = ~n35822 & ~n35844;
  assign n35846 = ~n2527 & ~n35845;
  assign n35847 = ~pi215 & ~n35846;
  assign n35848 = ~n35780 & n35847;
  assign n35849 = ~pi680 & n35531;
  assign n35850 = ~n16798 & n16952;
  assign n35851 = pi616 & ~n35850;
  assign n35852 = pi680 & ~n35851;
  assign n35853 = n16801 & n35852;
  assign n35854 = ~n35849 & ~n35853;
  assign n35855 = pi661 & n35854;
  assign n35856 = ~n35531 & n35674;
  assign n35857 = ~n35534 & ~n35856;
  assign n35858 = ~n35855 & n35857;
  assign n35859 = ~n6198 & ~n35858;
  assign n35860 = ~pi680 & n35537;
  assign n35861 = ~n16790 & n35813;
  assign n35862 = ~n35860 & ~n35861;
  assign n35863 = pi661 & n35862;
  assign n35864 = ~n35537 & n35674;
  assign n35865 = ~n35542 & ~n35864;
  assign n35866 = ~n35863 & n35865;
  assign n35867 = n6198 & ~n35866;
  assign n35868 = pi222 & ~n35867;
  assign n35869 = ~n35859 & n35868;
  assign n35870 = n16906 & n35632;
  assign n35871 = ~n35548 & ~n35870;
  assign n35872 = n6198 & ~n35871;
  assign n35873 = ~n16261 & n35524;
  assign n35874 = ~pi680 & n35873;
  assign n35875 = pi661 & ~n35874;
  assign n35876 = pi614 & ~pi616;
  assign n35877 = ~n16895 & n35876;
  assign n35878 = ~n16899 & ~n35877;
  assign n35879 = ~n16480 & ~n16978;
  assign n35880 = pi616 & n35879;
  assign n35881 = pi680 & ~n35880;
  assign n35882 = n35878 & n35881;
  assign n35883 = n35875 & ~n35882;
  assign n35884 = ~pi661 & ~n35873;
  assign n35885 = ~n16224 & n35524;
  assign n35886 = n6188 & ~n35885;
  assign n35887 = ~n35884 & ~n35886;
  assign n35888 = ~n35883 & n35887;
  assign n35889 = ~n6198 & n35888;
  assign n35890 = ~pi222 & ~n35889;
  assign n35891 = ~n35872 & n35890;
  assign n35892 = ~n35869 & ~n35891;
  assign n35893 = pi215 & n35892;
  assign n35894 = pi299 & ~n35893;
  assign n35895 = ~n35848 & n35894;
  assign n35896 = n35632 & ~n35778;
  assign n35897 = ~n35524 & ~n35632;
  assign n35898 = ~pi222 & ~n35897;
  assign n35899 = ~n35896 & n35898;
  assign n35900 = ~n3332 & ~n35899;
  assign n35901 = ~n6236 & n35828;
  assign n35902 = n6236 & n35841;
  assign n35903 = pi224 & ~n35902;
  assign n35904 = ~n35901 & n35903;
  assign n35905 = ~n35900 & ~n35904;
  assign n35906 = ~n6236 & n35809;
  assign n35907 = n6236 & n35819;
  assign n35908 = pi222 & ~n35907;
  assign n35909 = ~n35906 & n35908;
  assign n35910 = ~n35905 & ~n35909;
  assign n35911 = ~pi223 & ~n35910;
  assign n35912 = n6236 & ~n35871;
  assign n35913 = ~n6236 & n35888;
  assign n35914 = ~pi222 & ~n35913;
  assign n35915 = ~n35912 & n35914;
  assign n35916 = ~n6236 & ~n35858;
  assign n35917 = n6236 & ~n35866;
  assign n35918 = pi222 & ~n35917;
  assign n35919 = ~n35916 & n35918;
  assign n35920 = pi223 & ~n35919;
  assign n35921 = ~n35915 & n35920;
  assign n35922 = ~pi299 & ~n35921;
  assign n35923 = ~n35911 & n35922;
  assign n35924 = pi39 & ~n35923;
  assign n35925 = ~n35895 & n35924;
  assign n35926 = ~pi616 & n16458;
  assign n35927 = n18300 & ~n35632;
  assign n35928 = n16716 & ~n16810;
  assign n35929 = ~n35927 & ~n35928;
  assign n35930 = ~n35926 & n35929;
  assign n35931 = pi222 & ~n35930;
  assign n35932 = pi616 & n16458;
  assign n35933 = ~pi222 & ~n35932;
  assign n35934 = pi661 & n18301;
  assign n35935 = n35933 & ~n35934;
  assign n35936 = ~n35931 & ~n35935;
  assign n35937 = pi299 & ~n35936;
  assign n35938 = pi616 & n16453;
  assign n35939 = ~pi222 & ~n35938;
  assign n35940 = pi661 & n18293;
  assign n35941 = n35939 & ~n35940;
  assign n35942 = ~pi616 & n16453;
  assign n35943 = n18292 & ~n35632;
  assign n35944 = n16710 & ~n16810;
  assign n35945 = ~n35943 & ~n35944;
  assign n35946 = ~n35942 & n35945;
  assign n35947 = pi222 & ~n35946;
  assign n35948 = ~n35941 & ~n35947;
  assign n35949 = ~pi299 & ~n35948;
  assign n35950 = ~pi39 & ~n35949;
  assign n35951 = ~n35937 & n35950;
  assign n35952 = ~pi38 & ~n35951;
  assign n35953 = ~n35925 & n35952;
  assign n35954 = n16212 & n16952;
  assign n35955 = ~pi222 & ~pi616;
  assign n35956 = ~pi39 & pi616;
  assign n35957 = n35632 & n35956;
  assign n35958 = ~n35955 & ~n35957;
  assign n35959 = n35954 & ~n35958;
  assign n35960 = ~pi616 & ~n16814;
  assign n35961 = ~n35775 & ~n35960;
  assign n35962 = n16508 & n35961;
  assign n35963 = ~n35582 & ~n35962;
  assign n35964 = ~n35959 & ~n35963;
  assign n35965 = pi38 & ~n35964;
  assign n35966 = ~n35953 & ~n35965;
  assign n35967 = n10020 & n35966;
  assign n35968 = ~n35477 & ~n35967;
  assign n35969 = ~pi625 & n35968;
  assign n35970 = ~pi1153 & ~n35969;
  assign n35971 = ~n35774 & n35970;
  assign n35972 = ~pi608 & ~n35729;
  assign n35973 = ~n35971 & n35972;
  assign n35974 = ~pi625 & n35588;
  assign n35975 = pi625 & n35968;
  assign n35976 = ~n35974 & ~n35975;
  assign n35977 = pi1153 & n35976;
  assign n35978 = ~n35733 & ~n35977;
  assign n35979 = pi608 & n35978;
  assign n35980 = ~n35973 & ~n35979;
  assign n35981 = pi778 & ~n35980;
  assign n35982 = ~pi778 & n35968;
  assign n35983 = ~n35981 & ~n35982;
  assign n35984 = ~pi609 & ~n35983;
  assign n35985 = ~pi1155 & ~n35984;
  assign n35986 = ~n35773 & n35985;
  assign n35987 = ~pi660 & ~n35596;
  assign n35988 = ~n35986 & n35987;
  assign n35989 = ~pi609 & n35736;
  assign n35990 = pi609 & ~n35983;
  assign n35991 = ~n35989 & ~n35990;
  assign n35992 = pi1155 & n35991;
  assign n35993 = ~n35600 & ~n35992;
  assign n35994 = pi660 & n35993;
  assign n35995 = ~n35988 & ~n35994;
  assign n35996 = pi785 & ~n35995;
  assign n35997 = ~pi785 & ~n35983;
  assign n35998 = ~n35996 & ~n35997;
  assign n35999 = ~pi618 & ~n35998;
  assign n36000 = ~pi1154 & ~n35999;
  assign n36001 = ~n35772 & n36000;
  assign n36002 = ~pi627 & ~n35608;
  assign n36003 = ~n36001 & n36002;
  assign n36004 = ~pi618 & n35739;
  assign n36005 = pi618 & ~n35998;
  assign n36006 = ~n36004 & ~n36005;
  assign n36007 = pi1154 & n36006;
  assign n36008 = ~n35612 & ~n36007;
  assign n36009 = pi627 & n36008;
  assign n36010 = ~n36003 & ~n36009;
  assign n36011 = pi781 & ~n36010;
  assign n36012 = ~pi781 & ~n35998;
  assign n36013 = ~n36011 & ~n36012;
  assign n36014 = ~pi789 & n36013;
  assign n36015 = ~n35771 & ~n36014;
  assign n36016 = ~pi619 & ~n36013;
  assign n36017 = pi619 & n35742;
  assign n36018 = ~pi1159 & ~n36017;
  assign n36019 = ~n36016 & n36018;
  assign n36020 = ~pi648 & ~n36019;
  assign n36021 = ~n35620 & n36020;
  assign n36022 = ~pi619 & n35742;
  assign n36023 = pi619 & ~n36013;
  assign n36024 = ~n36022 & ~n36023;
  assign n36025 = pi1159 & n36024;
  assign n36026 = ~n35624 & ~n36025;
  assign n36027 = pi648 & n36026;
  assign n36028 = ~n36021 & ~n36027;
  assign n36029 = pi789 & n36028;
  assign n36030 = n36015 & ~n36029;
  assign n36031 = ~n35770 & ~n36030;
  assign n36032 = n19788 & n36031;
  assign n36033 = ~n35756 & ~n36032;
  assign n36034 = n19637 & ~n36033;
  assign n36035 = ~n18744 & ~n35745;
  assign n36036 = n17451 & ~n35475;
  assign n36037 = ~n36035 & ~n36036;
  assign n36038 = pi647 & ~n36037;
  assign n36039 = ~pi647 & ~n35475;
  assign n36040 = pi1157 & ~n36039;
  assign n36041 = ~n36038 & n36040;
  assign n36042 = ~pi630 & n36041;
  assign n36043 = ~n16124 & n35629;
  assign n36044 = n16124 & n35475;
  assign n36045 = ~n36043 & ~n36044;
  assign n36046 = ~n19987 & ~n36045;
  assign n36047 = ~pi647 & ~n36037;
  assign n36048 = pi647 & ~n35475;
  assign n36049 = ~pi1157 & ~n36048;
  assign n36050 = ~n36047 & n36049;
  assign n36051 = pi630 & n36050;
  assign n36052 = ~n36046 & ~n36051;
  assign n36053 = ~n36042 & n36052;
  assign n36054 = pi787 & ~n36053;
  assign n36055 = ~n36034 & ~n36054;
  assign n36056 = pi644 & n36055;
  assign n36057 = ~pi787 & n36037;
  assign n36058 = ~n36041 & ~n36050;
  assign n36059 = pi787 & ~n36058;
  assign n36060 = ~n36057 & ~n36059;
  assign n36061 = ~pi644 & n36060;
  assign n36062 = pi715 & ~n36061;
  assign n36063 = ~n36056 & n36062;
  assign n36064 = n17247 & ~n35475;
  assign n36065 = ~n17247 & n36045;
  assign n36066 = ~n36064 & ~n36065;
  assign n36067 = pi644 & ~n36066;
  assign n36068 = ~pi644 & ~n35475;
  assign n36069 = ~pi715 & ~n36068;
  assign n36070 = ~n36067 & n36069;
  assign n36071 = pi1160 & ~n36070;
  assign n36072 = ~n36063 & n36071;
  assign n36073 = pi644 & ~n35475;
  assign n36074 = ~pi644 & ~n36066;
  assign n36075 = pi715 & ~n36074;
  assign n36076 = ~n36073 & n36075;
  assign n36077 = pi644 & n36060;
  assign n36078 = ~pi644 & n36055;
  assign n36079 = ~pi715 & ~n36078;
  assign n36080 = ~n36077 & n36079;
  assign n36081 = ~pi1160 & ~n36080;
  assign n36082 = ~n36076 & n36081;
  assign n36083 = ~n36072 & ~n36082;
  assign n36084 = pi790 & ~n36083;
  assign n36085 = ~pi790 & n36055;
  assign n36086 = ~n36084 & ~n36085;
  assign n36087 = ~po1038 & ~n36086;
  assign n36088 = ~pi222 & po1038;
  assign po379 = ~n36087 & ~n36088;
  assign n36090 = ~pi299 & ~n16269;
  assign n36091 = ~n16354 & ~n36090;
  assign n36092 = pi39 & n36091;
  assign n36093 = ~n17520 & ~n36092;
  assign n36094 = n2575 & n36093;
  assign n36095 = n18119 & ~n36094;
  assign n36096 = pi223 & ~n36095;
  assign n36097 = ~n32843 & ~n36096;
  assign n36098 = n16593 & ~n36096;
  assign n36099 = pi223 & ~n10020;
  assign n36100 = pi680 & pi681;
  assign n36101 = n16728 & ~n36100;
  assign n36102 = pi223 & n16710;
  assign n36103 = ~pi223 & ~n16728;
  assign n36104 = ~pi299 & ~n36103;
  assign n36105 = ~n36102 & n36104;
  assign n36106 = ~n36101 & n36105;
  assign n36107 = ~pi39 & ~n36106;
  assign n36108 = n16733 & ~n36100;
  assign n36109 = pi223 & n16716;
  assign n36110 = ~pi223 & ~n16733;
  assign n36111 = pi299 & ~n36110;
  assign n36112 = ~n36109 & n36111;
  assign n36113 = ~n36108 & n36112;
  assign n36114 = n36107 & ~n36113;
  assign n36115 = pi223 & ~n16207;
  assign n36116 = n2527 & ~n36115;
  assign n36117 = pi681 & n16630;
  assign n36118 = n36116 & ~n36117;
  assign n36119 = pi681 & n35661;
  assign n36120 = ~n6198 & ~n36119;
  assign n36121 = ~n16607 & n36100;
  assign n36122 = n6198 & ~n36121;
  assign n36123 = ~pi223 & ~n36122;
  assign n36124 = ~n36120 & n36123;
  assign n36125 = pi681 & ~n16657;
  assign n36126 = ~n16326 & ~n36125;
  assign n36127 = n6198 & n36126;
  assign n36128 = ~pi681 & ~n16297;
  assign n36129 = pi681 & ~n35655;
  assign n36130 = ~n36128 & ~n36129;
  assign n36131 = ~n6198 & n36130;
  assign n36132 = pi223 & ~n36131;
  assign n36133 = ~n36127 & n36132;
  assign n36134 = ~n2527 & ~n36133;
  assign n36135 = ~n36124 & n36134;
  assign n36136 = ~n36118 & ~n36135;
  assign n36137 = ~pi215 & ~n36136;
  assign n36138 = ~pi223 & pi681;
  assign n36139 = n16634 & n36138;
  assign n36140 = pi681 & ~n16679;
  assign n36141 = ~n16266 & ~n36140;
  assign n36142 = ~n6198 & n36141;
  assign n36143 = pi681 & ~n35682;
  assign n36144 = ~n16249 & ~n36143;
  assign n36145 = n6198 & n36144;
  assign n36146 = pi223 & ~n36145;
  assign n36147 = ~n36142 & n36146;
  assign n36148 = pi215 & ~n36147;
  assign n36149 = ~n36139 & n36148;
  assign n36150 = pi299 & ~n36149;
  assign n36151 = ~n36137 & n36150;
  assign n36152 = n2607 & ~n36117;
  assign n36153 = ~n6236 & n36119;
  assign n36154 = n6236 & n36121;
  assign n36155 = ~n2607 & ~n36154;
  assign n36156 = ~n36153 & n36155;
  assign n36157 = ~n36152 & ~n36156;
  assign n36158 = ~pi223 & ~n36157;
  assign n36159 = ~n6236 & ~n36141;
  assign n36160 = n6236 & ~n36144;
  assign n36161 = ~n36159 & ~n36160;
  assign n36162 = pi223 & n36161;
  assign n36163 = ~pi299 & ~n36162;
  assign n36164 = ~n36158 & n36163;
  assign n36165 = pi39 & ~n36164;
  assign n36166 = ~n36151 & n36165;
  assign n36167 = ~n36114 & ~n36166;
  assign n36168 = ~pi38 & ~n36167;
  assign n36169 = pi681 & n16743;
  assign n36170 = pi223 & ~n16508;
  assign n36171 = pi38 & ~n36170;
  assign n36172 = ~n36169 & n36171;
  assign n36173 = ~n36168 & ~n36172;
  assign n36174 = n10020 & n36173;
  assign n36175 = ~n36099 & ~n36174;
  assign n36176 = ~pi778 & ~n36175;
  assign n36177 = pi625 & n36175;
  assign n36178 = ~pi625 & ~n36096;
  assign n36179 = pi1153 & ~n36178;
  assign n36180 = ~n36177 & n36179;
  assign n36181 = ~pi625 & n36175;
  assign n36182 = pi625 & ~n36096;
  assign n36183 = ~pi1153 & ~n36182;
  assign n36184 = ~n36181 & n36183;
  assign n36185 = ~n36180 & ~n36184;
  assign n36186 = pi778 & ~n36185;
  assign n36187 = ~n36176 & ~n36186;
  assign n36188 = ~n16593 & n36187;
  assign n36189 = ~n36098 & ~n36188;
  assign n36190 = ~n16589 & n36189;
  assign n36191 = n16589 & n36096;
  assign n36192 = ~n36190 & ~n36191;
  assign n36193 = ~n17159 & n36192;
  assign n36194 = ~n17183 & n36193;
  assign n36195 = ~n36097 & ~n36194;
  assign n36196 = ~n18744 & ~n36195;
  assign n36197 = n17451 & ~n36096;
  assign n36198 = ~n36196 & ~n36197;
  assign n36199 = pi647 & ~n36198;
  assign n36200 = ~pi647 & ~n36096;
  assign n36201 = pi1157 & ~n36200;
  assign n36202 = ~n36199 & n36201;
  assign n36203 = ~pi630 & n36202;
  assign n36204 = n17355 & ~n36096;
  assign n36205 = n16521 & ~n36096;
  assign n36206 = pi642 & n16465;
  assign n36207 = n36116 & ~n36206;
  assign n36208 = pi642 & n16393;
  assign n36209 = n35121 & ~n36208;
  assign n36210 = pi642 & ~n16394;
  assign n36211 = ~n16304 & ~n36210;
  assign n36212 = n6184 & n36211;
  assign n36213 = ~n36209 & ~n36212;
  assign n36214 = pi681 & n36213;
  assign n36215 = ~pi661 & n16253;
  assign n36216 = ~n36213 & ~n36215;
  assign n36217 = ~n16389 & ~n35119;
  assign n36218 = n36215 & ~n36217;
  assign n36219 = ~pi681 & ~n36218;
  assign n36220 = ~n36216 & n36219;
  assign n36221 = n6198 & ~n36220;
  assign n36222 = ~n36214 & n36221;
  assign n36223 = pi642 & ~n16861;
  assign n36224 = ~pi642 & n16294;
  assign n36225 = ~n36223 & ~n36224;
  assign n36226 = pi681 & ~n36225;
  assign n36227 = ~n36215 & n36225;
  assign n36228 = ~n16289 & ~n36208;
  assign n36229 = n36215 & n36228;
  assign n36230 = ~pi681 & ~n36229;
  assign n36231 = ~n36227 & n36230;
  assign n36232 = ~n6198 & ~n36231;
  assign n36233 = ~n36226 & n36232;
  assign n36234 = pi223 & ~n36233;
  assign n36235 = ~n36222 & n36234;
  assign n36236 = ~n16292 & n36208;
  assign n36237 = pi681 & ~n36236;
  assign n36238 = ~n36215 & n36236;
  assign n36239 = pi642 & n36215;
  assign n36240 = n16809 & n36239;
  assign n36241 = ~pi681 & ~n36240;
  assign n36242 = ~n36238 & n36241;
  assign n36243 = ~n36237 & ~n36242;
  assign n36244 = pi947 & ~n36243;
  assign n36245 = ~n20340 & n36243;
  assign n36246 = n36206 & ~n36215;
  assign n36247 = ~pi681 & ~n36246;
  assign n36248 = n16463 & n36239;
  assign n36249 = n36247 & ~n36248;
  assign n36250 = pi681 & ~n36206;
  assign n36251 = ~n36249 & ~n36250;
  assign n36252 = n20340 & n36251;
  assign n36253 = ~pi947 & ~n36252;
  assign n36254 = ~n36245 & n36253;
  assign n36255 = ~pi223 & ~n36254;
  assign n36256 = ~n36244 & n36255;
  assign n36257 = ~n2527 & ~n36256;
  assign n36258 = ~n36235 & n36257;
  assign n36259 = ~pi215 & ~n36258;
  assign n36260 = ~n36207 & n36259;
  assign n36261 = n16479 & n36239;
  assign n36262 = n36247 & ~n36261;
  assign n36263 = n6198 & ~n36262;
  assign n36264 = n36206 & n36263;
  assign n36265 = pi642 & ~n16420;
  assign n36266 = ~n16224 & ~n36265;
  assign n36267 = n36215 & n36266;
  assign n36268 = ~pi681 & ~n36267;
  assign n36269 = n16261 & n36268;
  assign n36270 = ~n36262 & ~n36269;
  assign n36271 = pi642 & n16480;
  assign n36272 = pi681 & ~n36271;
  assign n36273 = n36270 & ~n36272;
  assign n36274 = ~n20340 & n36273;
  assign n36275 = ~pi947 & ~n36274;
  assign n36276 = ~n36264 & n36275;
  assign n36277 = pi947 & ~n36273;
  assign n36278 = ~pi223 & ~n36277;
  assign n36279 = ~n36276 & n36278;
  assign n36280 = n16234 & ~n36206;
  assign n36281 = pi681 & ~n36280;
  assign n36282 = ~n36215 & n36280;
  assign n36283 = ~pi681 & ~n36282;
  assign n36284 = n16212 & ~n36208;
  assign n36285 = n16227 & n36284;
  assign n36286 = n36215 & n36285;
  assign n36287 = n36283 & ~n36286;
  assign n36288 = ~n36281 & ~n36287;
  assign n36289 = n6198 & n36288;
  assign n36290 = ~n16229 & n16392;
  assign n36291 = ~n16261 & ~n36290;
  assign n36292 = ~n36265 & n36291;
  assign n36293 = ~n36215 & n36292;
  assign n36294 = n36268 & ~n36293;
  assign n36295 = pi681 & ~n36292;
  assign n36296 = ~n36294 & ~n36295;
  assign n36297 = ~n6198 & n36296;
  assign n36298 = pi223 & ~n36297;
  assign n36299 = ~n36289 & n36298;
  assign n36300 = ~n36279 & ~n36299;
  assign n36301 = pi215 & ~n36300;
  assign n36302 = pi299 & ~n36301;
  assign n36303 = ~n36260 & n36302;
  assign n36304 = n6236 & n36251;
  assign n36305 = ~n6236 & n36243;
  assign n36306 = ~n2607 & ~n36305;
  assign n36307 = ~n36304 & n36306;
  assign n36308 = n2607 & ~n36206;
  assign n36309 = ~pi223 & ~n36308;
  assign n36310 = ~n36307 & n36309;
  assign n36311 = ~n6236 & n36296;
  assign n36312 = n6236 & n36288;
  assign n36313 = ~n36311 & ~n36312;
  assign n36314 = pi223 & n36313;
  assign n36315 = ~pi299 & ~n36314;
  assign n36316 = ~n36310 & n36315;
  assign n36317 = pi39 & ~n36316;
  assign n36318 = ~n36303 & n36317;
  assign n36319 = ~pi223 & pi642;
  assign n36320 = n16453 & n36319;
  assign n36321 = ~pi299 & ~n36320;
  assign n36322 = ~pi642 & n16453;
  assign n36323 = pi223 & ~n36322;
  assign n36324 = n16378 & n36323;
  assign n36325 = n36321 & ~n36324;
  assign n36326 = n16458 & n36319;
  assign n36327 = pi299 & ~n36326;
  assign n36328 = n6183 & n16457;
  assign n36329 = pi223 & ~n36328;
  assign n36330 = ~n16365 & n36329;
  assign n36331 = n36327 & ~n36330;
  assign n36332 = ~pi39 & ~n36331;
  assign n36333 = ~n36325 & n36332;
  assign n36334 = ~pi38 & ~n36333;
  assign n36335 = ~n36318 & n36334;
  assign n36336 = pi39 & pi223;
  assign n36337 = pi38 & ~n36336;
  assign n36338 = ~pi223 & ~n16212;
  assign n36339 = ~pi39 & ~n36338;
  assign n36340 = ~n36284 & n36339;
  assign n36341 = n36337 & ~n36340;
  assign n36342 = ~n36335 & ~n36341;
  assign n36343 = n10020 & n36342;
  assign n36344 = ~n36099 & ~n36343;
  assign n36345 = ~n16521 & n36344;
  assign n36346 = ~n36205 & ~n36345;
  assign n36347 = ~pi785 & n36346;
  assign n36348 = pi609 & ~n36346;
  assign n36349 = ~pi609 & ~n36096;
  assign n36350 = pi1155 & ~n36349;
  assign n36351 = ~n36348 & n36350;
  assign n36352 = ~pi609 & ~n36346;
  assign n36353 = pi609 & ~n36096;
  assign n36354 = ~pi1155 & ~n36353;
  assign n36355 = ~n36352 & n36354;
  assign n36356 = ~n36351 & ~n36355;
  assign n36357 = pi785 & ~n36356;
  assign n36358 = ~n36347 & ~n36357;
  assign n36359 = ~pi781 & ~n36358;
  assign n36360 = pi618 & n36358;
  assign n36361 = ~pi618 & ~n36096;
  assign n36362 = pi1154 & ~n36361;
  assign n36363 = ~n36360 & n36362;
  assign n36364 = ~pi618 & n36358;
  assign n36365 = pi618 & ~n36096;
  assign n36366 = ~pi1154 & ~n36365;
  assign n36367 = ~n36364 & n36366;
  assign n36368 = ~n36363 & ~n36367;
  assign n36369 = pi781 & ~n36368;
  assign n36370 = ~n36359 & ~n36369;
  assign n36371 = ~pi789 & ~n36370;
  assign n36372 = pi619 & n36370;
  assign n36373 = ~pi619 & ~n36096;
  assign n36374 = pi1159 & ~n36373;
  assign n36375 = ~n36372 & n36374;
  assign n36376 = ~pi619 & n36370;
  assign n36377 = pi619 & ~n36096;
  assign n36378 = ~pi1159 & ~n36377;
  assign n36379 = ~n36376 & n36378;
  assign n36380 = ~n36375 & ~n36379;
  assign n36381 = pi789 & ~n36380;
  assign n36382 = ~n36371 & ~n36381;
  assign n36383 = ~n17355 & n36382;
  assign n36384 = ~n36204 & ~n36383;
  assign n36385 = ~n16124 & n36384;
  assign n36386 = n16124 & n36096;
  assign n36387 = ~n36385 & ~n36386;
  assign n36388 = ~n19987 & ~n36387;
  assign n36389 = ~pi647 & ~n36198;
  assign n36390 = pi647 & ~n36096;
  assign n36391 = ~pi1157 & ~n36390;
  assign n36392 = ~n36389 & n36391;
  assign n36393 = pi630 & n36392;
  assign n36394 = ~n36388 & ~n36393;
  assign n36395 = ~n36203 & n36394;
  assign n36396 = pi787 & ~n36395;
  assign n36397 = ~n19999 & n36384;
  assign n36398 = pi628 & ~n36195;
  assign n36399 = ~pi628 & ~n36096;
  assign n36400 = n16121 & ~n36399;
  assign n36401 = ~n36398 & n36400;
  assign n36402 = ~pi628 & ~n36195;
  assign n36403 = pi628 & ~n36096;
  assign n36404 = n16122 & ~n36403;
  assign n36405 = ~n36402 & n36404;
  assign n36406 = ~n36401 & ~n36405;
  assign n36407 = ~n36397 & n36406;
  assign n36408 = ~n19788 & n36407;
  assign n36409 = pi792 & ~n36407;
  assign n36410 = n17159 & ~n36096;
  assign n36411 = ~n36193 & ~n36410;
  assign n36412 = n17350 & ~n36411;
  assign n36413 = pi626 & ~n36382;
  assign n36414 = ~pi626 & n36096;
  assign n36415 = n17180 & ~n36414;
  assign n36416 = ~n36413 & n36415;
  assign n36417 = ~n36412 & ~n36416;
  assign n36418 = ~pi626 & ~n36382;
  assign n36419 = pi626 & n36096;
  assign n36420 = n17181 & ~n36419;
  assign n36421 = ~n36418 & n36420;
  assign n36422 = n36417 & ~n36421;
  assign n36423 = pi788 & ~n36422;
  assign n36424 = pi618 & ~n36189;
  assign n36425 = pi609 & n36187;
  assign n36426 = pi625 & n36344;
  assign n36427 = ~n36100 & ~n36226;
  assign n36428 = n16392 & ~n35794;
  assign n36429 = pi642 & ~n35786;
  assign n36430 = ~pi642 & ~n6184;
  assign n36431 = n35788 & n36430;
  assign n36432 = pi680 & ~n36431;
  assign n36433 = ~n36429 & n36432;
  assign n36434 = ~n36428 & n36433;
  assign n36435 = ~n36427 & ~n36434;
  assign n36436 = n36232 & ~n36435;
  assign n36437 = ~n36100 & ~n36214;
  assign n36438 = pi642 & ~n17022;
  assign n36439 = ~n16820 & ~n36438;
  assign n36440 = n6184 & ~n36439;
  assign n36441 = ~pi642 & ~n16775;
  assign n36442 = ~n16952 & ~n36441;
  assign n36443 = n35121 & n36442;
  assign n36444 = pi680 & ~n36443;
  assign n36445 = ~n16208 & n36444;
  assign n36446 = ~n16231 & n36445;
  assign n36447 = ~n36440 & n36446;
  assign n36448 = ~n36437 & ~n36447;
  assign n36449 = n36221 & ~n36448;
  assign n36450 = pi223 & ~n36449;
  assign n36451 = ~n36436 & n36450;
  assign n36452 = ~pi680 & ~n36206;
  assign n36453 = pi642 & ~n16953;
  assign n36454 = n6184 & ~n36453;
  assign n36455 = ~pi642 & ~n16883;
  assign n36456 = n36454 & ~n36455;
  assign n36457 = n36444 & ~n36456;
  assign n36458 = ~n36452 & ~n36457;
  assign n36459 = pi681 & ~n36458;
  assign n36460 = ~n36249 & ~n36459;
  assign n36461 = n6198 & ~n36460;
  assign n36462 = ~n36100 & ~n36237;
  assign n36463 = pi642 & n16943;
  assign n36464 = pi680 & ~n36463;
  assign n36465 = ~n16867 & n36464;
  assign n36466 = ~n16862 & n36430;
  assign n36467 = n36465 & ~n36466;
  assign n36468 = ~n36462 & ~n36467;
  assign n36469 = ~n36242 & ~n36468;
  assign n36470 = ~n6198 & ~n36469;
  assign n36471 = ~pi223 & ~n36470;
  assign n36472 = ~n36461 & n36471;
  assign n36473 = ~n36451 & ~n36472;
  assign n36474 = ~n2527 & n36473;
  assign n36475 = ~n36100 & n36208;
  assign n36476 = ~n35954 & ~n36441;
  assign n36477 = n36100 & n36476;
  assign n36478 = ~n36475 & ~n36477;
  assign n36479 = n16207 & ~n36478;
  assign n36480 = n36116 & ~n36479;
  assign n36481 = ~pi215 & ~n36480;
  assign n36482 = ~n36474 & n36481;
  assign n36483 = ~n36100 & ~n36281;
  assign n36484 = ~pi614 & n16786;
  assign n36485 = ~n36438 & ~n36484;
  assign n36486 = ~pi616 & ~n36485;
  assign n36487 = n36446 & ~n36486;
  assign n36488 = ~n36483 & ~n36487;
  assign n36489 = ~n36287 & ~n36488;
  assign n36490 = n6198 & ~n36489;
  assign n36491 = ~n36100 & ~n36295;
  assign n36492 = ~n6184 & n16799;
  assign n36493 = pi642 & ~n35850;
  assign n36494 = pi680 & ~n36493;
  assign n36495 = ~n16800 & n36494;
  assign n36496 = ~n36492 & n36495;
  assign n36497 = ~n36491 & ~n36496;
  assign n36498 = ~n36294 & ~n36497;
  assign n36499 = ~n6198 & ~n36498;
  assign n36500 = pi223 & ~n36499;
  assign n36501 = ~n36490 & n36500;
  assign n36502 = ~n36100 & ~n36272;
  assign n36503 = pi642 & n35879;
  assign n36504 = ~n16895 & n36430;
  assign n36505 = n16896 & n16978;
  assign n36506 = n16392 & ~n36505;
  assign n36507 = pi680 & ~n36506;
  assign n36508 = ~n36504 & n36507;
  assign n36509 = ~n36503 & n36508;
  assign n36510 = ~n36502 & ~n36509;
  assign n36511 = ~n6198 & ~n36510;
  assign n36512 = n36270 & n36511;
  assign n36513 = ~n16897 & n36454;
  assign n36514 = n36444 & ~n36513;
  assign n36515 = ~n36452 & ~n36514;
  assign n36516 = pi681 & ~n36515;
  assign n36517 = n36263 & ~n36516;
  assign n36518 = ~pi223 & ~n36517;
  assign n36519 = ~n36512 & n36518;
  assign n36520 = ~n36501 & ~n36519;
  assign n36521 = pi215 & n36520;
  assign n36522 = pi299 & ~n36521;
  assign n36523 = ~n36482 & n36522;
  assign n36524 = ~n6236 & n36469;
  assign n36525 = n6236 & n36460;
  assign n36526 = ~n2607 & ~n36525;
  assign n36527 = ~n36524 & n36526;
  assign n36528 = n2607 & ~n36479;
  assign n36529 = ~pi223 & ~n36528;
  assign n36530 = ~n36527 & n36529;
  assign n36531 = ~n6236 & n36498;
  assign n36532 = n6236 & n36489;
  assign n36533 = ~n36531 & ~n36532;
  assign n36534 = pi223 & n36533;
  assign n36535 = ~pi299 & ~n36534;
  assign n36536 = ~n36530 & n36535;
  assign n36537 = pi39 & ~n36536;
  assign n36538 = ~n36523 & n36537;
  assign n36539 = n18301 & n36138;
  assign n36540 = n36327 & ~n36539;
  assign n36541 = n18300 & ~n36100;
  assign n36542 = ~n35928 & n36329;
  assign n36543 = ~n36541 & n36542;
  assign n36544 = n36540 & ~n36543;
  assign n36545 = n18293 & n36138;
  assign n36546 = n18292 & ~n36100;
  assign n36547 = ~n35944 & n36323;
  assign n36548 = ~n36546 & n36547;
  assign n36549 = ~n36545 & ~n36548;
  assign n36550 = n36321 & n36549;
  assign n36551 = ~pi39 & ~n36550;
  assign n36552 = ~n36544 & n36551;
  assign n36553 = ~pi38 & ~n36552;
  assign n36554 = ~n36538 & n36553;
  assign n36555 = ~n36170 & n36478;
  assign n36556 = n36339 & ~n36555;
  assign n36557 = n36337 & ~n36556;
  assign n36558 = ~n36554 & ~n36557;
  assign n36559 = n10020 & n36558;
  assign n36560 = ~n36099 & ~n36559;
  assign n36561 = ~pi625 & n36560;
  assign n36562 = ~pi1153 & ~n36561;
  assign n36563 = ~n36426 & n36562;
  assign n36564 = ~pi608 & ~n36563;
  assign n36565 = ~n36180 & n36564;
  assign n36566 = ~pi625 & n36344;
  assign n36567 = pi625 & n36560;
  assign n36568 = ~n36566 & ~n36567;
  assign n36569 = pi1153 & n36568;
  assign n36570 = ~n36184 & ~n36569;
  assign n36571 = pi608 & n36570;
  assign n36572 = ~n36565 & ~n36571;
  assign n36573 = pi778 & ~n36572;
  assign n36574 = ~pi778 & n36560;
  assign n36575 = ~n36573 & ~n36574;
  assign n36576 = ~pi609 & ~n36575;
  assign n36577 = ~pi1155 & ~n36576;
  assign n36578 = ~n36425 & n36577;
  assign n36579 = ~pi660 & ~n36351;
  assign n36580 = ~n36578 & n36579;
  assign n36581 = ~pi609 & n36187;
  assign n36582 = pi609 & ~n36575;
  assign n36583 = ~n36581 & ~n36582;
  assign n36584 = pi1155 & n36583;
  assign n36585 = ~n36355 & ~n36584;
  assign n36586 = pi660 & n36585;
  assign n36587 = ~n36580 & ~n36586;
  assign n36588 = pi785 & ~n36587;
  assign n36589 = ~pi785 & ~n36575;
  assign n36590 = ~n36588 & ~n36589;
  assign n36591 = ~pi618 & ~n36590;
  assign n36592 = ~pi1154 & ~n36591;
  assign n36593 = ~n36424 & n36592;
  assign n36594 = ~pi627 & ~n36363;
  assign n36595 = ~n36593 & n36594;
  assign n36596 = ~pi618 & ~n36189;
  assign n36597 = pi618 & ~n36590;
  assign n36598 = ~n36596 & ~n36597;
  assign n36599 = pi1154 & n36598;
  assign n36600 = ~n36367 & ~n36599;
  assign n36601 = pi627 & n36600;
  assign n36602 = ~n36595 & ~n36601;
  assign n36603 = pi781 & ~n36602;
  assign n36604 = ~pi781 & ~n36590;
  assign n36605 = ~n36603 & ~n36604;
  assign n36606 = ~pi619 & ~n36605;
  assign n36607 = pi619 & n36192;
  assign n36608 = ~pi1159 & ~n36607;
  assign n36609 = ~n36606 & n36608;
  assign n36610 = ~pi648 & ~n36609;
  assign n36611 = ~n36375 & n36610;
  assign n36612 = ~pi619 & n36192;
  assign n36613 = pi619 & ~n36605;
  assign n36614 = ~n36612 & ~n36613;
  assign n36615 = pi1159 & n36614;
  assign n36616 = ~n36379 & ~n36615;
  assign n36617 = pi648 & n36616;
  assign n36618 = ~n36611 & ~n36617;
  assign n36619 = pi789 & n36618;
  assign n36620 = ~pi789 & n36605;
  assign n36621 = n17356 & ~n36620;
  assign n36622 = ~n36619 & n36621;
  assign n36623 = ~n36423 & ~n36622;
  assign n36624 = ~n36409 & ~n36623;
  assign n36625 = ~n36408 & ~n36624;
  assign n36626 = n19637 & n36625;
  assign n36627 = ~n36396 & ~n36626;
  assign n36628 = pi644 & n36627;
  assign n36629 = ~pi787 & n36198;
  assign n36630 = ~n36202 & ~n36392;
  assign n36631 = pi787 & ~n36630;
  assign n36632 = ~n36629 & ~n36631;
  assign n36633 = ~pi644 & n36632;
  assign n36634 = pi715 & ~n36633;
  assign n36635 = ~n36628 & n36634;
  assign n36636 = n17247 & ~n36096;
  assign n36637 = ~n17247 & n36387;
  assign n36638 = ~n36636 & ~n36637;
  assign n36639 = pi644 & ~n36638;
  assign n36640 = ~pi644 & ~n36096;
  assign n36641 = ~pi715 & ~n36640;
  assign n36642 = ~n36639 & n36641;
  assign n36643 = pi1160 & ~n36642;
  assign n36644 = ~n36635 & n36643;
  assign n36645 = pi644 & ~n36096;
  assign n36646 = ~pi644 & ~n36638;
  assign n36647 = pi715 & ~n36646;
  assign n36648 = ~n36645 & n36647;
  assign n36649 = pi644 & n36632;
  assign n36650 = ~pi644 & n36627;
  assign n36651 = ~pi715 & ~n36650;
  assign n36652 = ~n36649 & n36651;
  assign n36653 = ~pi1160 & ~n36652;
  assign n36654 = ~n36648 & n36653;
  assign n36655 = ~n36644 & ~n36654;
  assign n36656 = pi790 & ~n36655;
  assign n36657 = ~pi790 & n36627;
  assign n36658 = ~n36656 & ~n36657;
  assign n36659 = ~po1038 & ~n36658;
  assign n36660 = ~pi223 & po1038;
  assign po380 = ~n36659 & ~n36660;
  assign n36662 = pi224 & ~n35474;
  assign n36663 = n17355 & ~n36662;
  assign n36664 = pi224 & ~n10020;
  assign n36665 = pi224 & ~n16508;
  assign n36666 = pi38 & ~n36665;
  assign n36667 = n16508 & n35782;
  assign n36668 = n36666 & ~n36667;
  assign n36669 = pi614 & n16458;
  assign n36670 = pi224 & n16363;
  assign n36671 = n36669 & ~n36670;
  assign n36672 = pi224 & ~n16195;
  assign n36673 = ~n36671 & ~n36672;
  assign n36674 = pi299 & n36673;
  assign n36675 = ~pi614 & n16453;
  assign n36676 = pi224 & ~n36675;
  assign n36677 = n16378 & n36676;
  assign n36678 = pi614 & n16453;
  assign n36679 = ~pi224 & n36678;
  assign n36680 = ~pi299 & ~n36679;
  assign n36681 = ~n36677 & n36680;
  assign n36682 = ~pi39 & ~n36681;
  assign n36683 = ~n36674 & n36682;
  assign n36684 = pi614 & ~n16421;
  assign n36685 = n16263 & ~n35876;
  assign n36686 = ~n36684 & ~n36685;
  assign n36687 = ~pi680 & ~n36686;
  assign n36688 = n16426 & ~n35228;
  assign n36689 = ~n36687 & ~n36688;
  assign n36690 = n6187 & ~n36689;
  assign n36691 = ~n6187 & ~n36686;
  assign n36692 = ~n36690 & ~n36691;
  assign n36693 = ~n6236 & n36692;
  assign n36694 = n16207 & ~n35782;
  assign n36695 = ~n6185 & ~n36694;
  assign n36696 = ~n16233 & ~n36695;
  assign n36697 = ~n6187 & ~n36696;
  assign n36698 = ~pi680 & ~n36696;
  assign n36699 = pi680 & n35782;
  assign n36700 = ~n16236 & ~n36699;
  assign n36701 = ~n36698 & n36700;
  assign n36702 = n6187 & ~n36701;
  assign n36703 = ~n36697 & ~n36702;
  assign n36704 = n6236 & n36703;
  assign n36705 = ~n36693 & ~n36704;
  assign n36706 = pi224 & n36705;
  assign n36707 = pi614 & ~n35547;
  assign n36708 = ~pi224 & n36707;
  assign n36709 = ~n16489 & n36708;
  assign n36710 = pi223 & ~n36709;
  assign n36711 = ~n36706 & n36710;
  assign n36712 = pi614 & ~n35519;
  assign n36713 = n6236 & ~n36712;
  assign n36714 = pi614 & n16809;
  assign n36715 = pi680 & ~n36714;
  assign n36716 = ~pi680 & ~n35783;
  assign n36717 = ~n36715 & ~n36716;
  assign n36718 = n6187 & ~n36717;
  assign n36719 = ~n6187 & ~n35783;
  assign n36720 = ~n36718 & ~n36719;
  assign n36721 = ~n6236 & ~n36720;
  assign n36722 = ~n36713 & ~n36721;
  assign n36723 = n5763 & n36722;
  assign n36724 = pi614 & n16497;
  assign n36725 = ~n16308 & ~n36695;
  assign n36726 = ~n6187 & ~n36725;
  assign n36727 = ~pi680 & ~n36725;
  assign n36728 = ~n16313 & ~n36727;
  assign n36729 = ~n36699 & n36728;
  assign n36730 = n6187 & ~n36729;
  assign n36731 = ~n36726 & ~n36730;
  assign n36732 = n6236 & n36731;
  assign n36733 = ~n16294 & ~n35782;
  assign n36734 = ~n6187 & ~n36733;
  assign n36735 = ~pi680 & ~n36733;
  assign n36736 = n16289 & n36715;
  assign n36737 = ~n36699 & ~n36736;
  assign n36738 = ~n36735 & n36737;
  assign n36739 = n6187 & ~n36738;
  assign n36740 = ~n36734 & ~n36739;
  assign n36741 = ~n6236 & n36740;
  assign n36742 = pi224 & ~n36741;
  assign n36743 = ~n36732 & n36742;
  assign n36744 = ~pi223 & ~n36743;
  assign n36745 = ~n36724 & n36744;
  assign n36746 = ~n36723 & n36745;
  assign n36747 = ~n36711 & ~n36746;
  assign n36748 = ~pi299 & ~n36747;
  assign n36749 = ~n16478 & n36708;
  assign n36750 = n6198 & n36703;
  assign n36751 = ~n6198 & n36692;
  assign n36752 = pi224 & ~n36751;
  assign n36753 = ~n36750 & n36752;
  assign n36754 = ~n36749 & ~n36753;
  assign n36755 = pi215 & ~n36754;
  assign n36756 = n6198 & n36731;
  assign n36757 = ~n6198 & n36740;
  assign n36758 = pi224 & ~n36757;
  assign n36759 = ~n36756 & n36758;
  assign n36760 = n6198 & ~n36712;
  assign n36761 = ~n6198 & ~n36720;
  assign n36762 = ~pi224 & ~n36761;
  assign n36763 = ~n36760 & n36762;
  assign n36764 = ~n2527 & ~n36763;
  assign n36765 = ~n36759 & n36764;
  assign n36766 = pi224 & ~n16207;
  assign n36767 = n2527 & ~n36766;
  assign n36768 = pi614 & n16465;
  assign n36769 = n36767 & ~n36768;
  assign n36770 = ~pi215 & ~n36769;
  assign n36771 = ~n36765 & n36770;
  assign n36772 = pi299 & ~n36771;
  assign n36773 = ~n36755 & n36772;
  assign n36774 = pi39 & ~n36773;
  assign n36775 = ~n36748 & n36774;
  assign n36776 = ~pi38 & ~n36775;
  assign n36777 = ~n36683 & n36776;
  assign n36778 = ~n36668 & ~n36777;
  assign n36779 = n10020 & n36778;
  assign n36780 = ~n36664 & ~n36779;
  assign n36781 = ~n16521 & ~n36780;
  assign n36782 = n16521 & n36662;
  assign n36783 = ~n36781 & ~n36782;
  assign n36784 = ~pi785 & ~n36783;
  assign n36785 = pi609 & n36783;
  assign n36786 = ~pi609 & ~n36662;
  assign n36787 = pi1155 & ~n36786;
  assign n36788 = ~n36785 & n36787;
  assign n36789 = ~pi609 & n36783;
  assign n36790 = pi609 & ~n36662;
  assign n36791 = ~pi1155 & ~n36790;
  assign n36792 = ~n36789 & n36791;
  assign n36793 = ~n36788 & ~n36792;
  assign n36794 = pi785 & ~n36793;
  assign n36795 = ~n36784 & ~n36794;
  assign n36796 = ~pi781 & ~n36795;
  assign n36797 = pi618 & n36795;
  assign n36798 = ~pi618 & ~n36662;
  assign n36799 = pi1154 & ~n36798;
  assign n36800 = ~n36797 & n36799;
  assign n36801 = ~pi618 & n36795;
  assign n36802 = pi618 & ~n36662;
  assign n36803 = ~pi1154 & ~n36802;
  assign n36804 = ~n36801 & n36803;
  assign n36805 = ~n36800 & ~n36804;
  assign n36806 = pi781 & ~n36805;
  assign n36807 = ~n36796 & ~n36806;
  assign n36808 = ~pi789 & ~n36807;
  assign n36809 = pi619 & n36807;
  assign n36810 = ~pi619 & ~n36662;
  assign n36811 = pi1159 & ~n36810;
  assign n36812 = ~n36809 & n36811;
  assign n36813 = ~pi619 & n36807;
  assign n36814 = pi619 & ~n36662;
  assign n36815 = ~pi1159 & ~n36814;
  assign n36816 = ~n36813 & n36815;
  assign n36817 = ~n36812 & ~n36816;
  assign n36818 = pi789 & ~n36817;
  assign n36819 = ~n36808 & ~n36818;
  assign n36820 = ~n17355 & n36819;
  assign n36821 = ~n36663 & ~n36820;
  assign n36822 = ~n19999 & n36821;
  assign n36823 = ~n32843 & ~n36662;
  assign n36824 = pi662 & pi680;
  assign n36825 = n16728 & ~n36824;
  assign n36826 = pi224 & n16710;
  assign n36827 = ~pi224 & ~n16728;
  assign n36828 = ~pi299 & ~n36827;
  assign n36829 = ~n36826 & n36828;
  assign n36830 = ~n36825 & n36829;
  assign n36831 = ~pi39 & ~n36830;
  assign n36832 = n16733 & ~n36824;
  assign n36833 = pi224 & n16716;
  assign n36834 = ~pi224 & ~n16733;
  assign n36835 = pi299 & ~n36834;
  assign n36836 = ~n36833 & n36835;
  assign n36837 = ~n36832 & n36836;
  assign n36838 = n36831 & ~n36837;
  assign n36839 = pi662 & n16630;
  assign n36840 = n36767 & ~n36839;
  assign n36841 = pi662 & n35661;
  assign n36842 = ~n6198 & ~n36841;
  assign n36843 = ~n16607 & n36824;
  assign n36844 = n6198 & ~n36843;
  assign n36845 = ~pi224 & ~n36844;
  assign n36846 = ~n36842 & n36845;
  assign n36847 = pi662 & ~n16657;
  assign n36848 = ~pi662 & ~n16327;
  assign n36849 = ~n36847 & ~n36848;
  assign n36850 = n6198 & n36849;
  assign n36851 = ~n16253 & ~n35655;
  assign n36852 = n16297 & ~n36851;
  assign n36853 = ~n6198 & n36852;
  assign n36854 = pi224 & ~n36853;
  assign n36855 = ~n36850 & n36854;
  assign n36856 = ~n2527 & ~n36855;
  assign n36857 = ~n36846 & n36856;
  assign n36858 = ~n36840 & ~n36857;
  assign n36859 = ~pi215 & ~n36858;
  assign n36860 = ~pi224 & pi662;
  assign n36861 = n16634 & n36860;
  assign n36862 = ~pi662 & ~n16267;
  assign n36863 = pi662 & ~n16679;
  assign n36864 = ~n36862 & ~n36863;
  assign n36865 = ~n6198 & n36864;
  assign n36866 = ~pi662 & ~n16250;
  assign n36867 = pi662 & ~n35682;
  assign n36868 = ~n36866 & ~n36867;
  assign n36869 = n6198 & n36868;
  assign n36870 = pi224 & ~n36869;
  assign n36871 = ~n36865 & n36870;
  assign n36872 = pi215 & ~n36871;
  assign n36873 = ~n36861 & n36872;
  assign n36874 = pi299 & ~n36873;
  assign n36875 = ~n36859 & n36874;
  assign n36876 = ~n6236 & ~n36841;
  assign n36877 = n6236 & ~n36843;
  assign n36878 = ~n36876 & ~n36877;
  assign n36879 = n5763 & n36878;
  assign n36880 = pi662 & n16597;
  assign n36881 = n6236 & n36849;
  assign n36882 = pi224 & ~n36881;
  assign n36883 = ~n6236 & n36852;
  assign n36884 = n36882 & ~n36883;
  assign n36885 = ~pi223 & ~n36884;
  assign n36886 = ~n36880 & n36885;
  assign n36887 = ~n36879 & n36886;
  assign n36888 = n16620 & n36860;
  assign n36889 = ~n6236 & n36864;
  assign n36890 = n6236 & n36868;
  assign n36891 = pi224 & ~n36890;
  assign n36892 = ~n36889 & n36891;
  assign n36893 = ~n36888 & ~n36892;
  assign n36894 = pi223 & n36893;
  assign n36895 = ~pi299 & ~n36894;
  assign n36896 = ~n36887 & n36895;
  assign n36897 = pi39 & ~n36896;
  assign n36898 = ~n36875 & n36897;
  assign n36899 = ~n36838 & ~n36898;
  assign n36900 = ~pi38 & ~n36899;
  assign n36901 = pi662 & n16743;
  assign n36902 = n36666 & ~n36901;
  assign n36903 = ~n36900 & ~n36902;
  assign n36904 = n10020 & n36903;
  assign n36905 = ~n36664 & ~n36904;
  assign n36906 = ~pi778 & ~n36905;
  assign n36907 = pi625 & n36905;
  assign n36908 = ~pi625 & ~n36662;
  assign n36909 = pi1153 & ~n36908;
  assign n36910 = ~n36907 & n36909;
  assign n36911 = ~pi625 & n36905;
  assign n36912 = pi625 & ~n36662;
  assign n36913 = ~pi1153 & ~n36912;
  assign n36914 = ~n36911 & n36913;
  assign n36915 = ~n36910 & ~n36914;
  assign n36916 = pi778 & ~n36915;
  assign n36917 = ~n36906 & ~n36916;
  assign n36918 = ~n16593 & ~n36917;
  assign n36919 = n16593 & n36662;
  assign n36920 = ~n36918 & ~n36919;
  assign n36921 = ~n16589 & ~n36920;
  assign n36922 = n16589 & n36662;
  assign n36923 = ~n36921 & ~n36922;
  assign n36924 = ~n17159 & n36923;
  assign n36925 = ~n17183 & n36924;
  assign n36926 = ~n36823 & ~n36925;
  assign n36927 = pi628 & ~n36926;
  assign n36928 = ~pi628 & ~n36662;
  assign n36929 = n16121 & ~n36928;
  assign n36930 = ~n36927 & n36929;
  assign n36931 = ~pi628 & ~n36926;
  assign n36932 = pi628 & ~n36662;
  assign n36933 = n16122 & ~n36932;
  assign n36934 = ~n36931 & n36933;
  assign n36935 = ~n36930 & ~n36934;
  assign n36936 = ~n36822 & n36935;
  assign n36937 = pi792 & ~n36936;
  assign n36938 = pi618 & n36920;
  assign n36939 = pi609 & n36917;
  assign n36940 = pi625 & n36780;
  assign n36941 = ~pi614 & ~n23427;
  assign n36942 = pi614 & ~n35954;
  assign n36943 = ~n36941 & ~n36942;
  assign n36944 = ~n16204 & n36943;
  assign n36945 = pi616 & ~n36944;
  assign n36946 = pi614 & ~n17022;
  assign n36947 = ~n16788 & ~n36946;
  assign n36948 = ~pi616 & ~n36947;
  assign n36949 = ~n36945 & ~n36948;
  assign n36950 = pi680 & ~n36949;
  assign n36951 = ~n36698 & ~n36950;
  assign n36952 = pi662 & ~n36951;
  assign n36953 = ~pi662 & ~n6186;
  assign n36954 = ~n36696 & n36953;
  assign n36955 = ~n36702 & ~n36954;
  assign n36956 = ~n36952 & n36955;
  assign n36957 = pi224 & n36956;
  assign n36958 = ~n16877 & n35798;
  assign n36959 = ~n35776 & ~n36958;
  assign n36960 = pi680 & ~n36959;
  assign n36961 = pi680 & ~n16907;
  assign n36962 = ~n36768 & ~n36961;
  assign n36963 = ~n36960 & ~n36962;
  assign n36964 = pi662 & ~n36963;
  assign n36965 = ~pi662 & ~n36707;
  assign n36966 = ~n36964 & ~n36965;
  assign n36967 = ~pi224 & ~n36966;
  assign n36968 = n6236 & ~n36967;
  assign n36969 = ~n36957 & n36968;
  assign n36970 = pi614 & ~n35850;
  assign n36971 = n16801 & ~n36970;
  assign n36972 = pi680 & ~n36971;
  assign n36973 = ~n36687 & ~n36972;
  assign n36974 = pi662 & ~n36973;
  assign n36975 = ~n36686 & n36953;
  assign n36976 = ~n36690 & ~n36975;
  assign n36977 = ~n36974 & n36976;
  assign n36978 = pi224 & n36977;
  assign n36979 = ~n16261 & n36707;
  assign n36980 = ~pi662 & ~n36979;
  assign n36981 = pi614 & n35879;
  assign n36982 = ~n16895 & n35798;
  assign n36983 = pi680 & ~n36982;
  assign n36984 = ~n36981 & n36983;
  assign n36985 = ~n16899 & n36984;
  assign n36986 = ~pi680 & ~n16261;
  assign n36987 = n36768 & n36986;
  assign n36988 = pi662 & ~n36987;
  assign n36989 = ~n36985 & n36988;
  assign n36990 = ~n36980 & ~n36989;
  assign n36991 = ~pi224 & ~n36990;
  assign n36992 = ~n6236 & ~n36991;
  assign n36993 = ~n36978 & n36992;
  assign n36994 = pi223 & ~n36993;
  assign n36995 = ~n36969 & n36994;
  assign n36996 = ~n35835 & ~n36768;
  assign n36997 = ~n36960 & ~n36996;
  assign n36998 = pi662 & ~n36997;
  assign n36999 = ~pi662 & ~n36712;
  assign n37000 = ~n36998 & ~n36999;
  assign n37001 = n6236 & ~n37000;
  assign n37002 = pi662 & n35823;
  assign n37003 = ~n36720 & ~n37002;
  assign n37004 = ~n6236 & n37003;
  assign n37005 = ~n37001 & ~n37004;
  assign n37006 = n5763 & n37005;
  assign n37007 = n16877 & n36824;
  assign n37008 = ~n36768 & ~n37007;
  assign n37009 = n2607 & ~n37008;
  assign n37010 = ~n16822 & ~n36946;
  assign n37011 = ~pi616 & ~n37010;
  assign n37012 = ~n36945 & ~n37011;
  assign n37013 = pi680 & ~n37012;
  assign n37014 = ~n36727 & ~n37013;
  assign n37015 = pi662 & ~n37014;
  assign n37016 = ~n36725 & n36953;
  assign n37017 = ~n36730 & ~n37016;
  assign n37018 = ~n37015 & n37017;
  assign n37019 = n6236 & n37018;
  assign n37020 = pi680 & ~n35801;
  assign n37021 = ~n36735 & ~n37020;
  assign n37022 = pi662 & ~n37021;
  assign n37023 = ~n36733 & n36953;
  assign n37024 = ~n36739 & ~n37023;
  assign n37025 = ~n37022 & n37024;
  assign n37026 = ~n6236 & n37025;
  assign n37027 = pi224 & ~n37026;
  assign n37028 = ~n37019 & n37027;
  assign n37029 = ~pi223 & ~n37028;
  assign n37030 = ~n37009 & n37029;
  assign n37031 = ~n37006 & n37030;
  assign n37032 = ~n36995 & ~n37031;
  assign n37033 = ~pi299 & ~n37032;
  assign n37034 = n6198 & ~n36956;
  assign n37035 = ~n6198 & ~n36977;
  assign n37036 = pi224 & ~n37035;
  assign n37037 = ~n37034 & n37036;
  assign n37038 = ~n6198 & n36990;
  assign n37039 = n6198 & n36966;
  assign n37040 = ~pi224 & ~n37039;
  assign n37041 = ~n37038 & n37040;
  assign n37042 = ~n37037 & ~n37041;
  assign n37043 = pi215 & n37042;
  assign n37044 = ~pi224 & n37003;
  assign n37045 = ~n6198 & ~n37044;
  assign n37046 = pi224 & n37025;
  assign n37047 = n37045 & ~n37046;
  assign n37048 = pi224 & n37018;
  assign n37049 = ~pi224 & ~n37000;
  assign n37050 = ~n37048 & ~n37049;
  assign n37051 = n6198 & n37050;
  assign n37052 = ~n2527 & ~n37051;
  assign n37053 = ~n37047 & n37052;
  assign n37054 = ~pi224 & ~n37008;
  assign n37055 = n36767 & ~n37054;
  assign n37056 = n36824 & n36943;
  assign n37057 = ~n35782 & ~n36824;
  assign n37058 = n16212 & n37057;
  assign n37059 = ~n37056 & ~n37058;
  assign n37060 = pi224 & n37059;
  assign n37061 = n37055 & ~n37060;
  assign n37062 = ~pi215 & ~n37061;
  assign n37063 = ~n37053 & n37062;
  assign n37064 = ~n37043 & ~n37063;
  assign n37065 = pi299 & n37064;
  assign n37066 = ~n37033 & ~n37065;
  assign n37067 = pi39 & n37066;
  assign n37068 = n18292 & n36824;
  assign n37069 = ~n36678 & ~n37068;
  assign n37070 = ~pi224 & ~n37069;
  assign n37071 = n18292 & ~n36824;
  assign n37072 = ~n35944 & ~n37071;
  assign n37073 = n36676 & n37072;
  assign n37074 = ~n37070 & ~n37073;
  assign n37075 = ~pi299 & ~n37074;
  assign n37076 = ~pi614 & n16458;
  assign n37077 = ~n35928 & ~n37076;
  assign n37078 = pi224 & ~n37077;
  assign n37079 = ~pi224 & ~n18300;
  assign n37080 = ~n36669 & n37079;
  assign n37081 = ~n37078 & ~n37080;
  assign n37082 = n36824 & ~n37081;
  assign n37083 = n36673 & ~n36824;
  assign n37084 = pi299 & ~n37083;
  assign n37085 = ~n37082 & n37084;
  assign n37086 = ~n37075 & ~n37085;
  assign n37087 = ~pi39 & ~n37086;
  assign n37088 = ~pi38 & ~n37087;
  assign n37089 = ~n37067 & n37088;
  assign n37090 = pi662 & n16814;
  assign n37091 = n16508 & n37090;
  assign n37092 = n36668 & ~n37091;
  assign n37093 = ~n37089 & ~n37092;
  assign n37094 = n10020 & n37093;
  assign n37095 = ~n36664 & ~n37094;
  assign n37096 = ~pi625 & n37095;
  assign n37097 = ~pi1153 & ~n37096;
  assign n37098 = ~n36940 & n37097;
  assign n37099 = ~pi608 & ~n36910;
  assign n37100 = ~n37098 & n37099;
  assign n37101 = ~pi625 & n36780;
  assign n37102 = pi625 & n37095;
  assign n37103 = ~n37101 & ~n37102;
  assign n37104 = pi1153 & n37103;
  assign n37105 = ~n36914 & ~n37104;
  assign n37106 = pi608 & n37105;
  assign n37107 = ~n37100 & ~n37106;
  assign n37108 = pi778 & ~n37107;
  assign n37109 = ~pi778 & n37095;
  assign n37110 = ~n37108 & ~n37109;
  assign n37111 = ~pi609 & ~n37110;
  assign n37112 = ~pi1155 & ~n37111;
  assign n37113 = ~n36939 & n37112;
  assign n37114 = ~pi660 & ~n36788;
  assign n37115 = ~n37113 & n37114;
  assign n37116 = ~pi609 & n36917;
  assign n37117 = pi609 & ~n37110;
  assign n37118 = ~n37116 & ~n37117;
  assign n37119 = pi1155 & n37118;
  assign n37120 = ~n36792 & ~n37119;
  assign n37121 = pi660 & n37120;
  assign n37122 = ~n37115 & ~n37121;
  assign n37123 = pi785 & ~n37122;
  assign n37124 = ~pi785 & ~n37110;
  assign n37125 = ~n37123 & ~n37124;
  assign n37126 = ~pi618 & ~n37125;
  assign n37127 = ~pi1154 & ~n37126;
  assign n37128 = ~n36938 & n37127;
  assign n37129 = ~pi627 & ~n36800;
  assign n37130 = ~n37128 & n37129;
  assign n37131 = ~pi618 & n36920;
  assign n37132 = pi618 & ~n37125;
  assign n37133 = ~n37131 & ~n37132;
  assign n37134 = pi1154 & n37133;
  assign n37135 = ~n36804 & ~n37134;
  assign n37136 = pi627 & n37135;
  assign n37137 = ~n37130 & ~n37136;
  assign n37138 = pi781 & ~n37137;
  assign n37139 = ~pi781 & ~n37125;
  assign n37140 = ~n37138 & ~n37139;
  assign n37141 = ~pi789 & n37140;
  assign n37142 = ~pi619 & ~n37140;
  assign n37143 = pi619 & n36923;
  assign n37144 = ~pi1159 & ~n37143;
  assign n37145 = ~n37142 & n37144;
  assign n37146 = ~pi648 & ~n37145;
  assign n37147 = ~n36812 & n37146;
  assign n37148 = ~pi619 & n36923;
  assign n37149 = pi619 & ~n37140;
  assign n37150 = ~n37148 & ~n37149;
  assign n37151 = pi1159 & n37150;
  assign n37152 = ~n36816 & ~n37151;
  assign n37153 = pi648 & n37152;
  assign n37154 = ~n37147 & ~n37153;
  assign n37155 = pi789 & n37154;
  assign n37156 = ~n37141 & ~n37155;
  assign n37157 = n17356 & n37156;
  assign n37158 = n17159 & ~n36662;
  assign n37159 = ~n36924 & ~n37158;
  assign n37160 = n17350 & ~n37159;
  assign n37161 = pi626 & ~n36819;
  assign n37162 = ~pi626 & n36662;
  assign n37163 = n17180 & ~n37162;
  assign n37164 = ~n37161 & n37163;
  assign n37165 = ~n37160 & ~n37164;
  assign n37166 = ~pi626 & ~n36819;
  assign n37167 = pi626 & n36662;
  assign n37168 = n17181 & ~n37167;
  assign n37169 = ~n37166 & n37168;
  assign n37170 = n37165 & ~n37169;
  assign n37171 = pi788 & ~n37170;
  assign n37172 = n19788 & ~n37171;
  assign n37173 = ~n37157 & n37172;
  assign n37174 = ~n36937 & ~n37173;
  assign n37175 = n19637 & ~n37174;
  assign n37176 = ~n18744 & ~n36926;
  assign n37177 = n17451 & ~n36662;
  assign n37178 = ~n37176 & ~n37177;
  assign n37179 = pi647 & ~n37178;
  assign n37180 = ~pi647 & ~n36662;
  assign n37181 = pi1157 & ~n37180;
  assign n37182 = ~n37179 & n37181;
  assign n37183 = ~pi630 & n37182;
  assign n37184 = ~n16124 & n36821;
  assign n37185 = n16124 & n36662;
  assign n37186 = ~n37184 & ~n37185;
  assign n37187 = ~n19987 & ~n37186;
  assign n37188 = ~pi647 & ~n37178;
  assign n37189 = pi647 & ~n36662;
  assign n37190 = ~pi1157 & ~n37189;
  assign n37191 = ~n37188 & n37190;
  assign n37192 = pi630 & n37191;
  assign n37193 = ~n37187 & ~n37192;
  assign n37194 = ~n37183 & n37193;
  assign n37195 = pi787 & ~n37194;
  assign n37196 = ~n37175 & ~n37195;
  assign n37197 = pi644 & n37196;
  assign n37198 = ~pi787 & n37178;
  assign n37199 = ~n37182 & ~n37191;
  assign n37200 = pi787 & ~n37199;
  assign n37201 = ~n37198 & ~n37200;
  assign n37202 = ~pi644 & n37201;
  assign n37203 = pi715 & ~n37202;
  assign n37204 = ~n37197 & n37203;
  assign n37205 = n17247 & ~n36662;
  assign n37206 = ~n17247 & n37186;
  assign n37207 = ~n37205 & ~n37206;
  assign n37208 = pi644 & ~n37207;
  assign n37209 = ~pi644 & ~n36662;
  assign n37210 = ~pi715 & ~n37209;
  assign n37211 = ~n37208 & n37210;
  assign n37212 = pi1160 & ~n37211;
  assign n37213 = ~n37204 & n37212;
  assign n37214 = pi644 & ~n36662;
  assign n37215 = ~pi644 & ~n37207;
  assign n37216 = pi715 & ~n37215;
  assign n37217 = ~n37214 & n37216;
  assign n37218 = pi644 & n37201;
  assign n37219 = ~pi644 & n37196;
  assign n37220 = ~pi715 & ~n37219;
  assign n37221 = ~n37218 & n37220;
  assign n37222 = ~pi1160 & ~n37221;
  assign n37223 = ~n37217 & n37222;
  assign n37224 = ~n37213 & ~n37223;
  assign n37225 = pi790 & ~n37224;
  assign n37226 = ~pi790 & n37196;
  assign n37227 = ~n37225 & ~n37226;
  assign n37228 = ~po1038 & ~n37227;
  assign n37229 = ~pi224 & po1038;
  assign po381 = ~n37228 & ~n37229;
  assign n37231 = n2553 & n2615;
  assign n37232 = n3314 & n37231;
  assign n37233 = pi62 & n37232;
  assign n37234 = ~pi54 & pi74;
  assign n37235 = n2535 & n37231;
  assign n37236 = ~pi92 & n37235;
  assign n37237 = n37234 & n37236;
  assign n37238 = pi54 & ~n37236;
  assign n37239 = pi92 & n37235;
  assign n37240 = ~n6106 & ~n6166;
  assign n37241 = ~pi137 & ~n37240;
  assign n37242 = n7252 & ~n37241;
  assign n37243 = pi75 & ~n37242;
  assign n37244 = n6099 & ~n37241;
  assign n37245 = pi38 & ~pi137;
  assign n37246 = pi39 & n2553;
  assign n37247 = ~n2895 & ~n11201;
  assign n37248 = n3065 & n37247;
  assign n37249 = n2740 & ~n37248;
  assign n37250 = n2738 & ~n37249;
  assign n37251 = ~n2923 & ~n37250;
  assign n37252 = ~pi95 & ~n37251;
  assign n37253 = ~n2907 & ~n37252;
  assign n37254 = pi137 & ~n37253;
  assign n37255 = n2968 & ~n11202;
  assign n37256 = n2928 & ~n37255;
  assign n37257 = pi1093 & ~n37256;
  assign n37258 = n2928 & n7447;
  assign n37259 = n2686 & ~n7406;
  assign n37260 = ~n2724 & n37259;
  assign n37261 = ~pi32 & ~n37260;
  assign n37262 = n37258 & ~n37261;
  assign n37263 = ~pi1093 & ~n37262;
  assign n37264 = ~n7447 & n37256;
  assign n37265 = n11200 & n37259;
  assign n37266 = n37258 & n37265;
  assign n37267 = ~n37264 & ~n37266;
  assign n37268 = n37263 & n37267;
  assign n37269 = ~n37257 & ~n37268;
  assign n37270 = n11401 & ~n37269;
  assign n37271 = n2995 & ~n7447;
  assign n37272 = n37263 & ~n37271;
  assign n37273 = ~n2948 & n37259;
  assign n37274 = ~pi32 & ~n37273;
  assign n37275 = n37258 & ~n37274;
  assign n37276 = ~n37271 & ~n37275;
  assign n37277 = pi1093 & n37276;
  assign n37278 = ~n37272 & ~n37277;
  assign n37279 = n11381 & ~n37278;
  assign n37280 = n37267 & n37279;
  assign n37281 = ~n37270 & ~n37280;
  assign n37282 = ~n37254 & n37281;
  assign n37283 = pi332 & ~n37282;
  assign n37284 = ~n2907 & ~n2925;
  assign n37285 = pi137 & ~n37284;
  assign n37286 = pi1093 & ~n2995;
  assign n37287 = ~n37272 & ~n37286;
  assign n37288 = n11401 & ~n37287;
  assign n37289 = ~n37279 & ~n37288;
  assign n37290 = ~n37285 & n37289;
  assign n37291 = ~pi332 & ~n37290;
  assign n37292 = ~n37283 & ~n37291;
  assign n37293 = ~n2628 & n37292;
  assign n37294 = ~pi137 & ~n37256;
  assign n37295 = ~n37254 & ~n37294;
  assign n37296 = pi332 & ~n37295;
  assign n37297 = ~n2996 & ~n37285;
  assign n37298 = ~pi332 & ~n37297;
  assign n37299 = ~n37296 & ~n37298;
  assign n37300 = n2628 & n37299;
  assign n37301 = ~pi210 & ~n37300;
  assign n37302 = ~n37293 & n37301;
  assign n37303 = ~n2906 & ~n2907;
  assign n37304 = pi137 & ~n37303;
  assign n37305 = ~n2970 & ~n37304;
  assign n37306 = ~pi332 & ~n37305;
  assign n37307 = ~n2702 & ~n37250;
  assign n37308 = ~pi95 & ~n37307;
  assign n37309 = n3221 & ~n37308;
  assign n37310 = pi332 & ~n37309;
  assign n37311 = ~pi137 & n2703;
  assign n37312 = ~n37255 & n37311;
  assign n37313 = n37310 & ~n37312;
  assign n37314 = ~n37306 & ~n37313;
  assign n37315 = pi210 & ~n37314;
  assign n37316 = pi299 & ~n37315;
  assign n37317 = ~n37302 & n37316;
  assign n37318 = n6498 & n37299;
  assign n37319 = ~n6498 & n37292;
  assign n37320 = ~pi198 & ~n37319;
  assign n37321 = ~n37318 & n37320;
  assign n37322 = pi198 & ~n37314;
  assign n37323 = ~pi299 & ~n37322;
  assign n37324 = ~n37321 & n37323;
  assign n37325 = ~n37317 & ~n37324;
  assign n37326 = ~pi39 & ~n37325;
  assign n37327 = ~pi38 & ~n37326;
  assign n37328 = ~n37246 & n37327;
  assign n37329 = ~n37245 & ~n37328;
  assign n37330 = n6134 & n37329;
  assign n37331 = ~n37244 & ~n37330;
  assign n37332 = ~pi87 & ~n37331;
  assign n37333 = pi87 & n37231;
  assign n37334 = ~pi75 & ~n37333;
  assign n37335 = ~n37332 & n37334;
  assign n37336 = ~pi92 & ~n37335;
  assign n37337 = ~n37243 & n37336;
  assign n37338 = ~pi54 & ~n37337;
  assign n37339 = ~n37239 & n37338;
  assign n37340 = ~pi74 & ~n37339;
  assign n37341 = ~n37238 & n37340;
  assign n37342 = ~pi55 & ~n37341;
  assign n37343 = ~n37237 & n37342;
  assign n37344 = ~pi56 & ~n7250;
  assign n37345 = ~n37343 & n37344;
  assign n37346 = pi56 & n2538;
  assign n37347 = n37231 & n37346;
  assign n37348 = ~n37345 & ~n37347;
  assign n37349 = ~pi62 & ~n37348;
  assign n37350 = ~n37233 & ~n37349;
  assign n37351 = n3327 & n37350;
  assign n37352 = ~pi62 & n37232;
  assign n37353 = ~n3327 & ~n37352;
  assign n37354 = ~n6084 & ~n37353;
  assign po382 = ~n37351 & n37354;
  assign n37356 = pi228 & pi231;
  assign n37357 = pi55 & ~n37356;
  assign n37358 = pi54 & ~n37356;
  assign n37359 = pi87 & ~n37356;
  assign n37360 = ~n7320 & n37359;
  assign n37361 = ~n7310 & ~n37356;
  assign n37362 = pi100 & ~n37361;
  assign n37363 = ~n2718 & ~n3060;
  assign n37364 = ~pi70 & ~n37363;
  assign n37365 = ~pi51 & ~n37364;
  assign n37366 = n2743 & ~n37365;
  assign n37367 = n3065 & ~n37366;
  assign n37368 = n2740 & ~n37367;
  assign n37369 = n2738 & ~n37368;
  assign n37370 = ~n6170 & ~n37369;
  assign n37371 = ~pi95 & ~n37370;
  assign n37372 = n2971 & ~n37371;
  assign n37373 = ~pi39 & ~n37372;
  assign n37374 = ~pi38 & ~n3366;
  assign n37375 = ~n37373 & n37374;
  assign n37376 = ~pi228 & n37375;
  assign n37377 = ~n37356 & ~n37376;
  assign n37378 = ~pi100 & ~n37377;
  assign n37379 = ~pi87 & ~n37378;
  assign n37380 = ~n37362 & n37379;
  assign n37381 = ~pi75 & ~n37380;
  assign n37382 = ~n37360 & n37381;
  assign n37383 = ~n7311 & ~n37356;
  assign n37384 = pi75 & ~n37383;
  assign n37385 = ~pi92 & ~n37384;
  assign n37386 = ~n37382 & n37385;
  assign n37387 = ~n7316 & ~n37356;
  assign n37388 = pi92 & n37387;
  assign n37389 = ~n37386 & ~n37388;
  assign n37390 = ~pi54 & ~n37389;
  assign n37391 = ~pi74 & ~n37390;
  assign n37392 = ~n37358 & n37391;
  assign n37393 = ~n6525 & ~n37356;
  assign n37394 = ~n37383 & ~n37393;
  assign n37395 = pi74 & n37394;
  assign n37396 = ~pi55 & ~n37395;
  assign n37397 = ~n37392 & n37396;
  assign n37398 = ~pi56 & ~n37397;
  assign n37399 = ~n37357 & n37398;
  assign n37400 = ~n7348 & ~n37356;
  assign n37401 = pi56 & ~n37400;
  assign n37402 = ~pi62 & ~n37401;
  assign n37403 = ~n37399 & n37402;
  assign n37404 = ~n7306 & ~n37356;
  assign n37405 = pi62 & n37404;
  assign n37406 = ~n37403 & ~n37405;
  assign n37407 = n3327 & ~n37406;
  assign n37408 = ~n3327 & ~n37356;
  assign po383 = ~n37407 & ~n37408;
  assign n37410 = n2698 & ~n6355;
  assign n37411 = ~pi91 & ~n2754;
  assign n37412 = ~n6120 & n10817;
  assign n37413 = n2725 & n10827;
  assign n37414 = n10825 & n37413;
  assign n37415 = ~n37412 & ~n37414;
  assign n37416 = n37411 & n37415;
  assign n37417 = n37410 & ~n37416;
  assign n37418 = ~pi72 & ~n37417;
  assign n37419 = n6367 & ~n37418;
  assign n37420 = n6208 & ~n37419;
  assign n37421 = n6367 & ~n12799;
  assign n37422 = n12774 & n37421;
  assign n37423 = ~n6447 & ~n37422;
  assign n37424 = pi1093 & ~n37423;
  assign n37425 = n37410 & ~n37411;
  assign n37426 = ~pi72 & ~n37425;
  assign n37427 = n10817 & n37410;
  assign n37428 = ~n7368 & n37427;
  assign n37429 = ~n8751 & ~n37428;
  assign n37430 = n37426 & n37429;
  assign n37431 = n6367 & ~n37430;
  assign n37432 = ~n37424 & ~n37431;
  assign n37433 = n37426 & ~n37427;
  assign n37434 = n6367 & ~n37433;
  assign n37435 = n6211 & ~n37434;
  assign n37436 = ~n37432 & ~n37435;
  assign n37437 = ~n37420 & n37436;
  assign n37438 = ~pi39 & ~n37437;
  assign po384 = ~n11255 | n37438;
  assign n37440 = ~pi39 & pi228;
  assign n37441 = ~n11206 & ~n11210;
  assign n37442 = pi39 & ~n37441;
  assign n37443 = n6455 & n37442;
  assign n37444 = ~n6210 & ~n8752;
  assign n37445 = n2731 & ~n37444;
  assign n37446 = ~n11276 & n37445;
  assign n37447 = n10016 & n37446;
  assign n37448 = ~n37443 & ~n37447;
  assign n37449 = n10024 & ~n37448;
  assign po385 = n37440 | n37449;
  assign n37451 = ~n6133 & n10021;
  assign n37452 = pi824 & ~n16181;
  assign n37453 = pi829 & pi1091;
  assign n37454 = n16186 & n37453;
  assign n37455 = ~pi824 & ~n37454;
  assign n37456 = ~n6451 & ~n37455;
  assign n37457 = ~n37452 & n37456;
  assign n37458 = ~n16148 & ~n37457;
  assign n37459 = ~n6166 & ~n6451;
  assign n37460 = n37453 & n37455;
  assign n37461 = ~n37452 & ~n37460;
  assign n37462 = ~n6451 & ~n37461;
  assign n37463 = n6120 & n37462;
  assign n37464 = ~n37459 & ~n37463;
  assign n37465 = ~n37458 & n37464;
  assign n37466 = ~n7368 & n16148;
  assign n37467 = ~n16165 & ~n37466;
  assign n37468 = n37459 & ~n37467;
  assign n37469 = pi1093 & ~n37468;
  assign n37470 = ~n37465 & n37469;
  assign n37471 = ~n6122 & n16148;
  assign n37472 = n16136 & ~n16138;
  assign n37473 = n2509 & n37472;
  assign n37474 = ~pi40 & ~n37473;
  assign n37475 = n10112 & ~n37474;
  assign n37476 = pi252 & ~n37475;
  assign n37477 = ~n16135 & ~n37476;
  assign n37478 = n6122 & n37477;
  assign n37479 = ~pi1093 & ~n37478;
  assign n37480 = ~n37471 & n37479;
  assign n37481 = ~pi39 & ~n37480;
  assign n37482 = ~n37470 & n37481;
  assign n37483 = ~n6121 & n7431;
  assign n37484 = n16203 & ~n37483;
  assign n37485 = n16273 & n37483;
  assign n37486 = pi1091 & ~n37485;
  assign n37487 = ~n37484 & n37486;
  assign n37488 = ~n6443 & n16203;
  assign n37489 = n6443 & n16273;
  assign n37490 = ~pi1091 & ~n37489;
  assign n37491 = ~n37488 & n37490;
  assign n37492 = ~n37487 & ~n37491;
  assign n37493 = ~pi120 & ~n37492;
  assign n37494 = ~n16205 & ~n37493;
  assign n37495 = ~n6215 & n37494;
  assign n37496 = ~n34901 & ~n37495;
  assign n37497 = ~n6236 & n37496;
  assign n37498 = ~n6191 & n16206;
  assign n37499 = n6191 & n37494;
  assign n37500 = ~n37498 & ~n37499;
  assign n37501 = n6236 & n37500;
  assign n37502 = ~n2607 & ~n37501;
  assign n37503 = ~n37497 & n37502;
  assign n37504 = ~pi223 & ~n37503;
  assign n37505 = ~n16664 & n37504;
  assign n37506 = pi120 & n6213;
  assign n37507 = n16206 & ~n37506;
  assign n37508 = ~n34901 & ~n37507;
  assign n37509 = ~n6236 & ~n37508;
  assign n37510 = pi223 & ~n37509;
  assign n37511 = ~n37498 & ~n37507;
  assign n37512 = n6236 & ~n37511;
  assign n37513 = n37510 & ~n37512;
  assign n37514 = ~pi299 & ~n37513;
  assign n37515 = ~n37505 & n37514;
  assign n37516 = ~n6198 & n37496;
  assign n37517 = n6198 & n37500;
  assign n37518 = ~n2527 & ~n37517;
  assign n37519 = ~n37516 & n37518;
  assign n37520 = ~pi215 & ~n37519;
  assign n37521 = ~n16965 & n37520;
  assign n37522 = ~n6198 & ~n37508;
  assign n37523 = pi215 & ~n37522;
  assign n37524 = n6198 & ~n37511;
  assign n37525 = n37523 & ~n37524;
  assign n37526 = pi299 & ~n37525;
  assign n37527 = ~n37521 & n37526;
  assign n37528 = ~n37515 & ~n37527;
  assign n37529 = pi39 & ~n37528;
  assign n37530 = ~pi38 & ~n37529;
  assign n37531 = ~n37482 & n37530;
  assign po387 = n37451 & ~n37531;
  assign n37533 = ~pi81 & ~n2857;
  assign n37534 = n6329 & ~n37533;
  assign n37535 = n2463 & ~n37534;
  assign n37536 = n2865 & ~n37535;
  assign n37537 = n2776 & ~n37536;
  assign n37538 = n2869 & ~n37537;
  assign n37539 = n2705 & ~n37538;
  assign n37540 = ~n2708 & ~n37539;
  assign n37541 = ~pi86 & ~n37540;
  assign n37542 = n2774 & ~n37541;
  assign n37543 = n2772 & ~n37542;
  assign n37544 = ~n2769 & ~n37543;
  assign n37545 = ~pi108 & ~n37544;
  assign n37546 = n2768 & ~n37545;
  assign n37547 = n2881 & ~n37546;
  assign n37548 = ~n2759 & ~n37547;
  assign n37549 = n2758 & ~n37548;
  assign n37550 = n2757 & ~n37549;
  assign n37551 = n2750 & ~n37550;
  assign n37552 = n3045 & ~n37551;
  assign n37553 = n2519 & ~n37552;
  assign n37554 = n15148 & ~n37553;
  assign n37555 = ~pi70 & ~n37554;
  assign n37556 = ~n3062 & ~n37555;
  assign n37557 = ~pi51 & ~n37556;
  assign n37558 = n2743 & ~n37557;
  assign n37559 = n3065 & ~n37558;
  assign n37560 = n2740 & ~n37559;
  assign n37561 = ~pi1082 & n2737;
  assign n37562 = ~pi32 & ~n37561;
  assign n37563 = ~n37560 & n37562;
  assign n37564 = ~n3376 & ~n37563;
  assign n37565 = ~pi95 & ~n37564;
  assign n37566 = ~n2907 & ~n37565;
  assign n37567 = ~pi39 & ~n37566;
  assign n37568 = ~n7263 & ~n11205;
  assign po950 = ~n6120 | ~n6212;
  assign n37570 = ~n37568 & ~po950;
  assign n37571 = n6441 & n37570;
  assign n37572 = n6179 & ~n37571;
  assign n37573 = n11152 & n37572;
  assign n37574 = ~n3366 & ~n37573;
  assign n37575 = ~n37567 & n37574;
  assign n37576 = ~pi38 & ~n37575;
  assign n37577 = n6134 & ~n37576;
  assign n37578 = ~pi87 & ~n6099;
  assign n37579 = ~n37577 & n37578;
  assign n37580 = ~n6095 & ~n37579;
  assign n37581 = n2573 & ~n37580;
  assign n37582 = n7259 & ~n37581;
  assign n37583 = ~pi54 & ~n37582;
  assign n37584 = ~n7295 & ~n37583;
  assign n37585 = n6262 & ~n37584;
  assign n37586 = n7251 & ~n37585;
  assign n37587 = ~pi56 & ~n37586;
  assign n37588 = ~n6264 & ~n37587;
  assign n37589 = ~pi62 & ~n37588;
  assign n37590 = ~n6268 & ~n37589;
  assign n37591 = n3327 & ~n37590;
  assign po389 = n6087 & ~n37591;
  assign n37593 = ~pi230 & ~pi233;
  assign n37594 = ~pi212 & pi214;
  assign n37595 = ~pi211 & pi1157;
  assign n37596 = pi211 & pi1156;
  assign n37597 = ~n37595 & ~n37596;
  assign n37598 = n37594 & ~n37597;
  assign n37599 = ~pi211 & pi1156;
  assign n37600 = pi211 & pi1155;
  assign n37601 = ~n37599 & ~n37600;
  assign n37602 = ~pi214 & n37601;
  assign n37603 = ~pi211 & pi1155;
  assign n37604 = pi211 & pi1154;
  assign n37605 = ~n37603 & ~n37604;
  assign n37606 = pi214 & n37605;
  assign n37607 = pi212 & ~n37606;
  assign n37608 = ~n37602 & n37607;
  assign n37609 = ~n37598 & ~n37608;
  assign n37610 = ~pi219 & n37609;
  assign n37611 = ~pi211 & pi1153;
  assign n37612 = n10468 & ~n37611;
  assign n37613 = ~pi211 & pi1154;
  assign n37614 = ~pi214 & ~n37613;
  assign n37615 = ~pi211 & pi214;
  assign n37616 = pi1155 & n37615;
  assign n37617 = ~pi212 & ~n37616;
  assign n37618 = ~n37614 & ~n37617;
  assign n37619 = ~n37612 & n37618;
  assign n37620 = pi219 & ~n37619;
  assign n37621 = ~n37610 & ~n37620;
  assign n37622 = po1038 & n37621;
  assign n37623 = ~pi213 & ~n37622;
  assign n37624 = pi199 & pi1142;
  assign n37625 = ~pi200 & ~n37624;
  assign n37626 = ~pi199 & pi1144;
  assign n37627 = n37625 & ~n37626;
  assign n37628 = ~pi199 & pi1143;
  assign n37629 = pi200 & ~n37628;
  assign n37630 = ~n37627 & ~n37629;
  assign n37631 = ~pi299 & ~n37630;
  assign n37632 = ~pi207 & ~n37631;
  assign n37633 = pi207 & ~pi299;
  assign n37634 = n37625 & ~n37628;
  assign n37635 = ~pi199 & pi1142;
  assign n37636 = pi200 & ~n37635;
  assign n37637 = ~n37634 & ~n37636;
  assign n37638 = n37633 & n37637;
  assign n37639 = ~n37632 & ~n37638;
  assign n37640 = pi208 & ~n37639;
  assign n37641 = pi207 & ~pi208;
  assign n37642 = n37630 & n37641;
  assign n37643 = ~n37640 & ~n37642;
  assign n37644 = ~pi299 & ~n37643;
  assign n37645 = ~pi219 & pi299;
  assign n37646 = ~n37609 & n37645;
  assign n37647 = pi299 & pi1155;
  assign n37648 = n37594 & n37647;
  assign n37649 = pi299 & pi1154;
  assign n37650 = ~pi214 & ~n37649;
  assign n37651 = pi299 & pi1153;
  assign n37652 = pi214 & ~n37651;
  assign n37653 = pi212 & ~n37652;
  assign n37654 = ~n37650 & n37653;
  assign n37655 = ~n37648 & ~n37654;
  assign n37656 = n10522 & ~n37655;
  assign n37657 = ~n37646 & ~n37656;
  assign n37658 = ~n37644 & n37657;
  assign n37659 = ~po1038 & ~n37658;
  assign n37660 = n37623 & ~n37659;
  assign n37661 = ~pi212 & ~pi214;
  assign n37662 = ~pi211 & ~n37661;
  assign n37663 = pi219 & ~n37662;
  assign n37664 = po1038 & ~n37663;
  assign n37665 = pi1142 & ~n10470;
  assign n37666 = pi211 & pi1143;
  assign n37667 = ~pi211 & pi1144;
  assign n37668 = ~n37666 & ~n37667;
  assign n37669 = pi212 & ~pi214;
  assign n37670 = ~n37594 & ~n37669;
  assign n37671 = ~n37668 & ~n37670;
  assign n37672 = ~pi211 & pi1143;
  assign n37673 = n10468 & n37672;
  assign n37674 = ~n37671 & ~n37673;
  assign n37675 = ~pi219 & ~n37674;
  assign n37676 = ~n37665 & ~n37675;
  assign n37677 = n37664 & ~n37676;
  assign n37678 = ~pi214 & ~n37644;
  assign n37679 = pi299 & ~n37668;
  assign n37680 = ~n37644 & ~n37679;
  assign n37681 = ~pi212 & ~n37680;
  assign n37682 = ~n37678 & n37681;
  assign n37683 = pi211 & pi1142;
  assign n37684 = ~n37672 & ~n37683;
  assign n37685 = pi299 & ~n37684;
  assign n37686 = ~n37644 & ~n37685;
  assign n37687 = pi214 & n37686;
  assign n37688 = n37678 & ~n37679;
  assign n37689 = pi212 & ~n37688;
  assign n37690 = ~n37687 & n37689;
  assign n37691 = ~pi219 & ~n37690;
  assign n37692 = ~n37682 & n37691;
  assign n37693 = pi299 & ~n37661;
  assign n37694 = ~pi211 & pi1142;
  assign n37695 = n37693 & n37694;
  assign n37696 = ~n37644 & ~n37695;
  assign n37697 = pi219 & n37696;
  assign n37698 = ~n37692 & ~n37697;
  assign n37699 = ~po1038 & n37698;
  assign n37700 = ~n37677 & ~n37699;
  assign n37701 = pi213 & n37700;
  assign n37702 = pi209 & ~n37701;
  assign n37703 = ~n37660 & n37702;
  assign n37704 = pi211 & pi214;
  assign n37705 = ~pi211 & ~pi214;
  assign n37706 = ~n37704 & ~n37705;
  assign n37707 = pi1155 & ~n11164;
  assign n37708 = pi199 & ~pi1153;
  assign n37709 = pi199 & pi200;
  assign n37710 = ~n10614 & ~n37709;
  assign n37711 = ~pi299 & n37710;
  assign n37712 = ~n37708 & n37711;
  assign n37713 = ~n37707 & ~n37712;
  assign n37714 = pi200 & ~pi299;
  assign n37715 = ~pi1154 & n37714;
  assign n37716 = ~n37713 & ~n37715;
  assign n37717 = pi207 & ~n37716;
  assign n37718 = ~pi199 & pi1155;
  assign n37719 = n37714 & n37718;
  assign n37720 = ~pi1154 & ~n37719;
  assign n37721 = pi200 & ~n37718;
  assign n37722 = n10615 & ~n37721;
  assign n37723 = ~n37720 & n37722;
  assign n37724 = pi200 & ~pi1155;
  assign n37725 = n11156 & ~n37724;
  assign n37726 = pi1156 & n37725;
  assign n37727 = ~n37723 & ~n37726;
  assign n37728 = ~pi207 & ~n37647;
  assign n37729 = n37727 & n37728;
  assign n37730 = ~n37717 & ~n37729;
  assign n37731 = pi208 & n37730;
  assign n37732 = ~pi208 & ~n37728;
  assign n37733 = ~pi200 & pi1155;
  assign n37734 = pi199 & n37733;
  assign n37735 = ~pi299 & n37734;
  assign n37736 = ~pi1156 & ~n37735;
  assign n37737 = ~pi299 & n37736;
  assign n37738 = ~pi299 & ~n37710;
  assign n37739 = ~pi1155 & ~n11156;
  assign n37740 = ~n37738 & ~n37739;
  assign n37741 = ~n37737 & n37740;
  assign n37742 = n37732 & n37741;
  assign n37743 = ~pi208 & pi1157;
  assign n37744 = pi1155 & ~n37714;
  assign n37745 = ~n11156 & ~n37744;
  assign n37746 = pi1156 & ~n37745;
  assign n37747 = pi199 & ~pi200;
  assign n37748 = ~pi299 & ~n37747;
  assign n37749 = ~pi1155 & ~n37748;
  assign n37750 = ~pi1156 & ~n37714;
  assign n37751 = ~n37749 & n37750;
  assign n37752 = ~n37746 & ~n37751;
  assign n37753 = n37743 & ~n37752;
  assign n37754 = ~n37728 & n37753;
  assign n37755 = ~n37742 & ~n37754;
  assign n37756 = ~n37731 & n37755;
  assign n37757 = n37706 & ~n37756;
  assign n37758 = ~pi207 & ~pi299;
  assign n37759 = ~pi208 & ~n37758;
  assign n37760 = ~pi299 & ~n11221;
  assign n37761 = pi1156 & ~n37734;
  assign n37762 = n37760 & n37761;
  assign n37763 = ~n37736 & ~n37762;
  assign n37764 = ~pi299 & ~n37763;
  assign n37765 = n37759 & ~n37764;
  assign n37766 = ~n37736 & n37765;
  assign n37767 = ~pi299 & ~n37709;
  assign n37768 = pi199 & ~pi1155;
  assign n37769 = pi1156 & ~n37768;
  assign n37770 = n37767 & n37769;
  assign n37771 = ~pi200 & ~pi299;
  assign n37772 = ~pi1156 & ~n37768;
  assign n37773 = n37771 & n37772;
  assign n37774 = ~n37770 & ~n37773;
  assign n37775 = pi207 & ~n37774;
  assign n37776 = pi299 & pi1156;
  assign n37777 = ~n37775 & ~n37776;
  assign n37778 = n37743 & ~n37777;
  assign n37779 = pi1153 & ~n37767;
  assign n37780 = pi1154 & ~n37779;
  assign n37781 = n11156 & n37733;
  assign n37782 = ~pi1153 & ~n11156;
  assign n37783 = pi1154 & ~n37782;
  assign n37784 = n37710 & n37783;
  assign n37785 = ~n37781 & ~n37784;
  assign n37786 = n37780 & ~n37785;
  assign n37787 = ~n37708 & n37771;
  assign n37788 = ~pi199 & ~pi1155;
  assign n37789 = ~pi1154 & ~n37788;
  assign n37790 = n37787 & n37789;
  assign n37791 = ~n37786 & ~n37790;
  assign n37792 = pi207 & ~n37791;
  assign n37793 = ~pi1155 & ~n10615;
  assign n37794 = ~n37707 & ~n37793;
  assign n37795 = pi1156 & ~n37794;
  assign n37796 = ~n37723 & ~n37795;
  assign n37797 = ~n37633 & ~n37796;
  assign n37798 = ~n37792 & ~n37797;
  assign n37799 = pi208 & ~n37798;
  assign n37800 = ~n37778 & ~n37799;
  assign n37801 = ~n37766 & n37800;
  assign n37802 = n37705 & ~n37801;
  assign n37803 = ~n37744 & ~n37793;
  assign n37804 = n11164 & ~n37733;
  assign n37805 = pi1156 & ~n37804;
  assign n37806 = n37803 & ~n37805;
  assign n37807 = pi207 & n37806;
  assign n37808 = n37759 & ~n37807;
  assign n37809 = pi299 & ~pi1154;
  assign n37810 = pi1157 & ~n37809;
  assign n37811 = n37808 & n37810;
  assign n37812 = n37711 & ~n37768;
  assign n37813 = ~n37736 & n37812;
  assign n37814 = pi207 & n37813;
  assign n37815 = ~n37649 & ~n37814;
  assign n37816 = ~pi208 & ~n37815;
  assign n37817 = ~pi1157 & n37816;
  assign n37818 = pi1155 & ~n37738;
  assign n37819 = ~n37749 & ~n37818;
  assign n37820 = pi1154 & ~n37819;
  assign n37821 = n37727 & ~n37820;
  assign n37822 = ~pi207 & ~n37821;
  assign n37823 = ~pi299 & n37713;
  assign n37824 = pi1154 & ~n37823;
  assign n37825 = ~n37790 & ~n37824;
  assign n37826 = pi207 & ~n37825;
  assign n37827 = ~n37822 & ~n37826;
  assign n37828 = pi208 & ~n37827;
  assign n37829 = ~n37817 & ~n37828;
  assign n37830 = ~n37811 & n37829;
  assign n37831 = n37704 & ~n37830;
  assign n37832 = ~n37802 & ~n37831;
  assign n37833 = ~n37757 & n37832;
  assign n37834 = pi212 & ~n37833;
  assign n37835 = ~pi208 & ~n37814;
  assign n37836 = pi207 & n37791;
  assign n37837 = ~n10302 & n37727;
  assign n37838 = ~n37836 & ~n37837;
  assign n37839 = pi208 & ~n37838;
  assign n37840 = ~n37835 & ~n37839;
  assign n37841 = ~pi1157 & ~n37840;
  assign n37842 = ~pi208 & ~n37775;
  assign n37843 = ~n37839 & ~n37842;
  assign n37844 = pi1157 & ~n37843;
  assign n37845 = ~n37841 & ~n37844;
  assign n37846 = ~pi214 & ~n37845;
  assign n37847 = ~pi212 & ~n37846;
  assign n37848 = pi211 & ~n37801;
  assign n37849 = pi1157 & ~n37808;
  assign n37850 = pi299 & ~pi1155;
  assign n37851 = pi1155 & ~n37760;
  assign n37852 = ~n37850 & ~n37851;
  assign n37853 = ~n37795 & n37852;
  assign n37854 = ~n37820 & n37853;
  assign n37855 = ~pi207 & n37854;
  assign n37856 = pi1153 & ~n37748;
  assign n37857 = n37785 & ~n37856;
  assign n37858 = n37633 & n37857;
  assign n37859 = ~n37855 & ~n37858;
  assign n37860 = pi208 & n37859;
  assign n37861 = n37849 & ~n37860;
  assign n37862 = ~pi211 & ~n37861;
  assign n37863 = ~n37841 & n37862;
  assign n37864 = ~n37848 & ~n37863;
  assign n37865 = pi214 & n37864;
  assign n37866 = n37847 & ~n37865;
  assign n37867 = ~pi219 & ~n37866;
  assign n37868 = ~n37834 & n37867;
  assign n37869 = pi211 & ~n37845;
  assign n37870 = n37615 & n37756;
  assign n37871 = n37847 & ~n37870;
  assign n37872 = pi207 & ~n37857;
  assign n37873 = pi299 & ~pi1153;
  assign n37874 = ~pi207 & ~n37873;
  assign n37875 = ~n37854 & n37874;
  assign n37876 = ~n37872 & ~n37875;
  assign n37877 = pi208 & ~n37876;
  assign n37878 = ~pi1157 & ~n37765;
  assign n37879 = ~n37849 & ~n37873;
  assign n37880 = ~n37878 & n37879;
  assign n37881 = ~n37877 & ~n37880;
  assign n37882 = n37615 & n37881;
  assign n37883 = n37705 & n37830;
  assign n37884 = pi212 & ~n37883;
  assign n37885 = ~n37882 & n37884;
  assign n37886 = ~n37871 & ~n37885;
  assign n37887 = ~n37869 & ~n37886;
  assign n37888 = pi219 & ~n37887;
  assign n37889 = ~po1038 & ~n37888;
  assign n37890 = ~n37868 & n37889;
  assign n37891 = n37623 & ~n37890;
  assign n37892 = ~pi209 & ~n37891;
  assign n37893 = pi299 & pi1144;
  assign n37894 = ~pi299 & ~n37796;
  assign n37895 = ~n37893 & ~n37894;
  assign n37896 = ~pi207 & n37895;
  assign n37897 = n37836 & ~n37893;
  assign n37898 = pi208 & ~n37897;
  assign n37899 = ~n37896 & n37898;
  assign n37900 = pi299 & ~pi1144;
  assign n37901 = ~pi1157 & n37765;
  assign n37902 = ~n37900 & n37901;
  assign n37903 = ~n37770 & n37803;
  assign n37904 = ~n37758 & ~n37900;
  assign n37905 = ~n37903 & n37904;
  assign n37906 = n37743 & n37905;
  assign n37907 = ~n37902 & ~n37906;
  assign n37908 = ~n37899 & n37907;
  assign n37909 = ~pi211 & ~n37908;
  assign n37910 = ~n37670 & ~n37909;
  assign n37911 = ~pi211 & n37910;
  assign n37912 = pi299 & pi1143;
  assign n37913 = ~n37894 & ~n37912;
  assign n37914 = ~pi207 & n37913;
  assign n37915 = n37836 & ~n37912;
  assign n37916 = pi208 & ~n37915;
  assign n37917 = ~n37914 & n37916;
  assign n37918 = ~pi211 & n10468;
  assign n37919 = ~n37910 & ~n37918;
  assign n37920 = pi299 & ~pi1143;
  assign n37921 = n37901 & ~n37920;
  assign n37922 = ~n37758 & ~n37920;
  assign n37923 = ~n37903 & n37922;
  assign n37924 = n37743 & n37923;
  assign n37925 = ~n37921 & ~n37924;
  assign n37926 = ~n37919 & n37925;
  assign n37927 = ~n37917 & n37926;
  assign n37928 = ~n37911 & ~n37927;
  assign n37929 = ~pi219 & ~n37928;
  assign n37930 = ~pi219 & ~n37661;
  assign n37931 = ~n37662 & ~n37930;
  assign n37932 = ~n37845 & n37931;
  assign n37933 = ~n37929 & ~n37932;
  assign n37934 = pi299 & ~pi1142;
  assign n37935 = ~n37878 & ~n37934;
  assign n37936 = ~n37849 & n37935;
  assign n37937 = pi299 & pi1142;
  assign n37938 = ~pi299 & n37716;
  assign n37939 = ~n37937 & ~n37938;
  assign n37940 = pi207 & n37939;
  assign n37941 = ~pi207 & ~n37937;
  assign n37942 = ~n37894 & n37941;
  assign n37943 = pi208 & ~n37942;
  assign n37944 = ~n37940 & n37943;
  assign n37945 = ~n10470 & ~n37944;
  assign n37946 = ~n37936 & n37945;
  assign n37947 = ~n37931 & n37946;
  assign n37948 = ~po1038 & ~n37947;
  assign n37949 = n37933 & n37948;
  assign n37950 = ~n37677 & ~n37949;
  assign n37951 = pi213 & n37950;
  assign n37952 = n37892 & ~n37951;
  assign n37953 = ~n37703 & ~n37952;
  assign n37954 = pi230 & ~n37953;
  assign po390 = n37593 | n37954;
  assign n37956 = ~pi207 & ~pi208;
  assign n37957 = ~n10302 & ~n37956;
  assign n37958 = ~pi1154 & ~n37781;
  assign n37959 = ~pi1155 & n10614;
  assign n37960 = ~n37709 & ~n37959;
  assign n37961 = ~n37958 & n37960;
  assign n37962 = n37633 & n37961;
  assign n37963 = ~n37957 & ~n37962;
  assign n37964 = ~n37837 & ~n37963;
  assign n37965 = ~n37662 & n37964;
  assign n37966 = pi219 & ~n37965;
  assign n37967 = ~pi207 & n37649;
  assign n37968 = pi207 & ~n37821;
  assign n37969 = ~n37967 & ~n37968;
  assign n37970 = ~pi208 & ~n37969;
  assign n37971 = ~pi299 & n37709;
  assign n37972 = pi207 & ~n37971;
  assign n37973 = ~pi299 & ~n37721;
  assign n37974 = pi1154 & ~n37973;
  assign n37975 = ~n37961 & ~n37974;
  assign n37976 = n37972 & ~n37975;
  assign n37977 = ~n37822 & ~n37976;
  assign n37978 = pi208 & ~n37977;
  assign n37979 = ~n37970 & ~n37978;
  assign n37980 = ~pi211 & ~n37979;
  assign n37981 = ~n37661 & n37980;
  assign n37982 = n37966 & ~n37981;
  assign n37983 = ~n37797 & ~n37962;
  assign n37984 = pi208 & ~n37983;
  assign n37985 = n37759 & ~n37796;
  assign n37986 = ~n37984 & ~n37985;
  assign n37987 = ~pi211 & ~n37986;
  assign n37988 = ~n37647 & ~n37964;
  assign n37989 = pi211 & ~n37988;
  assign n37990 = ~n37987 & ~n37989;
  assign n37991 = ~pi214 & n37990;
  assign n37992 = ~pi211 & ~n37988;
  assign n37993 = pi211 & ~n37979;
  assign n37994 = pi214 & ~n37993;
  assign n37995 = ~n37992 & n37994;
  assign n37996 = ~n37991 & ~n37995;
  assign n37997 = pi212 & n37996;
  assign n37998 = ~pi214 & ~n37964;
  assign n37999 = ~pi212 & ~n37998;
  assign n38000 = pi214 & n37990;
  assign n38001 = n37999 & ~n38000;
  assign n38002 = ~pi219 & ~n38001;
  assign n38003 = ~n37997 & n38002;
  assign n38004 = n35059 & ~n38003;
  assign n38005 = ~n37982 & n38004;
  assign n38006 = pi211 & pi1153;
  assign n38007 = ~n37613 & ~n38006;
  assign n38008 = ~n10468 & n38007;
  assign n38009 = n37930 & ~n38008;
  assign n38010 = ~n37612 & n38009;
  assign n38011 = po1038 & n38010;
  assign n38012 = ~pi1152 & ~n38011;
  assign n38013 = pi207 & n37853;
  assign n38014 = ~n37820 & n38013;
  assign n38015 = n37759 & ~n38014;
  assign n38016 = n37633 & ~n37961;
  assign n38017 = ~n37855 & ~n38016;
  assign n38018 = pi208 & n38017;
  assign n38019 = ~n38015 & ~n38018;
  assign n38020 = ~n37873 & ~n38019;
  assign n38021 = pi211 & n38020;
  assign n38022 = ~n37980 & ~n38021;
  assign n38023 = pi214 & n38022;
  assign n38024 = n37999 & ~n38023;
  assign n38025 = ~pi219 & ~n38024;
  assign n38026 = ~pi214 & ~n38022;
  assign n38027 = ~pi211 & ~n38020;
  assign n38028 = pi214 & ~n38027;
  assign n38029 = pi211 & ~n37964;
  assign n38030 = n38028 & ~n38029;
  assign n38031 = ~n38026 & ~n38030;
  assign n38032 = pi212 & ~n38031;
  assign n38033 = n38025 & ~n38032;
  assign n38034 = pi219 & ~n37964;
  assign n38035 = ~po1038 & ~n38034;
  assign n38036 = ~n38033 & n38035;
  assign n38037 = n38012 & ~n38036;
  assign n38038 = pi1153 & ~n37705;
  assign n38039 = ~n37614 & ~n37615;
  assign n38040 = ~n38038 & ~n38039;
  assign n38041 = pi212 & ~n38040;
  assign n38042 = n37594 & ~n38007;
  assign n38043 = ~pi219 & ~n38042;
  assign n38044 = ~n38041 & n38043;
  assign n38045 = n37664 & ~n38044;
  assign n38046 = pi1152 & ~n38045;
  assign n38047 = ~n38019 & n38028;
  assign n38048 = ~n38026 & ~n38047;
  assign n38049 = pi212 & ~n38048;
  assign n38050 = n38025 & ~n38049;
  assign n38051 = n37662 & ~n38019;
  assign n38052 = n37966 & ~n38051;
  assign n38053 = ~po1038 & ~n38052;
  assign n38054 = ~n38050 & n38053;
  assign n38055 = n38046 & ~n38054;
  assign n38056 = ~pi213 & ~n38055;
  assign n38057 = ~n38037 & n38056;
  assign n38058 = pi209 & ~n38057;
  assign n38059 = ~n38005 & n38058;
  assign n38060 = pi1154 & ~n37714;
  assign n38061 = pi1153 & n11221;
  assign n38062 = ~pi299 & n38061;
  assign n38063 = ~n38060 & ~n38062;
  assign n38064 = n37748 & n38063;
  assign n38065 = n37759 & ~n38064;
  assign n38066 = ~pi200 & ~pi1153;
  assign n38067 = ~pi199 & ~n38066;
  assign n38068 = ~pi299 & ~n38067;
  assign n38069 = ~n37747 & n38068;
  assign n38070 = pi207 & ~n38069;
  assign n38071 = ~pi207 & ~n38064;
  assign n38072 = ~n38070 & ~n38071;
  assign n38073 = pi208 & ~n38072;
  assign n38074 = ~n38065 & ~n38073;
  assign n38075 = ~pi211 & ~n38074;
  assign n38076 = ~pi299 & n10614;
  assign n38077 = ~pi1153 & ~n38076;
  assign n38078 = n37780 & ~n38077;
  assign n38079 = ~pi199 & ~pi1153;
  assign n38080 = n37711 & ~n38079;
  assign n38081 = ~n38078 & ~n38080;
  assign n38082 = ~n10302 & n38081;
  assign n38083 = ~pi1153 & n10614;
  assign n38084 = n37767 & ~n38083;
  assign n38085 = n10302 & ~n38084;
  assign n38086 = ~n37956 & ~n38085;
  assign n38087 = ~n38082 & n38086;
  assign n38088 = pi211 & n38087;
  assign n38089 = ~n38075 & ~n38088;
  assign n38090 = ~n37661 & ~n38089;
  assign n38091 = pi219 & ~n37661;
  assign n38092 = pi219 & ~n38087;
  assign n38093 = ~n38091 & ~n38092;
  assign n38094 = ~n38090 & ~n38093;
  assign n38095 = ~po1038 & ~n38094;
  assign n38096 = ~pi214 & ~n38087;
  assign n38097 = ~pi212 & ~n38096;
  assign n38098 = ~n37649 & ~n38087;
  assign n38099 = ~pi211 & ~n38098;
  assign n38100 = ~pi1153 & ~n37771;
  assign n38101 = ~n37738 & ~n38100;
  assign n38102 = pi1154 & ~n11164;
  assign n38103 = ~n38100 & n38102;
  assign n38104 = ~n38101 & ~n38103;
  assign n38105 = ~pi207 & ~n38104;
  assign n38106 = ~pi1153 & ~n10615;
  assign n38107 = n37972 & ~n38106;
  assign n38108 = ~n38105 & ~n38107;
  assign n38109 = pi208 & ~n38108;
  assign n38110 = n37767 & ~n37956;
  assign n38111 = ~pi299 & ~n38110;
  assign n38112 = ~pi208 & ~n38111;
  assign n38113 = ~n38104 & n38112;
  assign n38114 = ~n38109 & ~n38113;
  assign n38115 = pi211 & ~n38114;
  assign n38116 = ~n38099 & ~n38115;
  assign n38117 = pi214 & n38116;
  assign n38118 = n38097 & ~n38117;
  assign n38119 = ~pi214 & n38116;
  assign n38120 = pi211 & ~n38074;
  assign n38121 = ~pi211 & ~n38114;
  assign n38122 = ~n38120 & ~n38121;
  assign n38123 = pi214 & n38122;
  assign n38124 = ~n38119 & ~n38123;
  assign n38125 = pi212 & n38124;
  assign n38126 = ~pi219 & ~n38125;
  assign n38127 = ~n38118 & n38126;
  assign n38128 = n38095 & ~n38127;
  assign n38129 = n38046 & ~n38128;
  assign n38130 = ~pi1154 & ~n38062;
  assign n38131 = pi200 & ~pi1153;
  assign n38132 = n11156 & ~n38131;
  assign n38133 = ~n38130 & n38132;
  assign n38134 = n37957 & n38133;
  assign n38135 = pi208 & n37633;
  assign n38136 = pi1153 & ~n10615;
  assign n38137 = n38135 & n38136;
  assign n38138 = ~n38134 & ~n38137;
  assign n38139 = pi219 & n38138;
  assign n38140 = ~po1038 & ~n38139;
  assign n38141 = pi1153 & ~n11164;
  assign n38142 = ~n38106 & ~n38141;
  assign n38143 = pi1154 & ~n38142;
  assign n38144 = ~n38062 & ~n38143;
  assign n38145 = ~pi299 & n38144;
  assign n38146 = pi207 & n38145;
  assign n38147 = n37759 & ~n38146;
  assign n38148 = ~pi207 & n38145;
  assign n38149 = pi208 & ~n38148;
  assign n38150 = pi1153 & n38076;
  assign n38151 = n37633 & ~n38150;
  assign n38152 = n38149 & ~n38151;
  assign n38153 = ~n38147 & ~n38152;
  assign n38154 = ~n11164 & ~n38100;
  assign n38155 = ~n38153 & n38154;
  assign n38156 = n37918 & ~n38155;
  assign n38157 = ~n10468 & ~n37661;
  assign n38158 = ~n11164 & ~n37809;
  assign n38159 = ~n38153 & n38158;
  assign n38160 = ~pi211 & ~n38159;
  assign n38161 = pi211 & ~n38155;
  assign n38162 = ~n38160 & ~n38161;
  assign n38163 = n38157 & ~n38162;
  assign n38164 = ~n38156 & ~n38163;
  assign n38165 = ~pi219 & ~n38164;
  assign n38166 = ~n37615 & ~n38157;
  assign n38167 = n38138 & n38166;
  assign n38168 = ~n38165 & ~n38167;
  assign n38169 = n38140 & n38168;
  assign n38170 = n38012 & ~n38169;
  assign n38171 = ~n38129 & ~n38170;
  assign n38172 = ~pi213 & n38171;
  assign n38173 = ~pi1152 & ~po1038;
  assign n38174 = n37661 & ~n38138;
  assign n38175 = pi211 & ~n38159;
  assign n38176 = ~n11164 & ~n37739;
  assign n38177 = ~n38153 & n38176;
  assign n38178 = ~pi211 & ~n38177;
  assign n38179 = n10468 & ~n38178;
  assign n38180 = ~n38175 & n38179;
  assign n38181 = pi211 & ~n38177;
  assign n38182 = ~pi211 & ~n37776;
  assign n38183 = n38138 & n38182;
  assign n38184 = ~n37670 & ~n38183;
  assign n38185 = ~n38181 & n38184;
  assign n38186 = ~n38180 & ~n38185;
  assign n38187 = ~pi219 & ~n38186;
  assign n38188 = pi211 & n38138;
  assign n38189 = ~n38160 & ~n38188;
  assign n38190 = n38091 & n38189;
  assign n38191 = ~n38187 & ~n38190;
  assign n38192 = ~n38174 & n38191;
  assign n38193 = n38173 & ~n38192;
  assign n38194 = ~pi212 & n38096;
  assign n38195 = pi211 & ~n38110;
  assign n38196 = ~n38098 & ~n38195;
  assign n38197 = ~n38194 & n38196;
  assign n38198 = pi219 & n38197;
  assign n38199 = pi211 & ~n38098;
  assign n38200 = ~n37850 & ~n38074;
  assign n38201 = ~pi211 & n38200;
  assign n38202 = n10468 & ~n38201;
  assign n38203 = ~n38199 & n38202;
  assign n38204 = ~n37776 & n38081;
  assign n38205 = ~pi207 & ~n38204;
  assign n38206 = pi299 & ~pi1156;
  assign n38207 = n38070 & ~n38206;
  assign n38208 = pi208 & ~n38207;
  assign n38209 = ~n38205 & n38208;
  assign n38210 = ~pi208 & ~n37776;
  assign n38211 = ~n38087 & n38210;
  assign n38212 = ~n38209 & ~n38211;
  assign n38213 = ~pi211 & n38212;
  assign n38214 = pi211 & n38200;
  assign n38215 = ~n37670 & ~n38214;
  assign n38216 = ~n38213 & n38215;
  assign n38217 = ~pi219 & ~n38216;
  assign n38218 = ~n38203 & n38217;
  assign n38219 = ~n38194 & n38218;
  assign n38220 = ~n38198 & ~n38219;
  assign n38221 = ~po1038 & ~n38220;
  assign n38222 = pi1152 & n38221;
  assign n38223 = ~n38193 & ~n38222;
  assign n38224 = pi213 & ~n38223;
  assign n38225 = ~pi209 & ~n38224;
  assign n38226 = ~n38172 & n38225;
  assign n38227 = ~n38059 & ~n38226;
  assign n38228 = pi219 & ~n37613;
  assign n38229 = pi214 & ~n37601;
  assign n38230 = ~pi212 & n38229;
  assign n38231 = ~pi219 & ~n38230;
  assign n38232 = ~n37608 & n38231;
  assign n38233 = pi213 & ~n38232;
  assign n38234 = ~n38228 & n38233;
  assign n38235 = n37664 & n38234;
  assign n38236 = ~n38227 & ~n38235;
  assign n38237 = pi230 & ~n38236;
  assign n38238 = ~pi230 & pi234;
  assign po391 = n38237 | n38238;
  assign n38240 = ~pi1156 & n37719;
  assign n38241 = ~n37795 & ~n38240;
  assign n38242 = pi207 & ~n38241;
  assign n38243 = ~pi207 & n37763;
  assign n38244 = ~n38242 & ~n38243;
  assign n38245 = pi208 & ~n38244;
  assign n38246 = ~n37766 & ~n38245;
  assign n38247 = ~pi1157 & ~n38246;
  assign n38248 = pi208 & pi1157;
  assign n38249 = ~n37773 & ~n37805;
  assign n38250 = ~pi207 & ~n38249;
  assign n38251 = ~n38242 & ~n38250;
  assign n38252 = n38248 & ~n38251;
  assign n38253 = ~n37778 & ~n38252;
  assign n38254 = ~n38247 & n38253;
  assign n38255 = ~pi211 & ~n38254;
  assign n38256 = ~n37726 & ~n37851;
  assign n38257 = pi207 & ~n38256;
  assign n38258 = ~pi207 & n37741;
  assign n38259 = ~n38257 & ~n38258;
  assign n38260 = pi208 & ~n38259;
  assign n38261 = ~n37742 & ~n38260;
  assign n38262 = ~pi1157 & ~n38261;
  assign n38263 = ~pi207 & ~n37752;
  assign n38264 = ~n38257 & ~n38263;
  assign n38265 = n38248 & ~n38264;
  assign n38266 = ~n37754 & ~n38265;
  assign n38267 = ~n38262 & n38266;
  assign n38268 = pi211 & ~n38267;
  assign n38269 = n10468 & ~n38268;
  assign n38270 = ~n38255 & n38269;
  assign n38271 = ~pi207 & ~n37813;
  assign n38272 = n10302 & ~n37726;
  assign n38273 = ~n38240 & n38272;
  assign n38274 = ~n37835 & ~n38273;
  assign n38275 = ~n38271 & n38274;
  assign n38276 = n37957 & n38076;
  assign n38277 = pi1157 & n38276;
  assign n38278 = ~n38275 & ~n38277;
  assign n38279 = n37661 & n38278;
  assign n38280 = pi211 & ~n38254;
  assign n38281 = ~pi207 & n37806;
  assign n38282 = pi208 & ~n38281;
  assign n38283 = ~n38013 & n38282;
  assign n38284 = ~n37808 & ~n38283;
  assign n38285 = pi1157 & n38284;
  assign n38286 = ~pi1157 & ~n38275;
  assign n38287 = ~pi211 & ~n38286;
  assign n38288 = ~n38285 & n38287;
  assign n38289 = ~n38280 & ~n38288;
  assign n38290 = n38157 & n38289;
  assign n38291 = ~n38279 & ~n38290;
  assign n38292 = ~n38270 & n38291;
  assign n38293 = ~pi219 & ~n38292;
  assign n38294 = ~pi211 & n38267;
  assign n38295 = pi211 & n38278;
  assign n38296 = ~n37670 & ~n38295;
  assign n38297 = ~n38294 & n38296;
  assign n38298 = n37670 & ~n38278;
  assign n38299 = pi219 & ~n38298;
  assign n38300 = ~n38297 & n38299;
  assign n38301 = pi209 & ~n38300;
  assign n38302 = ~n38293 & n38301;
  assign n38303 = n10302 & ~n38133;
  assign n38304 = ~n37791 & ~n37956;
  assign n38305 = ~n10302 & ~n38304;
  assign n38306 = ~n38303 & ~n38305;
  assign n38307 = n37661 & ~n38306;
  assign n38308 = ~pi1157 & n38306;
  assign n38309 = n37759 & ~n37858;
  assign n38310 = n37758 & n37857;
  assign n38311 = ~n38146 & ~n38310;
  assign n38312 = pi208 & n38311;
  assign n38313 = ~n38309 & ~n38312;
  assign n38314 = pi1157 & ~n38313;
  assign n38315 = ~pi211 & ~n38314;
  assign n38316 = ~n38308 & n38315;
  assign n38317 = ~n37776 & ~n38306;
  assign n38318 = pi211 & n38317;
  assign n38319 = ~n38316 & ~n38318;
  assign n38320 = ~n37670 & ~n38319;
  assign n38321 = ~pi211 & ~n38317;
  assign n38322 = n37716 & n37732;
  assign n38323 = ~n37633 & ~n37716;
  assign n38324 = ~n38146 & ~n38323;
  assign n38325 = pi208 & n38324;
  assign n38326 = ~n38322 & ~n38325;
  assign n38327 = pi211 & ~n38326;
  assign n38328 = ~n38321 & ~n38327;
  assign n38329 = n10468 & n38328;
  assign n38330 = ~n38320 & ~n38329;
  assign n38331 = ~n38307 & n38330;
  assign n38332 = ~pi219 & ~n38331;
  assign n38333 = ~pi211 & n38326;
  assign n38334 = pi211 & ~n38306;
  assign n38335 = ~n37670 & ~n38334;
  assign n38336 = ~n38333 & n38335;
  assign n38337 = n37670 & n38306;
  assign n38338 = pi219 & ~n38337;
  assign n38339 = ~n38336 & n38338;
  assign n38340 = ~pi209 & ~n38339;
  assign n38341 = ~n38332 & n38340;
  assign n38342 = ~n38302 & ~n38341;
  assign n38343 = ~po1038 & ~n38342;
  assign n38344 = pi213 & ~n38343;
  assign n38345 = pi219 & ~n38157;
  assign n38346 = pi219 & ~n37603;
  assign n38347 = ~pi214 & ~n37597;
  assign n38348 = ~n38229 & ~n38347;
  assign n38349 = pi212 & ~n38348;
  assign n38350 = ~pi219 & ~n38349;
  assign n38351 = ~n37598 & n38350;
  assign n38352 = ~n38346 & ~n38351;
  assign n38353 = ~n38345 & n38352;
  assign n38354 = po1038 & n38353;
  assign n38355 = n38344 & ~n38354;
  assign n38356 = ~pi299 & ~pi1157;
  assign n38357 = ~n38247 & n38356;
  assign n38358 = ~n37873 & ~n38285;
  assign n38359 = ~n38357 & n38358;
  assign n38360 = ~pi211 & ~n38359;
  assign n38361 = n38296 & ~n38360;
  assign n38362 = n38299 & ~n38361;
  assign n38363 = pi211 & n38359;
  assign n38364 = ~n37720 & ~n37852;
  assign n38365 = ~n37726 & ~n38364;
  assign n38366 = pi207 & ~n38365;
  assign n38367 = pi1154 & ~n37762;
  assign n38368 = ~n37812 & ~n38367;
  assign n38369 = ~pi207 & ~n37737;
  assign n38370 = ~n38368 & n38369;
  assign n38371 = ~n38366 & ~n38370;
  assign n38372 = pi208 & ~n38371;
  assign n38373 = ~n37816 & ~n38372;
  assign n38374 = ~pi1157 & ~n38373;
  assign n38375 = n37810 & ~n38284;
  assign n38376 = ~n38374 & ~n38375;
  assign n38377 = ~pi211 & ~n38376;
  assign n38378 = n10468 & ~n38377;
  assign n38379 = ~n38363 & n38378;
  assign n38380 = pi211 & n38376;
  assign n38381 = ~n38294 & ~n38380;
  assign n38382 = n38157 & ~n38381;
  assign n38383 = ~n38279 & ~n38382;
  assign n38384 = ~n38379 & n38383;
  assign n38385 = ~pi219 & ~n38384;
  assign n38386 = ~n38362 & ~n38385;
  assign n38387 = pi209 & ~n38386;
  assign n38388 = pi1153 & ~n37738;
  assign n38389 = ~n38078 & ~n38388;
  assign n38390 = n37633 & n38389;
  assign n38391 = pi208 & ~n38390;
  assign n38392 = ~n38310 & n38391;
  assign n38393 = ~n38309 & ~n38392;
  assign n38394 = ~n37782 & ~n38310;
  assign n38395 = ~n38393 & n38394;
  assign n38396 = ~n38313 & n38395;
  assign n38397 = ~pi211 & ~n38396;
  assign n38398 = n38335 & ~n38397;
  assign n38399 = n38338 & ~n38398;
  assign n38400 = pi207 & ~n38144;
  assign n38401 = ~pi207 & ~n37825;
  assign n38402 = ~n38400 & ~n38401;
  assign n38403 = pi208 & ~n38402;
  assign n38404 = n37759 & ~n37825;
  assign n38405 = ~n38403 & ~n38404;
  assign n38406 = pi211 & n38405;
  assign n38407 = ~n38333 & ~n38406;
  assign n38408 = ~n37670 & ~n38407;
  assign n38409 = ~pi211 & ~n38405;
  assign n38410 = pi211 & n38396;
  assign n38411 = ~n38409 & ~n38410;
  assign n38412 = n10468 & n38411;
  assign n38413 = ~n38307 & ~n38412;
  assign n38414 = ~n38408 & n38413;
  assign n38415 = ~pi219 & ~n38414;
  assign n38416 = ~n38399 & ~n38415;
  assign n38417 = ~pi209 & ~n38416;
  assign n38418 = ~n38387 & ~n38417;
  assign n38419 = ~po1038 & n38418;
  assign n38420 = ~pi219 & po1038;
  assign n38421 = ~pi211 & po1038;
  assign n38422 = pi1153 & n38421;
  assign n38423 = ~n38420 & ~n38422;
  assign n38424 = n10468 & ~n38007;
  assign n38425 = ~pi219 & ~n38424;
  assign n38426 = ~n37605 & n38157;
  assign n38427 = n38425 & ~n38426;
  assign n38428 = ~n38345 & ~n38427;
  assign n38429 = ~n38423 & n38428;
  assign n38430 = ~pi213 & ~n38429;
  assign n38431 = ~n38419 & n38430;
  assign n38432 = ~n38355 & ~n38431;
  assign n38433 = pi230 & ~n38432;
  assign n38434 = ~pi230 & ~pi235;
  assign po392 = ~n38433 & ~n38434;
  assign n38436 = ~pi100 & n37375;
  assign n38437 = n37578 & ~n38436;
  assign n38438 = ~n6095 & ~n38437;
  assign n38439 = ~pi75 & ~n38438;
  assign n38440 = ~n7253 & ~n38439;
  assign n38441 = ~pi92 & ~n38440;
  assign n38442 = n15138 & ~n38441;
  assign n38443 = ~pi74 & ~n38442;
  assign n38444 = n6093 & ~n38443;
  assign n38445 = ~pi56 & ~n38444;
  assign n38446 = ~n6264 & ~n38445;
  assign n38447 = ~pi62 & ~n38446;
  assign po393 = n13319 & ~n38447;
  assign n38449 = pi211 & pi1157;
  assign n38450 = ~pi211 & pi1158;
  assign n38451 = ~n38449 & ~n38450;
  assign n38452 = n37594 & ~n38451;
  assign n38453 = n38350 & ~n38452;
  assign n38454 = po1038 & n37599;
  assign n38455 = n37594 & n38454;
  assign n38456 = ~n38420 & ~n38455;
  assign n38457 = ~pi214 & ~n37603;
  assign n38458 = pi212 & ~n38457;
  assign n38459 = pi214 & ~n37613;
  assign n38460 = po1038 & ~n38459;
  assign n38461 = n38458 & n38460;
  assign n38462 = n38456 & ~n38461;
  assign n38463 = ~n38453 & ~n38462;
  assign n38464 = ~pi213 & ~n38463;
  assign n38465 = pi199 & pi1143;
  assign n38466 = ~pi200 & ~n38465;
  assign n38467 = ~n37626 & n38466;
  assign n38468 = ~n37629 & n38135;
  assign n38469 = ~n38467 & n38468;
  assign n38470 = pi200 & ~n37626;
  assign n38471 = ~pi199 & pi1145;
  assign n38472 = n38466 & ~n38471;
  assign n38473 = ~n38470 & ~n38472;
  assign n38474 = n37957 & n38473;
  assign n38475 = ~n38469 & ~n38474;
  assign n38476 = ~pi299 & ~n38475;
  assign n38477 = n37645 & ~n38453;
  assign n38478 = n37594 & n37776;
  assign n38479 = ~pi214 & ~n37647;
  assign n38480 = pi214 & ~n37649;
  assign n38481 = pi212 & ~n38480;
  assign n38482 = ~n38479 & n38481;
  assign n38483 = ~n38478 & ~n38482;
  assign n38484 = n10522 & ~n38483;
  assign n38485 = ~n38477 & ~n38484;
  assign n38486 = ~n38476 & n38485;
  assign n38487 = ~po1038 & ~n38486;
  assign n38488 = n38464 & ~n38487;
  assign n38489 = ~pi211 & pi1145;
  assign n38490 = pi211 & pi1144;
  assign n38491 = ~n38489 & ~n38490;
  assign n38492 = ~n10468 & n38491;
  assign n38493 = pi212 & ~n37668;
  assign n38494 = n37670 & ~n38493;
  assign n38495 = ~n38492 & ~n38494;
  assign n38496 = ~pi219 & ~n38495;
  assign n38497 = pi219 & ~n37672;
  assign n38498 = n37664 & ~n38497;
  assign n38499 = ~n38496 & n38498;
  assign n38500 = n37645 & n38495;
  assign n38501 = pi299 & n38091;
  assign n38502 = n37672 & n38501;
  assign n38503 = ~n38476 & ~n38502;
  assign n38504 = ~n38500 & n38503;
  assign n38505 = ~po1038 & ~n38504;
  assign n38506 = ~n38499 & ~n38505;
  assign n38507 = pi213 & n38506;
  assign n38508 = pi209 & ~n38507;
  assign n38509 = ~n38488 & n38508;
  assign n38510 = pi1158 & n38076;
  assign n38511 = ~pi199 & ~pi1158;
  assign n38512 = pi1156 & ~n38511;
  assign n38513 = ~n38510 & ~n38512;
  assign n38514 = ~pi200 & pi207;
  assign n38515 = ~n38513 & n38514;
  assign n38516 = ~pi208 & ~pi299;
  assign n38517 = n38515 & n38516;
  assign n38518 = pi207 & n37727;
  assign n38519 = ~n38271 & ~n38518;
  assign n38520 = pi208 & n38519;
  assign n38521 = ~n38517 & ~n38520;
  assign n38522 = ~pi1157 & ~n38521;
  assign n38523 = pi1156 & n37747;
  assign n38524 = ~pi200 & ~pi1158;
  assign n38525 = ~pi199 & ~n38524;
  assign n38526 = ~n38523 & ~n38525;
  assign n38527 = n37633 & ~n38526;
  assign n38528 = ~pi208 & n38527;
  assign n38529 = ~pi207 & n37774;
  assign n38530 = ~n38518 & ~n38529;
  assign n38531 = pi208 & n38530;
  assign n38532 = ~n38528 & ~n38531;
  assign n38533 = pi1157 & ~n38532;
  assign n38534 = ~n38522 & ~n38533;
  assign n38535 = ~n37662 & n38534;
  assign n38536 = pi207 & ~n37796;
  assign n38537 = ~n38250 & ~n38536;
  assign n38538 = n38248 & ~n38537;
  assign n38539 = ~n37776 & ~n38527;
  assign n38540 = n37743 & ~n38539;
  assign n38541 = ~n38538 & ~n38540;
  assign n38542 = n38210 & ~n38515;
  assign n38543 = ~pi1157 & ~n38542;
  assign n38544 = ~n38243 & ~n38536;
  assign n38545 = pi208 & n38544;
  assign n38546 = n38543 & ~n38545;
  assign n38547 = n38541 & ~n38546;
  assign n38548 = n37594 & n38547;
  assign n38549 = ~n37647 & n37727;
  assign n38550 = pi207 & ~n38549;
  assign n38551 = ~n38263 & ~n38550;
  assign n38552 = n38248 & ~n38551;
  assign n38553 = ~n38515 & ~n38525;
  assign n38554 = n37633 & ~n38553;
  assign n38555 = ~n37647 & ~n38554;
  assign n38556 = n37743 & ~n38555;
  assign n38557 = ~n38552 & ~n38556;
  assign n38558 = ~pi208 & n37647;
  assign n38559 = ~n38258 & ~n38550;
  assign n38560 = pi208 & ~n38559;
  assign n38561 = ~n38517 & ~n38560;
  assign n38562 = ~n38558 & n38561;
  assign n38563 = ~pi1157 & ~n38562;
  assign n38564 = n38557 & ~n38563;
  assign n38565 = ~pi214 & ~n38564;
  assign n38566 = ~pi207 & ~n37806;
  assign n38567 = ~n37809 & n38566;
  assign n38568 = pi1157 & ~n38567;
  assign n38569 = ~pi1157 & ~n38517;
  assign n38570 = ~n38370 & n38569;
  assign n38571 = ~n38568 & ~n38570;
  assign n38572 = pi208 & ~n37968;
  assign n38573 = ~n38571 & n38572;
  assign n38574 = pi299 & pi1158;
  assign n38575 = ~n38517 & ~n38574;
  assign n38576 = ~n37743 & ~n38575;
  assign n38577 = ~n37743 & ~n38576;
  assign n38578 = n38554 & ~n38577;
  assign n38579 = ~pi208 & ~n38578;
  assign n38580 = ~n37649 & n38579;
  assign n38581 = ~n38573 & ~n38580;
  assign n38582 = pi214 & n38581;
  assign n38583 = pi212 & ~n38582;
  assign n38584 = ~n38565 & n38583;
  assign n38585 = ~n38548 & ~n38584;
  assign n38586 = ~pi211 & ~n38585;
  assign n38587 = ~n38535 & ~n38586;
  assign n38588 = pi219 & ~n38587;
  assign n38589 = n37706 & ~n38547;
  assign n38590 = n37704 & ~n38564;
  assign n38591 = ~pi299 & n38526;
  assign n38592 = n37759 & ~n38591;
  assign n38593 = ~n38014 & n38282;
  assign n38594 = ~n38592 & ~n38593;
  assign n38595 = pi1157 & ~n38594;
  assign n38596 = ~n38522 & ~n38595;
  assign n38597 = n37705 & ~n38596;
  assign n38598 = ~n38590 & ~n38597;
  assign n38599 = ~n38589 & n38598;
  assign n38600 = pi212 & ~n38599;
  assign n38601 = ~pi214 & n38534;
  assign n38602 = ~pi212 & ~n38601;
  assign n38603 = pi211 & n38596;
  assign n38604 = pi1158 & n37854;
  assign n38605 = ~pi1158 & n37727;
  assign n38606 = pi207 & ~n38605;
  assign n38607 = ~n38604 & n38606;
  assign n38608 = pi299 & ~pi1158;
  assign n38609 = n38566 & ~n38608;
  assign n38610 = ~n38607 & ~n38609;
  assign n38611 = n38248 & ~n38610;
  assign n38612 = pi207 & ~n10615;
  assign n38613 = ~pi299 & ~n38612;
  assign n38614 = pi1158 & ~n38613;
  assign n38615 = n37711 & ~n37750;
  assign n38616 = ~n38510 & ~n38615;
  assign n38617 = pi1157 & n38616;
  assign n38618 = pi207 & ~n38617;
  assign n38619 = ~n38614 & ~n38618;
  assign n38620 = n37743 & ~n38619;
  assign n38621 = ~pi211 & ~n38620;
  assign n38622 = ~n38611 & n38621;
  assign n38623 = ~pi207 & ~n38608;
  assign n38624 = ~n37764 & n38623;
  assign n38625 = ~n38607 & ~n38624;
  assign n38626 = pi208 & n38625;
  assign n38627 = ~pi1157 & ~n38626;
  assign n38628 = ~pi208 & ~n38614;
  assign n38629 = ~n38517 & n38628;
  assign n38630 = n38627 & ~n38629;
  assign n38631 = n38622 & ~n38630;
  assign n38632 = ~n38603 & ~n38631;
  assign n38633 = pi214 & ~n38632;
  assign n38634 = n38602 & ~n38633;
  assign n38635 = ~pi219 & ~n38634;
  assign n38636 = ~n38600 & n38635;
  assign n38637 = ~po1038 & ~n38636;
  assign n38638 = ~n38588 & n38637;
  assign n38639 = n38464 & ~n38638;
  assign n38640 = ~pi209 & ~n38639;
  assign n38641 = ~n37912 & n38579;
  assign n38642 = pi207 & ~n37913;
  assign n38643 = pi208 & ~n38642;
  assign n38644 = ~pi200 & pi1157;
  assign n38645 = ~pi199 & n38644;
  assign n38646 = n37764 & ~n38645;
  assign n38647 = ~pi207 & ~n37920;
  assign n38648 = ~n38646 & n38647;
  assign n38649 = n38643 & ~n38648;
  assign n38650 = ~n38641 & ~n38649;
  assign n38651 = n37662 & ~n38650;
  assign n38652 = ~n38535 & ~n38651;
  assign n38653 = pi219 & ~n38652;
  assign n38654 = pi299 & pi1145;
  assign n38655 = ~n37894 & ~n38654;
  assign n38656 = pi207 & ~n38655;
  assign n38657 = pi208 & ~n38656;
  assign n38658 = pi299 & ~pi1145;
  assign n38659 = ~pi207 & ~n38658;
  assign n38660 = ~n38646 & n38659;
  assign n38661 = n38657 & ~n38660;
  assign n38662 = ~pi208 & ~n38654;
  assign n38663 = ~pi1157 & ~n38514;
  assign n38664 = n38527 & ~n38663;
  assign n38665 = n38662 & ~n38664;
  assign n38666 = ~n38661 & ~n38665;
  assign n38667 = ~pi211 & ~n38666;
  assign n38668 = ~n37893 & n38579;
  assign n38669 = pi207 & ~n37895;
  assign n38670 = pi208 & ~n38669;
  assign n38671 = ~pi207 & ~n37900;
  assign n38672 = ~n38646 & n38671;
  assign n38673 = n38670 & ~n38672;
  assign n38674 = ~n38668 & ~n38673;
  assign n38675 = pi211 & ~n38674;
  assign n38676 = ~n38667 & ~n38675;
  assign n38677 = ~pi214 & ~n38676;
  assign n38678 = ~pi211 & n38674;
  assign n38679 = pi214 & ~n38678;
  assign n38680 = pi211 & n38650;
  assign n38681 = n38679 & ~n38680;
  assign n38682 = ~n38677 & ~n38681;
  assign n38683 = pi212 & n38682;
  assign n38684 = pi214 & ~n38676;
  assign n38685 = n38602 & ~n38684;
  assign n38686 = ~pi219 & ~n38685;
  assign n38687 = ~n38683 & n38686;
  assign n38688 = ~n38653 & ~n38687;
  assign n38689 = ~po1038 & n38688;
  assign n38690 = ~n38499 & ~n38689;
  assign n38691 = pi213 & n38690;
  assign n38692 = n38640 & ~n38691;
  assign n38693 = ~n38509 & ~n38692;
  assign n38694 = pi230 & ~n38693;
  assign n38695 = ~pi230 & ~pi237;
  assign po394 = n38694 | n38695;
  assign n38697 = pi1151 & ~po1038;
  assign n38698 = ~n37714 & n38112;
  assign n38699 = n37633 & ~n37710;
  assign n38700 = pi208 & ~n38699;
  assign n38701 = pi200 & n37758;
  assign n38702 = n38700 & ~n38701;
  assign n38703 = ~n38698 & ~n38702;
  assign n38704 = ~pi211 & ~n38703;
  assign n38705 = n37771 & n37957;
  assign n38706 = n37710 & n38135;
  assign n38707 = ~n38705 & ~n38706;
  assign n38708 = pi211 & ~n38707;
  assign n38709 = ~n38704 & ~n38708;
  assign n38710 = ~n38106 & ~n38709;
  assign n38711 = ~n38083 & ~n38707;
  assign n38712 = n37661 & ~n38711;
  assign n38713 = n38710 & ~n38712;
  assign n38714 = pi219 & ~n38713;
  assign n38715 = ~n38106 & ~n38703;
  assign n38716 = n37704 & ~n38715;
  assign n38717 = ~n37649 & n37706;
  assign n38718 = ~n38711 & n38717;
  assign n38719 = ~n37647 & ~n38711;
  assign n38720 = n37705 & n38719;
  assign n38721 = pi212 & ~n38720;
  assign n38722 = ~n38718 & n38721;
  assign n38723 = ~n38716 & n38722;
  assign n38724 = pi299 & ~n37605;
  assign n38725 = ~n38711 & ~n38724;
  assign n38726 = pi1153 & n38276;
  assign n38727 = n10614 & n37957;
  assign n38728 = n38110 & ~n38727;
  assign n38729 = ~pi214 & ~n38728;
  assign n38730 = ~n38726 & n38729;
  assign n38731 = ~pi212 & ~n38730;
  assign n38732 = ~n38725 & n38731;
  assign n38733 = ~n38723 & ~n38732;
  assign n38734 = ~pi219 & n38733;
  assign n38735 = ~n38714 & ~n38734;
  assign n38736 = n38697 & n38735;
  assign n38737 = ~pi1151 & ~po1038;
  assign n38738 = ~n37649 & ~n38726;
  assign n38739 = ~pi211 & ~n38738;
  assign n38740 = ~pi299 & ~n38727;
  assign n38741 = n38006 & ~n38740;
  assign n38742 = n10468 & ~n38741;
  assign n38743 = ~n38739 & n38742;
  assign n38744 = ~n37670 & ~n38724;
  assign n38745 = ~n38726 & n38744;
  assign n38746 = ~n38743 & ~n38745;
  assign n38747 = ~pi219 & ~n38746;
  assign n38748 = ~n12743 & ~n38740;
  assign n38749 = ~pi214 & ~n38276;
  assign n38750 = ~pi212 & n38749;
  assign n38751 = n38748 & ~n38750;
  assign n38752 = pi1153 & n38751;
  assign n38753 = ~n37930 & ~n38752;
  assign n38754 = ~n38747 & ~n38753;
  assign n38755 = n38737 & n38754;
  assign n38756 = ~pi1152 & ~n38755;
  assign n38757 = ~n38736 & n38756;
  assign n38758 = pi1153 & ~n38740;
  assign n38759 = ~n37957 & ~n38612;
  assign n38760 = ~n10302 & n37760;
  assign n38761 = ~n38759 & ~n38760;
  assign n38762 = n38740 & n38761;
  assign n38763 = ~n38758 & ~n38762;
  assign n38764 = pi211 & ~n38763;
  assign n38765 = n37759 & ~n38068;
  assign n38766 = pi208 & pi299;
  assign n38767 = ~n10302 & n38066;
  assign n38768 = pi200 & pi207;
  assign n38769 = ~pi199 & ~n38768;
  assign n38770 = ~pi299 & ~n38769;
  assign n38771 = pi208 & ~n38770;
  assign n38772 = ~pi299 & n38771;
  assign n38773 = ~n38767 & n38772;
  assign n38774 = ~n38766 & ~n38773;
  assign n38775 = ~n38765 & n38774;
  assign n38776 = ~pi211 & ~n37809;
  assign n38777 = ~n38775 & n38776;
  assign n38778 = ~n38764 & ~n38777;
  assign n38779 = n10468 & ~n38778;
  assign n38780 = pi299 & n37605;
  assign n38781 = ~n37670 & ~n38775;
  assign n38782 = ~n38780 & n38781;
  assign n38783 = ~n38779 & ~n38782;
  assign n38784 = ~pi219 & ~n38783;
  assign n38785 = n11156 & n37641;
  assign n38786 = ~n38772 & ~n38785;
  assign n38787 = ~n38767 & ~n38786;
  assign n38788 = ~pi211 & n37651;
  assign n38789 = ~n37661 & n38788;
  assign n38790 = ~n38787 & ~n38789;
  assign n38791 = ~n37930 & ~n38790;
  assign n38792 = ~n38784 & ~n38791;
  assign n38793 = n38737 & ~n38792;
  assign n38794 = pi219 & ~n38728;
  assign n38795 = ~n38752 & n38794;
  assign n38796 = ~n38741 & ~n38777;
  assign n38797 = ~n38728 & n38796;
  assign n38798 = n10468 & ~n38797;
  assign n38799 = ~n38726 & ~n38728;
  assign n38800 = n37661 & ~n38799;
  assign n38801 = n37748 & n38767;
  assign n38802 = ~n38111 & ~n38801;
  assign n38803 = ~pi211 & n38802;
  assign n38804 = ~n37850 & n38803;
  assign n38805 = pi211 & n38802;
  assign n38806 = ~n37809 & n38805;
  assign n38807 = ~n38804 & ~n38806;
  assign n38808 = ~n37670 & ~n38807;
  assign n38809 = ~pi219 & ~n38808;
  assign n38810 = ~n38800 & n38809;
  assign n38811 = ~n38798 & n38810;
  assign n38812 = ~n38795 & ~n38811;
  assign n38813 = n38697 & n38812;
  assign n38814 = pi1152 & ~n38813;
  assign n38815 = ~n38793 & n38814;
  assign n38816 = ~n38757 & ~n38815;
  assign n38817 = ~pi209 & ~n38816;
  assign n38818 = pi1153 & ~pi1154;
  assign n38819 = n37711 & n38818;
  assign n38820 = ~n38078 & ~n38819;
  assign n38821 = n10302 & n38820;
  assign n38822 = ~n38305 & ~n38821;
  assign n38823 = ~pi214 & ~n38822;
  assign n38824 = ~pi212 & n38823;
  assign n38825 = n37704 & n38395;
  assign n38826 = ~n38323 & n38391;
  assign n38827 = ~n38322 & ~n38826;
  assign n38828 = ~pi211 & ~n38827;
  assign n38829 = ~pi214 & n38828;
  assign n38830 = ~n37633 & n37825;
  assign n38831 = n38391 & ~n38830;
  assign n38832 = ~n38404 & ~n38831;
  assign n38833 = n37706 & ~n38832;
  assign n38834 = pi212 & ~n38833;
  assign n38835 = ~n38829 & n38834;
  assign n38836 = ~n38825 & n38835;
  assign n38837 = pi211 & ~n38832;
  assign n38838 = ~n38828 & ~n38837;
  assign n38839 = n37594 & n38838;
  assign n38840 = ~n38836 & ~n38839;
  assign n38841 = ~pi219 & ~n38840;
  assign n38842 = pi211 & n38822;
  assign n38843 = ~pi211 & n38395;
  assign n38844 = ~n38842 & ~n38843;
  assign n38845 = n38091 & n38844;
  assign n38846 = ~n38841 & ~n38845;
  assign n38847 = ~n38824 & n38846;
  assign n38848 = ~po1038 & n38847;
  assign n38849 = pi209 & ~n38848;
  assign n38850 = ~n38817 & ~n38849;
  assign n38851 = ~pi211 & ~pi1153;
  assign n38852 = pi219 & n38851;
  assign n38853 = ~n38427 & ~n38852;
  assign n38854 = n37664 & n38853;
  assign n38855 = ~n38850 & ~n38854;
  assign n38856 = pi213 & ~n38855;
  assign n38857 = ~n10469 & n37930;
  assign n38858 = po1038 & n38857;
  assign n38859 = ~n10524 & ~n37611;
  assign n38860 = n38858 & ~n38859;
  assign n38861 = ~n10470 & n37664;
  assign n38862 = pi1151 & ~n38861;
  assign n38863 = ~n38860 & n38862;
  assign n38864 = ~pi211 & ~n38393;
  assign n38865 = ~n38842 & ~n38864;
  assign n38866 = ~n37661 & n38865;
  assign n38867 = ~n38824 & ~n38866;
  assign n38868 = pi219 & ~n38867;
  assign n38869 = ~po1038 & ~n38868;
  assign n38870 = pi211 & ~n38393;
  assign n38871 = ~n38843 & ~n38870;
  assign n38872 = ~pi214 & ~n38871;
  assign n38873 = pi214 & ~n38393;
  assign n38874 = ~n38872 & ~n38873;
  assign n38875 = pi212 & ~n38874;
  assign n38876 = pi214 & n38871;
  assign n38877 = ~pi212 & ~n38823;
  assign n38878 = ~n38876 & n38877;
  assign n38879 = ~pi219 & ~n38878;
  assign n38880 = ~n38875 & n38879;
  assign n38881 = n38869 & ~n38880;
  assign n38882 = n38863 & ~n38881;
  assign n38883 = ~pi1151 & ~n38860;
  assign n38884 = pi214 & ~n38865;
  assign n38885 = ~n38872 & ~n38884;
  assign n38886 = pi212 & ~n38885;
  assign n38887 = n38879 & ~n38886;
  assign n38888 = pi219 & ~n38822;
  assign n38889 = ~po1038 & ~n38888;
  assign n38890 = ~n38887 & n38889;
  assign n38891 = n38883 & ~n38890;
  assign n38892 = pi1152 & ~n38891;
  assign n38893 = ~n38882 & n38892;
  assign n38894 = pi214 & n38844;
  assign n38895 = ~n38823 & ~n38894;
  assign n38896 = ~pi212 & ~n38895;
  assign n38897 = ~pi211 & n38822;
  assign n38898 = ~n38870 & ~n38897;
  assign n38899 = pi214 & ~n38898;
  assign n38900 = ~pi214 & ~n38844;
  assign n38901 = pi212 & ~n38900;
  assign n38902 = ~n38899 & n38901;
  assign n38903 = ~n38896 & ~n38902;
  assign n38904 = ~pi219 & ~n38903;
  assign n38905 = n38869 & ~n38904;
  assign n38906 = n10523 & n38858;
  assign n38907 = pi1153 & n38906;
  assign n38908 = n38862 & ~n38907;
  assign n38909 = ~n38905 & n38908;
  assign n38910 = ~pi1151 & ~n38907;
  assign n38911 = ~pi219 & n38157;
  assign n38912 = n38844 & n38911;
  assign n38913 = ~n38822 & ~n38911;
  assign n38914 = ~po1038 & ~n38913;
  assign n38915 = ~n38912 & n38914;
  assign n38916 = n38910 & ~n38915;
  assign n38917 = ~pi1152 & ~n38916;
  assign n38918 = ~n38909 & n38917;
  assign n38919 = ~n38893 & ~n38918;
  assign n38920 = pi209 & n38919;
  assign n38921 = ~pi211 & pi299;
  assign n38922 = ~n38711 & ~n38921;
  assign n38923 = ~n38712 & ~n38922;
  assign n38924 = pi219 & ~n38923;
  assign n38925 = ~pi214 & n38710;
  assign n38926 = ~n12743 & ~n38726;
  assign n38927 = ~n38711 & n38926;
  assign n38928 = pi214 & ~n38927;
  assign n38929 = pi212 & ~n38928;
  assign n38930 = ~n38925 & n38929;
  assign n38931 = ~pi212 & ~n38713;
  assign n38932 = ~n38930 & ~n38931;
  assign n38933 = ~pi219 & ~n38932;
  assign n38934 = ~po1038 & ~n38933;
  assign n38935 = ~n38924 & n38934;
  assign n38936 = n38908 & ~n38935;
  assign n38937 = pi219 & ~n38276;
  assign n38938 = ~po1038 & ~n38937;
  assign n38939 = n38751 & n38938;
  assign n38940 = ~n38749 & ~n38926;
  assign n38941 = pi212 & n38940;
  assign n38942 = ~pi219 & ~n38941;
  assign n38943 = ~n38276 & n38942;
  assign n38944 = pi214 & ~n38748;
  assign n38945 = pi212 & ~n38740;
  assign n38946 = ~pi211 & n38749;
  assign n38947 = n38945 & ~n38946;
  assign n38948 = ~n38944 & n38947;
  assign n38949 = n38751 & ~n38948;
  assign n38950 = n37651 & n38949;
  assign n38951 = n38943 & ~n38950;
  assign n38952 = pi1153 & ~n38951;
  assign n38953 = n38939 & n38952;
  assign n38954 = n38910 & ~n38953;
  assign n38955 = ~pi1152 & ~n38954;
  assign n38956 = ~n38936 & n38955;
  assign n38957 = n38799 & ~n38803;
  assign n38958 = pi214 & n38957;
  assign n38959 = ~n38730 & ~n38958;
  assign n38960 = ~pi212 & ~n38959;
  assign n38961 = ~n38957 & ~n38960;
  assign n38962 = pi219 & ~n38961;
  assign n38963 = ~po1038 & ~n38962;
  assign n38964 = ~n38758 & ~n38805;
  assign n38965 = pi214 & ~n38728;
  assign n38966 = n38964 & n38965;
  assign n38967 = n38731 & ~n38966;
  assign n38968 = ~n38959 & n38964;
  assign n38969 = pi212 & ~n38968;
  assign n38970 = ~pi219 & ~n38969;
  assign n38971 = ~n38967 & n38970;
  assign n38972 = n38963 & ~n38971;
  assign n38973 = n38863 & ~n38972;
  assign n38974 = pi219 & ~n38787;
  assign n38975 = ~po1038 & ~n38974;
  assign n38976 = n37670 & n38787;
  assign n38977 = n10468 & n38921;
  assign n38978 = ~pi211 & n38763;
  assign n38979 = n38781 & ~n38978;
  assign n38980 = ~pi219 & ~n38979;
  assign n38981 = ~n38977 & n38980;
  assign n38982 = ~n38976 & n38981;
  assign n38983 = n38975 & ~n38982;
  assign n38984 = n38883 & ~n38983;
  assign n38985 = pi1152 & ~n38984;
  assign n38986 = ~n38973 & n38985;
  assign n38987 = ~n38956 & ~n38986;
  assign n38988 = ~pi209 & n38987;
  assign n38989 = ~pi213 & ~n38988;
  assign n38990 = ~n38920 & n38989;
  assign n38991 = ~n38856 & ~n38990;
  assign n38992 = pi230 & ~n38991;
  assign n38993 = ~pi230 & pi238;
  assign po395 = n38992 | n38993;
  assign n38995 = ~pi219 & ~n38452;
  assign n38996 = ~n38456 & ~n38995;
  assign n38997 = pi212 & ~n38578;
  assign n38998 = ~po1038 & ~n38997;
  assign n38999 = ~pi214 & n38578;
  assign n39000 = ~pi212 & ~n38999;
  assign n39001 = pi219 & n39000;
  assign n39002 = pi211 & ~n38578;
  assign n39003 = n38182 & ~n38578;
  assign n39004 = pi214 & ~n39003;
  assign n39005 = ~n39002 & n39004;
  assign n39006 = n39001 & ~n39005;
  assign n39007 = pi209 & ~n39006;
  assign n39008 = ~pi219 & n39000;
  assign n39009 = pi1157 & ~n38766;
  assign n39010 = ~n38592 & n39009;
  assign n39011 = ~n38569 & ~n39010;
  assign n39012 = pi211 & ~n39011;
  assign n39013 = ~n38576 & n38621;
  assign n39014 = ~n39012 & ~n39013;
  assign n39015 = pi214 & n39014;
  assign n39016 = n39008 & ~n39015;
  assign n39017 = n39007 & ~n39016;
  assign n39018 = n38998 & n39017;
  assign n39019 = n37641 & ~n37727;
  assign n39020 = ~pi214 & n39019;
  assign n39021 = ~pi212 & ~n39020;
  assign n39022 = ~pi219 & n39021;
  assign n39023 = ~n37641 & n38574;
  assign n39024 = ~pi208 & n38607;
  assign n39025 = ~n39023 & ~n39024;
  assign n39026 = ~pi211 & ~n39025;
  assign n39027 = ~n38015 & n39009;
  assign n39028 = ~pi1157 & ~n39019;
  assign n39029 = pi211 & ~n39028;
  assign n39030 = ~n39027 & n39029;
  assign n39031 = ~n39026 & ~n39030;
  assign n39032 = pi214 & ~n39031;
  assign n39033 = n39022 & ~n39032;
  assign n39034 = pi219 & n39021;
  assign n39035 = pi211 & ~n39019;
  assign n39036 = pi214 & ~n39035;
  assign n39037 = ~n37985 & n38182;
  assign n39038 = n39036 & ~n39037;
  assign n39039 = n39034 & ~n39038;
  assign n39040 = pi212 & ~n39019;
  assign n39041 = ~po1038 & ~n39040;
  assign n39042 = ~n39039 & n39041;
  assign n39043 = ~pi209 & n39042;
  assign n39044 = ~n39033 & n39043;
  assign n39045 = pi213 & ~n39044;
  assign n39046 = ~n39018 & n39045;
  assign n39047 = ~n38996 & n39046;
  assign n39048 = ~n37649 & ~n37970;
  assign n39049 = n39036 & ~n39048;
  assign n39050 = n39034 & ~n39049;
  assign n39051 = pi211 & ~n37647;
  assign n39052 = ~n39019 & n39051;
  assign n39053 = ~n39037 & ~n39052;
  assign n39054 = pi214 & n39053;
  assign n39055 = n39022 & ~n39054;
  assign n39056 = ~n39050 & ~n39055;
  assign n39057 = n39041 & n39056;
  assign n39058 = ~pi209 & n39057;
  assign n39059 = ~pi213 & ~n39058;
  assign n39060 = ~n38578 & n39051;
  assign n39061 = n39004 & ~n39060;
  assign n39062 = n39008 & ~n39061;
  assign n39063 = ~pi211 & n37649;
  assign n39064 = ~n38578 & ~n39063;
  assign n39065 = pi214 & ~n39064;
  assign n39066 = n39001 & ~n39065;
  assign n39067 = ~n39062 & ~n39066;
  assign n39068 = n38998 & n39067;
  assign n39069 = pi209 & n39068;
  assign n39070 = n39059 & ~n39069;
  assign n39071 = po1038 & ~n38228;
  assign n39072 = n37594 & ~n38231;
  assign n39073 = n39071 & n39072;
  assign n39074 = n39070 & ~n39073;
  assign n39075 = ~n39047 & ~n39074;
  assign n39076 = pi230 & ~n39075;
  assign n39077 = ~pi230 & ~pi239;
  assign po396 = ~n39076 & ~n39077;
  assign n39079 = ~po1038 & ~n37663;
  assign n39080 = n37693 & n39079;
  assign n39081 = ~po1038 & n38110;
  assign n39082 = ~n39080 & ~n39081;
  assign n39083 = ~n37661 & n37664;
  assign n39084 = n39082 & ~n39083;
  assign n39085 = pi1147 & n39084;
  assign n39086 = pi1149 & ~n39085;
  assign n39087 = ~po1038 & ~n38786;
  assign n39088 = ~n38938 & ~n39087;
  assign n39089 = ~pi214 & n38786;
  assign n39090 = ~pi212 & ~n39089;
  assign n39091 = ~pi299 & n38786;
  assign n39092 = n39090 & ~n39091;
  assign n39093 = ~pi219 & ~n39092;
  assign n39094 = ~pi211 & ~n39091;
  assign n39095 = pi211 & ~n38786;
  assign n39096 = pi214 & ~n39095;
  assign n39097 = ~n39094 & n39096;
  assign n39098 = pi212 & ~n39097;
  assign n39099 = ~n39091 & n39098;
  assign n39100 = n39093 & ~n39099;
  assign n39101 = ~n39088 & ~n39100;
  assign n39102 = ~n38858 & ~n39101;
  assign n39103 = ~pi1147 & n39102;
  assign n39104 = n39086 & ~n39103;
  assign n39105 = ~n39080 & ~n39083;
  assign n39106 = pi212 & ~n37705;
  assign n39107 = pi211 & n37594;
  assign n39108 = ~pi219 & ~n39107;
  assign n39109 = ~n39106 & n39108;
  assign n39110 = ~n39105 & ~n39109;
  assign n39111 = ~po1038 & n38728;
  assign n39112 = ~n39110 & ~n39111;
  assign n39113 = pi1147 & n39112;
  assign n39114 = ~pi1149 & ~n39113;
  assign n39115 = pi212 & n37706;
  assign n39116 = ~n39107 & ~n39115;
  assign n39117 = n38420 & ~n39116;
  assign n39118 = pi299 & n37704;
  assign n39119 = ~n38762 & ~n39118;
  assign n39120 = ~pi212 & ~n39119;
  assign n39121 = ~pi219 & ~n39120;
  assign n39122 = ~pi299 & ~n38761;
  assign n39123 = pi214 & ~n39122;
  assign n39124 = ~pi214 & n38762;
  assign n39125 = ~pi212 & ~n39124;
  assign n39126 = ~n39123 & n39125;
  assign n39127 = ~pi211 & ~n39122;
  assign n39128 = ~n38762 & ~n39127;
  assign n39129 = pi214 & ~n39128;
  assign n39130 = pi212 & ~n39129;
  assign n39131 = ~pi214 & ~n39122;
  assign n39132 = n39130 & ~n39131;
  assign n39133 = ~n39126 & ~n39132;
  assign n39134 = pi212 & ~n39122;
  assign n39135 = ~n38949 & n39134;
  assign n39136 = n39133 & n39135;
  assign n39137 = n39121 & ~n39136;
  assign n39138 = pi219 & ~n38762;
  assign n39139 = ~po1038 & ~n39138;
  assign n39140 = ~n39137 & n39139;
  assign n39141 = ~n39117 & ~n39140;
  assign n39142 = ~pi1147 & n39141;
  assign n39143 = n39114 & ~n39142;
  assign n39144 = ~n39104 & ~n39143;
  assign n39145 = pi1148 & ~n39144;
  assign n39146 = pi211 & ~n38703;
  assign n39147 = ~pi211 & ~n38707;
  assign n39148 = pi214 & ~n39147;
  assign n39149 = ~n39146 & n39148;
  assign n39150 = n10468 & ~n39149;
  assign n39151 = ~pi214 & n38707;
  assign n39152 = ~pi212 & ~n39151;
  assign n39153 = pi214 & n38709;
  assign n39154 = n39152 & ~n39153;
  assign n39155 = ~pi219 & ~n39154;
  assign n39156 = pi212 & ~n39149;
  assign n39157 = ~n38709 & n39156;
  assign n39158 = n39155 & ~n39157;
  assign n39159 = ~n39150 & n39158;
  assign n39160 = pi212 & ~n38709;
  assign n39161 = ~n39154 & ~n39160;
  assign n39162 = pi219 & n39161;
  assign n39163 = ~po1038 & ~n39162;
  assign n39164 = ~n39159 & n39163;
  assign n39165 = ~n38861 & ~n38906;
  assign n39166 = ~n39164 & n39165;
  assign n39167 = pi1147 & n39166;
  assign n39168 = n15973 & n38727;
  assign n39169 = n10523 & n37930;
  assign n39170 = ~n15973 & n39169;
  assign n39171 = ~n39168 & ~n39170;
  assign n39172 = ~pi1147 & n39171;
  assign n39173 = pi1149 & ~n39172;
  assign n39174 = ~n39167 & n39173;
  assign n39175 = pi212 & n39118;
  assign n39176 = pi299 & n39106;
  assign n39177 = ~n39118 & ~n39176;
  assign n39178 = ~n39175 & ~n39177;
  assign n39179 = ~n38728 & ~n39178;
  assign n39180 = ~pi219 & n39179;
  assign n39181 = ~pi299 & n37747;
  assign n39182 = n37957 & n39181;
  assign n39183 = ~n38706 & ~n39182;
  assign n39184 = ~pi299 & n39183;
  assign n39185 = ~pi219 & n39184;
  assign n39186 = ~n39180 & ~n39185;
  assign n39187 = ~pi211 & ~n39186;
  assign n39188 = ~pi212 & ~n38740;
  assign n39189 = ~n38749 & n39188;
  assign n39190 = ~n38921 & n39189;
  assign n39191 = ~pi219 & ~n39190;
  assign n39192 = ~n38948 & n39191;
  assign n39193 = n38938 & ~n39192;
  assign n39194 = ~n39082 & ~n39193;
  assign n39195 = ~n39184 & n39194;
  assign n39196 = ~n39187 & n39195;
  assign n39197 = ~n38861 & ~n39196;
  assign n39198 = ~pi1149 & ~n39197;
  assign n39199 = pi1147 & n39198;
  assign n39200 = ~n39174 & ~n39199;
  assign n39201 = ~pi1148 & ~n39200;
  assign n39202 = ~n39145 & ~n39201;
  assign n39203 = pi213 & ~n39202;
  assign n39204 = ~pi211 & n38654;
  assign n39205 = pi219 & ~n39204;
  assign n39206 = n39079 & ~n39205;
  assign n39207 = pi219 & n38707;
  assign n39208 = ~po1038 & ~n39207;
  assign n39209 = ~n39206 & ~n39208;
  assign n39210 = ~pi211 & pi1146;
  assign n39211 = pi211 & pi1145;
  assign n39212 = ~n39210 & ~n39211;
  assign n39213 = pi299 & ~n39212;
  assign n39214 = pi214 & ~n39213;
  assign n39215 = n38707 & n39214;
  assign n39216 = pi299 & pi1146;
  assign n39217 = pi211 & n39216;
  assign n39218 = ~pi214 & n38709;
  assign n39219 = ~n39217 & n39218;
  assign n39220 = ~n39215 & ~n39219;
  assign n39221 = pi212 & n39220;
  assign n39222 = n39153 & ~n39217;
  assign n39223 = n39152 & ~n39222;
  assign n39224 = ~pi219 & ~n39223;
  assign n39225 = ~n39221 & n39224;
  assign n39226 = ~n39209 & ~n39225;
  assign n39227 = pi214 & ~n39212;
  assign n39228 = pi211 & pi1146;
  assign n39229 = ~pi214 & n39228;
  assign n39230 = ~n39227 & ~n39229;
  assign n39231 = pi212 & ~n39230;
  assign n39232 = n37594 & n39228;
  assign n39233 = ~n39231 & ~n39232;
  assign n39234 = ~n38091 & n39233;
  assign n39235 = po1038 & n38489;
  assign n39236 = ~n38420 & ~n39235;
  assign n39237 = ~n39234 & ~n39236;
  assign n39238 = pi1147 & ~n38906;
  assign n39239 = ~n39237 & n39238;
  assign n39240 = ~n39226 & n39239;
  assign n39241 = pi219 & n39206;
  assign n39242 = ~pi1147 & ~n39237;
  assign n39243 = pi299 & ~n39233;
  assign n39244 = n35335 & n39243;
  assign n39245 = n39242 & ~n39244;
  assign n39246 = ~n39241 & n39245;
  assign n39247 = ~n39168 & n39246;
  assign n39248 = ~pi1148 & ~n39247;
  assign n39249 = ~n39240 & n39248;
  assign n39250 = pi299 & n37662;
  assign n39251 = pi219 & ~n39250;
  assign n39252 = n38786 & n39251;
  assign n39253 = ~po1038 & ~n39252;
  assign n39254 = n11156 & n39253;
  assign n39255 = ~n39206 & ~n39254;
  assign n39256 = n39090 & n39217;
  assign n39257 = ~pi212 & ~n38786;
  assign n39258 = ~pi219 & ~n39257;
  assign n39259 = ~n39256 & n39258;
  assign n39260 = pi212 & ~n39091;
  assign n39261 = pi299 & n39230;
  assign n39262 = n39260 & ~n39261;
  assign n39263 = n39259 & ~n39262;
  assign n39264 = ~n39255 & ~n39263;
  assign n39265 = n39242 & ~n39264;
  assign n39266 = pi1148 & ~n39265;
  assign n39267 = pi219 & ~n38110;
  assign n39268 = ~po1038 & ~n39267;
  assign n39269 = pi212 & ~n38111;
  assign n39270 = pi214 & n38195;
  assign n39271 = n39269 & ~n39270;
  assign n39272 = pi214 & pi299;
  assign n39273 = ~n38110 & ~n39272;
  assign n39274 = ~pi212 & ~n39273;
  assign n39275 = ~pi219 & ~n39274;
  assign n39276 = ~n39271 & n39275;
  assign n39277 = n39268 & ~n39276;
  assign n39278 = ~n38195 & n39277;
  assign n39279 = ~n39176 & n39278;
  assign n39280 = n39239 & ~n39279;
  assign n39281 = ~n39241 & n39280;
  assign n39282 = ~n39244 & n39281;
  assign n39283 = n39266 & ~n39282;
  assign n39284 = pi1149 & ~n39283;
  assign n39285 = ~n39249 & n39284;
  assign n39286 = ~po1038 & n38762;
  assign n39287 = n39246 & ~n39286;
  assign n39288 = ~n39111 & ~n39206;
  assign n39289 = n37661 & n38728;
  assign n39290 = ~pi219 & ~n39289;
  assign n39291 = ~n38728 & ~n39213;
  assign n39292 = n10468 & ~n39291;
  assign n39293 = ~n38921 & ~n39217;
  assign n39294 = ~n38728 & n39293;
  assign n39295 = n38157 & ~n39294;
  assign n39296 = ~n39292 & ~n39295;
  assign n39297 = n39290 & n39296;
  assign n39298 = ~n39288 & ~n39297;
  assign n39299 = n39239 & ~n39298;
  assign n39300 = pi1148 & ~n39299;
  assign n39301 = ~n39287 & n39300;
  assign n39302 = ~pi1146 & n12743;
  assign n39303 = n38157 & ~n39302;
  assign n39304 = ~n39292 & ~n39303;
  assign n39305 = ~pi219 & ~n39184;
  assign n39306 = ~n39304 & n39305;
  assign n39307 = ~n37930 & ~n39183;
  assign n39308 = n38091 & n39204;
  assign n39309 = ~n39307 & ~n39308;
  assign n39310 = ~n39306 & n39309;
  assign n39311 = ~po1038 & ~n39310;
  assign n39312 = n39239 & ~n39311;
  assign n39313 = ~pi1148 & ~n39246;
  assign n39314 = ~n39312 & n39313;
  assign n39315 = ~n39301 & ~n39314;
  assign n39316 = ~pi1149 & n39315;
  assign n39317 = ~pi213 & ~n39316;
  assign n39318 = ~n39285 & n39317;
  assign n39319 = pi209 & ~n39318;
  assign n39320 = ~n39203 & n39319;
  assign n39321 = ~pi199 & pi1146;
  assign n39322 = pi200 & ~n39321;
  assign n39323 = ~pi299 & ~n39322;
  assign n39324 = pi199 & pi1145;
  assign n39325 = n37747 & ~n39324;
  assign n39326 = n39323 & ~n39325;
  assign n39327 = ~n10302 & ~n39326;
  assign n39328 = pi200 & ~n38471;
  assign n39329 = ~pi299 & ~n39328;
  assign n39330 = ~pi200 & ~n39324;
  assign n39331 = ~n39321 & n39330;
  assign n39332 = pi207 & ~n39331;
  assign n39333 = n39329 & n39332;
  assign n39334 = ~n37957 & ~n39333;
  assign n39335 = ~n39327 & ~n39334;
  assign n39336 = pi219 & ~n39308;
  assign n39337 = ~n39335 & n39336;
  assign n39338 = n39251 & n39337;
  assign n39339 = ~po1038 & ~n39338;
  assign n39340 = ~n39216 & ~n39335;
  assign n39341 = pi208 & ~n39340;
  assign n39342 = ~n39335 & ~n39341;
  assign n39343 = ~pi299 & n39342;
  assign n39344 = pi211 & ~n39343;
  assign n39345 = ~n37758 & n39341;
  assign n39346 = n39330 & ~n39345;
  assign n39347 = ~n39342 & ~n39346;
  assign n39348 = ~pi299 & ~n39347;
  assign n39349 = pi214 & ~n39348;
  assign n39350 = ~n39344 & ~n39349;
  assign n39351 = pi212 & ~n39350;
  assign n39352 = ~pi219 & ~n39335;
  assign n39353 = n37704 & ~n39343;
  assign n39354 = n39352 & ~n39353;
  assign n39355 = ~n39351 & n39354;
  assign n39356 = n39339 & ~n39355;
  assign n39357 = n37664 & ~n39109;
  assign n39358 = pi1147 & ~n39357;
  assign n39359 = ~n39356 & n39358;
  assign n39360 = ~pi1149 & ~n39359;
  assign n39361 = ~pi211 & ~n39343;
  assign n39362 = ~n39335 & ~n39361;
  assign n39363 = pi214 & n39362;
  assign n39364 = ~n39348 & ~n39363;
  assign n39365 = pi212 & ~n39364;
  assign n39366 = ~pi219 & n39365;
  assign n39367 = ~pi299 & n39347;
  assign n39368 = ~pi212 & ~n39272;
  assign n39369 = ~pi219 & ~n39368;
  assign n39370 = ~n39367 & ~n39369;
  assign n39371 = ~po1038 & ~n39370;
  assign n39372 = ~n39366 & n39371;
  assign n39373 = ~n39355 & n39372;
  assign n39374 = ~pi1147 & ~n39117;
  assign n39375 = ~n39373 & n39374;
  assign n39376 = n39360 & ~n39375;
  assign n39377 = ~pi1147 & ~n38858;
  assign n39378 = ~n39372 & n39377;
  assign n39379 = ~n37693 & n39352;
  assign n39380 = n39339 & ~n39379;
  assign n39381 = pi1147 & ~n39380;
  assign n39382 = ~n39083 & n39381;
  assign n39383 = pi1149 & ~n39382;
  assign n39384 = ~n39378 & n39383;
  assign n39385 = ~n39376 & ~n39384;
  assign n39386 = pi1148 & n39385;
  assign n39387 = pi214 & ~n39335;
  assign n39388 = ~n39344 & n39387;
  assign n39389 = ~pi214 & n39362;
  assign n39390 = ~n39388 & ~n39389;
  assign n39391 = pi212 & n39390;
  assign n39392 = ~pi214 & ~n39335;
  assign n39393 = ~pi212 & ~n39392;
  assign n39394 = ~n39362 & n39393;
  assign n39395 = ~pi219 & ~n39394;
  assign n39396 = ~n39391 & n39395;
  assign n39397 = n39339 & ~n39396;
  assign n39398 = n39165 & ~n39397;
  assign n39399 = pi1147 & ~n39398;
  assign n39400 = ~pi1147 & ~po1038;
  assign n39401 = n39367 & n39400;
  assign n39402 = ~pi1147 & n39169;
  assign n39403 = ~n39401 & ~n39402;
  assign n39404 = n39169 & ~n39347;
  assign n39405 = n15973 & n39404;
  assign n39406 = ~n39403 & ~n39405;
  assign n39407 = ~n39399 & ~n39406;
  assign n39408 = pi1149 & ~n39407;
  assign n39409 = n39356 & ~n39396;
  assign n39410 = ~n38861 & ~n39409;
  assign n39411 = pi1147 & ~n39410;
  assign n39412 = ~n39401 & ~n39411;
  assign n39413 = ~pi1149 & ~n39412;
  assign n39414 = ~pi1148 & ~n39413;
  assign n39415 = ~n39408 & n39414;
  assign n39416 = ~n39386 & ~n39415;
  assign n39417 = pi213 & n39416;
  assign n39418 = ~n39217 & ~n39367;
  assign n39419 = ~pi214 & ~n39367;
  assign n39420 = ~pi212 & ~n39419;
  assign n39421 = ~n39418 & n39420;
  assign n39422 = ~pi219 & ~n39421;
  assign n39423 = ~n39261 & ~n39348;
  assign n39424 = pi212 & n39423;
  assign n39425 = n39422 & ~n39424;
  assign n39426 = n39336 & ~n39367;
  assign n39427 = ~n39425 & ~n39426;
  assign n39428 = ~po1038 & n39427;
  assign n39429 = n39242 & ~n39428;
  assign n39430 = ~n38658 & n39344;
  assign n39431 = n39214 & n39342;
  assign n39432 = ~n39353 & ~n39431;
  assign n39433 = ~n39430 & ~n39432;
  assign n39434 = ~n39216 & n39389;
  assign n39435 = ~n39433 & ~n39434;
  assign n39436 = pi212 & n39435;
  assign n39437 = ~n39394 & ~n39436;
  assign n39438 = n39422 & n39437;
  assign n39439 = ~n39337 & ~n39438;
  assign n39440 = ~po1038 & n39439;
  assign n39441 = n39239 & ~n39440;
  assign n39442 = ~n39429 & ~n39441;
  assign n39443 = ~pi213 & n39442;
  assign n39444 = ~pi209 & ~n39443;
  assign n39445 = ~n39417 & n39444;
  assign n39446 = ~n39320 & ~n39445;
  assign n39447 = pi230 & ~n39446;
  assign n39448 = ~pi230 & ~pi240;
  assign po397 = ~n39447 & ~n39448;
  assign n39450 = n38862 & ~n38906;
  assign n39451 = ~pi214 & ~n38922;
  assign n39452 = n38929 & ~n39451;
  assign n39453 = ~pi212 & ~n38923;
  assign n39454 = ~n39452 & ~n39453;
  assign n39455 = ~pi219 & ~n39454;
  assign n39456 = n38173 & ~n38924;
  assign n39457 = ~n39455 & n39456;
  assign n39458 = n38802 & ~n39178;
  assign n39459 = ~n38960 & n39458;
  assign n39460 = ~pi219 & ~n39459;
  assign n39461 = pi1152 & ~n39460;
  assign n39462 = n38963 & n39461;
  assign n39463 = ~n39457 & ~n39462;
  assign n39464 = n39450 & n39463;
  assign n39465 = ~n38787 & n38942;
  assign n39466 = pi219 & ~n38921;
  assign n39467 = n39079 & ~n39466;
  assign n39468 = pi219 & ~n38726;
  assign n39469 = ~po1038 & ~n39468;
  assign n39470 = ~n39467 & ~n39469;
  assign n39471 = ~n38975 & n39470;
  assign n39472 = ~n39465 & ~n39471;
  assign n39473 = pi1152 & n39472;
  assign n39474 = ~pi1151 & ~n38861;
  assign n39475 = ~n38726 & n38942;
  assign n39476 = ~n39470 & ~n39475;
  assign n39477 = ~pi1152 & n39476;
  assign n39478 = n39474 & ~n39477;
  assign n39479 = ~n39473 & n39478;
  assign n39480 = ~pi1150 & ~n39479;
  assign n39481 = ~n39464 & n39480;
  assign n39482 = pi1151 & ~n39083;
  assign n39483 = ~pi299 & ~n38715;
  assign n39484 = ~n38712 & ~n39483;
  assign n39485 = ~pi219 & ~n39484;
  assign n39486 = n39456 & ~n39485;
  assign n39487 = n38731 & n38802;
  assign n39488 = ~pi219 & ~n39487;
  assign n39489 = pi212 & n38802;
  assign n39490 = n39488 & ~n39489;
  assign n39491 = pi1152 & ~n39490;
  assign n39492 = n38963 & n39491;
  assign n39493 = ~n39486 & ~n39492;
  assign n39494 = n39482 & n39493;
  assign n39495 = ~pi1151 & ~n39357;
  assign n39496 = n10468 & n38775;
  assign n39497 = ~n38750 & ~n38926;
  assign n39498 = ~n10468 & ~n38787;
  assign n39499 = ~n39497 & n39498;
  assign n39500 = ~n39496 & ~n39499;
  assign n39501 = ~pi219 & ~n39500;
  assign n39502 = ~n39471 & ~n39501;
  assign n39503 = pi1152 & ~n39502;
  assign n39504 = ~pi299 & n39475;
  assign n39505 = ~n39192 & ~n39504;
  assign n39506 = n39469 & n39505;
  assign n39507 = ~pi1152 & ~n39506;
  assign n39508 = ~n39476 & n39507;
  assign n39509 = ~n39503 & ~n39508;
  assign n39510 = n39495 & ~n39509;
  assign n39511 = pi1150 & ~n39510;
  assign n39512 = ~n39494 & n39511;
  assign n39513 = ~n39481 & ~n39512;
  assign n39514 = pi1149 & n39513;
  assign n39515 = po1038 & ~n39169;
  assign n39516 = pi1151 & ~n39515;
  assign n39517 = n38803 & n38911;
  assign n39518 = n38799 & ~n39517;
  assign n39519 = pi1152 & ~n39518;
  assign n39520 = ~po1038 & ~n39519;
  assign n39521 = n39516 & ~n39520;
  assign n39522 = n38726 & n38737;
  assign n39523 = n38911 & n38921;
  assign n39524 = ~n38711 & ~n39523;
  assign n39525 = n39516 & ~n39524;
  assign n39526 = ~n39522 & ~n39525;
  assign n39527 = ~pi1152 & ~n39526;
  assign n39528 = pi1152 & n38737;
  assign n39529 = n38787 & n39528;
  assign n39530 = ~n39527 & ~n39529;
  assign n39531 = ~n39521 & n39530;
  assign n39532 = ~pi1150 & ~n39531;
  assign n39533 = pi1151 & ~n38858;
  assign n39534 = ~n39111 & ~n39469;
  assign n39535 = ~pi214 & n38703;
  assign n39536 = pi212 & ~n39535;
  assign n39537 = ~n39153 & n39536;
  assign n39538 = n38731 & ~n39151;
  assign n39539 = ~n39537 & ~n39538;
  assign n39540 = ~n39483 & ~n39539;
  assign n39541 = ~pi219 & ~n39540;
  assign n39542 = ~pi1152 & ~n39207;
  assign n39543 = ~n39541 & n39542;
  assign n39544 = ~n39271 & n39488;
  assign n39545 = n39491 & ~n39544;
  assign n39546 = ~n39543 & ~n39545;
  assign n39547 = ~n39534 & ~n39546;
  assign n39548 = n39533 & ~n39547;
  assign n39549 = ~pi1151 & ~n39117;
  assign n39550 = ~n38787 & ~n39505;
  assign n39551 = n38975 & ~n39550;
  assign n39552 = pi1152 & ~n39551;
  assign n39553 = ~n39507 & ~n39552;
  assign n39554 = n39549 & ~n39553;
  assign n39555 = pi1150 & ~n39554;
  assign n39556 = ~n39548 & n39555;
  assign n39557 = ~n39532 & ~n39556;
  assign n39558 = ~pi1149 & n39557;
  assign n39559 = ~pi213 & ~n39558;
  assign n39560 = ~n39514 & n39559;
  assign n39561 = pi213 & ~n38987;
  assign n39562 = pi209 & ~n39561;
  assign n39563 = ~n39560 & n39562;
  assign n39564 = ~n37693 & n39183;
  assign n39565 = ~n37711 & n38859;
  assign n39566 = ~n39564 & ~n39565;
  assign n39567 = ~pi219 & ~n39566;
  assign n39568 = pi219 & n39183;
  assign n39569 = ~po1038 & ~n39568;
  assign n39570 = ~n39567 & n39569;
  assign n39571 = n38883 & ~n39570;
  assign n39572 = ~n39149 & ~n39151;
  assign n39573 = ~pi219 & ~n39572;
  assign n39574 = ~n38713 & n39573;
  assign n39575 = ~n39176 & n39574;
  assign n39576 = n39163 & ~n39575;
  assign n39577 = n38863 & ~n39576;
  assign n39578 = pi1152 & ~n39577;
  assign n39579 = ~n39571 & n39578;
  assign n39580 = pi299 & n38851;
  assign n39581 = n39183 & ~n39523;
  assign n39582 = ~po1038 & ~n39581;
  assign n39583 = ~n39580 & n39582;
  assign n39584 = n38910 & ~n39583;
  assign n39585 = ~n39152 & ~n39156;
  assign n39586 = ~n38705 & ~n38710;
  assign n39587 = ~n39150 & n39586;
  assign n39588 = ~n39585 & ~n39587;
  assign n39589 = ~pi219 & ~n39588;
  assign n39590 = n39163 & ~n39589;
  assign n39591 = n38908 & ~n39590;
  assign n39592 = ~pi1152 & ~n39591;
  assign n39593 = ~n39584 & n39592;
  assign n39594 = ~n39579 & ~n39593;
  assign n39595 = ~pi1150 & n39594;
  assign n39596 = ~pi219 & ~n38110;
  assign n39597 = ~n39176 & n39596;
  assign n39598 = ~pi1153 & n39597;
  assign n39599 = ~pi219 & ~n39175;
  assign n39600 = n39467 & ~n39599;
  assign n39601 = ~n39279 & ~n39600;
  assign n39602 = ~n39598 & ~n39601;
  assign n39603 = n38908 & ~n39602;
  assign n39604 = pi1153 & n39523;
  assign n39605 = n38910 & ~n39604;
  assign n39606 = ~pi1152 & ~n39605;
  assign n39607 = ~pi1151 & ~n39111;
  assign n39608 = ~pi1152 & ~n39607;
  assign n39609 = ~n39606 & ~n39608;
  assign n39610 = ~n39603 & ~n39609;
  assign n39611 = ~po1038 & ~n38794;
  assign n39612 = ~n38728 & ~n38921;
  assign n39613 = n10468 & ~n39612;
  assign n39614 = ~pi299 & ~n38728;
  assign n39615 = ~n37670 & ~n39580;
  assign n39616 = ~n39614 & n39615;
  assign n39617 = ~n39613 & ~n39616;
  assign n39618 = n39290 & n39617;
  assign n39619 = n39611 & ~n39618;
  assign n39620 = n38883 & ~n39619;
  assign n39621 = pi1152 & ~n39620;
  assign n39622 = ~pi211 & n39597;
  assign n39623 = ~n39082 & ~n39622;
  assign n39624 = ~n39602 & ~n39623;
  assign n39625 = n38863 & n39624;
  assign n39626 = n39621 & ~n39625;
  assign n39627 = ~n39610 & ~n39626;
  assign n39628 = pi1150 & n39627;
  assign n39629 = pi1149 & ~n39628;
  assign n39630 = ~n39595 & n39629;
  assign n39631 = ~n38947 & n38978;
  assign n39632 = n39133 & ~n39631;
  assign n39633 = ~pi219 & ~n39632;
  assign n39634 = n39139 & ~n39633;
  assign n39635 = n38883 & ~n39634;
  assign n39636 = pi211 & ~n39091;
  assign n39637 = n38786 & ~n39636;
  assign n39638 = ~pi214 & n39637;
  assign n39639 = n39098 & ~n39638;
  assign n39640 = ~pi219 & ~n39639;
  assign n39641 = ~n39089 & ~n39637;
  assign n39642 = n39640 & ~n39641;
  assign n39643 = n39253 & ~n39642;
  assign n39644 = n39090 & ~n39097;
  assign n39645 = pi214 & n39637;
  assign n39646 = n39089 & ~n39094;
  assign n39647 = pi212 & ~n39646;
  assign n39648 = ~n39645 & n39647;
  assign n39649 = ~pi219 & ~n39648;
  assign n39650 = ~n39644 & n39649;
  assign n39651 = n39253 & ~n39650;
  assign n39652 = ~pi1153 & n39642;
  assign n39653 = n39651 & ~n39652;
  assign n39654 = ~n39643 & ~n39653;
  assign n39655 = n38863 & n39654;
  assign n39656 = pi1152 & ~n39655;
  assign n39657 = ~n39635 & n39656;
  assign n39658 = n38908 & ~n39653;
  assign n39659 = ~po1038 & ~n38762;
  assign n39660 = n38911 & n39127;
  assign n39661 = n39659 & ~n39660;
  assign n39662 = ~n37873 & ~n39661;
  assign n39663 = ~po1038 & n39662;
  assign n39664 = n38910 & ~n39663;
  assign n39665 = ~pi1152 & ~n39664;
  assign n39666 = ~n39658 & n39665;
  assign n39667 = ~n39657 & ~n39666;
  assign n39668 = pi1150 & n39667;
  assign n39669 = ~n38938 & ~n39080;
  assign n39670 = ~n38951 & ~n39669;
  assign n39671 = n38908 & ~n39670;
  assign n39672 = n39606 & ~n39671;
  assign n39673 = pi299 & n38857;
  assign n39674 = ~n38859 & n39673;
  assign n39675 = n38883 & ~n39674;
  assign n39676 = pi1152 & ~n39675;
  assign n39677 = ~n38947 & n39191;
  assign n39678 = ~n39669 & ~n39677;
  assign n39679 = ~n39670 & ~n39678;
  assign n39680 = n38863 & n39679;
  assign n39681 = n39676 & ~n39680;
  assign n39682 = ~pi1150 & ~n39681;
  assign n39683 = ~n39672 & n39682;
  assign n39684 = ~pi1149 & ~n39683;
  assign n39685 = ~n39668 & n39684;
  assign n39686 = ~n39630 & ~n39685;
  assign n39687 = pi213 & ~n39686;
  assign n39688 = ~pi1150 & pi1151;
  assign n39689 = ~n39171 & n39688;
  assign n39690 = ~pi1149 & ~n39689;
  assign n39691 = ~n39140 & n39549;
  assign n39692 = ~n39101 & n39533;
  assign n39693 = ~n39691 & ~n39692;
  assign n39694 = pi1150 & n39693;
  assign n39695 = n39690 & ~n39694;
  assign n39696 = ~n39196 & n39474;
  assign n39697 = ~n39164 & n39450;
  assign n39698 = ~pi1150 & ~n39697;
  assign n39699 = ~n39696 & n39698;
  assign n39700 = ~n39110 & n39607;
  assign n39701 = n39082 & n39482;
  assign n39702 = pi1150 & ~n39701;
  assign n39703 = ~n39700 & n39702;
  assign n39704 = pi1149 & ~n39703;
  assign n39705 = ~n39699 & n39704;
  assign n39706 = ~n39695 & ~n39705;
  assign n39707 = ~pi213 & n39706;
  assign n39708 = ~pi209 & ~n39707;
  assign n39709 = ~n39687 & n39708;
  assign n39710 = ~n39563 & ~n39709;
  assign n39711 = pi230 & ~n39710;
  assign n39712 = ~pi230 & ~pi241;
  assign po398 = ~n39711 & ~n39712;
  assign n39714 = ~pi230 & ~pi242;
  assign n39715 = n37594 & ~n39212;
  assign n39716 = pi214 & ~n38491;
  assign n39717 = ~pi214 & ~n39212;
  assign n39718 = ~n39716 & ~n39717;
  assign n39719 = pi212 & ~n39718;
  assign n39720 = ~pi219 & ~n39719;
  assign n39721 = ~n39715 & n39720;
  assign n39722 = pi219 & ~n37667;
  assign n39723 = ~n37663 & ~n39722;
  assign n39724 = ~n39721 & n39723;
  assign n39725 = po1038 & n39724;
  assign n39726 = pi199 & pi1144;
  assign n39727 = ~pi200 & ~n39726;
  assign n39728 = ~n39321 & n39727;
  assign n39729 = n39329 & ~n39728;
  assign n39730 = n37957 & n39729;
  assign n39731 = ~pi299 & ~n38470;
  assign n39732 = ~n38471 & n39727;
  assign n39733 = n39731 & ~n39732;
  assign n39734 = pi207 & ~n39733;
  assign n39735 = ~pi207 & ~n39729;
  assign n39736 = pi208 & ~n39735;
  assign n39737 = ~n39734 & n39736;
  assign n39738 = ~n39730 & ~n39737;
  assign n39739 = ~n39213 & n39738;
  assign n39740 = ~pi214 & n39739;
  assign n39741 = pi211 & n37893;
  assign n39742 = ~n39204 & n39738;
  assign n39743 = pi214 & n39742;
  assign n39744 = ~n39741 & n39743;
  assign n39745 = ~n39740 & ~n39744;
  assign n39746 = pi212 & n39745;
  assign n39747 = ~pi214 & n39738;
  assign n39748 = ~pi212 & ~n39747;
  assign n39749 = ~n39739 & n39748;
  assign n39750 = ~pi219 & ~n39749;
  assign n39751 = ~n39746 & n39750;
  assign n39752 = ~n39251 & ~n39722;
  assign n39753 = n39738 & ~n39752;
  assign n39754 = ~n39751 & ~n39753;
  assign n39755 = ~po1038 & n39754;
  assign n39756 = ~n39725 & ~n39755;
  assign n39757 = pi213 & n39756;
  assign n39758 = n10468 & ~n37685;
  assign n39759 = ~n37679 & n38157;
  assign n39760 = ~n39758 & ~n39759;
  assign n39761 = n37641 & n39729;
  assign n39762 = ~pi219 & ~n39761;
  assign n39763 = ~n39760 & n39762;
  assign n39764 = n37661 & ~n39730;
  assign n39765 = pi211 & ~n39730;
  assign n39766 = ~n37937 & ~n39761;
  assign n39767 = n37662 & n39766;
  assign n39768 = ~n39765 & ~n39767;
  assign n39769 = pi219 & ~n39768;
  assign n39770 = ~n39764 & ~n39769;
  assign n39771 = ~n39763 & n39770;
  assign n39772 = ~n39737 & ~n39771;
  assign n39773 = ~po1038 & ~n39772;
  assign n39774 = ~pi213 & ~n37677;
  assign n39775 = ~n39773 & n39774;
  assign n39776 = ~n39757 & ~n39775;
  assign n39777 = pi209 & ~n39776;
  assign n39778 = ~pi213 & ~n37700;
  assign n39779 = ~n15973 & ~n39724;
  assign n39780 = pi213 & ~n39779;
  assign n39781 = n15973 & n37643;
  assign n39782 = n39780 & ~n39781;
  assign n39783 = ~pi209 & ~n39782;
  assign n39784 = ~n39778 & n39783;
  assign n39785 = ~n39777 & ~n39784;
  assign n39786 = pi230 & ~n39785;
  assign po399 = ~n39714 & ~n39786;
  assign n39788 = pi253 & pi254;
  assign n39789 = pi267 & n39788;
  assign n39790 = ~pi263 & n39789;
  assign n39791 = ~pi243 & ~pi1091;
  assign n39792 = ~pi299 & pi1091;
  assign n39793 = n37960 & n39792;
  assign n39794 = ~n39791 & ~n39793;
  assign n39795 = pi1156 & ~n39794;
  assign n39796 = pi1156 & ~n37971;
  assign n39797 = pi1091 & ~n38076;
  assign n39798 = n39796 & n39797;
  assign n39799 = ~n39795 & ~n39798;
  assign n39800 = pi243 & ~pi1091;
  assign n39801 = pi1091 & ~n39181;
  assign n39802 = ~n39800 & ~n39801;
  assign n39803 = pi1155 & ~n39800;
  assign n39804 = ~n39791 & ~n39803;
  assign n39805 = n37771 & ~n39804;
  assign n39806 = ~n39802 & ~n39805;
  assign n39807 = ~pi1156 & ~n39806;
  assign n39808 = n39799 & ~n39807;
  assign n39809 = pi1157 & ~n39808;
  assign n39810 = pi199 & pi1091;
  assign n39811 = ~pi299 & n39810;
  assign n39812 = n39803 & ~n39811;
  assign n39813 = pi1156 & ~n39812;
  assign n39814 = ~pi1155 & ~n39800;
  assign n39815 = ~n11221 & n39792;
  assign n39816 = n39814 & ~n39815;
  assign n39817 = n39813 & ~n39816;
  assign n39818 = ~n39797 & ~n39804;
  assign n39819 = ~pi1156 & ~n39818;
  assign n39820 = ~pi1157 & ~n39819;
  assign n39821 = ~n39817 & n39820;
  assign n39822 = ~n39809 & ~n39821;
  assign n39823 = pi211 & ~n39822;
  assign n39824 = pi200 & pi1091;
  assign n39825 = ~pi299 & n39824;
  assign n39826 = n39803 & ~n39825;
  assign n39827 = ~n39802 & ~n39826;
  assign n39828 = ~n39795 & n39827;
  assign n39829 = pi1157 & n39828;
  assign n39830 = pi1091 & ~n11222;
  assign n39831 = n39814 & ~n39830;
  assign n39832 = ~n39812 & ~n39831;
  assign n39833 = pi200 & ~pi1156;
  assign n39834 = n39792 & n39833;
  assign n39835 = ~n39832 & ~n39834;
  assign n39836 = ~pi1157 & ~n39835;
  assign n39837 = ~pi211 & ~n39836;
  assign n39838 = ~n39829 & n39837;
  assign n39839 = ~n39823 & ~n39838;
  assign n39840 = ~pi219 & ~n39839;
  assign n39841 = pi1091 & n37748;
  assign n39842 = n39814 & ~n39841;
  assign n39843 = ~n39826 & ~n39842;
  assign n39844 = ~pi1156 & ~n39843;
  assign n39845 = n37595 & ~n39844;
  assign n39846 = n39799 & n39845;
  assign n39847 = pi299 & pi1091;
  assign n39848 = n39835 & ~n39847;
  assign n39849 = ~pi1157 & ~n39848;
  assign n39850 = pi219 & ~n39849;
  assign n39851 = ~n39846 & n39850;
  assign n39852 = ~n39795 & ~n39807;
  assign n39853 = n38449 & n39852;
  assign n39854 = n39851 & ~n39853;
  assign n39855 = ~n39840 & ~n39854;
  assign n39856 = ~n39790 & ~n39855;
  assign n39857 = ~pi83 & ~pi85;
  assign n39858 = pi314 & ~n39857;
  assign n39859 = pi802 & n39858;
  assign n39860 = pi276 & n39859;
  assign n39861 = ~pi1091 & ~n39860;
  assign n39862 = pi271 & ~n39861;
  assign n39863 = ~pi1091 & ~n39862;
  assign n39864 = pi273 & ~n39863;
  assign n39865 = ~pi1091 & ~n39864;
  assign n39866 = pi299 & n39865;
  assign n39867 = ~pi200 & ~n39865;
  assign n39868 = pi199 & ~n39865;
  assign n39869 = ~pi81 & n39857;
  assign n39870 = pi314 & ~n39869;
  assign n39871 = pi802 & n39870;
  assign n39872 = pi276 & n39871;
  assign n39873 = ~pi1091 & n39872;
  assign n39874 = pi271 & n39873;
  assign n39875 = pi273 & n39874;
  assign n39876 = n39865 & ~n39875;
  assign n39877 = ~pi199 & ~n39876;
  assign n39878 = ~n39868 & ~n39877;
  assign n39879 = n39873 & ~n39878;
  assign n39880 = ~pi299 & ~n39879;
  assign n39881 = ~n39868 & n39880;
  assign n39882 = ~n39867 & n39881;
  assign n39883 = ~n39866 & ~n39882;
  assign n39884 = ~pi243 & n39883;
  assign n39885 = ~pi200 & ~n39873;
  assign n39886 = ~n39878 & ~n39885;
  assign n39887 = ~pi299 & ~n39886;
  assign n39888 = ~n39868 & n39887;
  assign n39889 = ~pi1091 & n39860;
  assign n39890 = pi271 & n39889;
  assign n39891 = pi273 & n39890;
  assign n39892 = pi299 & ~n39891;
  assign n39893 = ~n39867 & n39880;
  assign n39894 = ~n39877 & n39893;
  assign n39895 = ~n39892 & ~n39894;
  assign n39896 = ~n39888 & n39895;
  assign n39897 = pi243 & ~n39896;
  assign n39898 = ~n39884 & ~n39897;
  assign n39899 = ~n39877 & n39887;
  assign n39900 = ~n39866 & ~n39899;
  assign n39901 = ~pi243 & ~n39900;
  assign n39902 = ~pi1155 & ~n39901;
  assign n39903 = n39866 & ~n39875;
  assign n39904 = ~n39887 & ~n39903;
  assign n39905 = ~pi243 & ~n39904;
  assign n39906 = pi1155 & ~n39905;
  assign n39907 = pi243 & n39895;
  assign n39908 = n39906 & ~n39907;
  assign n39909 = ~n39902 & ~n39908;
  assign n39910 = ~n39898 & ~n39909;
  assign n39911 = pi1156 & ~n39910;
  assign n39912 = ~n39892 & ~n39893;
  assign n39913 = pi243 & n39912;
  assign n39914 = ~n39905 & ~n39913;
  assign n39915 = pi1155 & ~n39914;
  assign n39916 = pi243 & ~n39881;
  assign n39917 = n39912 & n39916;
  assign n39918 = ~n39915 & ~n39917;
  assign n39919 = ~n39901 & n39918;
  assign n39920 = ~pi1156 & ~n39919;
  assign n39921 = n38449 & ~n39920;
  assign n39922 = ~n39911 & n39921;
  assign n39923 = ~n39877 & n39880;
  assign n39924 = ~n39892 & ~n39923;
  assign n39925 = pi1155 & n39924;
  assign n39926 = ~n39887 & n39924;
  assign n39927 = ~n39925 & ~n39926;
  assign n39928 = pi243 & ~n39927;
  assign n39929 = pi299 & ~n39875;
  assign n39930 = ~n39893 & ~n39929;
  assign n39931 = ~pi1155 & n39930;
  assign n39932 = ~n39873 & n39931;
  assign n39933 = ~n39866 & ~n39881;
  assign n39934 = ~pi243 & ~n39933;
  assign n39935 = ~n39932 & n39934;
  assign n39936 = ~n39928 & ~n39935;
  assign n39937 = pi1156 & ~n39936;
  assign n39938 = ~n39880 & ~n39892;
  assign n39939 = n39791 & ~n39938;
  assign n39940 = ~pi1155 & ~n39939;
  assign n39941 = pi243 & n39938;
  assign n39942 = n39940 & ~n39941;
  assign n39943 = n39913 & ~n39923;
  assign n39944 = ~n39866 & ~n39888;
  assign n39945 = ~pi243 & ~n39944;
  assign n39946 = pi1155 & ~n39945;
  assign n39947 = ~n39943 & n39946;
  assign n39948 = ~pi1156 & ~n39947;
  assign n39949 = ~n39942 & n39948;
  assign n39950 = ~pi1157 & ~n39949;
  assign n39951 = ~n39937 & n39950;
  assign n39952 = ~n39922 & ~n39951;
  assign n39953 = ~n39887 & ~n39892;
  assign n39954 = n39884 & n39953;
  assign n39955 = ~n39866 & ~n39893;
  assign n39956 = pi243 & ~n39955;
  assign n39957 = ~n39896 & n39956;
  assign n39958 = pi1155 & ~n39957;
  assign n39959 = ~n39954 & n39958;
  assign n39960 = ~n39882 & ~n39929;
  assign n39961 = ~n39800 & ~n39960;
  assign n39962 = ~n39898 & ~n39961;
  assign n39963 = ~n39901 & n39962;
  assign n39964 = ~pi1155 & ~n39963;
  assign n39965 = ~n39959 & ~n39964;
  assign n39966 = pi1156 & ~n39965;
  assign n39967 = ~pi243 & pi1155;
  assign n39968 = n39953 & n39967;
  assign n39969 = ~pi1156 & ~n39968;
  assign n39970 = ~n39892 & ~n39916;
  assign n39971 = n39902 & n39970;
  assign n39972 = ~n39956 & ~n39971;
  assign n39973 = n39969 & n39972;
  assign n39974 = n37595 & ~n39973;
  assign n39975 = ~n39966 & n39974;
  assign n39976 = n39952 & ~n39975;
  assign n39977 = pi219 & ~n39976;
  assign n39978 = ~n39887 & ~n39929;
  assign n39979 = ~n39893 & ~n39903;
  assign n39980 = ~pi1155 & n39979;
  assign n39981 = ~n39978 & n39980;
  assign n39982 = pi1156 & ~n39932;
  assign n39983 = ~n39880 & ~n39929;
  assign n39984 = pi243 & n39983;
  assign n39985 = ~n39881 & ~n39929;
  assign n39986 = ~n39800 & ~n39985;
  assign n39987 = ~n39984 & ~n39986;
  assign n39988 = n39982 & ~n39987;
  assign n39989 = ~n39981 & n39988;
  assign n39990 = ~pi1155 & n39983;
  assign n39991 = ~n39940 & ~n39990;
  assign n39992 = ~n39984 & ~n39991;
  assign n39993 = ~pi1156 & ~n39992;
  assign n39994 = ~pi243 & n39978;
  assign n39995 = pi243 & ~n39979;
  assign n39996 = ~n39994 & ~n39995;
  assign n39997 = ~n39987 & n39996;
  assign n39998 = pi1155 & ~n39997;
  assign n39999 = n39993 & ~n39998;
  assign n40000 = ~pi1157 & ~n39999;
  assign n40001 = ~n39989 & n40000;
  assign n40002 = ~n39902 & ~n39990;
  assign n40003 = ~n39893 & n39985;
  assign n40004 = pi243 & n40003;
  assign n40005 = ~n40002 & ~n40004;
  assign n40006 = ~pi1156 & ~n40005;
  assign n40007 = n39996 & n40006;
  assign n40008 = ~n39894 & ~n39903;
  assign n40009 = pi1155 & n40008;
  assign n40010 = ~n39958 & ~n40009;
  assign n40011 = ~n39882 & n39994;
  assign n40012 = ~n40010 & ~n40011;
  assign n40013 = ~n39882 & ~n39899;
  assign n40014 = ~n39903 & n40013;
  assign n40015 = ~pi243 & ~n40014;
  assign n40016 = ~n39888 & ~n39929;
  assign n40017 = pi243 & ~n39894;
  assign n40018 = n40016 & n40017;
  assign n40019 = ~n40015 & ~n40018;
  assign n40020 = ~pi1155 & ~n40019;
  assign n40021 = ~n40012 & ~n40020;
  assign n40022 = pi1156 & ~n40021;
  assign n40023 = ~n40007 & ~n40022;
  assign n40024 = pi1157 & n40023;
  assign n40025 = ~pi211 & ~n40024;
  assign n40026 = ~n40001 & n40025;
  assign n40027 = pi243 & n39930;
  assign n40028 = n39906 & ~n40027;
  assign n40029 = n40006 & ~n40028;
  assign n40030 = ~n39961 & n40021;
  assign n40031 = pi1156 & ~n40030;
  assign n40032 = ~n40029 & ~n40031;
  assign n40033 = pi1157 & n40032;
  assign n40034 = n39803 & n39868;
  assign n40035 = ~n40028 & ~n40034;
  assign n40036 = n39993 & n40035;
  assign n40037 = ~pi1157 & ~n39988;
  assign n40038 = ~n40036 & n40037;
  assign n40039 = pi211 & ~n40038;
  assign n40040 = ~n40033 & n40039;
  assign n40041 = ~pi219 & ~n40040;
  assign n40042 = ~n40026 & n40041;
  assign n40043 = ~n39977 & ~n40042;
  assign n40044 = n39790 & n40043;
  assign n40045 = ~n39856 & ~n40044;
  assign n40046 = ~po1038 & n40045;
  assign n40047 = pi272 & pi283;
  assign n40048 = pi275 & n40047;
  assign n40049 = pi268 & n40048;
  assign n40050 = ~n37596 & ~n37603;
  assign n40051 = ~pi219 & ~n40050;
  assign n40052 = pi1157 & n10522;
  assign n40053 = ~n40051 & ~n40052;
  assign n40054 = pi1091 & ~n40053;
  assign n40055 = ~n39791 & ~n40054;
  assign n40056 = ~n39790 & ~n40055;
  assign n40057 = po1038 & ~n40056;
  assign n40058 = pi243 & n39891;
  assign n40059 = n37595 & ~n39889;
  assign n40060 = ~n39865 & ~n40059;
  assign n40061 = ~n39800 & ~n40060;
  assign n40062 = ~n40058 & ~n40061;
  assign n40063 = pi219 & ~n40062;
  assign n40064 = ~pi243 & n39875;
  assign n40065 = pi1091 & n40050;
  assign n40066 = pi243 & n39876;
  assign n40067 = ~pi219 & ~n40066;
  assign n40068 = ~n40065 & n40067;
  assign n40069 = ~n40064 & n40068;
  assign n40070 = ~n40063 & ~n40069;
  assign n40071 = n39790 & ~n40070;
  assign n40072 = n40057 & ~n40071;
  assign n40073 = n40049 & ~n40072;
  assign n40074 = ~n40046 & n40073;
  assign n40075 = ~po1038 & n39855;
  assign n40076 = po1038 & n40055;
  assign n40077 = ~n40049 & ~n40076;
  assign n40078 = ~n40075 & n40077;
  assign n40079 = ~pi230 & ~n40078;
  assign n40080 = ~n40074 & n40079;
  assign n40081 = pi199 & ~n38644;
  assign n40082 = n15973 & ~n40081;
  assign n40083 = ~n37959 & ~n39833;
  assign n40084 = n40082 & n40083;
  assign n40085 = ~n15973 & ~n40053;
  assign n40086 = pi230 & ~n40085;
  assign n40087 = ~n40084 & n40086;
  assign po400 = ~n40080 & ~n40087;
  assign n40089 = ~pi230 & ~pi244;
  assign n40090 = ~n39204 & ~n39741;
  assign n40091 = ~n39335 & n40090;
  assign n40092 = ~pi214 & n40091;
  assign n40093 = n37668 & n39272;
  assign n40094 = pi212 & ~n40093;
  assign n40095 = ~n40092 & n40094;
  assign n40096 = ~n39343 & n40095;
  assign n40097 = ~pi219 & ~n40096;
  assign n40098 = n39393 & ~n40091;
  assign n40099 = n40097 & ~n40098;
  assign n40100 = pi1147 & ~n40099;
  assign n40101 = pi299 & n38497;
  assign n40102 = n39339 & ~n40101;
  assign n40103 = n40100 & n40102;
  assign n40104 = ~n39348 & n40095;
  assign n40105 = ~n39348 & n40098;
  assign n40106 = ~pi219 & ~n40105;
  assign n40107 = ~n40104 & n40106;
  assign n40108 = pi219 & ~n38502;
  assign n40109 = ~n39367 & n40108;
  assign n40110 = ~n40107 & ~n40109;
  assign n40111 = n39400 & n40110;
  assign n40112 = ~n38499 & ~n40111;
  assign n40113 = ~n40103 & n40112;
  assign n40114 = ~pi213 & ~n40113;
  assign n40115 = pi213 & n39442;
  assign n40116 = pi209 & ~n40115;
  assign n40117 = ~n40114 & n40116;
  assign n40118 = ~n39239 & ~n39245;
  assign n40119 = ~n10468 & n39293;
  assign n40120 = pi212 & n39214;
  assign n40121 = n39242 & ~n39243;
  assign n40122 = n37930 & ~n40121;
  assign n40123 = ~n40120 & n40122;
  assign n40124 = ~n40119 & n40123;
  assign n40125 = ~n38476 & ~n39308;
  assign n40126 = ~n40124 & n40125;
  assign n40127 = ~po1038 & ~n40126;
  assign n40128 = ~n40118 & ~n40127;
  assign n40129 = pi213 & ~n40128;
  assign n40130 = ~pi213 & ~n38506;
  assign n40131 = ~pi209 & ~n40130;
  assign n40132 = ~n40129 & n40131;
  assign n40133 = ~n40117 & ~n40132;
  assign n40134 = pi230 & ~n40133;
  assign po401 = ~n40089 & ~n40134;
  assign n40136 = pi1146 & n38861;
  assign n40137 = pi1147 & ~n38858;
  assign n40138 = ~n40136 & n40137;
  assign n40139 = n37662 & n39216;
  assign n40140 = pi219 & ~n40139;
  assign n40141 = n39738 & n40140;
  assign n40142 = ~po1038 & ~n40141;
  assign n40143 = ~pi299 & n39738;
  assign n40144 = ~pi214 & n40143;
  assign n40145 = pi212 & ~n40144;
  assign n40146 = ~n38921 & n39738;
  assign n40147 = ~n39216 & n40146;
  assign n40148 = pi214 & n40147;
  assign n40149 = n40145 & ~n40148;
  assign n40150 = n39748 & ~n40143;
  assign n40151 = ~pi219 & ~n40150;
  assign n40152 = ~n40149 & n40151;
  assign n40153 = n40142 & ~n40152;
  assign n40154 = n40138 & ~n40153;
  assign n40155 = ~pi1147 & ~n40136;
  assign n40156 = ~n38906 & n40155;
  assign n40157 = pi214 & ~n39217;
  assign n40158 = n39738 & n40157;
  assign n40159 = pi212 & ~n40158;
  assign n40160 = ~pi214 & n40146;
  assign n40161 = n40159 & ~n40160;
  assign n40162 = n39748 & ~n40146;
  assign n40163 = ~pi219 & ~n40162;
  assign n40164 = ~n40161 & n40163;
  assign n40165 = n40142 & ~n40164;
  assign n40166 = n40156 & ~n40165;
  assign n40167 = pi1148 & ~n40166;
  assign n40168 = ~n40154 & n40167;
  assign n40169 = ~n39747 & n40159;
  assign n40170 = ~pi212 & ~n39738;
  assign n40171 = ~pi219 & ~n40170;
  assign n40172 = ~n40169 & n40171;
  assign n40173 = n40142 & ~n40172;
  assign n40174 = n40155 & ~n40173;
  assign n40175 = ~n39358 & ~n40138;
  assign n40176 = ~n12743 & n39738;
  assign n40177 = ~pi214 & n40176;
  assign n40178 = n40149 & ~n40177;
  assign n40179 = n39748 & ~n40176;
  assign n40180 = ~pi219 & ~n40179;
  assign n40181 = ~n40178 & n40180;
  assign n40182 = n40142 & ~n40181;
  assign n40183 = ~n40175 & ~n40182;
  assign n40184 = ~pi1148 & ~n40183;
  assign n40185 = ~n40174 & n40184;
  assign n40186 = ~n40168 & ~n40185;
  assign n40187 = pi213 & ~n40186;
  assign n40188 = ~pi213 & ~n39756;
  assign n40189 = ~pi209 & ~n40188;
  assign n40190 = ~n40187 & n40189;
  assign n40191 = pi199 & pi1146;
  assign n40192 = ~pi200 & ~n40191;
  assign n40193 = n39323 & ~n40192;
  assign n40194 = ~pi299 & ~n40193;
  assign n40195 = pi1146 & ~n38701;
  assign n40196 = ~n40194 & n40195;
  assign n40197 = ~n38516 & n40196;
  assign n40198 = n37747 & ~n40191;
  assign n40199 = n39323 & ~n40198;
  assign n40200 = n38705 & n40199;
  assign n40201 = ~n40197 & ~n40200;
  assign n40202 = ~pi299 & ~n40201;
  assign n40203 = ~pi214 & ~n40202;
  assign n40204 = ~pi212 & ~n40203;
  assign n40205 = ~n10302 & ~n38705;
  assign n40206 = n40193 & ~n40205;
  assign n40207 = pi211 & ~n40206;
  assign n40208 = ~n40194 & ~n40201;
  assign n40209 = ~pi299 & ~n40208;
  assign n40210 = ~pi211 & n40209;
  assign n40211 = ~n40207 & ~n40210;
  assign n40212 = ~n40202 & ~n40211;
  assign n40213 = n40204 & ~n40212;
  assign n40214 = ~pi219 & ~n40213;
  assign n40215 = n40157 & ~n40202;
  assign n40216 = ~pi214 & n40212;
  assign n40217 = pi212 & ~n40216;
  assign n40218 = ~n40215 & n40217;
  assign n40219 = n40214 & ~n40218;
  assign n40220 = ~n37662 & n40202;
  assign n40221 = pi219 & ~n40220;
  assign n40222 = n37662 & ~n40201;
  assign n40223 = n40221 & ~n40222;
  assign n40224 = ~po1038 & ~n40223;
  assign n40225 = ~n40219 & n40224;
  assign n40226 = n40156 & ~n40225;
  assign n40227 = pi207 & n40199;
  assign n40228 = ~n37957 & ~n40227;
  assign n40229 = n37767 & ~n40228;
  assign n40230 = ~n40198 & n40229;
  assign n40231 = ~pi214 & ~n40230;
  assign n40232 = ~pi212 & ~n40231;
  assign n40233 = ~pi299 & ~n40230;
  assign n40234 = n40232 & ~n40233;
  assign n40235 = ~pi219 & ~n40234;
  assign n40236 = pi212 & ~n40233;
  assign n40237 = ~pi1146 & ~n39271;
  assign n40238 = n40236 & ~n40237;
  assign n40239 = n40235 & ~n40238;
  assign n40240 = n40140 & ~n40230;
  assign n40241 = ~n40239 & ~n40240;
  assign n40242 = ~po1038 & n40241;
  assign n40243 = n40138 & ~n40242;
  assign n40244 = pi1148 & ~n40243;
  assign n40245 = ~n40226 & n40244;
  assign n40246 = ~n10302 & n40192;
  assign n40247 = n40229 & ~n40246;
  assign n40248 = ~n12743 & ~n40247;
  assign n40249 = pi214 & ~n40248;
  assign n40250 = ~pi214 & n40247;
  assign n40251 = ~pi212 & ~n40250;
  assign n40252 = ~n40249 & n40251;
  assign n40253 = ~pi214 & ~n40248;
  assign n40254 = ~pi299 & ~n40247;
  assign n40255 = pi214 & ~n40254;
  assign n40256 = ~n38195 & ~n40233;
  assign n40257 = n40255 & n40256;
  assign n40258 = pi212 & ~n40257;
  assign n40259 = ~n40253 & n40258;
  assign n40260 = ~n40252 & ~n40259;
  assign n40261 = ~pi219 & ~n40260;
  assign n40262 = ~pi1146 & ~n37706;
  assign n40263 = n39176 & ~n40262;
  assign n40264 = n40261 & ~n40263;
  assign n40265 = pi219 & ~n40247;
  assign n40266 = n40140 & n40265;
  assign n40267 = ~n40264 & ~n40266;
  assign n40268 = ~po1038 & n40267;
  assign n40269 = ~n40175 & ~n40268;
  assign n40270 = pi219 & ~n40206;
  assign n40271 = ~n38091 & ~n40270;
  assign n40272 = ~n37661 & ~n40207;
  assign n40273 = n40208 & n40272;
  assign n40274 = ~n40271 & ~n40273;
  assign n40275 = ~po1038 & ~n40274;
  assign n40276 = ~pi219 & ~n39228;
  assign n40277 = ~n39599 & ~n40276;
  assign n40278 = ~n40206 & ~n40277;
  assign n40279 = n40275 & ~n40278;
  assign n40280 = n40155 & ~n40279;
  assign n40281 = ~pi1148 & ~n40280;
  assign n40282 = ~n40269 & n40281;
  assign n40283 = ~n40245 & ~n40282;
  assign n40284 = pi213 & ~n40283;
  assign n40285 = ~pi299 & n40201;
  assign n40286 = n37662 & ~n40285;
  assign n40287 = ~n37900 & n40286;
  assign n40288 = n40221 & ~n40287;
  assign n40289 = n39400 & ~n40288;
  assign n40290 = ~n39213 & ~n40202;
  assign n40291 = n40204 & ~n40290;
  assign n40292 = pi299 & ~n39718;
  assign n40293 = ~n40202 & ~n40292;
  assign n40294 = pi212 & ~n40293;
  assign n40295 = ~pi219 & ~n40294;
  assign n40296 = ~n40291 & n40295;
  assign n40297 = n40289 & ~n40296;
  assign n40298 = pi1147 & ~po1038;
  assign n40299 = ~n39752 & ~n40230;
  assign n40300 = ~n40230 & ~n40292;
  assign n40301 = pi212 & ~n40300;
  assign n40302 = ~pi219 & ~n40301;
  assign n40303 = ~n39261 & n40234;
  assign n40304 = n40302 & ~n40303;
  assign n40305 = ~n40299 & ~n40304;
  assign n40306 = n40298 & n40305;
  assign n40307 = pi1148 & ~n40306;
  assign n40308 = ~n40297 & n40307;
  assign n40309 = ~n39725 & n40308;
  assign n40310 = ~n37661 & ~n37900;
  assign n40311 = n40211 & n40310;
  assign n40312 = ~n40271 & ~n40311;
  assign n40313 = ~pi214 & n40206;
  assign n40314 = pi214 & ~n40209;
  assign n40315 = ~n40290 & n40314;
  assign n40316 = ~n40313 & ~n40315;
  assign n40317 = ~pi212 & ~n40316;
  assign n40318 = ~n40194 & n40294;
  assign n40319 = ~pi219 & ~n40318;
  assign n40320 = ~n40317 & n40319;
  assign n40321 = ~n40312 & ~n40320;
  assign n40322 = n39400 & n40321;
  assign n40323 = n37661 & n40247;
  assign n40324 = ~n40254 & n40301;
  assign n40325 = ~pi219 & ~n40324;
  assign n40326 = n40255 & n40303;
  assign n40327 = n40325 & ~n40326;
  assign n40328 = ~n40265 & ~n40323;
  assign n40329 = ~n39752 & ~n40328;
  assign n40330 = ~n40327 & ~n40329;
  assign n40331 = ~n40323 & ~n40330;
  assign n40332 = n40298 & ~n40331;
  assign n40333 = ~pi1148 & ~n40332;
  assign n40334 = ~n39725 & n40333;
  assign n40335 = ~n40322 & n40334;
  assign n40336 = ~pi213 & ~n40335;
  assign n40337 = ~n40309 & n40336;
  assign n40338 = pi209 & ~n40337;
  assign n40339 = ~n40284 & n40338;
  assign n40340 = ~n40190 & ~n40339;
  assign n40341 = pi230 & ~n40340;
  assign n40342 = ~pi230 & ~pi245;
  assign po402 = ~n40341 & ~n40342;
  assign n40344 = ~n40138 & ~n40156;
  assign n40345 = ~po1038 & ~n40140;
  assign n40346 = ~po1038 & ~n39183;
  assign n40347 = ~n40345 & ~n40346;
  assign n40348 = ~n39184 & ~n39302;
  assign n40349 = n37670 & ~n40348;
  assign n40350 = ~n39564 & ~n40349;
  assign n40351 = ~pi219 & ~n40350;
  assign n40352 = ~n40347 & ~n40351;
  assign n40353 = ~n40344 & ~n40352;
  assign n40354 = ~n38948 & n39269;
  assign n40355 = ~n38729 & ~n39612;
  assign n40356 = ~pi212 & n40355;
  assign n40357 = ~pi219 & ~n40356;
  assign n40358 = ~n40354 & n40357;
  assign n40359 = ~n39185 & ~n40358;
  assign n40360 = n40156 & ~n40359;
  assign n40361 = ~pi1150 & ~n40360;
  assign n40362 = ~n40353 & n40361;
  assign n40363 = ~n39208 & ~n40345;
  assign n40364 = ~n39222 & n39536;
  assign n40365 = ~pi212 & ~n38707;
  assign n40366 = ~pi219 & ~n40365;
  assign n40367 = ~n39189 & n40366;
  assign n40368 = ~n40364 & n40367;
  assign n40369 = ~n40363 & ~n40368;
  assign n40370 = n40138 & ~n40369;
  assign n40371 = n38707 & n40157;
  assign n40372 = ~n39218 & ~n40371;
  assign n40373 = pi212 & n40372;
  assign n40374 = n39155 & ~n40373;
  assign n40375 = ~n40363 & ~n40374;
  assign n40376 = n40156 & ~n40375;
  assign n40377 = pi1150 & ~n40376;
  assign n40378 = ~n40370 & n40377;
  assign n40379 = ~n40362 & ~n40378;
  assign n40380 = pi1148 & ~n40379;
  assign n40381 = n40277 & n40345;
  assign n40382 = pi1150 & n39168;
  assign n40383 = ~n40175 & ~n40345;
  assign n40384 = ~n40155 & ~n40383;
  assign n40385 = ~n40382 & ~n40384;
  assign n40386 = ~n40381 & n40385;
  assign n40387 = pi1150 & n38276;
  assign n40388 = pi299 & n39107;
  assign n40389 = ~pi219 & ~n40388;
  assign n40390 = ~n40387 & n40389;
  assign n40391 = ~n40175 & ~n40263;
  assign n40392 = n40390 & n40391;
  assign n40393 = ~pi1148 & ~n40392;
  assign n40394 = ~n40386 & n40393;
  assign n40395 = ~n40380 & ~n40394;
  assign n40396 = ~pi1149 & ~n40395;
  assign n40397 = ~n39111 & ~n40345;
  assign n40398 = ~n39612 & n40354;
  assign n40399 = n39179 & ~n40398;
  assign n40400 = ~n40156 & ~n40399;
  assign n40401 = ~pi214 & n39612;
  assign n40402 = pi212 & ~n40401;
  assign n40403 = ~n38728 & n40157;
  assign n40404 = n40402 & ~n40403;
  assign n40405 = n40357 & ~n40404;
  assign n40406 = ~n40400 & n40405;
  assign n40407 = ~n40397 & ~n40406;
  assign n40408 = ~n40344 & ~n40407;
  assign n40409 = ~pi1150 & ~n40408;
  assign n40410 = pi1146 & n39080;
  assign n40411 = ~n39277 & ~n40410;
  assign n40412 = n40138 & n40411;
  assign n40413 = n40156 & ~n40381;
  assign n40414 = ~n39279 & n40413;
  assign n40415 = pi1150 & ~n40414;
  assign n40416 = ~n40412 & n40415;
  assign n40417 = pi1148 & ~n40416;
  assign n40418 = ~n40409 & n40417;
  assign n40419 = n39079 & ~n39122;
  assign n40420 = ~n39139 & ~n40419;
  assign n40421 = ~n38762 & n39599;
  assign n40422 = ~n40420 & ~n40421;
  assign n40423 = ~pi1146 & ~n38762;
  assign n40424 = n40422 & ~n40423;
  assign n40425 = n40155 & ~n40424;
  assign n40426 = ~pi1146 & n39138;
  assign n40427 = ~n40420 & ~n40426;
  assign n40428 = n39137 & ~n40277;
  assign n40429 = n40427 & ~n40428;
  assign n40430 = ~n40175 & ~n40429;
  assign n40431 = ~pi1150 & ~n40430;
  assign n40432 = ~n40425 & n40431;
  assign n40433 = ~n39254 & ~n40345;
  assign n40434 = ~n39642 & ~n40433;
  assign n40435 = ~n39100 & ~n39642;
  assign n40436 = ~n39216 & ~n40435;
  assign n40437 = n40434 & ~n40436;
  assign n40438 = ~n40175 & ~n40437;
  assign n40439 = n39651 & n40437;
  assign n40440 = n40155 & ~n40439;
  assign n40441 = pi1150 & ~n40440;
  assign n40442 = ~n40438 & n40441;
  assign n40443 = ~pi1148 & ~n40442;
  assign n40444 = ~n40432 & n40443;
  assign n40445 = pi1149 & ~n40444;
  assign n40446 = ~n40418 & n40445;
  assign n40447 = ~n40396 & ~n40446;
  assign n40448 = ~pi213 & ~n40447;
  assign n40449 = pi1150 & n39084;
  assign n40450 = ~pi1150 & n39112;
  assign n40451 = pi1149 & ~n40450;
  assign n40452 = ~n40449 & n40451;
  assign n40453 = pi1150 & n39165;
  assign n40454 = ~n39164 & n40453;
  assign n40455 = ~pi1149 & pi1150;
  assign n40456 = ~n39198 & ~n40455;
  assign n40457 = ~n40454 & ~n40456;
  assign n40458 = ~n40452 & ~n40457;
  assign n40459 = pi1148 & ~n40458;
  assign n40460 = ~n39171 & n40455;
  assign n40461 = ~pi1150 & ~n39117;
  assign n40462 = ~n39140 & n40461;
  assign n40463 = pi1150 & n39102;
  assign n40464 = pi1149 & ~n40463;
  assign n40465 = ~n40462 & n40464;
  assign n40466 = ~n40460 & ~n40465;
  assign n40467 = ~pi1148 & ~n40466;
  assign n40468 = ~n40459 & ~n40467;
  assign n40469 = pi213 & ~n40468;
  assign n40470 = pi209 & ~n40469;
  assign n40471 = ~n40448 & n40470;
  assign n40472 = n40221 & ~n40286;
  assign n40473 = n39400 & ~n40472;
  assign n40474 = ~n12743 & ~n40206;
  assign n40475 = ~n40202 & n40474;
  assign n40476 = pi214 & n40475;
  assign n40477 = n40217 & ~n40476;
  assign n40478 = n40214 & ~n40477;
  assign n40479 = n40473 & ~n40478;
  assign n40480 = n40232 & n40256;
  assign n40481 = ~n40229 & ~n40259;
  assign n40482 = n40236 & ~n40481;
  assign n40483 = ~pi219 & ~n40482;
  assign n40484 = ~n40480 & n40483;
  assign n40485 = n40298 & ~n40484;
  assign n40486 = n39251 & n40240;
  assign n40487 = n40485 & ~n40486;
  assign n40488 = ~n40479 & ~n40487;
  assign n40489 = n40453 & n40488;
  assign n40490 = n39599 & ~n40202;
  assign n40491 = n40473 & ~n40490;
  assign n40492 = ~pi1150 & ~n40491;
  assign n40493 = ~n12743 & ~n40230;
  assign n40494 = ~pi219 & n40493;
  assign n40495 = n40487 & ~n40494;
  assign n40496 = ~n38861 & ~n40495;
  assign n40497 = n40492 & n40496;
  assign n40498 = ~pi1149 & ~n40497;
  assign n40499 = ~n40489 & n40498;
  assign n40500 = ~n37930 & n40220;
  assign n40501 = n6274 & n40500;
  assign n40502 = n6274 & n40285;
  assign n40503 = ~n37931 & ~n40502;
  assign n40504 = ~pi1147 & ~n40503;
  assign n40505 = ~n40501 & n40504;
  assign n40506 = ~pi57 & ~n40505;
  assign n40507 = pi57 & ~n37931;
  assign n40508 = ~n40506 & ~n40507;
  assign n40509 = ~n6274 & ~n37931;
  assign n40510 = ~pi57 & pi1147;
  assign n40511 = n40235 & ~n40236;
  assign n40512 = n6274 & ~n40486;
  assign n40513 = ~n40511 & n40512;
  assign n40514 = n40510 & ~n40513;
  assign n40515 = ~n40509 & n40514;
  assign n40516 = ~n40508 & ~n40515;
  assign n40517 = pi1150 & ~n40516;
  assign n40518 = ~n39622 & n40513;
  assign n40519 = n40510 & n40518;
  assign n40520 = ~pi1150 & ~n40519;
  assign n40521 = ~n40314 & n40475;
  assign n40522 = pi212 & ~n40521;
  assign n40523 = n40204 & ~n40476;
  assign n40524 = ~pi219 & ~n40523;
  assign n40525 = ~n40522 & n40524;
  assign n40526 = n40473 & ~n40525;
  assign n40527 = ~n39357 & ~n40526;
  assign n40528 = n40520 & n40527;
  assign n40529 = pi1149 & ~n40528;
  assign n40530 = ~n40517 & n40529;
  assign n40531 = ~n40499 & ~n40530;
  assign n40532 = pi1148 & n40531;
  assign n40533 = ~pi212 & ~n40313;
  assign n40534 = pi214 & ~n40474;
  assign n40535 = n40533 & ~n40534;
  assign n40536 = ~pi214 & ~n40474;
  assign n40537 = pi214 & n40211;
  assign n40538 = pi212 & ~n40537;
  assign n40539 = ~n40536 & n40538;
  assign n40540 = ~n40535 & ~n40539;
  assign n40541 = ~pi219 & ~n40540;
  assign n40542 = ~n40270 & ~n40541;
  assign n40543 = n39400 & n40542;
  assign n40544 = ~n40261 & ~n40265;
  assign n40545 = n40298 & n40544;
  assign n40546 = n40461 & ~n40545;
  assign n40547 = ~n40543 & n40546;
  assign n40548 = ~n40314 & n40533;
  assign n40549 = ~pi214 & ~n40209;
  assign n40550 = n40538 & ~n40549;
  assign n40551 = ~n40548 & ~n40550;
  assign n40552 = ~pi219 & ~n40551;
  assign n40553 = ~n40270 & ~n40552;
  assign n40554 = ~pi1147 & ~n40553;
  assign n40555 = ~n39267 & ~n39276;
  assign n40556 = ~n40254 & n40555;
  assign n40557 = pi1147 & ~n40556;
  assign n40558 = ~n40554 & ~n40557;
  assign n40559 = ~po1038 & n40558;
  assign n40560 = ~n38858 & ~n40559;
  assign n40561 = pi1150 & n40560;
  assign n40562 = ~n40547 & ~n40561;
  assign n40563 = pi1149 & ~n40562;
  assign n40564 = pi1150 & n39169;
  assign n40565 = ~pi1147 & n40208;
  assign n40566 = n15973 & ~n40565;
  assign n40567 = n40564 & ~n40566;
  assign n40568 = pi1147 & ~n40247;
  assign n40569 = n40206 & ~n40564;
  assign n40570 = ~pi1147 & ~n40569;
  assign n40571 = ~n40568 & ~n40570;
  assign n40572 = ~po1038 & n40571;
  assign n40573 = ~pi1149 & ~n40572;
  assign n40574 = ~n40567 & n40573;
  assign n40575 = ~n40563 & ~n40574;
  assign n40576 = ~pi1148 & ~n40575;
  assign n40577 = ~n40532 & ~n40576;
  assign n40578 = pi213 & n40577;
  assign n40579 = ~pi213 & ~n40283;
  assign n40580 = ~pi209 & ~n40579;
  assign n40581 = ~n40578 & n40580;
  assign n40582 = ~n40471 & ~n40581;
  assign n40583 = pi230 & ~n40582;
  assign n40584 = ~pi230 & ~pi246;
  assign po403 = ~n40583 & ~n40584;
  assign n40586 = pi212 & ~n38703;
  assign n40587 = n40367 & ~n40586;
  assign n40588 = n39163 & ~n40587;
  assign n40589 = n39482 & ~n40588;
  assign n40590 = pi1147 & ~n40589;
  assign n40591 = ~pi1151 & ~n39083;
  assign n40592 = ~n39184 & n39569;
  assign n40593 = n37670 & ~n40355;
  assign n40594 = n40592 & ~n40593;
  assign n40595 = n40591 & ~n40594;
  assign n40596 = ~n39195 & n40595;
  assign n40597 = n40590 & ~n40596;
  assign n40598 = pi1149 & ~n40597;
  assign n40599 = ~pi1151 & ~n38858;
  assign n40600 = ~n40594 & n40599;
  assign n40601 = ~n39537 & n40367;
  assign n40602 = n39208 & ~n40601;
  assign n40603 = ~n38858 & ~n40602;
  assign n40604 = pi1151 & n40603;
  assign n40605 = ~pi1147 & ~n40604;
  assign n40606 = ~n40600 & n40605;
  assign n40607 = n40598 & ~n40606;
  assign n40608 = ~pi219 & ~n15973;
  assign n40609 = ~n39116 & n40608;
  assign n40610 = ~pi1151 & ~n40609;
  assign n40611 = ~pi1147 & ~n40610;
  assign n40612 = pi1151 & ~n39117;
  assign n40613 = ~n39193 & n40612;
  assign n40614 = n40611 & ~n40613;
  assign n40615 = pi1151 & ~n39357;
  assign n40616 = ~n39678 & n40615;
  assign n40617 = ~pi1151 & ~n39110;
  assign n40618 = ~n40616 & ~n40617;
  assign n40619 = pi1147 & n40618;
  assign n40620 = ~pi1149 & ~n40619;
  assign n40621 = ~n40614 & n40620;
  assign n40622 = ~pi1150 & ~n40621;
  assign n40623 = ~n40607 & n40622;
  assign n40624 = pi1147 & ~n39701;
  assign n40625 = n39105 & n39607;
  assign n40626 = n40624 & ~n40625;
  assign n40627 = n40357 & ~n40398;
  assign n40628 = n39611 & ~n40627;
  assign n40629 = ~n39180 & n39611;
  assign n40630 = ~n40628 & ~n40629;
  assign n40631 = n40599 & n40630;
  assign n40632 = ~n39277 & n39533;
  assign n40633 = ~pi1147 & ~n40632;
  assign n40634 = ~n40631 & n40633;
  assign n40635 = pi1149 & ~n40634;
  assign n40636 = ~n40626 & n40635;
  assign n40637 = ~pi1147 & ~n39691;
  assign n40638 = ~n39088 & n40435;
  assign n40639 = n40612 & ~n40638;
  assign n40640 = n40637 & ~n40639;
  assign n40641 = ~n39643 & n40615;
  assign n40642 = n39121 & ~n39135;
  assign n40643 = ~n40420 & ~n40642;
  assign n40644 = ~n39357 & ~n40643;
  assign n40645 = ~pi1151 & n40644;
  assign n40646 = ~n40641 & ~n40645;
  assign n40647 = pi1147 & n40646;
  assign n40648 = ~pi1149 & ~n40647;
  assign n40649 = ~n40640 & n40648;
  assign n40650 = pi1150 & ~n40649;
  assign n40651 = ~n40636 & n40650;
  assign n40652 = ~n40623 & ~n40651;
  assign n40653 = pi1148 & ~n40652;
  assign n40654 = pi1147 & ~n39697;
  assign n40655 = ~n38906 & n39474;
  assign n40656 = ~n39195 & n40655;
  assign n40657 = n40654 & ~n40656;
  assign n40658 = ~pi1150 & ~n40657;
  assign n40659 = ~pi1151 & ~n38906;
  assign n40660 = ~n39582 & n40659;
  assign n40661 = ~n39158 & n39208;
  assign n40662 = ~n38906 & ~n40661;
  assign n40663 = pi1151 & n40662;
  assign n40664 = ~pi1147 & ~n40663;
  assign n40665 = ~n40660 & n40664;
  assign n40666 = n40658 & ~n40665;
  assign n40667 = n39450 & n39601;
  assign n40668 = pi1147 & ~n40667;
  assign n40669 = ~n39194 & n40655;
  assign n40670 = n40668 & ~n40669;
  assign n40671 = pi1150 & ~n40670;
  assign n40672 = ~n40628 & n40659;
  assign n40673 = pi1151 & ~n38906;
  assign n40674 = ~n39279 & n40673;
  assign n40675 = ~pi1147 & ~n40674;
  assign n40676 = ~n40672 & n40675;
  assign n40677 = n40671 & ~n40676;
  assign n40678 = ~n40666 & ~n40677;
  assign n40679 = pi1149 & ~n40678;
  assign n40680 = ~pi1151 & ~n39286;
  assign n40681 = ~pi1147 & ~n40680;
  assign n40682 = pi1151 & ~n39087;
  assign n40683 = n40681 & ~n40682;
  assign n40684 = pi1150 & ~n40683;
  assign n40685 = n39643 & ~n39650;
  assign n40686 = n38862 & ~n40685;
  assign n40687 = ~n38861 & ~n40422;
  assign n40688 = ~pi1151 & n40687;
  assign n40689 = ~n40686 & ~n40688;
  assign n40690 = pi1147 & n40689;
  assign n40691 = n40684 & ~n40690;
  assign n40692 = ~pi1147 & pi1151;
  assign n40693 = n39168 & n40692;
  assign n40694 = ~pi1150 & ~n40693;
  assign n40695 = ~n38276 & n39599;
  assign n40696 = ~n39669 & ~n40695;
  assign n40697 = n38862 & ~n40696;
  assign n40698 = n39474 & ~n39600;
  assign n40699 = ~n40697 & ~n40698;
  assign n40700 = pi1147 & n40699;
  assign n40701 = n40694 & ~n40700;
  assign n40702 = ~n40691 & ~n40701;
  assign n40703 = ~pi1149 & ~n40702;
  assign n40704 = ~pi1148 & ~n40703;
  assign n40705 = ~n40679 & n40704;
  assign n40706 = ~n40653 & ~n40705;
  assign n40707 = ~pi213 & ~n40706;
  assign n40708 = pi213 & n39706;
  assign n40709 = pi209 & ~n40708;
  assign n40710 = ~n40707 & n40709;
  assign n40711 = ~n39515 & ~n39661;
  assign n40712 = n40681 & n40711;
  assign n40713 = ~pi1150 & ~n40712;
  assign n40714 = ~n40628 & n40673;
  assign n40715 = ~n39607 & ~n40714;
  assign n40716 = pi1147 & n40715;
  assign n40717 = n40713 & ~n40716;
  assign n40718 = n39133 & n39139;
  assign n40719 = n39533 & ~n40718;
  assign n40720 = n40637 & ~n40719;
  assign n40721 = pi1150 & ~n40720;
  assign n40722 = n39533 & n40630;
  assign n40723 = n39549 & ~n40629;
  assign n40724 = ~n40722 & ~n40723;
  assign n40725 = pi1147 & n40724;
  assign n40726 = n40721 & ~n40725;
  assign n40727 = ~n40717 & ~n40726;
  assign n40728 = ~pi1149 & ~n40727;
  assign n40729 = ~n39081 & n40698;
  assign n40730 = n40668 & ~n40729;
  assign n40731 = ~pi1150 & ~n40730;
  assign n40732 = n39474 & ~n40685;
  assign n40733 = n39165 & ~n39651;
  assign n40734 = ~pi1147 & ~n40733;
  assign n40735 = ~n40732 & n40734;
  assign n40736 = n40731 & ~n40735;
  assign n40737 = ~n39357 & ~n39623;
  assign n40738 = ~pi1151 & n40737;
  assign n40739 = n40624 & ~n40738;
  assign n40740 = pi1150 & ~n40739;
  assign n40741 = n39495 & ~n39643;
  assign n40742 = n39105 & n40682;
  assign n40743 = ~pi1147 & ~n40742;
  assign n40744 = ~n40741 & n40743;
  assign n40745 = n40740 & ~n40744;
  assign n40746 = ~n40736 & ~n40745;
  assign n40747 = pi1149 & ~n40746;
  assign n40748 = pi1148 & ~n40747;
  assign n40749 = ~n40728 & n40748;
  assign n40750 = ~n38947 & n39573;
  assign n40751 = n39163 & ~n40750;
  assign n40752 = ~n39159 & n40751;
  assign n40753 = n39474 & ~n40752;
  assign n40754 = n40654 & ~n40753;
  assign n40755 = ~pi1150 & ~n40754;
  assign n40756 = ~n10468 & n38939;
  assign n40757 = ~n40696 & ~n40756;
  assign n40758 = n39450 & n40757;
  assign n40759 = n39474 & ~n40696;
  assign n40760 = ~pi1147 & ~n40759;
  assign n40761 = ~n40758 & n40760;
  assign n40762 = n40755 & ~n40761;
  assign n40763 = ~n39357 & ~n40751;
  assign n40764 = ~pi1151 & n40763;
  assign n40765 = n40590 & ~n40764;
  assign n40766 = pi1150 & ~n40765;
  assign n40767 = n39495 & ~n39678;
  assign n40768 = ~n38939 & n39482;
  assign n40769 = ~n39678 & n40768;
  assign n40770 = ~pi1147 & ~n40769;
  assign n40771 = ~n40767 & n40770;
  assign n40772 = n40766 & ~n40771;
  assign n40773 = ~n40762 & ~n40772;
  assign n40774 = pi1149 & ~n40773;
  assign n40775 = ~n15973 & n38857;
  assign n40776 = pi1151 & ~n40775;
  assign n40777 = n40611 & ~n40776;
  assign n40778 = pi1150 & ~n40777;
  assign n40779 = n39533 & ~n40594;
  assign n40780 = n39186 & n39569;
  assign n40781 = ~n39117 & ~n40780;
  assign n40782 = ~pi1151 & n40781;
  assign n40783 = ~n40779 & ~n40782;
  assign n40784 = pi1147 & n40783;
  assign n40785 = n40778 & ~n40784;
  assign n40786 = n39170 & n40692;
  assign n40787 = ~pi1150 & ~n40786;
  assign n40788 = ~n38906 & ~n39582;
  assign n40789 = ~pi1151 & ~n40346;
  assign n40790 = ~n40788 & ~n40789;
  assign n40791 = pi1147 & n40790;
  assign n40792 = n40787 & ~n40791;
  assign n40793 = ~n40785 & ~n40792;
  assign n40794 = ~pi1149 & ~n40793;
  assign n40795 = ~pi1148 & ~n40794;
  assign n40796 = ~n40774 & n40795;
  assign n40797 = ~n40749 & ~n40796;
  assign n40798 = pi213 & ~n40797;
  assign n40799 = ~pi213 & ~n39202;
  assign n40800 = ~pi209 & ~n40799;
  assign n40801 = ~n40798 & n40800;
  assign n40802 = ~n40710 & ~n40801;
  assign n40803 = pi230 & ~n40802;
  assign n40804 = ~pi230 & ~pi247;
  assign po404 = ~n40803 & ~n40804;
  assign n40806 = pi1152 & ~n39701;
  assign n40807 = ~n40588 & n40591;
  assign n40808 = n40806 & ~n40807;
  assign n40809 = pi1150 & ~n40808;
  assign n40810 = pi1151 & ~n39111;
  assign n40811 = n39105 & n40810;
  assign n40812 = ~pi1152 & ~n40811;
  assign n40813 = ~n40596 & n40812;
  assign n40814 = n40809 & ~n40813;
  assign n40815 = ~pi1152 & ~n40617;
  assign n40816 = pi1151 & n40644;
  assign n40817 = n40815 & ~n40816;
  assign n40818 = ~n40641 & ~n40767;
  assign n40819 = pi1152 & n40818;
  assign n40820 = ~pi1150 & ~n40819;
  assign n40821 = ~n40817 & n40820;
  assign n40822 = pi1148 & ~n40821;
  assign n40823 = ~n40814 & n40822;
  assign n40824 = ~pi1151 & n40603;
  assign n40825 = ~n40632 & ~n40824;
  assign n40826 = pi1152 & n40825;
  assign n40827 = ~pi1152 & ~n40600;
  assign n40828 = ~n40722 & n40827;
  assign n40829 = pi1150 & ~n40828;
  assign n40830 = ~n40826 & n40829;
  assign n40831 = ~n39140 & n40612;
  assign n40832 = ~pi1152 & ~n40831;
  assign n40833 = ~n40610 & n40832;
  assign n40834 = ~n39193 & n39549;
  assign n40835 = ~n40639 & ~n40834;
  assign n40836 = pi1152 & n40835;
  assign n40837 = ~pi1150 & ~n40836;
  assign n40838 = ~n40833 & n40837;
  assign n40839 = ~pi1148 & ~n40838;
  assign n40840 = ~n40830 & n40839;
  assign n40841 = ~n40823 & ~n40840;
  assign n40842 = pi1149 & ~n40841;
  assign n40843 = ~n39164 & n40655;
  assign n40844 = pi1152 & ~n40843;
  assign n40845 = ~n40667 & n40844;
  assign n40846 = n39165 & ~n39194;
  assign n40847 = ~pi1152 & ~n40846;
  assign n40848 = ~n40656 & n40847;
  assign n40849 = ~n40845 & ~n40848;
  assign n40850 = pi1150 & ~n40849;
  assign n40851 = ~n40687 & ~n40698;
  assign n40852 = ~pi1152 & ~n40851;
  assign n40853 = ~n40686 & ~n40759;
  assign n40854 = pi1152 & ~n40853;
  assign n40855 = ~pi1150 & ~n40854;
  assign n40856 = ~n40852 & n40855;
  assign n40857 = ~n40850 & ~n40856;
  assign n40858 = pi1148 & n40857;
  assign n40859 = ~pi1151 & n40662;
  assign n40860 = ~n40674 & ~n40859;
  assign n40861 = pi1152 & n40860;
  assign n40862 = ~pi1152 & ~n40714;
  assign n40863 = ~n40660 & n40862;
  assign n40864 = pi1150 & ~n40863;
  assign n40865 = ~n40861 & n40864;
  assign n40866 = pi1151 & ~pi1152;
  assign n40867 = n39286 & n40866;
  assign n40868 = ~pi1150 & ~n40867;
  assign n40869 = ~pi1151 & ~n39168;
  assign n40870 = ~n40682 & ~n40869;
  assign n40871 = pi1152 & n40870;
  assign n40872 = n40868 & ~n40871;
  assign n40873 = ~n40865 & ~n40872;
  assign n40874 = ~pi1148 & ~n40873;
  assign n40875 = ~pi1149 & ~n40874;
  assign n40876 = ~n40858 & n40875;
  assign n40877 = ~n40842 & ~n40876;
  assign n40878 = ~pi213 & ~n40877;
  assign n40879 = ~n39141 & n40866;
  assign n40880 = ~pi1150 & ~n40879;
  assign n40881 = ~pi1151 & ~n39170;
  assign n40882 = ~n39168 & n40881;
  assign n40883 = ~n39692 & ~n40882;
  assign n40884 = pi1152 & n40883;
  assign n40885 = n40880 & ~n40884;
  assign n40886 = ~n39701 & n40844;
  assign n40887 = pi1151 & n39112;
  assign n40888 = ~pi1152 & ~n39696;
  assign n40889 = ~n40887 & n40888;
  assign n40890 = pi1150 & ~n40889;
  assign n40891 = ~n40886 & n40890;
  assign n40892 = ~n40885 & ~n40891;
  assign n40893 = pi213 & n40892;
  assign n40894 = pi209 & ~n40893;
  assign n40895 = ~n40878 & n40894;
  assign n40896 = ~n40589 & n40844;
  assign n40897 = pi1150 & ~n40896;
  assign n40898 = pi1151 & n40763;
  assign n40899 = ~pi1152 & ~n40898;
  assign n40900 = ~n40753 & n40899;
  assign n40901 = n40897 & ~n40900;
  assign n40902 = ~pi1152 & ~n40789;
  assign n40903 = pi1151 & n40781;
  assign n40904 = n40902 & ~n40903;
  assign n40905 = ~n40660 & ~n40779;
  assign n40906 = pi1152 & n40905;
  assign n40907 = ~pi1150 & ~n40906;
  assign n40908 = ~n40904 & n40907;
  assign n40909 = ~n40901 & ~n40908;
  assign n40910 = ~pi1149 & n40909;
  assign n40911 = n40612 & ~n40629;
  assign n40912 = n39608 & ~n40911;
  assign n40913 = ~pi1150 & ~n40912;
  assign n40914 = ~n40672 & ~n40722;
  assign n40915 = pi1152 & n40914;
  assign n40916 = n40913 & ~n40915;
  assign n40917 = pi1151 & n40737;
  assign n40918 = ~pi1152 & ~n40917;
  assign n40919 = ~n40729 & n40918;
  assign n40920 = n39601 & n40655;
  assign n40921 = n40806 & ~n40920;
  assign n40922 = pi1150 & ~n40921;
  assign n40923 = ~n40919 & n40922;
  assign n40924 = ~n40916 & ~n40923;
  assign n40925 = pi1149 & n40924;
  assign n40926 = pi1148 & ~n40925;
  assign n40927 = ~n40910 & n40926;
  assign n40928 = ~n39651 & n40655;
  assign n40929 = ~n40742 & ~n40928;
  assign n40930 = pi1152 & n40929;
  assign n40931 = ~pi1152 & ~n40641;
  assign n40932 = ~n40732 & n40931;
  assign n40933 = pi1150 & ~n40932;
  assign n40934 = ~n40930 & n40933;
  assign n40935 = ~n40680 & n40832;
  assign n40936 = ~pi1151 & ~n40711;
  assign n40937 = ~n40719 & ~n40936;
  assign n40938 = pi1152 & n40937;
  assign n40939 = ~pi1150 & ~n40938;
  assign n40940 = ~n40935 & n40939;
  assign n40941 = pi1149 & ~n40940;
  assign n40942 = ~n40934 & n40941;
  assign n40943 = n40655 & n40757;
  assign n40944 = ~n40769 & ~n40943;
  assign n40945 = pi1152 & n40944;
  assign n40946 = ~pi1152 & ~n40616;
  assign n40947 = ~n40759 & n40946;
  assign n40948 = pi1150 & ~n40947;
  assign n40949 = ~n40945 & n40948;
  assign n40950 = ~n40776 & ~n40881;
  assign n40951 = pi1152 & n40950;
  assign n40952 = n40609 & n40866;
  assign n40953 = ~pi1150 & ~n40952;
  assign n40954 = ~n40951 & n40953;
  assign n40955 = ~pi1149 & ~n40954;
  assign n40956 = ~n40949 & n40955;
  assign n40957 = ~n40942 & ~n40956;
  assign n40958 = ~pi1148 & n40957;
  assign n40959 = ~n40927 & ~n40958;
  assign n40960 = pi213 & n40959;
  assign n40961 = ~pi213 & ~n40468;
  assign n40962 = ~pi209 & ~n40961;
  assign n40963 = ~n40960 & n40962;
  assign n40964 = ~n40895 & ~n40963;
  assign n40965 = pi230 & ~n40964;
  assign n40966 = ~pi230 & ~pi248;
  assign po405 = ~n40965 & ~n40966;
  assign n40968 = ~pi213 & n40892;
  assign n40969 = pi299 & n38007;
  assign n40970 = ~n39614 & ~n40969;
  assign n40971 = ~pi214 & ~n40970;
  assign n40972 = ~n38788 & n38965;
  assign n40973 = ~n40971 & ~n40972;
  assign n40974 = pi212 & n40973;
  assign n40975 = ~pi219 & ~n40974;
  assign n40976 = n38731 & n40970;
  assign n40977 = n40975 & ~n40976;
  assign n40978 = ~n38794 & ~n40977;
  assign n40979 = n6274 & n40978;
  assign n40980 = ~pi57 & pi1151;
  assign n40981 = ~n6274 & n38010;
  assign n40982 = n40980 & ~n40981;
  assign n40983 = ~n40979 & n40982;
  assign n40984 = pi57 & ~n38010;
  assign n40985 = ~n39184 & ~n40969;
  assign n40986 = ~n38729 & n40985;
  assign n40987 = ~pi212 & ~n40986;
  assign n40988 = ~pi214 & n40985;
  assign n40989 = pi212 & ~n40988;
  assign n40990 = ~n38921 & n39183;
  assign n40991 = ~n39580 & ~n40990;
  assign n40992 = pi214 & n40991;
  assign n40993 = n40989 & ~n40992;
  assign n40994 = ~n40987 & ~n40993;
  assign n40995 = ~pi219 & ~n40994;
  assign n40996 = ~n39568 & ~n40995;
  assign n40997 = n6274 & n40996;
  assign n40998 = ~pi57 & ~pi1151;
  assign n40999 = ~n40981 & n40998;
  assign n41000 = ~n40997 & n40999;
  assign n41001 = ~n40984 & ~n41000;
  assign n41002 = ~n40983 & n41001;
  assign n41003 = ~pi1152 & ~n41002;
  assign n41004 = ~n38703 & ~n40969;
  assign n41005 = ~pi214 & ~n41004;
  assign n41006 = ~n38703 & ~n39580;
  assign n41007 = pi214 & ~n41006;
  assign n41008 = ~n41005 & ~n41007;
  assign n41009 = pi212 & n41008;
  assign n41010 = n39189 & ~n40969;
  assign n41011 = n40366 & ~n41010;
  assign n41012 = ~n41009 & n41011;
  assign n41013 = ~n39162 & ~n41012;
  assign n41014 = n38737 & n41013;
  assign n41015 = ~n39268 & ~n39467;
  assign n41016 = pi299 & ~n38007;
  assign n41017 = ~n10468 & n41016;
  assign n41018 = ~n38041 & ~n41017;
  assign n41019 = n37693 & ~n41018;
  assign n41020 = n39596 & ~n41019;
  assign n41021 = pi1151 & ~n41020;
  assign n41022 = ~n41015 & n41021;
  assign n41023 = n38046 & ~n41022;
  assign n41024 = ~n41014 & n41023;
  assign n41025 = pi1150 & ~n41024;
  assign n41026 = ~n41003 & n41025;
  assign n41027 = ~pi1151 & n40696;
  assign n41028 = ~n38788 & ~n41017;
  assign n41029 = n38009 & n38737;
  assign n41030 = ~n41028 & n41029;
  assign n41031 = ~n11164 & n37759;
  assign n41032 = ~n38771 & ~n41031;
  assign n41033 = ~pi211 & ~n41032;
  assign n41034 = ~n37873 & n41033;
  assign n41035 = ~n39636 & ~n41034;
  assign n41036 = pi214 & n41035;
  assign n41037 = n39089 & ~n41016;
  assign n41038 = ~n41036 & ~n41037;
  assign n41039 = pi212 & n41038;
  assign n41040 = ~n41010 & ~n41039;
  assign n41041 = n39258 & n41040;
  assign n41042 = pi1151 & ~n41041;
  assign n41043 = n39253 & n41042;
  assign n41044 = n38046 & ~n41043;
  assign n41045 = ~n41030 & n41044;
  assign n41046 = ~n41027 & n41045;
  assign n41047 = ~pi1150 & ~n41046;
  assign n41048 = ~n37873 & ~n39122;
  assign n41049 = pi211 & n41048;
  assign n41050 = ~n37670 & ~n41049;
  assign n41051 = ~n37809 & n39127;
  assign n41052 = n41050 & ~n41051;
  assign n41053 = n38166 & ~n38762;
  assign n41054 = n37918 & ~n41048;
  assign n41055 = ~n41053 & ~n41054;
  assign n41056 = ~n41052 & n41055;
  assign n41057 = ~pi219 & ~n41056;
  assign n41058 = pi1151 & ~n41057;
  assign n41059 = n39139 & n41058;
  assign n41060 = ~n41030 & ~n41059;
  assign n41061 = n38012 & n41060;
  assign n41062 = n41047 & ~n41061;
  assign n41063 = ~n41026 & ~n41062;
  assign n41064 = pi213 & ~n41063;
  assign n41065 = ~pi209 & ~n41064;
  assign n41066 = ~n40968 & n41065;
  assign n41067 = ~n37704 & ~n38138;
  assign n41068 = pi211 & ~n38153;
  assign n41069 = pi214 & n41068;
  assign n41070 = ~n41067 & ~n41069;
  assign n41071 = ~pi212 & ~n41070;
  assign n41072 = ~pi219 & ~n41071;
  assign n41073 = pi214 & n38153;
  assign n41074 = ~pi211 & ~n38138;
  assign n41075 = ~pi214 & ~n41074;
  assign n41076 = ~n41068 & n41075;
  assign n41077 = pi212 & ~n41076;
  assign n41078 = ~n41073 & n41077;
  assign n41079 = n41072 & ~n41078;
  assign n41080 = ~pi211 & n38153;
  assign n41081 = ~n38188 & ~n41080;
  assign n41082 = ~n37661 & n41081;
  assign n41083 = ~n38174 & ~n41082;
  assign n41084 = pi219 & n41083;
  assign n41085 = ~po1038 & ~n41084;
  assign n41086 = ~n41079 & n41085;
  assign n41087 = n40615 & ~n41086;
  assign n41088 = pi212 & ~n41070;
  assign n41089 = ~pi212 & ~n38138;
  assign n41090 = ~pi219 & ~n41089;
  assign n41091 = ~n41088 & n41090;
  assign n41092 = n41085 & ~n41091;
  assign n41093 = n39474 & ~n41092;
  assign n41094 = ~pi1152 & ~n41093;
  assign n41095 = ~n41087 & n41094;
  assign n41096 = pi214 & n38089;
  assign n41097 = ~n38096 & ~n41096;
  assign n41098 = ~pi212 & ~n41097;
  assign n41099 = ~pi214 & ~n38089;
  assign n41100 = ~pi211 & n38087;
  assign n41101 = ~n38120 & ~n41100;
  assign n41102 = pi214 & ~n41101;
  assign n41103 = pi212 & ~n41102;
  assign n41104 = ~n41099 & n41103;
  assign n41105 = ~n41098 & ~n41104;
  assign n41106 = ~pi219 & ~n41105;
  assign n41107 = n38095 & ~n41106;
  assign n41108 = n40655 & ~n41107;
  assign n41109 = pi214 & n38074;
  assign n41110 = n38097 & ~n41109;
  assign n41111 = ~pi219 & ~n41110;
  assign n41112 = pi212 & ~n38074;
  assign n41113 = n41111 & ~n41112;
  assign n41114 = n38095 & ~n41113;
  assign n41115 = n39482 & ~n41114;
  assign n41116 = pi1152 & ~n41115;
  assign n41117 = ~n41108 & n41116;
  assign n41118 = ~n41095 & ~n41117;
  assign n41119 = pi1150 & n41118;
  assign n41120 = pi214 & ~n41081;
  assign n41121 = n41077 & ~n41120;
  assign n41122 = n41072 & ~n41121;
  assign n41123 = n38140 & ~n41122;
  assign n41124 = n40612 & ~n41123;
  assign n41125 = ~n38138 & n38173;
  assign n41126 = ~n40866 & ~n41125;
  assign n41127 = ~n41124 & ~n41126;
  assign n41128 = ~pi214 & n38074;
  assign n41129 = ~n41096 & ~n41128;
  assign n41130 = pi212 & n41129;
  assign n41131 = n41111 & ~n41130;
  assign n41132 = ~n38092 & ~n41131;
  assign n41133 = ~po1038 & n41132;
  assign n41134 = n39533 & ~n41133;
  assign n41135 = n38089 & n38911;
  assign n41136 = ~n38087 & ~n38911;
  assign n41137 = ~po1038 & ~n41136;
  assign n41138 = ~n41135 & n41137;
  assign n41139 = n40659 & ~n41138;
  assign n41140 = pi1152 & ~n41139;
  assign n41141 = ~n41134 & n41140;
  assign n41142 = ~pi1150 & ~n41141;
  assign n41143 = ~n41127 & n41142;
  assign n41144 = ~pi213 & ~n41143;
  assign n41145 = ~n41119 & n41144;
  assign n41146 = pi213 & n38171;
  assign n41147 = pi209 & ~n41146;
  assign n41148 = ~n41145 & n41147;
  assign n41149 = ~n41066 & ~n41148;
  assign n41150 = pi230 & ~n41149;
  assign n41151 = ~pi230 & ~pi249;
  assign po406 = ~n41150 & ~n41151;
  assign n41153 = n2533 & n11307;
  assign n41154 = ~n6099 & ~n41153;
  assign n41155 = ~pi75 & ~n41154;
  assign n41156 = n7260 & n8821;
  assign n41157 = ~n41155 & ~n41156;
  assign n41158 = ~pi87 & ~n41157;
  assign n41159 = ~pi250 & n8739;
  assign po407 = n41158 & n41159;
  assign n41161 = pi897 & n10614;
  assign n41162 = ~pi476 & n11221;
  assign n41163 = ~n41161 & ~n41162;
  assign n41164 = pi200 & pi1039;
  assign n41165 = ~pi200 & pi1053;
  assign n41166 = ~pi199 & ~n41165;
  assign n41167 = ~n41164 & n41166;
  assign n41168 = ~n41163 & ~n41167;
  assign n41169 = pi251 & n41163;
  assign po408 = n41168 | n41169;
  assign n41171 = ~pi979 & ~pi984;
  assign n41172 = pi1001 & n41171;
  assign n41173 = n6180 & n41172;
  assign n41174 = ~n6121 & n41173;
  assign n41175 = n6440 & n41174;
  assign n41176 = ~pi252 & ~n41175;
  assign n41177 = pi1092 & ~n41176;
  assign n41178 = ~pi1093 & n41177;
  assign n41179 = n6456 & ~n41178;
  assign n41180 = n6455 & n41178;
  assign n41181 = ~n41179 & ~n41180;
  assign n41182 = ~n6215 & n41181;
  assign n41183 = n6215 & n11404;
  assign n41184 = ~n41182 & ~n41183;
  assign n41185 = ~n6198 & ~n41184;
  assign n41186 = pi299 & ~n41185;
  assign n41187 = ~n6191 & n11404;
  assign n41188 = n6191 & n41181;
  assign n41189 = ~n41187 & ~n41188;
  assign n41190 = n6198 & ~n41189;
  assign n41191 = n41186 & ~n41190;
  assign n41192 = n6236 & ~n41189;
  assign n41193 = ~n6236 & ~n41184;
  assign n41194 = ~pi299 & ~n41193;
  assign n41195 = ~n41192 & n41194;
  assign n41196 = n10780 & ~n41195;
  assign n41197 = ~n41191 & n41196;
  assign n41198 = ~n10780 & n11404;
  assign n41199 = ~n7588 & ~n41198;
  assign n41200 = ~n41197 & n41199;
  assign n41201 = pi57 & n11403;
  assign n41202 = n7588 & ~n41201;
  assign n41203 = n20537 & ~n37568;
  assign n41204 = n6212 & n41173;
  assign n41205 = n6440 & n41204;
  assign n41206 = n10779 & n41205;
  assign n41207 = n41203 & n41206;
  assign n41208 = ~pi252 & ~n41207;
  assign n41209 = ~pi57 & ~n41208;
  assign n41210 = pi1092 & n41209;
  assign n41211 = n41202 & ~n41210;
  assign po409 = ~n41200 & ~n41211;
  assign n41213 = ~n12743 & ~n37645;
  assign n41214 = ~n37748 & n41213;
  assign n41215 = ~po1038 & n41214;
  assign n41216 = pi219 & n38421;
  assign n41217 = ~n41215 & ~n41216;
  assign n41218 = pi1153 & ~n41217;
  assign n41219 = ~pi1151 & ~n41218;
  assign n41220 = ~n11223 & ~n38423;
  assign n41221 = pi1151 & ~n41220;
  assign n41222 = pi211 & ~n37787;
  assign n41223 = ~pi211 & ~pi219;
  assign n41224 = pi1153 & ~n37714;
  assign n41225 = ~n38106 & ~n41224;
  assign n41226 = n41223 & n41225;
  assign n41227 = ~n41222 & ~n41226;
  assign n41228 = ~n37714 & ~n37782;
  assign n41229 = n10522 & ~n41228;
  assign n41230 = ~po1038 & ~n41229;
  assign n41231 = n41227 & n41230;
  assign n41232 = n41221 & ~n41231;
  assign n41233 = ~n41219 & ~n41232;
  assign n41234 = ~pi1152 & ~n41233;
  assign n41235 = ~n37771 & ~n38921;
  assign n41236 = pi1153 & ~n41235;
  assign n41237 = ~n11156 & ~n37645;
  assign n41238 = pi1151 & n41237;
  assign n41239 = ~n41236 & n41238;
  assign n41240 = ~pi1151 & ~n37712;
  assign n41241 = n10522 & n38388;
  assign n41242 = ~n11224 & ~n41241;
  assign n41243 = n41240 & n41242;
  assign n41244 = ~po1038 & ~n41243;
  assign n41245 = ~n41239 & n41244;
  assign n41246 = ~pi1151 & n41223;
  assign n41247 = ~n38423 & ~n41246;
  assign n41248 = pi1152 & ~n41247;
  assign n41249 = ~n41245 & n41248;
  assign n41250 = ~n41234 & ~n41249;
  assign n41251 = pi230 & ~n41250;
  assign n41252 = ~pi1153 & ~n39933;
  assign n41253 = ~n39888 & ~n39903;
  assign n41254 = n38921 & ~n39875;
  assign n41255 = n41253 & ~n41254;
  assign n41256 = ~n39882 & n39900;
  assign n41257 = n41255 & n41256;
  assign n41258 = pi1153 & ~n41257;
  assign n41259 = ~n41252 & ~n41258;
  assign n41260 = pi219 & n41259;
  assign n41261 = ~pi219 & n39985;
  assign n41262 = pi1153 & ~n39904;
  assign n41263 = n41261 & ~n41262;
  assign n41264 = pi253 & ~n41263;
  assign n41265 = ~n41260 & n41264;
  assign n41266 = ~n39893 & n39933;
  assign n41267 = ~pi211 & n41266;
  assign n41268 = ~n39895 & ~n41267;
  assign n41269 = pi1153 & ~n41268;
  assign n41270 = ~n39924 & ~n41269;
  assign n41271 = pi219 & n41270;
  assign n41272 = ~n39903 & ~n39923;
  assign n41273 = pi1153 & n39955;
  assign n41274 = ~pi219 & ~n41273;
  assign n41275 = ~n41272 & n41274;
  assign n41276 = ~pi253 & ~n41275;
  assign n41277 = ~n41271 & n41276;
  assign n41278 = ~n41265 & ~n41277;
  assign n41279 = ~po1038 & ~n41278;
  assign n41280 = pi253 & po1038;
  assign n41281 = pi219 & pi1091;
  assign n41282 = ~n37611 & n41281;
  assign n41283 = ~pi219 & ~n39875;
  assign n41284 = ~pi211 & ~n39865;
  assign n41285 = pi219 & ~n39891;
  assign n41286 = ~n41284 & n41285;
  assign n41287 = po1038 & ~n41286;
  assign n41288 = ~n41283 & n41287;
  assign n41289 = ~n41282 & n41288;
  assign n41290 = ~n41280 & ~n41289;
  assign n41291 = ~pi219 & ~n39876;
  assign n41292 = ~n39891 & ~n41291;
  assign n41293 = ~n41282 & n41292;
  assign n41294 = pi253 & ~n41293;
  assign n41295 = ~n41290 & ~n41294;
  assign n41296 = ~pi211 & ~n39875;
  assign n41297 = n41291 & ~n41296;
  assign n41298 = ~pi219 & ~n41297;
  assign n41299 = po1038 & n41298;
  assign n41300 = ~n39865 & n41299;
  assign n41301 = pi1151 & ~n41300;
  assign n41302 = ~n41295 & n41301;
  assign n41303 = ~n41279 & n41302;
  assign n41304 = ~n39960 & ~n41267;
  assign n41305 = n41291 & ~n41304;
  assign n41306 = ~n39929 & n40013;
  assign n41307 = ~n39900 & ~n41306;
  assign n41308 = ~pi1153 & n41307;
  assign n41309 = ~n40013 & ~n41308;
  assign n41310 = n41305 & ~n41309;
  assign n41311 = pi219 & n39883;
  assign n41312 = ~n39892 & ~n39899;
  assign n41313 = n41258 & ~n41312;
  assign n41314 = n41311 & ~n41313;
  assign n41315 = ~n41310 & ~n41314;
  assign n41316 = pi253 & ~n41315;
  assign n41317 = pi219 & ~n41270;
  assign n41318 = ~n39881 & n41317;
  assign n41319 = ~pi253 & ~n41318;
  assign n41320 = n41255 & ~n41308;
  assign n41321 = ~n39894 & n41320;
  assign n41322 = ~n41271 & n41321;
  assign n41323 = n41319 & ~n41322;
  assign n41324 = ~n41316 & ~n41323;
  assign n41325 = ~po1038 & n41324;
  assign n41326 = ~pi1151 & ~n41325;
  assign n41327 = ~n41303 & ~n41326;
  assign n41328 = n41283 & ~n41284;
  assign n41329 = n41291 & ~n41328;
  assign n41330 = pi219 & ~n39865;
  assign n41331 = po1038 & ~n41330;
  assign n41332 = ~n41329 & n41331;
  assign n41333 = ~n39865 & n41332;
  assign n41334 = ~n41295 & ~n41333;
  assign n41335 = ~n41327 & n41334;
  assign n41336 = pi1152 & ~n41335;
  assign n41337 = ~n41275 & n41305;
  assign n41338 = ~n41317 & ~n41337;
  assign n41339 = ~n39893 & ~n41338;
  assign n41340 = ~pi253 & ~n41339;
  assign n41341 = n41255 & ~n41262;
  assign n41342 = n41291 & n41341;
  assign n41343 = ~n39953 & ~n41259;
  assign n41344 = pi219 & ~n41343;
  assign n41345 = ~n41342 & ~n41344;
  assign n41346 = pi253 & ~n41345;
  assign n41347 = ~po1038 & ~n41346;
  assign n41348 = ~n41340 & n41347;
  assign n41349 = n41302 & ~n41348;
  assign n41350 = ~pi1152 & ~n41349;
  assign n41351 = ~n41257 & ~n41312;
  assign n41352 = ~pi1091 & ~n39924;
  assign n41353 = ~pi1153 & ~n41352;
  assign n41354 = ~pi219 & ~n41307;
  assign n41355 = ~n41353 & ~n41354;
  assign n41356 = n41351 & n41355;
  assign n41357 = pi253 & ~n41356;
  assign n41358 = ~pi1153 & ~n39983;
  assign n41359 = ~n39893 & ~n41358;
  assign n41360 = n41261 & n41359;
  assign n41361 = n41319 & ~n41360;
  assign n41362 = ~n41357 & ~n41361;
  assign n41363 = ~po1038 & n41362;
  assign n41364 = ~pi1151 & ~n41295;
  assign n41365 = ~n41363 & n41364;
  assign n41366 = n41350 & ~n41365;
  assign n41367 = ~n41336 & ~n41366;
  assign n41368 = n40049 & ~n41367;
  assign n41369 = pi1091 & ~n41227;
  assign n41370 = pi1091 & n10522;
  assign n41371 = ~n38077 & ~n39825;
  assign n41372 = n41370 & ~n41371;
  assign n41373 = ~n41369 & ~n41372;
  assign n41374 = pi253 & ~n41373;
  assign n41375 = ~pi253 & ~pi1091;
  assign n41376 = ~po1038 & ~n41375;
  assign n41377 = ~n12746 & ~n41236;
  assign n41378 = ~pi253 & n41377;
  assign n41379 = n41376 & ~n41378;
  assign n41380 = ~n41374 & n41379;
  assign n41381 = pi1151 & ~n41380;
  assign n41382 = po1038 & ~n41375;
  assign n41383 = pi211 & pi1091;
  assign n41384 = pi1091 & ~pi1153;
  assign n41385 = pi219 & n41384;
  assign n41386 = ~n41383 & ~n41385;
  assign n41387 = n41382 & n41386;
  assign n41388 = n41381 & ~n41387;
  assign n41389 = pi1091 & pi1153;
  assign n41390 = n41215 & n41389;
  assign n41391 = ~pi1151 & ~n41390;
  assign n41392 = pi253 & ~pi1091;
  assign n41393 = ~n41282 & n41382;
  assign n41394 = pi219 & n41393;
  assign n41395 = ~n41392 & ~n41394;
  assign n41396 = n41391 & n41395;
  assign n41397 = ~n41388 & ~n41396;
  assign n41398 = ~pi1152 & ~n41397;
  assign n41399 = n41235 & ~n41392;
  assign n41400 = ~n41384 & ~n41399;
  assign n41401 = n41237 & ~n41400;
  assign n41402 = n41376 & ~n41401;
  assign n41403 = ~n41393 & ~n41402;
  assign n41404 = pi1151 & ~n41403;
  assign n41405 = ~pi211 & pi1091;
  assign n41406 = ~pi219 & n41405;
  assign n41407 = n41393 & ~n41406;
  assign n41408 = ~n37710 & n39792;
  assign n41409 = pi1153 & ~n41408;
  assign n41410 = n10522 & ~n41409;
  assign n41411 = n39830 & n41410;
  assign n41412 = pi253 & ~n41411;
  assign n41413 = n11223 & ~n37712;
  assign n41414 = n39792 & n41413;
  assign n41415 = n41412 & ~n41414;
  assign n41416 = pi1091 & n37712;
  assign n41417 = ~n39847 & ~n41416;
  assign n41418 = pi211 & n41417;
  assign n41419 = pi1091 & n38388;
  assign n41420 = n38079 & n39825;
  assign n41421 = n10522 & ~n41420;
  assign n41422 = ~n41419 & n41421;
  assign n41423 = ~pi253 & ~n41422;
  assign n41424 = ~n41418 & n41423;
  assign n41425 = ~n41415 & ~n41424;
  assign n41426 = n38737 & ~n41425;
  assign n41427 = ~n10522 & ~n11223;
  assign n41428 = ~n41392 & n41427;
  assign n41429 = ~n41416 & n41428;
  assign n41430 = n41426 & ~n41429;
  assign n41431 = pi1152 & ~n41430;
  assign n41432 = ~n41407 & n41431;
  assign n41433 = ~n41404 & n41432;
  assign n41434 = ~n41398 & ~n41433;
  assign n41435 = ~n40049 & n41434;
  assign n41436 = ~pi230 & ~n41435;
  assign n41437 = ~n41368 & n41436;
  assign po410 = ~n41251 & ~n41437;
  assign n41439 = ~pi1154 & n37760;
  assign n41440 = n38101 & ~n41439;
  assign n41441 = n11223 & n41440;
  assign n41442 = pi299 & n10522;
  assign n41443 = ~n11223 & n38080;
  assign n41444 = ~n41442 & ~n41443;
  assign n41445 = ~n38130 & ~n41444;
  assign n41446 = ~n41441 & ~n41445;
  assign n41447 = ~po1038 & ~n41446;
  assign n41448 = ~pi1152 & ~n41447;
  assign n41449 = ~pi219 & ~n38006;
  assign n41450 = ~n38228 & ~n41449;
  assign n41451 = po1038 & n41450;
  assign n41452 = n41448 & ~n41451;
  assign n41453 = n11223 & ~n38006;
  assign n41454 = n39071 & ~n41453;
  assign n41455 = pi1152 & ~n41454;
  assign n41456 = ~pi200 & pi1154;
  assign n41457 = n11164 & ~n41456;
  assign n41458 = n38100 & ~n38921;
  assign n41459 = ~n41457 & ~n41458;
  assign n41460 = ~pi219 & ~n41459;
  assign n41461 = ~n37779 & ~n38100;
  assign n41462 = n37604 & ~n41461;
  assign n41463 = n38063 & ~n38132;
  assign n41464 = ~n41462 & ~n41463;
  assign n41465 = pi219 & ~n41464;
  assign n41466 = ~po1038 & ~n41465;
  assign n41467 = ~n41460 & n41466;
  assign n41468 = n41455 & ~n41467;
  assign n41469 = ~n41452 & ~n41468;
  assign n41470 = pi230 & ~n41469;
  assign n41471 = pi1091 & ~n41450;
  assign n41472 = ~pi254 & ~pi1091;
  assign n41473 = po1038 & ~n41472;
  assign n41474 = ~n41471 & n41473;
  assign n41475 = ~n41280 & ~n41474;
  assign n41476 = n41328 & ~n41389;
  assign n41477 = pi1091 & n38228;
  assign n41478 = ~pi254 & ~n41477;
  assign n41479 = ~n41286 & n41478;
  assign n41480 = ~n41476 & n41479;
  assign n41481 = ~n41298 & n41480;
  assign n41482 = n11223 & n41384;
  assign n41483 = pi254 & ~n41477;
  assign n41484 = ~pi211 & ~n39889;
  assign n41485 = n41330 & ~n41484;
  assign n41486 = ~pi219 & n39875;
  assign n41487 = ~n41485 & ~n41486;
  assign n41488 = n41483 & n41487;
  assign n41489 = ~n41482 & n41488;
  assign n41490 = ~n41329 & n41489;
  assign n41491 = pi253 & ~n41490;
  assign n41492 = ~n41481 & n41491;
  assign n41493 = ~n41475 & ~n41492;
  assign n41494 = ~pi1152 & ~n41493;
  assign n41495 = pi1153 & ~n39811;
  assign n41496 = ~pi1154 & ~n41495;
  assign n41497 = pi211 & ~n41496;
  assign n41498 = ~pi1153 & ~n37748;
  assign n41499 = pi1091 & n41498;
  assign n41500 = ~n41419 & ~n41499;
  assign n41501 = ~n38106 & ~n41500;
  assign n41502 = n41497 & n41501;
  assign n41503 = pi1091 & n38080;
  assign n41504 = n11222 & n41389;
  assign n41505 = ~pi1154 & ~n41504;
  assign n41506 = ~pi211 & ~n41505;
  assign n41507 = n41503 & n41506;
  assign n41508 = ~n41502 & ~n41507;
  assign n41509 = ~pi219 & ~n41508;
  assign n41510 = n37613 & n41500;
  assign n41511 = n37604 & ~n41503;
  assign n41512 = ~n41505 & ~n41511;
  assign n41513 = pi219 & n41512;
  assign n41514 = ~n41510 & n41513;
  assign n41515 = ~n41509 & ~n41514;
  assign n41516 = ~pi254 & ~n41515;
  assign n41517 = pi1091 & ~n11223;
  assign n41518 = ~n38062 & n41517;
  assign n41519 = ~pi1154 & ~n41518;
  assign n41520 = pi1091 & ~n37711;
  assign n41521 = pi1091 & ~n41501;
  assign n41522 = ~n41520 & ~n41521;
  assign n41523 = n41427 & ~n41522;
  assign n41524 = n39841 & n41410;
  assign n41525 = pi1154 & ~n41524;
  assign n41526 = ~n41523 & n41525;
  assign n41527 = ~n41519 & ~n41526;
  assign n41528 = ~pi1154 & n39815;
  assign n41529 = ~n41521 & ~n41528;
  assign n41530 = n11223 & ~n41529;
  assign n41531 = pi254 & ~n41530;
  assign n41532 = ~n41527 & n41531;
  assign n41533 = ~n41516 & ~n41532;
  assign n41534 = ~pi253 & n41533;
  assign n41535 = n37613 & ~n41312;
  assign n41536 = pi219 & ~n41535;
  assign n41537 = ~n39881 & n39912;
  assign n41538 = ~pi1154 & n41537;
  assign n41539 = ~pi1153 & n39900;
  assign n41540 = ~n41256 & ~n41539;
  assign n41541 = ~n41538 & n41540;
  assign n41542 = n41536 & ~n41541;
  assign n41543 = n41304 & ~n41539;
  assign n41544 = pi1154 & n39899;
  assign n41545 = ~pi219 & ~n41544;
  assign n41546 = ~n41543 & n41545;
  assign n41547 = ~n41542 & ~n41546;
  assign n41548 = pi254 & ~n41547;
  assign n41549 = pi1154 & n39888;
  assign n41550 = ~n39929 & ~n41549;
  assign n41551 = ~pi211 & ~n41550;
  assign n41552 = ~pi219 & ~n41551;
  assign n41553 = ~n39894 & n39944;
  assign n41554 = pi1154 & n41553;
  assign n41555 = ~n41272 & ~n41554;
  assign n41556 = ~pi1153 & ~n39985;
  assign n41557 = ~n39888 & ~n41556;
  assign n41558 = ~n41555 & n41557;
  assign n41559 = n41552 & n41558;
  assign n41560 = ~pi254 & ~n41559;
  assign n41561 = ~n41252 & n41553;
  assign n41562 = n37613 & ~n41561;
  assign n41563 = ~pi1153 & ~n39938;
  assign n41564 = n39926 & ~n41563;
  assign n41565 = ~pi1154 & ~n41564;
  assign n41566 = n39896 & ~n41252;
  assign n41567 = n37604 & ~n41566;
  assign n41568 = pi219 & ~n41567;
  assign n41569 = ~n41565 & n41568;
  assign n41570 = ~n41562 & n41569;
  assign n41571 = n41560 & ~n41570;
  assign n41572 = ~n41548 & ~n41571;
  assign n41573 = pi253 & ~n41572;
  assign n41574 = ~po1038 & ~n41573;
  assign n41575 = ~n41534 & n41574;
  assign n41576 = n41494 & ~n41575;
  assign n41577 = ~pi1153 & ~n39797;
  assign n41578 = n41496 & ~n41577;
  assign n41579 = ~pi211 & n38106;
  assign n41580 = n41578 & ~n41579;
  assign n41581 = pi1091 & ~n38141;
  assign n41582 = ~n37771 & n41581;
  assign n41583 = n37604 & n41582;
  assign n41584 = ~n41580 & ~n41583;
  assign n41585 = ~pi219 & ~n41584;
  assign n41586 = pi1154 & n41405;
  assign n41587 = ~n41281 & ~n41586;
  assign n41588 = ~n41464 & ~n41587;
  assign n41589 = ~n41585 & ~n41588;
  assign n41590 = pi254 & ~n41589;
  assign n41591 = pi1154 & ~n41235;
  assign n41592 = ~n38132 & ~n41591;
  assign n41593 = pi219 & n41592;
  assign n41594 = ~n41460 & ~n41593;
  assign n41595 = ~pi254 & ~n41594;
  assign n41596 = ~n41472 & ~n41595;
  assign n41597 = ~n41590 & n41596;
  assign n41598 = ~pi253 & ~n41597;
  assign n41599 = ~n39953 & ~n41257;
  assign n41600 = ~n41258 & ~n41599;
  assign n41601 = pi1154 & n41600;
  assign n41602 = pi1153 & ~n39933;
  assign n41603 = ~pi1154 & n39944;
  assign n41604 = ~n41602 & n41603;
  assign n41605 = pi254 & ~n41604;
  assign n41606 = ~n41601 & n41605;
  assign n41607 = ~n39867 & n41562;
  assign n41608 = pi1153 & n39895;
  assign n41609 = n37604 & ~n39912;
  assign n41610 = ~n41608 & n41609;
  assign n41611 = ~n39893 & n39924;
  assign n41612 = n41565 & ~n41611;
  assign n41613 = ~pi254 & ~n41612;
  assign n41614 = ~n41610 & n41613;
  assign n41615 = ~n41607 & n41614;
  assign n41616 = ~n41606 & ~n41615;
  assign n41617 = pi219 & ~n41616;
  assign n41618 = n41341 & ~n41543;
  assign n41619 = ~n39985 & ~n41618;
  assign n41620 = ~pi1154 & ~n41619;
  assign n41621 = pi254 & ~n41620;
  assign n41622 = pi1154 & ~n39887;
  assign n41623 = n41618 & n41622;
  assign n41624 = n41621 & ~n41623;
  assign n41625 = ~pi254 & ~n41555;
  assign n41626 = ~pi1153 & ~n41254;
  assign n41627 = ~n39930 & n41626;
  assign n41628 = n41625 & ~n41627;
  assign n41629 = ~n41624 & ~n41628;
  assign n41630 = ~pi219 & ~n41629;
  assign n41631 = ~n41617 & ~n41630;
  assign n41632 = pi253 & n41631;
  assign n41633 = ~n41598 & ~n41632;
  assign n41634 = ~po1038 & n41633;
  assign n41635 = pi253 & ~n41489;
  assign n41636 = ~n41480 & n41635;
  assign n41637 = po1038 & n41406;
  assign n41638 = ~n41474 & ~n41637;
  assign n41639 = ~n41280 & n41638;
  assign n41640 = ~n41636 & ~n41639;
  assign n41641 = pi1152 & ~n41640;
  assign n41642 = ~n41634 & n41641;
  assign n41643 = ~n41576 & ~n41642;
  assign n41644 = n40049 & n41643;
  assign n41645 = ~po1038 & n41597;
  assign n41646 = n41638 & ~n41645;
  assign n41647 = pi1152 & n41646;
  assign n41648 = ~po1038 & ~n41533;
  assign n41649 = ~pi1152 & ~n41474;
  assign n41650 = ~n41648 & n41649;
  assign n41651 = ~n40049 & ~n41650;
  assign n41652 = ~n41647 & n41651;
  assign n41653 = ~pi230 & ~n41652;
  assign n41654 = ~n41644 & n41653;
  assign po411 = ~n41470 & ~n41654;
  assign n41656 = ~pi200 & pi1049;
  assign n41657 = pi200 & pi1036;
  assign n41658 = ~n41656 & ~n41657;
  assign n41659 = ~n41163 & n41658;
  assign n41660 = ~pi255 & n41163;
  assign po412 = ~n41659 & ~n41660;
  assign n41662 = ~pi200 & pi1048;
  assign n41663 = pi200 & pi1070;
  assign n41664 = ~n41662 & ~n41663;
  assign n41665 = ~n41163 & n41664;
  assign n41666 = ~pi256 & n41163;
  assign po413 = ~n41665 & ~n41666;
  assign n41668 = ~pi200 & pi1084;
  assign n41669 = pi200 & pi1065;
  assign n41670 = ~n41668 & ~n41669;
  assign n41671 = ~n41163 & n41670;
  assign n41672 = ~pi257 & n41163;
  assign po414 = ~n41671 & ~n41672;
  assign n41674 = ~pi200 & pi1072;
  assign n41675 = pi200 & pi1062;
  assign n41676 = ~n41674 & ~n41675;
  assign n41677 = ~n41163 & n41676;
  assign n41678 = ~pi258 & n41163;
  assign po415 = ~n41677 & ~n41678;
  assign n41680 = ~pi200 & pi1059;
  assign n41681 = pi200 & pi1069;
  assign n41682 = ~n41680 & ~n41681;
  assign n41683 = ~n41163 & n41682;
  assign n41684 = ~pi259 & n41163;
  assign po416 = ~n41683 & ~n41684;
  assign n41686 = pi200 & pi1067;
  assign n41687 = ~pi200 & pi1044;
  assign n41688 = ~pi199 & ~n41687;
  assign n41689 = ~n41686 & n41688;
  assign n41690 = ~n41163 & ~n41689;
  assign n41691 = pi260 & n41163;
  assign po417 = n41690 | n41691;
  assign n41693 = pi200 & pi1040;
  assign n41694 = ~pi200 & pi1037;
  assign n41695 = ~pi199 & ~n41694;
  assign n41696 = ~n41693 & n41695;
  assign n41697 = ~n41163 & ~n41696;
  assign n41698 = pi261 & n41163;
  assign po418 = n41697 | n41698;
  assign n41700 = pi1093 & pi1142;
  assign n41701 = ~pi262 & ~pi1093;
  assign n41702 = ~n41700 & ~n41701;
  assign n41703 = ~pi228 & ~n41702;
  assign n41704 = pi123 & pi262;
  assign n41705 = ~pi123 & ~pi1142;
  assign n41706 = pi228 & ~n41705;
  assign n41707 = ~n41704 & n41706;
  assign n41708 = ~n41703 & ~n41707;
  assign n41709 = ~pi228 & ~pi1093;
  assign n41710 = pi123 & pi228;
  assign n41711 = ~n41709 & ~n41710;
  assign n41712 = ~pi262 & ~n41711;
  assign n41713 = ~n39673 & ~n41712;
  assign n41714 = pi199 & n41711;
  assign n41715 = n37633 & ~n41714;
  assign n41716 = n41713 & ~n41715;
  assign n41717 = ~n41708 & ~n41716;
  assign n41718 = ~pi207 & n41712;
  assign n41719 = ~pi208 & ~n41718;
  assign n41720 = ~n39673 & ~n41719;
  assign n41721 = ~n41717 & ~n41720;
  assign n41722 = ~n38769 & n41711;
  assign n41723 = ~pi299 & ~n41722;
  assign n41724 = ~n41708 & n41723;
  assign n41725 = pi299 & ~n41713;
  assign n41726 = pi208 & ~n41725;
  assign n41727 = ~n41724 & n41726;
  assign n41728 = ~n41721 & ~n41727;
  assign n41729 = ~po1038 & n41728;
  assign n41730 = ~n38857 & n41711;
  assign n41731 = po1038 & ~n41708;
  assign n41732 = ~n41730 & n41731;
  assign po419 = n41729 | n41732;
  assign n41734 = ~n39925 & ~n39955;
  assign n41735 = ~n39896 & ~n41549;
  assign n41736 = ~n41734 & ~n41735;
  assign n41737 = n37596 & ~n41736;
  assign n41738 = ~n39923 & n41736;
  assign n41739 = ~pi1156 & ~n41738;
  assign n41740 = pi1154 & ~n41734;
  assign n41741 = ~pi1154 & ~n39990;
  assign n41742 = ~n39923 & n39978;
  assign n41743 = pi1155 & n41742;
  assign n41744 = n41741 & ~n41743;
  assign n41745 = ~n40003 & n41744;
  assign n41746 = ~pi299 & n41745;
  assign n41747 = n41603 & ~n41746;
  assign n41748 = n37599 & ~n41747;
  assign n41749 = ~n41740 & n41748;
  assign n41750 = pi219 & ~n41749;
  assign n41751 = ~n41739 & n41750;
  assign n41752 = ~n41737 & n41751;
  assign n41753 = pi263 & ~n41752;
  assign n41754 = pi1154 & ~n40009;
  assign n41755 = ~n39931 & n41754;
  assign n41756 = ~n39887 & n41272;
  assign n41757 = pi1155 & n41756;
  assign n41758 = n41741 & ~n41757;
  assign n41759 = ~n39980 & n41754;
  assign n41760 = ~pi1156 & ~n41544;
  assign n41761 = ~n41759 & n41760;
  assign n41762 = ~pi1156 & ~n41761;
  assign n41763 = ~n41758 & ~n41762;
  assign n41764 = pi1156 & n40003;
  assign n41765 = ~n41763 & ~n41764;
  assign n41766 = ~n41755 & ~n41765;
  assign n41767 = pi211 & ~n41766;
  assign n41768 = ~n41745 & ~n41759;
  assign n41769 = pi1156 & n41768;
  assign n41770 = ~n41744 & n41761;
  assign n41771 = ~pi211 & ~n41770;
  assign n41772 = ~n41769 & n41771;
  assign n41773 = ~pi219 & ~n41772;
  assign n41774 = ~n41767 & n41773;
  assign n41775 = n41753 & ~n41774;
  assign n41776 = ~pi1155 & n41352;
  assign n41777 = pi1155 & ~n39883;
  assign n41778 = ~pi1154 & ~n41777;
  assign n41779 = ~n41776 & n41778;
  assign n41780 = pi1155 & n39882;
  assign n41781 = pi1154 & ~n41780;
  assign n41782 = n39944 & n41781;
  assign n41783 = ~n41779 & ~n41782;
  assign n41784 = ~pi1156 & ~n41783;
  assign n41785 = n39900 & n41778;
  assign n41786 = ~n39887 & n41782;
  assign n41787 = ~n41785 & ~n41786;
  assign n41788 = n37596 & ~n41787;
  assign n41789 = pi219 & ~n41788;
  assign n41790 = ~pi1154 & n39924;
  assign n41791 = ~n39953 & ~n41790;
  assign n41792 = ~n41780 & ~n41791;
  assign n41793 = n37599 & n41792;
  assign n41794 = n41789 & ~n41793;
  assign n41795 = ~n41784 & n41794;
  assign n41796 = pi1155 & ~n39960;
  assign n41797 = ~pi1154 & ~n41796;
  assign n41798 = ~n41307 & n41797;
  assign n41799 = pi1156 & ~n41798;
  assign n41800 = pi1155 & ~n39985;
  assign n41801 = pi1154 & ~n41800;
  assign n41802 = n40016 & n41801;
  assign n41803 = ~n39885 & n41802;
  assign n41804 = ~n41785 & ~n41803;
  assign n41805 = n41799 & n41804;
  assign n41806 = ~n41272 & n41776;
  assign n41807 = n41797 & ~n41806;
  assign n41808 = ~pi1156 & ~n41807;
  assign n41809 = ~n41779 & ~n41802;
  assign n41810 = n41808 & n41809;
  assign n41811 = ~pi211 & ~n41810;
  assign n41812 = ~n41805 & n41811;
  assign n41813 = n41253 & n41801;
  assign n41814 = n41808 & ~n41813;
  assign n41815 = n39904 & n41801;
  assign n41816 = n41799 & ~n41815;
  assign n41817 = pi211 & ~n41816;
  assign n41818 = ~n41814 & n41817;
  assign n41819 = ~pi219 & ~n41818;
  assign n41820 = ~n41812 & n41819;
  assign n41821 = ~pi263 & ~n41820;
  assign n41822 = ~n41795 & n41821;
  assign n41823 = ~n41775 & ~n41822;
  assign n41824 = n39789 & n41823;
  assign n41825 = pi1155 & ~n37971;
  assign n41826 = n39825 & ~n41825;
  assign n41827 = ~pi1154 & n41520;
  assign n41828 = ~n41826 & ~n41827;
  assign n41829 = ~n39847 & n41828;
  assign n41830 = n37596 & ~n41829;
  assign n41831 = pi1091 & ~pi1154;
  assign n41832 = ~n39797 & ~n41831;
  assign n41833 = ~pi1156 & ~n41832;
  assign n41834 = ~n37719 & n41833;
  assign n41835 = pi219 & ~n41834;
  assign n41836 = pi1154 & ~n10615;
  assign n41837 = ~n37719 & ~n41836;
  assign n41838 = n37599 & n39841;
  assign n41839 = n41837 & n41838;
  assign n41840 = n41835 & ~n41839;
  assign n41841 = ~n41830 & n41840;
  assign n41842 = ~pi211 & ~n41828;
  assign n41843 = ~pi199 & ~pi1154;
  assign n41844 = n37771 & ~n41843;
  assign n41845 = ~n37851 & ~n41844;
  assign n41846 = n41383 & n41845;
  assign n41847 = ~n41842 & ~n41846;
  assign n41848 = pi1156 & ~n41847;
  assign n41849 = ~n37851 & ~n41832;
  assign n41850 = pi211 & n41849;
  assign n41851 = n41405 & n41837;
  assign n41852 = ~n41850 & ~n41851;
  assign n41853 = ~pi1156 & ~n41852;
  assign n41854 = ~pi219 & ~n41853;
  assign n41855 = ~n41848 & n41854;
  assign n41856 = ~n41841 & ~n41855;
  assign n41857 = ~pi263 & ~n41856;
  assign n41858 = pi1154 & ~n37721;
  assign n41859 = pi1156 & ~n41858;
  assign n41860 = ~pi299 & ~n41859;
  assign n41861 = ~n41837 & n41860;
  assign n41862 = ~n37722 & ~n38921;
  assign n41863 = ~n41860 & n41862;
  assign n41864 = pi1156 & ~n41863;
  assign n41865 = ~n41861 & ~n41864;
  assign n41866 = pi219 & n41865;
  assign n41867 = ~n37724 & n38615;
  assign n41868 = ~n41836 & ~n41867;
  assign n41869 = ~pi211 & ~n41868;
  assign n41870 = ~pi219 & ~n41869;
  assign n41871 = ~n37707 & ~n37771;
  assign n41872 = pi1154 & ~n41871;
  assign n41873 = ~pi1154 & ~n37819;
  assign n41874 = ~n37793 & n41873;
  assign n41875 = pi1156 & ~n41874;
  assign n41876 = ~n41872 & n41875;
  assign n41877 = ~pi1156 & n41849;
  assign n41878 = ~n41876 & ~n41877;
  assign n41879 = pi211 & n41878;
  assign n41880 = n41870 & ~n41879;
  assign n41881 = pi1091 & ~n41880;
  assign n41882 = pi263 & n41881;
  assign n41883 = ~n41866 & n41882;
  assign n41884 = ~n41857 & ~n41883;
  assign n41885 = ~n39789 & ~n41884;
  assign n41886 = ~po1038 & ~n41885;
  assign n41887 = ~n41824 & n41886;
  assign n41888 = pi211 & n39865;
  assign n41889 = ~pi211 & ~n41831;
  assign n41890 = ~n37600 & ~n41889;
  assign n41891 = ~n41888 & n41890;
  assign n41892 = ~n39875 & ~n41891;
  assign n41893 = ~pi219 & ~n41892;
  assign n41894 = ~pi263 & ~n41485;
  assign n41895 = ~n41893 & n41894;
  assign n41896 = ~n37600 & ~n41586;
  assign n41897 = ~n41888 & ~n41896;
  assign n41898 = n41283 & ~n41897;
  assign n41899 = ~n41286 & ~n41898;
  assign n41900 = pi263 & n41899;
  assign n41901 = ~n41895 & ~n41900;
  assign n41902 = n39789 & ~n41901;
  assign n41903 = pi219 & ~n37599;
  assign n41904 = pi1091 & n41903;
  assign n41905 = n41902 & ~n41904;
  assign n41906 = po1038 & ~n41905;
  assign n41907 = ~pi219 & ~n37600;
  assign n41908 = ~n37613 & n41907;
  assign n41909 = ~n41903 & ~n41908;
  assign n41910 = pi1091 & ~n41909;
  assign n41911 = pi263 & ~pi1091;
  assign n41912 = ~n41910 & ~n41911;
  assign n41913 = ~n39789 & n41912;
  assign n41914 = n41906 & ~n41913;
  assign n41915 = ~n41887 & ~n41914;
  assign n41916 = n40049 & n41915;
  assign n41917 = po1038 & ~n41912;
  assign n41918 = ~po1038 & n41884;
  assign n41919 = ~n40049 & ~n41918;
  assign n41920 = ~n41917 & n41919;
  assign n41921 = ~pi230 & ~n41920;
  assign n41922 = ~n41916 & n41921;
  assign n41923 = ~n37720 & n37725;
  assign n41924 = ~pi1156 & ~n41923;
  assign n41925 = ~pi200 & n41843;
  assign n41926 = n37973 & ~n41925;
  assign n41927 = ~n41924 & n41926;
  assign n41928 = ~n37647 & ~n41927;
  assign n41929 = pi211 & ~n41928;
  assign n41930 = n41870 & ~n41929;
  assign n41931 = pi1156 & n38921;
  assign n41932 = ~n41927 & ~n41931;
  assign n41933 = pi219 & n41932;
  assign n41934 = ~n41930 & ~n41933;
  assign n41935 = ~po1038 & n41934;
  assign n41936 = po1038 & n41909;
  assign n41937 = pi230 & ~n41936;
  assign n41938 = ~n41935 & n41937;
  assign po420 = ~n41922 & ~n41938;
  assign n41940 = pi219 & ~n41405;
  assign n41941 = ~n38497 & ~n41940;
  assign n41942 = pi264 & ~n39858;
  assign n41943 = ~pi796 & n39858;
  assign n41944 = ~pi1091 & ~n41943;
  assign n41945 = ~n41942 & n41944;
  assign n41946 = ~n41941 & ~n41945;
  assign n41947 = pi1091 & pi1141;
  assign n41948 = pi264 & ~n39870;
  assign n41949 = ~pi796 & n39870;
  assign n41950 = ~pi1091 & ~n41949;
  assign n41951 = ~n41948 & n41950;
  assign n41952 = ~n41947 & ~n41951;
  assign n41953 = ~pi211 & ~n41952;
  assign n41954 = pi1091 & pi1142;
  assign n41955 = ~n41951 & ~n41954;
  assign n41956 = pi211 & ~n41955;
  assign n41957 = ~pi219 & ~n41956;
  assign n41958 = ~n41953 & n41957;
  assign n41959 = ~n41946 & ~n41958;
  assign n41960 = ~n15973 & ~n41959;
  assign n41961 = ~pi230 & ~n41960;
  assign n41962 = pi1091 & pi1143;
  assign n41963 = ~pi200 & n41962;
  assign n41964 = pi199 & ~n41945;
  assign n41965 = ~n41963 & n41964;
  assign n41966 = ~pi200 & ~n41952;
  assign n41967 = pi200 & ~n41955;
  assign n41968 = ~pi199 & ~n41967;
  assign n41969 = ~n41966 & n41968;
  assign n41970 = ~n41965 & ~n41969;
  assign n41971 = n15973 & ~n41970;
  assign n41972 = n41961 & ~n41971;
  assign n41973 = ~pi199 & pi1141;
  assign n41974 = n38466 & ~n41973;
  assign n41975 = ~n37636 & ~n41974;
  assign n41976 = n15973 & ~n41975;
  assign n41977 = ~pi211 & pi1141;
  assign n41978 = ~pi219 & ~n37683;
  assign n41979 = ~n41977 & n41978;
  assign n41980 = ~n38497 & ~n41979;
  assign n41981 = ~n15973 & ~n41980;
  assign n41982 = pi230 & ~n41981;
  assign n41983 = ~n41976 & n41982;
  assign po421 = n41972 | n41983;
  assign n41985 = ~n39722 & ~n41940;
  assign n41986 = pi265 & ~n39858;
  assign n41987 = ~pi819 & n39858;
  assign n41988 = ~pi1091 & ~n41987;
  assign n41989 = ~n41986 & n41988;
  assign n41990 = ~n41985 & ~n41989;
  assign n41991 = pi265 & ~n39870;
  assign n41992 = ~pi819 & n39870;
  assign n41993 = ~pi1091 & ~n41992;
  assign n41994 = ~n41991 & n41993;
  assign n41995 = ~n41954 & ~n41994;
  assign n41996 = ~pi211 & ~n41995;
  assign n41997 = ~n41962 & ~n41994;
  assign n41998 = pi211 & ~n41997;
  assign n41999 = ~pi219 & ~n41998;
  assign n42000 = ~n41996 & n41999;
  assign n42001 = ~n41990 & ~n42000;
  assign n42002 = ~n15973 & ~n42001;
  assign n42003 = ~pi230 & ~n42002;
  assign n42004 = pi1091 & pi1144;
  assign n42005 = ~pi200 & n42004;
  assign n42006 = pi199 & ~n42005;
  assign n42007 = ~n41989 & n42006;
  assign n42008 = ~pi200 & ~n41995;
  assign n42009 = pi200 & ~n41997;
  assign n42010 = ~pi199 & ~n42009;
  assign n42011 = ~n42008 & n42010;
  assign n42012 = ~n42007 & ~n42011;
  assign n42013 = n15973 & ~n42012;
  assign n42014 = n42003 & ~n42013;
  assign n42015 = ~n37635 & n39727;
  assign n42016 = ~n37629 & ~n42015;
  assign n42017 = n15973 & ~n42016;
  assign n42018 = ~pi219 & ~n37666;
  assign n42019 = ~n37694 & n42018;
  assign n42020 = ~n39722 & ~n42019;
  assign n42021 = ~n15973 & ~n42020;
  assign n42022 = pi230 & ~n42021;
  assign n42023 = ~n42017 & n42022;
  assign po422 = n42014 | n42023;
  assign n42025 = ~pi211 & pi1136;
  assign n42026 = pi219 & ~n42025;
  assign n42027 = pi211 & ~pi1135;
  assign n42028 = ~n42026 & ~n42027;
  assign n42029 = ~n41223 & n42028;
  assign n42030 = pi299 & n42029;
  assign n42031 = pi199 & pi1136;
  assign n42032 = ~pi200 & ~n42031;
  assign n42033 = ~pi199 & pi1135;
  assign n42034 = pi200 & ~n42033;
  assign n42035 = ~pi299 & ~n42034;
  assign n42036 = ~n42032 & n42035;
  assign n42037 = ~n42030 & ~n42036;
  assign n42038 = ~po1038 & ~n42037;
  assign n42039 = po1038 & n42029;
  assign n42040 = pi230 & ~n42039;
  assign n42041 = ~n42038 & n42040;
  assign n42042 = ~pi948 & n39870;
  assign n42043 = ~pi266 & ~n39870;
  assign n42044 = ~pi1091 & ~n42043;
  assign n42045 = ~n42042 & n42044;
  assign n42046 = ~pi199 & ~n42045;
  assign n42047 = pi1091 & pi1136;
  assign n42048 = ~pi948 & n39858;
  assign n42049 = ~pi266 & ~n39858;
  assign n42050 = ~pi1091 & ~n42049;
  assign n42051 = ~n42048 & n42050;
  assign n42052 = pi199 & ~n42051;
  assign n42053 = ~n42047 & n42052;
  assign n42054 = ~n42046 & ~n42053;
  assign n42055 = ~pi200 & n42054;
  assign n42056 = pi1091 & pi1135;
  assign n42057 = n42046 & ~n42056;
  assign n42058 = pi200 & ~n42052;
  assign n42059 = ~n42057 & n42058;
  assign n42060 = ~n42055 & ~n42059;
  assign n42061 = n15973 & ~n42060;
  assign n42062 = ~n41940 & ~n42026;
  assign n42063 = ~n42051 & ~n42062;
  assign n42064 = ~n15973 & ~n42063;
  assign n42065 = ~pi219 & ~n42045;
  assign n42066 = pi1135 & n41383;
  assign n42067 = n42065 & ~n42066;
  assign n42068 = n42064 & ~n42067;
  assign n42069 = ~pi230 & ~n42068;
  assign n42070 = ~n42061 & n42069;
  assign n42071 = ~n42041 & ~n42070;
  assign n42072 = ~pi1134 & ~n42071;
  assign n42073 = ~n15973 & n42028;
  assign n42074 = pi230 & ~n42073;
  assign n42075 = n37747 & ~n42031;
  assign n42076 = ~n42034 & ~n42075;
  assign n42077 = n15973 & n42076;
  assign n42078 = n42074 & ~n42077;
  assign n42079 = ~pi199 & pi1091;
  assign n42080 = ~n42054 & ~n42079;
  assign n42081 = ~pi200 & ~n42080;
  assign n42082 = ~n42059 & ~n42081;
  assign n42083 = n15973 & ~n42082;
  assign n42084 = pi1091 & ~n42027;
  assign n42085 = n42065 & ~n42084;
  assign n42086 = n42064 & ~n42085;
  assign n42087 = ~pi230 & ~n42086;
  assign n42088 = ~n42083 & n42087;
  assign n42089 = ~n42078 & ~n42088;
  assign n42090 = pi1134 & ~n42089;
  assign po423 = ~n42072 & ~n42090;
  assign n42092 = pi1155 & n38084;
  assign n42093 = pi1154 & ~n42092;
  assign n42094 = pi1091 & ~n38136;
  assign n42095 = ~n11222 & n42094;
  assign n42096 = n42093 & n42095;
  assign n42097 = ~n37749 & ~n39801;
  assign n42098 = n42094 & ~n42097;
  assign n42099 = ~pi1154 & n42098;
  assign n42100 = ~pi219 & ~n42099;
  assign n42101 = ~n42096 & n42100;
  assign n42102 = ~n41224 & ~n41498;
  assign n42103 = ~n37749 & n41831;
  assign n42104 = ~n42102 & n42103;
  assign n42105 = n41831 & ~n42104;
  assign n42106 = pi219 & ~n42105;
  assign n42107 = pi1091 & n41825;
  assign n42108 = ~n41577 & n42107;
  assign n42109 = pi1154 & ~n42108;
  assign n42110 = ~pi299 & n38067;
  assign n42111 = pi1091 & ~n42110;
  assign n42112 = n42109 & n42111;
  assign n42113 = n42106 & ~n42112;
  assign n42114 = ~n42101 & ~n42113;
  assign n42115 = ~pi211 & ~n42114;
  assign n42116 = ~n38150 & n41831;
  assign n42117 = ~n42097 & n42116;
  assign n42118 = pi211 & ~n42117;
  assign n42119 = ~pi1155 & ~n38068;
  assign n42120 = ~n37818 & ~n42119;
  assign n42121 = ~n12744 & ~n42120;
  assign n42122 = pi1091 & ~n42121;
  assign n42123 = n42093 & n42122;
  assign n42124 = n42118 & ~n42123;
  assign n42125 = ~n42115 & ~n42124;
  assign n42126 = pi267 & ~n42125;
  assign n42127 = ~n37715 & ~n37804;
  assign n42128 = ~n38106 & n42127;
  assign n42129 = pi1091 & n42128;
  assign n42130 = ~pi211 & ~n42129;
  assign n42131 = ~pi219 & ~n42130;
  assign n42132 = pi1091 & ~pi1155;
  assign n42133 = ~n38068 & n42132;
  assign n42134 = ~n42108 & ~n42133;
  assign n42135 = n37604 & n42134;
  assign n42136 = n42131 & ~n42135;
  assign n42137 = n42110 & n42132;
  assign n42138 = n42109 & ~n42137;
  assign n42139 = pi1154 & ~n42138;
  assign n42140 = ~pi211 & ~n42104;
  assign n42141 = ~n42139 & n42140;
  assign n42142 = n41825 & n42093;
  assign n42143 = ~n42138 & ~n42142;
  assign n42144 = pi211 & ~n42143;
  assign n42145 = pi219 & ~n42144;
  assign n42146 = ~n42141 & n42145;
  assign n42147 = ~n42136 & ~n42146;
  assign n42148 = ~pi267 & ~n42147;
  assign n42149 = n39792 & ~n42098;
  assign n42150 = ~pi1154 & ~n42149;
  assign n42151 = pi211 & n42150;
  assign n42152 = n42148 & ~n42151;
  assign n42153 = ~n42126 & ~n42152;
  assign n42154 = ~n39788 & ~n42153;
  assign n42155 = ~n41563 & n41611;
  assign n42156 = ~pi1154 & ~n41537;
  assign n42157 = ~n42155 & n42156;
  assign n42158 = pi1154 & ~n41608;
  assign n42159 = ~n39896 & n42158;
  assign n42160 = pi1155 & n42159;
  assign n42161 = ~n42157 & ~n42160;
  assign n42162 = pi211 & ~n42161;
  assign n42163 = n37603 & ~n41554;
  assign n42164 = ~n41266 & ~n41273;
  assign n42165 = n42163 & n42164;
  assign n42166 = ~pi267 & ~n42165;
  assign n42167 = pi1154 & n39926;
  assign n42168 = ~pi1155 & ~n42167;
  assign n42169 = ~n42155 & n42168;
  assign n42170 = n42166 & ~n42169;
  assign n42171 = ~n42162 & n42170;
  assign n42172 = n39883 & ~n41602;
  assign n42173 = pi1154 & ~n42172;
  assign n42174 = ~pi1154 & ~n39944;
  assign n42175 = ~n41353 & n42174;
  assign n42176 = ~pi1155 & ~n42175;
  assign n42177 = ~n42173 & n42176;
  assign n42178 = pi267 & ~n42177;
  assign n42179 = pi1155 & ~n41262;
  assign n42180 = pi1154 & n39882;
  assign n42181 = ~n41351 & ~n42180;
  assign n42182 = n42179 & n42181;
  assign n42183 = n42178 & ~n42182;
  assign n42184 = ~n42171 & ~n42183;
  assign n42185 = pi219 & ~n42184;
  assign n42186 = pi1155 & ~n41553;
  assign n42187 = ~n40003 & ~n41273;
  assign n42188 = n42186 & n42187;
  assign n42189 = pi1154 & ~n42188;
  assign n42190 = ~pi1154 & ~n41556;
  assign n42191 = pi1155 & ~n42190;
  assign n42192 = n39930 & ~n42191;
  assign n42193 = ~n42189 & ~n42192;
  assign n42194 = pi211 & ~n42193;
  assign n42195 = ~pi1155 & ~n41756;
  assign n42196 = ~n42155 & n42195;
  assign n42197 = n42194 & ~n42196;
  assign n42198 = pi1153 & ~n41272;
  assign n42199 = ~pi1155 & ~n42198;
  assign n42200 = pi1153 & n42199;
  assign n42201 = pi1155 & ~n42187;
  assign n42202 = pi1154 & ~n42201;
  assign n42203 = ~n41742 & n42202;
  assign n42204 = ~n42200 & n42203;
  assign n42205 = n41359 & n42199;
  assign n42206 = ~pi1154 & ~n42205;
  assign n42207 = ~n42201 & n42206;
  assign n42208 = ~pi211 & ~n42207;
  assign n42209 = ~n42204 & n42208;
  assign n42210 = ~n42197 & ~n42209;
  assign n42211 = ~pi267 & n42210;
  assign n42212 = n41306 & n42179;
  assign n42213 = pi1154 & ~n42212;
  assign n42214 = ~pi1153 & n39979;
  assign n42215 = ~n39985 & ~n42214;
  assign n42216 = ~pi1155 & ~n42215;
  assign n42217 = n39960 & n42216;
  assign n42218 = n42213 & ~n42217;
  assign n42219 = ~pi1153 & n41272;
  assign n42220 = ~pi1154 & ~n42219;
  assign n42221 = ~n40016 & n42220;
  assign n42222 = ~pi1155 & ~n42221;
  assign n42223 = ~n39904 & n42220;
  assign n42224 = ~n42222 & n42223;
  assign n42225 = ~n42218 & ~n42224;
  assign n42226 = pi211 & ~n42225;
  assign n42227 = ~n39978 & ~n41539;
  assign n42228 = ~n42180 & ~n42227;
  assign n42229 = pi1155 & n42228;
  assign n42230 = pi1154 & n42215;
  assign n42231 = n42222 & ~n42230;
  assign n42232 = ~pi211 & ~n42231;
  assign n42233 = ~n42229 & n42232;
  assign n42234 = pi267 & ~n42233;
  assign n42235 = ~n42226 & n42234;
  assign n42236 = ~pi219 & ~n42235;
  assign n42237 = ~n42211 & n42236;
  assign n42238 = ~n42185 & ~n42237;
  assign n42239 = n39788 & ~n42238;
  assign n42240 = ~n42154 & ~n42239;
  assign n42241 = ~po1038 & n42240;
  assign n42242 = pi267 & n41487;
  assign n42243 = n39788 & ~n42242;
  assign n42244 = ~pi267 & ~n39876;
  assign n42245 = ~n41286 & n42244;
  assign n42246 = n42243 & ~n42245;
  assign n42247 = ~pi219 & ~n37604;
  assign n42248 = ~n37611 & n42247;
  assign n42249 = ~n38346 & ~n42248;
  assign n42250 = pi1091 & ~n42249;
  assign n42251 = ~pi267 & ~pi1091;
  assign n42252 = ~n39788 & n42251;
  assign n42253 = ~n42250 & ~n42252;
  assign n42254 = ~n42246 & n42253;
  assign n42255 = po1038 & ~n42254;
  assign n42256 = n40049 & ~n42255;
  assign n42257 = ~n42241 & n42256;
  assign n42258 = ~po1038 & n42153;
  assign n42259 = ~n42250 & ~n42251;
  assign n42260 = po1038 & ~n42259;
  assign n42261 = ~n40049 & ~n42260;
  assign n42262 = ~n42258 & n42261;
  assign n42263 = ~pi230 & ~n42262;
  assign n42264 = ~n42257 & n42263;
  assign n42265 = pi219 & ~n38084;
  assign n42266 = ~pi1155 & n38150;
  assign n42267 = ~pi1154 & ~n42266;
  assign n42268 = ~n38068 & ~n42267;
  assign n42269 = n37771 & ~n38079;
  assign n42270 = pi1155 & n42269;
  assign n42271 = ~n42268 & ~n42270;
  assign n42272 = ~n42265 & ~n42271;
  assign n42273 = pi211 & ~n42272;
  assign n42274 = ~pi219 & n42128;
  assign n42275 = ~pi199 & pi1154;
  assign n42276 = pi200 & ~n42275;
  assign n42277 = ~n37739 & ~n42276;
  assign n42278 = ~n38083 & n42277;
  assign n42279 = ~n37647 & ~n42278;
  assign n42280 = pi219 & ~n42279;
  assign n42281 = ~pi211 & ~n42280;
  assign n42282 = ~n42274 & n42281;
  assign n42283 = ~n42273 & ~n42282;
  assign n42284 = ~po1038 & n42283;
  assign n42285 = po1038 & n42249;
  assign n42286 = pi230 & ~n42285;
  assign n42287 = ~n42284 & n42286;
  assign po424 = ~n42264 & ~n42287;
  assign n42289 = ~pi199 & n15973;
  assign n42290 = ~n40608 & ~n42289;
  assign n42291 = ~pi211 & ~n15973;
  assign n42292 = ~po1038 & n37771;
  assign n42293 = ~n42291 & ~n42292;
  assign n42294 = pi1152 & ~n42293;
  assign n42295 = n42290 & ~n42294;
  assign n42296 = ~pi1151 & n42293;
  assign n42297 = pi1150 & ~n42296;
  assign n42298 = ~n42295 & n42297;
  assign n42299 = pi1152 & n42298;
  assign n42300 = pi1091 & ~n42299;
  assign n42301 = pi268 & ~n42300;
  assign n42302 = ~po1038 & ~n11225;
  assign n42303 = po1038 & n11223;
  assign n42304 = ~n42302 & ~n42303;
  assign n42305 = pi1151 & ~n42304;
  assign n42306 = ~pi1152 & ~n42305;
  assign n42307 = ~pi1151 & n41217;
  assign n42308 = ~n15973 & n41427;
  assign n42309 = ~po1038 & n37738;
  assign n42310 = ~n42308 & ~n42309;
  assign n42311 = pi1151 & ~n42310;
  assign n42312 = pi1152 & n42311;
  assign n42313 = ~pi1150 & ~n42312;
  assign n42314 = ~n42307 & n42313;
  assign n42315 = ~n42306 & n42314;
  assign n42316 = ~n42298 & ~n42315;
  assign n42317 = pi1091 & ~n42316;
  assign n42318 = ~n42301 & ~n42317;
  assign n42319 = ~n40048 & ~n42318;
  assign n42320 = ~n41297 & n41331;
  assign n42321 = ~po1038 & ~n41257;
  assign n42322 = pi219 & ~n41268;
  assign n42323 = ~n39888 & n42322;
  assign n42324 = ~pi219 & n40008;
  assign n42325 = n41255 & n42324;
  assign n42326 = ~n42323 & ~n42325;
  assign n42327 = n42321 & n42326;
  assign n42328 = ~n42320 & ~n42327;
  assign n42329 = ~pi1151 & ~n42328;
  assign n42330 = ~po1038 & ~n41261;
  assign n42331 = pi219 & n39933;
  assign n42332 = n42330 & ~n42331;
  assign n42333 = n41331 & ~n41486;
  assign n42334 = ~n42332 & ~n42333;
  assign n42335 = pi1151 & ~n42334;
  assign n42336 = ~n42329 & ~n42335;
  assign n42337 = pi268 & ~n42336;
  assign n42338 = n41287 & ~n41328;
  assign n42339 = po1038 & ~n41485;
  assign n42340 = ~n41291 & n42339;
  assign n42341 = n42338 & ~n42340;
  assign n42342 = pi219 & ~n39892;
  assign n42343 = ~n41305 & ~n42342;
  assign n42344 = ~n39893 & ~n42343;
  assign n42345 = ~po1038 & ~n39923;
  assign n42346 = n42344 & n42345;
  assign n42347 = ~n42341 & ~n42346;
  assign n42348 = ~pi1151 & n42347;
  assign n42349 = ~n39865 & ~n42334;
  assign n42350 = ~n39938 & n42330;
  assign n42351 = po1038 & n41285;
  assign n42352 = ~n41283 & ~n42351;
  assign n42353 = ~n42350 & n42352;
  assign n42354 = ~n42349 & ~n42353;
  assign n42355 = pi1151 & n42354;
  assign n42356 = ~pi268 & ~n42355;
  assign n42357 = ~n42348 & n42356;
  assign n42358 = ~n42337 & ~n42357;
  assign n42359 = ~pi1152 & ~n42358;
  assign n42360 = ~n39861 & n42321;
  assign n42361 = ~n42332 & ~n42360;
  assign n42362 = ~n41486 & n42339;
  assign n42363 = n42361 & ~n42362;
  assign n42364 = pi1151 & ~n42363;
  assign n42365 = ~n41297 & n42339;
  assign n42366 = ~n39953 & ~n41354;
  assign n42367 = ~n42326 & ~n42366;
  assign n42368 = ~po1038 & ~n42367;
  assign n42369 = ~n39891 & ~n41599;
  assign n42370 = n42368 & ~n42369;
  assign n42371 = ~n42365 & ~n42370;
  assign n42372 = ~pi1151 & ~n42371;
  assign n42373 = ~n42364 & ~n42372;
  assign n42374 = pi268 & n42373;
  assign n42375 = ~n42322 & ~n42324;
  assign n42376 = ~po1038 & ~n42375;
  assign n42377 = n41287 & ~n41298;
  assign n42378 = ~n42341 & ~n42377;
  assign n42379 = ~n42376 & n42378;
  assign n42380 = pi1151 & ~n42379;
  assign n42381 = ~n41267 & ~n42344;
  assign n42382 = ~po1038 & ~n42381;
  assign n42383 = ~n42338 & ~n42382;
  assign n42384 = ~pi1151 & ~n42383;
  assign n42385 = ~pi268 & ~n42384;
  assign n42386 = ~n42380 & n42385;
  assign n42387 = pi1152 & ~n42386;
  assign n42388 = ~n42374 & n42387;
  assign n42389 = ~n42359 & ~n42388;
  assign n42390 = pi1150 & ~n42389;
  assign n42391 = ~po1038 & ~n42326;
  assign n42392 = ~n42377 & ~n42391;
  assign n42393 = pi1151 & ~n42392;
  assign n42394 = ~pi219 & ~n39930;
  assign n42395 = ~n39881 & ~n42394;
  assign n42396 = n42376 & n42395;
  assign n42397 = ~n41288 & ~n42396;
  assign n42398 = ~pi1151 & ~n42397;
  assign n42399 = pi1152 & ~n42398;
  assign n42400 = ~n42393 & n42399;
  assign n42401 = ~n42351 & ~n42368;
  assign n42402 = ~n41299 & n42401;
  assign n42403 = pi1151 & n42402;
  assign n42404 = ~pi1151 & n42353;
  assign n42405 = ~pi1152 & ~n42404;
  assign n42406 = ~n42403 & n42405;
  assign n42407 = ~n42400 & ~n42406;
  assign n42408 = ~pi268 & ~n42407;
  assign n42409 = ~n41329 & n42339;
  assign n42410 = pi219 & ~n41351;
  assign n42411 = ~n41305 & ~n42410;
  assign n42412 = n40013 & ~n42411;
  assign n42413 = ~po1038 & ~n42412;
  assign n42414 = ~n42409 & ~n42413;
  assign n42415 = pi1151 & n42414;
  assign n42416 = ~po1038 & ~n41354;
  assign n42417 = ~n42410 & n42416;
  assign n42418 = ~n42340 & ~n42417;
  assign n42419 = ~pi1151 & n42418;
  assign n42420 = pi1152 & ~n42419;
  assign n42421 = ~n42415 & n42420;
  assign n42422 = n39865 & ~n42334;
  assign n42423 = ~pi1151 & ~n42422;
  assign n42424 = ~po1038 & ~n41305;
  assign n42425 = ~n41311 & n42424;
  assign n42426 = ~n41332 & ~n42425;
  assign n42427 = pi1151 & n42426;
  assign n42428 = ~pi1152 & ~n42427;
  assign n42429 = ~n42423 & n42428;
  assign n42430 = ~n42421 & ~n42429;
  assign n42431 = pi268 & n42430;
  assign n42432 = ~pi1150 & ~n42431;
  assign n42433 = ~n42408 & n42432;
  assign n42434 = ~n42390 & ~n42433;
  assign n42435 = n40048 & ~n42434;
  assign n42436 = ~n42319 & ~n42435;
  assign n42437 = ~pi230 & ~n42436;
  assign n42438 = pi230 & ~n42316;
  assign po425 = n42437 | n42438;
  assign n42440 = ~pi199 & pi1137;
  assign n42441 = pi200 & ~n42440;
  assign n42442 = ~pi199 & pi1136;
  assign n42443 = pi199 & pi1138;
  assign n42444 = ~pi200 & ~n42443;
  assign n42445 = ~n42442 & n42444;
  assign n42446 = ~n42441 & ~n42445;
  assign n42447 = n15973 & ~n42446;
  assign n42448 = pi1138 & n10522;
  assign n42449 = ~n15973 & ~n42448;
  assign n42450 = pi211 & pi1137;
  assign n42451 = ~n42025 & ~n42450;
  assign n42452 = ~pi219 & ~n42451;
  assign n42453 = n42449 & ~n42452;
  assign n42454 = ~n42447 & ~n42453;
  assign n42455 = pi230 & ~n42454;
  assign n42456 = pi1091 & ~n42451;
  assign n42457 = n40608 & ~n42456;
  assign n42458 = ~pi200 & pi1091;
  assign n42459 = pi1136 & n42458;
  assign n42460 = pi1137 & n39824;
  assign n42461 = ~n42459 & ~n42460;
  assign n42462 = n42289 & n42461;
  assign n42463 = ~n42457 & ~n42462;
  assign n42464 = pi269 & ~n39870;
  assign n42465 = ~pi817 & n39870;
  assign n42466 = ~pi1091 & ~n42465;
  assign n42467 = ~n42464 & n42466;
  assign n42468 = ~n42463 & ~n42467;
  assign n42469 = pi269 & ~n39858;
  assign n42470 = ~pi817 & n39858;
  assign n42471 = ~pi1091 & ~n42470;
  assign n42472 = ~n42469 & n42471;
  assign n42473 = pi219 & ~n15973;
  assign n42474 = pi1138 & n41405;
  assign n42475 = n42473 & ~n42474;
  assign n42476 = pi1138 & n42458;
  assign n42477 = pi199 & ~n42476;
  assign n42478 = n15973 & n42477;
  assign n42479 = ~n42475 & ~n42478;
  assign n42480 = ~n42472 & ~n42479;
  assign n42481 = ~n42468 & ~n42480;
  assign n42482 = ~pi230 & ~n42481;
  assign po426 = ~n42455 & ~n42482;
  assign n42484 = pi270 & ~n39870;
  assign n42485 = ~pi805 & n39870;
  assign n42486 = ~pi1091 & ~n42485;
  assign n42487 = ~n42484 & n42486;
  assign n42488 = ~pi211 & pi1139;
  assign n42489 = pi211 & pi1140;
  assign n42490 = ~n42488 & ~n42489;
  assign n42491 = pi1091 & ~n42490;
  assign n42492 = n40608 & ~n42491;
  assign n42493 = pi1139 & n42458;
  assign n42494 = pi1091 & pi1140;
  assign n42495 = pi200 & n42494;
  assign n42496 = ~n42493 & ~n42495;
  assign n42497 = n42289 & n42496;
  assign n42498 = ~n42492 & ~n42497;
  assign n42499 = ~n42487 & ~n42498;
  assign n42500 = pi270 & ~n39858;
  assign n42501 = ~pi805 & n39858;
  assign n42502 = ~pi1091 & ~n42501;
  assign n42503 = ~n42500 & n42502;
  assign n42504 = pi1091 & n41977;
  assign n42505 = n42473 & ~n42504;
  assign n42506 = ~pi200 & n41947;
  assign n42507 = pi199 & ~n42506;
  assign n42508 = n15973 & n42507;
  assign n42509 = ~n42505 & ~n42508;
  assign n42510 = ~n42503 & ~n42509;
  assign n42511 = ~pi230 & ~n42510;
  assign n42512 = ~n42499 & n42511;
  assign n42513 = ~pi199 & pi1140;
  assign n42514 = pi200 & ~n42513;
  assign n42515 = ~pi199 & pi1139;
  assign n42516 = pi199 & pi1141;
  assign n42517 = ~pi200 & ~n42516;
  assign n42518 = ~n42515 & n42517;
  assign n42519 = ~n42514 & ~n42518;
  assign n42520 = n15973 & ~n42519;
  assign n42521 = pi1141 & n10522;
  assign n42522 = ~pi219 & ~n42490;
  assign n42523 = ~n15973 & ~n42522;
  assign n42524 = ~n42521 & n42523;
  assign n42525 = pi230 & ~n42524;
  assign n42526 = ~n42520 & n42525;
  assign po427 = n42512 | n42526;
  assign n42528 = ~pi271 & ~n39889;
  assign n42529 = ~n39862 & ~n42528;
  assign n42530 = pi199 & ~n42529;
  assign n42531 = pi1091 & pi1146;
  assign n42532 = ~n39873 & ~n42529;
  assign n42533 = ~n39874 & ~n42532;
  assign n42534 = ~n42531 & ~n42533;
  assign n42535 = ~pi199 & n42534;
  assign n42536 = ~n42530 & ~n42535;
  assign n42537 = pi200 & ~n42536;
  assign n42538 = pi1091 & pi1145;
  assign n42539 = ~pi199 & ~n42538;
  assign n42540 = ~n42533 & n42539;
  assign n42541 = ~n42530 & ~n42540;
  assign n42542 = pi1147 & n39810;
  assign n42543 = ~pi200 & ~n42542;
  assign n42544 = ~n42541 & n42543;
  assign n42545 = ~n42537 & ~n42544;
  assign n42546 = n15973 & ~n42545;
  assign n42547 = pi219 & ~n42529;
  assign n42548 = ~pi211 & n42531;
  assign n42549 = ~n42534 & ~n42548;
  assign n42550 = pi1091 & n38489;
  assign n42551 = ~pi219 & ~n42550;
  assign n42552 = ~n42549 & n42551;
  assign n42553 = ~n42547 & ~n42552;
  assign n42554 = ~pi211 & pi1147;
  assign n42555 = n41281 & n42554;
  assign n42556 = ~n15973 & ~n42555;
  assign n42557 = ~n42553 & n42556;
  assign n42558 = ~n42546 & ~n42557;
  assign n42559 = ~pi230 & ~n42558;
  assign n42560 = ~n39204 & ~n39217;
  assign n42561 = ~pi219 & ~n42560;
  assign n42562 = pi1147 & n41214;
  assign n42563 = ~pi200 & ~n38471;
  assign n42564 = n39323 & ~n42563;
  assign n42565 = ~n42562 & ~n42564;
  assign n42566 = ~n42561 & n42565;
  assign n42567 = ~po1038 & ~n42566;
  assign n42568 = pi219 & ~n42554;
  assign n42569 = po1038 & ~n42568;
  assign n42570 = ~n38489 & n40276;
  assign n42571 = n42569 & ~n42570;
  assign n42572 = pi230 & ~n42571;
  assign n42573 = ~n42567 & n42572;
  assign po428 = ~n42559 & ~n42573;
  assign n42575 = pi1150 & ~n42379;
  assign n42576 = ~pi1150 & ~n42354;
  assign n42577 = pi1149 & ~n42576;
  assign n42578 = ~n42575 & n42577;
  assign n42579 = pi1150 & ~n42383;
  assign n42580 = ~pi1150 & ~n42347;
  assign n42581 = ~pi1149 & ~n42580;
  assign n42582 = ~n42579 & n42581;
  assign n42583 = ~n42578 & ~n42582;
  assign n42584 = pi1148 & ~n42583;
  assign n42585 = pi1150 & n42392;
  assign n42586 = ~pi1150 & ~n42402;
  assign n42587 = ~n42585 & ~n42586;
  assign n42588 = pi1149 & n42587;
  assign n42589 = ~pi1150 & ~n42353;
  assign n42590 = pi1150 & n42397;
  assign n42591 = ~pi1149 & ~n42590;
  assign n42592 = ~n42589 & n42591;
  assign n42593 = ~pi1148 & ~n42592;
  assign n42594 = ~n42588 & n42593;
  assign n42595 = ~n42584 & ~n42594;
  assign n42596 = pi283 & ~n42595;
  assign n42597 = pi1150 & ~n41217;
  assign n42598 = ~pi1149 & ~n42597;
  assign n42599 = ~pi1148 & ~n42598;
  assign n42600 = ~pi1150 & ~n42304;
  assign n42601 = pi1149 & ~pi1150;
  assign n42602 = pi1149 & ~n42310;
  assign n42603 = ~n42601 & ~n42602;
  assign n42604 = ~n42600 & ~n42603;
  assign n42605 = n42599 & ~n42604;
  assign n42606 = ~pi219 & n38421;
  assign n42607 = ~n12747 & ~n42606;
  assign n42608 = ~pi1150 & n42607;
  assign n42609 = ~n42293 & ~n42608;
  assign n42610 = ~pi1149 & ~n42609;
  assign n42611 = ~n42293 & ~n42601;
  assign n42612 = n42290 & ~n42611;
  assign n42613 = ~n42610 & ~n42612;
  assign n42614 = pi1148 & n42613;
  assign n42615 = ~n42605 & ~n42614;
  assign n42616 = pi1091 & ~n42615;
  assign n42617 = ~pi283 & ~n42616;
  assign n42618 = ~n42596 & ~n42617;
  assign n42619 = ~pi272 & n42618;
  assign n42620 = pi1150 & n42363;
  assign n42621 = ~pi1150 & n42334;
  assign n42622 = pi1149 & ~n42621;
  assign n42623 = ~n42620 & n42622;
  assign n42624 = pi1150 & n42371;
  assign n42625 = ~pi1150 & n42328;
  assign n42626 = ~pi1149 & ~n42625;
  assign n42627 = ~n42624 & n42626;
  assign n42628 = ~n42623 & ~n42627;
  assign n42629 = pi1148 & ~n42628;
  assign n42630 = pi1150 & n42418;
  assign n42631 = ~pi1150 & ~n42422;
  assign n42632 = ~pi1149 & ~n42631;
  assign n42633 = ~n42630 & n42632;
  assign n42634 = pi1150 & n42414;
  assign n42635 = ~pi1150 & n42426;
  assign n42636 = ~n42634 & ~n42635;
  assign n42637 = pi1149 & n42636;
  assign n42638 = ~n42633 & ~n42637;
  assign n42639 = ~pi1148 & ~n42638;
  assign n42640 = pi283 & ~n42639;
  assign n42641 = ~n42629 & n42640;
  assign n42642 = pi1091 & n42617;
  assign n42643 = ~n42641 & ~n42642;
  assign n42644 = pi272 & n42643;
  assign n42645 = ~pi230 & ~n42644;
  assign n42646 = ~n42619 & n42645;
  assign n42647 = pi230 & n42615;
  assign po429 = ~n42646 & ~n42647;
  assign n42649 = ~pi273 & ~n39890;
  assign n42650 = ~n39864 & ~n42649;
  assign n42651 = pi219 & ~n42650;
  assign n42652 = ~n39874 & ~n42650;
  assign n42653 = ~n39875 & ~n42652;
  assign n42654 = ~pi219 & ~n42548;
  assign n42655 = ~n42653 & n42654;
  assign n42656 = ~n42651 & ~n42655;
  assign n42657 = pi299 & n42656;
  assign n42658 = pi199 & ~n42650;
  assign n42659 = ~pi299 & ~n42658;
  assign n42660 = ~pi200 & n42531;
  assign n42661 = ~pi199 & ~n42660;
  assign n42662 = ~n42653 & n42661;
  assign n42663 = n42659 & ~n42662;
  assign n42664 = ~n42657 & ~n42663;
  assign n42665 = n39400 & ~n42664;
  assign n42666 = ~pi1148 & ~n42665;
  assign n42667 = ~n41370 & ~n42656;
  assign n42668 = pi299 & ~n42667;
  assign n42669 = n39811 & ~n42537;
  assign n42670 = ~n42668 & ~n42669;
  assign n42671 = ~n42663 & n42670;
  assign n42672 = ~po1038 & ~n42671;
  assign n42673 = n38421 & n41281;
  assign n42674 = ~n42672 & ~n42673;
  assign n42675 = pi1148 & n42674;
  assign n42676 = ~n42666 & ~n42675;
  assign n42677 = po1038 & n42656;
  assign n42678 = ~n11224 & ~n39926;
  assign n42679 = pi1091 & ~n42678;
  assign n42680 = n42664 & ~n42679;
  assign n42681 = ~po1038 & ~n42680;
  assign n42682 = pi1091 & n41332;
  assign n42683 = ~n42681 & ~n42682;
  assign n42684 = pi1147 & ~n42683;
  assign n42685 = ~n42677 & ~n42684;
  assign n42686 = ~n42676 & n42685;
  assign n42687 = ~pi230 & ~n42686;
  assign n42688 = ~pi1146 & n41223;
  assign n42689 = pi1147 & n40608;
  assign n42690 = ~n42291 & ~n42689;
  assign n42691 = ~n42688 & ~n42690;
  assign n42692 = pi1148 & ~n42691;
  assign n42693 = ~pi1146 & n10614;
  assign n42694 = ~pi199 & pi1147;
  assign n42695 = pi200 & ~n42694;
  assign n42696 = ~n42693 & ~n42695;
  assign n42697 = n15973 & n42696;
  assign n42698 = n42692 & ~n42697;
  assign n42699 = ~pi211 & ~n39216;
  assign n42700 = n40608 & ~n42699;
  assign n42701 = n42289 & ~n42693;
  assign n42702 = ~n42700 & ~n42701;
  assign n42703 = pi1147 & ~n42702;
  assign n42704 = ~n40298 & ~n42607;
  assign n42705 = pi1146 & n42704;
  assign n42706 = ~pi1148 & ~n42705;
  assign n42707 = ~n42703 & n42706;
  assign n42708 = pi230 & ~n42707;
  assign n42709 = ~n42698 & n42708;
  assign po430 = n42687 | n42709;
  assign n42711 = pi274 & ~n39858;
  assign n42712 = ~pi659 & n39858;
  assign n42713 = ~pi1091 & ~n42712;
  assign n42714 = ~n42711 & n42713;
  assign n42715 = ~pi200 & n42538;
  assign n42716 = ~n42714 & ~n42715;
  assign n42717 = pi199 & n42716;
  assign n42718 = pi274 & ~n39870;
  assign n42719 = ~pi659 & n39870;
  assign n42720 = ~pi1091 & ~n42719;
  assign n42721 = ~n42718 & n42720;
  assign n42722 = ~n41962 & ~n42721;
  assign n42723 = ~pi200 & ~n42722;
  assign n42724 = ~n42004 & ~n42721;
  assign n42725 = pi200 & ~n42724;
  assign n42726 = ~pi199 & ~n42725;
  assign n42727 = ~n42723 & n42726;
  assign n42728 = n15973 & ~n42727;
  assign n42729 = ~n42717 & n42728;
  assign n42730 = pi219 & ~n42550;
  assign n42731 = ~n42714 & n42730;
  assign n42732 = pi211 & ~n42724;
  assign n42733 = ~pi211 & ~n42722;
  assign n42734 = ~pi219 & ~n42733;
  assign n42735 = ~n42732 & n42734;
  assign n42736 = ~n15973 & ~n42735;
  assign n42737 = ~n42731 & n42736;
  assign n42738 = ~pi230 & ~n42737;
  assign n42739 = ~n42729 & n42738;
  assign n42740 = ~pi219 & ~n37672;
  assign n42741 = ~n38490 & n42740;
  assign n42742 = ~n39236 & ~n42741;
  assign n42743 = ~n37645 & ~n39204;
  assign n42744 = ~n42741 & ~n42743;
  assign n42745 = ~n37628 & n39330;
  assign n42746 = n39731 & ~n42745;
  assign n42747 = ~n42744 & ~n42746;
  assign n42748 = ~po1038 & ~n42747;
  assign n42749 = pi230 & ~n42748;
  assign n42750 = ~n42742 & n42749;
  assign po431 = ~n42739 & ~n42750;
  assign n42752 = ~pi1149 & n42311;
  assign n42753 = pi1151 & ~n42293;
  assign n42754 = pi1149 & n42290;
  assign n42755 = ~n42753 & n42754;
  assign n42756 = ~n42752 & ~n42755;
  assign n42757 = pi1150 & ~n42756;
  assign n42758 = n42607 & ~n42753;
  assign n42759 = pi1149 & ~n42758;
  assign n42760 = n39688 & ~n41217;
  assign n42761 = ~pi1149 & n42760;
  assign n42762 = ~pi1150 & ~n42761;
  assign n42763 = ~n42759 & n42762;
  assign n42764 = ~n42757 & ~n42763;
  assign n42765 = pi1091 & ~n42764;
  assign n42766 = ~pi1151 & n42304;
  assign n42767 = pi1091 & n40455;
  assign n42768 = n42766 & n42767;
  assign n42769 = ~n42765 & ~n42768;
  assign n42770 = pi275 & ~n42769;
  assign n42771 = ~n42311 & ~n42766;
  assign n42772 = pi1150 & n42771;
  assign n42773 = ~pi1149 & ~n42772;
  assign n42774 = ~n42760 & n42773;
  assign n42775 = n42293 & n42601;
  assign n42776 = ~n42755 & ~n42775;
  assign n42777 = ~n42774 & n42776;
  assign n42778 = pi1091 & n42777;
  assign n42779 = ~pi275 & ~n42778;
  assign n42780 = ~n40047 & ~n42779;
  assign n42781 = ~n42770 & n42780;
  assign n42782 = ~pi1150 & n42418;
  assign n42783 = ~n42634 & ~n42782;
  assign n42784 = pi1151 & ~n42783;
  assign n42785 = pi1150 & n42426;
  assign n42786 = ~n42631 & ~n42785;
  assign n42787 = ~pi1151 & ~n42786;
  assign n42788 = ~n42784 & ~n42787;
  assign n42789 = pi275 & n42788;
  assign n42790 = ~pi1150 & n42397;
  assign n42791 = pi1151 & ~n42585;
  assign n42792 = ~n42790 & n42791;
  assign n42793 = pi1150 & ~n42402;
  assign n42794 = ~pi1151 & ~n42589;
  assign n42795 = ~n42793 & n42794;
  assign n42796 = ~n42792 & ~n42795;
  assign n42797 = ~pi275 & ~n42796;
  assign n42798 = ~pi1149 & ~n42797;
  assign n42799 = ~n42789 & n42798;
  assign n42800 = pi1151 & ~n42371;
  assign n42801 = ~pi1150 & ~n42800;
  assign n42802 = ~n42329 & n42801;
  assign n42803 = ~pi1151 & ~n42334;
  assign n42804 = pi1150 & ~n42364;
  assign n42805 = ~n42803 & n42804;
  assign n42806 = pi275 & ~n42805;
  assign n42807 = ~n42802 & n42806;
  assign n42808 = ~pi1150 & ~n42383;
  assign n42809 = pi1151 & ~n42575;
  assign n42810 = ~n42808 & n42809;
  assign n42811 = pi1150 & ~n42354;
  assign n42812 = ~pi1151 & ~n42811;
  assign n42813 = ~n42580 & n42812;
  assign n42814 = ~pi275 & ~n42813;
  assign n42815 = ~n42810 & n42814;
  assign n42816 = pi1149 & ~n42815;
  assign n42817 = ~n42807 & n42816;
  assign n42818 = n40047 & ~n42817;
  assign n42819 = ~n42799 & n42818;
  assign n42820 = ~n42781 & ~n42819;
  assign n42821 = ~pi230 & ~n42820;
  assign n42822 = pi230 & n42777;
  assign po432 = n42821 | n42822;
  assign n42824 = ~pi276 & ~n39859;
  assign n42825 = n39861 & ~n42824;
  assign n42826 = n42473 & ~n42548;
  assign n42827 = pi199 & ~n42660;
  assign n42828 = n15973 & n42827;
  assign n42829 = ~n42826 & ~n42828;
  assign n42830 = ~n42825 & ~n42829;
  assign n42831 = ~n37667 & ~n39211;
  assign n42832 = pi1091 & ~n42831;
  assign n42833 = n40608 & ~n42832;
  assign n42834 = pi1145 & n39824;
  assign n42835 = ~n42005 & ~n42834;
  assign n42836 = n42289 & n42835;
  assign n42837 = ~n42833 & ~n42836;
  assign n42838 = ~pi276 & ~n39871;
  assign n42839 = ~pi1091 & ~n39872;
  assign n42840 = ~n42838 & n42839;
  assign n42841 = ~n42837 & ~n42840;
  assign n42842 = ~pi230 & ~n42841;
  assign n42843 = ~n42830 & n42842;
  assign n42844 = pi219 & n39210;
  assign n42845 = ~pi219 & ~n42831;
  assign n42846 = ~n15973 & ~n42845;
  assign n42847 = ~n42844 & n42846;
  assign n42848 = ~n37626 & n40192;
  assign n42849 = ~n39328 & ~n42848;
  assign n42850 = n15973 & ~n42849;
  assign n42851 = pi230 & ~n42850;
  assign n42852 = ~n42847 & n42851;
  assign po433 = n42843 | n42852;
  assign n42854 = pi219 & ~n37694;
  assign n42855 = ~n41940 & ~n42854;
  assign n42856 = pi277 & ~n39858;
  assign n42857 = ~pi820 & n39858;
  assign n42858 = ~pi1091 & ~n42857;
  assign n42859 = ~n42856 & n42858;
  assign n42860 = ~n42855 & ~n42859;
  assign n42861 = pi277 & ~n39870;
  assign n42862 = ~pi820 & n39870;
  assign n42863 = ~pi1091 & ~n42862;
  assign n42864 = ~n42861 & n42863;
  assign n42865 = ~n42494 & ~n42864;
  assign n42866 = ~pi211 & ~n42865;
  assign n42867 = ~n41947 & ~n42864;
  assign n42868 = pi211 & ~n42867;
  assign n42869 = ~pi219 & ~n42868;
  assign n42870 = ~n42866 & n42869;
  assign n42871 = ~n42860 & ~n42870;
  assign n42872 = ~n15973 & ~n42871;
  assign n42873 = ~pi230 & ~n42872;
  assign n42874 = ~pi200 & n41954;
  assign n42875 = pi199 & ~n42859;
  assign n42876 = ~n42874 & n42875;
  assign n42877 = ~pi200 & ~n42865;
  assign n42878 = pi200 & ~n42867;
  assign n42879 = ~pi199 & ~n42878;
  assign n42880 = ~n42877 & n42879;
  assign n42881 = ~n42876 & ~n42880;
  assign n42882 = n15973 & ~n42881;
  assign n42883 = n42873 & ~n42882;
  assign n42884 = n37625 & ~n42513;
  assign n42885 = pi200 & ~n41973;
  assign n42886 = ~n42884 & ~n42885;
  assign n42887 = n15973 & ~n42886;
  assign n42888 = ~pi211 & pi1140;
  assign n42889 = pi211 & pi1141;
  assign n42890 = ~pi219 & ~n42889;
  assign n42891 = ~n42888 & n42890;
  assign n42892 = ~n42854 & ~n42891;
  assign n42893 = ~n15973 & ~n42892;
  assign n42894 = pi230 & ~n42893;
  assign n42895 = ~n42887 & n42894;
  assign po434 = n42883 | n42895;
  assign n42897 = ~pi976 & n39858;
  assign n42898 = ~pi278 & ~n39858;
  assign n42899 = ~pi1091 & ~n42898;
  assign n42900 = ~n42897 & n42899;
  assign n42901 = pi199 & ~n42900;
  assign n42902 = pi1091 & ~pi1132;
  assign n42903 = pi278 & ~n39870;
  assign n42904 = pi976 & n39870;
  assign n42905 = ~pi1091 & ~n42904;
  assign n42906 = ~n42903 & n42905;
  assign n42907 = ~n42902 & ~n42906;
  assign n42908 = ~pi199 & ~n42907;
  assign n42909 = ~n42901 & ~n42908;
  assign n42910 = ~pi200 & ~n42909;
  assign n42911 = pi1091 & ~pi1133;
  assign n42912 = ~n42906 & ~n42911;
  assign n42913 = ~pi199 & ~n42912;
  assign n42914 = ~n42901 & ~n42913;
  assign n42915 = pi200 & ~n42914;
  assign n42916 = ~pi299 & ~n42915;
  assign n42917 = ~n42910 & n42916;
  assign n42918 = pi219 & ~n42900;
  assign n42919 = pi211 & ~pi1133;
  assign n42920 = ~pi211 & ~pi1132;
  assign n42921 = ~n42919 & ~n42920;
  assign n42922 = pi1091 & ~n42921;
  assign n42923 = ~n42906 & ~n42922;
  assign n42924 = ~pi219 & ~n42923;
  assign n42925 = ~n42918 & ~n42924;
  assign n42926 = pi299 & n42925;
  assign n42927 = ~n42917 & ~n42926;
  assign n42928 = ~po1038 & ~n42927;
  assign n42929 = po1038 & n42925;
  assign n42930 = ~pi230 & ~n42929;
  assign n42931 = ~n42928 & n42930;
  assign n42932 = ~pi199 & pi1132;
  assign n42933 = ~pi200 & ~n42932;
  assign n42934 = ~pi199 & pi1133;
  assign n42935 = pi200 & ~n42934;
  assign n42936 = ~pi299 & ~n42935;
  assign n42937 = ~n42933 & n42936;
  assign n42938 = n37645 & n42921;
  assign n42939 = ~n42937 & ~n42938;
  assign n42940 = ~po1038 & ~n42939;
  assign n42941 = n38420 & n42921;
  assign n42942 = ~n42940 & ~n42941;
  assign n42943 = pi230 & n42942;
  assign n42944 = ~n42931 & ~n42943;
  assign n42945 = ~pi1134 & ~n42944;
  assign n42946 = n10614 & ~n42932;
  assign n42947 = n42936 & ~n42946;
  assign n42948 = ~n41442 & ~n42938;
  assign n42949 = ~n42947 & n42948;
  assign n42950 = ~po1038 & ~n42949;
  assign n42951 = pi230 & ~n42950;
  assign n42952 = ~n41216 & ~n42941;
  assign n42953 = n42951 & n42952;
  assign n42954 = ~n39810 & n42910;
  assign n42955 = n42916 & ~n42954;
  assign n42956 = n12744 & n41405;
  assign n42957 = ~n42926 & ~n42956;
  assign n42958 = ~n42955 & n42957;
  assign n42959 = ~po1038 & ~n42958;
  assign n42960 = ~n42673 & ~n42959;
  assign n42961 = n42930 & n42960;
  assign n42962 = ~n42953 & ~n42961;
  assign n42963 = pi1134 & ~n42962;
  assign po435 = ~n42945 & ~n42963;
  assign n42965 = ~pi958 & n39858;
  assign n42966 = ~pi279 & ~n39858;
  assign n42967 = ~pi1091 & ~n42966;
  assign n42968 = ~n42965 & n42967;
  assign n42969 = pi1135 & n42458;
  assign n42970 = ~n42968 & ~n42969;
  assign n42971 = pi199 & ~n42970;
  assign n42972 = pi279 & ~n39870;
  assign n42973 = pi958 & n39870;
  assign n42974 = ~pi1091 & ~n42973;
  assign n42975 = ~n42972 & n42974;
  assign n42976 = ~pi1133 & n42458;
  assign n42977 = ~pi199 & ~n42976;
  assign n42978 = ~n42975 & n42977;
  assign n42979 = ~n42971 & ~n42978;
  assign n42980 = n15973 & ~n42979;
  assign n42981 = ~n39824 & n42980;
  assign n42982 = ~n41383 & ~n42975;
  assign n42983 = ~n42911 & n42982;
  assign n42984 = ~pi219 & ~n42983;
  assign n42985 = pi1135 & n41405;
  assign n42986 = ~n42968 & ~n42985;
  assign n42987 = pi219 & n42986;
  assign n42988 = ~n15973 & ~n42987;
  assign n42989 = ~n42984 & n42988;
  assign n42990 = ~pi230 & ~n42989;
  assign n42991 = ~n42981 & n42990;
  assign n42992 = pi199 & pi1135;
  assign n42993 = ~n42934 & ~n42992;
  assign n42994 = n37771 & ~n42993;
  assign n42995 = pi1135 & n10522;
  assign n42996 = ~pi211 & ~pi1133;
  assign n42997 = ~pi219 & ~n42996;
  assign n42998 = ~pi211 & n42997;
  assign n42999 = ~n42995 & ~n42998;
  assign n43000 = pi299 & ~n42999;
  assign n43001 = ~n42994 & ~n43000;
  assign n43002 = ~po1038 & ~n43001;
  assign n43003 = po1038 & ~n42999;
  assign n43004 = pi230 & ~n43003;
  assign n43005 = ~n43002 & n43004;
  assign n43006 = ~n42991 & ~n43005;
  assign n43007 = ~pi1134 & ~n43006;
  assign n43008 = ~pi1133 & n10614;
  assign n43009 = ~pi200 & pi1135;
  assign n43010 = pi199 & ~n43009;
  assign n43011 = ~n43008 & ~n43010;
  assign n43012 = n15973 & ~n43011;
  assign n43013 = ~n15973 & ~n42997;
  assign n43014 = ~n42995 & n43013;
  assign n43015 = ~n43012 & ~n43014;
  assign n43016 = pi230 & ~n43015;
  assign n43017 = pi1091 & ~n42996;
  assign n43018 = n40608 & n43017;
  assign n43019 = ~n42980 & ~n43018;
  assign n43020 = n42990 & n43019;
  assign n43021 = ~n43016 & ~n43020;
  assign n43022 = pi1134 & ~n43021;
  assign po436 = ~n43007 & ~n43022;
  assign n43024 = ~pi211 & pi1135;
  assign n43025 = pi211 & pi1136;
  assign n43026 = ~n43024 & ~n43025;
  assign n43027 = pi1091 & n43026;
  assign n43028 = pi914 & n39870;
  assign n43029 = ~pi280 & ~n39870;
  assign n43030 = ~pi1091 & ~n43029;
  assign n43031 = ~n43028 & n43030;
  assign n43032 = ~n43027 & ~n43031;
  assign n43033 = ~pi219 & ~n43032;
  assign n43034 = ~pi211 & pi1137;
  assign n43035 = pi219 & ~n43034;
  assign n43036 = ~n41940 & ~n43035;
  assign n43037 = pi280 & ~n39858;
  assign n43038 = ~pi914 & n39858;
  assign n43039 = ~pi1091 & ~n43038;
  assign n43040 = ~n43037 & n43039;
  assign n43041 = ~n43036 & ~n43040;
  assign n43042 = ~n43033 & ~n43041;
  assign n43043 = ~n15973 & ~n43042;
  assign n43044 = pi1137 & n42458;
  assign n43045 = ~n43040 & ~n43044;
  assign n43046 = pi199 & ~n43045;
  assign n43047 = n15973 & ~n43046;
  assign n43048 = pi200 & pi1136;
  assign n43049 = ~n43009 & ~n43048;
  assign n43050 = pi1091 & n43049;
  assign n43051 = ~pi199 & ~n43050;
  assign n43052 = ~n43031 & n43051;
  assign n43053 = n43047 & ~n43052;
  assign n43054 = ~n43043 & ~n43053;
  assign n43055 = ~pi230 & ~n43054;
  assign n43056 = ~pi219 & n43026;
  assign n43057 = ~n43035 & ~n43056;
  assign n43058 = ~n15973 & n43057;
  assign n43059 = pi200 & ~n42442;
  assign n43060 = pi199 & pi1137;
  assign n43061 = ~pi200 & ~n42033;
  assign n43062 = ~n43060 & n43061;
  assign n43063 = n15973 & ~n43062;
  assign n43064 = ~n43059 & n43063;
  assign n43065 = pi230 & ~n43064;
  assign n43066 = ~n43058 & n43065;
  assign po437 = ~n43055 & ~n43066;
  assign n43068 = ~pi199 & pi1138;
  assign n43069 = pi200 & ~n43068;
  assign n43070 = pi199 & pi1139;
  assign n43071 = ~pi200 & ~n42440;
  assign n43072 = ~n43070 & n43071;
  assign n43073 = ~n43069 & ~n43072;
  assign n43074 = n15973 & ~n43073;
  assign n43075 = pi1139 & n10522;
  assign n43076 = ~n15973 & ~n43075;
  assign n43077 = pi211 & pi1138;
  assign n43078 = ~n43034 & ~n43077;
  assign n43079 = ~pi219 & ~n43078;
  assign n43080 = n43076 & ~n43079;
  assign n43081 = ~n43074 & ~n43080;
  assign n43082 = pi230 & ~n43081;
  assign n43083 = pi281 & ~n39870;
  assign n43084 = ~pi830 & n39870;
  assign n43085 = ~pi1091 & ~n43084;
  assign n43086 = ~n43083 & n43085;
  assign n43087 = pi1091 & ~n43078;
  assign n43088 = n40608 & ~n43087;
  assign n43089 = pi1138 & n39824;
  assign n43090 = ~n43044 & ~n43089;
  assign n43091 = n42289 & n43090;
  assign n43092 = ~n43088 & ~n43091;
  assign n43093 = ~n43086 & ~n43092;
  assign n43094 = pi281 & ~n39858;
  assign n43095 = ~pi830 & n39858;
  assign n43096 = ~pi1091 & ~n43095;
  assign n43097 = ~n43094 & n43096;
  assign n43098 = pi1139 & n41405;
  assign n43099 = n42473 & ~n43098;
  assign n43100 = pi199 & ~n42493;
  assign n43101 = n15973 & n43100;
  assign n43102 = ~n43099 & ~n43101;
  assign n43103 = ~n43097 & ~n43102;
  assign n43104 = ~n43093 & ~n43103;
  assign n43105 = ~pi230 & ~n43104;
  assign po438 = ~n43082 & ~n43105;
  assign n43107 = pi200 & ~n42515;
  assign n43108 = pi199 & pi1140;
  assign n43109 = ~pi200 & ~n43068;
  assign n43110 = ~n43108 & n43109;
  assign n43111 = ~n43107 & ~n43110;
  assign n43112 = n15973 & ~n43111;
  assign n43113 = pi1140 & n10522;
  assign n43114 = ~n15973 & ~n43113;
  assign n43115 = ~pi211 & pi1138;
  assign n43116 = pi211 & pi1139;
  assign n43117 = ~n43115 & ~n43116;
  assign n43118 = ~pi219 & ~n43117;
  assign n43119 = n43114 & ~n43118;
  assign n43120 = ~n43112 & ~n43119;
  assign n43121 = pi230 & ~n43120;
  assign n43122 = pi282 & ~n39870;
  assign n43123 = ~pi836 & n39870;
  assign n43124 = ~pi1091 & ~n43123;
  assign n43125 = ~n43122 & n43124;
  assign n43126 = pi1091 & ~n43117;
  assign n43127 = n40608 & ~n43126;
  assign n43128 = pi1139 & n39824;
  assign n43129 = ~n42476 & ~n43128;
  assign n43130 = n42289 & n43129;
  assign n43131 = ~n43127 & ~n43130;
  assign n43132 = ~n43125 & ~n43131;
  assign n43133 = pi282 & ~n39858;
  assign n43134 = ~pi836 & n39858;
  assign n43135 = ~pi1091 & ~n43134;
  assign n43136 = ~n43133 & n43135;
  assign n43137 = pi1140 & n41405;
  assign n43138 = n42473 & ~n43137;
  assign n43139 = ~pi200 & n42494;
  assign n43140 = pi199 & ~n43139;
  assign n43141 = n15973 & n43140;
  assign n43142 = ~n43138 & ~n43141;
  assign n43143 = ~n43136 & ~n43142;
  assign n43144 = ~n43132 & ~n43143;
  assign n43145 = ~pi230 & ~n43144;
  assign po439 = ~n43121 & ~n43145;
  assign n43147 = pi1147 & ~n42607;
  assign n43148 = n42602 & ~n43147;
  assign n43149 = pi1147 & ~n42290;
  assign n43150 = ~pi1149 & n42304;
  assign n43151 = ~n43149 & n43150;
  assign n43152 = ~n43148 & ~n43151;
  assign n43153 = pi1148 & n43152;
  assign n43154 = pi1149 & ~n41217;
  assign n43155 = ~n43147 & ~n43154;
  assign n43156 = ~pi1148 & ~n43155;
  assign n43157 = pi230 & ~n43156;
  assign n43158 = ~n43153 & n43157;
  assign n43159 = pi1147 & n42383;
  assign n43160 = ~pi1147 & n42397;
  assign n43161 = pi1149 & ~n43160;
  assign n43162 = ~n43159 & n43161;
  assign n43163 = ~pi1147 & ~n42353;
  assign n43164 = pi1147 & n42347;
  assign n43165 = ~pi1149 & ~n43164;
  assign n43166 = ~n43163 & n43165;
  assign n43167 = ~n43162 & ~n43166;
  assign n43168 = ~pi1148 & n43167;
  assign n43169 = ~pi1147 & n42392;
  assign n43170 = pi1149 & ~n43169;
  assign n43171 = pi1147 & n42379;
  assign n43172 = n43170 & ~n43171;
  assign n43173 = pi1147 & n42354;
  assign n43174 = ~pi1147 & ~n42402;
  assign n43175 = ~pi1149 & ~n43174;
  assign n43176 = ~n43173 & n43175;
  assign n43177 = ~n43172 & ~n43176;
  assign n43178 = pi1148 & n43177;
  assign n43179 = ~pi283 & ~n43178;
  assign n43180 = ~n43168 & n43179;
  assign n43181 = ~pi1147 & n42414;
  assign n43182 = pi1148 & ~n43181;
  assign n43183 = pi1147 & n42363;
  assign n43184 = n43182 & ~n43183;
  assign n43185 = ~pi1147 & n42418;
  assign n43186 = pi1147 & n42371;
  assign n43187 = ~pi1148 & ~n43186;
  assign n43188 = ~n43185 & n43187;
  assign n43189 = pi1149 & ~n43188;
  assign n43190 = ~n43184 & n43189;
  assign n43191 = ~pi1147 & n42426;
  assign n43192 = pi1147 & n42334;
  assign n43193 = ~n43191 & ~n43192;
  assign n43194 = pi1148 & n43193;
  assign n43195 = pi1147 & n42328;
  assign n43196 = ~pi1147 & ~n42422;
  assign n43197 = ~pi1148 & ~n43196;
  assign n43198 = ~n43195 & n43197;
  assign n43199 = ~pi1149 & ~n43198;
  assign n43200 = ~n43194 & n43199;
  assign n43201 = ~n43190 & ~n43200;
  assign n43202 = pi283 & n43201;
  assign n43203 = ~pi230 & ~n43202;
  assign n43204 = ~n43180 & n43203;
  assign po440 = ~n43158 & ~n43204;
  assign n43206 = ~pi284 & ~n41711;
  assign n43207 = ~n39171 & n41711;
  assign n43208 = pi1143 & n43207;
  assign po441 = n43206 | n43208;
  assign n43210 = n2576 & ~n10188;
  assign n43211 = ~n7371 & n43210;
  assign n43212 = pi286 & n43211;
  assign n43213 = pi288 & pi289;
  assign n43214 = n43212 & n43213;
  assign n43215 = pi285 & n43214;
  assign po637 = ~po1038 & n43210;
  assign n43217 = ~pi285 & ~n43214;
  assign n43218 = po637 & ~n43217;
  assign n43219 = ~n43215 & n43218;
  assign n43220 = pi285 & ~pi289;
  assign n43221 = ~pi286 & ~pi288;
  assign n43222 = n7371 & n43221;
  assign n43223 = n43220 & n43222;
  assign n43224 = ~po1038 & n43214;
  assign n43225 = ~n43223 & ~n43224;
  assign n43226 = pi285 & n43225;
  assign n43227 = ~n43219 & ~n43226;
  assign po442 = ~pi793 & ~n43227;
  assign n43229 = ~pi286 & ~n43211;
  assign n43230 = pi288 & ~n43212;
  assign n43231 = ~n43229 & n43230;
  assign n43232 = ~pi288 & ~n7375;
  assign n43233 = n7371 & ~n43210;
  assign n43234 = pi286 & ~n43233;
  assign n43235 = ~pi286 & n43233;
  assign n43236 = ~n43234 & ~n43235;
  assign n43237 = n43232 & ~n43236;
  assign n43238 = ~n43231 & ~n43237;
  assign n43239 = ~po1038 & n43238;
  assign n43240 = n7371 & n43232;
  assign n43241 = ~pi286 & n43240;
  assign n43242 = pi286 & ~n43240;
  assign n43243 = po1038 & ~n43242;
  assign n43244 = ~n43241 & n43243;
  assign n43245 = ~pi793 & ~n43244;
  assign po443 = ~n43239 & n43245;
  assign n43247 = ~pi287 & pi457;
  assign po444 = ~pi332 & ~n43247;
  assign n43249 = pi288 & ~n7371;
  assign n43250 = ~n43240 & ~n43249;
  assign n43251 = ~po637 & n43250;
  assign n43252 = po637 & ~n43250;
  assign n43253 = ~n43251 & ~n43252;
  assign po445 = ~pi793 & n43253;
  assign n43255 = n43220 & n43235;
  assign n43256 = ~pi288 & ~n43255;
  assign n43257 = ~n43230 & ~n43256;
  assign n43258 = ~pi289 & ~n43257;
  assign n43259 = n43235 & n43256;
  assign n43260 = ~n43214 & ~n43259;
  assign n43261 = ~n43258 & n43260;
  assign n43262 = ~po1038 & ~n43261;
  assign n43263 = ~pi793 & ~n43262;
  assign n43264 = pi289 & ~n43222;
  assign n43265 = po1038 & ~n43223;
  assign n43266 = ~n43264 & n43265;
  assign po446 = n43263 & ~n43266;
  assign n43268 = ~pi290 & pi476;
  assign n43269 = ~pi476 & ~pi1048;
  assign po447 = ~n43268 & ~n43269;
  assign n43271 = ~pi291 & pi476;
  assign n43272 = ~pi476 & ~pi1049;
  assign po448 = ~n43271 & ~n43272;
  assign n43274 = ~pi292 & pi476;
  assign n43275 = ~pi476 & ~pi1084;
  assign po449 = ~n43274 & ~n43275;
  assign n43277 = ~pi293 & pi476;
  assign n43278 = ~pi476 & ~pi1059;
  assign po450 = ~n43277 & ~n43278;
  assign n43280 = ~pi294 & pi476;
  assign n43281 = ~pi476 & ~pi1072;
  assign po451 = ~n43280 & ~n43281;
  assign n43283 = ~pi295 & pi476;
  assign n43284 = ~pi476 & ~pi1053;
  assign po452 = ~n43283 & ~n43284;
  assign n43286 = ~pi296 & pi476;
  assign n43287 = ~pi476 & ~pi1037;
  assign po453 = ~n43286 & ~n43287;
  assign n43289 = ~pi297 & pi476;
  assign n43290 = ~pi476 & ~pi1044;
  assign po454 = ~n43289 & ~n43290;
  assign n43292 = ~pi478 & pi1044;
  assign n43293 = pi298 & pi478;
  assign po455 = n43292 | n43293;
  assign n43295 = pi54 & n2522;
  assign n43296 = ~pi54 & n12829;
  assign n43297 = n13082 & n43296;
  assign n43298 = ~n43295 & ~n43297;
  assign n43299 = n2574 & ~n43298;
  assign n43300 = n8738 & n43299;
  assign n43301 = ~pi39 & ~n43300;
  assign po456 = ~n11054 & ~n43301;
  assign n43303 = pi57 & ~pi59;
  assign n43304 = n9966 & n43303;
  assign n43305 = ~pi312 & n43304;
  assign n43306 = pi300 & ~n43305;
  assign n43307 = ~pi300 & n43305;
  assign n43308 = ~pi55 & ~n43307;
  assign po457 = n43306 | ~n43308;
  assign n43310 = ~pi301 & n43308;
  assign n43311 = ~pi300 & pi301;
  assign n43312 = ~pi55 & n43311;
  assign n43313 = n43305 & n43312;
  assign po458 = n43310 | n43313;
  assign n43315 = ~pi215 & n3300;
  assign n43316 = ~pi273 & n43315;
  assign n43317 = ~pi937 & n5746;
  assign n43318 = ~n43316 & ~n43317;
  assign n43319 = ~n15973 & ~n43318;
  assign n43320 = n5793 & ~po1038;
  assign n43321 = ~n2607 & n43320;
  assign n43322 = pi273 & n3332;
  assign n43323 = ~pi222 & ~pi223;
  assign n43324 = pi937 & ~n43323;
  assign n43325 = ~n43322 & ~n43324;
  assign n43326 = n43321 & n43325;
  assign n43327 = ~n5747 & ~n15973;
  assign n43328 = ~n43320 & ~n43327;
  assign n43329 = ~pi1148 & n43328;
  assign n43330 = n2528 & ~n15973;
  assign n43331 = ~po1038 & n12851;
  assign n43332 = ~n43330 & ~n43331;
  assign n43333 = ~n43326 & n43332;
  assign n43334 = pi237 & ~n43333;
  assign n43335 = ~n43329 & ~n43334;
  assign n43336 = ~n43326 & n43335;
  assign po459 = ~n43319 & n43336;
  assign n43338 = ~pi478 & pi1049;
  assign n43339 = pi303 & pi478;
  assign po460 = n43338 | n43339;
  assign n43341 = ~pi478 & pi1048;
  assign n43342 = pi304 & pi478;
  assign po461 = n43341 | n43342;
  assign n43344 = ~pi478 & pi1084;
  assign n43345 = pi305 & pi478;
  assign po462 = n43344 | n43345;
  assign n43347 = ~pi478 & pi1059;
  assign n43348 = pi306 & pi478;
  assign po463 = n43347 | n43348;
  assign n43350 = ~pi478 & pi1053;
  assign n43351 = pi307 & pi478;
  assign po464 = n43350 | n43351;
  assign n43353 = ~pi478 & pi1037;
  assign n43354 = pi308 & pi478;
  assign po465 = n43353 | n43354;
  assign n43356 = ~pi478 & pi1072;
  assign n43357 = pi309 & pi478;
  assign po466 = n43356 | n43357;
  assign n43359 = pi1147 & n43328;
  assign n43360 = ~n2527 & n43327;
  assign n43361 = pi934 & ~n3531;
  assign n43362 = pi271 & n3300;
  assign n43363 = ~n43361 & ~n43362;
  assign n43364 = n43360 & ~n43363;
  assign n43365 = pi222 & ~pi934;
  assign n43366 = ~pi271 & n3332;
  assign n43367 = ~n43365 & ~n43366;
  assign n43368 = n43320 & n43367;
  assign n43369 = ~n43330 & ~n43368;
  assign n43370 = ~n43364 & n43369;
  assign n43371 = ~n43359 & n43370;
  assign n43372 = ~pi233 & ~n43371;
  assign n43373 = n43320 & ~n43367;
  assign n43374 = pi1147 & ~n43331;
  assign n43375 = n43327 & n43363;
  assign n43376 = n43374 & ~n43375;
  assign n43377 = ~n43373 & n43376;
  assign n43378 = ~n43321 & ~n43360;
  assign n43379 = ~pi1147 & ~n43378;
  assign n43380 = ~n43370 & n43379;
  assign n43381 = ~n43377 & ~n43380;
  assign n43382 = pi233 & ~n43381;
  assign po467 = n43372 | n43382;
  assign n43384 = pi311 & ~n43313;
  assign n43385 = ~pi55 & ~n43313;
  assign n43386 = ~pi311 & ~n43385;
  assign po468 = ~n43384 & ~n43386;
  assign n43388 = pi312 & ~n43304;
  assign n43389 = ~n43305 & ~n43388;
  assign po469 = ~pi55 & ~n43389;
  assign n43391 = ~n10175 & ~n13115;
  assign n43392 = po740 & ~n13122;
  assign n43393 = n9988 & ~n43392;
  assign po634 = n43391 | ~n43393;
  assign n43395 = ~pi954 & po634;
  assign n43396 = pi313 & pi954;
  assign po470 = ~n43395 & ~n43396;
  assign n43398 = n2573 & n12806;
  assign n43399 = n14013 & ~n43398;
  assign n43400 = ~pi39 & ~n14083;
  assign n43401 = pi39 & ~n14543;
  assign n43402 = ~n43400 & ~n43401;
  assign n43403 = n2614 & n43402;
  assign n43404 = ~n15405 & ~n43403;
  assign n43405 = n2537 & ~n43404;
  assign n43406 = ~po1038 & n43405;
  assign n43407 = ~n43399 & ~n43406;
  assign n43408 = n14007 & n14008;
  assign po471 = ~n43407 & n43408;
  assign n43410 = ~pi340 & po637;
  assign n43411 = pi315 & ~n43410;
  assign n43412 = pi1080 & n43410;
  assign po472 = n43411 | n43412;
  assign n43414 = pi316 & ~n43410;
  assign n43415 = pi1047 & n43410;
  assign po473 = n43414 | n43415;
  assign n43417 = ~pi330 & po637;
  assign n43418 = pi317 & ~n43417;
  assign n43419 = pi1078 & n43417;
  assign po474 = n43418 | n43419;
  assign n43421 = ~pi341 & po637;
  assign n43422 = pi318 & ~n43421;
  assign n43423 = pi1074 & n43421;
  assign po475 = n43422 | n43423;
  assign n43425 = pi319 & ~n43421;
  assign n43426 = pi1072 & n43421;
  assign po476 = n43425 | n43426;
  assign n43428 = pi320 & ~n43410;
  assign n43429 = pi1048 & n43410;
  assign po477 = n43428 | n43429;
  assign n43431 = pi321 & ~n43410;
  assign n43432 = pi1058 & n43410;
  assign po478 = n43431 | n43432;
  assign n43434 = pi322 & ~n43410;
  assign n43435 = pi1051 & n43410;
  assign po479 = n43434 | n43435;
  assign n43437 = pi323 & ~n43410;
  assign n43438 = pi1065 & n43410;
  assign po480 = n43437 | n43438;
  assign n43440 = pi324 & ~n43421;
  assign n43441 = pi1086 & n43421;
  assign po481 = n43440 | n43441;
  assign n43443 = pi325 & ~n43421;
  assign n43444 = pi1063 & n43421;
  assign po482 = n43443 | n43444;
  assign n43446 = pi326 & ~n43421;
  assign n43447 = pi1057 & n43421;
  assign po483 = n43446 | n43447;
  assign n43449 = pi327 & ~n43410;
  assign n43450 = pi1040 & n43410;
  assign po484 = n43449 | n43450;
  assign n43452 = pi328 & ~n43421;
  assign n43453 = pi1058 & n43421;
  assign po485 = n43452 | n43453;
  assign n43455 = pi329 & ~n43421;
  assign n43456 = pi1043 & n43421;
  assign po486 = n43455 | n43456;
  assign n43458 = pi1092 & ~n6210;
  assign n43459 = po1038 & n43458;
  assign n43460 = pi340 & n43210;
  assign n43461 = ~po1038 & n43458;
  assign n43462 = ~n43460 & n43461;
  assign n43463 = ~n43459 & ~n43462;
  assign n43464 = ~pi330 & ~n43463;
  assign n43465 = n43210 & n43462;
  assign po487 = n43464 | n43465;
  assign n43467 = pi341 & n43210;
  assign n43468 = n43461 & ~n43467;
  assign n43469 = ~n43459 & ~n43468;
  assign n43470 = ~pi331 & ~n43469;
  assign n43471 = n43210 & n43468;
  assign po488 = n43470 | n43471;
  assign n43473 = n10798 & n12844;
  assign n43474 = ~n10798 & ~n12783;
  assign n43475 = n7394 & ~n43474;
  assign n43476 = ~pi70 & ~n43475;
  assign n43477 = pi332 & ~n43476;
  assign n43478 = n9427 & n43477;
  assign n43479 = ~n43473 & ~n43478;
  assign n43480 = ~pi39 & ~n43479;
  assign n43481 = pi39 & n10164;
  assign n43482 = ~pi38 & ~n43481;
  assign n43483 = ~n43480 & n43482;
  assign po489 = n37451 & ~n43483;
  assign n43485 = pi333 & ~n43421;
  assign n43486 = pi1040 & n43421;
  assign po490 = n43485 | n43486;
  assign n43488 = pi334 & ~n43421;
  assign n43489 = pi1065 & n43421;
  assign po491 = n43488 | n43489;
  assign n43491 = pi335 & ~n43421;
  assign n43492 = pi1069 & n43421;
  assign po492 = n43491 | n43492;
  assign n43494 = pi336 & ~n43417;
  assign n43495 = pi1070 & n43417;
  assign po493 = n43494 | n43495;
  assign n43497 = pi337 & ~n43417;
  assign n43498 = pi1044 & n43417;
  assign po494 = n43497 | n43498;
  assign n43500 = pi338 & ~n43417;
  assign n43501 = pi1072 & n43417;
  assign po495 = n43500 | n43501;
  assign n43503 = pi339 & ~n43417;
  assign n43504 = pi1086 & n43417;
  assign po496 = n43503 | n43504;
  assign n43506 = pi340 & n43459;
  assign n43507 = ~pi340 & ~n43210;
  assign n43508 = n43461 & ~n43507;
  assign n43509 = ~pi331 & n43210;
  assign n43510 = n43508 & ~n43509;
  assign po497 = ~n43506 & ~n43510;
  assign n43512 = ~pi341 & ~po637;
  assign n43513 = ~n43417 & ~n43512;
  assign po498 = n43458 & ~n43513;
  assign n43515 = pi342 & ~n43410;
  assign n43516 = pi1049 & n43410;
  assign po499 = n43515 | n43516;
  assign n43518 = pi343 & ~n43410;
  assign n43519 = pi1062 & n43410;
  assign po500 = n43518 | n43519;
  assign n43521 = pi344 & ~n43410;
  assign n43522 = pi1069 & n43410;
  assign po501 = n43521 | n43522;
  assign n43524 = pi345 & ~n43410;
  assign n43525 = pi1039 & n43410;
  assign po502 = n43524 | n43525;
  assign n43527 = pi346 & ~n43410;
  assign n43528 = pi1067 & n43410;
  assign po503 = n43527 | n43528;
  assign n43530 = pi347 & ~n43410;
  assign n43531 = pi1055 & n43410;
  assign po504 = n43530 | n43531;
  assign n43533 = pi348 & ~n43410;
  assign n43534 = pi1087 & n43410;
  assign po505 = n43533 | n43534;
  assign n43536 = pi349 & ~n43410;
  assign n43537 = pi1043 & n43410;
  assign po506 = n43536 | n43537;
  assign n43539 = pi350 & ~n43410;
  assign n43540 = pi1035 & n43410;
  assign po507 = n43539 | n43540;
  assign n43542 = pi351 & ~n43410;
  assign n43543 = pi1079 & n43410;
  assign po508 = n43542 | n43543;
  assign n43545 = pi352 & ~n43410;
  assign n43546 = pi1078 & n43410;
  assign po509 = n43545 | n43546;
  assign n43548 = pi353 & ~n43410;
  assign n43549 = pi1063 & n43410;
  assign po510 = n43548 | n43549;
  assign n43551 = pi354 & ~n43410;
  assign n43552 = pi1045 & n43410;
  assign po511 = n43551 | n43552;
  assign n43554 = pi355 & ~n43410;
  assign n43555 = pi1084 & n43410;
  assign po512 = n43554 | n43555;
  assign n43557 = pi356 & ~n43410;
  assign n43558 = pi1081 & n43410;
  assign po513 = n43557 | n43558;
  assign n43560 = pi357 & ~n43410;
  assign n43561 = pi1076 & n43410;
  assign po514 = n43560 | n43561;
  assign n43563 = pi358 & ~n43410;
  assign n43564 = pi1071 & n43410;
  assign po515 = n43563 | n43564;
  assign n43566 = pi359 & ~n43410;
  assign n43567 = pi1068 & n43410;
  assign po516 = n43566 | n43567;
  assign n43569 = pi360 & ~n43410;
  assign n43570 = pi1042 & n43410;
  assign po517 = n43569 | n43570;
  assign n43572 = pi361 & ~n43410;
  assign n43573 = pi1059 & n43410;
  assign po518 = n43572 | n43573;
  assign n43575 = pi362 & ~n43410;
  assign n43576 = pi1070 & n43410;
  assign po519 = n43575 | n43576;
  assign n43578 = pi363 & ~n43417;
  assign n43579 = pi1049 & n43417;
  assign po520 = n43578 | n43579;
  assign n43581 = pi364 & ~n43417;
  assign n43582 = pi1062 & n43417;
  assign po521 = n43581 | n43582;
  assign n43584 = pi365 & ~n43417;
  assign n43585 = pi1065 & n43417;
  assign po522 = n43584 | n43585;
  assign n43587 = pi366 & ~n43417;
  assign n43588 = pi1069 & n43417;
  assign po523 = n43587 | n43588;
  assign n43590 = pi367 & ~n43417;
  assign n43591 = pi1039 & n43417;
  assign po524 = n43590 | n43591;
  assign n43593 = pi368 & ~n43417;
  assign n43594 = pi1067 & n43417;
  assign po525 = n43593 | n43594;
  assign n43596 = pi369 & ~n43417;
  assign n43597 = pi1080 & n43417;
  assign po526 = n43596 | n43597;
  assign n43599 = pi370 & ~n43417;
  assign n43600 = pi1055 & n43417;
  assign po527 = n43599 | n43600;
  assign n43602 = pi371 & ~n43417;
  assign n43603 = pi1051 & n43417;
  assign po528 = n43602 | n43603;
  assign n43605 = pi372 & ~n43417;
  assign n43606 = pi1048 & n43417;
  assign po529 = n43605 | n43606;
  assign n43608 = pi373 & ~n43417;
  assign n43609 = pi1087 & n43417;
  assign po530 = n43608 | n43609;
  assign n43611 = pi374 & ~n43417;
  assign n43612 = pi1035 & n43417;
  assign po531 = n43611 | n43612;
  assign n43614 = pi375 & ~n43417;
  assign n43615 = pi1047 & n43417;
  assign po532 = n43614 | n43615;
  assign n43617 = pi376 & ~n43417;
  assign n43618 = pi1079 & n43417;
  assign po533 = n43617 | n43618;
  assign n43620 = pi377 & ~n43417;
  assign n43621 = pi1074 & n43417;
  assign po534 = n43620 | n43621;
  assign n43623 = pi378 & ~n43417;
  assign n43624 = pi1063 & n43417;
  assign po535 = n43623 | n43624;
  assign n43626 = pi379 & ~n43417;
  assign n43627 = pi1045 & n43417;
  assign po536 = n43626 | n43627;
  assign n43629 = pi380 & ~n43417;
  assign n43630 = pi1084 & n43417;
  assign po537 = n43629 | n43630;
  assign n43632 = pi381 & ~n43417;
  assign n43633 = pi1081 & n43417;
  assign po538 = n43632 | n43633;
  assign n43635 = pi382 & ~n43417;
  assign n43636 = pi1076 & n43417;
  assign po539 = n43635 | n43636;
  assign n43638 = pi383 & ~n43417;
  assign n43639 = pi1071 & n43417;
  assign po540 = n43638 | n43639;
  assign n43641 = pi384 & ~n43417;
  assign n43642 = pi1068 & n43417;
  assign po541 = n43641 | n43642;
  assign n43644 = pi385 & ~n43417;
  assign n43645 = pi1042 & n43417;
  assign po542 = n43644 | n43645;
  assign n43647 = pi386 & ~n43417;
  assign n43648 = pi1059 & n43417;
  assign po543 = n43647 | n43648;
  assign n43650 = pi387 & ~n43417;
  assign n43651 = pi1053 & n43417;
  assign po544 = n43650 | n43651;
  assign n43653 = pi388 & ~n43417;
  assign n43654 = pi1037 & n43417;
  assign po545 = n43653 | n43654;
  assign n43656 = pi389 & ~n43417;
  assign n43657 = pi1036 & n43417;
  assign po546 = n43656 | n43657;
  assign n43659 = pi390 & ~n43421;
  assign n43660 = pi1049 & n43421;
  assign po547 = n43659 | n43660;
  assign n43662 = pi391 & ~n43421;
  assign n43663 = pi1062 & n43421;
  assign po548 = n43662 | n43663;
  assign n43665 = pi392 & ~n43421;
  assign n43666 = pi1039 & n43421;
  assign po549 = n43665 | n43666;
  assign n43668 = pi393 & ~n43421;
  assign n43669 = pi1067 & n43421;
  assign po550 = n43668 | n43669;
  assign n43671 = pi394 & ~n43421;
  assign n43672 = pi1080 & n43421;
  assign po551 = n43671 | n43672;
  assign n43674 = pi395 & ~n43421;
  assign n43675 = pi1055 & n43421;
  assign po552 = n43674 | n43675;
  assign n43677 = pi396 & ~n43421;
  assign n43678 = pi1051 & n43421;
  assign po553 = n43677 | n43678;
  assign n43680 = pi397 & ~n43421;
  assign n43681 = pi1048 & n43421;
  assign po554 = n43680 | n43681;
  assign n43683 = pi398 & ~n43421;
  assign n43684 = pi1087 & n43421;
  assign po555 = n43683 | n43684;
  assign n43686 = pi399 & ~n43421;
  assign n43687 = pi1047 & n43421;
  assign po556 = n43686 | n43687;
  assign n43689 = pi400 & ~n43421;
  assign n43690 = pi1035 & n43421;
  assign po557 = n43689 | n43690;
  assign n43692 = pi401 & ~n43421;
  assign n43693 = pi1079 & n43421;
  assign po558 = n43692 | n43693;
  assign n43695 = pi402 & ~n43421;
  assign n43696 = pi1078 & n43421;
  assign po559 = n43695 | n43696;
  assign n43698 = pi403 & ~n43421;
  assign n43699 = pi1045 & n43421;
  assign po560 = n43698 | n43699;
  assign n43701 = pi404 & ~n43421;
  assign n43702 = pi1084 & n43421;
  assign po561 = n43701 | n43702;
  assign n43704 = pi405 & ~n43421;
  assign n43705 = pi1081 & n43421;
  assign po562 = n43704 | n43705;
  assign n43707 = pi406 & ~n43421;
  assign n43708 = pi1076 & n43421;
  assign po563 = n43707 | n43708;
  assign n43710 = pi407 & ~n43421;
  assign n43711 = pi1071 & n43421;
  assign po564 = n43710 | n43711;
  assign n43713 = pi408 & ~n43421;
  assign n43714 = pi1068 & n43421;
  assign po565 = n43713 | n43714;
  assign n43716 = pi409 & ~n43421;
  assign n43717 = pi1042 & n43421;
  assign po566 = n43716 | n43717;
  assign n43719 = pi410 & ~n43421;
  assign n43720 = pi1059 & n43421;
  assign po567 = n43719 | n43720;
  assign n43722 = pi411 & ~n43421;
  assign n43723 = pi1053 & n43421;
  assign po568 = n43722 | n43723;
  assign n43725 = pi412 & ~n43421;
  assign n43726 = pi1037 & n43421;
  assign po569 = n43725 | n43726;
  assign n43728 = pi413 & ~n43421;
  assign n43729 = pi1036 & n43421;
  assign po570 = n43728 | n43729;
  assign n43731 = ~po1038 & n43509;
  assign n43732 = pi414 & ~n43731;
  assign n43733 = pi1049 & n43731;
  assign po571 = n43732 | n43733;
  assign n43735 = pi415 & ~n43731;
  assign n43736 = pi1062 & n43731;
  assign po572 = n43735 | n43736;
  assign n43738 = pi416 & ~n43731;
  assign n43739 = pi1069 & n43731;
  assign po573 = n43738 | n43739;
  assign n43741 = pi417 & ~n43731;
  assign n43742 = pi1039 & n43731;
  assign po574 = n43741 | n43742;
  assign n43744 = pi418 & ~n43731;
  assign n43745 = pi1067 & n43731;
  assign po575 = n43744 | n43745;
  assign n43747 = pi419 & ~n43731;
  assign n43748 = pi1080 & n43731;
  assign po576 = n43747 | n43748;
  assign n43750 = pi420 & ~n43731;
  assign n43751 = pi1055 & n43731;
  assign po577 = n43750 | n43751;
  assign n43753 = pi421 & ~n43731;
  assign n43754 = pi1051 & n43731;
  assign po578 = n43753 | n43754;
  assign n43756 = pi422 & ~n43731;
  assign n43757 = pi1048 & n43731;
  assign po579 = n43756 | n43757;
  assign n43759 = pi423 & ~n43731;
  assign n43760 = pi1087 & n43731;
  assign po580 = n43759 | n43760;
  assign n43762 = pi424 & ~n43731;
  assign n43763 = pi1047 & n43731;
  assign po581 = n43762 | n43763;
  assign n43765 = pi425 & ~n43731;
  assign n43766 = pi1035 & n43731;
  assign po582 = n43765 | n43766;
  assign n43768 = pi426 & ~n43731;
  assign n43769 = pi1079 & n43731;
  assign po583 = n43768 | n43769;
  assign n43771 = pi427 & ~n43731;
  assign n43772 = pi1078 & n43731;
  assign po584 = n43771 | n43772;
  assign n43774 = pi428 & ~n43731;
  assign n43775 = pi1045 & n43731;
  assign po585 = n43774 | n43775;
  assign n43777 = pi429 & ~n43731;
  assign n43778 = pi1084 & n43731;
  assign po586 = n43777 | n43778;
  assign n43780 = pi430 & ~n43731;
  assign n43781 = pi1076 & n43731;
  assign po587 = n43780 | n43781;
  assign n43783 = pi431 & ~n43731;
  assign n43784 = pi1071 & n43731;
  assign po588 = n43783 | n43784;
  assign n43786 = pi432 & ~n43731;
  assign n43787 = pi1068 & n43731;
  assign po589 = n43786 | n43787;
  assign n43789 = pi433 & ~n43731;
  assign n43790 = pi1042 & n43731;
  assign po590 = n43789 | n43790;
  assign n43792 = pi434 & ~n43731;
  assign n43793 = pi1059 & n43731;
  assign po591 = n43792 | n43793;
  assign n43795 = pi435 & ~n43731;
  assign n43796 = pi1053 & n43731;
  assign po592 = n43795 | n43796;
  assign n43798 = pi436 & ~n43731;
  assign n43799 = pi1037 & n43731;
  assign po593 = n43798 | n43799;
  assign n43801 = pi437 & ~n43731;
  assign n43802 = pi1070 & n43731;
  assign po594 = n43801 | n43802;
  assign n43804 = pi438 & ~n43731;
  assign n43805 = pi1036 & n43731;
  assign po595 = n43804 | n43805;
  assign n43807 = pi439 & ~n43417;
  assign n43808 = pi1057 & n43417;
  assign po596 = n43807 | n43808;
  assign n43810 = pi440 & ~n43417;
  assign n43811 = pi1043 & n43417;
  assign po597 = n43810 | n43811;
  assign n43813 = pi441 & ~n43410;
  assign n43814 = pi1044 & n43410;
  assign po598 = n43813 | n43814;
  assign n43816 = pi442 & ~n43417;
  assign n43817 = pi1058 & n43417;
  assign po599 = n43816 | n43817;
  assign n43819 = pi443 & ~n43731;
  assign n43820 = pi1044 & n43731;
  assign po600 = n43819 | n43820;
  assign n43822 = pi444 & ~n43731;
  assign n43823 = pi1072 & n43731;
  assign po601 = n43822 | n43823;
  assign n43825 = pi445 & ~n43731;
  assign n43826 = pi1081 & n43731;
  assign po602 = n43825 | n43826;
  assign n43828 = pi446 & ~n43731;
  assign n43829 = pi1086 & n43731;
  assign po603 = n43828 | n43829;
  assign n43831 = pi447 & ~n43417;
  assign n43832 = pi1040 & n43417;
  assign po604 = n43831 | n43832;
  assign n43834 = pi448 & ~n43731;
  assign n43835 = pi1074 & n43731;
  assign po605 = n43834 | n43835;
  assign n43837 = pi449 & ~n43731;
  assign n43838 = pi1057 & n43731;
  assign po606 = n43837 | n43838;
  assign n43840 = pi450 & ~n43410;
  assign n43841 = pi1036 & n43410;
  assign po607 = n43840 | n43841;
  assign n43843 = pi451 & ~n43731;
  assign n43844 = pi1063 & n43731;
  assign po608 = n43843 | n43844;
  assign n43846 = pi452 & ~n43410;
  assign n43847 = pi1053 & n43410;
  assign po609 = n43846 | n43847;
  assign n43849 = pi453 & ~n43731;
  assign n43850 = pi1040 & n43731;
  assign po610 = n43849 | n43850;
  assign n43852 = pi454 & ~n43731;
  assign n43853 = pi1043 & n43731;
  assign po611 = n43852 | n43853;
  assign n43855 = pi455 & ~n43410;
  assign n43856 = pi1037 & n43410;
  assign po612 = n43855 | n43856;
  assign n43858 = pi456 & ~n43421;
  assign n43859 = pi1044 & n43421;
  assign po613 = n43858 | n43859;
  assign n43861 = ~pi804 & ~pi810;
  assign n43862 = ~pi595 & ~n43861;
  assign n43863 = pi594 & pi600;
  assign n43864 = pi597 & n43863;
  assign n43865 = pi601 & n43864;
  assign n43866 = ~pi599 & pi810;
  assign n43867 = pi596 & ~n43866;
  assign n43868 = pi804 & ~n43867;
  assign n43869 = pi815 & ~n43868;
  assign n43870 = pi595 & ~n43869;
  assign n43871 = n43865 & ~n43870;
  assign n43872 = ~n43862 & n43871;
  assign n43873 = ~pi601 & ~n43861;
  assign n43874 = pi600 & ~pi810;
  assign n43875 = pi804 & ~n43874;
  assign n43876 = ~pi815 & ~n43875;
  assign n43877 = ~n43873 & n43876;
  assign n43878 = ~n43872 & ~n43877;
  assign n43879 = pi605 & ~n43878;
  assign n43880 = pi990 & n43863;
  assign n43881 = ~pi815 & n43875;
  assign n43882 = n43880 & n43881;
  assign n43883 = ~n43879 & ~n43882;
  assign po614 = pi821 & ~n43883;
  assign n43885 = pi458 & ~n43410;
  assign n43886 = pi1072 & n43410;
  assign po615 = n43885 | n43886;
  assign n43888 = pi459 & ~n43731;
  assign n43889 = pi1058 & n43731;
  assign po616 = n43888 | n43889;
  assign n43891 = pi460 & ~n43410;
  assign n43892 = pi1086 & n43410;
  assign po617 = n43891 | n43892;
  assign n43894 = pi461 & ~n43410;
  assign n43895 = pi1057 & n43410;
  assign po618 = n43894 | n43895;
  assign n43897 = pi462 & ~n43410;
  assign n43898 = pi1074 & n43410;
  assign po619 = n43897 | n43898;
  assign n43900 = pi463 & ~n43421;
  assign n43901 = pi1070 & n43421;
  assign po620 = n43900 | n43901;
  assign n43903 = pi464 & ~n43731;
  assign n43904 = pi1065 & n43731;
  assign po621 = n43903 | n43904;
  assign n43906 = ~n11179 & ~n11182;
  assign n43907 = ~pi243 & ~n43906;
  assign n43908 = ~n5793 & ~n5810;
  assign n43909 = pi926 & ~n43908;
  assign n43910 = pi1157 & n43908;
  assign n43911 = ~n43909 & ~n43910;
  assign n43912 = ~n43907 & n43911;
  assign n43913 = ~pi299 & n43323;
  assign n43914 = pi299 & n3531;
  assign n43915 = ~n43913 & ~n43914;
  assign n43916 = ~pi243 & pi1157;
  assign n43917 = ~n43907 & ~n43916;
  assign n43918 = ~n43915 & n43917;
  assign n43919 = ~n11209 & ~n12851;
  assign n43920 = pi926 & ~n43919;
  assign n43921 = n43916 & n43920;
  assign n43922 = ~n43918 & ~n43921;
  assign n43923 = ~n43912 & n43922;
  assign n43924 = ~po1038 & ~n43923;
  assign n43925 = pi1157 & n5747;
  assign n43926 = ~pi243 & n43315;
  assign n43927 = pi926 & n5746;
  assign n43928 = po1038 & ~n43927;
  assign n43929 = ~n43926 & n43928;
  assign n43930 = ~n43925 & n43929;
  assign po622 = ~n43924 & ~n43930;
  assign n43932 = po1038 & ~n43315;
  assign n43933 = ~po1038 & n43906;
  assign n43934 = ~n43932 & ~n43933;
  assign n43935 = ~pi943 & ~n43934;
  assign n43936 = pi943 & n43378;
  assign n43937 = ~n43935 & ~n43936;
  assign n43938 = ~pi1151 & ~n43937;
  assign n43939 = ~n43328 & n43935;
  assign n43940 = ~po1038 & ~n43915;
  assign n43941 = n3531 & po1038;
  assign n43942 = ~n43940 & ~n43941;
  assign n43943 = ~pi275 & ~n43942;
  assign n43944 = ~n43939 & ~n43943;
  assign n43945 = pi943 & ~n43332;
  assign n43946 = pi1151 & n43945;
  assign n43947 = n43944 & ~n43946;
  assign po623 = ~n43938 & n43947;
  assign n43949 = pi40 & ~pi287;
  assign n43950 = n41172 & n43949;
  assign n43951 = po950 & n43950;
  assign n43952 = ~n9986 & ~n43951;
  assign n43953 = ~pi102 & ~n13058;
  assign n43954 = n16127 & ~n43953;
  assign n43955 = n11084 & n16129;
  assign n43956 = n43954 & n43955;
  assign n43957 = n43950 & ~n43956;
  assign n43958 = ~n43950 & n43956;
  assign n43959 = ~n43957 & ~n43958;
  assign n43960 = ~n6122 & ~n43959;
  assign n43961 = n6122 & n43956;
  assign n43962 = ~n43960 & ~n43961;
  assign n43963 = ~n7493 & ~n43962;
  assign n43964 = n7493 & ~n43959;
  assign n43965 = pi1091 & ~n43964;
  assign n43966 = ~n43963 & n43965;
  assign n43967 = ~n7368 & n43959;
  assign n43968 = n7368 & ~n43956;
  assign n43969 = ~n43967 & ~n43968;
  assign n43970 = pi1093 & n43969;
  assign n43971 = ~pi1093 & ~n43962;
  assign n43972 = ~pi1091 & ~n43971;
  assign n43973 = ~n43970 & n43972;
  assign n43974 = ~n43966 & ~n43973;
  assign n43975 = n12806 & ~n43974;
  assign n43976 = n3275 & n43975;
  assign po624 = ~n43952 & ~n43976;
  assign n43978 = n10024 & n11122;
  assign n43979 = n10021 & n18931;
  assign n43980 = n8817 & n43979;
  assign n43981 = pi468 & ~n43980;
  assign po625 = n43978 | n43981;
  assign n43983 = ~pi263 & ~n43906;
  assign n43984 = pi942 & ~n43908;
  assign n43985 = pi1156 & n43908;
  assign n43986 = ~n43984 & ~n43985;
  assign n43987 = ~n43983 & n43986;
  assign n43988 = ~pi263 & pi1156;
  assign n43989 = ~n43983 & ~n43988;
  assign n43990 = ~n43915 & n43989;
  assign n43991 = ~n43919 & n43988;
  assign n43992 = pi942 & n43991;
  assign n43993 = ~n43990 & ~n43992;
  assign n43994 = ~n43987 & n43993;
  assign n43995 = ~po1038 & ~n43994;
  assign n43996 = ~pi263 & n43315;
  assign n43997 = pi942 & n5746;
  assign n43998 = pi1156 & n5747;
  assign n43999 = po1038 & ~n43998;
  assign n44000 = ~n43997 & n43999;
  assign n44001 = ~n43996 & n44000;
  assign po626 = ~n43995 & ~n44001;
  assign n44003 = pi267 & ~n43906;
  assign n44004 = pi925 & ~n43908;
  assign n44005 = pi1155 & n43908;
  assign n44006 = ~n44004 & ~n44005;
  assign n44007 = ~n44003 & n44006;
  assign n44008 = pi267 & pi1155;
  assign n44009 = ~n44003 & ~n44008;
  assign n44010 = ~n43915 & n44009;
  assign n44011 = ~n43919 & n44008;
  assign n44012 = pi925 & n44011;
  assign n44013 = ~n44010 & ~n44012;
  assign n44014 = ~n44007 & n44013;
  assign n44015 = ~po1038 & ~n44014;
  assign n44016 = pi267 & n43315;
  assign n44017 = pi925 & n5746;
  assign n44018 = pi1155 & n5747;
  assign n44019 = po1038 & ~n44018;
  assign n44020 = ~n44017 & n44019;
  assign n44021 = ~n44016 & n44020;
  assign po627 = ~n44015 & ~n44021;
  assign n44023 = pi253 & ~n43906;
  assign n44024 = pi941 & ~n43908;
  assign n44025 = pi1153 & n43908;
  assign n44026 = ~n44024 & ~n44025;
  assign n44027 = ~n44023 & n44026;
  assign n44028 = pi253 & pi1153;
  assign n44029 = ~n44023 & ~n44028;
  assign n44030 = ~n43915 & n44029;
  assign n44031 = ~n43919 & n44028;
  assign n44032 = pi941 & n44031;
  assign n44033 = ~n44030 & ~n44032;
  assign n44034 = ~n44027 & n44033;
  assign n44035 = ~po1038 & ~n44034;
  assign n44036 = pi253 & n43315;
  assign n44037 = pi941 & n5746;
  assign n44038 = pi1153 & n5747;
  assign n44039 = po1038 & ~n44038;
  assign n44040 = ~n44037 & n44039;
  assign n44041 = ~n44036 & n44040;
  assign po628 = ~n44035 & ~n44041;
  assign n44043 = pi254 & ~n43906;
  assign n44044 = pi923 & ~n43908;
  assign n44045 = pi1154 & n43908;
  assign n44046 = ~n44044 & ~n44045;
  assign n44047 = ~n44043 & n44046;
  assign n44048 = pi254 & pi1154;
  assign n44049 = ~n44043 & ~n44048;
  assign n44050 = ~n43915 & n44049;
  assign n44051 = ~n43919 & n44048;
  assign n44052 = pi923 & n44051;
  assign n44053 = ~n44050 & ~n44052;
  assign n44054 = ~n44047 & n44053;
  assign n44055 = ~po1038 & ~n44054;
  assign n44056 = pi254 & n43315;
  assign n44057 = pi923 & n5746;
  assign n44058 = pi1154 & n5747;
  assign n44059 = po1038 & ~n44058;
  assign n44060 = ~n44057 & n44059;
  assign n44061 = ~n44056 & n44060;
  assign po629 = ~n44055 & ~n44061;
  assign n44063 = ~pi922 & ~n43934;
  assign n44064 = pi922 & n43378;
  assign n44065 = ~n44063 & ~n44064;
  assign n44066 = ~pi1152 & ~n44065;
  assign n44067 = ~n43328 & n44063;
  assign n44068 = ~pi268 & ~n43942;
  assign n44069 = ~n44067 & ~n44068;
  assign n44070 = pi922 & ~n43332;
  assign n44071 = pi1152 & n44070;
  assign n44072 = n44069 & ~n44071;
  assign po630 = ~n44066 & n44072;
  assign n44074 = ~pi931 & ~n43934;
  assign n44075 = pi931 & n43378;
  assign n44076 = ~n44074 & ~n44075;
  assign n44077 = ~pi1150 & ~n44076;
  assign n44078 = ~n43328 & n44074;
  assign n44079 = ~pi272 & ~n43942;
  assign n44080 = ~n44078 & ~n44079;
  assign n44081 = pi931 & ~n43332;
  assign n44082 = pi1150 & n44081;
  assign n44083 = n44080 & ~n44082;
  assign po631 = ~n44077 & n44083;
  assign n44085 = ~pi936 & ~n43934;
  assign n44086 = pi936 & n43378;
  assign n44087 = ~n44085 & ~n44086;
  assign n44088 = ~pi1149 & ~n44087;
  assign n44089 = ~n43328 & n44085;
  assign n44090 = ~pi283 & ~n43942;
  assign n44091 = ~n44089 & ~n44090;
  assign n44092 = pi936 & ~n43332;
  assign n44093 = pi1149 & n44092;
  assign n44094 = n44091 & ~n44093;
  assign po632 = ~n44088 & n44094;
  assign n44096 = pi71 & n42303;
  assign n44097 = pi71 & ~n11225;
  assign n44098 = n11225 & n12730;
  assign n44099 = n9975 & ~n11225;
  assign n44100 = n9971 & n44099;
  assign n44101 = ~n44098 & ~n44100;
  assign n44102 = n2576 & ~n44101;
  assign n44103 = n9987 & n44102;
  assign n44104 = n12734 & n44103;
  assign n44105 = ~n44097 & ~n44104;
  assign n44106 = ~po1038 & ~n44105;
  assign po633 = n44096 | n44106;
  assign po635 = pi71 & ~n42607;
  assign n44109 = pi481 & ~n34022;
  assign n44110 = pi248 & n34022;
  assign po638 = n44109 | n44110;
  assign n44112 = pi482 & ~n34038;
  assign n44113 = pi249 & n34038;
  assign po639 = n44112 | n44113;
  assign n44115 = pi483 & ~n34161;
  assign n44116 = pi242 & n34161;
  assign po640 = n44115 | n44116;
  assign n44118 = pi484 & ~n34161;
  assign n44119 = pi249 & n34161;
  assign po641 = n44118 | n44119;
  assign n44121 = pi485 & ~n35332;
  assign n44122 = pi234 & n35332;
  assign po642 = n44121 | n44122;
  assign n44124 = pi486 & ~n35332;
  assign n44125 = pi244 & n35332;
  assign po643 = n44124 | n44125;
  assign n44127 = pi487 & ~n34022;
  assign n44128 = pi246 & n34022;
  assign po644 = n44127 | n44128;
  assign n44130 = pi488 & ~n34022;
  assign n44131 = ~pi239 & n34022;
  assign po645 = ~n44130 & ~n44131;
  assign n44133 = pi489 & ~n35332;
  assign n44134 = pi242 & n35332;
  assign po646 = n44133 | n44134;
  assign n44136 = pi490 & ~n34161;
  assign n44137 = pi241 & n34161;
  assign po647 = n44136 | n44137;
  assign n44139 = pi491 & ~n34161;
  assign n44140 = pi238 & n34161;
  assign po648 = n44139 | n44140;
  assign n44142 = pi492 & ~n34161;
  assign n44143 = pi240 & n34161;
  assign po649 = n44142 | n44143;
  assign n44145 = pi493 & ~n34161;
  assign n44146 = pi244 & n34161;
  assign po650 = n44145 | n44146;
  assign n44148 = pi494 & ~n34161;
  assign n44149 = ~pi239 & n34161;
  assign po651 = ~n44148 & ~n44149;
  assign n44151 = pi495 & ~n34161;
  assign n44152 = pi235 & n34161;
  assign po652 = n44151 | n44152;
  assign n44154 = pi496 & ~n34153;
  assign n44155 = pi249 & n34153;
  assign po653 = n44154 | n44155;
  assign n44157 = pi497 & ~n34153;
  assign n44158 = ~pi239 & n34153;
  assign po654 = ~n44157 & ~n44158;
  assign n44160 = pi498 & ~n34038;
  assign n44161 = pi238 & n34038;
  assign po655 = n44160 | n44161;
  assign n44163 = pi499 & ~n34153;
  assign n44164 = pi246 & n34153;
  assign po656 = n44163 | n44164;
  assign n44166 = pi500 & ~n34153;
  assign n44167 = pi241 & n34153;
  assign po657 = n44166 | n44167;
  assign n44169 = pi501 & ~n34153;
  assign n44170 = pi248 & n34153;
  assign po658 = n44169 | n44170;
  assign n44172 = pi502 & ~n34153;
  assign n44173 = pi247 & n34153;
  assign po659 = n44172 | n44173;
  assign n44175 = pi503 & ~n34153;
  assign n44176 = pi245 & n34153;
  assign po660 = n44175 | n44176;
  assign n44178 = pi504 & ~n34146;
  assign n44179 = pi242 & n34146;
  assign po661 = n44178 | n44179;
  assign n44181 = pi505 & ~n34153;
  assign n44182 = pi234 & n34153;
  assign po662 = n44181 | n44182;
  assign n44184 = pi506 & ~n34146;
  assign n44185 = pi241 & n34146;
  assign po663 = n44184 | n44185;
  assign n44187 = pi507 & ~n34146;
  assign n44188 = pi238 & n34146;
  assign po664 = n44187 | n44188;
  assign n44190 = pi508 & ~n34146;
  assign n44191 = pi247 & n34146;
  assign po665 = n44190 | n44191;
  assign n44193 = pi509 & ~n34146;
  assign n44194 = pi245 & n34146;
  assign po666 = n44193 | n44194;
  assign n44196 = pi510 & ~n34022;
  assign n44197 = pi242 & n34022;
  assign po667 = n44196 | n44197;
  assign n44199 = pi511 & ~n34022;
  assign n44200 = pi234 & n34022;
  assign po668 = n44199 | n44200;
  assign n44202 = pi512 & ~n34022;
  assign n44203 = pi235 & n34022;
  assign po669 = n44202 | n44203;
  assign n44205 = pi513 & ~n34022;
  assign n44206 = pi244 & n34022;
  assign po670 = n44205 | n44206;
  assign n44208 = pi514 & ~n34022;
  assign n44209 = pi245 & n34022;
  assign po671 = n44208 | n44209;
  assign n44211 = pi515 & ~n34022;
  assign n44212 = pi240 & n34022;
  assign po672 = n44211 | n44212;
  assign n44214 = pi516 & ~n34022;
  assign n44215 = pi247 & n34022;
  assign po673 = n44214 | n44215;
  assign n44217 = pi517 & ~n34022;
  assign n44218 = pi238 & n34022;
  assign po674 = n44217 | n44218;
  assign n44220 = pi518 & ~n34030;
  assign n44221 = pi234 & n34030;
  assign po675 = n44220 | n44221;
  assign n44223 = pi519 & ~n34030;
  assign n44224 = ~pi239 & n34030;
  assign po676 = ~n44223 & ~n44224;
  assign n44226 = pi520 & ~n34030;
  assign n44227 = pi246 & n34030;
  assign po677 = n44226 | n44227;
  assign n44229 = pi521 & ~n34030;
  assign n44230 = pi248 & n34030;
  assign po678 = n44229 | n44230;
  assign n44232 = pi522 & ~n34030;
  assign n44233 = pi238 & n34030;
  assign po679 = n44232 | n44233;
  assign n44235 = pi523 & ~n35360;
  assign n44236 = pi234 & n35360;
  assign po680 = n44235 | n44236;
  assign n44238 = pi524 & ~n35360;
  assign n44239 = ~pi239 & n35360;
  assign po681 = ~n44238 & ~n44239;
  assign n44241 = pi525 & ~n35360;
  assign n44242 = pi245 & n35360;
  assign po682 = n44241 | n44242;
  assign n44244 = pi526 & ~n35360;
  assign n44245 = pi246 & n35360;
  assign po683 = n44244 | n44245;
  assign n44247 = pi527 & ~n35360;
  assign n44248 = pi247 & n35360;
  assign po684 = n44247 | n44248;
  assign n44250 = pi528 & ~n35360;
  assign n44251 = pi249 & n35360;
  assign po685 = n44250 | n44251;
  assign n44253 = pi529 & ~n35360;
  assign n44254 = pi238 & n35360;
  assign po686 = n44253 | n44254;
  assign n44256 = pi530 & ~n35360;
  assign n44257 = pi240 & n35360;
  assign po687 = n44256 | n44257;
  assign n44259 = pi531 & ~n34038;
  assign n44260 = pi235 & n34038;
  assign po688 = n44259 | n44260;
  assign n44262 = pi532 & ~n34038;
  assign n44263 = pi247 & n34038;
  assign po689 = n44262 | n44263;
  assign n44265 = pi533 & ~n34146;
  assign n44266 = pi235 & n34146;
  assign po690 = n44265 | n44266;
  assign n44268 = pi534 & ~n34146;
  assign n44269 = ~pi239 & n34146;
  assign po691 = ~n44268 & ~n44269;
  assign n44271 = pi535 & ~n34146;
  assign n44272 = pi240 & n34146;
  assign po692 = n44271 | n44272;
  assign n44274 = pi536 & ~n34146;
  assign n44275 = pi246 & n34146;
  assign po693 = n44274 | n44275;
  assign n44277 = pi537 & ~n34146;
  assign n44278 = pi248 & n34146;
  assign po694 = n44277 | n44278;
  assign n44280 = pi538 & ~n34146;
  assign n44281 = pi249 & n34146;
  assign po695 = n44280 | n44281;
  assign n44283 = pi539 & ~n34153;
  assign n44284 = pi242 & n34153;
  assign po696 = n44283 | n44284;
  assign n44286 = pi540 & ~n34153;
  assign n44287 = pi235 & n34153;
  assign po697 = n44286 | n44287;
  assign n44289 = pi541 & ~n34153;
  assign n44290 = pi244 & n34153;
  assign po698 = n44289 | n44290;
  assign n44292 = pi542 & ~n34153;
  assign n44293 = pi240 & n34153;
  assign po699 = n44292 | n44293;
  assign n44295 = pi543 & ~n34153;
  assign n44296 = pi238 & n34153;
  assign po700 = n44295 | n44296;
  assign n44298 = pi544 & ~n34161;
  assign n44299 = pi234 & n34161;
  assign po701 = n44298 | n44299;
  assign n44301 = pi545 & ~n34161;
  assign n44302 = pi245 & n34161;
  assign po702 = n44301 | n44302;
  assign n44304 = pi546 & ~n34161;
  assign n44305 = pi246 & n34161;
  assign po703 = n44304 | n44305;
  assign n44307 = pi547 & ~n34161;
  assign n44308 = pi247 & n34161;
  assign po704 = n44307 | n44308;
  assign n44310 = pi548 & ~n34161;
  assign n44311 = pi248 & n34161;
  assign po705 = n44310 | n44311;
  assign n44313 = pi549 & ~n35332;
  assign n44314 = pi235 & n35332;
  assign po706 = n44313 | n44314;
  assign n44316 = pi550 & ~n35332;
  assign n44317 = ~pi239 & n35332;
  assign po707 = ~n44316 & ~n44317;
  assign n44319 = pi551 & ~n35332;
  assign n44320 = pi240 & n35332;
  assign po708 = n44319 | n44320;
  assign n44322 = pi552 & ~n35332;
  assign n44323 = pi247 & n35332;
  assign po709 = n44322 | n44323;
  assign n44325 = pi553 & ~n35332;
  assign n44326 = pi241 & n35332;
  assign po710 = n44325 | n44326;
  assign n44328 = pi554 & ~n35332;
  assign n44329 = pi248 & n35332;
  assign po711 = n44328 | n44329;
  assign n44331 = pi555 & ~n35332;
  assign n44332 = pi249 & n35332;
  assign po712 = n44331 | n44332;
  assign n44334 = pi556 & ~n34038;
  assign n44335 = pi242 & n34038;
  assign po713 = n44334 | n44335;
  assign n44337 = pi557 & ~n34146;
  assign n44338 = pi234 & n34146;
  assign po714 = n44337 | n44338;
  assign n44340 = pi558 & ~n34146;
  assign n44341 = pi244 & n34146;
  assign po715 = n44340 | n44341;
  assign n44343 = pi559 & ~n34022;
  assign n44344 = pi241 & n34022;
  assign po716 = n44343 | n44344;
  assign n44346 = pi560 & ~n34038;
  assign n44347 = pi240 & n34038;
  assign po717 = n44346 | n44347;
  assign n44349 = pi561 & ~n34030;
  assign n44350 = pi247 & n34030;
  assign po718 = n44349 | n44350;
  assign n44352 = pi562 & ~n34038;
  assign n44353 = pi241 & n34038;
  assign po719 = n44352 | n44353;
  assign n44355 = pi563 & ~n35332;
  assign n44356 = pi246 & n35332;
  assign po720 = n44355 | n44356;
  assign n44358 = pi564 & ~n34038;
  assign n44359 = pi246 & n34038;
  assign po721 = n44358 | n44359;
  assign n44361 = pi565 & ~n34038;
  assign n44362 = pi248 & n34038;
  assign po722 = n44361 | n44362;
  assign n44364 = pi566 & ~n34038;
  assign n44365 = pi244 & n34038;
  assign po723 = n44364 | n44365;
  assign n44367 = ~pi567 & pi1092;
  assign n44368 = ~pi1093 & n44367;
  assign n44369 = n16124 & ~n44368;
  assign n44370 = pi603 & ~n19656;
  assign n44371 = n16420 & ~n19662;
  assign n44372 = ~n16521 & n44371;
  assign n44373 = n44370 & n44372;
  assign n44374 = ~pi619 & n44373;
  assign n44375 = ~n44368 & ~n44373;
  assign n44376 = ~n44374 & ~n44375;
  assign n44377 = pi1159 & n44376;
  assign n44378 = ~n44368 & ~n44374;
  assign n44379 = ~pi1159 & ~n44378;
  assign n44380 = pi789 & ~n44379;
  assign n44381 = ~n44377 & n44380;
  assign n44382 = ~n44375 & ~n44381;
  assign n44383 = ~n17355 & n44382;
  assign n44384 = n17355 & n44368;
  assign n44385 = ~n44383 & ~n44384;
  assign n44386 = ~n16124 & n44385;
  assign n44387 = ~n44369 & ~n44386;
  assign n44388 = pi647 & n44387;
  assign n44389 = pi680 & ~n18633;
  assign n44390 = n16665 & n44389;
  assign n44391 = ~n44368 & ~n44390;
  assign n44392 = n18716 & ~n44391;
  assign n44393 = ~n44382 & ~n44392;
  assign n44394 = n17356 & ~n44393;
  assign n44395 = n34457 & n44382;
  assign n44396 = ~pi641 & n44392;
  assign n44397 = ~n44368 & ~n44396;
  assign n44398 = n17345 & ~n44397;
  assign n44399 = pi641 & n44392;
  assign n44400 = ~n44368 & ~n44399;
  assign n44401 = n17344 & ~n44400;
  assign n44402 = ~n44398 & ~n44401;
  assign n44403 = ~n44395 & n44402;
  assign n44404 = pi788 & ~n44403;
  assign n44405 = ~n44394 & ~n44404;
  assign n44406 = n19788 & ~n44405;
  assign n44407 = n17448 & ~n44385;
  assign n44408 = n18717 & ~n44391;
  assign n44409 = ~pi628 & n44408;
  assign n44410 = ~n44368 & ~n44409;
  assign n44411 = ~pi1156 & ~n44410;
  assign n44412 = pi629 & ~n44411;
  assign n44413 = ~n44407 & n44412;
  assign n44414 = n17449 & ~n44385;
  assign n44415 = pi628 & n44408;
  assign n44416 = ~n44368 & ~n44415;
  assign n44417 = pi1156 & ~n44416;
  assign n44418 = ~pi629 & ~n44417;
  assign n44419 = ~n44414 & n44418;
  assign n44420 = pi792 & ~n44419;
  assign n44421 = ~n44413 & n44420;
  assign n44422 = ~n44406 & ~n44421;
  assign n44423 = ~pi647 & ~n44422;
  assign n44424 = ~pi1157 & ~n44423;
  assign n44425 = ~n44388 & n44424;
  assign n44426 = ~pi630 & ~n44425;
  assign n44427 = ~n18744 & n44408;
  assign n44428 = pi647 & n44427;
  assign n44429 = ~n44368 & ~n44428;
  assign n44430 = pi1157 & n44429;
  assign n44431 = n44426 & ~n44430;
  assign n44432 = ~pi647 & n44387;
  assign n44433 = pi647 & ~n44422;
  assign n44434 = ~n44432 & ~n44433;
  assign n44435 = pi1157 & n44434;
  assign n44436 = ~pi647 & n44427;
  assign n44437 = ~pi1157 & ~n44368;
  assign n44438 = ~n44436 & n44437;
  assign n44439 = pi630 & ~n44438;
  assign n44440 = ~n44435 & n44439;
  assign n44441 = ~n44431 & ~n44440;
  assign n44442 = pi787 & ~n44441;
  assign n44443 = ~pi787 & ~n44422;
  assign n44444 = ~n44442 & ~n44443;
  assign n44445 = ~pi790 & ~n44444;
  assign n44446 = ~pi644 & ~n44444;
  assign n44447 = ~n18767 & n44427;
  assign n44448 = ~n44368 & ~n44447;
  assign n44449 = pi644 & ~n44448;
  assign n44450 = ~pi715 & ~n44449;
  assign n44451 = ~n44446 & n44450;
  assign n44452 = n23049 & ~n44385;
  assign n44453 = ~pi644 & n44452;
  assign n44454 = ~n44368 & ~n44453;
  assign n44455 = pi715 & n44454;
  assign n44456 = ~n44451 & ~n44455;
  assign n44457 = ~pi1160 & ~n44456;
  assign n44458 = pi644 & n44452;
  assign n44459 = ~n44368 & ~n44458;
  assign n44460 = ~pi715 & ~n44459;
  assign n44461 = pi644 & n44444;
  assign n44462 = ~pi644 & n44448;
  assign n44463 = pi715 & ~n44462;
  assign n44464 = ~n44461 & n44463;
  assign n44465 = pi1160 & ~n44464;
  assign n44466 = ~n44460 & n44465;
  assign n44467 = ~n44457 & ~n44466;
  assign n44468 = pi790 & n44467;
  assign n44469 = ~n44445 & ~n44468;
  assign n44470 = pi230 & ~n44469;
  assign n44471 = ~pi230 & n44367;
  assign po724 = n44470 | n44471;
  assign n44473 = pi568 & ~n34038;
  assign n44474 = pi245 & n34038;
  assign po725 = n44473 | n44474;
  assign n44476 = pi569 & ~n34038;
  assign n44477 = ~pi239 & n34038;
  assign po726 = ~n44476 & ~n44477;
  assign n44479 = pi570 & ~n34038;
  assign n44480 = pi234 & n34038;
  assign po727 = n44479 | n44480;
  assign n44482 = pi571 & ~n35360;
  assign n44483 = pi241 & n35360;
  assign po728 = n44482 | n44483;
  assign n44485 = pi572 & ~n35360;
  assign n44486 = pi244 & n35360;
  assign po729 = n44485 | n44486;
  assign n44488 = pi573 & ~n35360;
  assign n44489 = pi242 & n35360;
  assign po730 = n44488 | n44489;
  assign n44491 = pi574 & ~n34030;
  assign n44492 = pi241 & n34030;
  assign po731 = n44491 | n44492;
  assign n44494 = pi575 & ~n35360;
  assign n44495 = pi235 & n35360;
  assign po732 = n44494 | n44495;
  assign n44497 = pi576 & ~n35360;
  assign n44498 = pi248 & n35360;
  assign po733 = n44497 | n44498;
  assign n44500 = pi577 & ~n35332;
  assign n44501 = pi238 & n35332;
  assign po734 = n44500 | n44501;
  assign n44503 = pi578 & ~n34030;
  assign n44504 = pi249 & n34030;
  assign po735 = n44503 | n44504;
  assign n44506 = pi579 & ~n34022;
  assign n44507 = pi249 & n34022;
  assign po736 = n44506 | n44507;
  assign n44509 = pi580 & ~n35332;
  assign n44510 = pi245 & n35332;
  assign po737 = n44509 | n44510;
  assign n44512 = pi581 & ~n34030;
  assign n44513 = pi235 & n34030;
  assign po738 = n44512 | n44513;
  assign n44515 = pi582 & ~n34030;
  assign n44516 = pi240 & n34030;
  assign po739 = n44515 | n44516;
  assign n44518 = pi584 & ~n34030;
  assign n44519 = pi245 & n34030;
  assign po741 = n44518 | n44519;
  assign n44521 = pi585 & ~n34030;
  assign n44522 = pi244 & n34030;
  assign po742 = n44521 | n44522;
  assign n44524 = pi586 & ~n34030;
  assign n44525 = pi242 & n34030;
  assign po743 = n44524 | n44525;
  assign n44527 = ~pi230 & pi587;
  assign n44528 = pi230 & ~n34837;
  assign n44529 = ~n19662 & n44528;
  assign n44530 = n19668 & n44529;
  assign n44531 = ~n16382 & n44530;
  assign n44532 = n30098 & n44531;
  assign n44533 = n44370 & n44532;
  assign po744 = n44527 | n44533;
  assign n44535 = ~pi123 & n12120;
  assign n44536 = ~pi591 & n44535;
  assign n44537 = ~pi588 & ~n44535;
  assign n44538 = n43458 & ~n44537;
  assign po745 = ~n44536 & n44538;
  assign n44540 = ~pi201 & n34017;
  assign n44541 = ~pi204 & ~n34144;
  assign n44542 = pi233 & ~n44541;
  assign n44543 = ~n44540 & n44542;
  assign n44544 = ~pi202 & n34017;
  assign n44545 = ~pi205 & ~n34144;
  assign n44546 = ~pi233 & ~n44545;
  assign n44547 = ~n44544 & n44546;
  assign n44548 = ~n44543 & ~n44547;
  assign n44549 = pi237 & ~n44548;
  assign n44550 = ~pi220 & n34017;
  assign n44551 = ~pi206 & ~n34144;
  assign n44552 = pi233 & ~n44551;
  assign n44553 = ~n44550 & n44552;
  assign n44554 = ~pi203 & n34017;
  assign n44555 = ~pi218 & ~n34144;
  assign n44556 = ~pi233 & ~n44555;
  assign n44557 = ~n44554 & n44556;
  assign n44558 = ~n44553 & ~n44557;
  assign n44559 = ~pi237 & ~n44558;
  assign po746 = ~n44549 & ~n44559;
  assign n44561 = pi590 & ~n44535;
  assign n44562 = pi588 & n44535;
  assign n44563 = n43458 & ~n44562;
  assign po747 = n44561 | ~n44563;
  assign n44565 = ~pi592 & n44535;
  assign n44566 = ~pi591 & ~n44535;
  assign n44567 = n43458 & ~n44566;
  assign po748 = ~n44565 & n44567;
  assign n44569 = ~pi590 & n44535;
  assign n44570 = ~pi592 & ~n44535;
  assign n44571 = n43458 & ~n44570;
  assign po749 = ~n44569 & n44571;
  assign n44573 = pi246 & pi536;
  assign n44574 = ~pi246 & ~pi536;
  assign n44575 = ~n44573 & ~n44574;
  assign n44576 = pi240 & pi535;
  assign n44577 = ~pi240 & ~pi535;
  assign n44578 = ~n44576 & ~n44577;
  assign n44579 = pi241 & pi506;
  assign n44580 = ~pi241 & ~pi506;
  assign n44581 = ~n44579 & ~n44580;
  assign n44582 = ~pi248 & ~pi537;
  assign n44583 = pi248 & pi537;
  assign n44584 = ~n44582 & ~n44583;
  assign n44585 = ~pi249 & ~pi538;
  assign n44586 = pi249 & pi538;
  assign n44587 = ~n44585 & ~n44586;
  assign n44588 = ~pi234 & ~n34144;
  assign n44589 = ~pi557 & ~n44588;
  assign n44590 = pi234 & ~n34144;
  assign n44591 = pi557 & ~n44590;
  assign n44592 = ~n44589 & ~n44591;
  assign n44593 = ~n44587 & n44592;
  assign n44594 = ~n44584 & n44593;
  assign n44595 = ~n44581 & n44594;
  assign n44596 = ~n44578 & n44595;
  assign n44597 = ~n44575 & n44596;
  assign n44598 = pi239 & ~pi534;
  assign n44599 = ~pi239 & pi534;
  assign n44600 = ~n44598 & ~n44599;
  assign n44601 = n44597 & ~n44600;
  assign n44602 = ~pi242 & ~pi504;
  assign n44603 = pi242 & pi504;
  assign n44604 = ~n44602 & ~n44603;
  assign n44605 = n44601 & ~n44604;
  assign n44606 = ~pi235 & ~pi533;
  assign n44607 = pi235 & pi533;
  assign n44608 = ~n44606 & ~n44607;
  assign n44609 = n44605 & ~n44608;
  assign n44610 = ~pi244 & ~pi558;
  assign n44611 = pi244 & pi558;
  assign n44612 = ~n44610 & ~n44611;
  assign n44613 = n44609 & ~n44612;
  assign n44614 = ~pi245 & ~pi509;
  assign n44615 = pi245 & pi509;
  assign n44616 = ~n44614 & ~n44615;
  assign n44617 = n44613 & ~n44616;
  assign n44618 = ~pi247 & ~pi508;
  assign n44619 = pi247 & pi508;
  assign n44620 = ~n44618 & ~n44619;
  assign n44621 = n44617 & ~n44620;
  assign n44622 = ~pi238 & n44621;
  assign n44623 = ~pi240 & ~pi515;
  assign n44624 = pi240 & pi515;
  assign n44625 = ~n44623 & ~n44624;
  assign n44626 = pi247 & pi516;
  assign n44627 = ~pi247 & ~pi516;
  assign n44628 = ~n44626 & ~n44627;
  assign n44629 = pi245 & pi514;
  assign n44630 = ~pi245 & ~pi514;
  assign n44631 = ~n44629 & ~n44630;
  assign n44632 = pi244 & pi513;
  assign n44633 = ~pi244 & ~pi513;
  assign n44634 = ~n44632 & ~n44633;
  assign n44635 = pi235 & pi512;
  assign n44636 = ~pi235 & ~pi512;
  assign n44637 = ~n44635 & ~n44636;
  assign n44638 = pi242 & pi510;
  assign n44639 = ~pi242 & ~pi510;
  assign n44640 = ~n44638 & ~n44639;
  assign n44641 = ~pi239 & pi488;
  assign n44642 = pi239 & ~pi488;
  assign n44643 = ~n44641 & ~n44642;
  assign n44644 = pi246 & pi487;
  assign n44645 = ~pi246 & ~pi487;
  assign n44646 = ~n44644 & ~n44645;
  assign n44647 = ~pi234 & n34017;
  assign n44648 = ~pi511 & ~n44647;
  assign n44649 = pi248 & pi481;
  assign n44650 = ~pi248 & ~pi481;
  assign n44651 = ~n44649 & ~n44650;
  assign n44652 = ~pi249 & ~pi579;
  assign n44653 = pi249 & pi579;
  assign n44654 = ~n44652 & ~n44653;
  assign n44655 = pi234 & n34017;
  assign n44656 = pi511 & ~n44655;
  assign n44657 = ~n44654 & ~n44656;
  assign n44658 = ~n44651 & n44657;
  assign n44659 = ~n44648 & n44658;
  assign n44660 = ~n44646 & n44659;
  assign n44661 = ~pi241 & ~pi559;
  assign n44662 = pi241 & pi559;
  assign n44663 = ~n44661 & ~n44662;
  assign n44664 = n44660 & ~n44663;
  assign n44665 = ~n44643 & n44664;
  assign n44666 = ~n44640 & n44665;
  assign n44667 = ~n44637 & n44666;
  assign n44668 = ~n44634 & n44667;
  assign n44669 = ~n44631 & n44668;
  assign n44670 = ~n44628 & n44669;
  assign n44671 = ~n44625 & n44670;
  assign n44672 = ~pi238 & n44671;
  assign n44673 = ~pi517 & ~n44672;
  assign n44674 = ~n44622 & n44673;
  assign n44675 = ~pi507 & ~n44674;
  assign n44676 = pi238 & n44671;
  assign n44677 = ~n44622 & ~n44676;
  assign n44678 = pi517 & n44677;
  assign n44679 = n44675 & ~n44678;
  assign n44680 = pi238 & n44621;
  assign n44681 = ~n44676 & ~n44680;
  assign n44682 = pi517 & n44681;
  assign n44683 = n44673 & ~n44680;
  assign n44684 = pi507 & ~n44683;
  assign n44685 = ~n44682 & n44684;
  assign n44686 = ~n44679 & ~n44685;
  assign n44687 = pi233 & ~n44686;
  assign n44688 = ~pi248 & ~pi501;
  assign n44689 = pi248 & pi501;
  assign n44690 = ~n44688 & ~n44689;
  assign n44691 = pi245 & pi503;
  assign n44692 = ~pi245 & ~pi503;
  assign n44693 = ~n44691 & ~n44692;
  assign n44694 = pi244 & pi541;
  assign n44695 = ~pi244 & ~pi541;
  assign n44696 = ~n44694 & ~n44695;
  assign n44697 = ~pi235 & ~pi540;
  assign n44698 = pi235 & pi540;
  assign n44699 = ~n44697 & ~n44698;
  assign n44700 = ~pi242 & ~pi539;
  assign n44701 = pi242 & pi539;
  assign n44702 = ~n44700 & ~n44701;
  assign n44703 = pi239 & ~pi497;
  assign n44704 = ~pi239 & pi497;
  assign n44705 = ~n44703 & ~n44704;
  assign n44706 = ~pi249 & ~pi496;
  assign n44707 = pi249 & pi496;
  assign n44708 = ~n44706 & ~n44707;
  assign n44709 = pi240 & pi542;
  assign n44710 = ~pi240 & ~pi542;
  assign n44711 = ~n44709 & ~n44710;
  assign n44712 = ~pi241 & ~pi500;
  assign n44713 = pi241 & pi500;
  assign n44714 = ~n44712 & ~n44713;
  assign n44715 = ~pi505 & ~n44588;
  assign n44716 = pi505 & ~n44590;
  assign n44717 = ~pi246 & ~pi499;
  assign n44718 = pi246 & pi499;
  assign n44719 = ~n44717 & ~n44718;
  assign n44720 = ~n44716 & ~n44719;
  assign n44721 = ~n44715 & n44720;
  assign n44722 = ~n44714 & n44721;
  assign n44723 = ~n44711 & n44722;
  assign n44724 = ~n44708 & n44723;
  assign n44725 = ~n44705 & n44724;
  assign n44726 = ~n44702 & n44725;
  assign n44727 = ~n44699 & n44726;
  assign n44728 = ~n44696 & n44727;
  assign n44729 = ~n44693 & n44728;
  assign n44730 = ~n44690 & n44729;
  assign n44731 = ~pi247 & ~pi502;
  assign n44732 = pi247 & pi502;
  assign n44733 = ~n44731 & ~n44732;
  assign n44734 = n44730 & ~n44733;
  assign n44735 = ~pi238 & n44734;
  assign n44736 = ~pi245 & ~pi584;
  assign n44737 = pi245 & pi584;
  assign n44738 = ~n44736 & ~n44737;
  assign n44739 = ~pi247 & ~pi561;
  assign n44740 = pi247 & pi561;
  assign n44741 = ~n44739 & ~n44740;
  assign n44742 = ~pi249 & pi578;
  assign n44743 = ~pi240 & ~pi582;
  assign n44744 = pi240 & pi582;
  assign n44745 = ~n44743 & ~n44744;
  assign n44746 = pi235 & pi581;
  assign n44747 = ~pi235 & ~pi581;
  assign n44748 = ~n44746 & ~n44747;
  assign n44749 = pi242 & pi586;
  assign n44750 = ~pi242 & ~pi586;
  assign n44751 = ~n44749 & ~n44750;
  assign n44752 = ~pi239 & pi519;
  assign n44753 = pi239 & ~pi519;
  assign n44754 = ~n44752 & ~n44753;
  assign n44755 = ~pi246 & ~pi520;
  assign n44756 = pi246 & pi520;
  assign n44757 = ~n44755 & ~n44756;
  assign n44758 = ~pi518 & ~n44647;
  assign n44759 = pi518 & ~n44655;
  assign n44760 = pi241 & pi574;
  assign n44761 = ~pi241 & ~pi574;
  assign n44762 = ~n44760 & ~n44761;
  assign n44763 = pi249 & ~pi578;
  assign n44764 = ~pi248 & ~pi521;
  assign n44765 = pi248 & pi521;
  assign n44766 = ~n44764 & ~n44765;
  assign n44767 = ~n44763 & ~n44766;
  assign n44768 = ~n44762 & n44767;
  assign n44769 = ~n44759 & n44768;
  assign n44770 = ~n44758 & n44769;
  assign n44771 = ~n44757 & n44770;
  assign n44772 = ~n44754 & n44771;
  assign n44773 = ~n44751 & n44772;
  assign n44774 = ~n44748 & n44773;
  assign n44775 = ~n44745 & n44774;
  assign n44776 = ~n44742 & n44775;
  assign n44777 = ~pi244 & ~pi585;
  assign n44778 = pi244 & pi585;
  assign n44779 = ~n44777 & ~n44778;
  assign n44780 = n44776 & ~n44779;
  assign n44781 = ~n44741 & n44780;
  assign n44782 = ~n44738 & n44781;
  assign n44783 = ~pi238 & n44782;
  assign n44784 = ~pi522 & ~n44783;
  assign n44785 = ~n44735 & n44784;
  assign n44786 = ~pi543 & ~n44785;
  assign n44787 = pi238 & n44782;
  assign n44788 = ~n44735 & ~n44787;
  assign n44789 = pi522 & n44788;
  assign n44790 = n44786 & ~n44789;
  assign n44791 = pi238 & n44734;
  assign n44792 = ~n44787 & ~n44791;
  assign n44793 = pi522 & n44792;
  assign n44794 = n44784 & ~n44791;
  assign n44795 = pi543 & ~n44794;
  assign n44796 = ~n44793 & n44795;
  assign n44797 = ~n44790 & ~n44796;
  assign n44798 = ~pi233 & ~n44797;
  assign n44799 = pi237 & ~n44798;
  assign n44800 = ~n44687 & n44799;
  assign n44801 = ~pi235 & ~pi495;
  assign n44802 = pi235 & pi495;
  assign n44803 = ~n44801 & ~n44802;
  assign n44804 = pi244 & pi493;
  assign n44805 = ~pi244 & ~pi493;
  assign n44806 = ~n44804 & ~n44805;
  assign n44807 = pi248 & pi548;
  assign n44808 = ~pi248 & ~pi548;
  assign n44809 = ~n44807 & ~n44808;
  assign n44810 = pi249 & pi484;
  assign n44811 = ~pi249 & ~pi484;
  assign n44812 = ~n44810 & ~n44811;
  assign n44813 = ~pi240 & ~pi492;
  assign n44814 = pi240 & pi492;
  assign n44815 = ~n44813 & ~n44814;
  assign n44816 = pi241 & pi490;
  assign n44817 = ~pi241 & ~pi490;
  assign n44818 = ~n44816 & ~n44817;
  assign n44819 = pi544 & ~n44590;
  assign n44820 = ~pi544 & ~n44588;
  assign n44821 = pi246 & pi546;
  assign n44822 = ~pi246 & ~pi546;
  assign n44823 = ~n44821 & ~n44822;
  assign n44824 = ~n44820 & ~n44823;
  assign n44825 = ~n44819 & n44824;
  assign n44826 = ~n44818 & n44825;
  assign n44827 = ~n44815 & n44826;
  assign n44828 = ~n44812 & n44827;
  assign n44829 = ~n44809 & n44828;
  assign n44830 = pi239 & ~pi494;
  assign n44831 = ~pi239 & pi494;
  assign n44832 = ~n44830 & ~n44831;
  assign n44833 = n44829 & ~n44832;
  assign n44834 = ~pi242 & ~pi483;
  assign n44835 = pi242 & pi483;
  assign n44836 = ~n44834 & ~n44835;
  assign n44837 = n44833 & ~n44836;
  assign n44838 = ~n44806 & n44837;
  assign n44839 = ~n44803 & n44838;
  assign n44840 = ~pi245 & ~pi545;
  assign n44841 = pi245 & pi545;
  assign n44842 = ~n44840 & ~n44841;
  assign n44843 = n44839 & ~n44842;
  assign n44844 = ~pi247 & ~pi547;
  assign n44845 = pi247 & pi547;
  assign n44846 = ~n44844 & ~n44845;
  assign n44847 = n44843 & ~n44846;
  assign n44848 = ~pi238 & n44847;
  assign n44849 = ~pi244 & ~pi572;
  assign n44850 = pi244 & pi572;
  assign n44851 = ~n44849 & ~n44850;
  assign n44852 = pi247 & pi527;
  assign n44853 = ~pi247 & ~pi527;
  assign n44854 = ~n44852 & ~n44853;
  assign n44855 = pi245 & pi525;
  assign n44856 = ~pi245 & ~pi525;
  assign n44857 = ~n44855 & ~n44856;
  assign n44858 = pi248 & pi576;
  assign n44859 = ~pi248 & ~pi576;
  assign n44860 = ~n44858 & ~n44859;
  assign n44861 = pi235 & pi575;
  assign n44862 = ~pi235 & ~pi575;
  assign n44863 = ~n44861 & ~n44862;
  assign n44864 = pi242 & pi573;
  assign n44865 = ~pi242 & ~pi573;
  assign n44866 = ~n44864 & ~n44865;
  assign n44867 = ~pi239 & pi524;
  assign n44868 = pi239 & ~pi524;
  assign n44869 = ~n44867 & ~n44868;
  assign n44870 = ~pi240 & ~pi530;
  assign n44871 = pi240 & pi530;
  assign n44872 = ~n44870 & ~n44871;
  assign n44873 = ~pi241 & ~pi571;
  assign n44874 = pi241 & pi571;
  assign n44875 = ~n44873 & ~n44874;
  assign n44876 = pi249 & pi528;
  assign n44877 = ~pi249 & ~pi528;
  assign n44878 = ~n44876 & ~n44877;
  assign n44879 = ~pi523 & ~n44647;
  assign n44880 = pi523 & ~n44655;
  assign n44881 = pi246 & pi526;
  assign n44882 = ~pi246 & ~pi526;
  assign n44883 = ~n44881 & ~n44882;
  assign n44884 = ~n44880 & ~n44883;
  assign n44885 = ~n44879 & n44884;
  assign n44886 = ~n44878 & n44885;
  assign n44887 = ~n44875 & n44886;
  assign n44888 = ~n44872 & n44887;
  assign n44889 = ~n44869 & n44888;
  assign n44890 = ~n44866 & n44889;
  assign n44891 = ~n44863 & n44890;
  assign n44892 = ~n44860 & n44891;
  assign n44893 = ~n44857 & n44892;
  assign n44894 = ~n44854 & n44893;
  assign n44895 = ~n44851 & n44894;
  assign n44896 = ~pi238 & n44895;
  assign n44897 = ~pi529 & ~n44896;
  assign n44898 = ~n44848 & n44897;
  assign n44899 = ~pi491 & ~n44898;
  assign n44900 = pi238 & n44895;
  assign n44901 = ~n44848 & ~n44900;
  assign n44902 = pi529 & n44901;
  assign n44903 = n44899 & ~n44902;
  assign n44904 = pi238 & n44847;
  assign n44905 = ~n44900 & ~n44904;
  assign n44906 = pi529 & n44905;
  assign n44907 = n44897 & ~n44904;
  assign n44908 = pi491 & ~n44907;
  assign n44909 = ~n44906 & n44908;
  assign n44910 = ~n44903 & ~n44909;
  assign n44911 = pi233 & ~n44910;
  assign n44912 = ~pi245 & ~pi568;
  assign n44913 = pi245 & pi568;
  assign n44914 = ~n44912 & ~n44913;
  assign n44915 = pi247 & pi532;
  assign n44916 = ~pi247 & ~pi532;
  assign n44917 = ~n44915 & ~n44916;
  assign n44918 = ~pi248 & ~pi565;
  assign n44919 = pi248 & pi565;
  assign n44920 = ~n44918 & ~n44919;
  assign n44921 = pi244 & pi566;
  assign n44922 = ~pi244 & ~pi566;
  assign n44923 = ~n44921 & ~n44922;
  assign n44924 = pi235 & pi531;
  assign n44925 = ~pi235 & ~pi531;
  assign n44926 = ~n44924 & ~n44925;
  assign n44927 = ~pi242 & ~pi556;
  assign n44928 = pi242 & pi556;
  assign n44929 = ~n44927 & ~n44928;
  assign n44930 = ~pi239 & pi569;
  assign n44931 = pi239 & ~pi569;
  assign n44932 = ~n44930 & ~n44931;
  assign n44933 = ~pi246 & pi564;
  assign n44934 = ~pi249 & ~pi482;
  assign n44935 = pi249 & pi482;
  assign n44936 = ~n44934 & ~n44935;
  assign n44937 = ~pi570 & ~n44647;
  assign n44938 = pi570 & ~n44655;
  assign n44939 = pi241 & pi562;
  assign n44940 = ~pi241 & ~pi562;
  assign n44941 = ~n44939 & ~n44940;
  assign n44942 = ~n44938 & ~n44941;
  assign n44943 = ~n44937 & n44942;
  assign n44944 = ~n44936 & n44943;
  assign n44945 = ~n44933 & n44944;
  assign n44946 = pi240 & pi560;
  assign n44947 = ~pi240 & ~pi560;
  assign n44948 = ~n44946 & ~n44947;
  assign n44949 = pi246 & ~pi564;
  assign n44950 = ~n44948 & ~n44949;
  assign n44951 = n44945 & n44950;
  assign n44952 = ~n44932 & n44951;
  assign n44953 = ~n44929 & n44952;
  assign n44954 = ~n44926 & n44953;
  assign n44955 = ~n44923 & n44954;
  assign n44956 = ~n44920 & n44955;
  assign n44957 = ~n44917 & n44956;
  assign n44958 = ~n44914 & n44957;
  assign n44959 = ~pi238 & n44958;
  assign n44960 = pi577 & ~n44959;
  assign n44961 = ~pi244 & ~pi486;
  assign n44962 = pi244 & pi486;
  assign n44963 = ~n44961 & ~n44962;
  assign n44964 = pi245 & pi580;
  assign n44965 = ~pi245 & ~pi580;
  assign n44966 = ~n44964 & ~n44965;
  assign n44967 = ~pi249 & ~pi555;
  assign n44968 = pi249 & pi555;
  assign n44969 = ~n44967 & ~n44968;
  assign n44970 = ~pi235 & ~pi549;
  assign n44971 = pi235 & pi549;
  assign n44972 = ~n44970 & ~n44971;
  assign n44973 = ~pi242 & ~pi489;
  assign n44974 = pi242 & pi489;
  assign n44975 = ~n44973 & ~n44974;
  assign n44976 = pi239 & ~pi550;
  assign n44977 = ~pi239 & pi550;
  assign n44978 = ~n44976 & ~n44977;
  assign n44979 = ~pi241 & ~pi553;
  assign n44980 = pi241 & pi553;
  assign n44981 = ~n44979 & ~n44980;
  assign n44982 = ~pi485 & ~n44588;
  assign n44983 = pi485 & ~n44590;
  assign n44984 = pi240 & pi551;
  assign n44985 = ~pi240 & ~pi551;
  assign n44986 = ~n44984 & ~n44985;
  assign n44987 = ~pi248 & pi554;
  assign n44988 = pi248 & ~pi554;
  assign n44989 = ~pi246 & ~pi563;
  assign n44990 = pi246 & pi563;
  assign n44991 = ~n44989 & ~n44990;
  assign n44992 = ~n44988 & ~n44991;
  assign n44993 = ~n44987 & n44992;
  assign n44994 = ~n44986 & n44993;
  assign n44995 = ~n44983 & n44994;
  assign n44996 = ~n44982 & n44995;
  assign n44997 = ~n44981 & n44996;
  assign n44998 = ~n44978 & n44997;
  assign n44999 = ~n44975 & n44998;
  assign n45000 = ~n44972 & n44999;
  assign n45001 = ~n44969 & n45000;
  assign n45002 = ~n44966 & n45001;
  assign n45003 = ~n44963 & n45002;
  assign n45004 = ~pi247 & ~pi552;
  assign n45005 = pi247 & pi552;
  assign n45006 = ~n45004 & ~n45005;
  assign n45007 = n45003 & ~n45006;
  assign n45008 = pi238 & n45007;
  assign n45009 = n44960 & ~n45008;
  assign n45010 = ~pi498 & ~n45009;
  assign n45011 = ~pi238 & n45007;
  assign n45012 = ~pi577 & ~n45011;
  assign n45013 = ~n44959 & n45012;
  assign n45014 = n45010 & ~n45013;
  assign n45015 = pi238 & n44958;
  assign n45016 = ~n45008 & ~n45015;
  assign n45017 = pi577 & n45016;
  assign n45018 = n45012 & ~n45015;
  assign n45019 = pi498 & ~n45018;
  assign n45020 = ~n45017 & n45019;
  assign n45021 = ~n45014 & ~n45020;
  assign n45022 = ~pi233 & ~n45021;
  assign n45023 = ~pi237 & ~n45022;
  assign n45024 = ~n44911 & n45023;
  assign po750 = ~n44800 & ~n45024;
  assign n45026 = ~pi806 & n43880;
  assign n45027 = ~pi332 & ~pi806;
  assign n45028 = pi990 & n45027;
  assign n45029 = pi600 & n45028;
  assign n45030 = ~pi332 & pi594;
  assign n45031 = ~n45029 & ~n45030;
  assign po751 = ~n45026 & ~n45031;
  assign n45033 = pi605 & ~pi806;
  assign n45034 = n43865 & n45033;
  assign n45035 = pi595 & n45034;
  assign n45036 = ~pi595 & ~n45034;
  assign n45037 = ~n45035 & ~n45036;
  assign po752 = ~pi332 & n45037;
  assign n45039 = ~pi332 & pi596;
  assign n45040 = pi595 & n43864;
  assign n45041 = n45028 & n45040;
  assign n45042 = ~n45039 & ~n45041;
  assign n45043 = pi596 & n45041;
  assign po753 = ~n45042 & ~n45043;
  assign n45045 = pi597 & n45026;
  assign n45046 = ~pi597 & ~n45026;
  assign n45047 = ~n45045 & ~n45046;
  assign po754 = ~pi332 & n45047;
  assign n45049 = ~pi882 & ~po1038;
  assign n45050 = pi947 & n45049;
  assign n45051 = pi598 & ~n45050;
  assign n45052 = pi740 & pi780;
  assign n45053 = n6185 & n45052;
  assign po755 = n45051 | n45053;
  assign n45055 = ~pi332 & pi599;
  assign n45056 = ~n45043 & ~n45055;
  assign n45057 = pi599 & n45043;
  assign po756 = ~n45056 & ~n45057;
  assign n45059 = ~pi332 & pi600;
  assign n45060 = ~n45028 & ~n45059;
  assign po757 = ~n45029 & ~n45060;
  assign n45062 = ~pi601 & pi806;
  assign n45063 = ~pi806 & ~pi989;
  assign n45064 = ~pi332 & ~n45063;
  assign po758 = ~n45062 & n45064;
  assign n45066 = ~pi230 & pi602;
  assign n45067 = ~n18633 & n18717;
  assign n45068 = pi715 & pi1160;
  assign n45069 = ~pi715 & ~pi1160;
  assign n45070 = pi790 & ~n45069;
  assign n45071 = ~n45068 & n45070;
  assign n45072 = pi230 & ~n45071;
  assign n45073 = ~n17451 & n45072;
  assign n45074 = n45067 & n45073;
  assign n45075 = ~n18767 & n45074;
  assign n45076 = n16596 & n45075;
  assign po759 = n45066 | n45076;
  assign n45078 = pi832 & ~pi1061;
  assign n45079 = ~pi980 & pi1038;
  assign n45080 = pi1060 & n45079;
  assign n45081 = pi952 & n45080;
  assign po897 = n45078 & n45081;
  assign n45083 = ~pi1100 & po897;
  assign n45084 = ~pi603 & ~po897;
  assign n45085 = ~pi966 & ~n45084;
  assign n45086 = ~n45083 & n45085;
  assign n45087 = pi872 & pi966;
  assign n45088 = pi871 & pi966;
  assign n45089 = ~n45087 & ~n45088;
  assign po760 = n45086 | ~n45089;
  assign n45091 = pi823 & n6187;
  assign n45092 = ~pi779 & n45091;
  assign n45093 = ~pi299 & pi983;
  assign n45094 = pi907 & n45093;
  assign n45095 = ~n45091 & ~n45094;
  assign n45096 = pi604 & n45095;
  assign po761 = n45092 | n45096;
  assign n45098 = ~pi605 & ~n45027;
  assign n45099 = ~pi332 & ~n45033;
  assign po762 = ~n45098 & n45099;
  assign n45101 = ~pi606 & ~po897;
  assign n45102 = ~pi1104 & po897;
  assign n45103 = ~n45101 & ~n45102;
  assign n45104 = ~pi966 & ~n45103;
  assign n45105 = ~pi837 & pi966;
  assign po763 = ~n45104 & ~n45105;
  assign n45107 = ~pi1107 & po897;
  assign n45108 = ~pi607 & ~po897;
  assign n45109 = ~pi966 & ~n45108;
  assign po764 = ~n45107 & n45109;
  assign n45111 = ~pi1116 & po897;
  assign n45112 = ~pi608 & ~po897;
  assign n45113 = ~pi966 & ~n45112;
  assign po765 = ~n45111 & n45113;
  assign n45115 = ~pi1118 & po897;
  assign n45116 = ~pi609 & ~po897;
  assign n45117 = ~pi966 & ~n45116;
  assign po766 = ~n45115 & n45117;
  assign n45119 = ~pi1113 & po897;
  assign n45120 = ~pi610 & ~po897;
  assign n45121 = ~pi966 & ~n45120;
  assign po767 = ~n45119 & n45121;
  assign n45123 = ~pi1114 & po897;
  assign n45124 = ~pi611 & ~po897;
  assign n45125 = ~pi966 & ~n45124;
  assign po768 = ~n45123 & n45125;
  assign n45127 = ~pi1111 & po897;
  assign n45128 = ~pi612 & ~po897;
  assign n45129 = ~pi966 & ~n45128;
  assign po769 = ~n45127 & n45129;
  assign n45131 = ~pi1115 & po897;
  assign n45132 = ~pi613 & ~po897;
  assign n45133 = ~pi966 & ~n45132;
  assign po770 = ~n45131 & n45133;
  assign n45135 = ~pi1102 & po897;
  assign n45136 = ~pi614 & ~po897;
  assign n45137 = ~pi966 & ~n45136;
  assign n45138 = ~n45135 & n45137;
  assign po771 = n45088 | n45138;
  assign n45140 = pi907 & n45049;
  assign n45141 = ~pi615 & ~n45140;
  assign n45142 = pi779 & pi797;
  assign n45143 = n6188 & n45142;
  assign po772 = n45141 | n45143;
  assign n45145 = ~pi1101 & po897;
  assign n45146 = ~pi616 & ~po897;
  assign n45147 = ~pi966 & ~n45146;
  assign n45148 = ~n45145 & n45147;
  assign po773 = n45087 | n45148;
  assign n45150 = ~pi617 & ~po897;
  assign n45151 = ~pi1105 & po897;
  assign n45152 = ~n45150 & ~n45151;
  assign n45153 = ~pi966 & ~n45152;
  assign n45154 = ~pi850 & pi966;
  assign po774 = ~n45153 & ~n45154;
  assign n45156 = ~pi1117 & po897;
  assign n45157 = ~pi618 & ~po897;
  assign n45158 = ~pi966 & ~n45157;
  assign po775 = ~n45156 & n45158;
  assign n45160 = ~pi1122 & po897;
  assign n45161 = ~pi619 & ~po897;
  assign n45162 = ~pi966 & ~n45161;
  assign po776 = ~n45160 & n45162;
  assign n45164 = ~pi1112 & po897;
  assign n45165 = ~pi620 & ~po897;
  assign n45166 = ~pi966 & ~n45165;
  assign po777 = ~n45164 & n45166;
  assign n45168 = ~pi1108 & po897;
  assign n45169 = ~pi621 & ~po897;
  assign n45170 = ~pi966 & ~n45169;
  assign po778 = ~n45168 & n45170;
  assign n45172 = ~pi1109 & po897;
  assign n45173 = ~pi622 & ~po897;
  assign n45174 = ~pi966 & ~n45173;
  assign po779 = ~n45172 & n45174;
  assign n45176 = ~pi1106 & po897;
  assign n45177 = ~pi623 & ~po897;
  assign n45178 = ~pi966 & ~n45177;
  assign po780 = ~n45176 & n45178;
  assign n45180 = pi831 & n16392;
  assign n45181 = ~pi780 & n45180;
  assign n45182 = pi947 & n45093;
  assign n45183 = ~n45180 & ~n45182;
  assign n45184 = pi624 & n45183;
  assign po781 = n45181 | n45184;
  assign n45186 = pi832 & ~pi973;
  assign n45187 = ~pi1054 & pi1066;
  assign n45188 = pi1088 & n45187;
  assign n45189 = n45186 & n45188;
  assign po954 = ~pi953 & n45189;
  assign n45191 = ~pi1116 & po954;
  assign n45192 = ~pi625 & ~po954;
  assign n45193 = ~pi962 & ~n45192;
  assign po782 = ~n45191 & n45193;
  assign n45195 = ~pi1121 & po897;
  assign n45196 = ~pi626 & ~po897;
  assign n45197 = ~pi966 & ~n45196;
  assign po783 = ~n45195 & n45197;
  assign n45199 = ~pi1117 & po954;
  assign n45200 = ~pi627 & ~po954;
  assign n45201 = ~pi962 & ~n45200;
  assign po784 = ~n45199 & n45201;
  assign n45203 = ~pi1119 & po954;
  assign n45204 = ~pi628 & ~po954;
  assign n45205 = ~pi962 & ~n45204;
  assign po785 = ~n45203 & n45205;
  assign n45207 = ~pi1119 & po897;
  assign n45208 = ~pi629 & ~po897;
  assign n45209 = ~pi966 & ~n45208;
  assign po786 = ~n45207 & n45209;
  assign n45211 = ~pi1120 & po897;
  assign n45212 = ~pi630 & ~po897;
  assign n45213 = ~pi966 & ~n45212;
  assign po787 = ~n45211 & n45213;
  assign n45215 = pi631 & ~po954;
  assign n45216 = ~pi1113 & po954;
  assign n45217 = ~pi962 & ~n45216;
  assign po788 = ~n45215 & n45217;
  assign n45219 = pi632 & ~po954;
  assign n45220 = ~pi1115 & po954;
  assign n45221 = ~pi962 & ~n45220;
  assign po789 = ~n45219 & n45221;
  assign n45223 = ~pi1110 & po897;
  assign n45224 = ~pi633 & ~po897;
  assign n45225 = ~pi966 & ~n45224;
  assign po790 = ~n45223 & n45225;
  assign n45227 = ~pi1110 & po954;
  assign n45228 = ~pi634 & ~po954;
  assign n45229 = ~pi962 & ~n45228;
  assign po791 = ~n45227 & n45229;
  assign n45231 = pi635 & ~po954;
  assign n45232 = ~pi1112 & po954;
  assign n45233 = ~pi962 & ~n45232;
  assign po792 = ~n45231 & n45233;
  assign n45235 = ~pi1127 & po897;
  assign n45236 = ~pi636 & ~po897;
  assign n45237 = ~pi966 & ~n45236;
  assign po793 = ~n45235 & n45237;
  assign n45239 = ~pi1105 & po954;
  assign n45240 = ~pi637 & ~po954;
  assign n45241 = ~pi962 & ~n45240;
  assign po794 = ~n45239 & n45241;
  assign n45243 = ~pi1107 & po954;
  assign n45244 = ~pi638 & ~po954;
  assign n45245 = ~pi962 & ~n45244;
  assign po795 = ~n45243 & n45245;
  assign n45247 = ~pi1109 & po954;
  assign n45248 = ~pi639 & ~po954;
  assign n45249 = ~pi962 & ~n45248;
  assign po796 = ~n45247 & n45249;
  assign n45251 = ~pi1128 & po897;
  assign n45252 = ~pi640 & ~po897;
  assign n45253 = ~pi966 & ~n45252;
  assign po797 = ~n45251 & n45253;
  assign n45255 = ~pi1121 & po954;
  assign n45256 = ~pi641 & ~po954;
  assign n45257 = ~pi962 & ~n45256;
  assign po798 = ~n45255 & n45257;
  assign n45259 = ~pi1103 & po897;
  assign n45260 = ~pi642 & ~po897;
  assign n45261 = ~pi966 & ~n45260;
  assign po799 = ~n45259 & n45261;
  assign n45263 = ~pi1104 & po954;
  assign n45264 = ~pi643 & ~po954;
  assign n45265 = ~pi962 & ~n45264;
  assign po800 = ~n45263 & n45265;
  assign n45267 = ~pi1123 & po897;
  assign n45268 = ~pi644 & ~po897;
  assign n45269 = ~pi966 & ~n45268;
  assign po801 = ~n45267 & n45269;
  assign n45271 = ~pi1125 & po897;
  assign n45272 = ~pi645 & ~po897;
  assign n45273 = ~pi966 & ~n45272;
  assign po802 = ~n45271 & n45273;
  assign n45275 = pi646 & ~po954;
  assign n45276 = ~pi1114 & po954;
  assign n45277 = ~pi962 & ~n45276;
  assign po803 = ~n45275 & n45277;
  assign n45279 = ~pi1120 & po954;
  assign n45280 = ~pi647 & ~po954;
  assign n45281 = ~pi962 & ~n45280;
  assign po804 = ~n45279 & n45281;
  assign n45283 = ~pi1122 & po954;
  assign n45284 = ~pi648 & ~po954;
  assign n45285 = ~pi962 & ~n45284;
  assign po805 = ~n45283 & n45285;
  assign n45287 = pi649 & ~po954;
  assign n45288 = ~pi1126 & po954;
  assign n45289 = ~pi962 & ~n45288;
  assign po806 = ~n45287 & n45289;
  assign n45291 = pi650 & ~po954;
  assign n45292 = ~pi1127 & po954;
  assign n45293 = ~pi962 & ~n45292;
  assign po807 = ~n45291 & n45293;
  assign n45295 = ~pi1130 & po897;
  assign n45296 = ~pi651 & ~po897;
  assign n45297 = ~pi966 & ~n45296;
  assign po808 = ~n45295 & n45297;
  assign n45299 = ~pi1131 & po897;
  assign n45300 = ~pi652 & ~po897;
  assign n45301 = ~pi966 & ~n45300;
  assign po809 = ~n45299 & n45301;
  assign n45303 = ~pi1129 & po897;
  assign n45304 = ~pi653 & ~po897;
  assign n45305 = ~pi966 & ~n45304;
  assign po810 = ~n45303 & n45305;
  assign n45307 = pi654 & ~po954;
  assign n45308 = ~pi1130 & po954;
  assign n45309 = ~pi962 & ~n45308;
  assign po811 = ~n45307 & n45309;
  assign n45311 = pi655 & ~po954;
  assign n45312 = ~pi1124 & po954;
  assign n45313 = ~pi962 & ~n45312;
  assign po812 = ~n45311 & n45313;
  assign n45315 = ~pi1126 & po897;
  assign n45316 = ~pi656 & ~po897;
  assign n45317 = ~pi966 & ~n45316;
  assign po813 = ~n45315 & n45317;
  assign n45319 = pi657 & ~po954;
  assign n45320 = ~pi1131 & po954;
  assign n45321 = ~pi962 & ~n45320;
  assign po814 = ~n45319 & n45321;
  assign n45323 = ~pi1124 & po897;
  assign n45324 = ~pi658 & ~po897;
  assign n45325 = ~pi966 & ~n45324;
  assign po815 = ~n45323 & n45325;
  assign n45327 = pi266 & pi992;
  assign n45328 = ~pi280 & n45327;
  assign n45329 = ~pi269 & n45328;
  assign n45330 = ~pi281 & n45329;
  assign n45331 = ~pi282 & n45330;
  assign n45332 = ~pi270 & n45331;
  assign n45333 = ~pi277 & n45332;
  assign n45334 = ~pi264 & n45333;
  assign n45335 = ~pi265 & n45334;
  assign po959 = ~pi274 & n45335;
  assign n45337 = pi274 & ~n45335;
  assign po816 = ~po959 & ~n45337;
  assign n45339 = ~pi1118 & po954;
  assign n45340 = ~pi660 & ~po954;
  assign n45341 = ~pi962 & ~n45340;
  assign po817 = ~n45339 & n45341;
  assign n45343 = ~pi1101 & po954;
  assign n45344 = ~pi661 & ~po954;
  assign n45345 = ~pi962 & ~n45344;
  assign po818 = ~n45343 & n45345;
  assign n45347 = ~pi1102 & po954;
  assign n45348 = ~pi662 & ~po954;
  assign n45349 = ~pi962 & ~n45348;
  assign po819 = ~n45347 & n45349;
  assign n45351 = ~pi1137 & ~pi1138;
  assign n45352 = ~pi1134 & n45351;
  assign n45353 = ~pi634 & pi1136;
  assign n45354 = ~pi784 & ~pi1136;
  assign n45355 = pi1135 & ~n45354;
  assign n45356 = ~n45353 & n45355;
  assign n45357 = ~pi633 & pi1136;
  assign n45358 = ~pi815 & ~pi1136;
  assign n45359 = ~pi1135 & ~n45358;
  assign n45360 = ~n45357 & n45359;
  assign n45361 = ~n45356 & ~n45360;
  assign n45362 = n45352 & ~n45361;
  assign n45363 = pi1135 & ~pi1136;
  assign n45364 = pi1134 & n45351;
  assign n45365 = ~n45363 & n45364;
  assign n45366 = ~pi700 & pi1135;
  assign n45367 = pi1135 & n45351;
  assign n45368 = pi1136 & ~n45367;
  assign n45369 = ~pi766 & n45368;
  assign n45370 = ~pi855 & ~pi1136;
  assign n45371 = ~n45369 & ~n45370;
  assign n45372 = ~n45366 & n45371;
  assign n45373 = n45365 & n45372;
  assign n45374 = ~n45362 & ~n45373;
  assign n45375 = ~n7588 & ~n45374;
  assign n45376 = ~pi223 & ~pi224;
  assign n45377 = ~pi199 & ~pi257;
  assign n45378 = pi199 & ~pi1065;
  assign n45379 = ~n45377 & ~n45378;
  assign n45380 = ~n45376 & ~n45379;
  assign n45381 = n7588 & ~n45380;
  assign n45382 = ~pi592 & n7958;
  assign n45383 = pi464 & n45382;
  assign n45384 = pi588 & ~n45383;
  assign n45385 = ~pi591 & ~pi592;
  assign n45386 = pi590 & n45385;
  assign n45387 = pi323 & n45386;
  assign n45388 = ~pi591 & pi592;
  assign n45389 = pi365 & n45388;
  assign n45390 = pi591 & ~pi592;
  assign n45391 = pi334 & n45390;
  assign n45392 = ~n45389 & ~n45391;
  assign n45393 = ~pi590 & ~n45392;
  assign n45394 = ~pi588 & ~n45393;
  assign n45395 = ~n45387 & n45394;
  assign n45396 = ~n45384 & ~n45395;
  assign n45397 = n45376 & ~n45396;
  assign n45398 = n45381 & ~n45397;
  assign po820 = n45375 | n45398;
  assign n45400 = pi429 & n45382;
  assign n45401 = pi588 & ~n45400;
  assign n45402 = ~pi590 & pi591;
  assign n45403 = pi404 & n45402;
  assign n45404 = ~pi590 & pi592;
  assign n45405 = ~pi588 & ~n45404;
  assign n45406 = ~n45403 & n45405;
  assign n45407 = pi380 & ~pi591;
  assign n45408 = pi592 & ~n45407;
  assign n45409 = ~n45406 & ~n45408;
  assign n45410 = pi355 & n45386;
  assign n45411 = ~n45409 & ~n45410;
  assign n45412 = ~n45401 & ~n45411;
  assign n45413 = n45376 & n45412;
  assign n45414 = pi199 & ~pi1084;
  assign n45415 = ~pi199 & ~pi292;
  assign n45416 = ~n45376 & ~n45415;
  assign n45417 = ~n45414 & n45416;
  assign n45418 = ~n45413 & ~n45417;
  assign n45419 = n7588 & ~n45418;
  assign n45420 = ~n7588 & n45351;
  assign n45421 = pi662 & pi1135;
  assign n45422 = pi614 & ~pi1135;
  assign n45423 = pi1136 & ~n45422;
  assign n45424 = ~n45421 & n45423;
  assign n45425 = pi785 & pi1135;
  assign n45426 = pi811 & ~pi1135;
  assign n45427 = ~pi1136 & ~n45426;
  assign n45428 = ~n45425 & n45427;
  assign n45429 = ~n45424 & ~n45428;
  assign n45430 = ~pi1134 & ~n45429;
  assign n45431 = ~pi1135 & ~pi1136;
  assign n45432 = pi872 & n45431;
  assign n45433 = ~pi727 & pi1135;
  assign n45434 = ~pi772 & ~pi1135;
  assign n45435 = pi1136 & ~n45434;
  assign n45436 = ~n45433 & n45435;
  assign n45437 = pi1134 & ~n45436;
  assign n45438 = ~n45432 & n45437;
  assign n45439 = ~n45430 & ~n45438;
  assign n45440 = n45420 & n45439;
  assign po821 = n45419 | n45440;
  assign n45442 = ~pi1108 & po954;
  assign n45443 = ~pi665 & ~po954;
  assign n45444 = ~pi962 & ~n45443;
  assign po822 = ~n45442 & n45444;
  assign n45446 = ~pi638 & pi1135;
  assign n45447 = ~pi607 & ~pi1135;
  assign n45448 = pi1136 & ~n45447;
  assign n45449 = ~n45446 & n45448;
  assign n45450 = pi799 & ~pi1135;
  assign n45451 = ~pi790 & pi1135;
  assign n45452 = ~pi1136 & ~n45451;
  assign n45453 = ~n45450 & n45452;
  assign n45454 = ~n45449 & ~n45453;
  assign n45455 = n45352 & ~n45454;
  assign n45456 = ~pi873 & ~pi1136;
  assign n45457 = ~pi764 & n45368;
  assign n45458 = ~pi691 & pi1135;
  assign n45459 = ~n45457 & ~n45458;
  assign n45460 = ~n45456 & n45459;
  assign n45461 = n45365 & n45460;
  assign n45462 = ~n45455 & ~n45461;
  assign n45463 = ~n7588 & ~n45462;
  assign n45464 = pi199 & ~pi1044;
  assign n45465 = ~pi199 & ~pi297;
  assign n45466 = ~n45376 & ~n45465;
  assign n45467 = ~n45464 & n45466;
  assign n45468 = pi456 & n45402;
  assign n45469 = n45405 & ~n45468;
  assign n45470 = pi337 & ~pi591;
  assign n45471 = pi592 & ~n45470;
  assign n45472 = ~n45469 & ~n45471;
  assign n45473 = pi441 & n45386;
  assign n45474 = ~n45472 & ~n45473;
  assign n45475 = pi443 & n45382;
  assign n45476 = pi588 & ~n45475;
  assign n45477 = n45376 & ~n45476;
  assign n45478 = ~n45474 & n45477;
  assign n45479 = ~n45467 & ~n45478;
  assign n45480 = n7588 & ~n45479;
  assign po823 = n45463 | n45480;
  assign n45482 = pi444 & n45382;
  assign n45483 = pi588 & ~n45482;
  assign n45484 = pi319 & n45402;
  assign n45485 = n45405 & ~n45484;
  assign n45486 = pi338 & ~pi591;
  assign n45487 = pi592 & ~n45486;
  assign n45488 = ~n45485 & ~n45487;
  assign n45489 = pi458 & n45386;
  assign n45490 = ~n45488 & ~n45489;
  assign n45491 = ~n45483 & ~n45490;
  assign n45492 = n45376 & n45491;
  assign n45493 = pi199 & ~pi1072;
  assign n45494 = ~pi199 & ~pi294;
  assign n45495 = ~n45376 & ~n45494;
  assign n45496 = ~n45493 & n45495;
  assign n45497 = ~n45492 & ~n45496;
  assign n45498 = n7588 & ~n45497;
  assign n45499 = pi681 & pi1136;
  assign n45500 = pi792 & ~pi1136;
  assign n45501 = pi1135 & ~n45500;
  assign n45502 = ~n45499 & n45501;
  assign n45503 = pi642 & pi1136;
  assign n45504 = ~pi809 & ~pi1136;
  assign n45505 = ~pi1135 & ~n45504;
  assign n45506 = ~n45503 & n45505;
  assign n45507 = ~n45502 & ~n45506;
  assign n45508 = ~pi1134 & ~n45507;
  assign n45509 = pi871 & n45431;
  assign n45510 = ~pi699 & pi1135;
  assign n45511 = ~pi763 & ~pi1135;
  assign n45512 = pi1136 & ~n45511;
  assign n45513 = ~n45510 & n45512;
  assign n45514 = pi1134 & ~n45513;
  assign n45515 = ~n45509 & n45514;
  assign n45516 = n45420 & ~n45515;
  assign n45517 = ~n45508 & n45516;
  assign po824 = n45498 | n45517;
  assign n45519 = ~pi680 & pi1135;
  assign n45520 = ~pi603 & ~pi1135;
  assign n45521 = pi1136 & ~n45520;
  assign n45522 = ~n45519 & n45521;
  assign n45523 = ~pi778 & pi1135;
  assign n45524 = ~pi981 & ~pi1135;
  assign n45525 = ~pi1136 & ~n45524;
  assign n45526 = ~n45523 & n45525;
  assign n45527 = ~n45522 & ~n45526;
  assign n45528 = n45352 & ~n45527;
  assign n45529 = ~pi837 & ~pi1136;
  assign n45530 = ~pi759 & n45368;
  assign n45531 = ~pi696 & pi1135;
  assign n45532 = ~n45530 & ~n45531;
  assign n45533 = ~n45529 & n45532;
  assign n45534 = n45365 & n45533;
  assign n45535 = ~n45528 & ~n45534;
  assign n45536 = ~n7588 & ~n45535;
  assign n45537 = pi199 & ~pi1049;
  assign n45538 = ~pi199 & ~pi291;
  assign n45539 = ~n45376 & ~n45538;
  assign n45540 = ~n45537 & n45539;
  assign n45541 = pi414 & n45382;
  assign n45542 = pi588 & ~n45541;
  assign n45543 = pi390 & n45402;
  assign n45544 = n45405 & ~n45543;
  assign n45545 = pi363 & ~pi591;
  assign n45546 = pi592 & ~n45545;
  assign n45547 = ~n45544 & ~n45546;
  assign n45548 = pi342 & n45386;
  assign n45549 = ~n45547 & ~n45548;
  assign n45550 = ~n45542 & ~n45549;
  assign n45551 = n45376 & n45550;
  assign n45552 = ~n45540 & ~n45551;
  assign n45553 = n7588 & ~n45552;
  assign po825 = n45536 | n45553;
  assign n45555 = pi669 & ~po954;
  assign n45556 = ~pi1125 & po954;
  assign n45557 = ~pi962 & ~n45556;
  assign po826 = ~n45555 & n45557;
  assign n45559 = pi199 & ~pi1062;
  assign n45560 = ~pi199 & ~pi258;
  assign n45561 = ~n45376 & ~n45560;
  assign n45562 = ~n45559 & n45561;
  assign n45563 = pi415 & n45382;
  assign n45564 = pi588 & ~n45563;
  assign n45565 = pi343 & n45386;
  assign n45566 = pi364 & n45388;
  assign n45567 = pi391 & n45390;
  assign n45568 = ~n45566 & ~n45567;
  assign n45569 = ~pi590 & ~n45568;
  assign n45570 = ~pi588 & ~n45569;
  assign n45571 = ~n45565 & n45570;
  assign n45572 = ~n45564 & ~n45571;
  assign n45573 = n45376 & n45572;
  assign n45574 = ~n45562 & ~n45573;
  assign n45575 = n7588 & ~n45574;
  assign n45576 = ~pi852 & ~pi1136;
  assign n45577 = pi745 & n45368;
  assign n45578 = pi723 & pi1135;
  assign n45579 = ~n45577 & ~n45578;
  assign n45580 = ~n45576 & n45579;
  assign n45581 = n45365 & n45580;
  assign n45582 = pi695 & pi1135;
  assign n45583 = ~pi612 & ~pi1135;
  assign n45584 = ~pi1134 & ~n45583;
  assign n45585 = pi1136 & n45351;
  assign n45586 = n45584 & n45585;
  assign n45587 = ~n45582 & n45586;
  assign n45588 = ~n45581 & ~n45587;
  assign n45589 = ~n7588 & ~n45588;
  assign po827 = n45575 | n45589;
  assign n45591 = pi199 & ~pi1040;
  assign n45592 = ~pi199 & ~pi261;
  assign n45593 = ~n45376 & ~n45592;
  assign n45594 = ~n45591 & n45593;
  assign n45595 = pi453 & n45382;
  assign n45596 = pi588 & ~n45595;
  assign n45597 = pi327 & n45386;
  assign n45598 = pi447 & n45388;
  assign n45599 = pi333 & n45390;
  assign n45600 = ~n45598 & ~n45599;
  assign n45601 = ~pi590 & ~n45600;
  assign n45602 = ~pi588 & ~n45601;
  assign n45603 = ~n45597 & n45602;
  assign n45604 = ~n45596 & ~n45603;
  assign n45605 = n45376 & n45604;
  assign n45606 = ~n45594 & ~n45605;
  assign n45607 = n7588 & ~n45606;
  assign n45608 = ~pi865 & ~pi1136;
  assign n45609 = pi741 & n45368;
  assign n45610 = pi724 & pi1135;
  assign n45611 = ~n45609 & ~n45610;
  assign n45612 = ~n45608 & n45611;
  assign n45613 = n45365 & n45612;
  assign n45614 = pi646 & pi1135;
  assign n45615 = ~pi611 & ~pi1135;
  assign n45616 = ~pi1134 & ~n45615;
  assign n45617 = n45585 & n45616;
  assign n45618 = ~n45614 & n45617;
  assign n45619 = ~n45613 & ~n45618;
  assign n45620 = ~n7588 & ~n45619;
  assign po828 = n45607 | n45620;
  assign n45622 = ~pi661 & pi1135;
  assign n45623 = ~pi616 & ~pi1135;
  assign n45624 = pi1136 & ~n45623;
  assign n45625 = ~n45622 & n45624;
  assign n45626 = ~pi781 & pi1135;
  assign n45627 = ~pi808 & ~pi1135;
  assign n45628 = ~pi1136 & ~n45627;
  assign n45629 = ~n45626 & n45628;
  assign n45630 = ~n45625 & ~n45629;
  assign n45631 = n45352 & ~n45630;
  assign n45632 = ~pi850 & ~pi1136;
  assign n45633 = ~pi758 & n45368;
  assign n45634 = ~pi736 & pi1135;
  assign n45635 = ~n45633 & ~n45634;
  assign n45636 = ~n45632 & n45635;
  assign n45637 = n45365 & n45636;
  assign n45638 = ~n45631 & ~n45637;
  assign n45639 = ~n7588 & ~n45638;
  assign n45640 = pi199 & ~pi1048;
  assign n45641 = ~pi199 & ~pi290;
  assign n45642 = ~n45376 & ~n45641;
  assign n45643 = ~n45640 & n45642;
  assign n45644 = pi422 & n45382;
  assign n45645 = pi588 & ~n45644;
  assign n45646 = pi397 & n45402;
  assign n45647 = n45405 & ~n45646;
  assign n45648 = pi372 & ~pi591;
  assign n45649 = pi592 & ~n45648;
  assign n45650 = ~n45647 & ~n45649;
  assign n45651 = pi320 & n45386;
  assign n45652 = ~n45650 & ~n45651;
  assign n45653 = ~n45645 & ~n45652;
  assign n45654 = n45376 & n45653;
  assign n45655 = ~n45643 & ~n45654;
  assign n45656 = n7588 & ~n45655;
  assign po829 = n45639 | n45656;
  assign n45658 = ~pi637 & pi1135;
  assign n45659 = ~pi617 & ~pi1135;
  assign n45660 = pi1136 & ~n45659;
  assign n45661 = ~n45658 & n45660;
  assign n45662 = pi814 & ~pi1135;
  assign n45663 = ~pi788 & pi1135;
  assign n45664 = ~pi1136 & ~n45663;
  assign n45665 = ~n45662 & n45664;
  assign n45666 = ~n45661 & ~n45665;
  assign n45667 = n45352 & ~n45666;
  assign n45668 = ~pi866 & ~pi1136;
  assign n45669 = ~pi749 & n45368;
  assign n45670 = ~pi706 & pi1135;
  assign n45671 = ~n45669 & ~n45670;
  assign n45672 = ~n45668 & n45671;
  assign n45673 = n45365 & n45672;
  assign n45674 = ~n45667 & ~n45673;
  assign n45675 = ~n7588 & ~n45674;
  assign n45676 = pi199 & ~pi1053;
  assign n45677 = ~pi199 & ~pi295;
  assign n45678 = ~n45376 & ~n45677;
  assign n45679 = ~n45676 & n45678;
  assign n45680 = pi435 & n45382;
  assign n45681 = pi588 & ~n45680;
  assign n45682 = pi411 & n45402;
  assign n45683 = n45405 & ~n45682;
  assign n45684 = pi387 & ~pi591;
  assign n45685 = pi592 & ~n45684;
  assign n45686 = ~n45683 & ~n45685;
  assign n45687 = pi452 & n45386;
  assign n45688 = ~n45686 & ~n45687;
  assign n45689 = ~n45681 & ~n45688;
  assign n45690 = n45376 & n45689;
  assign n45691 = ~n45679 & ~n45690;
  assign n45692 = n7588 & ~n45691;
  assign po830 = n45675 | n45692;
  assign n45694 = pi199 & ~pi1070;
  assign n45695 = ~pi199 & ~pi256;
  assign n45696 = ~n45376 & ~n45695;
  assign n45697 = ~n45694 & n45696;
  assign n45698 = pi437 & n45382;
  assign n45699 = pi588 & ~n45698;
  assign n45700 = pi362 & n45386;
  assign n45701 = pi336 & n45388;
  assign n45702 = pi463 & n45390;
  assign n45703 = ~n45701 & ~n45702;
  assign n45704 = ~pi590 & ~n45703;
  assign n45705 = ~pi588 & ~n45704;
  assign n45706 = ~n45700 & n45705;
  assign n45707 = ~n45699 & ~n45706;
  assign n45708 = n45376 & n45707;
  assign n45709 = ~n45697 & ~n45708;
  assign n45710 = n7588 & ~n45709;
  assign n45711 = pi639 & pi1135;
  assign n45712 = pi622 & ~pi1135;
  assign n45713 = pi1136 & ~n45712;
  assign n45714 = ~n45711 & n45713;
  assign n45715 = pi783 & pi1135;
  assign n45716 = pi804 & ~pi1135;
  assign n45717 = ~pi1136 & ~n45716;
  assign n45718 = ~n45715 & n45717;
  assign n45719 = ~n45714 & ~n45718;
  assign n45720 = ~pi1134 & ~n45719;
  assign n45721 = pi859 & n45431;
  assign n45722 = ~pi735 & pi1135;
  assign n45723 = ~pi743 & ~pi1135;
  assign n45724 = pi1136 & ~n45723;
  assign n45725 = ~n45722 & n45724;
  assign n45726 = pi1134 & ~n45725;
  assign n45727 = ~n45721 & n45726;
  assign n45728 = n45420 & ~n45727;
  assign n45729 = ~n45720 & n45728;
  assign po831 = n45710 | n45729;
  assign n45731 = pi876 & n45431;
  assign n45732 = ~pi730 & pi1135;
  assign n45733 = ~pi748 & ~pi1135;
  assign n45734 = pi1136 & ~n45733;
  assign n45735 = ~n45732 & n45734;
  assign n45736 = ~n45731 & ~n45735;
  assign n45737 = n45364 & ~n45736;
  assign n45738 = ~pi623 & n45368;
  assign n45739 = pi789 & n45363;
  assign n45740 = ~pi803 & ~pi1135;
  assign n45741 = ~pi710 & pi1135;
  assign n45742 = pi1136 & ~n45741;
  assign n45743 = ~n45740 & ~n45742;
  assign n45744 = ~n45739 & n45743;
  assign n45745 = ~n45738 & ~n45744;
  assign n45746 = n45352 & n45745;
  assign n45747 = ~n45737 & ~n45746;
  assign n45748 = ~n7588 & ~n45747;
  assign n45749 = pi199 & ~pi1037;
  assign n45750 = ~pi199 & ~pi296;
  assign n45751 = ~n45376 & ~n45750;
  assign n45752 = ~n45749 & n45751;
  assign n45753 = pi436 & n45382;
  assign n45754 = pi588 & ~n45753;
  assign n45755 = pi412 & n45402;
  assign n45756 = n45405 & ~n45755;
  assign n45757 = pi388 & ~pi591;
  assign n45758 = pi592 & ~n45757;
  assign n45759 = ~n45756 & ~n45758;
  assign n45760 = pi455 & n45386;
  assign n45761 = ~n45759 & ~n45760;
  assign n45762 = ~n45754 & ~n45761;
  assign n45763 = n45376 & n45762;
  assign n45764 = ~n45752 & ~n45763;
  assign n45765 = n7588 & ~n45764;
  assign po832 = n45748 | n45765;
  assign n45767 = ~pi643 & pi1135;
  assign n45768 = ~pi606 & ~pi1135;
  assign n45769 = pi1136 & ~n45768;
  assign n45770 = ~n45767 & n45769;
  assign n45771 = pi812 & ~pi1135;
  assign n45772 = ~pi787 & pi1135;
  assign n45773 = ~pi1136 & ~n45772;
  assign n45774 = ~n45771 & n45773;
  assign n45775 = ~n45770 & ~n45774;
  assign n45776 = n45352 & ~n45775;
  assign n45777 = ~pi881 & ~pi1136;
  assign n45778 = ~pi746 & n45368;
  assign n45779 = ~pi729 & pi1135;
  assign n45780 = ~n45778 & ~n45779;
  assign n45781 = ~n45777 & n45780;
  assign n45782 = n45365 & n45781;
  assign n45783 = ~n45776 & ~n45782;
  assign n45784 = ~n7588 & ~n45783;
  assign n45785 = pi199 & ~pi1059;
  assign n45786 = ~pi199 & ~pi293;
  assign n45787 = ~n45376 & ~n45786;
  assign n45788 = ~n45785 & n45787;
  assign n45789 = pi434 & n45382;
  assign n45790 = pi588 & ~n45789;
  assign n45791 = pi410 & n45402;
  assign n45792 = n45405 & ~n45791;
  assign n45793 = pi386 & ~pi591;
  assign n45794 = pi592 & ~n45793;
  assign n45795 = ~n45792 & ~n45794;
  assign n45796 = pi361 & n45386;
  assign n45797 = ~n45795 & ~n45796;
  assign n45798 = ~n45790 & ~n45797;
  assign n45799 = n45376 & n45798;
  assign n45800 = ~n45788 & ~n45799;
  assign n45801 = n7588 & ~n45800;
  assign po833 = n45784 | n45801;
  assign n45803 = pi199 & ~pi1069;
  assign n45804 = ~pi199 & ~pi259;
  assign n45805 = ~n45376 & ~n45804;
  assign n45806 = ~n45803 & n45805;
  assign n45807 = pi416 & n45382;
  assign n45808 = pi588 & ~n45807;
  assign n45809 = pi344 & n45386;
  assign n45810 = pi366 & n45388;
  assign n45811 = pi335 & n45390;
  assign n45812 = ~n45810 & ~n45811;
  assign n45813 = ~pi590 & ~n45812;
  assign n45814 = ~pi588 & ~n45813;
  assign n45815 = ~n45809 & n45814;
  assign n45816 = ~n45808 & ~n45815;
  assign n45817 = n45376 & n45816;
  assign n45818 = ~n45806 & ~n45817;
  assign n45819 = n7588 & ~n45818;
  assign n45820 = ~pi870 & ~pi1136;
  assign n45821 = pi742 & n45368;
  assign n45822 = pi704 & pi1135;
  assign n45823 = ~n45821 & ~n45822;
  assign n45824 = ~n45820 & n45823;
  assign n45825 = n45365 & n45824;
  assign n45826 = pi635 & pi1135;
  assign n45827 = ~pi620 & ~pi1135;
  assign n45828 = ~pi1134 & ~n45827;
  assign n45829 = n45585 & n45828;
  assign n45830 = ~n45826 & n45829;
  assign n45831 = ~n45825 & ~n45830;
  assign n45832 = ~n7588 & ~n45831;
  assign po834 = n45819 | n45832;
  assign n45834 = pi199 & ~pi1067;
  assign n45835 = ~pi199 & ~pi260;
  assign n45836 = ~n45376 & ~n45835;
  assign n45837 = ~n45834 & n45836;
  assign n45838 = pi418 & n45382;
  assign n45839 = pi588 & ~n45838;
  assign n45840 = pi346 & n45386;
  assign n45841 = pi368 & n45388;
  assign n45842 = pi393 & n45390;
  assign n45843 = ~n45841 & ~n45842;
  assign n45844 = ~pi590 & ~n45843;
  assign n45845 = ~pi588 & ~n45844;
  assign n45846 = ~n45840 & n45845;
  assign n45847 = ~n45839 & ~n45846;
  assign n45848 = n45376 & n45847;
  assign n45849 = ~n45837 & ~n45848;
  assign n45850 = n7588 & ~n45849;
  assign n45851 = ~pi856 & ~pi1136;
  assign n45852 = pi760 & n45368;
  assign n45853 = pi688 & pi1135;
  assign n45854 = ~n45852 & ~n45853;
  assign n45855 = ~n45851 & n45854;
  assign n45856 = n45365 & n45855;
  assign n45857 = pi632 & pi1135;
  assign n45858 = ~pi613 & ~pi1135;
  assign n45859 = ~pi1134 & ~n45858;
  assign n45860 = n45585 & n45859;
  assign n45861 = ~n45857 & n45860;
  assign n45862 = ~n45856 & ~n45861;
  assign n45863 = ~n7588 & ~n45862;
  assign po835 = n45850 | n45863;
  assign n45865 = pi199 & ~pi1036;
  assign n45866 = ~pi199 & ~pi255;
  assign n45867 = ~n45376 & ~n45866;
  assign n45868 = ~n45865 & n45867;
  assign n45869 = pi438 & n45382;
  assign n45870 = pi588 & ~n45869;
  assign n45871 = pi450 & n45386;
  assign n45872 = pi389 & n45388;
  assign n45873 = pi413 & n45390;
  assign n45874 = ~n45872 & ~n45873;
  assign n45875 = ~pi590 & ~n45874;
  assign n45876 = ~pi588 & ~n45875;
  assign n45877 = ~n45871 & n45876;
  assign n45878 = ~n45870 & ~n45877;
  assign n45879 = n45376 & n45878;
  assign n45880 = ~n45868 & ~n45879;
  assign n45881 = n7588 & ~n45880;
  assign n45882 = ~pi665 & pi1136;
  assign n45883 = ~pi791 & ~pi1136;
  assign n45884 = pi1135 & ~n45883;
  assign n45885 = ~n45882 & n45884;
  assign n45886 = ~pi621 & pi1136;
  assign n45887 = ~pi810 & ~pi1136;
  assign n45888 = ~pi1135 & ~n45887;
  assign n45889 = ~n45886 & n45888;
  assign n45890 = ~n45885 & ~n45889;
  assign n45891 = n45352 & ~n45890;
  assign n45892 = ~pi690 & pi1135;
  assign n45893 = ~pi739 & n45368;
  assign n45894 = ~pi874 & ~pi1136;
  assign n45895 = ~n45893 & ~n45894;
  assign n45896 = ~n45892 & n45895;
  assign n45897 = n45365 & n45896;
  assign n45898 = ~n45891 & ~n45897;
  assign n45899 = ~n7588 & ~n45898;
  assign po836 = n45881 | n45899;
  assign n45901 = ~pi1100 & po954;
  assign n45902 = ~pi680 & ~po954;
  assign n45903 = ~pi962 & ~n45902;
  assign po837 = ~n45901 & n45903;
  assign n45905 = ~pi1103 & po954;
  assign n45906 = ~pi681 & ~po954;
  assign n45907 = ~pi962 & ~n45906;
  assign po838 = ~n45905 & n45907;
  assign n45909 = pi199 & ~pi1039;
  assign n45910 = ~pi199 & ~pi251;
  assign n45911 = ~n45376 & ~n45910;
  assign n45912 = ~n45909 & n45911;
  assign n45913 = pi417 & n45382;
  assign n45914 = pi588 & ~n45913;
  assign n45915 = pi345 & n45386;
  assign n45916 = pi367 & n45388;
  assign n45917 = pi392 & n45390;
  assign n45918 = ~n45916 & ~n45917;
  assign n45919 = ~pi590 & ~n45918;
  assign n45920 = ~pi588 & ~n45919;
  assign n45921 = ~n45915 & n45920;
  assign n45922 = ~n45914 & ~n45921;
  assign n45923 = n45376 & n45922;
  assign n45924 = ~n45912 & ~n45923;
  assign n45925 = n7588 & ~n45924;
  assign n45926 = ~pi848 & ~pi1136;
  assign n45927 = pi757 & n45368;
  assign n45928 = pi686 & pi1135;
  assign n45929 = ~n45927 & ~n45928;
  assign n45930 = ~n45926 & n45929;
  assign n45931 = n45365 & n45930;
  assign n45932 = pi631 & pi1135;
  assign n45933 = ~pi610 & ~pi1135;
  assign n45934 = ~pi1134 & ~n45933;
  assign n45935 = n45585 & n45934;
  assign n45936 = ~n45932 & n45935;
  assign n45937 = ~n45931 & ~n45936;
  assign n45938 = ~n7588 & ~n45937;
  assign po839 = n45925 | n45938;
  assign po980 = pi953 & n45189;
  assign n45941 = pi684 & ~po980;
  assign n45942 = ~pi1130 & po980;
  assign n45943 = ~pi962 & ~n45942;
  assign po841 = ~n45941 & n45943;
  assign n45945 = pi590 & ~pi592;
  assign n45946 = pi357 & n45945;
  assign n45947 = pi382 & n45404;
  assign n45948 = ~n45946 & ~n45947;
  assign n45949 = ~pi591 & ~n45948;
  assign n45950 = ~pi590 & n45390;
  assign n45951 = pi406 & n45950;
  assign n45952 = ~n45949 & ~n45951;
  assign n45953 = ~pi588 & ~n45952;
  assign n45954 = pi588 & ~pi590;
  assign n45955 = pi430 & n45385;
  assign n45956 = n45954 & n45955;
  assign n45957 = ~n45953 & ~n45956;
  assign n45958 = n45376 & ~n45957;
  assign n45959 = pi199 & ~pi1076;
  assign n45960 = ~n45376 & ~n45959;
  assign n45961 = ~n41689 & n45960;
  assign n45962 = ~n45958 & ~n45961;
  assign n45963 = n7588 & ~n45962;
  assign n45964 = pi860 & n45431;
  assign n45965 = pi728 & pi1135;
  assign n45966 = pi744 & ~pi1135;
  assign n45967 = pi1136 & ~n45966;
  assign n45968 = ~n45965 & n45967;
  assign n45969 = ~n45964 & ~n45968;
  assign n45970 = n45364 & ~n45969;
  assign n45971 = pi1136 & ~n45351;
  assign n45972 = ~pi1134 & ~n45971;
  assign n45973 = pi657 & pi1135;
  assign n45974 = ~pi652 & ~pi1135;
  assign n45975 = pi1136 & ~n45974;
  assign n45976 = ~n45973 & n45975;
  assign n45977 = pi813 & n45351;
  assign n45978 = n45431 & n45977;
  assign n45979 = ~n45976 & ~n45978;
  assign n45980 = n45972 & ~n45979;
  assign n45981 = ~n45970 & ~n45980;
  assign n45982 = ~n7588 & ~n45981;
  assign po842 = n45963 | n45982;
  assign n45984 = pi686 & ~po980;
  assign n45985 = ~pi1113 & po980;
  assign n45986 = ~pi962 & ~n45985;
  assign po843 = ~n45984 & n45986;
  assign n45988 = ~pi1127 & po980;
  assign n45989 = ~pi687 & ~po980;
  assign n45990 = ~pi962 & ~n45989;
  assign po844 = ~n45988 & n45990;
  assign n45992 = pi688 & ~po980;
  assign n45993 = ~pi1115 & po980;
  assign n45994 = ~pi962 & ~n45993;
  assign po845 = ~n45992 & n45994;
  assign n45996 = pi351 & n45945;
  assign n45997 = pi376 & n45404;
  assign n45998 = ~n45996 & ~n45997;
  assign n45999 = ~pi591 & ~n45998;
  assign n46000 = pi401 & n45950;
  assign n46001 = ~n45999 & ~n46000;
  assign n46002 = ~pi588 & ~n46001;
  assign n46003 = pi426 & n45385;
  assign n46004 = n45954 & n46003;
  assign n46005 = ~n46002 & ~n46004;
  assign n46006 = n45376 & ~n46005;
  assign n46007 = ~pi199 & n41658;
  assign n46008 = pi199 & ~pi1079;
  assign n46009 = ~n45376 & ~n46008;
  assign n46010 = ~n46007 & n46009;
  assign n46011 = ~n46006 & ~n46010;
  assign n46012 = n7588 & ~n46011;
  assign n46013 = pi798 & n45431;
  assign n46014 = pi655 & pi1135;
  assign n46015 = ~pi658 & ~pi1135;
  assign n46016 = pi1136 & ~n46015;
  assign n46017 = ~n46014 & n46016;
  assign n46018 = ~n46013 & ~n46017;
  assign n46019 = n45352 & ~n46018;
  assign n46020 = ~pi843 & ~pi1136;
  assign n46021 = pi752 & n45368;
  assign n46022 = ~pi703 & pi1135;
  assign n46023 = ~n46021 & ~n46022;
  assign n46024 = ~n46020 & n46023;
  assign n46025 = n45365 & n46024;
  assign n46026 = ~n46019 & ~n46025;
  assign n46027 = ~n7588 & ~n46026;
  assign po846 = n46012 | n46027;
  assign n46029 = ~pi1108 & po980;
  assign n46030 = ~pi690 & ~po980;
  assign n46031 = ~pi962 & ~n46030;
  assign po847 = ~n46029 & n46031;
  assign n46033 = ~pi1107 & po980;
  assign n46034 = ~pi691 & ~po980;
  assign n46035 = ~pi962 & ~n46034;
  assign po848 = ~n46033 & n46035;
  assign n46037 = pi352 & n45945;
  assign n46038 = pi317 & n45404;
  assign n46039 = ~n46037 & ~n46038;
  assign n46040 = ~pi591 & ~n46039;
  assign n46041 = pi402 & n45950;
  assign n46042 = ~n46040 & ~n46041;
  assign n46043 = ~pi588 & ~n46042;
  assign n46044 = pi427 & n45385;
  assign n46045 = n45954 & n46044;
  assign n46046 = ~n46043 & ~n46045;
  assign n46047 = n45376 & ~n46046;
  assign n46048 = ~pi199 & n41670;
  assign n46049 = pi199 & ~pi1078;
  assign n46050 = ~n45376 & ~n46049;
  assign n46051 = ~n46048 & n46050;
  assign n46052 = ~n46047 & ~n46051;
  assign n46053 = n7588 & ~n46052;
  assign n46054 = pi844 & n45431;
  assign n46055 = pi770 & ~pi1135;
  assign n46056 = ~pi726 & pi1135;
  assign n46057 = pi1136 & ~n46056;
  assign n46058 = ~n46055 & n46057;
  assign n46059 = pi1134 & ~n46058;
  assign n46060 = ~n46054 & n46059;
  assign n46061 = pi801 & n45431;
  assign n46062 = ~pi656 & ~pi1135;
  assign n46063 = pi649 & pi1135;
  assign n46064 = ~n46062 & ~n46063;
  assign n46065 = pi1136 & n46064;
  assign n46066 = ~pi1134 & ~n46065;
  assign n46067 = ~n46061 & n46066;
  assign n46068 = ~n46060 & ~n46067;
  assign n46069 = n45420 & n46068;
  assign po849 = n46053 | n46069;
  assign n46071 = pi693 & ~po954;
  assign n46072 = ~pi1129 & po954;
  assign n46073 = ~pi962 & ~n46072;
  assign po850 = ~n46071 & n46073;
  assign n46075 = pi694 & ~po980;
  assign n46076 = ~pi1128 & po980;
  assign n46077 = ~pi962 & ~n46076;
  assign po851 = ~n46075 & n46077;
  assign n46079 = pi695 & ~po954;
  assign n46080 = ~pi1111 & po954;
  assign n46081 = ~pi962 & ~n46080;
  assign po852 = ~n46079 & n46081;
  assign n46083 = ~pi1100 & po980;
  assign n46084 = ~pi696 & ~po980;
  assign n46085 = ~pi962 & ~n46084;
  assign po853 = ~n46083 & n46085;
  assign n46087 = pi697 & ~po980;
  assign n46088 = ~pi1129 & po980;
  assign n46089 = ~pi962 & ~n46088;
  assign po854 = ~n46087 & n46089;
  assign n46091 = pi698 & ~po980;
  assign n46092 = ~pi1116 & po980;
  assign n46093 = ~pi962 & ~n46092;
  assign po855 = ~n46091 & n46093;
  assign n46095 = ~pi1103 & po980;
  assign n46096 = ~pi699 & ~po980;
  assign n46097 = ~pi962 & ~n46096;
  assign po856 = ~n46095 & n46097;
  assign n46099 = ~pi1110 & po980;
  assign n46100 = ~pi700 & ~po980;
  assign n46101 = ~pi962 & ~n46100;
  assign po857 = ~n46099 & n46101;
  assign n46103 = pi701 & ~po980;
  assign n46104 = ~pi1123 & po980;
  assign n46105 = ~pi962 & ~n46104;
  assign po858 = ~n46103 & n46105;
  assign n46107 = pi702 & ~po980;
  assign n46108 = ~pi1117 & po980;
  assign n46109 = ~pi962 & ~n46108;
  assign po859 = ~n46107 & n46109;
  assign n46111 = ~pi1124 & po980;
  assign n46112 = ~pi703 & ~po980;
  assign n46113 = ~pi962 & ~n46112;
  assign po860 = ~n46111 & n46113;
  assign n46115 = pi704 & ~po980;
  assign n46116 = ~pi1112 & po980;
  assign n46117 = ~pi962 & ~n46116;
  assign po861 = ~n46115 & n46117;
  assign n46119 = ~pi1125 & po980;
  assign n46120 = ~pi705 & ~po980;
  assign n46121 = ~pi962 & ~n46120;
  assign po862 = ~n46119 & n46121;
  assign n46123 = ~pi1105 & po980;
  assign n46124 = ~pi706 & ~po980;
  assign n46125 = ~pi962 & ~n46124;
  assign po863 = ~n46123 & n46125;
  assign n46127 = pi370 & n45388;
  assign n46128 = pi395 & n45390;
  assign n46129 = ~n46127 & ~n46128;
  assign n46130 = ~pi590 & ~n46129;
  assign n46131 = pi347 & n45386;
  assign n46132 = ~n46130 & ~n46131;
  assign n46133 = ~pi588 & n45376;
  assign n46134 = ~n46132 & n46133;
  assign n46135 = pi199 & ~pi1055;
  assign n46136 = pi200 & pi1048;
  assign n46137 = ~pi200 & pi304;
  assign n46138 = ~pi199 & ~n46137;
  assign n46139 = ~n46136 & n46138;
  assign n46140 = ~n46135 & ~n46139;
  assign n46141 = ~n45376 & n46140;
  assign n46142 = n45376 & n45382;
  assign n46143 = pi420 & pi588;
  assign n46144 = n46142 & n46143;
  assign n46145 = ~n46141 & ~n46144;
  assign n46146 = ~n46134 & n46145;
  assign n46147 = n7588 & ~n46146;
  assign n46148 = ~pi627 & pi1135;
  assign n46149 = ~pi618 & ~pi1135;
  assign n46150 = ~pi1134 & ~n46149;
  assign n46151 = n45585 & n46150;
  assign n46152 = ~n46148 & n46151;
  assign n46153 = ~pi847 & ~pi1136;
  assign n46154 = pi753 & n45368;
  assign n46155 = pi702 & pi1135;
  assign n46156 = ~n46154 & ~n46155;
  assign n46157 = ~n46153 & n46156;
  assign n46158 = n45365 & n46157;
  assign n46159 = ~n46152 & ~n46158;
  assign n46160 = ~n7588 & ~n46159;
  assign po864 = n46147 | n46160;
  assign n46162 = n45376 & n45388;
  assign n46163 = pi442 & n46162;
  assign n46164 = pi328 & n45390;
  assign n46165 = n45376 & n46164;
  assign n46166 = ~n46163 & ~n46165;
  assign n46167 = ~pi590 & ~n46166;
  assign n46168 = pi321 & n45376;
  assign n46169 = n45386 & n46168;
  assign n46170 = ~n46167 & ~n46169;
  assign n46171 = ~pi588 & ~n46170;
  assign n46172 = pi199 & ~pi1058;
  assign n46173 = pi200 & pi1084;
  assign n46174 = ~pi200 & pi305;
  assign n46175 = ~pi199 & ~n46174;
  assign n46176 = ~n46173 & n46175;
  assign n46177 = ~n45376 & ~n46176;
  assign n46178 = ~n46172 & n46177;
  assign n46179 = n45376 & n45385;
  assign n46180 = pi459 & n46179;
  assign n46181 = n45954 & n46180;
  assign n46182 = n7588 & ~n46181;
  assign n46183 = ~n46178 & n46182;
  assign n46184 = ~n46171 & n46183;
  assign n46185 = pi709 & pi1135;
  assign n46186 = pi754 & n45368;
  assign n46187 = ~pi857 & ~pi1136;
  assign n46188 = ~n46186 & ~n46187;
  assign n46189 = ~n46185 & n46188;
  assign n46190 = n45365 & n46189;
  assign n46191 = ~pi609 & ~pi1135;
  assign n46192 = ~pi1134 & ~n46191;
  assign n46193 = ~pi660 & pi1135;
  assign n46194 = n45585 & ~n46193;
  assign n46195 = n46192 & n46194;
  assign n46196 = ~n7588 & ~n46195;
  assign n46197 = ~n46190 & n46196;
  assign po865 = ~n46184 & ~n46197;
  assign n46199 = pi709 & ~po980;
  assign n46200 = ~pi1118 & po980;
  assign n46201 = ~pi962 & ~n46200;
  assign po866 = ~n46199 & n46201;
  assign n46203 = ~pi1106 & po954;
  assign n46204 = ~pi710 & ~po954;
  assign n46205 = ~pi962 & ~n46204;
  assign po867 = ~n46203 & n46205;
  assign n46207 = pi373 & n45388;
  assign n46208 = pi398 & n45390;
  assign n46209 = ~n46207 & ~n46208;
  assign n46210 = ~pi590 & ~n46209;
  assign n46211 = pi348 & n45386;
  assign n46212 = ~n46210 & ~n46211;
  assign n46213 = n46133 & ~n46212;
  assign n46214 = pi199 & ~pi1087;
  assign n46215 = pi200 & pi1059;
  assign n46216 = ~pi200 & pi306;
  assign n46217 = ~pi199 & ~n46216;
  assign n46218 = ~n46215 & n46217;
  assign n46219 = ~n46214 & ~n46218;
  assign n46220 = ~n45376 & n46219;
  assign n46221 = pi423 & pi588;
  assign n46222 = n46142 & n46221;
  assign n46223 = ~n46220 & ~n46222;
  assign n46224 = ~n46213 & n46223;
  assign n46225 = n7588 & ~n46224;
  assign n46226 = ~pi647 & pi1135;
  assign n46227 = ~pi630 & ~pi1135;
  assign n46228 = ~pi1134 & ~n46227;
  assign n46229 = n45585 & n46228;
  assign n46230 = ~n46226 & n46229;
  assign n46231 = ~pi858 & ~pi1136;
  assign n46232 = pi755 & n45368;
  assign n46233 = pi725 & pi1135;
  assign n46234 = ~n46232 & ~n46233;
  assign n46235 = ~n46231 & n46234;
  assign n46236 = n45365 & n46235;
  assign n46237 = ~n46230 & ~n46236;
  assign n46238 = ~n7588 & ~n46237;
  assign po868 = n46225 | n46238;
  assign n46240 = pi701 & pi1135;
  assign n46241 = pi751 & n45368;
  assign n46242 = ~pi842 & ~pi1136;
  assign n46243 = ~n46241 & ~n46242;
  assign n46244 = n45365 & n46243;
  assign n46245 = ~n46240 & n46244;
  assign n46246 = ~pi715 & pi1135;
  assign n46247 = ~pi644 & ~pi1135;
  assign n46248 = ~pi1134 & ~n46247;
  assign n46249 = n45585 & n46248;
  assign n46250 = ~n46246 & n46249;
  assign n46251 = ~n46245 & ~n46250;
  assign n46252 = ~n7588 & ~n46251;
  assign n46253 = pi298 & n10614;
  assign n46254 = pi199 & pi1035;
  assign n46255 = pi1044 & n11221;
  assign n46256 = ~n45376 & ~n46255;
  assign n46257 = ~n46254 & n46256;
  assign n46258 = ~n46253 & n46257;
  assign n46259 = n7588 & ~n46258;
  assign n46260 = pi374 & n45388;
  assign n46261 = pi400 & n45390;
  assign n46262 = ~n46260 & ~n46261;
  assign n46263 = ~pi590 & ~n46262;
  assign n46264 = pi350 & n45386;
  assign n46265 = ~n46263 & ~n46264;
  assign n46266 = ~pi588 & ~n46265;
  assign n46267 = n45376 & ~n46266;
  assign n46268 = pi425 & n45385;
  assign n46269 = n45954 & n46268;
  assign n46270 = n46267 & ~n46269;
  assign n46271 = n46259 & ~n46270;
  assign po869 = n46252 | n46271;
  assign n46273 = pi371 & n45388;
  assign n46274 = pi396 & n45390;
  assign n46275 = ~n46273 & ~n46274;
  assign n46276 = ~pi590 & ~n46275;
  assign n46277 = pi322 & n45386;
  assign n46278 = ~n46276 & ~n46277;
  assign n46279 = n46133 & ~n46278;
  assign n46280 = pi199 & ~pi1051;
  assign n46281 = pi200 & pi1072;
  assign n46282 = ~pi200 & pi309;
  assign n46283 = ~pi199 & ~n46282;
  assign n46284 = ~n46281 & n46283;
  assign n46285 = ~n46280 & ~n46284;
  assign n46286 = ~n45376 & n46285;
  assign n46287 = pi421 & pi588;
  assign n46288 = n46142 & n46287;
  assign n46289 = ~n46286 & ~n46288;
  assign n46290 = ~n46279 & n46289;
  assign n46291 = n7588 & ~n46290;
  assign n46292 = ~pi628 & pi1135;
  assign n46293 = ~pi629 & ~pi1135;
  assign n46294 = ~pi1134 & ~n46293;
  assign n46295 = n45585 & n46294;
  assign n46296 = ~n46292 & n46295;
  assign n46297 = ~pi854 & ~pi1136;
  assign n46298 = pi756 & n45368;
  assign n46299 = pi734 & pi1135;
  assign n46300 = ~n46298 & ~n46299;
  assign n46301 = ~n46297 & n46300;
  assign n46302 = n45365 & n46301;
  assign n46303 = ~n46296 & ~n46302;
  assign n46304 = ~n7588 & ~n46303;
  assign po870 = n46291 | n46304;
  assign n46306 = pi461 & n45945;
  assign n46307 = pi439 & n45404;
  assign n46308 = ~n46306 & ~n46307;
  assign n46309 = ~pi591 & ~n46308;
  assign n46310 = pi326 & n45950;
  assign n46311 = ~n46309 & ~n46310;
  assign n46312 = ~pi588 & ~n46311;
  assign n46313 = pi449 & n45385;
  assign n46314 = n45954 & n46313;
  assign n46315 = ~n46312 & ~n46314;
  assign n46316 = n45376 & ~n46315;
  assign n46317 = pi199 & ~pi1057;
  assign n46318 = ~n45376 & ~n46317;
  assign n46319 = ~n41167 & n46318;
  assign n46320 = ~n46316 & ~n46319;
  assign n46321 = n7588 & ~n46320;
  assign n46322 = pi867 & n45431;
  assign n46323 = pi697 & pi1135;
  assign n46324 = pi762 & ~pi1135;
  assign n46325 = pi1136 & ~n46324;
  assign n46326 = ~n46323 & n46325;
  assign n46327 = ~n46322 & ~n46326;
  assign n46328 = n45364 & ~n46327;
  assign n46329 = pi693 & pi1135;
  assign n46330 = ~pi653 & ~pi1135;
  assign n46331 = pi1136 & ~n46330;
  assign n46332 = ~n46329 & n46331;
  assign n46333 = pi816 & n45351;
  assign n46334 = n45431 & n46333;
  assign n46335 = ~n46332 & ~n46334;
  assign n46336 = n45972 & ~n46335;
  assign n46337 = ~n46328 & ~n46336;
  assign n46338 = ~n7588 & ~n46337;
  assign po871 = n46321 | n46338;
  assign n46340 = ~pi1123 & po954;
  assign n46341 = ~pi715 & ~po954;
  assign n46342 = ~pi962 & ~n46341;
  assign po872 = ~n46340 & n46342;
  assign n46344 = pi440 & n46162;
  assign n46345 = pi329 & n45390;
  assign n46346 = n45376 & n46345;
  assign n46347 = ~n46344 & ~n46346;
  assign n46348 = ~pi590 & ~n46347;
  assign n46349 = pi349 & n45376;
  assign n46350 = n45386 & n46349;
  assign n46351 = ~n46348 & ~n46350;
  assign n46352 = ~pi588 & ~n46351;
  assign n46353 = pi199 & ~pi1043;
  assign n46354 = pi200 & pi1053;
  assign n46355 = ~pi200 & pi307;
  assign n46356 = ~pi199 & ~n46355;
  assign n46357 = ~n46354 & n46356;
  assign n46358 = ~n45376 & ~n46357;
  assign n46359 = ~n46353 & n46358;
  assign n46360 = pi454 & n46179;
  assign n46361 = n45954 & n46360;
  assign n46362 = n7588 & ~n46361;
  assign n46363 = ~n46359 & n46362;
  assign n46364 = ~n46352 & n46363;
  assign n46365 = pi738 & pi1135;
  assign n46366 = pi761 & n45368;
  assign n46367 = ~pi845 & ~pi1136;
  assign n46368 = ~n46366 & ~n46367;
  assign n46369 = ~n46365 & n46368;
  assign n46370 = n45365 & n46369;
  assign n46371 = ~pi626 & ~pi1135;
  assign n46372 = ~pi1134 & ~n46371;
  assign n46373 = ~pi641 & pi1135;
  assign n46374 = n45585 & ~n46373;
  assign n46375 = n46372 & n46374;
  assign n46376 = ~n7588 & ~n46375;
  assign n46377 = ~n46370 & n46376;
  assign po873 = ~n46364 & ~n46377;
  assign n46379 = pi377 & n45388;
  assign n46380 = pi318 & n45390;
  assign n46381 = ~n46379 & ~n46380;
  assign n46382 = ~pi590 & ~n46381;
  assign n46383 = pi462 & n45386;
  assign n46384 = ~n46382 & ~n46383;
  assign n46385 = n46133 & ~n46384;
  assign n46386 = ~pi199 & n41664;
  assign n46387 = pi199 & ~pi1074;
  assign n46388 = ~n45376 & ~n46387;
  assign n46389 = ~n46386 & n46388;
  assign n46390 = pi448 & pi588;
  assign n46391 = n46142 & n46390;
  assign n46392 = ~n46389 & ~n46391;
  assign n46393 = ~n46385 & n46392;
  assign n46394 = n7588 & ~n46393;
  assign n46395 = pi800 & n45431;
  assign n46396 = pi669 & pi1135;
  assign n46397 = ~pi645 & ~pi1135;
  assign n46398 = pi1136 & ~n46397;
  assign n46399 = ~n46396 & n46398;
  assign n46400 = ~n46395 & ~n46399;
  assign n46401 = n45352 & ~n46400;
  assign n46402 = ~pi705 & pi1135;
  assign n46403 = pi768 & n45368;
  assign n46404 = ~pi839 & ~pi1136;
  assign n46405 = ~n46403 & ~n46404;
  assign n46406 = n45365 & n46405;
  assign n46407 = ~n46402 & n46406;
  assign n46408 = ~n46401 & ~n46407;
  assign n46409 = ~n7588 & ~n46408;
  assign po874 = n46394 | n46409;
  assign n46411 = pi369 & n46162;
  assign n46412 = pi394 & n45390;
  assign n46413 = n45376 & n46412;
  assign n46414 = ~n46411 & ~n46413;
  assign n46415 = ~pi590 & ~n46414;
  assign n46416 = pi315 & n45376;
  assign n46417 = n45386 & n46416;
  assign n46418 = ~n46415 & ~n46417;
  assign n46419 = ~pi588 & ~n46418;
  assign n46420 = pi199 & ~pi1080;
  assign n46421 = pi200 & pi1049;
  assign n46422 = ~pi200 & pi303;
  assign n46423 = ~pi199 & ~n46422;
  assign n46424 = ~n46421 & n46423;
  assign n46425 = ~n45376 & ~n46424;
  assign n46426 = ~n46420 & n46425;
  assign n46427 = pi419 & n46179;
  assign n46428 = n45954 & n46427;
  assign n46429 = n7588 & ~n46428;
  assign n46430 = ~n46426 & n46429;
  assign n46431 = ~n46419 & n46430;
  assign n46432 = pi698 & pi1135;
  assign n46433 = pi767 & n45368;
  assign n46434 = ~pi853 & ~pi1136;
  assign n46435 = ~n46433 & ~n46434;
  assign n46436 = ~n46432 & n46435;
  assign n46437 = n45365 & n46436;
  assign n46438 = ~pi608 & ~pi1135;
  assign n46439 = ~pi1134 & ~n46438;
  assign n46440 = ~pi625 & pi1135;
  assign n46441 = n45585 & ~n46440;
  assign n46442 = n46439 & n46441;
  assign n46443 = ~n7588 & ~n46442;
  assign n46444 = ~n46437 & n46443;
  assign po875 = ~n46431 & ~n46444;
  assign n46446 = pi378 & n45388;
  assign n46447 = pi325 & n45390;
  assign n46448 = ~n46446 & ~n46447;
  assign n46449 = ~pi590 & ~n46448;
  assign n46450 = pi353 & n45386;
  assign n46451 = ~n46449 & ~n46450;
  assign n46452 = n46133 & ~n46451;
  assign n46453 = ~pi199 & n41676;
  assign n46454 = pi199 & ~pi1063;
  assign n46455 = ~n45376 & ~n46454;
  assign n46456 = ~n46453 & n46455;
  assign n46457 = pi451 & pi588;
  assign n46458 = n46142 & n46457;
  assign n46459 = ~n46456 & ~n46458;
  assign n46460 = ~n46452 & n46459;
  assign n46461 = n7588 & ~n46460;
  assign n46462 = pi807 & n45431;
  assign n46463 = pi650 & pi1135;
  assign n46464 = ~pi636 & ~pi1135;
  assign n46465 = pi1136 & ~n46464;
  assign n46466 = ~n46463 & n46465;
  assign n46467 = ~n46462 & ~n46466;
  assign n46468 = n45352 & ~n46467;
  assign n46469 = ~pi687 & pi1135;
  assign n46470 = pi774 & n45368;
  assign n46471 = ~pi868 & ~pi1136;
  assign n46472 = ~n46470 & ~n46471;
  assign n46473 = n45365 & n46472;
  assign n46474 = ~n46469 & n46473;
  assign n46475 = ~n46468 & ~n46474;
  assign n46476 = ~n7588 & ~n46475;
  assign po876 = n46461 | n46476;
  assign n46478 = pi356 & n45945;
  assign n46479 = pi381 & n45404;
  assign n46480 = ~n46478 & ~n46479;
  assign n46481 = ~pi591 & ~n46480;
  assign n46482 = pi405 & n45950;
  assign n46483 = ~n46481 & ~n46482;
  assign n46484 = ~pi588 & ~n46483;
  assign n46485 = pi445 & n45385;
  assign n46486 = n45954 & n46485;
  assign n46487 = ~n46484 & ~n46486;
  assign n46488 = n45376 & ~n46487;
  assign n46489 = pi199 & ~pi1081;
  assign n46490 = ~n45376 & ~n46489;
  assign n46491 = ~n41696 & n46490;
  assign n46492 = ~n46488 & ~n46491;
  assign n46493 = n7588 & ~n46492;
  assign n46494 = pi880 & n45431;
  assign n46495 = pi684 & pi1135;
  assign n46496 = pi750 & ~pi1135;
  assign n46497 = pi1136 & ~n46496;
  assign n46498 = ~n46495 & n46497;
  assign n46499 = ~n46494 & ~n46498;
  assign n46500 = n45364 & ~n46499;
  assign n46501 = pi654 & pi1135;
  assign n46502 = ~pi651 & ~pi1135;
  assign n46503 = pi1136 & ~n46502;
  assign n46504 = ~n46501 & n46503;
  assign n46505 = pi794 & n45351;
  assign n46506 = n45431 & n46505;
  assign n46507 = ~n46504 & ~n46506;
  assign n46508 = n45972 & ~n46507;
  assign n46509 = ~n46500 & ~n46508;
  assign n46510 = ~n7588 & ~n46509;
  assign po877 = n46493 | n46510;
  assign n46512 = pi721 & ~pi775;
  assign n46513 = pi721 & pi813;
  assign n46514 = ~pi773 & ~pi801;
  assign n46515 = pi773 & pi801;
  assign n46516 = ~n46514 & ~n46515;
  assign n46517 = ~pi771 & ~pi800;
  assign n46518 = pi771 & pi800;
  assign n46519 = ~n46517 & ~n46518;
  assign n46520 = ~pi765 & ~pi798;
  assign n46521 = pi765 & pi798;
  assign n46522 = ~n46520 & ~n46521;
  assign n46523 = pi807 & ~n46522;
  assign n46524 = pi747 & n46523;
  assign n46525 = ~pi747 & ~pi807;
  assign n46526 = ~n46522 & n46525;
  assign n46527 = ~n46524 & ~n46526;
  assign n46528 = ~pi769 & ~pi794;
  assign n46529 = pi769 & pi794;
  assign n46530 = ~n46528 & ~n46529;
  assign n46531 = ~n46527 & ~n46530;
  assign n46532 = ~n46519 & n46531;
  assign n46533 = ~n46516 & n46532;
  assign n46534 = n46513 & n46533;
  assign n46535 = ~pi816 & n46534;
  assign n46536 = n46512 & ~n46535;
  assign n46537 = ~pi945 & pi988;
  assign n46538 = pi731 & n46537;
  assign n46539 = pi747 & pi773;
  assign n46540 = pi769 & n46539;
  assign n46541 = ~pi721 & ~n46540;
  assign n46542 = pi721 & n46540;
  assign n46543 = ~n46541 & ~n46542;
  assign n46544 = pi775 & n46543;
  assign n46545 = ~n46512 & ~n46544;
  assign n46546 = ~n46519 & n46523;
  assign n46547 = ~pi721 & ~pi813;
  assign n46548 = pi794 & n46547;
  assign n46549 = pi801 & n46548;
  assign n46550 = n46546 & n46549;
  assign n46551 = ~n46534 & ~n46550;
  assign n46552 = pi816 & ~n46551;
  assign n46553 = n46544 & ~n46552;
  assign n46554 = pi795 & ~n46553;
  assign n46555 = ~n46545 & ~n46554;
  assign n46556 = n46538 & n46555;
  assign n46557 = ~pi731 & ~pi795;
  assign n46558 = pi731 & pi795;
  assign n46559 = ~n46557 & ~n46558;
  assign n46560 = ~pi775 & ~pi816;
  assign n46561 = pi775 & pi816;
  assign n46562 = ~n46560 & ~n46561;
  assign n46563 = ~n46513 & ~n46547;
  assign n46564 = ~n46562 & ~n46563;
  assign n46565 = ~n46559 & n46564;
  assign po978 = n46533 & n46565;
  assign n46567 = ~n46538 & ~po978;
  assign n46568 = pi721 & n46567;
  assign n46569 = ~n46556 & ~n46568;
  assign po878 = n46536 | ~n46569;
  assign n46571 = pi379 & n45388;
  assign n46572 = pi403 & n45390;
  assign n46573 = ~n46571 & ~n46572;
  assign n46574 = ~pi590 & ~n46573;
  assign n46575 = pi354 & n45386;
  assign n46576 = ~n46574 & ~n46575;
  assign n46577 = n46133 & ~n46576;
  assign n46578 = ~pi199 & n41682;
  assign n46579 = pi199 & ~pi1045;
  assign n46580 = ~n45376 & ~n46579;
  assign n46581 = ~n46578 & n46580;
  assign n46582 = pi428 & pi588;
  assign n46583 = n46142 & n46582;
  assign n46584 = ~n46581 & ~n46583;
  assign n46585 = ~n46577 & n46584;
  assign n46586 = n7588 & ~n46585;
  assign n46587 = ~pi851 & pi1134;
  assign n46588 = ~pi795 & ~pi1134;
  assign n46589 = ~pi1136 & ~n46588;
  assign n46590 = ~n46587 & n46589;
  assign n46591 = pi776 & pi1134;
  assign n46592 = ~pi640 & ~pi1134;
  assign n46593 = pi1136 & ~n46592;
  assign n46594 = ~n46591 & n46593;
  assign n46595 = ~n46590 & ~n46594;
  assign n46596 = ~pi1135 & ~n46595;
  assign n46597 = pi732 & ~pi1134;
  assign n46598 = pi694 & pi1134;
  assign n46599 = pi1135 & ~n46598;
  assign n46600 = pi1136 & n46599;
  assign n46601 = ~n46597 & n46600;
  assign n46602 = ~n46596 & ~n46601;
  assign n46603 = n45420 & ~n46602;
  assign po879 = n46586 | n46603;
  assign n46605 = pi723 & ~po980;
  assign n46606 = ~pi1111 & po980;
  assign n46607 = ~pi962 & ~n46606;
  assign po880 = ~n46605 & n46607;
  assign n46609 = pi724 & ~po980;
  assign n46610 = ~pi1114 & po980;
  assign n46611 = ~pi962 & ~n46610;
  assign po881 = ~n46609 & n46611;
  assign n46613 = pi725 & ~po980;
  assign n46614 = ~pi1120 & po980;
  assign n46615 = ~pi962 & ~n46614;
  assign po882 = ~n46613 & n46615;
  assign n46617 = ~pi1126 & po980;
  assign n46618 = ~pi726 & ~po980;
  assign n46619 = ~pi962 & ~n46618;
  assign po883 = ~n46617 & n46619;
  assign n46621 = ~pi1102 & po980;
  assign n46622 = ~pi727 & ~po980;
  assign n46623 = ~pi962 & ~n46622;
  assign po884 = ~n46621 & n46623;
  assign n46625 = pi728 & ~po980;
  assign n46626 = ~pi1131 & po980;
  assign n46627 = ~pi962 & ~n46626;
  assign po885 = ~n46625 & n46627;
  assign n46629 = ~pi1104 & po980;
  assign n46630 = ~pi729 & ~po980;
  assign n46631 = ~pi962 & ~n46630;
  assign po886 = ~n46629 & n46631;
  assign n46633 = ~pi1106 & po980;
  assign n46634 = ~pi730 & ~po980;
  assign n46635 = ~pi962 & ~n46634;
  assign po887 = ~n46633 & n46635;
  assign n46637 = n46533 & ~n46563;
  assign n46638 = ~n46562 & n46637;
  assign n46639 = pi795 & n46638;
  assign n46640 = ~n46539 & ~n46639;
  assign n46641 = n46538 & ~n46640;
  assign n46642 = ~n46537 & n46639;
  assign n46643 = pi731 & ~n46642;
  assign n46644 = ~n46530 & n46564;
  assign n46645 = ~pi795 & n46644;
  assign n46646 = pi801 & n46645;
  assign n46647 = n46546 & n46646;
  assign n46648 = n46539 & ~n46647;
  assign n46649 = n46537 & n46648;
  assign n46650 = ~n46643 & ~n46649;
  assign po888 = ~n46641 & ~n46650;
  assign n46652 = pi732 & ~po954;
  assign n46653 = ~pi1128 & po954;
  assign n46654 = ~pi962 & ~n46653;
  assign po889 = ~n46652 & n46654;
  assign n46656 = pi375 & n46162;
  assign n46657 = pi399 & n45390;
  assign n46658 = n45376 & n46657;
  assign n46659 = ~n46656 & ~n46658;
  assign n46660 = ~pi590 & ~n46659;
  assign n46661 = pi316 & n45376;
  assign n46662 = n45386 & n46661;
  assign n46663 = ~n46660 & ~n46662;
  assign n46664 = ~pi588 & ~n46663;
  assign n46665 = pi199 & ~pi1047;
  assign n46666 = pi200 & pi1037;
  assign n46667 = ~pi200 & pi308;
  assign n46668 = ~pi199 & ~n46667;
  assign n46669 = ~n46666 & n46668;
  assign n46670 = ~n45376 & ~n46669;
  assign n46671 = ~n46665 & n46670;
  assign n46672 = pi424 & n46179;
  assign n46673 = n45954 & n46672;
  assign n46674 = n7588 & ~n46673;
  assign n46675 = ~n46671 & n46674;
  assign n46676 = ~n46664 & n46675;
  assign n46677 = ~pi619 & ~pi1135;
  assign n46678 = ~pi1134 & ~n46677;
  assign n46679 = ~pi648 & pi1135;
  assign n46680 = n45585 & ~n46679;
  assign n46681 = n46678 & n46680;
  assign n46682 = ~pi838 & ~pi1136;
  assign n46683 = pi737 & pi1135;
  assign n46684 = ~n46682 & ~n46683;
  assign n46685 = pi777 & n45368;
  assign n46686 = n45365 & ~n46685;
  assign n46687 = n46684 & n46686;
  assign n46688 = ~n7588 & ~n46687;
  assign n46689 = ~n46681 & n46688;
  assign po890 = ~n46676 & ~n46689;
  assign n46691 = pi734 & ~po980;
  assign n46692 = ~pi1119 & po980;
  assign n46693 = ~pi962 & ~n46692;
  assign po891 = ~n46691 & n46693;
  assign n46695 = ~pi1109 & po980;
  assign n46696 = ~pi735 & ~po980;
  assign n46697 = ~pi962 & ~n46696;
  assign po892 = ~n46695 & n46697;
  assign n46699 = ~pi1101 & po980;
  assign n46700 = ~pi736 & ~po980;
  assign n46701 = ~pi962 & ~n46700;
  assign po893 = ~n46699 & n46701;
  assign n46703 = pi737 & ~po980;
  assign n46704 = ~pi1122 & po980;
  assign n46705 = ~pi962 & ~n46704;
  assign po894 = ~n46703 & n46705;
  assign n46707 = pi738 & ~po980;
  assign n46708 = ~pi1121 & po980;
  assign n46709 = ~pi962 & ~n46708;
  assign po895 = ~n46707 & n46709;
  assign n46711 = ~pi952 & n45078;
  assign po988 = n45080 & n46711;
  assign n46713 = pi739 & ~po988;
  assign n46714 = pi1108 & po988;
  assign n46715 = ~pi966 & ~n46714;
  assign po896 = n46713 | ~n46715;
  assign n46717 = pi1114 & po988;
  assign n46718 = ~pi741 & ~po988;
  assign n46719 = ~pi966 & ~n46718;
  assign po898 = n46717 | ~n46719;
  assign n46721 = pi1112 & po988;
  assign n46722 = ~pi742 & ~po988;
  assign n46723 = ~pi966 & ~n46722;
  assign po899 = n46721 | ~n46723;
  assign n46725 = pi743 & ~po988;
  assign n46726 = pi1109 & po988;
  assign n46727 = ~pi966 & ~n46726;
  assign po900 = n46725 | ~n46727;
  assign n46729 = pi1131 & po988;
  assign n46730 = ~pi744 & ~po988;
  assign n46731 = ~pi966 & ~n46730;
  assign po901 = n46729 | ~n46731;
  assign n46733 = pi1111 & po988;
  assign n46734 = ~pi745 & ~po988;
  assign n46735 = ~pi966 & ~n46734;
  assign po902 = n46733 | ~n46735;
  assign n46737 = pi746 & ~po988;
  assign n46738 = pi1104 & po988;
  assign n46739 = ~pi966 & ~n46738;
  assign po903 = n46737 | ~n46739;
  assign n46741 = pi773 & n46537;
  assign n46742 = ~pi747 & ~n46741;
  assign n46743 = n46537 & n46539;
  assign n46744 = ~n46742 & ~n46743;
  assign n46745 = pi801 & n46526;
  assign n46746 = ~n46516 & ~n46741;
  assign n46747 = n46523 & n46746;
  assign n46748 = ~n46745 & ~n46747;
  assign n46749 = n46565 & ~n46748;
  assign n46750 = ~n46519 & n46749;
  assign n46751 = ~n46530 & n46750;
  assign po904 = n46744 & ~n46751;
  assign n46753 = pi748 & ~po988;
  assign n46754 = pi1106 & po988;
  assign n46755 = ~pi966 & ~n46754;
  assign po905 = n46753 | ~n46755;
  assign n46757 = pi749 & ~po988;
  assign n46758 = pi1105 & po988;
  assign n46759 = ~pi966 & ~n46758;
  assign po906 = n46757 | ~n46759;
  assign n46761 = pi1130 & po988;
  assign n46762 = ~pi750 & ~po988;
  assign n46763 = ~pi966 & ~n46762;
  assign po907 = n46761 | ~n46763;
  assign n46765 = pi1123 & po988;
  assign n46766 = ~pi751 & ~po988;
  assign n46767 = ~pi966 & ~n46766;
  assign po908 = n46765 | ~n46767;
  assign n46769 = pi1124 & po988;
  assign n46770 = ~pi752 & ~po988;
  assign n46771 = ~pi966 & ~n46770;
  assign po909 = n46769 | ~n46771;
  assign n46773 = pi1117 & po988;
  assign n46774 = ~pi753 & ~po988;
  assign n46775 = ~pi966 & ~n46774;
  assign po910 = n46773 | ~n46775;
  assign n46777 = pi1118 & po988;
  assign n46778 = ~pi754 & ~po988;
  assign n46779 = ~pi966 & ~n46778;
  assign po911 = n46777 | ~n46779;
  assign n46781 = pi1120 & po988;
  assign n46782 = ~pi755 & ~po988;
  assign n46783 = ~pi966 & ~n46782;
  assign po912 = n46781 | ~n46783;
  assign n46785 = pi1119 & po988;
  assign n46786 = ~pi756 & ~po988;
  assign n46787 = ~pi966 & ~n46786;
  assign po913 = n46785 | ~n46787;
  assign n46789 = pi1113 & po988;
  assign n46790 = ~pi757 & ~po988;
  assign n46791 = ~pi966 & ~n46790;
  assign po914 = n46789 | ~n46791;
  assign n46793 = pi758 & ~po988;
  assign n46794 = pi1101 & po988;
  assign n46795 = ~pi966 & ~n46794;
  assign po915 = n46793 | ~n46795;
  assign n46797 = pi1100 & po988;
  assign n46798 = pi759 & ~po988;
  assign n46799 = ~pi966 & ~n46798;
  assign po916 = n46797 | ~n46799;
  assign n46801 = pi1115 & po988;
  assign n46802 = ~pi760 & ~po988;
  assign n46803 = ~pi966 & ~n46802;
  assign po917 = n46801 | ~n46803;
  assign n46805 = pi1121 & po988;
  assign n46806 = ~pi761 & ~po988;
  assign n46807 = ~pi966 & ~n46806;
  assign po918 = n46805 | ~n46807;
  assign n46809 = pi1129 & po988;
  assign n46810 = ~pi762 & ~po988;
  assign n46811 = ~pi966 & ~n46810;
  assign po919 = n46809 | ~n46811;
  assign n46813 = pi763 & ~po988;
  assign n46814 = pi1103 & po988;
  assign n46815 = ~pi966 & ~n46814;
  assign po920 = n46813 | ~n46815;
  assign n46817 = pi764 & ~po988;
  assign n46818 = pi1107 & po988;
  assign n46819 = ~pi966 & ~n46818;
  assign po921 = n46817 | ~n46819;
  assign n46821 = pi765 & ~pi945;
  assign n46822 = pi765 & ~po978;
  assign n46823 = ~pi765 & ~n46529;
  assign n46824 = ~n46518 & n46823;
  assign n46825 = ~pi773 & n46824;
  assign n46826 = ~n46524 & n46825;
  assign n46827 = n46533 & ~n46826;
  assign n46828 = ~pi721 & ~n46827;
  assign n46829 = ~pi775 & n46828;
  assign n46830 = n46557 & ~n46829;
  assign n46831 = ~n46558 & ~n46830;
  assign po963 = n46638 & ~n46831;
  assign n46833 = pi765 & n46557;
  assign n46834 = ~pi945 & ~n46833;
  assign n46835 = ~po963 & n46834;
  assign n46836 = ~n46822 & ~n46835;
  assign po922 = ~n46821 & ~n46836;
  assign n46838 = pi766 & ~po988;
  assign n46839 = pi1110 & po988;
  assign n46840 = ~pi966 & ~n46839;
  assign po923 = n46838 | ~n46840;
  assign n46842 = pi1116 & po988;
  assign n46843 = ~pi767 & ~po988;
  assign n46844 = ~pi966 & ~n46843;
  assign po924 = n46842 | ~n46844;
  assign n46846 = pi1125 & po988;
  assign n46847 = ~pi768 & ~po988;
  assign n46848 = ~pi966 & ~n46847;
  assign po925 = n46846 | ~n46848;
  assign n46850 = n46561 & n46637;
  assign n46851 = pi794 & ~n46519;
  assign n46852 = ~n46527 & n46564;
  assign n46853 = ~n46516 & n46852;
  assign n46854 = n46851 & n46853;
  assign n46855 = ~pi775 & n46854;
  assign n46856 = ~n46850 & ~n46855;
  assign n46857 = pi795 & ~n46856;
  assign n46858 = n46538 & ~n46857;
  assign n46859 = pi775 & n46539;
  assign n46860 = ~pi769 & ~n46859;
  assign n46861 = pi769 & n46859;
  assign n46862 = ~n46860 & ~n46861;
  assign n46863 = n46858 & n46862;
  assign n46864 = pi769 & n46567;
  assign po926 = n46863 | n46864;
  assign n46866 = pi1126 & po988;
  assign n46867 = ~pi770 & ~po988;
  assign n46868 = ~pi966 & ~n46867;
  assign po927 = n46866 | ~n46868;
  assign n46870 = pi987 & ~po963;
  assign n46871 = ~pi945 & n46870;
  assign n46872 = pi771 & ~po978;
  assign n46873 = pi945 & n46872;
  assign po928 = n46871 | n46873;
  assign n46875 = pi772 & ~po988;
  assign n46876 = pi1102 & po988;
  assign n46877 = ~pi966 & ~n46876;
  assign po929 = n46875 | ~n46877;
  assign n46879 = pi773 & ~po978;
  assign n46880 = pi801 & ~n46563;
  assign n46881 = po963 & ~n46880;
  assign n46882 = n46537 & ~n46881;
  assign n46883 = ~n46879 & ~n46882;
  assign po930 = ~n46741 & ~n46883;
  assign n46885 = pi1127 & po988;
  assign n46886 = ~pi774 & ~po988;
  assign n46887 = ~pi966 & ~n46886;
  assign po931 = n46885 | ~n46887;
  assign n46889 = pi731 & ~pi945;
  assign n46890 = po978 & ~n46889;
  assign n46891 = pi775 & ~n46890;
  assign n46892 = pi765 & pi771;
  assign n46893 = n46539 & n46892;
  assign n46894 = pi795 & ~pi816;
  assign n46895 = n46531 & n46894;
  assign n46896 = pi800 & n46895;
  assign n46897 = n46880 & n46896;
  assign n46898 = n46889 & ~n46897;
  assign n46899 = n46893 & n46898;
  assign n46900 = ~n46891 & ~n46899;
  assign n46901 = ~n46639 & ~n46893;
  assign n46902 = pi775 & ~n46901;
  assign n46903 = n46889 & n46902;
  assign po932 = ~n46900 & ~n46903;
  assign n46905 = pi1128 & po988;
  assign n46906 = ~pi776 & ~po988;
  assign n46907 = ~pi966 & ~n46906;
  assign po933 = n46905 | ~n46907;
  assign n46909 = pi1122 & po988;
  assign n46910 = ~pi777 & ~po988;
  assign n46911 = ~pi966 & ~n46910;
  assign po934 = n46909 | ~n46911;
  assign n46913 = pi832 & pi956;
  assign n46914 = ~pi1046 & ~pi1083;
  assign n46915 = pi1085 & n46914;
  assign n46916 = n46913 & n46915;
  assign n46917 = ~pi968 & n46916;
  assign n46918 = pi778 & ~n46917;
  assign n46919 = pi1100 & n46917;
  assign po935 = n46918 | n46919;
  assign po936 = ~pi779 | n45140;
  assign po937 = ~pi780 | n45050;
  assign n46923 = pi781 & ~n46917;
  assign n46924 = pi1101 & n46917;
  assign po938 = n46923 | n46924;
  assign n46926 = ~n41171 & ~n45093;
  assign po939 = n45049 | ~n46926;
  assign n46928 = pi783 & ~n46917;
  assign n46929 = pi1109 & n46917;
  assign po940 = n46928 | n46929;
  assign n46931 = pi784 & ~n46917;
  assign n46932 = pi1110 & n46917;
  assign po941 = n46931 | n46932;
  assign n46934 = pi785 & ~n46917;
  assign n46935 = pi1102 & n46917;
  assign po942 = n46934 | n46935;
  assign n46937 = pi24 & ~pi954;
  assign n46938 = pi786 & pi954;
  assign po943 = ~n46937 & ~n46938;
  assign n46940 = pi787 & ~n46917;
  assign n46941 = pi1104 & n46917;
  assign po944 = n46940 | n46941;
  assign n46943 = pi788 & ~n46917;
  assign n46944 = pi1105 & n46917;
  assign po945 = n46943 | n46944;
  assign n46946 = pi789 & ~n46917;
  assign n46947 = pi1106 & n46917;
  assign po946 = n46946 | n46947;
  assign n46949 = pi790 & ~n46917;
  assign n46950 = pi1107 & n46917;
  assign po947 = n46949 | n46950;
  assign n46952 = pi791 & ~n46917;
  assign n46953 = pi1108 & n46917;
  assign po948 = n46952 | n46953;
  assign n46955 = pi792 & ~n46917;
  assign n46956 = pi1103 & n46917;
  assign po949 = n46955 | n46956;
  assign n46958 = pi968 & n46916;
  assign n46959 = pi794 & ~n46958;
  assign n46960 = pi1130 & n46958;
  assign po951 = n46959 | n46960;
  assign n46962 = pi795 & ~n46958;
  assign n46963 = pi1128 & n46958;
  assign po952 = n46962 | n46963;
  assign n46965 = pi266 & ~pi269;
  assign n46966 = pi278 & ~pi280;
  assign n46967 = pi279 & n46966;
  assign n46968 = n46965 & n46967;
  assign n46969 = ~pi281 & n46968;
  assign n46970 = ~pi282 & n46969;
  assign n46971 = ~pi270 & ~pi277;
  assign n46972 = n46970 & n46971;
  assign n46973 = pi264 & ~n46972;
  assign n46974 = ~pi264 & n46972;
  assign po953 = ~n46973 & ~n46974;
  assign n46976 = pi798 & ~n46958;
  assign n46977 = pi1124 & n46958;
  assign po955 = n46976 | n46977;
  assign n46979 = pi799 & ~n46958;
  assign n46980 = ~pi1107 & n46958;
  assign po956 = ~n46979 & ~n46980;
  assign n46982 = pi800 & ~n46958;
  assign n46983 = pi1125 & n46958;
  assign po957 = n46982 | n46983;
  assign n46985 = pi801 & ~n46958;
  assign n46986 = pi1126 & n46958;
  assign po958 = n46985 | n46986;
  assign n46988 = pi803 & ~n46958;
  assign n46989 = ~pi1106 & n46958;
  assign po960 = ~n46988 & ~n46989;
  assign n46991 = pi804 & ~n46958;
  assign n46992 = pi1109 & n46958;
  assign po961 = n46991 | n46992;
  assign n46994 = pi270 & ~n45331;
  assign po962 = ~n45332 & ~n46994;
  assign n46996 = pi807 & ~n46958;
  assign n46997 = pi1127 & n46958;
  assign po964 = n46996 | n46997;
  assign n46999 = pi808 & ~n46958;
  assign n47000 = pi1101 & n46958;
  assign po965 = n46999 | n47000;
  assign n47002 = pi809 & ~n46958;
  assign n47003 = ~pi1103 & n46958;
  assign po966 = ~n47002 & ~n47003;
  assign n47005 = pi810 & ~n46958;
  assign n47006 = pi1108 & n46958;
  assign po967 = n47005 | n47006;
  assign n47008 = pi811 & ~n46958;
  assign n47009 = pi1102 & n46958;
  assign po968 = n47008 | n47009;
  assign n47011 = pi812 & ~n46958;
  assign n47012 = ~pi1104 & n46958;
  assign po969 = ~n47011 & ~n47012;
  assign n47014 = pi813 & ~n46958;
  assign n47015 = pi1131 & n46958;
  assign po970 = n47014 | n47015;
  assign n47017 = pi814 & ~n46958;
  assign n47018 = ~pi1105 & n46958;
  assign po971 = ~n47017 & ~n47018;
  assign n47020 = pi815 & ~n46958;
  assign n47021 = pi1110 & n46958;
  assign po972 = n47020 | n47021;
  assign n47023 = pi816 & ~n46958;
  assign n47024 = pi1129 & n46958;
  assign po973 = n47023 | n47024;
  assign n47026 = pi269 & ~n45328;
  assign po974 = ~n45329 & ~n47026;
  assign n47028 = n7588 & n13780;
  assign po975 = n13669 | n47028;
  assign n47030 = pi265 & ~n45334;
  assign po976 = ~n45335 & ~n47030;
  assign n47032 = pi277 & ~n45332;
  assign po977 = ~n45333 & ~n47032;
  assign po979 = ~pi811 & ~pi893;
  assign n47035 = ~pi982 & ~n6211;
  assign n47036 = n7490 & n7588;
  assign n47037 = ~n47035 & ~n47036;
  assign po981 = n6120 & ~n47037;
  assign n47039 = pi1128 & ~pi1129;
  assign n47040 = ~pi1128 & pi1129;
  assign n47041 = ~n47039 & ~n47040;
  assign n47042 = pi1125 & ~pi1126;
  assign n47043 = ~pi1125 & pi1126;
  assign n47044 = ~n47042 & ~n47043;
  assign n47045 = pi1124 & ~pi1130;
  assign n47046 = ~pi1124 & pi1130;
  assign n47047 = ~n47045 & ~n47046;
  assign n47048 = n47044 & ~n47047;
  assign n47049 = ~n47044 & n47047;
  assign n47050 = ~n47048 & ~n47049;
  assign n47051 = n47041 & n47050;
  assign n47052 = ~n47041 & ~n47050;
  assign n47053 = ~n47051 & ~n47052;
  assign n47054 = pi123 & n2608;
  assign n47055 = pi825 & n47054;
  assign n47056 = pi1127 & ~n47054;
  assign n47057 = pi1131 & n47056;
  assign n47058 = pi1131 & ~n47054;
  assign n47059 = ~n47056 & ~n47058;
  assign n47060 = ~n47055 & n47059;
  assign n47061 = ~n47057 & ~n47060;
  assign n47062 = ~n47054 & ~n47061;
  assign n47063 = ~n47055 & ~n47062;
  assign n47064 = ~n47053 & ~n47063;
  assign n47065 = n47053 & n47061;
  assign po982 = ~n47064 & ~n47065;
  assign n47067 = pi1120 & ~pi1121;
  assign n47068 = ~pi1120 & pi1121;
  assign n47069 = ~n47067 & ~n47068;
  assign n47070 = pi1116 & ~pi1117;
  assign n47071 = ~pi1116 & pi1117;
  assign n47072 = ~n47070 & ~n47071;
  assign n47073 = pi1118 & ~pi1119;
  assign n47074 = ~pi1118 & pi1119;
  assign n47075 = ~n47073 & ~n47074;
  assign n47076 = n47072 & ~n47075;
  assign n47077 = ~n47072 & n47075;
  assign n47078 = ~n47076 & ~n47077;
  assign n47079 = n47069 & n47078;
  assign n47080 = ~n47069 & ~n47078;
  assign n47081 = ~n47079 & ~n47080;
  assign n47082 = pi826 & n47054;
  assign n47083 = pi1122 & ~n47054;
  assign n47084 = pi1123 & n47083;
  assign n47085 = pi1123 & ~n47054;
  assign n47086 = ~n47083 & ~n47085;
  assign n47087 = ~n47082 & n47086;
  assign n47088 = ~n47084 & ~n47087;
  assign n47089 = ~n47054 & ~n47088;
  assign n47090 = ~n47082 & ~n47089;
  assign n47091 = ~n47081 & ~n47090;
  assign n47092 = n47081 & n47088;
  assign po983 = ~n47091 & ~n47092;
  assign n47094 = pi1101 & ~pi1102;
  assign n47095 = ~pi1101 & pi1102;
  assign n47096 = ~n47094 & ~n47095;
  assign n47097 = pi1104 & ~pi1106;
  assign n47098 = ~pi1104 & pi1106;
  assign n47099 = ~n47097 & ~n47098;
  assign n47100 = pi1103 & ~pi1105;
  assign n47101 = ~pi1103 & pi1105;
  assign n47102 = ~n47100 & ~n47101;
  assign n47103 = n47099 & ~n47102;
  assign n47104 = ~n47099 & n47102;
  assign n47105 = ~n47103 & ~n47104;
  assign n47106 = n47096 & n47105;
  assign n47107 = ~n47096 & ~n47105;
  assign n47108 = ~n47106 & ~n47107;
  assign n47109 = pi827 & n47054;
  assign n47110 = pi1107 & ~n47054;
  assign n47111 = pi1100 & n47110;
  assign n47112 = pi1100 & ~n47054;
  assign n47113 = ~n47110 & ~n47112;
  assign n47114 = ~n47109 & n47113;
  assign n47115 = ~n47111 & ~n47114;
  assign n47116 = ~n47054 & ~n47115;
  assign n47117 = ~n47109 & ~n47116;
  assign n47118 = ~n47108 & ~n47117;
  assign n47119 = n47108 & n47115;
  assign po984 = ~n47118 & ~n47119;
  assign n47121 = pi1112 & ~pi1113;
  assign n47122 = ~pi1112 & pi1113;
  assign n47123 = ~n47121 & ~n47122;
  assign n47124 = pi1108 & ~pi1109;
  assign n47125 = ~pi1108 & pi1109;
  assign n47126 = ~n47124 & ~n47125;
  assign n47127 = pi1110 & ~pi1111;
  assign n47128 = ~pi1110 & pi1111;
  assign n47129 = ~n47127 & ~n47128;
  assign n47130 = n47126 & ~n47129;
  assign n47131 = ~n47126 & n47129;
  assign n47132 = ~n47130 & ~n47131;
  assign n47133 = n47123 & n47132;
  assign n47134 = ~n47123 & ~n47132;
  assign n47135 = ~n47133 & ~n47134;
  assign n47136 = pi828 & n47054;
  assign n47137 = pi1114 & ~n47054;
  assign n47138 = pi1115 & n47137;
  assign n47139 = pi1115 & ~n47054;
  assign n47140 = ~n47137 & ~n47139;
  assign n47141 = ~n47136 & n47140;
  assign n47142 = ~n47138 & ~n47141;
  assign n47143 = ~n47054 & ~n47142;
  assign n47144 = ~n47136 & ~n47143;
  assign n47145 = ~n47135 & ~n47144;
  assign n47146 = n47135 & n47142;
  assign po985 = ~n47145 & ~n47146;
  assign n47148 = n6210 & n7588;
  assign n47149 = pi951 & ~n47148;
  assign po986 = pi1092 & ~n47149;
  assign n47151 = pi281 & ~n46968;
  assign po987 = ~n46969 & ~n47151;
  assign n47153 = pi1091 & n8735;
  assign po989 = ~pi832 & n47153;
  assign n47155 = pi833 & ~n2934;
  assign po990 = n16169 | n47155;
  assign po991 = pi946 & n2934;
  assign n47158 = pi282 & ~n45330;
  assign po992 = ~n45331 & ~n47158;
  assign n47160 = ~pi955 & pi1049;
  assign n47161 = pi837 & pi955;
  assign po993 = n47160 | n47161;
  assign n47163 = ~pi955 & pi1047;
  assign n47164 = pi838 & pi955;
  assign po994 = n47163 | n47164;
  assign n47166 = ~pi955 & pi1074;
  assign n47167 = pi839 & pi955;
  assign po995 = n47166 | n47167;
  assign n47169 = pi840 & ~n2934;
  assign n47170 = pi1196 & n2934;
  assign po996 = n47169 | n47170;
  assign po997 = ~pi33 & n8834;
  assign n47173 = ~pi955 & pi1035;
  assign n47174 = pi842 & pi955;
  assign po998 = n47173 | n47174;
  assign n47176 = ~pi955 & pi1079;
  assign n47177 = pi843 & pi955;
  assign po999 = n47176 | n47177;
  assign n47179 = ~pi955 & pi1078;
  assign n47180 = pi844 & pi955;
  assign po1000 = n47179 | n47180;
  assign n47182 = ~pi955 & pi1043;
  assign n47183 = pi845 & pi955;
  assign po1001 = n47182 | n47183;
  assign n47185 = pi846 & ~n41711;
  assign n47186 = pi1134 & n41711;
  assign po1002 = n47185 | n47186;
  assign n47188 = ~pi955 & pi1055;
  assign n47189 = pi847 & pi955;
  assign po1003 = n47188 | n47189;
  assign n47191 = ~pi955 & pi1039;
  assign n47192 = pi848 & pi955;
  assign po1004 = n47191 | n47192;
  assign n47194 = pi849 & ~n2934;
  assign n47195 = pi1198 & n2934;
  assign po1005 = n47194 | n47195;
  assign n47197 = ~pi955 & pi1048;
  assign n47198 = pi850 & pi955;
  assign po1006 = n47197 | n47198;
  assign n47200 = ~pi955 & pi1045;
  assign n47201 = pi851 & pi955;
  assign po1007 = n47200 | n47201;
  assign n47203 = ~pi955 & pi1062;
  assign n47204 = pi852 & pi955;
  assign po1008 = n47203 | n47204;
  assign n47206 = ~pi955 & pi1080;
  assign n47207 = pi853 & pi955;
  assign po1009 = n47206 | n47207;
  assign n47209 = ~pi955 & pi1051;
  assign n47210 = pi854 & pi955;
  assign po1010 = n47209 | n47210;
  assign n47212 = ~pi955 & pi1065;
  assign n47213 = pi855 & pi955;
  assign po1011 = n47212 | n47213;
  assign n47215 = ~pi955 & pi1067;
  assign n47216 = pi856 & pi955;
  assign po1012 = n47215 | n47216;
  assign n47218 = ~pi955 & pi1058;
  assign n47219 = pi857 & pi955;
  assign po1013 = n47218 | n47219;
  assign n47221 = ~pi955 & pi1087;
  assign n47222 = pi858 & pi955;
  assign po1014 = n47221 | n47222;
  assign n47224 = ~pi955 & pi1070;
  assign n47225 = pi859 & pi955;
  assign po1015 = n47224 | n47225;
  assign n47227 = ~pi955 & pi1076;
  assign n47228 = pi860 & pi955;
  assign po1016 = n47227 | n47228;
  assign n47230 = pi1093 & pi1141;
  assign n47231 = pi861 & ~pi1093;
  assign n47232 = ~n47230 & ~n47231;
  assign n47233 = ~pi228 & ~n47232;
  assign n47234 = pi123 & ~pi861;
  assign n47235 = ~pi123 & ~pi1141;
  assign n47236 = pi228 & ~n47235;
  assign n47237 = ~n47234 & n47236;
  assign po1017 = n47233 | n47237;
  assign n47239 = pi862 & ~n41711;
  assign n47240 = pi1139 & n41711;
  assign po1018 = n47239 | n47240;
  assign n47242 = pi863 & ~n2934;
  assign n47243 = pi1199 & n2934;
  assign po1019 = n47242 | n47243;
  assign n47245 = pi864 & ~n2934;
  assign n47246 = pi1197 & n2934;
  assign po1020 = n47245 | n47246;
  assign n47248 = ~pi955 & pi1040;
  assign n47249 = pi865 & pi955;
  assign po1021 = n47248 | n47249;
  assign n47251 = ~pi955 & pi1053;
  assign n47252 = pi866 & pi955;
  assign po1022 = n47251 | n47252;
  assign n47254 = ~pi955 & pi1057;
  assign n47255 = pi867 & pi955;
  assign po1023 = n47254 | n47255;
  assign n47257 = ~pi955 & pi1063;
  assign n47258 = pi868 & pi955;
  assign po1024 = n47257 | n47258;
  assign n47260 = pi1093 & pi1140;
  assign n47261 = pi869 & ~pi1093;
  assign n47262 = ~n47260 & ~n47261;
  assign n47263 = ~pi228 & ~n47262;
  assign n47264 = pi123 & ~pi869;
  assign n47265 = ~pi123 & ~pi1140;
  assign n47266 = pi228 & ~n47265;
  assign n47267 = ~n47264 & n47266;
  assign po1025 = n47263 | n47267;
  assign n47269 = ~pi955 & pi1069;
  assign n47270 = pi870 & pi955;
  assign po1026 = n47269 | n47270;
  assign n47272 = ~pi955 & pi1072;
  assign n47273 = pi871 & pi955;
  assign po1027 = n47272 | n47273;
  assign n47275 = ~pi955 & pi1084;
  assign n47276 = pi872 & pi955;
  assign po1028 = n47275 | n47276;
  assign n47278 = ~pi955 & pi1044;
  assign n47279 = pi873 & pi955;
  assign po1029 = n47278 | n47279;
  assign n47281 = ~pi955 & pi1036;
  assign n47282 = pi874 & pi955;
  assign po1030 = n47281 | n47282;
  assign n47284 = pi1093 & ~pi1136;
  assign n47285 = ~pi875 & ~pi1093;
  assign n47286 = ~n47284 & ~n47285;
  assign n47287 = ~pi228 & ~n47286;
  assign n47288 = pi123 & pi875;
  assign n47289 = ~pi123 & pi1136;
  assign n47290 = pi228 & ~n47289;
  assign n47291 = ~n47288 & n47290;
  assign po1031 = ~n47287 & ~n47291;
  assign n47293 = ~pi955 & pi1037;
  assign n47294 = pi876 & pi955;
  assign po1032 = n47293 | n47294;
  assign n47296 = pi1093 & pi1138;
  assign n47297 = pi877 & ~pi1093;
  assign n47298 = ~n47296 & ~n47297;
  assign n47299 = ~pi228 & ~n47298;
  assign n47300 = pi123 & ~pi877;
  assign n47301 = ~pi123 & ~pi1138;
  assign n47302 = pi228 & ~n47301;
  assign n47303 = ~n47300 & n47302;
  assign po1033 = n47299 | n47303;
  assign n47305 = pi1093 & pi1137;
  assign n47306 = pi878 & ~pi1093;
  assign n47307 = ~n47305 & ~n47306;
  assign n47308 = ~pi228 & ~n47307;
  assign n47309 = pi123 & ~pi878;
  assign n47310 = ~pi123 & ~pi1137;
  assign n47311 = pi228 & ~n47310;
  assign n47312 = ~n47309 & n47311;
  assign po1034 = n47308 | n47312;
  assign n47314 = pi1093 & pi1135;
  assign n47315 = pi879 & ~pi1093;
  assign n47316 = ~n47314 & ~n47315;
  assign n47317 = ~pi228 & ~n47316;
  assign n47318 = pi123 & ~pi879;
  assign n47319 = ~pi123 & ~pi1135;
  assign n47320 = pi228 & ~n47319;
  assign n47321 = ~n47318 & n47320;
  assign po1035 = n47317 | n47321;
  assign n47323 = ~pi955 & pi1081;
  assign n47324 = pi880 & pi955;
  assign po1036 = n47323 | n47324;
  assign n47326 = ~pi955 & pi1059;
  assign n47327 = pi881 & pi955;
  assign po1037 = n47326 | n47327;
  assign n47329 = ~pi883 & n47054;
  assign po1039 = n47110 | n47329;
  assign n47331 = pi1124 & ~n47054;
  assign n47332 = ~pi884 & n47054;
  assign po1040 = n47331 | n47332;
  assign n47334 = pi1125 & ~n47054;
  assign n47335 = ~pi885 & n47054;
  assign po1041 = n47334 | n47335;
  assign n47337 = pi1109 & ~n47054;
  assign n47338 = ~pi886 & n47054;
  assign po1042 = n47337 | n47338;
  assign n47340 = ~pi887 & n47054;
  assign po1043 = n47112 | n47340;
  assign n47342 = pi1120 & ~n47054;
  assign n47343 = ~pi888 & n47054;
  assign po1044 = n47342 | n47343;
  assign n47345 = pi1103 & ~n47054;
  assign n47346 = ~pi889 & n47054;
  assign po1045 = n47345 | n47346;
  assign n47348 = pi1126 & ~n47054;
  assign n47349 = ~pi890 & n47054;
  assign po1046 = n47348 | n47349;
  assign n47351 = pi1116 & ~n47054;
  assign n47352 = ~pi891 & n47054;
  assign po1047 = n47351 | n47352;
  assign n47354 = pi1101 & ~n47054;
  assign n47355 = ~pi892 & n47054;
  assign po1048 = n47354 | n47355;
  assign n47357 = pi1119 & ~n47054;
  assign n47358 = ~pi894 & n47054;
  assign po1050 = n47357 | n47358;
  assign n47360 = pi1113 & ~n47054;
  assign n47361 = ~pi895 & n47054;
  assign po1051 = n47360 | n47361;
  assign n47363 = pi1118 & ~n47054;
  assign n47364 = ~pi896 & n47054;
  assign po1052 = n47363 | n47364;
  assign n47366 = pi1129 & ~n47054;
  assign n47367 = ~pi898 & n47054;
  assign po1054 = n47366 | n47367;
  assign n47369 = ~pi899 & n47054;
  assign po1055 = n47139 | n47369;
  assign n47371 = pi1110 & ~n47054;
  assign n47372 = ~pi900 & n47054;
  assign po1056 = n47371 | n47372;
  assign n47374 = pi1111 & ~n47054;
  assign n47375 = ~pi902 & n47054;
  assign po1058 = n47374 | n47375;
  assign n47377 = pi1121 & ~n47054;
  assign n47378 = ~pi903 & n47054;
  assign po1059 = n47377 | n47378;
  assign n47380 = ~pi904 & n47054;
  assign po1060 = n47056 | n47380;
  assign n47382 = ~pi905 & n47054;
  assign po1061 = n47058 | n47382;
  assign n47384 = pi1128 & ~n47054;
  assign n47385 = ~pi906 & n47054;
  assign po1062 = n47384 | n47385;
  assign n47387 = ~pi615 & pi979;
  assign n47388 = pi604 & ~pi979;
  assign n47389 = ~n47387 & ~n47388;
  assign n47390 = pi782 & n47389;
  assign n47391 = ~pi782 & ~pi907;
  assign n47392 = ~pi598 & pi979;
  assign n47393 = ~pi624 & ~pi979;
  assign n47394 = pi782 & ~n47393;
  assign n47395 = ~n47392 & n47394;
  assign n47396 = ~n47391 & ~n47395;
  assign po1063 = ~n47390 & n47396;
  assign n47398 = ~pi908 & n47054;
  assign po1064 = n47083 | n47398;
  assign n47400 = pi1105 & ~n47054;
  assign n47401 = ~pi909 & n47054;
  assign po1065 = n47400 | n47401;
  assign n47403 = pi1117 & ~n47054;
  assign n47404 = ~pi910 & n47054;
  assign po1066 = n47403 | n47404;
  assign n47406 = pi1130 & ~n47054;
  assign n47407 = ~pi911 & n47054;
  assign po1067 = n47406 | n47407;
  assign n47409 = ~pi912 & n47054;
  assign po1068 = n47137 | n47409;
  assign n47411 = pi1106 & ~n47054;
  assign n47412 = ~pi913 & n47054;
  assign po1069 = n47411 | n47412;
  assign n47414 = pi280 & ~n45327;
  assign po1070 = ~n45328 & ~n47414;
  assign n47416 = pi1108 & ~n47054;
  assign n47417 = ~pi915 & n47054;
  assign po1071 = n47416 | n47417;
  assign n47419 = ~pi916 & n47054;
  assign po1072 = n47085 | n47419;
  assign n47421 = pi1112 & ~n47054;
  assign n47422 = ~pi917 & n47054;
  assign po1073 = n47421 | n47422;
  assign n47424 = pi1104 & ~n47054;
  assign n47425 = ~pi918 & n47054;
  assign po1074 = n47424 | n47425;
  assign n47427 = pi1102 & ~n47054;
  assign n47428 = ~pi919 & n47054;
  assign po1075 = n47427 | n47428;
  assign n47430 = pi1093 & pi1139;
  assign n47431 = pi920 & ~pi1093;
  assign po1076 = n47430 | n47431;
  assign n47433 = pi921 & ~pi1093;
  assign po1077 = n47260 | n47433;
  assign n47435 = ~pi922 & ~pi1093;
  assign n47436 = pi1093 & ~pi1152;
  assign po1078 = ~n47435 & ~n47436;
  assign n47438 = ~pi923 & ~pi1093;
  assign n47439 = pi1093 & ~pi1154;
  assign po1079 = ~n47438 & ~n47439;
  assign n47441 = pi311 & ~pi312;
  assign po1080 = n43311 & n47441;
  assign n47443 = ~pi925 & ~pi1093;
  assign n47444 = pi1093 & ~pi1155;
  assign po1081 = ~n47443 & ~n47444;
  assign n47446 = ~pi926 & ~pi1093;
  assign n47447 = pi1093 & ~pi1157;
  assign po1082 = ~n47446 & ~n47447;
  assign n47449 = ~pi927 & ~pi1093;
  assign n47450 = pi1093 & ~pi1145;
  assign po1083 = ~n47449 & ~n47450;
  assign n47452 = ~pi928 & ~pi1093;
  assign po1084 = ~n47284 & ~n47452;
  assign n47454 = ~pi929 & ~pi1093;
  assign n47455 = pi1093 & ~pi1144;
  assign po1085 = ~n47454 & ~n47455;
  assign n47457 = ~pi930 & ~pi1093;
  assign n47458 = pi1093 & ~pi1134;
  assign po1086 = ~n47457 & ~n47458;
  assign n47460 = ~pi931 & ~pi1093;
  assign n47461 = pi1093 & ~pi1150;
  assign po1087 = ~n47460 & ~n47461;
  assign n47463 = pi932 & ~pi1093;
  assign po1088 = n41700 | n47463;
  assign n47465 = pi933 & ~pi1093;
  assign po1089 = n47305 | n47465;
  assign n47467 = ~pi934 & ~pi1093;
  assign n47468 = pi1093 & ~pi1147;
  assign po1090 = ~n47467 & ~n47468;
  assign n47470 = pi935 & ~pi1093;
  assign po1091 = n47230 | n47470;
  assign n47472 = ~pi936 & ~pi1093;
  assign n47473 = pi1093 & ~pi1149;
  assign po1092 = ~n47472 & ~n47473;
  assign n47475 = ~pi937 & ~pi1093;
  assign n47476 = pi1093 & ~pi1148;
  assign po1093 = ~n47475 & ~n47476;
  assign n47478 = pi938 & ~pi1093;
  assign po1094 = n47314 | n47478;
  assign n47480 = ~pi939 & ~pi1093;
  assign n47481 = pi1093 & ~pi1146;
  assign po1095 = ~n47480 & ~n47481;
  assign n47483 = pi940 & ~pi1093;
  assign po1096 = n47296 | n47483;
  assign n47485 = ~pi941 & ~pi1093;
  assign n47486 = pi1093 & ~pi1153;
  assign po1097 = ~n47485 & ~n47486;
  assign n47488 = ~pi942 & ~pi1093;
  assign n47489 = pi1093 & ~pi1156;
  assign po1098 = ~n47488 & ~n47489;
  assign n47491 = ~pi943 & ~pi1093;
  assign n47492 = pi1093 & ~pi1151;
  assign po1099 = ~n47491 & ~n47492;
  assign n47494 = pi1093 & pi1143;
  assign n47495 = pi944 & ~pi1093;
  assign po1100 = n47494 | n47495;
  assign po1102 = pi230 & n2934;
  assign n47498 = ~pi782 & pi947;
  assign po1103 = n47395 | n47498;
  assign n47500 = ~pi266 & ~pi992;
  assign po1104 = ~n45327 & ~n47500;
  assign n47502 = ~pi313 & ~pi954;
  assign n47503 = pi949 & pi954;
  assign po1105 = n47502 | n47503;
  assign po1107 = ~n7490 & n13822;
  assign n47506 = pi957 & pi1092;
  assign po1112 = pi31 | n47506;
  assign po1115 = ~pi782 & pi960;
  assign po1116 = ~pi230 & pi961;
  assign po1118 = ~pi782 & pi963;
  assign po1122 = ~pi230 & pi967;
  assign po1124 = ~pi230 & pi969;
  assign po1125 = ~pi782 & pi970;
  assign po1126 = ~pi230 & pi971;
  assign po1127 = ~pi782 & pi972;
  assign po1128 = ~pi230 & pi974;
  assign po1129 = ~pi782 & pi975;
  assign po1131 = ~pi230 & pi977;
  assign po1132 = ~pi782 & pi978;
  assign po1133 = pi598 | ~pi615;
  assign po1135 = pi824 & pi1092;
  assign po1137 = pi604 | pi624;
  assign po166 = 1'b1;
  assign po170 = ~pi1090;
  assign po1110 = ~pi954;
  assign po1130 = ~pi278;
  assign po1146 = ~pi915;
  assign po1147 = ~pi825;
  assign po1148 = ~pi826;
  assign po1149 = ~pi913;
  assign po1150 = ~pi894;
  assign po1151 = ~pi905;
  assign po1153 = ~pi890;
  assign po1155 = ~pi906;
  assign po1156 = ~pi896;
  assign po1157 = ~pi909;
  assign po1158 = ~pi911;
  assign po1159 = ~pi908;
  assign po1160 = ~pi891;
  assign po1161 = ~pi902;
  assign po1162 = ~pi903;
  assign po1163 = ~pi883;
  assign po1164 = ~pi888;
  assign po1165 = ~pi919;
  assign po1166 = ~pi886;
  assign po1167 = ~pi912;
  assign po1168 = ~pi895;
  assign po1169 = ~pi916;
  assign po1170 = ~pi889;
  assign po1171 = ~pi900;
  assign po1172 = ~pi885;
  assign po1173 = ~pi904;
  assign po1174 = ~pi899;
  assign po1175 = ~pi918;
  assign po1176 = ~pi898;
  assign po1177 = ~pi917;
  assign po1178 = ~pi827;
  assign po1179 = ~pi887;
  assign po1180 = ~pi884;
  assign po1181 = ~pi910;
  assign po1182 = ~pi828;
  assign po1183 = ~pi892;
  assign po0 = pi668;
  assign po1 = pi672;
  assign po2 = pi664;
  assign po3 = pi667;
  assign po4 = pi676;
  assign po5 = pi673;
  assign po6 = pi675;
  assign po7 = pi666;
  assign po8 = pi679;
  assign po9 = pi674;
  assign po10 = pi663;
  assign po11 = pi670;
  assign po12 = pi677;
  assign po13 = pi682;
  assign po14 = pi671;
  assign po15 = pi678;
  assign po16 = pi718;
  assign po17 = pi707;
  assign po18 = pi708;
  assign po19 = pi713;
  assign po20 = pi711;
  assign po21 = pi716;
  assign po22 = pi733;
  assign po23 = pi712;
  assign po24 = pi689;
  assign po25 = pi717;
  assign po26 = pi692;
  assign po27 = pi719;
  assign po28 = pi722;
  assign po29 = pi714;
  assign po30 = pi720;
  assign po31 = pi685;
  assign po32 = pi837;
  assign po33 = pi850;
  assign po34 = pi872;
  assign po35 = pi871;
  assign po36 = pi881;
  assign po37 = pi866;
  assign po38 = pi876;
  assign po39 = pi873;
  assign po40 = pi874;
  assign po41 = pi859;
  assign po42 = pi855;
  assign po43 = pi852;
  assign po44 = pi870;
  assign po45 = pi848;
  assign po46 = pi865;
  assign po47 = pi856;
  assign po48 = pi853;
  assign po49 = pi847;
  assign po50 = pi857;
  assign po51 = pi854;
  assign po52 = pi858;
  assign po53 = pi845;
  assign po54 = pi838;
  assign po55 = pi842;
  assign po56 = pi843;
  assign po57 = pi839;
  assign po58 = pi844;
  assign po59 = pi868;
  assign po60 = pi851;
  assign po61 = pi867;
  assign po62 = pi880;
  assign po63 = pi860;
  assign po64 = pi1030;
  assign po65 = pi1034;
  assign po66 = pi1015;
  assign po67 = pi1020;
  assign po68 = pi1025;
  assign po69 = pi1005;
  assign po70 = pi996;
  assign po71 = pi1012;
  assign po72 = pi993;
  assign po73 = pi1016;
  assign po74 = pi1021;
  assign po75 = pi1010;
  assign po76 = pi1027;
  assign po77 = pi1018;
  assign po78 = pi1017;
  assign po79 = pi1024;
  assign po80 = pi1009;
  assign po81 = pi1032;
  assign po82 = pi1003;
  assign po83 = pi997;
  assign po84 = pi1013;
  assign po85 = pi1011;
  assign po86 = pi1008;
  assign po87 = pi1019;
  assign po88 = pi1031;
  assign po89 = pi1022;
  assign po90 = pi1000;
  assign po91 = pi1023;
  assign po92 = pi1002;
  assign po93 = pi1026;
  assign po94 = pi1006;
  assign po95 = pi998;
  assign po96 = pi31;
  assign po97 = pi80;
  assign po98 = pi893;
  assign po99 = pi467;
  assign po100 = pi78;
  assign po101 = pi112;
  assign po102 = pi13;
  assign po103 = pi25;
  assign po104 = pi226;
  assign po105 = pi127;
  assign po106 = pi822;
  assign po107 = pi808;
  assign po108 = pi227;
  assign po109 = pi477;
  assign po110 = pi834;
  assign po111 = pi229;
  assign po112 = pi12;
  assign po113 = pi11;
  assign po114 = pi10;
  assign po115 = pi9;
  assign po116 = pi8;
  assign po117 = pi7;
  assign po118 = pi6;
  assign po119 = pi5;
  assign po120 = pi4;
  assign po121 = pi3;
  assign po122 = pi0;
  assign po123 = pi2;
  assign po124 = pi1;
  assign po125 = pi310;
  assign po126 = pi302;
  assign po127 = pi475;
  assign po128 = pi474;
  assign po129 = pi466;
  assign po130 = pi473;
  assign po131 = pi471;
  assign po132 = pi472;
  assign po133 = pi470;
  assign po134 = pi469;
  assign po135 = pi465;
  assign po136 = pi1028;
  assign po137 = pi1033;
  assign po138 = pi995;
  assign po139 = pi994;
  assign po140 = pi28;
  assign po141 = pi27;
  assign po142 = pi26;
  assign po143 = pi29;
  assign po144 = pi15;
  assign po145 = pi14;
  assign po146 = pi21;
  assign po147 = pi20;
  assign po148 = pi19;
  assign po149 = pi18;
  assign po150 = pi17;
  assign po151 = pi16;
  assign po152 = pi1096;
  assign po168 = pi228;
  assign po169 = pi22;
  assign po179 = pi1089;
  assign po180 = pi23;
  assign po181 = po167;
  assign po188 = pi37;
  assign po263 = pi117;
  assign po285 = pi131;
  assign po386 = pi232;
  assign po388 = pi236;
  assign po636 = pi583;
  assign po1053 = pi67;
  assign po1108 = pi1134;
  assign po1109 = pi964;
  assign po1111 = pi965;
  assign po1113 = pi991;
  assign po1114 = pi985;
  assign po1117 = pi1014;
  assign po1119 = pi1029;
  assign po1120 = pi1004;
  assign po1121 = pi1007;
  assign po1123 = pi1135;
  assign po1134 = pi1064;
  assign po1136 = pi299;
  assign po1138 = pi1075;
  assign po1139 = pi1052;
  assign po1140 = pi771;
  assign po1141 = pi765;
  assign po1142 = pi605;
  assign po1143 = pi601;
  assign po1144 = pi278;
  assign po1145 = pi279;
  assign po1152 = pi1095;
  assign po1154 = pi1094;
  assign po1184 = pi1187;
  assign po1185 = pi1172;
  assign po1186 = pi1170;
  assign po1187 = pi1138;
  assign po1188 = pi1177;
  assign po1189 = pi1178;
  assign po1190 = pi863;
  assign po1191 = pi1203;
  assign po1192 = pi1185;
  assign po1193 = pi1171;
  assign po1194 = pi1192;
  assign po1195 = pi1137;
  assign po1196 = pi1186;
  assign po1197 = pi1165;
  assign po1198 = pi1164;
  assign po1199 = pi1098;
  assign po1200 = pi1183;
  assign po1201 = pi230;
  assign po1202 = pi1169;
  assign po1203 = pi1136;
  assign po1204 = pi1181;
  assign po1205 = pi849;
  assign po1206 = pi1193;
  assign po1207 = pi1182;
  assign po1208 = pi1168;
  assign po1209 = pi1175;
  assign po1210 = pi1191;
  assign po1211 = pi1099;
  assign po1212 = pi1174;
  assign po1213 = pi1179;
  assign po1214 = pi1202;
  assign po1215 = pi1176;
  assign po1216 = pi1173;
  assign po1217 = pi1201;
  assign po1218 = pi1167;
  assign po1219 = pi840;
  assign po1220 = pi1189;
  assign po1221 = pi1195;
  assign po1222 = pi864;
  assign po1223 = pi1190;
  assign po1224 = pi1188;
  assign po1225 = pi1180;
  assign po1226 = pi1194;
  assign po1227 = pi1097;
  assign po1228 = pi1166;
  assign po1229 = pi1200;
  assign po1230 = pi1184;
endmodule
