module alu4_cl ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13,
    po0, po1, po2, po3, po4, po5, po6, po7  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13;
  output po0, po1, po2, po3, po4, po5, po6, po7;
  wire n23, n24, n25, n26, n27, n28, n29,
    n30, n31, n32, n33, n34, n35, n36, n37,
    n38, n39, n40, n41, n42, n43, n44, n45,
    n46, n47, n48, n49, n50, n51, n52, n53,
    n54, n55, n56, n57, n58, n59, n60, n61,
    n62, n63, n64, n65, n66, n67, n68, n69,
    n70, n71, n72, n73, n74, n75, n76, n77,
    n78, n79, n80, n81, n82, n83, n84, n85,
    n86, n87, n88, n89, n90, n91, n92, n93,
    n94, n95, n96, n97, n98, n99, n100,
    n101, n102, n103, n104, n105, n106, n107,
    n108, n109, n110, n111, n112, n113, n114,
    n115, n116, n117, n118, n119, n120, n121,
    n122, n123, n124, n125, n126, n127, n128,
    n129, n130, n131, n132, n133, n134, n135,
    n136, n137, n138, n139, n140, n141, n142,
    n143, n144, n145, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156,
    n157, n158, n159, n160, n161, n162, n163,
    n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177,
    n178, n179, n180, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192,
    n193, n194, n195, n196, n197, n198, n199,
    n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213,
    n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227,
    n228, n229, n230, n231, n232, n233, n234,
    n235, n236, n237, n238, n239, n240, n241,
    n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n323, n324, n325, n326,
    n327, n328, n329, n330, n331, n332, n333,
    n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403,
    n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416, n417,
    n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438,
    n439, n440, n441, n442, n443, n444, n445,
    n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n470, n472, n473, n474, n475,
    n476, n477, n478, n479, n480, n481, n482,
    n483, n484, n485, n486, n487, n488, n489,
    n490, n491, n492, n493, n494, n495, n496,
    n497, n498, n499, n500, n501, n502, n503,
    n504, n505, n506, n507, n508, n509, n510,
    n512, n513, n514, n515, n516, n517, n518,
    n519, n520, n521, n522, n523, n524, n525,
    n526, n527, n528, n529, n530, n531, n532,
    n533, n534, n535, n536, n537, n538, n539,
    n540, n541, n542, n543, n544, n545, n546,
    n547, n548, n549, n550, n551, n552, n553,
    n554, n555, n556, n557, n558, n559, n560,
    n561, n562, n563, n564, n565, n566, n567,
    n568, n569, n570, n571, n572, n573, n574,
    n575, n576, n577, n578, n579, n580, n581,
    n582, n583, n584, n585, n586, n587, n588,
    n589, n590, n591, n592, n593, n594, n595,
    n596, n597, n598, n599, n600, n601, n602,
    n603, n604, n605, n606, n607, n608, n609,
    n610, n611, n612, n613, n614, n615, n616,
    n617, n618, n619, n621, n622, n623, n624,
    n625, n626, n627, n628, n629, n630, n631,
    n632, n633, n634, n635, n636, n637, n638,
    n639, n640, n641, n642, n643, n644, n645,
    n647, n648;
  assign n23 = ~pi08 & ~pi09;
  assign n24 = ~pi10 & ~n23;
  assign n25 = pi00 & pi11;
  assign n26 = ~n24 & n25;
  assign n27 = ~pi08 & ~pi10;
  assign n28 = pi04 & n27;
  assign n29 = pi10 & ~pi11;
  assign n30 = pi08 & pi09;
  assign n31 = ~n24 & ~n30;
  assign n32 = ~n29 & n31;
  assign n33 = ~pi09 & n32;
  assign n34 = ~n28 & ~n33;
  assign n35 = ~pi00 & ~pi04;
  assign n36 = ~pi10 & ~pi11;
  assign n37 = ~pi13 & n36;
  assign n38 = pi10 & pi13;
  assign n39 = ~n37 & ~n38;
  assign n40 = pi08 & ~pi09;
  assign n41 = ~n39 & n40;
  assign n42 = ~n35 & n41;
  assign n43 = pi08 & ~pi10;
  assign n44 = ~pi08 & n29;
  assign n45 = ~n43 & ~n44;
  assign n46 = pi09 & ~n45;
  assign n47 = ~n36 & n46;
  assign n48 = pi11 & ~n24;
  assign n49 = ~n47 & ~n48;
  assign n50 = ~pi10 & pi13;
  assign n51 = ~n49 & n50;
  assign n52 = ~pi09 & ~pi11;
  assign n53 = ~pi08 & pi10;
  assign n54 = n52 & n53;
  assign n55 = ~n51 & ~n54;
  assign n56 = pi00 & pi04;
  assign n57 = ~n55 & n56;
  assign n58 = n29 & n30;
  assign n59 = pi08 & pi10;
  assign n60 = ~pi09 & pi11;
  assign n61 = ~pi13 & n60;
  assign n62 = n59 & n61;
  assign n63 = ~pi08 & pi09;
  assign n64 = pi13 & n63;
  assign n65 = ~n29 & n64;
  assign n66 = ~n58 & ~n62;
  assign n67 = ~n65 & n66;
  assign n68 = ~pi04 & ~n67;
  assign n69 = ~n37 & ~n61;
  assign n70 = ~pi10 & ~n69;
  assign n71 = ~pi08 & n70;
  assign n72 = ~pi00 & n71;
  assign n73 = ~n35 & ~n56;
  assign n74 = ~pi00 & ~n29;
  assign n75 = n64 & ~n74;
  assign n76 = n73 & n75;
  assign n77 = ~n42 & ~n76;
  assign n78 = ~n68 & n77;
  assign n79 = ~n72 & n78;
  assign n80 = ~n57 & n79;
  assign n81 = ~n34 & ~n80;
  assign n82 = n35 & n44;
  assign n83 = pi00 & ~n80;
  assign n84 = n59 & n83;
  assign n85 = ~pi08 & pi11;
  assign n86 = ~pi00 & ~n85;
  assign n87 = ~pi11 & ~n53;
  assign n88 = pi04 & ~n86;
  assign n89 = ~n87 & n88;
  assign n90 = pi09 & ~n82;
  assign n91 = ~n89 & n90;
  assign n92 = ~n84 & n91;
  assign n93 = pi08 & n29;
  assign n94 = ~n25 & ~n93;
  assign n95 = ~pi04 & ~n94;
  assign n96 = pi08 & n36;
  assign n97 = ~n53 & ~n96;
  assign n98 = n80 & ~n97;
  assign n99 = ~pi00 & pi04;
  assign n100 = pi11 & n43;
  assign n101 = n99 & n100;
  assign n102 = ~pi09 & ~n101;
  assign n103 = ~n95 & n102;
  assign n104 = ~n98 & n103;
  assign n105 = ~n92 & ~n104;
  assign n106 = ~n26 & ~n81;
  assign n107 = ~n105 & n106;
  assign n108 = ~pi13 & ~n107;
  assign n109 = ~pi09 & n43;
  assign n110 = n73 & n109;
  assign n111 = pi04 & n43;
  assign n112 = ~pi00 & n80;
  assign n113 = pi09 & pi13;
  assign n114 = n85 & n113;
  assign n115 = ~n112 & n114;
  assign n116 = pi13 & n29;
  assign n117 = n23 & n80;
  assign n118 = n30 & n83;
  assign n119 = n40 & n56;
  assign n120 = ~n117 & ~n119;
  assign n121 = ~n118 & n120;
  assign n122 = n116 & ~n121;
  assign n123 = ~n115 & ~n122;
  assign n124 = pi00 & ~pi08;
  assign n125 = n123 & n124;
  assign n126 = ~n111 & ~n125;
  assign n127 = n52 & ~n126;
  assign n128 = ~pi00 & n54;
  assign n129 = pi09 & n85;
  assign n130 = n50 & n129;
  assign n131 = n56 & n130;
  assign n132 = ~pi09 & n116;
  assign n133 = pi08 & n132;
  assign n134 = n123 & n133;
  assign n135 = ~n131 & ~n134;
  assign n136 = pi09 & n27;
  assign n137 = pi11 & n136;
  assign n138 = n135 & n137;
  assign n139 = ~n123 & ~n128;
  assign n140 = ~n138 & n139;
  assign n141 = ~n135 & n137;
  assign n142 = ~n58 & n123;
  assign n143 = ~n141 & n142;
  assign n144 = ~n140 & ~n143;
  assign n145 = ~pi00 & pi11;
  assign n146 = ~n24 & n145;
  assign n147 = n52 & n59;
  assign n148 = n135 & n147;
  assign n149 = ~n80 & ~n146;
  assign n150 = ~n148 & n149;
  assign n151 = n25 & ~n30;
  assign n152 = pi08 & n52;
  assign n153 = ~n135 & n152;
  assign n154 = ~n151 & ~n153;
  assign n155 = pi10 & ~n154;
  assign n156 = ~n47 & n80;
  assign n157 = ~n155 & n156;
  assign n158 = ~n150 & ~n157;
  assign n159 = pi10 & n30;
  assign n160 = n145 & n159;
  assign n161 = pi09 & ~n80;
  assign n162 = ~pi00 & ~n161;
  assign n163 = ~pi09 & n80;
  assign n164 = pi11 & ~n163;
  assign n165 = n27 & ~n162;
  assign n166 = ~n164 & n165;
  assign n167 = ~n110 & ~n160;
  assign n168 = ~n166 & n167;
  assign n169 = ~n127 & n168;
  assign n170 = ~n144 & n169;
  assign n171 = ~n158 & n170;
  assign n172 = pi13 & ~n171;
  assign n173 = pi12 & ~n172;
  assign n174 = ~pi12 & n172;
  assign n175 = pi13 & ~n174;
  assign n176 = ~n173 & n175;
  assign n177 = n53 & n61;
  assign n178 = n96 & n113;
  assign n179 = ~n177 & ~n178;
  assign n180 = ~n108 & n179;
  assign po0 = n176 | ~n180;
  assign n182 = ~pi08 & pi13;
  assign n183 = ~pi09 & pi10;
  assign n184 = n25 & n183;
  assign n185 = ~pi01 & ~pi05;
  assign n186 = n99 & n185;
  assign n187 = ~pi01 & ~n29;
  assign n188 = pi01 & pi05;
  assign n189 = ~n185 & ~n188;
  assign n190 = ~n99 & ~n187;
  assign n191 = n189 & n190;
  assign n192 = ~n186 & ~n191;
  assign n193 = pi09 & ~n192;
  assign n194 = ~n184 & ~n193;
  assign n195 = n182 & ~n194;
  assign n196 = n41 & ~n185;
  assign n197 = ~pi05 & ~n67;
  assign n198 = ~pi01 & n71;
  assign n199 = n55 & ~n132;
  assign n200 = n75 & n99;
  assign n201 = n199 & ~n200;
  assign n202 = n188 & ~n201;
  assign n203 = ~n196 & ~n197;
  assign n204 = ~n198 & n203;
  assign n205 = ~n195 & n204;
  assign n206 = ~n202 & n205;
  assign n207 = n83 & ~n206;
  assign n208 = ~n83 & n206;
  assign n209 = ~n207 & ~n208;
  assign n210 = pi11 & n31;
  assign n211 = n209 & n210;
  assign n212 = ~pi01 & n206;
  assign n213 = n114 & ~n212;
  assign n214 = pi09 & n206;
  assign n215 = ~pi05 & ~pi09;
  assign n216 = pi01 & pi08;
  assign n217 = ~n215 & n216;
  assign n218 = ~pi08 & n206;
  assign n219 = ~n217 & ~n218;
  assign n220 = n116 & ~n214;
  assign n221 = ~n219 & n220;
  assign n222 = ~n213 & ~n221;
  assign n223 = pi00 & ~n123;
  assign n224 = n222 & ~n223;
  assign n225 = ~n123 & ~n222;
  assign n226 = pi00 & n225;
  assign n227 = ~n224 & ~n226;
  assign n228 = n54 & n227;
  assign n229 = ~n211 & ~n228;
  assign n230 = ~pi01 & ~n229;
  assign n231 = n123 & n222;
  assign n232 = ~n225 & ~n231;
  assign n233 = n159 & ~n232;
  assign n234 = n136 & ~n206;
  assign n235 = ~n233 & ~n234;
  assign n236 = ~pi11 & ~n235;
  assign n237 = ~pi05 & ~n56;
  assign n238 = n109 & n237;
  assign n239 = n32 & ~n209;
  assign n240 = n25 & n159;
  assign n241 = ~n30 & n36;
  assign n242 = ~n238 & ~n241;
  assign n243 = ~n240 & n242;
  assign n244 = ~n239 & n243;
  assign n245 = pi01 & ~n244;
  assign n246 = ~pi11 & n136;
  assign n247 = ~n47 & ~n246;
  assign n248 = ~n80 & ~n247;
  assign n249 = ~n206 & n248;
  assign n250 = n80 & n206;
  assign n251 = n47 & n250;
  assign n252 = ~pi00 & ~pi01;
  assign n253 = n159 & n252;
  assign n254 = n56 & n185;
  assign n255 = n109 & n254;
  assign n256 = ~n253 & ~n255;
  assign n257 = pi11 & ~n256;
  assign n258 = ~pi01 & pi05;
  assign n259 = ~n56 & ~n258;
  assign n260 = n56 & ~n188;
  assign n261 = n109 & ~n259;
  assign n262 = ~n260 & n261;
  assign n263 = pi05 & n43;
  assign n264 = ~n80 & ~n135;
  assign n265 = n130 & n188;
  assign n266 = n133 & n222;
  assign n267 = ~n265 & ~n266;
  assign n268 = n264 & ~n267;
  assign n269 = ~n264 & n267;
  assign n270 = ~n268 & ~n269;
  assign n271 = ~n206 & ~n270;
  assign n272 = n206 & n270;
  assign n273 = ~n271 & ~n272;
  assign n274 = n59 & ~n273;
  assign n275 = pi01 & ~pi08;
  assign n276 = ~n227 & n275;
  assign n277 = ~n263 & ~n276;
  assign n278 = ~n274 & n277;
  assign n279 = n52 & ~n278;
  assign n280 = n131 & ~n267;
  assign n281 = ~n131 & n267;
  assign n282 = ~n280 & ~n281;
  assign n283 = ~n222 & ~n282;
  assign n284 = n222 & n282;
  assign n285 = ~n283 & ~n284;
  assign n286 = n137 & ~n285;
  assign n287 = ~n257 & ~n262;
  assign n288 = ~n249 & n287;
  assign n289 = ~n251 & n288;
  assign n290 = ~n245 & n289;
  assign n291 = ~n236 & n290;
  assign n292 = ~n230 & n291;
  assign n293 = ~n286 & n292;
  assign n294 = ~n279 & n293;
  assign n295 = n175 & ~n294;
  assign n296 = n174 & n294;
  assign n297 = pi01 & n48;
  assign n298 = n100 & n258;
  assign n299 = ~n97 & n206;
  assign n300 = pi01 & pi11;
  assign n301 = ~n93 & ~n300;
  assign n302 = ~pi05 & ~n301;
  assign n303 = ~n298 & ~n302;
  assign n304 = ~n299 & n303;
  assign n305 = ~pi09 & ~n304;
  assign n306 = pi05 & n85;
  assign n307 = ~n44 & ~n300;
  assign n308 = ~n189 & ~n307;
  assign n309 = ~n306 & ~n308;
  assign n310 = pi09 & ~n309;
  assign n311 = pi01 & n159;
  assign n312 = pi05 & n27;
  assign n313 = ~n311 & ~n312;
  assign n314 = ~n33 & n313;
  assign n315 = ~n206 & ~n314;
  assign n316 = ~n297 & ~n310;
  assign n317 = ~n315 & n316;
  assign n318 = ~n305 & n317;
  assign n319 = ~pi13 & ~n318;
  assign n320 = n179 & ~n319;
  assign n321 = ~n295 & n320;
  assign po1 = n296 | ~n321;
  assign n323 = ~pi02 & n71;
  assign n324 = n183 & n300;
  assign n325 = n99 & ~n189;
  assign n326 = ~n258 & ~n325;
  assign n327 = ~pi06 & n326;
  assign n328 = pi09 & n327;
  assign n329 = pi06 & n29;
  assign n330 = ~n326 & n329;
  assign n331 = ~n328 & ~n330;
  assign n332 = pi02 & ~n331;
  assign n333 = pi06 & ~n326;
  assign n334 = n326 & ~n329;
  assign n335 = ~pi02 & pi09;
  assign n336 = ~n333 & n335;
  assign n337 = ~n334 & n336;
  assign n338 = ~n324 & ~n337;
  assign n339 = ~n332 & n338;
  assign n340 = n182 & ~n339;
  assign n341 = pi02 & pi06;
  assign n342 = ~n199 & n341;
  assign n343 = ~pi02 & ~pi06;
  assign n344 = n41 & ~n343;
  assign n345 = ~pi06 & ~n67;
  assign n346 = ~n323 & ~n344;
  assign n347 = ~n345 & n346;
  assign n348 = ~n340 & n347;
  assign n349 = ~n342 & n348;
  assign n350 = ~n97 & n349;
  assign n351 = ~pi06 & n93;
  assign n352 = ~n350 & ~n351;
  assign n353 = ~pi09 & ~n352;
  assign n354 = n27 & ~n349;
  assign n355 = ~pi02 & n43;
  assign n356 = n60 & n355;
  assign n357 = ~n129 & ~n356;
  assign n358 = ~n354 & n357;
  assign n359 = pi06 & ~n358;
  assign n360 = pi02 & pi11;
  assign n361 = ~pi06 & ~pi09;
  assign n362 = n24 & ~n361;
  assign n363 = n360 & ~n362;
  assign n364 = pi02 & n159;
  assign n365 = ~n33 & ~n364;
  assign n366 = ~n349 & ~n365;
  assign n367 = ~n341 & ~n343;
  assign n368 = ~n44 & ~n360;
  assign n369 = pi09 & ~n367;
  assign n370 = ~n368 & n369;
  assign n371 = ~n363 & ~n370;
  assign n372 = ~n366 & n371;
  assign n373 = ~n353 & n372;
  assign n374 = ~n359 & n373;
  assign n375 = ~pi13 & ~n374;
  assign n376 = pi06 & n43;
  assign n377 = n130 & n341;
  assign n378 = ~pi02 & n349;
  assign n379 = n114 & ~n378;
  assign n380 = n23 & n349;
  assign n381 = pi09 & n349;
  assign n382 = pi02 & pi08;
  assign n383 = ~n361 & n382;
  assign n384 = ~n381 & n383;
  assign n385 = ~n380 & ~n384;
  assign n386 = n116 & ~n385;
  assign n387 = ~n379 & ~n386;
  assign n388 = n133 & n387;
  assign n389 = ~n377 & ~n388;
  assign n390 = n349 & n389;
  assign n391 = ~n349 & ~n389;
  assign n392 = ~n390 & ~n391;
  assign n393 = ~n269 & ~n272;
  assign n394 = ~n392 & n393;
  assign n395 = n392 & ~n393;
  assign n396 = ~n394 & ~n395;
  assign n397 = n59 & ~n396;
  assign n398 = pi01 & ~n224;
  assign n399 = ~n226 & ~n398;
  assign n400 = n387 & n399;
  assign n401 = ~n387 & ~n399;
  assign n402 = ~n400 & ~n401;
  assign n403 = pi02 & ~pi08;
  assign n404 = ~n402 & n403;
  assign n405 = ~n376 & ~n404;
  assign n406 = ~n397 & n405;
  assign n407 = n52 & ~n406;
  assign n408 = ~n281 & ~n284;
  assign n409 = n387 & ~n408;
  assign n410 = ~n387 & n408;
  assign n411 = ~n409 & ~n410;
  assign n412 = ~n389 & ~n411;
  assign n413 = n389 & n411;
  assign n414 = ~n412 & ~n413;
  assign n415 = n137 & ~n414;
  assign n416 = n54 & n402;
  assign n417 = pi01 & ~n208;
  assign n418 = ~n207 & ~n417;
  assign n419 = n210 & ~n349;
  assign n420 = n418 & n419;
  assign n421 = ~n416 & ~n420;
  assign n422 = ~pi02 & ~n421;
  assign n423 = pi02 & n32;
  assign n424 = n210 & ~n418;
  assign n425 = ~n423 & ~n424;
  assign n426 = pi02 & ~n418;
  assign n427 = n349 & ~n426;
  assign n428 = ~n425 & n427;
  assign n429 = n32 & ~n349;
  assign n430 = ~n418 & n429;
  assign n431 = ~n241 & ~n430;
  assign n432 = pi02 & ~n431;
  assign n433 = pi11 & n343;
  assign n434 = ~n341 & ~n433;
  assign n435 = ~n56 & ~n188;
  assign n436 = ~n185 & ~n435;
  assign n437 = ~n434 & n436;
  assign n438 = n367 & ~n436;
  assign n439 = ~n437 & ~n438;
  assign n440 = n109 & ~n439;
  assign n441 = n251 & n349;
  assign n442 = ~n246 & n250;
  assign n443 = ~n247 & ~n349;
  assign n444 = ~n442 & n443;
  assign n445 = n231 & n387;
  assign n446 = ~n231 & ~n387;
  assign n447 = ~pi11 & ~n445;
  assign n448 = ~n446 & n447;
  assign n449 = ~pi02 & n252;
  assign n450 = pi02 & ~n252;
  assign n451 = pi11 & ~n449;
  assign n452 = ~n450 & n451;
  assign n453 = n159 & ~n452;
  assign n454 = ~n448 & n453;
  assign n455 = ~n440 & ~n441;
  assign n456 = ~n444 & n455;
  assign n457 = ~n428 & n456;
  assign n458 = ~n432 & n457;
  assign n459 = ~n454 & n458;
  assign n460 = ~n422 & n459;
  assign n461 = ~n407 & n460;
  assign n462 = ~n415 & n461;
  assign n463 = pi13 & ~n462;
  assign n464 = n174 & ~n294;
  assign n465 = n463 & n464;
  assign n466 = ~n463 & ~n464;
  assign n467 = ~n465 & ~n466;
  assign n468 = n179 & ~n375;
  assign po2 = n467 | ~n468;
  assign n470 = ~n51 & ~n132;
  assign po5 = pi03 & pi07;
  assign n472 = ~n470 & po5;
  assign n473 = ~pi03 & ~pi07;
  assign n474 = n41 & ~n473;
  assign n475 = ~pi09 & n29;
  assign n476 = ~pi02 & ~n327;
  assign n477 = ~n333 & ~n476;
  assign n478 = n116 & ~n477;
  assign n479 = ~n475 & ~n478;
  assign n480 = po5 & ~n479;
  assign n481 = pi07 & n116;
  assign n482 = n479 & n481;
  assign n483 = ~n70 & ~n482;
  assign n484 = ~pi03 & ~n483;
  assign n485 = n183 & n360;
  assign n486 = pi09 & n473;
  assign n487 = ~n477 & n486;
  assign n488 = ~n485 & ~n487;
  assign n489 = pi13 & ~n488;
  assign n490 = ~n480 & ~n489;
  assign n491 = ~n484 & n490;
  assign n492 = ~pi08 & ~n491;
  assign n493 = pi03 & n64;
  assign n494 = n477 & n493;
  assign n495 = n67 & ~n494;
  assign n496 = ~pi07 & ~n495;
  assign n497 = ~n474 & ~n496;
  assign n498 = ~n492 & n497;
  assign n499 = ~n472 & n498;
  assign n500 = pi07 & n27;
  assign n501 = ~n33 & ~n500;
  assign n502 = ~n499 & ~n501;
  assign n503 = pi03 & pi11;
  assign n504 = ~pi07 & ~pi09;
  assign n505 = n24 & ~n504;
  assign n506 = n503 & ~n505;
  assign n507 = ~pi03 & n43;
  assign n508 = n60 & n507;
  assign n509 = ~n129 & ~n508;
  assign n510 = pi07 & ~n509;
  assign po4 = po5 | n473;
  assign n512 = ~n44 & ~n503;
  assign n513 = po4 & ~n512;
  assign n514 = pi03 & ~n499;
  assign n515 = n59 & n514;
  assign n516 = pi09 & ~n513;
  assign n517 = ~n515 & n516;
  assign n518 = ~pi07 & n93;
  assign n519 = ~n97 & n499;
  assign n520 = ~pi09 & ~n518;
  assign n521 = ~n519 & n520;
  assign n522 = ~n517 & ~n521;
  assign n523 = ~n506 & ~n510;
  assign n524 = ~n502 & n523;
  assign n525 = ~n522 & n524;
  assign n526 = ~pi13 & ~n525;
  assign n527 = ~n343 & ~n438;
  assign n528 = po5 & n527;
  assign n529 = ~po5 & ~n527;
  assign n530 = pi03 & n529;
  assign n531 = ~n528 & ~n530;
  assign n532 = n109 & ~n531;
  assign n533 = pi07 & n109;
  assign n534 = ~n527 & n533;
  assign n535 = ~pi02 & n418;
  assign n536 = ~n427 & ~n535;
  assign n537 = ~n499 & n536;
  assign n538 = n499 & ~n536;
  assign n539 = ~n537 & ~n538;
  assign n540 = n210 & n539;
  assign n541 = ~pi03 & ~n534;
  assign n542 = ~n540 & n541;
  assign n543 = n32 & ~n539;
  assign n544 = pi03 & ~n241;
  assign n545 = ~n543 & n544;
  assign n546 = ~n542 & ~n545;
  assign n547 = n159 & n503;
  assign n548 = ~n449 & n547;
  assign n549 = n441 & n499;
  assign n550 = ~n390 & ~n395;
  assign n551 = n130 & po5;
  assign n552 = ~pi03 & n498;
  assign n553 = n114 & ~n552;
  assign n554 = n23 & n499;
  assign n555 = n30 & n514;
  assign n556 = n40 & po5;
  assign n557 = ~n554 & ~n556;
  assign n558 = ~n555 & n557;
  assign n559 = n116 & ~n558;
  assign n560 = ~n553 & ~n559;
  assign n561 = n133 & n560;
  assign n562 = ~n551 & ~n561;
  assign n563 = n499 & n562;
  assign n564 = ~n499 & ~n562;
  assign n565 = ~n563 & ~n564;
  assign n566 = n550 & ~n565;
  assign n567 = ~n550 & n565;
  assign n568 = ~n566 & ~n567;
  assign n569 = pi08 & ~n568;
  assign n570 = pi02 & ~n400;
  assign n571 = ~n401 & ~n570;
  assign n572 = n560 & n571;
  assign n573 = ~pi08 & ~n572;
  assign n574 = ~n560 & ~n571;
  assign n575 = ~pi03 & ~n574;
  assign n576 = n573 & n575;
  assign n577 = ~n569 & ~n576;
  assign n578 = n475 & ~n577;
  assign n579 = ~n409 & ~n413;
  assign n580 = n560 & ~n579;
  assign n581 = ~n560 & n579;
  assign n582 = ~n580 & ~n581;
  assign n583 = ~n562 & ~n582;
  assign n584 = n562 & n582;
  assign n585 = ~n583 & ~n584;
  assign n586 = n136 & ~n585;
  assign n587 = ~pi03 & n159;
  assign n588 = n449 & n587;
  assign n589 = n109 & n473;
  assign n590 = n527 & n589;
  assign n591 = pi11 & ~n588;
  assign n592 = ~n590 & n591;
  assign n593 = ~n586 & n592;
  assign n594 = n445 & n560;
  assign n595 = ~n445 & ~n560;
  assign n596 = ~n594 & ~n595;
  assign n597 = n159 & ~n596;
  assign n598 = ~n572 & ~n574;
  assign n599 = pi03 & n23;
  assign n600 = ~n598 & n599;
  assign n601 = ~pi11 & ~n533;
  assign n602 = ~n597 & n601;
  assign n603 = ~n600 & n602;
  assign n604 = ~n593 & ~n603;
  assign n605 = n250 & n349;
  assign n606 = ~n246 & n605;
  assign n607 = ~n247 & ~n606;
  assign n608 = ~n499 & n607;
  assign n609 = ~n532 & ~n548;
  assign n610 = ~n549 & n609;
  assign n611 = ~n608 & n610;
  assign n612 = ~n546 & n611;
  assign n613 = ~n578 & n612;
  assign n614 = ~n604 & n613;
  assign n615 = pi13 & ~n614;
  assign n616 = ~n465 & ~n615;
  assign n617 = n465 & ~n614;
  assign n618 = ~n616 & ~n617;
  assign n619 = n179 & ~n526;
  assign po3 = n618 | ~n619;
  assign n621 = n109 & ~n473;
  assign n622 = ~n529 & n621;
  assign n623 = n536 & ~n552;
  assign n624 = ~n514 & ~n623;
  assign n625 = n31 & ~n624;
  assign n626 = n136 & ~n580;
  assign n627 = ~n584 & n626;
  assign n628 = ~n588 & ~n622;
  assign n629 = ~n625 & n628;
  assign n630 = ~n627 & n629;
  assign n631 = pi11 & ~n630;
  assign n632 = n46 & n605;
  assign n633 = n499 & n632;
  assign n634 = n573 & ~n575;
  assign n635 = pi08 & ~n563;
  assign n636 = ~n567 & n635;
  assign n637 = ~n634 & ~n636;
  assign n638 = n183 & ~n637;
  assign n639 = pi10 & ~n594;
  assign n640 = n30 & ~n639;
  assign n641 = ~n638 & ~n640;
  assign n642 = ~pi11 & ~n641;
  assign n643 = ~n633 & ~n642;
  assign n644 = ~n631 & n643;
  assign n645 = ~n617 & n644;
  assign po6 = pi13 & ~n645;
  assign n647 = ~n73 & ~n189;
  assign n648 = ~n367 & po4;
  assign po7 = n647 & n648;
endmodule
