module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 , pi32 ,
    pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 , pi40 ,
    pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 , pi56 ,
    pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 , pi64 ,
    pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 ,
    pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 ,
    pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 ,
    pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 ,
    pi97 , pi98 , pi99 , pi100 , pi101 , pi102 , pi103 ,
    pi104 , pi105 , pi106 , pi107 , pi108 , pi109 , pi110 ,
    pi111 , pi112 , pi113 , pi114 , pi115 , pi116 , pi117 ,
    pi118 , pi119 , pi120 , pi121 , pi122 , pi123 , pi124 ,
    pi125 , pi126 , pi127 ,
    po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7  );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    pi32 , pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 ,
    pi56 , pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 ,
    pi64 , pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 ,
    pi72 , pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 ,
    pi80 , pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 ,
    pi88 , pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 ,
    pi96 , pi97 , pi98 , pi99 , pi100 , pi101 , pi102 ,
    pi103 , pi104 , pi105 , pi106 , pi107 , pi108 , pi109 ,
    pi110 , pi111 , pi112 , pi113 , pi114 , pi115 , pi116 ,
    pi117 , pi118 , pi119 , pi120 , pi121 , pi122 , pi123 ,
    pi124 , pi125 , pi126 , pi127 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7;
  wire n137, n138, n139, n140, n141, n142, n143,
    n144, n145, n146, n147, n148, n149, n150,
    n151, n152, n153, n154, n155, n156, n157,
    n158, n159, n160, n161, n162, n163, n164,
    n165, n166, n167, n168, n169, n170, n171,
    n172, n173, n174, n175, n176, n177, n178,
    n179, n180, n181, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192,
    n193, n194, n195, n196, n197, n198, n199,
    n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213,
    n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227,
    n228, n229, n230, n231, n232, n233, n234,
    n235, n236, n237, n238, n239, n240, n241,
    n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n340,
    n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403,
    n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416, n417,
    n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438,
    n439, n440, n441, n442, n443, n444, n445,
    n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487,
    n488, n489, n491, n492, n493, n494, n495,
    n496, n497, n498, n499, n500, n501, n502,
    n503, n504, n505, n506, n507, n508, n509,
    n510, n512, n513, n514, n515, n516, n517,
    n518, n519, n520, n521, n522, n523, n524,
    n525, n526, n527, n528, n529, n530, n531,
    n532, n533, n534, n535, n536, n537, n538,
    n539, n540, n541, n542, n543, n544, n545,
    n546, n547, n548, n549, n550, n551, n552,
    n553, n554, n555, n556, n557, n558, n559,
    n560, n562, n563, n564, n565, n566, n567,
    n568, n569, n570, n571, n572, n573, n574,
    n575, n576, n577, n578, n579, n580, n581,
    n582, n584, n585, n586, n587, n588, n589,
    n590, n591, n593, n594, n596, n597, n598,
    n599, n600, n601;
  assign n137 = ~pi124  & ~pi125 ;
  assign n138 = ~pi126  & ~pi127 ;
  assign n139 = n137 & n138;
  assign n140 = ~pi122  & ~pi123 ;
  assign n141 = ~pi120  & ~pi121 ;
  assign n142 = n140 & n141;
  assign n143 = n139 & n142;
  assign n144 = pi125  & ~pi126 ;
  assign n145 = pi121  & ~pi122 ;
  assign n146 = ~pi123  & ~n145;
  assign n147 = n139 & ~n146;
  assign n148 = ~pi127  & ~n144;
  assign n149 = ~n147 & n148;
  assign n150 = ~n143 & n149;
  assign n151 = ~pi118  & ~n150;
  assign n152 = ~pi116  & n151;
  assign n153 = pi119  & n143;
  assign n154 = pi117  & n151;
  assign n155 = n149 & ~n153;
  assign n156 = ~n154 & n155;
  assign n157 = ~n152 & n156;
  assign n158 = ~pi114  & ~n157;
  assign n159 = ~pi112  & n158;
  assign n160 = ~pi110  & n159;
  assign n161 = pi115  & n152;
  assign n162 = pi111  & n159;
  assign n163 = pi113  & n158;
  assign n164 = n156 & ~n161;
  assign n165 = ~n163 & n164;
  assign n166 = ~n162 & n165;
  assign n167 = ~n160 & n166;
  assign n168 = ~pi108  & ~n167;
  assign n169 = ~pi106  & n168;
  assign n170 = pi109  & n160;
  assign n171 = pi107  & n168;
  assign n172 = n166 & ~n170;
  assign n173 = ~n171 & n172;
  assign n174 = ~n169 & n173;
  assign n175 = ~pi104  & ~n174;
  assign n176 = ~pi102  & n175;
  assign n177 = ~pi100  & n176;
  assign n178 = pi105  & n169;
  assign n179 = pi101  & n176;
  assign n180 = pi103  & n175;
  assign n181 = n173 & ~n178;
  assign n182 = ~n180 & n181;
  assign n183 = ~n179 & n182;
  assign n184 = ~n177 & n183;
  assign n185 = ~pi98  & ~n184;
  assign n186 = ~pi96  & n185;
  assign n187 = pi99  & n177;
  assign n188 = pi97  & n185;
  assign n189 = n183 & ~n187;
  assign n190 = ~n188 & n189;
  assign n191 = ~n186 & n190;
  assign n192 = ~pi94  & ~n191;
  assign n193 = ~pi92  & n192;
  assign n194 = ~pi90  & n193;
  assign n195 = pi95  & n186;
  assign n196 = pi91  & n193;
  assign n197 = pi93  & n192;
  assign n198 = n190 & ~n195;
  assign n199 = ~n197 & n198;
  assign n200 = ~n196 & n199;
  assign n201 = ~n194 & n200;
  assign n202 = ~pi88  & ~n201;
  assign n203 = ~pi86  & n202;
  assign n204 = pi89  & n194;
  assign n205 = pi87  & n202;
  assign n206 = n200 & ~n204;
  assign n207 = ~n205 & n206;
  assign n208 = ~n203 & n207;
  assign n209 = ~pi84  & ~n208;
  assign n210 = ~pi82  & n209;
  assign n211 = ~pi80  & n210;
  assign n212 = pi85  & n203;
  assign n213 = pi81  & n210;
  assign n214 = pi83  & n209;
  assign n215 = n207 & ~n212;
  assign n216 = ~n214 & n215;
  assign n217 = ~n213 & n216;
  assign n218 = ~n211 & n217;
  assign n219 = ~pi78  & ~n218;
  assign n220 = ~pi76  & n219;
  assign n221 = pi79  & n211;
  assign n222 = pi77  & n219;
  assign n223 = n217 & ~n221;
  assign n224 = ~n222 & n223;
  assign n225 = ~n220 & n224;
  assign n226 = ~pi74  & ~n225;
  assign n227 = ~pi72  & n226;
  assign n228 = ~pi70  & n227;
  assign n229 = pi75  & n220;
  assign n230 = pi71  & n227;
  assign n231 = pi73  & n226;
  assign n232 = n224 & ~n229;
  assign n233 = ~n231 & n232;
  assign n234 = ~n230 & n233;
  assign n235 = ~n228 & n234;
  assign n236 = ~pi68  & ~n235;
  assign n237 = ~pi66  & n236;
  assign n238 = pi69  & n228;
  assign n239 = pi67  & n236;
  assign n240 = n234 & ~n238;
  assign n241 = ~n239 & n240;
  assign n242 = ~n237 & n241;
  assign n243 = ~pi64  & ~n242;
  assign n244 = ~pi62  & n243;
  assign n245 = ~pi60  & n244;
  assign n246 = pi65  & n237;
  assign n247 = pi61  & n244;
  assign n248 = pi63  & n243;
  assign n249 = n241 & ~n246;
  assign n250 = ~n248 & n249;
  assign n251 = ~n247 & n250;
  assign n252 = ~n245 & n251;
  assign n253 = ~pi58  & ~n252;
  assign n254 = ~pi56  & n253;
  assign n255 = pi59  & n245;
  assign n256 = pi57  & n253;
  assign n257 = n251 & ~n255;
  assign n258 = ~n256 & n257;
  assign n259 = ~n254 & n258;
  assign n260 = ~pi54  & ~n259;
  assign n261 = ~pi52  & n260;
  assign n262 = ~pi50  & n261;
  assign n263 = pi55  & n254;
  assign n264 = pi51  & n261;
  assign n265 = pi53  & n260;
  assign n266 = n258 & ~n263;
  assign n267 = ~n265 & n266;
  assign n268 = ~n264 & n267;
  assign n269 = ~n262 & n268;
  assign n270 = ~pi48  & ~n269;
  assign n271 = ~pi46  & n270;
  assign n272 = pi49  & n262;
  assign n273 = pi47  & n270;
  assign n274 = n268 & ~n272;
  assign n275 = ~n273 & n274;
  assign n276 = ~n271 & n275;
  assign n277 = ~pi44  & ~n276;
  assign n278 = ~pi42  & n277;
  assign n279 = ~pi40  & n278;
  assign n280 = pi45  & n271;
  assign n281 = pi41  & n278;
  assign n282 = pi43  & n277;
  assign n283 = n275 & ~n280;
  assign n284 = ~n282 & n283;
  assign n285 = ~n281 & n284;
  assign n286 = ~n279 & n285;
  assign n287 = ~pi38  & ~n286;
  assign n288 = ~pi36  & n287;
  assign n289 = pi39  & n279;
  assign n290 = pi37  & n287;
  assign n291 = n285 & ~n289;
  assign n292 = ~n290 & n291;
  assign n293 = ~n288 & n292;
  assign n294 = ~pi34  & ~n293;
  assign n295 = ~pi32  & n294;
  assign n296 = ~pi30  & n295;
  assign n297 = pi35  & n288;
  assign n298 = pi31  & n295;
  assign n299 = pi33  & n294;
  assign n300 = n292 & ~n297;
  assign n301 = ~n299 & n300;
  assign n302 = ~n298 & n301;
  assign n303 = ~n296 & n302;
  assign n304 = ~pi28  & ~n303;
  assign n305 = ~pi26  & n304;
  assign n306 = pi25  & n305;
  assign n307 = pi29  & n296;
  assign n308 = pi27  & n304;
  assign n309 = n302 & ~n307;
  assign n310 = ~n308 & n309;
  assign n311 = ~n305 & n310;
  assign n312 = ~pi24  & ~n311;
  assign n313 = ~pi22  & n312;
  assign n314 = pi21  & n313;
  assign n315 = pi23  & n312;
  assign n316 = pi1  & ~pi2 ;
  assign n317 = ~pi3  & ~n316;
  assign n318 = ~pi4  & ~n317;
  assign n319 = ~pi5  & ~n318;
  assign n320 = ~pi6  & ~n319;
  assign n321 = ~pi7  & ~n320;
  assign n322 = ~pi8  & ~n321;
  assign n323 = ~pi9  & ~n322;
  assign n324 = ~pi10  & ~n323;
  assign n325 = ~pi11  & ~n324;
  assign n326 = ~pi12  & ~n325;
  assign n327 = ~pi13  & ~n326;
  assign n328 = ~pi14  & ~n327;
  assign n329 = ~pi15  & ~n328;
  assign n330 = ~pi16  & ~n329;
  assign n331 = ~pi17  & ~n330;
  assign n332 = ~pi18  & ~n331;
  assign n333 = ~pi19  & ~n332;
  assign n334 = ~pi20  & ~n333;
  assign n335 = n313 & n334;
  assign n336 = ~n306 & n310;
  assign n337 = ~n315 & n336;
  assign n338 = ~n314 & n337;
  assign po0  = n335 | ~n338;
  assign n340 = ~pi102  & ~pi103 ;
  assign n341 = ~pi114  & ~pi115 ;
  assign n342 = ~pi118  & ~pi119 ;
  assign n343 = ~pi116  & ~pi117 ;
  assign n344 = n342 & n343;
  assign n345 = ~pi112  & ~pi113 ;
  assign n346 = n341 & n345;
  assign n347 = n344 & n346;
  assign n348 = n143 & n347;
  assign n349 = ~pi110  & ~pi111 ;
  assign n350 = n348 & ~n349;
  assign n351 = ~pi106  & ~pi107 ;
  assign n352 = n137 & ~n140;
  assign n353 = ~n341 & n343;
  assign n354 = n342 & ~n353;
  assign n355 = n143 & ~n354;
  assign n356 = n138 & ~n352;
  assign n357 = ~n355 & n356;
  assign n358 = ~n350 & n351;
  assign n359 = n357 & n358;
  assign n360 = n340 & n359;
  assign n361 = ~pi98  & ~pi99 ;
  assign n362 = n360 & n361;
  assign n363 = ~pi94  & ~pi95 ;
  assign n364 = n362 & n363;
  assign n365 = ~pi92  & ~pi93 ;
  assign n366 = ~pi90  & ~pi91 ;
  assign n367 = ~pi88  & ~pi89 ;
  assign n368 = ~pi86  & ~pi87 ;
  assign n369 = ~pi84  & ~pi85 ;
  assign n370 = ~pi82  & ~pi83 ;
  assign n371 = ~pi80  & ~pi81 ;
  assign n372 = ~pi78  & ~pi79 ;
  assign n373 = ~pi76  & ~pi77 ;
  assign n374 = ~pi74  & ~pi75 ;
  assign n375 = n373 & ~n374;
  assign n376 = n372 & ~n375;
  assign n377 = n371 & ~n376;
  assign n378 = n370 & ~n377;
  assign n379 = n369 & ~n378;
  assign n380 = n368 & ~n379;
  assign n381 = n367 & ~n380;
  assign n382 = n366 & ~n381;
  assign n383 = n365 & ~n382;
  assign n384 = n364 & ~n383;
  assign n385 = ~pi104  & ~pi105 ;
  assign n386 = n359 & ~n385;
  assign n387 = ~pi96  & ~pi97 ;
  assign n388 = n362 & ~n387;
  assign n389 = ~pi100  & ~pi101 ;
  assign n390 = n360 & ~n389;
  assign n391 = ~pi108  & ~pi109 ;
  assign n392 = n349 & ~n391;
  assign n393 = n348 & ~n392;
  assign n394 = n357 & ~n393;
  assign n395 = ~n386 & ~n394;
  assign n396 = ~n390 & n395;
  assign n397 = ~n388 & n396;
  assign n398 = ~n384 & n397;
  assign n399 = n372 & n373;
  assign n400 = ~pi72  & ~pi73 ;
  assign n401 = n374 & n400;
  assign n402 = n399 & n401;
  assign n403 = ~pi70  & ~pi71 ;
  assign n404 = ~pi68  & ~pi69 ;
  assign n405 = n403 & ~n404;
  assign n406 = n364 & ~n365;
  assign n407 = n367 & n369;
  assign n408 = n371 & n407;
  assign n409 = ~n405 & n408;
  assign n410 = n402 & n409;
  assign n411 = n397 & n410;
  assign n412 = ~n406 & n411;
  assign n413 = ~n398 & ~n412;
  assign n414 = ~pi66  & ~pi67 ;
  assign n415 = n403 & n414;
  assign n416 = ~n398 & n415;
  assign n417 = ~n413 & ~n416;
  assign n418 = ~pi64  & ~pi65 ;
  assign n419 = ~pi62  & ~pi63 ;
  assign n420 = ~pi60  & ~pi61 ;
  assign n421 = n419 & ~n420;
  assign n422 = n418 & ~n421;
  assign n423 = ~n413 & n422;
  assign n424 = ~n417 & ~n423;
  assign n425 = ~pi56  & ~pi57 ;
  assign n426 = ~pi54  & ~pi55 ;
  assign n427 = n425 & ~n426;
  assign n428 = ~pi58  & ~pi59 ;
  assign n429 = n419 & n428;
  assign n430 = ~n417 & n429;
  assign n431 = ~pi50  & ~pi51 ;
  assign n432 = ~pi48  & ~pi49 ;
  assign n433 = ~pi46  & ~pi47 ;
  assign n434 = ~pi44  & ~pi45 ;
  assign n435 = n433 & ~n434;
  assign n436 = ~pi42  & ~pi43 ;
  assign n437 = ~pi38  & ~pi39 ;
  assign n438 = ~pi36  & ~pi37 ;
  assign n439 = n437 & ~n438;
  assign n440 = ~pi40  & ~pi41 ;
  assign n441 = ~pi32  & ~pi33 ;
  assign n442 = ~pi30  & ~pi31 ;
  assign n443 = n441 & ~n442;
  assign n444 = ~pi26  & ~pi27 ;
  assign n445 = ~pi28  & ~pi29 ;
  assign n446 = n441 & n445;
  assign n447 = ~n444 & n446;
  assign n448 = ~pi34  & ~pi35 ;
  assign n449 = ~pi22  & ~pi23 ;
  assign n450 = ~pi20  & ~pi21 ;
  assign n451 = ~pi18  & ~pi19 ;
  assign n452 = ~pi16  & ~pi17 ;
  assign n453 = ~pi14  & ~pi15 ;
  assign n454 = ~pi12  & ~pi13 ;
  assign n455 = ~pi10  & ~pi11 ;
  assign n456 = ~pi8  & ~pi9 ;
  assign n457 = ~pi6  & ~pi7 ;
  assign n458 = ~pi4  & ~pi5 ;
  assign n459 = ~pi2  & ~pi3 ;
  assign n460 = n458 & ~n459;
  assign n461 = n457 & ~n460;
  assign n462 = n456 & ~n461;
  assign n463 = n455 & ~n462;
  assign n464 = n454 & ~n463;
  assign n465 = n453 & ~n464;
  assign n466 = n452 & ~n465;
  assign n467 = n451 & ~n466;
  assign n468 = n450 & ~n467;
  assign n469 = n449 & ~n468;
  assign n470 = ~pi24  & ~pi25 ;
  assign n471 = n446 & n470;
  assign n472 = ~n469 & n471;
  assign n473 = n437 & n448;
  assign n474 = ~n443 & n473;
  assign n475 = ~n447 & n474;
  assign n476 = ~n472 & n475;
  assign n477 = ~n439 & n440;
  assign n478 = ~n476 & n477;
  assign n479 = n433 & n436;
  assign n480 = ~n478 & n479;
  assign n481 = n432 & ~n435;
  assign n482 = ~n480 & n481;
  assign n483 = n431 & ~n482;
  assign n484 = ~n425 & n430;
  assign n485 = ~pi52  & ~pi53 ;
  assign n486 = ~n483 & n485;
  assign n487 = ~n484 & n486;
  assign n488 = ~n427 & n430;
  assign n489 = ~n487 & n488;
  assign po1  = ~n424 & ~n489;
  assign n491 = n349 & n391;
  assign n492 = n351 & n385;
  assign n493 = n491 & n492;
  assign n494 = n340 & n389;
  assign n495 = n361 & n387;
  assign n496 = n494 & n495;
  assign n497 = n493 & n496;
  assign n498 = n348 & n497;
  assign n499 = n403 & n404;
  assign n500 = n414 & n418;
  assign n501 = n499 & n500;
  assign n502 = n402 & n501;
  assign n503 = n366 & n367;
  assign n504 = n363 & n365;
  assign n505 = n368 & n369;
  assign n506 = n370 & n371;
  assign n507 = n505 & n506;
  assign n508 = n503 & n504;
  assign n509 = n507 & n508;
  assign n510 = n502 & n509;
  assign po6  = ~n498 | ~n510;
  assign n512 = n419 & n420;
  assign n513 = n426 & n485;
  assign n514 = n425 & n428;
  assign n515 = ~n513 & n514;
  assign n516 = n512 & ~n515;
  assign n517 = ~po6  & ~n516;
  assign n518 = n142 & ~n344;
  assign n519 = n492 & ~n494;
  assign n520 = n401 & ~n499;
  assign n521 = n399 & ~n520;
  assign n522 = n506 & ~n521;
  assign n523 = n505 & ~n522;
  assign n524 = n503 & ~n523;
  assign n525 = n504 & ~n524;
  assign n526 = n497 & ~n525;
  assign n527 = n491 & ~n519;
  assign n528 = ~n526 & n527;
  assign n529 = n348 & ~n528;
  assign n530 = n139 & ~n518;
  assign n531 = ~n529 & n530;
  assign n532 = n431 & n432;
  assign n533 = n433 & n434;
  assign n534 = n436 & n440;
  assign n535 = n437 & n438;
  assign n536 = n441 & n448;
  assign n537 = n442 & n445;
  assign n538 = n444 & n470;
  assign n539 = n449 & n450;
  assign n540 = n451 & n452;
  assign n541 = n453 & n454;
  assign n542 = n455 & n456;
  assign n543 = n457 & n458;
  assign n544 = n542 & ~n543;
  assign n545 = n541 & ~n544;
  assign n546 = n540 & ~n545;
  assign n547 = n539 & ~n546;
  assign n548 = n538 & ~n547;
  assign n549 = n537 & ~n548;
  assign n550 = n536 & ~n549;
  assign n551 = n535 & ~n550;
  assign n552 = n534 & ~n551;
  assign n553 = n533 & ~n552;
  assign n554 = n532 & ~n553;
  assign n555 = ~n517 & n531;
  assign n556 = ~n554 & n555;
  assign n557 = n512 & ~n514;
  assign n558 = ~po6  & ~n557;
  assign n559 = n531 & ~n558;
  assign n560 = n554 & n559;
  assign po2  = ~n556 & ~n560;
  assign n562 = n347 & ~n493;
  assign n563 = n143 & ~n562;
  assign n564 = ~n498 & n563;
  assign n565 = n512 & n514;
  assign n566 = n513 & n532;
  assign n567 = n533 & n534;
  assign n568 = n535 & n536;
  assign n569 = n537 & n538;
  assign n570 = n539 & n540;
  assign n571 = n541 & n542;
  assign n572 = n570 & ~n571;
  assign n573 = n569 & ~n572;
  assign n574 = n568 & ~n573;
  assign n575 = n567 & ~n574;
  assign n576 = n566 & ~n575;
  assign n577 = n565 & ~n576;
  assign n578 = n501 & ~n577;
  assign n579 = n402 & ~n578;
  assign n580 = n507 & ~n579;
  assign n581 = n498 & n508;
  assign n582 = ~n580 & n581;
  assign po3  = ~n564 & ~n582;
  assign n584 = n565 & n566;
  assign n585 = n569 & n570;
  assign n586 = n567 & n568;
  assign n587 = ~n585 & n586;
  assign n588 = n584 & ~n587;
  assign n589 = n502 & ~n588;
  assign n590 = n509 & ~n589;
  assign n591 = n497 & ~n590;
  assign po4  = ~n348 | n591;
  assign n593 = n584 & n586;
  assign n594 = n510 & ~n593;
  assign po5  = ~n498 | n594;
  assign n596 = ~pi0  & ~pi1 ;
  assign n597 = n459 & n596;
  assign n598 = n543 & n597;
  assign n599 = n571 & n598;
  assign n600 = n585 & n599;
  assign n601 = n593 & n600;
  assign po7 = po6  | ~n601;
endmodule
