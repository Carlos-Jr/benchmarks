module i2c ( 
    pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8, pi9,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19,
    pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29,
    pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38, pi39,
    pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48, pi49,
    pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59,
    pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69,
    pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79,
    pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88, pi89,
    pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97, pi98, pi99,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146,
    po0, po1, po2, po3, po4, po5, po6, po7, po8, po9,
    po10, po11, po12, po13, po14, po15, po16, po17, po18, po19,
    po20, po21, po22, po23, po24, po25, po26, po27, po28, po29,
    po30, po31, po32, po33, po34, po35, po36, po37, po38, po39,
    po40, po41, po42, po43, po44, po45, po46, po47, po48, po49,
    po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66, po67, po68, po69,
    po70, po71, po72, po73, po74, po75, po76, po77, po78, po79,
    po80, po81, po82, po83, po84, po85, po86, po87, po88, po89,
    po90, po91, po92, po93, po94, po95, po96, po97, po98, po99,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141  );
  input  pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8,
    pi9, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18,
    pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28,
    pi29, pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38,
    pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48,
    pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58,
    pi59, pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68,
    pi69, pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78,
    pi79, pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88,
    pi89, pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97, pi98,
    pi99, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146;
  output po0, po1, po2, po3, po4, po5, po6, po7, po8, po9,
    po10, po11, po12, po13, po14, po15, po16, po17, po18, po19,
    po20, po21, po22, po23, po24, po25, po26, po27, po28, po29,
    po30, po31, po32, po33, po34, po35, po36, po37, po38, po39,
    po40, po41, po42, po43, po44, po45, po46, po47, po48, po49,
    po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66, po67, po68, po69,
    po70, po71, po72, po73, po74, po75, po76, po77, po78, po79,
    po80, po81, po82, po83, po84, po85, po86, po87, po88, po89,
    po90, po91, po92, po93, po94, po95, po96, po97, po98, po99,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141;
  wire n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n340,
    n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n375, n376,
    n377, n378, n379, n380, n381, n382, n383,
    n384, n385, n386, n387, n388, n389, n390,
    n391, n392, n393, n394, n395, n396, n397,
    n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n408, n409, n410, n411, n412,
    n413, n414, n415, n416, n417, n419, n420,
    n421, n422, n423, n424, n425, n426, n427,
    n428, n430, n431, n432, n433, n434, n435,
    n436, n437, n438, n439, n440, n442, n443,
    n444, n445, n446, n447, n448, n450, n451,
    n452, n453, n454, n455, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466,
    n468, n469, n470, n471, n472, n473, n475,
    n476, n477, n478, n479, n480, n481, n482,
    n483, n485, n486, n487, n488, n489, n490,
    n492, n493, n494, n495, n496, n497, n499,
    n500, n501, n502, n503, n504, n505, n506,
    n508, n509, n510, n511, n512, n513, n514,
    n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n542, n543, n544,
    n545, n546, n547, n549, n550, n551, n552,
    n553, n554, n555, n556, n558, n559, n560,
    n561, n562, n563, n565, n566, n567, n568,
    n569, n570, n572, n573, n574, n575, n576,
    n577, n578, n579, n580, n581, n582, n583,
    n584, n585, n586, n587, n588, n589, n591,
    n592, n593, n594, n595, n596, n597, n599,
    n600, n601, n602, n603, n604, n605, n606,
    n608, n609, n611, n612, n613, n614, n615,
    n616, n617, n618, n619, n620, n621, n622,
    n623, n624, n625, n626, n627, n628, n630,
    n631, n632, n633, n634, n635, n636, n637,
    n638, n639, n640, n641, n642, n643, n644,
    n645, n646, n647, n648, n649, n650, n651,
    n652, n653, n654, n655, n656, n657, n658,
    n659, n660, n661, n662, n663, n664, n665,
    n666, n667, n668, n669, n670, n671, n672,
    n673, n675, n676, n677, n678, n679, n680,
    n682, n683, n684, n685, n686, n687, n688,
    n689, n690, n692, n693, n694, n695, n696,
    n697, n698, n699, n700, n701, n702, n703,
    n704, n705, n706, n707, n708, n709, n710,
    n711, n712, n713, n714, n715, n716, n717,
    n718, n719, n720, n721, n722, n723, n724,
    n725, n726, n727, n728, n729, n730, n732,
    n733, n734, n735, n736, n737, n738, n739,
    n740, n741, n742, n743, n744, n745, n746,
    n747, n748, n749, n750, n751, n752, n753,
    n754, n755, n756, n757, n758, n759, n760,
    n761, n763, n764, n765, n766, n767, n768,
    n770, n771, n772, n773, n774, n775, n777,
    n778, n779, n780, n781, n782, n784, n785,
    n786, n787, n788, n789, n791, n792, n793,
    n794, n795, n796, n798, n799, n800, n801,
    n802, n803, n805, n806, n807, n808, n809,
    n810, n812, n813, n814, n815, n816, n817,
    n819, n820, n821, n822, n823, n824, n825,
    n826, n827, n828, n829, n830, n831, n832,
    n833, n834, n835, n836, n837, n838, n839,
    n840, n841, n843, n844, n845, n846, n847,
    n848, n850, n851, n852, n853, n854, n855,
    n856, n857, n858, n859, n860, n861, n862,
    n863, n864, n865, n867, n868, n869, n870,
    n871, n872, n873, n874, n875, n876, n877,
    n878, n879, n881, n882, n883, n884, n885,
    n886, n887, n888, n889, n890, n891, n892,
    n894, n895, n896, n897, n898, n899, n900,
    n901, n902, n903, n904, n905, n906, n907,
    n908, n909, n911, n912, n913, n914, n915,
    n916, n918, n919, n920, n921, n922, n923,
    n924, n925, n926, n927, n928, n929, n930,
    n931, n933, n934, n935, n936, n937, n938,
    n939, n940, n941, n942, n944, n945, n946,
    n947, n948, n949, n950, n951, n952, n953,
    n954, n955, n956, n958, n959, n960, n961,
    n962, n963, n964, n965, n966, n967, n968,
    n969, n970, n971, n973, n974, n975, n976,
    n977, n978, n979, n980, n981, n982, n983,
    n984, n985, n986, n988, n989, n990, n991,
    n992, n993, n994, n995, n996, n997, n998,
    n999, n1000, n1002, n1003, n1004, n1006,
    n1007, n1008, n1010, n1011, n1012, n1013,
    n1014, n1015, n1016, n1017, n1018, n1020,
    n1021, n1022, n1025, n1027, n1028, n1029,
    n1030, n1031, n1032, n1033, n1034, n1035,
    n1036, n1037, n1038, n1039, n1040, n1041,
    n1042, n1043, n1044, n1045, n1047, n1048,
    n1049, n1050, n1051, n1052, n1053, n1054,
    n1055, n1056, n1057, n1058, n1059, n1060,
    n1062, n1063, n1064, n1065, n1066, n1067,
    n1069, n1070, n1071, n1072, n1073, n1074,
    n1075, n1076, n1077, n1078, n1079, n1080,
    n1081, n1082, n1083, n1084, n1085, n1086,
    n1088, n1089, n1090, n1092, n1093, n1095,
    n1096, n1097, n1098, n1099, n1100, n1101,
    n1102, n1104, n1105, n1106, n1108, n1109,
    n1110, n1112, n1113, n1114, n1116, n1117,
    n1118, n1119, n1120, n1122, n1123, n1124,
    n1126, n1127, n1128, n1130, n1131, n1132,
    n1134, n1135, n1136, n1138, n1139, n1140,
    n1142, n1143, n1144, n1146, n1147, n1148,
    n1150, n1151, n1152, n1154, n1155, n1156,
    n1158, n1159, n1160, n1162, n1163, n1164,
    n1166, n1167, n1168, n1169, n1170, n1172,
    n1173, n1174, n1176, n1177, n1178, n1180,
    n1181, n1182, n1184, n1185, n1186, n1188,
    n1189, n1190, n1191, n1192, n1193, n1194,
    n1195, n1196, n1197, n1198, n1199, n1200,
    n1201, n1202, n1203, n1204, n1205, n1207,
    n1208, n1209, n1211, n1212, n1213, n1214,
    n1216, n1217, n1218, n1220, n1221, n1222,
    n1224, n1225, n1226, n1227, n1228, n1230,
    n1231, n1232, n1234, n1235, n1236, n1238,
    n1239, n1240, n1242, n1243, n1244, n1246,
    n1247, n1248, n1250, n1251, n1252, n1253,
    n1254, n1255, n1257, n1258, n1259, n1260,
    n1261, n1262, n1264, n1265, n1266, n1268,
    n1269, n1270, n1272, n1273, n1274, n1276,
    n1277, n1278, n1280, n1281, n1282, n1284,
    n1285, n1286, n1287, n1288, n1289, n1290,
    n1291, n1292, n1293, n1294, n1295, n1296,
    n1297, n1298, n1299, n1300, n1302, n1303,
    n1304, n1305, n1306, n1307, n1308, n1309,
    n1310, n1311, n1312, n1313, n1314, n1315,
    n1317, n1318, n1319, n1320, n1321, n1322,
    n1323, n1324, n1325, n1326, n1327, n1328,
    n1329, n1330, n1332, n1333, n1334, n1335,
    n1336, n1337, n1338, n1339, n1340, n1341,
    n1342, n1343, n1344, n1345, n1347, n1348,
    n1349, n1350, n1351, n1352, n1353, n1354,
    n1355, n1356, n1357, n1358, n1359, n1360,
    n1361, n1362, n1363, n1365, n1366, n1367,
    n1369, n1370, n1371, n1372, n1373, n1374,
    n1375, n1376, n1377, n1378, n1379, n1380,
    n1381, n1382, n1383, n1384, n1385, n1387,
    n1388, n1389, n1390, n1391, n1392, n1393,
    n1394, n1395, n1396, n1397, n1398, n1399,
    n1400, n1401, n1402, n1403, n1405, n1406,
    n1408, n1409, n1411, n1412, n1413, n1414,
    n1416, n1417, n1418, n1420, n1421, n1422,
    n1423, n1425, n1426, n1427, n1429, n1430,
    n1431, n1434, n1435, n1436, n1437, n1440,
    n1441, n1443, n1448, n1449, n1451;
  assign n291 = ~pi17 & ~pi21;
  assign n292 = ~pi8 & n291;
  assign n293 = ~pi4 & ~pi19;
  assign n294 = ~pi18 & n293;
  assign n295 = ~pi16 & n294;
  assign n296 = ~pi6 & ~pi12;
  assign n297 = ~pi5 & n296;
  assign n298 = ~pi7 & ~pi13;
  assign n299 = ~pi14 & ~pi22;
  assign n300 = ~pi9 & ~pi11;
  assign n301 = n298 & n299;
  assign n302 = n300 & n301;
  assign n303 = n292 & n297;
  assign n304 = n302 & n303;
  assign n305 = n295 & n304;
  assign n306 = pi54 & ~n305;
  assign n307 = ~pi0 & ~n306;
  assign n308 = ~pi5 & ~pi22;
  assign n309 = ~pi56 & ~n308;
  assign n310 = ~pi8 & ~pi21;
  assign n311 = ~pi7 & n310;
  assign n312 = pi8 & pi21;
  assign n313 = pi7 & ~n310;
  assign n314 = ~pi13 & ~n312;
  assign n315 = ~n313 & n314;
  assign n316 = ~n311 & ~n315;
  assign n317 = n298 & n310;
  assign n318 = ~n316 & ~n317;
  assign n319 = ~pi14 & ~n318;
  assign n320 = pi14 & ~n317;
  assign n321 = ~pi10 & ~n320;
  assign n322 = ~n319 & n321;
  assign n323 = ~pi14 & n310;
  assign n324 = pi10 & n298;
  assign n325 = n323 & n324;
  assign n326 = ~n322 & ~n325;
  assign n327 = ~pi17 & n296;
  assign n328 = n308 & n327;
  assign n329 = n295 & n328;
  assign n330 = ~n326 & n329;
  assign n331 = ~n309 & ~n330;
  assign n332 = n300 & ~n331;
  assign n333 = ~pi56 & ~n300;
  assign n334 = n308 & n333;
  assign n335 = ~n332 & ~n334;
  assign n336 = pi54 & ~n335;
  assign n337 = ~n307 & ~n336;
  assign n338 = ~pi3 & ~pi129;
  assign po15 = n337 | ~n338;
  assign n340 = ~pi17 & pi54;
  assign n341 = ~pi11 & ~pi12;
  assign n342 = ~pi10 & ~pi22;
  assign n343 = ~pi5 & ~pi6;
  assign n344 = n298 & n343;
  assign n345 = n295 & n344;
  assign n346 = n341 & n342;
  assign n347 = n323 & n346;
  assign n348 = n345 & n347;
  assign n349 = n340 & ~n348;
  assign n350 = ~pi1 & ~n349;
  assign n351 = ~pi5 & ~pi7;
  assign n352 = pi13 & n296;
  assign n353 = n351 & n352;
  assign n354 = ~pi7 & ~pi12;
  assign n355 = ~n343 & ~n354;
  assign n356 = n296 & n351;
  assign n357 = ~n296 & ~n351;
  assign n358 = ~pi13 & ~n355;
  assign n359 = ~n356 & ~n357;
  assign n360 = n358 & n359;
  assign n361 = ~pi9 & ~n353;
  assign n362 = ~n360 & n361;
  assign n363 = ~pi10 & pi54;
  assign n364 = n299 & n363;
  assign n365 = ~pi8 & ~pi11;
  assign n366 = n291 & n365;
  assign n367 = n297 & n298;
  assign n368 = pi9 & ~n367;
  assign n369 = n364 & n366;
  assign n370 = n295 & n369;
  assign n371 = ~n368 & n370;
  assign n372 = ~n362 & n371;
  assign n373 = ~n350 & ~n372;
  assign po16 = ~n338 | n373;
  assign n375 = ~pi15 & ~pi20;
  assign n376 = ~pi24 & ~pi49;
  assign n377 = ~pi45 & n375;
  assign n378 = n376 & n377;
  assign n379 = ~pi41 & ~pi43;
  assign n380 = ~pi42 & ~pi44;
  assign n381 = ~pi38 & ~pi50;
  assign n382 = ~pi46 & n381;
  assign n383 = ~pi40 & n382;
  assign n384 = n380 & n383;
  assign n385 = n379 & n384;
  assign n386 = ~pi47 & n385;
  assign n387 = ~pi48 & n386;
  assign n388 = pi82 & n378;
  assign n389 = n387 & n388;
  assign n390 = pi122 & pi127;
  assign n391 = ~pi82 & ~n390;
  assign n392 = pi2 & ~n391;
  assign n393 = ~n389 & n392;
  assign n394 = ~pi40 & n380;
  assign n395 = ~pi41 & ~pi46;
  assign n396 = n381 & n395;
  assign n397 = ~pi43 & ~pi47;
  assign n398 = ~pi48 & n397;
  assign n399 = ~pi2 & n398;
  assign n400 = n378 & n399;
  assign n401 = n396 & n400;
  assign n402 = n394 & n401;
  assign n403 = pi82 & ~n402;
  assign n404 = ~pi65 & ~n390;
  assign n405 = ~n403 & n404;
  assign n406 = ~n393 & ~n405;
  assign po17 = ~pi129 & ~n406;
  assign n408 = pi0 & ~pi113;
  assign n409 = ~pi123 & n408;
  assign n410 = ~pi9 & ~pi14;
  assign n411 = n342 & n410;
  assign n412 = ~pi12 & n366;
  assign n413 = n411 & n412;
  assign n414 = n345 & n413;
  assign n415 = ~pi61 & ~pi118;
  assign n416 = ~n414 & n415;
  assign n417 = ~n409 & ~n416;
  assign po18 = ~pi129 & ~n417;
  assign n419 = pi4 & ~pi54;
  assign n420 = ~pi16 & pi54;
  assign n421 = n291 & n420;
  assign n422 = n294 & n421;
  assign n423 = n365 & n422;
  assign n424 = n367 & n410;
  assign n425 = pi10 & ~pi22;
  assign n426 = n423 & n425;
  assign n427 = n424 & n426;
  assign n428 = ~n419 & ~n427;
  assign po19 = n338 & ~n428;
  assign n430 = pi5 & ~pi54;
  assign n431 = n356 & n420;
  assign n432 = ~pi13 & n411;
  assign n433 = ~pi59 & n366;
  assign n434 = n432 & n433;
  assign n435 = ~pi25 & pi28;
  assign n436 = ~pi29 & n435;
  assign n437 = n294 & n436;
  assign n438 = n431 & n437;
  assign n439 = n434 & n438;
  assign n440 = ~n430 & ~n439;
  assign po20 = n338 & ~n440;
  assign n442 = pi6 & ~pi54;
  assign n443 = ~pi28 & ~pi29;
  assign n444 = pi25 & n443;
  assign n445 = n294 & n444;
  assign n446 = n431 & n445;
  assign n447 = n434 & n446;
  assign n448 = ~n442 & ~n447;
  assign po21 = n338 & ~n448;
  assign n450 = pi7 & ~pi54;
  assign n451 = ~pi11 & n356;
  assign n452 = pi8 & n422;
  assign n453 = n432 & n451;
  assign n454 = n452 & n453;
  assign n455 = ~n450 & ~n454;
  assign po22 = n338 & ~n455;
  assign n457 = pi8 & ~pi54;
  assign n458 = ~pi17 & ~pi18;
  assign n459 = n365 & n458;
  assign n460 = n293 & n420;
  assign n461 = ~pi12 & n411;
  assign n462 = n344 & n461;
  assign n463 = pi21 & n459;
  assign n464 = n460 & n463;
  assign n465 = n462 & n464;
  assign n466 = ~n457 & ~n465;
  assign po23 = n338 & ~n466;
  assign n468 = pi9 & ~pi54;
  assign n469 = ~pi8 & n422;
  assign n470 = pi11 & n356;
  assign n471 = n432 & n470;
  assign n472 = n469 & n471;
  assign n473 = ~n468 & ~n472;
  assign po24 = n338 & ~n473;
  assign n475 = pi10 & ~pi54;
  assign n476 = ~pi9 & ~pi18;
  assign n477 = n292 & n476;
  assign n478 = n342 & n477;
  assign n479 = ~pi13 & pi14;
  assign n480 = n460 & n479;
  assign n481 = n451 & n480;
  assign n482 = n478 & n481;
  assign n483 = ~n475 & ~n482;
  assign po25 = n338 & ~n483;
  assign n485 = pi11 & ~pi54;
  assign n486 = ~pi10 & ~pi11;
  assign n487 = pi22 & n486;
  assign n488 = n424 & n487;
  assign n489 = n469 & n488;
  assign n490 = ~n485 & ~n489;
  assign po26 = n338 & ~n490;
  assign n492 = pi12 & ~pi54;
  assign n493 = pi18 & n344;
  assign n494 = n411 & n460;
  assign n495 = n493 & n494;
  assign n496 = n412 & n495;
  assign n497 = ~n492 & ~n496;
  assign po27 = n338 & ~n497;
  assign n499 = pi13 & ~pi54;
  assign n500 = ~pi25 & ~pi28;
  assign n501 = pi29 & n500;
  assign n502 = ~pi59 & n342;
  assign n503 = n501 & n502;
  assign n504 = n423 & n503;
  assign n505 = n424 & n504;
  assign n506 = ~n499 & ~n505;
  assign po28 = n338 & ~n506;
  assign n508 = pi14 & ~pi54;
  assign n509 = pi13 & ~pi16;
  assign n510 = n293 & n509;
  assign n511 = n364 & n510;
  assign n512 = n451 & n511;
  assign n513 = n477 & n512;
  assign n514 = ~n508 & ~n513;
  assign po29 = n338 & ~n514;
  assign n516 = ~pi82 & n390;
  assign n517 = pi15 & n516;
  assign n518 = ~pi45 & n376;
  assign n519 = n394 & n396;
  assign n520 = n398 & n518;
  assign n521 = n519 & n520;
  assign n522 = pi15 & ~n521;
  assign n523 = ~pi47 & ~pi48;
  assign n524 = ~pi45 & n523;
  assign n525 = ~pi2 & ~pi20;
  assign n526 = ~pi15 & n376;
  assign n527 = n524 & ~n525;
  assign n528 = n526 & n527;
  assign n529 = n385 & n528;
  assign n530 = ~n522 & ~n529;
  assign n531 = pi82 & ~n530;
  assign n532 = ~pi15 & n379;
  assign n533 = n523 & n532;
  assign n534 = n518 & n533;
  assign n535 = n384 & n534;
  assign n536 = pi82 & ~n535;
  assign n537 = ~pi70 & ~n390;
  assign n538 = ~n536 & n537;
  assign n539 = ~n517 & ~n538;
  assign n540 = ~n531 & n539;
  assign po30 = ~pi129 & ~n540;
  assign n542 = pi16 & ~pi54;
  assign n543 = pi6 & ~pi13;
  assign n544 = n351 & n543;
  assign n545 = n461 & n544;
  assign n546 = n423 & n545;
  assign n547 = ~n542 & ~n546;
  assign po31 = n338 & ~n547;
  assign n549 = pi17 & ~pi54;
  assign n550 = ~pi25 & pi59;
  assign n551 = n310 & n550;
  assign n552 = n340 & n443;
  assign n553 = n551 & n552;
  assign n554 = n295 & n553;
  assign n555 = n453 & n554;
  assign n556 = ~n549 & ~n555;
  assign po32 = n338 & ~n556;
  assign n558 = pi18 & ~pi54;
  assign n559 = n294 & n462;
  assign n560 = pi16 & pi54;
  assign n561 = n366 & n560;
  assign n562 = n559 & n561;
  assign n563 = ~n558 & ~n562;
  assign po33 = n338 & ~n563;
  assign n565 = pi19 & ~pi54;
  assign n566 = pi17 & ~pi21;
  assign n567 = n365 & n566;
  assign n568 = n420 & n567;
  assign n569 = n559 & n568;
  assign n570 = ~n565 & ~n569;
  assign po34 = n338 & ~n570;
  assign n572 = pi20 & n516;
  assign n573 = n379 & n524;
  assign n574 = ~pi38 & n394;
  assign n575 = ~pi50 & n574;
  assign n576 = ~pi46 & n575;
  assign n577 = n573 & n576;
  assign n578 = n376 & n577;
  assign n579 = n375 & n578;
  assign n580 = pi2 & n579;
  assign n581 = ~pi15 & n578;
  assign n582 = pi20 & ~n581;
  assign n583 = ~n580 & ~n582;
  assign n584 = pi82 & ~n583;
  assign n585 = pi82 & ~n579;
  assign n586 = ~pi71 & ~n390;
  assign n587 = ~n585 & n586;
  assign n588 = ~n572 & ~n587;
  assign n589 = ~n584 & n588;
  assign po35 = ~pi129 & ~n589;
  assign n591 = pi21 & ~pi54;
  assign n592 = ~pi4 & pi19;
  assign n593 = ~pi21 & n592;
  assign n594 = n420 & n593;
  assign n595 = n459 & n594;
  assign n596 = n462 & n595;
  assign n597 = ~n591 & ~n596;
  assign po36 = n338 & ~n597;
  assign n599 = pi22 & ~pi54;
  assign n600 = pi5 & ~pi6;
  assign n601 = ~pi14 & n600;
  assign n602 = n298 & n341;
  assign n603 = n601 & n602;
  assign n604 = n460 & n603;
  assign n605 = n478 & n604;
  assign n606 = ~n599 & ~n605;
  assign po37 = n338 & ~n606;
  assign n608 = ~pi23 & pi55;
  assign n609 = pi61 & ~pi129;
  assign po38 = ~n608 & n609;
  assign n611 = ~pi2 & n375;
  assign n612 = ~pi49 & n611;
  assign n613 = pi82 & ~n612;
  assign n614 = n390 & ~n613;
  assign n615 = n384 & n573;
  assign n616 = pi82 & ~n615;
  assign n617 = ~n614 & ~n616;
  assign n618 = ~pi24 & ~n617;
  assign n619 = pi24 & pi82;
  assign n620 = n577 & n619;
  assign n621 = ~pi45 & ~pi49;
  assign n622 = n611 & n621;
  assign n623 = n387 & n622;
  assign n624 = pi82 & ~n623;
  assign n625 = pi63 & ~n390;
  assign n626 = ~n624 & n625;
  assign n627 = ~pi129 & ~n620;
  assign n628 = ~n618 & n627;
  assign po39 = ~n626 & n628;
  assign n630 = ~pi53 & ~pi58;
  assign n631 = pi25 & ~pi116;
  assign n632 = ~pi27 & ~pi85;
  assign n633 = ~pi26 & n631;
  assign n634 = n632 & n633;
  assign n635 = ~n630 & ~n634;
  assign n636 = ~pi53 & pi58;
  assign n637 = pi53 & ~pi58;
  assign n638 = ~n636 & ~n637;
  assign n639 = pi85 & pi116;
  assign n640 = ~pi85 & ~pi110;
  assign n641 = ~pi96 & n640;
  assign n642 = ~n639 & ~n641;
  assign n643 = pi100 & ~n642;
  assign n644 = pi85 & ~pi116;
  assign n645 = pi25 & n644;
  assign n646 = ~n643 & ~n645;
  assign n647 = ~pi26 & ~n646;
  assign n648 = ~pi39 & ~pi52;
  assign n649 = ~pi51 & n648;
  assign n650 = pi116 & n649;
  assign n651 = ~pi85 & ~n650;
  assign n652 = pi26 & n651;
  assign n653 = ~pi25 & ~pi116;
  assign n654 = n652 & ~n653;
  assign n655 = ~n647 & ~n654;
  assign n656 = ~pi27 & ~n655;
  assign n657 = ~n631 & ~n650;
  assign n658 = pi27 & ~n657;
  assign n659 = ~pi95 & ~pi100;
  assign n660 = ~pi97 & n659;
  assign n661 = ~pi110 & ~n660;
  assign n662 = ~pi51 & ~pi52;
  assign n663 = ~pi39 & n662;
  assign n664 = pi27 & ~n663;
  assign n665 = pi25 & ~n661;
  assign n666 = ~n664 & n665;
  assign n667 = ~n658 & ~n666;
  assign n668 = ~pi26 & ~pi85;
  assign n669 = ~n667 & n668;
  assign n670 = ~n656 & ~n669;
  assign n671 = ~pi53 & ~n670;
  assign n672 = n638 & ~n671;
  assign n673 = n338 & ~n635;
  assign po40 = ~n672 & n673;
  assign n675 = ~pi27 & ~pi53;
  assign n676 = ~pi58 & n675;
  assign n677 = pi26 & pi116;
  assign n678 = n643 & ~n677;
  assign n679 = ~n652 & ~n678;
  assign n680 = n338 & n676;
  assign po41 = ~n679 & n680;
  assign n682 = ~pi26 & n338;
  assign n683 = pi27 & n651;
  assign n684 = pi95 & ~pi96;
  assign n685 = n640 & n684;
  assign n686 = ~n639 & ~n685;
  assign n687 = ~pi27 & ~pi100;
  assign n688 = ~n686 & n687;
  assign n689 = ~n683 & ~n688;
  assign n690 = n630 & n682;
  assign po42 = ~n689 & n690;
  assign n692 = ~pi26 & ~pi27;
  assign n693 = ~pi28 & ~pi116;
  assign n694 = pi100 & pi116;
  assign n695 = n692 & ~n693;
  assign n696 = ~n694 & n695;
  assign n697 = pi85 & ~n696;
  assign n698 = n649 & n677;
  assign n699 = ~pi26 & ~pi100;
  assign n700 = ~pi110 & n699;
  assign n701 = n684 & n700;
  assign n702 = ~n698 & ~n701;
  assign n703 = ~pi27 & ~n702;
  assign n704 = ~pi26 & ~n663;
  assign n705 = ~pi27 & n649;
  assign n706 = ~n704 & ~n705;
  assign n707 = ~n661 & ~n706;
  assign n708 = pi26 & pi27;
  assign n709 = ~n692 & ~n708;
  assign n710 = ~pi116 & n709;
  assign n711 = ~n707 & ~n710;
  assign n712 = pi28 & ~n711;
  assign n713 = ~pi26 & n664;
  assign n714 = pi116 & n713;
  assign n715 = ~pi85 & ~n703;
  assign n716 = ~n714 & n715;
  assign n717 = ~n712 & n716;
  assign n718 = ~pi53 & ~n697;
  assign n719 = ~n717 & n718;
  assign n720 = ~pi27 & pi28;
  assign n721 = ~pi116 & n720;
  assign n722 = pi53 & n668;
  assign n723 = n721 & n722;
  assign n724 = ~n719 & ~n723;
  assign n725 = ~pi58 & ~n724;
  assign n726 = ~pi26 & ~pi53;
  assign n727 = ~pi85 & n726;
  assign n728 = pi58 & n721;
  assign n729 = n727 & n728;
  assign n730 = ~n725 & ~n729;
  assign po43 = n338 & ~n730;
  assign n732 = ~pi96 & ~pi110;
  assign n733 = pi97 & ~n732;
  assign n734 = n659 & ~n733;
  assign n735 = pi97 & n734;
  assign n736 = ~pi110 & ~n734;
  assign n737 = pi29 & ~n736;
  assign n738 = ~pi58 & ~n735;
  assign n739 = ~n737 & n738;
  assign n740 = pi29 & ~pi116;
  assign n741 = pi97 & pi116;
  assign n742 = pi58 & ~n740;
  assign n743 = ~n741 & n742;
  assign n744 = ~pi53 & ~n743;
  assign n745 = ~n739 & n744;
  assign n746 = n637 & n740;
  assign n747 = ~n745 & ~n746;
  assign n748 = ~pi27 & ~n747;
  assign n749 = pi27 & n630;
  assign n750 = n740 & n749;
  assign n751 = ~n748 & ~n750;
  assign n752 = ~pi85 & ~n751;
  assign n753 = pi85 & n740;
  assign n754 = n676 & n753;
  assign n755 = ~n752 & ~n754;
  assign n756 = ~pi26 & ~n755;
  assign n757 = pi26 & ~pi27;
  assign n758 = ~pi85 & n630;
  assign n759 = n757 & n758;
  assign n760 = n740 & n759;
  assign n761 = ~n756 & ~n760;
  assign po44 = n338 & ~n761;
  assign n763 = ~pi88 & pi106;
  assign n764 = ~pi30 & ~pi109;
  assign n765 = ~pi60 & pi109;
  assign n766 = ~n764 & ~n765;
  assign n767 = ~pi106 & ~n766;
  assign n768 = ~pi129 & ~n763;
  assign po45 = ~n767 & n768;
  assign n770 = ~pi89 & pi106;
  assign n771 = ~pi31 & ~pi109;
  assign n772 = ~pi30 & pi109;
  assign n773 = ~n771 & ~n772;
  assign n774 = ~pi106 & ~n773;
  assign n775 = ~pi129 & ~n770;
  assign po46 = ~n774 & n775;
  assign n777 = ~pi99 & pi106;
  assign n778 = ~pi32 & ~pi109;
  assign n779 = ~pi31 & pi109;
  assign n780 = ~n778 & ~n779;
  assign n781 = ~pi106 & ~n780;
  assign n782 = ~pi129 & ~n777;
  assign po47 = ~n781 & n782;
  assign n784 = ~pi90 & pi106;
  assign n785 = ~pi33 & ~pi109;
  assign n786 = ~pi32 & pi109;
  assign n787 = ~n785 & ~n786;
  assign n788 = ~pi106 & ~n787;
  assign n789 = ~pi129 & ~n784;
  assign po48 = ~n788 & n789;
  assign n791 = ~pi91 & pi106;
  assign n792 = ~pi34 & ~pi109;
  assign n793 = ~pi33 & pi109;
  assign n794 = ~n792 & ~n793;
  assign n795 = ~pi106 & ~n794;
  assign n796 = ~pi129 & ~n791;
  assign po49 = ~n795 & n796;
  assign n798 = ~pi92 & pi106;
  assign n799 = ~pi35 & ~pi109;
  assign n800 = ~pi34 & pi109;
  assign n801 = ~n799 & ~n800;
  assign n802 = ~pi106 & ~n801;
  assign n803 = ~pi129 & ~n798;
  assign po50 = ~n802 & n803;
  assign n805 = ~pi98 & pi106;
  assign n806 = ~pi36 & ~pi109;
  assign n807 = ~pi35 & pi109;
  assign n808 = ~n806 & ~n807;
  assign n809 = ~pi106 & ~n808;
  assign n810 = ~pi129 & ~n805;
  assign po51 = ~n809 & n810;
  assign n812 = ~pi93 & pi106;
  assign n813 = ~pi37 & ~pi109;
  assign n814 = ~pi36 & pi109;
  assign n815 = ~n813 & ~n814;
  assign n816 = ~pi106 & ~n815;
  assign n817 = ~pi129 & ~n812;
  assign po52 = ~n816 & n817;
  assign n819 = ~pi40 & ~pi42;
  assign n820 = ~pi44 & pi82;
  assign n821 = pi38 & n819;
  assign n822 = n820 & n821;
  assign n823 = n518 & n611;
  assign n824 = ~pi48 & n823;
  assign n825 = n395 & n397;
  assign n826 = ~pi50 & n825;
  assign n827 = n824 & n826;
  assign n828 = n394 & n827;
  assign n829 = pi82 & ~n828;
  assign n830 = pi74 & ~n390;
  assign n831 = ~n829 & n830;
  assign n832 = pi82 & ~n394;
  assign n833 = n395 & n398;
  assign n834 = ~pi50 & n823;
  assign n835 = n833 & n834;
  assign n836 = pi82 & ~n835;
  assign n837 = n390 & ~n836;
  assign n838 = ~n832 & ~n837;
  assign n839 = ~pi38 & ~n838;
  assign n840 = ~pi129 & ~n822;
  assign n841 = ~n831 & n840;
  assign po53 = ~n839 & n841;
  assign n843 = pi109 & n662;
  assign n844 = pi39 & ~n843;
  assign n845 = ~pi51 & pi109;
  assign n846 = n648 & n845;
  assign n847 = ~pi106 & ~n846;
  assign n848 = ~n844 & n847;
  assign po54 = ~pi129 & ~n848;
  assign n850 = ~pi42 & n820;
  assign n851 = pi40 & n850;
  assign n852 = pi82 & ~n380;
  assign n853 = pi82 & ~n401;
  assign n854 = n390 & ~n853;
  assign n855 = ~n852 & ~n854;
  assign n856 = ~pi40 & ~n855;
  assign n857 = n523 & n823;
  assign n858 = n379 & n857;
  assign n859 = n382 & n858;
  assign n860 = n380 & n859;
  assign n861 = pi82 & ~n860;
  assign n862 = pi73 & ~n390;
  assign n863 = ~n861 & n862;
  assign n864 = ~pi129 & ~n851;
  assign n865 = ~n856 & n864;
  assign po55 = ~n863 & n865;
  assign n867 = pi41 & n850;
  assign n868 = n383 & n867;
  assign n869 = pi82 & ~n384;
  assign n870 = pi82 & ~n400;
  assign n871 = n390 & ~n870;
  assign n872 = ~n869 & ~n871;
  assign n873 = ~pi41 & ~n872;
  assign n874 = n400 & n576;
  assign n875 = pi82 & ~n874;
  assign n876 = pi76 & ~n390;
  assign n877 = ~n875 & n876;
  assign n878 = ~pi129 & ~n868;
  assign n879 = ~n873 & n878;
  assign po56 = ~n877 & n879;
  assign n881 = pi42 & n820;
  assign n882 = n819 & n859;
  assign n883 = ~n391 & ~n882;
  assign n884 = pi72 & ~n883;
  assign n885 = pi44 & pi82;
  assign n886 = ~pi40 & n859;
  assign n887 = pi82 & ~n886;
  assign n888 = n390 & ~n887;
  assign n889 = ~n885 & ~n888;
  assign n890 = ~pi42 & ~n889;
  assign n891 = ~pi129 & ~n881;
  assign n892 = ~n884 & n891;
  assign po57 = ~n890 & n892;
  assign n894 = n819 & n820;
  assign n895 = n396 & n894;
  assign n896 = pi43 & n895;
  assign n897 = pi82 & ~n519;
  assign n898 = n525 & n526;
  assign n899 = n524 & n898;
  assign n900 = pi82 & ~n899;
  assign n901 = n390 & ~n900;
  assign n902 = ~n897 & ~n901;
  assign n903 = ~pi43 & ~n902;
  assign n904 = n519 & n857;
  assign n905 = pi82 & ~n904;
  assign n906 = pi77 & ~n390;
  assign n907 = ~n905 & n906;
  assign n908 = ~pi129 & ~n896;
  assign n909 = ~n907 & n908;
  assign po58 = ~n903 & n909;
  assign n911 = pi82 & ~n882;
  assign n912 = ~pi67 & ~n390;
  assign n913 = pi44 & n390;
  assign n914 = ~n912 & ~n913;
  assign n915 = ~n911 & n914;
  assign n916 = ~pi129 & ~n885;
  assign po59 = ~n915 & n916;
  assign n918 = n575 & n833;
  assign n919 = pi45 & pi82;
  assign n920 = n918 & n919;
  assign n921 = pi82 & ~n898;
  assign n922 = n390 & ~n921;
  assign n923 = pi82 & ~n918;
  assign n924 = ~n922 & ~n923;
  assign n925 = ~pi45 & ~n924;
  assign n926 = n387 & n898;
  assign n927 = pi82 & ~n926;
  assign n928 = pi68 & ~n390;
  assign n929 = ~n927 & n928;
  assign n930 = ~pi129 & ~n920;
  assign n931 = ~n925 & n930;
  assign po60 = ~n929 & n931;
  assign n933 = ~pi75 & n391;
  assign n934 = ~pi75 & ~n390;
  assign n935 = pi82 & ~n858;
  assign n936 = ~n934 & ~n935;
  assign n937 = n576 & ~n936;
  assign n938 = pi82 & n575;
  assign n939 = pi46 & ~n391;
  assign n940 = ~n938 & n939;
  assign n941 = ~n933 & ~n940;
  assign n942 = ~n937 & n941;
  assign po61 = ~pi129 & ~n942;
  assign n944 = ~pi43 & pi47;
  assign n945 = n895 & n944;
  assign n946 = pi82 & ~n385;
  assign n947 = pi82 & ~n824;
  assign n948 = n390 & ~n947;
  assign n949 = ~n946 & ~n948;
  assign n950 = ~pi47 & ~n949;
  assign n951 = n385 & n824;
  assign n952 = pi82 & ~n951;
  assign n953 = pi64 & ~n390;
  assign n954 = ~n952 & n953;
  assign n955 = ~pi129 & ~n945;
  assign n956 = ~n950 & n955;
  assign po62 = ~n954 & n956;
  assign n958 = pi48 & n397;
  assign n959 = n895 & n958;
  assign n960 = pi82 & ~n823;
  assign n961 = n390 & ~n960;
  assign n962 = n575 & n825;
  assign n963 = pi82 & ~n962;
  assign n964 = ~n961 & ~n963;
  assign n965 = ~pi48 & ~n964;
  assign n966 = n386 & n823;
  assign n967 = pi82 & ~n966;
  assign n968 = pi62 & ~n390;
  assign n969 = ~n967 & n968;
  assign n970 = ~pi129 & ~n959;
  assign n971 = ~n965 & n970;
  assign po63 = ~n969 & n971;
  assign n973 = ~pi24 & ~pi40;
  assign n974 = n380 & n973;
  assign n975 = n382 & n974;
  assign n976 = n573 & n975;
  assign n977 = pi49 & ~n976;
  assign n978 = n578 & ~n611;
  assign n979 = ~n977 & ~n978;
  assign n980 = pi82 & ~n979;
  assign n981 = pi49 & n516;
  assign n982 = pi82 & ~n578;
  assign n983 = ~pi69 & ~n390;
  assign n984 = ~n982 & n983;
  assign n985 = ~n981 & ~n984;
  assign n986 = ~n980 & n985;
  assign po64 = ~pi129 & ~n986;
  assign n988 = pi50 & pi82;
  assign n989 = n574 & n988;
  assign n990 = pi82 & ~n574;
  assign n991 = n395 & n400;
  assign n992 = pi82 & ~n991;
  assign n993 = n390 & ~n992;
  assign n994 = ~n990 & ~n993;
  assign n995 = ~pi50 & ~n994;
  assign n996 = pi82 & ~n827;
  assign n997 = pi66 & ~n390;
  assign n998 = ~n996 & n997;
  assign n999 = ~pi129 & ~n989;
  assign n1000 = ~n998 & n999;
  assign po65 = ~n995 & n1000;
  assign n1002 = pi51 & ~pi109;
  assign n1003 = ~pi106 & ~n845;
  assign n1004 = ~n1002 & n1003;
  assign po66 = ~pi129 & ~n1004;
  assign n1006 = pi52 & ~n845;
  assign n1007 = ~pi106 & ~n843;
  assign n1008 = ~n1006 & n1007;
  assign po67 = ~pi129 & ~n1008;
  assign n1010 = ~pi116 & n637;
  assign n1011 = pi58 & pi116;
  assign n1012 = ~pi58 & n659;
  assign n1013 = n732 & n1012;
  assign n1014 = ~n1011 & ~n1013;
  assign n1015 = ~pi53 & pi97;
  assign n1016 = ~n1014 & n1015;
  assign n1017 = ~n1010 & ~n1016;
  assign n1018 = n632 & n682;
  assign po68 = ~n1017 & n1018;
  assign n1020 = ~n390 & n898;
  assign n1021 = n615 & n1020;
  assign n1022 = ~pi129 & ~n391;
  assign po69 = n1021 | ~n1022;
  assign po129 = pi123 | pi129;
  assign n1025 = pi114 & ~pi122;
  assign po70 = ~po129 & n1025;
  assign n1027 = ~pi26 & pi58;
  assign n1028 = ~pi58 & n677;
  assign n1029 = ~n1027 & ~n1028;
  assign n1030 = pi94 & ~n1029;
  assign n1031 = pi58 & ~pi116;
  assign n1032 = pi37 & ~pi116;
  assign n1033 = ~n1027 & ~n1032;
  assign n1034 = ~n1031 & ~n1033;
  assign n1035 = ~n1030 & ~n1034;
  assign n1036 = ~pi53 & ~n1035;
  assign n1037 = ~pi26 & pi37;
  assign n1038 = ~pi58 & n1037;
  assign n1039 = ~n1036 & ~n1038;
  assign n1040 = ~pi85 & ~n1039;
  assign n1041 = n630 & n1037;
  assign n1042 = ~n1040 & ~n1041;
  assign n1043 = ~pi27 & ~n1042;
  assign n1044 = n758 & n1037;
  assign n1045 = ~n1043 & ~n1044;
  assign po71 = n338 & ~n1045;
  assign n1047 = ~pi116 & n727;
  assign n1048 = pi85 & ~n726;
  assign n1049 = pi26 & pi53;
  assign n1050 = ~pi58 & ~n1049;
  assign n1051 = ~n1048 & n1050;
  assign n1052 = ~n1047 & ~n1051;
  assign n1053 = pi57 & ~n1052;
  assign n1054 = pi60 & n1011;
  assign n1055 = n727 & n1054;
  assign n1056 = ~n1053 & ~n1055;
  assign n1057 = ~pi27 & ~n1056;
  assign n1058 = pi57 & ~pi58;
  assign n1059 = n727 & n1058;
  assign n1060 = ~n1057 & ~n1059;
  assign po72 = n338 & ~n1060;
  assign n1062 = n692 & n1031;
  assign n1063 = ~pi58 & n709;
  assign n1064 = n650 & n1063;
  assign n1065 = ~n1062 & ~n1064;
  assign n1066 = ~pi53 & ~pi85;
  assign n1067 = n338 & n1066;
  assign po73 = ~n1065 & n1067;
  assign n1069 = ~pi59 & ~n661;
  assign n1070 = ~pi96 & n661;
  assign n1071 = n630 & ~n1069;
  assign n1072 = ~n1070 & n1071;
  assign n1073 = pi59 & ~pi116;
  assign n1074 = ~n638 & n1073;
  assign n1075 = ~n1072 & ~n1074;
  assign n1076 = ~pi85 & ~n1075;
  assign n1077 = pi85 & n630;
  assign n1078 = n1073 & n1077;
  assign n1079 = ~n1076 & ~n1078;
  assign n1080 = ~pi27 & ~n1079;
  assign n1081 = pi27 & n1073;
  assign n1082 = n758 & n1081;
  assign n1083 = ~n1080 & ~n1082;
  assign n1084 = ~pi26 & ~n1083;
  assign n1085 = n759 & n1073;
  assign n1086 = ~n1084 & ~n1085;
  assign po74 = n338 & ~n1086;
  assign n1088 = ~pi117 & ~pi122;
  assign n1089 = pi60 & ~n1088;
  assign n1090 = pi123 & n1088;
  assign po75 = n1089 | n1090;
  assign n1092 = ~pi114 & ~pi122;
  assign n1093 = pi123 & ~pi129;
  assign po76 = n1092 & n1093;
  assign n1095 = pi136 & ~pi137;
  assign n1096 = pi131 & pi132;
  assign n1097 = pi133 & n1096;
  assign n1098 = ~pi138 & n1097;
  assign n1099 = n1095 & n1098;
  assign n1100 = ~pi62 & ~n1099;
  assign n1101 = pi140 & n1099;
  assign n1102 = ~pi129 & ~n1100;
  assign po77 = n1101 | ~n1102;
  assign n1104 = ~pi63 & ~n1099;
  assign n1105 = pi142 & n1099;
  assign n1106 = ~pi129 & ~n1104;
  assign po78 = n1105 | ~n1106;
  assign n1108 = ~pi64 & ~n1099;
  assign n1109 = pi139 & n1099;
  assign n1110 = ~pi129 & ~n1108;
  assign po79 = n1109 | ~n1110;
  assign n1112 = ~pi65 & ~n1099;
  assign n1113 = pi146 & n1099;
  assign n1114 = ~pi129 & ~n1112;
  assign po80 = n1113 | ~n1114;
  assign n1116 = ~pi136 & ~pi137;
  assign n1117 = n1098 & n1116;
  assign n1118 = ~pi66 & ~n1117;
  assign n1119 = pi143 & n1117;
  assign n1120 = ~pi129 & ~n1118;
  assign po81 = n1119 | ~n1120;
  assign n1122 = ~pi67 & ~n1117;
  assign n1123 = pi139 & n1117;
  assign n1124 = ~pi129 & ~n1122;
  assign po82 = n1123 | ~n1124;
  assign n1126 = ~pi68 & ~n1099;
  assign n1127 = pi141 & n1099;
  assign n1128 = ~pi129 & ~n1126;
  assign po83 = n1127 | ~n1128;
  assign n1130 = ~pi69 & ~n1099;
  assign n1131 = pi143 & n1099;
  assign n1132 = ~pi129 & ~n1130;
  assign po84 = n1131 | ~n1132;
  assign n1134 = ~pi70 & ~n1099;
  assign n1135 = pi144 & n1099;
  assign n1136 = ~pi129 & ~n1134;
  assign po85 = n1135 | ~n1136;
  assign n1138 = ~pi71 & ~n1099;
  assign n1139 = pi145 & n1099;
  assign n1140 = ~pi129 & ~n1138;
  assign po86 = n1139 | ~n1140;
  assign n1142 = ~pi72 & ~n1117;
  assign n1143 = pi140 & n1117;
  assign n1144 = ~pi129 & ~n1142;
  assign po87 = n1143 | ~n1144;
  assign n1146 = ~pi73 & ~n1117;
  assign n1147 = pi141 & n1117;
  assign n1148 = ~pi129 & ~n1146;
  assign po88 = n1147 | ~n1148;
  assign n1150 = ~pi74 & ~n1117;
  assign n1151 = pi142 & n1117;
  assign n1152 = ~pi129 & ~n1150;
  assign po89 = n1151 | ~n1152;
  assign n1154 = ~pi75 & ~n1117;
  assign n1155 = pi144 & n1117;
  assign n1156 = ~pi129 & ~n1154;
  assign po90 = n1155 | ~n1156;
  assign n1158 = ~pi76 & ~n1117;
  assign n1159 = pi145 & n1117;
  assign n1160 = ~pi129 & ~n1158;
  assign po91 = n1159 | ~n1160;
  assign n1162 = ~pi77 & ~n1117;
  assign n1163 = pi146 & n1117;
  assign n1164 = ~pi129 & ~n1162;
  assign po92 = n1163 | ~n1164;
  assign n1166 = ~pi136 & pi137;
  assign n1167 = n1098 & n1166;
  assign n1168 = ~pi78 & ~n1167;
  assign n1169 = ~pi142 & n1167;
  assign n1170 = ~pi129 & ~n1168;
  assign po93 = ~n1169 & n1170;
  assign n1172 = ~pi79 & ~n1167;
  assign n1173 = ~pi143 & n1167;
  assign n1174 = ~pi129 & ~n1172;
  assign po94 = ~n1173 & n1174;
  assign n1176 = ~pi80 & ~n1167;
  assign n1177 = ~pi144 & n1167;
  assign n1178 = ~pi129 & ~n1176;
  assign po95 = ~n1177 & n1178;
  assign n1180 = ~pi81 & ~n1167;
  assign n1181 = ~pi145 & n1167;
  assign n1182 = ~pi129 & ~n1180;
  assign po96 = ~n1181 & n1182;
  assign n1184 = ~pi82 & ~n1167;
  assign n1185 = ~pi146 & n1167;
  assign n1186 = ~pi129 & ~n1184;
  assign po97 = ~n1185 & n1186;
  assign n1188 = pi136 & ~pi138;
  assign n1189 = pi31 & n1188;
  assign n1190 = ~pi87 & ~pi138;
  assign n1191 = pi115 & pi138;
  assign n1192 = ~pi136 & ~n1190;
  assign n1193 = ~n1191 & n1192;
  assign n1194 = ~n1189 & ~n1193;
  assign n1195 = pi137 & ~n1194;
  assign n1196 = ~pi89 & pi138;
  assign n1197 = pi62 & ~pi138;
  assign n1198 = pi136 & ~n1196;
  assign n1199 = ~n1197 & n1198;
  assign n1200 = ~pi119 & pi138;
  assign n1201 = pi72 & ~pi138;
  assign n1202 = ~pi136 & ~n1200;
  assign n1203 = ~n1201 & n1202;
  assign n1204 = ~n1199 & ~n1203;
  assign n1205 = ~pi137 & ~n1204;
  assign po98 = n1195 | n1205;
  assign n1207 = ~pi84 & ~n1167;
  assign n1208 = ~pi141 & n1167;
  assign n1209 = ~pi129 & ~n1207;
  assign po99 = ~n1208 & n1209;
  assign n1211 = n640 & ~n660;
  assign n1212 = pi96 & n1211;
  assign n1213 = ~n644 & ~n1212;
  assign n1214 = n676 & n682;
  assign po100 = ~n1213 & n1214;
  assign n1216 = ~pi86 & ~n1167;
  assign n1217 = ~pi139 & n1167;
  assign n1218 = ~pi129 & ~n1216;
  assign po101 = ~n1217 & n1218;
  assign n1220 = ~pi87 & ~n1167;
  assign n1221 = ~pi140 & n1167;
  assign n1222 = ~pi129 & ~n1220;
  assign po102 = ~n1221 & n1222;
  assign n1224 = pi137 & n1188;
  assign n1225 = n1097 & n1224;
  assign n1226 = ~pi88 & ~n1225;
  assign n1227 = ~pi139 & n1225;
  assign n1228 = ~pi129 & ~n1226;
  assign po103 = ~n1227 & n1228;
  assign n1230 = ~pi89 & ~n1225;
  assign n1231 = ~pi140 & n1225;
  assign n1232 = ~pi129 & ~n1230;
  assign po104 = ~n1231 & n1232;
  assign n1234 = ~pi90 & ~n1225;
  assign n1235 = ~pi142 & n1225;
  assign n1236 = ~pi129 & ~n1234;
  assign po105 = ~n1235 & n1236;
  assign n1238 = ~pi91 & ~n1225;
  assign n1239 = ~pi143 & n1225;
  assign n1240 = ~pi129 & ~n1238;
  assign po106 = ~n1239 & n1240;
  assign n1242 = ~pi92 & ~n1225;
  assign n1243 = ~pi144 & n1225;
  assign n1244 = ~pi129 & ~n1242;
  assign po107 = ~n1243 & n1244;
  assign n1246 = ~pi93 & ~n1225;
  assign n1247 = ~pi146 & n1225;
  assign n1248 = ~pi129 & ~n1246;
  assign po108 = ~n1247 & n1248;
  assign n1250 = pi82 & pi138;
  assign n1251 = n1116 & n1250;
  assign n1252 = n1097 & n1251;
  assign n1253 = ~pi94 & ~n1252;
  assign n1254 = ~pi142 & n1252;
  assign n1255 = ~pi129 & ~n1253;
  assign po109 = ~n1254 & n1255;
  assign n1257 = ~pi3 & ~pi110;
  assign n1258 = ~n1097 & ~n1257;
  assign n1259 = ~n1252 & ~n1258;
  assign n1260 = pi95 & n1259;
  assign n1261 = pi143 & n1252;
  assign n1262 = ~n1260 & ~n1261;
  assign po110 = ~pi129 & ~n1262;
  assign n1264 = pi96 & n1259;
  assign n1265 = pi146 & n1252;
  assign n1266 = ~n1264 & ~n1265;
  assign po111 = ~pi129 & ~n1266;
  assign n1268 = pi97 & n1259;
  assign n1269 = pi145 & n1252;
  assign n1270 = ~n1268 & ~n1269;
  assign po112 = ~pi129 & ~n1270;
  assign n1272 = ~pi98 & ~n1225;
  assign n1273 = ~pi145 & n1225;
  assign n1274 = ~pi129 & ~n1272;
  assign po113 = ~n1273 & n1274;
  assign n1276 = ~pi99 & ~n1225;
  assign n1277 = ~pi141 & n1225;
  assign n1278 = ~pi129 & ~n1276;
  assign po114 = ~n1277 & n1278;
  assign n1280 = pi100 & n1259;
  assign n1281 = pi144 & n1252;
  assign n1282 = ~n1280 & ~n1281;
  assign po115 = ~pi129 & ~n1282;
  assign n1284 = pi37 & n1188;
  assign n1285 = ~pi82 & ~pi138;
  assign n1286 = ~pi96 & pi138;
  assign n1287 = ~pi136 & ~n1285;
  assign n1288 = ~n1286 & n1287;
  assign n1289 = ~n1284 & ~n1288;
  assign n1290 = pi137 & ~n1289;
  assign n1291 = ~pi93 & pi138;
  assign n1292 = pi65 & ~pi138;
  assign n1293 = pi136 & ~n1291;
  assign n1294 = ~n1292 & n1293;
  assign n1295 = ~pi124 & pi138;
  assign n1296 = pi77 & ~pi138;
  assign n1297 = ~pi136 & ~n1295;
  assign n1298 = ~n1296 & n1297;
  assign n1299 = ~n1294 & ~n1298;
  assign n1300 = ~pi137 & ~n1299;
  assign po116 = n1290 | n1300;
  assign n1302 = pi91 & n1095;
  assign n1303 = pi95 & n1166;
  assign n1304 = ~n1302 & ~n1303;
  assign n1305 = pi138 & ~n1304;
  assign n1306 = ~pi79 & ~pi136;
  assign n1307 = ~pi34 & pi136;
  assign n1308 = pi137 & ~n1306;
  assign n1309 = ~n1307 & n1308;
  assign n1310 = pi66 & ~pi136;
  assign n1311 = pi69 & pi136;
  assign n1312 = ~pi137 & ~n1310;
  assign n1313 = ~n1311 & n1312;
  assign n1314 = ~n1309 & ~n1313;
  assign n1315 = ~pi138 & ~n1314;
  assign po117 = n1305 | n1315;
  assign n1317 = pi90 & n1095;
  assign n1318 = pi94 & n1166;
  assign n1319 = ~n1317 & ~n1318;
  assign n1320 = pi138 & ~n1319;
  assign n1321 = ~pi78 & ~pi136;
  assign n1322 = ~pi33 & pi136;
  assign n1323 = pi137 & ~n1321;
  assign n1324 = ~n1322 & n1323;
  assign n1325 = pi74 & ~pi136;
  assign n1326 = pi63 & pi136;
  assign n1327 = ~pi137 & ~n1325;
  assign n1328 = ~n1326 & n1327;
  assign n1329 = ~n1324 & ~n1328;
  assign n1330 = ~pi138 & ~n1329;
  assign po118 = n1320 | n1330;
  assign n1332 = pi99 & n1095;
  assign n1333 = ~pi112 & n1166;
  assign n1334 = ~n1332 & ~n1333;
  assign n1335 = pi138 & ~n1334;
  assign n1336 = ~pi84 & ~pi136;
  assign n1337 = ~pi32 & pi136;
  assign n1338 = pi137 & ~n1336;
  assign n1339 = ~n1337 & n1338;
  assign n1340 = pi73 & ~pi136;
  assign n1341 = pi68 & pi136;
  assign n1342 = ~pi137 & ~n1340;
  assign n1343 = ~n1341 & n1342;
  assign n1344 = ~n1339 & ~n1343;
  assign n1345 = ~pi138 & ~n1344;
  assign po119 = n1335 | n1345;
  assign n1347 = pi35 & n1188;
  assign n1348 = ~pi80 & ~pi138;
  assign n1349 = ~pi100 & pi138;
  assign n1350 = ~pi136 & ~n1348;
  assign n1351 = ~n1349 & n1350;
  assign n1352 = ~n1347 & ~n1351;
  assign n1353 = pi137 & ~n1352;
  assign n1354 = ~pi92 & pi138;
  assign n1355 = pi70 & ~pi138;
  assign n1356 = pi136 & ~n1354;
  assign n1357 = ~n1355 & n1356;
  assign n1358 = ~pi125 & pi138;
  assign n1359 = pi75 & ~pi138;
  assign n1360 = ~pi136 & ~n1358;
  assign n1361 = ~n1359 & n1360;
  assign n1362 = ~n1357 & ~n1361;
  assign n1363 = ~pi137 & ~n1362;
  assign po120 = n1353 | n1363;
  assign n1365 = ~pi26 & n676;
  assign n1366 = n1211 & n1365;
  assign n1367 = ~n639 & ~n1366;
  assign po121 = n338 & ~n1367;
  assign n1369 = pi36 & n1188;
  assign n1370 = ~pi81 & ~pi138;
  assign n1371 = ~pi97 & pi138;
  assign n1372 = ~pi136 & ~n1370;
  assign n1373 = ~n1371 & n1372;
  assign n1374 = ~n1369 & ~n1373;
  assign n1375 = pi137 & ~n1374;
  assign n1376 = ~pi98 & pi138;
  assign n1377 = pi71 & ~pi138;
  assign n1378 = pi136 & ~n1376;
  assign n1379 = ~n1377 & n1378;
  assign n1380 = ~pi23 & pi138;
  assign n1381 = pi76 & ~pi138;
  assign n1382 = ~pi136 & ~n1380;
  assign n1383 = ~n1381 & n1382;
  assign n1384 = ~n1379 & ~n1383;
  assign n1385 = ~pi137 & ~n1384;
  assign po122 = n1375 | n1385;
  assign n1387 = pi30 & n1188;
  assign n1388 = ~pi86 & ~pi138;
  assign n1389 = ~pi111 & pi138;
  assign n1390 = ~pi136 & ~n1388;
  assign n1391 = ~n1389 & n1390;
  assign n1392 = ~n1387 & ~n1391;
  assign n1393 = pi137 & ~n1392;
  assign n1394 = ~pi88 & pi138;
  assign n1395 = pi64 & ~pi138;
  assign n1396 = pi136 & ~n1394;
  assign n1397 = ~n1395 & n1396;
  assign n1398 = ~pi120 & pi138;
  assign n1399 = pi67 & ~pi138;
  assign n1400 = ~pi136 & ~n1398;
  assign n1401 = ~n1399 & n1400;
  assign n1402 = ~n1397 & ~n1401;
  assign n1403 = ~pi137 & ~n1402;
  assign po123 = n1393 | n1403;
  assign n1405 = ~n713 & ~n757;
  assign n1406 = pi116 & n338;
  assign po124 = ~n1405 & n1406;
  assign n1408 = ~pi97 & n636;
  assign n1409 = ~n637 & ~n1408;
  assign po125 = n1406 & ~n1409;
  assign n1411 = ~pi129 & n1097;
  assign n1412 = ~pi111 & ~n1251;
  assign n1413 = ~pi139 & n1251;
  assign n1414 = n1411 & ~n1412;
  assign po126 = ~n1413 & n1414;
  assign n1416 = ~pi141 & n1251;
  assign n1417 = pi112 & ~n1251;
  assign n1418 = n1411 & ~n1416;
  assign po127 = ~n1417 & n1418;
  assign n1420 = ~pi54 & pi113;
  assign n1421 = ~pi11 & ~pi22;
  assign n1422 = pi54 & n1421;
  assign n1423 = n338 & ~n1420;
  assign po128 = ~n1422 & n1423;
  assign n1425 = ~pi140 & n1251;
  assign n1426 = pi115 & ~n1251;
  assign n1427 = n1411 & ~n1425;
  assign po130 = ~n1426 & n1427;
  assign n1429 = ~pi4 & ~pi9;
  assign n1430 = n354 & n1429;
  assign n1431 = pi54 & n338;
  assign po131 = ~n1430 & n1431;
  assign po132 = ~pi122 | pi129;
  assign n1434 = ~pi54 & pi118;
  assign n1435 = pi54 & ~pi59;
  assign n1436 = n501 & n1435;
  assign n1437 = ~n1434 & ~n1436;
  assign po133 = ~pi129 & ~n1437;
  assign po134 = ~pi129 & ~n659;
  assign n1440 = ~pi120 & n1257;
  assign n1441 = ~pi111 & ~pi129;
  assign po135 = ~n1440 & n1441;
  assign n1443 = pi81 & pi120;
  assign po136 = ~pi129 & n1443;
  assign po137 = pi129 | pi134;
  assign po138 = pi129 | pi135;
  assign po139 = pi57 & ~pi129;
  assign n1448 = ~pi96 & pi125;
  assign n1449 = ~pi3 & ~n1448;
  assign po140 = ~pi129 & ~n1449;
  assign n1451 = ~pi126 & pi132;
  assign po141 = pi133 & n1451;
  assign po12 = 1'b1;
  assign po0 = pi108;
  assign po1 = pi83;
  assign po2 = pi104;
  assign po3 = pi103;
  assign po4 = pi102;
  assign po5 = pi105;
  assign po6 = pi107;
  assign po7 = pi101;
  assign po8 = pi126;
  assign po9 = pi121;
  assign po10 = pi1;
  assign po11 = pi0;
  assign po13 = pi130;
  assign po14 = pi128;
endmodule
