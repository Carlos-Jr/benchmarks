module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 , pi32 ,
    pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 , pi40 ,
    pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 , pi56 ,
    pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 , pi64 ,
    pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 ,
    pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 ,
    pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 ,
    pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 ,
    pi97 , pi98 , pi99 , pi100 , pi101 , pi102 , pi103 ,
    pi104 , pi105 , pi106 , pi107 , pi108 , pi109 , pi110 ,
    pi111 , pi112 , pi113 , pi114 , pi115 , pi116 , pi117 ,
    pi118 , pi119 , pi120 , pi121 , pi122 , pi123 , pi124 ,
    pi125 , pi126 , pi127 ,
    po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7  );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    pi32 , pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 ,
    pi56 , pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 ,
    pi64 , pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 ,
    pi72 , pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 ,
    pi80 , pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 ,
    pi88 , pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 ,
    pi96 , pi97 , pi98 , pi99 , pi100 , pi101 , pi102 ,
    pi103 , pi104 , pi105 , pi106 , pi107 , pi108 , pi109 ,
    pi110 , pi111 , pi112 , pi113 , pi114 , pi115 , pi116 ,
    pi117 , pi118 , pi119 , pi120 , pi121 , pi122 , pi123 ,
    pi124 , pi125 , pi126 , pi127 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7;
  wire n137, n138, n139, n140, n141, n142, n143,
    n144, n145, n146, n147, n148, n149, n150,
    n151, n152, n153, n154, n155, n156, n157,
    n158, n159, n160, n161, n162, n163, n164,
    n165, n166, n167, n168, n169, n170, n171,
    n172, n173, n174, n175, n176, n177, n178,
    n179, n180, n181, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192,
    n193, n194, n195, n196, n197, n198, n199,
    n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213,
    n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227,
    n228, n229, n230, n231, n232, n233, n234,
    n235, n236, n237, n238, n239, n240, n241,
    n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339,
    n340, n341, n342, n343, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403,
    n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416, n417,
    n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438,
    n439, n440, n441, n442, n443, n444, n445,
    n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487,
    n488, n489, n490, n491, n492, n493, n495,
    n496, n497, n498, n499, n500, n501, n502,
    n503, n504, n505, n506, n507, n508, n509,
    n510, n511, n512, n513, n514, n515, n516,
    n517, n518, n519, n520, n521, n522, n523,
    n524, n525, n526, n527, n528, n529, n530,
    n531, n532, n533, n534, n535, n536, n537,
    n538, n539, n540, n541, n542, n543, n544,
    n545, n546, n547, n548, n550, n551, n552,
    n553, n554, n555, n556, n557, n558, n559,
    n560, n561, n562, n563, n564, n565, n566,
    n568, n569, n570, n571, n572, n573, n574,
    n575, n576, n577, n578, n579, n580, n581,
    n582, n583, n584, n585, n586, n587, n588,
    n590, n591, n592, n593, n594, n595, n596,
    n597, n599, n600, n602, n603, n604, n605,
    n606, n607;
  assign n137 = ~pi124  & ~pi125 ;
  assign n138 = ~pi126  & ~pi127 ;
  assign n139 = n137 & n138;
  assign n140 = pi121  & ~pi122 ;
  assign n141 = ~pi123  & ~n140;
  assign n142 = n139 & ~n141;
  assign n143 = pi125  & ~pi126 ;
  assign n144 = ~pi127  & ~n143;
  assign n145 = ~n142 & n144;
  assign n146 = ~pi122  & ~pi123 ;
  assign n147 = ~pi120  & ~pi121 ;
  assign n148 = n146 & n147;
  assign n149 = n139 & n148;
  assign n150 = n145 & ~n149;
  assign n151 = ~pi118  & ~n150;
  assign n152 = ~pi116  & n151;
  assign n153 = pi117  & n151;
  assign n154 = pi119  & n149;
  assign n155 = n145 & ~n154;
  assign n156 = ~n153 & n155;
  assign n157 = ~n152 & n156;
  assign n158 = ~pi114  & ~n157;
  assign n159 = pi113  & n158;
  assign n160 = pi115  & n152;
  assign n161 = n156 & ~n160;
  assign n162 = ~n159 & n161;
  assign n163 = ~pi112  & n158;
  assign n164 = n162 & ~n163;
  assign n165 = ~pi110  & ~n164;
  assign n166 = ~pi108  & n165;
  assign n167 = pi109  & n165;
  assign n168 = pi111  & n163;
  assign n169 = n162 & ~n168;
  assign n170 = ~n167 & n169;
  assign n171 = ~n166 & n170;
  assign n172 = ~pi106  & ~n171;
  assign n173 = pi105  & n172;
  assign n174 = pi107  & n166;
  assign n175 = n170 & ~n174;
  assign n176 = ~n173 & n175;
  assign n177 = ~pi104  & n172;
  assign n178 = n176 & ~n177;
  assign n179 = ~pi102  & ~n178;
  assign n180 = ~pi100  & n179;
  assign n181 = pi101  & n179;
  assign n182 = pi103  & n177;
  assign n183 = n176 & ~n182;
  assign n184 = ~n181 & n183;
  assign n185 = ~n180 & n184;
  assign n186 = ~pi98  & ~n185;
  assign n187 = pi97  & n186;
  assign n188 = pi99  & n180;
  assign n189 = n184 & ~n188;
  assign n190 = ~n187 & n189;
  assign n191 = ~pi96  & n186;
  assign n192 = n190 & ~n191;
  assign n193 = ~pi94  & ~n192;
  assign n194 = ~pi92  & n193;
  assign n195 = pi93  & n193;
  assign n196 = pi95  & n191;
  assign n197 = n190 & ~n196;
  assign n198 = ~n195 & n197;
  assign n199 = ~n194 & n198;
  assign n200 = ~pi90  & ~n199;
  assign n201 = pi89  & n200;
  assign n202 = pi91  & n194;
  assign n203 = n198 & ~n202;
  assign n204 = ~n201 & n203;
  assign n205 = ~pi88  & n200;
  assign n206 = n204 & ~n205;
  assign n207 = ~pi86  & ~n206;
  assign n208 = ~pi84  & n207;
  assign n209 = pi85  & n207;
  assign n210 = pi87  & n205;
  assign n211 = n204 & ~n210;
  assign n212 = ~n209 & n211;
  assign n213 = ~n208 & n212;
  assign n214 = ~pi82  & ~n213;
  assign n215 = pi81  & n214;
  assign n216 = pi83  & n208;
  assign n217 = n212 & ~n216;
  assign n218 = ~n215 & n217;
  assign n219 = ~pi80  & n214;
  assign n220 = n218 & ~n219;
  assign n221 = ~pi78  & ~n220;
  assign n222 = ~pi76  & n221;
  assign n223 = pi77  & n221;
  assign n224 = pi79  & n219;
  assign n225 = n218 & ~n224;
  assign n226 = ~n223 & n225;
  assign n227 = ~n222 & n226;
  assign n228 = ~pi74  & ~n227;
  assign n229 = pi73  & n228;
  assign n230 = pi75  & n222;
  assign n231 = n226 & ~n230;
  assign n232 = ~n229 & n231;
  assign n233 = ~pi72  & n228;
  assign n234 = n232 & ~n233;
  assign n235 = ~pi70  & ~n234;
  assign n236 = ~pi68  & n235;
  assign n237 = pi69  & n235;
  assign n238 = pi71  & n233;
  assign n239 = n232 & ~n238;
  assign n240 = ~n237 & n239;
  assign n241 = ~n236 & n240;
  assign n242 = ~pi66  & ~n241;
  assign n243 = pi65  & n242;
  assign n244 = pi67  & n236;
  assign n245 = n240 & ~n244;
  assign n246 = ~n243 & n245;
  assign n247 = ~pi64  & n242;
  assign n248 = n246 & ~n247;
  assign n249 = ~pi62  & ~n248;
  assign n250 = ~pi60  & n249;
  assign n251 = pi61  & n249;
  assign n252 = pi63  & n247;
  assign n253 = n246 & ~n252;
  assign n254 = ~n251 & n253;
  assign n255 = ~n250 & n254;
  assign n256 = ~pi58  & ~n255;
  assign n257 = pi57  & n256;
  assign n258 = pi59  & n250;
  assign n259 = n254 & ~n258;
  assign n260 = ~n257 & n259;
  assign n261 = ~pi56  & n256;
  assign n262 = n260 & ~n261;
  assign n263 = ~pi54  & ~n262;
  assign n264 = ~pi52  & n263;
  assign n265 = pi53  & n263;
  assign n266 = pi55  & n261;
  assign n267 = n260 & ~n266;
  assign n268 = ~n265 & n267;
  assign n269 = ~n264 & n268;
  assign n270 = ~pi50  & ~n269;
  assign n271 = pi49  & n270;
  assign n272 = pi51  & n264;
  assign n273 = n268 & ~n272;
  assign n274 = ~n271 & n273;
  assign n275 = ~pi48  & n270;
  assign n276 = n274 & ~n275;
  assign n277 = ~pi46  & ~n276;
  assign n278 = ~pi44  & n277;
  assign n279 = pi45  & n277;
  assign n280 = pi47  & n275;
  assign n281 = n274 & ~n280;
  assign n282 = ~n279 & n281;
  assign n283 = ~n278 & n282;
  assign n284 = ~pi42  & ~n283;
  assign n285 = pi41  & n284;
  assign n286 = pi43  & n278;
  assign n287 = n282 & ~n286;
  assign n288 = ~n285 & n287;
  assign n289 = ~pi40  & n284;
  assign n290 = n288 & ~n289;
  assign n291 = ~pi38  & ~n290;
  assign n292 = ~pi36  & n291;
  assign n293 = pi37  & n291;
  assign n294 = pi39  & n289;
  assign n295 = n288 & ~n294;
  assign n296 = ~n293 & n295;
  assign n297 = ~n292 & n296;
  assign n298 = ~pi34  & ~n297;
  assign n299 = pi33  & n298;
  assign n300 = pi35  & n292;
  assign n301 = n296 & ~n300;
  assign n302 = ~n299 & n301;
  assign n303 = ~pi32  & n298;
  assign n304 = n302 & ~n303;
  assign n305 = ~pi30  & ~n304;
  assign n306 = ~pi28  & n305;
  assign n307 = pi29  & n305;
  assign n308 = pi31  & n303;
  assign n309 = n302 & ~n308;
  assign n310 = ~n307 & n309;
  assign n311 = ~n306 & n310;
  assign n312 = ~pi26  & ~n311;
  assign n313 = pi25  & n312;
  assign n314 = pi27  & n306;
  assign n315 = n310 & ~n314;
  assign n316 = ~n313 & n315;
  assign n317 = ~pi24  & n312;
  assign n318 = n316 & ~n317;
  assign n319 = ~pi22  & ~n318;
  assign n320 = pi21  & n319;
  assign n321 = pi23  & n317;
  assign n322 = pi1  & ~pi2 ;
  assign n323 = ~pi3  & ~n322;
  assign n324 = ~pi4  & ~n323;
  assign n325 = ~pi5  & ~n324;
  assign n326 = ~pi6  & ~n325;
  assign n327 = ~pi7  & ~n326;
  assign n328 = ~pi8  & ~n327;
  assign n329 = ~pi9  & ~n328;
  assign n330 = ~pi10  & ~n329;
  assign n331 = ~pi11  & ~n330;
  assign n332 = ~pi12  & ~n331;
  assign n333 = ~pi13  & ~n332;
  assign n334 = ~pi14  & ~n333;
  assign n335 = ~pi15  & ~n334;
  assign n336 = ~pi16  & ~n335;
  assign n337 = ~pi17  & ~n336;
  assign n338 = ~pi18  & ~n337;
  assign n339 = ~pi19  & ~n338;
  assign n340 = ~pi20  & ~n339;
  assign n341 = n319 & n340;
  assign n342 = n316 & ~n321;
  assign n343 = ~n320 & n342;
  assign po0  = n341 | ~n343;
  assign n345 = ~pi72  & ~pi73 ;
  assign n346 = ~pi84  & ~pi85 ;
  assign n347 = ~pi88  & ~pi89 ;
  assign n348 = ~pi92  & ~pi93 ;
  assign n349 = ~pi102  & ~pi103 ;
  assign n350 = ~pi114  & ~pi115 ;
  assign n351 = ~pi118  & ~pi119 ;
  assign n352 = ~pi116  & ~pi117 ;
  assign n353 = n351 & n352;
  assign n354 = ~pi112  & ~pi113 ;
  assign n355 = n350 & n354;
  assign n356 = n353 & n355;
  assign n357 = n149 & n356;
  assign n358 = ~pi110  & ~pi111 ;
  assign n359 = n357 & ~n358;
  assign n360 = ~pi106  & ~pi107 ;
  assign n361 = n137 & ~n146;
  assign n362 = ~n350 & n352;
  assign n363 = n351 & ~n362;
  assign n364 = n149 & ~n363;
  assign n365 = n138 & ~n361;
  assign n366 = ~n364 & n365;
  assign n367 = ~n359 & n360;
  assign n368 = n366 & n367;
  assign n369 = n349 & n368;
  assign n370 = ~pi98  & ~pi99 ;
  assign n371 = n369 & n370;
  assign n372 = ~pi94  & ~pi95 ;
  assign n373 = n371 & n372;
  assign n374 = ~n348 & n373;
  assign n375 = ~pi104  & ~pi105 ;
  assign n376 = n368 & ~n375;
  assign n377 = ~pi96  & ~pi97 ;
  assign n378 = n371 & ~n377;
  assign n379 = ~pi100  & ~pi101 ;
  assign n380 = n369 & ~n379;
  assign n381 = ~pi108  & ~pi109 ;
  assign n382 = n358 & ~n381;
  assign n383 = n357 & ~n382;
  assign n384 = n366 & ~n383;
  assign n385 = ~n376 & ~n384;
  assign n386 = ~n380 & n385;
  assign n387 = ~n378 & n386;
  assign n388 = n347 & ~n374;
  assign n389 = n387 & n388;
  assign n390 = n346 & n389;
  assign n391 = ~pi80  & ~pi81 ;
  assign n392 = n390 & n391;
  assign n393 = ~pi76  & ~pi77 ;
  assign n394 = n392 & n393;
  assign n395 = ~pi86  & ~pi87 ;
  assign n396 = n389 & ~n395;
  assign n397 = ~pi78  & ~pi79 ;
  assign n398 = n392 & ~n397;
  assign n399 = ~pi82  & ~pi83 ;
  assign n400 = n390 & ~n399;
  assign n401 = ~pi90  & ~pi91 ;
  assign n402 = n348 & ~n401;
  assign n403 = n373 & ~n402;
  assign n404 = n387 & ~n403;
  assign n405 = ~n396 & ~n404;
  assign n406 = ~n400 & n405;
  assign n407 = ~n398 & n406;
  assign n408 = ~n394 & n407;
  assign n409 = n345 & ~n408;
  assign n410 = ~pi66  & ~pi67 ;
  assign n411 = ~pi70  & ~pi71 ;
  assign n412 = ~pi68  & ~pi69 ;
  assign n413 = n411 & n412;
  assign n414 = ~pi64  & ~pi65 ;
  assign n415 = n410 & n414;
  assign n416 = n413 & n415;
  assign n417 = n409 & n416;
  assign n418 = ~pi60  & ~pi61 ;
  assign n419 = n417 & n418;
  assign n420 = ~pi58  & ~pi59 ;
  assign n421 = n419 & ~n420;
  assign n422 = ~pi74  & ~pi75 ;
  assign n423 = n394 & ~n422;
  assign n424 = ~pi62  & ~pi63 ;
  assign n425 = n417 & ~n424;
  assign n426 = ~n410 & n412;
  assign n427 = n411 & ~n426;
  assign n428 = n409 & ~n427;
  assign n429 = n407 & ~n423;
  assign n430 = ~n428 & n429;
  assign n431 = ~n425 & n430;
  assign n432 = ~pi56  & ~pi57 ;
  assign n433 = ~n419 & n431;
  assign n434 = n432 & ~n433;
  assign n435 = ~pi54  & ~pi55 ;
  assign n436 = n434 & ~n435;
  assign n437 = ~pi50  & ~pi51 ;
  assign n438 = ~pi46  & ~pi47 ;
  assign n439 = n437 & n438;
  assign n440 = ~pi44  & ~pi45 ;
  assign n441 = n439 & ~n440;
  assign n442 = ~pi52  & ~pi53 ;
  assign n443 = ~pi48  & ~pi49 ;
  assign n444 = n437 & ~n443;
  assign n445 = ~pi42  & ~pi43 ;
  assign n446 = ~pi40  & ~pi41 ;
  assign n447 = ~pi38  & ~pi39 ;
  assign n448 = ~pi36  & ~pi37 ;
  assign n449 = ~pi34  & ~pi35 ;
  assign n450 = ~pi32  & ~pi33 ;
  assign n451 = ~pi30  & ~pi31 ;
  assign n452 = n450 & ~n451;
  assign n453 = ~pi28  & ~pi29 ;
  assign n454 = ~pi24  & ~pi25 ;
  assign n455 = ~pi22  & ~pi23 ;
  assign n456 = ~pi20  & ~pi21 ;
  assign n457 = ~pi18  & ~pi19 ;
  assign n458 = ~pi16  & ~pi17 ;
  assign n459 = ~pi14  & ~pi15 ;
  assign n460 = ~pi12  & ~pi13 ;
  assign n461 = ~pi10  & ~pi11 ;
  assign n462 = ~pi8  & ~pi9 ;
  assign n463 = ~pi6  & ~pi7 ;
  assign n464 = ~pi4  & ~pi5 ;
  assign n465 = ~pi2  & ~pi3 ;
  assign n466 = n464 & ~n465;
  assign n467 = n463 & ~n466;
  assign n468 = n462 & ~n467;
  assign n469 = n461 & ~n468;
  assign n470 = n460 & ~n469;
  assign n471 = n459 & ~n470;
  assign n472 = n458 & ~n471;
  assign n473 = n457 & ~n472;
  assign n474 = n456 & ~n473;
  assign n475 = n455 & ~n474;
  assign n476 = n454 & ~n475;
  assign n477 = ~pi26  & ~pi27 ;
  assign n478 = ~n476 & n477;
  assign n479 = n450 & n453;
  assign n480 = ~n478 & n479;
  assign n481 = n449 & ~n452;
  assign n482 = ~n480 & n481;
  assign n483 = n448 & ~n482;
  assign n484 = n447 & ~n483;
  assign n485 = n446 & ~n484;
  assign n486 = n439 & n445;
  assign n487 = ~n485 & n486;
  assign n488 = n442 & ~n444;
  assign n489 = ~n441 & n488;
  assign n490 = ~n487 & n489;
  assign n491 = n434 & n490;
  assign n492 = ~n421 & n431;
  assign n493 = ~n436 & n492;
  assign po1  = n491 | ~n493;
  assign n495 = n358 & n381;
  assign n496 = n360 & n375;
  assign n497 = n349 & n379;
  assign n498 = n496 & ~n497;
  assign n499 = n348 & n372;
  assign n500 = n347 & n401;
  assign n501 = n346 & n395;
  assign n502 = n391 & n399;
  assign n503 = n393 & n397;
  assign n504 = n345 & n422;
  assign n505 = ~n413 & n504;
  assign n506 = n503 & ~n505;
  assign n507 = n502 & ~n506;
  assign n508 = n501 & ~n507;
  assign n509 = n500 & ~n508;
  assign n510 = n499 & ~n509;
  assign n511 = n495 & n496;
  assign n512 = n370 & n377;
  assign n513 = n497 & n512;
  assign n514 = n511 & n513;
  assign n515 = ~n510 & n514;
  assign n516 = n495 & ~n498;
  assign n517 = ~n515 & n516;
  assign n518 = n357 & ~n517;
  assign n519 = n438 & n440;
  assign n520 = n445 & n446;
  assign n521 = n447 & n448;
  assign n522 = n449 & n450;
  assign n523 = n451 & n453;
  assign n524 = n454 & n477;
  assign n525 = n455 & n456;
  assign n526 = n457 & n458;
  assign n527 = n459 & n460;
  assign n528 = n461 & n462;
  assign n529 = n463 & n464;
  assign n530 = n528 & ~n529;
  assign n531 = n527 & ~n530;
  assign n532 = n526 & ~n531;
  assign n533 = n525 & ~n532;
  assign n534 = n524 & ~n533;
  assign n535 = n523 & ~n534;
  assign n536 = n522 & ~n535;
  assign n537 = n521 & ~n536;
  assign n538 = n520 & ~n537;
  assign n539 = n519 & ~n538;
  assign n540 = n148 & ~n353;
  assign n541 = n139 & ~n540;
  assign n542 = n357 & n514;
  assign n543 = n503 & n504;
  assign n544 = n416 & n543;
  assign n545 = n501 & n502;
  assign n546 = n499 & n500;
  assign n547 = n545 & n546;
  assign n548 = n544 & n547;
  assign po6  = ~n542 | ~n548;
  assign n550 = n418 & n424;
  assign n551 = n435 & n442;
  assign n552 = n420 & n432;
  assign n553 = ~n551 & n552;
  assign n554 = n550 & ~n553;
  assign n555 = ~po6  & ~n554;
  assign n556 = n541 & ~n555;
  assign n557 = n539 & ~n556;
  assign n558 = n437 & n443;
  assign n559 = n556 & ~n558;
  assign n560 = n550 & ~n552;
  assign n561 = ~po6  & ~n560;
  assign n562 = n541 & n558;
  assign n563 = ~n561 & n562;
  assign n564 = ~n559 & ~n563;
  assign n565 = ~n539 & n564;
  assign n566 = ~n518 & ~n557;
  assign po2  = n565 | ~n566;
  assign n568 = n356 & ~n511;
  assign n569 = n149 & ~n568;
  assign n570 = ~n542 & n569;
  assign n571 = n550 & n552;
  assign n572 = n551 & n558;
  assign n573 = n519 & n520;
  assign n574 = n521 & n522;
  assign n575 = n523 & n524;
  assign n576 = n525 & n526;
  assign n577 = n527 & n528;
  assign n578 = n576 & ~n577;
  assign n579 = n575 & ~n578;
  assign n580 = n574 & ~n579;
  assign n581 = n573 & ~n580;
  assign n582 = n572 & ~n581;
  assign n583 = n571 & ~n582;
  assign n584 = n416 & ~n583;
  assign n585 = n543 & ~n584;
  assign n586 = n545 & ~n585;
  assign n587 = n542 & n546;
  assign n588 = ~n586 & n587;
  assign po3  = ~n570 & ~n588;
  assign n590 = n571 & n572;
  assign n591 = n575 & n576;
  assign n592 = n573 & n574;
  assign n593 = ~n591 & n592;
  assign n594 = n590 & ~n593;
  assign n595 = n544 & ~n594;
  assign n596 = n547 & ~n595;
  assign n597 = n514 & ~n596;
  assign po4  = ~n357 | n597;
  assign n599 = n590 & n592;
  assign n600 = n548 & ~n599;
  assign po5  = ~n542 | n600;
  assign n602 = ~pi0  & ~pi1 ;
  assign n603 = n465 & n602;
  assign n604 = n529 & n603;
  assign n605 = n577 & n604;
  assign n606 = n591 & n605;
  assign n607 = n599 & n606;
  assign po7 = po6  | ~n607;
endmodule
