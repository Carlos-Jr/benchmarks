module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 ,
    pi5 , pi6 , pi7 , pi8 , pi9 ,
    pi10 , pi11 , pi12 , pi13 , pi14 ,
    pi15 , pi16 , pi17 , pi18 , pi19 ,
    pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 ,
    pi30 , pi31 , pi32 , pi33 , pi34 ,
    pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 ,
    pi45 , pi46 , pi47 , pi48 , pi49 ,
    pi50 , pi51 , pi52 , pi53 , pi54 ,
    pi55 , pi56 , pi57 , pi58 , pi59 ,
    po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 ,
    po14 , po15 , po16 , po17 ,
    po18 , po19 , po20 , po21 ,
    po22 , po23 , po24 , po25 ,
    po26 , po27 , po28 , po29   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 ,
    pi5 , pi6 , pi7 , pi8 , pi9 ,
    pi10 , pi11 , pi12 , pi13 , pi14 ,
    pi15 , pi16 , pi17 , pi18 , pi19 ,
    pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 ,
    pi30 , pi31 , pi32 , pi33 , pi34 ,
    pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 ,
    pi45 , pi46 , pi47 , pi48 , pi49 ,
    pi50 , pi51 , pi52 , pi53 , pi54 ,
    pi55 , pi56 , pi57 , pi58 , pi59 ;
  output po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 ,
    po14 , po15 , po16 , po17 ,
    po18 , po19 , po20 , po21 ,
    po22 , po23 , po24 , po25 ,
    po26 , po27 , po28 , po29 ;
  wire n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105,
    n106, n107, n108, n109, n110, n111, n112,
    n113, n114, n115, n116, n117, n118, n119,
    n120, n121, n122, n123, n124, n125, n126,
    n127, n128, n129, n130, n131, n132, n133,
    n134, n135, n136, n137, n138, n139, n140,
    n141, n142, n143, n144, n145, n146, n147,
    n148, n149, n150, n151, n152, n153, n154,
    n155, n156, n157, n158, n159, n160, n161,
    n162, n163, n164, n165, n166, n167, n168,
    n169, n170, n171, n172, n173, n175, n176,
    n177, n178, n179, n180, n181, n182, n183,
    n184, n185, n186, n187, n188, n189, n190,
    n191, n192, n193, n194, n195, n196, n197,
    n198, n199, n200, n201, n202, n203, n204,
    n205, n206, n207, n208, n209, n210, n211,
    n212, n213, n214, n215, n216, n217, n218,
    n219, n220, n221, n222, n223, n224, n225,
    n226, n227, n228, n229, n230, n231, n232,
    n233, n234, n235, n236, n237, n238, n239,
    n240, n241, n242, n243, n244, n245, n246,
    n247, n248, n249, n250, n251, n252, n253,
    n254, n255, n256, n257, n258, n259, n260,
    n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n271, n272, n273;
  assign n92 = pi28  & pi29 ;
  assign n93 = pi24  & pi25 ;
  assign n94 = pi14  & pi15 ;
  assign n95 = ~pi9  & ~pi10 ;
  assign n96 = pi11  & ~n95;
  assign n97 = ~pi12  & ~pi13 ;
  assign n98 = ~n96 & n97;
  assign n99 = n94 & ~n98;
  assign n100 = ~pi16  & ~n99;
  assign n101 = pi17  & ~n100;
  assign n102 = ~pi18  & ~n101;
  assign n103 = pi19  & ~n102;
  assign n104 = pi20  & n103;
  assign n105 = ~pi21  & ~pi22 ;
  assign n106 = ~n104 & n105;
  assign n107 = pi23  & ~n106;
  assign n108 = n93 & n107;
  assign n109 = ~pi26  & ~n108;
  assign n110 = pi27  & n92;
  assign n111 = ~n109 & n110;
  assign n112 = pi18  & n101;
  assign n113 = ~n102 & ~n112;
  assign n114 = ~pi22  & pi23 ;
  assign n115 = ~pi19  & n102;
  assign n116 = ~pi17  & n100;
  assign n117 = pi16  & ~n99;
  assign n118 = ~pi16  & n99;
  assign n119 = ~n117 & ~n118;
  assign n120 = pi14  & ~n98;
  assign n121 = ~pi15  & ~n120;
  assign n122 = ~pi24  & ~n107;
  assign n123 = pi0  & pi1 ;
  assign n124 = pi2  & pi3 ;
  assign n125 = pi4  & pi5 ;
  assign n126 = pi6  & pi7 ;
  assign n127 = pi8  & pi11 ;
  assign n128 = pi14  & pi20 ;
  assign n129 = ~pi21  & pi25 ;
  assign n130 = ~pi26  & pi27 ;
  assign n131 = n129 & n130;
  assign n132 = n97 & n128;
  assign n133 = n126 & n127;
  assign n134 = n124 & n125;
  assign n135 = n92 & n123;
  assign n136 = n95 & n114;
  assign n137 = n135 & n136;
  assign n138 = n133 & n134;
  assign n139 = n131 & n132;
  assign n140 = n138 & n139;
  assign n141 = n137 & n140;
  assign n142 = ~n99 & n141;
  assign n143 = ~n121 & n142;
  assign n144 = ~n101 & ~n116;
  assign n145 = n119 & n144;
  assign n146 = n143 & n145;
  assign n147 = ~n103 & ~n113;
  assign n148 = ~n115 & n147;
  assign n149 = n146 & n148;
  assign n150 = ~n122 & n149;
  assign n151 = ~n111 & ~n150;
  assign n152 = ~pi1  & ~pi2 ;
  assign n153 = ~pi3  & ~pi4 ;
  assign n154 = ~pi5  & ~pi6 ;
  assign n155 = ~pi7  & ~pi8 ;
  assign n156 = ~pi10  & ~pi12 ;
  assign n157 = ~pi13  & pi17 ;
  assign n158 = ~pi18  & pi19 ;
  assign n159 = pi20  & ~pi21 ;
  assign n160 = ~pi26  & n159;
  assign n161 = n157 & n158;
  assign n162 = n155 & n156;
  assign n163 = n153 & n154;
  assign n164 = n93 & n152;
  assign n165 = n94 & n114;
  assign n166 = n164 & n165;
  assign n167 = n162 & n163;
  assign n168 = n160 & n161;
  assign n169 = n96 & n168;
  assign n170 = n166 & n167;
  assign n171 = n169 & n170;
  assign n172 = ~n119 & n171;
  assign n173 = n111 & ~n172;
  assign po0  = n151 | n173;
  assign n175 = ~pi39  & ~pi40 ;
  assign n176 = pi41  & ~n175;
  assign n177 = ~pi42  & ~n176;
  assign n178 = ~pi43  & n177;
  assign n179 = pi44  & ~n178;
  assign n180 = pi45  & n179;
  assign n181 = ~pi46  & ~n180;
  assign n182 = pi47  & ~n181;
  assign n183 = ~pi48  & ~n182;
  assign n184 = pi49  & ~n183;
  assign n185 = pi50  & n184;
  assign n186 = ~pi51  & ~n185;
  assign n187 = ~pi52  & n186;
  assign n188 = pi53  & ~n187;
  assign n189 = ~pi53  & n187;
  assign n190 = ~n188 & ~n189;
  assign n191 = pi46  & ~pi47 ;
  assign n192 = n179 & ~n191;
  assign n193 = ~pi46  & pi47 ;
  assign n194 = ~n179 & ~n193;
  assign n195 = pi48  & n182;
  assign n196 = ~pi49  & ~n195;
  assign n197 = pi30  & pi31 ;
  assign n198 = pi32  & pi33 ;
  assign n199 = pi34  & pi35 ;
  assign n200 = pi36  & pi37 ;
  assign n201 = pi38  & pi41 ;
  assign n202 = ~pi42  & ~pi43 ;
  assign n203 = pi44  & pi45 ;
  assign n204 = pi50  & ~pi51 ;
  assign n205 = ~pi52  & pi54 ;
  assign n206 = pi55  & ~pi56 ;
  assign n207 = pi57  & pi58 ;
  assign n208 = pi59  & n207;
  assign n209 = n205 & n206;
  assign n210 = n203 & n204;
  assign n211 = n201 & n202;
  assign n212 = n199 & n200;
  assign n213 = n197 & n198;
  assign n214 = n175 & n213;
  assign n215 = n211 & n212;
  assign n216 = n209 & n210;
  assign n217 = n208 & n216;
  assign n218 = n214 & n215;
  assign n219 = n217 & n218;
  assign n220 = ~n192 & n219;
  assign n221 = ~n194 & n220;
  assign n222 = ~n184 & n221;
  assign n223 = ~n196 & n222;
  assign n224 = n190 & n223;
  assign n225 = ~pi0  & n224;
  assign n226 = pi54  & n188;
  assign n227 = pi55  & n226;
  assign n228 = ~pi56  & ~n227;
  assign n229 = n208 & ~n228;
  assign n230 = ~n225 & ~n229;
  assign n231 = pi43  & ~n177;
  assign n232 = pi51  & n185;
  assign n233 = pi56  & n227;
  assign n234 = ~pi55  & ~n226;
  assign n235 = ~n227 & ~n234;
  assign n236 = ~pi54  & ~n188;
  assign n237 = ~n226 & ~n236;
  assign n238 = ~pi50  & ~n184;
  assign n239 = ~n185 & ~n238;
  assign n240 = ~pi31  & ~pi32 ;
  assign n241 = ~pi33  & ~pi34 ;
  assign n242 = ~pi35  & ~pi36 ;
  assign n243 = ~pi37  & ~pi38 ;
  assign n244 = pi39  & ~pi40 ;
  assign n245 = pi41  & ~pi42 ;
  assign n246 = pi49  & ~pi52 ;
  assign n247 = n245 & n246;
  assign n248 = n243 & n244;
  assign n249 = n241 & n242;
  assign n250 = n193 & n240;
  assign n251 = n249 & n250;
  assign n252 = n247 & n248;
  assign n253 = n251 & n252;
  assign n254 = ~n231 & n253;
  assign n255 = ~pi48  & n254;
  assign n256 = n180 & n255;
  assign n257 = ~n186 & n256;
  assign n258 = ~n232 & ~n239;
  assign n259 = n257 & n258;
  assign n260 = ~n190 & n259;
  assign n261 = ~n237 & n260;
  assign n262 = ~n228 & n261;
  assign n263 = ~n233 & ~n235;
  assign n264 = n262 & n263;
  assign n265 = ~pi0  & ~pi30 ;
  assign n266 = ~n224 & n265;
  assign n267 = n264 & n266;
  assign n268 = ~n151 & ~n230;
  assign n269 = ~n267 & n268;
  assign po1  = ~n173 & ~n269;
  assign n271 = pi0  & pi30 ;
  assign n272 = n264 & ~n271;
  assign n273 = ~po0  & n229;
  assign po2  = ~n272 & n273;
  assign po3  = 1'b0;
  assign po4  = 1'b0;
  assign po5  = 1'b0;
  assign po6  = 1'b0;
  assign po7  = 1'b0;
  assign po8  = 1'b0;
  assign po9  = 1'b0;
  assign po10  = 1'b0;
  assign po11  = 1'b0;
  assign po12  = 1'b0;
  assign po13  = 1'b0;
  assign po14  = 1'b0;
  assign po15  = 1'b0;
  assign po16  = 1'b0;
  assign po17  = 1'b0;
  assign po18  = 1'b0;
  assign po19  = 1'b0;
  assign po20  = 1'b0;
  assign po21  = 1'b0;
  assign po22  = 1'b0;
  assign po23  = 1'b0;
  assign po24  = 1'b0;
  assign po25  = 1'b0;
  assign po26  = 1'b0;
  assign po27  = 1'b0;
  assign po28  = 1'b0;
  assign po29  = 1'b0;
endmodule
