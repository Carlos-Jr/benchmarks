module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 ,
    po0 , po1 , po2 , po3 , po4 , po5 , po6   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 ;
  wire n19, n20, n21, n22, n23, n24, n25,
    n26, n27, n28, n29, n30, n31, n32, n33,
    n34, n35, n36, n37, n38, n39, n40, n41,
    n42, n43, n44, n45, n46, n47, n48, n49,
    n50, n51, n52, n53, n54, n55, n56, n57,
    n58, n59, n60, n61, n62, n63, n64, n65,
    n66, n67, n68, n69, n70, n71, n72, n73,
    n74, n75, n76, n77, n78, n79, n80, n81,
    n82, n83, n84, n85, n86, n87, n88, n89,
    n90, n91, n92, n93, n94, n95, n96, n97,
    n98, n99, n100, n101, n102, n103, n104,
    n105, n106, n107, n108, n109, n110, n111,
    n112, n113, n114, n115, n116, n117, n118,
    n119, n120, n121, n122, n123, n124, n125,
    n126, n127, n128, n129, n130, n131, n132,
    n133, n134, n135, n136, n137, n138, n139,
    n140, n141, n142, n143, n144, n145, n146,
    n147, n148, n149, n150, n151, n152, n153,
    n154, n155, n156, n157, n158, n159, n160,
    n161, n162, n163, n164, n165, n166, n167,
    n168, n169, n170, n171, n172, n173, n174,
    n175, n176, n177, n178, n179, n180, n181,
    n182, n183, n184, n185, n186, n187, n188,
    n189, n190, n191, n192, n193, n194, n195,
    n196, n197, n198, n199, n200, n201, n202,
    n203, n204, n205, n206, n207, n208, n209,
    n210, n211, n213, n214, n215, n216, n217,
    n218, n219, n220, n221, n222, n223, n224,
    n225, n226, n227, n228, n229, n230, n231,
    n232, n233, n234, n235, n236, n237, n238,
    n239, n240, n241, n242, n243, n244, n245,
    n246, n247, n248, n249, n250, n251, n252,
    n253, n254, n255, n256, n257, n258, n259,
    n260, n261, n262, n263, n264, n265, n266,
    n267, n268, n269, n270, n271, n272, n273,
    n274, n275, n276, n277, n278, n279, n280,
    n281, n282, n283, n284, n285, n286, n287,
    n288, n289, n290, n291, n292, n293, n294,
    n295, n296, n297, n298, n299, n300, n301,
    n302, n303, n304, n305, n306, n307, n308,
    n309, n310, n311, n312, n313, n314, n315,
    n316, n317, n318, n319, n320, n321, n322,
    n323, n324, n325, n326, n327, n328, n329,
    n330, n331, n332, n333, n334, n335, n336,
    n337, n338, n339, n340, n341, n342, n343,
    n344, n345, n346, n347, n348, n349, n350,
    n351, n352, n353, n354, n355, n356, n357,
    n358, n359, n360, n361, n362, n363, n364,
    n365, n366, n367, n368, n369, n370, n371,
    n372, n373, n374, n375, n376, n377, n378,
    n379, n380, n381, n382, n383, n384, n385,
    n386, n387, n388, n389, n390, n391, n392,
    n393, n394, n395, n396, n397, n398, n399,
    n400, n401, n402, n403, n404, n405, n406,
    n407, n408, n409, n410, n411, n412, n413,
    n414, n415, n416, n417, n418, n419, n420,
    n421, n422, n423, n424, n425, n426, n427,
    n428, n429, n430, n431;
  assign n19 = pi4  & pi8 ;
  assign n20 = pi1  & pi4 ;
  assign n21 = ~pi4  & pi8 ;
  assign n22 = ~pi1  & pi4 ;
  assign n23 = ~pi4  & ~pi8 ;
  assign n24 = ~n22 & ~n23;
  assign n25 = ~n20 & ~n21;
  assign n26 = pi0  & n383;
  assign n27 = ~pi6  & ~pi7 ;
  assign n28 = ~pi0  & ~n20;
  assign n29 = n27 & ~n28;
  assign n30 = pi0  & ~n383;
  assign n31 = ~pi0  & pi1 ;
  assign n32 = ~pi0  & n20;
  assign n33 = pi4  & n31;
  assign n34 = ~n30 & ~n384;
  assign n35 = ~pi6  & ~n34;
  assign n36 = ~pi7  & n35;
  assign n37 = n27 & ~n34;
  assign n38 = ~n26 & n29;
  assign n39 = ~n19 & ~n385;
  assign n40 = ~pi5  & ~n39;
  assign n41 = ~pi4  & pi7 ;
  assign n42 = ~pi2  & ~pi7 ;
  assign n43 = pi1  & pi5 ;
  assign n44 = pi1  & ~pi2 ;
  assign n45 = pi5  & ~pi7 ;
  assign n46 = n44 & n45;
  assign n47 = n42 & n43;
  assign n48 = ~n41 & ~n386;
  assign n49 = pi3  & ~n48;
  assign n50 = ~pi3  & pi4 ;
  assign n51 = pi4  & pi7 ;
  assign n52 = ~pi3  & n51;
  assign n53 = pi7  & n50;
  assign n54 = ~n49 & ~n387;
  assign n55 = ~pi8  & ~n54;
  assign n56 = ~pi4  & pi5 ;
  assign n57 = pi5  & pi8 ;
  assign n58 = ~pi4  & n57;
  assign n59 = pi8  & n56;
  assign n60 = ~n55 & ~n388;
  assign n61 = ~n40 & n60;
  assign n62 = ~pi9  & ~n61;
  assign n63 = ~pi5  & pi6 ;
  assign n64 = pi6  & pi9 ;
  assign n65 = ~pi5  & n64;
  assign n66 = pi9  & n63;
  assign n67 = pi5  & ~pi6 ;
  assign n68 = ~n41 & n44;
  assign n69 = pi3  & pi4 ;
  assign n70 = ~n19 & ~n69;
  assign n71 = pi4  & ~pi8 ;
  assign n72 = ~pi3  & n71;
  assign n73 = ~pi4  & ~pi7 ;
  assign n74 = ~n72 & ~n73;
  assign n75 = ~pi2  & ~n74;
  assign n76 = pi1  & n75;
  assign n77 = ~n19 & ~n41;
  assign n78 = n44 & ~n69;
  assign n79 = n77 & n78;
  assign n80 = n68 & n70;
  assign n81 = ~pi7  & ~pi8 ;
  assign n82 = ~pi1  & pi2 ;
  assign n83 = n81 & n82;
  assign n84 = ~pi9  & ~n83;
  assign n85 = ~n390 & n84;
  assign n86 = ~pi6  & ~n85;
  assign n87 = pi5  & n86;
  assign n88 = n67 & ~n85;
  assign n89 = ~n389 & ~n391;
  assign n90 = ~n62 & n89;
  assign n91 = ~pi10  & ~n90;
  assign n92 = ~pi6  & pi7 ;
  assign n93 = ~pi6  & pi10 ;
  assign n94 = pi7  & n93;
  assign n95 = pi10  & n92;
  assign n96 = ~pi2  & pi3 ;
  assign n97 = pi2  & ~pi3 ;
  assign n98 = ~n96 & ~n97;
  assign n99 = ~pi8  & ~pi9 ;
  assign n100 = ~pi9  & ~n98;
  assign n101 = ~pi8  & n100;
  assign n102 = ~n98 & n99;
  assign n103 = ~pi10  & ~n393;
  assign n104 = ~pi7  & ~n103;
  assign n105 = pi8  & pi10 ;
  assign n106 = pi9  & pi10 ;
  assign n107 = pi8  & n106;
  assign n108 = pi9  & n105;
  assign n109 = ~n104 & ~n394;
  assign n110 = pi6  & ~n109;
  assign n111 = ~n392 & ~n110;
  assign n112 = ~n91 & n111;
  assign n113 = pi1  & pi2 ;
  assign n114 = pi0  & ~n113;
  assign n115 = ~pi0  & pi2 ;
  assign n116 = pi4  & ~pi7 ;
  assign n117 = ~n115 & n116;
  assign n118 = pi0  & n113;
  assign n119 = ~pi0  & ~pi2 ;
  assign n120 = ~n118 & ~n119;
  assign n121 = ~pi7  & ~n120;
  assign n122 = pi4  & n121;
  assign n123 = ~n114 & n117;
  assign n124 = pi8  & ~pi9 ;
  assign n125 = ~pi4  & ~pi9 ;
  assign n126 = ~n42 & ~n125;
  assign n127 = ~pi1  & ~n126;
  assign n128 = ~n124 & ~n127;
  assign n129 = ~n395 & ~n124;
  assign n130 = ~n127 & n129;
  assign n131 = ~n395 & n128;
  assign n132 = ~pi6  & ~n396;
  assign n133 = ~pi7  & pi9 ;
  assign n134 = pi7  & ~n69;
  assign n135 = ~pi9  & n134;
  assign n136 = ~pi8  & n135;
  assign n137 = n99 & n134;
  assign n138 = ~n133 & ~n397;
  assign n139 = ~n132 & n138;
  assign n140 = ~pi5  & ~n139;
  assign n141 = ~pi4  & ~n27;
  assign n142 = pi3  & ~n141;
  assign n143 = ~pi7  & ~n113;
  assign n144 = pi4  & ~n99;
  assign n145 = ~n143 & ~n144;
  assign n146 = ~pi4  & ~pi6 ;
  assign n147 = ~pi4  & n27;
  assign n148 = ~pi7  & n146;
  assign n149 = pi4  & n99;
  assign n150 = ~n398 & ~n149;
  assign n151 = pi2  & ~n150;
  assign n152 = pi1  & n151;
  assign n153 = pi7  & ~pi9 ;
  assign n154 = n71 & n153;
  assign n155 = ~n152 & ~n154;
  assign n156 = pi3  & ~n155;
  assign n157 = pi3  & ~n143;
  assign n158 = ~n150 & n157;
  assign n159 = n142 & n145;
  assign n160 = pi6  & ~n99;
  assign n161 = ~n125 & ~n133;
  assign n162 = pi4  & n124;
  assign n163 = pi7  & pi9 ;
  assign n164 = ~n162 & ~n163;
  assign n165 = pi6  & ~n164;
  assign n166 = n160 & n161;
  assign n167 = ~n399 & ~n400;
  assign n168 = pi5  & ~n167;
  assign n169 = ~pi4  & n124;
  assign n170 = ~pi9  & n21;
  assign n171 = ~n133 & ~n401;
  assign n172 = ~pi6  & ~n171;
  assign n173 = ~n168 & ~n172;
  assign n174 = ~n140 & n173;
  assign n175 = ~pi10  & ~n174;
  assign n176 = pi6  & pi7 ;
  assign n177 = ~pi9  & n176;
  assign n178 = pi6  & pi10 ;
  assign n179 = pi7  & n178;
  assign n180 = n124 & n179;
  assign n181 = n105 & n177;
  assign n182 = pi6  & ~pi9 ;
  assign n183 = ~pi4  & n182;
  assign n184 = ~pi1  & n67;
  assign n185 = ~n183 & ~n184;
  assign n186 = ~pi3  & ~n185;
  assign n187 = ~pi3  & pi5 ;
  assign n188 = ~pi3  & n67;
  assign n189 = ~pi6  & n187;
  assign n190 = ~n183 & ~n403;
  assign n191 = ~pi2  & ~n190;
  assign n192 = pi2  & n69;
  assign n193 = pi2  & pi3 ;
  assign n194 = pi4  & n182;
  assign n195 = n193 & n194;
  assign n196 = n182 & n192;
  assign n197 = ~n191 & ~n404;
  assign n198 = ~n186 & n197;
  assign n199 = ~pi7  & ~n198;
  assign n200 = ~pi10  & ~n199;
  assign n201 = ~pi8  & ~n176;
  assign n202 = ~pi10  & ~n404;
  assign n203 = ~n191 & n202;
  assign n204 = ~n186 & n202;
  assign n205 = ~n191 & n204;
  assign n206 = ~n186 & n203;
  assign n207 = ~pi7  & ~n405;
  assign n208 = ~n93 & ~n207;
  assign n209 = ~pi8  & ~n208;
  assign n210 = ~n200 & n201;
  assign n211 = ~n402 & ~n406;
  assign po1  = ~n175 & n211;
  assign n213 = pi0  & ~pi6 ;
  assign n214 = pi4  & ~pi6 ;
  assign n215 = pi0  & ~pi3 ;
  assign n216 = n214 & n215;
  assign n217 = n50 & n213;
  assign n218 = pi3  & n56;
  assign n219 = ~n407 & ~n218;
  assign n220 = pi1  & ~n219;
  assign n221 = pi0  & pi1 ;
  assign n222 = pi4  & ~n221;
  assign n223 = pi3  & n222;
  assign n224 = n69 & ~n221;
  assign n225 = ~n146 & ~n408;
  assign n226 = ~pi5  & ~n225;
  assign n227 = ~n220 & ~n226;
  assign n228 = pi2  & ~n227;
  assign n229 = pi3  & ~pi6 ;
  assign n230 = ~pi2  & n229;
  assign n231 = ~pi6  & n96;
  assign n232 = ~n187 & ~n409;
  assign n233 = pi4  & ~n232;
  assign n234 = ~n228 & ~n233;
  assign n235 = ~pi7  & ~n234;
  assign n236 = pi5  & pi6 ;
  assign n237 = pi5  & ~n69;
  assign n238 = pi6  & n237;
  assign n239 = ~n69 & n236;
  assign n240 = pi2  & n63;
  assign n241 = ~n184 & ~n240;
  assign n242 = pi4  & ~n241;
  assign n243 = pi3  & n242;
  assign n244 = n69 & ~n241;
  assign n245 = ~n410 & ~n411;
  assign n246 = ~n235 & n245;
  assign n247 = ~pi8  & ~n246;
  assign n248 = pi4  & pi5 ;
  assign n249 = pi7  & ~n248;
  assign n250 = pi6  & n249;
  assign n251 = n176 & ~n248;
  assign n252 = pi3  & n92;
  assign n253 = pi6  & ~pi7 ;
  assign n254 = ~pi2  & n253;
  assign n255 = ~n252 & ~n254;
  assign n256 = pi5  & ~n255;
  assign n257 = pi4  & n256;
  assign n258 = n248 & ~n255;
  assign n259 = ~n412 & ~n413;
  assign n260 = ~n247 & n259;
  assign n261 = ~pi9  & ~n260;
  assign n262 = n116 & n236;
  assign n263 = pi4  & pi6 ;
  assign n264 = n45 & n263;
  assign n265 = n248 & n253;
  assign n266 = ~n92 & ~n414;
  assign n267 = pi8  & ~n266;
  assign n268 = ~n261 & ~n267;
  assign n269 = ~pi10  & ~n268;
  assign n270 = pi5  & ~pi8 ;
  assign n271 = ~pi8  & pi9 ;
  assign n272 = pi5  & n271;
  assign n273 = pi9  & n270;
  assign n274 = ~n105 & ~n415;
  assign n275 = pi7  & ~n274;
  assign n276 = pi6  & n275;
  assign n277 = n176 & ~n274;
  assign n278 = pi5  & pi7 ;
  assign n279 = pi8  & ~n278;
  assign n280 = ~pi10  & ~n279;
  assign n281 = pi9  & ~n280;
  assign n282 = ~n416 & ~n281;
  assign n283 = ~n269 & n282;
  assign n284 = pi7  & n236;
  assign n285 = pi9  & ~n284;
  assign n286 = pi8  & ~n285;
  assign n287 = pi5  & ~n113;
  assign n288 = ~pi7  & ~n287;
  assign n289 = ~n236 & ~n288;
  assign n290 = ~pi5  & ~pi6 ;
  assign n291 = n221 & n290;
  assign n292 = ~n414 & ~n291;
  assign n293 = pi3  & ~n292;
  assign n294 = pi2  & n293;
  assign n295 = n193 & ~n292;
  assign n296 = pi4  & ~pi5 ;
  assign n297 = ~pi6  & ~n69;
  assign n298 = ~n296 & n297;
  assign n299 = ~pi9  & ~n134;
  assign n300 = ~pi7  & ~n67;
  assign n301 = ~pi3  & ~n300;
  assign n302 = ~pi4  & ~n253;
  assign n303 = ~pi9  & ~n302;
  assign n304 = ~n301 & n303;
  assign n305 = ~n298 & n299;
  assign n306 = ~n417 & n418;
  assign n307 = pi7  & ~n236;
  assign n308 = ~pi6  & ~n113;
  assign n309 = pi5  & n308;
  assign n310 = ~pi9  & ~n309;
  assign n311 = ~n307 & n310;
  assign n312 = ~n301 & n311;
  assign n313 = ~n302 & n312;
  assign n314 = ~n289 & n418;
  assign n315 = ~n417 & n419;
  assign n316 = ~n289 & n306;
  assign n317 = ~n286 & ~n420;
  assign n318 = pi3  & pi8 ;
  assign n319 = ~n97 & ~n318;
  assign n320 = n177 & n248;
  assign n321 = pi6  & ~n319;
  assign n322 = pi5  & n321;
  assign n323 = pi7  & n322;
  assign n324 = ~pi9  & n323;
  assign n325 = pi4  & n324;
  assign n326 = ~n319 & n320;
  assign n327 = ~pi8  & ~n420;
  assign n328 = ~n285 & ~n421;
  assign n329 = ~n327 & n328;
  assign n330 = ~n317 & ~n421;
  assign n331 = ~pi10  & ~n422;
  assign n332 = pi6  & pi8 ;
  assign n333 = pi8  & n284;
  assign n334 = n278 & n332;
  assign n335 = pi3  & ~pi5 ;
  assign n336 = n81 & n335;
  assign n337 = pi1  & pi3 ;
  assign n338 = pi0  & n337;
  assign n339 = ~pi5  & ~pi7 ;
  assign n340 = ~pi8  & n339;
  assign n341 = n338 & n340;
  assign n342 = n221 & n336;
  assign n343 = ~n423 & ~n424;
  assign n344 = pi2  & ~n343;
  assign n345 = pi8  & n278;
  assign n346 = pi3  & pi6 ;
  assign n347 = n345 & n346;
  assign n348 = n284 & n318;
  assign n349 = ~n344 & ~n425;
  assign n350 = pi4  & ~n349;
  assign n351 = ~pi9  & ~pi10 ;
  assign n352 = n192 & n236;
  assign n353 = n81 & ~n290;
  assign n354 = n193 & n263;
  assign n355 = pi5  & ~n354;
  assign n356 = ~n63 & ~n355;
  assign n357 = ~pi7  & ~n356;
  assign n358 = ~pi8  & n357;
  assign n359 = ~n352 & n353;
  assign n360 = n351 & ~n426;
  assign n361 = ~n350 & n360;
  assign n362 = ~pi2  & n19;
  assign n363 = ~pi2  & n176;
  assign n364 = pi5  & n19;
  assign n365 = n363 & n364;
  assign n366 = n284 & n362;
  assign n367 = ~pi7  & n23;
  assign n368 = ~pi4  & n81;
  assign n369 = ~pi5  & n23;
  assign n370 = n27 & n369;
  assign n371 = n290 & n428;
  assign n372 = ~n427 & ~n429;
  assign n373 = ~pi3  & n351;
  assign n374 = ~pi9  & ~n372;
  assign n375 = ~pi10  & n374;
  assign n376 = ~pi3  & n375;
  assign n377 = ~n372 & n373;
  assign n378 = n81 & n351;
  assign n379 = ~pi9  & ~n352;
  assign n380 = ~pi10  & n379;
  assign n381 = n81 & n380;
  assign n382 = ~n352 & n378;
  assign n383 = n24 | ~n25;
  assign n384 = n32 | n33;
  assign n385 = n38 | n36 | n37;
  assign n386 = n46 | n47;
  assign n387 = n52 | n53;
  assign n388 = n58 | n59;
  assign n389 = n65 | n66;
  assign n390 = n80 | n76 | n79;
  assign n391 = n87 | n88;
  assign n392 = n94 | n95;
  assign n393 = n101 | n102;
  assign n394 = n107 | n108;
  assign n395 = n122 | n123;
  assign n396 = n130 | n131;
  assign n397 = n136 | n137;
  assign n398 = n147 | n148;
  assign n399 = n159 | n156 | n158;
  assign n400 = n165 | n166;
  assign n401 = n169 | n170;
  assign n402 = n180 | n181;
  assign n403 = n188 | n189;
  assign n404 = n195 | n196;
  assign n405 = n205 | n206;
  assign n406 = n209 | n210;
  assign n407 = n216 | n217;
  assign n408 = n223 | n224;
  assign n409 = n230 | n231;
  assign n410 = n238 | n239;
  assign n411 = n243 | n244;
  assign n412 = n250 | n251;
  assign n413 = n257 | n258;
  assign n414 = n265 | n262 | n264;
  assign n415 = n272 | n273;
  assign n416 = n276 | n277;
  assign n417 = n294 | n295;
  assign n418 = n304 | n305;
  assign n419 = n313 | n314;
  assign n420 = n315 | n316;
  assign n421 = n325 | n326;
  assign n422 = n329 | n330;
  assign n423 = n333 | n334;
  assign n424 = n341 | n342;
  assign n425 = n347 | n348;
  assign n426 = n358 | n359;
  assign n427 = n365 | n366;
  assign n428 = n367 | n368;
  assign n429 = n370 | n371;
  assign n430 = n376 | n377;
  assign n431 = n381 | n382;
  assign po0  = ~n112;
  assign po2  = ~n283;
  assign po3  = ~n430;
  assign po4  = ~n331;
  assign po5  = ~n361;
  assign po6  = ~n431;
endmodule
