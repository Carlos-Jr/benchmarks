module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 , pi32 ,
    pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 , pi40 ,
    pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 , pi56 ,
    pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 , pi64 ,
    pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 ,
    pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 ,
    pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 ,
    pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 ,
    pi97 , pi98 , pi99 , pi100 , pi101 , pi102 , pi103 ,
    pi104 , pi105 , pi106 , pi107 , pi108 , pi109 , pi110 ,
    pi111 , pi112 , pi113 , pi114 , pi115 , pi116 , pi117 ,
    pi118 , pi119 , pi120 , pi121 , pi122 , pi123 , pi124 ,
    pi125 , pi126 , pi127 ,
    po0 , po1 , po2 , po3 , po4 , po5 ,
    po6 , po7 , po8 , po9 , po10 ,
    po11 , po12 , po13 , po14 , po15 ,
    po16 , po17 , po18 , po19 , po20 ,
    po21 , po22 , po23 , po24 , po25 ,
    po26 , po27 , po28 , po29 , po30 ,
    po31 , po32 , po33 , po34 , po35 ,
    po36 , po37 , po38 , po39 , po40 ,
    po41 , po42 , po43 , po44 , po45 ,
    po46 , po47 , po48 , po49 , po50 ,
    po51 , po52 , po53 , po54 , po55 ,
    po56 , po57 , po58 , po59 , po60 ,
    po61 , po62 , po63   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    pi32 , pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 ,
    pi56 , pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 ,
    pi64 , pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 ,
    pi72 , pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 ,
    pi80 , pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 ,
    pi88 , pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 ,
    pi96 , pi97 , pi98 , pi99 , pi100 , pi101 , pi102 ,
    pi103 , pi104 , pi105 , pi106 , pi107 , pi108 , pi109 ,
    pi110 , pi111 , pi112 , pi113 , pi114 , pi115 , pi116 ,
    pi117 , pi118 , pi119 , pi120 , pi121 , pi122 , pi123 ,
    pi124 , pi125 , pi126 , pi127 ;
  output po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 , po14 ,
    po15 , po16 , po17 , po18 , po19 ,
    po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 ,
    po30 , po31 , po32 , po33 , po34 ,
    po35 , po36 , po37 , po38 , po39 ,
    po40 , po41 , po42 , po43 , po44 ,
    po45 , po46 , po47 , po48 , po49 ,
    po50 , po51 , po52 , po53 , po54 ,
    po55 , po56 , po57 , po58 , po59 ,
    po60 , po61 , po62 , po63 ;
  wire n193, n194, n195, n197, n198, n199, n201,
    n202, n203, n204, n205, n206, n207, n208,
    n209, n210, n211, n212, n214, n215, n216,
    n217, n218, n219, n220, n221, n222, n223,
    n224, n225, n226, n227, n228, n229, n230,
    n231, n232, n233, n234, n235, n236, n237,
    n238, n239, n240, n241, n242, n243, n244,
    n245, n247, n248, n249, n250, n251, n252,
    n253, n254, n255, n256, n257, n258, n259,
    n260, n261, n262, n263, n264, n265, n266,
    n267, n268, n269, n270, n271, n272, n273,
    n274, n275, n276, n277, n278, n279, n280,
    n281, n282, n283, n285, n286, n287, n288,
    n289, n290, n291, n292, n293, n294, n295,
    n296, n297, n298, n299, n300, n301, n302,
    n303, n304, n305, n306, n307, n308, n309,
    n310, n311, n312, n313, n314, n315, n316,
    n317, n318, n319, n320, n321, n322, n323,
    n324, n325, n326, n327, n328, n329, n330,
    n332, n333, n334, n335, n336, n337, n338,
    n339, n340, n341, n342, n343, n344, n345,
    n346, n347, n348, n349, n350, n351, n352,
    n353, n354, n355, n356, n357, n358, n359,
    n360, n361, n362, n363, n364, n365, n366,
    n367, n368, n369, n370, n371, n372, n373,
    n374, n375, n376, n377, n378, n379, n380,
    n381, n382, n383, n384, n385, n386, n387,
    n388, n390, n391, n392, n393, n394, n395,
    n396, n397, n398, n399, n400, n401, n402,
    n403, n404, n405, n406, n407, n408, n409,
    n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423,
    n424, n425, n426, n427, n428, n429, n430,
    n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444,
    n445, n446, n447, n448, n449, n450, n451,
    n452, n453, n454, n455, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487,
    n488, n489, n490, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501,
    n502, n503, n504, n505, n506, n507, n508,
    n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n533, n534, n535, n536, n537,
    n538, n539, n540, n541, n542, n543, n544,
    n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n557, n558,
    n559, n560, n561, n562, n563, n564, n565,
    n566, n567, n568, n569, n570, n571, n572,
    n573, n574, n575, n576, n577, n578, n579,
    n580, n581, n582, n583, n584, n585, n586,
    n587, n588, n589, n590, n591, n592, n593,
    n594, n595, n596, n597, n598, n599, n600,
    n601, n602, n603, n604, n605, n606, n607,
    n608, n609, n610, n611, n612, n613, n614,
    n615, n616, n618, n619, n620, n621, n622,
    n623, n624, n625, n626, n627, n628, n629,
    n630, n631, n632, n633, n634, n635, n636,
    n637, n638, n639, n640, n641, n642, n643,
    n644, n645, n646, n647, n648, n649, n650,
    n651, n652, n653, n654, n655, n656, n657,
    n658, n659, n660, n661, n662, n663, n664,
    n665, n666, n667, n668, n669, n670, n671,
    n672, n673, n674, n675, n676, n677, n678,
    n679, n680, n681, n682, n683, n684, n685,
    n686, n687, n688, n689, n690, n691, n692,
    n693, n694, n695, n696, n697, n698, n699,
    n700, n701, n702, n703, n704, n705, n706,
    n707, n708, n709, n710, n712, n713, n714,
    n715, n716, n717, n718, n719, n720, n721,
    n722, n723, n724, n725, n726, n727, n728,
    n729, n730, n731, n732, n733, n734, n735,
    n736, n737, n738, n739, n740, n741, n742,
    n743, n744, n745, n746, n747, n748, n749,
    n750, n751, n752, n753, n754, n755, n756,
    n757, n758, n759, n760, n761, n762, n763,
    n764, n765, n766, n767, n768, n769, n770,
    n771, n772, n773, n774, n775, n776, n777,
    n778, n779, n780, n781, n782, n783, n784,
    n785, n786, n787, n788, n789, n790, n791,
    n792, n793, n794, n795, n796, n797, n798,
    n799, n800, n801, n802, n803, n804, n805,
    n806, n807, n808, n809, n810, n811, n812,
    n813, n815, n816, n817, n818, n819, n820,
    n821, n822, n823, n824, n825, n826, n827,
    n828, n829, n830, n831, n832, n833, n834,
    n835, n836, n837, n838, n839, n840, n841,
    n842, n843, n844, n845, n846, n847, n848,
    n849, n850, n851, n852, n853, n854, n855,
    n856, n857, n858, n859, n860, n861, n862,
    n863, n864, n865, n866, n867, n868, n869,
    n870, n871, n872, n873, n874, n875, n876,
    n877, n878, n879, n880, n881, n882, n883,
    n884, n885, n886, n887, n888, n889, n890,
    n891, n892, n893, n894, n895, n896, n897,
    n898, n899, n900, n901, n902, n903, n904,
    n905, n906, n907, n908, n909, n910, n911,
    n912, n913, n914, n915, n916, n917, n918,
    n919, n920, n921, n922, n923, n924, n925,
    n927, n928, n929, n930, n931, n932, n933,
    n934, n935, n936, n937, n938, n939, n940,
    n941, n942, n943, n944, n945, n946, n947,
    n948, n949, n950, n951, n952, n953, n954,
    n955, n956, n957, n958, n959, n960, n961,
    n962, n963, n964, n965, n966, n967, n968,
    n969, n970, n971, n972, n973, n974, n975,
    n976, n977, n978, n979, n980, n981, n982,
    n983, n984, n985, n986, n987, n988, n989,
    n990, n991, n992, n993, n994, n995, n996,
    n997, n998, n999, n1000, n1001, n1002,
    n1003, n1004, n1005, n1006, n1007, n1008,
    n1009, n1010, n1011, n1012, n1013, n1014,
    n1015, n1016, n1017, n1018, n1019, n1020,
    n1021, n1022, n1023, n1024, n1025, n1026,
    n1027, n1028, n1029, n1030, n1031, n1032,
    n1033, n1034, n1035, n1036, n1037, n1038,
    n1039, n1040, n1041, n1042, n1043, n1044,
    n1045, n1046, n1048, n1049, n1050, n1051,
    n1052, n1053, n1054, n1055, n1056, n1057,
    n1058, n1059, n1060, n1061, n1062, n1063,
    n1064, n1065, n1066, n1067, n1068, n1069,
    n1070, n1071, n1072, n1073, n1074, n1075,
    n1076, n1077, n1078, n1079, n1080, n1081,
    n1082, n1083, n1084, n1085, n1086, n1087,
    n1088, n1089, n1090, n1091, n1092, n1093,
    n1094, n1095, n1096, n1097, n1098, n1099,
    n1100, n1101, n1102, n1103, n1104, n1105,
    n1106, n1107, n1108, n1109, n1110, n1111,
    n1112, n1113, n1114, n1115, n1116, n1117,
    n1118, n1119, n1120, n1121, n1122, n1123,
    n1124, n1125, n1126, n1127, n1128, n1129,
    n1130, n1131, n1132, n1133, n1134, n1135,
    n1136, n1137, n1138, n1139, n1140, n1141,
    n1142, n1143, n1144, n1145, n1146, n1147,
    n1148, n1149, n1150, n1151, n1152, n1153,
    n1154, n1155, n1156, n1157, n1158, n1159,
    n1160, n1161, n1162, n1163, n1164, n1165,
    n1166, n1167, n1168, n1169, n1170, n1171,
    n1172, n1173, n1174, n1175, n1176, n1178,
    n1179, n1180, n1181, n1182, n1183, n1184,
    n1185, n1186, n1187, n1188, n1189, n1190,
    n1191, n1192, n1193, n1194, n1195, n1196,
    n1197, n1198, n1199, n1200, n1201, n1202,
    n1203, n1204, n1205, n1206, n1207, n1208,
    n1209, n1210, n1211, n1212, n1213, n1214,
    n1215, n1216, n1217, n1218, n1219, n1220,
    n1221, n1222, n1223, n1224, n1225, n1226,
    n1227, n1228, n1229, n1230, n1231, n1232,
    n1233, n1234, n1235, n1236, n1237, n1238,
    n1239, n1240, n1241, n1242, n1243, n1244,
    n1245, n1246, n1247, n1248, n1249, n1250,
    n1251, n1252, n1253, n1254, n1255, n1256,
    n1257, n1258, n1259, n1260, n1261, n1262,
    n1263, n1264, n1265, n1266, n1267, n1268,
    n1269, n1270, n1271, n1272, n1273, n1274,
    n1275, n1276, n1277, n1278, n1279, n1280,
    n1281, n1282, n1283, n1284, n1285, n1286,
    n1287, n1288, n1289, n1290, n1291, n1292,
    n1293, n1294, n1295, n1296, n1297, n1298,
    n1299, n1300, n1301, n1302, n1303, n1304,
    n1305, n1306, n1307, n1308, n1309, n1310,
    n1311, n1312, n1313, n1314, n1315, n1317,
    n1318, n1319, n1320, n1321, n1322, n1323,
    n1324, n1325, n1326, n1327, n1328, n1329,
    n1330, n1331, n1332, n1333, n1334, n1335,
    n1336, n1337, n1338, n1339, n1340, n1341,
    n1342, n1343, n1344, n1345, n1346, n1347,
    n1348, n1349, n1350, n1351, n1352, n1353,
    n1354, n1355, n1356, n1357, n1358, n1359,
    n1360, n1361, n1362, n1363, n1364, n1365,
    n1366, n1367, n1368, n1369, n1370, n1371,
    n1372, n1373, n1374, n1375, n1376, n1377,
    n1378, n1379, n1380, n1381, n1382, n1383,
    n1384, n1385, n1386, n1387, n1388, n1389,
    n1390, n1391, n1392, n1393, n1394, n1395,
    n1396, n1397, n1398, n1399, n1400, n1401,
    n1402, n1403, n1404, n1405, n1406, n1407,
    n1408, n1409, n1410, n1411, n1412, n1413,
    n1414, n1415, n1416, n1417, n1418, n1419,
    n1420, n1421, n1422, n1423, n1424, n1425,
    n1426, n1427, n1428, n1429, n1430, n1431,
    n1432, n1433, n1434, n1435, n1436, n1437,
    n1438, n1439, n1440, n1441, n1442, n1443,
    n1444, n1445, n1446, n1447, n1448, n1449,
    n1450, n1451, n1452, n1453, n1454, n1455,
    n1456, n1457, n1458, n1459, n1460, n1461,
    n1462, n1463, n1465, n1466, n1467, n1468,
    n1469, n1470, n1471, n1472, n1473, n1474,
    n1475, n1476, n1477, n1478, n1479, n1480,
    n1481, n1482, n1483, n1484, n1485, n1486,
    n1487, n1488, n1489, n1490, n1491, n1492,
    n1493, n1494, n1495, n1496, n1497, n1498,
    n1499, n1500, n1501, n1502, n1503, n1504,
    n1505, n1506, n1507, n1508, n1509, n1510,
    n1511, n1512, n1513, n1514, n1515, n1516,
    n1517, n1518, n1519, n1520, n1521, n1522,
    n1523, n1524, n1525, n1526, n1527, n1528,
    n1529, n1530, n1531, n1532, n1533, n1534,
    n1535, n1536, n1537, n1538, n1539, n1540,
    n1541, n1542, n1543, n1544, n1545, n1546,
    n1547, n1548, n1549, n1550, n1551, n1552,
    n1553, n1554, n1555, n1556, n1557, n1558,
    n1559, n1560, n1561, n1562, n1563, n1564,
    n1565, n1566, n1567, n1568, n1569, n1570,
    n1571, n1572, n1573, n1574, n1575, n1576,
    n1577, n1578, n1579, n1580, n1581, n1582,
    n1583, n1584, n1585, n1586, n1587, n1588,
    n1589, n1590, n1591, n1592, n1593, n1594,
    n1595, n1596, n1597, n1598, n1599, n1600,
    n1601, n1602, n1603, n1604, n1605, n1606,
    n1607, n1608, n1609, n1610, n1611, n1612,
    n1613, n1614, n1615, n1616, n1617, n1618,
    n1619, n1620, n1622, n1623, n1624, n1625,
    n1626, n1627, n1628, n1629, n1630, n1631,
    n1632, n1633, n1634, n1635, n1636, n1637,
    n1638, n1639, n1640, n1641, n1642, n1643,
    n1644, n1645, n1646, n1647, n1648, n1649,
    n1650, n1651, n1652, n1653, n1654, n1655,
    n1656, n1657, n1658, n1659, n1660, n1661,
    n1662, n1663, n1664, n1665, n1666, n1667,
    n1668, n1669, n1670, n1671, n1672, n1673,
    n1674, n1675, n1676, n1677, n1678, n1679,
    n1680, n1681, n1682, n1683, n1684, n1685,
    n1686, n1687, n1688, n1689, n1690, n1691,
    n1692, n1693, n1694, n1695, n1696, n1697,
    n1698, n1699, n1700, n1701, n1702, n1703,
    n1704, n1705, n1706, n1707, n1708, n1709,
    n1710, n1711, n1712, n1713, n1714, n1715,
    n1716, n1717, n1718, n1719, n1720, n1721,
    n1722, n1723, n1724, n1725, n1726, n1727,
    n1728, n1729, n1730, n1731, n1732, n1733,
    n1734, n1735, n1736, n1737, n1738, n1739,
    n1740, n1741, n1742, n1743, n1744, n1745,
    n1746, n1747, n1748, n1749, n1750, n1751,
    n1752, n1753, n1754, n1755, n1756, n1757,
    n1758, n1759, n1760, n1761, n1762, n1763,
    n1764, n1765, n1766, n1767, n1768, n1769,
    n1770, n1771, n1772, n1773, n1774, n1775,
    n1776, n1777, n1778, n1779, n1780, n1781,
    n1782, n1783, n1784, n1785, n1786, n1788,
    n1789, n1790, n1791, n1792, n1793, n1794,
    n1795, n1796, n1797, n1798, n1799, n1800,
    n1801, n1802, n1803, n1804, n1805, n1806,
    n1807, n1808, n1809, n1810, n1811, n1812,
    n1813, n1814, n1815, n1816, n1817, n1818,
    n1819, n1820, n1821, n1822, n1823, n1824,
    n1825, n1826, n1827, n1828, n1829, n1830,
    n1831, n1832, n1833, n1834, n1835, n1836,
    n1837, n1838, n1839, n1840, n1841, n1842,
    n1843, n1844, n1845, n1846, n1847, n1848,
    n1849, n1850, n1851, n1852, n1853, n1854,
    n1855, n1856, n1857, n1858, n1859, n1860,
    n1861, n1862, n1863, n1864, n1865, n1866,
    n1867, n1868, n1869, n1870, n1871, n1872,
    n1873, n1874, n1875, n1876, n1877, n1878,
    n1879, n1880, n1881, n1882, n1883, n1884,
    n1885, n1886, n1887, n1888, n1889, n1890,
    n1891, n1892, n1893, n1894, n1895, n1896,
    n1897, n1898, n1899, n1900, n1901, n1902,
    n1903, n1904, n1905, n1906, n1907, n1908,
    n1909, n1910, n1911, n1912, n1913, n1914,
    n1915, n1916, n1917, n1918, n1919, n1920,
    n1921, n1922, n1923, n1924, n1925, n1926,
    n1927, n1928, n1929, n1930, n1931, n1932,
    n1933, n1934, n1935, n1936, n1937, n1938,
    n1939, n1940, n1941, n1942, n1943, n1944,
    n1945, n1946, n1947, n1948, n1949, n1950,
    n1951, n1952, n1953, n1954, n1955, n1956,
    n1957, n1958, n1959, n1960, n1961, n1963,
    n1964, n1965, n1966, n1967, n1968, n1969,
    n1970, n1971, n1972, n1973, n1974, n1975,
    n1976, n1977, n1978, n1979, n1980, n1981,
    n1982, n1983, n1984, n1985, n1986, n1987,
    n1988, n1989, n1990, n1991, n1992, n1993,
    n1994, n1995, n1996, n1997, n1998, n1999,
    n2000, n2001, n2002, n2003, n2004, n2005,
    n2006, n2007, n2008, n2009, n2010, n2011,
    n2012, n2013, n2014, n2015, n2016, n2017,
    n2018, n2019, n2020, n2021, n2022, n2023,
    n2024, n2025, n2026, n2027, n2028, n2029,
    n2030, n2031, n2032, n2033, n2034, n2035,
    n2036, n2037, n2038, n2039, n2040, n2041,
    n2042, n2043, n2044, n2045, n2046, n2047,
    n2048, n2049, n2050, n2051, n2052, n2053,
    n2054, n2055, n2056, n2057, n2058, n2059,
    n2060, n2061, n2062, n2063, n2064, n2065,
    n2066, n2067, n2068, n2069, n2070, n2071,
    n2072, n2073, n2074, n2075, n2076, n2077,
    n2078, n2079, n2080, n2081, n2082, n2083,
    n2084, n2085, n2086, n2087, n2088, n2089,
    n2090, n2091, n2092, n2093, n2094, n2095,
    n2096, n2097, n2098, n2099, n2100, n2101,
    n2102, n2103, n2104, n2105, n2106, n2107,
    n2108, n2109, n2110, n2111, n2112, n2113,
    n2114, n2115, n2116, n2117, n2118, n2119,
    n2120, n2121, n2122, n2123, n2124, n2125,
    n2126, n2127, n2128, n2129, n2130, n2131,
    n2132, n2133, n2134, n2135, n2136, n2137,
    n2138, n2139, n2140, n2141, n2142, n2143,
    n2144, n2145, n2147, n2148, n2149, n2150,
    n2151, n2152, n2153, n2154, n2155, n2156,
    n2157, n2158, n2159, n2160, n2161, n2162,
    n2163, n2164, n2165, n2166, n2167, n2168,
    n2169, n2170, n2171, n2172, n2173, n2174,
    n2175, n2176, n2177, n2178, n2179, n2180,
    n2181, n2182, n2183, n2184, n2185, n2186,
    n2187, n2188, n2189, n2190, n2191, n2192,
    n2193, n2194, n2195, n2196, n2197, n2198,
    n2199, n2200, n2201, n2202, n2203, n2204,
    n2205, n2206, n2207, n2208, n2209, n2210,
    n2211, n2212, n2213, n2214, n2215, n2216,
    n2217, n2218, n2219, n2220, n2221, n2222,
    n2223, n2224, n2225, n2226, n2227, n2228,
    n2229, n2230, n2231, n2232, n2233, n2234,
    n2235, n2236, n2237, n2238, n2239, n2240,
    n2241, n2242, n2243, n2244, n2245, n2246,
    n2247, n2248, n2249, n2250, n2251, n2252,
    n2253, n2254, n2255, n2256, n2257, n2258,
    n2259, n2260, n2261, n2262, n2263, n2264,
    n2265, n2266, n2267, n2268, n2269, n2270,
    n2271, n2272, n2273, n2274, n2275, n2276,
    n2277, n2278, n2279, n2280, n2281, n2282,
    n2283, n2284, n2285, n2286, n2287, n2288,
    n2289, n2290, n2291, n2292, n2293, n2294,
    n2295, n2296, n2297, n2298, n2299, n2300,
    n2301, n2302, n2303, n2304, n2305, n2306,
    n2307, n2308, n2309, n2310, n2311, n2312,
    n2313, n2314, n2315, n2316, n2317, n2318,
    n2319, n2320, n2321, n2322, n2323, n2324,
    n2325, n2326, n2327, n2328, n2329, n2330,
    n2331, n2332, n2333, n2334, n2335, n2336,
    n2337, n2338, n2340, n2341, n2342, n2343,
    n2344, n2345, n2346, n2347, n2348, n2349,
    n2350, n2351, n2352, n2353, n2354, n2355,
    n2356, n2357, n2358, n2359, n2360, n2361,
    n2362, n2363, n2364, n2365, n2366, n2367,
    n2368, n2369, n2370, n2371, n2372, n2373,
    n2374, n2375, n2376, n2377, n2378, n2379,
    n2380, n2381, n2382, n2383, n2384, n2385,
    n2386, n2387, n2388, n2389, n2390, n2391,
    n2392, n2393, n2394, n2395, n2396, n2397,
    n2398, n2399, n2400, n2401, n2402, n2403,
    n2404, n2405, n2406, n2407, n2408, n2409,
    n2410, n2411, n2412, n2413, n2414, n2415,
    n2416, n2417, n2418, n2419, n2420, n2421,
    n2422, n2423, n2424, n2425, n2426, n2427,
    n2428, n2429, n2430, n2431, n2432, n2433,
    n2434, n2435, n2436, n2437, n2438, n2439,
    n2440, n2441, n2442, n2443, n2444, n2445,
    n2446, n2447, n2448, n2449, n2450, n2451,
    n2452, n2453, n2454, n2455, n2456, n2457,
    n2458, n2459, n2460, n2461, n2462, n2463,
    n2464, n2465, n2466, n2467, n2468, n2469,
    n2470, n2471, n2472, n2473, n2474, n2475,
    n2476, n2477, n2478, n2479, n2480, n2481,
    n2482, n2483, n2484, n2485, n2486, n2487,
    n2488, n2489, n2490, n2491, n2492, n2493,
    n2494, n2495, n2496, n2497, n2498, n2499,
    n2500, n2501, n2502, n2503, n2504, n2505,
    n2506, n2507, n2508, n2509, n2510, n2511,
    n2512, n2513, n2514, n2515, n2516, n2517,
    n2518, n2519, n2520, n2521, n2522, n2523,
    n2524, n2525, n2526, n2527, n2528, n2529,
    n2530, n2531, n2532, n2533, n2534, n2535,
    n2536, n2537, n2538, n2539, n2540, n2542,
    n2543, n2544, n2545, n2546, n2547, n2548,
    n2549, n2550, n2551, n2552, n2553, n2554,
    n2555, n2556, n2557, n2558, n2559, n2560,
    n2561, n2562, n2563, n2564, n2565, n2566,
    n2567, n2568, n2569, n2570, n2571, n2572,
    n2573, n2574, n2575, n2576, n2577, n2578,
    n2579, n2580, n2581, n2582, n2583, n2584,
    n2585, n2586, n2587, n2588, n2589, n2590,
    n2591, n2592, n2593, n2594, n2595, n2596,
    n2597, n2598, n2599, n2600, n2601, n2602,
    n2603, n2604, n2605, n2606, n2607, n2608,
    n2609, n2610, n2611, n2612, n2613, n2614,
    n2615, n2616, n2617, n2618, n2619, n2620,
    n2621, n2622, n2623, n2624, n2625, n2626,
    n2627, n2628, n2629, n2630, n2631, n2632,
    n2633, n2634, n2635, n2636, n2637, n2638,
    n2639, n2640, n2641, n2642, n2643, n2644,
    n2645, n2646, n2647, n2648, n2649, n2650,
    n2651, n2652, n2653, n2654, n2655, n2656,
    n2657, n2658, n2659, n2660, n2661, n2662,
    n2663, n2664, n2665, n2666, n2667, n2668,
    n2669, n2670, n2671, n2672, n2673, n2674,
    n2675, n2676, n2677, n2678, n2679, n2680,
    n2681, n2682, n2683, n2684, n2685, n2686,
    n2687, n2688, n2689, n2690, n2691, n2692,
    n2693, n2694, n2695, n2696, n2697, n2698,
    n2699, n2700, n2701, n2702, n2703, n2704,
    n2705, n2706, n2707, n2708, n2709, n2710,
    n2711, n2712, n2713, n2714, n2715, n2716,
    n2717, n2718, n2719, n2720, n2721, n2722,
    n2723, n2724, n2725, n2726, n2727, n2728,
    n2729, n2730, n2731, n2732, n2733, n2734,
    n2735, n2736, n2737, n2738, n2739, n2740,
    n2741, n2742, n2743, n2744, n2745, n2746,
    n2747, n2748, n2749, n2750, n2751, n2753,
    n2754, n2755, n2756, n2757, n2758, n2759,
    n2760, n2761, n2762, n2763, n2764, n2765,
    n2766, n2767, n2768, n2769, n2770, n2771,
    n2772, n2773, n2774, n2775, n2776, n2777,
    n2778, n2779, n2780, n2781, n2782, n2783,
    n2784, n2785, n2786, n2787, n2788, n2789,
    n2790, n2791, n2792, n2793, n2794, n2795,
    n2796, n2797, n2798, n2799, n2800, n2801,
    n2802, n2803, n2804, n2805, n2806, n2807,
    n2808, n2809, n2810, n2811, n2812, n2813,
    n2814, n2815, n2816, n2817, n2818, n2819,
    n2820, n2821, n2822, n2823, n2824, n2825,
    n2826, n2827, n2828, n2829, n2830, n2831,
    n2832, n2833, n2834, n2835, n2836, n2837,
    n2838, n2839, n2840, n2841, n2842, n2843,
    n2844, n2845, n2846, n2847, n2848, n2849,
    n2850, n2851, n2852, n2853, n2854, n2855,
    n2856, n2857, n2858, n2859, n2860, n2861,
    n2862, n2863, n2864, n2865, n2866, n2867,
    n2868, n2869, n2870, n2871, n2872, n2873,
    n2874, n2875, n2876, n2877, n2878, n2879,
    n2880, n2881, n2882, n2883, n2884, n2885,
    n2886, n2887, n2888, n2889, n2890, n2891,
    n2892, n2893, n2894, n2895, n2896, n2897,
    n2898, n2899, n2900, n2901, n2902, n2903,
    n2904, n2905, n2906, n2907, n2908, n2909,
    n2910, n2911, n2912, n2913, n2914, n2915,
    n2916, n2917, n2918, n2919, n2920, n2921,
    n2922, n2923, n2924, n2925, n2926, n2927,
    n2928, n2929, n2930, n2931, n2932, n2933,
    n2934, n2935, n2936, n2937, n2938, n2939,
    n2940, n2941, n2942, n2943, n2944, n2945,
    n2946, n2947, n2948, n2949, n2950, n2951,
    n2952, n2953, n2954, n2955, n2956, n2957,
    n2958, n2959, n2960, n2961, n2962, n2963,
    n2964, n2965, n2966, n2967, n2968, n2969,
    n2970, n2971, n2973, n2974, n2975, n2976,
    n2977, n2978, n2979, n2980, n2981, n2982,
    n2983, n2984, n2985, n2986, n2987, n2988,
    n2989, n2990, n2991, n2992, n2993, n2994,
    n2995, n2996, n2997, n2998, n2999, n3000,
    n3001, n3002, n3003, n3004, n3005, n3006,
    n3007, n3008, n3009, n3010, n3011, n3012,
    n3013, n3014, n3015, n3016, n3017, n3018,
    n3019, n3020, n3021, n3022, n3023, n3024,
    n3025, n3026, n3027, n3028, n3029, n3030,
    n3031, n3032, n3033, n3034, n3035, n3036,
    n3037, n3038, n3039, n3040, n3041, n3042,
    n3043, n3044, n3045, n3046, n3047, n3048,
    n3049, n3050, n3051, n3052, n3053, n3054,
    n3055, n3056, n3057, n3058, n3059, n3060,
    n3061, n3062, n3063, n3064, n3065, n3066,
    n3067, n3068, n3069, n3070, n3071, n3072,
    n3073, n3074, n3075, n3076, n3077, n3078,
    n3079, n3080, n3081, n3082, n3083, n3084,
    n3085, n3086, n3087, n3088, n3089, n3090,
    n3091, n3092, n3093, n3094, n3095, n3096,
    n3097, n3098, n3099, n3100, n3101, n3102,
    n3103, n3104, n3105, n3106, n3107, n3108,
    n3109, n3110, n3111, n3112, n3113, n3114,
    n3115, n3116, n3117, n3118, n3119, n3120,
    n3121, n3122, n3123, n3124, n3125, n3126,
    n3127, n3128, n3129, n3130, n3131, n3132,
    n3133, n3134, n3135, n3136, n3137, n3138,
    n3139, n3140, n3141, n3142, n3143, n3144,
    n3145, n3146, n3147, n3148, n3149, n3150,
    n3151, n3152, n3153, n3154, n3155, n3156,
    n3157, n3158, n3159, n3160, n3161, n3162,
    n3163, n3164, n3165, n3166, n3167, n3168,
    n3169, n3170, n3171, n3172, n3173, n3174,
    n3175, n3176, n3177, n3178, n3179, n3180,
    n3181, n3182, n3183, n3184, n3185, n3186,
    n3187, n3188, n3189, n3190, n3191, n3192,
    n3193, n3194, n3195, n3196, n3197, n3198,
    n3199, n3200, n3202, n3203, n3204, n3205,
    n3206, n3207, n3208, n3209, n3210, n3211,
    n3212, n3213, n3214, n3215, n3216, n3217,
    n3218, n3219, n3220, n3221, n3222, n3223,
    n3224, n3225, n3226, n3227, n3228, n3229,
    n3230, n3231, n3232, n3233, n3234, n3235,
    n3236, n3237, n3238, n3239, n3240, n3241,
    n3242, n3243, n3244, n3245, n3246, n3247,
    n3248, n3249, n3250, n3251, n3252, n3253,
    n3254, n3255, n3256, n3257, n3258, n3259,
    n3260, n3261, n3262, n3263, n3264, n3265,
    n3266, n3267, n3268, n3269, n3270, n3271,
    n3272, n3273, n3274, n3275, n3276, n3277,
    n3278, n3279, n3280, n3281, n3282, n3283,
    n3284, n3285, n3286, n3287, n3288, n3289,
    n3290, n3291, n3292, n3293, n3294, n3295,
    n3296, n3297, n3298, n3299, n3300, n3301,
    n3302, n3303, n3304, n3305, n3306, n3307,
    n3308, n3309, n3310, n3311, n3312, n3313,
    n3314, n3315, n3316, n3317, n3318, n3319,
    n3320, n3321, n3322, n3323, n3324, n3325,
    n3326, n3327, n3328, n3329, n3330, n3331,
    n3332, n3333, n3334, n3335, n3336, n3337,
    n3338, n3339, n3340, n3341, n3342, n3343,
    n3344, n3345, n3346, n3347, n3348, n3349,
    n3350, n3351, n3352, n3353, n3354, n3355,
    n3356, n3357, n3358, n3359, n3360, n3361,
    n3362, n3363, n3364, n3365, n3366, n3367,
    n3368, n3369, n3370, n3371, n3372, n3373,
    n3374, n3375, n3376, n3377, n3378, n3379,
    n3380, n3381, n3382, n3383, n3384, n3385,
    n3386, n3387, n3388, n3389, n3390, n3391,
    n3392, n3393, n3394, n3395, n3396, n3397,
    n3398, n3399, n3400, n3401, n3402, n3403,
    n3404, n3405, n3406, n3407, n3408, n3409,
    n3410, n3411, n3412, n3413, n3414, n3415,
    n3416, n3417, n3418, n3419, n3420, n3421,
    n3422, n3423, n3424, n3425, n3426, n3427,
    n3428, n3429, n3430, n3431, n3432, n3433,
    n3434, n3435, n3436, n3437, n3438, n3440,
    n3441, n3442, n3443, n3444, n3445, n3446,
    n3447, n3448, n3449, n3450, n3451, n3452,
    n3453, n3454, n3455, n3456, n3457, n3458,
    n3459, n3460, n3461, n3462, n3463, n3464,
    n3465, n3466, n3467, n3468, n3469, n3470,
    n3471, n3472, n3473, n3474, n3475, n3476,
    n3477, n3478, n3479, n3480, n3481, n3482,
    n3483, n3484, n3485, n3486, n3487, n3488,
    n3489, n3490, n3491, n3492, n3493, n3494,
    n3495, n3496, n3497, n3498, n3499, n3500,
    n3501, n3502, n3503, n3504, n3505, n3506,
    n3507, n3508, n3509, n3510, n3511, n3512,
    n3513, n3514, n3515, n3516, n3517, n3518,
    n3519, n3520, n3521, n3522, n3523, n3524,
    n3525, n3526, n3527, n3528, n3529, n3530,
    n3531, n3532, n3533, n3534, n3535, n3536,
    n3537, n3538, n3539, n3540, n3541, n3542,
    n3543, n3544, n3545, n3546, n3547, n3548,
    n3549, n3550, n3551, n3552, n3553, n3554,
    n3555, n3556, n3557, n3558, n3559, n3560,
    n3561, n3562, n3563, n3564, n3565, n3566,
    n3567, n3568, n3569, n3570, n3571, n3572,
    n3573, n3574, n3575, n3576, n3577, n3578,
    n3579, n3580, n3581, n3582, n3583, n3584,
    n3585, n3586, n3587, n3588, n3589, n3590,
    n3591, n3592, n3593, n3594, n3595, n3596,
    n3597, n3598, n3599, n3600, n3601, n3602,
    n3603, n3604, n3605, n3606, n3607, n3608,
    n3609, n3610, n3611, n3612, n3613, n3614,
    n3615, n3616, n3617, n3618, n3619, n3620,
    n3621, n3622, n3623, n3624, n3625, n3626,
    n3627, n3628, n3629, n3630, n3631, n3632,
    n3633, n3634, n3635, n3636, n3637, n3638,
    n3639, n3640, n3641, n3642, n3643, n3644,
    n3645, n3646, n3647, n3648, n3649, n3650,
    n3651, n3652, n3653, n3654, n3655, n3656,
    n3657, n3658, n3659, n3660, n3661, n3662,
    n3663, n3664, n3665, n3666, n3667, n3668,
    n3669, n3670, n3671, n3672, n3673, n3674,
    n3675, n3676, n3677, n3678, n3679, n3680,
    n3681, n3682, n3683, n3684, n3685, n3687,
    n3688, n3689, n3690, n3691, n3692, n3693,
    n3694, n3695, n3696, n3697, n3698, n3699,
    n3700, n3701, n3702, n3703, n3704, n3705,
    n3706, n3707, n3708, n3709, n3710, n3711,
    n3712, n3713, n3714, n3715, n3716, n3717,
    n3718, n3719, n3720, n3721, n3722, n3723,
    n3724, n3725, n3726, n3727, n3728, n3729,
    n3730, n3731, n3732, n3733, n3734, n3735,
    n3736, n3737, n3738, n3739, n3740, n3741,
    n3742, n3743, n3744, n3745, n3746, n3747,
    n3748, n3749, n3750, n3751, n3752, n3753,
    n3754, n3755, n3756, n3757, n3758, n3759,
    n3760, n3761, n3762, n3763, n3764, n3765,
    n3766, n3767, n3768, n3769, n3770, n3771,
    n3772, n3773, n3774, n3775, n3776, n3777,
    n3778, n3779, n3780, n3781, n3782, n3783,
    n3784, n3785, n3786, n3787, n3788, n3789,
    n3790, n3791, n3792, n3793, n3794, n3795,
    n3796, n3797, n3798, n3799, n3800, n3801,
    n3802, n3803, n3804, n3805, n3806, n3807,
    n3808, n3809, n3810, n3811, n3812, n3813,
    n3814, n3815, n3816, n3817, n3818, n3819,
    n3820, n3821, n3822, n3823, n3824, n3825,
    n3826, n3827, n3828, n3829, n3830, n3831,
    n3832, n3833, n3834, n3835, n3836, n3837,
    n3838, n3839, n3840, n3841, n3842, n3843,
    n3844, n3845, n3846, n3847, n3848, n3849,
    n3850, n3851, n3852, n3853, n3854, n3855,
    n3856, n3857, n3858, n3859, n3860, n3861,
    n3862, n3863, n3864, n3865, n3866, n3867,
    n3868, n3869, n3870, n3871, n3872, n3873,
    n3874, n3875, n3876, n3877, n3878, n3879,
    n3880, n3881, n3882, n3883, n3884, n3885,
    n3886, n3887, n3888, n3889, n3890, n3891,
    n3892, n3893, n3894, n3895, n3896, n3897,
    n3898, n3899, n3900, n3901, n3902, n3903,
    n3904, n3905, n3906, n3907, n3908, n3909,
    n3910, n3911, n3912, n3913, n3914, n3915,
    n3916, n3917, n3918, n3919, n3920, n3921,
    n3922, n3923, n3924, n3925, n3926, n3927,
    n3928, n3929, n3930, n3931, n3932, n3933,
    n3934, n3935, n3936, n3937, n3938, n3939,
    n3940, n3941, n3943, n3944, n3945, n3946,
    n3947, n3948, n3949, n3950, n3951, n3952,
    n3953, n3954, n3955, n3956, n3957, n3958,
    n3959, n3960, n3961, n3962, n3963, n3964,
    n3965, n3966, n3967, n3968, n3969, n3970,
    n3971, n3972, n3973, n3974, n3975, n3976,
    n3977, n3978, n3979, n3980, n3981, n3982,
    n3983, n3984, n3985, n3986, n3987, n3988,
    n3989, n3990, n3991, n3992, n3993, n3994,
    n3995, n3996, n3997, n3998, n3999, n4000,
    n4001, n4002, n4003, n4004, n4005, n4006,
    n4007, n4008, n4009, n4010, n4011, n4012,
    n4013, n4014, n4015, n4016, n4017, n4018,
    n4019, n4020, n4021, n4022, n4023, n4024,
    n4025, n4026, n4027, n4028, n4029, n4030,
    n4031, n4032, n4033, n4034, n4035, n4036,
    n4037, n4038, n4039, n4040, n4041, n4042,
    n4043, n4044, n4045, n4046, n4047, n4048,
    n4049, n4050, n4051, n4052, n4053, n4054,
    n4055, n4056, n4057, n4058, n4059, n4060,
    n4061, n4062, n4063, n4064, n4065, n4066,
    n4067, n4068, n4069, n4070, n4071, n4072,
    n4073, n4074, n4075, n4076, n4077, n4078,
    n4079, n4080, n4081, n4082, n4083, n4084,
    n4085, n4086, n4087, n4088, n4089, n4090,
    n4091, n4092, n4093, n4094, n4095, n4096,
    n4097, n4098, n4099, n4100, n4101, n4102,
    n4103, n4104, n4105, n4106, n4107, n4108,
    n4109, n4110, n4111, n4112, n4113, n4114,
    n4115, n4116, n4117, n4118, n4119, n4120,
    n4121, n4122, n4123, n4124, n4125, n4126,
    n4127, n4128, n4129, n4130, n4131, n4132,
    n4133, n4134, n4135, n4136, n4137, n4138,
    n4139, n4140, n4141, n4142, n4143, n4144,
    n4145, n4146, n4147, n4148, n4149, n4150,
    n4151, n4152, n4153, n4154, n4155, n4156,
    n4157, n4158, n4159, n4160, n4161, n4162,
    n4163, n4164, n4165, n4166, n4167, n4168,
    n4169, n4170, n4171, n4172, n4173, n4174,
    n4175, n4176, n4177, n4178, n4179, n4180,
    n4181, n4182, n4183, n4184, n4185, n4186,
    n4187, n4188, n4189, n4190, n4191, n4192,
    n4193, n4194, n4195, n4196, n4197, n4198,
    n4199, n4200, n4201, n4202, n4203, n4204,
    n4205, n4206, n4208, n4209, n4210, n4211,
    n4212, n4213, n4214, n4215, n4216, n4217,
    n4218, n4219, n4220, n4221, n4222, n4223,
    n4224, n4225, n4226, n4227, n4228, n4229,
    n4230, n4231, n4232, n4233, n4234, n4235,
    n4236, n4237, n4238, n4239, n4240, n4241,
    n4242, n4243, n4244, n4245, n4246, n4247,
    n4248, n4249, n4250, n4251, n4252, n4253,
    n4254, n4255, n4256, n4257, n4258, n4259,
    n4260, n4261, n4262, n4263, n4264, n4265,
    n4266, n4267, n4268, n4269, n4270, n4271,
    n4272, n4273, n4274, n4275, n4276, n4277,
    n4278, n4279, n4280, n4281, n4282, n4283,
    n4284, n4285, n4286, n4287, n4288, n4289,
    n4290, n4291, n4292, n4293, n4294, n4295,
    n4296, n4297, n4298, n4299, n4300, n4301,
    n4302, n4303, n4304, n4305, n4306, n4307,
    n4308, n4309, n4310, n4311, n4312, n4313,
    n4314, n4315, n4316, n4317, n4318, n4319,
    n4320, n4321, n4322, n4323, n4324, n4325,
    n4326, n4327, n4328, n4329, n4330, n4331,
    n4332, n4333, n4334, n4335, n4336, n4337,
    n4338, n4339, n4340, n4341, n4342, n4343,
    n4344, n4345, n4346, n4347, n4348, n4349,
    n4350, n4351, n4352, n4353, n4354, n4355,
    n4356, n4357, n4358, n4359, n4360, n4361,
    n4362, n4363, n4364, n4365, n4366, n4367,
    n4368, n4369, n4370, n4371, n4372, n4373,
    n4374, n4375, n4376, n4377, n4378, n4379,
    n4380, n4381, n4382, n4383, n4384, n4385,
    n4386, n4387, n4388, n4389, n4390, n4391,
    n4392, n4393, n4394, n4395, n4396, n4397,
    n4398, n4399, n4400, n4401, n4402, n4403,
    n4404, n4405, n4406, n4407, n4408, n4409,
    n4410, n4411, n4412, n4413, n4414, n4415,
    n4416, n4417, n4418, n4419, n4420, n4421,
    n4422, n4423, n4424, n4425, n4426, n4427,
    n4428, n4429, n4430, n4431, n4432, n4433,
    n4434, n4435, n4436, n4437, n4438, n4439,
    n4440, n4441, n4442, n4443, n4444, n4445,
    n4446, n4447, n4448, n4449, n4450, n4451,
    n4452, n4453, n4454, n4455, n4456, n4457,
    n4458, n4459, n4460, n4461, n4462, n4463,
    n4464, n4465, n4466, n4467, n4468, n4469,
    n4470, n4471, n4472, n4473, n4474, n4475,
    n4476, n4477, n4478, n4479, n4480, n4482,
    n4483, n4484, n4485, n4486, n4487, n4488,
    n4489, n4490, n4491, n4492, n4493, n4494,
    n4495, n4496, n4497, n4498, n4499, n4500,
    n4501, n4502, n4503, n4504, n4505, n4506,
    n4507, n4508, n4509, n4510, n4511, n4512,
    n4513, n4514, n4515, n4516, n4517, n4518,
    n4519, n4520, n4521, n4522, n4523, n4524,
    n4525, n4526, n4527, n4528, n4529, n4530,
    n4531, n4532, n4533, n4534, n4535, n4536,
    n4537, n4538, n4539, n4540, n4541, n4542,
    n4543, n4544, n4545, n4546, n4547, n4548,
    n4549, n4550, n4551, n4552, n4553, n4554,
    n4555, n4556, n4557, n4558, n4559, n4560,
    n4561, n4562, n4563, n4564, n4565, n4566,
    n4567, n4568, n4569, n4570, n4571, n4572,
    n4573, n4574, n4575, n4576, n4577, n4578,
    n4579, n4580, n4581, n4582, n4583, n4584,
    n4585, n4586, n4587, n4588, n4589, n4590,
    n4591, n4592, n4593, n4594, n4595, n4596,
    n4597, n4598, n4599, n4600, n4601, n4602,
    n4603, n4604, n4605, n4606, n4607, n4608,
    n4609, n4610, n4611, n4612, n4613, n4614,
    n4615, n4616, n4617, n4618, n4619, n4620,
    n4621, n4622, n4623, n4624, n4625, n4626,
    n4627, n4628, n4629, n4630, n4631, n4632,
    n4633, n4634, n4635, n4636, n4637, n4638,
    n4639, n4640, n4641, n4642, n4643, n4644,
    n4645, n4646, n4647, n4648, n4649, n4650,
    n4651, n4652, n4653, n4654, n4655, n4656,
    n4657, n4658, n4659, n4660, n4661, n4662,
    n4663, n4664, n4665, n4666, n4667, n4668,
    n4669, n4670, n4671, n4672, n4673, n4674,
    n4675, n4676, n4677, n4678, n4679, n4680,
    n4681, n4682, n4683, n4684, n4685, n4686,
    n4687, n4688, n4689, n4690, n4691, n4692,
    n4693, n4694, n4695, n4696, n4697, n4698,
    n4699, n4700, n4701, n4702, n4703, n4704,
    n4705, n4706, n4707, n4708, n4709, n4710,
    n4711, n4712, n4713, n4714, n4715, n4716,
    n4717, n4718, n4719, n4720, n4721, n4722,
    n4723, n4724, n4725, n4726, n4727, n4728,
    n4729, n4730, n4731, n4732, n4733, n4734,
    n4735, n4736, n4737, n4738, n4739, n4740,
    n4741, n4742, n4743, n4744, n4745, n4746,
    n4747, n4748, n4749, n4750, n4751, n4752,
    n4753, n4754, n4755, n4756, n4757, n4758,
    n4759, n4760, n4761, n4762, n4763, n4765,
    n4766, n4767, n4768, n4769, n4770, n4771,
    n4772, n4773, n4774, n4775, n4776, n4777,
    n4778, n4779, n4780, n4781, n4782, n4783,
    n4784, n4785, n4786, n4787, n4788, n4789,
    n4790, n4791, n4792, n4793, n4794, n4795,
    n4796, n4797, n4798, n4799, n4800, n4801,
    n4802, n4803, n4804, n4805, n4806, n4807,
    n4808, n4809, n4810, n4811, n4812, n4813,
    n4814, n4815, n4816, n4817, n4818, n4819,
    n4820, n4821, n4822, n4823, n4824, n4825,
    n4826, n4827, n4828, n4829, n4830, n4831,
    n4832, n4833, n4834, n4835, n4836, n4837,
    n4838, n4839, n4840, n4841, n4842, n4843,
    n4844, n4845, n4846, n4847, n4848, n4849,
    n4850, n4851, n4852, n4853, n4854, n4855,
    n4856, n4857, n4858, n4859, n4860, n4861,
    n4862, n4863, n4864, n4865, n4866, n4867,
    n4868, n4869, n4870, n4871, n4872, n4873,
    n4874, n4875, n4876, n4877, n4878, n4879,
    n4880, n4881, n4882, n4883, n4884, n4885,
    n4886, n4887, n4888, n4889, n4890, n4891,
    n4892, n4893, n4894, n4895, n4896, n4897,
    n4898, n4899, n4900, n4901, n4902, n4903,
    n4904, n4905, n4906, n4907, n4908, n4909,
    n4910, n4911, n4912, n4913, n4914, n4915,
    n4916, n4917, n4918, n4919, n4920, n4921,
    n4922, n4923, n4924, n4925, n4926, n4927,
    n4928, n4929, n4930, n4931, n4932, n4933,
    n4934, n4935, n4936, n4937, n4938, n4939,
    n4940, n4941, n4942, n4943, n4944, n4945,
    n4946, n4947, n4948, n4949, n4950, n4951,
    n4952, n4953, n4954, n4955, n4956, n4957,
    n4958, n4959, n4960, n4961, n4962, n4963,
    n4964, n4965, n4966, n4967, n4968, n4969,
    n4970, n4971, n4972, n4973, n4974, n4975,
    n4976, n4977, n4978, n4979, n4980, n4981,
    n4982, n4983, n4984, n4985, n4986, n4987,
    n4988, n4989, n4990, n4991, n4992, n4993,
    n4994, n4995, n4996, n4997, n4998, n4999,
    n5000, n5001, n5002, n5003, n5004, n5005,
    n5006, n5007, n5008, n5009, n5010, n5011,
    n5012, n5013, n5014, n5015, n5016, n5017,
    n5018, n5019, n5020, n5021, n5022, n5023,
    n5024, n5025, n5026, n5027, n5028, n5029,
    n5030, n5031, n5032, n5033, n5034, n5035,
    n5036, n5037, n5038, n5039, n5040, n5041,
    n5042, n5043, n5044, n5045, n5046, n5047,
    n5048, n5049, n5050, n5051, n5052, n5053,
    n5054, n5055, n5057, n5058, n5059, n5060,
    n5061, n5062, n5063, n5064, n5065, n5066,
    n5067, n5068, n5069, n5070, n5071, n5072,
    n5073, n5074, n5075, n5076, n5077, n5078,
    n5079, n5080, n5081, n5082, n5083, n5084,
    n5085, n5086, n5087, n5088, n5089, n5090,
    n5091, n5092, n5093, n5094, n5095, n5096,
    n5097, n5098, n5099, n5100, n5101, n5102,
    n5103, n5104, n5105, n5106, n5107, n5108,
    n5109, n5110, n5111, n5112, n5113, n5114,
    n5115, n5116, n5117, n5118, n5119, n5120,
    n5121, n5122, n5123, n5124, n5125, n5126,
    n5127, n5128, n5129, n5130, n5131, n5132,
    n5133, n5134, n5135, n5136, n5137, n5138,
    n5139, n5140, n5141, n5142, n5143, n5144,
    n5145, n5146, n5147, n5148, n5149, n5150,
    n5151, n5152, n5153, n5154, n5155, n5156,
    n5157, n5158, n5159, n5160, n5161, n5162,
    n5163, n5164, n5165, n5166, n5167, n5168,
    n5169, n5170, n5171, n5172, n5173, n5174,
    n5175, n5176, n5177, n5178, n5179, n5180,
    n5181, n5182, n5183, n5184, n5185, n5186,
    n5187, n5188, n5189, n5190, n5191, n5192,
    n5193, n5194, n5195, n5196, n5197, n5198,
    n5199, n5200, n5201, n5202, n5203, n5204,
    n5205, n5206, n5207, n5208, n5209, n5210,
    n5211, n5212, n5213, n5214, n5215, n5216,
    n5217, n5218, n5219, n5220, n5221, n5222,
    n5223, n5224, n5225, n5226, n5227, n5228,
    n5229, n5230, n5231, n5232, n5233, n5234,
    n5235, n5236, n5237, n5238, n5239, n5240,
    n5241, n5242, n5243, n5244, n5245, n5246,
    n5247, n5248, n5249, n5250, n5251, n5252,
    n5253, n5254, n5255, n5256, n5257, n5258,
    n5259, n5260, n5261, n5262, n5263, n5264,
    n5265, n5266, n5267, n5268, n5269, n5270,
    n5271, n5272, n5273, n5274, n5275, n5276,
    n5277, n5278, n5279, n5280, n5281, n5282,
    n5283, n5284, n5285, n5286, n5287, n5288,
    n5289, n5290, n5291, n5292, n5293, n5294,
    n5295, n5296, n5297, n5298, n5299, n5300,
    n5301, n5302, n5303, n5304, n5305, n5306,
    n5307, n5308, n5309, n5310, n5311, n5312,
    n5313, n5314, n5315, n5316, n5317, n5318,
    n5319, n5320, n5321, n5322, n5323, n5324,
    n5325, n5326, n5327, n5328, n5329, n5330,
    n5331, n5332, n5333, n5334, n5335, n5336,
    n5337, n5338, n5339, n5340, n5341, n5342,
    n5343, n5344, n5345, n5346, n5347, n5348,
    n5349, n5350, n5351, n5352, n5353, n5354,
    n5355, n5356, n5358, n5359, n5360, n5361,
    n5362, n5363, n5364, n5365, n5366, n5367,
    n5368, n5369, n5370, n5371, n5372, n5373,
    n5374, n5375, n5376, n5377, n5378, n5379,
    n5380, n5381, n5382, n5383, n5384, n5385,
    n5386, n5387, n5388, n5389, n5390, n5391,
    n5392, n5393, n5394, n5395, n5396, n5397,
    n5398, n5399, n5400, n5401, n5402, n5403,
    n5404, n5405, n5406, n5407, n5408, n5409,
    n5410, n5411, n5412, n5413, n5414, n5415,
    n5416, n5417, n5418, n5419, n5420, n5421,
    n5422, n5423, n5424, n5425, n5426, n5427,
    n5428, n5429, n5430, n5431, n5432, n5433,
    n5434, n5435, n5436, n5437, n5438, n5439,
    n5440, n5441, n5442, n5443, n5444, n5445,
    n5446, n5447, n5448, n5449, n5450, n5451,
    n5452, n5453, n5454, n5455, n5456, n5457,
    n5458, n5459, n5460, n5461, n5462, n5463,
    n5464, n5465, n5466, n5467, n5468, n5469,
    n5470, n5471, n5472, n5473, n5474, n5475,
    n5476, n5477, n5478, n5479, n5480, n5481,
    n5482, n5483, n5484, n5485, n5486, n5487,
    n5488, n5489, n5490, n5491, n5492, n5493,
    n5494, n5495, n5496, n5497, n5498, n5499,
    n5500, n5501, n5502, n5503, n5504, n5505,
    n5506, n5507, n5508, n5509, n5510, n5511,
    n5512, n5513, n5514, n5515, n5516, n5517,
    n5518, n5519, n5520, n5521, n5522, n5523,
    n5524, n5525, n5526, n5527, n5528, n5529,
    n5530, n5531, n5532, n5533, n5534, n5535,
    n5536, n5537, n5538, n5539, n5540, n5541,
    n5542, n5543, n5544, n5545, n5546, n5547,
    n5548, n5549, n5550, n5551, n5552, n5553,
    n5554, n5555, n5556, n5557, n5558, n5559,
    n5560, n5561, n5562, n5563, n5564, n5565,
    n5566, n5567, n5568, n5569, n5570, n5571,
    n5572, n5573, n5574, n5575, n5576, n5577,
    n5578, n5579, n5580, n5581, n5582, n5583,
    n5584, n5585, n5586, n5587, n5588, n5589,
    n5590, n5591, n5592, n5593, n5594, n5595,
    n5596, n5597, n5598, n5599, n5600, n5601,
    n5602, n5603, n5604, n5605, n5606, n5607,
    n5608, n5609, n5610, n5611, n5612, n5613,
    n5614, n5615, n5616, n5617, n5618, n5619,
    n5620, n5621, n5622, n5623, n5624, n5625,
    n5626, n5627, n5628, n5629, n5630, n5631,
    n5632, n5633, n5634, n5635, n5636, n5637,
    n5638, n5639, n5640, n5641, n5642, n5643,
    n5644, n5645, n5646, n5647, n5648, n5649,
    n5650, n5651, n5652, n5653, n5654, n5655,
    n5656, n5657, n5658, n5659, n5660, n5661,
    n5662, n5663, n5664, n5665, n5666, n5668,
    n5669, n5670, n5671, n5672, n5673, n5674,
    n5675, n5676, n5677, n5678, n5679, n5680,
    n5681, n5682, n5683, n5684, n5685, n5686,
    n5687, n5688, n5689, n5690, n5691, n5692,
    n5693, n5694, n5695, n5696, n5697, n5698,
    n5699, n5700, n5701, n5702, n5703, n5704,
    n5705, n5706, n5707, n5708, n5709, n5710,
    n5711, n5712, n5713, n5714, n5715, n5716,
    n5717, n5718, n5719, n5720, n5721, n5722,
    n5723, n5724, n5725, n5726, n5727, n5728,
    n5729, n5730, n5731, n5732, n5733, n5734,
    n5735, n5736, n5737, n5738, n5739, n5740,
    n5741, n5742, n5743, n5744, n5745, n5746,
    n5747, n5748, n5749, n5750, n5751, n5752,
    n5753, n5754, n5755, n5756, n5757, n5758,
    n5759, n5760, n5761, n5762, n5763, n5764,
    n5765, n5766, n5767, n5768, n5769, n5770,
    n5771, n5772, n5773, n5774, n5775, n5776,
    n5777, n5778, n5779, n5780, n5781, n5782,
    n5783, n5784, n5785, n5786, n5787, n5788,
    n5789, n5790, n5791, n5792, n5793, n5794,
    n5795, n5796, n5797, n5798, n5799, n5800,
    n5801, n5802, n5803, n5804, n5805, n5806,
    n5807, n5808, n5809, n5810, n5811, n5812,
    n5813, n5814, n5815, n5816, n5817, n5818,
    n5819, n5820, n5821, n5822, n5823, n5824,
    n5825, n5826, n5827, n5828, n5829, n5830,
    n5831, n5832, n5833, n5834, n5835, n5836,
    n5837, n5838, n5839, n5840, n5841, n5842,
    n5843, n5844, n5845, n5846, n5847, n5848,
    n5849, n5850, n5851, n5852, n5853, n5854,
    n5855, n5856, n5857, n5858, n5859, n5860,
    n5861, n5862, n5863, n5864, n5865, n5866,
    n5867, n5868, n5869, n5870, n5871, n5872,
    n5873, n5874, n5875, n5876, n5877, n5878,
    n5879, n5880, n5881, n5882, n5883, n5884,
    n5885, n5886, n5887, n5888, n5889, n5890,
    n5891, n5892, n5893, n5894, n5895, n5896,
    n5897, n5898, n5899, n5900, n5901, n5902,
    n5903, n5904, n5905, n5906, n5907, n5908,
    n5909, n5910, n5911, n5912, n5913, n5914,
    n5915, n5916, n5917, n5918, n5919, n5920,
    n5921, n5922, n5923, n5924, n5925, n5926,
    n5927, n5928, n5929, n5930, n5931, n5932,
    n5933, n5934, n5935, n5936, n5937, n5938,
    n5939, n5940, n5941, n5942, n5943, n5944,
    n5945, n5946, n5947, n5948, n5949, n5950,
    n5951, n5952, n5953, n5954, n5955, n5956,
    n5957, n5958, n5959, n5960, n5961, n5962,
    n5963, n5964, n5965, n5966, n5967, n5968,
    n5969, n5970, n5971, n5972, n5973, n5974,
    n5975, n5976, n5977, n5978, n5979, n5980,
    n5981, n5982, n5983, n5984, n5985, n5987,
    n5988, n5989, n5990, n5991, n5992, n5993,
    n5994, n5995, n5996, n5997, n5998, n5999,
    n6000, n6001, n6002, n6003, n6004, n6005,
    n6006, n6007, n6008, n6009, n6010, n6011,
    n6012, n6013, n6014, n6015, n6016, n6017,
    n6018, n6019, n6020, n6021, n6022, n6023,
    n6024, n6025, n6026, n6027, n6028, n6029,
    n6030, n6031, n6032, n6033, n6034, n6035,
    n6036, n6037, n6038, n6039, n6040, n6041,
    n6042, n6043, n6044, n6045, n6046, n6047,
    n6048, n6049, n6050, n6051, n6052, n6053,
    n6054, n6055, n6056, n6057, n6058, n6059,
    n6060, n6061, n6062, n6063, n6064, n6065,
    n6066, n6067, n6068, n6069, n6070, n6071,
    n6072, n6073, n6074, n6075, n6076, n6077,
    n6078, n6079, n6080, n6081, n6082, n6083,
    n6084, n6085, n6086, n6087, n6088, n6089,
    n6090, n6091, n6092, n6093, n6094, n6095,
    n6096, n6097, n6098, n6099, n6100, n6101,
    n6102, n6103, n6104, n6105, n6106, n6107,
    n6108, n6109, n6110, n6111, n6112, n6113,
    n6114, n6115, n6116, n6117, n6118, n6119,
    n6120, n6121, n6122, n6123, n6124, n6125,
    n6126, n6127, n6128, n6129, n6130, n6131,
    n6132, n6133, n6134, n6135, n6136, n6137,
    n6138, n6139, n6140, n6141, n6142, n6143,
    n6144, n6145, n6146, n6147, n6148, n6149,
    n6150, n6151, n6152, n6153, n6154, n6155,
    n6156, n6157, n6158, n6159, n6160, n6161,
    n6162, n6163, n6164, n6165, n6166, n6167,
    n6168, n6169, n6170, n6171, n6172, n6173,
    n6174, n6175, n6176, n6177, n6178, n6179,
    n6180, n6181, n6182, n6183, n6184, n6185,
    n6186, n6187, n6188, n6189, n6190, n6191,
    n6192, n6193, n6194, n6195, n6196, n6197,
    n6198, n6199, n6200, n6201, n6202, n6203,
    n6204, n6205, n6206, n6207, n6208, n6209,
    n6210, n6211, n6212, n6213, n6214, n6215,
    n6216, n6217, n6218, n6219, n6220, n6221,
    n6222, n6223, n6224, n6225, n6226, n6227,
    n6228, n6229, n6230, n6231, n6232, n6233,
    n6234, n6235, n6236, n6237, n6238, n6239,
    n6240, n6241, n6242, n6243, n6244, n6245,
    n6246, n6247, n6248, n6249, n6250, n6251,
    n6252, n6253, n6254, n6255, n6256, n6257,
    n6258, n6259, n6260, n6261, n6262, n6263,
    n6264, n6265, n6266, n6267, n6268, n6269,
    n6270, n6271, n6272, n6273, n6274, n6275,
    n6276, n6277, n6278, n6279, n6280, n6281,
    n6282, n6283, n6284, n6285, n6286, n6287,
    n6288, n6289, n6290, n6291, n6292, n6293,
    n6294, n6295, n6296, n6297, n6298, n6299,
    n6300, n6301, n6302, n6303, n6304, n6305,
    n6306, n6307, n6308, n6309, n6310, n6311,
    n6312, n6313, n6315, n6316, n6317, n6318,
    n6319, n6320, n6321, n6322, n6323, n6324,
    n6325, n6326, n6327, n6328, n6329, n6330,
    n6331, n6332, n6333, n6334, n6335, n6336,
    n6337, n6338, n6339, n6340, n6341, n6342,
    n6343, n6344, n6345, n6346, n6347, n6348,
    n6349, n6350, n6351, n6352, n6353, n6354,
    n6355, n6356, n6357, n6358, n6359, n6360,
    n6361, n6362, n6363, n6364, n6365, n6366,
    n6367, n6368, n6369, n6370, n6371, n6372,
    n6373, n6374, n6375, n6376, n6377, n6378,
    n6379, n6380, n6381, n6382, n6383, n6384,
    n6385, n6386, n6387, n6388, n6389, n6390,
    n6391, n6392, n6393, n6394, n6395, n6396,
    n6397, n6398, n6399, n6400, n6401, n6402,
    n6403, n6404, n6405, n6406, n6407, n6408,
    n6409, n6410, n6411, n6412, n6413, n6414,
    n6415, n6416, n6417, n6418, n6419, n6420,
    n6421, n6422, n6423, n6424, n6425, n6426,
    n6427, n6428, n6429, n6430, n6431, n6432,
    n6433, n6434, n6435, n6436, n6437, n6438,
    n6439, n6440, n6441, n6442, n6443, n6444,
    n6445, n6446, n6447, n6448, n6449, n6450,
    n6451, n6452, n6453, n6454, n6455, n6456,
    n6457, n6458, n6459, n6460, n6461, n6462,
    n6463, n6464, n6465, n6466, n6467, n6468,
    n6469, n6470, n6471, n6472, n6473, n6474,
    n6475, n6476, n6477, n6478, n6479, n6480,
    n6481, n6482, n6483, n6484, n6485, n6486,
    n6487, n6488, n6489, n6490, n6491, n6492,
    n6493, n6494, n6495, n6496, n6497, n6498,
    n6499, n6500, n6501, n6502, n6503, n6504,
    n6505, n6506, n6507, n6508, n6509, n6510,
    n6511, n6512, n6513, n6514, n6515, n6516,
    n6517, n6518, n6519, n6520, n6521, n6522,
    n6523, n6524, n6525, n6526, n6527, n6528,
    n6529, n6530, n6531, n6532, n6533, n6534,
    n6535, n6536, n6537, n6538, n6539, n6540,
    n6541, n6542, n6543, n6544, n6545, n6546,
    n6547, n6548, n6549, n6550, n6551, n6552,
    n6553, n6554, n6555, n6556, n6557, n6558,
    n6559, n6560, n6561, n6562, n6563, n6564,
    n6565, n6566, n6567, n6568, n6569, n6570,
    n6571, n6572, n6573, n6574, n6575, n6576,
    n6577, n6578, n6579, n6580, n6581, n6582,
    n6583, n6584, n6585, n6586, n6587, n6588,
    n6589, n6590, n6591, n6592, n6593, n6594,
    n6595, n6596, n6597, n6598, n6599, n6600,
    n6601, n6602, n6603, n6604, n6605, n6606,
    n6607, n6608, n6609, n6610, n6611, n6612,
    n6613, n6614, n6615, n6616, n6617, n6618,
    n6619, n6620, n6621, n6622, n6623, n6624,
    n6625, n6626, n6627, n6628, n6629, n6630,
    n6631, n6632, n6633, n6634, n6635, n6636,
    n6637, n6638, n6639, n6640, n6641, n6642,
    n6643, n6644, n6645, n6646, n6647, n6648,
    n6649, n6650, n6652, n6653, n6654, n6655,
    n6656, n6657, n6658, n6659, n6660, n6661,
    n6662, n6663, n6664, n6665, n6666, n6667,
    n6668, n6669, n6670, n6671, n6672, n6673,
    n6674, n6675, n6676, n6677, n6678, n6679,
    n6680, n6681, n6682, n6683, n6684, n6685,
    n6686, n6687, n6688, n6689, n6690, n6691,
    n6692, n6693, n6694, n6695, n6696, n6697,
    n6698, n6699, n6700, n6701, n6702, n6703,
    n6704, n6705, n6706, n6707, n6708, n6709,
    n6710, n6711, n6712, n6713, n6714, n6715,
    n6716, n6717, n6718, n6719, n6720, n6721,
    n6722, n6723, n6724, n6725, n6726, n6727,
    n6728, n6729, n6730, n6731, n6732, n6733,
    n6734, n6735, n6736, n6737, n6738, n6739,
    n6740, n6741, n6742, n6743, n6744, n6745,
    n6746, n6747, n6748, n6749, n6750, n6751,
    n6752, n6753, n6754, n6755, n6756, n6757,
    n6758, n6759, n6760, n6761, n6762, n6763,
    n6764, n6765, n6766, n6767, n6768, n6769,
    n6770, n6771, n6772, n6773, n6774, n6775,
    n6776, n6777, n6778, n6779, n6780, n6781,
    n6782, n6783, n6784, n6785, n6786, n6787,
    n6788, n6789, n6790, n6791, n6792, n6793,
    n6794, n6795, n6796, n6797, n6798, n6799,
    n6800, n6801, n6802, n6803, n6804, n6805,
    n6806, n6807, n6808, n6809, n6810, n6811,
    n6812, n6813, n6814, n6815, n6816, n6817,
    n6818, n6819, n6820, n6821, n6822, n6823,
    n6824, n6825, n6826, n6827, n6828, n6829,
    n6830, n6831, n6832, n6833, n6834, n6835,
    n6836, n6837, n6838, n6839, n6840, n6841,
    n6842, n6843, n6844, n6845, n6846, n6847,
    n6848, n6849, n6850, n6851, n6852, n6853,
    n6854, n6855, n6856, n6857, n6858, n6859,
    n6860, n6861, n6862, n6863, n6864, n6865,
    n6866, n6867, n6868, n6869, n6870, n6871,
    n6872, n6873, n6874, n6875, n6876, n6877,
    n6878, n6879, n6880, n6881, n6882, n6883,
    n6884, n6885, n6886, n6887, n6888, n6889,
    n6890, n6891, n6892, n6893, n6894, n6895,
    n6896, n6897, n6898, n6899, n6900, n6901,
    n6902, n6903, n6904, n6905, n6906, n6907,
    n6908, n6909, n6910, n6911, n6912, n6913,
    n6914, n6915, n6916, n6917, n6918, n6919,
    n6920, n6921, n6922, n6923, n6924, n6925,
    n6926, n6927, n6928, n6929, n6930, n6931,
    n6932, n6933, n6934, n6935, n6936, n6937,
    n6938, n6939, n6940, n6941, n6942, n6943,
    n6944, n6945, n6946, n6947, n6948, n6949,
    n6950, n6951, n6952, n6953, n6954, n6955,
    n6956, n6957, n6958, n6959, n6960, n6961,
    n6962, n6963, n6964, n6965, n6966, n6967,
    n6968, n6969, n6970, n6971, n6972, n6973,
    n6974, n6975, n6976, n6977, n6978, n6979,
    n6980, n6981, n6982, n6983, n6984, n6985,
    n6986, n6987, n6988, n6989, n6990, n6991,
    n6992, n6993, n6994, n6995, n6996, n6998,
    n6999, n7000, n7001, n7002, n7003, n7004,
    n7005, n7006, n7007, n7008, n7009, n7010,
    n7011, n7012, n7013, n7014, n7015, n7016,
    n7017, n7018, n7019, n7020, n7021, n7022,
    n7023, n7024, n7025, n7026, n7027, n7028,
    n7029, n7030, n7031, n7032, n7033, n7034,
    n7035, n7036, n7037, n7038, n7039, n7040,
    n7041, n7042, n7043, n7044, n7045, n7046,
    n7047, n7048, n7049, n7050, n7051, n7052,
    n7053, n7054, n7055, n7056, n7057, n7058,
    n7059, n7060, n7061, n7062, n7063, n7064,
    n7065, n7066, n7067, n7068, n7069, n7070,
    n7071, n7072, n7073, n7074, n7075, n7076,
    n7077, n7078, n7079, n7080, n7081, n7082,
    n7083, n7084, n7085, n7086, n7087, n7088,
    n7089, n7090, n7091, n7092, n7093, n7094,
    n7095, n7096, n7097, n7098, n7099, n7100,
    n7101, n7102, n7103, n7104, n7105, n7106,
    n7107, n7108, n7109, n7110, n7111, n7112,
    n7113, n7114, n7115, n7116, n7117, n7118,
    n7119, n7120, n7121, n7122, n7123, n7124,
    n7125, n7126, n7127, n7128, n7129, n7130,
    n7131, n7132, n7133, n7134, n7135, n7136,
    n7137, n7138, n7139, n7140, n7141, n7142,
    n7143, n7144, n7145, n7146, n7147, n7148,
    n7149, n7150, n7151, n7152, n7153, n7154,
    n7155, n7156, n7157, n7158, n7159, n7160,
    n7161, n7162, n7163, n7164, n7165, n7166,
    n7167, n7168, n7169, n7170, n7171, n7172,
    n7173, n7174, n7175, n7176, n7177, n7178,
    n7179, n7180, n7181, n7182, n7183, n7184,
    n7185, n7186, n7187, n7188, n7189, n7190,
    n7191, n7192, n7193, n7194, n7195, n7196,
    n7197, n7198, n7199, n7200, n7201, n7202,
    n7203, n7204, n7205, n7206, n7207, n7208,
    n7209, n7210, n7211, n7212, n7213, n7214,
    n7215, n7216, n7217, n7218, n7219, n7220,
    n7221, n7222, n7223, n7224, n7225, n7226,
    n7227, n7228, n7229, n7230, n7231, n7232,
    n7233, n7234, n7235, n7236, n7237, n7238,
    n7239, n7240, n7241, n7242, n7243, n7244,
    n7245, n7246, n7247, n7248, n7249, n7250,
    n7251, n7252, n7253, n7254, n7255, n7256,
    n7257, n7258, n7259, n7260, n7261, n7262,
    n7263, n7264, n7265, n7266, n7267, n7268,
    n7269, n7270, n7271, n7272, n7273, n7274,
    n7275, n7276, n7277, n7278, n7279, n7280,
    n7281, n7282, n7283, n7284, n7285, n7286,
    n7287, n7288, n7289, n7290, n7291, n7292,
    n7293, n7294, n7295, n7296, n7297, n7298,
    n7299, n7300, n7301, n7302, n7303, n7304,
    n7305, n7306, n7307, n7308, n7309, n7310,
    n7311, n7312, n7313, n7314, n7315, n7316,
    n7317, n7318, n7319, n7320, n7321, n7322,
    n7323, n7324, n7325, n7326, n7327, n7328,
    n7329, n7330, n7331, n7332, n7333, n7334,
    n7335, n7336, n7337, n7338, n7339, n7340,
    n7341, n7342, n7343, n7344, n7345, n7346,
    n7347, n7348, n7349, n7350, n7351, n7353,
    n7354, n7355, n7356, n7357, n7358, n7359,
    n7360, n7361, n7362, n7363, n7364, n7365,
    n7366, n7367, n7368, n7369, n7370, n7371,
    n7372, n7373, n7374, n7375, n7376, n7377,
    n7378, n7379, n7380, n7381, n7382, n7383,
    n7384, n7385, n7386, n7387, n7388, n7389,
    n7390, n7391, n7392, n7393, n7394, n7395,
    n7396, n7397, n7398, n7399, n7400, n7401,
    n7402, n7403, n7404, n7405, n7406, n7407,
    n7408, n7409, n7410, n7411, n7412, n7413,
    n7414, n7415, n7416, n7417, n7418, n7419,
    n7420, n7421, n7422, n7423, n7424, n7425,
    n7426, n7427, n7428, n7429, n7430, n7431,
    n7432, n7433, n7434, n7435, n7436, n7437,
    n7438, n7439, n7440, n7441, n7442, n7443,
    n7444, n7445, n7446, n7447, n7448, n7449,
    n7450, n7451, n7452, n7453, n7454, n7455,
    n7456, n7457, n7458, n7459, n7460, n7461,
    n7462, n7463, n7464, n7465, n7466, n7467,
    n7468, n7469, n7470, n7471, n7472, n7473,
    n7474, n7475, n7476, n7477, n7478, n7479,
    n7480, n7481, n7482, n7483, n7484, n7485,
    n7486, n7487, n7488, n7489, n7490, n7491,
    n7492, n7493, n7494, n7495, n7496, n7497,
    n7498, n7499, n7500, n7501, n7502, n7503,
    n7504, n7505, n7506, n7507, n7508, n7509,
    n7510, n7511, n7512, n7513, n7514, n7515,
    n7516, n7517, n7518, n7519, n7520, n7521,
    n7522, n7523, n7524, n7525, n7526, n7527,
    n7528, n7529, n7530, n7531, n7532, n7533,
    n7534, n7535, n7536, n7537, n7538, n7539,
    n7540, n7541, n7542, n7543, n7544, n7545,
    n7546, n7547, n7548, n7549, n7550, n7551,
    n7552, n7553, n7554, n7555, n7556, n7557,
    n7558, n7559, n7560, n7561, n7562, n7563,
    n7564, n7565, n7566, n7567, n7568, n7569,
    n7570, n7571, n7572, n7573, n7574, n7575,
    n7576, n7577, n7578, n7579, n7580, n7581,
    n7582, n7583, n7584, n7585, n7586, n7587,
    n7588, n7589, n7590, n7591, n7592, n7593,
    n7594, n7595, n7596, n7597, n7598, n7599,
    n7600, n7601, n7602, n7603, n7604, n7605,
    n7606, n7607, n7608, n7609, n7610, n7611,
    n7612, n7613, n7614, n7615, n7616, n7617,
    n7618, n7619, n7620, n7621, n7622, n7623,
    n7624, n7625, n7626, n7627, n7628, n7629,
    n7630, n7631, n7632, n7633, n7634, n7635,
    n7636, n7637, n7638, n7639, n7640, n7641,
    n7642, n7643, n7644, n7645, n7646, n7647,
    n7648, n7649, n7650, n7651, n7652, n7653,
    n7654, n7655, n7656, n7657, n7658, n7659,
    n7660, n7661, n7662, n7663, n7664, n7665,
    n7666, n7667, n7668, n7669, n7670, n7671,
    n7672, n7673, n7674, n7675, n7676, n7677,
    n7678, n7679, n7680, n7681, n7682, n7683,
    n7684, n7685, n7686, n7687, n7688, n7689,
    n7690, n7691, n7692, n7693, n7694, n7695,
    n7696, n7697, n7698, n7699, n7700, n7701,
    n7702, n7703, n7704, n7705, n7706, n7707,
    n7708, n7709, n7710, n7711, n7712, n7713,
    n7714, n7715, n7717, n7718, n7719, n7720,
    n7721, n7722, n7723, n7724, n7725, n7726,
    n7727, n7728, n7729, n7730, n7731, n7732,
    n7733, n7734, n7735, n7736, n7737, n7738,
    n7739, n7740, n7741, n7742, n7743, n7744,
    n7745, n7746, n7747, n7748, n7749, n7750,
    n7751, n7752, n7753, n7754, n7755, n7756,
    n7757, n7758, n7759, n7760, n7761, n7762,
    n7763, n7764, n7765, n7766, n7767, n7768,
    n7769, n7770, n7771, n7772, n7773, n7774,
    n7775, n7776, n7777, n7778, n7779, n7780,
    n7781, n7782, n7783, n7784, n7785, n7786,
    n7787, n7788, n7789, n7790, n7791, n7792,
    n7793, n7794, n7795, n7796, n7797, n7798,
    n7799, n7800, n7801, n7802, n7803, n7804,
    n7805, n7806, n7807, n7808, n7809, n7810,
    n7811, n7812, n7813, n7814, n7815, n7816,
    n7817, n7818, n7819, n7820, n7821, n7822,
    n7823, n7824, n7825, n7826, n7827, n7828,
    n7829, n7830, n7831, n7832, n7833, n7834,
    n7835, n7836, n7837, n7838, n7839, n7840,
    n7841, n7842, n7843, n7844, n7845, n7846,
    n7847, n7848, n7849, n7850, n7851, n7852,
    n7853, n7854, n7855, n7856, n7857, n7858,
    n7859, n7860, n7861, n7862, n7863, n7864,
    n7865, n7866, n7867, n7868, n7869, n7870,
    n7871, n7872, n7873, n7874, n7875, n7876,
    n7877, n7878, n7879, n7880, n7881, n7882,
    n7883, n7884, n7885, n7886, n7887, n7888,
    n7889, n7890, n7891, n7892, n7893, n7894,
    n7895, n7896, n7897, n7898, n7899, n7900,
    n7901, n7902, n7903, n7904, n7905, n7906,
    n7907, n7908, n7909, n7910, n7911, n7912,
    n7913, n7914, n7915, n7916, n7917, n7918,
    n7919, n7920, n7921, n7922, n7923, n7924,
    n7925, n7926, n7927, n7928, n7929, n7930,
    n7931, n7932, n7933, n7934, n7935, n7936,
    n7937, n7938, n7939, n7940, n7941, n7942,
    n7943, n7944, n7945, n7946, n7947, n7948,
    n7949, n7950, n7951, n7952, n7953, n7954,
    n7955, n7956, n7957, n7958, n7959, n7960,
    n7961, n7962, n7963, n7964, n7965, n7966,
    n7967, n7968, n7969, n7970, n7971, n7972,
    n7973, n7974, n7975, n7976, n7977, n7978,
    n7979, n7980, n7981, n7982, n7983, n7984,
    n7985, n7986, n7987, n7988, n7989, n7990,
    n7991, n7992, n7993, n7994, n7995, n7996,
    n7997, n7998, n7999, n8000, n8001, n8002,
    n8003, n8004, n8005, n8006, n8007, n8008,
    n8009, n8010, n8011, n8012, n8013, n8014,
    n8015, n8016, n8017, n8018, n8019, n8020,
    n8021, n8022, n8023, n8024, n8025, n8026,
    n8027, n8028, n8029, n8030, n8031, n8032,
    n8033, n8034, n8035, n8036, n8037, n8038,
    n8039, n8040, n8041, n8042, n8043, n8044,
    n8045, n8046, n8047, n8048, n8049, n8050,
    n8051, n8052, n8053, n8054, n8055, n8056,
    n8057, n8058, n8059, n8060, n8061, n8062,
    n8063, n8064, n8065, n8066, n8067, n8068,
    n8069, n8070, n8071, n8072, n8073, n8074,
    n8075, n8076, n8077, n8078, n8079, n8080,
    n8081, n8082, n8083, n8084, n8085, n8086,
    n8087, n8088, n8090, n8091, n8092, n8093,
    n8094, n8095, n8096, n8097, n8098, n8099,
    n8100, n8101, n8102, n8103, n8104, n8105,
    n8106, n8107, n8108, n8109, n8110, n8111,
    n8112, n8113, n8114, n8115, n8116, n8117,
    n8118, n8119, n8120, n8121, n8122, n8123,
    n8124, n8125, n8126, n8127, n8128, n8129,
    n8130, n8131, n8132, n8133, n8134, n8135,
    n8136, n8137, n8138, n8139, n8140, n8141,
    n8142, n8143, n8144, n8145, n8146, n8147,
    n8148, n8149, n8150, n8151, n8152, n8153,
    n8154, n8155, n8156, n8157, n8158, n8159,
    n8160, n8161, n8162, n8163, n8164, n8165,
    n8166, n8167, n8168, n8169, n8170, n8171,
    n8172, n8173, n8174, n8175, n8176, n8177,
    n8178, n8179, n8180, n8181, n8182, n8183,
    n8184, n8185, n8186, n8187, n8188, n8189,
    n8190, n8191, n8192, n8193, n8194, n8195,
    n8196, n8197, n8198, n8199, n8200, n8201,
    n8202, n8203, n8204, n8205, n8206, n8207,
    n8208, n8209, n8210, n8211, n8212, n8213,
    n8214, n8215, n8216, n8217, n8218, n8219,
    n8220, n8221, n8222, n8223, n8224, n8225,
    n8226, n8227, n8228, n8229, n8230, n8231,
    n8232, n8233, n8234, n8235, n8236, n8237,
    n8238, n8239, n8240, n8241, n8242, n8243,
    n8244, n8245, n8246, n8247, n8248, n8249,
    n8250, n8251, n8252, n8253, n8254, n8255,
    n8256, n8257, n8258, n8259, n8260, n8261,
    n8262, n8263, n8264, n8265, n8266, n8267,
    n8268, n8269, n8270, n8271, n8272, n8273,
    n8274, n8275, n8276, n8277, n8278, n8279,
    n8280, n8281, n8282, n8283, n8284, n8285,
    n8286, n8287, n8288, n8289, n8290, n8291,
    n8292, n8293, n8294, n8295, n8296, n8297,
    n8298, n8299, n8300, n8301, n8302, n8303,
    n8304, n8305, n8306, n8307, n8308, n8309,
    n8310, n8311, n8312, n8313, n8314, n8315,
    n8316, n8317, n8318, n8319, n8320, n8321,
    n8322, n8323, n8324, n8325, n8326, n8327,
    n8328, n8329, n8330, n8331, n8332, n8333,
    n8334, n8335, n8336, n8337, n8338, n8339,
    n8340, n8341, n8342, n8343, n8344, n8345,
    n8346, n8347, n8348, n8349, n8350, n8351,
    n8352, n8353, n8354, n8355, n8356, n8357,
    n8358, n8359, n8360, n8361, n8362, n8363,
    n8364, n8365, n8366, n8367, n8368, n8369,
    n8370, n8371, n8372, n8373, n8374, n8375,
    n8376, n8377, n8378, n8379, n8380, n8381,
    n8382, n8383, n8384, n8385, n8386, n8387,
    n8388, n8389, n8390, n8391, n8392, n8393,
    n8394, n8395, n8396, n8397, n8398, n8399,
    n8400, n8401, n8402, n8403, n8404, n8405,
    n8406, n8407, n8408, n8409, n8410, n8411,
    n8412, n8413, n8414, n8415, n8416, n8417,
    n8418, n8419, n8420, n8421, n8422, n8423,
    n8424, n8425, n8426, n8427, n8428, n8429,
    n8430, n8431, n8432, n8433, n8434, n8435,
    n8436, n8437, n8438, n8439, n8440, n8441,
    n8442, n8443, n8444, n8445, n8446, n8447,
    n8448, n8449, n8450, n8451, n8452, n8453,
    n8454, n8455, n8456, n8457, n8458, n8459,
    n8460, n8461, n8462, n8463, n8464, n8465,
    n8466, n8467, n8468, n8469, n8470, n8472,
    n8473, n8474, n8475, n8476, n8477, n8478,
    n8479, n8480, n8481, n8482, n8483, n8484,
    n8485, n8486, n8487, n8488, n8489, n8490,
    n8491, n8492, n8493, n8494, n8495, n8496,
    n8497, n8498, n8499, n8500, n8501, n8502,
    n8503, n8504, n8505, n8506, n8507, n8508,
    n8509, n8510, n8511, n8512, n8513, n8514,
    n8515, n8516, n8517, n8518, n8519, n8520,
    n8521, n8522, n8523, n8524, n8525, n8526,
    n8527, n8528, n8529, n8530, n8531, n8532,
    n8533, n8534, n8535, n8536, n8537, n8538,
    n8539, n8540, n8541, n8542, n8543, n8544,
    n8545, n8546, n8547, n8548, n8549, n8550,
    n8551, n8552, n8553, n8554, n8555, n8556,
    n8557, n8558, n8559, n8560, n8561, n8562,
    n8563, n8564, n8565, n8566, n8567, n8568,
    n8569, n8570, n8571, n8572, n8573, n8574,
    n8575, n8576, n8577, n8578, n8579, n8580,
    n8581, n8582, n8583, n8584, n8585, n8586,
    n8587, n8588, n8589, n8590, n8591, n8592,
    n8593, n8594, n8595, n8596, n8597, n8598,
    n8599, n8600, n8601, n8602, n8603, n8604,
    n8605, n8606, n8607, n8608, n8609, n8610,
    n8611, n8612, n8613, n8614, n8615, n8616,
    n8617, n8618, n8619, n8620, n8621, n8622,
    n8623, n8624, n8625, n8626, n8627, n8628,
    n8629, n8630, n8631, n8632, n8633, n8634,
    n8635, n8636, n8637, n8638, n8639, n8640,
    n8641, n8642, n8643, n8644, n8645, n8646,
    n8647, n8648, n8649, n8650, n8651, n8652,
    n8653, n8654, n8655, n8656, n8657, n8658,
    n8659, n8660, n8661, n8662, n8663, n8664,
    n8665, n8666, n8667, n8668, n8669, n8670,
    n8671, n8672, n8673, n8674, n8675, n8676,
    n8677, n8678, n8679, n8680, n8681, n8682,
    n8683, n8684, n8685, n8686, n8687, n8688,
    n8689, n8690, n8691, n8692, n8693, n8694,
    n8695, n8696, n8697, n8698, n8699, n8700,
    n8701, n8702, n8703, n8704, n8705, n8706,
    n8707, n8708, n8709, n8710, n8711, n8712,
    n8713, n8714, n8715, n8716, n8717, n8718,
    n8719, n8720, n8721, n8722, n8723, n8724,
    n8725, n8726, n8727, n8728, n8729, n8730,
    n8731, n8732, n8733, n8734, n8735, n8736,
    n8737, n8738, n8739, n8740, n8741, n8742,
    n8743, n8744, n8745, n8746, n8747, n8748,
    n8749, n8750, n8751, n8752, n8753, n8754,
    n8755, n8756, n8757, n8758, n8759, n8760,
    n8761, n8762, n8763, n8764, n8765, n8766,
    n8767, n8768, n8769, n8770, n8771, n8772,
    n8773, n8774, n8775, n8776, n8777, n8778,
    n8779, n8780, n8781, n8782, n8783, n8784,
    n8785, n8786, n8787, n8788, n8789, n8790,
    n8791, n8792, n8793, n8794, n8795, n8796,
    n8797, n8798, n8799, n8800, n8801, n8802,
    n8803, n8804, n8805, n8806, n8807, n8808,
    n8809, n8810, n8811, n8812, n8813, n8814,
    n8815, n8816, n8817, n8818, n8819, n8820,
    n8821, n8822, n8823, n8824, n8825, n8826,
    n8827, n8828, n8829, n8830, n8831, n8832,
    n8833, n8834, n8835, n8836, n8837, n8838,
    n8839, n8840, n8841, n8842, n8843, n8844,
    n8845, n8846, n8847, n8848, n8849, n8850,
    n8851, n8852, n8853, n8854, n8855, n8856,
    n8857, n8858, n8859, n8860, n8861, n8863,
    n8864, n8865, n8866, n8867, n8868, n8869,
    n8870, n8871, n8872, n8873, n8874, n8875,
    n8876, n8877, n8878, n8879, n8880, n8881,
    n8882, n8883, n8884, n8885, n8886, n8887,
    n8888, n8889, n8890, n8891, n8892, n8893,
    n8894, n8895, n8896, n8897, n8898, n8899,
    n8900, n8901, n8902, n8903, n8904, n8905,
    n8906, n8907, n8908, n8909, n8910, n8911,
    n8912, n8913, n8914, n8915, n8916, n8917,
    n8918, n8919, n8920, n8921, n8922, n8923,
    n8924, n8925, n8926, n8927, n8928, n8929,
    n8930, n8931, n8932, n8933, n8934, n8935,
    n8936, n8937, n8938, n8939, n8940, n8941,
    n8942, n8943, n8944, n8945, n8946, n8947,
    n8948, n8949, n8950, n8951, n8952, n8953,
    n8954, n8955, n8956, n8957, n8958, n8959,
    n8960, n8961, n8962, n8963, n8964, n8965,
    n8966, n8967, n8968, n8969, n8970, n8971,
    n8972, n8973, n8974, n8975, n8976, n8977,
    n8978, n8979, n8980, n8981, n8982, n8983,
    n8984, n8985, n8986, n8987, n8988, n8989,
    n8990, n8991, n8992, n8993, n8994, n8995,
    n8996, n8997, n8998, n8999, n9000, n9001,
    n9002, n9003, n9004, n9005, n9006, n9007,
    n9008, n9009, n9010, n9011, n9012, n9013,
    n9014, n9015, n9016, n9017, n9018, n9019,
    n9020, n9021, n9022, n9023, n9024, n9025,
    n9026, n9027, n9028, n9029, n9030, n9031,
    n9032, n9033, n9034, n9035, n9036, n9037,
    n9038, n9039, n9040, n9041, n9042, n9043,
    n9044, n9045, n9046, n9047, n9048, n9049,
    n9050, n9051, n9052, n9053, n9054, n9055,
    n9056, n9057, n9058, n9059, n9060, n9061,
    n9062, n9063, n9064, n9065, n9066, n9067,
    n9068, n9069, n9070, n9071, n9072, n9073,
    n9074, n9075, n9076, n9077, n9078, n9079,
    n9080, n9081, n9082, n9083, n9084, n9085,
    n9086, n9087, n9088, n9089, n9090, n9091,
    n9092, n9093, n9094, n9095, n9096, n9097,
    n9098, n9099, n9100, n9101, n9102, n9103,
    n9104, n9105, n9106, n9107, n9108, n9109,
    n9110, n9111, n9112, n9113, n9114, n9115,
    n9116, n9117, n9118, n9119, n9120, n9121,
    n9122, n9123, n9124, n9125, n9126, n9127,
    n9128, n9129, n9130, n9131, n9132, n9133,
    n9134, n9135, n9136, n9137, n9138, n9139,
    n9140, n9141, n9142, n9143, n9144, n9145,
    n9146, n9147, n9148, n9149, n9150, n9151,
    n9152, n9153, n9154, n9155, n9156, n9157,
    n9158, n9159, n9160, n9161, n9162, n9163,
    n9164, n9165, n9166, n9167, n9168, n9169,
    n9170, n9171, n9172, n9173, n9174, n9175,
    n9176, n9177, n9178, n9179, n9180, n9181,
    n9182, n9183, n9184, n9185, n9186, n9187,
    n9188, n9189, n9190, n9191, n9192, n9193,
    n9194, n9195, n9196, n9197, n9198, n9199,
    n9200, n9201, n9202, n9203, n9204, n9205,
    n9206, n9207, n9208, n9209, n9210, n9211,
    n9212, n9213, n9214, n9215, n9216, n9217,
    n9218, n9219, n9220, n9221, n9222, n9223,
    n9224, n9225, n9226, n9227, n9228, n9229,
    n9230, n9231, n9232, n9233, n9234, n9235,
    n9236, n9237, n9238, n9239, n9240, n9241,
    n9242, n9243, n9244, n9245, n9246, n9247,
    n9248, n9249, n9250, n9251, n9252, n9253,
    n9254, n9255, n9256, n9257, n9258, n9259,
    n9260, n9261, n9263, n9264, n9265, n9266,
    n9267, n9268, n9269, n9270, n9271, n9272,
    n9273, n9274, n9275, n9276, n9277, n9278,
    n9279, n9280, n9281, n9282, n9283, n9284,
    n9285, n9286, n9287, n9288, n9289, n9290,
    n9291, n9292, n9293, n9294, n9295, n9296,
    n9297, n9298, n9299, n9300, n9301, n9302,
    n9303, n9304, n9305, n9306, n9307, n9308,
    n9309, n9310, n9311, n9312, n9313, n9314,
    n9315, n9316, n9317, n9318, n9319, n9320,
    n9321, n9322, n9323, n9324, n9325, n9326,
    n9327, n9328, n9329, n9330, n9331, n9332,
    n9333, n9334, n9335, n9336, n9337, n9338,
    n9339, n9340, n9341, n9342, n9343, n9344,
    n9345, n9346, n9347, n9348, n9349, n9350,
    n9351, n9352, n9353, n9354, n9355, n9356,
    n9357, n9358, n9359, n9360, n9361, n9362,
    n9363, n9364, n9365, n9366, n9367, n9368,
    n9369, n9370, n9371, n9372, n9373, n9374,
    n9375, n9376, n9377, n9378, n9379, n9380,
    n9381, n9382, n9383, n9384, n9385, n9386,
    n9387, n9388, n9389, n9390, n9391, n9392,
    n9393, n9394, n9395, n9396, n9397, n9398,
    n9399, n9400, n9401, n9402, n9403, n9404,
    n9405, n9406, n9407, n9408, n9409, n9410,
    n9411, n9412, n9413, n9414, n9415, n9416,
    n9417, n9418, n9419, n9420, n9421, n9422,
    n9423, n9424, n9425, n9426, n9427, n9428,
    n9429, n9430, n9431, n9432, n9433, n9434,
    n9435, n9436, n9437, n9438, n9439, n9440,
    n9441, n9442, n9443, n9444, n9445, n9446,
    n9447, n9448, n9449, n9450, n9451, n9452,
    n9453, n9454, n9455, n9456, n9457, n9458,
    n9459, n9460, n9461, n9462, n9463, n9464,
    n9465, n9466, n9467, n9468, n9469, n9470,
    n9471, n9472, n9473, n9474, n9475, n9476,
    n9477, n9478, n9479, n9480, n9481, n9482,
    n9483, n9484, n9485, n9486, n9487, n9488,
    n9489, n9490, n9491, n9492, n9493, n9494,
    n9495, n9496, n9497, n9498, n9499, n9500,
    n9501, n9502, n9503, n9504, n9505, n9506,
    n9507, n9508, n9509, n9510, n9511, n9512,
    n9513, n9514, n9515, n9516, n9517, n9518,
    n9519, n9520, n9521, n9522, n9523, n9524,
    n9525, n9526, n9527, n9528, n9529, n9530,
    n9531, n9532, n9533, n9534, n9535, n9536,
    n9537, n9538, n9539, n9540, n9541, n9542,
    n9543, n9544, n9545, n9546, n9547, n9548,
    n9549, n9550, n9551, n9552, n9553, n9554,
    n9555, n9556, n9557, n9558, n9559, n9560,
    n9561, n9562, n9563, n9564, n9565, n9566,
    n9567, n9568, n9569, n9570, n9571, n9572,
    n9573, n9574, n9575, n9576, n9577, n9578,
    n9579, n9580, n9581, n9582, n9583, n9584,
    n9585, n9586, n9587, n9588, n9589, n9590,
    n9591, n9592, n9593, n9594, n9595, n9596,
    n9597, n9598, n9599, n9600, n9601, n9602,
    n9603, n9604, n9605, n9606, n9607, n9608,
    n9609, n9610, n9611, n9612, n9613, n9614,
    n9615, n9616, n9617, n9618, n9619, n9620,
    n9621, n9622, n9623, n9624, n9625, n9626,
    n9627, n9628, n9629, n9630, n9631, n9632,
    n9633, n9634, n9635, n9636, n9637, n9638,
    n9639, n9640, n9641, n9642, n9643, n9644,
    n9645, n9646, n9647, n9648, n9649, n9650,
    n9651, n9652, n9653, n9654, n9655, n9656,
    n9657, n9658, n9659, n9660, n9661, n9662,
    n9663, n9664, n9665, n9666, n9667, n9668,
    n9669, n9670, n9672, n9673, n9674, n9675,
    n9676, n9677, n9678, n9679, n9680, n9681,
    n9682, n9683, n9684, n9685, n9686, n9687,
    n9688, n9689, n9690, n9691, n9692, n9693,
    n9694, n9695, n9696, n9697, n9698, n9699,
    n9700, n9701, n9702, n9703, n9704, n9705,
    n9706, n9707, n9708, n9709, n9710, n9711,
    n9712, n9713, n9714, n9715, n9716, n9717,
    n9718, n9719, n9720, n9721, n9722, n9723,
    n9724, n9725, n9726, n9727, n9728, n9729,
    n9730, n9731, n9732, n9733, n9734, n9735,
    n9736, n9737, n9738, n9739, n9740, n9741,
    n9742, n9743, n9744, n9745, n9746, n9747,
    n9748, n9749, n9750, n9751, n9752, n9753,
    n9754, n9755, n9756, n9757, n9758, n9759,
    n9760, n9761, n9762, n9763, n9764, n9765,
    n9766, n9767, n9768, n9769, n9770, n9771,
    n9772, n9773, n9774, n9775, n9776, n9777,
    n9778, n9779, n9780, n9781, n9782, n9783,
    n9784, n9785, n9786, n9787, n9788, n9789,
    n9790, n9791, n9792, n9793, n9794, n9795,
    n9796, n9797, n9798, n9799, n9800, n9801,
    n9802, n9803, n9804, n9805, n9806, n9807,
    n9808, n9809, n9810, n9811, n9812, n9813,
    n9814, n9815, n9816, n9817, n9818, n9819,
    n9820, n9821, n9822, n9823, n9824, n9825,
    n9826, n9827, n9828, n9829, n9830, n9831,
    n9832, n9833, n9834, n9835, n9836, n9837,
    n9838, n9839, n9840, n9841, n9842, n9843,
    n9844, n9845, n9846, n9847, n9848, n9849,
    n9850, n9851, n9852, n9853, n9854, n9855,
    n9856, n9857, n9858, n9859, n9860, n9861,
    n9862, n9863, n9864, n9865, n9866, n9867,
    n9868, n9869, n9870, n9871, n9872, n9873,
    n9874, n9875, n9876, n9877, n9878, n9879,
    n9880, n9881, n9882, n9883, n9884, n9885,
    n9886, n9887, n9888, n9889, n9890, n9891,
    n9892, n9893, n9894, n9895, n9896, n9897,
    n9898, n9899, n9900, n9901, n9902, n9903,
    n9904, n9905, n9906, n9907, n9908, n9909,
    n9910, n9911, n9912, n9913, n9914, n9915,
    n9916, n9917, n9918, n9919, n9920, n9921,
    n9922, n9923, n9924, n9925, n9926, n9927,
    n9928, n9929, n9930, n9931, n9932, n9933,
    n9934, n9935, n9936, n9937, n9938, n9939,
    n9940, n9941, n9942, n9943, n9944, n9945,
    n9946, n9947, n9948, n9949, n9950, n9951,
    n9952, n9953, n9954, n9955, n9956, n9957,
    n9958, n9959, n9960, n9961, n9962, n9963,
    n9964, n9965, n9966, n9967, n9968, n9969,
    n9970, n9971, n9972, n9973, n9974, n9975,
    n9976, n9977, n9978, n9979, n9980, n9981,
    n9982, n9983, n9984, n9985, n9986, n9987,
    n9988, n9989, n9990, n9991, n9992, n9993,
    n9994, n9995, n9996, n9997, n9998, n9999,
    n10000, n10001, n10002, n10003, n10004, n10005,
    n10006, n10007, n10008, n10009, n10010, n10011,
    n10012, n10013, n10014, n10015, n10016, n10017,
    n10018, n10019, n10020, n10021, n10022, n10023,
    n10024, n10025, n10026, n10027, n10028, n10029,
    n10030, n10031, n10032, n10033, n10034, n10035,
    n10036, n10037, n10038, n10039, n10040, n10041,
    n10042, n10043, n10044, n10045, n10046, n10047,
    n10048, n10049, n10050, n10051, n10052, n10053,
    n10054, n10055, n10056, n10057, n10058, n10059,
    n10060, n10061, n10062, n10063, n10064, n10065,
    n10066, n10067, n10068, n10069, n10070, n10071,
    n10072, n10073, n10074, n10075, n10076, n10077,
    n10078, n10079, n10080, n10081, n10082, n10083,
    n10084, n10085, n10086, n10087, n10088, n10090,
    n10091, n10092, n10093, n10094, n10095, n10096,
    n10097, n10098, n10099, n10100, n10101, n10102,
    n10103, n10104, n10105, n10106, n10107, n10108,
    n10109, n10110, n10111, n10112, n10113, n10114,
    n10115, n10116, n10117, n10118, n10119, n10120,
    n10121, n10122, n10123, n10124, n10125, n10126,
    n10127, n10128, n10129, n10130, n10131, n10132,
    n10133, n10134, n10135, n10136, n10137, n10138,
    n10139, n10140, n10141, n10142, n10143, n10144,
    n10145, n10146, n10147, n10148, n10149, n10150,
    n10151, n10152, n10153, n10154, n10155, n10156,
    n10157, n10158, n10159, n10160, n10161, n10162,
    n10163, n10164, n10165, n10166, n10167, n10168,
    n10169, n10170, n10171, n10172, n10173, n10174,
    n10175, n10176, n10177, n10178, n10179, n10180,
    n10181, n10182, n10183, n10184, n10185, n10186,
    n10187, n10188, n10189, n10190, n10191, n10192,
    n10193, n10194, n10195, n10196, n10197, n10198,
    n10199, n10200, n10201, n10202, n10203, n10204,
    n10205, n10206, n10207, n10208, n10209, n10210,
    n10211, n10212, n10213, n10214, n10215, n10216,
    n10217, n10218, n10219, n10220, n10221, n10222,
    n10223, n10224, n10225, n10226, n10227, n10228,
    n10229, n10230, n10231, n10232, n10233, n10234,
    n10235, n10236, n10237, n10238, n10239, n10240,
    n10241, n10242, n10243, n10244, n10245, n10246,
    n10247, n10248, n10249, n10250, n10251, n10252,
    n10253, n10254, n10255, n10256, n10257, n10258,
    n10259, n10260, n10261, n10262, n10263, n10264,
    n10265, n10266, n10267, n10268, n10269, n10270,
    n10271, n10272, n10273, n10274, n10275, n10276,
    n10277, n10278, n10279, n10280, n10281, n10282,
    n10283, n10284, n10285, n10286, n10287, n10288,
    n10289, n10290, n10291, n10292, n10293, n10294,
    n10295, n10296, n10297, n10298, n10299, n10300,
    n10301, n10302, n10303, n10304, n10305, n10306,
    n10307, n10308, n10309, n10310, n10311, n10312,
    n10313, n10314, n10315, n10316, n10317, n10318,
    n10319, n10320, n10321, n10322, n10323, n10324,
    n10325, n10326, n10327, n10328, n10329, n10330,
    n10331, n10332, n10333, n10334, n10335, n10336,
    n10337, n10338, n10339, n10340, n10341, n10342,
    n10343, n10344, n10345, n10346, n10347, n10348,
    n10349, n10350, n10351, n10352, n10353, n10354,
    n10355, n10356, n10357, n10358, n10359, n10360,
    n10361, n10362, n10363, n10364, n10365, n10366,
    n10367, n10368, n10369, n10370, n10371, n10372,
    n10373, n10374, n10375, n10376, n10377, n10378,
    n10379, n10380, n10381, n10382, n10383, n10384,
    n10385, n10386, n10387, n10388, n10389, n10390,
    n10391, n10392, n10393, n10394, n10395, n10396,
    n10397, n10398, n10399, n10400, n10401, n10402,
    n10403, n10404, n10405, n10406, n10407, n10408,
    n10409, n10410, n10411, n10412, n10413, n10414,
    n10415, n10416, n10417, n10418, n10419, n10420,
    n10421, n10422, n10423, n10424, n10425, n10426,
    n10427, n10428, n10429, n10430, n10431, n10432,
    n10433, n10434, n10435, n10436, n10437, n10438,
    n10439, n10440, n10441, n10442, n10443, n10444,
    n10445, n10446, n10447, n10448, n10449, n10450,
    n10451, n10452, n10453, n10454, n10455, n10456,
    n10457, n10458, n10459, n10460, n10461, n10462,
    n10463, n10464, n10465, n10466, n10467, n10468,
    n10469, n10470, n10471, n10472, n10473, n10474,
    n10475, n10476, n10477, n10478, n10479, n10480,
    n10481, n10482, n10483, n10484, n10485, n10486,
    n10487, n10488, n10489, n10490, n10491, n10492,
    n10493, n10494, n10495, n10496, n10497, n10498,
    n10499, n10500, n10501, n10502, n10503, n10504,
    n10505, n10506, n10507, n10508, n10509, n10510,
    n10511, n10512, n10513, n10514, n10515, n10517,
    n10518, n10519, n10520, n10521, n10522, n10523,
    n10524, n10525, n10526, n10527, n10528, n10529,
    n10530, n10531, n10532, n10533, n10534, n10535,
    n10536, n10537, n10538, n10539, n10540, n10541,
    n10542, n10543, n10544, n10545, n10546, n10547,
    n10548, n10549, n10550, n10551, n10552, n10553,
    n10554, n10555, n10556, n10557, n10558, n10559,
    n10560, n10561, n10562, n10563, n10564, n10565,
    n10566, n10567, n10568, n10569, n10570, n10571,
    n10572, n10573, n10574, n10575, n10576, n10577,
    n10578, n10579, n10580, n10581, n10582, n10583,
    n10584, n10585, n10586, n10587, n10588, n10589,
    n10590, n10591, n10592, n10593, n10594, n10595,
    n10596, n10597, n10598, n10599, n10600, n10601,
    n10602, n10603, n10604, n10605, n10606, n10607,
    n10608, n10609, n10610, n10611, n10612, n10613,
    n10614, n10615, n10616, n10617, n10618, n10619,
    n10620, n10621, n10622, n10623, n10624, n10625,
    n10626, n10627, n10628, n10629, n10630, n10631,
    n10632, n10633, n10634, n10635, n10636, n10637,
    n10638, n10639, n10640, n10641, n10642, n10643,
    n10644, n10645, n10646, n10647, n10648, n10649,
    n10650, n10651, n10652, n10653, n10654, n10655,
    n10656, n10657, n10658, n10659, n10660, n10661,
    n10662, n10663, n10664, n10665, n10666, n10667,
    n10668, n10669, n10670, n10671, n10672, n10673,
    n10674, n10675, n10676, n10677, n10678, n10679,
    n10680, n10681, n10682, n10683, n10684, n10685,
    n10686, n10687, n10688, n10689, n10690, n10691,
    n10692, n10693, n10694, n10695, n10696, n10697,
    n10698, n10699, n10700, n10701, n10702, n10703,
    n10704, n10705, n10706, n10707, n10708, n10709,
    n10710, n10711, n10712, n10713, n10714, n10715,
    n10716, n10717, n10718, n10719, n10720, n10721,
    n10722, n10723, n10724, n10725, n10726, n10727,
    n10728, n10729, n10730, n10731, n10732, n10733,
    n10734, n10735, n10736, n10737, n10738, n10739,
    n10740, n10741, n10742, n10743, n10744, n10745,
    n10746, n10747, n10748, n10749, n10750, n10751,
    n10752, n10753, n10754, n10755, n10756, n10757,
    n10758, n10759, n10760, n10761, n10762, n10763,
    n10764, n10765, n10766, n10767, n10768, n10769,
    n10770, n10771, n10772, n10773, n10774, n10775,
    n10776, n10777, n10778, n10779, n10780, n10781,
    n10782, n10783, n10784, n10785, n10786, n10787,
    n10788, n10789, n10790, n10791, n10792, n10793,
    n10794, n10795, n10796, n10797, n10798, n10799,
    n10800, n10801, n10802, n10803, n10804, n10805,
    n10806, n10807, n10808, n10809, n10810, n10811,
    n10812, n10813, n10814, n10815, n10816, n10817,
    n10818, n10819, n10820, n10821, n10822, n10823,
    n10824, n10825, n10826, n10827, n10828, n10829,
    n10830, n10831, n10832, n10833, n10834, n10835,
    n10836, n10837, n10838, n10839, n10840, n10841,
    n10842, n10843, n10844, n10845, n10846, n10847,
    n10848, n10849, n10850, n10851, n10852, n10853,
    n10854, n10855, n10856, n10857, n10858, n10859,
    n10860, n10861, n10862, n10863, n10864, n10865,
    n10866, n10867, n10868, n10869, n10870, n10871,
    n10872, n10873, n10874, n10875, n10876, n10877,
    n10878, n10879, n10880, n10881, n10882, n10883,
    n10884, n10885, n10886, n10887, n10888, n10889,
    n10890, n10891, n10892, n10893, n10894, n10895,
    n10896, n10897, n10898, n10899, n10900, n10901,
    n10902, n10903, n10904, n10905, n10906, n10907,
    n10908, n10909, n10910, n10911, n10912, n10913,
    n10914, n10915, n10916, n10917, n10918, n10919,
    n10920, n10921, n10922, n10923, n10924, n10925,
    n10926, n10927, n10928, n10929, n10930, n10931,
    n10932, n10933, n10934, n10935, n10936, n10937,
    n10938, n10939, n10940, n10941, n10942, n10943,
    n10944, n10945, n10946, n10947, n10948, n10949,
    n10950, n10951, n10953, n10954, n10955, n10956,
    n10957, n10958, n10959, n10960, n10961, n10962,
    n10963, n10964, n10965, n10966, n10967, n10968,
    n10969, n10970, n10971, n10972, n10973, n10974,
    n10975, n10976, n10977, n10978, n10979, n10980,
    n10981, n10982, n10983, n10984, n10985, n10986,
    n10987, n10988, n10989, n10990, n10991, n10992,
    n10993, n10994, n10995, n10996, n10997, n10998,
    n10999, n11000, n11001, n11002, n11003, n11004,
    n11005, n11006, n11007, n11008, n11009, n11010,
    n11011, n11012, n11013, n11014, n11015, n11016,
    n11017, n11018, n11019, n11020, n11021, n11022,
    n11023, n11024, n11025, n11026, n11027, n11028,
    n11029, n11030, n11031, n11032, n11033, n11034,
    n11035, n11036, n11037, n11038, n11039, n11040,
    n11041, n11042, n11043, n11044, n11045, n11046,
    n11047, n11048, n11049, n11050, n11051, n11052,
    n11053, n11054, n11055, n11056, n11057, n11058,
    n11059, n11060, n11061, n11062, n11063, n11064,
    n11065, n11066, n11067, n11068, n11069, n11070,
    n11071, n11072, n11073, n11074, n11075, n11076,
    n11077, n11078, n11079, n11080, n11081, n11082,
    n11083, n11084, n11085, n11086, n11087, n11088,
    n11089, n11090, n11091, n11092, n11093, n11094,
    n11095, n11096, n11097, n11098, n11099, n11100,
    n11101, n11102, n11103, n11104, n11105, n11106,
    n11107, n11108, n11109, n11110, n11111, n11112,
    n11113, n11114, n11115, n11116, n11117, n11118,
    n11119, n11120, n11121, n11122, n11123, n11124,
    n11125, n11126, n11127, n11128, n11129, n11130,
    n11131, n11132, n11133, n11134, n11135, n11136,
    n11137, n11138, n11139, n11140, n11141, n11142,
    n11143, n11144, n11145, n11146, n11147, n11148,
    n11149, n11150, n11151, n11152, n11153, n11154,
    n11155, n11156, n11157, n11158, n11159, n11160,
    n11161, n11162, n11163, n11164, n11165, n11166,
    n11167, n11168, n11169, n11170, n11171, n11172,
    n11173, n11174, n11175, n11176, n11177, n11178,
    n11179, n11180, n11181, n11182, n11183, n11184,
    n11185, n11186, n11187, n11188, n11189, n11190,
    n11191, n11192, n11193, n11194, n11195, n11196,
    n11197, n11198, n11199, n11200, n11201, n11202,
    n11203, n11204, n11205, n11206, n11207, n11208,
    n11209, n11210, n11211, n11212, n11213, n11214,
    n11215, n11216, n11217, n11218, n11219, n11220,
    n11221, n11222, n11223, n11224, n11225, n11226,
    n11227, n11228, n11229, n11230, n11231, n11232,
    n11233, n11234, n11235, n11236, n11237, n11238,
    n11239, n11240, n11241, n11242, n11243, n11244,
    n11245, n11246, n11247, n11248, n11249, n11250,
    n11251, n11252, n11253, n11254, n11255, n11256,
    n11257, n11258, n11259, n11260, n11261, n11262,
    n11263, n11264, n11265, n11266, n11267, n11268,
    n11269, n11270, n11271, n11272, n11273, n11274,
    n11275, n11276, n11277, n11278, n11279, n11280,
    n11281, n11282, n11283, n11284, n11285, n11286,
    n11287, n11288, n11289, n11290, n11291, n11292,
    n11293, n11294, n11295, n11296, n11297, n11298,
    n11299, n11300, n11301, n11302, n11303, n11304,
    n11305, n11306, n11307, n11308, n11309, n11310,
    n11311, n11312, n11313, n11314, n11315, n11316,
    n11317, n11318, n11319, n11320, n11321, n11322,
    n11323, n11324, n11325, n11326, n11327, n11328,
    n11329, n11330, n11331, n11332, n11333, n11334,
    n11335, n11336, n11337, n11338, n11339, n11340,
    n11341, n11342, n11343, n11344, n11345, n11346,
    n11347, n11348, n11349, n11350, n11351, n11352,
    n11353, n11354, n11355, n11356, n11357, n11358,
    n11359, n11360, n11361, n11362, n11363, n11364,
    n11365, n11366, n11367, n11368, n11369, n11370,
    n11371, n11372, n11373, n11374, n11375, n11376,
    n11377, n11378, n11379, n11380, n11381, n11382,
    n11383, n11384, n11385, n11386, n11387, n11388,
    n11389, n11390, n11391, n11392, n11393, n11394,
    n11395, n11396, n11398, n11399, n11400, n11401,
    n11402, n11403, n11404, n11405, n11406, n11407,
    n11408, n11409, n11410, n11411, n11412, n11413,
    n11414, n11415, n11416, n11417, n11418, n11419,
    n11420, n11421, n11422, n11423, n11424, n11425,
    n11426, n11427, n11428, n11429, n11430, n11431,
    n11432, n11433, n11434, n11435, n11436, n11437,
    n11438, n11439, n11440, n11441, n11442, n11443,
    n11444, n11445, n11446, n11447, n11448, n11449,
    n11450, n11451, n11452, n11453, n11454, n11455,
    n11456, n11457, n11458, n11459, n11460, n11461,
    n11462, n11463, n11464, n11465, n11466, n11467,
    n11468, n11469, n11470, n11471, n11472, n11473,
    n11474, n11475, n11476, n11477, n11478, n11479,
    n11480, n11481, n11482, n11483, n11484, n11485,
    n11486, n11487, n11488, n11489, n11490, n11491,
    n11492, n11493, n11494, n11495, n11496, n11497,
    n11498, n11499, n11500, n11501, n11502, n11503,
    n11504, n11505, n11506, n11507, n11508, n11509,
    n11510, n11511, n11512, n11513, n11514, n11515,
    n11516, n11517, n11518, n11519, n11520, n11521,
    n11522, n11523, n11524, n11525, n11526, n11527,
    n11528, n11529, n11530, n11531, n11532, n11533,
    n11534, n11535, n11536, n11537, n11538, n11539,
    n11540, n11541, n11542, n11543, n11544, n11545,
    n11546, n11547, n11548, n11549, n11550, n11551,
    n11552, n11553, n11554, n11555, n11556, n11557,
    n11558, n11559, n11560, n11561, n11562, n11563,
    n11564, n11565, n11566, n11567, n11568, n11569,
    n11570, n11571, n11572, n11573, n11574, n11575,
    n11576, n11577, n11578, n11579, n11580, n11581,
    n11582, n11583, n11584, n11585, n11586, n11587,
    n11588, n11589, n11590, n11591, n11592, n11593,
    n11594, n11595, n11596, n11597, n11598, n11599,
    n11600, n11601, n11602, n11603, n11604, n11605,
    n11606, n11607, n11608, n11609, n11610, n11611,
    n11612, n11613, n11614, n11615, n11616, n11617,
    n11618, n11619, n11620, n11621, n11622, n11623,
    n11624, n11625, n11626, n11627, n11628, n11629,
    n11630, n11631, n11632, n11633, n11634, n11635,
    n11636, n11637, n11638, n11639, n11640, n11641,
    n11642, n11643, n11644, n11645, n11646, n11647,
    n11648, n11649, n11650, n11651, n11652, n11653,
    n11654, n11655, n11656, n11657, n11658, n11659,
    n11660, n11661, n11662, n11663, n11664, n11665,
    n11666, n11667, n11668, n11669, n11670, n11671,
    n11672, n11673, n11674, n11675, n11676, n11677,
    n11678, n11679, n11680, n11681, n11682, n11683,
    n11684, n11685, n11686, n11687, n11688, n11689,
    n11690, n11691, n11692, n11693, n11694, n11695,
    n11696, n11697, n11698, n11699, n11700, n11701,
    n11702, n11703, n11704, n11705, n11706, n11707,
    n11708, n11709, n11710, n11711, n11712, n11713,
    n11714, n11715, n11716, n11717, n11718, n11719,
    n11720, n11721, n11722, n11723, n11724, n11725,
    n11726, n11727, n11728, n11729, n11730, n11731,
    n11732, n11733, n11734, n11735, n11736, n11737,
    n11738, n11739, n11740, n11741, n11742, n11743,
    n11744, n11745, n11746, n11747, n11748, n11749,
    n11750, n11751, n11752, n11753, n11754, n11755,
    n11756, n11757, n11758, n11759, n11760, n11761,
    n11762, n11763, n11764, n11765, n11766, n11767,
    n11768, n11769, n11770, n11771, n11772, n11773,
    n11774, n11775, n11776, n11777, n11778, n11779,
    n11780, n11781, n11782, n11783, n11784, n11785,
    n11786, n11787, n11788, n11789, n11790, n11791,
    n11792, n11793, n11794, n11795, n11796, n11797,
    n11798, n11799, n11800, n11801, n11802, n11803,
    n11804, n11805, n11806, n11807, n11808, n11809,
    n11810, n11811, n11812, n11813, n11814, n11815,
    n11816, n11817, n11818, n11819, n11820, n11821,
    n11822, n11823, n11824, n11825, n11826, n11827,
    n11828, n11829, n11830, n11831, n11832, n11833,
    n11834, n11835, n11836, n11837, n11838, n11839,
    n11840, n11841, n11842, n11843, n11844, n11845,
    n11846, n11847, n11848, n11849, n11850, n11852,
    n11853, n11854, n11855, n11856, n11857, n11858,
    n11859, n11860, n11861, n11862, n11863, n11864,
    n11865, n11866, n11867, n11868, n11869, n11870,
    n11871, n11872, n11873, n11874, n11875, n11876,
    n11877, n11878, n11879, n11880, n11881, n11882,
    n11883, n11884, n11885, n11886, n11887, n11888,
    n11889, n11890, n11891, n11892, n11893, n11894,
    n11895, n11896, n11897, n11898, n11899, n11900,
    n11901, n11902, n11903, n11904, n11905, n11906,
    n11907, n11908, n11909, n11910, n11911, n11912,
    n11913, n11914, n11915, n11916, n11917, n11918,
    n11919, n11920, n11921, n11922, n11923, n11924,
    n11925, n11926, n11927, n11928, n11929, n11930,
    n11931, n11932, n11933, n11934, n11935, n11936,
    n11937, n11938, n11939, n11940, n11941, n11942,
    n11943, n11944, n11945, n11946, n11947, n11948,
    n11949, n11950, n11951, n11952, n11953, n11954,
    n11955, n11956, n11957, n11958, n11959, n11960,
    n11961, n11962, n11963, n11964, n11965, n11966,
    n11967, n11968, n11969, n11970, n11971, n11972,
    n11973, n11974, n11975, n11976, n11977, n11978,
    n11979, n11980, n11981, n11982, n11983, n11984,
    n11985, n11986, n11987, n11988, n11989, n11990,
    n11991, n11992, n11993, n11994, n11995, n11996,
    n11997, n11998, n11999, n12000, n12001, n12002,
    n12003, n12004, n12005, n12006, n12007, n12008,
    n12009, n12010, n12011, n12012, n12013, n12014,
    n12015, n12016, n12017, n12018, n12019, n12020,
    n12021, n12022, n12023, n12024, n12025, n12026,
    n12027, n12028, n12029, n12030, n12031, n12032,
    n12033, n12034, n12035, n12036, n12037, n12038,
    n12039, n12040, n12041, n12042, n12043, n12044,
    n12045, n12046, n12047, n12048, n12049, n12050,
    n12051, n12052, n12053, n12054, n12055, n12056,
    n12057, n12058, n12059, n12060, n12061, n12062,
    n12063, n12064, n12065, n12066, n12067, n12068,
    n12069, n12070, n12071, n12072, n12073, n12074,
    n12075, n12076, n12077, n12078, n12079, n12080,
    n12081, n12082, n12083, n12084, n12085, n12086,
    n12087, n12088, n12089, n12090, n12091, n12092,
    n12093, n12094, n12095, n12096, n12097, n12098,
    n12099, n12100, n12101, n12102, n12103, n12104,
    n12105, n12106, n12107, n12108, n12109, n12110,
    n12111, n12112, n12113, n12114, n12115, n12116,
    n12117, n12118, n12119, n12120, n12121, n12122,
    n12123, n12124, n12125, n12126, n12127, n12128,
    n12129, n12130, n12131, n12132, n12133, n12134,
    n12135, n12136, n12137, n12138, n12139, n12140,
    n12141, n12142, n12143, n12144, n12145, n12146,
    n12147, n12148, n12149, n12150, n12151, n12152,
    n12153, n12154, n12155, n12156, n12157, n12158,
    n12159, n12160, n12161, n12162, n12163, n12164,
    n12165, n12166, n12167, n12168, n12169, n12170,
    n12171, n12172, n12173, n12174, n12175, n12176,
    n12177, n12178, n12179, n12180, n12181, n12182,
    n12183, n12184, n12185, n12186, n12187, n12188,
    n12189, n12190, n12191, n12192, n12193, n12194,
    n12195, n12196, n12197, n12198, n12199, n12200,
    n12201, n12202, n12203, n12204, n12205, n12206,
    n12207, n12208, n12209, n12210, n12211, n12212,
    n12213, n12214, n12215, n12216, n12217, n12218,
    n12219, n12220, n12221, n12222, n12223, n12224,
    n12225, n12226, n12227, n12228, n12229, n12230,
    n12231, n12232, n12233, n12234, n12235, n12236,
    n12237, n12238, n12239, n12240, n12241, n12242,
    n12243, n12244, n12245, n12246, n12247, n12248,
    n12249, n12250, n12251, n12252, n12253, n12254,
    n12255, n12256, n12257, n12258, n12259, n12260,
    n12261, n12262, n12263, n12264, n12265, n12266,
    n12267, n12268, n12269, n12270, n12271, n12272,
    n12273, n12274, n12275, n12276, n12277, n12278,
    n12279, n12280, n12281, n12282, n12283, n12284,
    n12285, n12286, n12287, n12288, n12289, n12290,
    n12291, n12292, n12293, n12294, n12295, n12296,
    n12297, n12298, n12299, n12300, n12301, n12302,
    n12303, n12304, n12305, n12306, n12307, n12308,
    n12309, n12310, n12311, n12312, n12313, n12315,
    n12316, n12317, n12318, n12319, n12320, n12321,
    n12322, n12323, n12324, n12325, n12326, n12327,
    n12328, n12329, n12330, n12331, n12332, n12333,
    n12334, n12335, n12336, n12337, n12338, n12339,
    n12340, n12341, n12342, n12343, n12344, n12345,
    n12346, n12347, n12348, n12349, n12350, n12351,
    n12352, n12353, n12354, n12355, n12356, n12357,
    n12358, n12359, n12360, n12361, n12362, n12363,
    n12364, n12365, n12366, n12367, n12368, n12369,
    n12370, n12371, n12372, n12373, n12374, n12375,
    n12376, n12377, n12378, n12379, n12380, n12381,
    n12382, n12383, n12384, n12385, n12386, n12387,
    n12388, n12389, n12390, n12391, n12392, n12393,
    n12394, n12395, n12396, n12397, n12398, n12399,
    n12400, n12401, n12402, n12403, n12404, n12405,
    n12406, n12407, n12408, n12409, n12410, n12411,
    n12412, n12413, n12414, n12415, n12416, n12417,
    n12418, n12419, n12420, n12421, n12422, n12423,
    n12424, n12425, n12426, n12427, n12428, n12429,
    n12430, n12431, n12432, n12433, n12434, n12435,
    n12436, n12437, n12438, n12439, n12440, n12441,
    n12442, n12443, n12444, n12445, n12446, n12447,
    n12448, n12449, n12450, n12451, n12452, n12453,
    n12454, n12455, n12456, n12457, n12458, n12459,
    n12460, n12461, n12462, n12463, n12464, n12465,
    n12466, n12467, n12468, n12469, n12470, n12471,
    n12472, n12473, n12474, n12475, n12476, n12477,
    n12478, n12479, n12480, n12481, n12482, n12483,
    n12484, n12485, n12486, n12487, n12488, n12489,
    n12490, n12491, n12492, n12493, n12494, n12495,
    n12496, n12497, n12498, n12499, n12500, n12501,
    n12502, n12503, n12504, n12505, n12506, n12507,
    n12508, n12509, n12510, n12511, n12512, n12513,
    n12514, n12515, n12516, n12517, n12518, n12519,
    n12520, n12521, n12522, n12523, n12524, n12525,
    n12526, n12527, n12528, n12529, n12530, n12531,
    n12532, n12533, n12534, n12535, n12536, n12537,
    n12538, n12539, n12540, n12541, n12542, n12543,
    n12544, n12545, n12546, n12547, n12548, n12549,
    n12550, n12551, n12552, n12553, n12554, n12555,
    n12556, n12557, n12558, n12559, n12560, n12561,
    n12562, n12563, n12564, n12565, n12566, n12567,
    n12568, n12569, n12570, n12571, n12572, n12573,
    n12574, n12575, n12576, n12577, n12578, n12579,
    n12580, n12581, n12582, n12583, n12584, n12585,
    n12586, n12587, n12588, n12589, n12590, n12591,
    n12592, n12593, n12594, n12595, n12596, n12597,
    n12598, n12599, n12600, n12601, n12602, n12603,
    n12604, n12605, n12606, n12607, n12608, n12609,
    n12610, n12611, n12612, n12613, n12614, n12615,
    n12616, n12617, n12618, n12619, n12620, n12621,
    n12622, n12623, n12624, n12625, n12626, n12627,
    n12628, n12629, n12630, n12631, n12632, n12633,
    n12634, n12635, n12636, n12637, n12638, n12639,
    n12640, n12641, n12642, n12643, n12644, n12645,
    n12646, n12647, n12648, n12649, n12650, n12651,
    n12652, n12653, n12654, n12655, n12656, n12657,
    n12658, n12659, n12660, n12661, n12662, n12663,
    n12664, n12665, n12666, n12667, n12668, n12669,
    n12670, n12671, n12672, n12673, n12674, n12675,
    n12676, n12677, n12678, n12679, n12680, n12681,
    n12682, n12683, n12684, n12685, n12686, n12687,
    n12688, n12689, n12690, n12691, n12692, n12693,
    n12694, n12695, n12696, n12697, n12698, n12699,
    n12700, n12701, n12702, n12703, n12704, n12705,
    n12706, n12707, n12708, n12709, n12710, n12711,
    n12712, n12713, n12714, n12715, n12716, n12717,
    n12718, n12719, n12720, n12721, n12722, n12723,
    n12724, n12725, n12726, n12727, n12728, n12729,
    n12730, n12731, n12732, n12733, n12734, n12735,
    n12736, n12737, n12738, n12739, n12740, n12741,
    n12742, n12743, n12744, n12745, n12746, n12747,
    n12748, n12749, n12750, n12751, n12752, n12753,
    n12754, n12755, n12756, n12757, n12758, n12759,
    n12760, n12761, n12762, n12763, n12764, n12765,
    n12766, n12767, n12768, n12769, n12770, n12771,
    n12772, n12773, n12774, n12775, n12776, n12777,
    n12778, n12779, n12780, n12781, n12782, n12783,
    n12784, n12785, n12787, n12788, n12789, n12790,
    n12791, n12792, n12793, n12794, n12795, n12796,
    n12797, n12798, n12799, n12800, n12801, n12802,
    n12803, n12804, n12805, n12806, n12807, n12808,
    n12809, n12810, n12811, n12812, n12813, n12814,
    n12815, n12816, n12817, n12818, n12819, n12820,
    n12821, n12822, n12823, n12824, n12825, n12826,
    n12827, n12828, n12829, n12830, n12831, n12832,
    n12833, n12834, n12835, n12836, n12837, n12838,
    n12839, n12840, n12841, n12842, n12843, n12844,
    n12845, n12846, n12847, n12848, n12849, n12850,
    n12851, n12852, n12853, n12854, n12855, n12856,
    n12857, n12858, n12859, n12860, n12861, n12862,
    n12863, n12864, n12865, n12866, n12867, n12868,
    n12869, n12870, n12871, n12872, n12873, n12874,
    n12875, n12876, n12877, n12878, n12879, n12880,
    n12881, n12882, n12883, n12884, n12885, n12886,
    n12887, n12888, n12889, n12890, n12891, n12892,
    n12893, n12894, n12895, n12896, n12897, n12898,
    n12899, n12900, n12901, n12902, n12903, n12904,
    n12905, n12906, n12907, n12908, n12909, n12910,
    n12911, n12912, n12913, n12914, n12915, n12916,
    n12917, n12918, n12919, n12920, n12921, n12922,
    n12923, n12924, n12925, n12926, n12927, n12928,
    n12929, n12930, n12931, n12932, n12933, n12934,
    n12935, n12936, n12937, n12938, n12939, n12940,
    n12941, n12942, n12943, n12944, n12945, n12946,
    n12947, n12948, n12949, n12950, n12951, n12952,
    n12953, n12954, n12955, n12956, n12957, n12958,
    n12959, n12960, n12961, n12962, n12963, n12964,
    n12965, n12966, n12967, n12968, n12969, n12970,
    n12971, n12972, n12973, n12974, n12975, n12976,
    n12977, n12978, n12979, n12980, n12981, n12982,
    n12983, n12984, n12985, n12986, n12987, n12988,
    n12989, n12990, n12991, n12992, n12993, n12994,
    n12995, n12996, n12997, n12998, n12999, n13000,
    n13001, n13002, n13003, n13004, n13005, n13006,
    n13007, n13008, n13009, n13010, n13011, n13012,
    n13013, n13014, n13015, n13016, n13017, n13018,
    n13019, n13020, n13021, n13022, n13023, n13024,
    n13025, n13026, n13027, n13028, n13029, n13030,
    n13031, n13032, n13033, n13034, n13035, n13036,
    n13037, n13038, n13039, n13040, n13041, n13042,
    n13043, n13044, n13045, n13046, n13047, n13048,
    n13049, n13050, n13051, n13052, n13053, n13054,
    n13055, n13056, n13057, n13058, n13059, n13060,
    n13061, n13062, n13063, n13064, n13065, n13066,
    n13067, n13068, n13069, n13070, n13071, n13072,
    n13073, n13074, n13075, n13076, n13077, n13078,
    n13079, n13080, n13081, n13082, n13083, n13084,
    n13085, n13086, n13087, n13088, n13089, n13090,
    n13091, n13092, n13093, n13094, n13095, n13096,
    n13097, n13098, n13099, n13100, n13101, n13102,
    n13103, n13104, n13105, n13106, n13107, n13108,
    n13109, n13110, n13111, n13112, n13113, n13114,
    n13115, n13116, n13117, n13118, n13119, n13120,
    n13121, n13122, n13123, n13124, n13125, n13126,
    n13127, n13128, n13129, n13130, n13131, n13132,
    n13133, n13134, n13135, n13136, n13137, n13138,
    n13139, n13140, n13141, n13142, n13143, n13144,
    n13145, n13146, n13147, n13148, n13149, n13150,
    n13151, n13152, n13153, n13154, n13155, n13156,
    n13157, n13158, n13159, n13160, n13161, n13162,
    n13163, n13164, n13165, n13166, n13167, n13168,
    n13169, n13170, n13171, n13172, n13173, n13174,
    n13175, n13176, n13177, n13178, n13179, n13180,
    n13181, n13182, n13183, n13184, n13185, n13186,
    n13187, n13188, n13189, n13190, n13191, n13192,
    n13193, n13194, n13195, n13196, n13197, n13198,
    n13199, n13200, n13201, n13202, n13203, n13204,
    n13205, n13206, n13207, n13208, n13209, n13210,
    n13211, n13212, n13213, n13214, n13215, n13216,
    n13217, n13218, n13219, n13220, n13221, n13222,
    n13223, n13224, n13225, n13226, n13227, n13228,
    n13229, n13230, n13231, n13232, n13233, n13234,
    n13235, n13236, n13237, n13238, n13239, n13240,
    n13241, n13242, n13243, n13244, n13245, n13246,
    n13247, n13248, n13249, n13250, n13251, n13252,
    n13253, n13254, n13255, n13256, n13257, n13258,
    n13259, n13260, n13261, n13262, n13263, n13264,
    n13265, n13266, n13268, n13269, n13270, n13271,
    n13272, n13273, n13274, n13275, n13276, n13277,
    n13278, n13279, n13280, n13281, n13282, n13283,
    n13284, n13285, n13286, n13287, n13288, n13289,
    n13290, n13291, n13292, n13293, n13294, n13295,
    n13296, n13297, n13298, n13299, n13300, n13301,
    n13302, n13303, n13304, n13305, n13306, n13307,
    n13308, n13309, n13310, n13311, n13312, n13313,
    n13314, n13315, n13316, n13317, n13318, n13319,
    n13320, n13321, n13322, n13323, n13324, n13325,
    n13326, n13327, n13328, n13329, n13330, n13331,
    n13332, n13333, n13334, n13335, n13336, n13337,
    n13338, n13339, n13340, n13341, n13342, n13343,
    n13344, n13345, n13346, n13347, n13348, n13349,
    n13350, n13351, n13352, n13353, n13354, n13355,
    n13356, n13357, n13358, n13359, n13360, n13361,
    n13362, n13363, n13364, n13365, n13366, n13367,
    n13368, n13369, n13370, n13371, n13372, n13373,
    n13374, n13375, n13376, n13377, n13378, n13379,
    n13380, n13381, n13382, n13383, n13384, n13385,
    n13386, n13387, n13388, n13389, n13390, n13391,
    n13392, n13393, n13394, n13395, n13396, n13397,
    n13398, n13399, n13400, n13401, n13402, n13403,
    n13404, n13405, n13406, n13407, n13408, n13409,
    n13410, n13411, n13412, n13413, n13414, n13415,
    n13416, n13417, n13418, n13419, n13420, n13421,
    n13422, n13423, n13424, n13425, n13426, n13427,
    n13428, n13429, n13430, n13431, n13432, n13433,
    n13434, n13435, n13436, n13437, n13438, n13439,
    n13440, n13441, n13442, n13443, n13444, n13445,
    n13446, n13447, n13448, n13449, n13450, n13451,
    n13452, n13453, n13454, n13455, n13456, n13457,
    n13458, n13459, n13460, n13461, n13462, n13463,
    n13464, n13465, n13466, n13467, n13468, n13469,
    n13470, n13471, n13472, n13473, n13474, n13475,
    n13476, n13477, n13478, n13479, n13480, n13481,
    n13482, n13483, n13484, n13485, n13486, n13487,
    n13488, n13489, n13490, n13491, n13492, n13493,
    n13494, n13495, n13496, n13497, n13498, n13499,
    n13500, n13501, n13502, n13503, n13504, n13505,
    n13506, n13507, n13508, n13509, n13510, n13511,
    n13512, n13513, n13514, n13515, n13516, n13517,
    n13518, n13519, n13520, n13521, n13522, n13523,
    n13524, n13525, n13526, n13527, n13528, n13529,
    n13530, n13531, n13532, n13533, n13534, n13535,
    n13536, n13537, n13538, n13539, n13540, n13541,
    n13542, n13543, n13544, n13545, n13546, n13547,
    n13548, n13549, n13550, n13551, n13552, n13553,
    n13554, n13555, n13556, n13557, n13558, n13559,
    n13560, n13561, n13562, n13563, n13564, n13565,
    n13566, n13567, n13568, n13569, n13570, n13571,
    n13572, n13573, n13574, n13575, n13576, n13577,
    n13578, n13579, n13580, n13581, n13582, n13583,
    n13584, n13585, n13586, n13587, n13588, n13589,
    n13590, n13591, n13592, n13593, n13594, n13595,
    n13596, n13597, n13598, n13599, n13600, n13601,
    n13602, n13603, n13604, n13605, n13606, n13607,
    n13608, n13609, n13610, n13611, n13612, n13613,
    n13614, n13615, n13616, n13617, n13618, n13619,
    n13620, n13621, n13622, n13623, n13624, n13625,
    n13626, n13627, n13628, n13629, n13630, n13631,
    n13632, n13633, n13634, n13635, n13636, n13637,
    n13638, n13639, n13640, n13641, n13642, n13643,
    n13644, n13645, n13646, n13647, n13648, n13649,
    n13650, n13651, n13652, n13653, n13654, n13655,
    n13656, n13657, n13658, n13659, n13660, n13661,
    n13662, n13663, n13664, n13665, n13666, n13667,
    n13668, n13669, n13670, n13671, n13672, n13673,
    n13674, n13675, n13676, n13677, n13678, n13679,
    n13680, n13681, n13682, n13683, n13684, n13685,
    n13686, n13687, n13688, n13689, n13690, n13691,
    n13692, n13693, n13694, n13695, n13696, n13697,
    n13698, n13699, n13700, n13701, n13702, n13703,
    n13704, n13705, n13706, n13707, n13708, n13709,
    n13710, n13711, n13712, n13713, n13714, n13715,
    n13716, n13717, n13718, n13719, n13720, n13721,
    n13722, n13723, n13724, n13725, n13726, n13727,
    n13728, n13729, n13730, n13731, n13732, n13733,
    n13734, n13735, n13736, n13737, n13738, n13739,
    n13740, n13741, n13742, n13743, n13744, n13745,
    n13746, n13747, n13748, n13749, n13750, n13751,
    n13752, n13753, n13754, n13755, n13756, n13758,
    n13759, n13760, n13761, n13762, n13763, n13764,
    n13765, n13766, n13767, n13768, n13769, n13770,
    n13771, n13772, n13773, n13774, n13775, n13776,
    n13777, n13778, n13779, n13780, n13781, n13782,
    n13783, n13784, n13785, n13786, n13787, n13788,
    n13789, n13790, n13791, n13792, n13793, n13794,
    n13795, n13796, n13797, n13798, n13799, n13800,
    n13801, n13802, n13803, n13804, n13805, n13806,
    n13807, n13808, n13809, n13810, n13811, n13812,
    n13813, n13814, n13815, n13816, n13817, n13818,
    n13819, n13820, n13821, n13822, n13823, n13824,
    n13825, n13826, n13827, n13828, n13829, n13830,
    n13831, n13832, n13833, n13834, n13835, n13836,
    n13837, n13838, n13839, n13840, n13841, n13842,
    n13843, n13844, n13845, n13846, n13847, n13848,
    n13849, n13850, n13851, n13852, n13853, n13854,
    n13855, n13856, n13857, n13858, n13859, n13860,
    n13861, n13862, n13863, n13864, n13865, n13866,
    n13867, n13868, n13869, n13870, n13871, n13872,
    n13873, n13874, n13875, n13876, n13877, n13878,
    n13879, n13880, n13881, n13882, n13883, n13884,
    n13885, n13886, n13887, n13888, n13889, n13890,
    n13891, n13892, n13893, n13894, n13895, n13896,
    n13897, n13898, n13899, n13900, n13901, n13902,
    n13903, n13904, n13905, n13906, n13907, n13908,
    n13909, n13910, n13911, n13912, n13913, n13914,
    n13915, n13916, n13917, n13918, n13919, n13920,
    n13921, n13922, n13923, n13924, n13925, n13926,
    n13927, n13928, n13929, n13930, n13931, n13932,
    n13933, n13934, n13935, n13936, n13937, n13938,
    n13939, n13940, n13941, n13942, n13943, n13944,
    n13945, n13946, n13947, n13948, n13949, n13950,
    n13951, n13952, n13953, n13954, n13955, n13956,
    n13957, n13958, n13959, n13960, n13961, n13962,
    n13963, n13964, n13965, n13966, n13967, n13968,
    n13969, n13970, n13971, n13972, n13973, n13974,
    n13975, n13976, n13977, n13978, n13979, n13980,
    n13981, n13982, n13983, n13984, n13985, n13986,
    n13987, n13988, n13989, n13990, n13991, n13992,
    n13993, n13994, n13995, n13996, n13997, n13998,
    n13999, n14000, n14001, n14002, n14003, n14004,
    n14005, n14006, n14007, n14008, n14009, n14010,
    n14011, n14012, n14013, n14014, n14015, n14016,
    n14017, n14018, n14019, n14020, n14021, n14022,
    n14023, n14024, n14025, n14026, n14027, n14028,
    n14029, n14030, n14031, n14032, n14033, n14034,
    n14035, n14036, n14037, n14038, n14039, n14040,
    n14041, n14042, n14043, n14044, n14045, n14046,
    n14047, n14048, n14049, n14050, n14051, n14052,
    n14053, n14054, n14055, n14056, n14057, n14058,
    n14059, n14060, n14061, n14062, n14063, n14064,
    n14065, n14066, n14067, n14068, n14069, n14070,
    n14071, n14072, n14073, n14074, n14075, n14076,
    n14077, n14078, n14079, n14080, n14081, n14082,
    n14083, n14084, n14085, n14086, n14087, n14088,
    n14089, n14090, n14091, n14092, n14093, n14094,
    n14095, n14096, n14097, n14098, n14099, n14100,
    n14101, n14102, n14103, n14104, n14105, n14106,
    n14107, n14108, n14109, n14110, n14111, n14112,
    n14113, n14114, n14115, n14116, n14117, n14118,
    n14119, n14120, n14121, n14122, n14123, n14124,
    n14125, n14126, n14127, n14128, n14129, n14130,
    n14131, n14132, n14133, n14134, n14135, n14136,
    n14137, n14138, n14139, n14140, n14141, n14142,
    n14143, n14144, n14145, n14146, n14147, n14148,
    n14149, n14150, n14151, n14152, n14153, n14154,
    n14155, n14156, n14157, n14158, n14159, n14160,
    n14161, n14162, n14163, n14164, n14165, n14166,
    n14167, n14168, n14169, n14170, n14171, n14172,
    n14173, n14174, n14175, n14176, n14177, n14178,
    n14179, n14180, n14181, n14182, n14183, n14184,
    n14185, n14186, n14187, n14188, n14189, n14190,
    n14191, n14192, n14193, n14194, n14195, n14196,
    n14197, n14198, n14199, n14200, n14201, n14202,
    n14203, n14204, n14205, n14206, n14207, n14208,
    n14209, n14210, n14211, n14212, n14213, n14214,
    n14215, n14216, n14217, n14218, n14219, n14220,
    n14221, n14222, n14223, n14224, n14225, n14226,
    n14227, n14228, n14229, n14230, n14231, n14232,
    n14233, n14234, n14235, n14236, n14237, n14238,
    n14239, n14240, n14241, n14242, n14243, n14244,
    n14245, n14246, n14247, n14248, n14249, n14250,
    n14251, n14252, n14253, n14254, n14255, n14257,
    n14258, n14259, n14260, n14261, n14262, n14263,
    n14264, n14265, n14266, n14267, n14268, n14269,
    n14270, n14271, n14272, n14273, n14274, n14275,
    n14276, n14277, n14278, n14279, n14280, n14281,
    n14282, n14283, n14284, n14285, n14286, n14287,
    n14288, n14289, n14290, n14291, n14292, n14293,
    n14294, n14295, n14296, n14297, n14298, n14299,
    n14300, n14301, n14302, n14303, n14304, n14305,
    n14306, n14307, n14308, n14309, n14310, n14311,
    n14312, n14313, n14314, n14315, n14316, n14317,
    n14318, n14319, n14320, n14321, n14322, n14323,
    n14324, n14325, n14326, n14327, n14328, n14329,
    n14330, n14331, n14332, n14333, n14334, n14335,
    n14336, n14337, n14338, n14339, n14340, n14341,
    n14342, n14343, n14344, n14345, n14346, n14347,
    n14348, n14349, n14350, n14351, n14352, n14353,
    n14354, n14355, n14356, n14357, n14358, n14359,
    n14360, n14361, n14362, n14363, n14364, n14365,
    n14366, n14367, n14368, n14369, n14370, n14371,
    n14372, n14373, n14374, n14375, n14376, n14377,
    n14378, n14379, n14380, n14381, n14382, n14383,
    n14384, n14385, n14386, n14387, n14388, n14389,
    n14390, n14391, n14392, n14393, n14394, n14395,
    n14396, n14397, n14398, n14399, n14400, n14401,
    n14402, n14403, n14404, n14405, n14406, n14407,
    n14408, n14409, n14410, n14411, n14412, n14413,
    n14414, n14415, n14416, n14417, n14418, n14419,
    n14420, n14421, n14422, n14423, n14424, n14425,
    n14426, n14427, n14428, n14429, n14430, n14431,
    n14432, n14433, n14434, n14435, n14436, n14437,
    n14438, n14439, n14440, n14441, n14442, n14443,
    n14444, n14445, n14446, n14447, n14448, n14449,
    n14450, n14451, n14452, n14453, n14454, n14455,
    n14456, n14457, n14458, n14459, n14460, n14461,
    n14462, n14463, n14464, n14465, n14466, n14467,
    n14468, n14469, n14470, n14471, n14472, n14473,
    n14474, n14475, n14476, n14477, n14478, n14479,
    n14480, n14481, n14482, n14483, n14484, n14485,
    n14486, n14487, n14488, n14489, n14490, n14491,
    n14492, n14493, n14494, n14495, n14496, n14497,
    n14498, n14499, n14500, n14501, n14502, n14503,
    n14504, n14505, n14506, n14507, n14508, n14509,
    n14510, n14511, n14512, n14513, n14514, n14515,
    n14516, n14517, n14518, n14519, n14520, n14521,
    n14522, n14523, n14524, n14525, n14526, n14527,
    n14528, n14529, n14530, n14531, n14532, n14533,
    n14534, n14535, n14536, n14537, n14538, n14539,
    n14540, n14541, n14542, n14543, n14544, n14545,
    n14546, n14547, n14548, n14549, n14550, n14551,
    n14552, n14553, n14554, n14555, n14556, n14557,
    n14558, n14559, n14560, n14561, n14562, n14563,
    n14564, n14565, n14566, n14567, n14568, n14569,
    n14570, n14571, n14572, n14573, n14574, n14575,
    n14576, n14577, n14578, n14579, n14580, n14581,
    n14582, n14583, n14584, n14585, n14586, n14587,
    n14588, n14589, n14590, n14591, n14592, n14593,
    n14594, n14595, n14596, n14597, n14598, n14599,
    n14600, n14601, n14602, n14603, n14604, n14605,
    n14606, n14607, n14608, n14609, n14610, n14611,
    n14612, n14613, n14614, n14615, n14616, n14617,
    n14618, n14619, n14620, n14621, n14622, n14623,
    n14624, n14625, n14626, n14627, n14628, n14629,
    n14630, n14631, n14632, n14633, n14634, n14635,
    n14636, n14637, n14638, n14639, n14640, n14641,
    n14642, n14643, n14644, n14645, n14646, n14647,
    n14648, n14649, n14650, n14651, n14652, n14653,
    n14654, n14655, n14656, n14657, n14658, n14659,
    n14660, n14661, n14662, n14663, n14664, n14665,
    n14666, n14667, n14668, n14669, n14670, n14671,
    n14672, n14673, n14674, n14675, n14676, n14677,
    n14678, n14679, n14680, n14681, n14682, n14683,
    n14684, n14685, n14686, n14687, n14688, n14689,
    n14690, n14691, n14692, n14693, n14694, n14695,
    n14696, n14697, n14698, n14699, n14700, n14701,
    n14702, n14703, n14704, n14705, n14706, n14707,
    n14708, n14709, n14710, n14711, n14712, n14713,
    n14714, n14715, n14716, n14717, n14718, n14719,
    n14720, n14721, n14722, n14723, n14724, n14725,
    n14726, n14727, n14728, n14729, n14730, n14731,
    n14732, n14733, n14734, n14735, n14736, n14737,
    n14738, n14739, n14740, n14741, n14742, n14743,
    n14744, n14745, n14746, n14747, n14748, n14749,
    n14750, n14751, n14752, n14753, n14754, n14755,
    n14756, n14757, n14758, n14759, n14760, n14761,
    n14762, n14763, n14765, n14766, n14767, n14768,
    n14769, n14770, n14771, n14772, n14773, n14774,
    n14775, n14776, n14777, n14778, n14779, n14780,
    n14781, n14782, n14783, n14784, n14785, n14786,
    n14787, n14788, n14789, n14790, n14791, n14792,
    n14793, n14794, n14795, n14796, n14797, n14798,
    n14799, n14800, n14801, n14802, n14803, n14804,
    n14805, n14806, n14807, n14808, n14809, n14810,
    n14811, n14812, n14813, n14814, n14815, n14816,
    n14817, n14818, n14819, n14820, n14821, n14822,
    n14823, n14824, n14825, n14826, n14827, n14828,
    n14829, n14830, n14831, n14832, n14833, n14834,
    n14835, n14836, n14837, n14838, n14839, n14840,
    n14841, n14842, n14843, n14844, n14845, n14846,
    n14847, n14848, n14849, n14850, n14851, n14852,
    n14853, n14854, n14855, n14856, n14857, n14858,
    n14859, n14860, n14861, n14862, n14863, n14864,
    n14865, n14866, n14867, n14868, n14869, n14870,
    n14871, n14872, n14873, n14874, n14875, n14876,
    n14877, n14878, n14879, n14880, n14881, n14882,
    n14883, n14884, n14885, n14886, n14887, n14888,
    n14889, n14890, n14891, n14892, n14893, n14894,
    n14895, n14896, n14897, n14898, n14899, n14900,
    n14901, n14902, n14903, n14904, n14905, n14906,
    n14907, n14908, n14909, n14910, n14911, n14912,
    n14913, n14914, n14915, n14916, n14917, n14918,
    n14919, n14920, n14921, n14922, n14923, n14924,
    n14925, n14926, n14927, n14928, n14929, n14930,
    n14931, n14932, n14933, n14934, n14935, n14936,
    n14937, n14938, n14939, n14940, n14941, n14942,
    n14943, n14944, n14945, n14946, n14947, n14948,
    n14949, n14950, n14951, n14952, n14953, n14954,
    n14955, n14956, n14957, n14958, n14959, n14960,
    n14961, n14962, n14963, n14964, n14965, n14966,
    n14967, n14968, n14969, n14970, n14971, n14972,
    n14973, n14974, n14975, n14976, n14977, n14978,
    n14979, n14980, n14981, n14982, n14983, n14984,
    n14985, n14986, n14987, n14988, n14989, n14990,
    n14991, n14992, n14993, n14994, n14995, n14996,
    n14997, n14998, n14999, n15000, n15001, n15002,
    n15003, n15004, n15005, n15006, n15007, n15008,
    n15009, n15010, n15011, n15012, n15013, n15014,
    n15015, n15016, n15017, n15018, n15019, n15020,
    n15021, n15022, n15023, n15024, n15025, n15026,
    n15027, n15028, n15029, n15030, n15031, n15032,
    n15033, n15034, n15035, n15036, n15037, n15038,
    n15039, n15040, n15041, n15042, n15043, n15044,
    n15045, n15046, n15047, n15048, n15049, n15050,
    n15051, n15052, n15053, n15054, n15055, n15056,
    n15057, n15058, n15059, n15060, n15061, n15062,
    n15063, n15064, n15065, n15066, n15067, n15068,
    n15069, n15070, n15071, n15072, n15073, n15074,
    n15075, n15076, n15077, n15078, n15079, n15080,
    n15081, n15082, n15083, n15084, n15085, n15086,
    n15087, n15088, n15089, n15090, n15091, n15092,
    n15093, n15094, n15095, n15096, n15097, n15098,
    n15099, n15100, n15101, n15102, n15103, n15104,
    n15105, n15106, n15107, n15108, n15109, n15110,
    n15111, n15112, n15113, n15114, n15115, n15116,
    n15117, n15118, n15119, n15120, n15121, n15122,
    n15123, n15124, n15125, n15126, n15127, n15128,
    n15129, n15130, n15131, n15132, n15133, n15134,
    n15135, n15136, n15137, n15138, n15139, n15140,
    n15141, n15142, n15143, n15144, n15145, n15146,
    n15147, n15148, n15149, n15150, n15151, n15152,
    n15153, n15154, n15155, n15156, n15157, n15158,
    n15159, n15160, n15161, n15162, n15163, n15164,
    n15165, n15166, n15167, n15168, n15169, n15170,
    n15171, n15172, n15173, n15174, n15175, n15176,
    n15177, n15178, n15179, n15180, n15181, n15182,
    n15183, n15184, n15185, n15186, n15187, n15188,
    n15189, n15190, n15191, n15192, n15193, n15194,
    n15195, n15196, n15197, n15198, n15199, n15200,
    n15201, n15202, n15203, n15204, n15205, n15206,
    n15207, n15208, n15209, n15210, n15211, n15212,
    n15213, n15214, n15215, n15216, n15217, n15218,
    n15219, n15220, n15221, n15222, n15223, n15224,
    n15225, n15226, n15227, n15228, n15229, n15230,
    n15231, n15232, n15233, n15234, n15235, n15236,
    n15237, n15238, n15239, n15240, n15241, n15242,
    n15243, n15244, n15245, n15246, n15247, n15248,
    n15249, n15250, n15251, n15252, n15253, n15254,
    n15255, n15256, n15257, n15258, n15259, n15260,
    n15261, n15262, n15263, n15264, n15265, n15266,
    n15267, n15268, n15269, n15270, n15271, n15272,
    n15273, n15274, n15275, n15276, n15277, n15278,
    n15279, n15280, n15282, n15283, n15284, n15285,
    n15286, n15287, n15288, n15289, n15290, n15291,
    n15292, n15293, n15294, n15295, n15296, n15297,
    n15298, n15299, n15300, n15301, n15302, n15303,
    n15304, n15305, n15306, n15307, n15308, n15309,
    n15310, n15311, n15312, n15313, n15314, n15315,
    n15316, n15317, n15318, n15319, n15320, n15321,
    n15322, n15323, n15324, n15325, n15326, n15327,
    n15328, n15329, n15330, n15331, n15332, n15333,
    n15334, n15335, n15336, n15337, n15338, n15339,
    n15340, n15341, n15342, n15343, n15344, n15345,
    n15346, n15347, n15348, n15349, n15350, n15351,
    n15352, n15353, n15354, n15355, n15356, n15357,
    n15358, n15359, n15360, n15361, n15362, n15363,
    n15364, n15365, n15366, n15367, n15368, n15369,
    n15370, n15371, n15372, n15373, n15374, n15375,
    n15376, n15377, n15378, n15379, n15380, n15381,
    n15382, n15383, n15384, n15385, n15386, n15387,
    n15388, n15389, n15390, n15391, n15392, n15393,
    n15394, n15395, n15396, n15397, n15398, n15399,
    n15400, n15401, n15402, n15403, n15404, n15405,
    n15406, n15407, n15408, n15409, n15410, n15411,
    n15412, n15413, n15414, n15415, n15416, n15417,
    n15418, n15419, n15420, n15421, n15422, n15423,
    n15424, n15425, n15426, n15427, n15428, n15429,
    n15430, n15431, n15432, n15433, n15434, n15435,
    n15436, n15437, n15438, n15439, n15440, n15441,
    n15442, n15443, n15444, n15445, n15446, n15447,
    n15448, n15449, n15450, n15451, n15452, n15453,
    n15454, n15455, n15456, n15457, n15458, n15459,
    n15460, n15461, n15462, n15463, n15464, n15465,
    n15466, n15467, n15468, n15469, n15470, n15471,
    n15472, n15473, n15474, n15475, n15476, n15477,
    n15478, n15479, n15480, n15481, n15482, n15483,
    n15484, n15485, n15486, n15487, n15488, n15489,
    n15490, n15491, n15492, n15493, n15494, n15495,
    n15496, n15497, n15498, n15499, n15500, n15501,
    n15502, n15503, n15504, n15505, n15506, n15507,
    n15508, n15509, n15510, n15511, n15512, n15513,
    n15514, n15515, n15516, n15517, n15518, n15519,
    n15520, n15521, n15522, n15523, n15524, n15525,
    n15526, n15527, n15528, n15529, n15530, n15531,
    n15532, n15533, n15534, n15535, n15536, n15537,
    n15538, n15539, n15540, n15541, n15542, n15543,
    n15544, n15545, n15546, n15547, n15548, n15549,
    n15550, n15551, n15552, n15553, n15554, n15555,
    n15556, n15557, n15558, n15559, n15560, n15561,
    n15562, n15563, n15564, n15565, n15566, n15567,
    n15568, n15569, n15570, n15571, n15572, n15573,
    n15574, n15575, n15576, n15577, n15578, n15579,
    n15580, n15581, n15582, n15583, n15584, n15585,
    n15586, n15587, n15588, n15589, n15590, n15591,
    n15592, n15593, n15594, n15595, n15596, n15597,
    n15598, n15599, n15600, n15601, n15602, n15603,
    n15604, n15605, n15606, n15607, n15608, n15609,
    n15610, n15611, n15612, n15613, n15614, n15615,
    n15616, n15617, n15618, n15619, n15620, n15621,
    n15622, n15623, n15624, n15625, n15626, n15627,
    n15628, n15629, n15630, n15631, n15632, n15633,
    n15634, n15635, n15636, n15637, n15638, n15639,
    n15640, n15641, n15642, n15643, n15644, n15645,
    n15646, n15647, n15648, n15649, n15650, n15651,
    n15652, n15653, n15654, n15655, n15656, n15657,
    n15658, n15659, n15660, n15661, n15662, n15663,
    n15664, n15665, n15666, n15667, n15668, n15669,
    n15670, n15671, n15672, n15673, n15674, n15675,
    n15676, n15677, n15678, n15679, n15680, n15681,
    n15682, n15683, n15684, n15685, n15686, n15687,
    n15688, n15689, n15690, n15691, n15692, n15693,
    n15694, n15695, n15696, n15697, n15698, n15699,
    n15700, n15701, n15702, n15703, n15704, n15705,
    n15706, n15707, n15708, n15709, n15710, n15711,
    n15712, n15713, n15714, n15715, n15716, n15717,
    n15718, n15719, n15720, n15721, n15722, n15723,
    n15724, n15725, n15726, n15727, n15728, n15729,
    n15730, n15731, n15732, n15733, n15734, n15735,
    n15736, n15737, n15738, n15739, n15740, n15741,
    n15742, n15743, n15744, n15745, n15746, n15747,
    n15748, n15749, n15750, n15751, n15752, n15753,
    n15754, n15755, n15756, n15757, n15758, n15759,
    n15760, n15761, n15762, n15763, n15764, n15765,
    n15766, n15767, n15768, n15769, n15770, n15771,
    n15772, n15773, n15774, n15775, n15776, n15777,
    n15778, n15779, n15780, n15781, n15782, n15783,
    n15784, n15785, n15786, n15787, n15788, n15789,
    n15790, n15791, n15792, n15793, n15794, n15795,
    n15796, n15797, n15798, n15799, n15800, n15801,
    n15802, n15803, n15804, n15806, n15807, n15808,
    n15809, n15810, n15811, n15812, n15813, n15814,
    n15815, n15816, n15817, n15818, n15819, n15820,
    n15821, n15822, n15823, n15824, n15825, n15826,
    n15827, n15828, n15829, n15830, n15831, n15832,
    n15833, n15834, n15835, n15836, n15837, n15838,
    n15839, n15840, n15841, n15842, n15843, n15844,
    n15845, n15846, n15847, n15848, n15849, n15850,
    n15851, n15852, n15853, n15854, n15855, n15856,
    n15857, n15858, n15859, n15860, n15861, n15862,
    n15863, n15864, n15865, n15866, n15867, n15868,
    n15869, n15870, n15871, n15872, n15873, n15874,
    n15875, n15876, n15877, n15878, n15879, n15880,
    n15881, n15882, n15883, n15884, n15885, n15886,
    n15887, n15888, n15889, n15890, n15891, n15892,
    n15893, n15894, n15895, n15896, n15897, n15898,
    n15899, n15900, n15901, n15902, n15903, n15904,
    n15905, n15906, n15907, n15908, n15909, n15910,
    n15911, n15912, n15913, n15914, n15915, n15916,
    n15917, n15918, n15919, n15920, n15921, n15922,
    n15923, n15924, n15925, n15926, n15927, n15928,
    n15929, n15930, n15931, n15932, n15933, n15934,
    n15935, n15936, n15937, n15938, n15939, n15940,
    n15941, n15942, n15943, n15944, n15945, n15946,
    n15947, n15948, n15949, n15950, n15951, n15952,
    n15953, n15954, n15955, n15956, n15957, n15958,
    n15959, n15960, n15961, n15962, n15963, n15964,
    n15965, n15966, n15967, n15968, n15969, n15970,
    n15971, n15972, n15973, n15974, n15975, n15976,
    n15977, n15978, n15979, n15980, n15981, n15982,
    n15983, n15984, n15985, n15986, n15987, n15988,
    n15989, n15990, n15991, n15992, n15993, n15994,
    n15995, n15996, n15997, n15998, n15999, n16000,
    n16001, n16002, n16003, n16004, n16005, n16006,
    n16007, n16008, n16009, n16010, n16011, n16012,
    n16013, n16014, n16015, n16016, n16017, n16018,
    n16019, n16020, n16021, n16022, n16023, n16024,
    n16025, n16026, n16027, n16028, n16029, n16030,
    n16031, n16032, n16033, n16034, n16035, n16036,
    n16037, n16038, n16039, n16040, n16041, n16042,
    n16043, n16044, n16045, n16046, n16047, n16048,
    n16049, n16050, n16051, n16052, n16053, n16054,
    n16055, n16056, n16057, n16058, n16059, n16060,
    n16061, n16062, n16063, n16064, n16065, n16066,
    n16067, n16068, n16069, n16070, n16071, n16072,
    n16073, n16074, n16075, n16076, n16077, n16078,
    n16079, n16080, n16081, n16082, n16083, n16084,
    n16085, n16086, n16087, n16088, n16089, n16090,
    n16091, n16092, n16093, n16094, n16095, n16096,
    n16097, n16098, n16099, n16100, n16101, n16102,
    n16103, n16104, n16105, n16106, n16107, n16108,
    n16109, n16110, n16111, n16112, n16113, n16114,
    n16115, n16116, n16117, n16118, n16119, n16120,
    n16121, n16122, n16123, n16124, n16125, n16126,
    n16127, n16128, n16129, n16130, n16131, n16132,
    n16133, n16134, n16135, n16136, n16137, n16138,
    n16139, n16140, n16141, n16142, n16143, n16144,
    n16145, n16146, n16147, n16148, n16149, n16150,
    n16151, n16152, n16153, n16154, n16155, n16156,
    n16157, n16158, n16159, n16160, n16161, n16162,
    n16163, n16164, n16165, n16166, n16167, n16168,
    n16169, n16170, n16171, n16172, n16173, n16174,
    n16175, n16176, n16177, n16178, n16179, n16180,
    n16181, n16182, n16183, n16184, n16185, n16186,
    n16187, n16188, n16189, n16190, n16191, n16192,
    n16193, n16194, n16195, n16196, n16197, n16198,
    n16199, n16200, n16201, n16202, n16203, n16204,
    n16205, n16206, n16207, n16208, n16209, n16210,
    n16211, n16212, n16213, n16214, n16215, n16216,
    n16217, n16218, n16219, n16220, n16221, n16222,
    n16223, n16224, n16225, n16226, n16227, n16228,
    n16229, n16230, n16231, n16232, n16233, n16234,
    n16235, n16236, n16237, n16238, n16239, n16240,
    n16241, n16242, n16243, n16244, n16245, n16246,
    n16247, n16248, n16249, n16250, n16251, n16252,
    n16253, n16254, n16255, n16256, n16257, n16258,
    n16259, n16260, n16261, n16262, n16263, n16264,
    n16265, n16266, n16267, n16268, n16269, n16270,
    n16271, n16272, n16273, n16274, n16275, n16276,
    n16277, n16278, n16279, n16280, n16281, n16282,
    n16283, n16284, n16285, n16286, n16287, n16288,
    n16289, n16290, n16291, n16292, n16293, n16294,
    n16295, n16296, n16297, n16298, n16299, n16300,
    n16301, n16302, n16303, n16304, n16305, n16306,
    n16307, n16308, n16309, n16310, n16311, n16312,
    n16313, n16314, n16315, n16316, n16317, n16318,
    n16319, n16320, n16321, n16322, n16323, n16324,
    n16325, n16326, n16327, n16328, n16329, n16330,
    n16331, n16332, n16333, n16334, n16335, n16336,
    n16337, n16339, n16340, n16341, n16342, n16343,
    n16344, n16345, n16346, n16347, n16348, n16349,
    n16350, n16351, n16352, n16353, n16354, n16355,
    n16356, n16357, n16358, n16359, n16360, n16361,
    n16362, n16363, n16364, n16365, n16366, n16367,
    n16368, n16369, n16370, n16371, n16372, n16373,
    n16374, n16375, n16376, n16377, n16378, n16379,
    n16380, n16381, n16382, n16383, n16384, n16385,
    n16386, n16387, n16388, n16389, n16390, n16391,
    n16392, n16393, n16394, n16395, n16396, n16397,
    n16398, n16399, n16400, n16401, n16402, n16403,
    n16404, n16405, n16406, n16407, n16408, n16409,
    n16410, n16411, n16412, n16413, n16414, n16415,
    n16416, n16417, n16418, n16419, n16420, n16421,
    n16422, n16423, n16424, n16425, n16426, n16427,
    n16428, n16429, n16430, n16431, n16432, n16433,
    n16434, n16435, n16436, n16437, n16438, n16439,
    n16440, n16441, n16442, n16443, n16444, n16445,
    n16446, n16447, n16448, n16449, n16450, n16451,
    n16452, n16453, n16454, n16455, n16456, n16457,
    n16458, n16459, n16460, n16461, n16462, n16463,
    n16464, n16465, n16466, n16467, n16468, n16469,
    n16470, n16471, n16472, n16473, n16474, n16475,
    n16476, n16477, n16478, n16479, n16480, n16481,
    n16482, n16483, n16484, n16485, n16486, n16487,
    n16488, n16489, n16490, n16491, n16492, n16493,
    n16494, n16495, n16496, n16497, n16498, n16499,
    n16500, n16501, n16502, n16503, n16504, n16505,
    n16506, n16507, n16508, n16509, n16510, n16511,
    n16512, n16513, n16514, n16515, n16516, n16517,
    n16518, n16519, n16520, n16521, n16522, n16523,
    n16524, n16525, n16526, n16527, n16528, n16529,
    n16530, n16531, n16532, n16533, n16534, n16535,
    n16536, n16537, n16538, n16539, n16540, n16541,
    n16542, n16543, n16544, n16545, n16546, n16547,
    n16548, n16549, n16550, n16551, n16552, n16553,
    n16554, n16555, n16556, n16557, n16558, n16559,
    n16560, n16561, n16562, n16563, n16564, n16565,
    n16566, n16567, n16568, n16569, n16570, n16571,
    n16572, n16573, n16574, n16575, n16576, n16577,
    n16578, n16579, n16580, n16581, n16582, n16583,
    n16584, n16585, n16586, n16587, n16588, n16589,
    n16590, n16591, n16592, n16593, n16594, n16595,
    n16596, n16597, n16598, n16599, n16600, n16601,
    n16602, n16603, n16604, n16605, n16606, n16607,
    n16608, n16609, n16610, n16611, n16612, n16613,
    n16614, n16615, n16616, n16617, n16618, n16619,
    n16620, n16621, n16622, n16623, n16624, n16625,
    n16626, n16627, n16628, n16629, n16630, n16631,
    n16632, n16633, n16634, n16635, n16636, n16637,
    n16638, n16639, n16640, n16641, n16642, n16643,
    n16644, n16645, n16646, n16647, n16648, n16649,
    n16650, n16651, n16652, n16653, n16654, n16655,
    n16656, n16657, n16658, n16659, n16660, n16661,
    n16662, n16663, n16664, n16665, n16666, n16667,
    n16668, n16669, n16670, n16671, n16672, n16673,
    n16674, n16675, n16676, n16677, n16678, n16679,
    n16680, n16681, n16682, n16683, n16684, n16685,
    n16686, n16687, n16688, n16689, n16690, n16691,
    n16692, n16693, n16694, n16695, n16696, n16697,
    n16698, n16699, n16700, n16701, n16702, n16703,
    n16704, n16705, n16706, n16707, n16708, n16709,
    n16710, n16711, n16712, n16713, n16714, n16715,
    n16716, n16717, n16718, n16719, n16720, n16721,
    n16722, n16723, n16724, n16725, n16726, n16727,
    n16728, n16729, n16730, n16731, n16732, n16733,
    n16734, n16735, n16736, n16737, n16738, n16739,
    n16740, n16741, n16742, n16743, n16744, n16745,
    n16746, n16747, n16748, n16749, n16750, n16751,
    n16752, n16753, n16754, n16755, n16756, n16757,
    n16758, n16759, n16760, n16761, n16762, n16763,
    n16764, n16765, n16766, n16767, n16768, n16769,
    n16770, n16771, n16772, n16773, n16774, n16775,
    n16776, n16777, n16778, n16779, n16780, n16781,
    n16782, n16783, n16784, n16785, n16786, n16787,
    n16788, n16789, n16790, n16791, n16792, n16793,
    n16794, n16795, n16796, n16797, n16798, n16799,
    n16800, n16801, n16802, n16803, n16804, n16805,
    n16806, n16807, n16808, n16809, n16810, n16811,
    n16812, n16813, n16814, n16815, n16816, n16817,
    n16818, n16819, n16820, n16821, n16822, n16823,
    n16824, n16825, n16826, n16827, n16828, n16829,
    n16830, n16831, n16832, n16833, n16834, n16835,
    n16836, n16837, n16838, n16839, n16840, n16841,
    n16842, n16843, n16844, n16845, n16846, n16847,
    n16848, n16849, n16850, n16851, n16852, n16853,
    n16854, n16855, n16856, n16857, n16858, n16859,
    n16860, n16861, n16862, n16863, n16864, n16865,
    n16866, n16867, n16868, n16869, n16870, n16871,
    n16872, n16873, n16874, n16875, n16876, n16877,
    n16878, n16879, n16881, n16882, n16883, n16884,
    n16885, n16886, n16887, n16888, n16889, n16890,
    n16891, n16892, n16893, n16894, n16895, n16896,
    n16897, n16898, n16899, n16900, n16901, n16902,
    n16903, n16904, n16905, n16906, n16907, n16908,
    n16909, n16910, n16911, n16912, n16913, n16914,
    n16915, n16916, n16917, n16918, n16919, n16920,
    n16921, n16922, n16923, n16924, n16925, n16926,
    n16927, n16928, n16929, n16930, n16931, n16932,
    n16933, n16934, n16935, n16936, n16937, n16938,
    n16939, n16940, n16941, n16942, n16943, n16944,
    n16945, n16946, n16947, n16948, n16949, n16950,
    n16951, n16952, n16953, n16954, n16955, n16956,
    n16957, n16958, n16959, n16960, n16961, n16962,
    n16963, n16964, n16965, n16966, n16967, n16968,
    n16969, n16970, n16971, n16972, n16973, n16974,
    n16975, n16976, n16977, n16978, n16979, n16980,
    n16981, n16982, n16983, n16984, n16985, n16986,
    n16987, n16988, n16989, n16990, n16991, n16992,
    n16993, n16994, n16995, n16996, n16997, n16998,
    n16999, n17000, n17001, n17002, n17003, n17004,
    n17005, n17006, n17007, n17008, n17009, n17010,
    n17011, n17012, n17013, n17014, n17015, n17016,
    n17017, n17018, n17019, n17020, n17021, n17022,
    n17023, n17024, n17025, n17026, n17027, n17028,
    n17029, n17030, n17031, n17032, n17033, n17034,
    n17035, n17036, n17037, n17038, n17039, n17040,
    n17041, n17042, n17043, n17044, n17045, n17046,
    n17047, n17048, n17049, n17050, n17051, n17052,
    n17053, n17054, n17055, n17056, n17057, n17058,
    n17059, n17060, n17061, n17062, n17063, n17064,
    n17065, n17066, n17067, n17068, n17069, n17070,
    n17071, n17072, n17073, n17074, n17075, n17076,
    n17077, n17078, n17079, n17080, n17081, n17082,
    n17083, n17084, n17085, n17086, n17087, n17088,
    n17089, n17090, n17091, n17092, n17093, n17094,
    n17095, n17096, n17097, n17098, n17099, n17100,
    n17101, n17102, n17103, n17104, n17105, n17106,
    n17107, n17108, n17109, n17110, n17111, n17112,
    n17113, n17114, n17115, n17116, n17117, n17118,
    n17119, n17120, n17121, n17122, n17123, n17124,
    n17125, n17126, n17127, n17128, n17129, n17130,
    n17131, n17132, n17133, n17134, n17135, n17136,
    n17137, n17138, n17139, n17140, n17141, n17142,
    n17143, n17144, n17145, n17146, n17147, n17148,
    n17149, n17150, n17151, n17152, n17153, n17154,
    n17155, n17156, n17157, n17158, n17159, n17160,
    n17161, n17162, n17163, n17164, n17165, n17166,
    n17167, n17168, n17169, n17170, n17171, n17172,
    n17173, n17174, n17175, n17176, n17177, n17178,
    n17179, n17180, n17181, n17182, n17183, n17184,
    n17185, n17186, n17187, n17188, n17189, n17190,
    n17191, n17192, n17193, n17194, n17195, n17196,
    n17197, n17198, n17199, n17200, n17201, n17202,
    n17203, n17204, n17205, n17206, n17207, n17208,
    n17209, n17210, n17211, n17212, n17213, n17214,
    n17215, n17216, n17217, n17218, n17219, n17220,
    n17221, n17222, n17223, n17224, n17225, n17226,
    n17227, n17228, n17229, n17230, n17231, n17232,
    n17233, n17234, n17235, n17236, n17237, n17238,
    n17239, n17240, n17241, n17242, n17243, n17244,
    n17245, n17246, n17247, n17248, n17249, n17250,
    n17251, n17252, n17253, n17254, n17255, n17256,
    n17257, n17258, n17259, n17260, n17261, n17262,
    n17263, n17264, n17265, n17266, n17267, n17268,
    n17269, n17270, n17271, n17272, n17273, n17274,
    n17275, n17276, n17277, n17278, n17279, n17280,
    n17281, n17282, n17283, n17284, n17285, n17286,
    n17287, n17288, n17289, n17290, n17291, n17292,
    n17293, n17294, n17295, n17296, n17297, n17298,
    n17299, n17300, n17301, n17302, n17303, n17304,
    n17305, n17306, n17307, n17308, n17309, n17310,
    n17311, n17312, n17313, n17314, n17315, n17316,
    n17317, n17318, n17319, n17320, n17321, n17322,
    n17323, n17324, n17325, n17326, n17327, n17328,
    n17329, n17330, n17331, n17332, n17333, n17334,
    n17335, n17336, n17337, n17338, n17339, n17340,
    n17341, n17342, n17343, n17344, n17345, n17346,
    n17347, n17348, n17349, n17350, n17351, n17352,
    n17353, n17354, n17355, n17356, n17357, n17358,
    n17359, n17360, n17361, n17362, n17363, n17364,
    n17365, n17366, n17367, n17368, n17369, n17370,
    n17371, n17372, n17373, n17374, n17375, n17376,
    n17377, n17378, n17379, n17380, n17381, n17382,
    n17383, n17384, n17385, n17386, n17387, n17388,
    n17389, n17390, n17391, n17392, n17393, n17394,
    n17395, n17396, n17397, n17398, n17399, n17400,
    n17401, n17402, n17403, n17404, n17405, n17406,
    n17407, n17408, n17409, n17410, n17411, n17412,
    n17413, n17414, n17415, n17416, n17417, n17418,
    n17419, n17420, n17421, n17422, n17423, n17424,
    n17425, n17426, n17427, n17428, n17429, n17430,
    n17432, n17433, n17434, n17435, n17436, n17437,
    n17438, n17439, n17440, n17441, n17442, n17443,
    n17444, n17445, n17446, n17447, n17448, n17449,
    n17450, n17451, n17452, n17453, n17454, n17455,
    n17456, n17457, n17458, n17459, n17460, n17461,
    n17462, n17463, n17464, n17465, n17466, n17467,
    n17468, n17469, n17470, n17471, n17472, n17473,
    n17474, n17475, n17476, n17477, n17478, n17479,
    n17480, n17481, n17482, n17483, n17484, n17485,
    n17486, n17487, n17488, n17489, n17490, n17491,
    n17492, n17493, n17494, n17495, n17496, n17497,
    n17498, n17499, n17500, n17501, n17502, n17503,
    n17504, n17505, n17506, n17507, n17508, n17509,
    n17510, n17511, n17512, n17513, n17514, n17515,
    n17516, n17517, n17518, n17519, n17520, n17521,
    n17522, n17523, n17524, n17525, n17526, n17527,
    n17528, n17529, n17530, n17531, n17532, n17533,
    n17534, n17535, n17536, n17537, n17538, n17539,
    n17540, n17541, n17542, n17543, n17544, n17545,
    n17546, n17547, n17548, n17549, n17550, n17551,
    n17552, n17553, n17554, n17555, n17556, n17557,
    n17558, n17559, n17560, n17561, n17562, n17563,
    n17564, n17565, n17566, n17567, n17568, n17569,
    n17570, n17571, n17572, n17573, n17574, n17575,
    n17576, n17577, n17578, n17579, n17580, n17581,
    n17582, n17583, n17584, n17585, n17586, n17587,
    n17588, n17589, n17590, n17591, n17592, n17593,
    n17594, n17595, n17596, n17597, n17598, n17599,
    n17600, n17601, n17602, n17603, n17604, n17605,
    n17606, n17607, n17608, n17609, n17610, n17611,
    n17612, n17613, n17614, n17615, n17616, n17617,
    n17618, n17619, n17620, n17621, n17622, n17623,
    n17624, n17625, n17626, n17627, n17628, n17629,
    n17630, n17631, n17632, n17633, n17634, n17635,
    n17636, n17637, n17638, n17639, n17640, n17641,
    n17642, n17643, n17644, n17645, n17646, n17647,
    n17648, n17649, n17650, n17651, n17652, n17653,
    n17654, n17655, n17656, n17657, n17658, n17659,
    n17660, n17661, n17662, n17663, n17664, n17665,
    n17666, n17667, n17668, n17669, n17670, n17671,
    n17672, n17673, n17674, n17675, n17676, n17677,
    n17678, n17679, n17680, n17681, n17682, n17683,
    n17684, n17685, n17686, n17687, n17688, n17689,
    n17690, n17691, n17692, n17693, n17694, n17695,
    n17696, n17697, n17698, n17699, n17700, n17701,
    n17702, n17703, n17704, n17705, n17706, n17707,
    n17708, n17709, n17710, n17711, n17712, n17713,
    n17714, n17715, n17716, n17717, n17718, n17719,
    n17720, n17721, n17722, n17723, n17724, n17725,
    n17726, n17727, n17728, n17729, n17730, n17731,
    n17732, n17733, n17734, n17735, n17736, n17737,
    n17738, n17739, n17740, n17741, n17742, n17743,
    n17744, n17745, n17746, n17747, n17748, n17749,
    n17750, n17751, n17752, n17753, n17754, n17755,
    n17756, n17757, n17758, n17759, n17760, n17761,
    n17762, n17763, n17764, n17765, n17766, n17767,
    n17768, n17769, n17770, n17771, n17772, n17773,
    n17774, n17775, n17776, n17777, n17778, n17779,
    n17780, n17781, n17782, n17783, n17784, n17785,
    n17786, n17787, n17788, n17789, n17790, n17791,
    n17792, n17793, n17794, n17795, n17796, n17797,
    n17798, n17799, n17800, n17801, n17802, n17803,
    n17804, n17805, n17806, n17807, n17808, n17809,
    n17810, n17811, n17812, n17813, n17814, n17815,
    n17816, n17817, n17818, n17819, n17820, n17821,
    n17822, n17823, n17824, n17825, n17826, n17827,
    n17828, n17829, n17830, n17831, n17832, n17833,
    n17834, n17835, n17836, n17837, n17838, n17839,
    n17840, n17841, n17842, n17843, n17844, n17845,
    n17846, n17847, n17848, n17849, n17850, n17851,
    n17852, n17853, n17854, n17855, n17856, n17857,
    n17858, n17859, n17860, n17861, n17862, n17863,
    n17864, n17865, n17866, n17867, n17868, n17869,
    n17870, n17871, n17872, n17873, n17874, n17875,
    n17876, n17877, n17878, n17879, n17880, n17881,
    n17882, n17883, n17884, n17885, n17886, n17887,
    n17888, n17889, n17890, n17891, n17892, n17893,
    n17894, n17895, n17896, n17897, n17898, n17899,
    n17900, n17901, n17902, n17903, n17904, n17905,
    n17906, n17907, n17908, n17909, n17910, n17911,
    n17912, n17913, n17914, n17915, n17916, n17917,
    n17918, n17919, n17920, n17921, n17922, n17923,
    n17924, n17925, n17926, n17927, n17928, n17929,
    n17930, n17931, n17932, n17933, n17934, n17935,
    n17936, n17937, n17938, n17939, n17940, n17941,
    n17942, n17943, n17944, n17945, n17946, n17947,
    n17948, n17949, n17950, n17951, n17952, n17953,
    n17954, n17955, n17956, n17957, n17958, n17959,
    n17960, n17961, n17962, n17963, n17964, n17965,
    n17966, n17967, n17968, n17969, n17970, n17971,
    n17972, n17973, n17974, n17975, n17976, n17977,
    n17978, n17979, n17980, n17981, n17982, n17983,
    n17984, n17985, n17986, n17987, n17988, n17989,
    n17990, n17992, n17993, n17994, n17995, n17996,
    n17997, n17998, n17999, n18000, n18001, n18002,
    n18003, n18004, n18005, n18006, n18007, n18008,
    n18009, n18010, n18011, n18012, n18013, n18014,
    n18015, n18016, n18017, n18018, n18019, n18020,
    n18021, n18022, n18023, n18024, n18025, n18026,
    n18027, n18028, n18029, n18030, n18031, n18032,
    n18033, n18034, n18035, n18036, n18037, n18038,
    n18039, n18040, n18041, n18042, n18043, n18044,
    n18045, n18046, n18047, n18048, n18049, n18050,
    n18051, n18052, n18053, n18054, n18055, n18056,
    n18057, n18058, n18059, n18060, n18061, n18062,
    n18063, n18064, n18065, n18066, n18067, n18068,
    n18069, n18070, n18071, n18072, n18073, n18074,
    n18075, n18076, n18077, n18078, n18079, n18080,
    n18081, n18082, n18083, n18084, n18085, n18086,
    n18087, n18088, n18089, n18090, n18091, n18092,
    n18093, n18094, n18095, n18096, n18097, n18098,
    n18099, n18100, n18101, n18102, n18103, n18104,
    n18105, n18106, n18107, n18108, n18109, n18110,
    n18111, n18112, n18113, n18114, n18115, n18116,
    n18117, n18118, n18119, n18120, n18121, n18122,
    n18123, n18124, n18125, n18126, n18127, n18128,
    n18129, n18130, n18131, n18132, n18133, n18134,
    n18135, n18136, n18137, n18138, n18139, n18140,
    n18141, n18142, n18143, n18144, n18145, n18146,
    n18147, n18148, n18149, n18150, n18151, n18152,
    n18153, n18154, n18155, n18156, n18157, n18158,
    n18159, n18160, n18161, n18162, n18163, n18164,
    n18165, n18166, n18167, n18168, n18169, n18170,
    n18171, n18172, n18173, n18174, n18175, n18176,
    n18177, n18178, n18179, n18180, n18181, n18182,
    n18183, n18184, n18185, n18186, n18187, n18188,
    n18189, n18190, n18191, n18192, n18193, n18194,
    n18195, n18196, n18197, n18198, n18199, n18200,
    n18201, n18202, n18203, n18204, n18205, n18206,
    n18207, n18208, n18209, n18210, n18211, n18212,
    n18213, n18214, n18215, n18216, n18217, n18218,
    n18219, n18220, n18221, n18222, n18223, n18224,
    n18225, n18226, n18227, n18228, n18229, n18230,
    n18231, n18232, n18233, n18234, n18235, n18236,
    n18237, n18238, n18239, n18240, n18241, n18242,
    n18243, n18244, n18245, n18246, n18247, n18248,
    n18249, n18250, n18251, n18252, n18253, n18254,
    n18255, n18256, n18257, n18258, n18259, n18260,
    n18261, n18262, n18263, n18264, n18265, n18266,
    n18267, n18268, n18269, n18270, n18271, n18272,
    n18273, n18274, n18275, n18276, n18277, n18278,
    n18279, n18280, n18281, n18282, n18283, n18284,
    n18285, n18286, n18287, n18288, n18289, n18290,
    n18291, n18292, n18293, n18294, n18295, n18296,
    n18297, n18298, n18299, n18300, n18301, n18302,
    n18303, n18304, n18305, n18306, n18307, n18308,
    n18309, n18310, n18311, n18312, n18313, n18314,
    n18315, n18316, n18317, n18318, n18319, n18320,
    n18321, n18322, n18323, n18324, n18325, n18326,
    n18327, n18328, n18329, n18330, n18331, n18332,
    n18333, n18334, n18335, n18336, n18337, n18338,
    n18339, n18340, n18341, n18342, n18343, n18344,
    n18345, n18346, n18347, n18348, n18349, n18350,
    n18351, n18352, n18353, n18354, n18355, n18356,
    n18357, n18358, n18359, n18360, n18361, n18362,
    n18363, n18364, n18365, n18366, n18367, n18368,
    n18369, n18370, n18371, n18372, n18373, n18374,
    n18375, n18376, n18377, n18378, n18379, n18380,
    n18381, n18382, n18383, n18384, n18385, n18386,
    n18387, n18388, n18389, n18390, n18391, n18392,
    n18393, n18394, n18395, n18396, n18397, n18398,
    n18399, n18400, n18401, n18402, n18403, n18404,
    n18405, n18406, n18407, n18408, n18409, n18410,
    n18411, n18412, n18413, n18414, n18415, n18416,
    n18417, n18418, n18419, n18420, n18421, n18422,
    n18423, n18424, n18425, n18426, n18427, n18428,
    n18429, n18430, n18431, n18432, n18433, n18434,
    n18435, n18436, n18437, n18438, n18439, n18440,
    n18441, n18442, n18443, n18444, n18445, n18446,
    n18447, n18448, n18449, n18450, n18451, n18452,
    n18453, n18454, n18455, n18456, n18457, n18458,
    n18459, n18460, n18461, n18462, n18463, n18464,
    n18465, n18466, n18467, n18468, n18469, n18470,
    n18471, n18472, n18473, n18474, n18475, n18476,
    n18477, n18478, n18479, n18480, n18481, n18482,
    n18483, n18484, n18485, n18486, n18487, n18488,
    n18489, n18490, n18491, n18492, n18493, n18494,
    n18495, n18496, n18497, n18498, n18499, n18500,
    n18501, n18502, n18503, n18504, n18505, n18506,
    n18507, n18508, n18509, n18510, n18511, n18512,
    n18513, n18514, n18515, n18516, n18517, n18518,
    n18519, n18520, n18521, n18522, n18523, n18524,
    n18525, n18526, n18527, n18528, n18529, n18530,
    n18531, n18532, n18533, n18534, n18535, n18536,
    n18537, n18538, n18539, n18540, n18541, n18542,
    n18543, n18544, n18545, n18546, n18547, n18548,
    n18549, n18550, n18551, n18552, n18553, n18554,
    n18555, n18556, n18557, n18558, n18559;
  assign n193 = pi126  & pi127 ;
  assign n194 = ~pi124  & ~pi125 ;
  assign n195 = ~pi126  & ~n194;
  assign po62  = n193 | n195;
  assign n197 = pi126  & n194;
  assign n198 = pi127  & ~n195;
  assign n199 = ~n197 & n198;
  assign po63  = pi126  | pi127 ;
  assign n201 = ~pi124  & po62 ;
  assign n202 = pi125  & ~n201;
  assign n203 = n193 & n194;
  assign n204 = ~n202 & ~n203;
  assign n205 = pi124  & po62 ;
  assign n206 = ~pi122  & ~pi123 ;
  assign n207 = ~pi124  & n206;
  assign n208 = ~n205 & ~n207;
  assign n209 = n204 & ~n208;
  assign n210 = ~po63  & ~n209;
  assign n211 = ~n204 & n208;
  assign n212 = ~n199 & ~n211;
  assign po61  = n210 | ~n212;
  assign n214 = po62  & ~po61 ;
  assign n215 = ~pi122  & po61 ;
  assign n216 = ~pi123  & n215;
  assign n217 = ~n214 & ~n216;
  assign n218 = pi124  & ~n217;
  assign n219 = ~pi124  & n217;
  assign n220 = ~n218 & ~n219;
  assign n221 = pi122  & po61 ;
  assign n222 = ~pi120  & ~pi121 ;
  assign n223 = ~pi122  & n222;
  assign n224 = ~n221 & ~n223;
  assign n225 = po62  & ~n224;
  assign n226 = ~po62  & n224;
  assign n227 = pi123  & ~n215;
  assign n228 = ~n216 & ~n227;
  assign n229 = ~n226 & n228;
  assign n230 = ~n225 & ~n229;
  assign n231 = n220 & n230;
  assign n232 = ~n220 & ~n230;
  assign n233 = po63  & ~n231;
  assign n234 = ~n232 & n233;
  assign n235 = ~n204 & ~po61 ;
  assign n236 = n204 & po61 ;
  assign n237 = ~n208 & n236;
  assign n238 = ~n211 & ~n237;
  assign n239 = n232 & n238;
  assign n240 = ~po63  & ~n239;
  assign n241 = n208 & ~n236;
  assign n242 = po63  & ~n209;
  assign n243 = ~n241 & n242;
  assign n244 = ~n231 & ~n243;
  assign n245 = ~n240 & n244;
  assign po60  = n235 | ~n245;
  assign n247 = pi120  & po60 ;
  assign n248 = ~pi118  & ~pi119 ;
  assign n249 = ~pi120  & n248;
  assign n250 = ~n247 & ~n249;
  assign n251 = po61  & ~n250;
  assign n252 = ~po61  & n250;
  assign n253 = ~pi120  & po60 ;
  assign n254 = pi121  & ~n253;
  assign n255 = ~pi121  & n253;
  assign n256 = ~n254 & ~n255;
  assign n257 = ~n252 & n256;
  assign n258 = ~n251 & ~n257;
  assign n259 = po62  & ~n258;
  assign n260 = ~po62  & n258;
  assign n261 = po61  & n245;
  assign n262 = ~n255 & ~n261;
  assign n263 = pi122  & ~n262;
  assign n264 = ~pi122  & n262;
  assign n265 = ~n263 & ~n264;
  assign n266 = ~n260 & ~n265;
  assign n267 = ~n259 & ~n266;
  assign n268 = ~n225 & ~n226;
  assign n269 = po60  & n268;
  assign n270 = n228 & ~n269;
  assign n271 = ~n228 & n269;
  assign n272 = ~n270 & ~n271;
  assign n273 = n267 & n272;
  assign n274 = po63  & ~n273;
  assign n275 = n232 & po60 ;
  assign n276 = ~n267 & ~n272;
  assign n277 = ~n231 & ~n275;
  assign n278 = n276 & n277;
  assign n279 = ~n274 & ~n278;
  assign n280 = ~n234 & po60 ;
  assign n281 = ~n279 & n280;
  assign n282 = ~n220 & ~po60 ;
  assign n283 = ~n279 & n282;
  assign po59  = ~n281 & ~n283;
  assign n285 = ~pi118  & po59 ;
  assign n286 = ~pi119  & n285;
  assign n287 = ~n281 & ~n286;
  assign n288 = pi120  & ~n287;
  assign n289 = ~pi120  & n287;
  assign n290 = ~n288 & ~n289;
  assign n291 = pi118  & ~po59 ;
  assign n292 = ~pi116  & ~pi117 ;
  assign n293 = ~pi118  & ~n292;
  assign n294 = ~n291 & ~n293;
  assign n295 = po60  & n294;
  assign n296 = ~po60  & ~n294;
  assign n297 = pi119  & ~n285;
  assign n298 = ~n286 & ~n297;
  assign n299 = ~n296 & n298;
  assign n300 = ~n295 & ~n299;
  assign n301 = po61  & ~n300;
  assign n302 = ~po61  & n300;
  assign n303 = n272 & ~po59 ;
  assign n304 = ~n272 & ~po59 ;
  assign n305 = n274 & ~n276;
  assign n306 = ~n304 & n305;
  assign n307 = ~n259 & ~n260;
  assign n308 = po59  & n307;
  assign n309 = ~n265 & ~n308;
  assign n310 = n265 & n308;
  assign n311 = ~n309 & ~n310;
  assign n312 = ~n290 & ~n302;
  assign n313 = ~n301 & ~n312;
  assign n314 = po62  & ~n313;
  assign n315 = ~po62  & n313;
  assign n316 = ~n251 & ~n252;
  assign n317 = po59  & n316;
  assign n318 = n256 & ~n317;
  assign n319 = ~n256 & n317;
  assign n320 = ~n318 & ~n319;
  assign n321 = ~n315 & ~n320;
  assign n322 = ~n314 & ~n321;
  assign n323 = n311 & n322;
  assign n324 = ~n311 & ~n322;
  assign n325 = n276 & po59 ;
  assign n326 = ~n273 & ~n325;
  assign n327 = n324 & n326;
  assign n328 = ~po63  & ~n327;
  assign n329 = ~n306 & ~n323;
  assign n330 = ~n328 & n329;
  assign po58  = n303 | ~n330;
  assign n332 = ~n301 & ~n302;
  assign n333 = po58  & n332;
  assign n334 = ~n290 & ~n333;
  assign n335 = n290 & n333;
  assign n336 = ~n334 & ~n335;
  assign n337 = pi116  & po58 ;
  assign n338 = ~pi114  & ~pi115 ;
  assign n339 = ~pi116  & n338;
  assign n340 = ~n337 & ~n339;
  assign n341 = po59  & ~n340;
  assign n342 = ~po59  & n340;
  assign n343 = ~pi116  & po58 ;
  assign n344 = pi117  & ~n343;
  assign n345 = n292 & po58 ;
  assign n346 = ~n344 & ~n345;
  assign n347 = ~n342 & n346;
  assign n348 = ~n341 & ~n347;
  assign n349 = po60  & ~n348;
  assign n350 = ~po60  & n348;
  assign n351 = po59  & n330;
  assign n352 = ~n345 & ~n351;
  assign n353 = pi118  & ~n352;
  assign n354 = ~pi118  & n352;
  assign n355 = ~n353 & ~n354;
  assign n356 = ~n350 & ~n355;
  assign n357 = ~n349 & ~n356;
  assign n358 = po61  & ~n357;
  assign n359 = ~po61  & n357;
  assign n360 = ~n295 & ~n296;
  assign n361 = po58  & n360;
  assign n362 = n298 & ~n361;
  assign n363 = ~n298 & n361;
  assign n364 = ~n362 & ~n363;
  assign n365 = ~n359 & ~n364;
  assign n366 = ~n358 & ~n365;
  assign n367 = po62  & ~n366;
  assign n368 = ~po62  & n366;
  assign n369 = n311 & ~po58 ;
  assign n370 = ~n336 & ~n368;
  assign n371 = ~n367 & ~n370;
  assign n372 = ~n314 & ~n315;
  assign n373 = po58  & n372;
  assign n374 = n320 & n373;
  assign n375 = ~n320 & ~n373;
  assign n376 = ~n374 & ~n375;
  assign n377 = n371 & n376;
  assign n378 = ~n371 & ~n376;
  assign n379 = n324 & po58 ;
  assign n380 = ~n323 & ~n379;
  assign n381 = n378 & n380;
  assign n382 = ~po63  & ~n381;
  assign n383 = ~n311 & po58 ;
  assign n384 = n322 & ~n383;
  assign n385 = po63  & ~n324;
  assign n386 = ~n384 & n385;
  assign n387 = ~n377 & ~n386;
  assign n388 = ~n382 & n387;
  assign po57  = n369 | ~n388;
  assign n390 = ~n367 & ~n368;
  assign n391 = po57  & n390;
  assign n392 = ~n336 & ~n391;
  assign n393 = n336 & n391;
  assign n394 = ~n392 & ~n393;
  assign n395 = n376 & ~po57 ;
  assign n396 = pi114  & po57 ;
  assign n397 = ~pi112  & ~pi113 ;
  assign n398 = ~pi114  & n397;
  assign n399 = ~n396 & ~n398;
  assign n400 = po58  & ~n399;
  assign n401 = ~po58  & n399;
  assign n402 = ~pi114  & po57 ;
  assign n403 = pi115  & ~n402;
  assign n404 = ~pi115  & n402;
  assign n405 = ~n403 & ~n404;
  assign n406 = ~n401 & n405;
  assign n407 = ~n400 & ~n406;
  assign n408 = po59  & ~n407;
  assign n409 = ~po59  & n407;
  assign n410 = po58  & n388;
  assign n411 = ~n404 & ~n410;
  assign n412 = pi116  & ~n411;
  assign n413 = ~pi116  & n411;
  assign n414 = ~n412 & ~n413;
  assign n415 = ~n409 & ~n414;
  assign n416 = ~n408 & ~n415;
  assign n417 = po60  & ~n416;
  assign n418 = ~po60  & n416;
  assign n419 = ~n341 & ~n342;
  assign n420 = po57  & n419;
  assign n421 = n346 & ~n420;
  assign n422 = ~n346 & n420;
  assign n423 = ~n421 & ~n422;
  assign n424 = ~n418 & ~n423;
  assign n425 = ~n417 & ~n424;
  assign n426 = po61  & ~n425;
  assign n427 = ~po61  & n425;
  assign n428 = ~n349 & ~n350;
  assign n429 = po57  & n428;
  assign n430 = ~n355 & ~n429;
  assign n431 = n355 & n429;
  assign n432 = ~n430 & ~n431;
  assign n433 = ~n427 & ~n432;
  assign n434 = ~n426 & ~n433;
  assign n435 = po62  & ~n434;
  assign n436 = ~po62  & n434;
  assign n437 = ~n358 & ~n359;
  assign n438 = po57  & n437;
  assign n439 = n364 & n438;
  assign n440 = ~n364 & ~n438;
  assign n441 = ~n439 & ~n440;
  assign n442 = ~n436 & ~n441;
  assign n443 = ~n435 & ~n442;
  assign n444 = n394 & n443;
  assign n445 = ~n394 & ~n443;
  assign n446 = n378 & po57 ;
  assign n447 = ~n377 & ~n446;
  assign n448 = n445 & n447;
  assign n449 = ~po63  & ~n448;
  assign n450 = ~n376 & po57 ;
  assign n451 = n371 & ~n450;
  assign n452 = po63  & ~n378;
  assign n453 = ~n451 & n452;
  assign n454 = ~n444 & ~n453;
  assign n455 = ~n449 & n454;
  assign po56  = n395 | ~n455;
  assign n457 = n394 & ~po56 ;
  assign n458 = ~n435 & ~n436;
  assign n459 = po56  & n458;
  assign n460 = ~n441 & ~n459;
  assign n461 = n441 & n459;
  assign n462 = ~n460 & ~n461;
  assign n463 = pi112  & po56 ;
  assign n464 = ~pi110  & ~pi111 ;
  assign n465 = ~pi112  & n464;
  assign n466 = ~n463 & ~n465;
  assign n467 = po57  & ~n466;
  assign n468 = ~po57  & n466;
  assign n469 = ~pi112  & po56 ;
  assign n470 = pi113  & ~n469;
  assign n471 = ~pi113  & n469;
  assign n472 = ~n470 & ~n471;
  assign n473 = ~n468 & n472;
  assign n474 = ~n467 & ~n473;
  assign n475 = po58  & ~n474;
  assign n476 = ~po58  & n474;
  assign n477 = po57  & n455;
  assign n478 = ~n471 & ~n477;
  assign n479 = pi114  & ~n478;
  assign n480 = ~pi114  & n478;
  assign n481 = ~n479 & ~n480;
  assign n482 = ~n476 & ~n481;
  assign n483 = ~n475 & ~n482;
  assign n484 = po59  & ~n483;
  assign n485 = ~po59  & n483;
  assign n486 = ~n400 & ~n401;
  assign n487 = po56  & n486;
  assign n488 = n405 & ~n487;
  assign n489 = ~n405 & n487;
  assign n490 = ~n488 & ~n489;
  assign n491 = ~n485 & ~n490;
  assign n492 = ~n484 & ~n491;
  assign n493 = po60  & ~n492;
  assign n494 = ~po60  & n492;
  assign n495 = ~n408 & ~n409;
  assign n496 = po56  & n495;
  assign n497 = ~n414 & ~n496;
  assign n498 = n414 & n496;
  assign n499 = ~n497 & ~n498;
  assign n500 = ~n494 & ~n499;
  assign n501 = ~n493 & ~n500;
  assign n502 = po61  & ~n501;
  assign n503 = ~po61  & n501;
  assign n504 = ~n417 & ~n418;
  assign n505 = po56  & n504;
  assign n506 = n423 & n505;
  assign n507 = ~n423 & ~n505;
  assign n508 = ~n506 & ~n507;
  assign n509 = ~n503 & ~n508;
  assign n510 = ~n502 & ~n509;
  assign n511 = po62  & ~n510;
  assign n512 = ~po62  & n510;
  assign n513 = ~n426 & ~n427;
  assign n514 = po56  & n513;
  assign n515 = ~n432 & ~n514;
  assign n516 = n432 & n514;
  assign n517 = ~n515 & ~n516;
  assign n518 = ~n512 & ~n517;
  assign n519 = ~n511 & ~n518;
  assign n520 = n462 & n519;
  assign n521 = ~n462 & ~n519;
  assign n522 = n445 & po56 ;
  assign n523 = ~n444 & ~n522;
  assign n524 = n521 & n523;
  assign n525 = ~po63  & ~n524;
  assign n526 = ~n394 & po56 ;
  assign n527 = n443 & ~n526;
  assign n528 = po63  & ~n445;
  assign n529 = ~n527 & n528;
  assign n530 = ~n520 & ~n529;
  assign n531 = ~n525 & n530;
  assign po55  = n457 | ~n531;
  assign n533 = ~pi110  & po55 ;
  assign n534 = ~pi111  & n533;
  assign n535 = po56  & n531;
  assign n536 = ~n534 & ~n535;
  assign n537 = pi112  & ~n536;
  assign n538 = ~pi112  & n536;
  assign n539 = ~n537 & ~n538;
  assign n540 = pi110  & po55 ;
  assign n541 = ~pi108  & ~pi109 ;
  assign n542 = ~pi110  & n541;
  assign n543 = ~n540 & ~n542;
  assign n544 = po56  & ~n543;
  assign n545 = ~po56  & n543;
  assign n546 = pi111  & ~n533;
  assign n547 = ~n534 & ~n546;
  assign n548 = ~n545 & n547;
  assign n549 = ~n544 & ~n548;
  assign n550 = po57  & ~n549;
  assign n551 = ~po57  & n549;
  assign n552 = n462 & ~po55 ;
  assign n553 = ~n511 & ~n512;
  assign n554 = po55  & n553;
  assign n555 = ~n517 & ~n554;
  assign n556 = n517 & n554;
  assign n557 = ~n555 & ~n556;
  assign n558 = ~n539 & ~n551;
  assign n559 = ~n550 & ~n558;
  assign n560 = po58  & ~n559;
  assign n561 = ~po58  & n559;
  assign n562 = ~n467 & ~n468;
  assign n563 = po55  & n562;
  assign n564 = n472 & ~n563;
  assign n565 = ~n472 & n563;
  assign n566 = ~n564 & ~n565;
  assign n567 = ~n561 & ~n566;
  assign n568 = ~n560 & ~n567;
  assign n569 = po59  & ~n568;
  assign n570 = ~po59  & n568;
  assign n571 = ~n475 & ~n476;
  assign n572 = po55  & n571;
  assign n573 = ~n481 & ~n572;
  assign n574 = n481 & n572;
  assign n575 = ~n573 & ~n574;
  assign n576 = ~n570 & ~n575;
  assign n577 = ~n569 & ~n576;
  assign n578 = po60  & ~n577;
  assign n579 = ~po60  & n577;
  assign n580 = ~n484 & ~n485;
  assign n581 = po55  & n580;
  assign n582 = n490 & n581;
  assign n583 = ~n490 & ~n581;
  assign n584 = ~n582 & ~n583;
  assign n585 = ~n579 & ~n584;
  assign n586 = ~n578 & ~n585;
  assign n587 = po61  & ~n586;
  assign n588 = ~po61  & n586;
  assign n589 = ~n493 & ~n494;
  assign n590 = po55  & n589;
  assign n591 = ~n499 & ~n590;
  assign n592 = n499 & n590;
  assign n593 = ~n591 & ~n592;
  assign n594 = ~n588 & ~n593;
  assign n595 = ~n587 & ~n594;
  assign n596 = po62  & ~n595;
  assign n597 = ~po62  & n595;
  assign n598 = ~n502 & ~n503;
  assign n599 = po55  & n598;
  assign n600 = ~n508 & ~n599;
  assign n601 = n508 & n599;
  assign n602 = ~n600 & ~n601;
  assign n603 = ~n597 & ~n602;
  assign n604 = ~n596 & ~n603;
  assign n605 = n557 & n604;
  assign n606 = ~n557 & ~n604;
  assign n607 = n521 & po55 ;
  assign n608 = ~n520 & ~n607;
  assign n609 = n606 & n608;
  assign n610 = ~po63  & ~n609;
  assign n611 = ~n462 & po55 ;
  assign n612 = n519 & ~n611;
  assign n613 = po63  & ~n521;
  assign n614 = ~n612 & n613;
  assign n615 = ~n605 & ~n614;
  assign n616 = ~n610 & n615;
  assign po54  = n552 | ~n616;
  assign n618 = ~n550 & ~n551;
  assign n619 = po54  & n618;
  assign n620 = ~n539 & ~n619;
  assign n621 = n539 & n619;
  assign n622 = ~n620 & ~n621;
  assign n623 = pi108  & po54 ;
  assign n624 = ~pi106  & ~pi107 ;
  assign n625 = ~pi108  & n624;
  assign n626 = ~n623 & ~n625;
  assign n627 = po55  & ~n626;
  assign n628 = ~po55  & n626;
  assign n629 = ~pi108  & po54 ;
  assign n630 = pi109  & ~n629;
  assign n631 = ~pi109  & n629;
  assign n632 = ~n630 & ~n631;
  assign n633 = ~n628 & n632;
  assign n634 = ~n627 & ~n633;
  assign n635 = po56  & ~n634;
  assign n636 = ~po56  & n634;
  assign n637 = po55  & n616;
  assign n638 = ~n631 & ~n637;
  assign n639 = pi110  & ~n638;
  assign n640 = ~pi110  & n638;
  assign n641 = ~n639 & ~n640;
  assign n642 = ~n636 & ~n641;
  assign n643 = ~n635 & ~n642;
  assign n644 = po57  & ~n643;
  assign n645 = ~po57  & n643;
  assign n646 = ~n544 & ~n545;
  assign n647 = po54  & n646;
  assign n648 = n547 & ~n647;
  assign n649 = ~n547 & n647;
  assign n650 = ~n648 & ~n649;
  assign n651 = ~n645 & ~n650;
  assign n652 = ~n644 & ~n651;
  assign n653 = po58  & ~n652;
  assign n654 = ~po58  & n652;
  assign n655 = n557 & ~po54 ;
  assign n656 = ~n596 & ~n597;
  assign n657 = po54  & n656;
  assign n658 = ~n602 & ~n657;
  assign n659 = n602 & n657;
  assign n660 = ~n658 & ~n659;
  assign n661 = ~n622 & ~n654;
  assign n662 = ~n653 & ~n661;
  assign n663 = po59  & ~n662;
  assign n664 = ~po59  & n662;
  assign n665 = ~n560 & ~n561;
  assign n666 = po54  & n665;
  assign n667 = n566 & n666;
  assign n668 = ~n566 & ~n666;
  assign n669 = ~n667 & ~n668;
  assign n670 = ~n664 & ~n669;
  assign n671 = ~n663 & ~n670;
  assign n672 = po60  & ~n671;
  assign n673 = ~po60  & n671;
  assign n674 = ~n569 & ~n570;
  assign n675 = po54  & n674;
  assign n676 = ~n575 & ~n675;
  assign n677 = n575 & n675;
  assign n678 = ~n676 & ~n677;
  assign n679 = ~n673 & ~n678;
  assign n680 = ~n672 & ~n679;
  assign n681 = po61  & ~n680;
  assign n682 = ~po61  & n680;
  assign n683 = ~n578 & ~n579;
  assign n684 = po54  & n683;
  assign n685 = ~n584 & ~n684;
  assign n686 = n584 & n684;
  assign n687 = ~n685 & ~n686;
  assign n688 = ~n682 & ~n687;
  assign n689 = ~n681 & ~n688;
  assign n690 = po62  & ~n689;
  assign n691 = ~po62  & n689;
  assign n692 = ~n587 & ~n588;
  assign n693 = po54  & n692;
  assign n694 = ~n593 & ~n693;
  assign n695 = n593 & n693;
  assign n696 = ~n694 & ~n695;
  assign n697 = ~n691 & ~n696;
  assign n698 = ~n690 & ~n697;
  assign n699 = n660 & n698;
  assign n700 = ~n660 & ~n698;
  assign n701 = n606 & po54 ;
  assign n702 = ~n605 & ~n701;
  assign n703 = n700 & n702;
  assign n704 = ~po63  & ~n703;
  assign n705 = ~n557 & po54 ;
  assign n706 = n604 & ~n705;
  assign n707 = po63  & ~n606;
  assign n708 = ~n706 & n707;
  assign n709 = ~n699 & ~n708;
  assign n710 = ~n704 & n709;
  assign po53  = n655 | ~n710;
  assign n712 = ~n653 & ~n654;
  assign n713 = po53  & n712;
  assign n714 = ~n622 & ~n713;
  assign n715 = n622 & n713;
  assign n716 = ~n714 & ~n715;
  assign n717 = pi106  & po53 ;
  assign n718 = ~pi104  & ~pi105 ;
  assign n719 = ~pi106  & n718;
  assign n720 = ~n717 & ~n719;
  assign n721 = po54  & ~n720;
  assign n722 = ~po54  & n720;
  assign n723 = ~pi106  & po53 ;
  assign n724 = pi107  & ~n723;
  assign n725 = ~pi107  & n723;
  assign n726 = ~n724 & ~n725;
  assign n727 = ~n722 & n726;
  assign n728 = ~n721 & ~n727;
  assign n729 = po55  & ~n728;
  assign n730 = ~po55  & n728;
  assign n731 = po54  & n710;
  assign n732 = ~n725 & ~n731;
  assign n733 = pi108  & ~n732;
  assign n734 = ~pi108  & n732;
  assign n735 = ~n733 & ~n734;
  assign n736 = ~n730 & ~n735;
  assign n737 = ~n729 & ~n736;
  assign n738 = po56  & ~n737;
  assign n739 = ~po56  & n737;
  assign n740 = ~n627 & ~n628;
  assign n741 = po53  & n740;
  assign n742 = n632 & ~n741;
  assign n743 = ~n632 & n741;
  assign n744 = ~n742 & ~n743;
  assign n745 = ~n739 & ~n744;
  assign n746 = ~n738 & ~n745;
  assign n747 = po57  & ~n746;
  assign n748 = ~po57  & n746;
  assign n749 = ~n635 & ~n636;
  assign n750 = po53  & n749;
  assign n751 = ~n641 & ~n750;
  assign n752 = n641 & n750;
  assign n753 = ~n751 & ~n752;
  assign n754 = ~n748 & ~n753;
  assign n755 = ~n747 & ~n754;
  assign n756 = po58  & ~n755;
  assign n757 = ~po58  & n755;
  assign n758 = ~n644 & ~n645;
  assign n759 = po53  & n758;
  assign n760 = n650 & n759;
  assign n761 = ~n650 & ~n759;
  assign n762 = ~n760 & ~n761;
  assign n763 = ~n757 & ~n762;
  assign n764 = ~n756 & ~n763;
  assign n765 = po59  & ~n764;
  assign n766 = ~po59  & n764;
  assign n767 = n660 & ~po53 ;
  assign n768 = ~n690 & ~n691;
  assign n769 = po53  & n768;
  assign n770 = ~n696 & ~n769;
  assign n771 = n696 & n769;
  assign n772 = ~n770 & ~n771;
  assign n773 = ~n716 & ~n766;
  assign n774 = ~n765 & ~n773;
  assign n775 = po60  & ~n774;
  assign n776 = ~po60  & n774;
  assign n777 = ~n663 & ~n664;
  assign n778 = po53  & n777;
  assign n779 = ~n669 & ~n778;
  assign n780 = n669 & n778;
  assign n781 = ~n779 & ~n780;
  assign n782 = ~n776 & ~n781;
  assign n783 = ~n775 & ~n782;
  assign n784 = po61  & ~n783;
  assign n785 = ~po61  & n783;
  assign n786 = ~n672 & ~n673;
  assign n787 = po53  & n786;
  assign n788 = ~n678 & ~n787;
  assign n789 = n678 & n787;
  assign n790 = ~n788 & ~n789;
  assign n791 = ~n785 & ~n790;
  assign n792 = ~n784 & ~n791;
  assign n793 = po62  & ~n792;
  assign n794 = ~po62  & n792;
  assign n795 = ~n681 & ~n682;
  assign n796 = po53  & n795;
  assign n797 = ~n687 & ~n796;
  assign n798 = n687 & n796;
  assign n799 = ~n797 & ~n798;
  assign n800 = ~n794 & ~n799;
  assign n801 = ~n793 & ~n800;
  assign n802 = n772 & n801;
  assign n803 = ~n772 & ~n801;
  assign n804 = n700 & po53 ;
  assign n805 = ~n699 & ~n804;
  assign n806 = n803 & n805;
  assign n807 = ~po63  & ~n806;
  assign n808 = ~n660 & po53 ;
  assign n809 = n698 & ~n808;
  assign n810 = po63  & ~n700;
  assign n811 = ~n809 & n810;
  assign n812 = ~n802 & ~n811;
  assign n813 = ~n807 & n812;
  assign po52  = n767 | ~n813;
  assign n815 = ~n765 & ~n766;
  assign n816 = po52  & n815;
  assign n817 = ~n716 & ~n816;
  assign n818 = n716 & n816;
  assign n819 = ~n817 & ~n818;
  assign n820 = pi104  & po52 ;
  assign n821 = ~pi102  & ~pi103 ;
  assign n822 = ~pi104  & n821;
  assign n823 = ~n820 & ~n822;
  assign n824 = po53  & ~n823;
  assign n825 = ~po53  & n823;
  assign n826 = ~pi104  & po52 ;
  assign n827 = pi105  & ~n826;
  assign n828 = ~pi105  & n826;
  assign n829 = ~n827 & ~n828;
  assign n830 = ~n825 & n829;
  assign n831 = ~n824 & ~n830;
  assign n832 = po54  & ~n831;
  assign n833 = ~po54  & n831;
  assign n834 = po53  & n813;
  assign n835 = ~n828 & ~n834;
  assign n836 = pi106  & ~n835;
  assign n837 = ~pi106  & n835;
  assign n838 = ~n836 & ~n837;
  assign n839 = ~n833 & ~n838;
  assign n840 = ~n832 & ~n839;
  assign n841 = po55  & ~n840;
  assign n842 = ~po55  & n840;
  assign n843 = ~n721 & ~n722;
  assign n844 = po52  & n843;
  assign n845 = n726 & ~n844;
  assign n846 = ~n726 & n844;
  assign n847 = ~n845 & ~n846;
  assign n848 = ~n842 & ~n847;
  assign n849 = ~n841 & ~n848;
  assign n850 = po56  & ~n849;
  assign n851 = ~po56  & n849;
  assign n852 = ~n729 & ~n730;
  assign n853 = po52  & n852;
  assign n854 = ~n735 & ~n853;
  assign n855 = n735 & n853;
  assign n856 = ~n854 & ~n855;
  assign n857 = ~n851 & ~n856;
  assign n858 = ~n850 & ~n857;
  assign n859 = po57  & ~n858;
  assign n860 = ~po57  & n858;
  assign n861 = ~n738 & ~n739;
  assign n862 = po52  & n861;
  assign n863 = n744 & n862;
  assign n864 = ~n744 & ~n862;
  assign n865 = ~n863 & ~n864;
  assign n866 = ~n860 & ~n865;
  assign n867 = ~n859 & ~n866;
  assign n868 = po58  & ~n867;
  assign n869 = ~po58  & n867;
  assign n870 = ~n747 & ~n748;
  assign n871 = po52  & n870;
  assign n872 = ~n753 & ~n871;
  assign n873 = n753 & n871;
  assign n874 = ~n872 & ~n873;
  assign n875 = ~n869 & ~n874;
  assign n876 = ~n868 & ~n875;
  assign n877 = po59  & ~n876;
  assign n878 = ~po59  & n876;
  assign n879 = ~n756 & ~n757;
  assign n880 = po52  & n879;
  assign n881 = ~n762 & ~n880;
  assign n882 = n762 & n880;
  assign n883 = ~n881 & ~n882;
  assign n884 = ~n878 & ~n883;
  assign n885 = ~n877 & ~n884;
  assign n886 = po60  & ~n885;
  assign n887 = ~po60  & n885;
  assign n888 = n772 & ~po52 ;
  assign n889 = ~n793 & ~n794;
  assign n890 = po52  & n889;
  assign n891 = ~n799 & ~n890;
  assign n892 = n799 & n890;
  assign n893 = ~n891 & ~n892;
  assign n894 = ~n819 & ~n887;
  assign n895 = ~n886 & ~n894;
  assign n896 = po61  & ~n895;
  assign n897 = ~po61  & n895;
  assign n898 = ~n775 & ~n776;
  assign n899 = po52  & n898;
  assign n900 = ~n781 & ~n899;
  assign n901 = n781 & n899;
  assign n902 = ~n900 & ~n901;
  assign n903 = ~n897 & ~n902;
  assign n904 = ~n896 & ~n903;
  assign n905 = po62  & ~n904;
  assign n906 = ~po62  & n904;
  assign n907 = ~n784 & ~n785;
  assign n908 = po52  & n907;
  assign n909 = ~n790 & ~n908;
  assign n910 = n790 & n908;
  assign n911 = ~n909 & ~n910;
  assign n912 = ~n906 & ~n911;
  assign n913 = ~n905 & ~n912;
  assign n914 = n893 & n913;
  assign n915 = ~n893 & ~n913;
  assign n916 = n803 & po52 ;
  assign n917 = ~n802 & ~n916;
  assign n918 = n915 & n917;
  assign n919 = ~po63  & ~n918;
  assign n920 = ~n772 & po52 ;
  assign n921 = n801 & ~n920;
  assign n922 = po63  & ~n803;
  assign n923 = ~n921 & n922;
  assign n924 = ~n914 & ~n923;
  assign n925 = ~n919 & n924;
  assign po51  = n888 | ~n925;
  assign n927 = ~n886 & ~n887;
  assign n928 = po51  & n927;
  assign n929 = ~n819 & ~n928;
  assign n930 = n819 & n928;
  assign n931 = ~n929 & ~n930;
  assign n932 = pi102  & po51 ;
  assign n933 = ~pi100  & ~pi101 ;
  assign n934 = ~pi102  & n933;
  assign n935 = ~n932 & ~n934;
  assign n936 = po52  & ~n935;
  assign n937 = ~po52  & n935;
  assign n938 = ~pi102  & po51 ;
  assign n939 = pi103  & ~n938;
  assign n940 = ~pi103  & n938;
  assign n941 = ~n939 & ~n940;
  assign n942 = ~n937 & n941;
  assign n943 = ~n936 & ~n942;
  assign n944 = po53  & ~n943;
  assign n945 = ~po53  & n943;
  assign n946 = po52  & n925;
  assign n947 = ~n940 & ~n946;
  assign n948 = pi104  & ~n947;
  assign n949 = ~pi104  & n947;
  assign n950 = ~n948 & ~n949;
  assign n951 = ~n945 & ~n950;
  assign n952 = ~n944 & ~n951;
  assign n953 = po54  & ~n952;
  assign n954 = ~po54  & n952;
  assign n955 = ~n824 & ~n825;
  assign n956 = po51  & n955;
  assign n957 = n829 & ~n956;
  assign n958 = ~n829 & n956;
  assign n959 = ~n957 & ~n958;
  assign n960 = ~n954 & ~n959;
  assign n961 = ~n953 & ~n960;
  assign n962 = po55  & ~n961;
  assign n963 = ~po55  & n961;
  assign n964 = ~n832 & ~n833;
  assign n965 = po51  & n964;
  assign n966 = ~n838 & ~n965;
  assign n967 = n838 & n965;
  assign n968 = ~n966 & ~n967;
  assign n969 = ~n963 & ~n968;
  assign n970 = ~n962 & ~n969;
  assign n971 = po56  & ~n970;
  assign n972 = ~po56  & n970;
  assign n973 = ~n841 & ~n842;
  assign n974 = po51  & n973;
  assign n975 = n847 & n974;
  assign n976 = ~n847 & ~n974;
  assign n977 = ~n975 & ~n976;
  assign n978 = ~n972 & ~n977;
  assign n979 = ~n971 & ~n978;
  assign n980 = po57  & ~n979;
  assign n981 = ~po57  & n979;
  assign n982 = ~n850 & ~n851;
  assign n983 = po51  & n982;
  assign n984 = ~n856 & ~n983;
  assign n985 = n856 & n983;
  assign n986 = ~n984 & ~n985;
  assign n987 = ~n981 & ~n986;
  assign n988 = ~n980 & ~n987;
  assign n989 = po58  & ~n988;
  assign n990 = ~po58  & n988;
  assign n991 = ~n859 & ~n860;
  assign n992 = po51  & n991;
  assign n993 = ~n865 & ~n992;
  assign n994 = n865 & n992;
  assign n995 = ~n993 & ~n994;
  assign n996 = ~n990 & ~n995;
  assign n997 = ~n989 & ~n996;
  assign n998 = po59  & ~n997;
  assign n999 = ~po59  & n997;
  assign n1000 = ~n868 & ~n869;
  assign n1001 = po51  & n1000;
  assign n1002 = ~n874 & ~n1001;
  assign n1003 = n874 & n1001;
  assign n1004 = ~n1002 & ~n1003;
  assign n1005 = ~n999 & ~n1004;
  assign n1006 = ~n998 & ~n1005;
  assign n1007 = po60  & ~n1006;
  assign n1008 = ~po60  & n1006;
  assign n1009 = ~n877 & ~n878;
  assign n1010 = po51  & n1009;
  assign n1011 = ~n883 & ~n1010;
  assign n1012 = n883 & n1010;
  assign n1013 = ~n1011 & ~n1012;
  assign n1014 = ~n1008 & ~n1013;
  assign n1015 = ~n1007 & ~n1014;
  assign n1016 = po61  & ~n1015;
  assign n1017 = ~po61  & n1015;
  assign n1018 = n893 & ~po51 ;
  assign n1019 = ~n905 & ~n906;
  assign n1020 = po51  & n1019;
  assign n1021 = ~n911 & ~n1020;
  assign n1022 = n911 & n1020;
  assign n1023 = ~n1021 & ~n1022;
  assign n1024 = ~n931 & ~n1017;
  assign n1025 = ~n1016 & ~n1024;
  assign n1026 = po62  & ~n1025;
  assign n1027 = ~po62  & n1025;
  assign n1028 = ~n896 & ~n897;
  assign n1029 = po51  & n1028;
  assign n1030 = ~n902 & ~n1029;
  assign n1031 = n902 & n1029;
  assign n1032 = ~n1030 & ~n1031;
  assign n1033 = ~n1027 & ~n1032;
  assign n1034 = ~n1026 & ~n1033;
  assign n1035 = n1023 & n1034;
  assign n1036 = ~n1023 & ~n1034;
  assign n1037 = n915 & po51 ;
  assign n1038 = ~n914 & ~n1037;
  assign n1039 = n1036 & n1038;
  assign n1040 = ~po63  & ~n1039;
  assign n1041 = ~n893 & po51 ;
  assign n1042 = n913 & ~n1041;
  assign n1043 = po63  & ~n915;
  assign n1044 = ~n1042 & n1043;
  assign n1045 = ~n1035 & ~n1044;
  assign n1046 = ~n1040 & n1045;
  assign po50  = n1018 | ~n1046;
  assign n1048 = ~n1016 & ~n1017;
  assign n1049 = po50  & n1048;
  assign n1050 = ~n931 & ~n1049;
  assign n1051 = n931 & n1049;
  assign n1052 = ~n1050 & ~n1051;
  assign n1053 = pi100  & po50 ;
  assign n1054 = ~pi98  & ~pi99 ;
  assign n1055 = ~pi100  & n1054;
  assign n1056 = ~n1053 & ~n1055;
  assign n1057 = po51  & ~n1056;
  assign n1058 = ~po51  & n1056;
  assign n1059 = ~pi100  & po50 ;
  assign n1060 = pi101  & ~n1059;
  assign n1061 = ~pi101  & n1059;
  assign n1062 = ~n1060 & ~n1061;
  assign n1063 = ~n1058 & n1062;
  assign n1064 = ~n1057 & ~n1063;
  assign n1065 = po52  & ~n1064;
  assign n1066 = ~po52  & n1064;
  assign n1067 = po51  & n1046;
  assign n1068 = ~n1061 & ~n1067;
  assign n1069 = pi102  & ~n1068;
  assign n1070 = ~pi102  & n1068;
  assign n1071 = ~n1069 & ~n1070;
  assign n1072 = ~n1066 & ~n1071;
  assign n1073 = ~n1065 & ~n1072;
  assign n1074 = po53  & ~n1073;
  assign n1075 = ~po53  & n1073;
  assign n1076 = ~n936 & ~n937;
  assign n1077 = po50  & n1076;
  assign n1078 = n941 & ~n1077;
  assign n1079 = ~n941 & n1077;
  assign n1080 = ~n1078 & ~n1079;
  assign n1081 = ~n1075 & ~n1080;
  assign n1082 = ~n1074 & ~n1081;
  assign n1083 = po54  & ~n1082;
  assign n1084 = ~po54  & n1082;
  assign n1085 = ~n944 & ~n945;
  assign n1086 = po50  & n1085;
  assign n1087 = ~n950 & ~n1086;
  assign n1088 = n950 & n1086;
  assign n1089 = ~n1087 & ~n1088;
  assign n1090 = ~n1084 & ~n1089;
  assign n1091 = ~n1083 & ~n1090;
  assign n1092 = po55  & ~n1091;
  assign n1093 = ~po55  & n1091;
  assign n1094 = ~n953 & ~n954;
  assign n1095 = po50  & n1094;
  assign n1096 = n959 & n1095;
  assign n1097 = ~n959 & ~n1095;
  assign n1098 = ~n1096 & ~n1097;
  assign n1099 = ~n1093 & ~n1098;
  assign n1100 = ~n1092 & ~n1099;
  assign n1101 = po56  & ~n1100;
  assign n1102 = ~po56  & n1100;
  assign n1103 = ~n962 & ~n963;
  assign n1104 = po50  & n1103;
  assign n1105 = ~n968 & ~n1104;
  assign n1106 = n968 & n1104;
  assign n1107 = ~n1105 & ~n1106;
  assign n1108 = ~n1102 & ~n1107;
  assign n1109 = ~n1101 & ~n1108;
  assign n1110 = po57  & ~n1109;
  assign n1111 = ~po57  & n1109;
  assign n1112 = ~n971 & ~n972;
  assign n1113 = po50  & n1112;
  assign n1114 = ~n977 & ~n1113;
  assign n1115 = n977 & n1113;
  assign n1116 = ~n1114 & ~n1115;
  assign n1117 = ~n1111 & ~n1116;
  assign n1118 = ~n1110 & ~n1117;
  assign n1119 = po58  & ~n1118;
  assign n1120 = ~po58  & n1118;
  assign n1121 = ~n980 & ~n981;
  assign n1122 = po50  & n1121;
  assign n1123 = ~n986 & ~n1122;
  assign n1124 = n986 & n1122;
  assign n1125 = ~n1123 & ~n1124;
  assign n1126 = ~n1120 & ~n1125;
  assign n1127 = ~n1119 & ~n1126;
  assign n1128 = po59  & ~n1127;
  assign n1129 = ~po59  & n1127;
  assign n1130 = ~n989 & ~n990;
  assign n1131 = po50  & n1130;
  assign n1132 = ~n995 & ~n1131;
  assign n1133 = n995 & n1131;
  assign n1134 = ~n1132 & ~n1133;
  assign n1135 = ~n1129 & ~n1134;
  assign n1136 = ~n1128 & ~n1135;
  assign n1137 = po60  & ~n1136;
  assign n1138 = ~po60  & n1136;
  assign n1139 = ~n998 & ~n999;
  assign n1140 = po50  & n1139;
  assign n1141 = ~n1004 & ~n1140;
  assign n1142 = n1004 & n1140;
  assign n1143 = ~n1141 & ~n1142;
  assign n1144 = ~n1138 & ~n1143;
  assign n1145 = ~n1137 & ~n1144;
  assign n1146 = po61  & ~n1145;
  assign n1147 = ~po61  & n1145;
  assign n1148 = ~n1007 & ~n1008;
  assign n1149 = po50  & n1148;
  assign n1150 = ~n1013 & ~n1149;
  assign n1151 = n1013 & n1149;
  assign n1152 = ~n1150 & ~n1151;
  assign n1153 = ~n1147 & ~n1152;
  assign n1154 = ~n1146 & ~n1153;
  assign n1155 = po62  & ~n1154;
  assign n1156 = ~po62  & n1154;
  assign n1157 = n1023 & ~po50 ;
  assign n1158 = ~n1026 & ~n1027;
  assign n1159 = po50  & n1158;
  assign n1160 = ~n1032 & ~n1159;
  assign n1161 = n1032 & n1159;
  assign n1162 = ~n1160 & ~n1161;
  assign n1163 = ~n1052 & ~n1156;
  assign n1164 = ~n1155 & ~n1163;
  assign n1165 = n1162 & n1164;
  assign n1166 = ~n1162 & ~n1164;
  assign n1167 = n1036 & po50 ;
  assign n1168 = ~n1035 & ~n1167;
  assign n1169 = n1166 & n1168;
  assign n1170 = ~po63  & ~n1169;
  assign n1171 = ~n1023 & po50 ;
  assign n1172 = n1034 & ~n1171;
  assign n1173 = po63  & ~n1036;
  assign n1174 = ~n1172 & n1173;
  assign n1175 = ~n1165 & ~n1174;
  assign n1176 = ~n1170 & n1175;
  assign po49  = n1157 | ~n1176;
  assign n1178 = ~n1155 & ~n1156;
  assign n1179 = po49  & n1178;
  assign n1180 = ~n1052 & ~n1179;
  assign n1181 = n1052 & n1179;
  assign n1182 = ~n1180 & ~n1181;
  assign n1183 = n1162 & ~po49 ;
  assign n1184 = pi98  & po49 ;
  assign n1185 = ~pi96  & ~pi97 ;
  assign n1186 = ~pi98  & n1185;
  assign n1187 = ~n1184 & ~n1186;
  assign n1188 = po50  & ~n1187;
  assign n1189 = ~po50  & n1187;
  assign n1190 = ~pi98  & po49 ;
  assign n1191 = pi99  & ~n1190;
  assign n1192 = ~pi99  & n1190;
  assign n1193 = ~n1191 & ~n1192;
  assign n1194 = ~n1189 & n1193;
  assign n1195 = ~n1188 & ~n1194;
  assign n1196 = po51  & ~n1195;
  assign n1197 = ~po51  & n1195;
  assign n1198 = po50  & n1176;
  assign n1199 = ~n1192 & ~n1198;
  assign n1200 = pi100  & ~n1199;
  assign n1201 = ~pi100  & n1199;
  assign n1202 = ~n1200 & ~n1201;
  assign n1203 = ~n1197 & ~n1202;
  assign n1204 = ~n1196 & ~n1203;
  assign n1205 = po52  & ~n1204;
  assign n1206 = ~po52  & n1204;
  assign n1207 = ~n1057 & ~n1058;
  assign n1208 = po49  & n1207;
  assign n1209 = n1062 & ~n1208;
  assign n1210 = ~n1062 & n1208;
  assign n1211 = ~n1209 & ~n1210;
  assign n1212 = ~n1206 & ~n1211;
  assign n1213 = ~n1205 & ~n1212;
  assign n1214 = po53  & ~n1213;
  assign n1215 = ~po53  & n1213;
  assign n1216 = ~n1065 & ~n1066;
  assign n1217 = po49  & n1216;
  assign n1218 = ~n1071 & ~n1217;
  assign n1219 = n1071 & n1217;
  assign n1220 = ~n1218 & ~n1219;
  assign n1221 = ~n1215 & ~n1220;
  assign n1222 = ~n1214 & ~n1221;
  assign n1223 = po54  & ~n1222;
  assign n1224 = ~po54  & n1222;
  assign n1225 = ~n1074 & ~n1075;
  assign n1226 = po49  & n1225;
  assign n1227 = n1080 & n1226;
  assign n1228 = ~n1080 & ~n1226;
  assign n1229 = ~n1227 & ~n1228;
  assign n1230 = ~n1224 & ~n1229;
  assign n1231 = ~n1223 & ~n1230;
  assign n1232 = po55  & ~n1231;
  assign n1233 = ~po55  & n1231;
  assign n1234 = ~n1083 & ~n1084;
  assign n1235 = po49  & n1234;
  assign n1236 = ~n1089 & ~n1235;
  assign n1237 = n1089 & n1235;
  assign n1238 = ~n1236 & ~n1237;
  assign n1239 = ~n1233 & ~n1238;
  assign n1240 = ~n1232 & ~n1239;
  assign n1241 = po56  & ~n1240;
  assign n1242 = ~po56  & n1240;
  assign n1243 = ~n1092 & ~n1093;
  assign n1244 = po49  & n1243;
  assign n1245 = ~n1098 & ~n1244;
  assign n1246 = n1098 & n1244;
  assign n1247 = ~n1245 & ~n1246;
  assign n1248 = ~n1242 & ~n1247;
  assign n1249 = ~n1241 & ~n1248;
  assign n1250 = po57  & ~n1249;
  assign n1251 = ~po57  & n1249;
  assign n1252 = ~n1101 & ~n1102;
  assign n1253 = po49  & n1252;
  assign n1254 = ~n1107 & ~n1253;
  assign n1255 = n1107 & n1253;
  assign n1256 = ~n1254 & ~n1255;
  assign n1257 = ~n1251 & ~n1256;
  assign n1258 = ~n1250 & ~n1257;
  assign n1259 = po58  & ~n1258;
  assign n1260 = ~po58  & n1258;
  assign n1261 = ~n1110 & ~n1111;
  assign n1262 = po49  & n1261;
  assign n1263 = ~n1116 & ~n1262;
  assign n1264 = n1116 & n1262;
  assign n1265 = ~n1263 & ~n1264;
  assign n1266 = ~n1260 & ~n1265;
  assign n1267 = ~n1259 & ~n1266;
  assign n1268 = po59  & ~n1267;
  assign n1269 = ~po59  & n1267;
  assign n1270 = ~n1119 & ~n1120;
  assign n1271 = po49  & n1270;
  assign n1272 = ~n1125 & ~n1271;
  assign n1273 = n1125 & n1271;
  assign n1274 = ~n1272 & ~n1273;
  assign n1275 = ~n1269 & ~n1274;
  assign n1276 = ~n1268 & ~n1275;
  assign n1277 = po60  & ~n1276;
  assign n1278 = ~po60  & n1276;
  assign n1279 = ~n1128 & ~n1129;
  assign n1280 = po49  & n1279;
  assign n1281 = ~n1134 & ~n1280;
  assign n1282 = n1134 & n1280;
  assign n1283 = ~n1281 & ~n1282;
  assign n1284 = ~n1278 & ~n1283;
  assign n1285 = ~n1277 & ~n1284;
  assign n1286 = po61  & ~n1285;
  assign n1287 = ~po61  & n1285;
  assign n1288 = ~n1137 & ~n1138;
  assign n1289 = po49  & n1288;
  assign n1290 = ~n1143 & ~n1289;
  assign n1291 = n1143 & n1289;
  assign n1292 = ~n1290 & ~n1291;
  assign n1293 = ~n1287 & ~n1292;
  assign n1294 = ~n1286 & ~n1293;
  assign n1295 = po62  & ~n1294;
  assign n1296 = ~po62  & n1294;
  assign n1297 = ~n1146 & ~n1147;
  assign n1298 = po49  & n1297;
  assign n1299 = ~n1152 & ~n1298;
  assign n1300 = n1152 & n1298;
  assign n1301 = ~n1299 & ~n1300;
  assign n1302 = ~n1296 & ~n1301;
  assign n1303 = ~n1295 & ~n1302;
  assign n1304 = n1182 & n1303;
  assign n1305 = ~n1182 & ~n1303;
  assign n1306 = n1166 & po49 ;
  assign n1307 = ~n1165 & ~n1306;
  assign n1308 = n1305 & n1307;
  assign n1309 = ~po63  & ~n1308;
  assign n1310 = ~n1162 & po49 ;
  assign n1311 = n1164 & ~n1310;
  assign n1312 = po63  & ~n1166;
  assign n1313 = ~n1311 & n1312;
  assign n1314 = ~n1304 & ~n1313;
  assign n1315 = ~n1309 & n1314;
  assign po48  = n1183 | ~n1315;
  assign n1317 = n1182 & ~po48 ;
  assign n1318 = ~n1295 & ~n1296;
  assign n1319 = po48  & n1318;
  assign n1320 = ~n1301 & ~n1319;
  assign n1321 = n1301 & n1319;
  assign n1322 = ~n1320 & ~n1321;
  assign n1323 = pi96  & po48 ;
  assign n1324 = ~pi94  & ~pi95 ;
  assign n1325 = ~pi96  & n1324;
  assign n1326 = ~n1323 & ~n1325;
  assign n1327 = po49  & ~n1326;
  assign n1328 = ~po49  & n1326;
  assign n1329 = ~pi96  & po48 ;
  assign n1330 = pi97  & ~n1329;
  assign n1331 = ~pi97  & n1329;
  assign n1332 = ~n1330 & ~n1331;
  assign n1333 = ~n1328 & n1332;
  assign n1334 = ~n1327 & ~n1333;
  assign n1335 = po50  & ~n1334;
  assign n1336 = ~po50  & n1334;
  assign n1337 = po49  & n1315;
  assign n1338 = ~n1331 & ~n1337;
  assign n1339 = pi98  & ~n1338;
  assign n1340 = ~pi98  & n1338;
  assign n1341 = ~n1339 & ~n1340;
  assign n1342 = ~n1336 & ~n1341;
  assign n1343 = ~n1335 & ~n1342;
  assign n1344 = po51  & ~n1343;
  assign n1345 = ~po51  & n1343;
  assign n1346 = ~n1188 & ~n1189;
  assign n1347 = po48  & n1346;
  assign n1348 = n1193 & ~n1347;
  assign n1349 = ~n1193 & n1347;
  assign n1350 = ~n1348 & ~n1349;
  assign n1351 = ~n1345 & ~n1350;
  assign n1352 = ~n1344 & ~n1351;
  assign n1353 = po52  & ~n1352;
  assign n1354 = ~po52  & n1352;
  assign n1355 = ~n1196 & ~n1197;
  assign n1356 = po48  & n1355;
  assign n1357 = ~n1202 & ~n1356;
  assign n1358 = n1202 & n1356;
  assign n1359 = ~n1357 & ~n1358;
  assign n1360 = ~n1354 & ~n1359;
  assign n1361 = ~n1353 & ~n1360;
  assign n1362 = po53  & ~n1361;
  assign n1363 = ~po53  & n1361;
  assign n1364 = ~n1205 & ~n1206;
  assign n1365 = po48  & n1364;
  assign n1366 = n1211 & n1365;
  assign n1367 = ~n1211 & ~n1365;
  assign n1368 = ~n1366 & ~n1367;
  assign n1369 = ~n1363 & ~n1368;
  assign n1370 = ~n1362 & ~n1369;
  assign n1371 = po54  & ~n1370;
  assign n1372 = ~po54  & n1370;
  assign n1373 = ~n1214 & ~n1215;
  assign n1374 = po48  & n1373;
  assign n1375 = ~n1220 & ~n1374;
  assign n1376 = n1220 & n1374;
  assign n1377 = ~n1375 & ~n1376;
  assign n1378 = ~n1372 & ~n1377;
  assign n1379 = ~n1371 & ~n1378;
  assign n1380 = po55  & ~n1379;
  assign n1381 = ~po55  & n1379;
  assign n1382 = ~n1223 & ~n1224;
  assign n1383 = po48  & n1382;
  assign n1384 = ~n1229 & ~n1383;
  assign n1385 = n1229 & n1383;
  assign n1386 = ~n1384 & ~n1385;
  assign n1387 = ~n1381 & ~n1386;
  assign n1388 = ~n1380 & ~n1387;
  assign n1389 = po56  & ~n1388;
  assign n1390 = ~po56  & n1388;
  assign n1391 = ~n1232 & ~n1233;
  assign n1392 = po48  & n1391;
  assign n1393 = ~n1238 & ~n1392;
  assign n1394 = n1238 & n1392;
  assign n1395 = ~n1393 & ~n1394;
  assign n1396 = ~n1390 & ~n1395;
  assign n1397 = ~n1389 & ~n1396;
  assign n1398 = po57  & ~n1397;
  assign n1399 = ~po57  & n1397;
  assign n1400 = ~n1241 & ~n1242;
  assign n1401 = po48  & n1400;
  assign n1402 = ~n1247 & ~n1401;
  assign n1403 = n1247 & n1401;
  assign n1404 = ~n1402 & ~n1403;
  assign n1405 = ~n1399 & ~n1404;
  assign n1406 = ~n1398 & ~n1405;
  assign n1407 = po58  & ~n1406;
  assign n1408 = ~po58  & n1406;
  assign n1409 = ~n1250 & ~n1251;
  assign n1410 = po48  & n1409;
  assign n1411 = ~n1256 & ~n1410;
  assign n1412 = n1256 & n1410;
  assign n1413 = ~n1411 & ~n1412;
  assign n1414 = ~n1408 & ~n1413;
  assign n1415 = ~n1407 & ~n1414;
  assign n1416 = po59  & ~n1415;
  assign n1417 = ~po59  & n1415;
  assign n1418 = ~n1259 & ~n1260;
  assign n1419 = po48  & n1418;
  assign n1420 = ~n1265 & ~n1419;
  assign n1421 = n1265 & n1419;
  assign n1422 = ~n1420 & ~n1421;
  assign n1423 = ~n1417 & ~n1422;
  assign n1424 = ~n1416 & ~n1423;
  assign n1425 = po60  & ~n1424;
  assign n1426 = ~po60  & n1424;
  assign n1427 = ~n1268 & ~n1269;
  assign n1428 = po48  & n1427;
  assign n1429 = ~n1274 & ~n1428;
  assign n1430 = n1274 & n1428;
  assign n1431 = ~n1429 & ~n1430;
  assign n1432 = ~n1426 & ~n1431;
  assign n1433 = ~n1425 & ~n1432;
  assign n1434 = po61  & ~n1433;
  assign n1435 = ~po61  & n1433;
  assign n1436 = ~n1277 & ~n1278;
  assign n1437 = po48  & n1436;
  assign n1438 = ~n1283 & ~n1437;
  assign n1439 = n1283 & n1437;
  assign n1440 = ~n1438 & ~n1439;
  assign n1441 = ~n1435 & ~n1440;
  assign n1442 = ~n1434 & ~n1441;
  assign n1443 = po62  & ~n1442;
  assign n1444 = ~po62  & n1442;
  assign n1445 = ~n1286 & ~n1287;
  assign n1446 = po48  & n1445;
  assign n1447 = ~n1292 & ~n1446;
  assign n1448 = n1292 & n1446;
  assign n1449 = ~n1447 & ~n1448;
  assign n1450 = ~n1444 & ~n1449;
  assign n1451 = ~n1443 & ~n1450;
  assign n1452 = n1322 & n1451;
  assign n1453 = ~n1322 & ~n1451;
  assign n1454 = n1305 & po48 ;
  assign n1455 = ~n1304 & ~n1454;
  assign n1456 = n1453 & n1455;
  assign n1457 = ~po63  & ~n1456;
  assign n1458 = ~n1182 & po48 ;
  assign n1459 = n1303 & ~n1458;
  assign n1460 = po63  & ~n1305;
  assign n1461 = ~n1459 & n1460;
  assign n1462 = ~n1452 & ~n1461;
  assign n1463 = ~n1457 & n1462;
  assign po47  = n1317 | ~n1463;
  assign n1465 = ~pi94  & po47 ;
  assign n1466 = ~pi95  & n1465;
  assign n1467 = po48  & n1463;
  assign n1468 = ~n1466 & ~n1467;
  assign n1469 = pi96  & ~n1468;
  assign n1470 = ~pi96  & n1468;
  assign n1471 = ~n1469 & ~n1470;
  assign n1472 = pi94  & po47 ;
  assign n1473 = ~pi92  & ~pi93 ;
  assign n1474 = ~pi94  & n1473;
  assign n1475 = ~n1472 & ~n1474;
  assign n1476 = po48  & ~n1475;
  assign n1477 = ~po48  & n1475;
  assign n1478 = pi95  & ~n1465;
  assign n1479 = ~n1466 & ~n1478;
  assign n1480 = ~n1477 & n1479;
  assign n1481 = ~n1476 & ~n1480;
  assign n1482 = po49  & ~n1481;
  assign n1483 = ~po49  & n1481;
  assign n1484 = n1322 & ~po47 ;
  assign n1485 = ~n1443 & ~n1444;
  assign n1486 = po47  & n1485;
  assign n1487 = ~n1449 & ~n1486;
  assign n1488 = n1449 & n1486;
  assign n1489 = ~n1487 & ~n1488;
  assign n1490 = ~n1471 & ~n1483;
  assign n1491 = ~n1482 & ~n1490;
  assign n1492 = po50  & ~n1491;
  assign n1493 = ~po50  & n1491;
  assign n1494 = ~n1327 & ~n1328;
  assign n1495 = po47  & n1494;
  assign n1496 = n1332 & ~n1495;
  assign n1497 = ~n1332 & n1495;
  assign n1498 = ~n1496 & ~n1497;
  assign n1499 = ~n1493 & ~n1498;
  assign n1500 = ~n1492 & ~n1499;
  assign n1501 = po51  & ~n1500;
  assign n1502 = ~po51  & n1500;
  assign n1503 = ~n1335 & ~n1336;
  assign n1504 = po47  & n1503;
  assign n1505 = ~n1341 & ~n1504;
  assign n1506 = n1341 & n1504;
  assign n1507 = ~n1505 & ~n1506;
  assign n1508 = ~n1502 & ~n1507;
  assign n1509 = ~n1501 & ~n1508;
  assign n1510 = po52  & ~n1509;
  assign n1511 = ~po52  & n1509;
  assign n1512 = ~n1344 & ~n1345;
  assign n1513 = po47  & n1512;
  assign n1514 = n1350 & n1513;
  assign n1515 = ~n1350 & ~n1513;
  assign n1516 = ~n1514 & ~n1515;
  assign n1517 = ~n1511 & ~n1516;
  assign n1518 = ~n1510 & ~n1517;
  assign n1519 = po53  & ~n1518;
  assign n1520 = ~po53  & n1518;
  assign n1521 = ~n1353 & ~n1354;
  assign n1522 = po47  & n1521;
  assign n1523 = ~n1359 & ~n1522;
  assign n1524 = n1359 & n1522;
  assign n1525 = ~n1523 & ~n1524;
  assign n1526 = ~n1520 & ~n1525;
  assign n1527 = ~n1519 & ~n1526;
  assign n1528 = po54  & ~n1527;
  assign n1529 = ~po54  & n1527;
  assign n1530 = ~n1362 & ~n1363;
  assign n1531 = po47  & n1530;
  assign n1532 = ~n1368 & ~n1531;
  assign n1533 = n1368 & n1531;
  assign n1534 = ~n1532 & ~n1533;
  assign n1535 = ~n1529 & ~n1534;
  assign n1536 = ~n1528 & ~n1535;
  assign n1537 = po55  & ~n1536;
  assign n1538 = ~po55  & n1536;
  assign n1539 = ~n1371 & ~n1372;
  assign n1540 = po47  & n1539;
  assign n1541 = ~n1377 & ~n1540;
  assign n1542 = n1377 & n1540;
  assign n1543 = ~n1541 & ~n1542;
  assign n1544 = ~n1538 & ~n1543;
  assign n1545 = ~n1537 & ~n1544;
  assign n1546 = po56  & ~n1545;
  assign n1547 = ~po56  & n1545;
  assign n1548 = ~n1380 & ~n1381;
  assign n1549 = po47  & n1548;
  assign n1550 = ~n1386 & ~n1549;
  assign n1551 = n1386 & n1549;
  assign n1552 = ~n1550 & ~n1551;
  assign n1553 = ~n1547 & ~n1552;
  assign n1554 = ~n1546 & ~n1553;
  assign n1555 = po57  & ~n1554;
  assign n1556 = ~po57  & n1554;
  assign n1557 = ~n1389 & ~n1390;
  assign n1558 = po47  & n1557;
  assign n1559 = ~n1395 & ~n1558;
  assign n1560 = n1395 & n1558;
  assign n1561 = ~n1559 & ~n1560;
  assign n1562 = ~n1556 & ~n1561;
  assign n1563 = ~n1555 & ~n1562;
  assign n1564 = po58  & ~n1563;
  assign n1565 = ~po58  & n1563;
  assign n1566 = ~n1398 & ~n1399;
  assign n1567 = po47  & n1566;
  assign n1568 = ~n1404 & ~n1567;
  assign n1569 = n1404 & n1567;
  assign n1570 = ~n1568 & ~n1569;
  assign n1571 = ~n1565 & ~n1570;
  assign n1572 = ~n1564 & ~n1571;
  assign n1573 = po59  & ~n1572;
  assign n1574 = ~po59  & n1572;
  assign n1575 = ~n1407 & ~n1408;
  assign n1576 = po47  & n1575;
  assign n1577 = ~n1413 & ~n1576;
  assign n1578 = n1413 & n1576;
  assign n1579 = ~n1577 & ~n1578;
  assign n1580 = ~n1574 & ~n1579;
  assign n1581 = ~n1573 & ~n1580;
  assign n1582 = po60  & ~n1581;
  assign n1583 = ~po60  & n1581;
  assign n1584 = ~n1416 & ~n1417;
  assign n1585 = po47  & n1584;
  assign n1586 = ~n1422 & ~n1585;
  assign n1587 = n1422 & n1585;
  assign n1588 = ~n1586 & ~n1587;
  assign n1589 = ~n1583 & ~n1588;
  assign n1590 = ~n1582 & ~n1589;
  assign n1591 = po61  & ~n1590;
  assign n1592 = ~po61  & n1590;
  assign n1593 = ~n1425 & ~n1426;
  assign n1594 = po47  & n1593;
  assign n1595 = ~n1431 & ~n1594;
  assign n1596 = n1431 & n1594;
  assign n1597 = ~n1595 & ~n1596;
  assign n1598 = ~n1592 & ~n1597;
  assign n1599 = ~n1591 & ~n1598;
  assign n1600 = po62  & ~n1599;
  assign n1601 = ~po62  & n1599;
  assign n1602 = ~n1434 & ~n1435;
  assign n1603 = po47  & n1602;
  assign n1604 = ~n1440 & ~n1603;
  assign n1605 = n1440 & n1603;
  assign n1606 = ~n1604 & ~n1605;
  assign n1607 = ~n1601 & ~n1606;
  assign n1608 = ~n1600 & ~n1607;
  assign n1609 = n1489 & n1608;
  assign n1610 = ~n1489 & ~n1608;
  assign n1611 = n1453 & po47 ;
  assign n1612 = ~n1452 & ~n1611;
  assign n1613 = n1610 & n1612;
  assign n1614 = ~po63  & ~n1613;
  assign n1615 = ~n1322 & po47 ;
  assign n1616 = n1451 & ~n1615;
  assign n1617 = po63  & ~n1453;
  assign n1618 = ~n1616 & n1617;
  assign n1619 = ~n1609 & ~n1618;
  assign n1620 = ~n1614 & n1619;
  assign po46  = n1484 | ~n1620;
  assign n1622 = ~n1482 & ~n1483;
  assign n1623 = po46  & n1622;
  assign n1624 = ~n1471 & ~n1623;
  assign n1625 = n1471 & n1623;
  assign n1626 = ~n1624 & ~n1625;
  assign n1627 = pi92  & po46 ;
  assign n1628 = ~pi90  & ~pi91 ;
  assign n1629 = ~pi92  & n1628;
  assign n1630 = ~n1627 & ~n1629;
  assign n1631 = po47  & ~n1630;
  assign n1632 = ~po47  & n1630;
  assign n1633 = ~pi92  & po46 ;
  assign n1634 = pi93  & ~n1633;
  assign n1635 = ~pi93  & n1633;
  assign n1636 = ~n1634 & ~n1635;
  assign n1637 = ~n1632 & n1636;
  assign n1638 = ~n1631 & ~n1637;
  assign n1639 = po48  & ~n1638;
  assign n1640 = ~po48  & n1638;
  assign n1641 = po47  & n1620;
  assign n1642 = ~n1635 & ~n1641;
  assign n1643 = pi94  & ~n1642;
  assign n1644 = ~pi94  & n1642;
  assign n1645 = ~n1643 & ~n1644;
  assign n1646 = ~n1640 & ~n1645;
  assign n1647 = ~n1639 & ~n1646;
  assign n1648 = po49  & ~n1647;
  assign n1649 = ~po49  & n1647;
  assign n1650 = ~n1476 & ~n1477;
  assign n1651 = po46  & n1650;
  assign n1652 = n1479 & ~n1651;
  assign n1653 = ~n1479 & n1651;
  assign n1654 = ~n1652 & ~n1653;
  assign n1655 = ~n1649 & ~n1654;
  assign n1656 = ~n1648 & ~n1655;
  assign n1657 = po50  & ~n1656;
  assign n1658 = ~po50  & n1656;
  assign n1659 = n1489 & ~po46 ;
  assign n1660 = ~n1600 & ~n1601;
  assign n1661 = po46  & n1660;
  assign n1662 = ~n1606 & ~n1661;
  assign n1663 = n1606 & n1661;
  assign n1664 = ~n1662 & ~n1663;
  assign n1665 = ~n1626 & ~n1658;
  assign n1666 = ~n1657 & ~n1665;
  assign n1667 = po51  & ~n1666;
  assign n1668 = ~po51  & n1666;
  assign n1669 = ~n1492 & ~n1493;
  assign n1670 = po46  & n1669;
  assign n1671 = n1498 & n1670;
  assign n1672 = ~n1498 & ~n1670;
  assign n1673 = ~n1671 & ~n1672;
  assign n1674 = ~n1668 & ~n1673;
  assign n1675 = ~n1667 & ~n1674;
  assign n1676 = po52  & ~n1675;
  assign n1677 = ~po52  & n1675;
  assign n1678 = ~n1501 & ~n1502;
  assign n1679 = po46  & n1678;
  assign n1680 = ~n1507 & ~n1679;
  assign n1681 = n1507 & n1679;
  assign n1682 = ~n1680 & ~n1681;
  assign n1683 = ~n1677 & ~n1682;
  assign n1684 = ~n1676 & ~n1683;
  assign n1685 = po53  & ~n1684;
  assign n1686 = ~po53  & n1684;
  assign n1687 = ~n1510 & ~n1511;
  assign n1688 = po46  & n1687;
  assign n1689 = ~n1516 & ~n1688;
  assign n1690 = n1516 & n1688;
  assign n1691 = ~n1689 & ~n1690;
  assign n1692 = ~n1686 & ~n1691;
  assign n1693 = ~n1685 & ~n1692;
  assign n1694 = po54  & ~n1693;
  assign n1695 = ~po54  & n1693;
  assign n1696 = ~n1519 & ~n1520;
  assign n1697 = po46  & n1696;
  assign n1698 = ~n1525 & ~n1697;
  assign n1699 = n1525 & n1697;
  assign n1700 = ~n1698 & ~n1699;
  assign n1701 = ~n1695 & ~n1700;
  assign n1702 = ~n1694 & ~n1701;
  assign n1703 = po55  & ~n1702;
  assign n1704 = ~po55  & n1702;
  assign n1705 = ~n1528 & ~n1529;
  assign n1706 = po46  & n1705;
  assign n1707 = ~n1534 & ~n1706;
  assign n1708 = n1534 & n1706;
  assign n1709 = ~n1707 & ~n1708;
  assign n1710 = ~n1704 & ~n1709;
  assign n1711 = ~n1703 & ~n1710;
  assign n1712 = po56  & ~n1711;
  assign n1713 = ~po56  & n1711;
  assign n1714 = ~n1537 & ~n1538;
  assign n1715 = po46  & n1714;
  assign n1716 = ~n1543 & ~n1715;
  assign n1717 = n1543 & n1715;
  assign n1718 = ~n1716 & ~n1717;
  assign n1719 = ~n1713 & ~n1718;
  assign n1720 = ~n1712 & ~n1719;
  assign n1721 = po57  & ~n1720;
  assign n1722 = ~po57  & n1720;
  assign n1723 = ~n1546 & ~n1547;
  assign n1724 = po46  & n1723;
  assign n1725 = ~n1552 & ~n1724;
  assign n1726 = n1552 & n1724;
  assign n1727 = ~n1725 & ~n1726;
  assign n1728 = ~n1722 & ~n1727;
  assign n1729 = ~n1721 & ~n1728;
  assign n1730 = po58  & ~n1729;
  assign n1731 = ~po58  & n1729;
  assign n1732 = ~n1555 & ~n1556;
  assign n1733 = po46  & n1732;
  assign n1734 = ~n1561 & ~n1733;
  assign n1735 = n1561 & n1733;
  assign n1736 = ~n1734 & ~n1735;
  assign n1737 = ~n1731 & ~n1736;
  assign n1738 = ~n1730 & ~n1737;
  assign n1739 = po59  & ~n1738;
  assign n1740 = ~po59  & n1738;
  assign n1741 = ~n1564 & ~n1565;
  assign n1742 = po46  & n1741;
  assign n1743 = ~n1570 & ~n1742;
  assign n1744 = n1570 & n1742;
  assign n1745 = ~n1743 & ~n1744;
  assign n1746 = ~n1740 & ~n1745;
  assign n1747 = ~n1739 & ~n1746;
  assign n1748 = po60  & ~n1747;
  assign n1749 = ~po60  & n1747;
  assign n1750 = ~n1573 & ~n1574;
  assign n1751 = po46  & n1750;
  assign n1752 = ~n1579 & ~n1751;
  assign n1753 = n1579 & n1751;
  assign n1754 = ~n1752 & ~n1753;
  assign n1755 = ~n1749 & ~n1754;
  assign n1756 = ~n1748 & ~n1755;
  assign n1757 = po61  & ~n1756;
  assign n1758 = ~po61  & n1756;
  assign n1759 = ~n1582 & ~n1583;
  assign n1760 = po46  & n1759;
  assign n1761 = ~n1588 & ~n1760;
  assign n1762 = n1588 & n1760;
  assign n1763 = ~n1761 & ~n1762;
  assign n1764 = ~n1758 & ~n1763;
  assign n1765 = ~n1757 & ~n1764;
  assign n1766 = po62  & ~n1765;
  assign n1767 = ~po62  & n1765;
  assign n1768 = ~n1591 & ~n1592;
  assign n1769 = po46  & n1768;
  assign n1770 = ~n1597 & ~n1769;
  assign n1771 = n1597 & n1769;
  assign n1772 = ~n1770 & ~n1771;
  assign n1773 = ~n1767 & ~n1772;
  assign n1774 = ~n1766 & ~n1773;
  assign n1775 = n1664 & n1774;
  assign n1776 = ~n1664 & ~n1774;
  assign n1777 = n1610 & po46 ;
  assign n1778 = ~n1609 & ~n1777;
  assign n1779 = n1776 & n1778;
  assign n1780 = ~po63  & ~n1779;
  assign n1781 = ~n1489 & po46 ;
  assign n1782 = n1608 & ~n1781;
  assign n1783 = po63  & ~n1610;
  assign n1784 = ~n1782 & n1783;
  assign n1785 = ~n1775 & ~n1784;
  assign n1786 = ~n1780 & n1785;
  assign po45  = n1659 | ~n1786;
  assign n1788 = ~n1657 & ~n1658;
  assign n1789 = po45  & n1788;
  assign n1790 = ~n1626 & ~n1789;
  assign n1791 = n1626 & n1789;
  assign n1792 = ~n1790 & ~n1791;
  assign n1793 = pi90  & po45 ;
  assign n1794 = ~pi88  & ~pi89 ;
  assign n1795 = ~pi90  & n1794;
  assign n1796 = ~n1793 & ~n1795;
  assign n1797 = po46  & ~n1796;
  assign n1798 = ~po46  & n1796;
  assign n1799 = ~pi90  & po45 ;
  assign n1800 = pi91  & ~n1799;
  assign n1801 = ~pi91  & n1799;
  assign n1802 = ~n1800 & ~n1801;
  assign n1803 = ~n1798 & n1802;
  assign n1804 = ~n1797 & ~n1803;
  assign n1805 = po47  & ~n1804;
  assign n1806 = ~po47  & n1804;
  assign n1807 = po46  & n1786;
  assign n1808 = ~n1801 & ~n1807;
  assign n1809 = pi92  & ~n1808;
  assign n1810 = ~pi92  & n1808;
  assign n1811 = ~n1809 & ~n1810;
  assign n1812 = ~n1806 & ~n1811;
  assign n1813 = ~n1805 & ~n1812;
  assign n1814 = po48  & ~n1813;
  assign n1815 = ~po48  & n1813;
  assign n1816 = ~n1631 & ~n1632;
  assign n1817 = po45  & n1816;
  assign n1818 = n1636 & ~n1817;
  assign n1819 = ~n1636 & n1817;
  assign n1820 = ~n1818 & ~n1819;
  assign n1821 = ~n1815 & ~n1820;
  assign n1822 = ~n1814 & ~n1821;
  assign n1823 = po49  & ~n1822;
  assign n1824 = ~po49  & n1822;
  assign n1825 = ~n1639 & ~n1640;
  assign n1826 = po45  & n1825;
  assign n1827 = ~n1645 & ~n1826;
  assign n1828 = n1645 & n1826;
  assign n1829 = ~n1827 & ~n1828;
  assign n1830 = ~n1824 & ~n1829;
  assign n1831 = ~n1823 & ~n1830;
  assign n1832 = po50  & ~n1831;
  assign n1833 = ~po50  & n1831;
  assign n1834 = ~n1648 & ~n1649;
  assign n1835 = po45  & n1834;
  assign n1836 = n1654 & n1835;
  assign n1837 = ~n1654 & ~n1835;
  assign n1838 = ~n1836 & ~n1837;
  assign n1839 = ~n1833 & ~n1838;
  assign n1840 = ~n1832 & ~n1839;
  assign n1841 = po51  & ~n1840;
  assign n1842 = ~po51  & n1840;
  assign n1843 = n1664 & ~po45 ;
  assign n1844 = ~n1766 & ~n1767;
  assign n1845 = po45  & n1844;
  assign n1846 = ~n1772 & ~n1845;
  assign n1847 = n1772 & n1845;
  assign n1848 = ~n1846 & ~n1847;
  assign n1849 = ~n1792 & ~n1842;
  assign n1850 = ~n1841 & ~n1849;
  assign n1851 = po52  & ~n1850;
  assign n1852 = ~po52  & n1850;
  assign n1853 = ~n1667 & ~n1668;
  assign n1854 = po45  & n1853;
  assign n1855 = ~n1673 & ~n1854;
  assign n1856 = n1673 & n1854;
  assign n1857 = ~n1855 & ~n1856;
  assign n1858 = ~n1852 & ~n1857;
  assign n1859 = ~n1851 & ~n1858;
  assign n1860 = po53  & ~n1859;
  assign n1861 = ~po53  & n1859;
  assign n1862 = ~n1676 & ~n1677;
  assign n1863 = po45  & n1862;
  assign n1864 = ~n1682 & ~n1863;
  assign n1865 = n1682 & n1863;
  assign n1866 = ~n1864 & ~n1865;
  assign n1867 = ~n1861 & ~n1866;
  assign n1868 = ~n1860 & ~n1867;
  assign n1869 = po54  & ~n1868;
  assign n1870 = ~po54  & n1868;
  assign n1871 = ~n1685 & ~n1686;
  assign n1872 = po45  & n1871;
  assign n1873 = ~n1691 & ~n1872;
  assign n1874 = n1691 & n1872;
  assign n1875 = ~n1873 & ~n1874;
  assign n1876 = ~n1870 & ~n1875;
  assign n1877 = ~n1869 & ~n1876;
  assign n1878 = po55  & ~n1877;
  assign n1879 = ~po55  & n1877;
  assign n1880 = ~n1694 & ~n1695;
  assign n1881 = po45  & n1880;
  assign n1882 = ~n1700 & ~n1881;
  assign n1883 = n1700 & n1881;
  assign n1884 = ~n1882 & ~n1883;
  assign n1885 = ~n1879 & ~n1884;
  assign n1886 = ~n1878 & ~n1885;
  assign n1887 = po56  & ~n1886;
  assign n1888 = ~po56  & n1886;
  assign n1889 = ~n1703 & ~n1704;
  assign n1890 = po45  & n1889;
  assign n1891 = ~n1709 & ~n1890;
  assign n1892 = n1709 & n1890;
  assign n1893 = ~n1891 & ~n1892;
  assign n1894 = ~n1888 & ~n1893;
  assign n1895 = ~n1887 & ~n1894;
  assign n1896 = po57  & ~n1895;
  assign n1897 = ~po57  & n1895;
  assign n1898 = ~n1712 & ~n1713;
  assign n1899 = po45  & n1898;
  assign n1900 = ~n1718 & ~n1899;
  assign n1901 = n1718 & n1899;
  assign n1902 = ~n1900 & ~n1901;
  assign n1903 = ~n1897 & ~n1902;
  assign n1904 = ~n1896 & ~n1903;
  assign n1905 = po58  & ~n1904;
  assign n1906 = ~po58  & n1904;
  assign n1907 = ~n1721 & ~n1722;
  assign n1908 = po45  & n1907;
  assign n1909 = ~n1727 & ~n1908;
  assign n1910 = n1727 & n1908;
  assign n1911 = ~n1909 & ~n1910;
  assign n1912 = ~n1906 & ~n1911;
  assign n1913 = ~n1905 & ~n1912;
  assign n1914 = po59  & ~n1913;
  assign n1915 = ~po59  & n1913;
  assign n1916 = ~n1730 & ~n1731;
  assign n1917 = po45  & n1916;
  assign n1918 = ~n1736 & ~n1917;
  assign n1919 = n1736 & n1917;
  assign n1920 = ~n1918 & ~n1919;
  assign n1921 = ~n1915 & ~n1920;
  assign n1922 = ~n1914 & ~n1921;
  assign n1923 = po60  & ~n1922;
  assign n1924 = ~po60  & n1922;
  assign n1925 = ~n1739 & ~n1740;
  assign n1926 = po45  & n1925;
  assign n1927 = ~n1745 & ~n1926;
  assign n1928 = n1745 & n1926;
  assign n1929 = ~n1927 & ~n1928;
  assign n1930 = ~n1924 & ~n1929;
  assign n1931 = ~n1923 & ~n1930;
  assign n1932 = po61  & ~n1931;
  assign n1933 = ~po61  & n1931;
  assign n1934 = ~n1748 & ~n1749;
  assign n1935 = po45  & n1934;
  assign n1936 = ~n1754 & ~n1935;
  assign n1937 = n1754 & n1935;
  assign n1938 = ~n1936 & ~n1937;
  assign n1939 = ~n1933 & ~n1938;
  assign n1940 = ~n1932 & ~n1939;
  assign n1941 = po62  & ~n1940;
  assign n1942 = ~po62  & n1940;
  assign n1943 = ~n1757 & ~n1758;
  assign n1944 = po45  & n1943;
  assign n1945 = ~n1763 & ~n1944;
  assign n1946 = n1763 & n1944;
  assign n1947 = ~n1945 & ~n1946;
  assign n1948 = ~n1942 & ~n1947;
  assign n1949 = ~n1941 & ~n1948;
  assign n1950 = n1848 & n1949;
  assign n1951 = ~n1848 & ~n1949;
  assign n1952 = n1776 & po45 ;
  assign n1953 = ~n1775 & ~n1952;
  assign n1954 = n1951 & n1953;
  assign n1955 = ~po63  & ~n1954;
  assign n1956 = ~n1664 & po45 ;
  assign n1957 = n1774 & ~n1956;
  assign n1958 = po63  & ~n1776;
  assign n1959 = ~n1957 & n1958;
  assign n1960 = ~n1950 & ~n1959;
  assign n1961 = ~n1955 & n1960;
  assign po44  = n1843 | ~n1961;
  assign n1963 = ~n1841 & ~n1842;
  assign n1964 = po44  & n1963;
  assign n1965 = ~n1792 & ~n1964;
  assign n1966 = n1792 & n1964;
  assign n1967 = ~n1965 & ~n1966;
  assign n1968 = pi88  & po44 ;
  assign n1969 = ~pi86  & ~pi87 ;
  assign n1970 = ~pi88  & n1969;
  assign n1971 = ~n1968 & ~n1970;
  assign n1972 = po45  & ~n1971;
  assign n1973 = ~po45  & n1971;
  assign n1974 = ~pi88  & po44 ;
  assign n1975 = pi89  & ~n1974;
  assign n1976 = ~pi89  & n1974;
  assign n1977 = ~n1975 & ~n1976;
  assign n1978 = ~n1973 & n1977;
  assign n1979 = ~n1972 & ~n1978;
  assign n1980 = po46  & ~n1979;
  assign n1981 = ~po46  & n1979;
  assign n1982 = po45  & n1961;
  assign n1983 = ~n1976 & ~n1982;
  assign n1984 = pi90  & ~n1983;
  assign n1985 = ~pi90  & n1983;
  assign n1986 = ~n1984 & ~n1985;
  assign n1987 = ~n1981 & ~n1986;
  assign n1988 = ~n1980 & ~n1987;
  assign n1989 = po47  & ~n1988;
  assign n1990 = ~po47  & n1988;
  assign n1991 = ~n1797 & ~n1798;
  assign n1992 = po44  & n1991;
  assign n1993 = n1802 & ~n1992;
  assign n1994 = ~n1802 & n1992;
  assign n1995 = ~n1993 & ~n1994;
  assign n1996 = ~n1990 & ~n1995;
  assign n1997 = ~n1989 & ~n1996;
  assign n1998 = po48  & ~n1997;
  assign n1999 = ~po48  & n1997;
  assign n2000 = ~n1805 & ~n1806;
  assign n2001 = po44  & n2000;
  assign n2002 = ~n1811 & ~n2001;
  assign n2003 = n1811 & n2001;
  assign n2004 = ~n2002 & ~n2003;
  assign n2005 = ~n1999 & ~n2004;
  assign n2006 = ~n1998 & ~n2005;
  assign n2007 = po49  & ~n2006;
  assign n2008 = ~po49  & n2006;
  assign n2009 = ~n1814 & ~n1815;
  assign n2010 = po44  & n2009;
  assign n2011 = n1820 & n2010;
  assign n2012 = ~n1820 & ~n2010;
  assign n2013 = ~n2011 & ~n2012;
  assign n2014 = ~n2008 & ~n2013;
  assign n2015 = ~n2007 & ~n2014;
  assign n2016 = po50  & ~n2015;
  assign n2017 = ~po50  & n2015;
  assign n2018 = ~n1823 & ~n1824;
  assign n2019 = po44  & n2018;
  assign n2020 = ~n1829 & ~n2019;
  assign n2021 = n1829 & n2019;
  assign n2022 = ~n2020 & ~n2021;
  assign n2023 = ~n2017 & ~n2022;
  assign n2024 = ~n2016 & ~n2023;
  assign n2025 = po51  & ~n2024;
  assign n2026 = ~po51  & n2024;
  assign n2027 = ~n1832 & ~n1833;
  assign n2028 = po44  & n2027;
  assign n2029 = ~n1838 & ~n2028;
  assign n2030 = n1838 & n2028;
  assign n2031 = ~n2029 & ~n2030;
  assign n2032 = ~n2026 & ~n2031;
  assign n2033 = ~n2025 & ~n2032;
  assign n2034 = po52  & ~n2033;
  assign n2035 = ~po52  & n2033;
  assign n2036 = n1848 & ~po44 ;
  assign n2037 = ~n1941 & ~n1942;
  assign n2038 = po44  & n2037;
  assign n2039 = ~n1947 & ~n2038;
  assign n2040 = n1947 & n2038;
  assign n2041 = ~n2039 & ~n2040;
  assign n2042 = ~n1967 & ~n2035;
  assign n2043 = ~n2034 & ~n2042;
  assign n2044 = po53  & ~n2043;
  assign n2045 = ~po53  & n2043;
  assign n2046 = ~n1851 & ~n1852;
  assign n2047 = po44  & n2046;
  assign n2048 = ~n1857 & ~n2047;
  assign n2049 = n1857 & n2047;
  assign n2050 = ~n2048 & ~n2049;
  assign n2051 = ~n2045 & ~n2050;
  assign n2052 = ~n2044 & ~n2051;
  assign n2053 = po54  & ~n2052;
  assign n2054 = ~po54  & n2052;
  assign n2055 = ~n1860 & ~n1861;
  assign n2056 = po44  & n2055;
  assign n2057 = ~n1866 & ~n2056;
  assign n2058 = n1866 & n2056;
  assign n2059 = ~n2057 & ~n2058;
  assign n2060 = ~n2054 & ~n2059;
  assign n2061 = ~n2053 & ~n2060;
  assign n2062 = po55  & ~n2061;
  assign n2063 = ~po55  & n2061;
  assign n2064 = ~n1869 & ~n1870;
  assign n2065 = po44  & n2064;
  assign n2066 = ~n1875 & ~n2065;
  assign n2067 = n1875 & n2065;
  assign n2068 = ~n2066 & ~n2067;
  assign n2069 = ~n2063 & ~n2068;
  assign n2070 = ~n2062 & ~n2069;
  assign n2071 = po56  & ~n2070;
  assign n2072 = ~po56  & n2070;
  assign n2073 = ~n1878 & ~n1879;
  assign n2074 = po44  & n2073;
  assign n2075 = ~n1884 & ~n2074;
  assign n2076 = n1884 & n2074;
  assign n2077 = ~n2075 & ~n2076;
  assign n2078 = ~n2072 & ~n2077;
  assign n2079 = ~n2071 & ~n2078;
  assign n2080 = po57  & ~n2079;
  assign n2081 = ~po57  & n2079;
  assign n2082 = ~n1887 & ~n1888;
  assign n2083 = po44  & n2082;
  assign n2084 = ~n1893 & ~n2083;
  assign n2085 = n1893 & n2083;
  assign n2086 = ~n2084 & ~n2085;
  assign n2087 = ~n2081 & ~n2086;
  assign n2088 = ~n2080 & ~n2087;
  assign n2089 = po58  & ~n2088;
  assign n2090 = ~po58  & n2088;
  assign n2091 = ~n1896 & ~n1897;
  assign n2092 = po44  & n2091;
  assign n2093 = ~n1902 & ~n2092;
  assign n2094 = n1902 & n2092;
  assign n2095 = ~n2093 & ~n2094;
  assign n2096 = ~n2090 & ~n2095;
  assign n2097 = ~n2089 & ~n2096;
  assign n2098 = po59  & ~n2097;
  assign n2099 = ~po59  & n2097;
  assign n2100 = ~n1905 & ~n1906;
  assign n2101 = po44  & n2100;
  assign n2102 = ~n1911 & ~n2101;
  assign n2103 = n1911 & n2101;
  assign n2104 = ~n2102 & ~n2103;
  assign n2105 = ~n2099 & ~n2104;
  assign n2106 = ~n2098 & ~n2105;
  assign n2107 = po60  & ~n2106;
  assign n2108 = ~po60  & n2106;
  assign n2109 = ~n1914 & ~n1915;
  assign n2110 = po44  & n2109;
  assign n2111 = ~n1920 & ~n2110;
  assign n2112 = n1920 & n2110;
  assign n2113 = ~n2111 & ~n2112;
  assign n2114 = ~n2108 & ~n2113;
  assign n2115 = ~n2107 & ~n2114;
  assign n2116 = po61  & ~n2115;
  assign n2117 = ~po61  & n2115;
  assign n2118 = ~n1923 & ~n1924;
  assign n2119 = po44  & n2118;
  assign n2120 = ~n1929 & ~n2119;
  assign n2121 = n1929 & n2119;
  assign n2122 = ~n2120 & ~n2121;
  assign n2123 = ~n2117 & ~n2122;
  assign n2124 = ~n2116 & ~n2123;
  assign n2125 = po62  & ~n2124;
  assign n2126 = ~po62  & n2124;
  assign n2127 = ~n1932 & ~n1933;
  assign n2128 = po44  & n2127;
  assign n2129 = ~n1938 & ~n2128;
  assign n2130 = n1938 & n2128;
  assign n2131 = ~n2129 & ~n2130;
  assign n2132 = ~n2126 & ~n2131;
  assign n2133 = ~n2125 & ~n2132;
  assign n2134 = n2041 & n2133;
  assign n2135 = ~n2041 & ~n2133;
  assign n2136 = n1951 & po44 ;
  assign n2137 = ~n1950 & ~n2136;
  assign n2138 = n2135 & n2137;
  assign n2139 = ~po63  & ~n2138;
  assign n2140 = ~n1848 & po44 ;
  assign n2141 = n1949 & ~n2140;
  assign n2142 = po63  & ~n1951;
  assign n2143 = ~n2141 & n2142;
  assign n2144 = ~n2134 & ~n2143;
  assign n2145 = ~n2139 & n2144;
  assign po43  = n2036 | ~n2145;
  assign n2147 = ~n2034 & ~n2035;
  assign n2148 = po43  & n2147;
  assign n2149 = ~n1967 & ~n2148;
  assign n2150 = n1967 & n2148;
  assign n2151 = ~n2149 & ~n2150;
  assign n2152 = pi86  & po43 ;
  assign n2153 = ~pi84  & ~pi85 ;
  assign n2154 = ~pi86  & n2153;
  assign n2155 = ~n2152 & ~n2154;
  assign n2156 = po44  & ~n2155;
  assign n2157 = ~po44  & n2155;
  assign n2158 = ~pi86  & po43 ;
  assign n2159 = pi87  & ~n2158;
  assign n2160 = ~pi87  & n2158;
  assign n2161 = ~n2159 & ~n2160;
  assign n2162 = ~n2157 & n2161;
  assign n2163 = ~n2156 & ~n2162;
  assign n2164 = po45  & ~n2163;
  assign n2165 = ~po45  & n2163;
  assign n2166 = po44  & n2145;
  assign n2167 = ~n2160 & ~n2166;
  assign n2168 = pi88  & ~n2167;
  assign n2169 = ~pi88  & n2167;
  assign n2170 = ~n2168 & ~n2169;
  assign n2171 = ~n2165 & ~n2170;
  assign n2172 = ~n2164 & ~n2171;
  assign n2173 = po46  & ~n2172;
  assign n2174 = ~po46  & n2172;
  assign n2175 = ~n1972 & ~n1973;
  assign n2176 = po43  & n2175;
  assign n2177 = n1977 & ~n2176;
  assign n2178 = ~n1977 & n2176;
  assign n2179 = ~n2177 & ~n2178;
  assign n2180 = ~n2174 & ~n2179;
  assign n2181 = ~n2173 & ~n2180;
  assign n2182 = po47  & ~n2181;
  assign n2183 = ~po47  & n2181;
  assign n2184 = ~n1980 & ~n1981;
  assign n2185 = po43  & n2184;
  assign n2186 = ~n1986 & ~n2185;
  assign n2187 = n1986 & n2185;
  assign n2188 = ~n2186 & ~n2187;
  assign n2189 = ~n2183 & ~n2188;
  assign n2190 = ~n2182 & ~n2189;
  assign n2191 = po48  & ~n2190;
  assign n2192 = ~po48  & n2190;
  assign n2193 = ~n1989 & ~n1990;
  assign n2194 = po43  & n2193;
  assign n2195 = n1995 & n2194;
  assign n2196 = ~n1995 & ~n2194;
  assign n2197 = ~n2195 & ~n2196;
  assign n2198 = ~n2192 & ~n2197;
  assign n2199 = ~n2191 & ~n2198;
  assign n2200 = po49  & ~n2199;
  assign n2201 = ~po49  & n2199;
  assign n2202 = ~n1998 & ~n1999;
  assign n2203 = po43  & n2202;
  assign n2204 = ~n2004 & ~n2203;
  assign n2205 = n2004 & n2203;
  assign n2206 = ~n2204 & ~n2205;
  assign n2207 = ~n2201 & ~n2206;
  assign n2208 = ~n2200 & ~n2207;
  assign n2209 = po50  & ~n2208;
  assign n2210 = ~po50  & n2208;
  assign n2211 = ~n2007 & ~n2008;
  assign n2212 = po43  & n2211;
  assign n2213 = ~n2013 & ~n2212;
  assign n2214 = n2013 & n2212;
  assign n2215 = ~n2213 & ~n2214;
  assign n2216 = ~n2210 & ~n2215;
  assign n2217 = ~n2209 & ~n2216;
  assign n2218 = po51  & ~n2217;
  assign n2219 = ~po51  & n2217;
  assign n2220 = ~n2016 & ~n2017;
  assign n2221 = po43  & n2220;
  assign n2222 = ~n2022 & ~n2221;
  assign n2223 = n2022 & n2221;
  assign n2224 = ~n2222 & ~n2223;
  assign n2225 = ~n2219 & ~n2224;
  assign n2226 = ~n2218 & ~n2225;
  assign n2227 = po52  & ~n2226;
  assign n2228 = ~po52  & n2226;
  assign n2229 = ~n2025 & ~n2026;
  assign n2230 = po43  & n2229;
  assign n2231 = ~n2031 & ~n2230;
  assign n2232 = n2031 & n2230;
  assign n2233 = ~n2231 & ~n2232;
  assign n2234 = ~n2228 & ~n2233;
  assign n2235 = ~n2227 & ~n2234;
  assign n2236 = po53  & ~n2235;
  assign n2237 = ~po53  & n2235;
  assign n2238 = n2041 & ~po43 ;
  assign n2239 = ~n2125 & ~n2126;
  assign n2240 = po43  & n2239;
  assign n2241 = ~n2131 & ~n2240;
  assign n2242 = n2131 & n2240;
  assign n2243 = ~n2241 & ~n2242;
  assign n2244 = ~n2151 & ~n2237;
  assign n2245 = ~n2236 & ~n2244;
  assign n2246 = po54  & ~n2245;
  assign n2247 = ~po54  & n2245;
  assign n2248 = ~n2044 & ~n2045;
  assign n2249 = po43  & n2248;
  assign n2250 = ~n2050 & ~n2249;
  assign n2251 = n2050 & n2249;
  assign n2252 = ~n2250 & ~n2251;
  assign n2253 = ~n2247 & ~n2252;
  assign n2254 = ~n2246 & ~n2253;
  assign n2255 = po55  & ~n2254;
  assign n2256 = ~po55  & n2254;
  assign n2257 = ~n2053 & ~n2054;
  assign n2258 = po43  & n2257;
  assign n2259 = ~n2059 & ~n2258;
  assign n2260 = n2059 & n2258;
  assign n2261 = ~n2259 & ~n2260;
  assign n2262 = ~n2256 & ~n2261;
  assign n2263 = ~n2255 & ~n2262;
  assign n2264 = po56  & ~n2263;
  assign n2265 = ~po56  & n2263;
  assign n2266 = ~n2062 & ~n2063;
  assign n2267 = po43  & n2266;
  assign n2268 = ~n2068 & ~n2267;
  assign n2269 = n2068 & n2267;
  assign n2270 = ~n2268 & ~n2269;
  assign n2271 = ~n2265 & ~n2270;
  assign n2272 = ~n2264 & ~n2271;
  assign n2273 = po57  & ~n2272;
  assign n2274 = ~po57  & n2272;
  assign n2275 = ~n2071 & ~n2072;
  assign n2276 = po43  & n2275;
  assign n2277 = ~n2077 & ~n2276;
  assign n2278 = n2077 & n2276;
  assign n2279 = ~n2277 & ~n2278;
  assign n2280 = ~n2274 & ~n2279;
  assign n2281 = ~n2273 & ~n2280;
  assign n2282 = po58  & ~n2281;
  assign n2283 = ~po58  & n2281;
  assign n2284 = ~n2080 & ~n2081;
  assign n2285 = po43  & n2284;
  assign n2286 = ~n2086 & ~n2285;
  assign n2287 = n2086 & n2285;
  assign n2288 = ~n2286 & ~n2287;
  assign n2289 = ~n2283 & ~n2288;
  assign n2290 = ~n2282 & ~n2289;
  assign n2291 = po59  & ~n2290;
  assign n2292 = ~po59  & n2290;
  assign n2293 = ~n2089 & ~n2090;
  assign n2294 = po43  & n2293;
  assign n2295 = ~n2095 & ~n2294;
  assign n2296 = n2095 & n2294;
  assign n2297 = ~n2295 & ~n2296;
  assign n2298 = ~n2292 & ~n2297;
  assign n2299 = ~n2291 & ~n2298;
  assign n2300 = po60  & ~n2299;
  assign n2301 = ~po60  & n2299;
  assign n2302 = ~n2098 & ~n2099;
  assign n2303 = po43  & n2302;
  assign n2304 = ~n2104 & ~n2303;
  assign n2305 = n2104 & n2303;
  assign n2306 = ~n2304 & ~n2305;
  assign n2307 = ~n2301 & ~n2306;
  assign n2308 = ~n2300 & ~n2307;
  assign n2309 = po61  & ~n2308;
  assign n2310 = ~po61  & n2308;
  assign n2311 = ~n2107 & ~n2108;
  assign n2312 = po43  & n2311;
  assign n2313 = ~n2113 & ~n2312;
  assign n2314 = n2113 & n2312;
  assign n2315 = ~n2313 & ~n2314;
  assign n2316 = ~n2310 & ~n2315;
  assign n2317 = ~n2309 & ~n2316;
  assign n2318 = po62  & ~n2317;
  assign n2319 = ~po62  & n2317;
  assign n2320 = ~n2116 & ~n2117;
  assign n2321 = po43  & n2320;
  assign n2322 = ~n2122 & ~n2321;
  assign n2323 = n2122 & n2321;
  assign n2324 = ~n2322 & ~n2323;
  assign n2325 = ~n2319 & ~n2324;
  assign n2326 = ~n2318 & ~n2325;
  assign n2327 = n2243 & n2326;
  assign n2328 = ~n2243 & ~n2326;
  assign n2329 = n2135 & po43 ;
  assign n2330 = ~n2134 & ~n2329;
  assign n2331 = n2328 & n2330;
  assign n2332 = ~po63  & ~n2331;
  assign n2333 = ~n2041 & po43 ;
  assign n2334 = n2133 & ~n2333;
  assign n2335 = po63  & ~n2135;
  assign n2336 = ~n2334 & n2335;
  assign n2337 = ~n2327 & ~n2336;
  assign n2338 = ~n2332 & n2337;
  assign po42  = n2238 | ~n2338;
  assign n2340 = ~n2236 & ~n2237;
  assign n2341 = po42  & n2340;
  assign n2342 = ~n2151 & ~n2341;
  assign n2343 = n2151 & n2341;
  assign n2344 = ~n2342 & ~n2343;
  assign n2345 = pi84  & po42 ;
  assign n2346 = ~pi82  & ~pi83 ;
  assign n2347 = ~pi84  & n2346;
  assign n2348 = ~n2345 & ~n2347;
  assign n2349 = po43  & ~n2348;
  assign n2350 = ~po43  & n2348;
  assign n2351 = ~pi84  & po42 ;
  assign n2352 = pi85  & ~n2351;
  assign n2353 = ~pi85  & n2351;
  assign n2354 = ~n2352 & ~n2353;
  assign n2355 = ~n2350 & n2354;
  assign n2356 = ~n2349 & ~n2355;
  assign n2357 = po44  & ~n2356;
  assign n2358 = ~po44  & n2356;
  assign n2359 = po43  & n2338;
  assign n2360 = ~n2353 & ~n2359;
  assign n2361 = pi86  & ~n2360;
  assign n2362 = ~pi86  & n2360;
  assign n2363 = ~n2361 & ~n2362;
  assign n2364 = ~n2358 & ~n2363;
  assign n2365 = ~n2357 & ~n2364;
  assign n2366 = po45  & ~n2365;
  assign n2367 = ~po45  & n2365;
  assign n2368 = ~n2156 & ~n2157;
  assign n2369 = po42  & n2368;
  assign n2370 = n2161 & ~n2369;
  assign n2371 = ~n2161 & n2369;
  assign n2372 = ~n2370 & ~n2371;
  assign n2373 = ~n2367 & ~n2372;
  assign n2374 = ~n2366 & ~n2373;
  assign n2375 = po46  & ~n2374;
  assign n2376 = ~po46  & n2374;
  assign n2377 = ~n2164 & ~n2165;
  assign n2378 = po42  & n2377;
  assign n2379 = ~n2170 & ~n2378;
  assign n2380 = n2170 & n2378;
  assign n2381 = ~n2379 & ~n2380;
  assign n2382 = ~n2376 & ~n2381;
  assign n2383 = ~n2375 & ~n2382;
  assign n2384 = po47  & ~n2383;
  assign n2385 = ~po47  & n2383;
  assign n2386 = ~n2173 & ~n2174;
  assign n2387 = po42  & n2386;
  assign n2388 = n2179 & n2387;
  assign n2389 = ~n2179 & ~n2387;
  assign n2390 = ~n2388 & ~n2389;
  assign n2391 = ~n2385 & ~n2390;
  assign n2392 = ~n2384 & ~n2391;
  assign n2393 = po48  & ~n2392;
  assign n2394 = ~po48  & n2392;
  assign n2395 = ~n2182 & ~n2183;
  assign n2396 = po42  & n2395;
  assign n2397 = ~n2188 & ~n2396;
  assign n2398 = n2188 & n2396;
  assign n2399 = ~n2397 & ~n2398;
  assign n2400 = ~n2394 & ~n2399;
  assign n2401 = ~n2393 & ~n2400;
  assign n2402 = po49  & ~n2401;
  assign n2403 = ~po49  & n2401;
  assign n2404 = ~n2191 & ~n2192;
  assign n2405 = po42  & n2404;
  assign n2406 = ~n2197 & ~n2405;
  assign n2407 = n2197 & n2405;
  assign n2408 = ~n2406 & ~n2407;
  assign n2409 = ~n2403 & ~n2408;
  assign n2410 = ~n2402 & ~n2409;
  assign n2411 = po50  & ~n2410;
  assign n2412 = ~po50  & n2410;
  assign n2413 = ~n2200 & ~n2201;
  assign n2414 = po42  & n2413;
  assign n2415 = ~n2206 & ~n2414;
  assign n2416 = n2206 & n2414;
  assign n2417 = ~n2415 & ~n2416;
  assign n2418 = ~n2412 & ~n2417;
  assign n2419 = ~n2411 & ~n2418;
  assign n2420 = po51  & ~n2419;
  assign n2421 = ~po51  & n2419;
  assign n2422 = ~n2209 & ~n2210;
  assign n2423 = po42  & n2422;
  assign n2424 = ~n2215 & ~n2423;
  assign n2425 = n2215 & n2423;
  assign n2426 = ~n2424 & ~n2425;
  assign n2427 = ~n2421 & ~n2426;
  assign n2428 = ~n2420 & ~n2427;
  assign n2429 = po52  & ~n2428;
  assign n2430 = ~po52  & n2428;
  assign n2431 = ~n2218 & ~n2219;
  assign n2432 = po42  & n2431;
  assign n2433 = ~n2224 & ~n2432;
  assign n2434 = n2224 & n2432;
  assign n2435 = ~n2433 & ~n2434;
  assign n2436 = ~n2430 & ~n2435;
  assign n2437 = ~n2429 & ~n2436;
  assign n2438 = po53  & ~n2437;
  assign n2439 = ~po53  & n2437;
  assign n2440 = ~n2227 & ~n2228;
  assign n2441 = po42  & n2440;
  assign n2442 = ~n2233 & ~n2441;
  assign n2443 = n2233 & n2441;
  assign n2444 = ~n2442 & ~n2443;
  assign n2445 = ~n2439 & ~n2444;
  assign n2446 = ~n2438 & ~n2445;
  assign n2447 = po54  & ~n2446;
  assign n2448 = ~po54  & n2446;
  assign n2449 = n2243 & ~po42 ;
  assign n2450 = ~n2318 & ~n2319;
  assign n2451 = po42  & n2450;
  assign n2452 = ~n2324 & ~n2451;
  assign n2453 = n2324 & n2451;
  assign n2454 = ~n2452 & ~n2453;
  assign n2455 = ~n2344 & ~n2448;
  assign n2456 = ~n2447 & ~n2455;
  assign n2457 = po55  & ~n2456;
  assign n2458 = ~po55  & n2456;
  assign n2459 = ~n2246 & ~n2247;
  assign n2460 = po42  & n2459;
  assign n2461 = ~n2252 & ~n2460;
  assign n2462 = n2252 & n2460;
  assign n2463 = ~n2461 & ~n2462;
  assign n2464 = ~n2458 & ~n2463;
  assign n2465 = ~n2457 & ~n2464;
  assign n2466 = po56  & ~n2465;
  assign n2467 = ~po56  & n2465;
  assign n2468 = ~n2255 & ~n2256;
  assign n2469 = po42  & n2468;
  assign n2470 = ~n2261 & ~n2469;
  assign n2471 = n2261 & n2469;
  assign n2472 = ~n2470 & ~n2471;
  assign n2473 = ~n2467 & ~n2472;
  assign n2474 = ~n2466 & ~n2473;
  assign n2475 = po57  & ~n2474;
  assign n2476 = ~po57  & n2474;
  assign n2477 = ~n2264 & ~n2265;
  assign n2478 = po42  & n2477;
  assign n2479 = ~n2270 & ~n2478;
  assign n2480 = n2270 & n2478;
  assign n2481 = ~n2479 & ~n2480;
  assign n2482 = ~n2476 & ~n2481;
  assign n2483 = ~n2475 & ~n2482;
  assign n2484 = po58  & ~n2483;
  assign n2485 = ~po58  & n2483;
  assign n2486 = ~n2273 & ~n2274;
  assign n2487 = po42  & n2486;
  assign n2488 = ~n2279 & ~n2487;
  assign n2489 = n2279 & n2487;
  assign n2490 = ~n2488 & ~n2489;
  assign n2491 = ~n2485 & ~n2490;
  assign n2492 = ~n2484 & ~n2491;
  assign n2493 = po59  & ~n2492;
  assign n2494 = ~po59  & n2492;
  assign n2495 = ~n2282 & ~n2283;
  assign n2496 = po42  & n2495;
  assign n2497 = ~n2288 & ~n2496;
  assign n2498 = n2288 & n2496;
  assign n2499 = ~n2497 & ~n2498;
  assign n2500 = ~n2494 & ~n2499;
  assign n2501 = ~n2493 & ~n2500;
  assign n2502 = po60  & ~n2501;
  assign n2503 = ~po60  & n2501;
  assign n2504 = ~n2291 & ~n2292;
  assign n2505 = po42  & n2504;
  assign n2506 = ~n2297 & ~n2505;
  assign n2507 = n2297 & n2505;
  assign n2508 = ~n2506 & ~n2507;
  assign n2509 = ~n2503 & ~n2508;
  assign n2510 = ~n2502 & ~n2509;
  assign n2511 = po61  & ~n2510;
  assign n2512 = ~po61  & n2510;
  assign n2513 = ~n2300 & ~n2301;
  assign n2514 = po42  & n2513;
  assign n2515 = ~n2306 & ~n2514;
  assign n2516 = n2306 & n2514;
  assign n2517 = ~n2515 & ~n2516;
  assign n2518 = ~n2512 & ~n2517;
  assign n2519 = ~n2511 & ~n2518;
  assign n2520 = po62  & ~n2519;
  assign n2521 = ~po62  & n2519;
  assign n2522 = ~n2309 & ~n2310;
  assign n2523 = po42  & n2522;
  assign n2524 = ~n2315 & ~n2523;
  assign n2525 = n2315 & n2523;
  assign n2526 = ~n2524 & ~n2525;
  assign n2527 = ~n2521 & ~n2526;
  assign n2528 = ~n2520 & ~n2527;
  assign n2529 = n2454 & n2528;
  assign n2530 = ~n2454 & ~n2528;
  assign n2531 = n2328 & po42 ;
  assign n2532 = ~n2327 & ~n2531;
  assign n2533 = n2530 & n2532;
  assign n2534 = ~po63  & ~n2533;
  assign n2535 = ~n2243 & po42 ;
  assign n2536 = n2326 & ~n2535;
  assign n2537 = po63  & ~n2328;
  assign n2538 = ~n2536 & n2537;
  assign n2539 = ~n2529 & ~n2538;
  assign n2540 = ~n2534 & n2539;
  assign po41  = n2449 | ~n2540;
  assign n2542 = ~n2447 & ~n2448;
  assign n2543 = po41  & n2542;
  assign n2544 = ~n2344 & ~n2543;
  assign n2545 = n2344 & n2543;
  assign n2546 = ~n2544 & ~n2545;
  assign n2547 = pi82  & po41 ;
  assign n2548 = ~pi80  & ~pi81 ;
  assign n2549 = ~pi82  & n2548;
  assign n2550 = ~n2547 & ~n2549;
  assign n2551 = po42  & ~n2550;
  assign n2552 = ~po42  & n2550;
  assign n2553 = ~pi82  & po41 ;
  assign n2554 = pi83  & ~n2553;
  assign n2555 = ~pi83  & n2553;
  assign n2556 = ~n2554 & ~n2555;
  assign n2557 = ~n2552 & n2556;
  assign n2558 = ~n2551 & ~n2557;
  assign n2559 = po43  & ~n2558;
  assign n2560 = ~po43  & n2558;
  assign n2561 = po42  & n2540;
  assign n2562 = ~n2555 & ~n2561;
  assign n2563 = pi84  & ~n2562;
  assign n2564 = ~pi84  & n2562;
  assign n2565 = ~n2563 & ~n2564;
  assign n2566 = ~n2560 & ~n2565;
  assign n2567 = ~n2559 & ~n2566;
  assign n2568 = po44  & ~n2567;
  assign n2569 = ~po44  & n2567;
  assign n2570 = ~n2349 & ~n2350;
  assign n2571 = po41  & n2570;
  assign n2572 = n2354 & ~n2571;
  assign n2573 = ~n2354 & n2571;
  assign n2574 = ~n2572 & ~n2573;
  assign n2575 = ~n2569 & ~n2574;
  assign n2576 = ~n2568 & ~n2575;
  assign n2577 = po45  & ~n2576;
  assign n2578 = ~po45  & n2576;
  assign n2579 = ~n2357 & ~n2358;
  assign n2580 = po41  & n2579;
  assign n2581 = ~n2363 & ~n2580;
  assign n2582 = n2363 & n2580;
  assign n2583 = ~n2581 & ~n2582;
  assign n2584 = ~n2578 & ~n2583;
  assign n2585 = ~n2577 & ~n2584;
  assign n2586 = po46  & ~n2585;
  assign n2587 = ~po46  & n2585;
  assign n2588 = ~n2366 & ~n2367;
  assign n2589 = po41  & n2588;
  assign n2590 = n2372 & n2589;
  assign n2591 = ~n2372 & ~n2589;
  assign n2592 = ~n2590 & ~n2591;
  assign n2593 = ~n2587 & ~n2592;
  assign n2594 = ~n2586 & ~n2593;
  assign n2595 = po47  & ~n2594;
  assign n2596 = ~po47  & n2594;
  assign n2597 = ~n2375 & ~n2376;
  assign n2598 = po41  & n2597;
  assign n2599 = ~n2381 & ~n2598;
  assign n2600 = n2381 & n2598;
  assign n2601 = ~n2599 & ~n2600;
  assign n2602 = ~n2596 & ~n2601;
  assign n2603 = ~n2595 & ~n2602;
  assign n2604 = po48  & ~n2603;
  assign n2605 = ~po48  & n2603;
  assign n2606 = ~n2384 & ~n2385;
  assign n2607 = po41  & n2606;
  assign n2608 = ~n2390 & ~n2607;
  assign n2609 = n2390 & n2607;
  assign n2610 = ~n2608 & ~n2609;
  assign n2611 = ~n2605 & ~n2610;
  assign n2612 = ~n2604 & ~n2611;
  assign n2613 = po49  & ~n2612;
  assign n2614 = ~po49  & n2612;
  assign n2615 = ~n2393 & ~n2394;
  assign n2616 = po41  & n2615;
  assign n2617 = ~n2399 & ~n2616;
  assign n2618 = n2399 & n2616;
  assign n2619 = ~n2617 & ~n2618;
  assign n2620 = ~n2614 & ~n2619;
  assign n2621 = ~n2613 & ~n2620;
  assign n2622 = po50  & ~n2621;
  assign n2623 = ~po50  & n2621;
  assign n2624 = ~n2402 & ~n2403;
  assign n2625 = po41  & n2624;
  assign n2626 = ~n2408 & ~n2625;
  assign n2627 = n2408 & n2625;
  assign n2628 = ~n2626 & ~n2627;
  assign n2629 = ~n2623 & ~n2628;
  assign n2630 = ~n2622 & ~n2629;
  assign n2631 = po51  & ~n2630;
  assign n2632 = ~po51  & n2630;
  assign n2633 = ~n2411 & ~n2412;
  assign n2634 = po41  & n2633;
  assign n2635 = ~n2417 & ~n2634;
  assign n2636 = n2417 & n2634;
  assign n2637 = ~n2635 & ~n2636;
  assign n2638 = ~n2632 & ~n2637;
  assign n2639 = ~n2631 & ~n2638;
  assign n2640 = po52  & ~n2639;
  assign n2641 = ~po52  & n2639;
  assign n2642 = ~n2420 & ~n2421;
  assign n2643 = po41  & n2642;
  assign n2644 = ~n2426 & ~n2643;
  assign n2645 = n2426 & n2643;
  assign n2646 = ~n2644 & ~n2645;
  assign n2647 = ~n2641 & ~n2646;
  assign n2648 = ~n2640 & ~n2647;
  assign n2649 = po53  & ~n2648;
  assign n2650 = ~po53  & n2648;
  assign n2651 = ~n2429 & ~n2430;
  assign n2652 = po41  & n2651;
  assign n2653 = ~n2435 & ~n2652;
  assign n2654 = n2435 & n2652;
  assign n2655 = ~n2653 & ~n2654;
  assign n2656 = ~n2650 & ~n2655;
  assign n2657 = ~n2649 & ~n2656;
  assign n2658 = po54  & ~n2657;
  assign n2659 = ~po54  & n2657;
  assign n2660 = ~n2438 & ~n2439;
  assign n2661 = po41  & n2660;
  assign n2662 = ~n2444 & ~n2661;
  assign n2663 = n2444 & n2661;
  assign n2664 = ~n2662 & ~n2663;
  assign n2665 = ~n2659 & ~n2664;
  assign n2666 = ~n2658 & ~n2665;
  assign n2667 = po55  & ~n2666;
  assign n2668 = ~po55  & n2666;
  assign n2669 = n2454 & ~po41 ;
  assign n2670 = ~n2520 & ~n2521;
  assign n2671 = po41  & n2670;
  assign n2672 = ~n2526 & ~n2671;
  assign n2673 = n2526 & n2671;
  assign n2674 = ~n2672 & ~n2673;
  assign n2675 = ~n2546 & ~n2668;
  assign n2676 = ~n2667 & ~n2675;
  assign n2677 = po56  & ~n2676;
  assign n2678 = ~po56  & n2676;
  assign n2679 = ~n2457 & ~n2458;
  assign n2680 = po41  & n2679;
  assign n2681 = ~n2463 & ~n2680;
  assign n2682 = n2463 & n2680;
  assign n2683 = ~n2681 & ~n2682;
  assign n2684 = ~n2678 & ~n2683;
  assign n2685 = ~n2677 & ~n2684;
  assign n2686 = po57  & ~n2685;
  assign n2687 = ~po57  & n2685;
  assign n2688 = ~n2466 & ~n2467;
  assign n2689 = po41  & n2688;
  assign n2690 = ~n2472 & ~n2689;
  assign n2691 = n2472 & n2689;
  assign n2692 = ~n2690 & ~n2691;
  assign n2693 = ~n2687 & ~n2692;
  assign n2694 = ~n2686 & ~n2693;
  assign n2695 = po58  & ~n2694;
  assign n2696 = ~po58  & n2694;
  assign n2697 = ~n2475 & ~n2476;
  assign n2698 = po41  & n2697;
  assign n2699 = ~n2481 & ~n2698;
  assign n2700 = n2481 & n2698;
  assign n2701 = ~n2699 & ~n2700;
  assign n2702 = ~n2696 & ~n2701;
  assign n2703 = ~n2695 & ~n2702;
  assign n2704 = po59  & ~n2703;
  assign n2705 = ~po59  & n2703;
  assign n2706 = ~n2484 & ~n2485;
  assign n2707 = po41  & n2706;
  assign n2708 = ~n2490 & ~n2707;
  assign n2709 = n2490 & n2707;
  assign n2710 = ~n2708 & ~n2709;
  assign n2711 = ~n2705 & ~n2710;
  assign n2712 = ~n2704 & ~n2711;
  assign n2713 = po60  & ~n2712;
  assign n2714 = ~po60  & n2712;
  assign n2715 = ~n2493 & ~n2494;
  assign n2716 = po41  & n2715;
  assign n2717 = ~n2499 & ~n2716;
  assign n2718 = n2499 & n2716;
  assign n2719 = ~n2717 & ~n2718;
  assign n2720 = ~n2714 & ~n2719;
  assign n2721 = ~n2713 & ~n2720;
  assign n2722 = po61  & ~n2721;
  assign n2723 = ~po61  & n2721;
  assign n2724 = ~n2502 & ~n2503;
  assign n2725 = po41  & n2724;
  assign n2726 = ~n2508 & ~n2725;
  assign n2727 = n2508 & n2725;
  assign n2728 = ~n2726 & ~n2727;
  assign n2729 = ~n2723 & ~n2728;
  assign n2730 = ~n2722 & ~n2729;
  assign n2731 = po62  & ~n2730;
  assign n2732 = ~po62  & n2730;
  assign n2733 = ~n2511 & ~n2512;
  assign n2734 = po41  & n2733;
  assign n2735 = ~n2517 & ~n2734;
  assign n2736 = n2517 & n2734;
  assign n2737 = ~n2735 & ~n2736;
  assign n2738 = ~n2732 & ~n2737;
  assign n2739 = ~n2731 & ~n2738;
  assign n2740 = n2674 & n2739;
  assign n2741 = ~n2674 & ~n2739;
  assign n2742 = n2530 & po41 ;
  assign n2743 = ~n2529 & ~n2742;
  assign n2744 = n2741 & n2743;
  assign n2745 = ~po63  & ~n2744;
  assign n2746 = ~n2454 & po41 ;
  assign n2747 = n2528 & ~n2746;
  assign n2748 = po63  & ~n2530;
  assign n2749 = ~n2747 & n2748;
  assign n2750 = ~n2740 & ~n2749;
  assign n2751 = ~n2745 & n2750;
  assign po40  = n2669 | ~n2751;
  assign n2753 = ~n2667 & ~n2668;
  assign n2754 = po40  & n2753;
  assign n2755 = ~n2546 & ~n2754;
  assign n2756 = n2546 & n2754;
  assign n2757 = ~n2755 & ~n2756;
  assign n2758 = pi80  & po40 ;
  assign n2759 = ~pi78  & ~pi79 ;
  assign n2760 = ~pi80  & n2759;
  assign n2761 = ~n2758 & ~n2760;
  assign n2762 = po41  & ~n2761;
  assign n2763 = ~po41  & n2761;
  assign n2764 = ~pi80  & po40 ;
  assign n2765 = pi81  & ~n2764;
  assign n2766 = ~pi81  & n2764;
  assign n2767 = ~n2765 & ~n2766;
  assign n2768 = ~n2763 & n2767;
  assign n2769 = ~n2762 & ~n2768;
  assign n2770 = po42  & ~n2769;
  assign n2771 = ~po42  & n2769;
  assign n2772 = po41  & n2751;
  assign n2773 = ~n2766 & ~n2772;
  assign n2774 = pi82  & ~n2773;
  assign n2775 = ~pi82  & n2773;
  assign n2776 = ~n2774 & ~n2775;
  assign n2777 = ~n2771 & ~n2776;
  assign n2778 = ~n2770 & ~n2777;
  assign n2779 = po43  & ~n2778;
  assign n2780 = ~po43  & n2778;
  assign n2781 = ~n2551 & ~n2552;
  assign n2782 = po40  & n2781;
  assign n2783 = n2556 & ~n2782;
  assign n2784 = ~n2556 & n2782;
  assign n2785 = ~n2783 & ~n2784;
  assign n2786 = ~n2780 & ~n2785;
  assign n2787 = ~n2779 & ~n2786;
  assign n2788 = po44  & ~n2787;
  assign n2789 = ~po44  & n2787;
  assign n2790 = ~n2559 & ~n2560;
  assign n2791 = po40  & n2790;
  assign n2792 = ~n2565 & ~n2791;
  assign n2793 = n2565 & n2791;
  assign n2794 = ~n2792 & ~n2793;
  assign n2795 = ~n2789 & ~n2794;
  assign n2796 = ~n2788 & ~n2795;
  assign n2797 = po45  & ~n2796;
  assign n2798 = ~po45  & n2796;
  assign n2799 = ~n2568 & ~n2569;
  assign n2800 = po40  & n2799;
  assign n2801 = n2574 & n2800;
  assign n2802 = ~n2574 & ~n2800;
  assign n2803 = ~n2801 & ~n2802;
  assign n2804 = ~n2798 & ~n2803;
  assign n2805 = ~n2797 & ~n2804;
  assign n2806 = po46  & ~n2805;
  assign n2807 = ~po46  & n2805;
  assign n2808 = ~n2577 & ~n2578;
  assign n2809 = po40  & n2808;
  assign n2810 = ~n2583 & ~n2809;
  assign n2811 = n2583 & n2809;
  assign n2812 = ~n2810 & ~n2811;
  assign n2813 = ~n2807 & ~n2812;
  assign n2814 = ~n2806 & ~n2813;
  assign n2815 = po47  & ~n2814;
  assign n2816 = ~po47  & n2814;
  assign n2817 = ~n2586 & ~n2587;
  assign n2818 = po40  & n2817;
  assign n2819 = ~n2592 & ~n2818;
  assign n2820 = n2592 & n2818;
  assign n2821 = ~n2819 & ~n2820;
  assign n2822 = ~n2816 & ~n2821;
  assign n2823 = ~n2815 & ~n2822;
  assign n2824 = po48  & ~n2823;
  assign n2825 = ~po48  & n2823;
  assign n2826 = ~n2595 & ~n2596;
  assign n2827 = po40  & n2826;
  assign n2828 = ~n2601 & ~n2827;
  assign n2829 = n2601 & n2827;
  assign n2830 = ~n2828 & ~n2829;
  assign n2831 = ~n2825 & ~n2830;
  assign n2832 = ~n2824 & ~n2831;
  assign n2833 = po49  & ~n2832;
  assign n2834 = ~po49  & n2832;
  assign n2835 = ~n2604 & ~n2605;
  assign n2836 = po40  & n2835;
  assign n2837 = ~n2610 & ~n2836;
  assign n2838 = n2610 & n2836;
  assign n2839 = ~n2837 & ~n2838;
  assign n2840 = ~n2834 & ~n2839;
  assign n2841 = ~n2833 & ~n2840;
  assign n2842 = po50  & ~n2841;
  assign n2843 = ~po50  & n2841;
  assign n2844 = ~n2613 & ~n2614;
  assign n2845 = po40  & n2844;
  assign n2846 = ~n2619 & ~n2845;
  assign n2847 = n2619 & n2845;
  assign n2848 = ~n2846 & ~n2847;
  assign n2849 = ~n2843 & ~n2848;
  assign n2850 = ~n2842 & ~n2849;
  assign n2851 = po51  & ~n2850;
  assign n2852 = ~po51  & n2850;
  assign n2853 = ~n2622 & ~n2623;
  assign n2854 = po40  & n2853;
  assign n2855 = ~n2628 & ~n2854;
  assign n2856 = n2628 & n2854;
  assign n2857 = ~n2855 & ~n2856;
  assign n2858 = ~n2852 & ~n2857;
  assign n2859 = ~n2851 & ~n2858;
  assign n2860 = po52  & ~n2859;
  assign n2861 = ~po52  & n2859;
  assign n2862 = ~n2631 & ~n2632;
  assign n2863 = po40  & n2862;
  assign n2864 = ~n2637 & ~n2863;
  assign n2865 = n2637 & n2863;
  assign n2866 = ~n2864 & ~n2865;
  assign n2867 = ~n2861 & ~n2866;
  assign n2868 = ~n2860 & ~n2867;
  assign n2869 = po53  & ~n2868;
  assign n2870 = ~po53  & n2868;
  assign n2871 = ~n2640 & ~n2641;
  assign n2872 = po40  & n2871;
  assign n2873 = ~n2646 & ~n2872;
  assign n2874 = n2646 & n2872;
  assign n2875 = ~n2873 & ~n2874;
  assign n2876 = ~n2870 & ~n2875;
  assign n2877 = ~n2869 & ~n2876;
  assign n2878 = po54  & ~n2877;
  assign n2879 = ~po54  & n2877;
  assign n2880 = ~n2649 & ~n2650;
  assign n2881 = po40  & n2880;
  assign n2882 = ~n2655 & ~n2881;
  assign n2883 = n2655 & n2881;
  assign n2884 = ~n2882 & ~n2883;
  assign n2885 = ~n2879 & ~n2884;
  assign n2886 = ~n2878 & ~n2885;
  assign n2887 = po55  & ~n2886;
  assign n2888 = ~po55  & n2886;
  assign n2889 = ~n2658 & ~n2659;
  assign n2890 = po40  & n2889;
  assign n2891 = ~n2664 & ~n2890;
  assign n2892 = n2664 & n2890;
  assign n2893 = ~n2891 & ~n2892;
  assign n2894 = ~n2888 & ~n2893;
  assign n2895 = ~n2887 & ~n2894;
  assign n2896 = po56  & ~n2895;
  assign n2897 = ~po56  & n2895;
  assign n2898 = n2674 & ~po40 ;
  assign n2899 = ~n2731 & ~n2732;
  assign n2900 = po40  & n2899;
  assign n2901 = ~n2737 & ~n2900;
  assign n2902 = n2737 & n2900;
  assign n2903 = ~n2901 & ~n2902;
  assign n2904 = ~n2757 & ~n2897;
  assign n2905 = ~n2896 & ~n2904;
  assign n2906 = po57  & ~n2905;
  assign n2907 = ~po57  & n2905;
  assign n2908 = ~n2677 & ~n2678;
  assign n2909 = po40  & n2908;
  assign n2910 = ~n2683 & ~n2909;
  assign n2911 = n2683 & n2909;
  assign n2912 = ~n2910 & ~n2911;
  assign n2913 = ~n2907 & ~n2912;
  assign n2914 = ~n2906 & ~n2913;
  assign n2915 = po58  & ~n2914;
  assign n2916 = ~po58  & n2914;
  assign n2917 = ~n2686 & ~n2687;
  assign n2918 = po40  & n2917;
  assign n2919 = ~n2692 & ~n2918;
  assign n2920 = n2692 & n2918;
  assign n2921 = ~n2919 & ~n2920;
  assign n2922 = ~n2916 & ~n2921;
  assign n2923 = ~n2915 & ~n2922;
  assign n2924 = po59  & ~n2923;
  assign n2925 = ~po59  & n2923;
  assign n2926 = ~n2695 & ~n2696;
  assign n2927 = po40  & n2926;
  assign n2928 = ~n2701 & ~n2927;
  assign n2929 = n2701 & n2927;
  assign n2930 = ~n2928 & ~n2929;
  assign n2931 = ~n2925 & ~n2930;
  assign n2932 = ~n2924 & ~n2931;
  assign n2933 = po60  & ~n2932;
  assign n2934 = ~po60  & n2932;
  assign n2935 = ~n2704 & ~n2705;
  assign n2936 = po40  & n2935;
  assign n2937 = ~n2710 & ~n2936;
  assign n2938 = n2710 & n2936;
  assign n2939 = ~n2937 & ~n2938;
  assign n2940 = ~n2934 & ~n2939;
  assign n2941 = ~n2933 & ~n2940;
  assign n2942 = po61  & ~n2941;
  assign n2943 = ~po61  & n2941;
  assign n2944 = ~n2713 & ~n2714;
  assign n2945 = po40  & n2944;
  assign n2946 = ~n2719 & ~n2945;
  assign n2947 = n2719 & n2945;
  assign n2948 = ~n2946 & ~n2947;
  assign n2949 = ~n2943 & ~n2948;
  assign n2950 = ~n2942 & ~n2949;
  assign n2951 = po62  & ~n2950;
  assign n2952 = ~po62  & n2950;
  assign n2953 = ~n2722 & ~n2723;
  assign n2954 = po40  & n2953;
  assign n2955 = ~n2728 & ~n2954;
  assign n2956 = n2728 & n2954;
  assign n2957 = ~n2955 & ~n2956;
  assign n2958 = ~n2952 & ~n2957;
  assign n2959 = ~n2951 & ~n2958;
  assign n2960 = n2903 & n2959;
  assign n2961 = ~n2903 & ~n2959;
  assign n2962 = n2741 & po40 ;
  assign n2963 = ~n2740 & ~n2962;
  assign n2964 = n2961 & n2963;
  assign n2965 = ~po63  & ~n2964;
  assign n2966 = ~n2674 & po40 ;
  assign n2967 = n2739 & ~n2966;
  assign n2968 = po63  & ~n2741;
  assign n2969 = ~n2967 & n2968;
  assign n2970 = ~n2960 & ~n2969;
  assign n2971 = ~n2965 & n2970;
  assign po39  = n2898 | ~n2971;
  assign n2973 = ~n2896 & ~n2897;
  assign n2974 = po39  & n2973;
  assign n2975 = ~n2757 & ~n2974;
  assign n2976 = n2757 & n2974;
  assign n2977 = ~n2975 & ~n2976;
  assign n2978 = pi78  & po39 ;
  assign n2979 = ~pi76  & ~pi77 ;
  assign n2980 = ~pi78  & n2979;
  assign n2981 = ~n2978 & ~n2980;
  assign n2982 = po40  & ~n2981;
  assign n2983 = ~po40  & n2981;
  assign n2984 = ~pi78  & po39 ;
  assign n2985 = pi79  & ~n2984;
  assign n2986 = ~pi79  & n2984;
  assign n2987 = ~n2985 & ~n2986;
  assign n2988 = ~n2983 & n2987;
  assign n2989 = ~n2982 & ~n2988;
  assign n2990 = po41  & ~n2989;
  assign n2991 = ~po41  & n2989;
  assign n2992 = po40  & n2971;
  assign n2993 = ~n2986 & ~n2992;
  assign n2994 = pi80  & ~n2993;
  assign n2995 = ~pi80  & n2993;
  assign n2996 = ~n2994 & ~n2995;
  assign n2997 = ~n2991 & ~n2996;
  assign n2998 = ~n2990 & ~n2997;
  assign n2999 = po42  & ~n2998;
  assign n3000 = ~po42  & n2998;
  assign n3001 = ~n2762 & ~n2763;
  assign n3002 = po39  & n3001;
  assign n3003 = n2767 & ~n3002;
  assign n3004 = ~n2767 & n3002;
  assign n3005 = ~n3003 & ~n3004;
  assign n3006 = ~n3000 & ~n3005;
  assign n3007 = ~n2999 & ~n3006;
  assign n3008 = po43  & ~n3007;
  assign n3009 = ~po43  & n3007;
  assign n3010 = ~n2770 & ~n2771;
  assign n3011 = po39  & n3010;
  assign n3012 = ~n2776 & ~n3011;
  assign n3013 = n2776 & n3011;
  assign n3014 = ~n3012 & ~n3013;
  assign n3015 = ~n3009 & ~n3014;
  assign n3016 = ~n3008 & ~n3015;
  assign n3017 = po44  & ~n3016;
  assign n3018 = ~po44  & n3016;
  assign n3019 = ~n2779 & ~n2780;
  assign n3020 = po39  & n3019;
  assign n3021 = n2785 & n3020;
  assign n3022 = ~n2785 & ~n3020;
  assign n3023 = ~n3021 & ~n3022;
  assign n3024 = ~n3018 & ~n3023;
  assign n3025 = ~n3017 & ~n3024;
  assign n3026 = po45  & ~n3025;
  assign n3027 = ~po45  & n3025;
  assign n3028 = ~n2788 & ~n2789;
  assign n3029 = po39  & n3028;
  assign n3030 = ~n2794 & ~n3029;
  assign n3031 = n2794 & n3029;
  assign n3032 = ~n3030 & ~n3031;
  assign n3033 = ~n3027 & ~n3032;
  assign n3034 = ~n3026 & ~n3033;
  assign n3035 = po46  & ~n3034;
  assign n3036 = ~po46  & n3034;
  assign n3037 = ~n2797 & ~n2798;
  assign n3038 = po39  & n3037;
  assign n3039 = ~n2803 & ~n3038;
  assign n3040 = n2803 & n3038;
  assign n3041 = ~n3039 & ~n3040;
  assign n3042 = ~n3036 & ~n3041;
  assign n3043 = ~n3035 & ~n3042;
  assign n3044 = po47  & ~n3043;
  assign n3045 = ~po47  & n3043;
  assign n3046 = ~n2806 & ~n2807;
  assign n3047 = po39  & n3046;
  assign n3048 = ~n2812 & ~n3047;
  assign n3049 = n2812 & n3047;
  assign n3050 = ~n3048 & ~n3049;
  assign n3051 = ~n3045 & ~n3050;
  assign n3052 = ~n3044 & ~n3051;
  assign n3053 = po48  & ~n3052;
  assign n3054 = ~po48  & n3052;
  assign n3055 = ~n2815 & ~n2816;
  assign n3056 = po39  & n3055;
  assign n3057 = ~n2821 & ~n3056;
  assign n3058 = n2821 & n3056;
  assign n3059 = ~n3057 & ~n3058;
  assign n3060 = ~n3054 & ~n3059;
  assign n3061 = ~n3053 & ~n3060;
  assign n3062 = po49  & ~n3061;
  assign n3063 = ~po49  & n3061;
  assign n3064 = ~n2824 & ~n2825;
  assign n3065 = po39  & n3064;
  assign n3066 = ~n2830 & ~n3065;
  assign n3067 = n2830 & n3065;
  assign n3068 = ~n3066 & ~n3067;
  assign n3069 = ~n3063 & ~n3068;
  assign n3070 = ~n3062 & ~n3069;
  assign n3071 = po50  & ~n3070;
  assign n3072 = ~po50  & n3070;
  assign n3073 = ~n2833 & ~n2834;
  assign n3074 = po39  & n3073;
  assign n3075 = ~n2839 & ~n3074;
  assign n3076 = n2839 & n3074;
  assign n3077 = ~n3075 & ~n3076;
  assign n3078 = ~n3072 & ~n3077;
  assign n3079 = ~n3071 & ~n3078;
  assign n3080 = po51  & ~n3079;
  assign n3081 = ~po51  & n3079;
  assign n3082 = ~n2842 & ~n2843;
  assign n3083 = po39  & n3082;
  assign n3084 = ~n2848 & ~n3083;
  assign n3085 = n2848 & n3083;
  assign n3086 = ~n3084 & ~n3085;
  assign n3087 = ~n3081 & ~n3086;
  assign n3088 = ~n3080 & ~n3087;
  assign n3089 = po52  & ~n3088;
  assign n3090 = ~po52  & n3088;
  assign n3091 = ~n2851 & ~n2852;
  assign n3092 = po39  & n3091;
  assign n3093 = ~n2857 & ~n3092;
  assign n3094 = n2857 & n3092;
  assign n3095 = ~n3093 & ~n3094;
  assign n3096 = ~n3090 & ~n3095;
  assign n3097 = ~n3089 & ~n3096;
  assign n3098 = po53  & ~n3097;
  assign n3099 = ~po53  & n3097;
  assign n3100 = ~n2860 & ~n2861;
  assign n3101 = po39  & n3100;
  assign n3102 = ~n2866 & ~n3101;
  assign n3103 = n2866 & n3101;
  assign n3104 = ~n3102 & ~n3103;
  assign n3105 = ~n3099 & ~n3104;
  assign n3106 = ~n3098 & ~n3105;
  assign n3107 = po54  & ~n3106;
  assign n3108 = ~po54  & n3106;
  assign n3109 = ~n2869 & ~n2870;
  assign n3110 = po39  & n3109;
  assign n3111 = ~n2875 & ~n3110;
  assign n3112 = n2875 & n3110;
  assign n3113 = ~n3111 & ~n3112;
  assign n3114 = ~n3108 & ~n3113;
  assign n3115 = ~n3107 & ~n3114;
  assign n3116 = po55  & ~n3115;
  assign n3117 = ~po55  & n3115;
  assign n3118 = ~n2878 & ~n2879;
  assign n3119 = po39  & n3118;
  assign n3120 = ~n2884 & ~n3119;
  assign n3121 = n2884 & n3119;
  assign n3122 = ~n3120 & ~n3121;
  assign n3123 = ~n3117 & ~n3122;
  assign n3124 = ~n3116 & ~n3123;
  assign n3125 = po56  & ~n3124;
  assign n3126 = ~po56  & n3124;
  assign n3127 = ~n2887 & ~n2888;
  assign n3128 = po39  & n3127;
  assign n3129 = ~n2893 & ~n3128;
  assign n3130 = n2893 & n3128;
  assign n3131 = ~n3129 & ~n3130;
  assign n3132 = ~n3126 & ~n3131;
  assign n3133 = ~n3125 & ~n3132;
  assign n3134 = po57  & ~n3133;
  assign n3135 = ~po57  & n3133;
  assign n3136 = n2903 & ~po39 ;
  assign n3137 = ~n2951 & ~n2952;
  assign n3138 = po39  & n3137;
  assign n3139 = ~n2957 & ~n3138;
  assign n3140 = n2957 & n3138;
  assign n3141 = ~n3139 & ~n3140;
  assign n3142 = ~n2977 & ~n3135;
  assign n3143 = ~n3134 & ~n3142;
  assign n3144 = po58  & ~n3143;
  assign n3145 = ~po58  & n3143;
  assign n3146 = ~n2906 & ~n2907;
  assign n3147 = po39  & n3146;
  assign n3148 = ~n2912 & ~n3147;
  assign n3149 = n2912 & n3147;
  assign n3150 = ~n3148 & ~n3149;
  assign n3151 = ~n3145 & ~n3150;
  assign n3152 = ~n3144 & ~n3151;
  assign n3153 = po59  & ~n3152;
  assign n3154 = ~po59  & n3152;
  assign n3155 = ~n2915 & ~n2916;
  assign n3156 = po39  & n3155;
  assign n3157 = ~n2921 & ~n3156;
  assign n3158 = n2921 & n3156;
  assign n3159 = ~n3157 & ~n3158;
  assign n3160 = ~n3154 & ~n3159;
  assign n3161 = ~n3153 & ~n3160;
  assign n3162 = po60  & ~n3161;
  assign n3163 = ~po60  & n3161;
  assign n3164 = ~n2924 & ~n2925;
  assign n3165 = po39  & n3164;
  assign n3166 = ~n2930 & ~n3165;
  assign n3167 = n2930 & n3165;
  assign n3168 = ~n3166 & ~n3167;
  assign n3169 = ~n3163 & ~n3168;
  assign n3170 = ~n3162 & ~n3169;
  assign n3171 = po61  & ~n3170;
  assign n3172 = ~po61  & n3170;
  assign n3173 = ~n2933 & ~n2934;
  assign n3174 = po39  & n3173;
  assign n3175 = ~n2939 & ~n3174;
  assign n3176 = n2939 & n3174;
  assign n3177 = ~n3175 & ~n3176;
  assign n3178 = ~n3172 & ~n3177;
  assign n3179 = ~n3171 & ~n3178;
  assign n3180 = po62  & ~n3179;
  assign n3181 = ~po62  & n3179;
  assign n3182 = ~n2942 & ~n2943;
  assign n3183 = po39  & n3182;
  assign n3184 = ~n2948 & ~n3183;
  assign n3185 = n2948 & n3183;
  assign n3186 = ~n3184 & ~n3185;
  assign n3187 = ~n3181 & ~n3186;
  assign n3188 = ~n3180 & ~n3187;
  assign n3189 = n3141 & n3188;
  assign n3190 = ~n3141 & ~n3188;
  assign n3191 = n2961 & po39 ;
  assign n3192 = ~n2960 & ~n3191;
  assign n3193 = n3190 & n3192;
  assign n3194 = ~po63  & ~n3193;
  assign n3195 = ~n2903 & po39 ;
  assign n3196 = n2959 & ~n3195;
  assign n3197 = po63  & ~n2961;
  assign n3198 = ~n3196 & n3197;
  assign n3199 = ~n3189 & ~n3198;
  assign n3200 = ~n3194 & n3199;
  assign po38  = n3136 | ~n3200;
  assign n3202 = ~n3134 & ~n3135;
  assign n3203 = po38  & n3202;
  assign n3204 = ~n2977 & ~n3203;
  assign n3205 = n2977 & n3203;
  assign n3206 = ~n3204 & ~n3205;
  assign n3207 = pi76  & po38 ;
  assign n3208 = ~pi74  & ~pi75 ;
  assign n3209 = ~pi76  & n3208;
  assign n3210 = ~n3207 & ~n3209;
  assign n3211 = po39  & ~n3210;
  assign n3212 = ~po39  & n3210;
  assign n3213 = ~pi76  & po38 ;
  assign n3214 = pi77  & ~n3213;
  assign n3215 = ~pi77  & n3213;
  assign n3216 = ~n3214 & ~n3215;
  assign n3217 = ~n3212 & n3216;
  assign n3218 = ~n3211 & ~n3217;
  assign n3219 = po40  & ~n3218;
  assign n3220 = ~po40  & n3218;
  assign n3221 = po39  & n3200;
  assign n3222 = ~n3215 & ~n3221;
  assign n3223 = pi78  & ~n3222;
  assign n3224 = ~pi78  & n3222;
  assign n3225 = ~n3223 & ~n3224;
  assign n3226 = ~n3220 & ~n3225;
  assign n3227 = ~n3219 & ~n3226;
  assign n3228 = po41  & ~n3227;
  assign n3229 = ~po41  & n3227;
  assign n3230 = ~n2982 & ~n2983;
  assign n3231 = po38  & n3230;
  assign n3232 = n2987 & ~n3231;
  assign n3233 = ~n2987 & n3231;
  assign n3234 = ~n3232 & ~n3233;
  assign n3235 = ~n3229 & ~n3234;
  assign n3236 = ~n3228 & ~n3235;
  assign n3237 = po42  & ~n3236;
  assign n3238 = ~po42  & n3236;
  assign n3239 = ~n2990 & ~n2991;
  assign n3240 = po38  & n3239;
  assign n3241 = ~n2996 & ~n3240;
  assign n3242 = n2996 & n3240;
  assign n3243 = ~n3241 & ~n3242;
  assign n3244 = ~n3238 & ~n3243;
  assign n3245 = ~n3237 & ~n3244;
  assign n3246 = po43  & ~n3245;
  assign n3247 = ~po43  & n3245;
  assign n3248 = ~n2999 & ~n3000;
  assign n3249 = po38  & n3248;
  assign n3250 = n3005 & n3249;
  assign n3251 = ~n3005 & ~n3249;
  assign n3252 = ~n3250 & ~n3251;
  assign n3253 = ~n3247 & ~n3252;
  assign n3254 = ~n3246 & ~n3253;
  assign n3255 = po44  & ~n3254;
  assign n3256 = ~po44  & n3254;
  assign n3257 = ~n3008 & ~n3009;
  assign n3258 = po38  & n3257;
  assign n3259 = ~n3014 & ~n3258;
  assign n3260 = n3014 & n3258;
  assign n3261 = ~n3259 & ~n3260;
  assign n3262 = ~n3256 & ~n3261;
  assign n3263 = ~n3255 & ~n3262;
  assign n3264 = po45  & ~n3263;
  assign n3265 = ~po45  & n3263;
  assign n3266 = ~n3017 & ~n3018;
  assign n3267 = po38  & n3266;
  assign n3268 = ~n3023 & ~n3267;
  assign n3269 = n3023 & n3267;
  assign n3270 = ~n3268 & ~n3269;
  assign n3271 = ~n3265 & ~n3270;
  assign n3272 = ~n3264 & ~n3271;
  assign n3273 = po46  & ~n3272;
  assign n3274 = ~po46  & n3272;
  assign n3275 = ~n3026 & ~n3027;
  assign n3276 = po38  & n3275;
  assign n3277 = ~n3032 & ~n3276;
  assign n3278 = n3032 & n3276;
  assign n3279 = ~n3277 & ~n3278;
  assign n3280 = ~n3274 & ~n3279;
  assign n3281 = ~n3273 & ~n3280;
  assign n3282 = po47  & ~n3281;
  assign n3283 = ~po47  & n3281;
  assign n3284 = ~n3035 & ~n3036;
  assign n3285 = po38  & n3284;
  assign n3286 = ~n3041 & ~n3285;
  assign n3287 = n3041 & n3285;
  assign n3288 = ~n3286 & ~n3287;
  assign n3289 = ~n3283 & ~n3288;
  assign n3290 = ~n3282 & ~n3289;
  assign n3291 = po48  & ~n3290;
  assign n3292 = ~po48  & n3290;
  assign n3293 = ~n3044 & ~n3045;
  assign n3294 = po38  & n3293;
  assign n3295 = ~n3050 & ~n3294;
  assign n3296 = n3050 & n3294;
  assign n3297 = ~n3295 & ~n3296;
  assign n3298 = ~n3292 & ~n3297;
  assign n3299 = ~n3291 & ~n3298;
  assign n3300 = po49  & ~n3299;
  assign n3301 = ~po49  & n3299;
  assign n3302 = ~n3053 & ~n3054;
  assign n3303 = po38  & n3302;
  assign n3304 = ~n3059 & ~n3303;
  assign n3305 = n3059 & n3303;
  assign n3306 = ~n3304 & ~n3305;
  assign n3307 = ~n3301 & ~n3306;
  assign n3308 = ~n3300 & ~n3307;
  assign n3309 = po50  & ~n3308;
  assign n3310 = ~po50  & n3308;
  assign n3311 = ~n3062 & ~n3063;
  assign n3312 = po38  & n3311;
  assign n3313 = ~n3068 & ~n3312;
  assign n3314 = n3068 & n3312;
  assign n3315 = ~n3313 & ~n3314;
  assign n3316 = ~n3310 & ~n3315;
  assign n3317 = ~n3309 & ~n3316;
  assign n3318 = po51  & ~n3317;
  assign n3319 = ~po51  & n3317;
  assign n3320 = ~n3071 & ~n3072;
  assign n3321 = po38  & n3320;
  assign n3322 = ~n3077 & ~n3321;
  assign n3323 = n3077 & n3321;
  assign n3324 = ~n3322 & ~n3323;
  assign n3325 = ~n3319 & ~n3324;
  assign n3326 = ~n3318 & ~n3325;
  assign n3327 = po52  & ~n3326;
  assign n3328 = ~po52  & n3326;
  assign n3329 = ~n3080 & ~n3081;
  assign n3330 = po38  & n3329;
  assign n3331 = ~n3086 & ~n3330;
  assign n3332 = n3086 & n3330;
  assign n3333 = ~n3331 & ~n3332;
  assign n3334 = ~n3328 & ~n3333;
  assign n3335 = ~n3327 & ~n3334;
  assign n3336 = po53  & ~n3335;
  assign n3337 = ~po53  & n3335;
  assign n3338 = ~n3089 & ~n3090;
  assign n3339 = po38  & n3338;
  assign n3340 = ~n3095 & ~n3339;
  assign n3341 = n3095 & n3339;
  assign n3342 = ~n3340 & ~n3341;
  assign n3343 = ~n3337 & ~n3342;
  assign n3344 = ~n3336 & ~n3343;
  assign n3345 = po54  & ~n3344;
  assign n3346 = ~po54  & n3344;
  assign n3347 = ~n3098 & ~n3099;
  assign n3348 = po38  & n3347;
  assign n3349 = ~n3104 & ~n3348;
  assign n3350 = n3104 & n3348;
  assign n3351 = ~n3349 & ~n3350;
  assign n3352 = ~n3346 & ~n3351;
  assign n3353 = ~n3345 & ~n3352;
  assign n3354 = po55  & ~n3353;
  assign n3355 = ~po55  & n3353;
  assign n3356 = ~n3107 & ~n3108;
  assign n3357 = po38  & n3356;
  assign n3358 = ~n3113 & ~n3357;
  assign n3359 = n3113 & n3357;
  assign n3360 = ~n3358 & ~n3359;
  assign n3361 = ~n3355 & ~n3360;
  assign n3362 = ~n3354 & ~n3361;
  assign n3363 = po56  & ~n3362;
  assign n3364 = ~po56  & n3362;
  assign n3365 = ~n3116 & ~n3117;
  assign n3366 = po38  & n3365;
  assign n3367 = ~n3122 & ~n3366;
  assign n3368 = n3122 & n3366;
  assign n3369 = ~n3367 & ~n3368;
  assign n3370 = ~n3364 & ~n3369;
  assign n3371 = ~n3363 & ~n3370;
  assign n3372 = po57  & ~n3371;
  assign n3373 = ~po57  & n3371;
  assign n3374 = ~n3125 & ~n3126;
  assign n3375 = po38  & n3374;
  assign n3376 = ~n3131 & ~n3375;
  assign n3377 = n3131 & n3375;
  assign n3378 = ~n3376 & ~n3377;
  assign n3379 = ~n3373 & ~n3378;
  assign n3380 = ~n3372 & ~n3379;
  assign n3381 = po58  & ~n3380;
  assign n3382 = ~po58  & n3380;
  assign n3383 = n3141 & ~po38 ;
  assign n3384 = ~n3180 & ~n3181;
  assign n3385 = po38  & n3384;
  assign n3386 = ~n3186 & ~n3385;
  assign n3387 = n3186 & n3385;
  assign n3388 = ~n3386 & ~n3387;
  assign n3389 = ~n3206 & ~n3382;
  assign n3390 = ~n3381 & ~n3389;
  assign n3391 = po59  & ~n3390;
  assign n3392 = ~po59  & n3390;
  assign n3393 = ~n3144 & ~n3145;
  assign n3394 = po38  & n3393;
  assign n3395 = ~n3150 & ~n3394;
  assign n3396 = n3150 & n3394;
  assign n3397 = ~n3395 & ~n3396;
  assign n3398 = ~n3392 & ~n3397;
  assign n3399 = ~n3391 & ~n3398;
  assign n3400 = po60  & ~n3399;
  assign n3401 = ~po60  & n3399;
  assign n3402 = ~n3153 & ~n3154;
  assign n3403 = po38  & n3402;
  assign n3404 = ~n3159 & ~n3403;
  assign n3405 = n3159 & n3403;
  assign n3406 = ~n3404 & ~n3405;
  assign n3407 = ~n3401 & ~n3406;
  assign n3408 = ~n3400 & ~n3407;
  assign n3409 = po61  & ~n3408;
  assign n3410 = ~po61  & n3408;
  assign n3411 = ~n3162 & ~n3163;
  assign n3412 = po38  & n3411;
  assign n3413 = ~n3168 & ~n3412;
  assign n3414 = n3168 & n3412;
  assign n3415 = ~n3413 & ~n3414;
  assign n3416 = ~n3410 & ~n3415;
  assign n3417 = ~n3409 & ~n3416;
  assign n3418 = po62  & ~n3417;
  assign n3419 = ~po62  & n3417;
  assign n3420 = ~n3171 & ~n3172;
  assign n3421 = po38  & n3420;
  assign n3422 = ~n3177 & ~n3421;
  assign n3423 = n3177 & n3421;
  assign n3424 = ~n3422 & ~n3423;
  assign n3425 = ~n3419 & ~n3424;
  assign n3426 = ~n3418 & ~n3425;
  assign n3427 = n3388 & n3426;
  assign n3428 = ~n3388 & ~n3426;
  assign n3429 = n3190 & po38 ;
  assign n3430 = ~n3189 & ~n3429;
  assign n3431 = n3428 & n3430;
  assign n3432 = ~po63  & ~n3431;
  assign n3433 = ~n3141 & po38 ;
  assign n3434 = n3188 & ~n3433;
  assign n3435 = po63  & ~n3190;
  assign n3436 = ~n3434 & n3435;
  assign n3437 = ~n3427 & ~n3436;
  assign n3438 = ~n3432 & n3437;
  assign po37  = n3383 | ~n3438;
  assign n3440 = ~n3381 & ~n3382;
  assign n3441 = po37  & n3440;
  assign n3442 = ~n3206 & ~n3441;
  assign n3443 = n3206 & n3441;
  assign n3444 = ~n3442 & ~n3443;
  assign n3445 = pi74  & po37 ;
  assign n3446 = ~pi72  & ~pi73 ;
  assign n3447 = ~pi74  & n3446;
  assign n3448 = ~n3445 & ~n3447;
  assign n3449 = po38  & ~n3448;
  assign n3450 = ~po38  & n3448;
  assign n3451 = ~pi74  & po37 ;
  assign n3452 = pi75  & ~n3451;
  assign n3453 = ~pi75  & n3451;
  assign n3454 = ~n3452 & ~n3453;
  assign n3455 = ~n3450 & n3454;
  assign n3456 = ~n3449 & ~n3455;
  assign n3457 = po39  & ~n3456;
  assign n3458 = ~po39  & n3456;
  assign n3459 = po38  & n3438;
  assign n3460 = ~n3453 & ~n3459;
  assign n3461 = pi76  & ~n3460;
  assign n3462 = ~pi76  & n3460;
  assign n3463 = ~n3461 & ~n3462;
  assign n3464 = ~n3458 & ~n3463;
  assign n3465 = ~n3457 & ~n3464;
  assign n3466 = po40  & ~n3465;
  assign n3467 = ~po40  & n3465;
  assign n3468 = ~n3211 & ~n3212;
  assign n3469 = po37  & n3468;
  assign n3470 = n3216 & ~n3469;
  assign n3471 = ~n3216 & n3469;
  assign n3472 = ~n3470 & ~n3471;
  assign n3473 = ~n3467 & ~n3472;
  assign n3474 = ~n3466 & ~n3473;
  assign n3475 = po41  & ~n3474;
  assign n3476 = ~po41  & n3474;
  assign n3477 = ~n3219 & ~n3220;
  assign n3478 = po37  & n3477;
  assign n3479 = ~n3225 & ~n3478;
  assign n3480 = n3225 & n3478;
  assign n3481 = ~n3479 & ~n3480;
  assign n3482 = ~n3476 & ~n3481;
  assign n3483 = ~n3475 & ~n3482;
  assign n3484 = po42  & ~n3483;
  assign n3485 = ~po42  & n3483;
  assign n3486 = ~n3228 & ~n3229;
  assign n3487 = po37  & n3486;
  assign n3488 = n3234 & n3487;
  assign n3489 = ~n3234 & ~n3487;
  assign n3490 = ~n3488 & ~n3489;
  assign n3491 = ~n3485 & ~n3490;
  assign n3492 = ~n3484 & ~n3491;
  assign n3493 = po43  & ~n3492;
  assign n3494 = ~po43  & n3492;
  assign n3495 = ~n3237 & ~n3238;
  assign n3496 = po37  & n3495;
  assign n3497 = ~n3243 & ~n3496;
  assign n3498 = n3243 & n3496;
  assign n3499 = ~n3497 & ~n3498;
  assign n3500 = ~n3494 & ~n3499;
  assign n3501 = ~n3493 & ~n3500;
  assign n3502 = po44  & ~n3501;
  assign n3503 = ~po44  & n3501;
  assign n3504 = ~n3246 & ~n3247;
  assign n3505 = po37  & n3504;
  assign n3506 = ~n3252 & ~n3505;
  assign n3507 = n3252 & n3505;
  assign n3508 = ~n3506 & ~n3507;
  assign n3509 = ~n3503 & ~n3508;
  assign n3510 = ~n3502 & ~n3509;
  assign n3511 = po45  & ~n3510;
  assign n3512 = ~po45  & n3510;
  assign n3513 = ~n3255 & ~n3256;
  assign n3514 = po37  & n3513;
  assign n3515 = ~n3261 & ~n3514;
  assign n3516 = n3261 & n3514;
  assign n3517 = ~n3515 & ~n3516;
  assign n3518 = ~n3512 & ~n3517;
  assign n3519 = ~n3511 & ~n3518;
  assign n3520 = po46  & ~n3519;
  assign n3521 = ~po46  & n3519;
  assign n3522 = ~n3264 & ~n3265;
  assign n3523 = po37  & n3522;
  assign n3524 = ~n3270 & ~n3523;
  assign n3525 = n3270 & n3523;
  assign n3526 = ~n3524 & ~n3525;
  assign n3527 = ~n3521 & ~n3526;
  assign n3528 = ~n3520 & ~n3527;
  assign n3529 = po47  & ~n3528;
  assign n3530 = ~po47  & n3528;
  assign n3531 = ~n3273 & ~n3274;
  assign n3532 = po37  & n3531;
  assign n3533 = ~n3279 & ~n3532;
  assign n3534 = n3279 & n3532;
  assign n3535 = ~n3533 & ~n3534;
  assign n3536 = ~n3530 & ~n3535;
  assign n3537 = ~n3529 & ~n3536;
  assign n3538 = po48  & ~n3537;
  assign n3539 = ~po48  & n3537;
  assign n3540 = ~n3282 & ~n3283;
  assign n3541 = po37  & n3540;
  assign n3542 = ~n3288 & ~n3541;
  assign n3543 = n3288 & n3541;
  assign n3544 = ~n3542 & ~n3543;
  assign n3545 = ~n3539 & ~n3544;
  assign n3546 = ~n3538 & ~n3545;
  assign n3547 = po49  & ~n3546;
  assign n3548 = ~po49  & n3546;
  assign n3549 = ~n3291 & ~n3292;
  assign n3550 = po37  & n3549;
  assign n3551 = ~n3297 & ~n3550;
  assign n3552 = n3297 & n3550;
  assign n3553 = ~n3551 & ~n3552;
  assign n3554 = ~n3548 & ~n3553;
  assign n3555 = ~n3547 & ~n3554;
  assign n3556 = po50  & ~n3555;
  assign n3557 = ~po50  & n3555;
  assign n3558 = ~n3300 & ~n3301;
  assign n3559 = po37  & n3558;
  assign n3560 = ~n3306 & ~n3559;
  assign n3561 = n3306 & n3559;
  assign n3562 = ~n3560 & ~n3561;
  assign n3563 = ~n3557 & ~n3562;
  assign n3564 = ~n3556 & ~n3563;
  assign n3565 = po51  & ~n3564;
  assign n3566 = ~po51  & n3564;
  assign n3567 = ~n3309 & ~n3310;
  assign n3568 = po37  & n3567;
  assign n3569 = ~n3315 & ~n3568;
  assign n3570 = n3315 & n3568;
  assign n3571 = ~n3569 & ~n3570;
  assign n3572 = ~n3566 & ~n3571;
  assign n3573 = ~n3565 & ~n3572;
  assign n3574 = po52  & ~n3573;
  assign n3575 = ~po52  & n3573;
  assign n3576 = ~n3318 & ~n3319;
  assign n3577 = po37  & n3576;
  assign n3578 = ~n3324 & ~n3577;
  assign n3579 = n3324 & n3577;
  assign n3580 = ~n3578 & ~n3579;
  assign n3581 = ~n3575 & ~n3580;
  assign n3582 = ~n3574 & ~n3581;
  assign n3583 = po53  & ~n3582;
  assign n3584 = ~po53  & n3582;
  assign n3585 = ~n3327 & ~n3328;
  assign n3586 = po37  & n3585;
  assign n3587 = ~n3333 & ~n3586;
  assign n3588 = n3333 & n3586;
  assign n3589 = ~n3587 & ~n3588;
  assign n3590 = ~n3584 & ~n3589;
  assign n3591 = ~n3583 & ~n3590;
  assign n3592 = po54  & ~n3591;
  assign n3593 = ~po54  & n3591;
  assign n3594 = ~n3336 & ~n3337;
  assign n3595 = po37  & n3594;
  assign n3596 = ~n3342 & ~n3595;
  assign n3597 = n3342 & n3595;
  assign n3598 = ~n3596 & ~n3597;
  assign n3599 = ~n3593 & ~n3598;
  assign n3600 = ~n3592 & ~n3599;
  assign n3601 = po55  & ~n3600;
  assign n3602 = ~po55  & n3600;
  assign n3603 = ~n3345 & ~n3346;
  assign n3604 = po37  & n3603;
  assign n3605 = ~n3351 & ~n3604;
  assign n3606 = n3351 & n3604;
  assign n3607 = ~n3605 & ~n3606;
  assign n3608 = ~n3602 & ~n3607;
  assign n3609 = ~n3601 & ~n3608;
  assign n3610 = po56  & ~n3609;
  assign n3611 = ~po56  & n3609;
  assign n3612 = ~n3354 & ~n3355;
  assign n3613 = po37  & n3612;
  assign n3614 = ~n3360 & ~n3613;
  assign n3615 = n3360 & n3613;
  assign n3616 = ~n3614 & ~n3615;
  assign n3617 = ~n3611 & ~n3616;
  assign n3618 = ~n3610 & ~n3617;
  assign n3619 = po57  & ~n3618;
  assign n3620 = ~po57  & n3618;
  assign n3621 = ~n3363 & ~n3364;
  assign n3622 = po37  & n3621;
  assign n3623 = ~n3369 & ~n3622;
  assign n3624 = n3369 & n3622;
  assign n3625 = ~n3623 & ~n3624;
  assign n3626 = ~n3620 & ~n3625;
  assign n3627 = ~n3619 & ~n3626;
  assign n3628 = po58  & ~n3627;
  assign n3629 = ~po58  & n3627;
  assign n3630 = ~n3372 & ~n3373;
  assign n3631 = po37  & n3630;
  assign n3632 = ~n3378 & ~n3631;
  assign n3633 = n3378 & n3631;
  assign n3634 = ~n3632 & ~n3633;
  assign n3635 = ~n3629 & ~n3634;
  assign n3636 = ~n3628 & ~n3635;
  assign n3637 = po59  & ~n3636;
  assign n3638 = ~po59  & n3636;
  assign n3639 = n3388 & ~po37 ;
  assign n3640 = ~n3418 & ~n3419;
  assign n3641 = po37  & n3640;
  assign n3642 = ~n3424 & ~n3641;
  assign n3643 = n3424 & n3641;
  assign n3644 = ~n3642 & ~n3643;
  assign n3645 = ~n3444 & ~n3638;
  assign n3646 = ~n3637 & ~n3645;
  assign n3647 = po60  & ~n3646;
  assign n3648 = ~po60  & n3646;
  assign n3649 = ~n3391 & ~n3392;
  assign n3650 = po37  & n3649;
  assign n3651 = ~n3397 & ~n3650;
  assign n3652 = n3397 & n3650;
  assign n3653 = ~n3651 & ~n3652;
  assign n3654 = ~n3648 & ~n3653;
  assign n3655 = ~n3647 & ~n3654;
  assign n3656 = po61  & ~n3655;
  assign n3657 = ~po61  & n3655;
  assign n3658 = ~n3400 & ~n3401;
  assign n3659 = po37  & n3658;
  assign n3660 = ~n3406 & ~n3659;
  assign n3661 = n3406 & n3659;
  assign n3662 = ~n3660 & ~n3661;
  assign n3663 = ~n3657 & ~n3662;
  assign n3664 = ~n3656 & ~n3663;
  assign n3665 = po62  & ~n3664;
  assign n3666 = ~po62  & n3664;
  assign n3667 = ~n3409 & ~n3410;
  assign n3668 = po37  & n3667;
  assign n3669 = ~n3415 & ~n3668;
  assign n3670 = n3415 & n3668;
  assign n3671 = ~n3669 & ~n3670;
  assign n3672 = ~n3666 & ~n3671;
  assign n3673 = ~n3665 & ~n3672;
  assign n3674 = n3644 & n3673;
  assign n3675 = ~n3644 & ~n3673;
  assign n3676 = n3428 & po37 ;
  assign n3677 = ~n3427 & ~n3676;
  assign n3678 = n3675 & n3677;
  assign n3679 = ~po63  & ~n3678;
  assign n3680 = ~n3388 & po37 ;
  assign n3681 = n3426 & ~n3680;
  assign n3682 = po63  & ~n3428;
  assign n3683 = ~n3681 & n3682;
  assign n3684 = ~n3674 & ~n3683;
  assign n3685 = ~n3679 & n3684;
  assign po36  = n3639 | ~n3685;
  assign n3687 = ~n3637 & ~n3638;
  assign n3688 = po36  & n3687;
  assign n3689 = ~n3444 & ~n3688;
  assign n3690 = n3444 & n3688;
  assign n3691 = ~n3689 & ~n3690;
  assign n3692 = pi72  & po36 ;
  assign n3693 = ~pi70  & ~pi71 ;
  assign n3694 = ~pi72  & n3693;
  assign n3695 = ~n3692 & ~n3694;
  assign n3696 = po37  & ~n3695;
  assign n3697 = ~po37  & n3695;
  assign n3698 = ~pi72  & po36 ;
  assign n3699 = pi73  & ~n3698;
  assign n3700 = ~pi73  & n3698;
  assign n3701 = ~n3699 & ~n3700;
  assign n3702 = ~n3697 & n3701;
  assign n3703 = ~n3696 & ~n3702;
  assign n3704 = po38  & ~n3703;
  assign n3705 = ~po38  & n3703;
  assign n3706 = po37  & n3685;
  assign n3707 = ~n3700 & ~n3706;
  assign n3708 = pi74  & ~n3707;
  assign n3709 = ~pi74  & n3707;
  assign n3710 = ~n3708 & ~n3709;
  assign n3711 = ~n3705 & ~n3710;
  assign n3712 = ~n3704 & ~n3711;
  assign n3713 = po39  & ~n3712;
  assign n3714 = ~po39  & n3712;
  assign n3715 = ~n3449 & ~n3450;
  assign n3716 = po36  & n3715;
  assign n3717 = n3454 & ~n3716;
  assign n3718 = ~n3454 & n3716;
  assign n3719 = ~n3717 & ~n3718;
  assign n3720 = ~n3714 & ~n3719;
  assign n3721 = ~n3713 & ~n3720;
  assign n3722 = po40  & ~n3721;
  assign n3723 = ~po40  & n3721;
  assign n3724 = ~n3457 & ~n3458;
  assign n3725 = po36  & n3724;
  assign n3726 = ~n3463 & ~n3725;
  assign n3727 = n3463 & n3725;
  assign n3728 = ~n3726 & ~n3727;
  assign n3729 = ~n3723 & ~n3728;
  assign n3730 = ~n3722 & ~n3729;
  assign n3731 = po41  & ~n3730;
  assign n3732 = ~po41  & n3730;
  assign n3733 = ~n3466 & ~n3467;
  assign n3734 = po36  & n3733;
  assign n3735 = n3472 & n3734;
  assign n3736 = ~n3472 & ~n3734;
  assign n3737 = ~n3735 & ~n3736;
  assign n3738 = ~n3732 & ~n3737;
  assign n3739 = ~n3731 & ~n3738;
  assign n3740 = po42  & ~n3739;
  assign n3741 = ~po42  & n3739;
  assign n3742 = ~n3475 & ~n3476;
  assign n3743 = po36  & n3742;
  assign n3744 = ~n3481 & ~n3743;
  assign n3745 = n3481 & n3743;
  assign n3746 = ~n3744 & ~n3745;
  assign n3747 = ~n3741 & ~n3746;
  assign n3748 = ~n3740 & ~n3747;
  assign n3749 = po43  & ~n3748;
  assign n3750 = ~po43  & n3748;
  assign n3751 = ~n3484 & ~n3485;
  assign n3752 = po36  & n3751;
  assign n3753 = ~n3490 & ~n3752;
  assign n3754 = n3490 & n3752;
  assign n3755 = ~n3753 & ~n3754;
  assign n3756 = ~n3750 & ~n3755;
  assign n3757 = ~n3749 & ~n3756;
  assign n3758 = po44  & ~n3757;
  assign n3759 = ~po44  & n3757;
  assign n3760 = ~n3493 & ~n3494;
  assign n3761 = po36  & n3760;
  assign n3762 = ~n3499 & ~n3761;
  assign n3763 = n3499 & n3761;
  assign n3764 = ~n3762 & ~n3763;
  assign n3765 = ~n3759 & ~n3764;
  assign n3766 = ~n3758 & ~n3765;
  assign n3767 = po45  & ~n3766;
  assign n3768 = ~po45  & n3766;
  assign n3769 = ~n3502 & ~n3503;
  assign n3770 = po36  & n3769;
  assign n3771 = ~n3508 & ~n3770;
  assign n3772 = n3508 & n3770;
  assign n3773 = ~n3771 & ~n3772;
  assign n3774 = ~n3768 & ~n3773;
  assign n3775 = ~n3767 & ~n3774;
  assign n3776 = po46  & ~n3775;
  assign n3777 = ~po46  & n3775;
  assign n3778 = ~n3511 & ~n3512;
  assign n3779 = po36  & n3778;
  assign n3780 = ~n3517 & ~n3779;
  assign n3781 = n3517 & n3779;
  assign n3782 = ~n3780 & ~n3781;
  assign n3783 = ~n3777 & ~n3782;
  assign n3784 = ~n3776 & ~n3783;
  assign n3785 = po47  & ~n3784;
  assign n3786 = ~po47  & n3784;
  assign n3787 = ~n3520 & ~n3521;
  assign n3788 = po36  & n3787;
  assign n3789 = ~n3526 & ~n3788;
  assign n3790 = n3526 & n3788;
  assign n3791 = ~n3789 & ~n3790;
  assign n3792 = ~n3786 & ~n3791;
  assign n3793 = ~n3785 & ~n3792;
  assign n3794 = po48  & ~n3793;
  assign n3795 = ~po48  & n3793;
  assign n3796 = ~n3529 & ~n3530;
  assign n3797 = po36  & n3796;
  assign n3798 = ~n3535 & ~n3797;
  assign n3799 = n3535 & n3797;
  assign n3800 = ~n3798 & ~n3799;
  assign n3801 = ~n3795 & ~n3800;
  assign n3802 = ~n3794 & ~n3801;
  assign n3803 = po49  & ~n3802;
  assign n3804 = ~po49  & n3802;
  assign n3805 = ~n3538 & ~n3539;
  assign n3806 = po36  & n3805;
  assign n3807 = ~n3544 & ~n3806;
  assign n3808 = n3544 & n3806;
  assign n3809 = ~n3807 & ~n3808;
  assign n3810 = ~n3804 & ~n3809;
  assign n3811 = ~n3803 & ~n3810;
  assign n3812 = po50  & ~n3811;
  assign n3813 = ~po50  & n3811;
  assign n3814 = ~n3547 & ~n3548;
  assign n3815 = po36  & n3814;
  assign n3816 = ~n3553 & ~n3815;
  assign n3817 = n3553 & n3815;
  assign n3818 = ~n3816 & ~n3817;
  assign n3819 = ~n3813 & ~n3818;
  assign n3820 = ~n3812 & ~n3819;
  assign n3821 = po51  & ~n3820;
  assign n3822 = ~po51  & n3820;
  assign n3823 = ~n3556 & ~n3557;
  assign n3824 = po36  & n3823;
  assign n3825 = ~n3562 & ~n3824;
  assign n3826 = n3562 & n3824;
  assign n3827 = ~n3825 & ~n3826;
  assign n3828 = ~n3822 & ~n3827;
  assign n3829 = ~n3821 & ~n3828;
  assign n3830 = po52  & ~n3829;
  assign n3831 = ~po52  & n3829;
  assign n3832 = ~n3565 & ~n3566;
  assign n3833 = po36  & n3832;
  assign n3834 = ~n3571 & ~n3833;
  assign n3835 = n3571 & n3833;
  assign n3836 = ~n3834 & ~n3835;
  assign n3837 = ~n3831 & ~n3836;
  assign n3838 = ~n3830 & ~n3837;
  assign n3839 = po53  & ~n3838;
  assign n3840 = ~po53  & n3838;
  assign n3841 = ~n3574 & ~n3575;
  assign n3842 = po36  & n3841;
  assign n3843 = ~n3580 & ~n3842;
  assign n3844 = n3580 & n3842;
  assign n3845 = ~n3843 & ~n3844;
  assign n3846 = ~n3840 & ~n3845;
  assign n3847 = ~n3839 & ~n3846;
  assign n3848 = po54  & ~n3847;
  assign n3849 = ~po54  & n3847;
  assign n3850 = ~n3583 & ~n3584;
  assign n3851 = po36  & n3850;
  assign n3852 = ~n3589 & ~n3851;
  assign n3853 = n3589 & n3851;
  assign n3854 = ~n3852 & ~n3853;
  assign n3855 = ~n3849 & ~n3854;
  assign n3856 = ~n3848 & ~n3855;
  assign n3857 = po55  & ~n3856;
  assign n3858 = ~po55  & n3856;
  assign n3859 = ~n3592 & ~n3593;
  assign n3860 = po36  & n3859;
  assign n3861 = ~n3598 & ~n3860;
  assign n3862 = n3598 & n3860;
  assign n3863 = ~n3861 & ~n3862;
  assign n3864 = ~n3858 & ~n3863;
  assign n3865 = ~n3857 & ~n3864;
  assign n3866 = po56  & ~n3865;
  assign n3867 = ~po56  & n3865;
  assign n3868 = ~n3601 & ~n3602;
  assign n3869 = po36  & n3868;
  assign n3870 = ~n3607 & ~n3869;
  assign n3871 = n3607 & n3869;
  assign n3872 = ~n3870 & ~n3871;
  assign n3873 = ~n3867 & ~n3872;
  assign n3874 = ~n3866 & ~n3873;
  assign n3875 = po57  & ~n3874;
  assign n3876 = ~po57  & n3874;
  assign n3877 = ~n3610 & ~n3611;
  assign n3878 = po36  & n3877;
  assign n3879 = ~n3616 & ~n3878;
  assign n3880 = n3616 & n3878;
  assign n3881 = ~n3879 & ~n3880;
  assign n3882 = ~n3876 & ~n3881;
  assign n3883 = ~n3875 & ~n3882;
  assign n3884 = po58  & ~n3883;
  assign n3885 = ~po58  & n3883;
  assign n3886 = ~n3619 & ~n3620;
  assign n3887 = po36  & n3886;
  assign n3888 = ~n3625 & ~n3887;
  assign n3889 = n3625 & n3887;
  assign n3890 = ~n3888 & ~n3889;
  assign n3891 = ~n3885 & ~n3890;
  assign n3892 = ~n3884 & ~n3891;
  assign n3893 = po59  & ~n3892;
  assign n3894 = ~po59  & n3892;
  assign n3895 = ~n3628 & ~n3629;
  assign n3896 = po36  & n3895;
  assign n3897 = ~n3634 & ~n3896;
  assign n3898 = n3634 & n3896;
  assign n3899 = ~n3897 & ~n3898;
  assign n3900 = ~n3894 & ~n3899;
  assign n3901 = ~n3893 & ~n3900;
  assign n3902 = po60  & ~n3901;
  assign n3903 = ~po60  & n3901;
  assign n3904 = n3644 & ~po36 ;
  assign n3905 = ~n3665 & ~n3666;
  assign n3906 = po36  & n3905;
  assign n3907 = ~n3671 & ~n3906;
  assign n3908 = n3671 & n3906;
  assign n3909 = ~n3907 & ~n3908;
  assign n3910 = ~n3691 & ~n3903;
  assign n3911 = ~n3902 & ~n3910;
  assign n3912 = po61  & ~n3911;
  assign n3913 = ~po61  & n3911;
  assign n3914 = ~n3647 & ~n3648;
  assign n3915 = po36  & n3914;
  assign n3916 = ~n3653 & ~n3915;
  assign n3917 = n3653 & n3915;
  assign n3918 = ~n3916 & ~n3917;
  assign n3919 = ~n3913 & ~n3918;
  assign n3920 = ~n3912 & ~n3919;
  assign n3921 = po62  & ~n3920;
  assign n3922 = ~po62  & n3920;
  assign n3923 = ~n3656 & ~n3657;
  assign n3924 = po36  & n3923;
  assign n3925 = ~n3662 & ~n3924;
  assign n3926 = n3662 & n3924;
  assign n3927 = ~n3925 & ~n3926;
  assign n3928 = ~n3922 & ~n3927;
  assign n3929 = ~n3921 & ~n3928;
  assign n3930 = n3909 & n3929;
  assign n3931 = ~n3909 & ~n3929;
  assign n3932 = n3675 & po36 ;
  assign n3933 = ~n3674 & ~n3932;
  assign n3934 = n3931 & n3933;
  assign n3935 = ~po63  & ~n3934;
  assign n3936 = ~n3644 & po36 ;
  assign n3937 = n3673 & ~n3936;
  assign n3938 = po63  & ~n3675;
  assign n3939 = ~n3937 & n3938;
  assign n3940 = ~n3930 & ~n3939;
  assign n3941 = ~n3935 & n3940;
  assign po35  = n3904 | ~n3941;
  assign n3943 = ~n3902 & ~n3903;
  assign n3944 = po35  & n3943;
  assign n3945 = ~n3691 & ~n3944;
  assign n3946 = n3691 & n3944;
  assign n3947 = ~n3945 & ~n3946;
  assign n3948 = pi70  & po35 ;
  assign n3949 = ~pi68  & ~pi69 ;
  assign n3950 = ~pi70  & n3949;
  assign n3951 = ~n3948 & ~n3950;
  assign n3952 = po36  & ~n3951;
  assign n3953 = ~po36  & n3951;
  assign n3954 = ~pi70  & po35 ;
  assign n3955 = pi71  & ~n3954;
  assign n3956 = ~pi71  & n3954;
  assign n3957 = ~n3955 & ~n3956;
  assign n3958 = ~n3953 & n3957;
  assign n3959 = ~n3952 & ~n3958;
  assign n3960 = po37  & ~n3959;
  assign n3961 = ~po37  & n3959;
  assign n3962 = po36  & n3941;
  assign n3963 = ~n3956 & ~n3962;
  assign n3964 = pi72  & ~n3963;
  assign n3965 = ~pi72  & n3963;
  assign n3966 = ~n3964 & ~n3965;
  assign n3967 = ~n3961 & ~n3966;
  assign n3968 = ~n3960 & ~n3967;
  assign n3969 = po38  & ~n3968;
  assign n3970 = ~po38  & n3968;
  assign n3971 = ~n3696 & ~n3697;
  assign n3972 = po35  & n3971;
  assign n3973 = n3701 & ~n3972;
  assign n3974 = ~n3701 & n3972;
  assign n3975 = ~n3973 & ~n3974;
  assign n3976 = ~n3970 & ~n3975;
  assign n3977 = ~n3969 & ~n3976;
  assign n3978 = po39  & ~n3977;
  assign n3979 = ~po39  & n3977;
  assign n3980 = ~n3704 & ~n3705;
  assign n3981 = po35  & n3980;
  assign n3982 = ~n3710 & ~n3981;
  assign n3983 = n3710 & n3981;
  assign n3984 = ~n3982 & ~n3983;
  assign n3985 = ~n3979 & ~n3984;
  assign n3986 = ~n3978 & ~n3985;
  assign n3987 = po40  & ~n3986;
  assign n3988 = ~po40  & n3986;
  assign n3989 = ~n3713 & ~n3714;
  assign n3990 = po35  & n3989;
  assign n3991 = n3719 & n3990;
  assign n3992 = ~n3719 & ~n3990;
  assign n3993 = ~n3991 & ~n3992;
  assign n3994 = ~n3988 & ~n3993;
  assign n3995 = ~n3987 & ~n3994;
  assign n3996 = po41  & ~n3995;
  assign n3997 = ~po41  & n3995;
  assign n3998 = ~n3722 & ~n3723;
  assign n3999 = po35  & n3998;
  assign n4000 = ~n3728 & ~n3999;
  assign n4001 = n3728 & n3999;
  assign n4002 = ~n4000 & ~n4001;
  assign n4003 = ~n3997 & ~n4002;
  assign n4004 = ~n3996 & ~n4003;
  assign n4005 = po42  & ~n4004;
  assign n4006 = ~po42  & n4004;
  assign n4007 = ~n3731 & ~n3732;
  assign n4008 = po35  & n4007;
  assign n4009 = ~n3737 & ~n4008;
  assign n4010 = n3737 & n4008;
  assign n4011 = ~n4009 & ~n4010;
  assign n4012 = ~n4006 & ~n4011;
  assign n4013 = ~n4005 & ~n4012;
  assign n4014 = po43  & ~n4013;
  assign n4015 = ~po43  & n4013;
  assign n4016 = ~n3740 & ~n3741;
  assign n4017 = po35  & n4016;
  assign n4018 = ~n3746 & ~n4017;
  assign n4019 = n3746 & n4017;
  assign n4020 = ~n4018 & ~n4019;
  assign n4021 = ~n4015 & ~n4020;
  assign n4022 = ~n4014 & ~n4021;
  assign n4023 = po44  & ~n4022;
  assign n4024 = ~po44  & n4022;
  assign n4025 = ~n3749 & ~n3750;
  assign n4026 = po35  & n4025;
  assign n4027 = ~n3755 & ~n4026;
  assign n4028 = n3755 & n4026;
  assign n4029 = ~n4027 & ~n4028;
  assign n4030 = ~n4024 & ~n4029;
  assign n4031 = ~n4023 & ~n4030;
  assign n4032 = po45  & ~n4031;
  assign n4033 = ~po45  & n4031;
  assign n4034 = ~n3758 & ~n3759;
  assign n4035 = po35  & n4034;
  assign n4036 = ~n3764 & ~n4035;
  assign n4037 = n3764 & n4035;
  assign n4038 = ~n4036 & ~n4037;
  assign n4039 = ~n4033 & ~n4038;
  assign n4040 = ~n4032 & ~n4039;
  assign n4041 = po46  & ~n4040;
  assign n4042 = ~po46  & n4040;
  assign n4043 = ~n3767 & ~n3768;
  assign n4044 = po35  & n4043;
  assign n4045 = ~n3773 & ~n4044;
  assign n4046 = n3773 & n4044;
  assign n4047 = ~n4045 & ~n4046;
  assign n4048 = ~n4042 & ~n4047;
  assign n4049 = ~n4041 & ~n4048;
  assign n4050 = po47  & ~n4049;
  assign n4051 = ~po47  & n4049;
  assign n4052 = ~n3776 & ~n3777;
  assign n4053 = po35  & n4052;
  assign n4054 = ~n3782 & ~n4053;
  assign n4055 = n3782 & n4053;
  assign n4056 = ~n4054 & ~n4055;
  assign n4057 = ~n4051 & ~n4056;
  assign n4058 = ~n4050 & ~n4057;
  assign n4059 = po48  & ~n4058;
  assign n4060 = ~po48  & n4058;
  assign n4061 = ~n3785 & ~n3786;
  assign n4062 = po35  & n4061;
  assign n4063 = ~n3791 & ~n4062;
  assign n4064 = n3791 & n4062;
  assign n4065 = ~n4063 & ~n4064;
  assign n4066 = ~n4060 & ~n4065;
  assign n4067 = ~n4059 & ~n4066;
  assign n4068 = po49  & ~n4067;
  assign n4069 = ~po49  & n4067;
  assign n4070 = ~n3794 & ~n3795;
  assign n4071 = po35  & n4070;
  assign n4072 = ~n3800 & ~n4071;
  assign n4073 = n3800 & n4071;
  assign n4074 = ~n4072 & ~n4073;
  assign n4075 = ~n4069 & ~n4074;
  assign n4076 = ~n4068 & ~n4075;
  assign n4077 = po50  & ~n4076;
  assign n4078 = ~po50  & n4076;
  assign n4079 = ~n3803 & ~n3804;
  assign n4080 = po35  & n4079;
  assign n4081 = ~n3809 & ~n4080;
  assign n4082 = n3809 & n4080;
  assign n4083 = ~n4081 & ~n4082;
  assign n4084 = ~n4078 & ~n4083;
  assign n4085 = ~n4077 & ~n4084;
  assign n4086 = po51  & ~n4085;
  assign n4087 = ~po51  & n4085;
  assign n4088 = ~n3812 & ~n3813;
  assign n4089 = po35  & n4088;
  assign n4090 = ~n3818 & ~n4089;
  assign n4091 = n3818 & n4089;
  assign n4092 = ~n4090 & ~n4091;
  assign n4093 = ~n4087 & ~n4092;
  assign n4094 = ~n4086 & ~n4093;
  assign n4095 = po52  & ~n4094;
  assign n4096 = ~po52  & n4094;
  assign n4097 = ~n3821 & ~n3822;
  assign n4098 = po35  & n4097;
  assign n4099 = ~n3827 & ~n4098;
  assign n4100 = n3827 & n4098;
  assign n4101 = ~n4099 & ~n4100;
  assign n4102 = ~n4096 & ~n4101;
  assign n4103 = ~n4095 & ~n4102;
  assign n4104 = po53  & ~n4103;
  assign n4105 = ~po53  & n4103;
  assign n4106 = ~n3830 & ~n3831;
  assign n4107 = po35  & n4106;
  assign n4108 = ~n3836 & ~n4107;
  assign n4109 = n3836 & n4107;
  assign n4110 = ~n4108 & ~n4109;
  assign n4111 = ~n4105 & ~n4110;
  assign n4112 = ~n4104 & ~n4111;
  assign n4113 = po54  & ~n4112;
  assign n4114 = ~po54  & n4112;
  assign n4115 = ~n3839 & ~n3840;
  assign n4116 = po35  & n4115;
  assign n4117 = ~n3845 & ~n4116;
  assign n4118 = n3845 & n4116;
  assign n4119 = ~n4117 & ~n4118;
  assign n4120 = ~n4114 & ~n4119;
  assign n4121 = ~n4113 & ~n4120;
  assign n4122 = po55  & ~n4121;
  assign n4123 = ~po55  & n4121;
  assign n4124 = ~n3848 & ~n3849;
  assign n4125 = po35  & n4124;
  assign n4126 = ~n3854 & ~n4125;
  assign n4127 = n3854 & n4125;
  assign n4128 = ~n4126 & ~n4127;
  assign n4129 = ~n4123 & ~n4128;
  assign n4130 = ~n4122 & ~n4129;
  assign n4131 = po56  & ~n4130;
  assign n4132 = ~po56  & n4130;
  assign n4133 = ~n3857 & ~n3858;
  assign n4134 = po35  & n4133;
  assign n4135 = ~n3863 & ~n4134;
  assign n4136 = n3863 & n4134;
  assign n4137 = ~n4135 & ~n4136;
  assign n4138 = ~n4132 & ~n4137;
  assign n4139 = ~n4131 & ~n4138;
  assign n4140 = po57  & ~n4139;
  assign n4141 = ~po57  & n4139;
  assign n4142 = ~n3866 & ~n3867;
  assign n4143 = po35  & n4142;
  assign n4144 = ~n3872 & ~n4143;
  assign n4145 = n3872 & n4143;
  assign n4146 = ~n4144 & ~n4145;
  assign n4147 = ~n4141 & ~n4146;
  assign n4148 = ~n4140 & ~n4147;
  assign n4149 = po58  & ~n4148;
  assign n4150 = ~po58  & n4148;
  assign n4151 = ~n3875 & ~n3876;
  assign n4152 = po35  & n4151;
  assign n4153 = ~n3881 & ~n4152;
  assign n4154 = n3881 & n4152;
  assign n4155 = ~n4153 & ~n4154;
  assign n4156 = ~n4150 & ~n4155;
  assign n4157 = ~n4149 & ~n4156;
  assign n4158 = po59  & ~n4157;
  assign n4159 = ~po59  & n4157;
  assign n4160 = ~n3884 & ~n3885;
  assign n4161 = po35  & n4160;
  assign n4162 = ~n3890 & ~n4161;
  assign n4163 = n3890 & n4161;
  assign n4164 = ~n4162 & ~n4163;
  assign n4165 = ~n4159 & ~n4164;
  assign n4166 = ~n4158 & ~n4165;
  assign n4167 = po60  & ~n4166;
  assign n4168 = ~po60  & n4166;
  assign n4169 = ~n3893 & ~n3894;
  assign n4170 = po35  & n4169;
  assign n4171 = ~n3899 & ~n4170;
  assign n4172 = n3899 & n4170;
  assign n4173 = ~n4171 & ~n4172;
  assign n4174 = ~n4168 & ~n4173;
  assign n4175 = ~n4167 & ~n4174;
  assign n4176 = po61  & ~n4175;
  assign n4177 = ~po61  & n4175;
  assign n4178 = n3909 & ~po35 ;
  assign n4179 = ~n3921 & ~n3922;
  assign n4180 = po35  & n4179;
  assign n4181 = ~n3927 & ~n4180;
  assign n4182 = n3927 & n4180;
  assign n4183 = ~n4181 & ~n4182;
  assign n4184 = ~n3947 & ~n4177;
  assign n4185 = ~n4176 & ~n4184;
  assign n4186 = po62  & ~n4185;
  assign n4187 = ~po62  & n4185;
  assign n4188 = ~n3912 & ~n3913;
  assign n4189 = po35  & n4188;
  assign n4190 = ~n3918 & ~n4189;
  assign n4191 = n3918 & n4189;
  assign n4192 = ~n4190 & ~n4191;
  assign n4193 = ~n4187 & ~n4192;
  assign n4194 = ~n4186 & ~n4193;
  assign n4195 = n4183 & n4194;
  assign n4196 = ~n4183 & ~n4194;
  assign n4197 = n3931 & po35 ;
  assign n4198 = ~n3930 & ~n4197;
  assign n4199 = n4196 & n4198;
  assign n4200 = ~po63  & ~n4199;
  assign n4201 = ~n3909 & po35 ;
  assign n4202 = n3929 & ~n4201;
  assign n4203 = po63  & ~n3931;
  assign n4204 = ~n4202 & n4203;
  assign n4205 = ~n4195 & ~n4204;
  assign n4206 = ~n4200 & n4205;
  assign po34  = n4178 | ~n4206;
  assign n4208 = ~n4176 & ~n4177;
  assign n4209 = po34  & n4208;
  assign n4210 = ~n3947 & ~n4209;
  assign n4211 = n3947 & n4209;
  assign n4212 = ~n4210 & ~n4211;
  assign n4213 = pi68  & po34 ;
  assign n4214 = ~pi66  & ~pi67 ;
  assign n4215 = ~pi68  & n4214;
  assign n4216 = ~n4213 & ~n4215;
  assign n4217 = po35  & ~n4216;
  assign n4218 = ~po35  & n4216;
  assign n4219 = ~pi68  & po34 ;
  assign n4220 = pi69  & ~n4219;
  assign n4221 = ~pi69  & n4219;
  assign n4222 = ~n4220 & ~n4221;
  assign n4223 = ~n4218 & n4222;
  assign n4224 = ~n4217 & ~n4223;
  assign n4225 = po36  & ~n4224;
  assign n4226 = ~po36  & n4224;
  assign n4227 = po35  & n4206;
  assign n4228 = ~n4221 & ~n4227;
  assign n4229 = pi70  & ~n4228;
  assign n4230 = ~pi70  & n4228;
  assign n4231 = ~n4229 & ~n4230;
  assign n4232 = ~n4226 & ~n4231;
  assign n4233 = ~n4225 & ~n4232;
  assign n4234 = po37  & ~n4233;
  assign n4235 = ~po37  & n4233;
  assign n4236 = ~n3952 & ~n3953;
  assign n4237 = po34  & n4236;
  assign n4238 = n3957 & ~n4237;
  assign n4239 = ~n3957 & n4237;
  assign n4240 = ~n4238 & ~n4239;
  assign n4241 = ~n4235 & ~n4240;
  assign n4242 = ~n4234 & ~n4241;
  assign n4243 = po38  & ~n4242;
  assign n4244 = ~po38  & n4242;
  assign n4245 = ~n3960 & ~n3961;
  assign n4246 = po34  & n4245;
  assign n4247 = ~n3966 & ~n4246;
  assign n4248 = n3966 & n4246;
  assign n4249 = ~n4247 & ~n4248;
  assign n4250 = ~n4244 & ~n4249;
  assign n4251 = ~n4243 & ~n4250;
  assign n4252 = po39  & ~n4251;
  assign n4253 = ~po39  & n4251;
  assign n4254 = ~n3969 & ~n3970;
  assign n4255 = po34  & n4254;
  assign n4256 = n3975 & n4255;
  assign n4257 = ~n3975 & ~n4255;
  assign n4258 = ~n4256 & ~n4257;
  assign n4259 = ~n4253 & ~n4258;
  assign n4260 = ~n4252 & ~n4259;
  assign n4261 = po40  & ~n4260;
  assign n4262 = ~po40  & n4260;
  assign n4263 = ~n3978 & ~n3979;
  assign n4264 = po34  & n4263;
  assign n4265 = ~n3984 & ~n4264;
  assign n4266 = n3984 & n4264;
  assign n4267 = ~n4265 & ~n4266;
  assign n4268 = ~n4262 & ~n4267;
  assign n4269 = ~n4261 & ~n4268;
  assign n4270 = po41  & ~n4269;
  assign n4271 = ~po41  & n4269;
  assign n4272 = ~n3987 & ~n3988;
  assign n4273 = po34  & n4272;
  assign n4274 = ~n3993 & ~n4273;
  assign n4275 = n3993 & n4273;
  assign n4276 = ~n4274 & ~n4275;
  assign n4277 = ~n4271 & ~n4276;
  assign n4278 = ~n4270 & ~n4277;
  assign n4279 = po42  & ~n4278;
  assign n4280 = ~po42  & n4278;
  assign n4281 = ~n3996 & ~n3997;
  assign n4282 = po34  & n4281;
  assign n4283 = ~n4002 & ~n4282;
  assign n4284 = n4002 & n4282;
  assign n4285 = ~n4283 & ~n4284;
  assign n4286 = ~n4280 & ~n4285;
  assign n4287 = ~n4279 & ~n4286;
  assign n4288 = po43  & ~n4287;
  assign n4289 = ~po43  & n4287;
  assign n4290 = ~n4005 & ~n4006;
  assign n4291 = po34  & n4290;
  assign n4292 = ~n4011 & ~n4291;
  assign n4293 = n4011 & n4291;
  assign n4294 = ~n4292 & ~n4293;
  assign n4295 = ~n4289 & ~n4294;
  assign n4296 = ~n4288 & ~n4295;
  assign n4297 = po44  & ~n4296;
  assign n4298 = ~po44  & n4296;
  assign n4299 = ~n4014 & ~n4015;
  assign n4300 = po34  & n4299;
  assign n4301 = ~n4020 & ~n4300;
  assign n4302 = n4020 & n4300;
  assign n4303 = ~n4301 & ~n4302;
  assign n4304 = ~n4298 & ~n4303;
  assign n4305 = ~n4297 & ~n4304;
  assign n4306 = po45  & ~n4305;
  assign n4307 = ~po45  & n4305;
  assign n4308 = ~n4023 & ~n4024;
  assign n4309 = po34  & n4308;
  assign n4310 = ~n4029 & ~n4309;
  assign n4311 = n4029 & n4309;
  assign n4312 = ~n4310 & ~n4311;
  assign n4313 = ~n4307 & ~n4312;
  assign n4314 = ~n4306 & ~n4313;
  assign n4315 = po46  & ~n4314;
  assign n4316 = ~po46  & n4314;
  assign n4317 = ~n4032 & ~n4033;
  assign n4318 = po34  & n4317;
  assign n4319 = ~n4038 & ~n4318;
  assign n4320 = n4038 & n4318;
  assign n4321 = ~n4319 & ~n4320;
  assign n4322 = ~n4316 & ~n4321;
  assign n4323 = ~n4315 & ~n4322;
  assign n4324 = po47  & ~n4323;
  assign n4325 = ~po47  & n4323;
  assign n4326 = ~n4041 & ~n4042;
  assign n4327 = po34  & n4326;
  assign n4328 = ~n4047 & ~n4327;
  assign n4329 = n4047 & n4327;
  assign n4330 = ~n4328 & ~n4329;
  assign n4331 = ~n4325 & ~n4330;
  assign n4332 = ~n4324 & ~n4331;
  assign n4333 = po48  & ~n4332;
  assign n4334 = ~po48  & n4332;
  assign n4335 = ~n4050 & ~n4051;
  assign n4336 = po34  & n4335;
  assign n4337 = ~n4056 & ~n4336;
  assign n4338 = n4056 & n4336;
  assign n4339 = ~n4337 & ~n4338;
  assign n4340 = ~n4334 & ~n4339;
  assign n4341 = ~n4333 & ~n4340;
  assign n4342 = po49  & ~n4341;
  assign n4343 = ~po49  & n4341;
  assign n4344 = ~n4059 & ~n4060;
  assign n4345 = po34  & n4344;
  assign n4346 = ~n4065 & ~n4345;
  assign n4347 = n4065 & n4345;
  assign n4348 = ~n4346 & ~n4347;
  assign n4349 = ~n4343 & ~n4348;
  assign n4350 = ~n4342 & ~n4349;
  assign n4351 = po50  & ~n4350;
  assign n4352 = ~po50  & n4350;
  assign n4353 = ~n4068 & ~n4069;
  assign n4354 = po34  & n4353;
  assign n4355 = ~n4074 & ~n4354;
  assign n4356 = n4074 & n4354;
  assign n4357 = ~n4355 & ~n4356;
  assign n4358 = ~n4352 & ~n4357;
  assign n4359 = ~n4351 & ~n4358;
  assign n4360 = po51  & ~n4359;
  assign n4361 = ~po51  & n4359;
  assign n4362 = ~n4077 & ~n4078;
  assign n4363 = po34  & n4362;
  assign n4364 = ~n4083 & ~n4363;
  assign n4365 = n4083 & n4363;
  assign n4366 = ~n4364 & ~n4365;
  assign n4367 = ~n4361 & ~n4366;
  assign n4368 = ~n4360 & ~n4367;
  assign n4369 = po52  & ~n4368;
  assign n4370 = ~po52  & n4368;
  assign n4371 = ~n4086 & ~n4087;
  assign n4372 = po34  & n4371;
  assign n4373 = ~n4092 & ~n4372;
  assign n4374 = n4092 & n4372;
  assign n4375 = ~n4373 & ~n4374;
  assign n4376 = ~n4370 & ~n4375;
  assign n4377 = ~n4369 & ~n4376;
  assign n4378 = po53  & ~n4377;
  assign n4379 = ~po53  & n4377;
  assign n4380 = ~n4095 & ~n4096;
  assign n4381 = po34  & n4380;
  assign n4382 = ~n4101 & ~n4381;
  assign n4383 = n4101 & n4381;
  assign n4384 = ~n4382 & ~n4383;
  assign n4385 = ~n4379 & ~n4384;
  assign n4386 = ~n4378 & ~n4385;
  assign n4387 = po54  & ~n4386;
  assign n4388 = ~po54  & n4386;
  assign n4389 = ~n4104 & ~n4105;
  assign n4390 = po34  & n4389;
  assign n4391 = ~n4110 & ~n4390;
  assign n4392 = n4110 & n4390;
  assign n4393 = ~n4391 & ~n4392;
  assign n4394 = ~n4388 & ~n4393;
  assign n4395 = ~n4387 & ~n4394;
  assign n4396 = po55  & ~n4395;
  assign n4397 = ~po55  & n4395;
  assign n4398 = ~n4113 & ~n4114;
  assign n4399 = po34  & n4398;
  assign n4400 = ~n4119 & ~n4399;
  assign n4401 = n4119 & n4399;
  assign n4402 = ~n4400 & ~n4401;
  assign n4403 = ~n4397 & ~n4402;
  assign n4404 = ~n4396 & ~n4403;
  assign n4405 = po56  & ~n4404;
  assign n4406 = ~po56  & n4404;
  assign n4407 = ~n4122 & ~n4123;
  assign n4408 = po34  & n4407;
  assign n4409 = ~n4128 & ~n4408;
  assign n4410 = n4128 & n4408;
  assign n4411 = ~n4409 & ~n4410;
  assign n4412 = ~n4406 & ~n4411;
  assign n4413 = ~n4405 & ~n4412;
  assign n4414 = po57  & ~n4413;
  assign n4415 = ~po57  & n4413;
  assign n4416 = ~n4131 & ~n4132;
  assign n4417 = po34  & n4416;
  assign n4418 = ~n4137 & ~n4417;
  assign n4419 = n4137 & n4417;
  assign n4420 = ~n4418 & ~n4419;
  assign n4421 = ~n4415 & ~n4420;
  assign n4422 = ~n4414 & ~n4421;
  assign n4423 = po58  & ~n4422;
  assign n4424 = ~po58  & n4422;
  assign n4425 = ~n4140 & ~n4141;
  assign n4426 = po34  & n4425;
  assign n4427 = ~n4146 & ~n4426;
  assign n4428 = n4146 & n4426;
  assign n4429 = ~n4427 & ~n4428;
  assign n4430 = ~n4424 & ~n4429;
  assign n4431 = ~n4423 & ~n4430;
  assign n4432 = po59  & ~n4431;
  assign n4433 = ~po59  & n4431;
  assign n4434 = ~n4149 & ~n4150;
  assign n4435 = po34  & n4434;
  assign n4436 = ~n4155 & ~n4435;
  assign n4437 = n4155 & n4435;
  assign n4438 = ~n4436 & ~n4437;
  assign n4439 = ~n4433 & ~n4438;
  assign n4440 = ~n4432 & ~n4439;
  assign n4441 = po60  & ~n4440;
  assign n4442 = ~po60  & n4440;
  assign n4443 = ~n4158 & ~n4159;
  assign n4444 = po34  & n4443;
  assign n4445 = ~n4164 & ~n4444;
  assign n4446 = n4164 & n4444;
  assign n4447 = ~n4445 & ~n4446;
  assign n4448 = ~n4442 & ~n4447;
  assign n4449 = ~n4441 & ~n4448;
  assign n4450 = po61  & ~n4449;
  assign n4451 = ~po61  & n4449;
  assign n4452 = ~n4167 & ~n4168;
  assign n4453 = po34  & n4452;
  assign n4454 = ~n4173 & ~n4453;
  assign n4455 = n4173 & n4453;
  assign n4456 = ~n4454 & ~n4455;
  assign n4457 = ~n4451 & ~n4456;
  assign n4458 = ~n4450 & ~n4457;
  assign n4459 = po62  & ~n4458;
  assign n4460 = ~po62  & n4458;
  assign n4461 = n4183 & ~po34 ;
  assign n4462 = ~n4186 & ~n4187;
  assign n4463 = po34  & n4462;
  assign n4464 = ~n4192 & ~n4463;
  assign n4465 = n4192 & n4463;
  assign n4466 = ~n4464 & ~n4465;
  assign n4467 = ~n4212 & ~n4460;
  assign n4468 = ~n4459 & ~n4467;
  assign n4469 = n4466 & n4468;
  assign n4470 = ~n4466 & ~n4468;
  assign n4471 = n4196 & po34 ;
  assign n4472 = ~n4195 & ~n4471;
  assign n4473 = n4470 & n4472;
  assign n4474 = ~po63  & ~n4473;
  assign n4475 = ~n4183 & po34 ;
  assign n4476 = n4194 & ~n4475;
  assign n4477 = po63  & ~n4196;
  assign n4478 = ~n4476 & n4477;
  assign n4479 = ~n4469 & ~n4478;
  assign n4480 = ~n4474 & n4479;
  assign po33  = n4461 | ~n4480;
  assign n4482 = ~n4459 & ~n4460;
  assign n4483 = po33  & n4482;
  assign n4484 = ~n4212 & ~n4483;
  assign n4485 = n4212 & n4483;
  assign n4486 = ~n4484 & ~n4485;
  assign n4487 = n4466 & ~po33 ;
  assign n4488 = pi66  & po33 ;
  assign n4489 = ~pi64  & ~pi65 ;
  assign n4490 = ~pi66  & n4489;
  assign n4491 = ~n4488 & ~n4490;
  assign n4492 = po34  & ~n4491;
  assign n4493 = ~po34  & n4491;
  assign n4494 = ~pi66  & po33 ;
  assign n4495 = pi67  & ~n4494;
  assign n4496 = ~pi67  & n4494;
  assign n4497 = ~n4495 & ~n4496;
  assign n4498 = ~n4493 & n4497;
  assign n4499 = ~n4492 & ~n4498;
  assign n4500 = po35  & ~n4499;
  assign n4501 = ~po35  & n4499;
  assign n4502 = po34  & n4480;
  assign n4503 = ~n4496 & ~n4502;
  assign n4504 = pi68  & ~n4503;
  assign n4505 = ~pi68  & n4503;
  assign n4506 = ~n4504 & ~n4505;
  assign n4507 = ~n4501 & ~n4506;
  assign n4508 = ~n4500 & ~n4507;
  assign n4509 = po36  & ~n4508;
  assign n4510 = ~po36  & n4508;
  assign n4511 = ~n4217 & ~n4218;
  assign n4512 = po33  & n4511;
  assign n4513 = n4222 & ~n4512;
  assign n4514 = ~n4222 & n4512;
  assign n4515 = ~n4513 & ~n4514;
  assign n4516 = ~n4510 & ~n4515;
  assign n4517 = ~n4509 & ~n4516;
  assign n4518 = po37  & ~n4517;
  assign n4519 = ~po37  & n4517;
  assign n4520 = ~n4225 & ~n4226;
  assign n4521 = po33  & n4520;
  assign n4522 = ~n4231 & ~n4521;
  assign n4523 = n4231 & n4521;
  assign n4524 = ~n4522 & ~n4523;
  assign n4525 = ~n4519 & ~n4524;
  assign n4526 = ~n4518 & ~n4525;
  assign n4527 = po38  & ~n4526;
  assign n4528 = ~po38  & n4526;
  assign n4529 = ~n4234 & ~n4235;
  assign n4530 = po33  & n4529;
  assign n4531 = n4240 & n4530;
  assign n4532 = ~n4240 & ~n4530;
  assign n4533 = ~n4531 & ~n4532;
  assign n4534 = ~n4528 & ~n4533;
  assign n4535 = ~n4527 & ~n4534;
  assign n4536 = po39  & ~n4535;
  assign n4537 = ~po39  & n4535;
  assign n4538 = ~n4243 & ~n4244;
  assign n4539 = po33  & n4538;
  assign n4540 = ~n4249 & ~n4539;
  assign n4541 = n4249 & n4539;
  assign n4542 = ~n4540 & ~n4541;
  assign n4543 = ~n4537 & ~n4542;
  assign n4544 = ~n4536 & ~n4543;
  assign n4545 = po40  & ~n4544;
  assign n4546 = ~po40  & n4544;
  assign n4547 = ~n4252 & ~n4253;
  assign n4548 = po33  & n4547;
  assign n4549 = ~n4258 & ~n4548;
  assign n4550 = n4258 & n4548;
  assign n4551 = ~n4549 & ~n4550;
  assign n4552 = ~n4546 & ~n4551;
  assign n4553 = ~n4545 & ~n4552;
  assign n4554 = po41  & ~n4553;
  assign n4555 = ~po41  & n4553;
  assign n4556 = ~n4261 & ~n4262;
  assign n4557 = po33  & n4556;
  assign n4558 = ~n4267 & ~n4557;
  assign n4559 = n4267 & n4557;
  assign n4560 = ~n4558 & ~n4559;
  assign n4561 = ~n4555 & ~n4560;
  assign n4562 = ~n4554 & ~n4561;
  assign n4563 = po42  & ~n4562;
  assign n4564 = ~po42  & n4562;
  assign n4565 = ~n4270 & ~n4271;
  assign n4566 = po33  & n4565;
  assign n4567 = ~n4276 & ~n4566;
  assign n4568 = n4276 & n4566;
  assign n4569 = ~n4567 & ~n4568;
  assign n4570 = ~n4564 & ~n4569;
  assign n4571 = ~n4563 & ~n4570;
  assign n4572 = po43  & ~n4571;
  assign n4573 = ~po43  & n4571;
  assign n4574 = ~n4279 & ~n4280;
  assign n4575 = po33  & n4574;
  assign n4576 = ~n4285 & ~n4575;
  assign n4577 = n4285 & n4575;
  assign n4578 = ~n4576 & ~n4577;
  assign n4579 = ~n4573 & ~n4578;
  assign n4580 = ~n4572 & ~n4579;
  assign n4581 = po44  & ~n4580;
  assign n4582 = ~po44  & n4580;
  assign n4583 = ~n4288 & ~n4289;
  assign n4584 = po33  & n4583;
  assign n4585 = ~n4294 & ~n4584;
  assign n4586 = n4294 & n4584;
  assign n4587 = ~n4585 & ~n4586;
  assign n4588 = ~n4582 & ~n4587;
  assign n4589 = ~n4581 & ~n4588;
  assign n4590 = po45  & ~n4589;
  assign n4591 = ~po45  & n4589;
  assign n4592 = ~n4297 & ~n4298;
  assign n4593 = po33  & n4592;
  assign n4594 = ~n4303 & ~n4593;
  assign n4595 = n4303 & n4593;
  assign n4596 = ~n4594 & ~n4595;
  assign n4597 = ~n4591 & ~n4596;
  assign n4598 = ~n4590 & ~n4597;
  assign n4599 = po46  & ~n4598;
  assign n4600 = ~po46  & n4598;
  assign n4601 = ~n4306 & ~n4307;
  assign n4602 = po33  & n4601;
  assign n4603 = ~n4312 & ~n4602;
  assign n4604 = n4312 & n4602;
  assign n4605 = ~n4603 & ~n4604;
  assign n4606 = ~n4600 & ~n4605;
  assign n4607 = ~n4599 & ~n4606;
  assign n4608 = po47  & ~n4607;
  assign n4609 = ~po47  & n4607;
  assign n4610 = ~n4315 & ~n4316;
  assign n4611 = po33  & n4610;
  assign n4612 = ~n4321 & ~n4611;
  assign n4613 = n4321 & n4611;
  assign n4614 = ~n4612 & ~n4613;
  assign n4615 = ~n4609 & ~n4614;
  assign n4616 = ~n4608 & ~n4615;
  assign n4617 = po48  & ~n4616;
  assign n4618 = ~po48  & n4616;
  assign n4619 = ~n4324 & ~n4325;
  assign n4620 = po33  & n4619;
  assign n4621 = ~n4330 & ~n4620;
  assign n4622 = n4330 & n4620;
  assign n4623 = ~n4621 & ~n4622;
  assign n4624 = ~n4618 & ~n4623;
  assign n4625 = ~n4617 & ~n4624;
  assign n4626 = po49  & ~n4625;
  assign n4627 = ~po49  & n4625;
  assign n4628 = ~n4333 & ~n4334;
  assign n4629 = po33  & n4628;
  assign n4630 = ~n4339 & ~n4629;
  assign n4631 = n4339 & n4629;
  assign n4632 = ~n4630 & ~n4631;
  assign n4633 = ~n4627 & ~n4632;
  assign n4634 = ~n4626 & ~n4633;
  assign n4635 = po50  & ~n4634;
  assign n4636 = ~po50  & n4634;
  assign n4637 = ~n4342 & ~n4343;
  assign n4638 = po33  & n4637;
  assign n4639 = ~n4348 & ~n4638;
  assign n4640 = n4348 & n4638;
  assign n4641 = ~n4639 & ~n4640;
  assign n4642 = ~n4636 & ~n4641;
  assign n4643 = ~n4635 & ~n4642;
  assign n4644 = po51  & ~n4643;
  assign n4645 = ~po51  & n4643;
  assign n4646 = ~n4351 & ~n4352;
  assign n4647 = po33  & n4646;
  assign n4648 = ~n4357 & ~n4647;
  assign n4649 = n4357 & n4647;
  assign n4650 = ~n4648 & ~n4649;
  assign n4651 = ~n4645 & ~n4650;
  assign n4652 = ~n4644 & ~n4651;
  assign n4653 = po52  & ~n4652;
  assign n4654 = ~po52  & n4652;
  assign n4655 = ~n4360 & ~n4361;
  assign n4656 = po33  & n4655;
  assign n4657 = ~n4366 & ~n4656;
  assign n4658 = n4366 & n4656;
  assign n4659 = ~n4657 & ~n4658;
  assign n4660 = ~n4654 & ~n4659;
  assign n4661 = ~n4653 & ~n4660;
  assign n4662 = po53  & ~n4661;
  assign n4663 = ~po53  & n4661;
  assign n4664 = ~n4369 & ~n4370;
  assign n4665 = po33  & n4664;
  assign n4666 = ~n4375 & ~n4665;
  assign n4667 = n4375 & n4665;
  assign n4668 = ~n4666 & ~n4667;
  assign n4669 = ~n4663 & ~n4668;
  assign n4670 = ~n4662 & ~n4669;
  assign n4671 = po54  & ~n4670;
  assign n4672 = ~po54  & n4670;
  assign n4673 = ~n4378 & ~n4379;
  assign n4674 = po33  & n4673;
  assign n4675 = ~n4384 & ~n4674;
  assign n4676 = n4384 & n4674;
  assign n4677 = ~n4675 & ~n4676;
  assign n4678 = ~n4672 & ~n4677;
  assign n4679 = ~n4671 & ~n4678;
  assign n4680 = po55  & ~n4679;
  assign n4681 = ~po55  & n4679;
  assign n4682 = ~n4387 & ~n4388;
  assign n4683 = po33  & n4682;
  assign n4684 = ~n4393 & ~n4683;
  assign n4685 = n4393 & n4683;
  assign n4686 = ~n4684 & ~n4685;
  assign n4687 = ~n4681 & ~n4686;
  assign n4688 = ~n4680 & ~n4687;
  assign n4689 = po56  & ~n4688;
  assign n4690 = ~po56  & n4688;
  assign n4691 = ~n4396 & ~n4397;
  assign n4692 = po33  & n4691;
  assign n4693 = ~n4402 & ~n4692;
  assign n4694 = n4402 & n4692;
  assign n4695 = ~n4693 & ~n4694;
  assign n4696 = ~n4690 & ~n4695;
  assign n4697 = ~n4689 & ~n4696;
  assign n4698 = po57  & ~n4697;
  assign n4699 = ~po57  & n4697;
  assign n4700 = ~n4405 & ~n4406;
  assign n4701 = po33  & n4700;
  assign n4702 = ~n4411 & ~n4701;
  assign n4703 = n4411 & n4701;
  assign n4704 = ~n4702 & ~n4703;
  assign n4705 = ~n4699 & ~n4704;
  assign n4706 = ~n4698 & ~n4705;
  assign n4707 = po58  & ~n4706;
  assign n4708 = ~po58  & n4706;
  assign n4709 = ~n4414 & ~n4415;
  assign n4710 = po33  & n4709;
  assign n4711 = ~n4420 & ~n4710;
  assign n4712 = n4420 & n4710;
  assign n4713 = ~n4711 & ~n4712;
  assign n4714 = ~n4708 & ~n4713;
  assign n4715 = ~n4707 & ~n4714;
  assign n4716 = po59  & ~n4715;
  assign n4717 = ~po59  & n4715;
  assign n4718 = ~n4423 & ~n4424;
  assign n4719 = po33  & n4718;
  assign n4720 = ~n4429 & ~n4719;
  assign n4721 = n4429 & n4719;
  assign n4722 = ~n4720 & ~n4721;
  assign n4723 = ~n4717 & ~n4722;
  assign n4724 = ~n4716 & ~n4723;
  assign n4725 = po60  & ~n4724;
  assign n4726 = ~po60  & n4724;
  assign n4727 = ~n4432 & ~n4433;
  assign n4728 = po33  & n4727;
  assign n4729 = ~n4438 & ~n4728;
  assign n4730 = n4438 & n4728;
  assign n4731 = ~n4729 & ~n4730;
  assign n4732 = ~n4726 & ~n4731;
  assign n4733 = ~n4725 & ~n4732;
  assign n4734 = po61  & ~n4733;
  assign n4735 = ~po61  & n4733;
  assign n4736 = ~n4441 & ~n4442;
  assign n4737 = po33  & n4736;
  assign n4738 = ~n4447 & ~n4737;
  assign n4739 = n4447 & n4737;
  assign n4740 = ~n4738 & ~n4739;
  assign n4741 = ~n4735 & ~n4740;
  assign n4742 = ~n4734 & ~n4741;
  assign n4743 = po62  & ~n4742;
  assign n4744 = ~po62  & n4742;
  assign n4745 = ~n4450 & ~n4451;
  assign n4746 = po33  & n4745;
  assign n4747 = ~n4456 & ~n4746;
  assign n4748 = n4456 & n4746;
  assign n4749 = ~n4747 & ~n4748;
  assign n4750 = ~n4744 & ~n4749;
  assign n4751 = ~n4743 & ~n4750;
  assign n4752 = n4486 & n4751;
  assign n4753 = ~n4486 & ~n4751;
  assign n4754 = n4470 & po33 ;
  assign n4755 = ~n4469 & ~n4754;
  assign n4756 = n4753 & n4755;
  assign n4757 = ~po63  & ~n4756;
  assign n4758 = ~n4466 & po33 ;
  assign n4759 = n4468 & ~n4758;
  assign n4760 = po63  & ~n4470;
  assign n4761 = ~n4759 & n4760;
  assign n4762 = ~n4752 & ~n4761;
  assign n4763 = ~n4757 & n4762;
  assign po32  = n4487 | ~n4763;
  assign n4765 = n4486 & ~po32 ;
  assign n4766 = ~n4743 & ~n4744;
  assign n4767 = po32  & n4766;
  assign n4768 = ~n4749 & ~n4767;
  assign n4769 = n4749 & n4767;
  assign n4770 = ~n4768 & ~n4769;
  assign n4771 = pi64  & po32 ;
  assign n4772 = ~pi62  & ~pi63 ;
  assign n4773 = ~pi64  & n4772;
  assign n4774 = ~n4771 & ~n4773;
  assign n4775 = po33  & ~n4774;
  assign n4776 = ~po33  & n4774;
  assign n4777 = ~pi64  & po32 ;
  assign n4778 = pi65  & ~n4777;
  assign n4779 = ~pi65  & n4777;
  assign n4780 = ~n4778 & ~n4779;
  assign n4781 = ~n4776 & n4780;
  assign n4782 = ~n4775 & ~n4781;
  assign n4783 = po34  & ~n4782;
  assign n4784 = ~po34  & n4782;
  assign n4785 = po33  & n4763;
  assign n4786 = ~n4779 & ~n4785;
  assign n4787 = pi66  & ~n4786;
  assign n4788 = ~pi66  & n4786;
  assign n4789 = ~n4787 & ~n4788;
  assign n4790 = ~n4784 & ~n4789;
  assign n4791 = ~n4783 & ~n4790;
  assign n4792 = po35  & ~n4791;
  assign n4793 = ~po35  & n4791;
  assign n4794 = ~n4492 & ~n4493;
  assign n4795 = po32  & n4794;
  assign n4796 = n4497 & ~n4795;
  assign n4797 = ~n4497 & n4795;
  assign n4798 = ~n4796 & ~n4797;
  assign n4799 = ~n4793 & ~n4798;
  assign n4800 = ~n4792 & ~n4799;
  assign n4801 = po36  & ~n4800;
  assign n4802 = ~po36  & n4800;
  assign n4803 = ~n4500 & ~n4501;
  assign n4804 = po32  & n4803;
  assign n4805 = ~n4506 & ~n4804;
  assign n4806 = n4506 & n4804;
  assign n4807 = ~n4805 & ~n4806;
  assign n4808 = ~n4802 & ~n4807;
  assign n4809 = ~n4801 & ~n4808;
  assign n4810 = po37  & ~n4809;
  assign n4811 = ~po37  & n4809;
  assign n4812 = ~n4509 & ~n4510;
  assign n4813 = po32  & n4812;
  assign n4814 = n4515 & n4813;
  assign n4815 = ~n4515 & ~n4813;
  assign n4816 = ~n4814 & ~n4815;
  assign n4817 = ~n4811 & ~n4816;
  assign n4818 = ~n4810 & ~n4817;
  assign n4819 = po38  & ~n4818;
  assign n4820 = ~po38  & n4818;
  assign n4821 = ~n4518 & ~n4519;
  assign n4822 = po32  & n4821;
  assign n4823 = ~n4524 & ~n4822;
  assign n4824 = n4524 & n4822;
  assign n4825 = ~n4823 & ~n4824;
  assign n4826 = ~n4820 & ~n4825;
  assign n4827 = ~n4819 & ~n4826;
  assign n4828 = po39  & ~n4827;
  assign n4829 = ~po39  & n4827;
  assign n4830 = ~n4527 & ~n4528;
  assign n4831 = po32  & n4830;
  assign n4832 = ~n4533 & ~n4831;
  assign n4833 = n4533 & n4831;
  assign n4834 = ~n4832 & ~n4833;
  assign n4835 = ~n4829 & ~n4834;
  assign n4836 = ~n4828 & ~n4835;
  assign n4837 = po40  & ~n4836;
  assign n4838 = ~po40  & n4836;
  assign n4839 = ~n4536 & ~n4537;
  assign n4840 = po32  & n4839;
  assign n4841 = ~n4542 & ~n4840;
  assign n4842 = n4542 & n4840;
  assign n4843 = ~n4841 & ~n4842;
  assign n4844 = ~n4838 & ~n4843;
  assign n4845 = ~n4837 & ~n4844;
  assign n4846 = po41  & ~n4845;
  assign n4847 = ~po41  & n4845;
  assign n4848 = ~n4545 & ~n4546;
  assign n4849 = po32  & n4848;
  assign n4850 = ~n4551 & ~n4849;
  assign n4851 = n4551 & n4849;
  assign n4852 = ~n4850 & ~n4851;
  assign n4853 = ~n4847 & ~n4852;
  assign n4854 = ~n4846 & ~n4853;
  assign n4855 = po42  & ~n4854;
  assign n4856 = ~po42  & n4854;
  assign n4857 = ~n4554 & ~n4555;
  assign n4858 = po32  & n4857;
  assign n4859 = ~n4560 & ~n4858;
  assign n4860 = n4560 & n4858;
  assign n4861 = ~n4859 & ~n4860;
  assign n4862 = ~n4856 & ~n4861;
  assign n4863 = ~n4855 & ~n4862;
  assign n4864 = po43  & ~n4863;
  assign n4865 = ~po43  & n4863;
  assign n4866 = ~n4563 & ~n4564;
  assign n4867 = po32  & n4866;
  assign n4868 = ~n4569 & ~n4867;
  assign n4869 = n4569 & n4867;
  assign n4870 = ~n4868 & ~n4869;
  assign n4871 = ~n4865 & ~n4870;
  assign n4872 = ~n4864 & ~n4871;
  assign n4873 = po44  & ~n4872;
  assign n4874 = ~po44  & n4872;
  assign n4875 = ~n4572 & ~n4573;
  assign n4876 = po32  & n4875;
  assign n4877 = ~n4578 & ~n4876;
  assign n4878 = n4578 & n4876;
  assign n4879 = ~n4877 & ~n4878;
  assign n4880 = ~n4874 & ~n4879;
  assign n4881 = ~n4873 & ~n4880;
  assign n4882 = po45  & ~n4881;
  assign n4883 = ~po45  & n4881;
  assign n4884 = ~n4581 & ~n4582;
  assign n4885 = po32  & n4884;
  assign n4886 = ~n4587 & ~n4885;
  assign n4887 = n4587 & n4885;
  assign n4888 = ~n4886 & ~n4887;
  assign n4889 = ~n4883 & ~n4888;
  assign n4890 = ~n4882 & ~n4889;
  assign n4891 = po46  & ~n4890;
  assign n4892 = ~po46  & n4890;
  assign n4893 = ~n4590 & ~n4591;
  assign n4894 = po32  & n4893;
  assign n4895 = ~n4596 & ~n4894;
  assign n4896 = n4596 & n4894;
  assign n4897 = ~n4895 & ~n4896;
  assign n4898 = ~n4892 & ~n4897;
  assign n4899 = ~n4891 & ~n4898;
  assign n4900 = po47  & ~n4899;
  assign n4901 = ~po47  & n4899;
  assign n4902 = ~n4599 & ~n4600;
  assign n4903 = po32  & n4902;
  assign n4904 = ~n4605 & ~n4903;
  assign n4905 = n4605 & n4903;
  assign n4906 = ~n4904 & ~n4905;
  assign n4907 = ~n4901 & ~n4906;
  assign n4908 = ~n4900 & ~n4907;
  assign n4909 = po48  & ~n4908;
  assign n4910 = ~po48  & n4908;
  assign n4911 = ~n4608 & ~n4609;
  assign n4912 = po32  & n4911;
  assign n4913 = ~n4614 & ~n4912;
  assign n4914 = n4614 & n4912;
  assign n4915 = ~n4913 & ~n4914;
  assign n4916 = ~n4910 & ~n4915;
  assign n4917 = ~n4909 & ~n4916;
  assign n4918 = po49  & ~n4917;
  assign n4919 = ~po49  & n4917;
  assign n4920 = ~n4617 & ~n4618;
  assign n4921 = po32  & n4920;
  assign n4922 = ~n4623 & ~n4921;
  assign n4923 = n4623 & n4921;
  assign n4924 = ~n4922 & ~n4923;
  assign n4925 = ~n4919 & ~n4924;
  assign n4926 = ~n4918 & ~n4925;
  assign n4927 = po50  & ~n4926;
  assign n4928 = ~po50  & n4926;
  assign n4929 = ~n4626 & ~n4627;
  assign n4930 = po32  & n4929;
  assign n4931 = ~n4632 & ~n4930;
  assign n4932 = n4632 & n4930;
  assign n4933 = ~n4931 & ~n4932;
  assign n4934 = ~n4928 & ~n4933;
  assign n4935 = ~n4927 & ~n4934;
  assign n4936 = po51  & ~n4935;
  assign n4937 = ~po51  & n4935;
  assign n4938 = ~n4635 & ~n4636;
  assign n4939 = po32  & n4938;
  assign n4940 = ~n4641 & ~n4939;
  assign n4941 = n4641 & n4939;
  assign n4942 = ~n4940 & ~n4941;
  assign n4943 = ~n4937 & ~n4942;
  assign n4944 = ~n4936 & ~n4943;
  assign n4945 = po52  & ~n4944;
  assign n4946 = ~po52  & n4944;
  assign n4947 = ~n4644 & ~n4645;
  assign n4948 = po32  & n4947;
  assign n4949 = ~n4650 & ~n4948;
  assign n4950 = n4650 & n4948;
  assign n4951 = ~n4949 & ~n4950;
  assign n4952 = ~n4946 & ~n4951;
  assign n4953 = ~n4945 & ~n4952;
  assign n4954 = po53  & ~n4953;
  assign n4955 = ~po53  & n4953;
  assign n4956 = ~n4653 & ~n4654;
  assign n4957 = po32  & n4956;
  assign n4958 = ~n4659 & ~n4957;
  assign n4959 = n4659 & n4957;
  assign n4960 = ~n4958 & ~n4959;
  assign n4961 = ~n4955 & ~n4960;
  assign n4962 = ~n4954 & ~n4961;
  assign n4963 = po54  & ~n4962;
  assign n4964 = ~po54  & n4962;
  assign n4965 = ~n4662 & ~n4663;
  assign n4966 = po32  & n4965;
  assign n4967 = ~n4668 & ~n4966;
  assign n4968 = n4668 & n4966;
  assign n4969 = ~n4967 & ~n4968;
  assign n4970 = ~n4964 & ~n4969;
  assign n4971 = ~n4963 & ~n4970;
  assign n4972 = po55  & ~n4971;
  assign n4973 = ~po55  & n4971;
  assign n4974 = ~n4671 & ~n4672;
  assign n4975 = po32  & n4974;
  assign n4976 = ~n4677 & ~n4975;
  assign n4977 = n4677 & n4975;
  assign n4978 = ~n4976 & ~n4977;
  assign n4979 = ~n4973 & ~n4978;
  assign n4980 = ~n4972 & ~n4979;
  assign n4981 = po56  & ~n4980;
  assign n4982 = ~po56  & n4980;
  assign n4983 = ~n4680 & ~n4681;
  assign n4984 = po32  & n4983;
  assign n4985 = ~n4686 & ~n4984;
  assign n4986 = n4686 & n4984;
  assign n4987 = ~n4985 & ~n4986;
  assign n4988 = ~n4982 & ~n4987;
  assign n4989 = ~n4981 & ~n4988;
  assign n4990 = po57  & ~n4989;
  assign n4991 = ~po57  & n4989;
  assign n4992 = ~n4689 & ~n4690;
  assign n4993 = po32  & n4992;
  assign n4994 = ~n4695 & ~n4993;
  assign n4995 = n4695 & n4993;
  assign n4996 = ~n4994 & ~n4995;
  assign n4997 = ~n4991 & ~n4996;
  assign n4998 = ~n4990 & ~n4997;
  assign n4999 = po58  & ~n4998;
  assign n5000 = ~po58  & n4998;
  assign n5001 = ~n4698 & ~n4699;
  assign n5002 = po32  & n5001;
  assign n5003 = ~n4704 & ~n5002;
  assign n5004 = n4704 & n5002;
  assign n5005 = ~n5003 & ~n5004;
  assign n5006 = ~n5000 & ~n5005;
  assign n5007 = ~n4999 & ~n5006;
  assign n5008 = po59  & ~n5007;
  assign n5009 = ~po59  & n5007;
  assign n5010 = ~n4707 & ~n4708;
  assign n5011 = po32  & n5010;
  assign n5012 = ~n4713 & ~n5011;
  assign n5013 = n4713 & n5011;
  assign n5014 = ~n5012 & ~n5013;
  assign n5015 = ~n5009 & ~n5014;
  assign n5016 = ~n5008 & ~n5015;
  assign n5017 = po60  & ~n5016;
  assign n5018 = ~po60  & n5016;
  assign n5019 = ~n4716 & ~n4717;
  assign n5020 = po32  & n5019;
  assign n5021 = ~n4722 & ~n5020;
  assign n5022 = n4722 & n5020;
  assign n5023 = ~n5021 & ~n5022;
  assign n5024 = ~n5018 & ~n5023;
  assign n5025 = ~n5017 & ~n5024;
  assign n5026 = po61  & ~n5025;
  assign n5027 = ~po61  & n5025;
  assign n5028 = ~n4725 & ~n4726;
  assign n5029 = po32  & n5028;
  assign n5030 = ~n4731 & ~n5029;
  assign n5031 = n4731 & n5029;
  assign n5032 = ~n5030 & ~n5031;
  assign n5033 = ~n5027 & ~n5032;
  assign n5034 = ~n5026 & ~n5033;
  assign n5035 = po62  & ~n5034;
  assign n5036 = ~po62  & n5034;
  assign n5037 = ~n4734 & ~n4735;
  assign n5038 = po32  & n5037;
  assign n5039 = ~n4740 & ~n5038;
  assign n5040 = n4740 & n5038;
  assign n5041 = ~n5039 & ~n5040;
  assign n5042 = ~n5036 & ~n5041;
  assign n5043 = ~n5035 & ~n5042;
  assign n5044 = n4770 & n5043;
  assign n5045 = ~n4770 & ~n5043;
  assign n5046 = n4753 & po32 ;
  assign n5047 = ~n4752 & ~n5046;
  assign n5048 = n5045 & n5047;
  assign n5049 = ~po63  & ~n5048;
  assign n5050 = ~n4486 & po32 ;
  assign n5051 = n4751 & ~n5050;
  assign n5052 = po63  & ~n4753;
  assign n5053 = ~n5051 & n5052;
  assign n5054 = ~n5044 & ~n5053;
  assign n5055 = ~n5049 & n5054;
  assign po31  = n4765 | ~n5055;
  assign n5057 = ~pi62  & po31 ;
  assign n5058 = ~pi63  & n5057;
  assign n5059 = po32  & n5055;
  assign n5060 = ~n5058 & ~n5059;
  assign n5061 = pi64  & ~n5060;
  assign n5062 = ~pi64  & n5060;
  assign n5063 = ~n5061 & ~n5062;
  assign n5064 = pi62  & po31 ;
  assign n5065 = ~pi60  & ~pi61 ;
  assign n5066 = ~pi62  & n5065;
  assign n5067 = ~n5064 & ~n5066;
  assign n5068 = po32  & ~n5067;
  assign n5069 = pi63  & ~n5057;
  assign n5070 = ~n5058 & ~n5069;
  assign n5071 = ~po32  & n5067;
  assign n5072 = n5070 & ~n5071;
  assign n5073 = ~n5068 & ~n5072;
  assign n5074 = po33  & ~n5073;
  assign n5075 = ~po33  & n5073;
  assign n5076 = n4770 & ~po31 ;
  assign n5077 = ~n5035 & ~n5036;
  assign n5078 = po31  & n5077;
  assign n5079 = ~n5041 & ~n5078;
  assign n5080 = n5041 & n5078;
  assign n5081 = ~n5079 & ~n5080;
  assign n5082 = ~n5063 & ~n5075;
  assign n5083 = ~n5074 & ~n5082;
  assign n5084 = po34  & ~n5083;
  assign n5085 = ~po34  & n5083;
  assign n5086 = ~n4775 & ~n4776;
  assign n5087 = po31  & n5086;
  assign n5088 = n4780 & ~n5087;
  assign n5089 = ~n4780 & n5087;
  assign n5090 = ~n5088 & ~n5089;
  assign n5091 = ~n5085 & ~n5090;
  assign n5092 = ~n5084 & ~n5091;
  assign n5093 = po35  & ~n5092;
  assign n5094 = ~po35  & n5092;
  assign n5095 = ~n4783 & ~n4784;
  assign n5096 = po31  & n5095;
  assign n5097 = ~n4789 & ~n5096;
  assign n5098 = n4789 & n5096;
  assign n5099 = ~n5097 & ~n5098;
  assign n5100 = ~n5094 & ~n5099;
  assign n5101 = ~n5093 & ~n5100;
  assign n5102 = po36  & ~n5101;
  assign n5103 = ~po36  & n5101;
  assign n5104 = ~n4792 & ~n4793;
  assign n5105 = po31  & n5104;
  assign n5106 = n4798 & n5105;
  assign n5107 = ~n4798 & ~n5105;
  assign n5108 = ~n5106 & ~n5107;
  assign n5109 = ~n5103 & ~n5108;
  assign n5110 = ~n5102 & ~n5109;
  assign n5111 = po37  & ~n5110;
  assign n5112 = ~po37  & n5110;
  assign n5113 = ~n4801 & ~n4802;
  assign n5114 = po31  & n5113;
  assign n5115 = ~n4807 & ~n5114;
  assign n5116 = n4807 & n5114;
  assign n5117 = ~n5115 & ~n5116;
  assign n5118 = ~n5112 & ~n5117;
  assign n5119 = ~n5111 & ~n5118;
  assign n5120 = po38  & ~n5119;
  assign n5121 = ~po38  & n5119;
  assign n5122 = ~n4810 & ~n4811;
  assign n5123 = po31  & n5122;
  assign n5124 = ~n4816 & ~n5123;
  assign n5125 = n4816 & n5123;
  assign n5126 = ~n5124 & ~n5125;
  assign n5127 = ~n5121 & ~n5126;
  assign n5128 = ~n5120 & ~n5127;
  assign n5129 = po39  & ~n5128;
  assign n5130 = ~po39  & n5128;
  assign n5131 = ~n4819 & ~n4820;
  assign n5132 = po31  & n5131;
  assign n5133 = ~n4825 & ~n5132;
  assign n5134 = n4825 & n5132;
  assign n5135 = ~n5133 & ~n5134;
  assign n5136 = ~n5130 & ~n5135;
  assign n5137 = ~n5129 & ~n5136;
  assign n5138 = po40  & ~n5137;
  assign n5139 = ~po40  & n5137;
  assign n5140 = ~n4828 & ~n4829;
  assign n5141 = po31  & n5140;
  assign n5142 = ~n4834 & ~n5141;
  assign n5143 = n4834 & n5141;
  assign n5144 = ~n5142 & ~n5143;
  assign n5145 = ~n5139 & ~n5144;
  assign n5146 = ~n5138 & ~n5145;
  assign n5147 = po41  & ~n5146;
  assign n5148 = ~po41  & n5146;
  assign n5149 = ~n4837 & ~n4838;
  assign n5150 = po31  & n5149;
  assign n5151 = ~n4843 & ~n5150;
  assign n5152 = n4843 & n5150;
  assign n5153 = ~n5151 & ~n5152;
  assign n5154 = ~n5148 & ~n5153;
  assign n5155 = ~n5147 & ~n5154;
  assign n5156 = po42  & ~n5155;
  assign n5157 = ~po42  & n5155;
  assign n5158 = ~n4846 & ~n4847;
  assign n5159 = po31  & n5158;
  assign n5160 = ~n4852 & ~n5159;
  assign n5161 = n4852 & n5159;
  assign n5162 = ~n5160 & ~n5161;
  assign n5163 = ~n5157 & ~n5162;
  assign n5164 = ~n5156 & ~n5163;
  assign n5165 = po43  & ~n5164;
  assign n5166 = ~po43  & n5164;
  assign n5167 = ~n4855 & ~n4856;
  assign n5168 = po31  & n5167;
  assign n5169 = ~n4861 & ~n5168;
  assign n5170 = n4861 & n5168;
  assign n5171 = ~n5169 & ~n5170;
  assign n5172 = ~n5166 & ~n5171;
  assign n5173 = ~n5165 & ~n5172;
  assign n5174 = po44  & ~n5173;
  assign n5175 = ~po44  & n5173;
  assign n5176 = ~n4864 & ~n4865;
  assign n5177 = po31  & n5176;
  assign n5178 = ~n4870 & ~n5177;
  assign n5179 = n4870 & n5177;
  assign n5180 = ~n5178 & ~n5179;
  assign n5181 = ~n5175 & ~n5180;
  assign n5182 = ~n5174 & ~n5181;
  assign n5183 = po45  & ~n5182;
  assign n5184 = ~po45  & n5182;
  assign n5185 = ~n4873 & ~n4874;
  assign n5186 = po31  & n5185;
  assign n5187 = ~n4879 & ~n5186;
  assign n5188 = n4879 & n5186;
  assign n5189 = ~n5187 & ~n5188;
  assign n5190 = ~n5184 & ~n5189;
  assign n5191 = ~n5183 & ~n5190;
  assign n5192 = po46  & ~n5191;
  assign n5193 = ~po46  & n5191;
  assign n5194 = ~n4882 & ~n4883;
  assign n5195 = po31  & n5194;
  assign n5196 = ~n4888 & ~n5195;
  assign n5197 = n4888 & n5195;
  assign n5198 = ~n5196 & ~n5197;
  assign n5199 = ~n5193 & ~n5198;
  assign n5200 = ~n5192 & ~n5199;
  assign n5201 = po47  & ~n5200;
  assign n5202 = ~po47  & n5200;
  assign n5203 = ~n4891 & ~n4892;
  assign n5204 = po31  & n5203;
  assign n5205 = ~n4897 & ~n5204;
  assign n5206 = n4897 & n5204;
  assign n5207 = ~n5205 & ~n5206;
  assign n5208 = ~n5202 & ~n5207;
  assign n5209 = ~n5201 & ~n5208;
  assign n5210 = po48  & ~n5209;
  assign n5211 = ~po48  & n5209;
  assign n5212 = ~n4900 & ~n4901;
  assign n5213 = po31  & n5212;
  assign n5214 = ~n4906 & ~n5213;
  assign n5215 = n4906 & n5213;
  assign n5216 = ~n5214 & ~n5215;
  assign n5217 = ~n5211 & ~n5216;
  assign n5218 = ~n5210 & ~n5217;
  assign n5219 = po49  & ~n5218;
  assign n5220 = ~po49  & n5218;
  assign n5221 = ~n4909 & ~n4910;
  assign n5222 = po31  & n5221;
  assign n5223 = ~n4915 & ~n5222;
  assign n5224 = n4915 & n5222;
  assign n5225 = ~n5223 & ~n5224;
  assign n5226 = ~n5220 & ~n5225;
  assign n5227 = ~n5219 & ~n5226;
  assign n5228 = po50  & ~n5227;
  assign n5229 = ~po50  & n5227;
  assign n5230 = ~n4918 & ~n4919;
  assign n5231 = po31  & n5230;
  assign n5232 = ~n4924 & ~n5231;
  assign n5233 = n4924 & n5231;
  assign n5234 = ~n5232 & ~n5233;
  assign n5235 = ~n5229 & ~n5234;
  assign n5236 = ~n5228 & ~n5235;
  assign n5237 = po51  & ~n5236;
  assign n5238 = ~po51  & n5236;
  assign n5239 = ~n4927 & ~n4928;
  assign n5240 = po31  & n5239;
  assign n5241 = ~n4933 & ~n5240;
  assign n5242 = n4933 & n5240;
  assign n5243 = ~n5241 & ~n5242;
  assign n5244 = ~n5238 & ~n5243;
  assign n5245 = ~n5237 & ~n5244;
  assign n5246 = po52  & ~n5245;
  assign n5247 = ~po52  & n5245;
  assign n5248 = ~n4936 & ~n4937;
  assign n5249 = po31  & n5248;
  assign n5250 = ~n4942 & ~n5249;
  assign n5251 = n4942 & n5249;
  assign n5252 = ~n5250 & ~n5251;
  assign n5253 = ~n5247 & ~n5252;
  assign n5254 = ~n5246 & ~n5253;
  assign n5255 = po53  & ~n5254;
  assign n5256 = ~po53  & n5254;
  assign n5257 = ~n4945 & ~n4946;
  assign n5258 = po31  & n5257;
  assign n5259 = ~n4951 & ~n5258;
  assign n5260 = n4951 & n5258;
  assign n5261 = ~n5259 & ~n5260;
  assign n5262 = ~n5256 & ~n5261;
  assign n5263 = ~n5255 & ~n5262;
  assign n5264 = po54  & ~n5263;
  assign n5265 = ~po54  & n5263;
  assign n5266 = ~n4954 & ~n4955;
  assign n5267 = po31  & n5266;
  assign n5268 = ~n4960 & ~n5267;
  assign n5269 = n4960 & n5267;
  assign n5270 = ~n5268 & ~n5269;
  assign n5271 = ~n5265 & ~n5270;
  assign n5272 = ~n5264 & ~n5271;
  assign n5273 = po55  & ~n5272;
  assign n5274 = ~po55  & n5272;
  assign n5275 = ~n4963 & ~n4964;
  assign n5276 = po31  & n5275;
  assign n5277 = ~n4969 & ~n5276;
  assign n5278 = n4969 & n5276;
  assign n5279 = ~n5277 & ~n5278;
  assign n5280 = ~n5274 & ~n5279;
  assign n5281 = ~n5273 & ~n5280;
  assign n5282 = po56  & ~n5281;
  assign n5283 = ~po56  & n5281;
  assign n5284 = ~n4972 & ~n4973;
  assign n5285 = po31  & n5284;
  assign n5286 = ~n4978 & ~n5285;
  assign n5287 = n4978 & n5285;
  assign n5288 = ~n5286 & ~n5287;
  assign n5289 = ~n5283 & ~n5288;
  assign n5290 = ~n5282 & ~n5289;
  assign n5291 = po57  & ~n5290;
  assign n5292 = ~po57  & n5290;
  assign n5293 = ~n4981 & ~n4982;
  assign n5294 = po31  & n5293;
  assign n5295 = ~n4987 & ~n5294;
  assign n5296 = n4987 & n5294;
  assign n5297 = ~n5295 & ~n5296;
  assign n5298 = ~n5292 & ~n5297;
  assign n5299 = ~n5291 & ~n5298;
  assign n5300 = po58  & ~n5299;
  assign n5301 = ~po58  & n5299;
  assign n5302 = ~n4990 & ~n4991;
  assign n5303 = po31  & n5302;
  assign n5304 = ~n4996 & ~n5303;
  assign n5305 = n4996 & n5303;
  assign n5306 = ~n5304 & ~n5305;
  assign n5307 = ~n5301 & ~n5306;
  assign n5308 = ~n5300 & ~n5307;
  assign n5309 = po59  & ~n5308;
  assign n5310 = ~po59  & n5308;
  assign n5311 = ~n4999 & ~n5000;
  assign n5312 = po31  & n5311;
  assign n5313 = ~n5005 & ~n5312;
  assign n5314 = n5005 & n5312;
  assign n5315 = ~n5313 & ~n5314;
  assign n5316 = ~n5310 & ~n5315;
  assign n5317 = ~n5309 & ~n5316;
  assign n5318 = po60  & ~n5317;
  assign n5319 = ~po60  & n5317;
  assign n5320 = ~n5008 & ~n5009;
  assign n5321 = po31  & n5320;
  assign n5322 = ~n5014 & ~n5321;
  assign n5323 = n5014 & n5321;
  assign n5324 = ~n5322 & ~n5323;
  assign n5325 = ~n5319 & ~n5324;
  assign n5326 = ~n5318 & ~n5325;
  assign n5327 = po61  & ~n5326;
  assign n5328 = ~po61  & n5326;
  assign n5329 = ~n5017 & ~n5018;
  assign n5330 = po31  & n5329;
  assign n5331 = ~n5023 & ~n5330;
  assign n5332 = n5023 & n5330;
  assign n5333 = ~n5331 & ~n5332;
  assign n5334 = ~n5328 & ~n5333;
  assign n5335 = ~n5327 & ~n5334;
  assign n5336 = po62  & ~n5335;
  assign n5337 = ~po62  & n5335;
  assign n5338 = ~n5026 & ~n5027;
  assign n5339 = po31  & n5338;
  assign n5340 = ~n5032 & ~n5339;
  assign n5341 = n5032 & n5339;
  assign n5342 = ~n5340 & ~n5341;
  assign n5343 = ~n5337 & ~n5342;
  assign n5344 = ~n5336 & ~n5343;
  assign n5345 = n5081 & n5344;
  assign n5346 = ~n5081 & ~n5344;
  assign n5347 = n5045 & po31 ;
  assign n5348 = ~n5044 & ~n5347;
  assign n5349 = n5346 & n5348;
  assign n5350 = ~po63  & ~n5349;
  assign n5351 = ~n4770 & po31 ;
  assign n5352 = n5043 & ~n5351;
  assign n5353 = po63  & ~n5045;
  assign n5354 = ~n5352 & n5353;
  assign n5355 = ~n5345 & ~n5354;
  assign n5356 = ~n5350 & n5355;
  assign po30  = n5076 | ~n5356;
  assign n5358 = ~n5074 & ~n5075;
  assign n5359 = po30  & n5358;
  assign n5360 = ~n5063 & ~n5359;
  assign n5361 = n5063 & n5359;
  assign n5362 = ~n5360 & ~n5361;
  assign n5363 = pi60  & po30 ;
  assign n5364 = ~pi58  & ~pi59 ;
  assign n5365 = ~pi60  & n5364;
  assign n5366 = ~n5363 & ~n5365;
  assign n5367 = po31  & ~n5366;
  assign n5368 = ~po31  & n5366;
  assign n5369 = ~pi60  & po30 ;
  assign n5370 = pi61  & ~n5369;
  assign n5371 = ~pi61  & n5369;
  assign n5372 = ~n5370 & ~n5371;
  assign n5373 = ~n5368 & n5372;
  assign n5374 = ~n5367 & ~n5373;
  assign n5375 = po32  & ~n5374;
  assign n5376 = ~po32  & n5374;
  assign n5377 = po31  & n5356;
  assign n5378 = ~n5371 & ~n5377;
  assign n5379 = pi62  & ~n5378;
  assign n5380 = ~pi62  & n5378;
  assign n5381 = ~n5379 & ~n5380;
  assign n5382 = ~n5376 & ~n5381;
  assign n5383 = ~n5375 & ~n5382;
  assign n5384 = po33  & ~n5383;
  assign n5385 = ~po33  & n5383;
  assign n5386 = ~n5068 & ~n5071;
  assign n5387 = po30  & n5386;
  assign n5388 = n5070 & ~n5387;
  assign n5389 = ~n5070 & n5387;
  assign n5390 = ~n5388 & ~n5389;
  assign n5391 = ~n5385 & ~n5390;
  assign n5392 = ~n5384 & ~n5391;
  assign n5393 = po34  & ~n5392;
  assign n5394 = ~po34  & n5392;
  assign n5395 = n5081 & ~po30 ;
  assign n5396 = ~n5336 & ~n5337;
  assign n5397 = po30  & n5396;
  assign n5398 = ~n5342 & ~n5397;
  assign n5399 = n5342 & n5397;
  assign n5400 = ~n5398 & ~n5399;
  assign n5401 = ~n5362 & ~n5394;
  assign n5402 = ~n5393 & ~n5401;
  assign n5403 = po35  & ~n5402;
  assign n5404 = ~po35  & n5402;
  assign n5405 = ~n5084 & ~n5085;
  assign n5406 = po30  & n5405;
  assign n5407 = n5090 & n5406;
  assign n5408 = ~n5090 & ~n5406;
  assign n5409 = ~n5407 & ~n5408;
  assign n5410 = ~n5404 & ~n5409;
  assign n5411 = ~n5403 & ~n5410;
  assign n5412 = po36  & ~n5411;
  assign n5413 = ~po36  & n5411;
  assign n5414 = ~n5093 & ~n5094;
  assign n5415 = po30  & n5414;
  assign n5416 = ~n5099 & ~n5415;
  assign n5417 = n5099 & n5415;
  assign n5418 = ~n5416 & ~n5417;
  assign n5419 = ~n5413 & ~n5418;
  assign n5420 = ~n5412 & ~n5419;
  assign n5421 = po37  & ~n5420;
  assign n5422 = ~po37  & n5420;
  assign n5423 = ~n5102 & ~n5103;
  assign n5424 = po30  & n5423;
  assign n5425 = ~n5108 & ~n5424;
  assign n5426 = n5108 & n5424;
  assign n5427 = ~n5425 & ~n5426;
  assign n5428 = ~n5422 & ~n5427;
  assign n5429 = ~n5421 & ~n5428;
  assign n5430 = po38  & ~n5429;
  assign n5431 = ~po38  & n5429;
  assign n5432 = ~n5111 & ~n5112;
  assign n5433 = po30  & n5432;
  assign n5434 = ~n5117 & ~n5433;
  assign n5435 = n5117 & n5433;
  assign n5436 = ~n5434 & ~n5435;
  assign n5437 = ~n5431 & ~n5436;
  assign n5438 = ~n5430 & ~n5437;
  assign n5439 = po39  & ~n5438;
  assign n5440 = ~po39  & n5438;
  assign n5441 = ~n5120 & ~n5121;
  assign n5442 = po30  & n5441;
  assign n5443 = ~n5126 & ~n5442;
  assign n5444 = n5126 & n5442;
  assign n5445 = ~n5443 & ~n5444;
  assign n5446 = ~n5440 & ~n5445;
  assign n5447 = ~n5439 & ~n5446;
  assign n5448 = po40  & ~n5447;
  assign n5449 = ~po40  & n5447;
  assign n5450 = ~n5129 & ~n5130;
  assign n5451 = po30  & n5450;
  assign n5452 = ~n5135 & ~n5451;
  assign n5453 = n5135 & n5451;
  assign n5454 = ~n5452 & ~n5453;
  assign n5455 = ~n5449 & ~n5454;
  assign n5456 = ~n5448 & ~n5455;
  assign n5457 = po41  & ~n5456;
  assign n5458 = ~po41  & n5456;
  assign n5459 = ~n5138 & ~n5139;
  assign n5460 = po30  & n5459;
  assign n5461 = ~n5144 & ~n5460;
  assign n5462 = n5144 & n5460;
  assign n5463 = ~n5461 & ~n5462;
  assign n5464 = ~n5458 & ~n5463;
  assign n5465 = ~n5457 & ~n5464;
  assign n5466 = po42  & ~n5465;
  assign n5467 = ~po42  & n5465;
  assign n5468 = ~n5147 & ~n5148;
  assign n5469 = po30  & n5468;
  assign n5470 = ~n5153 & ~n5469;
  assign n5471 = n5153 & n5469;
  assign n5472 = ~n5470 & ~n5471;
  assign n5473 = ~n5467 & ~n5472;
  assign n5474 = ~n5466 & ~n5473;
  assign n5475 = po43  & ~n5474;
  assign n5476 = ~po43  & n5474;
  assign n5477 = ~n5156 & ~n5157;
  assign n5478 = po30  & n5477;
  assign n5479 = ~n5162 & ~n5478;
  assign n5480 = n5162 & n5478;
  assign n5481 = ~n5479 & ~n5480;
  assign n5482 = ~n5476 & ~n5481;
  assign n5483 = ~n5475 & ~n5482;
  assign n5484 = po44  & ~n5483;
  assign n5485 = ~po44  & n5483;
  assign n5486 = ~n5165 & ~n5166;
  assign n5487 = po30  & n5486;
  assign n5488 = ~n5171 & ~n5487;
  assign n5489 = n5171 & n5487;
  assign n5490 = ~n5488 & ~n5489;
  assign n5491 = ~n5485 & ~n5490;
  assign n5492 = ~n5484 & ~n5491;
  assign n5493 = po45  & ~n5492;
  assign n5494 = ~po45  & n5492;
  assign n5495 = ~n5174 & ~n5175;
  assign n5496 = po30  & n5495;
  assign n5497 = ~n5180 & ~n5496;
  assign n5498 = n5180 & n5496;
  assign n5499 = ~n5497 & ~n5498;
  assign n5500 = ~n5494 & ~n5499;
  assign n5501 = ~n5493 & ~n5500;
  assign n5502 = po46  & ~n5501;
  assign n5503 = ~po46  & n5501;
  assign n5504 = ~n5183 & ~n5184;
  assign n5505 = po30  & n5504;
  assign n5506 = ~n5189 & ~n5505;
  assign n5507 = n5189 & n5505;
  assign n5508 = ~n5506 & ~n5507;
  assign n5509 = ~n5503 & ~n5508;
  assign n5510 = ~n5502 & ~n5509;
  assign n5511 = po47  & ~n5510;
  assign n5512 = ~po47  & n5510;
  assign n5513 = ~n5192 & ~n5193;
  assign n5514 = po30  & n5513;
  assign n5515 = ~n5198 & ~n5514;
  assign n5516 = n5198 & n5514;
  assign n5517 = ~n5515 & ~n5516;
  assign n5518 = ~n5512 & ~n5517;
  assign n5519 = ~n5511 & ~n5518;
  assign n5520 = po48  & ~n5519;
  assign n5521 = ~po48  & n5519;
  assign n5522 = ~n5201 & ~n5202;
  assign n5523 = po30  & n5522;
  assign n5524 = ~n5207 & ~n5523;
  assign n5525 = n5207 & n5523;
  assign n5526 = ~n5524 & ~n5525;
  assign n5527 = ~n5521 & ~n5526;
  assign n5528 = ~n5520 & ~n5527;
  assign n5529 = po49  & ~n5528;
  assign n5530 = ~po49  & n5528;
  assign n5531 = ~n5210 & ~n5211;
  assign n5532 = po30  & n5531;
  assign n5533 = ~n5216 & ~n5532;
  assign n5534 = n5216 & n5532;
  assign n5535 = ~n5533 & ~n5534;
  assign n5536 = ~n5530 & ~n5535;
  assign n5537 = ~n5529 & ~n5536;
  assign n5538 = po50  & ~n5537;
  assign n5539 = ~po50  & n5537;
  assign n5540 = ~n5219 & ~n5220;
  assign n5541 = po30  & n5540;
  assign n5542 = ~n5225 & ~n5541;
  assign n5543 = n5225 & n5541;
  assign n5544 = ~n5542 & ~n5543;
  assign n5545 = ~n5539 & ~n5544;
  assign n5546 = ~n5538 & ~n5545;
  assign n5547 = po51  & ~n5546;
  assign n5548 = ~po51  & n5546;
  assign n5549 = ~n5228 & ~n5229;
  assign n5550 = po30  & n5549;
  assign n5551 = ~n5234 & ~n5550;
  assign n5552 = n5234 & n5550;
  assign n5553 = ~n5551 & ~n5552;
  assign n5554 = ~n5548 & ~n5553;
  assign n5555 = ~n5547 & ~n5554;
  assign n5556 = po52  & ~n5555;
  assign n5557 = ~po52  & n5555;
  assign n5558 = ~n5237 & ~n5238;
  assign n5559 = po30  & n5558;
  assign n5560 = ~n5243 & ~n5559;
  assign n5561 = n5243 & n5559;
  assign n5562 = ~n5560 & ~n5561;
  assign n5563 = ~n5557 & ~n5562;
  assign n5564 = ~n5556 & ~n5563;
  assign n5565 = po53  & ~n5564;
  assign n5566 = ~po53  & n5564;
  assign n5567 = ~n5246 & ~n5247;
  assign n5568 = po30  & n5567;
  assign n5569 = ~n5252 & ~n5568;
  assign n5570 = n5252 & n5568;
  assign n5571 = ~n5569 & ~n5570;
  assign n5572 = ~n5566 & ~n5571;
  assign n5573 = ~n5565 & ~n5572;
  assign n5574 = po54  & ~n5573;
  assign n5575 = ~po54  & n5573;
  assign n5576 = ~n5255 & ~n5256;
  assign n5577 = po30  & n5576;
  assign n5578 = ~n5261 & ~n5577;
  assign n5579 = n5261 & n5577;
  assign n5580 = ~n5578 & ~n5579;
  assign n5581 = ~n5575 & ~n5580;
  assign n5582 = ~n5574 & ~n5581;
  assign n5583 = po55  & ~n5582;
  assign n5584 = ~po55  & n5582;
  assign n5585 = ~n5264 & ~n5265;
  assign n5586 = po30  & n5585;
  assign n5587 = ~n5270 & ~n5586;
  assign n5588 = n5270 & n5586;
  assign n5589 = ~n5587 & ~n5588;
  assign n5590 = ~n5584 & ~n5589;
  assign n5591 = ~n5583 & ~n5590;
  assign n5592 = po56  & ~n5591;
  assign n5593 = ~po56  & n5591;
  assign n5594 = ~n5273 & ~n5274;
  assign n5595 = po30  & n5594;
  assign n5596 = ~n5279 & ~n5595;
  assign n5597 = n5279 & n5595;
  assign n5598 = ~n5596 & ~n5597;
  assign n5599 = ~n5593 & ~n5598;
  assign n5600 = ~n5592 & ~n5599;
  assign n5601 = po57  & ~n5600;
  assign n5602 = ~po57  & n5600;
  assign n5603 = ~n5282 & ~n5283;
  assign n5604 = po30  & n5603;
  assign n5605 = ~n5288 & ~n5604;
  assign n5606 = n5288 & n5604;
  assign n5607 = ~n5605 & ~n5606;
  assign n5608 = ~n5602 & ~n5607;
  assign n5609 = ~n5601 & ~n5608;
  assign n5610 = po58  & ~n5609;
  assign n5611 = ~po58  & n5609;
  assign n5612 = ~n5291 & ~n5292;
  assign n5613 = po30  & n5612;
  assign n5614 = ~n5297 & ~n5613;
  assign n5615 = n5297 & n5613;
  assign n5616 = ~n5614 & ~n5615;
  assign n5617 = ~n5611 & ~n5616;
  assign n5618 = ~n5610 & ~n5617;
  assign n5619 = po59  & ~n5618;
  assign n5620 = ~po59  & n5618;
  assign n5621 = ~n5300 & ~n5301;
  assign n5622 = po30  & n5621;
  assign n5623 = ~n5306 & ~n5622;
  assign n5624 = n5306 & n5622;
  assign n5625 = ~n5623 & ~n5624;
  assign n5626 = ~n5620 & ~n5625;
  assign n5627 = ~n5619 & ~n5626;
  assign n5628 = po60  & ~n5627;
  assign n5629 = ~po60  & n5627;
  assign n5630 = ~n5309 & ~n5310;
  assign n5631 = po30  & n5630;
  assign n5632 = ~n5315 & ~n5631;
  assign n5633 = n5315 & n5631;
  assign n5634 = ~n5632 & ~n5633;
  assign n5635 = ~n5629 & ~n5634;
  assign n5636 = ~n5628 & ~n5635;
  assign n5637 = po61  & ~n5636;
  assign n5638 = ~po61  & n5636;
  assign n5639 = ~n5318 & ~n5319;
  assign n5640 = po30  & n5639;
  assign n5641 = ~n5324 & ~n5640;
  assign n5642 = n5324 & n5640;
  assign n5643 = ~n5641 & ~n5642;
  assign n5644 = ~n5638 & ~n5643;
  assign n5645 = ~n5637 & ~n5644;
  assign n5646 = po62  & ~n5645;
  assign n5647 = ~po62  & n5645;
  assign n5648 = ~n5327 & ~n5328;
  assign n5649 = po30  & n5648;
  assign n5650 = ~n5333 & ~n5649;
  assign n5651 = n5333 & n5649;
  assign n5652 = ~n5650 & ~n5651;
  assign n5653 = ~n5647 & ~n5652;
  assign n5654 = ~n5646 & ~n5653;
  assign n5655 = n5400 & n5654;
  assign n5656 = ~n5400 & ~n5654;
  assign n5657 = n5346 & po30 ;
  assign n5658 = ~n5345 & ~n5657;
  assign n5659 = n5656 & n5658;
  assign n5660 = ~po63  & ~n5659;
  assign n5661 = ~n5081 & po30 ;
  assign n5662 = n5344 & ~n5661;
  assign n5663 = po63  & ~n5346;
  assign n5664 = ~n5662 & n5663;
  assign n5665 = ~n5655 & ~n5664;
  assign n5666 = ~n5660 & n5665;
  assign po29  = n5395 | ~n5666;
  assign n5668 = ~n5393 & ~n5394;
  assign n5669 = po29  & n5668;
  assign n5670 = ~n5362 & ~n5669;
  assign n5671 = n5362 & n5669;
  assign n5672 = ~n5670 & ~n5671;
  assign n5673 = pi58  & po29 ;
  assign n5674 = ~pi56  & ~pi57 ;
  assign n5675 = ~pi58  & n5674;
  assign n5676 = ~n5673 & ~n5675;
  assign n5677 = po30  & ~n5676;
  assign n5678 = ~po30  & n5676;
  assign n5679 = ~pi58  & po29 ;
  assign n5680 = pi59  & ~n5679;
  assign n5681 = ~pi59  & n5679;
  assign n5682 = ~n5680 & ~n5681;
  assign n5683 = ~n5678 & n5682;
  assign n5684 = ~n5677 & ~n5683;
  assign n5685 = po31  & ~n5684;
  assign n5686 = ~po31  & n5684;
  assign n5687 = po30  & n5666;
  assign n5688 = ~n5681 & ~n5687;
  assign n5689 = pi60  & ~n5688;
  assign n5690 = ~pi60  & n5688;
  assign n5691 = ~n5689 & ~n5690;
  assign n5692 = ~n5686 & ~n5691;
  assign n5693 = ~n5685 & ~n5692;
  assign n5694 = po32  & ~n5693;
  assign n5695 = ~po32  & n5693;
  assign n5696 = ~n5367 & ~n5368;
  assign n5697 = po29  & n5696;
  assign n5698 = n5372 & ~n5697;
  assign n5699 = ~n5372 & n5697;
  assign n5700 = ~n5698 & ~n5699;
  assign n5701 = ~n5695 & ~n5700;
  assign n5702 = ~n5694 & ~n5701;
  assign n5703 = po33  & ~n5702;
  assign n5704 = ~po33  & n5702;
  assign n5705 = ~n5375 & ~n5376;
  assign n5706 = po29  & n5705;
  assign n5707 = ~n5381 & ~n5706;
  assign n5708 = n5381 & n5706;
  assign n5709 = ~n5707 & ~n5708;
  assign n5710 = ~n5704 & ~n5709;
  assign n5711 = ~n5703 & ~n5710;
  assign n5712 = po34  & ~n5711;
  assign n5713 = ~po34  & n5711;
  assign n5714 = ~n5384 & ~n5385;
  assign n5715 = po29  & n5714;
  assign n5716 = n5390 & n5715;
  assign n5717 = ~n5390 & ~n5715;
  assign n5718 = ~n5716 & ~n5717;
  assign n5719 = ~n5713 & ~n5718;
  assign n5720 = ~n5712 & ~n5719;
  assign n5721 = po35  & ~n5720;
  assign n5722 = ~po35  & n5720;
  assign n5723 = n5400 & ~po29 ;
  assign n5724 = ~n5646 & ~n5647;
  assign n5725 = po29  & n5724;
  assign n5726 = ~n5652 & ~n5725;
  assign n5727 = n5652 & n5725;
  assign n5728 = ~n5726 & ~n5727;
  assign n5729 = ~n5672 & ~n5722;
  assign n5730 = ~n5721 & ~n5729;
  assign n5731 = po36  & ~n5730;
  assign n5732 = ~po36  & n5730;
  assign n5733 = ~n5403 & ~n5404;
  assign n5734 = po29  & n5733;
  assign n5735 = ~n5409 & ~n5734;
  assign n5736 = n5409 & n5734;
  assign n5737 = ~n5735 & ~n5736;
  assign n5738 = ~n5732 & ~n5737;
  assign n5739 = ~n5731 & ~n5738;
  assign n5740 = po37  & ~n5739;
  assign n5741 = ~po37  & n5739;
  assign n5742 = ~n5412 & ~n5413;
  assign n5743 = po29  & n5742;
  assign n5744 = ~n5418 & ~n5743;
  assign n5745 = n5418 & n5743;
  assign n5746 = ~n5744 & ~n5745;
  assign n5747 = ~n5741 & ~n5746;
  assign n5748 = ~n5740 & ~n5747;
  assign n5749 = po38  & ~n5748;
  assign n5750 = ~po38  & n5748;
  assign n5751 = ~n5421 & ~n5422;
  assign n5752 = po29  & n5751;
  assign n5753 = ~n5427 & ~n5752;
  assign n5754 = n5427 & n5752;
  assign n5755 = ~n5753 & ~n5754;
  assign n5756 = ~n5750 & ~n5755;
  assign n5757 = ~n5749 & ~n5756;
  assign n5758 = po39  & ~n5757;
  assign n5759 = ~po39  & n5757;
  assign n5760 = ~n5430 & ~n5431;
  assign n5761 = po29  & n5760;
  assign n5762 = ~n5436 & ~n5761;
  assign n5763 = n5436 & n5761;
  assign n5764 = ~n5762 & ~n5763;
  assign n5765 = ~n5759 & ~n5764;
  assign n5766 = ~n5758 & ~n5765;
  assign n5767 = po40  & ~n5766;
  assign n5768 = ~po40  & n5766;
  assign n5769 = ~n5439 & ~n5440;
  assign n5770 = po29  & n5769;
  assign n5771 = ~n5445 & ~n5770;
  assign n5772 = n5445 & n5770;
  assign n5773 = ~n5771 & ~n5772;
  assign n5774 = ~n5768 & ~n5773;
  assign n5775 = ~n5767 & ~n5774;
  assign n5776 = po41  & ~n5775;
  assign n5777 = ~po41  & n5775;
  assign n5778 = ~n5448 & ~n5449;
  assign n5779 = po29  & n5778;
  assign n5780 = ~n5454 & ~n5779;
  assign n5781 = n5454 & n5779;
  assign n5782 = ~n5780 & ~n5781;
  assign n5783 = ~n5777 & ~n5782;
  assign n5784 = ~n5776 & ~n5783;
  assign n5785 = po42  & ~n5784;
  assign n5786 = ~po42  & n5784;
  assign n5787 = ~n5457 & ~n5458;
  assign n5788 = po29  & n5787;
  assign n5789 = ~n5463 & ~n5788;
  assign n5790 = n5463 & n5788;
  assign n5791 = ~n5789 & ~n5790;
  assign n5792 = ~n5786 & ~n5791;
  assign n5793 = ~n5785 & ~n5792;
  assign n5794 = po43  & ~n5793;
  assign n5795 = ~po43  & n5793;
  assign n5796 = ~n5466 & ~n5467;
  assign n5797 = po29  & n5796;
  assign n5798 = ~n5472 & ~n5797;
  assign n5799 = n5472 & n5797;
  assign n5800 = ~n5798 & ~n5799;
  assign n5801 = ~n5795 & ~n5800;
  assign n5802 = ~n5794 & ~n5801;
  assign n5803 = po44  & ~n5802;
  assign n5804 = ~po44  & n5802;
  assign n5805 = ~n5475 & ~n5476;
  assign n5806 = po29  & n5805;
  assign n5807 = ~n5481 & ~n5806;
  assign n5808 = n5481 & n5806;
  assign n5809 = ~n5807 & ~n5808;
  assign n5810 = ~n5804 & ~n5809;
  assign n5811 = ~n5803 & ~n5810;
  assign n5812 = po45  & ~n5811;
  assign n5813 = ~po45  & n5811;
  assign n5814 = ~n5484 & ~n5485;
  assign n5815 = po29  & n5814;
  assign n5816 = ~n5490 & ~n5815;
  assign n5817 = n5490 & n5815;
  assign n5818 = ~n5816 & ~n5817;
  assign n5819 = ~n5813 & ~n5818;
  assign n5820 = ~n5812 & ~n5819;
  assign n5821 = po46  & ~n5820;
  assign n5822 = ~po46  & n5820;
  assign n5823 = ~n5493 & ~n5494;
  assign n5824 = po29  & n5823;
  assign n5825 = ~n5499 & ~n5824;
  assign n5826 = n5499 & n5824;
  assign n5827 = ~n5825 & ~n5826;
  assign n5828 = ~n5822 & ~n5827;
  assign n5829 = ~n5821 & ~n5828;
  assign n5830 = po47  & ~n5829;
  assign n5831 = ~po47  & n5829;
  assign n5832 = ~n5502 & ~n5503;
  assign n5833 = po29  & n5832;
  assign n5834 = ~n5508 & ~n5833;
  assign n5835 = n5508 & n5833;
  assign n5836 = ~n5834 & ~n5835;
  assign n5837 = ~n5831 & ~n5836;
  assign n5838 = ~n5830 & ~n5837;
  assign n5839 = po48  & ~n5838;
  assign n5840 = ~po48  & n5838;
  assign n5841 = ~n5511 & ~n5512;
  assign n5842 = po29  & n5841;
  assign n5843 = ~n5517 & ~n5842;
  assign n5844 = n5517 & n5842;
  assign n5845 = ~n5843 & ~n5844;
  assign n5846 = ~n5840 & ~n5845;
  assign n5847 = ~n5839 & ~n5846;
  assign n5848 = po49  & ~n5847;
  assign n5849 = ~po49  & n5847;
  assign n5850 = ~n5520 & ~n5521;
  assign n5851 = po29  & n5850;
  assign n5852 = ~n5526 & ~n5851;
  assign n5853 = n5526 & n5851;
  assign n5854 = ~n5852 & ~n5853;
  assign n5855 = ~n5849 & ~n5854;
  assign n5856 = ~n5848 & ~n5855;
  assign n5857 = po50  & ~n5856;
  assign n5858 = ~po50  & n5856;
  assign n5859 = ~n5529 & ~n5530;
  assign n5860 = po29  & n5859;
  assign n5861 = ~n5535 & ~n5860;
  assign n5862 = n5535 & n5860;
  assign n5863 = ~n5861 & ~n5862;
  assign n5864 = ~n5858 & ~n5863;
  assign n5865 = ~n5857 & ~n5864;
  assign n5866 = po51  & ~n5865;
  assign n5867 = ~po51  & n5865;
  assign n5868 = ~n5538 & ~n5539;
  assign n5869 = po29  & n5868;
  assign n5870 = ~n5544 & ~n5869;
  assign n5871 = n5544 & n5869;
  assign n5872 = ~n5870 & ~n5871;
  assign n5873 = ~n5867 & ~n5872;
  assign n5874 = ~n5866 & ~n5873;
  assign n5875 = po52  & ~n5874;
  assign n5876 = ~po52  & n5874;
  assign n5877 = ~n5547 & ~n5548;
  assign n5878 = po29  & n5877;
  assign n5879 = ~n5553 & ~n5878;
  assign n5880 = n5553 & n5878;
  assign n5881 = ~n5879 & ~n5880;
  assign n5882 = ~n5876 & ~n5881;
  assign n5883 = ~n5875 & ~n5882;
  assign n5884 = po53  & ~n5883;
  assign n5885 = ~po53  & n5883;
  assign n5886 = ~n5556 & ~n5557;
  assign n5887 = po29  & n5886;
  assign n5888 = ~n5562 & ~n5887;
  assign n5889 = n5562 & n5887;
  assign n5890 = ~n5888 & ~n5889;
  assign n5891 = ~n5885 & ~n5890;
  assign n5892 = ~n5884 & ~n5891;
  assign n5893 = po54  & ~n5892;
  assign n5894 = ~po54  & n5892;
  assign n5895 = ~n5565 & ~n5566;
  assign n5896 = po29  & n5895;
  assign n5897 = ~n5571 & ~n5896;
  assign n5898 = n5571 & n5896;
  assign n5899 = ~n5897 & ~n5898;
  assign n5900 = ~n5894 & ~n5899;
  assign n5901 = ~n5893 & ~n5900;
  assign n5902 = po55  & ~n5901;
  assign n5903 = ~po55  & n5901;
  assign n5904 = ~n5574 & ~n5575;
  assign n5905 = po29  & n5904;
  assign n5906 = ~n5580 & ~n5905;
  assign n5907 = n5580 & n5905;
  assign n5908 = ~n5906 & ~n5907;
  assign n5909 = ~n5903 & ~n5908;
  assign n5910 = ~n5902 & ~n5909;
  assign n5911 = po56  & ~n5910;
  assign n5912 = ~po56  & n5910;
  assign n5913 = ~n5583 & ~n5584;
  assign n5914 = po29  & n5913;
  assign n5915 = ~n5589 & ~n5914;
  assign n5916 = n5589 & n5914;
  assign n5917 = ~n5915 & ~n5916;
  assign n5918 = ~n5912 & ~n5917;
  assign n5919 = ~n5911 & ~n5918;
  assign n5920 = po57  & ~n5919;
  assign n5921 = ~po57  & n5919;
  assign n5922 = ~n5592 & ~n5593;
  assign n5923 = po29  & n5922;
  assign n5924 = ~n5598 & ~n5923;
  assign n5925 = n5598 & n5923;
  assign n5926 = ~n5924 & ~n5925;
  assign n5927 = ~n5921 & ~n5926;
  assign n5928 = ~n5920 & ~n5927;
  assign n5929 = po58  & ~n5928;
  assign n5930 = ~po58  & n5928;
  assign n5931 = ~n5601 & ~n5602;
  assign n5932 = po29  & n5931;
  assign n5933 = ~n5607 & ~n5932;
  assign n5934 = n5607 & n5932;
  assign n5935 = ~n5933 & ~n5934;
  assign n5936 = ~n5930 & ~n5935;
  assign n5937 = ~n5929 & ~n5936;
  assign n5938 = po59  & ~n5937;
  assign n5939 = ~po59  & n5937;
  assign n5940 = ~n5610 & ~n5611;
  assign n5941 = po29  & n5940;
  assign n5942 = ~n5616 & ~n5941;
  assign n5943 = n5616 & n5941;
  assign n5944 = ~n5942 & ~n5943;
  assign n5945 = ~n5939 & ~n5944;
  assign n5946 = ~n5938 & ~n5945;
  assign n5947 = po60  & ~n5946;
  assign n5948 = ~po60  & n5946;
  assign n5949 = ~n5619 & ~n5620;
  assign n5950 = po29  & n5949;
  assign n5951 = ~n5625 & ~n5950;
  assign n5952 = n5625 & n5950;
  assign n5953 = ~n5951 & ~n5952;
  assign n5954 = ~n5948 & ~n5953;
  assign n5955 = ~n5947 & ~n5954;
  assign n5956 = po61  & ~n5955;
  assign n5957 = ~po61  & n5955;
  assign n5958 = ~n5628 & ~n5629;
  assign n5959 = po29  & n5958;
  assign n5960 = ~n5634 & ~n5959;
  assign n5961 = n5634 & n5959;
  assign n5962 = ~n5960 & ~n5961;
  assign n5963 = ~n5957 & ~n5962;
  assign n5964 = ~n5956 & ~n5963;
  assign n5965 = po62  & ~n5964;
  assign n5966 = ~po62  & n5964;
  assign n5967 = ~n5637 & ~n5638;
  assign n5968 = po29  & n5967;
  assign n5969 = ~n5643 & ~n5968;
  assign n5970 = n5643 & n5968;
  assign n5971 = ~n5969 & ~n5970;
  assign n5972 = ~n5966 & ~n5971;
  assign n5973 = ~n5965 & ~n5972;
  assign n5974 = n5728 & n5973;
  assign n5975 = ~n5728 & ~n5973;
  assign n5976 = n5656 & po29 ;
  assign n5977 = ~n5655 & ~n5976;
  assign n5978 = n5975 & n5977;
  assign n5979 = ~po63  & ~n5978;
  assign n5980 = ~n5400 & po29 ;
  assign n5981 = n5654 & ~n5980;
  assign n5982 = po63  & ~n5656;
  assign n5983 = ~n5981 & n5982;
  assign n5984 = ~n5974 & ~n5983;
  assign n5985 = ~n5979 & n5984;
  assign po28  = n5723 | ~n5985;
  assign n5987 = ~n5721 & ~n5722;
  assign n5988 = po28  & n5987;
  assign n5989 = ~n5672 & ~n5988;
  assign n5990 = n5672 & n5988;
  assign n5991 = ~n5989 & ~n5990;
  assign n5992 = pi56  & po28 ;
  assign n5993 = ~pi54  & ~pi55 ;
  assign n5994 = ~pi56  & n5993;
  assign n5995 = ~n5992 & ~n5994;
  assign n5996 = po29  & ~n5995;
  assign n5997 = ~po29  & n5995;
  assign n5998 = ~pi56  & po28 ;
  assign n5999 = pi57  & ~n5998;
  assign n6000 = ~pi57  & n5998;
  assign n6001 = ~n5999 & ~n6000;
  assign n6002 = ~n5997 & n6001;
  assign n6003 = ~n5996 & ~n6002;
  assign n6004 = po30  & ~n6003;
  assign n6005 = ~po30  & n6003;
  assign n6006 = po29  & n5985;
  assign n6007 = ~n6000 & ~n6006;
  assign n6008 = pi58  & ~n6007;
  assign n6009 = ~pi58  & n6007;
  assign n6010 = ~n6008 & ~n6009;
  assign n6011 = ~n6005 & ~n6010;
  assign n6012 = ~n6004 & ~n6011;
  assign n6013 = po31  & ~n6012;
  assign n6014 = ~po31  & n6012;
  assign n6015 = ~n5677 & ~n5678;
  assign n6016 = po28  & n6015;
  assign n6017 = n5682 & ~n6016;
  assign n6018 = ~n5682 & n6016;
  assign n6019 = ~n6017 & ~n6018;
  assign n6020 = ~n6014 & ~n6019;
  assign n6021 = ~n6013 & ~n6020;
  assign n6022 = po32  & ~n6021;
  assign n6023 = ~po32  & n6021;
  assign n6024 = ~n5685 & ~n5686;
  assign n6025 = po28  & n6024;
  assign n6026 = ~n5691 & ~n6025;
  assign n6027 = n5691 & n6025;
  assign n6028 = ~n6026 & ~n6027;
  assign n6029 = ~n6023 & ~n6028;
  assign n6030 = ~n6022 & ~n6029;
  assign n6031 = po33  & ~n6030;
  assign n6032 = ~po33  & n6030;
  assign n6033 = ~n5694 & ~n5695;
  assign n6034 = po28  & n6033;
  assign n6035 = n5700 & n6034;
  assign n6036 = ~n5700 & ~n6034;
  assign n6037 = ~n6035 & ~n6036;
  assign n6038 = ~n6032 & ~n6037;
  assign n6039 = ~n6031 & ~n6038;
  assign n6040 = po34  & ~n6039;
  assign n6041 = ~po34  & n6039;
  assign n6042 = ~n5703 & ~n5704;
  assign n6043 = po28  & n6042;
  assign n6044 = ~n5709 & ~n6043;
  assign n6045 = n5709 & n6043;
  assign n6046 = ~n6044 & ~n6045;
  assign n6047 = ~n6041 & ~n6046;
  assign n6048 = ~n6040 & ~n6047;
  assign n6049 = po35  & ~n6048;
  assign n6050 = ~n5712 & ~n5713;
  assign n6051 = po28  & n6050;
  assign n6052 = ~n5718 & ~n6051;
  assign n6053 = n5718 & n6051;
  assign n6054 = ~n6052 & ~n6053;
  assign n6055 = ~po35  & n6048;
  assign n6056 = ~n6054 & ~n6055;
  assign n6057 = ~n6049 & ~n6056;
  assign n6058 = po36  & ~n6057;
  assign n6059 = ~po36  & n6057;
  assign n6060 = n5728 & ~po28 ;
  assign n6061 = ~n5965 & ~n5966;
  assign n6062 = po28  & n6061;
  assign n6063 = ~n5971 & ~n6062;
  assign n6064 = n5971 & n6062;
  assign n6065 = ~n6063 & ~n6064;
  assign n6066 = ~n5991 & ~n6059;
  assign n6067 = ~n6058 & ~n6066;
  assign n6068 = po37  & ~n6067;
  assign n6069 = ~po37  & n6067;
  assign n6070 = ~n5731 & ~n5732;
  assign n6071 = po28  & n6070;
  assign n6072 = ~n5737 & ~n6071;
  assign n6073 = n5737 & n6071;
  assign n6074 = ~n6072 & ~n6073;
  assign n6075 = ~n6069 & ~n6074;
  assign n6076 = ~n6068 & ~n6075;
  assign n6077 = po38  & ~n6076;
  assign n6078 = ~po38  & n6076;
  assign n6079 = ~n5740 & ~n5741;
  assign n6080 = po28  & n6079;
  assign n6081 = ~n5746 & ~n6080;
  assign n6082 = n5746 & n6080;
  assign n6083 = ~n6081 & ~n6082;
  assign n6084 = ~n6078 & ~n6083;
  assign n6085 = ~n6077 & ~n6084;
  assign n6086 = po39  & ~n6085;
  assign n6087 = ~po39  & n6085;
  assign n6088 = ~n5749 & ~n5750;
  assign n6089 = po28  & n6088;
  assign n6090 = ~n5755 & ~n6089;
  assign n6091 = n5755 & n6089;
  assign n6092 = ~n6090 & ~n6091;
  assign n6093 = ~n6087 & ~n6092;
  assign n6094 = ~n6086 & ~n6093;
  assign n6095 = po40  & ~n6094;
  assign n6096 = ~po40  & n6094;
  assign n6097 = ~n5758 & ~n5759;
  assign n6098 = po28  & n6097;
  assign n6099 = ~n5764 & ~n6098;
  assign n6100 = n5764 & n6098;
  assign n6101 = ~n6099 & ~n6100;
  assign n6102 = ~n6096 & ~n6101;
  assign n6103 = ~n6095 & ~n6102;
  assign n6104 = po41  & ~n6103;
  assign n6105 = ~po41  & n6103;
  assign n6106 = ~n5767 & ~n5768;
  assign n6107 = po28  & n6106;
  assign n6108 = ~n5773 & ~n6107;
  assign n6109 = n5773 & n6107;
  assign n6110 = ~n6108 & ~n6109;
  assign n6111 = ~n6105 & ~n6110;
  assign n6112 = ~n6104 & ~n6111;
  assign n6113 = po42  & ~n6112;
  assign n6114 = ~po42  & n6112;
  assign n6115 = ~n5776 & ~n5777;
  assign n6116 = po28  & n6115;
  assign n6117 = ~n5782 & ~n6116;
  assign n6118 = n5782 & n6116;
  assign n6119 = ~n6117 & ~n6118;
  assign n6120 = ~n6114 & ~n6119;
  assign n6121 = ~n6113 & ~n6120;
  assign n6122 = po43  & ~n6121;
  assign n6123 = ~po43  & n6121;
  assign n6124 = ~n5785 & ~n5786;
  assign n6125 = po28  & n6124;
  assign n6126 = ~n5791 & ~n6125;
  assign n6127 = n5791 & n6125;
  assign n6128 = ~n6126 & ~n6127;
  assign n6129 = ~n6123 & ~n6128;
  assign n6130 = ~n6122 & ~n6129;
  assign n6131 = po44  & ~n6130;
  assign n6132 = ~po44  & n6130;
  assign n6133 = ~n5794 & ~n5795;
  assign n6134 = po28  & n6133;
  assign n6135 = ~n5800 & ~n6134;
  assign n6136 = n5800 & n6134;
  assign n6137 = ~n6135 & ~n6136;
  assign n6138 = ~n6132 & ~n6137;
  assign n6139 = ~n6131 & ~n6138;
  assign n6140 = po45  & ~n6139;
  assign n6141 = ~po45  & n6139;
  assign n6142 = ~n5803 & ~n5804;
  assign n6143 = po28  & n6142;
  assign n6144 = ~n5809 & ~n6143;
  assign n6145 = n5809 & n6143;
  assign n6146 = ~n6144 & ~n6145;
  assign n6147 = ~n6141 & ~n6146;
  assign n6148 = ~n6140 & ~n6147;
  assign n6149 = po46  & ~n6148;
  assign n6150 = ~po46  & n6148;
  assign n6151 = ~n5812 & ~n5813;
  assign n6152 = po28  & n6151;
  assign n6153 = ~n5818 & ~n6152;
  assign n6154 = n5818 & n6152;
  assign n6155 = ~n6153 & ~n6154;
  assign n6156 = ~n6150 & ~n6155;
  assign n6157 = ~n6149 & ~n6156;
  assign n6158 = po47  & ~n6157;
  assign n6159 = ~po47  & n6157;
  assign n6160 = ~n5821 & ~n5822;
  assign n6161 = po28  & n6160;
  assign n6162 = ~n5827 & ~n6161;
  assign n6163 = n5827 & n6161;
  assign n6164 = ~n6162 & ~n6163;
  assign n6165 = ~n6159 & ~n6164;
  assign n6166 = ~n6158 & ~n6165;
  assign n6167 = po48  & ~n6166;
  assign n6168 = ~po48  & n6166;
  assign n6169 = ~n5830 & ~n5831;
  assign n6170 = po28  & n6169;
  assign n6171 = ~n5836 & ~n6170;
  assign n6172 = n5836 & n6170;
  assign n6173 = ~n6171 & ~n6172;
  assign n6174 = ~n6168 & ~n6173;
  assign n6175 = ~n6167 & ~n6174;
  assign n6176 = po49  & ~n6175;
  assign n6177 = ~po49  & n6175;
  assign n6178 = ~n5839 & ~n5840;
  assign n6179 = po28  & n6178;
  assign n6180 = ~n5845 & ~n6179;
  assign n6181 = n5845 & n6179;
  assign n6182 = ~n6180 & ~n6181;
  assign n6183 = ~n6177 & ~n6182;
  assign n6184 = ~n6176 & ~n6183;
  assign n6185 = po50  & ~n6184;
  assign n6186 = ~po50  & n6184;
  assign n6187 = ~n5848 & ~n5849;
  assign n6188 = po28  & n6187;
  assign n6189 = ~n5854 & ~n6188;
  assign n6190 = n5854 & n6188;
  assign n6191 = ~n6189 & ~n6190;
  assign n6192 = ~n6186 & ~n6191;
  assign n6193 = ~n6185 & ~n6192;
  assign n6194 = po51  & ~n6193;
  assign n6195 = ~po51  & n6193;
  assign n6196 = ~n5857 & ~n5858;
  assign n6197 = po28  & n6196;
  assign n6198 = ~n5863 & ~n6197;
  assign n6199 = n5863 & n6197;
  assign n6200 = ~n6198 & ~n6199;
  assign n6201 = ~n6195 & ~n6200;
  assign n6202 = ~n6194 & ~n6201;
  assign n6203 = po52  & ~n6202;
  assign n6204 = ~po52  & n6202;
  assign n6205 = ~n5866 & ~n5867;
  assign n6206 = po28  & n6205;
  assign n6207 = ~n5872 & ~n6206;
  assign n6208 = n5872 & n6206;
  assign n6209 = ~n6207 & ~n6208;
  assign n6210 = ~n6204 & ~n6209;
  assign n6211 = ~n6203 & ~n6210;
  assign n6212 = po53  & ~n6211;
  assign n6213 = ~po53  & n6211;
  assign n6214 = ~n5875 & ~n5876;
  assign n6215 = po28  & n6214;
  assign n6216 = ~n5881 & ~n6215;
  assign n6217 = n5881 & n6215;
  assign n6218 = ~n6216 & ~n6217;
  assign n6219 = ~n6213 & ~n6218;
  assign n6220 = ~n6212 & ~n6219;
  assign n6221 = po54  & ~n6220;
  assign n6222 = ~po54  & n6220;
  assign n6223 = ~n5884 & ~n5885;
  assign n6224 = po28  & n6223;
  assign n6225 = ~n5890 & ~n6224;
  assign n6226 = n5890 & n6224;
  assign n6227 = ~n6225 & ~n6226;
  assign n6228 = ~n6222 & ~n6227;
  assign n6229 = ~n6221 & ~n6228;
  assign n6230 = po55  & ~n6229;
  assign n6231 = ~po55  & n6229;
  assign n6232 = ~n5893 & ~n5894;
  assign n6233 = po28  & n6232;
  assign n6234 = ~n5899 & ~n6233;
  assign n6235 = n5899 & n6233;
  assign n6236 = ~n6234 & ~n6235;
  assign n6237 = ~n6231 & ~n6236;
  assign n6238 = ~n6230 & ~n6237;
  assign n6239 = po56  & ~n6238;
  assign n6240 = ~po56  & n6238;
  assign n6241 = ~n5902 & ~n5903;
  assign n6242 = po28  & n6241;
  assign n6243 = ~n5908 & ~n6242;
  assign n6244 = n5908 & n6242;
  assign n6245 = ~n6243 & ~n6244;
  assign n6246 = ~n6240 & ~n6245;
  assign n6247 = ~n6239 & ~n6246;
  assign n6248 = po57  & ~n6247;
  assign n6249 = ~po57  & n6247;
  assign n6250 = ~n5911 & ~n5912;
  assign n6251 = po28  & n6250;
  assign n6252 = ~n5917 & ~n6251;
  assign n6253 = n5917 & n6251;
  assign n6254 = ~n6252 & ~n6253;
  assign n6255 = ~n6249 & ~n6254;
  assign n6256 = ~n6248 & ~n6255;
  assign n6257 = po58  & ~n6256;
  assign n6258 = ~po58  & n6256;
  assign n6259 = ~n5920 & ~n5921;
  assign n6260 = po28  & n6259;
  assign n6261 = ~n5926 & ~n6260;
  assign n6262 = n5926 & n6260;
  assign n6263 = ~n6261 & ~n6262;
  assign n6264 = ~n6258 & ~n6263;
  assign n6265 = ~n6257 & ~n6264;
  assign n6266 = po59  & ~n6265;
  assign n6267 = ~po59  & n6265;
  assign n6268 = ~n5929 & ~n5930;
  assign n6269 = po28  & n6268;
  assign n6270 = ~n5935 & ~n6269;
  assign n6271 = n5935 & n6269;
  assign n6272 = ~n6270 & ~n6271;
  assign n6273 = ~n6267 & ~n6272;
  assign n6274 = ~n6266 & ~n6273;
  assign n6275 = po60  & ~n6274;
  assign n6276 = ~po60  & n6274;
  assign n6277 = ~n5938 & ~n5939;
  assign n6278 = po28  & n6277;
  assign n6279 = ~n5944 & ~n6278;
  assign n6280 = n5944 & n6278;
  assign n6281 = ~n6279 & ~n6280;
  assign n6282 = ~n6276 & ~n6281;
  assign n6283 = ~n6275 & ~n6282;
  assign n6284 = po61  & ~n6283;
  assign n6285 = ~po61  & n6283;
  assign n6286 = ~n5947 & ~n5948;
  assign n6287 = po28  & n6286;
  assign n6288 = ~n5953 & ~n6287;
  assign n6289 = n5953 & n6287;
  assign n6290 = ~n6288 & ~n6289;
  assign n6291 = ~n6285 & ~n6290;
  assign n6292 = ~n6284 & ~n6291;
  assign n6293 = po62  & ~n6292;
  assign n6294 = ~po62  & n6292;
  assign n6295 = ~n5956 & ~n5957;
  assign n6296 = po28  & n6295;
  assign n6297 = ~n5962 & ~n6296;
  assign n6298 = n5962 & n6296;
  assign n6299 = ~n6297 & ~n6298;
  assign n6300 = ~n6294 & ~n6299;
  assign n6301 = ~n6293 & ~n6300;
  assign n6302 = n6065 & n6301;
  assign n6303 = ~n6065 & ~n6301;
  assign n6304 = n5975 & po28 ;
  assign n6305 = ~n5974 & ~n6304;
  assign n6306 = n6303 & n6305;
  assign n6307 = ~po63  & ~n6306;
  assign n6308 = ~n5728 & po28 ;
  assign n6309 = n5973 & ~n6308;
  assign n6310 = po63  & ~n5975;
  assign n6311 = ~n6309 & n6310;
  assign n6312 = ~n6302 & ~n6311;
  assign n6313 = ~n6307 & n6312;
  assign po27  = n6060 | ~n6313;
  assign n6315 = ~n6058 & ~n6059;
  assign n6316 = po27  & n6315;
  assign n6317 = ~n5991 & ~n6316;
  assign n6318 = n5991 & n6316;
  assign n6319 = ~n6317 & ~n6318;
  assign n6320 = pi54  & po27 ;
  assign n6321 = ~pi52  & ~pi53 ;
  assign n6322 = ~pi54  & n6321;
  assign n6323 = ~n6320 & ~n6322;
  assign n6324 = po28  & ~n6323;
  assign n6325 = ~po28  & n6323;
  assign n6326 = ~pi54  & po27 ;
  assign n6327 = pi55  & ~n6326;
  assign n6328 = ~pi55  & n6326;
  assign n6329 = ~n6327 & ~n6328;
  assign n6330 = ~n6325 & n6329;
  assign n6331 = ~n6324 & ~n6330;
  assign n6332 = po29  & ~n6331;
  assign n6333 = ~po29  & n6331;
  assign n6334 = po28  & n6313;
  assign n6335 = ~n6328 & ~n6334;
  assign n6336 = pi56  & ~n6335;
  assign n6337 = ~pi56  & n6335;
  assign n6338 = ~n6336 & ~n6337;
  assign n6339 = ~n6333 & ~n6338;
  assign n6340 = ~n6332 & ~n6339;
  assign n6341 = po30  & ~n6340;
  assign n6342 = ~po30  & n6340;
  assign n6343 = ~n5996 & ~n5997;
  assign n6344 = po27  & n6343;
  assign n6345 = n6001 & ~n6344;
  assign n6346 = ~n6001 & n6344;
  assign n6347 = ~n6345 & ~n6346;
  assign n6348 = ~n6342 & ~n6347;
  assign n6349 = ~n6341 & ~n6348;
  assign n6350 = po31  & ~n6349;
  assign n6351 = ~po31  & n6349;
  assign n6352 = ~n6004 & ~n6005;
  assign n6353 = po27  & n6352;
  assign n6354 = ~n6010 & ~n6353;
  assign n6355 = n6010 & n6353;
  assign n6356 = ~n6354 & ~n6355;
  assign n6357 = ~n6351 & ~n6356;
  assign n6358 = ~n6350 & ~n6357;
  assign n6359 = po32  & ~n6358;
  assign n6360 = ~po32  & n6358;
  assign n6361 = ~n6013 & ~n6014;
  assign n6362 = po27  & n6361;
  assign n6363 = n6019 & n6362;
  assign n6364 = ~n6019 & ~n6362;
  assign n6365 = ~n6363 & ~n6364;
  assign n6366 = ~n6360 & ~n6365;
  assign n6367 = ~n6359 & ~n6366;
  assign n6368 = po33  & ~n6367;
  assign n6369 = ~po33  & n6367;
  assign n6370 = ~n6022 & ~n6023;
  assign n6371 = po27  & n6370;
  assign n6372 = ~n6028 & ~n6371;
  assign n6373 = n6028 & n6371;
  assign n6374 = ~n6372 & ~n6373;
  assign n6375 = ~n6369 & ~n6374;
  assign n6376 = ~n6368 & ~n6375;
  assign n6377 = po34  & ~n6376;
  assign n6378 = ~po34  & n6376;
  assign n6379 = ~n6031 & ~n6032;
  assign n6380 = po27  & n6379;
  assign n6381 = ~n6037 & ~n6380;
  assign n6382 = n6037 & n6380;
  assign n6383 = ~n6381 & ~n6382;
  assign n6384 = ~n6378 & ~n6383;
  assign n6385 = ~n6377 & ~n6384;
  assign n6386 = po35  & ~n6385;
  assign n6387 = ~po35  & n6385;
  assign n6388 = ~n6040 & ~n6041;
  assign n6389 = po27  & n6388;
  assign n6390 = ~n6046 & ~n6389;
  assign n6391 = n6046 & n6389;
  assign n6392 = ~n6390 & ~n6391;
  assign n6393 = ~n6387 & ~n6392;
  assign n6394 = ~n6386 & ~n6393;
  assign n6395 = po36  & ~n6394;
  assign n6396 = ~n6049 & ~n6055;
  assign n6397 = po27  & n6396;
  assign n6398 = ~n6054 & ~n6397;
  assign n6399 = n6054 & n6397;
  assign n6400 = ~n6398 & ~n6399;
  assign n6401 = ~po36  & n6394;
  assign n6402 = ~n6400 & ~n6401;
  assign n6403 = ~n6395 & ~n6402;
  assign n6404 = po37  & ~n6403;
  assign n6405 = ~po37  & n6403;
  assign n6406 = n6065 & ~po27 ;
  assign n6407 = ~n6293 & ~n6294;
  assign n6408 = po27  & n6407;
  assign n6409 = ~n6299 & ~n6408;
  assign n6410 = n6299 & n6408;
  assign n6411 = ~n6409 & ~n6410;
  assign n6412 = ~n6319 & ~n6405;
  assign n6413 = ~n6404 & ~n6412;
  assign n6414 = po38  & ~n6413;
  assign n6415 = ~po38  & n6413;
  assign n6416 = ~n6068 & ~n6069;
  assign n6417 = po27  & n6416;
  assign n6418 = ~n6074 & ~n6417;
  assign n6419 = n6074 & n6417;
  assign n6420 = ~n6418 & ~n6419;
  assign n6421 = ~n6415 & ~n6420;
  assign n6422 = ~n6414 & ~n6421;
  assign n6423 = po39  & ~n6422;
  assign n6424 = ~po39  & n6422;
  assign n6425 = ~n6077 & ~n6078;
  assign n6426 = po27  & n6425;
  assign n6427 = ~n6083 & ~n6426;
  assign n6428 = n6083 & n6426;
  assign n6429 = ~n6427 & ~n6428;
  assign n6430 = ~n6424 & ~n6429;
  assign n6431 = ~n6423 & ~n6430;
  assign n6432 = po40  & ~n6431;
  assign n6433 = ~po40  & n6431;
  assign n6434 = ~n6086 & ~n6087;
  assign n6435 = po27  & n6434;
  assign n6436 = ~n6092 & ~n6435;
  assign n6437 = n6092 & n6435;
  assign n6438 = ~n6436 & ~n6437;
  assign n6439 = ~n6433 & ~n6438;
  assign n6440 = ~n6432 & ~n6439;
  assign n6441 = po41  & ~n6440;
  assign n6442 = ~po41  & n6440;
  assign n6443 = ~n6095 & ~n6096;
  assign n6444 = po27  & n6443;
  assign n6445 = ~n6101 & ~n6444;
  assign n6446 = n6101 & n6444;
  assign n6447 = ~n6445 & ~n6446;
  assign n6448 = ~n6442 & ~n6447;
  assign n6449 = ~n6441 & ~n6448;
  assign n6450 = po42  & ~n6449;
  assign n6451 = ~po42  & n6449;
  assign n6452 = ~n6104 & ~n6105;
  assign n6453 = po27  & n6452;
  assign n6454 = ~n6110 & ~n6453;
  assign n6455 = n6110 & n6453;
  assign n6456 = ~n6454 & ~n6455;
  assign n6457 = ~n6451 & ~n6456;
  assign n6458 = ~n6450 & ~n6457;
  assign n6459 = po43  & ~n6458;
  assign n6460 = ~po43  & n6458;
  assign n6461 = ~n6113 & ~n6114;
  assign n6462 = po27  & n6461;
  assign n6463 = ~n6119 & ~n6462;
  assign n6464 = n6119 & n6462;
  assign n6465 = ~n6463 & ~n6464;
  assign n6466 = ~n6460 & ~n6465;
  assign n6467 = ~n6459 & ~n6466;
  assign n6468 = po44  & ~n6467;
  assign n6469 = ~po44  & n6467;
  assign n6470 = ~n6122 & ~n6123;
  assign n6471 = po27  & n6470;
  assign n6472 = ~n6128 & ~n6471;
  assign n6473 = n6128 & n6471;
  assign n6474 = ~n6472 & ~n6473;
  assign n6475 = ~n6469 & ~n6474;
  assign n6476 = ~n6468 & ~n6475;
  assign n6477 = po45  & ~n6476;
  assign n6478 = ~po45  & n6476;
  assign n6479 = ~n6131 & ~n6132;
  assign n6480 = po27  & n6479;
  assign n6481 = ~n6137 & ~n6480;
  assign n6482 = n6137 & n6480;
  assign n6483 = ~n6481 & ~n6482;
  assign n6484 = ~n6478 & ~n6483;
  assign n6485 = ~n6477 & ~n6484;
  assign n6486 = po46  & ~n6485;
  assign n6487 = ~po46  & n6485;
  assign n6488 = ~n6140 & ~n6141;
  assign n6489 = po27  & n6488;
  assign n6490 = ~n6146 & ~n6489;
  assign n6491 = n6146 & n6489;
  assign n6492 = ~n6490 & ~n6491;
  assign n6493 = ~n6487 & ~n6492;
  assign n6494 = ~n6486 & ~n6493;
  assign n6495 = po47  & ~n6494;
  assign n6496 = ~po47  & n6494;
  assign n6497 = ~n6149 & ~n6150;
  assign n6498 = po27  & n6497;
  assign n6499 = ~n6155 & ~n6498;
  assign n6500 = n6155 & n6498;
  assign n6501 = ~n6499 & ~n6500;
  assign n6502 = ~n6496 & ~n6501;
  assign n6503 = ~n6495 & ~n6502;
  assign n6504 = po48  & ~n6503;
  assign n6505 = ~po48  & n6503;
  assign n6506 = ~n6158 & ~n6159;
  assign n6507 = po27  & n6506;
  assign n6508 = ~n6164 & ~n6507;
  assign n6509 = n6164 & n6507;
  assign n6510 = ~n6508 & ~n6509;
  assign n6511 = ~n6505 & ~n6510;
  assign n6512 = ~n6504 & ~n6511;
  assign n6513 = po49  & ~n6512;
  assign n6514 = ~po49  & n6512;
  assign n6515 = ~n6167 & ~n6168;
  assign n6516 = po27  & n6515;
  assign n6517 = ~n6173 & ~n6516;
  assign n6518 = n6173 & n6516;
  assign n6519 = ~n6517 & ~n6518;
  assign n6520 = ~n6514 & ~n6519;
  assign n6521 = ~n6513 & ~n6520;
  assign n6522 = po50  & ~n6521;
  assign n6523 = ~po50  & n6521;
  assign n6524 = ~n6176 & ~n6177;
  assign n6525 = po27  & n6524;
  assign n6526 = ~n6182 & ~n6525;
  assign n6527 = n6182 & n6525;
  assign n6528 = ~n6526 & ~n6527;
  assign n6529 = ~n6523 & ~n6528;
  assign n6530 = ~n6522 & ~n6529;
  assign n6531 = po51  & ~n6530;
  assign n6532 = ~po51  & n6530;
  assign n6533 = ~n6185 & ~n6186;
  assign n6534 = po27  & n6533;
  assign n6535 = ~n6191 & ~n6534;
  assign n6536 = n6191 & n6534;
  assign n6537 = ~n6535 & ~n6536;
  assign n6538 = ~n6532 & ~n6537;
  assign n6539 = ~n6531 & ~n6538;
  assign n6540 = po52  & ~n6539;
  assign n6541 = ~po52  & n6539;
  assign n6542 = ~n6194 & ~n6195;
  assign n6543 = po27  & n6542;
  assign n6544 = ~n6200 & ~n6543;
  assign n6545 = n6200 & n6543;
  assign n6546 = ~n6544 & ~n6545;
  assign n6547 = ~n6541 & ~n6546;
  assign n6548 = ~n6540 & ~n6547;
  assign n6549 = po53  & ~n6548;
  assign n6550 = ~po53  & n6548;
  assign n6551 = ~n6203 & ~n6204;
  assign n6552 = po27  & n6551;
  assign n6553 = ~n6209 & ~n6552;
  assign n6554 = n6209 & n6552;
  assign n6555 = ~n6553 & ~n6554;
  assign n6556 = ~n6550 & ~n6555;
  assign n6557 = ~n6549 & ~n6556;
  assign n6558 = po54  & ~n6557;
  assign n6559 = ~po54  & n6557;
  assign n6560 = ~n6212 & ~n6213;
  assign n6561 = po27  & n6560;
  assign n6562 = ~n6218 & ~n6561;
  assign n6563 = n6218 & n6561;
  assign n6564 = ~n6562 & ~n6563;
  assign n6565 = ~n6559 & ~n6564;
  assign n6566 = ~n6558 & ~n6565;
  assign n6567 = po55  & ~n6566;
  assign n6568 = ~po55  & n6566;
  assign n6569 = ~n6221 & ~n6222;
  assign n6570 = po27  & n6569;
  assign n6571 = ~n6227 & ~n6570;
  assign n6572 = n6227 & n6570;
  assign n6573 = ~n6571 & ~n6572;
  assign n6574 = ~n6568 & ~n6573;
  assign n6575 = ~n6567 & ~n6574;
  assign n6576 = po56  & ~n6575;
  assign n6577 = ~po56  & n6575;
  assign n6578 = ~n6230 & ~n6231;
  assign n6579 = po27  & n6578;
  assign n6580 = ~n6236 & ~n6579;
  assign n6581 = n6236 & n6579;
  assign n6582 = ~n6580 & ~n6581;
  assign n6583 = ~n6577 & ~n6582;
  assign n6584 = ~n6576 & ~n6583;
  assign n6585 = po57  & ~n6584;
  assign n6586 = ~po57  & n6584;
  assign n6587 = ~n6239 & ~n6240;
  assign n6588 = po27  & n6587;
  assign n6589 = ~n6245 & ~n6588;
  assign n6590 = n6245 & n6588;
  assign n6591 = ~n6589 & ~n6590;
  assign n6592 = ~n6586 & ~n6591;
  assign n6593 = ~n6585 & ~n6592;
  assign n6594 = po58  & ~n6593;
  assign n6595 = ~po58  & n6593;
  assign n6596 = ~n6248 & ~n6249;
  assign n6597 = po27  & n6596;
  assign n6598 = ~n6254 & ~n6597;
  assign n6599 = n6254 & n6597;
  assign n6600 = ~n6598 & ~n6599;
  assign n6601 = ~n6595 & ~n6600;
  assign n6602 = ~n6594 & ~n6601;
  assign n6603 = po59  & ~n6602;
  assign n6604 = ~po59  & n6602;
  assign n6605 = ~n6257 & ~n6258;
  assign n6606 = po27  & n6605;
  assign n6607 = ~n6263 & ~n6606;
  assign n6608 = n6263 & n6606;
  assign n6609 = ~n6607 & ~n6608;
  assign n6610 = ~n6604 & ~n6609;
  assign n6611 = ~n6603 & ~n6610;
  assign n6612 = po60  & ~n6611;
  assign n6613 = ~po60  & n6611;
  assign n6614 = ~n6266 & ~n6267;
  assign n6615 = po27  & n6614;
  assign n6616 = ~n6272 & ~n6615;
  assign n6617 = n6272 & n6615;
  assign n6618 = ~n6616 & ~n6617;
  assign n6619 = ~n6613 & ~n6618;
  assign n6620 = ~n6612 & ~n6619;
  assign n6621 = po61  & ~n6620;
  assign n6622 = ~po61  & n6620;
  assign n6623 = ~n6275 & ~n6276;
  assign n6624 = po27  & n6623;
  assign n6625 = ~n6281 & ~n6624;
  assign n6626 = n6281 & n6624;
  assign n6627 = ~n6625 & ~n6626;
  assign n6628 = ~n6622 & ~n6627;
  assign n6629 = ~n6621 & ~n6628;
  assign n6630 = po62  & ~n6629;
  assign n6631 = ~po62  & n6629;
  assign n6632 = ~n6284 & ~n6285;
  assign n6633 = po27  & n6632;
  assign n6634 = ~n6290 & ~n6633;
  assign n6635 = n6290 & n6633;
  assign n6636 = ~n6634 & ~n6635;
  assign n6637 = ~n6631 & ~n6636;
  assign n6638 = ~n6630 & ~n6637;
  assign n6639 = n6411 & n6638;
  assign n6640 = ~n6411 & ~n6638;
  assign n6641 = n6303 & po27 ;
  assign n6642 = ~n6302 & ~n6641;
  assign n6643 = n6640 & n6642;
  assign n6644 = ~po63  & ~n6643;
  assign n6645 = ~n6065 & po27 ;
  assign n6646 = n6301 & ~n6645;
  assign n6647 = po63  & ~n6303;
  assign n6648 = ~n6646 & n6647;
  assign n6649 = ~n6639 & ~n6648;
  assign n6650 = ~n6644 & n6649;
  assign po26  = n6406 | ~n6650;
  assign n6652 = ~n6404 & ~n6405;
  assign n6653 = po26  & n6652;
  assign n6654 = ~n6319 & ~n6653;
  assign n6655 = n6319 & n6653;
  assign n6656 = ~n6654 & ~n6655;
  assign n6657 = pi52  & po26 ;
  assign n6658 = ~pi50  & ~pi51 ;
  assign n6659 = ~pi52  & n6658;
  assign n6660 = ~n6657 & ~n6659;
  assign n6661 = po27  & ~n6660;
  assign n6662 = ~po27  & n6660;
  assign n6663 = ~pi52  & po26 ;
  assign n6664 = pi53  & ~n6663;
  assign n6665 = ~pi53  & n6663;
  assign n6666 = ~n6664 & ~n6665;
  assign n6667 = ~n6662 & n6666;
  assign n6668 = ~n6661 & ~n6667;
  assign n6669 = po28  & ~n6668;
  assign n6670 = ~po28  & n6668;
  assign n6671 = po27  & n6650;
  assign n6672 = ~n6665 & ~n6671;
  assign n6673 = pi54  & ~n6672;
  assign n6674 = ~pi54  & n6672;
  assign n6675 = ~n6673 & ~n6674;
  assign n6676 = ~n6670 & ~n6675;
  assign n6677 = ~n6669 & ~n6676;
  assign n6678 = po29  & ~n6677;
  assign n6679 = ~po29  & n6677;
  assign n6680 = ~n6324 & ~n6325;
  assign n6681 = po26  & n6680;
  assign n6682 = n6329 & ~n6681;
  assign n6683 = ~n6329 & n6681;
  assign n6684 = ~n6682 & ~n6683;
  assign n6685 = ~n6679 & ~n6684;
  assign n6686 = ~n6678 & ~n6685;
  assign n6687 = po30  & ~n6686;
  assign n6688 = ~po30  & n6686;
  assign n6689 = ~n6332 & ~n6333;
  assign n6690 = po26  & n6689;
  assign n6691 = ~n6338 & ~n6690;
  assign n6692 = n6338 & n6690;
  assign n6693 = ~n6691 & ~n6692;
  assign n6694 = ~n6688 & ~n6693;
  assign n6695 = ~n6687 & ~n6694;
  assign n6696 = po31  & ~n6695;
  assign n6697 = ~po31  & n6695;
  assign n6698 = ~n6341 & ~n6342;
  assign n6699 = po26  & n6698;
  assign n6700 = n6347 & n6699;
  assign n6701 = ~n6347 & ~n6699;
  assign n6702 = ~n6700 & ~n6701;
  assign n6703 = ~n6697 & ~n6702;
  assign n6704 = ~n6696 & ~n6703;
  assign n6705 = po32  & ~n6704;
  assign n6706 = ~po32  & n6704;
  assign n6707 = ~n6350 & ~n6351;
  assign n6708 = po26  & n6707;
  assign n6709 = ~n6356 & ~n6708;
  assign n6710 = n6356 & n6708;
  assign n6711 = ~n6709 & ~n6710;
  assign n6712 = ~n6706 & ~n6711;
  assign n6713 = ~n6705 & ~n6712;
  assign n6714 = po33  & ~n6713;
  assign n6715 = ~po33  & n6713;
  assign n6716 = ~n6359 & ~n6360;
  assign n6717 = po26  & n6716;
  assign n6718 = ~n6365 & ~n6717;
  assign n6719 = n6365 & n6717;
  assign n6720 = ~n6718 & ~n6719;
  assign n6721 = ~n6715 & ~n6720;
  assign n6722 = ~n6714 & ~n6721;
  assign n6723 = po34  & ~n6722;
  assign n6724 = ~po34  & n6722;
  assign n6725 = ~n6368 & ~n6369;
  assign n6726 = po26  & n6725;
  assign n6727 = ~n6374 & ~n6726;
  assign n6728 = n6374 & n6726;
  assign n6729 = ~n6727 & ~n6728;
  assign n6730 = ~n6724 & ~n6729;
  assign n6731 = ~n6723 & ~n6730;
  assign n6732 = po35  & ~n6731;
  assign n6733 = ~po35  & n6731;
  assign n6734 = ~n6377 & ~n6378;
  assign n6735 = po26  & n6734;
  assign n6736 = ~n6383 & ~n6735;
  assign n6737 = n6383 & n6735;
  assign n6738 = ~n6736 & ~n6737;
  assign n6739 = ~n6733 & ~n6738;
  assign n6740 = ~n6732 & ~n6739;
  assign n6741 = po36  & ~n6740;
  assign n6742 = ~po36  & n6740;
  assign n6743 = ~n6386 & ~n6387;
  assign n6744 = po26  & n6743;
  assign n6745 = ~n6392 & ~n6744;
  assign n6746 = n6392 & n6744;
  assign n6747 = ~n6745 & ~n6746;
  assign n6748 = ~n6742 & ~n6747;
  assign n6749 = ~n6741 & ~n6748;
  assign n6750 = po37  & ~n6749;
  assign n6751 = ~n6395 & ~n6401;
  assign n6752 = po26  & n6751;
  assign n6753 = ~n6400 & ~n6752;
  assign n6754 = n6400 & n6752;
  assign n6755 = ~n6753 & ~n6754;
  assign n6756 = ~po37  & n6749;
  assign n6757 = ~n6755 & ~n6756;
  assign n6758 = ~n6750 & ~n6757;
  assign n6759 = po38  & ~n6758;
  assign n6760 = ~po38  & n6758;
  assign n6761 = n6411 & ~po26 ;
  assign n6762 = ~n6630 & ~n6631;
  assign n6763 = po26  & n6762;
  assign n6764 = ~n6636 & ~n6763;
  assign n6765 = n6636 & n6763;
  assign n6766 = ~n6764 & ~n6765;
  assign n6767 = ~n6656 & ~n6760;
  assign n6768 = ~n6759 & ~n6767;
  assign n6769 = po39  & ~n6768;
  assign n6770 = ~po39  & n6768;
  assign n6771 = ~n6414 & ~n6415;
  assign n6772 = po26  & n6771;
  assign n6773 = ~n6420 & ~n6772;
  assign n6774 = n6420 & n6772;
  assign n6775 = ~n6773 & ~n6774;
  assign n6776 = ~n6770 & ~n6775;
  assign n6777 = ~n6769 & ~n6776;
  assign n6778 = po40  & ~n6777;
  assign n6779 = ~po40  & n6777;
  assign n6780 = ~n6423 & ~n6424;
  assign n6781 = po26  & n6780;
  assign n6782 = ~n6429 & ~n6781;
  assign n6783 = n6429 & n6781;
  assign n6784 = ~n6782 & ~n6783;
  assign n6785 = ~n6779 & ~n6784;
  assign n6786 = ~n6778 & ~n6785;
  assign n6787 = po41  & ~n6786;
  assign n6788 = ~po41  & n6786;
  assign n6789 = ~n6432 & ~n6433;
  assign n6790 = po26  & n6789;
  assign n6791 = ~n6438 & ~n6790;
  assign n6792 = n6438 & n6790;
  assign n6793 = ~n6791 & ~n6792;
  assign n6794 = ~n6788 & ~n6793;
  assign n6795 = ~n6787 & ~n6794;
  assign n6796 = po42  & ~n6795;
  assign n6797 = ~po42  & n6795;
  assign n6798 = ~n6441 & ~n6442;
  assign n6799 = po26  & n6798;
  assign n6800 = ~n6447 & ~n6799;
  assign n6801 = n6447 & n6799;
  assign n6802 = ~n6800 & ~n6801;
  assign n6803 = ~n6797 & ~n6802;
  assign n6804 = ~n6796 & ~n6803;
  assign n6805 = po43  & ~n6804;
  assign n6806 = ~po43  & n6804;
  assign n6807 = ~n6450 & ~n6451;
  assign n6808 = po26  & n6807;
  assign n6809 = ~n6456 & ~n6808;
  assign n6810 = n6456 & n6808;
  assign n6811 = ~n6809 & ~n6810;
  assign n6812 = ~n6806 & ~n6811;
  assign n6813 = ~n6805 & ~n6812;
  assign n6814 = po44  & ~n6813;
  assign n6815 = ~po44  & n6813;
  assign n6816 = ~n6459 & ~n6460;
  assign n6817 = po26  & n6816;
  assign n6818 = ~n6465 & ~n6817;
  assign n6819 = n6465 & n6817;
  assign n6820 = ~n6818 & ~n6819;
  assign n6821 = ~n6815 & ~n6820;
  assign n6822 = ~n6814 & ~n6821;
  assign n6823 = po45  & ~n6822;
  assign n6824 = ~po45  & n6822;
  assign n6825 = ~n6468 & ~n6469;
  assign n6826 = po26  & n6825;
  assign n6827 = ~n6474 & ~n6826;
  assign n6828 = n6474 & n6826;
  assign n6829 = ~n6827 & ~n6828;
  assign n6830 = ~n6824 & ~n6829;
  assign n6831 = ~n6823 & ~n6830;
  assign n6832 = po46  & ~n6831;
  assign n6833 = ~po46  & n6831;
  assign n6834 = ~n6477 & ~n6478;
  assign n6835 = po26  & n6834;
  assign n6836 = ~n6483 & ~n6835;
  assign n6837 = n6483 & n6835;
  assign n6838 = ~n6836 & ~n6837;
  assign n6839 = ~n6833 & ~n6838;
  assign n6840 = ~n6832 & ~n6839;
  assign n6841 = po47  & ~n6840;
  assign n6842 = ~po47  & n6840;
  assign n6843 = ~n6486 & ~n6487;
  assign n6844 = po26  & n6843;
  assign n6845 = ~n6492 & ~n6844;
  assign n6846 = n6492 & n6844;
  assign n6847 = ~n6845 & ~n6846;
  assign n6848 = ~n6842 & ~n6847;
  assign n6849 = ~n6841 & ~n6848;
  assign n6850 = po48  & ~n6849;
  assign n6851 = ~po48  & n6849;
  assign n6852 = ~n6495 & ~n6496;
  assign n6853 = po26  & n6852;
  assign n6854 = ~n6501 & ~n6853;
  assign n6855 = n6501 & n6853;
  assign n6856 = ~n6854 & ~n6855;
  assign n6857 = ~n6851 & ~n6856;
  assign n6858 = ~n6850 & ~n6857;
  assign n6859 = po49  & ~n6858;
  assign n6860 = ~po49  & n6858;
  assign n6861 = ~n6504 & ~n6505;
  assign n6862 = po26  & n6861;
  assign n6863 = ~n6510 & ~n6862;
  assign n6864 = n6510 & n6862;
  assign n6865 = ~n6863 & ~n6864;
  assign n6866 = ~n6860 & ~n6865;
  assign n6867 = ~n6859 & ~n6866;
  assign n6868 = po50  & ~n6867;
  assign n6869 = ~po50  & n6867;
  assign n6870 = ~n6513 & ~n6514;
  assign n6871 = po26  & n6870;
  assign n6872 = ~n6519 & ~n6871;
  assign n6873 = n6519 & n6871;
  assign n6874 = ~n6872 & ~n6873;
  assign n6875 = ~n6869 & ~n6874;
  assign n6876 = ~n6868 & ~n6875;
  assign n6877 = po51  & ~n6876;
  assign n6878 = ~po51  & n6876;
  assign n6879 = ~n6522 & ~n6523;
  assign n6880 = po26  & n6879;
  assign n6881 = ~n6528 & ~n6880;
  assign n6882 = n6528 & n6880;
  assign n6883 = ~n6881 & ~n6882;
  assign n6884 = ~n6878 & ~n6883;
  assign n6885 = ~n6877 & ~n6884;
  assign n6886 = po52  & ~n6885;
  assign n6887 = ~po52  & n6885;
  assign n6888 = ~n6531 & ~n6532;
  assign n6889 = po26  & n6888;
  assign n6890 = ~n6537 & ~n6889;
  assign n6891 = n6537 & n6889;
  assign n6892 = ~n6890 & ~n6891;
  assign n6893 = ~n6887 & ~n6892;
  assign n6894 = ~n6886 & ~n6893;
  assign n6895 = po53  & ~n6894;
  assign n6896 = ~po53  & n6894;
  assign n6897 = ~n6540 & ~n6541;
  assign n6898 = po26  & n6897;
  assign n6899 = ~n6546 & ~n6898;
  assign n6900 = n6546 & n6898;
  assign n6901 = ~n6899 & ~n6900;
  assign n6902 = ~n6896 & ~n6901;
  assign n6903 = ~n6895 & ~n6902;
  assign n6904 = po54  & ~n6903;
  assign n6905 = ~po54  & n6903;
  assign n6906 = ~n6549 & ~n6550;
  assign n6907 = po26  & n6906;
  assign n6908 = ~n6555 & ~n6907;
  assign n6909 = n6555 & n6907;
  assign n6910 = ~n6908 & ~n6909;
  assign n6911 = ~n6905 & ~n6910;
  assign n6912 = ~n6904 & ~n6911;
  assign n6913 = po55  & ~n6912;
  assign n6914 = ~po55  & n6912;
  assign n6915 = ~n6558 & ~n6559;
  assign n6916 = po26  & n6915;
  assign n6917 = ~n6564 & ~n6916;
  assign n6918 = n6564 & n6916;
  assign n6919 = ~n6917 & ~n6918;
  assign n6920 = ~n6914 & ~n6919;
  assign n6921 = ~n6913 & ~n6920;
  assign n6922 = po56  & ~n6921;
  assign n6923 = ~po56  & n6921;
  assign n6924 = ~n6567 & ~n6568;
  assign n6925 = po26  & n6924;
  assign n6926 = ~n6573 & ~n6925;
  assign n6927 = n6573 & n6925;
  assign n6928 = ~n6926 & ~n6927;
  assign n6929 = ~n6923 & ~n6928;
  assign n6930 = ~n6922 & ~n6929;
  assign n6931 = po57  & ~n6930;
  assign n6932 = ~po57  & n6930;
  assign n6933 = ~n6576 & ~n6577;
  assign n6934 = po26  & n6933;
  assign n6935 = ~n6582 & ~n6934;
  assign n6936 = n6582 & n6934;
  assign n6937 = ~n6935 & ~n6936;
  assign n6938 = ~n6932 & ~n6937;
  assign n6939 = ~n6931 & ~n6938;
  assign n6940 = po58  & ~n6939;
  assign n6941 = ~po58  & n6939;
  assign n6942 = ~n6585 & ~n6586;
  assign n6943 = po26  & n6942;
  assign n6944 = ~n6591 & ~n6943;
  assign n6945 = n6591 & n6943;
  assign n6946 = ~n6944 & ~n6945;
  assign n6947 = ~n6941 & ~n6946;
  assign n6948 = ~n6940 & ~n6947;
  assign n6949 = po59  & ~n6948;
  assign n6950 = ~po59  & n6948;
  assign n6951 = ~n6594 & ~n6595;
  assign n6952 = po26  & n6951;
  assign n6953 = ~n6600 & ~n6952;
  assign n6954 = n6600 & n6952;
  assign n6955 = ~n6953 & ~n6954;
  assign n6956 = ~n6950 & ~n6955;
  assign n6957 = ~n6949 & ~n6956;
  assign n6958 = po60  & ~n6957;
  assign n6959 = ~po60  & n6957;
  assign n6960 = ~n6603 & ~n6604;
  assign n6961 = po26  & n6960;
  assign n6962 = ~n6609 & ~n6961;
  assign n6963 = n6609 & n6961;
  assign n6964 = ~n6962 & ~n6963;
  assign n6965 = ~n6959 & ~n6964;
  assign n6966 = ~n6958 & ~n6965;
  assign n6967 = po61  & ~n6966;
  assign n6968 = ~po61  & n6966;
  assign n6969 = ~n6612 & ~n6613;
  assign n6970 = po26  & n6969;
  assign n6971 = ~n6618 & ~n6970;
  assign n6972 = n6618 & n6970;
  assign n6973 = ~n6971 & ~n6972;
  assign n6974 = ~n6968 & ~n6973;
  assign n6975 = ~n6967 & ~n6974;
  assign n6976 = po62  & ~n6975;
  assign n6977 = ~po62  & n6975;
  assign n6978 = ~n6621 & ~n6622;
  assign n6979 = po26  & n6978;
  assign n6980 = ~n6627 & ~n6979;
  assign n6981 = n6627 & n6979;
  assign n6982 = ~n6980 & ~n6981;
  assign n6983 = ~n6977 & ~n6982;
  assign n6984 = ~n6976 & ~n6983;
  assign n6985 = n6766 & n6984;
  assign n6986 = ~n6766 & ~n6984;
  assign n6987 = n6640 & po26 ;
  assign n6988 = ~n6639 & ~n6987;
  assign n6989 = n6986 & n6988;
  assign n6990 = ~po63  & ~n6989;
  assign n6991 = ~n6411 & po26 ;
  assign n6992 = n6638 & ~n6991;
  assign n6993 = po63  & ~n6640;
  assign n6994 = ~n6992 & n6993;
  assign n6995 = ~n6985 & ~n6994;
  assign n6996 = ~n6990 & n6995;
  assign po25  = n6761 | ~n6996;
  assign n6998 = ~n6759 & ~n6760;
  assign n6999 = po25  & n6998;
  assign n7000 = ~n6656 & ~n6999;
  assign n7001 = n6656 & n6999;
  assign n7002 = ~n7000 & ~n7001;
  assign n7003 = pi50  & po25 ;
  assign n7004 = ~pi48  & ~pi49 ;
  assign n7005 = ~pi50  & n7004;
  assign n7006 = ~n7003 & ~n7005;
  assign n7007 = po26  & ~n7006;
  assign n7008 = ~po26  & n7006;
  assign n7009 = ~pi50  & po25 ;
  assign n7010 = pi51  & ~n7009;
  assign n7011 = ~pi51  & n7009;
  assign n7012 = ~n7010 & ~n7011;
  assign n7013 = ~n7008 & n7012;
  assign n7014 = ~n7007 & ~n7013;
  assign n7015 = po27  & ~n7014;
  assign n7016 = ~po27  & n7014;
  assign n7017 = po26  & n6996;
  assign n7018 = ~n7011 & ~n7017;
  assign n7019 = pi52  & ~n7018;
  assign n7020 = ~pi52  & n7018;
  assign n7021 = ~n7019 & ~n7020;
  assign n7022 = ~n7016 & ~n7021;
  assign n7023 = ~n7015 & ~n7022;
  assign n7024 = po28  & ~n7023;
  assign n7025 = ~po28  & n7023;
  assign n7026 = ~n6661 & ~n6662;
  assign n7027 = po25  & n7026;
  assign n7028 = n6666 & ~n7027;
  assign n7029 = ~n6666 & n7027;
  assign n7030 = ~n7028 & ~n7029;
  assign n7031 = ~n7025 & ~n7030;
  assign n7032 = ~n7024 & ~n7031;
  assign n7033 = po29  & ~n7032;
  assign n7034 = ~po29  & n7032;
  assign n7035 = ~n6669 & ~n6670;
  assign n7036 = po25  & n7035;
  assign n7037 = ~n6675 & ~n7036;
  assign n7038 = n6675 & n7036;
  assign n7039 = ~n7037 & ~n7038;
  assign n7040 = ~n7034 & ~n7039;
  assign n7041 = ~n7033 & ~n7040;
  assign n7042 = po30  & ~n7041;
  assign n7043 = ~po30  & n7041;
  assign n7044 = ~n6678 & ~n6679;
  assign n7045 = po25  & n7044;
  assign n7046 = n6684 & n7045;
  assign n7047 = ~n6684 & ~n7045;
  assign n7048 = ~n7046 & ~n7047;
  assign n7049 = ~n7043 & ~n7048;
  assign n7050 = ~n7042 & ~n7049;
  assign n7051 = po31  & ~n7050;
  assign n7052 = ~po31  & n7050;
  assign n7053 = ~n6687 & ~n6688;
  assign n7054 = po25  & n7053;
  assign n7055 = ~n6693 & ~n7054;
  assign n7056 = n6693 & n7054;
  assign n7057 = ~n7055 & ~n7056;
  assign n7058 = ~n7052 & ~n7057;
  assign n7059 = ~n7051 & ~n7058;
  assign n7060 = po32  & ~n7059;
  assign n7061 = ~po32  & n7059;
  assign n7062 = ~n6696 & ~n6697;
  assign n7063 = po25  & n7062;
  assign n7064 = ~n6702 & ~n7063;
  assign n7065 = n6702 & n7063;
  assign n7066 = ~n7064 & ~n7065;
  assign n7067 = ~n7061 & ~n7066;
  assign n7068 = ~n7060 & ~n7067;
  assign n7069 = po33  & ~n7068;
  assign n7070 = ~po33  & n7068;
  assign n7071 = ~n6705 & ~n6706;
  assign n7072 = po25  & n7071;
  assign n7073 = ~n6711 & ~n7072;
  assign n7074 = n6711 & n7072;
  assign n7075 = ~n7073 & ~n7074;
  assign n7076 = ~n7070 & ~n7075;
  assign n7077 = ~n7069 & ~n7076;
  assign n7078 = po34  & ~n7077;
  assign n7079 = ~po34  & n7077;
  assign n7080 = ~n6714 & ~n6715;
  assign n7081 = po25  & n7080;
  assign n7082 = ~n6720 & ~n7081;
  assign n7083 = n6720 & n7081;
  assign n7084 = ~n7082 & ~n7083;
  assign n7085 = ~n7079 & ~n7084;
  assign n7086 = ~n7078 & ~n7085;
  assign n7087 = po35  & ~n7086;
  assign n7088 = ~po35  & n7086;
  assign n7089 = ~n6723 & ~n6724;
  assign n7090 = po25  & n7089;
  assign n7091 = ~n6729 & ~n7090;
  assign n7092 = n6729 & n7090;
  assign n7093 = ~n7091 & ~n7092;
  assign n7094 = ~n7088 & ~n7093;
  assign n7095 = ~n7087 & ~n7094;
  assign n7096 = po36  & ~n7095;
  assign n7097 = ~po36  & n7095;
  assign n7098 = ~n6732 & ~n6733;
  assign n7099 = po25  & n7098;
  assign n7100 = ~n6738 & ~n7099;
  assign n7101 = n6738 & n7099;
  assign n7102 = ~n7100 & ~n7101;
  assign n7103 = ~n7097 & ~n7102;
  assign n7104 = ~n7096 & ~n7103;
  assign n7105 = po37  & ~n7104;
  assign n7106 = ~po37  & n7104;
  assign n7107 = ~n6741 & ~n6742;
  assign n7108 = po25  & n7107;
  assign n7109 = ~n6747 & ~n7108;
  assign n7110 = n6747 & n7108;
  assign n7111 = ~n7109 & ~n7110;
  assign n7112 = ~n7106 & ~n7111;
  assign n7113 = ~n7105 & ~n7112;
  assign n7114 = po38  & ~n7113;
  assign n7115 = ~n6750 & ~n6756;
  assign n7116 = po25  & n7115;
  assign n7117 = ~n6755 & ~n7116;
  assign n7118 = n6755 & n7116;
  assign n7119 = ~n7117 & ~n7118;
  assign n7120 = ~po38  & n7113;
  assign n7121 = ~n7119 & ~n7120;
  assign n7122 = ~n7114 & ~n7121;
  assign n7123 = po39  & ~n7122;
  assign n7124 = ~po39  & n7122;
  assign n7125 = n6766 & ~po25 ;
  assign n7126 = ~n6976 & ~n6977;
  assign n7127 = po25  & n7126;
  assign n7128 = ~n6982 & ~n7127;
  assign n7129 = n6982 & n7127;
  assign n7130 = ~n7128 & ~n7129;
  assign n7131 = ~n7002 & ~n7124;
  assign n7132 = ~n7123 & ~n7131;
  assign n7133 = po40  & ~n7132;
  assign n7134 = ~po40  & n7132;
  assign n7135 = ~n6769 & ~n6770;
  assign n7136 = po25  & n7135;
  assign n7137 = ~n6775 & ~n7136;
  assign n7138 = n6775 & n7136;
  assign n7139 = ~n7137 & ~n7138;
  assign n7140 = ~n7134 & ~n7139;
  assign n7141 = ~n7133 & ~n7140;
  assign n7142 = po41  & ~n7141;
  assign n7143 = ~po41  & n7141;
  assign n7144 = ~n6778 & ~n6779;
  assign n7145 = po25  & n7144;
  assign n7146 = ~n6784 & ~n7145;
  assign n7147 = n6784 & n7145;
  assign n7148 = ~n7146 & ~n7147;
  assign n7149 = ~n7143 & ~n7148;
  assign n7150 = ~n7142 & ~n7149;
  assign n7151 = po42  & ~n7150;
  assign n7152 = ~po42  & n7150;
  assign n7153 = ~n6787 & ~n6788;
  assign n7154 = po25  & n7153;
  assign n7155 = ~n6793 & ~n7154;
  assign n7156 = n6793 & n7154;
  assign n7157 = ~n7155 & ~n7156;
  assign n7158 = ~n7152 & ~n7157;
  assign n7159 = ~n7151 & ~n7158;
  assign n7160 = po43  & ~n7159;
  assign n7161 = ~po43  & n7159;
  assign n7162 = ~n6796 & ~n6797;
  assign n7163 = po25  & n7162;
  assign n7164 = ~n6802 & ~n7163;
  assign n7165 = n6802 & n7163;
  assign n7166 = ~n7164 & ~n7165;
  assign n7167 = ~n7161 & ~n7166;
  assign n7168 = ~n7160 & ~n7167;
  assign n7169 = po44  & ~n7168;
  assign n7170 = ~po44  & n7168;
  assign n7171 = ~n6805 & ~n6806;
  assign n7172 = po25  & n7171;
  assign n7173 = ~n6811 & ~n7172;
  assign n7174 = n6811 & n7172;
  assign n7175 = ~n7173 & ~n7174;
  assign n7176 = ~n7170 & ~n7175;
  assign n7177 = ~n7169 & ~n7176;
  assign n7178 = po45  & ~n7177;
  assign n7179 = ~po45  & n7177;
  assign n7180 = ~n6814 & ~n6815;
  assign n7181 = po25  & n7180;
  assign n7182 = ~n6820 & ~n7181;
  assign n7183 = n6820 & n7181;
  assign n7184 = ~n7182 & ~n7183;
  assign n7185 = ~n7179 & ~n7184;
  assign n7186 = ~n7178 & ~n7185;
  assign n7187 = po46  & ~n7186;
  assign n7188 = ~po46  & n7186;
  assign n7189 = ~n6823 & ~n6824;
  assign n7190 = po25  & n7189;
  assign n7191 = ~n6829 & ~n7190;
  assign n7192 = n6829 & n7190;
  assign n7193 = ~n7191 & ~n7192;
  assign n7194 = ~n7188 & ~n7193;
  assign n7195 = ~n7187 & ~n7194;
  assign n7196 = po47  & ~n7195;
  assign n7197 = ~po47  & n7195;
  assign n7198 = ~n6832 & ~n6833;
  assign n7199 = po25  & n7198;
  assign n7200 = ~n6838 & ~n7199;
  assign n7201 = n6838 & n7199;
  assign n7202 = ~n7200 & ~n7201;
  assign n7203 = ~n7197 & ~n7202;
  assign n7204 = ~n7196 & ~n7203;
  assign n7205 = po48  & ~n7204;
  assign n7206 = ~po48  & n7204;
  assign n7207 = ~n6841 & ~n6842;
  assign n7208 = po25  & n7207;
  assign n7209 = ~n6847 & ~n7208;
  assign n7210 = n6847 & n7208;
  assign n7211 = ~n7209 & ~n7210;
  assign n7212 = ~n7206 & ~n7211;
  assign n7213 = ~n7205 & ~n7212;
  assign n7214 = po49  & ~n7213;
  assign n7215 = ~po49  & n7213;
  assign n7216 = ~n6850 & ~n6851;
  assign n7217 = po25  & n7216;
  assign n7218 = ~n6856 & ~n7217;
  assign n7219 = n6856 & n7217;
  assign n7220 = ~n7218 & ~n7219;
  assign n7221 = ~n7215 & ~n7220;
  assign n7222 = ~n7214 & ~n7221;
  assign n7223 = po50  & ~n7222;
  assign n7224 = ~po50  & n7222;
  assign n7225 = ~n6859 & ~n6860;
  assign n7226 = po25  & n7225;
  assign n7227 = ~n6865 & ~n7226;
  assign n7228 = n6865 & n7226;
  assign n7229 = ~n7227 & ~n7228;
  assign n7230 = ~n7224 & ~n7229;
  assign n7231 = ~n7223 & ~n7230;
  assign n7232 = po51  & ~n7231;
  assign n7233 = ~po51  & n7231;
  assign n7234 = ~n6868 & ~n6869;
  assign n7235 = po25  & n7234;
  assign n7236 = ~n6874 & ~n7235;
  assign n7237 = n6874 & n7235;
  assign n7238 = ~n7236 & ~n7237;
  assign n7239 = ~n7233 & ~n7238;
  assign n7240 = ~n7232 & ~n7239;
  assign n7241 = po52  & ~n7240;
  assign n7242 = ~po52  & n7240;
  assign n7243 = ~n6877 & ~n6878;
  assign n7244 = po25  & n7243;
  assign n7245 = ~n6883 & ~n7244;
  assign n7246 = n6883 & n7244;
  assign n7247 = ~n7245 & ~n7246;
  assign n7248 = ~n7242 & ~n7247;
  assign n7249 = ~n7241 & ~n7248;
  assign n7250 = po53  & ~n7249;
  assign n7251 = ~po53  & n7249;
  assign n7252 = ~n6886 & ~n6887;
  assign n7253 = po25  & n7252;
  assign n7254 = ~n6892 & ~n7253;
  assign n7255 = n6892 & n7253;
  assign n7256 = ~n7254 & ~n7255;
  assign n7257 = ~n7251 & ~n7256;
  assign n7258 = ~n7250 & ~n7257;
  assign n7259 = po54  & ~n7258;
  assign n7260 = ~po54  & n7258;
  assign n7261 = ~n6895 & ~n6896;
  assign n7262 = po25  & n7261;
  assign n7263 = ~n6901 & ~n7262;
  assign n7264 = n6901 & n7262;
  assign n7265 = ~n7263 & ~n7264;
  assign n7266 = ~n7260 & ~n7265;
  assign n7267 = ~n7259 & ~n7266;
  assign n7268 = po55  & ~n7267;
  assign n7269 = ~po55  & n7267;
  assign n7270 = ~n6904 & ~n6905;
  assign n7271 = po25  & n7270;
  assign n7272 = ~n6910 & ~n7271;
  assign n7273 = n6910 & n7271;
  assign n7274 = ~n7272 & ~n7273;
  assign n7275 = ~n7269 & ~n7274;
  assign n7276 = ~n7268 & ~n7275;
  assign n7277 = po56  & ~n7276;
  assign n7278 = ~po56  & n7276;
  assign n7279 = ~n6913 & ~n6914;
  assign n7280 = po25  & n7279;
  assign n7281 = ~n6919 & ~n7280;
  assign n7282 = n6919 & n7280;
  assign n7283 = ~n7281 & ~n7282;
  assign n7284 = ~n7278 & ~n7283;
  assign n7285 = ~n7277 & ~n7284;
  assign n7286 = po57  & ~n7285;
  assign n7287 = ~po57  & n7285;
  assign n7288 = ~n6922 & ~n6923;
  assign n7289 = po25  & n7288;
  assign n7290 = ~n6928 & ~n7289;
  assign n7291 = n6928 & n7289;
  assign n7292 = ~n7290 & ~n7291;
  assign n7293 = ~n7287 & ~n7292;
  assign n7294 = ~n7286 & ~n7293;
  assign n7295 = po58  & ~n7294;
  assign n7296 = ~po58  & n7294;
  assign n7297 = ~n6931 & ~n6932;
  assign n7298 = po25  & n7297;
  assign n7299 = ~n6937 & ~n7298;
  assign n7300 = n6937 & n7298;
  assign n7301 = ~n7299 & ~n7300;
  assign n7302 = ~n7296 & ~n7301;
  assign n7303 = ~n7295 & ~n7302;
  assign n7304 = po59  & ~n7303;
  assign n7305 = ~po59  & n7303;
  assign n7306 = ~n6940 & ~n6941;
  assign n7307 = po25  & n7306;
  assign n7308 = ~n6946 & ~n7307;
  assign n7309 = n6946 & n7307;
  assign n7310 = ~n7308 & ~n7309;
  assign n7311 = ~n7305 & ~n7310;
  assign n7312 = ~n7304 & ~n7311;
  assign n7313 = po60  & ~n7312;
  assign n7314 = ~po60  & n7312;
  assign n7315 = ~n6949 & ~n6950;
  assign n7316 = po25  & n7315;
  assign n7317 = ~n6955 & ~n7316;
  assign n7318 = n6955 & n7316;
  assign n7319 = ~n7317 & ~n7318;
  assign n7320 = ~n7314 & ~n7319;
  assign n7321 = ~n7313 & ~n7320;
  assign n7322 = po61  & ~n7321;
  assign n7323 = ~po61  & n7321;
  assign n7324 = ~n6958 & ~n6959;
  assign n7325 = po25  & n7324;
  assign n7326 = ~n6964 & ~n7325;
  assign n7327 = n6964 & n7325;
  assign n7328 = ~n7326 & ~n7327;
  assign n7329 = ~n7323 & ~n7328;
  assign n7330 = ~n7322 & ~n7329;
  assign n7331 = po62  & ~n7330;
  assign n7332 = ~po62  & n7330;
  assign n7333 = ~n6967 & ~n6968;
  assign n7334 = po25  & n7333;
  assign n7335 = ~n6973 & ~n7334;
  assign n7336 = n6973 & n7334;
  assign n7337 = ~n7335 & ~n7336;
  assign n7338 = ~n7332 & ~n7337;
  assign n7339 = ~n7331 & ~n7338;
  assign n7340 = n7130 & n7339;
  assign n7341 = ~n7130 & ~n7339;
  assign n7342 = n6986 & po25 ;
  assign n7343 = ~n6985 & ~n7342;
  assign n7344 = n7341 & n7343;
  assign n7345 = ~po63  & ~n7344;
  assign n7346 = ~n6766 & po25 ;
  assign n7347 = n6984 & ~n7346;
  assign n7348 = po63  & ~n6986;
  assign n7349 = ~n7347 & n7348;
  assign n7350 = ~n7340 & ~n7349;
  assign n7351 = ~n7345 & n7350;
  assign po24  = n7125 | ~n7351;
  assign n7353 = ~n7123 & ~n7124;
  assign n7354 = po24  & n7353;
  assign n7355 = ~n7002 & ~n7354;
  assign n7356 = n7002 & n7354;
  assign n7357 = ~n7355 & ~n7356;
  assign n7358 = pi48  & po24 ;
  assign n7359 = ~pi46  & ~pi47 ;
  assign n7360 = ~pi48  & n7359;
  assign n7361 = ~n7358 & ~n7360;
  assign n7362 = po25  & ~n7361;
  assign n7363 = ~po25  & n7361;
  assign n7364 = ~pi48  & po24 ;
  assign n7365 = pi49  & ~n7364;
  assign n7366 = ~pi49  & n7364;
  assign n7367 = ~n7365 & ~n7366;
  assign n7368 = ~n7363 & n7367;
  assign n7369 = ~n7362 & ~n7368;
  assign n7370 = po26  & ~n7369;
  assign n7371 = ~po26  & n7369;
  assign n7372 = po25  & n7351;
  assign n7373 = ~n7366 & ~n7372;
  assign n7374 = pi50  & ~n7373;
  assign n7375 = ~pi50  & n7373;
  assign n7376 = ~n7374 & ~n7375;
  assign n7377 = ~n7371 & ~n7376;
  assign n7378 = ~n7370 & ~n7377;
  assign n7379 = po27  & ~n7378;
  assign n7380 = ~po27  & n7378;
  assign n7381 = ~n7007 & ~n7008;
  assign n7382 = po24  & n7381;
  assign n7383 = n7012 & ~n7382;
  assign n7384 = ~n7012 & n7382;
  assign n7385 = ~n7383 & ~n7384;
  assign n7386 = ~n7380 & ~n7385;
  assign n7387 = ~n7379 & ~n7386;
  assign n7388 = po28  & ~n7387;
  assign n7389 = ~po28  & n7387;
  assign n7390 = ~n7015 & ~n7016;
  assign n7391 = po24  & n7390;
  assign n7392 = ~n7021 & ~n7391;
  assign n7393 = n7021 & n7391;
  assign n7394 = ~n7392 & ~n7393;
  assign n7395 = ~n7389 & ~n7394;
  assign n7396 = ~n7388 & ~n7395;
  assign n7397 = po29  & ~n7396;
  assign n7398 = ~po29  & n7396;
  assign n7399 = ~n7024 & ~n7025;
  assign n7400 = po24  & n7399;
  assign n7401 = n7030 & n7400;
  assign n7402 = ~n7030 & ~n7400;
  assign n7403 = ~n7401 & ~n7402;
  assign n7404 = ~n7398 & ~n7403;
  assign n7405 = ~n7397 & ~n7404;
  assign n7406 = po30  & ~n7405;
  assign n7407 = ~po30  & n7405;
  assign n7408 = ~n7033 & ~n7034;
  assign n7409 = po24  & n7408;
  assign n7410 = ~n7039 & ~n7409;
  assign n7411 = n7039 & n7409;
  assign n7412 = ~n7410 & ~n7411;
  assign n7413 = ~n7407 & ~n7412;
  assign n7414 = ~n7406 & ~n7413;
  assign n7415 = po31  & ~n7414;
  assign n7416 = ~po31  & n7414;
  assign n7417 = ~n7042 & ~n7043;
  assign n7418 = po24  & n7417;
  assign n7419 = ~n7048 & ~n7418;
  assign n7420 = n7048 & n7418;
  assign n7421 = ~n7419 & ~n7420;
  assign n7422 = ~n7416 & ~n7421;
  assign n7423 = ~n7415 & ~n7422;
  assign n7424 = po32  & ~n7423;
  assign n7425 = ~po32  & n7423;
  assign n7426 = ~n7051 & ~n7052;
  assign n7427 = po24  & n7426;
  assign n7428 = ~n7057 & ~n7427;
  assign n7429 = n7057 & n7427;
  assign n7430 = ~n7428 & ~n7429;
  assign n7431 = ~n7425 & ~n7430;
  assign n7432 = ~n7424 & ~n7431;
  assign n7433 = po33  & ~n7432;
  assign n7434 = ~po33  & n7432;
  assign n7435 = ~n7060 & ~n7061;
  assign n7436 = po24  & n7435;
  assign n7437 = ~n7066 & ~n7436;
  assign n7438 = n7066 & n7436;
  assign n7439 = ~n7437 & ~n7438;
  assign n7440 = ~n7434 & ~n7439;
  assign n7441 = ~n7433 & ~n7440;
  assign n7442 = po34  & ~n7441;
  assign n7443 = ~po34  & n7441;
  assign n7444 = ~n7069 & ~n7070;
  assign n7445 = po24  & n7444;
  assign n7446 = ~n7075 & ~n7445;
  assign n7447 = n7075 & n7445;
  assign n7448 = ~n7446 & ~n7447;
  assign n7449 = ~n7443 & ~n7448;
  assign n7450 = ~n7442 & ~n7449;
  assign n7451 = po35  & ~n7450;
  assign n7452 = ~po35  & n7450;
  assign n7453 = ~n7078 & ~n7079;
  assign n7454 = po24  & n7453;
  assign n7455 = ~n7084 & ~n7454;
  assign n7456 = n7084 & n7454;
  assign n7457 = ~n7455 & ~n7456;
  assign n7458 = ~n7452 & ~n7457;
  assign n7459 = ~n7451 & ~n7458;
  assign n7460 = po36  & ~n7459;
  assign n7461 = ~po36  & n7459;
  assign n7462 = ~n7087 & ~n7088;
  assign n7463 = po24  & n7462;
  assign n7464 = ~n7093 & ~n7463;
  assign n7465 = n7093 & n7463;
  assign n7466 = ~n7464 & ~n7465;
  assign n7467 = ~n7461 & ~n7466;
  assign n7468 = ~n7460 & ~n7467;
  assign n7469 = po37  & ~n7468;
  assign n7470 = ~po37  & n7468;
  assign n7471 = ~n7096 & ~n7097;
  assign n7472 = po24  & n7471;
  assign n7473 = ~n7102 & ~n7472;
  assign n7474 = n7102 & n7472;
  assign n7475 = ~n7473 & ~n7474;
  assign n7476 = ~n7470 & ~n7475;
  assign n7477 = ~n7469 & ~n7476;
  assign n7478 = po38  & ~n7477;
  assign n7479 = ~po38  & n7477;
  assign n7480 = ~n7105 & ~n7106;
  assign n7481 = po24  & n7480;
  assign n7482 = ~n7111 & ~n7481;
  assign n7483 = n7111 & n7481;
  assign n7484 = ~n7482 & ~n7483;
  assign n7485 = ~n7479 & ~n7484;
  assign n7486 = ~n7478 & ~n7485;
  assign n7487 = po39  & ~n7486;
  assign n7488 = ~n7114 & ~n7120;
  assign n7489 = po24  & n7488;
  assign n7490 = ~n7119 & ~n7489;
  assign n7491 = n7119 & n7489;
  assign n7492 = ~n7490 & ~n7491;
  assign n7493 = ~po39  & n7486;
  assign n7494 = ~n7492 & ~n7493;
  assign n7495 = ~n7487 & ~n7494;
  assign n7496 = po40  & ~n7495;
  assign n7497 = ~po40  & n7495;
  assign n7498 = n7130 & ~po24 ;
  assign n7499 = ~n7331 & ~n7332;
  assign n7500 = po24  & n7499;
  assign n7501 = ~n7337 & ~n7500;
  assign n7502 = n7337 & n7500;
  assign n7503 = ~n7501 & ~n7502;
  assign n7504 = ~n7357 & ~n7497;
  assign n7505 = ~n7496 & ~n7504;
  assign n7506 = po41  & ~n7505;
  assign n7507 = ~po41  & n7505;
  assign n7508 = ~n7133 & ~n7134;
  assign n7509 = po24  & n7508;
  assign n7510 = ~n7139 & ~n7509;
  assign n7511 = n7139 & n7509;
  assign n7512 = ~n7510 & ~n7511;
  assign n7513 = ~n7507 & ~n7512;
  assign n7514 = ~n7506 & ~n7513;
  assign n7515 = po42  & ~n7514;
  assign n7516 = ~po42  & n7514;
  assign n7517 = ~n7142 & ~n7143;
  assign n7518 = po24  & n7517;
  assign n7519 = ~n7148 & ~n7518;
  assign n7520 = n7148 & n7518;
  assign n7521 = ~n7519 & ~n7520;
  assign n7522 = ~n7516 & ~n7521;
  assign n7523 = ~n7515 & ~n7522;
  assign n7524 = po43  & ~n7523;
  assign n7525 = ~po43  & n7523;
  assign n7526 = ~n7151 & ~n7152;
  assign n7527 = po24  & n7526;
  assign n7528 = ~n7157 & ~n7527;
  assign n7529 = n7157 & n7527;
  assign n7530 = ~n7528 & ~n7529;
  assign n7531 = ~n7525 & ~n7530;
  assign n7532 = ~n7524 & ~n7531;
  assign n7533 = po44  & ~n7532;
  assign n7534 = ~po44  & n7532;
  assign n7535 = ~n7160 & ~n7161;
  assign n7536 = po24  & n7535;
  assign n7537 = ~n7166 & ~n7536;
  assign n7538 = n7166 & n7536;
  assign n7539 = ~n7537 & ~n7538;
  assign n7540 = ~n7534 & ~n7539;
  assign n7541 = ~n7533 & ~n7540;
  assign n7542 = po45  & ~n7541;
  assign n7543 = ~po45  & n7541;
  assign n7544 = ~n7169 & ~n7170;
  assign n7545 = po24  & n7544;
  assign n7546 = ~n7175 & ~n7545;
  assign n7547 = n7175 & n7545;
  assign n7548 = ~n7546 & ~n7547;
  assign n7549 = ~n7543 & ~n7548;
  assign n7550 = ~n7542 & ~n7549;
  assign n7551 = po46  & ~n7550;
  assign n7552 = ~po46  & n7550;
  assign n7553 = ~n7178 & ~n7179;
  assign n7554 = po24  & n7553;
  assign n7555 = ~n7184 & ~n7554;
  assign n7556 = n7184 & n7554;
  assign n7557 = ~n7555 & ~n7556;
  assign n7558 = ~n7552 & ~n7557;
  assign n7559 = ~n7551 & ~n7558;
  assign n7560 = po47  & ~n7559;
  assign n7561 = ~po47  & n7559;
  assign n7562 = ~n7187 & ~n7188;
  assign n7563 = po24  & n7562;
  assign n7564 = ~n7193 & ~n7563;
  assign n7565 = n7193 & n7563;
  assign n7566 = ~n7564 & ~n7565;
  assign n7567 = ~n7561 & ~n7566;
  assign n7568 = ~n7560 & ~n7567;
  assign n7569 = po48  & ~n7568;
  assign n7570 = ~po48  & n7568;
  assign n7571 = ~n7196 & ~n7197;
  assign n7572 = po24  & n7571;
  assign n7573 = ~n7202 & ~n7572;
  assign n7574 = n7202 & n7572;
  assign n7575 = ~n7573 & ~n7574;
  assign n7576 = ~n7570 & ~n7575;
  assign n7577 = ~n7569 & ~n7576;
  assign n7578 = po49  & ~n7577;
  assign n7579 = ~po49  & n7577;
  assign n7580 = ~n7205 & ~n7206;
  assign n7581 = po24  & n7580;
  assign n7582 = ~n7211 & ~n7581;
  assign n7583 = n7211 & n7581;
  assign n7584 = ~n7582 & ~n7583;
  assign n7585 = ~n7579 & ~n7584;
  assign n7586 = ~n7578 & ~n7585;
  assign n7587 = po50  & ~n7586;
  assign n7588 = ~po50  & n7586;
  assign n7589 = ~n7214 & ~n7215;
  assign n7590 = po24  & n7589;
  assign n7591 = ~n7220 & ~n7590;
  assign n7592 = n7220 & n7590;
  assign n7593 = ~n7591 & ~n7592;
  assign n7594 = ~n7588 & ~n7593;
  assign n7595 = ~n7587 & ~n7594;
  assign n7596 = po51  & ~n7595;
  assign n7597 = ~po51  & n7595;
  assign n7598 = ~n7223 & ~n7224;
  assign n7599 = po24  & n7598;
  assign n7600 = ~n7229 & ~n7599;
  assign n7601 = n7229 & n7599;
  assign n7602 = ~n7600 & ~n7601;
  assign n7603 = ~n7597 & ~n7602;
  assign n7604 = ~n7596 & ~n7603;
  assign n7605 = po52  & ~n7604;
  assign n7606 = ~po52  & n7604;
  assign n7607 = ~n7232 & ~n7233;
  assign n7608 = po24  & n7607;
  assign n7609 = ~n7238 & ~n7608;
  assign n7610 = n7238 & n7608;
  assign n7611 = ~n7609 & ~n7610;
  assign n7612 = ~n7606 & ~n7611;
  assign n7613 = ~n7605 & ~n7612;
  assign n7614 = po53  & ~n7613;
  assign n7615 = ~po53  & n7613;
  assign n7616 = ~n7241 & ~n7242;
  assign n7617 = po24  & n7616;
  assign n7618 = ~n7247 & ~n7617;
  assign n7619 = n7247 & n7617;
  assign n7620 = ~n7618 & ~n7619;
  assign n7621 = ~n7615 & ~n7620;
  assign n7622 = ~n7614 & ~n7621;
  assign n7623 = po54  & ~n7622;
  assign n7624 = ~po54  & n7622;
  assign n7625 = ~n7250 & ~n7251;
  assign n7626 = po24  & n7625;
  assign n7627 = ~n7256 & ~n7626;
  assign n7628 = n7256 & n7626;
  assign n7629 = ~n7627 & ~n7628;
  assign n7630 = ~n7624 & ~n7629;
  assign n7631 = ~n7623 & ~n7630;
  assign n7632 = po55  & ~n7631;
  assign n7633 = ~po55  & n7631;
  assign n7634 = ~n7259 & ~n7260;
  assign n7635 = po24  & n7634;
  assign n7636 = ~n7265 & ~n7635;
  assign n7637 = n7265 & n7635;
  assign n7638 = ~n7636 & ~n7637;
  assign n7639 = ~n7633 & ~n7638;
  assign n7640 = ~n7632 & ~n7639;
  assign n7641 = po56  & ~n7640;
  assign n7642 = ~po56  & n7640;
  assign n7643 = ~n7268 & ~n7269;
  assign n7644 = po24  & n7643;
  assign n7645 = ~n7274 & ~n7644;
  assign n7646 = n7274 & n7644;
  assign n7647 = ~n7645 & ~n7646;
  assign n7648 = ~n7642 & ~n7647;
  assign n7649 = ~n7641 & ~n7648;
  assign n7650 = po57  & ~n7649;
  assign n7651 = ~po57  & n7649;
  assign n7652 = ~n7277 & ~n7278;
  assign n7653 = po24  & n7652;
  assign n7654 = ~n7283 & ~n7653;
  assign n7655 = n7283 & n7653;
  assign n7656 = ~n7654 & ~n7655;
  assign n7657 = ~n7651 & ~n7656;
  assign n7658 = ~n7650 & ~n7657;
  assign n7659 = po58  & ~n7658;
  assign n7660 = ~po58  & n7658;
  assign n7661 = ~n7286 & ~n7287;
  assign n7662 = po24  & n7661;
  assign n7663 = ~n7292 & ~n7662;
  assign n7664 = n7292 & n7662;
  assign n7665 = ~n7663 & ~n7664;
  assign n7666 = ~n7660 & ~n7665;
  assign n7667 = ~n7659 & ~n7666;
  assign n7668 = po59  & ~n7667;
  assign n7669 = ~po59  & n7667;
  assign n7670 = ~n7295 & ~n7296;
  assign n7671 = po24  & n7670;
  assign n7672 = ~n7301 & ~n7671;
  assign n7673 = n7301 & n7671;
  assign n7674 = ~n7672 & ~n7673;
  assign n7675 = ~n7669 & ~n7674;
  assign n7676 = ~n7668 & ~n7675;
  assign n7677 = po60  & ~n7676;
  assign n7678 = ~po60  & n7676;
  assign n7679 = ~n7304 & ~n7305;
  assign n7680 = po24  & n7679;
  assign n7681 = ~n7310 & ~n7680;
  assign n7682 = n7310 & n7680;
  assign n7683 = ~n7681 & ~n7682;
  assign n7684 = ~n7678 & ~n7683;
  assign n7685 = ~n7677 & ~n7684;
  assign n7686 = po61  & ~n7685;
  assign n7687 = ~po61  & n7685;
  assign n7688 = ~n7313 & ~n7314;
  assign n7689 = po24  & n7688;
  assign n7690 = ~n7319 & ~n7689;
  assign n7691 = n7319 & n7689;
  assign n7692 = ~n7690 & ~n7691;
  assign n7693 = ~n7687 & ~n7692;
  assign n7694 = ~n7686 & ~n7693;
  assign n7695 = po62  & ~n7694;
  assign n7696 = ~po62  & n7694;
  assign n7697 = ~n7322 & ~n7323;
  assign n7698 = po24  & n7697;
  assign n7699 = ~n7328 & ~n7698;
  assign n7700 = n7328 & n7698;
  assign n7701 = ~n7699 & ~n7700;
  assign n7702 = ~n7696 & ~n7701;
  assign n7703 = ~n7695 & ~n7702;
  assign n7704 = n7503 & n7703;
  assign n7705 = ~n7503 & ~n7703;
  assign n7706 = n7341 & po24 ;
  assign n7707 = ~n7340 & ~n7706;
  assign n7708 = n7705 & n7707;
  assign n7709 = ~po63  & ~n7708;
  assign n7710 = ~n7130 & po24 ;
  assign n7711 = n7339 & ~n7710;
  assign n7712 = po63  & ~n7341;
  assign n7713 = ~n7711 & n7712;
  assign n7714 = ~n7704 & ~n7713;
  assign n7715 = ~n7709 & n7714;
  assign po23  = n7498 | ~n7715;
  assign n7717 = ~n7496 & ~n7497;
  assign n7718 = po23  & n7717;
  assign n7719 = ~n7357 & ~n7718;
  assign n7720 = n7357 & n7718;
  assign n7721 = ~n7719 & ~n7720;
  assign n7722 = pi46  & po23 ;
  assign n7723 = ~pi44  & ~pi45 ;
  assign n7724 = ~pi46  & n7723;
  assign n7725 = ~n7722 & ~n7724;
  assign n7726 = po24  & ~n7725;
  assign n7727 = ~po24  & n7725;
  assign n7728 = ~pi46  & po23 ;
  assign n7729 = pi47  & ~n7728;
  assign n7730 = ~pi47  & n7728;
  assign n7731 = ~n7729 & ~n7730;
  assign n7732 = ~n7727 & n7731;
  assign n7733 = ~n7726 & ~n7732;
  assign n7734 = po25  & ~n7733;
  assign n7735 = ~po25  & n7733;
  assign n7736 = po24  & n7715;
  assign n7737 = ~n7730 & ~n7736;
  assign n7738 = pi48  & ~n7737;
  assign n7739 = ~pi48  & n7737;
  assign n7740 = ~n7738 & ~n7739;
  assign n7741 = ~n7735 & ~n7740;
  assign n7742 = ~n7734 & ~n7741;
  assign n7743 = po26  & ~n7742;
  assign n7744 = ~po26  & n7742;
  assign n7745 = ~n7362 & ~n7363;
  assign n7746 = po23  & n7745;
  assign n7747 = n7367 & ~n7746;
  assign n7748 = ~n7367 & n7746;
  assign n7749 = ~n7747 & ~n7748;
  assign n7750 = ~n7744 & ~n7749;
  assign n7751 = ~n7743 & ~n7750;
  assign n7752 = po27  & ~n7751;
  assign n7753 = ~po27  & n7751;
  assign n7754 = ~n7370 & ~n7371;
  assign n7755 = po23  & n7754;
  assign n7756 = ~n7376 & ~n7755;
  assign n7757 = n7376 & n7755;
  assign n7758 = ~n7756 & ~n7757;
  assign n7759 = ~n7753 & ~n7758;
  assign n7760 = ~n7752 & ~n7759;
  assign n7761 = po28  & ~n7760;
  assign n7762 = ~po28  & n7760;
  assign n7763 = ~n7379 & ~n7380;
  assign n7764 = po23  & n7763;
  assign n7765 = n7385 & n7764;
  assign n7766 = ~n7385 & ~n7764;
  assign n7767 = ~n7765 & ~n7766;
  assign n7768 = ~n7762 & ~n7767;
  assign n7769 = ~n7761 & ~n7768;
  assign n7770 = po29  & ~n7769;
  assign n7771 = ~po29  & n7769;
  assign n7772 = ~n7388 & ~n7389;
  assign n7773 = po23  & n7772;
  assign n7774 = ~n7394 & ~n7773;
  assign n7775 = n7394 & n7773;
  assign n7776 = ~n7774 & ~n7775;
  assign n7777 = ~n7771 & ~n7776;
  assign n7778 = ~n7770 & ~n7777;
  assign n7779 = po30  & ~n7778;
  assign n7780 = ~po30  & n7778;
  assign n7781 = ~n7397 & ~n7398;
  assign n7782 = po23  & n7781;
  assign n7783 = ~n7403 & ~n7782;
  assign n7784 = n7403 & n7782;
  assign n7785 = ~n7783 & ~n7784;
  assign n7786 = ~n7780 & ~n7785;
  assign n7787 = ~n7779 & ~n7786;
  assign n7788 = po31  & ~n7787;
  assign n7789 = ~po31  & n7787;
  assign n7790 = ~n7406 & ~n7407;
  assign n7791 = po23  & n7790;
  assign n7792 = ~n7412 & ~n7791;
  assign n7793 = n7412 & n7791;
  assign n7794 = ~n7792 & ~n7793;
  assign n7795 = ~n7789 & ~n7794;
  assign n7796 = ~n7788 & ~n7795;
  assign n7797 = po32  & ~n7796;
  assign n7798 = ~po32  & n7796;
  assign n7799 = ~n7415 & ~n7416;
  assign n7800 = po23  & n7799;
  assign n7801 = ~n7421 & ~n7800;
  assign n7802 = n7421 & n7800;
  assign n7803 = ~n7801 & ~n7802;
  assign n7804 = ~n7798 & ~n7803;
  assign n7805 = ~n7797 & ~n7804;
  assign n7806 = po33  & ~n7805;
  assign n7807 = ~po33  & n7805;
  assign n7808 = ~n7424 & ~n7425;
  assign n7809 = po23  & n7808;
  assign n7810 = ~n7430 & ~n7809;
  assign n7811 = n7430 & n7809;
  assign n7812 = ~n7810 & ~n7811;
  assign n7813 = ~n7807 & ~n7812;
  assign n7814 = ~n7806 & ~n7813;
  assign n7815 = po34  & ~n7814;
  assign n7816 = ~po34  & n7814;
  assign n7817 = ~n7433 & ~n7434;
  assign n7818 = po23  & n7817;
  assign n7819 = ~n7439 & ~n7818;
  assign n7820 = n7439 & n7818;
  assign n7821 = ~n7819 & ~n7820;
  assign n7822 = ~n7816 & ~n7821;
  assign n7823 = ~n7815 & ~n7822;
  assign n7824 = po35  & ~n7823;
  assign n7825 = ~po35  & n7823;
  assign n7826 = ~n7442 & ~n7443;
  assign n7827 = po23  & n7826;
  assign n7828 = ~n7448 & ~n7827;
  assign n7829 = n7448 & n7827;
  assign n7830 = ~n7828 & ~n7829;
  assign n7831 = ~n7825 & ~n7830;
  assign n7832 = ~n7824 & ~n7831;
  assign n7833 = po36  & ~n7832;
  assign n7834 = ~po36  & n7832;
  assign n7835 = ~n7451 & ~n7452;
  assign n7836 = po23  & n7835;
  assign n7837 = ~n7457 & ~n7836;
  assign n7838 = n7457 & n7836;
  assign n7839 = ~n7837 & ~n7838;
  assign n7840 = ~n7834 & ~n7839;
  assign n7841 = ~n7833 & ~n7840;
  assign n7842 = po37  & ~n7841;
  assign n7843 = ~po37  & n7841;
  assign n7844 = ~n7460 & ~n7461;
  assign n7845 = po23  & n7844;
  assign n7846 = ~n7466 & ~n7845;
  assign n7847 = n7466 & n7845;
  assign n7848 = ~n7846 & ~n7847;
  assign n7849 = ~n7843 & ~n7848;
  assign n7850 = ~n7842 & ~n7849;
  assign n7851 = po38  & ~n7850;
  assign n7852 = ~po38  & n7850;
  assign n7853 = ~n7469 & ~n7470;
  assign n7854 = po23  & n7853;
  assign n7855 = ~n7475 & ~n7854;
  assign n7856 = n7475 & n7854;
  assign n7857 = ~n7855 & ~n7856;
  assign n7858 = ~n7852 & ~n7857;
  assign n7859 = ~n7851 & ~n7858;
  assign n7860 = po39  & ~n7859;
  assign n7861 = ~po39  & n7859;
  assign n7862 = ~n7478 & ~n7479;
  assign n7863 = po23  & n7862;
  assign n7864 = ~n7484 & ~n7863;
  assign n7865 = n7484 & n7863;
  assign n7866 = ~n7864 & ~n7865;
  assign n7867 = ~n7861 & ~n7866;
  assign n7868 = ~n7860 & ~n7867;
  assign n7869 = po40  & ~n7868;
  assign n7870 = ~n7487 & ~n7493;
  assign n7871 = po23  & n7870;
  assign n7872 = ~n7492 & ~n7871;
  assign n7873 = n7492 & n7871;
  assign n7874 = ~n7872 & ~n7873;
  assign n7875 = ~po40  & n7868;
  assign n7876 = ~n7874 & ~n7875;
  assign n7877 = ~n7869 & ~n7876;
  assign n7878 = po41  & ~n7877;
  assign n7879 = ~po41  & n7877;
  assign n7880 = n7503 & ~po23 ;
  assign n7881 = ~n7695 & ~n7696;
  assign n7882 = po23  & n7881;
  assign n7883 = ~n7701 & ~n7882;
  assign n7884 = n7701 & n7882;
  assign n7885 = ~n7883 & ~n7884;
  assign n7886 = ~n7721 & ~n7879;
  assign n7887 = ~n7878 & ~n7886;
  assign n7888 = po42  & ~n7887;
  assign n7889 = ~po42  & n7887;
  assign n7890 = ~n7506 & ~n7507;
  assign n7891 = po23  & n7890;
  assign n7892 = ~n7512 & ~n7891;
  assign n7893 = n7512 & n7891;
  assign n7894 = ~n7892 & ~n7893;
  assign n7895 = ~n7889 & ~n7894;
  assign n7896 = ~n7888 & ~n7895;
  assign n7897 = po43  & ~n7896;
  assign n7898 = ~po43  & n7896;
  assign n7899 = ~n7515 & ~n7516;
  assign n7900 = po23  & n7899;
  assign n7901 = ~n7521 & ~n7900;
  assign n7902 = n7521 & n7900;
  assign n7903 = ~n7901 & ~n7902;
  assign n7904 = ~n7898 & ~n7903;
  assign n7905 = ~n7897 & ~n7904;
  assign n7906 = po44  & ~n7905;
  assign n7907 = ~po44  & n7905;
  assign n7908 = ~n7524 & ~n7525;
  assign n7909 = po23  & n7908;
  assign n7910 = ~n7530 & ~n7909;
  assign n7911 = n7530 & n7909;
  assign n7912 = ~n7910 & ~n7911;
  assign n7913 = ~n7907 & ~n7912;
  assign n7914 = ~n7906 & ~n7913;
  assign n7915 = po45  & ~n7914;
  assign n7916 = ~po45  & n7914;
  assign n7917 = ~n7533 & ~n7534;
  assign n7918 = po23  & n7917;
  assign n7919 = ~n7539 & ~n7918;
  assign n7920 = n7539 & n7918;
  assign n7921 = ~n7919 & ~n7920;
  assign n7922 = ~n7916 & ~n7921;
  assign n7923 = ~n7915 & ~n7922;
  assign n7924 = po46  & ~n7923;
  assign n7925 = ~po46  & n7923;
  assign n7926 = ~n7542 & ~n7543;
  assign n7927 = po23  & n7926;
  assign n7928 = ~n7548 & ~n7927;
  assign n7929 = n7548 & n7927;
  assign n7930 = ~n7928 & ~n7929;
  assign n7931 = ~n7925 & ~n7930;
  assign n7932 = ~n7924 & ~n7931;
  assign n7933 = po47  & ~n7932;
  assign n7934 = ~po47  & n7932;
  assign n7935 = ~n7551 & ~n7552;
  assign n7936 = po23  & n7935;
  assign n7937 = ~n7557 & ~n7936;
  assign n7938 = n7557 & n7936;
  assign n7939 = ~n7937 & ~n7938;
  assign n7940 = ~n7934 & ~n7939;
  assign n7941 = ~n7933 & ~n7940;
  assign n7942 = po48  & ~n7941;
  assign n7943 = ~po48  & n7941;
  assign n7944 = ~n7560 & ~n7561;
  assign n7945 = po23  & n7944;
  assign n7946 = ~n7566 & ~n7945;
  assign n7947 = n7566 & n7945;
  assign n7948 = ~n7946 & ~n7947;
  assign n7949 = ~n7943 & ~n7948;
  assign n7950 = ~n7942 & ~n7949;
  assign n7951 = po49  & ~n7950;
  assign n7952 = ~po49  & n7950;
  assign n7953 = ~n7569 & ~n7570;
  assign n7954 = po23  & n7953;
  assign n7955 = ~n7575 & ~n7954;
  assign n7956 = n7575 & n7954;
  assign n7957 = ~n7955 & ~n7956;
  assign n7958 = ~n7952 & ~n7957;
  assign n7959 = ~n7951 & ~n7958;
  assign n7960 = po50  & ~n7959;
  assign n7961 = ~po50  & n7959;
  assign n7962 = ~n7578 & ~n7579;
  assign n7963 = po23  & n7962;
  assign n7964 = ~n7584 & ~n7963;
  assign n7965 = n7584 & n7963;
  assign n7966 = ~n7964 & ~n7965;
  assign n7967 = ~n7961 & ~n7966;
  assign n7968 = ~n7960 & ~n7967;
  assign n7969 = po51  & ~n7968;
  assign n7970 = ~po51  & n7968;
  assign n7971 = ~n7587 & ~n7588;
  assign n7972 = po23  & n7971;
  assign n7973 = ~n7593 & ~n7972;
  assign n7974 = n7593 & n7972;
  assign n7975 = ~n7973 & ~n7974;
  assign n7976 = ~n7970 & ~n7975;
  assign n7977 = ~n7969 & ~n7976;
  assign n7978 = po52  & ~n7977;
  assign n7979 = ~po52  & n7977;
  assign n7980 = ~n7596 & ~n7597;
  assign n7981 = po23  & n7980;
  assign n7982 = ~n7602 & ~n7981;
  assign n7983 = n7602 & n7981;
  assign n7984 = ~n7982 & ~n7983;
  assign n7985 = ~n7979 & ~n7984;
  assign n7986 = ~n7978 & ~n7985;
  assign n7987 = po53  & ~n7986;
  assign n7988 = ~po53  & n7986;
  assign n7989 = ~n7605 & ~n7606;
  assign n7990 = po23  & n7989;
  assign n7991 = ~n7611 & ~n7990;
  assign n7992 = n7611 & n7990;
  assign n7993 = ~n7991 & ~n7992;
  assign n7994 = ~n7988 & ~n7993;
  assign n7995 = ~n7987 & ~n7994;
  assign n7996 = po54  & ~n7995;
  assign n7997 = ~po54  & n7995;
  assign n7998 = ~n7614 & ~n7615;
  assign n7999 = po23  & n7998;
  assign n8000 = ~n7620 & ~n7999;
  assign n8001 = n7620 & n7999;
  assign n8002 = ~n8000 & ~n8001;
  assign n8003 = ~n7997 & ~n8002;
  assign n8004 = ~n7996 & ~n8003;
  assign n8005 = po55  & ~n8004;
  assign n8006 = ~po55  & n8004;
  assign n8007 = ~n7623 & ~n7624;
  assign n8008 = po23  & n8007;
  assign n8009 = ~n7629 & ~n8008;
  assign n8010 = n7629 & n8008;
  assign n8011 = ~n8009 & ~n8010;
  assign n8012 = ~n8006 & ~n8011;
  assign n8013 = ~n8005 & ~n8012;
  assign n8014 = po56  & ~n8013;
  assign n8015 = ~po56  & n8013;
  assign n8016 = ~n7632 & ~n7633;
  assign n8017 = po23  & n8016;
  assign n8018 = ~n7638 & ~n8017;
  assign n8019 = n7638 & n8017;
  assign n8020 = ~n8018 & ~n8019;
  assign n8021 = ~n8015 & ~n8020;
  assign n8022 = ~n8014 & ~n8021;
  assign n8023 = po57  & ~n8022;
  assign n8024 = ~po57  & n8022;
  assign n8025 = ~n7641 & ~n7642;
  assign n8026 = po23  & n8025;
  assign n8027 = ~n7647 & ~n8026;
  assign n8028 = n7647 & n8026;
  assign n8029 = ~n8027 & ~n8028;
  assign n8030 = ~n8024 & ~n8029;
  assign n8031 = ~n8023 & ~n8030;
  assign n8032 = po58  & ~n8031;
  assign n8033 = ~po58  & n8031;
  assign n8034 = ~n7650 & ~n7651;
  assign n8035 = po23  & n8034;
  assign n8036 = ~n7656 & ~n8035;
  assign n8037 = n7656 & n8035;
  assign n8038 = ~n8036 & ~n8037;
  assign n8039 = ~n8033 & ~n8038;
  assign n8040 = ~n8032 & ~n8039;
  assign n8041 = po59  & ~n8040;
  assign n8042 = ~po59  & n8040;
  assign n8043 = ~n7659 & ~n7660;
  assign n8044 = po23  & n8043;
  assign n8045 = ~n7665 & ~n8044;
  assign n8046 = n7665 & n8044;
  assign n8047 = ~n8045 & ~n8046;
  assign n8048 = ~n8042 & ~n8047;
  assign n8049 = ~n8041 & ~n8048;
  assign n8050 = po60  & ~n8049;
  assign n8051 = ~po60  & n8049;
  assign n8052 = ~n7668 & ~n7669;
  assign n8053 = po23  & n8052;
  assign n8054 = ~n7674 & ~n8053;
  assign n8055 = n7674 & n8053;
  assign n8056 = ~n8054 & ~n8055;
  assign n8057 = ~n8051 & ~n8056;
  assign n8058 = ~n8050 & ~n8057;
  assign n8059 = po61  & ~n8058;
  assign n8060 = ~po61  & n8058;
  assign n8061 = ~n7677 & ~n7678;
  assign n8062 = po23  & n8061;
  assign n8063 = ~n7683 & ~n8062;
  assign n8064 = n7683 & n8062;
  assign n8065 = ~n8063 & ~n8064;
  assign n8066 = ~n8060 & ~n8065;
  assign n8067 = ~n8059 & ~n8066;
  assign n8068 = po62  & ~n8067;
  assign n8069 = ~po62  & n8067;
  assign n8070 = ~n7686 & ~n7687;
  assign n8071 = po23  & n8070;
  assign n8072 = ~n7692 & ~n8071;
  assign n8073 = n7692 & n8071;
  assign n8074 = ~n8072 & ~n8073;
  assign n8075 = ~n8069 & ~n8074;
  assign n8076 = ~n8068 & ~n8075;
  assign n8077 = n7885 & n8076;
  assign n8078 = ~n7885 & ~n8076;
  assign n8079 = n7705 & po23 ;
  assign n8080 = ~n7704 & ~n8079;
  assign n8081 = n8078 & n8080;
  assign n8082 = ~po63  & ~n8081;
  assign n8083 = ~n7503 & po23 ;
  assign n8084 = n7703 & ~n8083;
  assign n8085 = po63  & ~n7705;
  assign n8086 = ~n8084 & n8085;
  assign n8087 = ~n8077 & ~n8086;
  assign n8088 = ~n8082 & n8087;
  assign po22  = n7880 | ~n8088;
  assign n8090 = ~n7878 & ~n7879;
  assign n8091 = po22  & n8090;
  assign n8092 = ~n7721 & ~n8091;
  assign n8093 = n7721 & n8091;
  assign n8094 = ~n8092 & ~n8093;
  assign n8095 = pi44  & po22 ;
  assign n8096 = ~pi42  & ~pi43 ;
  assign n8097 = ~pi44  & n8096;
  assign n8098 = ~n8095 & ~n8097;
  assign n8099 = po23  & ~n8098;
  assign n8100 = ~po23  & n8098;
  assign n8101 = ~pi44  & po22 ;
  assign n8102 = pi45  & ~n8101;
  assign n8103 = ~pi45  & n8101;
  assign n8104 = ~n8102 & ~n8103;
  assign n8105 = ~n8100 & n8104;
  assign n8106 = ~n8099 & ~n8105;
  assign n8107 = po24  & ~n8106;
  assign n8108 = ~po24  & n8106;
  assign n8109 = po23  & n8088;
  assign n8110 = ~n8103 & ~n8109;
  assign n8111 = pi46  & ~n8110;
  assign n8112 = ~pi46  & n8110;
  assign n8113 = ~n8111 & ~n8112;
  assign n8114 = ~n8108 & ~n8113;
  assign n8115 = ~n8107 & ~n8114;
  assign n8116 = po25  & ~n8115;
  assign n8117 = ~po25  & n8115;
  assign n8118 = ~n7726 & ~n7727;
  assign n8119 = po22  & n8118;
  assign n8120 = n7731 & ~n8119;
  assign n8121 = ~n7731 & n8119;
  assign n8122 = ~n8120 & ~n8121;
  assign n8123 = ~n8117 & ~n8122;
  assign n8124 = ~n8116 & ~n8123;
  assign n8125 = po26  & ~n8124;
  assign n8126 = ~po26  & n8124;
  assign n8127 = ~n7734 & ~n7735;
  assign n8128 = po22  & n8127;
  assign n8129 = ~n7740 & ~n8128;
  assign n8130 = n7740 & n8128;
  assign n8131 = ~n8129 & ~n8130;
  assign n8132 = ~n8126 & ~n8131;
  assign n8133 = ~n8125 & ~n8132;
  assign n8134 = po27  & ~n8133;
  assign n8135 = ~po27  & n8133;
  assign n8136 = ~n7743 & ~n7744;
  assign n8137 = po22  & n8136;
  assign n8138 = n7749 & n8137;
  assign n8139 = ~n7749 & ~n8137;
  assign n8140 = ~n8138 & ~n8139;
  assign n8141 = ~n8135 & ~n8140;
  assign n8142 = ~n8134 & ~n8141;
  assign n8143 = po28  & ~n8142;
  assign n8144 = ~po28  & n8142;
  assign n8145 = ~n7752 & ~n7753;
  assign n8146 = po22  & n8145;
  assign n8147 = ~n7758 & ~n8146;
  assign n8148 = n7758 & n8146;
  assign n8149 = ~n8147 & ~n8148;
  assign n8150 = ~n8144 & ~n8149;
  assign n8151 = ~n8143 & ~n8150;
  assign n8152 = po29  & ~n8151;
  assign n8153 = ~po29  & n8151;
  assign n8154 = ~n7761 & ~n7762;
  assign n8155 = po22  & n8154;
  assign n8156 = ~n7767 & ~n8155;
  assign n8157 = n7767 & n8155;
  assign n8158 = ~n8156 & ~n8157;
  assign n8159 = ~n8153 & ~n8158;
  assign n8160 = ~n8152 & ~n8159;
  assign n8161 = po30  & ~n8160;
  assign n8162 = ~po30  & n8160;
  assign n8163 = ~n7770 & ~n7771;
  assign n8164 = po22  & n8163;
  assign n8165 = ~n7776 & ~n8164;
  assign n8166 = n7776 & n8164;
  assign n8167 = ~n8165 & ~n8166;
  assign n8168 = ~n8162 & ~n8167;
  assign n8169 = ~n8161 & ~n8168;
  assign n8170 = po31  & ~n8169;
  assign n8171 = ~po31  & n8169;
  assign n8172 = ~n7779 & ~n7780;
  assign n8173 = po22  & n8172;
  assign n8174 = ~n7785 & ~n8173;
  assign n8175 = n7785 & n8173;
  assign n8176 = ~n8174 & ~n8175;
  assign n8177 = ~n8171 & ~n8176;
  assign n8178 = ~n8170 & ~n8177;
  assign n8179 = po32  & ~n8178;
  assign n8180 = ~po32  & n8178;
  assign n8181 = ~n7788 & ~n7789;
  assign n8182 = po22  & n8181;
  assign n8183 = ~n7794 & ~n8182;
  assign n8184 = n7794 & n8182;
  assign n8185 = ~n8183 & ~n8184;
  assign n8186 = ~n8180 & ~n8185;
  assign n8187 = ~n8179 & ~n8186;
  assign n8188 = po33  & ~n8187;
  assign n8189 = ~po33  & n8187;
  assign n8190 = ~n7797 & ~n7798;
  assign n8191 = po22  & n8190;
  assign n8192 = ~n7803 & ~n8191;
  assign n8193 = n7803 & n8191;
  assign n8194 = ~n8192 & ~n8193;
  assign n8195 = ~n8189 & ~n8194;
  assign n8196 = ~n8188 & ~n8195;
  assign n8197 = po34  & ~n8196;
  assign n8198 = ~po34  & n8196;
  assign n8199 = ~n7806 & ~n7807;
  assign n8200 = po22  & n8199;
  assign n8201 = ~n7812 & ~n8200;
  assign n8202 = n7812 & n8200;
  assign n8203 = ~n8201 & ~n8202;
  assign n8204 = ~n8198 & ~n8203;
  assign n8205 = ~n8197 & ~n8204;
  assign n8206 = po35  & ~n8205;
  assign n8207 = ~po35  & n8205;
  assign n8208 = ~n7815 & ~n7816;
  assign n8209 = po22  & n8208;
  assign n8210 = ~n7821 & ~n8209;
  assign n8211 = n7821 & n8209;
  assign n8212 = ~n8210 & ~n8211;
  assign n8213 = ~n8207 & ~n8212;
  assign n8214 = ~n8206 & ~n8213;
  assign n8215 = po36  & ~n8214;
  assign n8216 = ~po36  & n8214;
  assign n8217 = ~n7824 & ~n7825;
  assign n8218 = po22  & n8217;
  assign n8219 = ~n7830 & ~n8218;
  assign n8220 = n7830 & n8218;
  assign n8221 = ~n8219 & ~n8220;
  assign n8222 = ~n8216 & ~n8221;
  assign n8223 = ~n8215 & ~n8222;
  assign n8224 = po37  & ~n8223;
  assign n8225 = ~po37  & n8223;
  assign n8226 = ~n7833 & ~n7834;
  assign n8227 = po22  & n8226;
  assign n8228 = ~n7839 & ~n8227;
  assign n8229 = n7839 & n8227;
  assign n8230 = ~n8228 & ~n8229;
  assign n8231 = ~n8225 & ~n8230;
  assign n8232 = ~n8224 & ~n8231;
  assign n8233 = po38  & ~n8232;
  assign n8234 = ~po38  & n8232;
  assign n8235 = ~n7842 & ~n7843;
  assign n8236 = po22  & n8235;
  assign n8237 = ~n7848 & ~n8236;
  assign n8238 = n7848 & n8236;
  assign n8239 = ~n8237 & ~n8238;
  assign n8240 = ~n8234 & ~n8239;
  assign n8241 = ~n8233 & ~n8240;
  assign n8242 = po39  & ~n8241;
  assign n8243 = ~po39  & n8241;
  assign n8244 = ~n7851 & ~n7852;
  assign n8245 = po22  & n8244;
  assign n8246 = ~n7857 & ~n8245;
  assign n8247 = n7857 & n8245;
  assign n8248 = ~n8246 & ~n8247;
  assign n8249 = ~n8243 & ~n8248;
  assign n8250 = ~n8242 & ~n8249;
  assign n8251 = po40  & ~n8250;
  assign n8252 = ~po40  & n8250;
  assign n8253 = ~n7860 & ~n7861;
  assign n8254 = po22  & n8253;
  assign n8255 = ~n7866 & ~n8254;
  assign n8256 = n7866 & n8254;
  assign n8257 = ~n8255 & ~n8256;
  assign n8258 = ~n8252 & ~n8257;
  assign n8259 = ~n8251 & ~n8258;
  assign n8260 = po41  & ~n8259;
  assign n8261 = ~n7869 & ~n7875;
  assign n8262 = po22  & n8261;
  assign n8263 = ~n7874 & ~n8262;
  assign n8264 = n7874 & n8262;
  assign n8265 = ~n8263 & ~n8264;
  assign n8266 = ~po41  & n8259;
  assign n8267 = ~n8265 & ~n8266;
  assign n8268 = ~n8260 & ~n8267;
  assign n8269 = po42  & ~n8268;
  assign n8270 = ~po42  & n8268;
  assign n8271 = n7885 & ~po22 ;
  assign n8272 = ~n8068 & ~n8069;
  assign n8273 = po22  & n8272;
  assign n8274 = ~n8074 & ~n8273;
  assign n8275 = n8074 & n8273;
  assign n8276 = ~n8274 & ~n8275;
  assign n8277 = ~n8094 & ~n8270;
  assign n8278 = ~n8269 & ~n8277;
  assign n8279 = po43  & ~n8278;
  assign n8280 = ~po43  & n8278;
  assign n8281 = ~n7888 & ~n7889;
  assign n8282 = po22  & n8281;
  assign n8283 = ~n7894 & ~n8282;
  assign n8284 = n7894 & n8282;
  assign n8285 = ~n8283 & ~n8284;
  assign n8286 = ~n8280 & ~n8285;
  assign n8287 = ~n8279 & ~n8286;
  assign n8288 = po44  & ~n8287;
  assign n8289 = ~po44  & n8287;
  assign n8290 = ~n7897 & ~n7898;
  assign n8291 = po22  & n8290;
  assign n8292 = ~n7903 & ~n8291;
  assign n8293 = n7903 & n8291;
  assign n8294 = ~n8292 & ~n8293;
  assign n8295 = ~n8289 & ~n8294;
  assign n8296 = ~n8288 & ~n8295;
  assign n8297 = po45  & ~n8296;
  assign n8298 = ~po45  & n8296;
  assign n8299 = ~n7906 & ~n7907;
  assign n8300 = po22  & n8299;
  assign n8301 = ~n7912 & ~n8300;
  assign n8302 = n7912 & n8300;
  assign n8303 = ~n8301 & ~n8302;
  assign n8304 = ~n8298 & ~n8303;
  assign n8305 = ~n8297 & ~n8304;
  assign n8306 = po46  & ~n8305;
  assign n8307 = ~po46  & n8305;
  assign n8308 = ~n7915 & ~n7916;
  assign n8309 = po22  & n8308;
  assign n8310 = ~n7921 & ~n8309;
  assign n8311 = n7921 & n8309;
  assign n8312 = ~n8310 & ~n8311;
  assign n8313 = ~n8307 & ~n8312;
  assign n8314 = ~n8306 & ~n8313;
  assign n8315 = po47  & ~n8314;
  assign n8316 = ~po47  & n8314;
  assign n8317 = ~n7924 & ~n7925;
  assign n8318 = po22  & n8317;
  assign n8319 = ~n7930 & ~n8318;
  assign n8320 = n7930 & n8318;
  assign n8321 = ~n8319 & ~n8320;
  assign n8322 = ~n8316 & ~n8321;
  assign n8323 = ~n8315 & ~n8322;
  assign n8324 = po48  & ~n8323;
  assign n8325 = ~po48  & n8323;
  assign n8326 = ~n7933 & ~n7934;
  assign n8327 = po22  & n8326;
  assign n8328 = ~n7939 & ~n8327;
  assign n8329 = n7939 & n8327;
  assign n8330 = ~n8328 & ~n8329;
  assign n8331 = ~n8325 & ~n8330;
  assign n8332 = ~n8324 & ~n8331;
  assign n8333 = po49  & ~n8332;
  assign n8334 = ~po49  & n8332;
  assign n8335 = ~n7942 & ~n7943;
  assign n8336 = po22  & n8335;
  assign n8337 = ~n7948 & ~n8336;
  assign n8338 = n7948 & n8336;
  assign n8339 = ~n8337 & ~n8338;
  assign n8340 = ~n8334 & ~n8339;
  assign n8341 = ~n8333 & ~n8340;
  assign n8342 = po50  & ~n8341;
  assign n8343 = ~po50  & n8341;
  assign n8344 = ~n7951 & ~n7952;
  assign n8345 = po22  & n8344;
  assign n8346 = ~n7957 & ~n8345;
  assign n8347 = n7957 & n8345;
  assign n8348 = ~n8346 & ~n8347;
  assign n8349 = ~n8343 & ~n8348;
  assign n8350 = ~n8342 & ~n8349;
  assign n8351 = po51  & ~n8350;
  assign n8352 = ~po51  & n8350;
  assign n8353 = ~n7960 & ~n7961;
  assign n8354 = po22  & n8353;
  assign n8355 = ~n7966 & ~n8354;
  assign n8356 = n7966 & n8354;
  assign n8357 = ~n8355 & ~n8356;
  assign n8358 = ~n8352 & ~n8357;
  assign n8359 = ~n8351 & ~n8358;
  assign n8360 = po52  & ~n8359;
  assign n8361 = ~po52  & n8359;
  assign n8362 = ~n7969 & ~n7970;
  assign n8363 = po22  & n8362;
  assign n8364 = ~n7975 & ~n8363;
  assign n8365 = n7975 & n8363;
  assign n8366 = ~n8364 & ~n8365;
  assign n8367 = ~n8361 & ~n8366;
  assign n8368 = ~n8360 & ~n8367;
  assign n8369 = po53  & ~n8368;
  assign n8370 = ~po53  & n8368;
  assign n8371 = ~n7978 & ~n7979;
  assign n8372 = po22  & n8371;
  assign n8373 = ~n7984 & ~n8372;
  assign n8374 = n7984 & n8372;
  assign n8375 = ~n8373 & ~n8374;
  assign n8376 = ~n8370 & ~n8375;
  assign n8377 = ~n8369 & ~n8376;
  assign n8378 = po54  & ~n8377;
  assign n8379 = ~po54  & n8377;
  assign n8380 = ~n7987 & ~n7988;
  assign n8381 = po22  & n8380;
  assign n8382 = ~n7993 & ~n8381;
  assign n8383 = n7993 & n8381;
  assign n8384 = ~n8382 & ~n8383;
  assign n8385 = ~n8379 & ~n8384;
  assign n8386 = ~n8378 & ~n8385;
  assign n8387 = po55  & ~n8386;
  assign n8388 = ~po55  & n8386;
  assign n8389 = ~n7996 & ~n7997;
  assign n8390 = po22  & n8389;
  assign n8391 = ~n8002 & ~n8390;
  assign n8392 = n8002 & n8390;
  assign n8393 = ~n8391 & ~n8392;
  assign n8394 = ~n8388 & ~n8393;
  assign n8395 = ~n8387 & ~n8394;
  assign n8396 = po56  & ~n8395;
  assign n8397 = ~po56  & n8395;
  assign n8398 = ~n8005 & ~n8006;
  assign n8399 = po22  & n8398;
  assign n8400 = ~n8011 & ~n8399;
  assign n8401 = n8011 & n8399;
  assign n8402 = ~n8400 & ~n8401;
  assign n8403 = ~n8397 & ~n8402;
  assign n8404 = ~n8396 & ~n8403;
  assign n8405 = po57  & ~n8404;
  assign n8406 = ~po57  & n8404;
  assign n8407 = ~n8014 & ~n8015;
  assign n8408 = po22  & n8407;
  assign n8409 = ~n8020 & ~n8408;
  assign n8410 = n8020 & n8408;
  assign n8411 = ~n8409 & ~n8410;
  assign n8412 = ~n8406 & ~n8411;
  assign n8413 = ~n8405 & ~n8412;
  assign n8414 = po58  & ~n8413;
  assign n8415 = ~po58  & n8413;
  assign n8416 = ~n8023 & ~n8024;
  assign n8417 = po22  & n8416;
  assign n8418 = ~n8029 & ~n8417;
  assign n8419 = n8029 & n8417;
  assign n8420 = ~n8418 & ~n8419;
  assign n8421 = ~n8415 & ~n8420;
  assign n8422 = ~n8414 & ~n8421;
  assign n8423 = po59  & ~n8422;
  assign n8424 = ~po59  & n8422;
  assign n8425 = ~n8032 & ~n8033;
  assign n8426 = po22  & n8425;
  assign n8427 = ~n8038 & ~n8426;
  assign n8428 = n8038 & n8426;
  assign n8429 = ~n8427 & ~n8428;
  assign n8430 = ~n8424 & ~n8429;
  assign n8431 = ~n8423 & ~n8430;
  assign n8432 = po60  & ~n8431;
  assign n8433 = ~po60  & n8431;
  assign n8434 = ~n8041 & ~n8042;
  assign n8435 = po22  & n8434;
  assign n8436 = ~n8047 & ~n8435;
  assign n8437 = n8047 & n8435;
  assign n8438 = ~n8436 & ~n8437;
  assign n8439 = ~n8433 & ~n8438;
  assign n8440 = ~n8432 & ~n8439;
  assign n8441 = po61  & ~n8440;
  assign n8442 = ~po61  & n8440;
  assign n8443 = ~n8050 & ~n8051;
  assign n8444 = po22  & n8443;
  assign n8445 = ~n8056 & ~n8444;
  assign n8446 = n8056 & n8444;
  assign n8447 = ~n8445 & ~n8446;
  assign n8448 = ~n8442 & ~n8447;
  assign n8449 = ~n8441 & ~n8448;
  assign n8450 = po62  & ~n8449;
  assign n8451 = ~po62  & n8449;
  assign n8452 = ~n8059 & ~n8060;
  assign n8453 = po22  & n8452;
  assign n8454 = ~n8065 & ~n8453;
  assign n8455 = n8065 & n8453;
  assign n8456 = ~n8454 & ~n8455;
  assign n8457 = ~n8451 & ~n8456;
  assign n8458 = ~n8450 & ~n8457;
  assign n8459 = n8276 & n8458;
  assign n8460 = ~n8276 & ~n8458;
  assign n8461 = n8078 & po22 ;
  assign n8462 = ~n8077 & ~n8461;
  assign n8463 = n8460 & n8462;
  assign n8464 = ~po63  & ~n8463;
  assign n8465 = ~n7885 & po22 ;
  assign n8466 = n8076 & ~n8465;
  assign n8467 = po63  & ~n8078;
  assign n8468 = ~n8466 & n8467;
  assign n8469 = ~n8459 & ~n8468;
  assign n8470 = ~n8464 & n8469;
  assign po21  = n8271 | ~n8470;
  assign n8472 = ~n8269 & ~n8270;
  assign n8473 = po21  & n8472;
  assign n8474 = ~n8094 & ~n8473;
  assign n8475 = n8094 & n8473;
  assign n8476 = ~n8474 & ~n8475;
  assign n8477 = pi42  & po21 ;
  assign n8478 = ~pi40  & ~pi41 ;
  assign n8479 = ~pi42  & n8478;
  assign n8480 = ~n8477 & ~n8479;
  assign n8481 = po22  & ~n8480;
  assign n8482 = ~po22  & n8480;
  assign n8483 = ~pi42  & po21 ;
  assign n8484 = pi43  & ~n8483;
  assign n8485 = ~pi43  & n8483;
  assign n8486 = ~n8484 & ~n8485;
  assign n8487 = ~n8482 & n8486;
  assign n8488 = ~n8481 & ~n8487;
  assign n8489 = po23  & ~n8488;
  assign n8490 = ~po23  & n8488;
  assign n8491 = po22  & n8470;
  assign n8492 = ~n8485 & ~n8491;
  assign n8493 = pi44  & ~n8492;
  assign n8494 = ~pi44  & n8492;
  assign n8495 = ~n8493 & ~n8494;
  assign n8496 = ~n8490 & ~n8495;
  assign n8497 = ~n8489 & ~n8496;
  assign n8498 = po24  & ~n8497;
  assign n8499 = ~po24  & n8497;
  assign n8500 = ~n8099 & ~n8100;
  assign n8501 = po21  & n8500;
  assign n8502 = n8104 & ~n8501;
  assign n8503 = ~n8104 & n8501;
  assign n8504 = ~n8502 & ~n8503;
  assign n8505 = ~n8499 & ~n8504;
  assign n8506 = ~n8498 & ~n8505;
  assign n8507 = po25  & ~n8506;
  assign n8508 = ~po25  & n8506;
  assign n8509 = ~n8107 & ~n8108;
  assign n8510 = po21  & n8509;
  assign n8511 = ~n8113 & ~n8510;
  assign n8512 = n8113 & n8510;
  assign n8513 = ~n8511 & ~n8512;
  assign n8514 = ~n8508 & ~n8513;
  assign n8515 = ~n8507 & ~n8514;
  assign n8516 = po26  & ~n8515;
  assign n8517 = ~po26  & n8515;
  assign n8518 = ~n8116 & ~n8117;
  assign n8519 = po21  & n8518;
  assign n8520 = n8122 & n8519;
  assign n8521 = ~n8122 & ~n8519;
  assign n8522 = ~n8520 & ~n8521;
  assign n8523 = ~n8517 & ~n8522;
  assign n8524 = ~n8516 & ~n8523;
  assign n8525 = po27  & ~n8524;
  assign n8526 = ~po27  & n8524;
  assign n8527 = ~n8125 & ~n8126;
  assign n8528 = po21  & n8527;
  assign n8529 = ~n8131 & ~n8528;
  assign n8530 = n8131 & n8528;
  assign n8531 = ~n8529 & ~n8530;
  assign n8532 = ~n8526 & ~n8531;
  assign n8533 = ~n8525 & ~n8532;
  assign n8534 = po28  & ~n8533;
  assign n8535 = ~po28  & n8533;
  assign n8536 = ~n8134 & ~n8135;
  assign n8537 = po21  & n8536;
  assign n8538 = ~n8140 & ~n8537;
  assign n8539 = n8140 & n8537;
  assign n8540 = ~n8538 & ~n8539;
  assign n8541 = ~n8535 & ~n8540;
  assign n8542 = ~n8534 & ~n8541;
  assign n8543 = po29  & ~n8542;
  assign n8544 = ~po29  & n8542;
  assign n8545 = ~n8143 & ~n8144;
  assign n8546 = po21  & n8545;
  assign n8547 = ~n8149 & ~n8546;
  assign n8548 = n8149 & n8546;
  assign n8549 = ~n8547 & ~n8548;
  assign n8550 = ~n8544 & ~n8549;
  assign n8551 = ~n8543 & ~n8550;
  assign n8552 = po30  & ~n8551;
  assign n8553 = ~po30  & n8551;
  assign n8554 = ~n8152 & ~n8153;
  assign n8555 = po21  & n8554;
  assign n8556 = ~n8158 & ~n8555;
  assign n8557 = n8158 & n8555;
  assign n8558 = ~n8556 & ~n8557;
  assign n8559 = ~n8553 & ~n8558;
  assign n8560 = ~n8552 & ~n8559;
  assign n8561 = po31  & ~n8560;
  assign n8562 = ~po31  & n8560;
  assign n8563 = ~n8161 & ~n8162;
  assign n8564 = po21  & n8563;
  assign n8565 = ~n8167 & ~n8564;
  assign n8566 = n8167 & n8564;
  assign n8567 = ~n8565 & ~n8566;
  assign n8568 = ~n8562 & ~n8567;
  assign n8569 = ~n8561 & ~n8568;
  assign n8570 = po32  & ~n8569;
  assign n8571 = ~po32  & n8569;
  assign n8572 = ~n8170 & ~n8171;
  assign n8573 = po21  & n8572;
  assign n8574 = ~n8176 & ~n8573;
  assign n8575 = n8176 & n8573;
  assign n8576 = ~n8574 & ~n8575;
  assign n8577 = ~n8571 & ~n8576;
  assign n8578 = ~n8570 & ~n8577;
  assign n8579 = po33  & ~n8578;
  assign n8580 = ~po33  & n8578;
  assign n8581 = ~n8179 & ~n8180;
  assign n8582 = po21  & n8581;
  assign n8583 = ~n8185 & ~n8582;
  assign n8584 = n8185 & n8582;
  assign n8585 = ~n8583 & ~n8584;
  assign n8586 = ~n8580 & ~n8585;
  assign n8587 = ~n8579 & ~n8586;
  assign n8588 = po34  & ~n8587;
  assign n8589 = ~po34  & n8587;
  assign n8590 = ~n8188 & ~n8189;
  assign n8591 = po21  & n8590;
  assign n8592 = ~n8194 & ~n8591;
  assign n8593 = n8194 & n8591;
  assign n8594 = ~n8592 & ~n8593;
  assign n8595 = ~n8589 & ~n8594;
  assign n8596 = ~n8588 & ~n8595;
  assign n8597 = po35  & ~n8596;
  assign n8598 = ~po35  & n8596;
  assign n8599 = ~n8197 & ~n8198;
  assign n8600 = po21  & n8599;
  assign n8601 = ~n8203 & ~n8600;
  assign n8602 = n8203 & n8600;
  assign n8603 = ~n8601 & ~n8602;
  assign n8604 = ~n8598 & ~n8603;
  assign n8605 = ~n8597 & ~n8604;
  assign n8606 = po36  & ~n8605;
  assign n8607 = ~po36  & n8605;
  assign n8608 = ~n8206 & ~n8207;
  assign n8609 = po21  & n8608;
  assign n8610 = ~n8212 & ~n8609;
  assign n8611 = n8212 & n8609;
  assign n8612 = ~n8610 & ~n8611;
  assign n8613 = ~n8607 & ~n8612;
  assign n8614 = ~n8606 & ~n8613;
  assign n8615 = po37  & ~n8614;
  assign n8616 = ~po37  & n8614;
  assign n8617 = ~n8215 & ~n8216;
  assign n8618 = po21  & n8617;
  assign n8619 = ~n8221 & ~n8618;
  assign n8620 = n8221 & n8618;
  assign n8621 = ~n8619 & ~n8620;
  assign n8622 = ~n8616 & ~n8621;
  assign n8623 = ~n8615 & ~n8622;
  assign n8624 = po38  & ~n8623;
  assign n8625 = ~po38  & n8623;
  assign n8626 = ~n8224 & ~n8225;
  assign n8627 = po21  & n8626;
  assign n8628 = ~n8230 & ~n8627;
  assign n8629 = n8230 & n8627;
  assign n8630 = ~n8628 & ~n8629;
  assign n8631 = ~n8625 & ~n8630;
  assign n8632 = ~n8624 & ~n8631;
  assign n8633 = po39  & ~n8632;
  assign n8634 = ~po39  & n8632;
  assign n8635 = ~n8233 & ~n8234;
  assign n8636 = po21  & n8635;
  assign n8637 = ~n8239 & ~n8636;
  assign n8638 = n8239 & n8636;
  assign n8639 = ~n8637 & ~n8638;
  assign n8640 = ~n8634 & ~n8639;
  assign n8641 = ~n8633 & ~n8640;
  assign n8642 = po40  & ~n8641;
  assign n8643 = ~po40  & n8641;
  assign n8644 = ~n8242 & ~n8243;
  assign n8645 = po21  & n8644;
  assign n8646 = ~n8248 & ~n8645;
  assign n8647 = n8248 & n8645;
  assign n8648 = ~n8646 & ~n8647;
  assign n8649 = ~n8643 & ~n8648;
  assign n8650 = ~n8642 & ~n8649;
  assign n8651 = po41  & ~n8650;
  assign n8652 = ~po41  & n8650;
  assign n8653 = ~n8251 & ~n8252;
  assign n8654 = po21  & n8653;
  assign n8655 = ~n8257 & ~n8654;
  assign n8656 = n8257 & n8654;
  assign n8657 = ~n8655 & ~n8656;
  assign n8658 = ~n8652 & ~n8657;
  assign n8659 = ~n8651 & ~n8658;
  assign n8660 = po42  & ~n8659;
  assign n8661 = ~n8260 & ~n8266;
  assign n8662 = po21  & n8661;
  assign n8663 = ~n8265 & ~n8662;
  assign n8664 = n8265 & n8662;
  assign n8665 = ~n8663 & ~n8664;
  assign n8666 = ~po42  & n8659;
  assign n8667 = ~n8665 & ~n8666;
  assign n8668 = ~n8660 & ~n8667;
  assign n8669 = po43  & ~n8668;
  assign n8670 = ~po43  & n8668;
  assign n8671 = n8276 & ~po21 ;
  assign n8672 = ~n8450 & ~n8451;
  assign n8673 = po21  & n8672;
  assign n8674 = ~n8456 & ~n8673;
  assign n8675 = n8456 & n8673;
  assign n8676 = ~n8674 & ~n8675;
  assign n8677 = ~n8476 & ~n8670;
  assign n8678 = ~n8669 & ~n8677;
  assign n8679 = po44  & ~n8678;
  assign n8680 = ~po44  & n8678;
  assign n8681 = ~n8279 & ~n8280;
  assign n8682 = po21  & n8681;
  assign n8683 = ~n8285 & ~n8682;
  assign n8684 = n8285 & n8682;
  assign n8685 = ~n8683 & ~n8684;
  assign n8686 = ~n8680 & ~n8685;
  assign n8687 = ~n8679 & ~n8686;
  assign n8688 = po45  & ~n8687;
  assign n8689 = ~po45  & n8687;
  assign n8690 = ~n8288 & ~n8289;
  assign n8691 = po21  & n8690;
  assign n8692 = ~n8294 & ~n8691;
  assign n8693 = n8294 & n8691;
  assign n8694 = ~n8692 & ~n8693;
  assign n8695 = ~n8689 & ~n8694;
  assign n8696 = ~n8688 & ~n8695;
  assign n8697 = po46  & ~n8696;
  assign n8698 = ~po46  & n8696;
  assign n8699 = ~n8297 & ~n8298;
  assign n8700 = po21  & n8699;
  assign n8701 = ~n8303 & ~n8700;
  assign n8702 = n8303 & n8700;
  assign n8703 = ~n8701 & ~n8702;
  assign n8704 = ~n8698 & ~n8703;
  assign n8705 = ~n8697 & ~n8704;
  assign n8706 = po47  & ~n8705;
  assign n8707 = ~po47  & n8705;
  assign n8708 = ~n8306 & ~n8307;
  assign n8709 = po21  & n8708;
  assign n8710 = ~n8312 & ~n8709;
  assign n8711 = n8312 & n8709;
  assign n8712 = ~n8710 & ~n8711;
  assign n8713 = ~n8707 & ~n8712;
  assign n8714 = ~n8706 & ~n8713;
  assign n8715 = po48  & ~n8714;
  assign n8716 = ~po48  & n8714;
  assign n8717 = ~n8315 & ~n8316;
  assign n8718 = po21  & n8717;
  assign n8719 = ~n8321 & ~n8718;
  assign n8720 = n8321 & n8718;
  assign n8721 = ~n8719 & ~n8720;
  assign n8722 = ~n8716 & ~n8721;
  assign n8723 = ~n8715 & ~n8722;
  assign n8724 = po49  & ~n8723;
  assign n8725 = ~po49  & n8723;
  assign n8726 = ~n8324 & ~n8325;
  assign n8727 = po21  & n8726;
  assign n8728 = ~n8330 & ~n8727;
  assign n8729 = n8330 & n8727;
  assign n8730 = ~n8728 & ~n8729;
  assign n8731 = ~n8725 & ~n8730;
  assign n8732 = ~n8724 & ~n8731;
  assign n8733 = po50  & ~n8732;
  assign n8734 = ~po50  & n8732;
  assign n8735 = ~n8333 & ~n8334;
  assign n8736 = po21  & n8735;
  assign n8737 = ~n8339 & ~n8736;
  assign n8738 = n8339 & n8736;
  assign n8739 = ~n8737 & ~n8738;
  assign n8740 = ~n8734 & ~n8739;
  assign n8741 = ~n8733 & ~n8740;
  assign n8742 = po51  & ~n8741;
  assign n8743 = ~po51  & n8741;
  assign n8744 = ~n8342 & ~n8343;
  assign n8745 = po21  & n8744;
  assign n8746 = ~n8348 & ~n8745;
  assign n8747 = n8348 & n8745;
  assign n8748 = ~n8746 & ~n8747;
  assign n8749 = ~n8743 & ~n8748;
  assign n8750 = ~n8742 & ~n8749;
  assign n8751 = po52  & ~n8750;
  assign n8752 = ~po52  & n8750;
  assign n8753 = ~n8351 & ~n8352;
  assign n8754 = po21  & n8753;
  assign n8755 = ~n8357 & ~n8754;
  assign n8756 = n8357 & n8754;
  assign n8757 = ~n8755 & ~n8756;
  assign n8758 = ~n8752 & ~n8757;
  assign n8759 = ~n8751 & ~n8758;
  assign n8760 = po53  & ~n8759;
  assign n8761 = ~po53  & n8759;
  assign n8762 = ~n8360 & ~n8361;
  assign n8763 = po21  & n8762;
  assign n8764 = ~n8366 & ~n8763;
  assign n8765 = n8366 & n8763;
  assign n8766 = ~n8764 & ~n8765;
  assign n8767 = ~n8761 & ~n8766;
  assign n8768 = ~n8760 & ~n8767;
  assign n8769 = po54  & ~n8768;
  assign n8770 = ~po54  & n8768;
  assign n8771 = ~n8369 & ~n8370;
  assign n8772 = po21  & n8771;
  assign n8773 = ~n8375 & ~n8772;
  assign n8774 = n8375 & n8772;
  assign n8775 = ~n8773 & ~n8774;
  assign n8776 = ~n8770 & ~n8775;
  assign n8777 = ~n8769 & ~n8776;
  assign n8778 = po55  & ~n8777;
  assign n8779 = ~po55  & n8777;
  assign n8780 = ~n8378 & ~n8379;
  assign n8781 = po21  & n8780;
  assign n8782 = ~n8384 & ~n8781;
  assign n8783 = n8384 & n8781;
  assign n8784 = ~n8782 & ~n8783;
  assign n8785 = ~n8779 & ~n8784;
  assign n8786 = ~n8778 & ~n8785;
  assign n8787 = po56  & ~n8786;
  assign n8788 = ~po56  & n8786;
  assign n8789 = ~n8387 & ~n8388;
  assign n8790 = po21  & n8789;
  assign n8791 = ~n8393 & ~n8790;
  assign n8792 = n8393 & n8790;
  assign n8793 = ~n8791 & ~n8792;
  assign n8794 = ~n8788 & ~n8793;
  assign n8795 = ~n8787 & ~n8794;
  assign n8796 = po57  & ~n8795;
  assign n8797 = ~po57  & n8795;
  assign n8798 = ~n8396 & ~n8397;
  assign n8799 = po21  & n8798;
  assign n8800 = ~n8402 & ~n8799;
  assign n8801 = n8402 & n8799;
  assign n8802 = ~n8800 & ~n8801;
  assign n8803 = ~n8797 & ~n8802;
  assign n8804 = ~n8796 & ~n8803;
  assign n8805 = po58  & ~n8804;
  assign n8806 = ~po58  & n8804;
  assign n8807 = ~n8405 & ~n8406;
  assign n8808 = po21  & n8807;
  assign n8809 = ~n8411 & ~n8808;
  assign n8810 = n8411 & n8808;
  assign n8811 = ~n8809 & ~n8810;
  assign n8812 = ~n8806 & ~n8811;
  assign n8813 = ~n8805 & ~n8812;
  assign n8814 = po59  & ~n8813;
  assign n8815 = ~po59  & n8813;
  assign n8816 = ~n8414 & ~n8415;
  assign n8817 = po21  & n8816;
  assign n8818 = ~n8420 & ~n8817;
  assign n8819 = n8420 & n8817;
  assign n8820 = ~n8818 & ~n8819;
  assign n8821 = ~n8815 & ~n8820;
  assign n8822 = ~n8814 & ~n8821;
  assign n8823 = po60  & ~n8822;
  assign n8824 = ~po60  & n8822;
  assign n8825 = ~n8423 & ~n8424;
  assign n8826 = po21  & n8825;
  assign n8827 = ~n8429 & ~n8826;
  assign n8828 = n8429 & n8826;
  assign n8829 = ~n8827 & ~n8828;
  assign n8830 = ~n8824 & ~n8829;
  assign n8831 = ~n8823 & ~n8830;
  assign n8832 = po61  & ~n8831;
  assign n8833 = ~po61  & n8831;
  assign n8834 = ~n8432 & ~n8433;
  assign n8835 = po21  & n8834;
  assign n8836 = ~n8438 & ~n8835;
  assign n8837 = n8438 & n8835;
  assign n8838 = ~n8836 & ~n8837;
  assign n8839 = ~n8833 & ~n8838;
  assign n8840 = ~n8832 & ~n8839;
  assign n8841 = po62  & ~n8840;
  assign n8842 = ~po62  & n8840;
  assign n8843 = ~n8441 & ~n8442;
  assign n8844 = po21  & n8843;
  assign n8845 = ~n8447 & ~n8844;
  assign n8846 = n8447 & n8844;
  assign n8847 = ~n8845 & ~n8846;
  assign n8848 = ~n8842 & ~n8847;
  assign n8849 = ~n8841 & ~n8848;
  assign n8850 = n8676 & n8849;
  assign n8851 = ~n8676 & ~n8849;
  assign n8852 = n8460 & po21 ;
  assign n8853 = ~n8459 & ~n8852;
  assign n8854 = n8851 & n8853;
  assign n8855 = ~po63  & ~n8854;
  assign n8856 = ~n8276 & po21 ;
  assign n8857 = n8458 & ~n8856;
  assign n8858 = po63  & ~n8460;
  assign n8859 = ~n8857 & n8858;
  assign n8860 = ~n8850 & ~n8859;
  assign n8861 = ~n8855 & n8860;
  assign po20  = n8671 | ~n8861;
  assign n8863 = ~n8669 & ~n8670;
  assign n8864 = po20  & n8863;
  assign n8865 = ~n8476 & ~n8864;
  assign n8866 = n8476 & n8864;
  assign n8867 = ~n8865 & ~n8866;
  assign n8868 = pi40  & po20 ;
  assign n8869 = ~pi38  & ~pi39 ;
  assign n8870 = ~pi40  & n8869;
  assign n8871 = ~n8868 & ~n8870;
  assign n8872 = po21  & ~n8871;
  assign n8873 = ~po21  & n8871;
  assign n8874 = ~pi40  & po20 ;
  assign n8875 = pi41  & ~n8874;
  assign n8876 = ~pi41  & n8874;
  assign n8877 = ~n8875 & ~n8876;
  assign n8878 = ~n8873 & n8877;
  assign n8879 = ~n8872 & ~n8878;
  assign n8880 = po22  & ~n8879;
  assign n8881 = ~po22  & n8879;
  assign n8882 = po21  & n8861;
  assign n8883 = ~n8876 & ~n8882;
  assign n8884 = pi42  & ~n8883;
  assign n8885 = ~pi42  & n8883;
  assign n8886 = ~n8884 & ~n8885;
  assign n8887 = ~n8881 & ~n8886;
  assign n8888 = ~n8880 & ~n8887;
  assign n8889 = po23  & ~n8888;
  assign n8890 = ~po23  & n8888;
  assign n8891 = ~n8481 & ~n8482;
  assign n8892 = po20  & n8891;
  assign n8893 = n8486 & ~n8892;
  assign n8894 = ~n8486 & n8892;
  assign n8895 = ~n8893 & ~n8894;
  assign n8896 = ~n8890 & ~n8895;
  assign n8897 = ~n8889 & ~n8896;
  assign n8898 = po24  & ~n8897;
  assign n8899 = ~po24  & n8897;
  assign n8900 = ~n8489 & ~n8490;
  assign n8901 = po20  & n8900;
  assign n8902 = ~n8495 & ~n8901;
  assign n8903 = n8495 & n8901;
  assign n8904 = ~n8902 & ~n8903;
  assign n8905 = ~n8899 & ~n8904;
  assign n8906 = ~n8898 & ~n8905;
  assign n8907 = po25  & ~n8906;
  assign n8908 = ~po25  & n8906;
  assign n8909 = ~n8498 & ~n8499;
  assign n8910 = po20  & n8909;
  assign n8911 = n8504 & n8910;
  assign n8912 = ~n8504 & ~n8910;
  assign n8913 = ~n8911 & ~n8912;
  assign n8914 = ~n8908 & ~n8913;
  assign n8915 = ~n8907 & ~n8914;
  assign n8916 = po26  & ~n8915;
  assign n8917 = ~po26  & n8915;
  assign n8918 = ~n8507 & ~n8508;
  assign n8919 = po20  & n8918;
  assign n8920 = ~n8513 & ~n8919;
  assign n8921 = n8513 & n8919;
  assign n8922 = ~n8920 & ~n8921;
  assign n8923 = ~n8917 & ~n8922;
  assign n8924 = ~n8916 & ~n8923;
  assign n8925 = po27  & ~n8924;
  assign n8926 = ~po27  & n8924;
  assign n8927 = ~n8516 & ~n8517;
  assign n8928 = po20  & n8927;
  assign n8929 = ~n8522 & ~n8928;
  assign n8930 = n8522 & n8928;
  assign n8931 = ~n8929 & ~n8930;
  assign n8932 = ~n8926 & ~n8931;
  assign n8933 = ~n8925 & ~n8932;
  assign n8934 = po28  & ~n8933;
  assign n8935 = ~po28  & n8933;
  assign n8936 = ~n8525 & ~n8526;
  assign n8937 = po20  & n8936;
  assign n8938 = ~n8531 & ~n8937;
  assign n8939 = n8531 & n8937;
  assign n8940 = ~n8938 & ~n8939;
  assign n8941 = ~n8935 & ~n8940;
  assign n8942 = ~n8934 & ~n8941;
  assign n8943 = po29  & ~n8942;
  assign n8944 = ~po29  & n8942;
  assign n8945 = ~n8534 & ~n8535;
  assign n8946 = po20  & n8945;
  assign n8947 = ~n8540 & ~n8946;
  assign n8948 = n8540 & n8946;
  assign n8949 = ~n8947 & ~n8948;
  assign n8950 = ~n8944 & ~n8949;
  assign n8951 = ~n8943 & ~n8950;
  assign n8952 = po30  & ~n8951;
  assign n8953 = ~po30  & n8951;
  assign n8954 = ~n8543 & ~n8544;
  assign n8955 = po20  & n8954;
  assign n8956 = ~n8549 & ~n8955;
  assign n8957 = n8549 & n8955;
  assign n8958 = ~n8956 & ~n8957;
  assign n8959 = ~n8953 & ~n8958;
  assign n8960 = ~n8952 & ~n8959;
  assign n8961 = po31  & ~n8960;
  assign n8962 = ~po31  & n8960;
  assign n8963 = ~n8552 & ~n8553;
  assign n8964 = po20  & n8963;
  assign n8965 = ~n8558 & ~n8964;
  assign n8966 = n8558 & n8964;
  assign n8967 = ~n8965 & ~n8966;
  assign n8968 = ~n8962 & ~n8967;
  assign n8969 = ~n8961 & ~n8968;
  assign n8970 = po32  & ~n8969;
  assign n8971 = ~po32  & n8969;
  assign n8972 = ~n8561 & ~n8562;
  assign n8973 = po20  & n8972;
  assign n8974 = ~n8567 & ~n8973;
  assign n8975 = n8567 & n8973;
  assign n8976 = ~n8974 & ~n8975;
  assign n8977 = ~n8971 & ~n8976;
  assign n8978 = ~n8970 & ~n8977;
  assign n8979 = po33  & ~n8978;
  assign n8980 = ~po33  & n8978;
  assign n8981 = ~n8570 & ~n8571;
  assign n8982 = po20  & n8981;
  assign n8983 = ~n8576 & ~n8982;
  assign n8984 = n8576 & n8982;
  assign n8985 = ~n8983 & ~n8984;
  assign n8986 = ~n8980 & ~n8985;
  assign n8987 = ~n8979 & ~n8986;
  assign n8988 = po34  & ~n8987;
  assign n8989 = ~po34  & n8987;
  assign n8990 = ~n8579 & ~n8580;
  assign n8991 = po20  & n8990;
  assign n8992 = ~n8585 & ~n8991;
  assign n8993 = n8585 & n8991;
  assign n8994 = ~n8992 & ~n8993;
  assign n8995 = ~n8989 & ~n8994;
  assign n8996 = ~n8988 & ~n8995;
  assign n8997 = po35  & ~n8996;
  assign n8998 = ~po35  & n8996;
  assign n8999 = ~n8588 & ~n8589;
  assign n9000 = po20  & n8999;
  assign n9001 = ~n8594 & ~n9000;
  assign n9002 = n8594 & n9000;
  assign n9003 = ~n9001 & ~n9002;
  assign n9004 = ~n8998 & ~n9003;
  assign n9005 = ~n8997 & ~n9004;
  assign n9006 = po36  & ~n9005;
  assign n9007 = ~po36  & n9005;
  assign n9008 = ~n8597 & ~n8598;
  assign n9009 = po20  & n9008;
  assign n9010 = ~n8603 & ~n9009;
  assign n9011 = n8603 & n9009;
  assign n9012 = ~n9010 & ~n9011;
  assign n9013 = ~n9007 & ~n9012;
  assign n9014 = ~n9006 & ~n9013;
  assign n9015 = po37  & ~n9014;
  assign n9016 = ~po37  & n9014;
  assign n9017 = ~n8606 & ~n8607;
  assign n9018 = po20  & n9017;
  assign n9019 = ~n8612 & ~n9018;
  assign n9020 = n8612 & n9018;
  assign n9021 = ~n9019 & ~n9020;
  assign n9022 = ~n9016 & ~n9021;
  assign n9023 = ~n9015 & ~n9022;
  assign n9024 = po38  & ~n9023;
  assign n9025 = ~po38  & n9023;
  assign n9026 = ~n8615 & ~n8616;
  assign n9027 = po20  & n9026;
  assign n9028 = ~n8621 & ~n9027;
  assign n9029 = n8621 & n9027;
  assign n9030 = ~n9028 & ~n9029;
  assign n9031 = ~n9025 & ~n9030;
  assign n9032 = ~n9024 & ~n9031;
  assign n9033 = po39  & ~n9032;
  assign n9034 = ~po39  & n9032;
  assign n9035 = ~n8624 & ~n8625;
  assign n9036 = po20  & n9035;
  assign n9037 = ~n8630 & ~n9036;
  assign n9038 = n8630 & n9036;
  assign n9039 = ~n9037 & ~n9038;
  assign n9040 = ~n9034 & ~n9039;
  assign n9041 = ~n9033 & ~n9040;
  assign n9042 = po40  & ~n9041;
  assign n9043 = ~po40  & n9041;
  assign n9044 = ~n8633 & ~n8634;
  assign n9045 = po20  & n9044;
  assign n9046 = ~n8639 & ~n9045;
  assign n9047 = n8639 & n9045;
  assign n9048 = ~n9046 & ~n9047;
  assign n9049 = ~n9043 & ~n9048;
  assign n9050 = ~n9042 & ~n9049;
  assign n9051 = po41  & ~n9050;
  assign n9052 = ~po41  & n9050;
  assign n9053 = ~n8642 & ~n8643;
  assign n9054 = po20  & n9053;
  assign n9055 = ~n8648 & ~n9054;
  assign n9056 = n8648 & n9054;
  assign n9057 = ~n9055 & ~n9056;
  assign n9058 = ~n9052 & ~n9057;
  assign n9059 = ~n9051 & ~n9058;
  assign n9060 = po42  & ~n9059;
  assign n9061 = ~po42  & n9059;
  assign n9062 = ~n8651 & ~n8652;
  assign n9063 = po20  & n9062;
  assign n9064 = ~n8657 & ~n9063;
  assign n9065 = n8657 & n9063;
  assign n9066 = ~n9064 & ~n9065;
  assign n9067 = ~n9061 & ~n9066;
  assign n9068 = ~n9060 & ~n9067;
  assign n9069 = po43  & ~n9068;
  assign n9070 = ~n8660 & ~n8666;
  assign n9071 = po20  & n9070;
  assign n9072 = ~n8665 & ~n9071;
  assign n9073 = n8665 & n9071;
  assign n9074 = ~n9072 & ~n9073;
  assign n9075 = ~po43  & n9068;
  assign n9076 = ~n9074 & ~n9075;
  assign n9077 = ~n9069 & ~n9076;
  assign n9078 = po44  & ~n9077;
  assign n9079 = ~po44  & n9077;
  assign n9080 = n8676 & ~po20 ;
  assign n9081 = ~n8841 & ~n8842;
  assign n9082 = po20  & n9081;
  assign n9083 = ~n8847 & ~n9082;
  assign n9084 = n8847 & n9082;
  assign n9085 = ~n9083 & ~n9084;
  assign n9086 = ~n8867 & ~n9079;
  assign n9087 = ~n9078 & ~n9086;
  assign n9088 = po45  & ~n9087;
  assign n9089 = ~po45  & n9087;
  assign n9090 = ~n8679 & ~n8680;
  assign n9091 = po20  & n9090;
  assign n9092 = ~n8685 & ~n9091;
  assign n9093 = n8685 & n9091;
  assign n9094 = ~n9092 & ~n9093;
  assign n9095 = ~n9089 & ~n9094;
  assign n9096 = ~n9088 & ~n9095;
  assign n9097 = po46  & ~n9096;
  assign n9098 = ~po46  & n9096;
  assign n9099 = ~n8688 & ~n8689;
  assign n9100 = po20  & n9099;
  assign n9101 = ~n8694 & ~n9100;
  assign n9102 = n8694 & n9100;
  assign n9103 = ~n9101 & ~n9102;
  assign n9104 = ~n9098 & ~n9103;
  assign n9105 = ~n9097 & ~n9104;
  assign n9106 = po47  & ~n9105;
  assign n9107 = ~po47  & n9105;
  assign n9108 = ~n8697 & ~n8698;
  assign n9109 = po20  & n9108;
  assign n9110 = ~n8703 & ~n9109;
  assign n9111 = n8703 & n9109;
  assign n9112 = ~n9110 & ~n9111;
  assign n9113 = ~n9107 & ~n9112;
  assign n9114 = ~n9106 & ~n9113;
  assign n9115 = po48  & ~n9114;
  assign n9116 = ~po48  & n9114;
  assign n9117 = ~n8706 & ~n8707;
  assign n9118 = po20  & n9117;
  assign n9119 = ~n8712 & ~n9118;
  assign n9120 = n8712 & n9118;
  assign n9121 = ~n9119 & ~n9120;
  assign n9122 = ~n9116 & ~n9121;
  assign n9123 = ~n9115 & ~n9122;
  assign n9124 = po49  & ~n9123;
  assign n9125 = ~po49  & n9123;
  assign n9126 = ~n8715 & ~n8716;
  assign n9127 = po20  & n9126;
  assign n9128 = ~n8721 & ~n9127;
  assign n9129 = n8721 & n9127;
  assign n9130 = ~n9128 & ~n9129;
  assign n9131 = ~n9125 & ~n9130;
  assign n9132 = ~n9124 & ~n9131;
  assign n9133 = po50  & ~n9132;
  assign n9134 = ~po50  & n9132;
  assign n9135 = ~n8724 & ~n8725;
  assign n9136 = po20  & n9135;
  assign n9137 = ~n8730 & ~n9136;
  assign n9138 = n8730 & n9136;
  assign n9139 = ~n9137 & ~n9138;
  assign n9140 = ~n9134 & ~n9139;
  assign n9141 = ~n9133 & ~n9140;
  assign n9142 = po51  & ~n9141;
  assign n9143 = ~po51  & n9141;
  assign n9144 = ~n8733 & ~n8734;
  assign n9145 = po20  & n9144;
  assign n9146 = ~n8739 & ~n9145;
  assign n9147 = n8739 & n9145;
  assign n9148 = ~n9146 & ~n9147;
  assign n9149 = ~n9143 & ~n9148;
  assign n9150 = ~n9142 & ~n9149;
  assign n9151 = po52  & ~n9150;
  assign n9152 = ~po52  & n9150;
  assign n9153 = ~n8742 & ~n8743;
  assign n9154 = po20  & n9153;
  assign n9155 = ~n8748 & ~n9154;
  assign n9156 = n8748 & n9154;
  assign n9157 = ~n9155 & ~n9156;
  assign n9158 = ~n9152 & ~n9157;
  assign n9159 = ~n9151 & ~n9158;
  assign n9160 = po53  & ~n9159;
  assign n9161 = ~po53  & n9159;
  assign n9162 = ~n8751 & ~n8752;
  assign n9163 = po20  & n9162;
  assign n9164 = ~n8757 & ~n9163;
  assign n9165 = n8757 & n9163;
  assign n9166 = ~n9164 & ~n9165;
  assign n9167 = ~n9161 & ~n9166;
  assign n9168 = ~n9160 & ~n9167;
  assign n9169 = po54  & ~n9168;
  assign n9170 = ~po54  & n9168;
  assign n9171 = ~n8760 & ~n8761;
  assign n9172 = po20  & n9171;
  assign n9173 = ~n8766 & ~n9172;
  assign n9174 = n8766 & n9172;
  assign n9175 = ~n9173 & ~n9174;
  assign n9176 = ~n9170 & ~n9175;
  assign n9177 = ~n9169 & ~n9176;
  assign n9178 = po55  & ~n9177;
  assign n9179 = ~po55  & n9177;
  assign n9180 = ~n8769 & ~n8770;
  assign n9181 = po20  & n9180;
  assign n9182 = ~n8775 & ~n9181;
  assign n9183 = n8775 & n9181;
  assign n9184 = ~n9182 & ~n9183;
  assign n9185 = ~n9179 & ~n9184;
  assign n9186 = ~n9178 & ~n9185;
  assign n9187 = po56  & ~n9186;
  assign n9188 = ~po56  & n9186;
  assign n9189 = ~n8778 & ~n8779;
  assign n9190 = po20  & n9189;
  assign n9191 = ~n8784 & ~n9190;
  assign n9192 = n8784 & n9190;
  assign n9193 = ~n9191 & ~n9192;
  assign n9194 = ~n9188 & ~n9193;
  assign n9195 = ~n9187 & ~n9194;
  assign n9196 = po57  & ~n9195;
  assign n9197 = ~po57  & n9195;
  assign n9198 = ~n8787 & ~n8788;
  assign n9199 = po20  & n9198;
  assign n9200 = ~n8793 & ~n9199;
  assign n9201 = n8793 & n9199;
  assign n9202 = ~n9200 & ~n9201;
  assign n9203 = ~n9197 & ~n9202;
  assign n9204 = ~n9196 & ~n9203;
  assign n9205 = po58  & ~n9204;
  assign n9206 = ~po58  & n9204;
  assign n9207 = ~n8796 & ~n8797;
  assign n9208 = po20  & n9207;
  assign n9209 = ~n8802 & ~n9208;
  assign n9210 = n8802 & n9208;
  assign n9211 = ~n9209 & ~n9210;
  assign n9212 = ~n9206 & ~n9211;
  assign n9213 = ~n9205 & ~n9212;
  assign n9214 = po59  & ~n9213;
  assign n9215 = ~po59  & n9213;
  assign n9216 = ~n8805 & ~n8806;
  assign n9217 = po20  & n9216;
  assign n9218 = ~n8811 & ~n9217;
  assign n9219 = n8811 & n9217;
  assign n9220 = ~n9218 & ~n9219;
  assign n9221 = ~n9215 & ~n9220;
  assign n9222 = ~n9214 & ~n9221;
  assign n9223 = po60  & ~n9222;
  assign n9224 = ~po60  & n9222;
  assign n9225 = ~n8814 & ~n8815;
  assign n9226 = po20  & n9225;
  assign n9227 = ~n8820 & ~n9226;
  assign n9228 = n8820 & n9226;
  assign n9229 = ~n9227 & ~n9228;
  assign n9230 = ~n9224 & ~n9229;
  assign n9231 = ~n9223 & ~n9230;
  assign n9232 = po61  & ~n9231;
  assign n9233 = ~po61  & n9231;
  assign n9234 = ~n8823 & ~n8824;
  assign n9235 = po20  & n9234;
  assign n9236 = ~n8829 & ~n9235;
  assign n9237 = n8829 & n9235;
  assign n9238 = ~n9236 & ~n9237;
  assign n9239 = ~n9233 & ~n9238;
  assign n9240 = ~n9232 & ~n9239;
  assign n9241 = po62  & ~n9240;
  assign n9242 = ~po62  & n9240;
  assign n9243 = ~n8832 & ~n8833;
  assign n9244 = po20  & n9243;
  assign n9245 = ~n8838 & ~n9244;
  assign n9246 = n8838 & n9244;
  assign n9247 = ~n9245 & ~n9246;
  assign n9248 = ~n9242 & ~n9247;
  assign n9249 = ~n9241 & ~n9248;
  assign n9250 = n9085 & n9249;
  assign n9251 = ~n9085 & ~n9249;
  assign n9252 = n8851 & po20 ;
  assign n9253 = ~n8850 & ~n9252;
  assign n9254 = n9251 & n9253;
  assign n9255 = ~po63  & ~n9254;
  assign n9256 = ~n8676 & po20 ;
  assign n9257 = n8849 & ~n9256;
  assign n9258 = po63  & ~n8851;
  assign n9259 = ~n9257 & n9258;
  assign n9260 = ~n9250 & ~n9259;
  assign n9261 = ~n9255 & n9260;
  assign po19  = n9080 | ~n9261;
  assign n9263 = ~n9078 & ~n9079;
  assign n9264 = po19  & n9263;
  assign n9265 = ~n8867 & ~n9264;
  assign n9266 = n8867 & n9264;
  assign n9267 = ~n9265 & ~n9266;
  assign n9268 = pi38  & po19 ;
  assign n9269 = ~pi36  & ~pi37 ;
  assign n9270 = ~pi38  & n9269;
  assign n9271 = ~n9268 & ~n9270;
  assign n9272 = po20  & ~n9271;
  assign n9273 = ~po20  & n9271;
  assign n9274 = ~pi38  & po19 ;
  assign n9275 = pi39  & ~n9274;
  assign n9276 = ~pi39  & n9274;
  assign n9277 = ~n9275 & ~n9276;
  assign n9278 = ~n9273 & n9277;
  assign n9279 = ~n9272 & ~n9278;
  assign n9280 = po21  & ~n9279;
  assign n9281 = ~po21  & n9279;
  assign n9282 = po20  & n9261;
  assign n9283 = ~n9276 & ~n9282;
  assign n9284 = pi40  & ~n9283;
  assign n9285 = ~pi40  & n9283;
  assign n9286 = ~n9284 & ~n9285;
  assign n9287 = ~n9281 & ~n9286;
  assign n9288 = ~n9280 & ~n9287;
  assign n9289 = po22  & ~n9288;
  assign n9290 = ~po22  & n9288;
  assign n9291 = ~n8872 & ~n8873;
  assign n9292 = po19  & n9291;
  assign n9293 = n8877 & ~n9292;
  assign n9294 = ~n8877 & n9292;
  assign n9295 = ~n9293 & ~n9294;
  assign n9296 = ~n9290 & ~n9295;
  assign n9297 = ~n9289 & ~n9296;
  assign n9298 = po23  & ~n9297;
  assign n9299 = ~po23  & n9297;
  assign n9300 = ~n8880 & ~n8881;
  assign n9301 = po19  & n9300;
  assign n9302 = ~n8886 & ~n9301;
  assign n9303 = n8886 & n9301;
  assign n9304 = ~n9302 & ~n9303;
  assign n9305 = ~n9299 & ~n9304;
  assign n9306 = ~n9298 & ~n9305;
  assign n9307 = po24  & ~n9306;
  assign n9308 = ~po24  & n9306;
  assign n9309 = ~n8889 & ~n8890;
  assign n9310 = po19  & n9309;
  assign n9311 = n8895 & n9310;
  assign n9312 = ~n8895 & ~n9310;
  assign n9313 = ~n9311 & ~n9312;
  assign n9314 = ~n9308 & ~n9313;
  assign n9315 = ~n9307 & ~n9314;
  assign n9316 = po25  & ~n9315;
  assign n9317 = ~po25  & n9315;
  assign n9318 = ~n8898 & ~n8899;
  assign n9319 = po19  & n9318;
  assign n9320 = ~n8904 & ~n9319;
  assign n9321 = n8904 & n9319;
  assign n9322 = ~n9320 & ~n9321;
  assign n9323 = ~n9317 & ~n9322;
  assign n9324 = ~n9316 & ~n9323;
  assign n9325 = po26  & ~n9324;
  assign n9326 = ~po26  & n9324;
  assign n9327 = ~n8907 & ~n8908;
  assign n9328 = po19  & n9327;
  assign n9329 = ~n8913 & ~n9328;
  assign n9330 = n8913 & n9328;
  assign n9331 = ~n9329 & ~n9330;
  assign n9332 = ~n9326 & ~n9331;
  assign n9333 = ~n9325 & ~n9332;
  assign n9334 = po27  & ~n9333;
  assign n9335 = ~po27  & n9333;
  assign n9336 = ~n8916 & ~n8917;
  assign n9337 = po19  & n9336;
  assign n9338 = ~n8922 & ~n9337;
  assign n9339 = n8922 & n9337;
  assign n9340 = ~n9338 & ~n9339;
  assign n9341 = ~n9335 & ~n9340;
  assign n9342 = ~n9334 & ~n9341;
  assign n9343 = po28  & ~n9342;
  assign n9344 = ~po28  & n9342;
  assign n9345 = ~n8925 & ~n8926;
  assign n9346 = po19  & n9345;
  assign n9347 = ~n8931 & ~n9346;
  assign n9348 = n8931 & n9346;
  assign n9349 = ~n9347 & ~n9348;
  assign n9350 = ~n9344 & ~n9349;
  assign n9351 = ~n9343 & ~n9350;
  assign n9352 = po29  & ~n9351;
  assign n9353 = ~po29  & n9351;
  assign n9354 = ~n8934 & ~n8935;
  assign n9355 = po19  & n9354;
  assign n9356 = ~n8940 & ~n9355;
  assign n9357 = n8940 & n9355;
  assign n9358 = ~n9356 & ~n9357;
  assign n9359 = ~n9353 & ~n9358;
  assign n9360 = ~n9352 & ~n9359;
  assign n9361 = po30  & ~n9360;
  assign n9362 = ~po30  & n9360;
  assign n9363 = ~n8943 & ~n8944;
  assign n9364 = po19  & n9363;
  assign n9365 = ~n8949 & ~n9364;
  assign n9366 = n8949 & n9364;
  assign n9367 = ~n9365 & ~n9366;
  assign n9368 = ~n9362 & ~n9367;
  assign n9369 = ~n9361 & ~n9368;
  assign n9370 = po31  & ~n9369;
  assign n9371 = ~po31  & n9369;
  assign n9372 = ~n8952 & ~n8953;
  assign n9373 = po19  & n9372;
  assign n9374 = ~n8958 & ~n9373;
  assign n9375 = n8958 & n9373;
  assign n9376 = ~n9374 & ~n9375;
  assign n9377 = ~n9371 & ~n9376;
  assign n9378 = ~n9370 & ~n9377;
  assign n9379 = po32  & ~n9378;
  assign n9380 = ~po32  & n9378;
  assign n9381 = ~n8961 & ~n8962;
  assign n9382 = po19  & n9381;
  assign n9383 = ~n8967 & ~n9382;
  assign n9384 = n8967 & n9382;
  assign n9385 = ~n9383 & ~n9384;
  assign n9386 = ~n9380 & ~n9385;
  assign n9387 = ~n9379 & ~n9386;
  assign n9388 = po33  & ~n9387;
  assign n9389 = ~po33  & n9387;
  assign n9390 = ~n8970 & ~n8971;
  assign n9391 = po19  & n9390;
  assign n9392 = ~n8976 & ~n9391;
  assign n9393 = n8976 & n9391;
  assign n9394 = ~n9392 & ~n9393;
  assign n9395 = ~n9389 & ~n9394;
  assign n9396 = ~n9388 & ~n9395;
  assign n9397 = po34  & ~n9396;
  assign n9398 = ~po34  & n9396;
  assign n9399 = ~n8979 & ~n8980;
  assign n9400 = po19  & n9399;
  assign n9401 = ~n8985 & ~n9400;
  assign n9402 = n8985 & n9400;
  assign n9403 = ~n9401 & ~n9402;
  assign n9404 = ~n9398 & ~n9403;
  assign n9405 = ~n9397 & ~n9404;
  assign n9406 = po35  & ~n9405;
  assign n9407 = ~po35  & n9405;
  assign n9408 = ~n8988 & ~n8989;
  assign n9409 = po19  & n9408;
  assign n9410 = ~n8994 & ~n9409;
  assign n9411 = n8994 & n9409;
  assign n9412 = ~n9410 & ~n9411;
  assign n9413 = ~n9407 & ~n9412;
  assign n9414 = ~n9406 & ~n9413;
  assign n9415 = po36  & ~n9414;
  assign n9416 = ~po36  & n9414;
  assign n9417 = ~n8997 & ~n8998;
  assign n9418 = po19  & n9417;
  assign n9419 = ~n9003 & ~n9418;
  assign n9420 = n9003 & n9418;
  assign n9421 = ~n9419 & ~n9420;
  assign n9422 = ~n9416 & ~n9421;
  assign n9423 = ~n9415 & ~n9422;
  assign n9424 = po37  & ~n9423;
  assign n9425 = ~po37  & n9423;
  assign n9426 = ~n9006 & ~n9007;
  assign n9427 = po19  & n9426;
  assign n9428 = ~n9012 & ~n9427;
  assign n9429 = n9012 & n9427;
  assign n9430 = ~n9428 & ~n9429;
  assign n9431 = ~n9425 & ~n9430;
  assign n9432 = ~n9424 & ~n9431;
  assign n9433 = po38  & ~n9432;
  assign n9434 = ~po38  & n9432;
  assign n9435 = ~n9015 & ~n9016;
  assign n9436 = po19  & n9435;
  assign n9437 = ~n9021 & ~n9436;
  assign n9438 = n9021 & n9436;
  assign n9439 = ~n9437 & ~n9438;
  assign n9440 = ~n9434 & ~n9439;
  assign n9441 = ~n9433 & ~n9440;
  assign n9442 = po39  & ~n9441;
  assign n9443 = ~po39  & n9441;
  assign n9444 = ~n9024 & ~n9025;
  assign n9445 = po19  & n9444;
  assign n9446 = ~n9030 & ~n9445;
  assign n9447 = n9030 & n9445;
  assign n9448 = ~n9446 & ~n9447;
  assign n9449 = ~n9443 & ~n9448;
  assign n9450 = ~n9442 & ~n9449;
  assign n9451 = po40  & ~n9450;
  assign n9452 = ~po40  & n9450;
  assign n9453 = ~n9033 & ~n9034;
  assign n9454 = po19  & n9453;
  assign n9455 = ~n9039 & ~n9454;
  assign n9456 = n9039 & n9454;
  assign n9457 = ~n9455 & ~n9456;
  assign n9458 = ~n9452 & ~n9457;
  assign n9459 = ~n9451 & ~n9458;
  assign n9460 = po41  & ~n9459;
  assign n9461 = ~po41  & n9459;
  assign n9462 = ~n9042 & ~n9043;
  assign n9463 = po19  & n9462;
  assign n9464 = ~n9048 & ~n9463;
  assign n9465 = n9048 & n9463;
  assign n9466 = ~n9464 & ~n9465;
  assign n9467 = ~n9461 & ~n9466;
  assign n9468 = ~n9460 & ~n9467;
  assign n9469 = po42  & ~n9468;
  assign n9470 = ~po42  & n9468;
  assign n9471 = ~n9051 & ~n9052;
  assign n9472 = po19  & n9471;
  assign n9473 = ~n9057 & ~n9472;
  assign n9474 = n9057 & n9472;
  assign n9475 = ~n9473 & ~n9474;
  assign n9476 = ~n9470 & ~n9475;
  assign n9477 = ~n9469 & ~n9476;
  assign n9478 = po43  & ~n9477;
  assign n9479 = ~po43  & n9477;
  assign n9480 = ~n9060 & ~n9061;
  assign n9481 = po19  & n9480;
  assign n9482 = ~n9066 & ~n9481;
  assign n9483 = n9066 & n9481;
  assign n9484 = ~n9482 & ~n9483;
  assign n9485 = ~n9479 & ~n9484;
  assign n9486 = ~n9478 & ~n9485;
  assign n9487 = po44  & ~n9486;
  assign n9488 = ~n9069 & ~n9075;
  assign n9489 = po19  & n9488;
  assign n9490 = ~n9074 & ~n9489;
  assign n9491 = n9074 & n9489;
  assign n9492 = ~n9490 & ~n9491;
  assign n9493 = ~po44  & n9486;
  assign n9494 = ~n9492 & ~n9493;
  assign n9495 = ~n9487 & ~n9494;
  assign n9496 = po45  & ~n9495;
  assign n9497 = ~po45  & n9495;
  assign n9498 = n9085 & ~po19 ;
  assign n9499 = ~n9241 & ~n9242;
  assign n9500 = po19  & n9499;
  assign n9501 = ~n9247 & ~n9500;
  assign n9502 = n9247 & n9500;
  assign n9503 = ~n9501 & ~n9502;
  assign n9504 = ~n9267 & ~n9497;
  assign n9505 = ~n9496 & ~n9504;
  assign n9506 = po46  & ~n9505;
  assign n9507 = ~po46  & n9505;
  assign n9508 = ~n9088 & ~n9089;
  assign n9509 = po19  & n9508;
  assign n9510 = ~n9094 & ~n9509;
  assign n9511 = n9094 & n9509;
  assign n9512 = ~n9510 & ~n9511;
  assign n9513 = ~n9507 & ~n9512;
  assign n9514 = ~n9506 & ~n9513;
  assign n9515 = po47  & ~n9514;
  assign n9516 = ~po47  & n9514;
  assign n9517 = ~n9097 & ~n9098;
  assign n9518 = po19  & n9517;
  assign n9519 = ~n9103 & ~n9518;
  assign n9520 = n9103 & n9518;
  assign n9521 = ~n9519 & ~n9520;
  assign n9522 = ~n9516 & ~n9521;
  assign n9523 = ~n9515 & ~n9522;
  assign n9524 = po48  & ~n9523;
  assign n9525 = ~po48  & n9523;
  assign n9526 = ~n9106 & ~n9107;
  assign n9527 = po19  & n9526;
  assign n9528 = ~n9112 & ~n9527;
  assign n9529 = n9112 & n9527;
  assign n9530 = ~n9528 & ~n9529;
  assign n9531 = ~n9525 & ~n9530;
  assign n9532 = ~n9524 & ~n9531;
  assign n9533 = po49  & ~n9532;
  assign n9534 = ~po49  & n9532;
  assign n9535 = ~n9115 & ~n9116;
  assign n9536 = po19  & n9535;
  assign n9537 = ~n9121 & ~n9536;
  assign n9538 = n9121 & n9536;
  assign n9539 = ~n9537 & ~n9538;
  assign n9540 = ~n9534 & ~n9539;
  assign n9541 = ~n9533 & ~n9540;
  assign n9542 = po50  & ~n9541;
  assign n9543 = ~po50  & n9541;
  assign n9544 = ~n9124 & ~n9125;
  assign n9545 = po19  & n9544;
  assign n9546 = ~n9130 & ~n9545;
  assign n9547 = n9130 & n9545;
  assign n9548 = ~n9546 & ~n9547;
  assign n9549 = ~n9543 & ~n9548;
  assign n9550 = ~n9542 & ~n9549;
  assign n9551 = po51  & ~n9550;
  assign n9552 = ~po51  & n9550;
  assign n9553 = ~n9133 & ~n9134;
  assign n9554 = po19  & n9553;
  assign n9555 = ~n9139 & ~n9554;
  assign n9556 = n9139 & n9554;
  assign n9557 = ~n9555 & ~n9556;
  assign n9558 = ~n9552 & ~n9557;
  assign n9559 = ~n9551 & ~n9558;
  assign n9560 = po52  & ~n9559;
  assign n9561 = ~po52  & n9559;
  assign n9562 = ~n9142 & ~n9143;
  assign n9563 = po19  & n9562;
  assign n9564 = ~n9148 & ~n9563;
  assign n9565 = n9148 & n9563;
  assign n9566 = ~n9564 & ~n9565;
  assign n9567 = ~n9561 & ~n9566;
  assign n9568 = ~n9560 & ~n9567;
  assign n9569 = po53  & ~n9568;
  assign n9570 = ~po53  & n9568;
  assign n9571 = ~n9151 & ~n9152;
  assign n9572 = po19  & n9571;
  assign n9573 = ~n9157 & ~n9572;
  assign n9574 = n9157 & n9572;
  assign n9575 = ~n9573 & ~n9574;
  assign n9576 = ~n9570 & ~n9575;
  assign n9577 = ~n9569 & ~n9576;
  assign n9578 = po54  & ~n9577;
  assign n9579 = ~po54  & n9577;
  assign n9580 = ~n9160 & ~n9161;
  assign n9581 = po19  & n9580;
  assign n9582 = ~n9166 & ~n9581;
  assign n9583 = n9166 & n9581;
  assign n9584 = ~n9582 & ~n9583;
  assign n9585 = ~n9579 & ~n9584;
  assign n9586 = ~n9578 & ~n9585;
  assign n9587 = po55  & ~n9586;
  assign n9588 = ~po55  & n9586;
  assign n9589 = ~n9169 & ~n9170;
  assign n9590 = po19  & n9589;
  assign n9591 = ~n9175 & ~n9590;
  assign n9592 = n9175 & n9590;
  assign n9593 = ~n9591 & ~n9592;
  assign n9594 = ~n9588 & ~n9593;
  assign n9595 = ~n9587 & ~n9594;
  assign n9596 = po56  & ~n9595;
  assign n9597 = ~po56  & n9595;
  assign n9598 = ~n9178 & ~n9179;
  assign n9599 = po19  & n9598;
  assign n9600 = ~n9184 & ~n9599;
  assign n9601 = n9184 & n9599;
  assign n9602 = ~n9600 & ~n9601;
  assign n9603 = ~n9597 & ~n9602;
  assign n9604 = ~n9596 & ~n9603;
  assign n9605 = po57  & ~n9604;
  assign n9606 = ~po57  & n9604;
  assign n9607 = ~n9187 & ~n9188;
  assign n9608 = po19  & n9607;
  assign n9609 = ~n9193 & ~n9608;
  assign n9610 = n9193 & n9608;
  assign n9611 = ~n9609 & ~n9610;
  assign n9612 = ~n9606 & ~n9611;
  assign n9613 = ~n9605 & ~n9612;
  assign n9614 = po58  & ~n9613;
  assign n9615 = ~po58  & n9613;
  assign n9616 = ~n9196 & ~n9197;
  assign n9617 = po19  & n9616;
  assign n9618 = ~n9202 & ~n9617;
  assign n9619 = n9202 & n9617;
  assign n9620 = ~n9618 & ~n9619;
  assign n9621 = ~n9615 & ~n9620;
  assign n9622 = ~n9614 & ~n9621;
  assign n9623 = po59  & ~n9622;
  assign n9624 = ~po59  & n9622;
  assign n9625 = ~n9205 & ~n9206;
  assign n9626 = po19  & n9625;
  assign n9627 = ~n9211 & ~n9626;
  assign n9628 = n9211 & n9626;
  assign n9629 = ~n9627 & ~n9628;
  assign n9630 = ~n9624 & ~n9629;
  assign n9631 = ~n9623 & ~n9630;
  assign n9632 = po60  & ~n9631;
  assign n9633 = ~po60  & n9631;
  assign n9634 = ~n9214 & ~n9215;
  assign n9635 = po19  & n9634;
  assign n9636 = ~n9220 & ~n9635;
  assign n9637 = n9220 & n9635;
  assign n9638 = ~n9636 & ~n9637;
  assign n9639 = ~n9633 & ~n9638;
  assign n9640 = ~n9632 & ~n9639;
  assign n9641 = po61  & ~n9640;
  assign n9642 = ~po61  & n9640;
  assign n9643 = ~n9223 & ~n9224;
  assign n9644 = po19  & n9643;
  assign n9645 = ~n9229 & ~n9644;
  assign n9646 = n9229 & n9644;
  assign n9647 = ~n9645 & ~n9646;
  assign n9648 = ~n9642 & ~n9647;
  assign n9649 = ~n9641 & ~n9648;
  assign n9650 = po62  & ~n9649;
  assign n9651 = ~po62  & n9649;
  assign n9652 = ~n9232 & ~n9233;
  assign n9653 = po19  & n9652;
  assign n9654 = ~n9238 & ~n9653;
  assign n9655 = n9238 & n9653;
  assign n9656 = ~n9654 & ~n9655;
  assign n9657 = ~n9651 & ~n9656;
  assign n9658 = ~n9650 & ~n9657;
  assign n9659 = n9503 & n9658;
  assign n9660 = ~n9503 & ~n9658;
  assign n9661 = n9251 & po19 ;
  assign n9662 = ~n9250 & ~n9661;
  assign n9663 = n9660 & n9662;
  assign n9664 = ~po63  & ~n9663;
  assign n9665 = ~n9085 & po19 ;
  assign n9666 = n9249 & ~n9665;
  assign n9667 = po63  & ~n9251;
  assign n9668 = ~n9666 & n9667;
  assign n9669 = ~n9659 & ~n9668;
  assign n9670 = ~n9664 & n9669;
  assign po18  = n9498 | ~n9670;
  assign n9672 = ~n9496 & ~n9497;
  assign n9673 = po18  & n9672;
  assign n9674 = ~n9267 & ~n9673;
  assign n9675 = n9267 & n9673;
  assign n9676 = ~n9674 & ~n9675;
  assign n9677 = pi36  & po18 ;
  assign n9678 = ~pi34  & ~pi35 ;
  assign n9679 = ~pi36  & n9678;
  assign n9680 = ~n9677 & ~n9679;
  assign n9681 = po19  & ~n9680;
  assign n9682 = ~po19  & n9680;
  assign n9683 = ~pi36  & po18 ;
  assign n9684 = pi37  & ~n9683;
  assign n9685 = ~pi37  & n9683;
  assign n9686 = ~n9684 & ~n9685;
  assign n9687 = ~n9682 & n9686;
  assign n9688 = ~n9681 & ~n9687;
  assign n9689 = po20  & ~n9688;
  assign n9690 = ~po20  & n9688;
  assign n9691 = po19  & n9670;
  assign n9692 = ~n9685 & ~n9691;
  assign n9693 = pi38  & ~n9692;
  assign n9694 = ~pi38  & n9692;
  assign n9695 = ~n9693 & ~n9694;
  assign n9696 = ~n9690 & ~n9695;
  assign n9697 = ~n9689 & ~n9696;
  assign n9698 = po21  & ~n9697;
  assign n9699 = ~po21  & n9697;
  assign n9700 = ~n9272 & ~n9273;
  assign n9701 = po18  & n9700;
  assign n9702 = n9277 & ~n9701;
  assign n9703 = ~n9277 & n9701;
  assign n9704 = ~n9702 & ~n9703;
  assign n9705 = ~n9699 & ~n9704;
  assign n9706 = ~n9698 & ~n9705;
  assign n9707 = po22  & ~n9706;
  assign n9708 = ~po22  & n9706;
  assign n9709 = ~n9280 & ~n9281;
  assign n9710 = po18  & n9709;
  assign n9711 = ~n9286 & ~n9710;
  assign n9712 = n9286 & n9710;
  assign n9713 = ~n9711 & ~n9712;
  assign n9714 = ~n9708 & ~n9713;
  assign n9715 = ~n9707 & ~n9714;
  assign n9716 = po23  & ~n9715;
  assign n9717 = ~po23  & n9715;
  assign n9718 = ~n9289 & ~n9290;
  assign n9719 = po18  & n9718;
  assign n9720 = n9295 & n9719;
  assign n9721 = ~n9295 & ~n9719;
  assign n9722 = ~n9720 & ~n9721;
  assign n9723 = ~n9717 & ~n9722;
  assign n9724 = ~n9716 & ~n9723;
  assign n9725 = po24  & ~n9724;
  assign n9726 = ~po24  & n9724;
  assign n9727 = ~n9298 & ~n9299;
  assign n9728 = po18  & n9727;
  assign n9729 = ~n9304 & ~n9728;
  assign n9730 = n9304 & n9728;
  assign n9731 = ~n9729 & ~n9730;
  assign n9732 = ~n9726 & ~n9731;
  assign n9733 = ~n9725 & ~n9732;
  assign n9734 = po25  & ~n9733;
  assign n9735 = ~po25  & n9733;
  assign n9736 = ~n9307 & ~n9308;
  assign n9737 = po18  & n9736;
  assign n9738 = ~n9313 & ~n9737;
  assign n9739 = n9313 & n9737;
  assign n9740 = ~n9738 & ~n9739;
  assign n9741 = ~n9735 & ~n9740;
  assign n9742 = ~n9734 & ~n9741;
  assign n9743 = po26  & ~n9742;
  assign n9744 = ~po26  & n9742;
  assign n9745 = ~n9316 & ~n9317;
  assign n9746 = po18  & n9745;
  assign n9747 = ~n9322 & ~n9746;
  assign n9748 = n9322 & n9746;
  assign n9749 = ~n9747 & ~n9748;
  assign n9750 = ~n9744 & ~n9749;
  assign n9751 = ~n9743 & ~n9750;
  assign n9752 = po27  & ~n9751;
  assign n9753 = ~po27  & n9751;
  assign n9754 = ~n9325 & ~n9326;
  assign n9755 = po18  & n9754;
  assign n9756 = ~n9331 & ~n9755;
  assign n9757 = n9331 & n9755;
  assign n9758 = ~n9756 & ~n9757;
  assign n9759 = ~n9753 & ~n9758;
  assign n9760 = ~n9752 & ~n9759;
  assign n9761 = po28  & ~n9760;
  assign n9762 = ~po28  & n9760;
  assign n9763 = ~n9334 & ~n9335;
  assign n9764 = po18  & n9763;
  assign n9765 = ~n9340 & ~n9764;
  assign n9766 = n9340 & n9764;
  assign n9767 = ~n9765 & ~n9766;
  assign n9768 = ~n9762 & ~n9767;
  assign n9769 = ~n9761 & ~n9768;
  assign n9770 = po29  & ~n9769;
  assign n9771 = ~po29  & n9769;
  assign n9772 = ~n9343 & ~n9344;
  assign n9773 = po18  & n9772;
  assign n9774 = ~n9349 & ~n9773;
  assign n9775 = n9349 & n9773;
  assign n9776 = ~n9774 & ~n9775;
  assign n9777 = ~n9771 & ~n9776;
  assign n9778 = ~n9770 & ~n9777;
  assign n9779 = po30  & ~n9778;
  assign n9780 = ~po30  & n9778;
  assign n9781 = ~n9352 & ~n9353;
  assign n9782 = po18  & n9781;
  assign n9783 = ~n9358 & ~n9782;
  assign n9784 = n9358 & n9782;
  assign n9785 = ~n9783 & ~n9784;
  assign n9786 = ~n9780 & ~n9785;
  assign n9787 = ~n9779 & ~n9786;
  assign n9788 = po31  & ~n9787;
  assign n9789 = ~po31  & n9787;
  assign n9790 = ~n9361 & ~n9362;
  assign n9791 = po18  & n9790;
  assign n9792 = ~n9367 & ~n9791;
  assign n9793 = n9367 & n9791;
  assign n9794 = ~n9792 & ~n9793;
  assign n9795 = ~n9789 & ~n9794;
  assign n9796 = ~n9788 & ~n9795;
  assign n9797 = po32  & ~n9796;
  assign n9798 = ~po32  & n9796;
  assign n9799 = ~n9370 & ~n9371;
  assign n9800 = po18  & n9799;
  assign n9801 = ~n9376 & ~n9800;
  assign n9802 = n9376 & n9800;
  assign n9803 = ~n9801 & ~n9802;
  assign n9804 = ~n9798 & ~n9803;
  assign n9805 = ~n9797 & ~n9804;
  assign n9806 = po33  & ~n9805;
  assign n9807 = ~po33  & n9805;
  assign n9808 = ~n9379 & ~n9380;
  assign n9809 = po18  & n9808;
  assign n9810 = ~n9385 & ~n9809;
  assign n9811 = n9385 & n9809;
  assign n9812 = ~n9810 & ~n9811;
  assign n9813 = ~n9807 & ~n9812;
  assign n9814 = ~n9806 & ~n9813;
  assign n9815 = po34  & ~n9814;
  assign n9816 = ~po34  & n9814;
  assign n9817 = ~n9388 & ~n9389;
  assign n9818 = po18  & n9817;
  assign n9819 = ~n9394 & ~n9818;
  assign n9820 = n9394 & n9818;
  assign n9821 = ~n9819 & ~n9820;
  assign n9822 = ~n9816 & ~n9821;
  assign n9823 = ~n9815 & ~n9822;
  assign n9824 = po35  & ~n9823;
  assign n9825 = ~po35  & n9823;
  assign n9826 = ~n9397 & ~n9398;
  assign n9827 = po18  & n9826;
  assign n9828 = ~n9403 & ~n9827;
  assign n9829 = n9403 & n9827;
  assign n9830 = ~n9828 & ~n9829;
  assign n9831 = ~n9825 & ~n9830;
  assign n9832 = ~n9824 & ~n9831;
  assign n9833 = po36  & ~n9832;
  assign n9834 = ~po36  & n9832;
  assign n9835 = ~n9406 & ~n9407;
  assign n9836 = po18  & n9835;
  assign n9837 = ~n9412 & ~n9836;
  assign n9838 = n9412 & n9836;
  assign n9839 = ~n9837 & ~n9838;
  assign n9840 = ~n9834 & ~n9839;
  assign n9841 = ~n9833 & ~n9840;
  assign n9842 = po37  & ~n9841;
  assign n9843 = ~po37  & n9841;
  assign n9844 = ~n9415 & ~n9416;
  assign n9845 = po18  & n9844;
  assign n9846 = ~n9421 & ~n9845;
  assign n9847 = n9421 & n9845;
  assign n9848 = ~n9846 & ~n9847;
  assign n9849 = ~n9843 & ~n9848;
  assign n9850 = ~n9842 & ~n9849;
  assign n9851 = po38  & ~n9850;
  assign n9852 = ~po38  & n9850;
  assign n9853 = ~n9424 & ~n9425;
  assign n9854 = po18  & n9853;
  assign n9855 = ~n9430 & ~n9854;
  assign n9856 = n9430 & n9854;
  assign n9857 = ~n9855 & ~n9856;
  assign n9858 = ~n9852 & ~n9857;
  assign n9859 = ~n9851 & ~n9858;
  assign n9860 = po39  & ~n9859;
  assign n9861 = ~po39  & n9859;
  assign n9862 = ~n9433 & ~n9434;
  assign n9863 = po18  & n9862;
  assign n9864 = ~n9439 & ~n9863;
  assign n9865 = n9439 & n9863;
  assign n9866 = ~n9864 & ~n9865;
  assign n9867 = ~n9861 & ~n9866;
  assign n9868 = ~n9860 & ~n9867;
  assign n9869 = po40  & ~n9868;
  assign n9870 = ~po40  & n9868;
  assign n9871 = ~n9442 & ~n9443;
  assign n9872 = po18  & n9871;
  assign n9873 = ~n9448 & ~n9872;
  assign n9874 = n9448 & n9872;
  assign n9875 = ~n9873 & ~n9874;
  assign n9876 = ~n9870 & ~n9875;
  assign n9877 = ~n9869 & ~n9876;
  assign n9878 = po41  & ~n9877;
  assign n9879 = ~po41  & n9877;
  assign n9880 = ~n9451 & ~n9452;
  assign n9881 = po18  & n9880;
  assign n9882 = ~n9457 & ~n9881;
  assign n9883 = n9457 & n9881;
  assign n9884 = ~n9882 & ~n9883;
  assign n9885 = ~n9879 & ~n9884;
  assign n9886 = ~n9878 & ~n9885;
  assign n9887 = po42  & ~n9886;
  assign n9888 = ~po42  & n9886;
  assign n9889 = ~n9460 & ~n9461;
  assign n9890 = po18  & n9889;
  assign n9891 = ~n9466 & ~n9890;
  assign n9892 = n9466 & n9890;
  assign n9893 = ~n9891 & ~n9892;
  assign n9894 = ~n9888 & ~n9893;
  assign n9895 = ~n9887 & ~n9894;
  assign n9896 = po43  & ~n9895;
  assign n9897 = ~po43  & n9895;
  assign n9898 = ~n9469 & ~n9470;
  assign n9899 = po18  & n9898;
  assign n9900 = ~n9475 & ~n9899;
  assign n9901 = n9475 & n9899;
  assign n9902 = ~n9900 & ~n9901;
  assign n9903 = ~n9897 & ~n9902;
  assign n9904 = ~n9896 & ~n9903;
  assign n9905 = po44  & ~n9904;
  assign n9906 = ~po44  & n9904;
  assign n9907 = ~n9478 & ~n9479;
  assign n9908 = po18  & n9907;
  assign n9909 = ~n9484 & ~n9908;
  assign n9910 = n9484 & n9908;
  assign n9911 = ~n9909 & ~n9910;
  assign n9912 = ~n9906 & ~n9911;
  assign n9913 = ~n9905 & ~n9912;
  assign n9914 = po45  & ~n9913;
  assign n9915 = ~n9487 & ~n9493;
  assign n9916 = po18  & n9915;
  assign n9917 = ~n9492 & ~n9916;
  assign n9918 = n9492 & n9916;
  assign n9919 = ~n9917 & ~n9918;
  assign n9920 = ~po45  & n9913;
  assign n9921 = ~n9919 & ~n9920;
  assign n9922 = ~n9914 & ~n9921;
  assign n9923 = po46  & ~n9922;
  assign n9924 = ~po46  & n9922;
  assign n9925 = n9503 & ~po18 ;
  assign n9926 = ~n9650 & ~n9651;
  assign n9927 = po18  & n9926;
  assign n9928 = ~n9656 & ~n9927;
  assign n9929 = n9656 & n9927;
  assign n9930 = ~n9928 & ~n9929;
  assign n9931 = ~n9676 & ~n9924;
  assign n9932 = ~n9923 & ~n9931;
  assign n9933 = po47  & ~n9932;
  assign n9934 = ~po47  & n9932;
  assign n9935 = ~n9506 & ~n9507;
  assign n9936 = po18  & n9935;
  assign n9937 = ~n9512 & ~n9936;
  assign n9938 = n9512 & n9936;
  assign n9939 = ~n9937 & ~n9938;
  assign n9940 = ~n9934 & ~n9939;
  assign n9941 = ~n9933 & ~n9940;
  assign n9942 = po48  & ~n9941;
  assign n9943 = ~po48  & n9941;
  assign n9944 = ~n9515 & ~n9516;
  assign n9945 = po18  & n9944;
  assign n9946 = ~n9521 & ~n9945;
  assign n9947 = n9521 & n9945;
  assign n9948 = ~n9946 & ~n9947;
  assign n9949 = ~n9943 & ~n9948;
  assign n9950 = ~n9942 & ~n9949;
  assign n9951 = po49  & ~n9950;
  assign n9952 = ~po49  & n9950;
  assign n9953 = ~n9524 & ~n9525;
  assign n9954 = po18  & n9953;
  assign n9955 = ~n9530 & ~n9954;
  assign n9956 = n9530 & n9954;
  assign n9957 = ~n9955 & ~n9956;
  assign n9958 = ~n9952 & ~n9957;
  assign n9959 = ~n9951 & ~n9958;
  assign n9960 = po50  & ~n9959;
  assign n9961 = ~po50  & n9959;
  assign n9962 = ~n9533 & ~n9534;
  assign n9963 = po18  & n9962;
  assign n9964 = ~n9539 & ~n9963;
  assign n9965 = n9539 & n9963;
  assign n9966 = ~n9964 & ~n9965;
  assign n9967 = ~n9961 & ~n9966;
  assign n9968 = ~n9960 & ~n9967;
  assign n9969 = po51  & ~n9968;
  assign n9970 = ~po51  & n9968;
  assign n9971 = ~n9542 & ~n9543;
  assign n9972 = po18  & n9971;
  assign n9973 = ~n9548 & ~n9972;
  assign n9974 = n9548 & n9972;
  assign n9975 = ~n9973 & ~n9974;
  assign n9976 = ~n9970 & ~n9975;
  assign n9977 = ~n9969 & ~n9976;
  assign n9978 = po52  & ~n9977;
  assign n9979 = ~po52  & n9977;
  assign n9980 = ~n9551 & ~n9552;
  assign n9981 = po18  & n9980;
  assign n9982 = ~n9557 & ~n9981;
  assign n9983 = n9557 & n9981;
  assign n9984 = ~n9982 & ~n9983;
  assign n9985 = ~n9979 & ~n9984;
  assign n9986 = ~n9978 & ~n9985;
  assign n9987 = po53  & ~n9986;
  assign n9988 = ~po53  & n9986;
  assign n9989 = ~n9560 & ~n9561;
  assign n9990 = po18  & n9989;
  assign n9991 = ~n9566 & ~n9990;
  assign n9992 = n9566 & n9990;
  assign n9993 = ~n9991 & ~n9992;
  assign n9994 = ~n9988 & ~n9993;
  assign n9995 = ~n9987 & ~n9994;
  assign n9996 = po54  & ~n9995;
  assign n9997 = ~po54  & n9995;
  assign n9998 = ~n9569 & ~n9570;
  assign n9999 = po18  & n9998;
  assign n10000 = ~n9575 & ~n9999;
  assign n10001 = n9575 & n9999;
  assign n10002 = ~n10000 & ~n10001;
  assign n10003 = ~n9997 & ~n10002;
  assign n10004 = ~n9996 & ~n10003;
  assign n10005 = po55  & ~n10004;
  assign n10006 = ~po55  & n10004;
  assign n10007 = ~n9578 & ~n9579;
  assign n10008 = po18  & n10007;
  assign n10009 = ~n9584 & ~n10008;
  assign n10010 = n9584 & n10008;
  assign n10011 = ~n10009 & ~n10010;
  assign n10012 = ~n10006 & ~n10011;
  assign n10013 = ~n10005 & ~n10012;
  assign n10014 = po56  & ~n10013;
  assign n10015 = ~po56  & n10013;
  assign n10016 = ~n9587 & ~n9588;
  assign n10017 = po18  & n10016;
  assign n10018 = ~n9593 & ~n10017;
  assign n10019 = n9593 & n10017;
  assign n10020 = ~n10018 & ~n10019;
  assign n10021 = ~n10015 & ~n10020;
  assign n10022 = ~n10014 & ~n10021;
  assign n10023 = po57  & ~n10022;
  assign n10024 = ~po57  & n10022;
  assign n10025 = ~n9596 & ~n9597;
  assign n10026 = po18  & n10025;
  assign n10027 = ~n9602 & ~n10026;
  assign n10028 = n9602 & n10026;
  assign n10029 = ~n10027 & ~n10028;
  assign n10030 = ~n10024 & ~n10029;
  assign n10031 = ~n10023 & ~n10030;
  assign n10032 = po58  & ~n10031;
  assign n10033 = ~po58  & n10031;
  assign n10034 = ~n9605 & ~n9606;
  assign n10035 = po18  & n10034;
  assign n10036 = ~n9611 & ~n10035;
  assign n10037 = n9611 & n10035;
  assign n10038 = ~n10036 & ~n10037;
  assign n10039 = ~n10033 & ~n10038;
  assign n10040 = ~n10032 & ~n10039;
  assign n10041 = po59  & ~n10040;
  assign n10042 = ~po59  & n10040;
  assign n10043 = ~n9614 & ~n9615;
  assign n10044 = po18  & n10043;
  assign n10045 = ~n9620 & ~n10044;
  assign n10046 = n9620 & n10044;
  assign n10047 = ~n10045 & ~n10046;
  assign n10048 = ~n10042 & ~n10047;
  assign n10049 = ~n10041 & ~n10048;
  assign n10050 = po60  & ~n10049;
  assign n10051 = ~po60  & n10049;
  assign n10052 = ~n9623 & ~n9624;
  assign n10053 = po18  & n10052;
  assign n10054 = ~n9629 & ~n10053;
  assign n10055 = n9629 & n10053;
  assign n10056 = ~n10054 & ~n10055;
  assign n10057 = ~n10051 & ~n10056;
  assign n10058 = ~n10050 & ~n10057;
  assign n10059 = po61  & ~n10058;
  assign n10060 = ~po61  & n10058;
  assign n10061 = ~n9632 & ~n9633;
  assign n10062 = po18  & n10061;
  assign n10063 = ~n9638 & ~n10062;
  assign n10064 = n9638 & n10062;
  assign n10065 = ~n10063 & ~n10064;
  assign n10066 = ~n10060 & ~n10065;
  assign n10067 = ~n10059 & ~n10066;
  assign n10068 = po62  & ~n10067;
  assign n10069 = ~po62  & n10067;
  assign n10070 = ~n9641 & ~n9642;
  assign n10071 = po18  & n10070;
  assign n10072 = ~n9647 & ~n10071;
  assign n10073 = n9647 & n10071;
  assign n10074 = ~n10072 & ~n10073;
  assign n10075 = ~n10069 & ~n10074;
  assign n10076 = ~n10068 & ~n10075;
  assign n10077 = n9930 & n10076;
  assign n10078 = ~n9930 & ~n10076;
  assign n10079 = n9660 & po18 ;
  assign n10080 = ~n9659 & ~n10079;
  assign n10081 = n10078 & n10080;
  assign n10082 = ~po63  & ~n10081;
  assign n10083 = ~n9503 & po18 ;
  assign n10084 = n9658 & ~n10083;
  assign n10085 = po63  & ~n9660;
  assign n10086 = ~n10084 & n10085;
  assign n10087 = ~n10077 & ~n10086;
  assign n10088 = ~n10082 & n10087;
  assign po17  = n9925 | ~n10088;
  assign n10090 = ~n9923 & ~n9924;
  assign n10091 = po17  & n10090;
  assign n10092 = ~n9676 & ~n10091;
  assign n10093 = n9676 & n10091;
  assign n10094 = ~n10092 & ~n10093;
  assign n10095 = pi34  & po17 ;
  assign n10096 = ~pi32  & ~pi33 ;
  assign n10097 = ~pi34  & n10096;
  assign n10098 = ~n10095 & ~n10097;
  assign n10099 = po18  & ~n10098;
  assign n10100 = ~po18  & n10098;
  assign n10101 = ~pi34  & po17 ;
  assign n10102 = pi35  & ~n10101;
  assign n10103 = ~pi35  & n10101;
  assign n10104 = ~n10102 & ~n10103;
  assign n10105 = ~n10100 & n10104;
  assign n10106 = ~n10099 & ~n10105;
  assign n10107 = po19  & ~n10106;
  assign n10108 = ~po19  & n10106;
  assign n10109 = po18  & n10088;
  assign n10110 = ~n10103 & ~n10109;
  assign n10111 = pi36  & ~n10110;
  assign n10112 = ~pi36  & n10110;
  assign n10113 = ~n10111 & ~n10112;
  assign n10114 = ~n10108 & ~n10113;
  assign n10115 = ~n10107 & ~n10114;
  assign n10116 = po20  & ~n10115;
  assign n10117 = ~po20  & n10115;
  assign n10118 = ~n9681 & ~n9682;
  assign n10119 = po17  & n10118;
  assign n10120 = n9686 & ~n10119;
  assign n10121 = ~n9686 & n10119;
  assign n10122 = ~n10120 & ~n10121;
  assign n10123 = ~n10117 & ~n10122;
  assign n10124 = ~n10116 & ~n10123;
  assign n10125 = po21  & ~n10124;
  assign n10126 = ~po21  & n10124;
  assign n10127 = ~n9689 & ~n9690;
  assign n10128 = po17  & n10127;
  assign n10129 = ~n9695 & ~n10128;
  assign n10130 = n9695 & n10128;
  assign n10131 = ~n10129 & ~n10130;
  assign n10132 = ~n10126 & ~n10131;
  assign n10133 = ~n10125 & ~n10132;
  assign n10134 = po22  & ~n10133;
  assign n10135 = ~po22  & n10133;
  assign n10136 = ~n9698 & ~n9699;
  assign n10137 = po17  & n10136;
  assign n10138 = n9704 & n10137;
  assign n10139 = ~n9704 & ~n10137;
  assign n10140 = ~n10138 & ~n10139;
  assign n10141 = ~n10135 & ~n10140;
  assign n10142 = ~n10134 & ~n10141;
  assign n10143 = po23  & ~n10142;
  assign n10144 = ~po23  & n10142;
  assign n10145 = ~n9707 & ~n9708;
  assign n10146 = po17  & n10145;
  assign n10147 = ~n9713 & ~n10146;
  assign n10148 = n9713 & n10146;
  assign n10149 = ~n10147 & ~n10148;
  assign n10150 = ~n10144 & ~n10149;
  assign n10151 = ~n10143 & ~n10150;
  assign n10152 = po24  & ~n10151;
  assign n10153 = ~po24  & n10151;
  assign n10154 = ~n9716 & ~n9717;
  assign n10155 = po17  & n10154;
  assign n10156 = ~n9722 & ~n10155;
  assign n10157 = n9722 & n10155;
  assign n10158 = ~n10156 & ~n10157;
  assign n10159 = ~n10153 & ~n10158;
  assign n10160 = ~n10152 & ~n10159;
  assign n10161 = po25  & ~n10160;
  assign n10162 = ~po25  & n10160;
  assign n10163 = ~n9725 & ~n9726;
  assign n10164 = po17  & n10163;
  assign n10165 = ~n9731 & ~n10164;
  assign n10166 = n9731 & n10164;
  assign n10167 = ~n10165 & ~n10166;
  assign n10168 = ~n10162 & ~n10167;
  assign n10169 = ~n10161 & ~n10168;
  assign n10170 = po26  & ~n10169;
  assign n10171 = ~po26  & n10169;
  assign n10172 = ~n9734 & ~n9735;
  assign n10173 = po17  & n10172;
  assign n10174 = ~n9740 & ~n10173;
  assign n10175 = n9740 & n10173;
  assign n10176 = ~n10174 & ~n10175;
  assign n10177 = ~n10171 & ~n10176;
  assign n10178 = ~n10170 & ~n10177;
  assign n10179 = po27  & ~n10178;
  assign n10180 = ~po27  & n10178;
  assign n10181 = ~n9743 & ~n9744;
  assign n10182 = po17  & n10181;
  assign n10183 = ~n9749 & ~n10182;
  assign n10184 = n9749 & n10182;
  assign n10185 = ~n10183 & ~n10184;
  assign n10186 = ~n10180 & ~n10185;
  assign n10187 = ~n10179 & ~n10186;
  assign n10188 = po28  & ~n10187;
  assign n10189 = ~po28  & n10187;
  assign n10190 = ~n9752 & ~n9753;
  assign n10191 = po17  & n10190;
  assign n10192 = ~n9758 & ~n10191;
  assign n10193 = n9758 & n10191;
  assign n10194 = ~n10192 & ~n10193;
  assign n10195 = ~n10189 & ~n10194;
  assign n10196 = ~n10188 & ~n10195;
  assign n10197 = po29  & ~n10196;
  assign n10198 = ~po29  & n10196;
  assign n10199 = ~n9761 & ~n9762;
  assign n10200 = po17  & n10199;
  assign n10201 = ~n9767 & ~n10200;
  assign n10202 = n9767 & n10200;
  assign n10203 = ~n10201 & ~n10202;
  assign n10204 = ~n10198 & ~n10203;
  assign n10205 = ~n10197 & ~n10204;
  assign n10206 = po30  & ~n10205;
  assign n10207 = ~po30  & n10205;
  assign n10208 = ~n9770 & ~n9771;
  assign n10209 = po17  & n10208;
  assign n10210 = ~n9776 & ~n10209;
  assign n10211 = n9776 & n10209;
  assign n10212 = ~n10210 & ~n10211;
  assign n10213 = ~n10207 & ~n10212;
  assign n10214 = ~n10206 & ~n10213;
  assign n10215 = po31  & ~n10214;
  assign n10216 = ~po31  & n10214;
  assign n10217 = ~n9779 & ~n9780;
  assign n10218 = po17  & n10217;
  assign n10219 = ~n9785 & ~n10218;
  assign n10220 = n9785 & n10218;
  assign n10221 = ~n10219 & ~n10220;
  assign n10222 = ~n10216 & ~n10221;
  assign n10223 = ~n10215 & ~n10222;
  assign n10224 = po32  & ~n10223;
  assign n10225 = ~po32  & n10223;
  assign n10226 = ~n9788 & ~n9789;
  assign n10227 = po17  & n10226;
  assign n10228 = ~n9794 & ~n10227;
  assign n10229 = n9794 & n10227;
  assign n10230 = ~n10228 & ~n10229;
  assign n10231 = ~n10225 & ~n10230;
  assign n10232 = ~n10224 & ~n10231;
  assign n10233 = po33  & ~n10232;
  assign n10234 = ~po33  & n10232;
  assign n10235 = ~n9797 & ~n9798;
  assign n10236 = po17  & n10235;
  assign n10237 = ~n9803 & ~n10236;
  assign n10238 = n9803 & n10236;
  assign n10239 = ~n10237 & ~n10238;
  assign n10240 = ~n10234 & ~n10239;
  assign n10241 = ~n10233 & ~n10240;
  assign n10242 = po34  & ~n10241;
  assign n10243 = ~po34  & n10241;
  assign n10244 = ~n9806 & ~n9807;
  assign n10245 = po17  & n10244;
  assign n10246 = ~n9812 & ~n10245;
  assign n10247 = n9812 & n10245;
  assign n10248 = ~n10246 & ~n10247;
  assign n10249 = ~n10243 & ~n10248;
  assign n10250 = ~n10242 & ~n10249;
  assign n10251 = po35  & ~n10250;
  assign n10252 = ~po35  & n10250;
  assign n10253 = ~n9815 & ~n9816;
  assign n10254 = po17  & n10253;
  assign n10255 = ~n9821 & ~n10254;
  assign n10256 = n9821 & n10254;
  assign n10257 = ~n10255 & ~n10256;
  assign n10258 = ~n10252 & ~n10257;
  assign n10259 = ~n10251 & ~n10258;
  assign n10260 = po36  & ~n10259;
  assign n10261 = ~po36  & n10259;
  assign n10262 = ~n9824 & ~n9825;
  assign n10263 = po17  & n10262;
  assign n10264 = ~n9830 & ~n10263;
  assign n10265 = n9830 & n10263;
  assign n10266 = ~n10264 & ~n10265;
  assign n10267 = ~n10261 & ~n10266;
  assign n10268 = ~n10260 & ~n10267;
  assign n10269 = po37  & ~n10268;
  assign n10270 = ~po37  & n10268;
  assign n10271 = ~n9833 & ~n9834;
  assign n10272 = po17  & n10271;
  assign n10273 = ~n9839 & ~n10272;
  assign n10274 = n9839 & n10272;
  assign n10275 = ~n10273 & ~n10274;
  assign n10276 = ~n10270 & ~n10275;
  assign n10277 = ~n10269 & ~n10276;
  assign n10278 = po38  & ~n10277;
  assign n10279 = ~po38  & n10277;
  assign n10280 = ~n9842 & ~n9843;
  assign n10281 = po17  & n10280;
  assign n10282 = ~n9848 & ~n10281;
  assign n10283 = n9848 & n10281;
  assign n10284 = ~n10282 & ~n10283;
  assign n10285 = ~n10279 & ~n10284;
  assign n10286 = ~n10278 & ~n10285;
  assign n10287 = po39  & ~n10286;
  assign n10288 = ~po39  & n10286;
  assign n10289 = ~n9851 & ~n9852;
  assign n10290 = po17  & n10289;
  assign n10291 = ~n9857 & ~n10290;
  assign n10292 = n9857 & n10290;
  assign n10293 = ~n10291 & ~n10292;
  assign n10294 = ~n10288 & ~n10293;
  assign n10295 = ~n10287 & ~n10294;
  assign n10296 = po40  & ~n10295;
  assign n10297 = ~po40  & n10295;
  assign n10298 = ~n9860 & ~n9861;
  assign n10299 = po17  & n10298;
  assign n10300 = ~n9866 & ~n10299;
  assign n10301 = n9866 & n10299;
  assign n10302 = ~n10300 & ~n10301;
  assign n10303 = ~n10297 & ~n10302;
  assign n10304 = ~n10296 & ~n10303;
  assign n10305 = po41  & ~n10304;
  assign n10306 = ~po41  & n10304;
  assign n10307 = ~n9869 & ~n9870;
  assign n10308 = po17  & n10307;
  assign n10309 = ~n9875 & ~n10308;
  assign n10310 = n9875 & n10308;
  assign n10311 = ~n10309 & ~n10310;
  assign n10312 = ~n10306 & ~n10311;
  assign n10313 = ~n10305 & ~n10312;
  assign n10314 = po42  & ~n10313;
  assign n10315 = ~po42  & n10313;
  assign n10316 = ~n9878 & ~n9879;
  assign n10317 = po17  & n10316;
  assign n10318 = ~n9884 & ~n10317;
  assign n10319 = n9884 & n10317;
  assign n10320 = ~n10318 & ~n10319;
  assign n10321 = ~n10315 & ~n10320;
  assign n10322 = ~n10314 & ~n10321;
  assign n10323 = po43  & ~n10322;
  assign n10324 = ~po43  & n10322;
  assign n10325 = ~n9887 & ~n9888;
  assign n10326 = po17  & n10325;
  assign n10327 = ~n9893 & ~n10326;
  assign n10328 = n9893 & n10326;
  assign n10329 = ~n10327 & ~n10328;
  assign n10330 = ~n10324 & ~n10329;
  assign n10331 = ~n10323 & ~n10330;
  assign n10332 = po44  & ~n10331;
  assign n10333 = ~po44  & n10331;
  assign n10334 = ~n9896 & ~n9897;
  assign n10335 = po17  & n10334;
  assign n10336 = ~n9902 & ~n10335;
  assign n10337 = n9902 & n10335;
  assign n10338 = ~n10336 & ~n10337;
  assign n10339 = ~n10333 & ~n10338;
  assign n10340 = ~n10332 & ~n10339;
  assign n10341 = po45  & ~n10340;
  assign n10342 = ~po45  & n10340;
  assign n10343 = ~n9905 & ~n9906;
  assign n10344 = po17  & n10343;
  assign n10345 = ~n9911 & ~n10344;
  assign n10346 = n9911 & n10344;
  assign n10347 = ~n10345 & ~n10346;
  assign n10348 = ~n10342 & ~n10347;
  assign n10349 = ~n10341 & ~n10348;
  assign n10350 = po46  & ~n10349;
  assign n10351 = ~n9914 & ~n9920;
  assign n10352 = po17  & n10351;
  assign n10353 = ~n9919 & ~n10352;
  assign n10354 = n9919 & n10352;
  assign n10355 = ~n10353 & ~n10354;
  assign n10356 = ~po46  & n10349;
  assign n10357 = ~n10355 & ~n10356;
  assign n10358 = ~n10350 & ~n10357;
  assign n10359 = po47  & ~n10358;
  assign n10360 = ~po47  & n10358;
  assign n10361 = n9930 & ~po17 ;
  assign n10362 = ~n10068 & ~n10069;
  assign n10363 = po17  & n10362;
  assign n10364 = ~n10074 & ~n10363;
  assign n10365 = n10074 & n10363;
  assign n10366 = ~n10364 & ~n10365;
  assign n10367 = ~n10094 & ~n10360;
  assign n10368 = ~n10359 & ~n10367;
  assign n10369 = po48  & ~n10368;
  assign n10370 = ~po48  & n10368;
  assign n10371 = ~n9933 & ~n9934;
  assign n10372 = po17  & n10371;
  assign n10373 = ~n9939 & ~n10372;
  assign n10374 = n9939 & n10372;
  assign n10375 = ~n10373 & ~n10374;
  assign n10376 = ~n10370 & ~n10375;
  assign n10377 = ~n10369 & ~n10376;
  assign n10378 = po49  & ~n10377;
  assign n10379 = ~po49  & n10377;
  assign n10380 = ~n9942 & ~n9943;
  assign n10381 = po17  & n10380;
  assign n10382 = ~n9948 & ~n10381;
  assign n10383 = n9948 & n10381;
  assign n10384 = ~n10382 & ~n10383;
  assign n10385 = ~n10379 & ~n10384;
  assign n10386 = ~n10378 & ~n10385;
  assign n10387 = po50  & ~n10386;
  assign n10388 = ~po50  & n10386;
  assign n10389 = ~n9951 & ~n9952;
  assign n10390 = po17  & n10389;
  assign n10391 = ~n9957 & ~n10390;
  assign n10392 = n9957 & n10390;
  assign n10393 = ~n10391 & ~n10392;
  assign n10394 = ~n10388 & ~n10393;
  assign n10395 = ~n10387 & ~n10394;
  assign n10396 = po51  & ~n10395;
  assign n10397 = ~po51  & n10395;
  assign n10398 = ~n9960 & ~n9961;
  assign n10399 = po17  & n10398;
  assign n10400 = ~n9966 & ~n10399;
  assign n10401 = n9966 & n10399;
  assign n10402 = ~n10400 & ~n10401;
  assign n10403 = ~n10397 & ~n10402;
  assign n10404 = ~n10396 & ~n10403;
  assign n10405 = po52  & ~n10404;
  assign n10406 = ~po52  & n10404;
  assign n10407 = ~n9969 & ~n9970;
  assign n10408 = po17  & n10407;
  assign n10409 = ~n9975 & ~n10408;
  assign n10410 = n9975 & n10408;
  assign n10411 = ~n10409 & ~n10410;
  assign n10412 = ~n10406 & ~n10411;
  assign n10413 = ~n10405 & ~n10412;
  assign n10414 = po53  & ~n10413;
  assign n10415 = ~po53  & n10413;
  assign n10416 = ~n9978 & ~n9979;
  assign n10417 = po17  & n10416;
  assign n10418 = ~n9984 & ~n10417;
  assign n10419 = n9984 & n10417;
  assign n10420 = ~n10418 & ~n10419;
  assign n10421 = ~n10415 & ~n10420;
  assign n10422 = ~n10414 & ~n10421;
  assign n10423 = po54  & ~n10422;
  assign n10424 = ~po54  & n10422;
  assign n10425 = ~n9987 & ~n9988;
  assign n10426 = po17  & n10425;
  assign n10427 = ~n9993 & ~n10426;
  assign n10428 = n9993 & n10426;
  assign n10429 = ~n10427 & ~n10428;
  assign n10430 = ~n10424 & ~n10429;
  assign n10431 = ~n10423 & ~n10430;
  assign n10432 = po55  & ~n10431;
  assign n10433 = ~po55  & n10431;
  assign n10434 = ~n9996 & ~n9997;
  assign n10435 = po17  & n10434;
  assign n10436 = ~n10002 & ~n10435;
  assign n10437 = n10002 & n10435;
  assign n10438 = ~n10436 & ~n10437;
  assign n10439 = ~n10433 & ~n10438;
  assign n10440 = ~n10432 & ~n10439;
  assign n10441 = po56  & ~n10440;
  assign n10442 = ~po56  & n10440;
  assign n10443 = ~n10005 & ~n10006;
  assign n10444 = po17  & n10443;
  assign n10445 = ~n10011 & ~n10444;
  assign n10446 = n10011 & n10444;
  assign n10447 = ~n10445 & ~n10446;
  assign n10448 = ~n10442 & ~n10447;
  assign n10449 = ~n10441 & ~n10448;
  assign n10450 = po57  & ~n10449;
  assign n10451 = ~po57  & n10449;
  assign n10452 = ~n10014 & ~n10015;
  assign n10453 = po17  & n10452;
  assign n10454 = ~n10020 & ~n10453;
  assign n10455 = n10020 & n10453;
  assign n10456 = ~n10454 & ~n10455;
  assign n10457 = ~n10451 & ~n10456;
  assign n10458 = ~n10450 & ~n10457;
  assign n10459 = po58  & ~n10458;
  assign n10460 = ~po58  & n10458;
  assign n10461 = ~n10023 & ~n10024;
  assign n10462 = po17  & n10461;
  assign n10463 = ~n10029 & ~n10462;
  assign n10464 = n10029 & n10462;
  assign n10465 = ~n10463 & ~n10464;
  assign n10466 = ~n10460 & ~n10465;
  assign n10467 = ~n10459 & ~n10466;
  assign n10468 = po59  & ~n10467;
  assign n10469 = ~po59  & n10467;
  assign n10470 = ~n10032 & ~n10033;
  assign n10471 = po17  & n10470;
  assign n10472 = ~n10038 & ~n10471;
  assign n10473 = n10038 & n10471;
  assign n10474 = ~n10472 & ~n10473;
  assign n10475 = ~n10469 & ~n10474;
  assign n10476 = ~n10468 & ~n10475;
  assign n10477 = po60  & ~n10476;
  assign n10478 = ~po60  & n10476;
  assign n10479 = ~n10041 & ~n10042;
  assign n10480 = po17  & n10479;
  assign n10481 = ~n10047 & ~n10480;
  assign n10482 = n10047 & n10480;
  assign n10483 = ~n10481 & ~n10482;
  assign n10484 = ~n10478 & ~n10483;
  assign n10485 = ~n10477 & ~n10484;
  assign n10486 = po61  & ~n10485;
  assign n10487 = ~po61  & n10485;
  assign n10488 = ~n10050 & ~n10051;
  assign n10489 = po17  & n10488;
  assign n10490 = ~n10056 & ~n10489;
  assign n10491 = n10056 & n10489;
  assign n10492 = ~n10490 & ~n10491;
  assign n10493 = ~n10487 & ~n10492;
  assign n10494 = ~n10486 & ~n10493;
  assign n10495 = po62  & ~n10494;
  assign n10496 = ~po62  & n10494;
  assign n10497 = ~n10059 & ~n10060;
  assign n10498 = po17  & n10497;
  assign n10499 = ~n10065 & ~n10498;
  assign n10500 = n10065 & n10498;
  assign n10501 = ~n10499 & ~n10500;
  assign n10502 = ~n10496 & ~n10501;
  assign n10503 = ~n10495 & ~n10502;
  assign n10504 = n10366 & n10503;
  assign n10505 = ~n10366 & ~n10503;
  assign n10506 = n10078 & po17 ;
  assign n10507 = ~n10077 & ~n10506;
  assign n10508 = n10505 & n10507;
  assign n10509 = ~po63  & ~n10508;
  assign n10510 = ~n9930 & po17 ;
  assign n10511 = n10076 & ~n10510;
  assign n10512 = po63  & ~n10078;
  assign n10513 = ~n10511 & n10512;
  assign n10514 = ~n10504 & ~n10513;
  assign n10515 = ~n10509 & n10514;
  assign po16  = n10361 | ~n10515;
  assign n10517 = ~n10359 & ~n10360;
  assign n10518 = po16  & n10517;
  assign n10519 = ~n10094 & ~n10518;
  assign n10520 = n10094 & n10518;
  assign n10521 = ~n10519 & ~n10520;
  assign n10522 = pi32  & po16 ;
  assign n10523 = ~pi30  & ~pi31 ;
  assign n10524 = ~pi32  & n10523;
  assign n10525 = ~n10522 & ~n10524;
  assign n10526 = po17  & ~n10525;
  assign n10527 = ~po17  & n10525;
  assign n10528 = ~pi32  & po16 ;
  assign n10529 = pi33  & ~n10528;
  assign n10530 = ~pi33  & n10528;
  assign n10531 = ~n10529 & ~n10530;
  assign n10532 = ~n10527 & n10531;
  assign n10533 = ~n10526 & ~n10532;
  assign n10534 = po18  & ~n10533;
  assign n10535 = ~po18  & n10533;
  assign n10536 = po17  & n10515;
  assign n10537 = ~n10530 & ~n10536;
  assign n10538 = pi34  & ~n10537;
  assign n10539 = ~pi34  & n10537;
  assign n10540 = ~n10538 & ~n10539;
  assign n10541 = ~n10535 & ~n10540;
  assign n10542 = ~n10534 & ~n10541;
  assign n10543 = po19  & ~n10542;
  assign n10544 = ~po19  & n10542;
  assign n10545 = ~n10099 & ~n10100;
  assign n10546 = po16  & n10545;
  assign n10547 = n10104 & ~n10546;
  assign n10548 = ~n10104 & n10546;
  assign n10549 = ~n10547 & ~n10548;
  assign n10550 = ~n10544 & ~n10549;
  assign n10551 = ~n10543 & ~n10550;
  assign n10552 = po20  & ~n10551;
  assign n10553 = ~po20  & n10551;
  assign n10554 = ~n10107 & ~n10108;
  assign n10555 = po16  & n10554;
  assign n10556 = ~n10113 & ~n10555;
  assign n10557 = n10113 & n10555;
  assign n10558 = ~n10556 & ~n10557;
  assign n10559 = ~n10553 & ~n10558;
  assign n10560 = ~n10552 & ~n10559;
  assign n10561 = po21  & ~n10560;
  assign n10562 = ~po21  & n10560;
  assign n10563 = ~n10116 & ~n10117;
  assign n10564 = po16  & n10563;
  assign n10565 = n10122 & n10564;
  assign n10566 = ~n10122 & ~n10564;
  assign n10567 = ~n10565 & ~n10566;
  assign n10568 = ~n10562 & ~n10567;
  assign n10569 = ~n10561 & ~n10568;
  assign n10570 = po22  & ~n10569;
  assign n10571 = ~po22  & n10569;
  assign n10572 = ~n10125 & ~n10126;
  assign n10573 = po16  & n10572;
  assign n10574 = ~n10131 & ~n10573;
  assign n10575 = n10131 & n10573;
  assign n10576 = ~n10574 & ~n10575;
  assign n10577 = ~n10571 & ~n10576;
  assign n10578 = ~n10570 & ~n10577;
  assign n10579 = po23  & ~n10578;
  assign n10580 = ~po23  & n10578;
  assign n10581 = ~n10134 & ~n10135;
  assign n10582 = po16  & n10581;
  assign n10583 = ~n10140 & ~n10582;
  assign n10584 = n10140 & n10582;
  assign n10585 = ~n10583 & ~n10584;
  assign n10586 = ~n10580 & ~n10585;
  assign n10587 = ~n10579 & ~n10586;
  assign n10588 = po24  & ~n10587;
  assign n10589 = ~po24  & n10587;
  assign n10590 = ~n10143 & ~n10144;
  assign n10591 = po16  & n10590;
  assign n10592 = ~n10149 & ~n10591;
  assign n10593 = n10149 & n10591;
  assign n10594 = ~n10592 & ~n10593;
  assign n10595 = ~n10589 & ~n10594;
  assign n10596 = ~n10588 & ~n10595;
  assign n10597 = po25  & ~n10596;
  assign n10598 = ~po25  & n10596;
  assign n10599 = ~n10152 & ~n10153;
  assign n10600 = po16  & n10599;
  assign n10601 = ~n10158 & ~n10600;
  assign n10602 = n10158 & n10600;
  assign n10603 = ~n10601 & ~n10602;
  assign n10604 = ~n10598 & ~n10603;
  assign n10605 = ~n10597 & ~n10604;
  assign n10606 = po26  & ~n10605;
  assign n10607 = ~po26  & n10605;
  assign n10608 = ~n10161 & ~n10162;
  assign n10609 = po16  & n10608;
  assign n10610 = ~n10167 & ~n10609;
  assign n10611 = n10167 & n10609;
  assign n10612 = ~n10610 & ~n10611;
  assign n10613 = ~n10607 & ~n10612;
  assign n10614 = ~n10606 & ~n10613;
  assign n10615 = po27  & ~n10614;
  assign n10616 = ~po27  & n10614;
  assign n10617 = ~n10170 & ~n10171;
  assign n10618 = po16  & n10617;
  assign n10619 = ~n10176 & ~n10618;
  assign n10620 = n10176 & n10618;
  assign n10621 = ~n10619 & ~n10620;
  assign n10622 = ~n10616 & ~n10621;
  assign n10623 = ~n10615 & ~n10622;
  assign n10624 = po28  & ~n10623;
  assign n10625 = ~po28  & n10623;
  assign n10626 = ~n10179 & ~n10180;
  assign n10627 = po16  & n10626;
  assign n10628 = ~n10185 & ~n10627;
  assign n10629 = n10185 & n10627;
  assign n10630 = ~n10628 & ~n10629;
  assign n10631 = ~n10625 & ~n10630;
  assign n10632 = ~n10624 & ~n10631;
  assign n10633 = po29  & ~n10632;
  assign n10634 = ~po29  & n10632;
  assign n10635 = ~n10188 & ~n10189;
  assign n10636 = po16  & n10635;
  assign n10637 = ~n10194 & ~n10636;
  assign n10638 = n10194 & n10636;
  assign n10639 = ~n10637 & ~n10638;
  assign n10640 = ~n10634 & ~n10639;
  assign n10641 = ~n10633 & ~n10640;
  assign n10642 = po30  & ~n10641;
  assign n10643 = ~po30  & n10641;
  assign n10644 = ~n10197 & ~n10198;
  assign n10645 = po16  & n10644;
  assign n10646 = ~n10203 & ~n10645;
  assign n10647 = n10203 & n10645;
  assign n10648 = ~n10646 & ~n10647;
  assign n10649 = ~n10643 & ~n10648;
  assign n10650 = ~n10642 & ~n10649;
  assign n10651 = po31  & ~n10650;
  assign n10652 = ~po31  & n10650;
  assign n10653 = ~n10206 & ~n10207;
  assign n10654 = po16  & n10653;
  assign n10655 = ~n10212 & ~n10654;
  assign n10656 = n10212 & n10654;
  assign n10657 = ~n10655 & ~n10656;
  assign n10658 = ~n10652 & ~n10657;
  assign n10659 = ~n10651 & ~n10658;
  assign n10660 = po32  & ~n10659;
  assign n10661 = ~po32  & n10659;
  assign n10662 = ~n10215 & ~n10216;
  assign n10663 = po16  & n10662;
  assign n10664 = ~n10221 & ~n10663;
  assign n10665 = n10221 & n10663;
  assign n10666 = ~n10664 & ~n10665;
  assign n10667 = ~n10661 & ~n10666;
  assign n10668 = ~n10660 & ~n10667;
  assign n10669 = po33  & ~n10668;
  assign n10670 = ~po33  & n10668;
  assign n10671 = ~n10224 & ~n10225;
  assign n10672 = po16  & n10671;
  assign n10673 = ~n10230 & ~n10672;
  assign n10674 = n10230 & n10672;
  assign n10675 = ~n10673 & ~n10674;
  assign n10676 = ~n10670 & ~n10675;
  assign n10677 = ~n10669 & ~n10676;
  assign n10678 = po34  & ~n10677;
  assign n10679 = ~po34  & n10677;
  assign n10680 = ~n10233 & ~n10234;
  assign n10681 = po16  & n10680;
  assign n10682 = ~n10239 & ~n10681;
  assign n10683 = n10239 & n10681;
  assign n10684 = ~n10682 & ~n10683;
  assign n10685 = ~n10679 & ~n10684;
  assign n10686 = ~n10678 & ~n10685;
  assign n10687 = po35  & ~n10686;
  assign n10688 = ~po35  & n10686;
  assign n10689 = ~n10242 & ~n10243;
  assign n10690 = po16  & n10689;
  assign n10691 = ~n10248 & ~n10690;
  assign n10692 = n10248 & n10690;
  assign n10693 = ~n10691 & ~n10692;
  assign n10694 = ~n10688 & ~n10693;
  assign n10695 = ~n10687 & ~n10694;
  assign n10696 = po36  & ~n10695;
  assign n10697 = ~po36  & n10695;
  assign n10698 = ~n10251 & ~n10252;
  assign n10699 = po16  & n10698;
  assign n10700 = ~n10257 & ~n10699;
  assign n10701 = n10257 & n10699;
  assign n10702 = ~n10700 & ~n10701;
  assign n10703 = ~n10697 & ~n10702;
  assign n10704 = ~n10696 & ~n10703;
  assign n10705 = po37  & ~n10704;
  assign n10706 = ~po37  & n10704;
  assign n10707 = ~n10260 & ~n10261;
  assign n10708 = po16  & n10707;
  assign n10709 = ~n10266 & ~n10708;
  assign n10710 = n10266 & n10708;
  assign n10711 = ~n10709 & ~n10710;
  assign n10712 = ~n10706 & ~n10711;
  assign n10713 = ~n10705 & ~n10712;
  assign n10714 = po38  & ~n10713;
  assign n10715 = ~po38  & n10713;
  assign n10716 = ~n10269 & ~n10270;
  assign n10717 = po16  & n10716;
  assign n10718 = ~n10275 & ~n10717;
  assign n10719 = n10275 & n10717;
  assign n10720 = ~n10718 & ~n10719;
  assign n10721 = ~n10715 & ~n10720;
  assign n10722 = ~n10714 & ~n10721;
  assign n10723 = po39  & ~n10722;
  assign n10724 = ~po39  & n10722;
  assign n10725 = ~n10278 & ~n10279;
  assign n10726 = po16  & n10725;
  assign n10727 = ~n10284 & ~n10726;
  assign n10728 = n10284 & n10726;
  assign n10729 = ~n10727 & ~n10728;
  assign n10730 = ~n10724 & ~n10729;
  assign n10731 = ~n10723 & ~n10730;
  assign n10732 = po40  & ~n10731;
  assign n10733 = ~po40  & n10731;
  assign n10734 = ~n10287 & ~n10288;
  assign n10735 = po16  & n10734;
  assign n10736 = ~n10293 & ~n10735;
  assign n10737 = n10293 & n10735;
  assign n10738 = ~n10736 & ~n10737;
  assign n10739 = ~n10733 & ~n10738;
  assign n10740 = ~n10732 & ~n10739;
  assign n10741 = po41  & ~n10740;
  assign n10742 = ~po41  & n10740;
  assign n10743 = ~n10296 & ~n10297;
  assign n10744 = po16  & n10743;
  assign n10745 = ~n10302 & ~n10744;
  assign n10746 = n10302 & n10744;
  assign n10747 = ~n10745 & ~n10746;
  assign n10748 = ~n10742 & ~n10747;
  assign n10749 = ~n10741 & ~n10748;
  assign n10750 = po42  & ~n10749;
  assign n10751 = ~po42  & n10749;
  assign n10752 = ~n10305 & ~n10306;
  assign n10753 = po16  & n10752;
  assign n10754 = ~n10311 & ~n10753;
  assign n10755 = n10311 & n10753;
  assign n10756 = ~n10754 & ~n10755;
  assign n10757 = ~n10751 & ~n10756;
  assign n10758 = ~n10750 & ~n10757;
  assign n10759 = po43  & ~n10758;
  assign n10760 = ~po43  & n10758;
  assign n10761 = ~n10314 & ~n10315;
  assign n10762 = po16  & n10761;
  assign n10763 = ~n10320 & ~n10762;
  assign n10764 = n10320 & n10762;
  assign n10765 = ~n10763 & ~n10764;
  assign n10766 = ~n10760 & ~n10765;
  assign n10767 = ~n10759 & ~n10766;
  assign n10768 = po44  & ~n10767;
  assign n10769 = ~po44  & n10767;
  assign n10770 = ~n10323 & ~n10324;
  assign n10771 = po16  & n10770;
  assign n10772 = ~n10329 & ~n10771;
  assign n10773 = n10329 & n10771;
  assign n10774 = ~n10772 & ~n10773;
  assign n10775 = ~n10769 & ~n10774;
  assign n10776 = ~n10768 & ~n10775;
  assign n10777 = po45  & ~n10776;
  assign n10778 = ~po45  & n10776;
  assign n10779 = ~n10332 & ~n10333;
  assign n10780 = po16  & n10779;
  assign n10781 = ~n10338 & ~n10780;
  assign n10782 = n10338 & n10780;
  assign n10783 = ~n10781 & ~n10782;
  assign n10784 = ~n10778 & ~n10783;
  assign n10785 = ~n10777 & ~n10784;
  assign n10786 = po46  & ~n10785;
  assign n10787 = ~po46  & n10785;
  assign n10788 = ~n10341 & ~n10342;
  assign n10789 = po16  & n10788;
  assign n10790 = ~n10347 & ~n10789;
  assign n10791 = n10347 & n10789;
  assign n10792 = ~n10790 & ~n10791;
  assign n10793 = ~n10787 & ~n10792;
  assign n10794 = ~n10786 & ~n10793;
  assign n10795 = po47  & ~n10794;
  assign n10796 = ~n10350 & ~n10356;
  assign n10797 = po16  & n10796;
  assign n10798 = ~n10355 & ~n10797;
  assign n10799 = n10355 & n10797;
  assign n10800 = ~n10798 & ~n10799;
  assign n10801 = ~po47  & n10794;
  assign n10802 = ~n10800 & ~n10801;
  assign n10803 = ~n10795 & ~n10802;
  assign n10804 = po48  & ~n10803;
  assign n10805 = ~po48  & n10803;
  assign n10806 = n10366 & ~po16 ;
  assign n10807 = ~n10495 & ~n10496;
  assign n10808 = po16  & n10807;
  assign n10809 = ~n10501 & ~n10808;
  assign n10810 = n10501 & n10808;
  assign n10811 = ~n10809 & ~n10810;
  assign n10812 = ~n10521 & ~n10805;
  assign n10813 = ~n10804 & ~n10812;
  assign n10814 = po49  & ~n10813;
  assign n10815 = ~po49  & n10813;
  assign n10816 = ~n10369 & ~n10370;
  assign n10817 = po16  & n10816;
  assign n10818 = ~n10375 & ~n10817;
  assign n10819 = n10375 & n10817;
  assign n10820 = ~n10818 & ~n10819;
  assign n10821 = ~n10815 & ~n10820;
  assign n10822 = ~n10814 & ~n10821;
  assign n10823 = po50  & ~n10822;
  assign n10824 = ~po50  & n10822;
  assign n10825 = ~n10378 & ~n10379;
  assign n10826 = po16  & n10825;
  assign n10827 = ~n10384 & ~n10826;
  assign n10828 = n10384 & n10826;
  assign n10829 = ~n10827 & ~n10828;
  assign n10830 = ~n10824 & ~n10829;
  assign n10831 = ~n10823 & ~n10830;
  assign n10832 = po51  & ~n10831;
  assign n10833 = ~po51  & n10831;
  assign n10834 = ~n10387 & ~n10388;
  assign n10835 = po16  & n10834;
  assign n10836 = ~n10393 & ~n10835;
  assign n10837 = n10393 & n10835;
  assign n10838 = ~n10836 & ~n10837;
  assign n10839 = ~n10833 & ~n10838;
  assign n10840 = ~n10832 & ~n10839;
  assign n10841 = po52  & ~n10840;
  assign n10842 = ~po52  & n10840;
  assign n10843 = ~n10396 & ~n10397;
  assign n10844 = po16  & n10843;
  assign n10845 = ~n10402 & ~n10844;
  assign n10846 = n10402 & n10844;
  assign n10847 = ~n10845 & ~n10846;
  assign n10848 = ~n10842 & ~n10847;
  assign n10849 = ~n10841 & ~n10848;
  assign n10850 = po53  & ~n10849;
  assign n10851 = ~po53  & n10849;
  assign n10852 = ~n10405 & ~n10406;
  assign n10853 = po16  & n10852;
  assign n10854 = ~n10411 & ~n10853;
  assign n10855 = n10411 & n10853;
  assign n10856 = ~n10854 & ~n10855;
  assign n10857 = ~n10851 & ~n10856;
  assign n10858 = ~n10850 & ~n10857;
  assign n10859 = po54  & ~n10858;
  assign n10860 = ~po54  & n10858;
  assign n10861 = ~n10414 & ~n10415;
  assign n10862 = po16  & n10861;
  assign n10863 = ~n10420 & ~n10862;
  assign n10864 = n10420 & n10862;
  assign n10865 = ~n10863 & ~n10864;
  assign n10866 = ~n10860 & ~n10865;
  assign n10867 = ~n10859 & ~n10866;
  assign n10868 = po55  & ~n10867;
  assign n10869 = ~po55  & n10867;
  assign n10870 = ~n10423 & ~n10424;
  assign n10871 = po16  & n10870;
  assign n10872 = ~n10429 & ~n10871;
  assign n10873 = n10429 & n10871;
  assign n10874 = ~n10872 & ~n10873;
  assign n10875 = ~n10869 & ~n10874;
  assign n10876 = ~n10868 & ~n10875;
  assign n10877 = po56  & ~n10876;
  assign n10878 = ~po56  & n10876;
  assign n10879 = ~n10432 & ~n10433;
  assign n10880 = po16  & n10879;
  assign n10881 = ~n10438 & ~n10880;
  assign n10882 = n10438 & n10880;
  assign n10883 = ~n10881 & ~n10882;
  assign n10884 = ~n10878 & ~n10883;
  assign n10885 = ~n10877 & ~n10884;
  assign n10886 = po57  & ~n10885;
  assign n10887 = ~po57  & n10885;
  assign n10888 = ~n10441 & ~n10442;
  assign n10889 = po16  & n10888;
  assign n10890 = ~n10447 & ~n10889;
  assign n10891 = n10447 & n10889;
  assign n10892 = ~n10890 & ~n10891;
  assign n10893 = ~n10887 & ~n10892;
  assign n10894 = ~n10886 & ~n10893;
  assign n10895 = po58  & ~n10894;
  assign n10896 = ~po58  & n10894;
  assign n10897 = ~n10450 & ~n10451;
  assign n10898 = po16  & n10897;
  assign n10899 = ~n10456 & ~n10898;
  assign n10900 = n10456 & n10898;
  assign n10901 = ~n10899 & ~n10900;
  assign n10902 = ~n10896 & ~n10901;
  assign n10903 = ~n10895 & ~n10902;
  assign n10904 = po59  & ~n10903;
  assign n10905 = ~po59  & n10903;
  assign n10906 = ~n10459 & ~n10460;
  assign n10907 = po16  & n10906;
  assign n10908 = ~n10465 & ~n10907;
  assign n10909 = n10465 & n10907;
  assign n10910 = ~n10908 & ~n10909;
  assign n10911 = ~n10905 & ~n10910;
  assign n10912 = ~n10904 & ~n10911;
  assign n10913 = po60  & ~n10912;
  assign n10914 = ~po60  & n10912;
  assign n10915 = ~n10468 & ~n10469;
  assign n10916 = po16  & n10915;
  assign n10917 = ~n10474 & ~n10916;
  assign n10918 = n10474 & n10916;
  assign n10919 = ~n10917 & ~n10918;
  assign n10920 = ~n10914 & ~n10919;
  assign n10921 = ~n10913 & ~n10920;
  assign n10922 = po61  & ~n10921;
  assign n10923 = ~po61  & n10921;
  assign n10924 = ~n10477 & ~n10478;
  assign n10925 = po16  & n10924;
  assign n10926 = ~n10483 & ~n10925;
  assign n10927 = n10483 & n10925;
  assign n10928 = ~n10926 & ~n10927;
  assign n10929 = ~n10923 & ~n10928;
  assign n10930 = ~n10922 & ~n10929;
  assign n10931 = po62  & ~n10930;
  assign n10932 = ~po62  & n10930;
  assign n10933 = ~n10486 & ~n10487;
  assign n10934 = po16  & n10933;
  assign n10935 = ~n10492 & ~n10934;
  assign n10936 = n10492 & n10934;
  assign n10937 = ~n10935 & ~n10936;
  assign n10938 = ~n10932 & ~n10937;
  assign n10939 = ~n10931 & ~n10938;
  assign n10940 = n10811 & n10939;
  assign n10941 = ~n10811 & ~n10939;
  assign n10942 = n10505 & po16 ;
  assign n10943 = ~n10504 & ~n10942;
  assign n10944 = n10941 & n10943;
  assign n10945 = ~po63  & ~n10944;
  assign n10946 = ~n10366 & po16 ;
  assign n10947 = n10503 & ~n10946;
  assign n10948 = po63  & ~n10505;
  assign n10949 = ~n10947 & n10948;
  assign n10950 = ~n10940 & ~n10949;
  assign n10951 = ~n10945 & n10950;
  assign po15  = n10806 | ~n10951;
  assign n10953 = ~n10804 & ~n10805;
  assign n10954 = po15  & n10953;
  assign n10955 = ~n10521 & ~n10954;
  assign n10956 = n10521 & n10954;
  assign n10957 = ~n10955 & ~n10956;
  assign n10958 = pi30  & po15 ;
  assign n10959 = ~pi28  & ~pi29 ;
  assign n10960 = ~pi30  & n10959;
  assign n10961 = ~n10958 & ~n10960;
  assign n10962 = po16  & ~n10961;
  assign n10963 = ~po16  & n10961;
  assign n10964 = ~pi30  & po15 ;
  assign n10965 = pi31  & ~n10964;
  assign n10966 = ~pi31  & n10964;
  assign n10967 = ~n10965 & ~n10966;
  assign n10968 = ~n10963 & n10967;
  assign n10969 = ~n10962 & ~n10968;
  assign n10970 = po17  & ~n10969;
  assign n10971 = ~po17  & n10969;
  assign n10972 = po16  & n10951;
  assign n10973 = ~n10966 & ~n10972;
  assign n10974 = pi32  & ~n10973;
  assign n10975 = ~pi32  & n10973;
  assign n10976 = ~n10974 & ~n10975;
  assign n10977 = ~n10971 & ~n10976;
  assign n10978 = ~n10970 & ~n10977;
  assign n10979 = po18  & ~n10978;
  assign n10980 = ~po18  & n10978;
  assign n10981 = ~n10526 & ~n10527;
  assign n10982 = po15  & n10981;
  assign n10983 = n10531 & ~n10982;
  assign n10984 = ~n10531 & n10982;
  assign n10985 = ~n10983 & ~n10984;
  assign n10986 = ~n10980 & ~n10985;
  assign n10987 = ~n10979 & ~n10986;
  assign n10988 = po19  & ~n10987;
  assign n10989 = ~po19  & n10987;
  assign n10990 = ~n10534 & ~n10535;
  assign n10991 = po15  & n10990;
  assign n10992 = ~n10540 & ~n10991;
  assign n10993 = n10540 & n10991;
  assign n10994 = ~n10992 & ~n10993;
  assign n10995 = ~n10989 & ~n10994;
  assign n10996 = ~n10988 & ~n10995;
  assign n10997 = po20  & ~n10996;
  assign n10998 = ~po20  & n10996;
  assign n10999 = ~n10543 & ~n10544;
  assign n11000 = po15  & n10999;
  assign n11001 = n10549 & n11000;
  assign n11002 = ~n10549 & ~n11000;
  assign n11003 = ~n11001 & ~n11002;
  assign n11004 = ~n10998 & ~n11003;
  assign n11005 = ~n10997 & ~n11004;
  assign n11006 = po21  & ~n11005;
  assign n11007 = ~po21  & n11005;
  assign n11008 = ~n10552 & ~n10553;
  assign n11009 = po15  & n11008;
  assign n11010 = ~n10558 & ~n11009;
  assign n11011 = n10558 & n11009;
  assign n11012 = ~n11010 & ~n11011;
  assign n11013 = ~n11007 & ~n11012;
  assign n11014 = ~n11006 & ~n11013;
  assign n11015 = po22  & ~n11014;
  assign n11016 = ~po22  & n11014;
  assign n11017 = ~n10561 & ~n10562;
  assign n11018 = po15  & n11017;
  assign n11019 = ~n10567 & ~n11018;
  assign n11020 = n10567 & n11018;
  assign n11021 = ~n11019 & ~n11020;
  assign n11022 = ~n11016 & ~n11021;
  assign n11023 = ~n11015 & ~n11022;
  assign n11024 = po23  & ~n11023;
  assign n11025 = ~po23  & n11023;
  assign n11026 = ~n10570 & ~n10571;
  assign n11027 = po15  & n11026;
  assign n11028 = ~n10576 & ~n11027;
  assign n11029 = n10576 & n11027;
  assign n11030 = ~n11028 & ~n11029;
  assign n11031 = ~n11025 & ~n11030;
  assign n11032 = ~n11024 & ~n11031;
  assign n11033 = po24  & ~n11032;
  assign n11034 = ~po24  & n11032;
  assign n11035 = ~n10579 & ~n10580;
  assign n11036 = po15  & n11035;
  assign n11037 = ~n10585 & ~n11036;
  assign n11038 = n10585 & n11036;
  assign n11039 = ~n11037 & ~n11038;
  assign n11040 = ~n11034 & ~n11039;
  assign n11041 = ~n11033 & ~n11040;
  assign n11042 = po25  & ~n11041;
  assign n11043 = ~po25  & n11041;
  assign n11044 = ~n10588 & ~n10589;
  assign n11045 = po15  & n11044;
  assign n11046 = ~n10594 & ~n11045;
  assign n11047 = n10594 & n11045;
  assign n11048 = ~n11046 & ~n11047;
  assign n11049 = ~n11043 & ~n11048;
  assign n11050 = ~n11042 & ~n11049;
  assign n11051 = po26  & ~n11050;
  assign n11052 = ~po26  & n11050;
  assign n11053 = ~n10597 & ~n10598;
  assign n11054 = po15  & n11053;
  assign n11055 = ~n10603 & ~n11054;
  assign n11056 = n10603 & n11054;
  assign n11057 = ~n11055 & ~n11056;
  assign n11058 = ~n11052 & ~n11057;
  assign n11059 = ~n11051 & ~n11058;
  assign n11060 = po27  & ~n11059;
  assign n11061 = ~po27  & n11059;
  assign n11062 = ~n10606 & ~n10607;
  assign n11063 = po15  & n11062;
  assign n11064 = ~n10612 & ~n11063;
  assign n11065 = n10612 & n11063;
  assign n11066 = ~n11064 & ~n11065;
  assign n11067 = ~n11061 & ~n11066;
  assign n11068 = ~n11060 & ~n11067;
  assign n11069 = po28  & ~n11068;
  assign n11070 = ~po28  & n11068;
  assign n11071 = ~n10615 & ~n10616;
  assign n11072 = po15  & n11071;
  assign n11073 = ~n10621 & ~n11072;
  assign n11074 = n10621 & n11072;
  assign n11075 = ~n11073 & ~n11074;
  assign n11076 = ~n11070 & ~n11075;
  assign n11077 = ~n11069 & ~n11076;
  assign n11078 = po29  & ~n11077;
  assign n11079 = ~po29  & n11077;
  assign n11080 = ~n10624 & ~n10625;
  assign n11081 = po15  & n11080;
  assign n11082 = ~n10630 & ~n11081;
  assign n11083 = n10630 & n11081;
  assign n11084 = ~n11082 & ~n11083;
  assign n11085 = ~n11079 & ~n11084;
  assign n11086 = ~n11078 & ~n11085;
  assign n11087 = po30  & ~n11086;
  assign n11088 = ~po30  & n11086;
  assign n11089 = ~n10633 & ~n10634;
  assign n11090 = po15  & n11089;
  assign n11091 = ~n10639 & ~n11090;
  assign n11092 = n10639 & n11090;
  assign n11093 = ~n11091 & ~n11092;
  assign n11094 = ~n11088 & ~n11093;
  assign n11095 = ~n11087 & ~n11094;
  assign n11096 = po31  & ~n11095;
  assign n11097 = ~po31  & n11095;
  assign n11098 = ~n10642 & ~n10643;
  assign n11099 = po15  & n11098;
  assign n11100 = ~n10648 & ~n11099;
  assign n11101 = n10648 & n11099;
  assign n11102 = ~n11100 & ~n11101;
  assign n11103 = ~n11097 & ~n11102;
  assign n11104 = ~n11096 & ~n11103;
  assign n11105 = po32  & ~n11104;
  assign n11106 = ~po32  & n11104;
  assign n11107 = ~n10651 & ~n10652;
  assign n11108 = po15  & n11107;
  assign n11109 = ~n10657 & ~n11108;
  assign n11110 = n10657 & n11108;
  assign n11111 = ~n11109 & ~n11110;
  assign n11112 = ~n11106 & ~n11111;
  assign n11113 = ~n11105 & ~n11112;
  assign n11114 = po33  & ~n11113;
  assign n11115 = ~po33  & n11113;
  assign n11116 = ~n10660 & ~n10661;
  assign n11117 = po15  & n11116;
  assign n11118 = ~n10666 & ~n11117;
  assign n11119 = n10666 & n11117;
  assign n11120 = ~n11118 & ~n11119;
  assign n11121 = ~n11115 & ~n11120;
  assign n11122 = ~n11114 & ~n11121;
  assign n11123 = po34  & ~n11122;
  assign n11124 = ~po34  & n11122;
  assign n11125 = ~n10669 & ~n10670;
  assign n11126 = po15  & n11125;
  assign n11127 = ~n10675 & ~n11126;
  assign n11128 = n10675 & n11126;
  assign n11129 = ~n11127 & ~n11128;
  assign n11130 = ~n11124 & ~n11129;
  assign n11131 = ~n11123 & ~n11130;
  assign n11132 = po35  & ~n11131;
  assign n11133 = ~po35  & n11131;
  assign n11134 = ~n10678 & ~n10679;
  assign n11135 = po15  & n11134;
  assign n11136 = ~n10684 & ~n11135;
  assign n11137 = n10684 & n11135;
  assign n11138 = ~n11136 & ~n11137;
  assign n11139 = ~n11133 & ~n11138;
  assign n11140 = ~n11132 & ~n11139;
  assign n11141 = po36  & ~n11140;
  assign n11142 = ~po36  & n11140;
  assign n11143 = ~n10687 & ~n10688;
  assign n11144 = po15  & n11143;
  assign n11145 = ~n10693 & ~n11144;
  assign n11146 = n10693 & n11144;
  assign n11147 = ~n11145 & ~n11146;
  assign n11148 = ~n11142 & ~n11147;
  assign n11149 = ~n11141 & ~n11148;
  assign n11150 = po37  & ~n11149;
  assign n11151 = ~po37  & n11149;
  assign n11152 = ~n10696 & ~n10697;
  assign n11153 = po15  & n11152;
  assign n11154 = ~n10702 & ~n11153;
  assign n11155 = n10702 & n11153;
  assign n11156 = ~n11154 & ~n11155;
  assign n11157 = ~n11151 & ~n11156;
  assign n11158 = ~n11150 & ~n11157;
  assign n11159 = po38  & ~n11158;
  assign n11160 = ~po38  & n11158;
  assign n11161 = ~n10705 & ~n10706;
  assign n11162 = po15  & n11161;
  assign n11163 = ~n10711 & ~n11162;
  assign n11164 = n10711 & n11162;
  assign n11165 = ~n11163 & ~n11164;
  assign n11166 = ~n11160 & ~n11165;
  assign n11167 = ~n11159 & ~n11166;
  assign n11168 = po39  & ~n11167;
  assign n11169 = ~po39  & n11167;
  assign n11170 = ~n10714 & ~n10715;
  assign n11171 = po15  & n11170;
  assign n11172 = ~n10720 & ~n11171;
  assign n11173 = n10720 & n11171;
  assign n11174 = ~n11172 & ~n11173;
  assign n11175 = ~n11169 & ~n11174;
  assign n11176 = ~n11168 & ~n11175;
  assign n11177 = po40  & ~n11176;
  assign n11178 = ~po40  & n11176;
  assign n11179 = ~n10723 & ~n10724;
  assign n11180 = po15  & n11179;
  assign n11181 = ~n10729 & ~n11180;
  assign n11182 = n10729 & n11180;
  assign n11183 = ~n11181 & ~n11182;
  assign n11184 = ~n11178 & ~n11183;
  assign n11185 = ~n11177 & ~n11184;
  assign n11186 = po41  & ~n11185;
  assign n11187 = ~po41  & n11185;
  assign n11188 = ~n10732 & ~n10733;
  assign n11189 = po15  & n11188;
  assign n11190 = ~n10738 & ~n11189;
  assign n11191 = n10738 & n11189;
  assign n11192 = ~n11190 & ~n11191;
  assign n11193 = ~n11187 & ~n11192;
  assign n11194 = ~n11186 & ~n11193;
  assign n11195 = po42  & ~n11194;
  assign n11196 = ~po42  & n11194;
  assign n11197 = ~n10741 & ~n10742;
  assign n11198 = po15  & n11197;
  assign n11199 = ~n10747 & ~n11198;
  assign n11200 = n10747 & n11198;
  assign n11201 = ~n11199 & ~n11200;
  assign n11202 = ~n11196 & ~n11201;
  assign n11203 = ~n11195 & ~n11202;
  assign n11204 = po43  & ~n11203;
  assign n11205 = ~po43  & n11203;
  assign n11206 = ~n10750 & ~n10751;
  assign n11207 = po15  & n11206;
  assign n11208 = ~n10756 & ~n11207;
  assign n11209 = n10756 & n11207;
  assign n11210 = ~n11208 & ~n11209;
  assign n11211 = ~n11205 & ~n11210;
  assign n11212 = ~n11204 & ~n11211;
  assign n11213 = po44  & ~n11212;
  assign n11214 = ~po44  & n11212;
  assign n11215 = ~n10759 & ~n10760;
  assign n11216 = po15  & n11215;
  assign n11217 = ~n10765 & ~n11216;
  assign n11218 = n10765 & n11216;
  assign n11219 = ~n11217 & ~n11218;
  assign n11220 = ~n11214 & ~n11219;
  assign n11221 = ~n11213 & ~n11220;
  assign n11222 = po45  & ~n11221;
  assign n11223 = ~po45  & n11221;
  assign n11224 = ~n10768 & ~n10769;
  assign n11225 = po15  & n11224;
  assign n11226 = ~n10774 & ~n11225;
  assign n11227 = n10774 & n11225;
  assign n11228 = ~n11226 & ~n11227;
  assign n11229 = ~n11223 & ~n11228;
  assign n11230 = ~n11222 & ~n11229;
  assign n11231 = po46  & ~n11230;
  assign n11232 = ~po46  & n11230;
  assign n11233 = ~n10777 & ~n10778;
  assign n11234 = po15  & n11233;
  assign n11235 = ~n10783 & ~n11234;
  assign n11236 = n10783 & n11234;
  assign n11237 = ~n11235 & ~n11236;
  assign n11238 = ~n11232 & ~n11237;
  assign n11239 = ~n11231 & ~n11238;
  assign n11240 = po47  & ~n11239;
  assign n11241 = ~po47  & n11239;
  assign n11242 = ~n10786 & ~n10787;
  assign n11243 = po15  & n11242;
  assign n11244 = ~n10792 & ~n11243;
  assign n11245 = n10792 & n11243;
  assign n11246 = ~n11244 & ~n11245;
  assign n11247 = ~n11241 & ~n11246;
  assign n11248 = ~n11240 & ~n11247;
  assign n11249 = po48  & ~n11248;
  assign n11250 = ~n10795 & ~n10801;
  assign n11251 = po15  & n11250;
  assign n11252 = ~n10800 & ~n11251;
  assign n11253 = n10800 & n11251;
  assign n11254 = ~n11252 & ~n11253;
  assign n11255 = ~po48  & n11248;
  assign n11256 = ~n11254 & ~n11255;
  assign n11257 = ~n11249 & ~n11256;
  assign n11258 = po49  & ~n11257;
  assign n11259 = ~po49  & n11257;
  assign n11260 = n10811 & ~po15 ;
  assign n11261 = ~n10931 & ~n10932;
  assign n11262 = po15  & n11261;
  assign n11263 = ~n10937 & ~n11262;
  assign n11264 = n10937 & n11262;
  assign n11265 = ~n11263 & ~n11264;
  assign n11266 = ~n10957 & ~n11259;
  assign n11267 = ~n11258 & ~n11266;
  assign n11268 = po50  & ~n11267;
  assign n11269 = ~po50  & n11267;
  assign n11270 = ~n10814 & ~n10815;
  assign n11271 = po15  & n11270;
  assign n11272 = ~n10820 & ~n11271;
  assign n11273 = n10820 & n11271;
  assign n11274 = ~n11272 & ~n11273;
  assign n11275 = ~n11269 & ~n11274;
  assign n11276 = ~n11268 & ~n11275;
  assign n11277 = po51  & ~n11276;
  assign n11278 = ~po51  & n11276;
  assign n11279 = ~n10823 & ~n10824;
  assign n11280 = po15  & n11279;
  assign n11281 = ~n10829 & ~n11280;
  assign n11282 = n10829 & n11280;
  assign n11283 = ~n11281 & ~n11282;
  assign n11284 = ~n11278 & ~n11283;
  assign n11285 = ~n11277 & ~n11284;
  assign n11286 = po52  & ~n11285;
  assign n11287 = ~po52  & n11285;
  assign n11288 = ~n10832 & ~n10833;
  assign n11289 = po15  & n11288;
  assign n11290 = ~n10838 & ~n11289;
  assign n11291 = n10838 & n11289;
  assign n11292 = ~n11290 & ~n11291;
  assign n11293 = ~n11287 & ~n11292;
  assign n11294 = ~n11286 & ~n11293;
  assign n11295 = po53  & ~n11294;
  assign n11296 = ~po53  & n11294;
  assign n11297 = ~n10841 & ~n10842;
  assign n11298 = po15  & n11297;
  assign n11299 = ~n10847 & ~n11298;
  assign n11300 = n10847 & n11298;
  assign n11301 = ~n11299 & ~n11300;
  assign n11302 = ~n11296 & ~n11301;
  assign n11303 = ~n11295 & ~n11302;
  assign n11304 = po54  & ~n11303;
  assign n11305 = ~po54  & n11303;
  assign n11306 = ~n10850 & ~n10851;
  assign n11307 = po15  & n11306;
  assign n11308 = ~n10856 & ~n11307;
  assign n11309 = n10856 & n11307;
  assign n11310 = ~n11308 & ~n11309;
  assign n11311 = ~n11305 & ~n11310;
  assign n11312 = ~n11304 & ~n11311;
  assign n11313 = po55  & ~n11312;
  assign n11314 = ~po55  & n11312;
  assign n11315 = ~n10859 & ~n10860;
  assign n11316 = po15  & n11315;
  assign n11317 = ~n10865 & ~n11316;
  assign n11318 = n10865 & n11316;
  assign n11319 = ~n11317 & ~n11318;
  assign n11320 = ~n11314 & ~n11319;
  assign n11321 = ~n11313 & ~n11320;
  assign n11322 = po56  & ~n11321;
  assign n11323 = ~po56  & n11321;
  assign n11324 = ~n10868 & ~n10869;
  assign n11325 = po15  & n11324;
  assign n11326 = ~n10874 & ~n11325;
  assign n11327 = n10874 & n11325;
  assign n11328 = ~n11326 & ~n11327;
  assign n11329 = ~n11323 & ~n11328;
  assign n11330 = ~n11322 & ~n11329;
  assign n11331 = po57  & ~n11330;
  assign n11332 = ~po57  & n11330;
  assign n11333 = ~n10877 & ~n10878;
  assign n11334 = po15  & n11333;
  assign n11335 = ~n10883 & ~n11334;
  assign n11336 = n10883 & n11334;
  assign n11337 = ~n11335 & ~n11336;
  assign n11338 = ~n11332 & ~n11337;
  assign n11339 = ~n11331 & ~n11338;
  assign n11340 = po58  & ~n11339;
  assign n11341 = ~po58  & n11339;
  assign n11342 = ~n10886 & ~n10887;
  assign n11343 = po15  & n11342;
  assign n11344 = ~n10892 & ~n11343;
  assign n11345 = n10892 & n11343;
  assign n11346 = ~n11344 & ~n11345;
  assign n11347 = ~n11341 & ~n11346;
  assign n11348 = ~n11340 & ~n11347;
  assign n11349 = po59  & ~n11348;
  assign n11350 = ~po59  & n11348;
  assign n11351 = ~n10895 & ~n10896;
  assign n11352 = po15  & n11351;
  assign n11353 = ~n10901 & ~n11352;
  assign n11354 = n10901 & n11352;
  assign n11355 = ~n11353 & ~n11354;
  assign n11356 = ~n11350 & ~n11355;
  assign n11357 = ~n11349 & ~n11356;
  assign n11358 = po60  & ~n11357;
  assign n11359 = ~po60  & n11357;
  assign n11360 = ~n10904 & ~n10905;
  assign n11361 = po15  & n11360;
  assign n11362 = ~n10910 & ~n11361;
  assign n11363 = n10910 & n11361;
  assign n11364 = ~n11362 & ~n11363;
  assign n11365 = ~n11359 & ~n11364;
  assign n11366 = ~n11358 & ~n11365;
  assign n11367 = po61  & ~n11366;
  assign n11368 = ~po61  & n11366;
  assign n11369 = ~n10913 & ~n10914;
  assign n11370 = po15  & n11369;
  assign n11371 = ~n10919 & ~n11370;
  assign n11372 = n10919 & n11370;
  assign n11373 = ~n11371 & ~n11372;
  assign n11374 = ~n11368 & ~n11373;
  assign n11375 = ~n11367 & ~n11374;
  assign n11376 = po62  & ~n11375;
  assign n11377 = ~po62  & n11375;
  assign n11378 = ~n10922 & ~n10923;
  assign n11379 = po15  & n11378;
  assign n11380 = ~n10928 & ~n11379;
  assign n11381 = n10928 & n11379;
  assign n11382 = ~n11380 & ~n11381;
  assign n11383 = ~n11377 & ~n11382;
  assign n11384 = ~n11376 & ~n11383;
  assign n11385 = n11265 & n11384;
  assign n11386 = ~n11265 & ~n11384;
  assign n11387 = n10941 & po15 ;
  assign n11388 = ~n10940 & ~n11387;
  assign n11389 = n11386 & n11388;
  assign n11390 = ~po63  & ~n11389;
  assign n11391 = ~n10811 & po15 ;
  assign n11392 = n10939 & ~n11391;
  assign n11393 = po63  & ~n10941;
  assign n11394 = ~n11392 & n11393;
  assign n11395 = ~n11385 & ~n11394;
  assign n11396 = ~n11390 & n11395;
  assign po14  = n11260 | ~n11396;
  assign n11398 = ~n11258 & ~n11259;
  assign n11399 = po14  & n11398;
  assign n11400 = ~n10957 & ~n11399;
  assign n11401 = n10957 & n11399;
  assign n11402 = ~n11400 & ~n11401;
  assign n11403 = pi28  & po14 ;
  assign n11404 = ~pi26  & ~pi27 ;
  assign n11405 = ~pi28  & n11404;
  assign n11406 = ~n11403 & ~n11405;
  assign n11407 = po15  & ~n11406;
  assign n11408 = ~po15  & n11406;
  assign n11409 = ~pi28  & po14 ;
  assign n11410 = pi29  & ~n11409;
  assign n11411 = ~pi29  & n11409;
  assign n11412 = ~n11410 & ~n11411;
  assign n11413 = ~n11408 & n11412;
  assign n11414 = ~n11407 & ~n11413;
  assign n11415 = po16  & ~n11414;
  assign n11416 = ~po16  & n11414;
  assign n11417 = po15  & n11396;
  assign n11418 = ~n11411 & ~n11417;
  assign n11419 = pi30  & ~n11418;
  assign n11420 = ~pi30  & n11418;
  assign n11421 = ~n11419 & ~n11420;
  assign n11422 = ~n11416 & ~n11421;
  assign n11423 = ~n11415 & ~n11422;
  assign n11424 = po17  & ~n11423;
  assign n11425 = ~po17  & n11423;
  assign n11426 = ~n10962 & ~n10963;
  assign n11427 = po14  & n11426;
  assign n11428 = n10967 & ~n11427;
  assign n11429 = ~n10967 & n11427;
  assign n11430 = ~n11428 & ~n11429;
  assign n11431 = ~n11425 & ~n11430;
  assign n11432 = ~n11424 & ~n11431;
  assign n11433 = po18  & ~n11432;
  assign n11434 = ~po18  & n11432;
  assign n11435 = ~n10970 & ~n10971;
  assign n11436 = po14  & n11435;
  assign n11437 = ~n10976 & ~n11436;
  assign n11438 = n10976 & n11436;
  assign n11439 = ~n11437 & ~n11438;
  assign n11440 = ~n11434 & ~n11439;
  assign n11441 = ~n11433 & ~n11440;
  assign n11442 = po19  & ~n11441;
  assign n11443 = ~po19  & n11441;
  assign n11444 = ~n10979 & ~n10980;
  assign n11445 = po14  & n11444;
  assign n11446 = n10985 & n11445;
  assign n11447 = ~n10985 & ~n11445;
  assign n11448 = ~n11446 & ~n11447;
  assign n11449 = ~n11443 & ~n11448;
  assign n11450 = ~n11442 & ~n11449;
  assign n11451 = po20  & ~n11450;
  assign n11452 = ~po20  & n11450;
  assign n11453 = ~n10988 & ~n10989;
  assign n11454 = po14  & n11453;
  assign n11455 = ~n10994 & ~n11454;
  assign n11456 = n10994 & n11454;
  assign n11457 = ~n11455 & ~n11456;
  assign n11458 = ~n11452 & ~n11457;
  assign n11459 = ~n11451 & ~n11458;
  assign n11460 = po21  & ~n11459;
  assign n11461 = ~po21  & n11459;
  assign n11462 = ~n10997 & ~n10998;
  assign n11463 = po14  & n11462;
  assign n11464 = ~n11003 & ~n11463;
  assign n11465 = n11003 & n11463;
  assign n11466 = ~n11464 & ~n11465;
  assign n11467 = ~n11461 & ~n11466;
  assign n11468 = ~n11460 & ~n11467;
  assign n11469 = po22  & ~n11468;
  assign n11470 = ~po22  & n11468;
  assign n11471 = ~n11006 & ~n11007;
  assign n11472 = po14  & n11471;
  assign n11473 = ~n11012 & ~n11472;
  assign n11474 = n11012 & n11472;
  assign n11475 = ~n11473 & ~n11474;
  assign n11476 = ~n11470 & ~n11475;
  assign n11477 = ~n11469 & ~n11476;
  assign n11478 = po23  & ~n11477;
  assign n11479 = ~po23  & n11477;
  assign n11480 = ~n11015 & ~n11016;
  assign n11481 = po14  & n11480;
  assign n11482 = ~n11021 & ~n11481;
  assign n11483 = n11021 & n11481;
  assign n11484 = ~n11482 & ~n11483;
  assign n11485 = ~n11479 & ~n11484;
  assign n11486 = ~n11478 & ~n11485;
  assign n11487 = po24  & ~n11486;
  assign n11488 = ~po24  & n11486;
  assign n11489 = ~n11024 & ~n11025;
  assign n11490 = po14  & n11489;
  assign n11491 = ~n11030 & ~n11490;
  assign n11492 = n11030 & n11490;
  assign n11493 = ~n11491 & ~n11492;
  assign n11494 = ~n11488 & ~n11493;
  assign n11495 = ~n11487 & ~n11494;
  assign n11496 = po25  & ~n11495;
  assign n11497 = ~po25  & n11495;
  assign n11498 = ~n11033 & ~n11034;
  assign n11499 = po14  & n11498;
  assign n11500 = ~n11039 & ~n11499;
  assign n11501 = n11039 & n11499;
  assign n11502 = ~n11500 & ~n11501;
  assign n11503 = ~n11497 & ~n11502;
  assign n11504 = ~n11496 & ~n11503;
  assign n11505 = po26  & ~n11504;
  assign n11506 = ~po26  & n11504;
  assign n11507 = ~n11042 & ~n11043;
  assign n11508 = po14  & n11507;
  assign n11509 = ~n11048 & ~n11508;
  assign n11510 = n11048 & n11508;
  assign n11511 = ~n11509 & ~n11510;
  assign n11512 = ~n11506 & ~n11511;
  assign n11513 = ~n11505 & ~n11512;
  assign n11514 = po27  & ~n11513;
  assign n11515 = ~po27  & n11513;
  assign n11516 = ~n11051 & ~n11052;
  assign n11517 = po14  & n11516;
  assign n11518 = ~n11057 & ~n11517;
  assign n11519 = n11057 & n11517;
  assign n11520 = ~n11518 & ~n11519;
  assign n11521 = ~n11515 & ~n11520;
  assign n11522 = ~n11514 & ~n11521;
  assign n11523 = po28  & ~n11522;
  assign n11524 = ~po28  & n11522;
  assign n11525 = ~n11060 & ~n11061;
  assign n11526 = po14  & n11525;
  assign n11527 = ~n11066 & ~n11526;
  assign n11528 = n11066 & n11526;
  assign n11529 = ~n11527 & ~n11528;
  assign n11530 = ~n11524 & ~n11529;
  assign n11531 = ~n11523 & ~n11530;
  assign n11532 = po29  & ~n11531;
  assign n11533 = ~po29  & n11531;
  assign n11534 = ~n11069 & ~n11070;
  assign n11535 = po14  & n11534;
  assign n11536 = ~n11075 & ~n11535;
  assign n11537 = n11075 & n11535;
  assign n11538 = ~n11536 & ~n11537;
  assign n11539 = ~n11533 & ~n11538;
  assign n11540 = ~n11532 & ~n11539;
  assign n11541 = po30  & ~n11540;
  assign n11542 = ~po30  & n11540;
  assign n11543 = ~n11078 & ~n11079;
  assign n11544 = po14  & n11543;
  assign n11545 = ~n11084 & ~n11544;
  assign n11546 = n11084 & n11544;
  assign n11547 = ~n11545 & ~n11546;
  assign n11548 = ~n11542 & ~n11547;
  assign n11549 = ~n11541 & ~n11548;
  assign n11550 = po31  & ~n11549;
  assign n11551 = ~po31  & n11549;
  assign n11552 = ~n11087 & ~n11088;
  assign n11553 = po14  & n11552;
  assign n11554 = ~n11093 & ~n11553;
  assign n11555 = n11093 & n11553;
  assign n11556 = ~n11554 & ~n11555;
  assign n11557 = ~n11551 & ~n11556;
  assign n11558 = ~n11550 & ~n11557;
  assign n11559 = po32  & ~n11558;
  assign n11560 = ~po32  & n11558;
  assign n11561 = ~n11096 & ~n11097;
  assign n11562 = po14  & n11561;
  assign n11563 = ~n11102 & ~n11562;
  assign n11564 = n11102 & n11562;
  assign n11565 = ~n11563 & ~n11564;
  assign n11566 = ~n11560 & ~n11565;
  assign n11567 = ~n11559 & ~n11566;
  assign n11568 = po33  & ~n11567;
  assign n11569 = ~po33  & n11567;
  assign n11570 = ~n11105 & ~n11106;
  assign n11571 = po14  & n11570;
  assign n11572 = ~n11111 & ~n11571;
  assign n11573 = n11111 & n11571;
  assign n11574 = ~n11572 & ~n11573;
  assign n11575 = ~n11569 & ~n11574;
  assign n11576 = ~n11568 & ~n11575;
  assign n11577 = po34  & ~n11576;
  assign n11578 = ~po34  & n11576;
  assign n11579 = ~n11114 & ~n11115;
  assign n11580 = po14  & n11579;
  assign n11581 = ~n11120 & ~n11580;
  assign n11582 = n11120 & n11580;
  assign n11583 = ~n11581 & ~n11582;
  assign n11584 = ~n11578 & ~n11583;
  assign n11585 = ~n11577 & ~n11584;
  assign n11586 = po35  & ~n11585;
  assign n11587 = ~po35  & n11585;
  assign n11588 = ~n11123 & ~n11124;
  assign n11589 = po14  & n11588;
  assign n11590 = ~n11129 & ~n11589;
  assign n11591 = n11129 & n11589;
  assign n11592 = ~n11590 & ~n11591;
  assign n11593 = ~n11587 & ~n11592;
  assign n11594 = ~n11586 & ~n11593;
  assign n11595 = po36  & ~n11594;
  assign n11596 = ~po36  & n11594;
  assign n11597 = ~n11132 & ~n11133;
  assign n11598 = po14  & n11597;
  assign n11599 = ~n11138 & ~n11598;
  assign n11600 = n11138 & n11598;
  assign n11601 = ~n11599 & ~n11600;
  assign n11602 = ~n11596 & ~n11601;
  assign n11603 = ~n11595 & ~n11602;
  assign n11604 = po37  & ~n11603;
  assign n11605 = ~po37  & n11603;
  assign n11606 = ~n11141 & ~n11142;
  assign n11607 = po14  & n11606;
  assign n11608 = ~n11147 & ~n11607;
  assign n11609 = n11147 & n11607;
  assign n11610 = ~n11608 & ~n11609;
  assign n11611 = ~n11605 & ~n11610;
  assign n11612 = ~n11604 & ~n11611;
  assign n11613 = po38  & ~n11612;
  assign n11614 = ~po38  & n11612;
  assign n11615 = ~n11150 & ~n11151;
  assign n11616 = po14  & n11615;
  assign n11617 = ~n11156 & ~n11616;
  assign n11618 = n11156 & n11616;
  assign n11619 = ~n11617 & ~n11618;
  assign n11620 = ~n11614 & ~n11619;
  assign n11621 = ~n11613 & ~n11620;
  assign n11622 = po39  & ~n11621;
  assign n11623 = ~po39  & n11621;
  assign n11624 = ~n11159 & ~n11160;
  assign n11625 = po14  & n11624;
  assign n11626 = ~n11165 & ~n11625;
  assign n11627 = n11165 & n11625;
  assign n11628 = ~n11626 & ~n11627;
  assign n11629 = ~n11623 & ~n11628;
  assign n11630 = ~n11622 & ~n11629;
  assign n11631 = po40  & ~n11630;
  assign n11632 = ~po40  & n11630;
  assign n11633 = ~n11168 & ~n11169;
  assign n11634 = po14  & n11633;
  assign n11635 = ~n11174 & ~n11634;
  assign n11636 = n11174 & n11634;
  assign n11637 = ~n11635 & ~n11636;
  assign n11638 = ~n11632 & ~n11637;
  assign n11639 = ~n11631 & ~n11638;
  assign n11640 = po41  & ~n11639;
  assign n11641 = ~po41  & n11639;
  assign n11642 = ~n11177 & ~n11178;
  assign n11643 = po14  & n11642;
  assign n11644 = ~n11183 & ~n11643;
  assign n11645 = n11183 & n11643;
  assign n11646 = ~n11644 & ~n11645;
  assign n11647 = ~n11641 & ~n11646;
  assign n11648 = ~n11640 & ~n11647;
  assign n11649 = po42  & ~n11648;
  assign n11650 = ~po42  & n11648;
  assign n11651 = ~n11186 & ~n11187;
  assign n11652 = po14  & n11651;
  assign n11653 = ~n11192 & ~n11652;
  assign n11654 = n11192 & n11652;
  assign n11655 = ~n11653 & ~n11654;
  assign n11656 = ~n11650 & ~n11655;
  assign n11657 = ~n11649 & ~n11656;
  assign n11658 = po43  & ~n11657;
  assign n11659 = ~po43  & n11657;
  assign n11660 = ~n11195 & ~n11196;
  assign n11661 = po14  & n11660;
  assign n11662 = ~n11201 & ~n11661;
  assign n11663 = n11201 & n11661;
  assign n11664 = ~n11662 & ~n11663;
  assign n11665 = ~n11659 & ~n11664;
  assign n11666 = ~n11658 & ~n11665;
  assign n11667 = po44  & ~n11666;
  assign n11668 = ~po44  & n11666;
  assign n11669 = ~n11204 & ~n11205;
  assign n11670 = po14  & n11669;
  assign n11671 = ~n11210 & ~n11670;
  assign n11672 = n11210 & n11670;
  assign n11673 = ~n11671 & ~n11672;
  assign n11674 = ~n11668 & ~n11673;
  assign n11675 = ~n11667 & ~n11674;
  assign n11676 = po45  & ~n11675;
  assign n11677 = ~po45  & n11675;
  assign n11678 = ~n11213 & ~n11214;
  assign n11679 = po14  & n11678;
  assign n11680 = ~n11219 & ~n11679;
  assign n11681 = n11219 & n11679;
  assign n11682 = ~n11680 & ~n11681;
  assign n11683 = ~n11677 & ~n11682;
  assign n11684 = ~n11676 & ~n11683;
  assign n11685 = po46  & ~n11684;
  assign n11686 = ~po46  & n11684;
  assign n11687 = ~n11222 & ~n11223;
  assign n11688 = po14  & n11687;
  assign n11689 = ~n11228 & ~n11688;
  assign n11690 = n11228 & n11688;
  assign n11691 = ~n11689 & ~n11690;
  assign n11692 = ~n11686 & ~n11691;
  assign n11693 = ~n11685 & ~n11692;
  assign n11694 = po47  & ~n11693;
  assign n11695 = ~po47  & n11693;
  assign n11696 = ~n11231 & ~n11232;
  assign n11697 = po14  & n11696;
  assign n11698 = ~n11237 & ~n11697;
  assign n11699 = n11237 & n11697;
  assign n11700 = ~n11698 & ~n11699;
  assign n11701 = ~n11695 & ~n11700;
  assign n11702 = ~n11694 & ~n11701;
  assign n11703 = po48  & ~n11702;
  assign n11704 = ~po48  & n11702;
  assign n11705 = ~n11240 & ~n11241;
  assign n11706 = po14  & n11705;
  assign n11707 = ~n11246 & ~n11706;
  assign n11708 = n11246 & n11706;
  assign n11709 = ~n11707 & ~n11708;
  assign n11710 = ~n11704 & ~n11709;
  assign n11711 = ~n11703 & ~n11710;
  assign n11712 = po49  & ~n11711;
  assign n11713 = ~n11249 & ~n11255;
  assign n11714 = po14  & n11713;
  assign n11715 = ~n11254 & ~n11714;
  assign n11716 = n11254 & n11714;
  assign n11717 = ~n11715 & ~n11716;
  assign n11718 = ~po49  & n11711;
  assign n11719 = ~n11717 & ~n11718;
  assign n11720 = ~n11712 & ~n11719;
  assign n11721 = po50  & ~n11720;
  assign n11722 = ~po50  & n11720;
  assign n11723 = n11265 & ~po14 ;
  assign n11724 = ~n11376 & ~n11377;
  assign n11725 = po14  & n11724;
  assign n11726 = ~n11382 & ~n11725;
  assign n11727 = n11382 & n11725;
  assign n11728 = ~n11726 & ~n11727;
  assign n11729 = ~n11402 & ~n11722;
  assign n11730 = ~n11721 & ~n11729;
  assign n11731 = po51  & ~n11730;
  assign n11732 = ~po51  & n11730;
  assign n11733 = ~n11268 & ~n11269;
  assign n11734 = po14  & n11733;
  assign n11735 = ~n11274 & ~n11734;
  assign n11736 = n11274 & n11734;
  assign n11737 = ~n11735 & ~n11736;
  assign n11738 = ~n11732 & ~n11737;
  assign n11739 = ~n11731 & ~n11738;
  assign n11740 = po52  & ~n11739;
  assign n11741 = ~po52  & n11739;
  assign n11742 = ~n11277 & ~n11278;
  assign n11743 = po14  & n11742;
  assign n11744 = ~n11283 & ~n11743;
  assign n11745 = n11283 & n11743;
  assign n11746 = ~n11744 & ~n11745;
  assign n11747 = ~n11741 & ~n11746;
  assign n11748 = ~n11740 & ~n11747;
  assign n11749 = po53  & ~n11748;
  assign n11750 = ~po53  & n11748;
  assign n11751 = ~n11286 & ~n11287;
  assign n11752 = po14  & n11751;
  assign n11753 = ~n11292 & ~n11752;
  assign n11754 = n11292 & n11752;
  assign n11755 = ~n11753 & ~n11754;
  assign n11756 = ~n11750 & ~n11755;
  assign n11757 = ~n11749 & ~n11756;
  assign n11758 = po54  & ~n11757;
  assign n11759 = ~po54  & n11757;
  assign n11760 = ~n11295 & ~n11296;
  assign n11761 = po14  & n11760;
  assign n11762 = ~n11301 & ~n11761;
  assign n11763 = n11301 & n11761;
  assign n11764 = ~n11762 & ~n11763;
  assign n11765 = ~n11759 & ~n11764;
  assign n11766 = ~n11758 & ~n11765;
  assign n11767 = po55  & ~n11766;
  assign n11768 = ~po55  & n11766;
  assign n11769 = ~n11304 & ~n11305;
  assign n11770 = po14  & n11769;
  assign n11771 = ~n11310 & ~n11770;
  assign n11772 = n11310 & n11770;
  assign n11773 = ~n11771 & ~n11772;
  assign n11774 = ~n11768 & ~n11773;
  assign n11775 = ~n11767 & ~n11774;
  assign n11776 = po56  & ~n11775;
  assign n11777 = ~po56  & n11775;
  assign n11778 = ~n11313 & ~n11314;
  assign n11779 = po14  & n11778;
  assign n11780 = ~n11319 & ~n11779;
  assign n11781 = n11319 & n11779;
  assign n11782 = ~n11780 & ~n11781;
  assign n11783 = ~n11777 & ~n11782;
  assign n11784 = ~n11776 & ~n11783;
  assign n11785 = po57  & ~n11784;
  assign n11786 = ~po57  & n11784;
  assign n11787 = ~n11322 & ~n11323;
  assign n11788 = po14  & n11787;
  assign n11789 = ~n11328 & ~n11788;
  assign n11790 = n11328 & n11788;
  assign n11791 = ~n11789 & ~n11790;
  assign n11792 = ~n11786 & ~n11791;
  assign n11793 = ~n11785 & ~n11792;
  assign n11794 = po58  & ~n11793;
  assign n11795 = ~po58  & n11793;
  assign n11796 = ~n11331 & ~n11332;
  assign n11797 = po14  & n11796;
  assign n11798 = ~n11337 & ~n11797;
  assign n11799 = n11337 & n11797;
  assign n11800 = ~n11798 & ~n11799;
  assign n11801 = ~n11795 & ~n11800;
  assign n11802 = ~n11794 & ~n11801;
  assign n11803 = po59  & ~n11802;
  assign n11804 = ~po59  & n11802;
  assign n11805 = ~n11340 & ~n11341;
  assign n11806 = po14  & n11805;
  assign n11807 = ~n11346 & ~n11806;
  assign n11808 = n11346 & n11806;
  assign n11809 = ~n11807 & ~n11808;
  assign n11810 = ~n11804 & ~n11809;
  assign n11811 = ~n11803 & ~n11810;
  assign n11812 = po60  & ~n11811;
  assign n11813 = ~po60  & n11811;
  assign n11814 = ~n11349 & ~n11350;
  assign n11815 = po14  & n11814;
  assign n11816 = ~n11355 & ~n11815;
  assign n11817 = n11355 & n11815;
  assign n11818 = ~n11816 & ~n11817;
  assign n11819 = ~n11813 & ~n11818;
  assign n11820 = ~n11812 & ~n11819;
  assign n11821 = po61  & ~n11820;
  assign n11822 = ~po61  & n11820;
  assign n11823 = ~n11358 & ~n11359;
  assign n11824 = po14  & n11823;
  assign n11825 = ~n11364 & ~n11824;
  assign n11826 = n11364 & n11824;
  assign n11827 = ~n11825 & ~n11826;
  assign n11828 = ~n11822 & ~n11827;
  assign n11829 = ~n11821 & ~n11828;
  assign n11830 = po62  & ~n11829;
  assign n11831 = ~po62  & n11829;
  assign n11832 = ~n11367 & ~n11368;
  assign n11833 = po14  & n11832;
  assign n11834 = ~n11373 & ~n11833;
  assign n11835 = n11373 & n11833;
  assign n11836 = ~n11834 & ~n11835;
  assign n11837 = ~n11831 & ~n11836;
  assign n11838 = ~n11830 & ~n11837;
  assign n11839 = n11728 & n11838;
  assign n11840 = ~n11728 & ~n11838;
  assign n11841 = n11386 & po14 ;
  assign n11842 = ~n11385 & ~n11841;
  assign n11843 = n11840 & n11842;
  assign n11844 = ~po63  & ~n11843;
  assign n11845 = ~n11265 & po14 ;
  assign n11846 = n11384 & ~n11845;
  assign n11847 = po63  & ~n11386;
  assign n11848 = ~n11846 & n11847;
  assign n11849 = ~n11839 & ~n11848;
  assign n11850 = ~n11844 & n11849;
  assign po13  = n11723 | ~n11850;
  assign n11852 = ~n11721 & ~n11722;
  assign n11853 = po13  & n11852;
  assign n11854 = ~n11402 & ~n11853;
  assign n11855 = n11402 & n11853;
  assign n11856 = ~n11854 & ~n11855;
  assign n11857 = pi26  & po13 ;
  assign n11858 = ~pi24  & ~pi25 ;
  assign n11859 = ~pi26  & n11858;
  assign n11860 = ~n11857 & ~n11859;
  assign n11861 = po14  & ~n11860;
  assign n11862 = ~po14  & n11860;
  assign n11863 = ~pi26  & po13 ;
  assign n11864 = pi27  & ~n11863;
  assign n11865 = ~pi27  & n11863;
  assign n11866 = ~n11864 & ~n11865;
  assign n11867 = ~n11862 & n11866;
  assign n11868 = ~n11861 & ~n11867;
  assign n11869 = po15  & ~n11868;
  assign n11870 = ~po15  & n11868;
  assign n11871 = po14  & n11850;
  assign n11872 = ~n11865 & ~n11871;
  assign n11873 = pi28  & ~n11872;
  assign n11874 = ~pi28  & n11872;
  assign n11875 = ~n11873 & ~n11874;
  assign n11876 = ~n11870 & ~n11875;
  assign n11877 = ~n11869 & ~n11876;
  assign n11878 = po16  & ~n11877;
  assign n11879 = ~po16  & n11877;
  assign n11880 = ~n11407 & ~n11408;
  assign n11881 = po13  & n11880;
  assign n11882 = n11412 & ~n11881;
  assign n11883 = ~n11412 & n11881;
  assign n11884 = ~n11882 & ~n11883;
  assign n11885 = ~n11879 & ~n11884;
  assign n11886 = ~n11878 & ~n11885;
  assign n11887 = po17  & ~n11886;
  assign n11888 = ~po17  & n11886;
  assign n11889 = ~n11415 & ~n11416;
  assign n11890 = po13  & n11889;
  assign n11891 = ~n11421 & ~n11890;
  assign n11892 = n11421 & n11890;
  assign n11893 = ~n11891 & ~n11892;
  assign n11894 = ~n11888 & ~n11893;
  assign n11895 = ~n11887 & ~n11894;
  assign n11896 = po18  & ~n11895;
  assign n11897 = ~po18  & n11895;
  assign n11898 = ~n11424 & ~n11425;
  assign n11899 = po13  & n11898;
  assign n11900 = n11430 & n11899;
  assign n11901 = ~n11430 & ~n11899;
  assign n11902 = ~n11900 & ~n11901;
  assign n11903 = ~n11897 & ~n11902;
  assign n11904 = ~n11896 & ~n11903;
  assign n11905 = po19  & ~n11904;
  assign n11906 = ~po19  & n11904;
  assign n11907 = ~n11433 & ~n11434;
  assign n11908 = po13  & n11907;
  assign n11909 = ~n11439 & ~n11908;
  assign n11910 = n11439 & n11908;
  assign n11911 = ~n11909 & ~n11910;
  assign n11912 = ~n11906 & ~n11911;
  assign n11913 = ~n11905 & ~n11912;
  assign n11914 = po20  & ~n11913;
  assign n11915 = ~po20  & n11913;
  assign n11916 = ~n11442 & ~n11443;
  assign n11917 = po13  & n11916;
  assign n11918 = ~n11448 & ~n11917;
  assign n11919 = n11448 & n11917;
  assign n11920 = ~n11918 & ~n11919;
  assign n11921 = ~n11915 & ~n11920;
  assign n11922 = ~n11914 & ~n11921;
  assign n11923 = po21  & ~n11922;
  assign n11924 = ~po21  & n11922;
  assign n11925 = ~n11451 & ~n11452;
  assign n11926 = po13  & n11925;
  assign n11927 = ~n11457 & ~n11926;
  assign n11928 = n11457 & n11926;
  assign n11929 = ~n11927 & ~n11928;
  assign n11930 = ~n11924 & ~n11929;
  assign n11931 = ~n11923 & ~n11930;
  assign n11932 = po22  & ~n11931;
  assign n11933 = ~po22  & n11931;
  assign n11934 = ~n11460 & ~n11461;
  assign n11935 = po13  & n11934;
  assign n11936 = ~n11466 & ~n11935;
  assign n11937 = n11466 & n11935;
  assign n11938 = ~n11936 & ~n11937;
  assign n11939 = ~n11933 & ~n11938;
  assign n11940 = ~n11932 & ~n11939;
  assign n11941 = po23  & ~n11940;
  assign n11942 = ~po23  & n11940;
  assign n11943 = ~n11469 & ~n11470;
  assign n11944 = po13  & n11943;
  assign n11945 = ~n11475 & ~n11944;
  assign n11946 = n11475 & n11944;
  assign n11947 = ~n11945 & ~n11946;
  assign n11948 = ~n11942 & ~n11947;
  assign n11949 = ~n11941 & ~n11948;
  assign n11950 = po24  & ~n11949;
  assign n11951 = ~po24  & n11949;
  assign n11952 = ~n11478 & ~n11479;
  assign n11953 = po13  & n11952;
  assign n11954 = ~n11484 & ~n11953;
  assign n11955 = n11484 & n11953;
  assign n11956 = ~n11954 & ~n11955;
  assign n11957 = ~n11951 & ~n11956;
  assign n11958 = ~n11950 & ~n11957;
  assign n11959 = po25  & ~n11958;
  assign n11960 = ~po25  & n11958;
  assign n11961 = ~n11487 & ~n11488;
  assign n11962 = po13  & n11961;
  assign n11963 = ~n11493 & ~n11962;
  assign n11964 = n11493 & n11962;
  assign n11965 = ~n11963 & ~n11964;
  assign n11966 = ~n11960 & ~n11965;
  assign n11967 = ~n11959 & ~n11966;
  assign n11968 = po26  & ~n11967;
  assign n11969 = ~po26  & n11967;
  assign n11970 = ~n11496 & ~n11497;
  assign n11971 = po13  & n11970;
  assign n11972 = ~n11502 & ~n11971;
  assign n11973 = n11502 & n11971;
  assign n11974 = ~n11972 & ~n11973;
  assign n11975 = ~n11969 & ~n11974;
  assign n11976 = ~n11968 & ~n11975;
  assign n11977 = po27  & ~n11976;
  assign n11978 = ~po27  & n11976;
  assign n11979 = ~n11505 & ~n11506;
  assign n11980 = po13  & n11979;
  assign n11981 = ~n11511 & ~n11980;
  assign n11982 = n11511 & n11980;
  assign n11983 = ~n11981 & ~n11982;
  assign n11984 = ~n11978 & ~n11983;
  assign n11985 = ~n11977 & ~n11984;
  assign n11986 = po28  & ~n11985;
  assign n11987 = ~po28  & n11985;
  assign n11988 = ~n11514 & ~n11515;
  assign n11989 = po13  & n11988;
  assign n11990 = ~n11520 & ~n11989;
  assign n11991 = n11520 & n11989;
  assign n11992 = ~n11990 & ~n11991;
  assign n11993 = ~n11987 & ~n11992;
  assign n11994 = ~n11986 & ~n11993;
  assign n11995 = po29  & ~n11994;
  assign n11996 = ~po29  & n11994;
  assign n11997 = ~n11523 & ~n11524;
  assign n11998 = po13  & n11997;
  assign n11999 = ~n11529 & ~n11998;
  assign n12000 = n11529 & n11998;
  assign n12001 = ~n11999 & ~n12000;
  assign n12002 = ~n11996 & ~n12001;
  assign n12003 = ~n11995 & ~n12002;
  assign n12004 = po30  & ~n12003;
  assign n12005 = ~po30  & n12003;
  assign n12006 = ~n11532 & ~n11533;
  assign n12007 = po13  & n12006;
  assign n12008 = ~n11538 & ~n12007;
  assign n12009 = n11538 & n12007;
  assign n12010 = ~n12008 & ~n12009;
  assign n12011 = ~n12005 & ~n12010;
  assign n12012 = ~n12004 & ~n12011;
  assign n12013 = po31  & ~n12012;
  assign n12014 = ~po31  & n12012;
  assign n12015 = ~n11541 & ~n11542;
  assign n12016 = po13  & n12015;
  assign n12017 = ~n11547 & ~n12016;
  assign n12018 = n11547 & n12016;
  assign n12019 = ~n12017 & ~n12018;
  assign n12020 = ~n12014 & ~n12019;
  assign n12021 = ~n12013 & ~n12020;
  assign n12022 = po32  & ~n12021;
  assign n12023 = ~po32  & n12021;
  assign n12024 = ~n11550 & ~n11551;
  assign n12025 = po13  & n12024;
  assign n12026 = ~n11556 & ~n12025;
  assign n12027 = n11556 & n12025;
  assign n12028 = ~n12026 & ~n12027;
  assign n12029 = ~n12023 & ~n12028;
  assign n12030 = ~n12022 & ~n12029;
  assign n12031 = po33  & ~n12030;
  assign n12032 = ~po33  & n12030;
  assign n12033 = ~n11559 & ~n11560;
  assign n12034 = po13  & n12033;
  assign n12035 = ~n11565 & ~n12034;
  assign n12036 = n11565 & n12034;
  assign n12037 = ~n12035 & ~n12036;
  assign n12038 = ~n12032 & ~n12037;
  assign n12039 = ~n12031 & ~n12038;
  assign n12040 = po34  & ~n12039;
  assign n12041 = ~po34  & n12039;
  assign n12042 = ~n11568 & ~n11569;
  assign n12043 = po13  & n12042;
  assign n12044 = ~n11574 & ~n12043;
  assign n12045 = n11574 & n12043;
  assign n12046 = ~n12044 & ~n12045;
  assign n12047 = ~n12041 & ~n12046;
  assign n12048 = ~n12040 & ~n12047;
  assign n12049 = po35  & ~n12048;
  assign n12050 = ~po35  & n12048;
  assign n12051 = ~n11577 & ~n11578;
  assign n12052 = po13  & n12051;
  assign n12053 = ~n11583 & ~n12052;
  assign n12054 = n11583 & n12052;
  assign n12055 = ~n12053 & ~n12054;
  assign n12056 = ~n12050 & ~n12055;
  assign n12057 = ~n12049 & ~n12056;
  assign n12058 = po36  & ~n12057;
  assign n12059 = ~po36  & n12057;
  assign n12060 = ~n11586 & ~n11587;
  assign n12061 = po13  & n12060;
  assign n12062 = ~n11592 & ~n12061;
  assign n12063 = n11592 & n12061;
  assign n12064 = ~n12062 & ~n12063;
  assign n12065 = ~n12059 & ~n12064;
  assign n12066 = ~n12058 & ~n12065;
  assign n12067 = po37  & ~n12066;
  assign n12068 = ~po37  & n12066;
  assign n12069 = ~n11595 & ~n11596;
  assign n12070 = po13  & n12069;
  assign n12071 = ~n11601 & ~n12070;
  assign n12072 = n11601 & n12070;
  assign n12073 = ~n12071 & ~n12072;
  assign n12074 = ~n12068 & ~n12073;
  assign n12075 = ~n12067 & ~n12074;
  assign n12076 = po38  & ~n12075;
  assign n12077 = ~po38  & n12075;
  assign n12078 = ~n11604 & ~n11605;
  assign n12079 = po13  & n12078;
  assign n12080 = ~n11610 & ~n12079;
  assign n12081 = n11610 & n12079;
  assign n12082 = ~n12080 & ~n12081;
  assign n12083 = ~n12077 & ~n12082;
  assign n12084 = ~n12076 & ~n12083;
  assign n12085 = po39  & ~n12084;
  assign n12086 = ~po39  & n12084;
  assign n12087 = ~n11613 & ~n11614;
  assign n12088 = po13  & n12087;
  assign n12089 = ~n11619 & ~n12088;
  assign n12090 = n11619 & n12088;
  assign n12091 = ~n12089 & ~n12090;
  assign n12092 = ~n12086 & ~n12091;
  assign n12093 = ~n12085 & ~n12092;
  assign n12094 = po40  & ~n12093;
  assign n12095 = ~po40  & n12093;
  assign n12096 = ~n11622 & ~n11623;
  assign n12097 = po13  & n12096;
  assign n12098 = ~n11628 & ~n12097;
  assign n12099 = n11628 & n12097;
  assign n12100 = ~n12098 & ~n12099;
  assign n12101 = ~n12095 & ~n12100;
  assign n12102 = ~n12094 & ~n12101;
  assign n12103 = po41  & ~n12102;
  assign n12104 = ~po41  & n12102;
  assign n12105 = ~n11631 & ~n11632;
  assign n12106 = po13  & n12105;
  assign n12107 = ~n11637 & ~n12106;
  assign n12108 = n11637 & n12106;
  assign n12109 = ~n12107 & ~n12108;
  assign n12110 = ~n12104 & ~n12109;
  assign n12111 = ~n12103 & ~n12110;
  assign n12112 = po42  & ~n12111;
  assign n12113 = ~po42  & n12111;
  assign n12114 = ~n11640 & ~n11641;
  assign n12115 = po13  & n12114;
  assign n12116 = ~n11646 & ~n12115;
  assign n12117 = n11646 & n12115;
  assign n12118 = ~n12116 & ~n12117;
  assign n12119 = ~n12113 & ~n12118;
  assign n12120 = ~n12112 & ~n12119;
  assign n12121 = po43  & ~n12120;
  assign n12122 = ~po43  & n12120;
  assign n12123 = ~n11649 & ~n11650;
  assign n12124 = po13  & n12123;
  assign n12125 = ~n11655 & ~n12124;
  assign n12126 = n11655 & n12124;
  assign n12127 = ~n12125 & ~n12126;
  assign n12128 = ~n12122 & ~n12127;
  assign n12129 = ~n12121 & ~n12128;
  assign n12130 = po44  & ~n12129;
  assign n12131 = ~po44  & n12129;
  assign n12132 = ~n11658 & ~n11659;
  assign n12133 = po13  & n12132;
  assign n12134 = ~n11664 & ~n12133;
  assign n12135 = n11664 & n12133;
  assign n12136 = ~n12134 & ~n12135;
  assign n12137 = ~n12131 & ~n12136;
  assign n12138 = ~n12130 & ~n12137;
  assign n12139 = po45  & ~n12138;
  assign n12140 = ~po45  & n12138;
  assign n12141 = ~n11667 & ~n11668;
  assign n12142 = po13  & n12141;
  assign n12143 = ~n11673 & ~n12142;
  assign n12144 = n11673 & n12142;
  assign n12145 = ~n12143 & ~n12144;
  assign n12146 = ~n12140 & ~n12145;
  assign n12147 = ~n12139 & ~n12146;
  assign n12148 = po46  & ~n12147;
  assign n12149 = ~po46  & n12147;
  assign n12150 = ~n11676 & ~n11677;
  assign n12151 = po13  & n12150;
  assign n12152 = ~n11682 & ~n12151;
  assign n12153 = n11682 & n12151;
  assign n12154 = ~n12152 & ~n12153;
  assign n12155 = ~n12149 & ~n12154;
  assign n12156 = ~n12148 & ~n12155;
  assign n12157 = po47  & ~n12156;
  assign n12158 = ~po47  & n12156;
  assign n12159 = ~n11685 & ~n11686;
  assign n12160 = po13  & n12159;
  assign n12161 = ~n11691 & ~n12160;
  assign n12162 = n11691 & n12160;
  assign n12163 = ~n12161 & ~n12162;
  assign n12164 = ~n12158 & ~n12163;
  assign n12165 = ~n12157 & ~n12164;
  assign n12166 = po48  & ~n12165;
  assign n12167 = ~po48  & n12165;
  assign n12168 = ~n11694 & ~n11695;
  assign n12169 = po13  & n12168;
  assign n12170 = ~n11700 & ~n12169;
  assign n12171 = n11700 & n12169;
  assign n12172 = ~n12170 & ~n12171;
  assign n12173 = ~n12167 & ~n12172;
  assign n12174 = ~n12166 & ~n12173;
  assign n12175 = po49  & ~n12174;
  assign n12176 = ~po49  & n12174;
  assign n12177 = ~n11703 & ~n11704;
  assign n12178 = po13  & n12177;
  assign n12179 = ~n11709 & ~n12178;
  assign n12180 = n11709 & n12178;
  assign n12181 = ~n12179 & ~n12180;
  assign n12182 = ~n12176 & ~n12181;
  assign n12183 = ~n12175 & ~n12182;
  assign n12184 = po50  & ~n12183;
  assign n12185 = ~n11712 & ~n11718;
  assign n12186 = po13  & n12185;
  assign n12187 = ~n11717 & ~n12186;
  assign n12188 = n11717 & n12186;
  assign n12189 = ~n12187 & ~n12188;
  assign n12190 = ~po50  & n12183;
  assign n12191 = ~n12189 & ~n12190;
  assign n12192 = ~n12184 & ~n12191;
  assign n12193 = po51  & ~n12192;
  assign n12194 = ~po51  & n12192;
  assign n12195 = n11728 & ~po13 ;
  assign n12196 = ~n11830 & ~n11831;
  assign n12197 = po13  & n12196;
  assign n12198 = ~n11836 & ~n12197;
  assign n12199 = n11836 & n12197;
  assign n12200 = ~n12198 & ~n12199;
  assign n12201 = ~n11856 & ~n12194;
  assign n12202 = ~n12193 & ~n12201;
  assign n12203 = po52  & ~n12202;
  assign n12204 = ~po52  & n12202;
  assign n12205 = ~n11731 & ~n11732;
  assign n12206 = po13  & n12205;
  assign n12207 = ~n11737 & ~n12206;
  assign n12208 = n11737 & n12206;
  assign n12209 = ~n12207 & ~n12208;
  assign n12210 = ~n12204 & ~n12209;
  assign n12211 = ~n12203 & ~n12210;
  assign n12212 = po53  & ~n12211;
  assign n12213 = ~po53  & n12211;
  assign n12214 = ~n11740 & ~n11741;
  assign n12215 = po13  & n12214;
  assign n12216 = ~n11746 & ~n12215;
  assign n12217 = n11746 & n12215;
  assign n12218 = ~n12216 & ~n12217;
  assign n12219 = ~n12213 & ~n12218;
  assign n12220 = ~n12212 & ~n12219;
  assign n12221 = po54  & ~n12220;
  assign n12222 = ~po54  & n12220;
  assign n12223 = ~n11749 & ~n11750;
  assign n12224 = po13  & n12223;
  assign n12225 = ~n11755 & ~n12224;
  assign n12226 = n11755 & n12224;
  assign n12227 = ~n12225 & ~n12226;
  assign n12228 = ~n12222 & ~n12227;
  assign n12229 = ~n12221 & ~n12228;
  assign n12230 = po55  & ~n12229;
  assign n12231 = ~po55  & n12229;
  assign n12232 = ~n11758 & ~n11759;
  assign n12233 = po13  & n12232;
  assign n12234 = ~n11764 & ~n12233;
  assign n12235 = n11764 & n12233;
  assign n12236 = ~n12234 & ~n12235;
  assign n12237 = ~n12231 & ~n12236;
  assign n12238 = ~n12230 & ~n12237;
  assign n12239 = po56  & ~n12238;
  assign n12240 = ~po56  & n12238;
  assign n12241 = ~n11767 & ~n11768;
  assign n12242 = po13  & n12241;
  assign n12243 = ~n11773 & ~n12242;
  assign n12244 = n11773 & n12242;
  assign n12245 = ~n12243 & ~n12244;
  assign n12246 = ~n12240 & ~n12245;
  assign n12247 = ~n12239 & ~n12246;
  assign n12248 = po57  & ~n12247;
  assign n12249 = ~po57  & n12247;
  assign n12250 = ~n11776 & ~n11777;
  assign n12251 = po13  & n12250;
  assign n12252 = ~n11782 & ~n12251;
  assign n12253 = n11782 & n12251;
  assign n12254 = ~n12252 & ~n12253;
  assign n12255 = ~n12249 & ~n12254;
  assign n12256 = ~n12248 & ~n12255;
  assign n12257 = po58  & ~n12256;
  assign n12258 = ~po58  & n12256;
  assign n12259 = ~n11785 & ~n11786;
  assign n12260 = po13  & n12259;
  assign n12261 = ~n11791 & ~n12260;
  assign n12262 = n11791 & n12260;
  assign n12263 = ~n12261 & ~n12262;
  assign n12264 = ~n12258 & ~n12263;
  assign n12265 = ~n12257 & ~n12264;
  assign n12266 = po59  & ~n12265;
  assign n12267 = ~po59  & n12265;
  assign n12268 = ~n11794 & ~n11795;
  assign n12269 = po13  & n12268;
  assign n12270 = ~n11800 & ~n12269;
  assign n12271 = n11800 & n12269;
  assign n12272 = ~n12270 & ~n12271;
  assign n12273 = ~n12267 & ~n12272;
  assign n12274 = ~n12266 & ~n12273;
  assign n12275 = po60  & ~n12274;
  assign n12276 = ~po60  & n12274;
  assign n12277 = ~n11803 & ~n11804;
  assign n12278 = po13  & n12277;
  assign n12279 = ~n11809 & ~n12278;
  assign n12280 = n11809 & n12278;
  assign n12281 = ~n12279 & ~n12280;
  assign n12282 = ~n12276 & ~n12281;
  assign n12283 = ~n12275 & ~n12282;
  assign n12284 = po61  & ~n12283;
  assign n12285 = ~po61  & n12283;
  assign n12286 = ~n11812 & ~n11813;
  assign n12287 = po13  & n12286;
  assign n12288 = ~n11818 & ~n12287;
  assign n12289 = n11818 & n12287;
  assign n12290 = ~n12288 & ~n12289;
  assign n12291 = ~n12285 & ~n12290;
  assign n12292 = ~n12284 & ~n12291;
  assign n12293 = po62  & ~n12292;
  assign n12294 = ~po62  & n12292;
  assign n12295 = ~n11821 & ~n11822;
  assign n12296 = po13  & n12295;
  assign n12297 = ~n11827 & ~n12296;
  assign n12298 = n11827 & n12296;
  assign n12299 = ~n12297 & ~n12298;
  assign n12300 = ~n12294 & ~n12299;
  assign n12301 = ~n12293 & ~n12300;
  assign n12302 = n12200 & n12301;
  assign n12303 = ~n12200 & ~n12301;
  assign n12304 = n11840 & po13 ;
  assign n12305 = ~n11839 & ~n12304;
  assign n12306 = n12303 & n12305;
  assign n12307 = ~po63  & ~n12306;
  assign n12308 = ~n11728 & po13 ;
  assign n12309 = n11838 & ~n12308;
  assign n12310 = po63  & ~n11840;
  assign n12311 = ~n12309 & n12310;
  assign n12312 = ~n12302 & ~n12311;
  assign n12313 = ~n12307 & n12312;
  assign po12  = n12195 | ~n12313;
  assign n12315 = ~n12193 & ~n12194;
  assign n12316 = po12  & n12315;
  assign n12317 = ~n11856 & ~n12316;
  assign n12318 = n11856 & n12316;
  assign n12319 = ~n12317 & ~n12318;
  assign n12320 = pi24  & po12 ;
  assign n12321 = ~pi22  & ~pi23 ;
  assign n12322 = ~pi24  & n12321;
  assign n12323 = ~n12320 & ~n12322;
  assign n12324 = po13  & ~n12323;
  assign n12325 = ~po13  & n12323;
  assign n12326 = ~pi24  & po12 ;
  assign n12327 = pi25  & ~n12326;
  assign n12328 = ~pi25  & n12326;
  assign n12329 = ~n12327 & ~n12328;
  assign n12330 = ~n12325 & n12329;
  assign n12331 = ~n12324 & ~n12330;
  assign n12332 = po14  & ~n12331;
  assign n12333 = ~po14  & n12331;
  assign n12334 = po13  & n12313;
  assign n12335 = ~n12328 & ~n12334;
  assign n12336 = pi26  & ~n12335;
  assign n12337 = ~pi26  & n12335;
  assign n12338 = ~n12336 & ~n12337;
  assign n12339 = ~n12333 & ~n12338;
  assign n12340 = ~n12332 & ~n12339;
  assign n12341 = po15  & ~n12340;
  assign n12342 = ~po15  & n12340;
  assign n12343 = ~n11861 & ~n11862;
  assign n12344 = po12  & n12343;
  assign n12345 = n11866 & ~n12344;
  assign n12346 = ~n11866 & n12344;
  assign n12347 = ~n12345 & ~n12346;
  assign n12348 = ~n12342 & ~n12347;
  assign n12349 = ~n12341 & ~n12348;
  assign n12350 = po16  & ~n12349;
  assign n12351 = ~po16  & n12349;
  assign n12352 = ~n11869 & ~n11870;
  assign n12353 = po12  & n12352;
  assign n12354 = ~n11875 & ~n12353;
  assign n12355 = n11875 & n12353;
  assign n12356 = ~n12354 & ~n12355;
  assign n12357 = ~n12351 & ~n12356;
  assign n12358 = ~n12350 & ~n12357;
  assign n12359 = po17  & ~n12358;
  assign n12360 = ~po17  & n12358;
  assign n12361 = ~n11878 & ~n11879;
  assign n12362 = po12  & n12361;
  assign n12363 = n11884 & n12362;
  assign n12364 = ~n11884 & ~n12362;
  assign n12365 = ~n12363 & ~n12364;
  assign n12366 = ~n12360 & ~n12365;
  assign n12367 = ~n12359 & ~n12366;
  assign n12368 = po18  & ~n12367;
  assign n12369 = ~po18  & n12367;
  assign n12370 = ~n11887 & ~n11888;
  assign n12371 = po12  & n12370;
  assign n12372 = ~n11893 & ~n12371;
  assign n12373 = n11893 & n12371;
  assign n12374 = ~n12372 & ~n12373;
  assign n12375 = ~n12369 & ~n12374;
  assign n12376 = ~n12368 & ~n12375;
  assign n12377 = po19  & ~n12376;
  assign n12378 = ~po19  & n12376;
  assign n12379 = ~n11896 & ~n11897;
  assign n12380 = po12  & n12379;
  assign n12381 = ~n11902 & ~n12380;
  assign n12382 = n11902 & n12380;
  assign n12383 = ~n12381 & ~n12382;
  assign n12384 = ~n12378 & ~n12383;
  assign n12385 = ~n12377 & ~n12384;
  assign n12386 = po20  & ~n12385;
  assign n12387 = ~po20  & n12385;
  assign n12388 = ~n11905 & ~n11906;
  assign n12389 = po12  & n12388;
  assign n12390 = ~n11911 & ~n12389;
  assign n12391 = n11911 & n12389;
  assign n12392 = ~n12390 & ~n12391;
  assign n12393 = ~n12387 & ~n12392;
  assign n12394 = ~n12386 & ~n12393;
  assign n12395 = po21  & ~n12394;
  assign n12396 = ~po21  & n12394;
  assign n12397 = ~n11914 & ~n11915;
  assign n12398 = po12  & n12397;
  assign n12399 = ~n11920 & ~n12398;
  assign n12400 = n11920 & n12398;
  assign n12401 = ~n12399 & ~n12400;
  assign n12402 = ~n12396 & ~n12401;
  assign n12403 = ~n12395 & ~n12402;
  assign n12404 = po22  & ~n12403;
  assign n12405 = ~po22  & n12403;
  assign n12406 = ~n11923 & ~n11924;
  assign n12407 = po12  & n12406;
  assign n12408 = ~n11929 & ~n12407;
  assign n12409 = n11929 & n12407;
  assign n12410 = ~n12408 & ~n12409;
  assign n12411 = ~n12405 & ~n12410;
  assign n12412 = ~n12404 & ~n12411;
  assign n12413 = po23  & ~n12412;
  assign n12414 = ~po23  & n12412;
  assign n12415 = ~n11932 & ~n11933;
  assign n12416 = po12  & n12415;
  assign n12417 = ~n11938 & ~n12416;
  assign n12418 = n11938 & n12416;
  assign n12419 = ~n12417 & ~n12418;
  assign n12420 = ~n12414 & ~n12419;
  assign n12421 = ~n12413 & ~n12420;
  assign n12422 = po24  & ~n12421;
  assign n12423 = ~po24  & n12421;
  assign n12424 = ~n11941 & ~n11942;
  assign n12425 = po12  & n12424;
  assign n12426 = ~n11947 & ~n12425;
  assign n12427 = n11947 & n12425;
  assign n12428 = ~n12426 & ~n12427;
  assign n12429 = ~n12423 & ~n12428;
  assign n12430 = ~n12422 & ~n12429;
  assign n12431 = po25  & ~n12430;
  assign n12432 = ~po25  & n12430;
  assign n12433 = ~n11950 & ~n11951;
  assign n12434 = po12  & n12433;
  assign n12435 = ~n11956 & ~n12434;
  assign n12436 = n11956 & n12434;
  assign n12437 = ~n12435 & ~n12436;
  assign n12438 = ~n12432 & ~n12437;
  assign n12439 = ~n12431 & ~n12438;
  assign n12440 = po26  & ~n12439;
  assign n12441 = ~po26  & n12439;
  assign n12442 = ~n11959 & ~n11960;
  assign n12443 = po12  & n12442;
  assign n12444 = ~n11965 & ~n12443;
  assign n12445 = n11965 & n12443;
  assign n12446 = ~n12444 & ~n12445;
  assign n12447 = ~n12441 & ~n12446;
  assign n12448 = ~n12440 & ~n12447;
  assign n12449 = po27  & ~n12448;
  assign n12450 = ~po27  & n12448;
  assign n12451 = ~n11968 & ~n11969;
  assign n12452 = po12  & n12451;
  assign n12453 = ~n11974 & ~n12452;
  assign n12454 = n11974 & n12452;
  assign n12455 = ~n12453 & ~n12454;
  assign n12456 = ~n12450 & ~n12455;
  assign n12457 = ~n12449 & ~n12456;
  assign n12458 = po28  & ~n12457;
  assign n12459 = ~po28  & n12457;
  assign n12460 = ~n11977 & ~n11978;
  assign n12461 = po12  & n12460;
  assign n12462 = ~n11983 & ~n12461;
  assign n12463 = n11983 & n12461;
  assign n12464 = ~n12462 & ~n12463;
  assign n12465 = ~n12459 & ~n12464;
  assign n12466 = ~n12458 & ~n12465;
  assign n12467 = po29  & ~n12466;
  assign n12468 = ~po29  & n12466;
  assign n12469 = ~n11986 & ~n11987;
  assign n12470 = po12  & n12469;
  assign n12471 = ~n11992 & ~n12470;
  assign n12472 = n11992 & n12470;
  assign n12473 = ~n12471 & ~n12472;
  assign n12474 = ~n12468 & ~n12473;
  assign n12475 = ~n12467 & ~n12474;
  assign n12476 = po30  & ~n12475;
  assign n12477 = ~po30  & n12475;
  assign n12478 = ~n11995 & ~n11996;
  assign n12479 = po12  & n12478;
  assign n12480 = ~n12001 & ~n12479;
  assign n12481 = n12001 & n12479;
  assign n12482 = ~n12480 & ~n12481;
  assign n12483 = ~n12477 & ~n12482;
  assign n12484 = ~n12476 & ~n12483;
  assign n12485 = po31  & ~n12484;
  assign n12486 = ~po31  & n12484;
  assign n12487 = ~n12004 & ~n12005;
  assign n12488 = po12  & n12487;
  assign n12489 = ~n12010 & ~n12488;
  assign n12490 = n12010 & n12488;
  assign n12491 = ~n12489 & ~n12490;
  assign n12492 = ~n12486 & ~n12491;
  assign n12493 = ~n12485 & ~n12492;
  assign n12494 = po32  & ~n12493;
  assign n12495 = ~po32  & n12493;
  assign n12496 = ~n12013 & ~n12014;
  assign n12497 = po12  & n12496;
  assign n12498 = ~n12019 & ~n12497;
  assign n12499 = n12019 & n12497;
  assign n12500 = ~n12498 & ~n12499;
  assign n12501 = ~n12495 & ~n12500;
  assign n12502 = ~n12494 & ~n12501;
  assign n12503 = po33  & ~n12502;
  assign n12504 = ~po33  & n12502;
  assign n12505 = ~n12022 & ~n12023;
  assign n12506 = po12  & n12505;
  assign n12507 = ~n12028 & ~n12506;
  assign n12508 = n12028 & n12506;
  assign n12509 = ~n12507 & ~n12508;
  assign n12510 = ~n12504 & ~n12509;
  assign n12511 = ~n12503 & ~n12510;
  assign n12512 = po34  & ~n12511;
  assign n12513 = ~po34  & n12511;
  assign n12514 = ~n12031 & ~n12032;
  assign n12515 = po12  & n12514;
  assign n12516 = ~n12037 & ~n12515;
  assign n12517 = n12037 & n12515;
  assign n12518 = ~n12516 & ~n12517;
  assign n12519 = ~n12513 & ~n12518;
  assign n12520 = ~n12512 & ~n12519;
  assign n12521 = po35  & ~n12520;
  assign n12522 = ~po35  & n12520;
  assign n12523 = ~n12040 & ~n12041;
  assign n12524 = po12  & n12523;
  assign n12525 = ~n12046 & ~n12524;
  assign n12526 = n12046 & n12524;
  assign n12527 = ~n12525 & ~n12526;
  assign n12528 = ~n12522 & ~n12527;
  assign n12529 = ~n12521 & ~n12528;
  assign n12530 = po36  & ~n12529;
  assign n12531 = ~po36  & n12529;
  assign n12532 = ~n12049 & ~n12050;
  assign n12533 = po12  & n12532;
  assign n12534 = ~n12055 & ~n12533;
  assign n12535 = n12055 & n12533;
  assign n12536 = ~n12534 & ~n12535;
  assign n12537 = ~n12531 & ~n12536;
  assign n12538 = ~n12530 & ~n12537;
  assign n12539 = po37  & ~n12538;
  assign n12540 = ~po37  & n12538;
  assign n12541 = ~n12058 & ~n12059;
  assign n12542 = po12  & n12541;
  assign n12543 = ~n12064 & ~n12542;
  assign n12544 = n12064 & n12542;
  assign n12545 = ~n12543 & ~n12544;
  assign n12546 = ~n12540 & ~n12545;
  assign n12547 = ~n12539 & ~n12546;
  assign n12548 = po38  & ~n12547;
  assign n12549 = ~po38  & n12547;
  assign n12550 = ~n12067 & ~n12068;
  assign n12551 = po12  & n12550;
  assign n12552 = ~n12073 & ~n12551;
  assign n12553 = n12073 & n12551;
  assign n12554 = ~n12552 & ~n12553;
  assign n12555 = ~n12549 & ~n12554;
  assign n12556 = ~n12548 & ~n12555;
  assign n12557 = po39  & ~n12556;
  assign n12558 = ~po39  & n12556;
  assign n12559 = ~n12076 & ~n12077;
  assign n12560 = po12  & n12559;
  assign n12561 = ~n12082 & ~n12560;
  assign n12562 = n12082 & n12560;
  assign n12563 = ~n12561 & ~n12562;
  assign n12564 = ~n12558 & ~n12563;
  assign n12565 = ~n12557 & ~n12564;
  assign n12566 = po40  & ~n12565;
  assign n12567 = ~po40  & n12565;
  assign n12568 = ~n12085 & ~n12086;
  assign n12569 = po12  & n12568;
  assign n12570 = ~n12091 & ~n12569;
  assign n12571 = n12091 & n12569;
  assign n12572 = ~n12570 & ~n12571;
  assign n12573 = ~n12567 & ~n12572;
  assign n12574 = ~n12566 & ~n12573;
  assign n12575 = po41  & ~n12574;
  assign n12576 = ~po41  & n12574;
  assign n12577 = ~n12094 & ~n12095;
  assign n12578 = po12  & n12577;
  assign n12579 = ~n12100 & ~n12578;
  assign n12580 = n12100 & n12578;
  assign n12581 = ~n12579 & ~n12580;
  assign n12582 = ~n12576 & ~n12581;
  assign n12583 = ~n12575 & ~n12582;
  assign n12584 = po42  & ~n12583;
  assign n12585 = ~po42  & n12583;
  assign n12586 = ~n12103 & ~n12104;
  assign n12587 = po12  & n12586;
  assign n12588 = ~n12109 & ~n12587;
  assign n12589 = n12109 & n12587;
  assign n12590 = ~n12588 & ~n12589;
  assign n12591 = ~n12585 & ~n12590;
  assign n12592 = ~n12584 & ~n12591;
  assign n12593 = po43  & ~n12592;
  assign n12594 = ~po43  & n12592;
  assign n12595 = ~n12112 & ~n12113;
  assign n12596 = po12  & n12595;
  assign n12597 = ~n12118 & ~n12596;
  assign n12598 = n12118 & n12596;
  assign n12599 = ~n12597 & ~n12598;
  assign n12600 = ~n12594 & ~n12599;
  assign n12601 = ~n12593 & ~n12600;
  assign n12602 = po44  & ~n12601;
  assign n12603 = ~po44  & n12601;
  assign n12604 = ~n12121 & ~n12122;
  assign n12605 = po12  & n12604;
  assign n12606 = ~n12127 & ~n12605;
  assign n12607 = n12127 & n12605;
  assign n12608 = ~n12606 & ~n12607;
  assign n12609 = ~n12603 & ~n12608;
  assign n12610 = ~n12602 & ~n12609;
  assign n12611 = po45  & ~n12610;
  assign n12612 = ~po45  & n12610;
  assign n12613 = ~n12130 & ~n12131;
  assign n12614 = po12  & n12613;
  assign n12615 = ~n12136 & ~n12614;
  assign n12616 = n12136 & n12614;
  assign n12617 = ~n12615 & ~n12616;
  assign n12618 = ~n12612 & ~n12617;
  assign n12619 = ~n12611 & ~n12618;
  assign n12620 = po46  & ~n12619;
  assign n12621 = ~po46  & n12619;
  assign n12622 = ~n12139 & ~n12140;
  assign n12623 = po12  & n12622;
  assign n12624 = ~n12145 & ~n12623;
  assign n12625 = n12145 & n12623;
  assign n12626 = ~n12624 & ~n12625;
  assign n12627 = ~n12621 & ~n12626;
  assign n12628 = ~n12620 & ~n12627;
  assign n12629 = po47  & ~n12628;
  assign n12630 = ~po47  & n12628;
  assign n12631 = ~n12148 & ~n12149;
  assign n12632 = po12  & n12631;
  assign n12633 = ~n12154 & ~n12632;
  assign n12634 = n12154 & n12632;
  assign n12635 = ~n12633 & ~n12634;
  assign n12636 = ~n12630 & ~n12635;
  assign n12637 = ~n12629 & ~n12636;
  assign n12638 = po48  & ~n12637;
  assign n12639 = ~po48  & n12637;
  assign n12640 = ~n12157 & ~n12158;
  assign n12641 = po12  & n12640;
  assign n12642 = ~n12163 & ~n12641;
  assign n12643 = n12163 & n12641;
  assign n12644 = ~n12642 & ~n12643;
  assign n12645 = ~n12639 & ~n12644;
  assign n12646 = ~n12638 & ~n12645;
  assign n12647 = po49  & ~n12646;
  assign n12648 = ~po49  & n12646;
  assign n12649 = ~n12166 & ~n12167;
  assign n12650 = po12  & n12649;
  assign n12651 = ~n12172 & ~n12650;
  assign n12652 = n12172 & n12650;
  assign n12653 = ~n12651 & ~n12652;
  assign n12654 = ~n12648 & ~n12653;
  assign n12655 = ~n12647 & ~n12654;
  assign n12656 = po50  & ~n12655;
  assign n12657 = ~po50  & n12655;
  assign n12658 = ~n12175 & ~n12176;
  assign n12659 = po12  & n12658;
  assign n12660 = ~n12181 & ~n12659;
  assign n12661 = n12181 & n12659;
  assign n12662 = ~n12660 & ~n12661;
  assign n12663 = ~n12657 & ~n12662;
  assign n12664 = ~n12656 & ~n12663;
  assign n12665 = po51  & ~n12664;
  assign n12666 = ~n12184 & ~n12190;
  assign n12667 = po12  & n12666;
  assign n12668 = ~n12189 & ~n12667;
  assign n12669 = n12189 & n12667;
  assign n12670 = ~n12668 & ~n12669;
  assign n12671 = ~po51  & n12664;
  assign n12672 = ~n12670 & ~n12671;
  assign n12673 = ~n12665 & ~n12672;
  assign n12674 = po52  & ~n12673;
  assign n12675 = ~po52  & n12673;
  assign n12676 = n12200 & ~po12 ;
  assign n12677 = ~n12293 & ~n12294;
  assign n12678 = po12  & n12677;
  assign n12679 = ~n12299 & ~n12678;
  assign n12680 = n12299 & n12678;
  assign n12681 = ~n12679 & ~n12680;
  assign n12682 = ~n12319 & ~n12675;
  assign n12683 = ~n12674 & ~n12682;
  assign n12684 = po53  & ~n12683;
  assign n12685 = ~po53  & n12683;
  assign n12686 = ~n12203 & ~n12204;
  assign n12687 = po12  & n12686;
  assign n12688 = ~n12209 & ~n12687;
  assign n12689 = n12209 & n12687;
  assign n12690 = ~n12688 & ~n12689;
  assign n12691 = ~n12685 & ~n12690;
  assign n12692 = ~n12684 & ~n12691;
  assign n12693 = po54  & ~n12692;
  assign n12694 = ~po54  & n12692;
  assign n12695 = ~n12212 & ~n12213;
  assign n12696 = po12  & n12695;
  assign n12697 = ~n12218 & ~n12696;
  assign n12698 = n12218 & n12696;
  assign n12699 = ~n12697 & ~n12698;
  assign n12700 = ~n12694 & ~n12699;
  assign n12701 = ~n12693 & ~n12700;
  assign n12702 = po55  & ~n12701;
  assign n12703 = ~po55  & n12701;
  assign n12704 = ~n12221 & ~n12222;
  assign n12705 = po12  & n12704;
  assign n12706 = ~n12227 & ~n12705;
  assign n12707 = n12227 & n12705;
  assign n12708 = ~n12706 & ~n12707;
  assign n12709 = ~n12703 & ~n12708;
  assign n12710 = ~n12702 & ~n12709;
  assign n12711 = po56  & ~n12710;
  assign n12712 = ~po56  & n12710;
  assign n12713 = ~n12230 & ~n12231;
  assign n12714 = po12  & n12713;
  assign n12715 = ~n12236 & ~n12714;
  assign n12716 = n12236 & n12714;
  assign n12717 = ~n12715 & ~n12716;
  assign n12718 = ~n12712 & ~n12717;
  assign n12719 = ~n12711 & ~n12718;
  assign n12720 = po57  & ~n12719;
  assign n12721 = ~po57  & n12719;
  assign n12722 = ~n12239 & ~n12240;
  assign n12723 = po12  & n12722;
  assign n12724 = ~n12245 & ~n12723;
  assign n12725 = n12245 & n12723;
  assign n12726 = ~n12724 & ~n12725;
  assign n12727 = ~n12721 & ~n12726;
  assign n12728 = ~n12720 & ~n12727;
  assign n12729 = po58  & ~n12728;
  assign n12730 = ~po58  & n12728;
  assign n12731 = ~n12248 & ~n12249;
  assign n12732 = po12  & n12731;
  assign n12733 = ~n12254 & ~n12732;
  assign n12734 = n12254 & n12732;
  assign n12735 = ~n12733 & ~n12734;
  assign n12736 = ~n12730 & ~n12735;
  assign n12737 = ~n12729 & ~n12736;
  assign n12738 = po59  & ~n12737;
  assign n12739 = ~po59  & n12737;
  assign n12740 = ~n12257 & ~n12258;
  assign n12741 = po12  & n12740;
  assign n12742 = ~n12263 & ~n12741;
  assign n12743 = n12263 & n12741;
  assign n12744 = ~n12742 & ~n12743;
  assign n12745 = ~n12739 & ~n12744;
  assign n12746 = ~n12738 & ~n12745;
  assign n12747 = po60  & ~n12746;
  assign n12748 = ~po60  & n12746;
  assign n12749 = ~n12266 & ~n12267;
  assign n12750 = po12  & n12749;
  assign n12751 = ~n12272 & ~n12750;
  assign n12752 = n12272 & n12750;
  assign n12753 = ~n12751 & ~n12752;
  assign n12754 = ~n12748 & ~n12753;
  assign n12755 = ~n12747 & ~n12754;
  assign n12756 = po61  & ~n12755;
  assign n12757 = ~po61  & n12755;
  assign n12758 = ~n12275 & ~n12276;
  assign n12759 = po12  & n12758;
  assign n12760 = ~n12281 & ~n12759;
  assign n12761 = n12281 & n12759;
  assign n12762 = ~n12760 & ~n12761;
  assign n12763 = ~n12757 & ~n12762;
  assign n12764 = ~n12756 & ~n12763;
  assign n12765 = po62  & ~n12764;
  assign n12766 = ~po62  & n12764;
  assign n12767 = ~n12284 & ~n12285;
  assign n12768 = po12  & n12767;
  assign n12769 = ~n12290 & ~n12768;
  assign n12770 = n12290 & n12768;
  assign n12771 = ~n12769 & ~n12770;
  assign n12772 = ~n12766 & ~n12771;
  assign n12773 = ~n12765 & ~n12772;
  assign n12774 = n12681 & n12773;
  assign n12775 = ~n12681 & ~n12773;
  assign n12776 = n12303 & po12 ;
  assign n12777 = ~n12302 & ~n12776;
  assign n12778 = n12775 & n12777;
  assign n12779 = ~po63  & ~n12778;
  assign n12780 = ~n12200 & po12 ;
  assign n12781 = n12301 & ~n12780;
  assign n12782 = po63  & ~n12303;
  assign n12783 = ~n12781 & n12782;
  assign n12784 = ~n12774 & ~n12783;
  assign n12785 = ~n12779 & n12784;
  assign po11  = n12676 | ~n12785;
  assign n12787 = ~n12674 & ~n12675;
  assign n12788 = po11  & n12787;
  assign n12789 = ~n12319 & ~n12788;
  assign n12790 = n12319 & n12788;
  assign n12791 = ~n12789 & ~n12790;
  assign n12792 = pi22  & po11 ;
  assign n12793 = ~pi20  & ~pi21 ;
  assign n12794 = ~pi22  & n12793;
  assign n12795 = ~n12792 & ~n12794;
  assign n12796 = po12  & ~n12795;
  assign n12797 = ~po12  & n12795;
  assign n12798 = ~pi22  & po11 ;
  assign n12799 = pi23  & ~n12798;
  assign n12800 = ~pi23  & n12798;
  assign n12801 = ~n12799 & ~n12800;
  assign n12802 = ~n12797 & n12801;
  assign n12803 = ~n12796 & ~n12802;
  assign n12804 = po13  & ~n12803;
  assign n12805 = ~po13  & n12803;
  assign n12806 = po12  & n12785;
  assign n12807 = ~n12800 & ~n12806;
  assign n12808 = pi24  & ~n12807;
  assign n12809 = ~pi24  & n12807;
  assign n12810 = ~n12808 & ~n12809;
  assign n12811 = ~n12805 & ~n12810;
  assign n12812 = ~n12804 & ~n12811;
  assign n12813 = po14  & ~n12812;
  assign n12814 = ~po14  & n12812;
  assign n12815 = ~n12324 & ~n12325;
  assign n12816 = po11  & n12815;
  assign n12817 = n12329 & ~n12816;
  assign n12818 = ~n12329 & n12816;
  assign n12819 = ~n12817 & ~n12818;
  assign n12820 = ~n12814 & ~n12819;
  assign n12821 = ~n12813 & ~n12820;
  assign n12822 = po15  & ~n12821;
  assign n12823 = ~po15  & n12821;
  assign n12824 = ~n12332 & ~n12333;
  assign n12825 = po11  & n12824;
  assign n12826 = ~n12338 & ~n12825;
  assign n12827 = n12338 & n12825;
  assign n12828 = ~n12826 & ~n12827;
  assign n12829 = ~n12823 & ~n12828;
  assign n12830 = ~n12822 & ~n12829;
  assign n12831 = po16  & ~n12830;
  assign n12832 = ~po16  & n12830;
  assign n12833 = ~n12341 & ~n12342;
  assign n12834 = po11  & n12833;
  assign n12835 = n12347 & n12834;
  assign n12836 = ~n12347 & ~n12834;
  assign n12837 = ~n12835 & ~n12836;
  assign n12838 = ~n12832 & ~n12837;
  assign n12839 = ~n12831 & ~n12838;
  assign n12840 = po17  & ~n12839;
  assign n12841 = ~po17  & n12839;
  assign n12842 = ~n12350 & ~n12351;
  assign n12843 = po11  & n12842;
  assign n12844 = ~n12356 & ~n12843;
  assign n12845 = n12356 & n12843;
  assign n12846 = ~n12844 & ~n12845;
  assign n12847 = ~n12841 & ~n12846;
  assign n12848 = ~n12840 & ~n12847;
  assign n12849 = po18  & ~n12848;
  assign n12850 = ~po18  & n12848;
  assign n12851 = ~n12359 & ~n12360;
  assign n12852 = po11  & n12851;
  assign n12853 = ~n12365 & ~n12852;
  assign n12854 = n12365 & n12852;
  assign n12855 = ~n12853 & ~n12854;
  assign n12856 = ~n12850 & ~n12855;
  assign n12857 = ~n12849 & ~n12856;
  assign n12858 = po19  & ~n12857;
  assign n12859 = ~po19  & n12857;
  assign n12860 = ~n12368 & ~n12369;
  assign n12861 = po11  & n12860;
  assign n12862 = ~n12374 & ~n12861;
  assign n12863 = n12374 & n12861;
  assign n12864 = ~n12862 & ~n12863;
  assign n12865 = ~n12859 & ~n12864;
  assign n12866 = ~n12858 & ~n12865;
  assign n12867 = po20  & ~n12866;
  assign n12868 = ~po20  & n12866;
  assign n12869 = ~n12377 & ~n12378;
  assign n12870 = po11  & n12869;
  assign n12871 = ~n12383 & ~n12870;
  assign n12872 = n12383 & n12870;
  assign n12873 = ~n12871 & ~n12872;
  assign n12874 = ~n12868 & ~n12873;
  assign n12875 = ~n12867 & ~n12874;
  assign n12876 = po21  & ~n12875;
  assign n12877 = ~po21  & n12875;
  assign n12878 = ~n12386 & ~n12387;
  assign n12879 = po11  & n12878;
  assign n12880 = ~n12392 & ~n12879;
  assign n12881 = n12392 & n12879;
  assign n12882 = ~n12880 & ~n12881;
  assign n12883 = ~n12877 & ~n12882;
  assign n12884 = ~n12876 & ~n12883;
  assign n12885 = po22  & ~n12884;
  assign n12886 = ~po22  & n12884;
  assign n12887 = ~n12395 & ~n12396;
  assign n12888 = po11  & n12887;
  assign n12889 = ~n12401 & ~n12888;
  assign n12890 = n12401 & n12888;
  assign n12891 = ~n12889 & ~n12890;
  assign n12892 = ~n12886 & ~n12891;
  assign n12893 = ~n12885 & ~n12892;
  assign n12894 = po23  & ~n12893;
  assign n12895 = ~po23  & n12893;
  assign n12896 = ~n12404 & ~n12405;
  assign n12897 = po11  & n12896;
  assign n12898 = ~n12410 & ~n12897;
  assign n12899 = n12410 & n12897;
  assign n12900 = ~n12898 & ~n12899;
  assign n12901 = ~n12895 & ~n12900;
  assign n12902 = ~n12894 & ~n12901;
  assign n12903 = po24  & ~n12902;
  assign n12904 = ~po24  & n12902;
  assign n12905 = ~n12413 & ~n12414;
  assign n12906 = po11  & n12905;
  assign n12907 = ~n12419 & ~n12906;
  assign n12908 = n12419 & n12906;
  assign n12909 = ~n12907 & ~n12908;
  assign n12910 = ~n12904 & ~n12909;
  assign n12911 = ~n12903 & ~n12910;
  assign n12912 = po25  & ~n12911;
  assign n12913 = ~po25  & n12911;
  assign n12914 = ~n12422 & ~n12423;
  assign n12915 = po11  & n12914;
  assign n12916 = ~n12428 & ~n12915;
  assign n12917 = n12428 & n12915;
  assign n12918 = ~n12916 & ~n12917;
  assign n12919 = ~n12913 & ~n12918;
  assign n12920 = ~n12912 & ~n12919;
  assign n12921 = po26  & ~n12920;
  assign n12922 = ~po26  & n12920;
  assign n12923 = ~n12431 & ~n12432;
  assign n12924 = po11  & n12923;
  assign n12925 = ~n12437 & ~n12924;
  assign n12926 = n12437 & n12924;
  assign n12927 = ~n12925 & ~n12926;
  assign n12928 = ~n12922 & ~n12927;
  assign n12929 = ~n12921 & ~n12928;
  assign n12930 = po27  & ~n12929;
  assign n12931 = ~po27  & n12929;
  assign n12932 = ~n12440 & ~n12441;
  assign n12933 = po11  & n12932;
  assign n12934 = ~n12446 & ~n12933;
  assign n12935 = n12446 & n12933;
  assign n12936 = ~n12934 & ~n12935;
  assign n12937 = ~n12931 & ~n12936;
  assign n12938 = ~n12930 & ~n12937;
  assign n12939 = po28  & ~n12938;
  assign n12940 = ~po28  & n12938;
  assign n12941 = ~n12449 & ~n12450;
  assign n12942 = po11  & n12941;
  assign n12943 = ~n12455 & ~n12942;
  assign n12944 = n12455 & n12942;
  assign n12945 = ~n12943 & ~n12944;
  assign n12946 = ~n12940 & ~n12945;
  assign n12947 = ~n12939 & ~n12946;
  assign n12948 = po29  & ~n12947;
  assign n12949 = ~po29  & n12947;
  assign n12950 = ~n12458 & ~n12459;
  assign n12951 = po11  & n12950;
  assign n12952 = ~n12464 & ~n12951;
  assign n12953 = n12464 & n12951;
  assign n12954 = ~n12952 & ~n12953;
  assign n12955 = ~n12949 & ~n12954;
  assign n12956 = ~n12948 & ~n12955;
  assign n12957 = po30  & ~n12956;
  assign n12958 = ~po30  & n12956;
  assign n12959 = ~n12467 & ~n12468;
  assign n12960 = po11  & n12959;
  assign n12961 = ~n12473 & ~n12960;
  assign n12962 = n12473 & n12960;
  assign n12963 = ~n12961 & ~n12962;
  assign n12964 = ~n12958 & ~n12963;
  assign n12965 = ~n12957 & ~n12964;
  assign n12966 = po31  & ~n12965;
  assign n12967 = ~po31  & n12965;
  assign n12968 = ~n12476 & ~n12477;
  assign n12969 = po11  & n12968;
  assign n12970 = ~n12482 & ~n12969;
  assign n12971 = n12482 & n12969;
  assign n12972 = ~n12970 & ~n12971;
  assign n12973 = ~n12967 & ~n12972;
  assign n12974 = ~n12966 & ~n12973;
  assign n12975 = po32  & ~n12974;
  assign n12976 = ~po32  & n12974;
  assign n12977 = ~n12485 & ~n12486;
  assign n12978 = po11  & n12977;
  assign n12979 = ~n12491 & ~n12978;
  assign n12980 = n12491 & n12978;
  assign n12981 = ~n12979 & ~n12980;
  assign n12982 = ~n12976 & ~n12981;
  assign n12983 = ~n12975 & ~n12982;
  assign n12984 = po33  & ~n12983;
  assign n12985 = ~po33  & n12983;
  assign n12986 = ~n12494 & ~n12495;
  assign n12987 = po11  & n12986;
  assign n12988 = ~n12500 & ~n12987;
  assign n12989 = n12500 & n12987;
  assign n12990 = ~n12988 & ~n12989;
  assign n12991 = ~n12985 & ~n12990;
  assign n12992 = ~n12984 & ~n12991;
  assign n12993 = po34  & ~n12992;
  assign n12994 = ~po34  & n12992;
  assign n12995 = ~n12503 & ~n12504;
  assign n12996 = po11  & n12995;
  assign n12997 = ~n12509 & ~n12996;
  assign n12998 = n12509 & n12996;
  assign n12999 = ~n12997 & ~n12998;
  assign n13000 = ~n12994 & ~n12999;
  assign n13001 = ~n12993 & ~n13000;
  assign n13002 = po35  & ~n13001;
  assign n13003 = ~po35  & n13001;
  assign n13004 = ~n12512 & ~n12513;
  assign n13005 = po11  & n13004;
  assign n13006 = ~n12518 & ~n13005;
  assign n13007 = n12518 & n13005;
  assign n13008 = ~n13006 & ~n13007;
  assign n13009 = ~n13003 & ~n13008;
  assign n13010 = ~n13002 & ~n13009;
  assign n13011 = po36  & ~n13010;
  assign n13012 = ~po36  & n13010;
  assign n13013 = ~n12521 & ~n12522;
  assign n13014 = po11  & n13013;
  assign n13015 = ~n12527 & ~n13014;
  assign n13016 = n12527 & n13014;
  assign n13017 = ~n13015 & ~n13016;
  assign n13018 = ~n13012 & ~n13017;
  assign n13019 = ~n13011 & ~n13018;
  assign n13020 = po37  & ~n13019;
  assign n13021 = ~po37  & n13019;
  assign n13022 = ~n12530 & ~n12531;
  assign n13023 = po11  & n13022;
  assign n13024 = ~n12536 & ~n13023;
  assign n13025 = n12536 & n13023;
  assign n13026 = ~n13024 & ~n13025;
  assign n13027 = ~n13021 & ~n13026;
  assign n13028 = ~n13020 & ~n13027;
  assign n13029 = po38  & ~n13028;
  assign n13030 = ~po38  & n13028;
  assign n13031 = ~n12539 & ~n12540;
  assign n13032 = po11  & n13031;
  assign n13033 = ~n12545 & ~n13032;
  assign n13034 = n12545 & n13032;
  assign n13035 = ~n13033 & ~n13034;
  assign n13036 = ~n13030 & ~n13035;
  assign n13037 = ~n13029 & ~n13036;
  assign n13038 = po39  & ~n13037;
  assign n13039 = ~po39  & n13037;
  assign n13040 = ~n12548 & ~n12549;
  assign n13041 = po11  & n13040;
  assign n13042 = ~n12554 & ~n13041;
  assign n13043 = n12554 & n13041;
  assign n13044 = ~n13042 & ~n13043;
  assign n13045 = ~n13039 & ~n13044;
  assign n13046 = ~n13038 & ~n13045;
  assign n13047 = po40  & ~n13046;
  assign n13048 = ~po40  & n13046;
  assign n13049 = ~n12557 & ~n12558;
  assign n13050 = po11  & n13049;
  assign n13051 = ~n12563 & ~n13050;
  assign n13052 = n12563 & n13050;
  assign n13053 = ~n13051 & ~n13052;
  assign n13054 = ~n13048 & ~n13053;
  assign n13055 = ~n13047 & ~n13054;
  assign n13056 = po41  & ~n13055;
  assign n13057 = ~po41  & n13055;
  assign n13058 = ~n12566 & ~n12567;
  assign n13059 = po11  & n13058;
  assign n13060 = ~n12572 & ~n13059;
  assign n13061 = n12572 & n13059;
  assign n13062 = ~n13060 & ~n13061;
  assign n13063 = ~n13057 & ~n13062;
  assign n13064 = ~n13056 & ~n13063;
  assign n13065 = po42  & ~n13064;
  assign n13066 = ~po42  & n13064;
  assign n13067 = ~n12575 & ~n12576;
  assign n13068 = po11  & n13067;
  assign n13069 = ~n12581 & ~n13068;
  assign n13070 = n12581 & n13068;
  assign n13071 = ~n13069 & ~n13070;
  assign n13072 = ~n13066 & ~n13071;
  assign n13073 = ~n13065 & ~n13072;
  assign n13074 = po43  & ~n13073;
  assign n13075 = ~po43  & n13073;
  assign n13076 = ~n12584 & ~n12585;
  assign n13077 = po11  & n13076;
  assign n13078 = ~n12590 & ~n13077;
  assign n13079 = n12590 & n13077;
  assign n13080 = ~n13078 & ~n13079;
  assign n13081 = ~n13075 & ~n13080;
  assign n13082 = ~n13074 & ~n13081;
  assign n13083 = po44  & ~n13082;
  assign n13084 = ~po44  & n13082;
  assign n13085 = ~n12593 & ~n12594;
  assign n13086 = po11  & n13085;
  assign n13087 = ~n12599 & ~n13086;
  assign n13088 = n12599 & n13086;
  assign n13089 = ~n13087 & ~n13088;
  assign n13090 = ~n13084 & ~n13089;
  assign n13091 = ~n13083 & ~n13090;
  assign n13092 = po45  & ~n13091;
  assign n13093 = ~po45  & n13091;
  assign n13094 = ~n12602 & ~n12603;
  assign n13095 = po11  & n13094;
  assign n13096 = ~n12608 & ~n13095;
  assign n13097 = n12608 & n13095;
  assign n13098 = ~n13096 & ~n13097;
  assign n13099 = ~n13093 & ~n13098;
  assign n13100 = ~n13092 & ~n13099;
  assign n13101 = po46  & ~n13100;
  assign n13102 = ~po46  & n13100;
  assign n13103 = ~n12611 & ~n12612;
  assign n13104 = po11  & n13103;
  assign n13105 = ~n12617 & ~n13104;
  assign n13106 = n12617 & n13104;
  assign n13107 = ~n13105 & ~n13106;
  assign n13108 = ~n13102 & ~n13107;
  assign n13109 = ~n13101 & ~n13108;
  assign n13110 = po47  & ~n13109;
  assign n13111 = ~po47  & n13109;
  assign n13112 = ~n12620 & ~n12621;
  assign n13113 = po11  & n13112;
  assign n13114 = ~n12626 & ~n13113;
  assign n13115 = n12626 & n13113;
  assign n13116 = ~n13114 & ~n13115;
  assign n13117 = ~n13111 & ~n13116;
  assign n13118 = ~n13110 & ~n13117;
  assign n13119 = po48  & ~n13118;
  assign n13120 = ~po48  & n13118;
  assign n13121 = ~n12629 & ~n12630;
  assign n13122 = po11  & n13121;
  assign n13123 = ~n12635 & ~n13122;
  assign n13124 = n12635 & n13122;
  assign n13125 = ~n13123 & ~n13124;
  assign n13126 = ~n13120 & ~n13125;
  assign n13127 = ~n13119 & ~n13126;
  assign n13128 = po49  & ~n13127;
  assign n13129 = ~po49  & n13127;
  assign n13130 = ~n12638 & ~n12639;
  assign n13131 = po11  & n13130;
  assign n13132 = ~n12644 & ~n13131;
  assign n13133 = n12644 & n13131;
  assign n13134 = ~n13132 & ~n13133;
  assign n13135 = ~n13129 & ~n13134;
  assign n13136 = ~n13128 & ~n13135;
  assign n13137 = po50  & ~n13136;
  assign n13138 = ~po50  & n13136;
  assign n13139 = ~n12647 & ~n12648;
  assign n13140 = po11  & n13139;
  assign n13141 = ~n12653 & ~n13140;
  assign n13142 = n12653 & n13140;
  assign n13143 = ~n13141 & ~n13142;
  assign n13144 = ~n13138 & ~n13143;
  assign n13145 = ~n13137 & ~n13144;
  assign n13146 = po51  & ~n13145;
  assign n13147 = ~po51  & n13145;
  assign n13148 = ~n12656 & ~n12657;
  assign n13149 = po11  & n13148;
  assign n13150 = ~n12662 & ~n13149;
  assign n13151 = n12662 & n13149;
  assign n13152 = ~n13150 & ~n13151;
  assign n13153 = ~n13147 & ~n13152;
  assign n13154 = ~n13146 & ~n13153;
  assign n13155 = po52  & ~n13154;
  assign n13156 = ~n12665 & ~n12671;
  assign n13157 = po11  & n13156;
  assign n13158 = ~n12670 & ~n13157;
  assign n13159 = n12670 & n13157;
  assign n13160 = ~n13158 & ~n13159;
  assign n13161 = ~po52  & n13154;
  assign n13162 = ~n13160 & ~n13161;
  assign n13163 = ~n13155 & ~n13162;
  assign n13164 = po53  & ~n13163;
  assign n13165 = ~po53  & n13163;
  assign n13166 = n12681 & ~po11 ;
  assign n13167 = ~n12765 & ~n12766;
  assign n13168 = po11  & n13167;
  assign n13169 = ~n12771 & ~n13168;
  assign n13170 = n12771 & n13168;
  assign n13171 = ~n13169 & ~n13170;
  assign n13172 = ~n12791 & ~n13165;
  assign n13173 = ~n13164 & ~n13172;
  assign n13174 = po54  & ~n13173;
  assign n13175 = ~po54  & n13173;
  assign n13176 = ~n12684 & ~n12685;
  assign n13177 = po11  & n13176;
  assign n13178 = ~n12690 & ~n13177;
  assign n13179 = n12690 & n13177;
  assign n13180 = ~n13178 & ~n13179;
  assign n13181 = ~n13175 & ~n13180;
  assign n13182 = ~n13174 & ~n13181;
  assign n13183 = po55  & ~n13182;
  assign n13184 = ~po55  & n13182;
  assign n13185 = ~n12693 & ~n12694;
  assign n13186 = po11  & n13185;
  assign n13187 = ~n12699 & ~n13186;
  assign n13188 = n12699 & n13186;
  assign n13189 = ~n13187 & ~n13188;
  assign n13190 = ~n13184 & ~n13189;
  assign n13191 = ~n13183 & ~n13190;
  assign n13192 = po56  & ~n13191;
  assign n13193 = ~po56  & n13191;
  assign n13194 = ~n12702 & ~n12703;
  assign n13195 = po11  & n13194;
  assign n13196 = ~n12708 & ~n13195;
  assign n13197 = n12708 & n13195;
  assign n13198 = ~n13196 & ~n13197;
  assign n13199 = ~n13193 & ~n13198;
  assign n13200 = ~n13192 & ~n13199;
  assign n13201 = po57  & ~n13200;
  assign n13202 = ~po57  & n13200;
  assign n13203 = ~n12711 & ~n12712;
  assign n13204 = po11  & n13203;
  assign n13205 = ~n12717 & ~n13204;
  assign n13206 = n12717 & n13204;
  assign n13207 = ~n13205 & ~n13206;
  assign n13208 = ~n13202 & ~n13207;
  assign n13209 = ~n13201 & ~n13208;
  assign n13210 = po58  & ~n13209;
  assign n13211 = ~po58  & n13209;
  assign n13212 = ~n12720 & ~n12721;
  assign n13213 = po11  & n13212;
  assign n13214 = ~n12726 & ~n13213;
  assign n13215 = n12726 & n13213;
  assign n13216 = ~n13214 & ~n13215;
  assign n13217 = ~n13211 & ~n13216;
  assign n13218 = ~n13210 & ~n13217;
  assign n13219 = po59  & ~n13218;
  assign n13220 = ~po59  & n13218;
  assign n13221 = ~n12729 & ~n12730;
  assign n13222 = po11  & n13221;
  assign n13223 = ~n12735 & ~n13222;
  assign n13224 = n12735 & n13222;
  assign n13225 = ~n13223 & ~n13224;
  assign n13226 = ~n13220 & ~n13225;
  assign n13227 = ~n13219 & ~n13226;
  assign n13228 = po60  & ~n13227;
  assign n13229 = ~po60  & n13227;
  assign n13230 = ~n12738 & ~n12739;
  assign n13231 = po11  & n13230;
  assign n13232 = ~n12744 & ~n13231;
  assign n13233 = n12744 & n13231;
  assign n13234 = ~n13232 & ~n13233;
  assign n13235 = ~n13229 & ~n13234;
  assign n13236 = ~n13228 & ~n13235;
  assign n13237 = po61  & ~n13236;
  assign n13238 = ~po61  & n13236;
  assign n13239 = ~n12747 & ~n12748;
  assign n13240 = po11  & n13239;
  assign n13241 = ~n12753 & ~n13240;
  assign n13242 = n12753 & n13240;
  assign n13243 = ~n13241 & ~n13242;
  assign n13244 = ~n13238 & ~n13243;
  assign n13245 = ~n13237 & ~n13244;
  assign n13246 = po62  & ~n13245;
  assign n13247 = ~po62  & n13245;
  assign n13248 = ~n12756 & ~n12757;
  assign n13249 = po11  & n13248;
  assign n13250 = ~n12762 & ~n13249;
  assign n13251 = n12762 & n13249;
  assign n13252 = ~n13250 & ~n13251;
  assign n13253 = ~n13247 & ~n13252;
  assign n13254 = ~n13246 & ~n13253;
  assign n13255 = n13171 & n13254;
  assign n13256 = ~n13171 & ~n13254;
  assign n13257 = n12775 & po11 ;
  assign n13258 = ~n12774 & ~n13257;
  assign n13259 = n13256 & n13258;
  assign n13260 = ~po63  & ~n13259;
  assign n13261 = ~n12681 & po11 ;
  assign n13262 = n12773 & ~n13261;
  assign n13263 = po63  & ~n12775;
  assign n13264 = ~n13262 & n13263;
  assign n13265 = ~n13255 & ~n13264;
  assign n13266 = ~n13260 & n13265;
  assign po10  = n13166 | ~n13266;
  assign n13268 = ~n13164 & ~n13165;
  assign n13269 = po10  & n13268;
  assign n13270 = ~n12791 & ~n13269;
  assign n13271 = n12791 & n13269;
  assign n13272 = ~n13270 & ~n13271;
  assign n13273 = pi20  & po10 ;
  assign n13274 = ~pi18  & ~pi19 ;
  assign n13275 = ~pi20  & n13274;
  assign n13276 = ~n13273 & ~n13275;
  assign n13277 = po11  & ~n13276;
  assign n13278 = ~po11  & n13276;
  assign n13279 = ~pi20  & po10 ;
  assign n13280 = pi21  & ~n13279;
  assign n13281 = ~pi21  & n13279;
  assign n13282 = ~n13280 & ~n13281;
  assign n13283 = ~n13278 & n13282;
  assign n13284 = ~n13277 & ~n13283;
  assign n13285 = po12  & ~n13284;
  assign n13286 = ~po12  & n13284;
  assign n13287 = po11  & n13266;
  assign n13288 = ~n13281 & ~n13287;
  assign n13289 = pi22  & ~n13288;
  assign n13290 = ~pi22  & n13288;
  assign n13291 = ~n13289 & ~n13290;
  assign n13292 = ~n13286 & ~n13291;
  assign n13293 = ~n13285 & ~n13292;
  assign n13294 = po13  & ~n13293;
  assign n13295 = ~po13  & n13293;
  assign n13296 = ~n12796 & ~n12797;
  assign n13297 = po10  & n13296;
  assign n13298 = n12801 & ~n13297;
  assign n13299 = ~n12801 & n13297;
  assign n13300 = ~n13298 & ~n13299;
  assign n13301 = ~n13295 & ~n13300;
  assign n13302 = ~n13294 & ~n13301;
  assign n13303 = po14  & ~n13302;
  assign n13304 = ~po14  & n13302;
  assign n13305 = ~n12804 & ~n12805;
  assign n13306 = po10  & n13305;
  assign n13307 = ~n12810 & ~n13306;
  assign n13308 = n12810 & n13306;
  assign n13309 = ~n13307 & ~n13308;
  assign n13310 = ~n13304 & ~n13309;
  assign n13311 = ~n13303 & ~n13310;
  assign n13312 = po15  & ~n13311;
  assign n13313 = ~po15  & n13311;
  assign n13314 = ~n12813 & ~n12814;
  assign n13315 = po10  & n13314;
  assign n13316 = n12819 & n13315;
  assign n13317 = ~n12819 & ~n13315;
  assign n13318 = ~n13316 & ~n13317;
  assign n13319 = ~n13313 & ~n13318;
  assign n13320 = ~n13312 & ~n13319;
  assign n13321 = po16  & ~n13320;
  assign n13322 = ~po16  & n13320;
  assign n13323 = ~n12822 & ~n12823;
  assign n13324 = po10  & n13323;
  assign n13325 = ~n12828 & ~n13324;
  assign n13326 = n12828 & n13324;
  assign n13327 = ~n13325 & ~n13326;
  assign n13328 = ~n13322 & ~n13327;
  assign n13329 = ~n13321 & ~n13328;
  assign n13330 = po17  & ~n13329;
  assign n13331 = ~po17  & n13329;
  assign n13332 = ~n12831 & ~n12832;
  assign n13333 = po10  & n13332;
  assign n13334 = ~n12837 & ~n13333;
  assign n13335 = n12837 & n13333;
  assign n13336 = ~n13334 & ~n13335;
  assign n13337 = ~n13331 & ~n13336;
  assign n13338 = ~n13330 & ~n13337;
  assign n13339 = po18  & ~n13338;
  assign n13340 = ~po18  & n13338;
  assign n13341 = ~n12840 & ~n12841;
  assign n13342 = po10  & n13341;
  assign n13343 = ~n12846 & ~n13342;
  assign n13344 = n12846 & n13342;
  assign n13345 = ~n13343 & ~n13344;
  assign n13346 = ~n13340 & ~n13345;
  assign n13347 = ~n13339 & ~n13346;
  assign n13348 = po19  & ~n13347;
  assign n13349 = ~po19  & n13347;
  assign n13350 = ~n12849 & ~n12850;
  assign n13351 = po10  & n13350;
  assign n13352 = ~n12855 & ~n13351;
  assign n13353 = n12855 & n13351;
  assign n13354 = ~n13352 & ~n13353;
  assign n13355 = ~n13349 & ~n13354;
  assign n13356 = ~n13348 & ~n13355;
  assign n13357 = po20  & ~n13356;
  assign n13358 = ~po20  & n13356;
  assign n13359 = ~n12858 & ~n12859;
  assign n13360 = po10  & n13359;
  assign n13361 = ~n12864 & ~n13360;
  assign n13362 = n12864 & n13360;
  assign n13363 = ~n13361 & ~n13362;
  assign n13364 = ~n13358 & ~n13363;
  assign n13365 = ~n13357 & ~n13364;
  assign n13366 = po21  & ~n13365;
  assign n13367 = ~po21  & n13365;
  assign n13368 = ~n12867 & ~n12868;
  assign n13369 = po10  & n13368;
  assign n13370 = ~n12873 & ~n13369;
  assign n13371 = n12873 & n13369;
  assign n13372 = ~n13370 & ~n13371;
  assign n13373 = ~n13367 & ~n13372;
  assign n13374 = ~n13366 & ~n13373;
  assign n13375 = po22  & ~n13374;
  assign n13376 = ~po22  & n13374;
  assign n13377 = ~n12876 & ~n12877;
  assign n13378 = po10  & n13377;
  assign n13379 = ~n12882 & ~n13378;
  assign n13380 = n12882 & n13378;
  assign n13381 = ~n13379 & ~n13380;
  assign n13382 = ~n13376 & ~n13381;
  assign n13383 = ~n13375 & ~n13382;
  assign n13384 = po23  & ~n13383;
  assign n13385 = ~po23  & n13383;
  assign n13386 = ~n12885 & ~n12886;
  assign n13387 = po10  & n13386;
  assign n13388 = ~n12891 & ~n13387;
  assign n13389 = n12891 & n13387;
  assign n13390 = ~n13388 & ~n13389;
  assign n13391 = ~n13385 & ~n13390;
  assign n13392 = ~n13384 & ~n13391;
  assign n13393 = po24  & ~n13392;
  assign n13394 = ~po24  & n13392;
  assign n13395 = ~n12894 & ~n12895;
  assign n13396 = po10  & n13395;
  assign n13397 = ~n12900 & ~n13396;
  assign n13398 = n12900 & n13396;
  assign n13399 = ~n13397 & ~n13398;
  assign n13400 = ~n13394 & ~n13399;
  assign n13401 = ~n13393 & ~n13400;
  assign n13402 = po25  & ~n13401;
  assign n13403 = ~po25  & n13401;
  assign n13404 = ~n12903 & ~n12904;
  assign n13405 = po10  & n13404;
  assign n13406 = ~n12909 & ~n13405;
  assign n13407 = n12909 & n13405;
  assign n13408 = ~n13406 & ~n13407;
  assign n13409 = ~n13403 & ~n13408;
  assign n13410 = ~n13402 & ~n13409;
  assign n13411 = po26  & ~n13410;
  assign n13412 = ~po26  & n13410;
  assign n13413 = ~n12912 & ~n12913;
  assign n13414 = po10  & n13413;
  assign n13415 = ~n12918 & ~n13414;
  assign n13416 = n12918 & n13414;
  assign n13417 = ~n13415 & ~n13416;
  assign n13418 = ~n13412 & ~n13417;
  assign n13419 = ~n13411 & ~n13418;
  assign n13420 = po27  & ~n13419;
  assign n13421 = ~po27  & n13419;
  assign n13422 = ~n12921 & ~n12922;
  assign n13423 = po10  & n13422;
  assign n13424 = ~n12927 & ~n13423;
  assign n13425 = n12927 & n13423;
  assign n13426 = ~n13424 & ~n13425;
  assign n13427 = ~n13421 & ~n13426;
  assign n13428 = ~n13420 & ~n13427;
  assign n13429 = po28  & ~n13428;
  assign n13430 = ~po28  & n13428;
  assign n13431 = ~n12930 & ~n12931;
  assign n13432 = po10  & n13431;
  assign n13433 = ~n12936 & ~n13432;
  assign n13434 = n12936 & n13432;
  assign n13435 = ~n13433 & ~n13434;
  assign n13436 = ~n13430 & ~n13435;
  assign n13437 = ~n13429 & ~n13436;
  assign n13438 = po29  & ~n13437;
  assign n13439 = ~po29  & n13437;
  assign n13440 = ~n12939 & ~n12940;
  assign n13441 = po10  & n13440;
  assign n13442 = ~n12945 & ~n13441;
  assign n13443 = n12945 & n13441;
  assign n13444 = ~n13442 & ~n13443;
  assign n13445 = ~n13439 & ~n13444;
  assign n13446 = ~n13438 & ~n13445;
  assign n13447 = po30  & ~n13446;
  assign n13448 = ~po30  & n13446;
  assign n13449 = ~n12948 & ~n12949;
  assign n13450 = po10  & n13449;
  assign n13451 = ~n12954 & ~n13450;
  assign n13452 = n12954 & n13450;
  assign n13453 = ~n13451 & ~n13452;
  assign n13454 = ~n13448 & ~n13453;
  assign n13455 = ~n13447 & ~n13454;
  assign n13456 = po31  & ~n13455;
  assign n13457 = ~po31  & n13455;
  assign n13458 = ~n12957 & ~n12958;
  assign n13459 = po10  & n13458;
  assign n13460 = ~n12963 & ~n13459;
  assign n13461 = n12963 & n13459;
  assign n13462 = ~n13460 & ~n13461;
  assign n13463 = ~n13457 & ~n13462;
  assign n13464 = ~n13456 & ~n13463;
  assign n13465 = po32  & ~n13464;
  assign n13466 = ~po32  & n13464;
  assign n13467 = ~n12966 & ~n12967;
  assign n13468 = po10  & n13467;
  assign n13469 = ~n12972 & ~n13468;
  assign n13470 = n12972 & n13468;
  assign n13471 = ~n13469 & ~n13470;
  assign n13472 = ~n13466 & ~n13471;
  assign n13473 = ~n13465 & ~n13472;
  assign n13474 = po33  & ~n13473;
  assign n13475 = ~po33  & n13473;
  assign n13476 = ~n12975 & ~n12976;
  assign n13477 = po10  & n13476;
  assign n13478 = ~n12981 & ~n13477;
  assign n13479 = n12981 & n13477;
  assign n13480 = ~n13478 & ~n13479;
  assign n13481 = ~n13475 & ~n13480;
  assign n13482 = ~n13474 & ~n13481;
  assign n13483 = po34  & ~n13482;
  assign n13484 = ~po34  & n13482;
  assign n13485 = ~n12984 & ~n12985;
  assign n13486 = po10  & n13485;
  assign n13487 = ~n12990 & ~n13486;
  assign n13488 = n12990 & n13486;
  assign n13489 = ~n13487 & ~n13488;
  assign n13490 = ~n13484 & ~n13489;
  assign n13491 = ~n13483 & ~n13490;
  assign n13492 = po35  & ~n13491;
  assign n13493 = ~po35  & n13491;
  assign n13494 = ~n12993 & ~n12994;
  assign n13495 = po10  & n13494;
  assign n13496 = ~n12999 & ~n13495;
  assign n13497 = n12999 & n13495;
  assign n13498 = ~n13496 & ~n13497;
  assign n13499 = ~n13493 & ~n13498;
  assign n13500 = ~n13492 & ~n13499;
  assign n13501 = po36  & ~n13500;
  assign n13502 = ~po36  & n13500;
  assign n13503 = ~n13002 & ~n13003;
  assign n13504 = po10  & n13503;
  assign n13505 = ~n13008 & ~n13504;
  assign n13506 = n13008 & n13504;
  assign n13507 = ~n13505 & ~n13506;
  assign n13508 = ~n13502 & ~n13507;
  assign n13509 = ~n13501 & ~n13508;
  assign n13510 = po37  & ~n13509;
  assign n13511 = ~po37  & n13509;
  assign n13512 = ~n13011 & ~n13012;
  assign n13513 = po10  & n13512;
  assign n13514 = ~n13017 & ~n13513;
  assign n13515 = n13017 & n13513;
  assign n13516 = ~n13514 & ~n13515;
  assign n13517 = ~n13511 & ~n13516;
  assign n13518 = ~n13510 & ~n13517;
  assign n13519 = po38  & ~n13518;
  assign n13520 = ~po38  & n13518;
  assign n13521 = ~n13020 & ~n13021;
  assign n13522 = po10  & n13521;
  assign n13523 = ~n13026 & ~n13522;
  assign n13524 = n13026 & n13522;
  assign n13525 = ~n13523 & ~n13524;
  assign n13526 = ~n13520 & ~n13525;
  assign n13527 = ~n13519 & ~n13526;
  assign n13528 = po39  & ~n13527;
  assign n13529 = ~po39  & n13527;
  assign n13530 = ~n13029 & ~n13030;
  assign n13531 = po10  & n13530;
  assign n13532 = ~n13035 & ~n13531;
  assign n13533 = n13035 & n13531;
  assign n13534 = ~n13532 & ~n13533;
  assign n13535 = ~n13529 & ~n13534;
  assign n13536 = ~n13528 & ~n13535;
  assign n13537 = po40  & ~n13536;
  assign n13538 = ~po40  & n13536;
  assign n13539 = ~n13038 & ~n13039;
  assign n13540 = po10  & n13539;
  assign n13541 = ~n13044 & ~n13540;
  assign n13542 = n13044 & n13540;
  assign n13543 = ~n13541 & ~n13542;
  assign n13544 = ~n13538 & ~n13543;
  assign n13545 = ~n13537 & ~n13544;
  assign n13546 = po41  & ~n13545;
  assign n13547 = ~po41  & n13545;
  assign n13548 = ~n13047 & ~n13048;
  assign n13549 = po10  & n13548;
  assign n13550 = ~n13053 & ~n13549;
  assign n13551 = n13053 & n13549;
  assign n13552 = ~n13550 & ~n13551;
  assign n13553 = ~n13547 & ~n13552;
  assign n13554 = ~n13546 & ~n13553;
  assign n13555 = po42  & ~n13554;
  assign n13556 = ~po42  & n13554;
  assign n13557 = ~n13056 & ~n13057;
  assign n13558 = po10  & n13557;
  assign n13559 = ~n13062 & ~n13558;
  assign n13560 = n13062 & n13558;
  assign n13561 = ~n13559 & ~n13560;
  assign n13562 = ~n13556 & ~n13561;
  assign n13563 = ~n13555 & ~n13562;
  assign n13564 = po43  & ~n13563;
  assign n13565 = ~po43  & n13563;
  assign n13566 = ~n13065 & ~n13066;
  assign n13567 = po10  & n13566;
  assign n13568 = ~n13071 & ~n13567;
  assign n13569 = n13071 & n13567;
  assign n13570 = ~n13568 & ~n13569;
  assign n13571 = ~n13565 & ~n13570;
  assign n13572 = ~n13564 & ~n13571;
  assign n13573 = po44  & ~n13572;
  assign n13574 = ~po44  & n13572;
  assign n13575 = ~n13074 & ~n13075;
  assign n13576 = po10  & n13575;
  assign n13577 = ~n13080 & ~n13576;
  assign n13578 = n13080 & n13576;
  assign n13579 = ~n13577 & ~n13578;
  assign n13580 = ~n13574 & ~n13579;
  assign n13581 = ~n13573 & ~n13580;
  assign n13582 = po45  & ~n13581;
  assign n13583 = ~po45  & n13581;
  assign n13584 = ~n13083 & ~n13084;
  assign n13585 = po10  & n13584;
  assign n13586 = ~n13089 & ~n13585;
  assign n13587 = n13089 & n13585;
  assign n13588 = ~n13586 & ~n13587;
  assign n13589 = ~n13583 & ~n13588;
  assign n13590 = ~n13582 & ~n13589;
  assign n13591 = po46  & ~n13590;
  assign n13592 = ~po46  & n13590;
  assign n13593 = ~n13092 & ~n13093;
  assign n13594 = po10  & n13593;
  assign n13595 = ~n13098 & ~n13594;
  assign n13596 = n13098 & n13594;
  assign n13597 = ~n13595 & ~n13596;
  assign n13598 = ~n13592 & ~n13597;
  assign n13599 = ~n13591 & ~n13598;
  assign n13600 = po47  & ~n13599;
  assign n13601 = ~po47  & n13599;
  assign n13602 = ~n13101 & ~n13102;
  assign n13603 = po10  & n13602;
  assign n13604 = ~n13107 & ~n13603;
  assign n13605 = n13107 & n13603;
  assign n13606 = ~n13604 & ~n13605;
  assign n13607 = ~n13601 & ~n13606;
  assign n13608 = ~n13600 & ~n13607;
  assign n13609 = po48  & ~n13608;
  assign n13610 = ~po48  & n13608;
  assign n13611 = ~n13110 & ~n13111;
  assign n13612 = po10  & n13611;
  assign n13613 = ~n13116 & ~n13612;
  assign n13614 = n13116 & n13612;
  assign n13615 = ~n13613 & ~n13614;
  assign n13616 = ~n13610 & ~n13615;
  assign n13617 = ~n13609 & ~n13616;
  assign n13618 = po49  & ~n13617;
  assign n13619 = ~po49  & n13617;
  assign n13620 = ~n13119 & ~n13120;
  assign n13621 = po10  & n13620;
  assign n13622 = ~n13125 & ~n13621;
  assign n13623 = n13125 & n13621;
  assign n13624 = ~n13622 & ~n13623;
  assign n13625 = ~n13619 & ~n13624;
  assign n13626 = ~n13618 & ~n13625;
  assign n13627 = po50  & ~n13626;
  assign n13628 = ~po50  & n13626;
  assign n13629 = ~n13128 & ~n13129;
  assign n13630 = po10  & n13629;
  assign n13631 = ~n13134 & ~n13630;
  assign n13632 = n13134 & n13630;
  assign n13633 = ~n13631 & ~n13632;
  assign n13634 = ~n13628 & ~n13633;
  assign n13635 = ~n13627 & ~n13634;
  assign n13636 = po51  & ~n13635;
  assign n13637 = ~po51  & n13635;
  assign n13638 = ~n13137 & ~n13138;
  assign n13639 = po10  & n13638;
  assign n13640 = ~n13143 & ~n13639;
  assign n13641 = n13143 & n13639;
  assign n13642 = ~n13640 & ~n13641;
  assign n13643 = ~n13637 & ~n13642;
  assign n13644 = ~n13636 & ~n13643;
  assign n13645 = po52  & ~n13644;
  assign n13646 = ~po52  & n13644;
  assign n13647 = ~n13146 & ~n13147;
  assign n13648 = po10  & n13647;
  assign n13649 = ~n13152 & ~n13648;
  assign n13650 = n13152 & n13648;
  assign n13651 = ~n13649 & ~n13650;
  assign n13652 = ~n13646 & ~n13651;
  assign n13653 = ~n13645 & ~n13652;
  assign n13654 = po53  & ~n13653;
  assign n13655 = ~n13155 & ~n13161;
  assign n13656 = po10  & n13655;
  assign n13657 = ~n13160 & ~n13656;
  assign n13658 = n13160 & n13656;
  assign n13659 = ~n13657 & ~n13658;
  assign n13660 = ~po53  & n13653;
  assign n13661 = ~n13659 & ~n13660;
  assign n13662 = ~n13654 & ~n13661;
  assign n13663 = po54  & ~n13662;
  assign n13664 = ~po54  & n13662;
  assign n13665 = n13171 & ~po10 ;
  assign n13666 = ~n13246 & ~n13247;
  assign n13667 = po10  & n13666;
  assign n13668 = ~n13252 & ~n13667;
  assign n13669 = n13252 & n13667;
  assign n13670 = ~n13668 & ~n13669;
  assign n13671 = ~n13272 & ~n13664;
  assign n13672 = ~n13663 & ~n13671;
  assign n13673 = po55  & ~n13672;
  assign n13674 = ~po55  & n13672;
  assign n13675 = ~n13174 & ~n13175;
  assign n13676 = po10  & n13675;
  assign n13677 = ~n13180 & ~n13676;
  assign n13678 = n13180 & n13676;
  assign n13679 = ~n13677 & ~n13678;
  assign n13680 = ~n13674 & ~n13679;
  assign n13681 = ~n13673 & ~n13680;
  assign n13682 = po56  & ~n13681;
  assign n13683 = ~po56  & n13681;
  assign n13684 = ~n13183 & ~n13184;
  assign n13685 = po10  & n13684;
  assign n13686 = ~n13189 & ~n13685;
  assign n13687 = n13189 & n13685;
  assign n13688 = ~n13686 & ~n13687;
  assign n13689 = ~n13683 & ~n13688;
  assign n13690 = ~n13682 & ~n13689;
  assign n13691 = po57  & ~n13690;
  assign n13692 = ~po57  & n13690;
  assign n13693 = ~n13192 & ~n13193;
  assign n13694 = po10  & n13693;
  assign n13695 = ~n13198 & ~n13694;
  assign n13696 = n13198 & n13694;
  assign n13697 = ~n13695 & ~n13696;
  assign n13698 = ~n13692 & ~n13697;
  assign n13699 = ~n13691 & ~n13698;
  assign n13700 = po58  & ~n13699;
  assign n13701 = ~po58  & n13699;
  assign n13702 = ~n13201 & ~n13202;
  assign n13703 = po10  & n13702;
  assign n13704 = ~n13207 & ~n13703;
  assign n13705 = n13207 & n13703;
  assign n13706 = ~n13704 & ~n13705;
  assign n13707 = ~n13701 & ~n13706;
  assign n13708 = ~n13700 & ~n13707;
  assign n13709 = po59  & ~n13708;
  assign n13710 = ~po59  & n13708;
  assign n13711 = ~n13210 & ~n13211;
  assign n13712 = po10  & n13711;
  assign n13713 = ~n13216 & ~n13712;
  assign n13714 = n13216 & n13712;
  assign n13715 = ~n13713 & ~n13714;
  assign n13716 = ~n13710 & ~n13715;
  assign n13717 = ~n13709 & ~n13716;
  assign n13718 = po60  & ~n13717;
  assign n13719 = ~po60  & n13717;
  assign n13720 = ~n13219 & ~n13220;
  assign n13721 = po10  & n13720;
  assign n13722 = ~n13225 & ~n13721;
  assign n13723 = n13225 & n13721;
  assign n13724 = ~n13722 & ~n13723;
  assign n13725 = ~n13719 & ~n13724;
  assign n13726 = ~n13718 & ~n13725;
  assign n13727 = po61  & ~n13726;
  assign n13728 = ~po61  & n13726;
  assign n13729 = ~n13228 & ~n13229;
  assign n13730 = po10  & n13729;
  assign n13731 = ~n13234 & ~n13730;
  assign n13732 = n13234 & n13730;
  assign n13733 = ~n13731 & ~n13732;
  assign n13734 = ~n13728 & ~n13733;
  assign n13735 = ~n13727 & ~n13734;
  assign n13736 = po62  & ~n13735;
  assign n13737 = ~po62  & n13735;
  assign n13738 = ~n13237 & ~n13238;
  assign n13739 = po10  & n13738;
  assign n13740 = ~n13243 & ~n13739;
  assign n13741 = n13243 & n13739;
  assign n13742 = ~n13740 & ~n13741;
  assign n13743 = ~n13737 & ~n13742;
  assign n13744 = ~n13736 & ~n13743;
  assign n13745 = n13670 & n13744;
  assign n13746 = ~n13670 & ~n13744;
  assign n13747 = n13256 & po10 ;
  assign n13748 = ~n13255 & ~n13747;
  assign n13749 = n13746 & n13748;
  assign n13750 = ~po63  & ~n13749;
  assign n13751 = ~n13171 & po10 ;
  assign n13752 = n13254 & ~n13751;
  assign n13753 = po63  & ~n13256;
  assign n13754 = ~n13752 & n13753;
  assign n13755 = ~n13745 & ~n13754;
  assign n13756 = ~n13750 & n13755;
  assign po9  = n13665 | ~n13756;
  assign n13758 = ~n13663 & ~n13664;
  assign n13759 = po9  & n13758;
  assign n13760 = ~n13272 & ~n13759;
  assign n13761 = n13272 & n13759;
  assign n13762 = ~n13760 & ~n13761;
  assign n13763 = pi18  & po9 ;
  assign n13764 = ~pi16  & ~pi17 ;
  assign n13765 = ~pi18  & n13764;
  assign n13766 = ~n13763 & ~n13765;
  assign n13767 = po10  & ~n13766;
  assign n13768 = ~po10  & n13766;
  assign n13769 = ~pi18  & po9 ;
  assign n13770 = pi19  & ~n13769;
  assign n13771 = ~pi19  & n13769;
  assign n13772 = ~n13770 & ~n13771;
  assign n13773 = ~n13768 & n13772;
  assign n13774 = ~n13767 & ~n13773;
  assign n13775 = po11  & ~n13774;
  assign n13776 = ~po11  & n13774;
  assign n13777 = po10  & n13756;
  assign n13778 = ~n13771 & ~n13777;
  assign n13779 = pi20  & ~n13778;
  assign n13780 = ~pi20  & n13778;
  assign n13781 = ~n13779 & ~n13780;
  assign n13782 = ~n13776 & ~n13781;
  assign n13783 = ~n13775 & ~n13782;
  assign n13784 = po12  & ~n13783;
  assign n13785 = ~po12  & n13783;
  assign n13786 = ~n13277 & ~n13278;
  assign n13787 = po9  & n13786;
  assign n13788 = n13282 & ~n13787;
  assign n13789 = ~n13282 & n13787;
  assign n13790 = ~n13788 & ~n13789;
  assign n13791 = ~n13785 & ~n13790;
  assign n13792 = ~n13784 & ~n13791;
  assign n13793 = po13  & ~n13792;
  assign n13794 = ~po13  & n13792;
  assign n13795 = ~n13285 & ~n13286;
  assign n13796 = po9  & n13795;
  assign n13797 = ~n13291 & ~n13796;
  assign n13798 = n13291 & n13796;
  assign n13799 = ~n13797 & ~n13798;
  assign n13800 = ~n13794 & ~n13799;
  assign n13801 = ~n13793 & ~n13800;
  assign n13802 = po14  & ~n13801;
  assign n13803 = ~po14  & n13801;
  assign n13804 = ~n13294 & ~n13295;
  assign n13805 = po9  & n13804;
  assign n13806 = n13300 & n13805;
  assign n13807 = ~n13300 & ~n13805;
  assign n13808 = ~n13806 & ~n13807;
  assign n13809 = ~n13803 & ~n13808;
  assign n13810 = ~n13802 & ~n13809;
  assign n13811 = po15  & ~n13810;
  assign n13812 = ~po15  & n13810;
  assign n13813 = ~n13303 & ~n13304;
  assign n13814 = po9  & n13813;
  assign n13815 = ~n13309 & ~n13814;
  assign n13816 = n13309 & n13814;
  assign n13817 = ~n13815 & ~n13816;
  assign n13818 = ~n13812 & ~n13817;
  assign n13819 = ~n13811 & ~n13818;
  assign n13820 = po16  & ~n13819;
  assign n13821 = ~po16  & n13819;
  assign n13822 = ~n13312 & ~n13313;
  assign n13823 = po9  & n13822;
  assign n13824 = ~n13318 & ~n13823;
  assign n13825 = n13318 & n13823;
  assign n13826 = ~n13824 & ~n13825;
  assign n13827 = ~n13821 & ~n13826;
  assign n13828 = ~n13820 & ~n13827;
  assign n13829 = po17  & ~n13828;
  assign n13830 = ~po17  & n13828;
  assign n13831 = ~n13321 & ~n13322;
  assign n13832 = po9  & n13831;
  assign n13833 = ~n13327 & ~n13832;
  assign n13834 = n13327 & n13832;
  assign n13835 = ~n13833 & ~n13834;
  assign n13836 = ~n13830 & ~n13835;
  assign n13837 = ~n13829 & ~n13836;
  assign n13838 = po18  & ~n13837;
  assign n13839 = ~po18  & n13837;
  assign n13840 = ~n13330 & ~n13331;
  assign n13841 = po9  & n13840;
  assign n13842 = ~n13336 & ~n13841;
  assign n13843 = n13336 & n13841;
  assign n13844 = ~n13842 & ~n13843;
  assign n13845 = ~n13839 & ~n13844;
  assign n13846 = ~n13838 & ~n13845;
  assign n13847 = po19  & ~n13846;
  assign n13848 = ~po19  & n13846;
  assign n13849 = ~n13339 & ~n13340;
  assign n13850 = po9  & n13849;
  assign n13851 = ~n13345 & ~n13850;
  assign n13852 = n13345 & n13850;
  assign n13853 = ~n13851 & ~n13852;
  assign n13854 = ~n13848 & ~n13853;
  assign n13855 = ~n13847 & ~n13854;
  assign n13856 = po20  & ~n13855;
  assign n13857 = ~po20  & n13855;
  assign n13858 = ~n13348 & ~n13349;
  assign n13859 = po9  & n13858;
  assign n13860 = ~n13354 & ~n13859;
  assign n13861 = n13354 & n13859;
  assign n13862 = ~n13860 & ~n13861;
  assign n13863 = ~n13857 & ~n13862;
  assign n13864 = ~n13856 & ~n13863;
  assign n13865 = po21  & ~n13864;
  assign n13866 = ~po21  & n13864;
  assign n13867 = ~n13357 & ~n13358;
  assign n13868 = po9  & n13867;
  assign n13869 = ~n13363 & ~n13868;
  assign n13870 = n13363 & n13868;
  assign n13871 = ~n13869 & ~n13870;
  assign n13872 = ~n13866 & ~n13871;
  assign n13873 = ~n13865 & ~n13872;
  assign n13874 = po22  & ~n13873;
  assign n13875 = ~po22  & n13873;
  assign n13876 = ~n13366 & ~n13367;
  assign n13877 = po9  & n13876;
  assign n13878 = ~n13372 & ~n13877;
  assign n13879 = n13372 & n13877;
  assign n13880 = ~n13878 & ~n13879;
  assign n13881 = ~n13875 & ~n13880;
  assign n13882 = ~n13874 & ~n13881;
  assign n13883 = po23  & ~n13882;
  assign n13884 = ~po23  & n13882;
  assign n13885 = ~n13375 & ~n13376;
  assign n13886 = po9  & n13885;
  assign n13887 = ~n13381 & ~n13886;
  assign n13888 = n13381 & n13886;
  assign n13889 = ~n13887 & ~n13888;
  assign n13890 = ~n13884 & ~n13889;
  assign n13891 = ~n13883 & ~n13890;
  assign n13892 = po24  & ~n13891;
  assign n13893 = ~po24  & n13891;
  assign n13894 = ~n13384 & ~n13385;
  assign n13895 = po9  & n13894;
  assign n13896 = ~n13390 & ~n13895;
  assign n13897 = n13390 & n13895;
  assign n13898 = ~n13896 & ~n13897;
  assign n13899 = ~n13893 & ~n13898;
  assign n13900 = ~n13892 & ~n13899;
  assign n13901 = po25  & ~n13900;
  assign n13902 = ~po25  & n13900;
  assign n13903 = ~n13393 & ~n13394;
  assign n13904 = po9  & n13903;
  assign n13905 = ~n13399 & ~n13904;
  assign n13906 = n13399 & n13904;
  assign n13907 = ~n13905 & ~n13906;
  assign n13908 = ~n13902 & ~n13907;
  assign n13909 = ~n13901 & ~n13908;
  assign n13910 = po26  & ~n13909;
  assign n13911 = ~po26  & n13909;
  assign n13912 = ~n13402 & ~n13403;
  assign n13913 = po9  & n13912;
  assign n13914 = ~n13408 & ~n13913;
  assign n13915 = n13408 & n13913;
  assign n13916 = ~n13914 & ~n13915;
  assign n13917 = ~n13911 & ~n13916;
  assign n13918 = ~n13910 & ~n13917;
  assign n13919 = po27  & ~n13918;
  assign n13920 = ~po27  & n13918;
  assign n13921 = ~n13411 & ~n13412;
  assign n13922 = po9  & n13921;
  assign n13923 = ~n13417 & ~n13922;
  assign n13924 = n13417 & n13922;
  assign n13925 = ~n13923 & ~n13924;
  assign n13926 = ~n13920 & ~n13925;
  assign n13927 = ~n13919 & ~n13926;
  assign n13928 = po28  & ~n13927;
  assign n13929 = ~po28  & n13927;
  assign n13930 = ~n13420 & ~n13421;
  assign n13931 = po9  & n13930;
  assign n13932 = ~n13426 & ~n13931;
  assign n13933 = n13426 & n13931;
  assign n13934 = ~n13932 & ~n13933;
  assign n13935 = ~n13929 & ~n13934;
  assign n13936 = ~n13928 & ~n13935;
  assign n13937 = po29  & ~n13936;
  assign n13938 = ~po29  & n13936;
  assign n13939 = ~n13429 & ~n13430;
  assign n13940 = po9  & n13939;
  assign n13941 = ~n13435 & ~n13940;
  assign n13942 = n13435 & n13940;
  assign n13943 = ~n13941 & ~n13942;
  assign n13944 = ~n13938 & ~n13943;
  assign n13945 = ~n13937 & ~n13944;
  assign n13946 = po30  & ~n13945;
  assign n13947 = ~po30  & n13945;
  assign n13948 = ~n13438 & ~n13439;
  assign n13949 = po9  & n13948;
  assign n13950 = ~n13444 & ~n13949;
  assign n13951 = n13444 & n13949;
  assign n13952 = ~n13950 & ~n13951;
  assign n13953 = ~n13947 & ~n13952;
  assign n13954 = ~n13946 & ~n13953;
  assign n13955 = po31  & ~n13954;
  assign n13956 = ~po31  & n13954;
  assign n13957 = ~n13447 & ~n13448;
  assign n13958 = po9  & n13957;
  assign n13959 = ~n13453 & ~n13958;
  assign n13960 = n13453 & n13958;
  assign n13961 = ~n13959 & ~n13960;
  assign n13962 = ~n13956 & ~n13961;
  assign n13963 = ~n13955 & ~n13962;
  assign n13964 = po32  & ~n13963;
  assign n13965 = ~po32  & n13963;
  assign n13966 = ~n13456 & ~n13457;
  assign n13967 = po9  & n13966;
  assign n13968 = ~n13462 & ~n13967;
  assign n13969 = n13462 & n13967;
  assign n13970 = ~n13968 & ~n13969;
  assign n13971 = ~n13965 & ~n13970;
  assign n13972 = ~n13964 & ~n13971;
  assign n13973 = po33  & ~n13972;
  assign n13974 = ~po33  & n13972;
  assign n13975 = ~n13465 & ~n13466;
  assign n13976 = po9  & n13975;
  assign n13977 = ~n13471 & ~n13976;
  assign n13978 = n13471 & n13976;
  assign n13979 = ~n13977 & ~n13978;
  assign n13980 = ~n13974 & ~n13979;
  assign n13981 = ~n13973 & ~n13980;
  assign n13982 = po34  & ~n13981;
  assign n13983 = ~po34  & n13981;
  assign n13984 = ~n13474 & ~n13475;
  assign n13985 = po9  & n13984;
  assign n13986 = ~n13480 & ~n13985;
  assign n13987 = n13480 & n13985;
  assign n13988 = ~n13986 & ~n13987;
  assign n13989 = ~n13983 & ~n13988;
  assign n13990 = ~n13982 & ~n13989;
  assign n13991 = po35  & ~n13990;
  assign n13992 = ~po35  & n13990;
  assign n13993 = ~n13483 & ~n13484;
  assign n13994 = po9  & n13993;
  assign n13995 = ~n13489 & ~n13994;
  assign n13996 = n13489 & n13994;
  assign n13997 = ~n13995 & ~n13996;
  assign n13998 = ~n13992 & ~n13997;
  assign n13999 = ~n13991 & ~n13998;
  assign n14000 = po36  & ~n13999;
  assign n14001 = ~po36  & n13999;
  assign n14002 = ~n13492 & ~n13493;
  assign n14003 = po9  & n14002;
  assign n14004 = ~n13498 & ~n14003;
  assign n14005 = n13498 & n14003;
  assign n14006 = ~n14004 & ~n14005;
  assign n14007 = ~n14001 & ~n14006;
  assign n14008 = ~n14000 & ~n14007;
  assign n14009 = po37  & ~n14008;
  assign n14010 = ~po37  & n14008;
  assign n14011 = ~n13501 & ~n13502;
  assign n14012 = po9  & n14011;
  assign n14013 = ~n13507 & ~n14012;
  assign n14014 = n13507 & n14012;
  assign n14015 = ~n14013 & ~n14014;
  assign n14016 = ~n14010 & ~n14015;
  assign n14017 = ~n14009 & ~n14016;
  assign n14018 = po38  & ~n14017;
  assign n14019 = ~po38  & n14017;
  assign n14020 = ~n13510 & ~n13511;
  assign n14021 = po9  & n14020;
  assign n14022 = ~n13516 & ~n14021;
  assign n14023 = n13516 & n14021;
  assign n14024 = ~n14022 & ~n14023;
  assign n14025 = ~n14019 & ~n14024;
  assign n14026 = ~n14018 & ~n14025;
  assign n14027 = po39  & ~n14026;
  assign n14028 = ~po39  & n14026;
  assign n14029 = ~n13519 & ~n13520;
  assign n14030 = po9  & n14029;
  assign n14031 = ~n13525 & ~n14030;
  assign n14032 = n13525 & n14030;
  assign n14033 = ~n14031 & ~n14032;
  assign n14034 = ~n14028 & ~n14033;
  assign n14035 = ~n14027 & ~n14034;
  assign n14036 = po40  & ~n14035;
  assign n14037 = ~po40  & n14035;
  assign n14038 = ~n13528 & ~n13529;
  assign n14039 = po9  & n14038;
  assign n14040 = ~n13534 & ~n14039;
  assign n14041 = n13534 & n14039;
  assign n14042 = ~n14040 & ~n14041;
  assign n14043 = ~n14037 & ~n14042;
  assign n14044 = ~n14036 & ~n14043;
  assign n14045 = po41  & ~n14044;
  assign n14046 = ~po41  & n14044;
  assign n14047 = ~n13537 & ~n13538;
  assign n14048 = po9  & n14047;
  assign n14049 = ~n13543 & ~n14048;
  assign n14050 = n13543 & n14048;
  assign n14051 = ~n14049 & ~n14050;
  assign n14052 = ~n14046 & ~n14051;
  assign n14053 = ~n14045 & ~n14052;
  assign n14054 = po42  & ~n14053;
  assign n14055 = ~po42  & n14053;
  assign n14056 = ~n13546 & ~n13547;
  assign n14057 = po9  & n14056;
  assign n14058 = ~n13552 & ~n14057;
  assign n14059 = n13552 & n14057;
  assign n14060 = ~n14058 & ~n14059;
  assign n14061 = ~n14055 & ~n14060;
  assign n14062 = ~n14054 & ~n14061;
  assign n14063 = po43  & ~n14062;
  assign n14064 = ~po43  & n14062;
  assign n14065 = ~n13555 & ~n13556;
  assign n14066 = po9  & n14065;
  assign n14067 = ~n13561 & ~n14066;
  assign n14068 = n13561 & n14066;
  assign n14069 = ~n14067 & ~n14068;
  assign n14070 = ~n14064 & ~n14069;
  assign n14071 = ~n14063 & ~n14070;
  assign n14072 = po44  & ~n14071;
  assign n14073 = ~po44  & n14071;
  assign n14074 = ~n13564 & ~n13565;
  assign n14075 = po9  & n14074;
  assign n14076 = ~n13570 & ~n14075;
  assign n14077 = n13570 & n14075;
  assign n14078 = ~n14076 & ~n14077;
  assign n14079 = ~n14073 & ~n14078;
  assign n14080 = ~n14072 & ~n14079;
  assign n14081 = po45  & ~n14080;
  assign n14082 = ~po45  & n14080;
  assign n14083 = ~n13573 & ~n13574;
  assign n14084 = po9  & n14083;
  assign n14085 = ~n13579 & ~n14084;
  assign n14086 = n13579 & n14084;
  assign n14087 = ~n14085 & ~n14086;
  assign n14088 = ~n14082 & ~n14087;
  assign n14089 = ~n14081 & ~n14088;
  assign n14090 = po46  & ~n14089;
  assign n14091 = ~po46  & n14089;
  assign n14092 = ~n13582 & ~n13583;
  assign n14093 = po9  & n14092;
  assign n14094 = ~n13588 & ~n14093;
  assign n14095 = n13588 & n14093;
  assign n14096 = ~n14094 & ~n14095;
  assign n14097 = ~n14091 & ~n14096;
  assign n14098 = ~n14090 & ~n14097;
  assign n14099 = po47  & ~n14098;
  assign n14100 = ~po47  & n14098;
  assign n14101 = ~n13591 & ~n13592;
  assign n14102 = po9  & n14101;
  assign n14103 = ~n13597 & ~n14102;
  assign n14104 = n13597 & n14102;
  assign n14105 = ~n14103 & ~n14104;
  assign n14106 = ~n14100 & ~n14105;
  assign n14107 = ~n14099 & ~n14106;
  assign n14108 = po48  & ~n14107;
  assign n14109 = ~po48  & n14107;
  assign n14110 = ~n13600 & ~n13601;
  assign n14111 = po9  & n14110;
  assign n14112 = ~n13606 & ~n14111;
  assign n14113 = n13606 & n14111;
  assign n14114 = ~n14112 & ~n14113;
  assign n14115 = ~n14109 & ~n14114;
  assign n14116 = ~n14108 & ~n14115;
  assign n14117 = po49  & ~n14116;
  assign n14118 = ~po49  & n14116;
  assign n14119 = ~n13609 & ~n13610;
  assign n14120 = po9  & n14119;
  assign n14121 = ~n13615 & ~n14120;
  assign n14122 = n13615 & n14120;
  assign n14123 = ~n14121 & ~n14122;
  assign n14124 = ~n14118 & ~n14123;
  assign n14125 = ~n14117 & ~n14124;
  assign n14126 = po50  & ~n14125;
  assign n14127 = ~po50  & n14125;
  assign n14128 = ~n13618 & ~n13619;
  assign n14129 = po9  & n14128;
  assign n14130 = ~n13624 & ~n14129;
  assign n14131 = n13624 & n14129;
  assign n14132 = ~n14130 & ~n14131;
  assign n14133 = ~n14127 & ~n14132;
  assign n14134 = ~n14126 & ~n14133;
  assign n14135 = po51  & ~n14134;
  assign n14136 = ~po51  & n14134;
  assign n14137 = ~n13627 & ~n13628;
  assign n14138 = po9  & n14137;
  assign n14139 = ~n13633 & ~n14138;
  assign n14140 = n13633 & n14138;
  assign n14141 = ~n14139 & ~n14140;
  assign n14142 = ~n14136 & ~n14141;
  assign n14143 = ~n14135 & ~n14142;
  assign n14144 = po52  & ~n14143;
  assign n14145 = ~po52  & n14143;
  assign n14146 = ~n13636 & ~n13637;
  assign n14147 = po9  & n14146;
  assign n14148 = ~n13642 & ~n14147;
  assign n14149 = n13642 & n14147;
  assign n14150 = ~n14148 & ~n14149;
  assign n14151 = ~n14145 & ~n14150;
  assign n14152 = ~n14144 & ~n14151;
  assign n14153 = po53  & ~n14152;
  assign n14154 = ~po53  & n14152;
  assign n14155 = ~n13645 & ~n13646;
  assign n14156 = po9  & n14155;
  assign n14157 = ~n13651 & ~n14156;
  assign n14158 = n13651 & n14156;
  assign n14159 = ~n14157 & ~n14158;
  assign n14160 = ~n14154 & ~n14159;
  assign n14161 = ~n14153 & ~n14160;
  assign n14162 = po54  & ~n14161;
  assign n14163 = ~n13654 & ~n13660;
  assign n14164 = po9  & n14163;
  assign n14165 = ~n13659 & ~n14164;
  assign n14166 = n13659 & n14164;
  assign n14167 = ~n14165 & ~n14166;
  assign n14168 = ~po54  & n14161;
  assign n14169 = ~n14167 & ~n14168;
  assign n14170 = ~n14162 & ~n14169;
  assign n14171 = po55  & ~n14170;
  assign n14172 = ~po55  & n14170;
  assign n14173 = n13670 & ~po9 ;
  assign n14174 = ~n13736 & ~n13737;
  assign n14175 = po9  & n14174;
  assign n14176 = ~n13742 & ~n14175;
  assign n14177 = n13742 & n14175;
  assign n14178 = ~n14176 & ~n14177;
  assign n14179 = ~n13762 & ~n14172;
  assign n14180 = ~n14171 & ~n14179;
  assign n14181 = po56  & ~n14180;
  assign n14182 = ~po56  & n14180;
  assign n14183 = ~n13673 & ~n13674;
  assign n14184 = po9  & n14183;
  assign n14185 = ~n13679 & ~n14184;
  assign n14186 = n13679 & n14184;
  assign n14187 = ~n14185 & ~n14186;
  assign n14188 = ~n14182 & ~n14187;
  assign n14189 = ~n14181 & ~n14188;
  assign n14190 = po57  & ~n14189;
  assign n14191 = ~po57  & n14189;
  assign n14192 = ~n13682 & ~n13683;
  assign n14193 = po9  & n14192;
  assign n14194 = ~n13688 & ~n14193;
  assign n14195 = n13688 & n14193;
  assign n14196 = ~n14194 & ~n14195;
  assign n14197 = ~n14191 & ~n14196;
  assign n14198 = ~n14190 & ~n14197;
  assign n14199 = po58  & ~n14198;
  assign n14200 = ~po58  & n14198;
  assign n14201 = ~n13691 & ~n13692;
  assign n14202 = po9  & n14201;
  assign n14203 = ~n13697 & ~n14202;
  assign n14204 = n13697 & n14202;
  assign n14205 = ~n14203 & ~n14204;
  assign n14206 = ~n14200 & ~n14205;
  assign n14207 = ~n14199 & ~n14206;
  assign n14208 = po59  & ~n14207;
  assign n14209 = ~po59  & n14207;
  assign n14210 = ~n13700 & ~n13701;
  assign n14211 = po9  & n14210;
  assign n14212 = ~n13706 & ~n14211;
  assign n14213 = n13706 & n14211;
  assign n14214 = ~n14212 & ~n14213;
  assign n14215 = ~n14209 & ~n14214;
  assign n14216 = ~n14208 & ~n14215;
  assign n14217 = po60  & ~n14216;
  assign n14218 = ~po60  & n14216;
  assign n14219 = ~n13709 & ~n13710;
  assign n14220 = po9  & n14219;
  assign n14221 = ~n13715 & ~n14220;
  assign n14222 = n13715 & n14220;
  assign n14223 = ~n14221 & ~n14222;
  assign n14224 = ~n14218 & ~n14223;
  assign n14225 = ~n14217 & ~n14224;
  assign n14226 = po61  & ~n14225;
  assign n14227 = ~po61  & n14225;
  assign n14228 = ~n13718 & ~n13719;
  assign n14229 = po9  & n14228;
  assign n14230 = ~n13724 & ~n14229;
  assign n14231 = n13724 & n14229;
  assign n14232 = ~n14230 & ~n14231;
  assign n14233 = ~n14227 & ~n14232;
  assign n14234 = ~n14226 & ~n14233;
  assign n14235 = po62  & ~n14234;
  assign n14236 = ~po62  & n14234;
  assign n14237 = ~n13727 & ~n13728;
  assign n14238 = po9  & n14237;
  assign n14239 = ~n13733 & ~n14238;
  assign n14240 = n13733 & n14238;
  assign n14241 = ~n14239 & ~n14240;
  assign n14242 = ~n14236 & ~n14241;
  assign n14243 = ~n14235 & ~n14242;
  assign n14244 = n14178 & n14243;
  assign n14245 = ~n14178 & ~n14243;
  assign n14246 = n13746 & po9 ;
  assign n14247 = ~n13745 & ~n14246;
  assign n14248 = n14245 & n14247;
  assign n14249 = ~po63  & ~n14248;
  assign n14250 = ~n13670 & po9 ;
  assign n14251 = n13744 & ~n14250;
  assign n14252 = po63  & ~n13746;
  assign n14253 = ~n14251 & n14252;
  assign n14254 = ~n14244 & ~n14253;
  assign n14255 = ~n14249 & n14254;
  assign po8  = n14173 | ~n14255;
  assign n14257 = ~n14171 & ~n14172;
  assign n14258 = po8  & n14257;
  assign n14259 = ~n13762 & ~n14258;
  assign n14260 = n13762 & n14258;
  assign n14261 = ~n14259 & ~n14260;
  assign n14262 = pi16  & po8 ;
  assign n14263 = ~pi14  & ~pi15 ;
  assign n14264 = ~pi16  & n14263;
  assign n14265 = ~n14262 & ~n14264;
  assign n14266 = po9  & ~n14265;
  assign n14267 = ~po9  & n14265;
  assign n14268 = ~pi16  & po8 ;
  assign n14269 = pi17  & ~n14268;
  assign n14270 = ~pi17  & n14268;
  assign n14271 = ~n14269 & ~n14270;
  assign n14272 = ~n14267 & n14271;
  assign n14273 = ~n14266 & ~n14272;
  assign n14274 = po10  & ~n14273;
  assign n14275 = ~po10  & n14273;
  assign n14276 = po9  & n14255;
  assign n14277 = ~n14270 & ~n14276;
  assign n14278 = pi18  & ~n14277;
  assign n14279 = ~pi18  & n14277;
  assign n14280 = ~n14278 & ~n14279;
  assign n14281 = ~n14275 & ~n14280;
  assign n14282 = ~n14274 & ~n14281;
  assign n14283 = po11  & ~n14282;
  assign n14284 = ~po11  & n14282;
  assign n14285 = ~n13767 & ~n13768;
  assign n14286 = po8  & n14285;
  assign n14287 = n13772 & ~n14286;
  assign n14288 = ~n13772 & n14286;
  assign n14289 = ~n14287 & ~n14288;
  assign n14290 = ~n14284 & ~n14289;
  assign n14291 = ~n14283 & ~n14290;
  assign n14292 = po12  & ~n14291;
  assign n14293 = ~po12  & n14291;
  assign n14294 = ~n13775 & ~n13776;
  assign n14295 = po8  & n14294;
  assign n14296 = ~n13781 & ~n14295;
  assign n14297 = n13781 & n14295;
  assign n14298 = ~n14296 & ~n14297;
  assign n14299 = ~n14293 & ~n14298;
  assign n14300 = ~n14292 & ~n14299;
  assign n14301 = po13  & ~n14300;
  assign n14302 = ~po13  & n14300;
  assign n14303 = ~n13784 & ~n13785;
  assign n14304 = po8  & n14303;
  assign n14305 = n13790 & n14304;
  assign n14306 = ~n13790 & ~n14304;
  assign n14307 = ~n14305 & ~n14306;
  assign n14308 = ~n14302 & ~n14307;
  assign n14309 = ~n14301 & ~n14308;
  assign n14310 = po14  & ~n14309;
  assign n14311 = ~po14  & n14309;
  assign n14312 = ~n13793 & ~n13794;
  assign n14313 = po8  & n14312;
  assign n14314 = ~n13799 & ~n14313;
  assign n14315 = n13799 & n14313;
  assign n14316 = ~n14314 & ~n14315;
  assign n14317 = ~n14311 & ~n14316;
  assign n14318 = ~n14310 & ~n14317;
  assign n14319 = po15  & ~n14318;
  assign n14320 = ~po15  & n14318;
  assign n14321 = ~n13802 & ~n13803;
  assign n14322 = po8  & n14321;
  assign n14323 = ~n13808 & ~n14322;
  assign n14324 = n13808 & n14322;
  assign n14325 = ~n14323 & ~n14324;
  assign n14326 = ~n14320 & ~n14325;
  assign n14327 = ~n14319 & ~n14326;
  assign n14328 = po16  & ~n14327;
  assign n14329 = ~po16  & n14327;
  assign n14330 = ~n13811 & ~n13812;
  assign n14331 = po8  & n14330;
  assign n14332 = ~n13817 & ~n14331;
  assign n14333 = n13817 & n14331;
  assign n14334 = ~n14332 & ~n14333;
  assign n14335 = ~n14329 & ~n14334;
  assign n14336 = ~n14328 & ~n14335;
  assign n14337 = po17  & ~n14336;
  assign n14338 = ~po17  & n14336;
  assign n14339 = ~n13820 & ~n13821;
  assign n14340 = po8  & n14339;
  assign n14341 = ~n13826 & ~n14340;
  assign n14342 = n13826 & n14340;
  assign n14343 = ~n14341 & ~n14342;
  assign n14344 = ~n14338 & ~n14343;
  assign n14345 = ~n14337 & ~n14344;
  assign n14346 = po18  & ~n14345;
  assign n14347 = ~po18  & n14345;
  assign n14348 = ~n13829 & ~n13830;
  assign n14349 = po8  & n14348;
  assign n14350 = ~n13835 & ~n14349;
  assign n14351 = n13835 & n14349;
  assign n14352 = ~n14350 & ~n14351;
  assign n14353 = ~n14347 & ~n14352;
  assign n14354 = ~n14346 & ~n14353;
  assign n14355 = po19  & ~n14354;
  assign n14356 = ~po19  & n14354;
  assign n14357 = ~n13838 & ~n13839;
  assign n14358 = po8  & n14357;
  assign n14359 = ~n13844 & ~n14358;
  assign n14360 = n13844 & n14358;
  assign n14361 = ~n14359 & ~n14360;
  assign n14362 = ~n14356 & ~n14361;
  assign n14363 = ~n14355 & ~n14362;
  assign n14364 = po20  & ~n14363;
  assign n14365 = ~po20  & n14363;
  assign n14366 = ~n13847 & ~n13848;
  assign n14367 = po8  & n14366;
  assign n14368 = ~n13853 & ~n14367;
  assign n14369 = n13853 & n14367;
  assign n14370 = ~n14368 & ~n14369;
  assign n14371 = ~n14365 & ~n14370;
  assign n14372 = ~n14364 & ~n14371;
  assign n14373 = po21  & ~n14372;
  assign n14374 = ~po21  & n14372;
  assign n14375 = ~n13856 & ~n13857;
  assign n14376 = po8  & n14375;
  assign n14377 = ~n13862 & ~n14376;
  assign n14378 = n13862 & n14376;
  assign n14379 = ~n14377 & ~n14378;
  assign n14380 = ~n14374 & ~n14379;
  assign n14381 = ~n14373 & ~n14380;
  assign n14382 = po22  & ~n14381;
  assign n14383 = ~po22  & n14381;
  assign n14384 = ~n13865 & ~n13866;
  assign n14385 = po8  & n14384;
  assign n14386 = ~n13871 & ~n14385;
  assign n14387 = n13871 & n14385;
  assign n14388 = ~n14386 & ~n14387;
  assign n14389 = ~n14383 & ~n14388;
  assign n14390 = ~n14382 & ~n14389;
  assign n14391 = po23  & ~n14390;
  assign n14392 = ~po23  & n14390;
  assign n14393 = ~n13874 & ~n13875;
  assign n14394 = po8  & n14393;
  assign n14395 = ~n13880 & ~n14394;
  assign n14396 = n13880 & n14394;
  assign n14397 = ~n14395 & ~n14396;
  assign n14398 = ~n14392 & ~n14397;
  assign n14399 = ~n14391 & ~n14398;
  assign n14400 = po24  & ~n14399;
  assign n14401 = ~po24  & n14399;
  assign n14402 = ~n13883 & ~n13884;
  assign n14403 = po8  & n14402;
  assign n14404 = ~n13889 & ~n14403;
  assign n14405 = n13889 & n14403;
  assign n14406 = ~n14404 & ~n14405;
  assign n14407 = ~n14401 & ~n14406;
  assign n14408 = ~n14400 & ~n14407;
  assign n14409 = po25  & ~n14408;
  assign n14410 = ~po25  & n14408;
  assign n14411 = ~n13892 & ~n13893;
  assign n14412 = po8  & n14411;
  assign n14413 = ~n13898 & ~n14412;
  assign n14414 = n13898 & n14412;
  assign n14415 = ~n14413 & ~n14414;
  assign n14416 = ~n14410 & ~n14415;
  assign n14417 = ~n14409 & ~n14416;
  assign n14418 = po26  & ~n14417;
  assign n14419 = ~po26  & n14417;
  assign n14420 = ~n13901 & ~n13902;
  assign n14421 = po8  & n14420;
  assign n14422 = ~n13907 & ~n14421;
  assign n14423 = n13907 & n14421;
  assign n14424 = ~n14422 & ~n14423;
  assign n14425 = ~n14419 & ~n14424;
  assign n14426 = ~n14418 & ~n14425;
  assign n14427 = po27  & ~n14426;
  assign n14428 = ~po27  & n14426;
  assign n14429 = ~n13910 & ~n13911;
  assign n14430 = po8  & n14429;
  assign n14431 = ~n13916 & ~n14430;
  assign n14432 = n13916 & n14430;
  assign n14433 = ~n14431 & ~n14432;
  assign n14434 = ~n14428 & ~n14433;
  assign n14435 = ~n14427 & ~n14434;
  assign n14436 = po28  & ~n14435;
  assign n14437 = ~po28  & n14435;
  assign n14438 = ~n13919 & ~n13920;
  assign n14439 = po8  & n14438;
  assign n14440 = ~n13925 & ~n14439;
  assign n14441 = n13925 & n14439;
  assign n14442 = ~n14440 & ~n14441;
  assign n14443 = ~n14437 & ~n14442;
  assign n14444 = ~n14436 & ~n14443;
  assign n14445 = po29  & ~n14444;
  assign n14446 = ~po29  & n14444;
  assign n14447 = ~n13928 & ~n13929;
  assign n14448 = po8  & n14447;
  assign n14449 = ~n13934 & ~n14448;
  assign n14450 = n13934 & n14448;
  assign n14451 = ~n14449 & ~n14450;
  assign n14452 = ~n14446 & ~n14451;
  assign n14453 = ~n14445 & ~n14452;
  assign n14454 = po30  & ~n14453;
  assign n14455 = ~po30  & n14453;
  assign n14456 = ~n13937 & ~n13938;
  assign n14457 = po8  & n14456;
  assign n14458 = ~n13943 & ~n14457;
  assign n14459 = n13943 & n14457;
  assign n14460 = ~n14458 & ~n14459;
  assign n14461 = ~n14455 & ~n14460;
  assign n14462 = ~n14454 & ~n14461;
  assign n14463 = po31  & ~n14462;
  assign n14464 = ~po31  & n14462;
  assign n14465 = ~n13946 & ~n13947;
  assign n14466 = po8  & n14465;
  assign n14467 = ~n13952 & ~n14466;
  assign n14468 = n13952 & n14466;
  assign n14469 = ~n14467 & ~n14468;
  assign n14470 = ~n14464 & ~n14469;
  assign n14471 = ~n14463 & ~n14470;
  assign n14472 = po32  & ~n14471;
  assign n14473 = ~po32  & n14471;
  assign n14474 = ~n13955 & ~n13956;
  assign n14475 = po8  & n14474;
  assign n14476 = ~n13961 & ~n14475;
  assign n14477 = n13961 & n14475;
  assign n14478 = ~n14476 & ~n14477;
  assign n14479 = ~n14473 & ~n14478;
  assign n14480 = ~n14472 & ~n14479;
  assign n14481 = po33  & ~n14480;
  assign n14482 = ~po33  & n14480;
  assign n14483 = ~n13964 & ~n13965;
  assign n14484 = po8  & n14483;
  assign n14485 = ~n13970 & ~n14484;
  assign n14486 = n13970 & n14484;
  assign n14487 = ~n14485 & ~n14486;
  assign n14488 = ~n14482 & ~n14487;
  assign n14489 = ~n14481 & ~n14488;
  assign n14490 = po34  & ~n14489;
  assign n14491 = ~po34  & n14489;
  assign n14492 = ~n13973 & ~n13974;
  assign n14493 = po8  & n14492;
  assign n14494 = ~n13979 & ~n14493;
  assign n14495 = n13979 & n14493;
  assign n14496 = ~n14494 & ~n14495;
  assign n14497 = ~n14491 & ~n14496;
  assign n14498 = ~n14490 & ~n14497;
  assign n14499 = po35  & ~n14498;
  assign n14500 = ~po35  & n14498;
  assign n14501 = ~n13982 & ~n13983;
  assign n14502 = po8  & n14501;
  assign n14503 = ~n13988 & ~n14502;
  assign n14504 = n13988 & n14502;
  assign n14505 = ~n14503 & ~n14504;
  assign n14506 = ~n14500 & ~n14505;
  assign n14507 = ~n14499 & ~n14506;
  assign n14508 = po36  & ~n14507;
  assign n14509 = ~po36  & n14507;
  assign n14510 = ~n13991 & ~n13992;
  assign n14511 = po8  & n14510;
  assign n14512 = ~n13997 & ~n14511;
  assign n14513 = n13997 & n14511;
  assign n14514 = ~n14512 & ~n14513;
  assign n14515 = ~n14509 & ~n14514;
  assign n14516 = ~n14508 & ~n14515;
  assign n14517 = po37  & ~n14516;
  assign n14518 = ~po37  & n14516;
  assign n14519 = ~n14000 & ~n14001;
  assign n14520 = po8  & n14519;
  assign n14521 = ~n14006 & ~n14520;
  assign n14522 = n14006 & n14520;
  assign n14523 = ~n14521 & ~n14522;
  assign n14524 = ~n14518 & ~n14523;
  assign n14525 = ~n14517 & ~n14524;
  assign n14526 = po38  & ~n14525;
  assign n14527 = ~po38  & n14525;
  assign n14528 = ~n14009 & ~n14010;
  assign n14529 = po8  & n14528;
  assign n14530 = ~n14015 & ~n14529;
  assign n14531 = n14015 & n14529;
  assign n14532 = ~n14530 & ~n14531;
  assign n14533 = ~n14527 & ~n14532;
  assign n14534 = ~n14526 & ~n14533;
  assign n14535 = po39  & ~n14534;
  assign n14536 = ~po39  & n14534;
  assign n14537 = ~n14018 & ~n14019;
  assign n14538 = po8  & n14537;
  assign n14539 = ~n14024 & ~n14538;
  assign n14540 = n14024 & n14538;
  assign n14541 = ~n14539 & ~n14540;
  assign n14542 = ~n14536 & ~n14541;
  assign n14543 = ~n14535 & ~n14542;
  assign n14544 = po40  & ~n14543;
  assign n14545 = ~po40  & n14543;
  assign n14546 = ~n14027 & ~n14028;
  assign n14547 = po8  & n14546;
  assign n14548 = ~n14033 & ~n14547;
  assign n14549 = n14033 & n14547;
  assign n14550 = ~n14548 & ~n14549;
  assign n14551 = ~n14545 & ~n14550;
  assign n14552 = ~n14544 & ~n14551;
  assign n14553 = po41  & ~n14552;
  assign n14554 = ~po41  & n14552;
  assign n14555 = ~n14036 & ~n14037;
  assign n14556 = po8  & n14555;
  assign n14557 = ~n14042 & ~n14556;
  assign n14558 = n14042 & n14556;
  assign n14559 = ~n14557 & ~n14558;
  assign n14560 = ~n14554 & ~n14559;
  assign n14561 = ~n14553 & ~n14560;
  assign n14562 = po42  & ~n14561;
  assign n14563 = ~po42  & n14561;
  assign n14564 = ~n14045 & ~n14046;
  assign n14565 = po8  & n14564;
  assign n14566 = ~n14051 & ~n14565;
  assign n14567 = n14051 & n14565;
  assign n14568 = ~n14566 & ~n14567;
  assign n14569 = ~n14563 & ~n14568;
  assign n14570 = ~n14562 & ~n14569;
  assign n14571 = po43  & ~n14570;
  assign n14572 = ~po43  & n14570;
  assign n14573 = ~n14054 & ~n14055;
  assign n14574 = po8  & n14573;
  assign n14575 = ~n14060 & ~n14574;
  assign n14576 = n14060 & n14574;
  assign n14577 = ~n14575 & ~n14576;
  assign n14578 = ~n14572 & ~n14577;
  assign n14579 = ~n14571 & ~n14578;
  assign n14580 = po44  & ~n14579;
  assign n14581 = ~po44  & n14579;
  assign n14582 = ~n14063 & ~n14064;
  assign n14583 = po8  & n14582;
  assign n14584 = ~n14069 & ~n14583;
  assign n14585 = n14069 & n14583;
  assign n14586 = ~n14584 & ~n14585;
  assign n14587 = ~n14581 & ~n14586;
  assign n14588 = ~n14580 & ~n14587;
  assign n14589 = po45  & ~n14588;
  assign n14590 = ~po45  & n14588;
  assign n14591 = ~n14072 & ~n14073;
  assign n14592 = po8  & n14591;
  assign n14593 = ~n14078 & ~n14592;
  assign n14594 = n14078 & n14592;
  assign n14595 = ~n14593 & ~n14594;
  assign n14596 = ~n14590 & ~n14595;
  assign n14597 = ~n14589 & ~n14596;
  assign n14598 = po46  & ~n14597;
  assign n14599 = ~po46  & n14597;
  assign n14600 = ~n14081 & ~n14082;
  assign n14601 = po8  & n14600;
  assign n14602 = ~n14087 & ~n14601;
  assign n14603 = n14087 & n14601;
  assign n14604 = ~n14602 & ~n14603;
  assign n14605 = ~n14599 & ~n14604;
  assign n14606 = ~n14598 & ~n14605;
  assign n14607 = po47  & ~n14606;
  assign n14608 = ~po47  & n14606;
  assign n14609 = ~n14090 & ~n14091;
  assign n14610 = po8  & n14609;
  assign n14611 = ~n14096 & ~n14610;
  assign n14612 = n14096 & n14610;
  assign n14613 = ~n14611 & ~n14612;
  assign n14614 = ~n14608 & ~n14613;
  assign n14615 = ~n14607 & ~n14614;
  assign n14616 = po48  & ~n14615;
  assign n14617 = ~po48  & n14615;
  assign n14618 = ~n14099 & ~n14100;
  assign n14619 = po8  & n14618;
  assign n14620 = ~n14105 & ~n14619;
  assign n14621 = n14105 & n14619;
  assign n14622 = ~n14620 & ~n14621;
  assign n14623 = ~n14617 & ~n14622;
  assign n14624 = ~n14616 & ~n14623;
  assign n14625 = po49  & ~n14624;
  assign n14626 = ~po49  & n14624;
  assign n14627 = ~n14108 & ~n14109;
  assign n14628 = po8  & n14627;
  assign n14629 = ~n14114 & ~n14628;
  assign n14630 = n14114 & n14628;
  assign n14631 = ~n14629 & ~n14630;
  assign n14632 = ~n14626 & ~n14631;
  assign n14633 = ~n14625 & ~n14632;
  assign n14634 = po50  & ~n14633;
  assign n14635 = ~po50  & n14633;
  assign n14636 = ~n14117 & ~n14118;
  assign n14637 = po8  & n14636;
  assign n14638 = ~n14123 & ~n14637;
  assign n14639 = n14123 & n14637;
  assign n14640 = ~n14638 & ~n14639;
  assign n14641 = ~n14635 & ~n14640;
  assign n14642 = ~n14634 & ~n14641;
  assign n14643 = po51  & ~n14642;
  assign n14644 = ~po51  & n14642;
  assign n14645 = ~n14126 & ~n14127;
  assign n14646 = po8  & n14645;
  assign n14647 = ~n14132 & ~n14646;
  assign n14648 = n14132 & n14646;
  assign n14649 = ~n14647 & ~n14648;
  assign n14650 = ~n14644 & ~n14649;
  assign n14651 = ~n14643 & ~n14650;
  assign n14652 = po52  & ~n14651;
  assign n14653 = ~po52  & n14651;
  assign n14654 = ~n14135 & ~n14136;
  assign n14655 = po8  & n14654;
  assign n14656 = ~n14141 & ~n14655;
  assign n14657 = n14141 & n14655;
  assign n14658 = ~n14656 & ~n14657;
  assign n14659 = ~n14653 & ~n14658;
  assign n14660 = ~n14652 & ~n14659;
  assign n14661 = po53  & ~n14660;
  assign n14662 = ~po53  & n14660;
  assign n14663 = ~n14144 & ~n14145;
  assign n14664 = po8  & n14663;
  assign n14665 = ~n14150 & ~n14664;
  assign n14666 = n14150 & n14664;
  assign n14667 = ~n14665 & ~n14666;
  assign n14668 = ~n14662 & ~n14667;
  assign n14669 = ~n14661 & ~n14668;
  assign n14670 = po54  & ~n14669;
  assign n14671 = ~po54  & n14669;
  assign n14672 = ~n14153 & ~n14154;
  assign n14673 = po8  & n14672;
  assign n14674 = ~n14159 & ~n14673;
  assign n14675 = n14159 & n14673;
  assign n14676 = ~n14674 & ~n14675;
  assign n14677 = ~n14671 & ~n14676;
  assign n14678 = ~n14670 & ~n14677;
  assign n14679 = po55  & ~n14678;
  assign n14680 = ~n14162 & ~n14168;
  assign n14681 = po8  & n14680;
  assign n14682 = ~n14167 & ~n14681;
  assign n14683 = n14167 & n14681;
  assign n14684 = ~n14682 & ~n14683;
  assign n14685 = ~po55  & n14678;
  assign n14686 = ~n14684 & ~n14685;
  assign n14687 = ~n14679 & ~n14686;
  assign n14688 = po56  & ~n14687;
  assign n14689 = ~po56  & n14687;
  assign n14690 = n14178 & ~po8 ;
  assign n14691 = ~n14235 & ~n14236;
  assign n14692 = po8  & n14691;
  assign n14693 = ~n14241 & ~n14692;
  assign n14694 = n14241 & n14692;
  assign n14695 = ~n14693 & ~n14694;
  assign n14696 = ~n14261 & ~n14689;
  assign n14697 = ~n14688 & ~n14696;
  assign n14698 = po57  & ~n14697;
  assign n14699 = ~po57  & n14697;
  assign n14700 = ~n14181 & ~n14182;
  assign n14701 = po8  & n14700;
  assign n14702 = ~n14187 & ~n14701;
  assign n14703 = n14187 & n14701;
  assign n14704 = ~n14702 & ~n14703;
  assign n14705 = ~n14699 & ~n14704;
  assign n14706 = ~n14698 & ~n14705;
  assign n14707 = po58  & ~n14706;
  assign n14708 = ~po58  & n14706;
  assign n14709 = ~n14190 & ~n14191;
  assign n14710 = po8  & n14709;
  assign n14711 = ~n14196 & ~n14710;
  assign n14712 = n14196 & n14710;
  assign n14713 = ~n14711 & ~n14712;
  assign n14714 = ~n14708 & ~n14713;
  assign n14715 = ~n14707 & ~n14714;
  assign n14716 = po59  & ~n14715;
  assign n14717 = ~po59  & n14715;
  assign n14718 = ~n14199 & ~n14200;
  assign n14719 = po8  & n14718;
  assign n14720 = ~n14205 & ~n14719;
  assign n14721 = n14205 & n14719;
  assign n14722 = ~n14720 & ~n14721;
  assign n14723 = ~n14717 & ~n14722;
  assign n14724 = ~n14716 & ~n14723;
  assign n14725 = po60  & ~n14724;
  assign n14726 = ~po60  & n14724;
  assign n14727 = ~n14208 & ~n14209;
  assign n14728 = po8  & n14727;
  assign n14729 = ~n14214 & ~n14728;
  assign n14730 = n14214 & n14728;
  assign n14731 = ~n14729 & ~n14730;
  assign n14732 = ~n14726 & ~n14731;
  assign n14733 = ~n14725 & ~n14732;
  assign n14734 = po61  & ~n14733;
  assign n14735 = ~po61  & n14733;
  assign n14736 = ~n14217 & ~n14218;
  assign n14737 = po8  & n14736;
  assign n14738 = ~n14223 & ~n14737;
  assign n14739 = n14223 & n14737;
  assign n14740 = ~n14738 & ~n14739;
  assign n14741 = ~n14735 & ~n14740;
  assign n14742 = ~n14734 & ~n14741;
  assign n14743 = po62  & ~n14742;
  assign n14744 = ~po62  & n14742;
  assign n14745 = ~n14226 & ~n14227;
  assign n14746 = po8  & n14745;
  assign n14747 = ~n14232 & ~n14746;
  assign n14748 = n14232 & n14746;
  assign n14749 = ~n14747 & ~n14748;
  assign n14750 = ~n14744 & ~n14749;
  assign n14751 = ~n14743 & ~n14750;
  assign n14752 = n14695 & n14751;
  assign n14753 = ~n14695 & ~n14751;
  assign n14754 = n14245 & po8 ;
  assign n14755 = ~n14244 & ~n14754;
  assign n14756 = n14753 & n14755;
  assign n14757 = ~po63  & ~n14756;
  assign n14758 = ~n14178 & po8 ;
  assign n14759 = n14243 & ~n14758;
  assign n14760 = po63  & ~n14245;
  assign n14761 = ~n14759 & n14760;
  assign n14762 = ~n14752 & ~n14761;
  assign n14763 = ~n14757 & n14762;
  assign po7  = n14690 | ~n14763;
  assign n14765 = ~n14688 & ~n14689;
  assign n14766 = po7  & n14765;
  assign n14767 = ~n14261 & ~n14766;
  assign n14768 = n14261 & n14766;
  assign n14769 = ~n14767 & ~n14768;
  assign n14770 = pi14  & po7 ;
  assign n14771 = ~pi12  & ~pi13 ;
  assign n14772 = ~pi14  & n14771;
  assign n14773 = ~n14770 & ~n14772;
  assign n14774 = po8  & ~n14773;
  assign n14775 = ~po8  & n14773;
  assign n14776 = ~pi14  & po7 ;
  assign n14777 = pi15  & ~n14776;
  assign n14778 = ~pi15  & n14776;
  assign n14779 = ~n14777 & ~n14778;
  assign n14780 = ~n14775 & n14779;
  assign n14781 = ~n14774 & ~n14780;
  assign n14782 = po9  & ~n14781;
  assign n14783 = ~po9  & n14781;
  assign n14784 = po8  & n14763;
  assign n14785 = ~n14778 & ~n14784;
  assign n14786 = pi16  & ~n14785;
  assign n14787 = ~pi16  & n14785;
  assign n14788 = ~n14786 & ~n14787;
  assign n14789 = ~n14783 & ~n14788;
  assign n14790 = ~n14782 & ~n14789;
  assign n14791 = po10  & ~n14790;
  assign n14792 = ~po10  & n14790;
  assign n14793 = ~n14266 & ~n14267;
  assign n14794 = po7  & n14793;
  assign n14795 = n14271 & ~n14794;
  assign n14796 = ~n14271 & n14794;
  assign n14797 = ~n14795 & ~n14796;
  assign n14798 = ~n14792 & ~n14797;
  assign n14799 = ~n14791 & ~n14798;
  assign n14800 = po11  & ~n14799;
  assign n14801 = ~po11  & n14799;
  assign n14802 = ~n14274 & ~n14275;
  assign n14803 = po7  & n14802;
  assign n14804 = ~n14280 & ~n14803;
  assign n14805 = n14280 & n14803;
  assign n14806 = ~n14804 & ~n14805;
  assign n14807 = ~n14801 & ~n14806;
  assign n14808 = ~n14800 & ~n14807;
  assign n14809 = po12  & ~n14808;
  assign n14810 = ~po12  & n14808;
  assign n14811 = ~n14283 & ~n14284;
  assign n14812 = po7  & n14811;
  assign n14813 = n14289 & n14812;
  assign n14814 = ~n14289 & ~n14812;
  assign n14815 = ~n14813 & ~n14814;
  assign n14816 = ~n14810 & ~n14815;
  assign n14817 = ~n14809 & ~n14816;
  assign n14818 = po13  & ~n14817;
  assign n14819 = ~po13  & n14817;
  assign n14820 = ~n14292 & ~n14293;
  assign n14821 = po7  & n14820;
  assign n14822 = ~n14298 & ~n14821;
  assign n14823 = n14298 & n14821;
  assign n14824 = ~n14822 & ~n14823;
  assign n14825 = ~n14819 & ~n14824;
  assign n14826 = ~n14818 & ~n14825;
  assign n14827 = po14  & ~n14826;
  assign n14828 = ~po14  & n14826;
  assign n14829 = ~n14301 & ~n14302;
  assign n14830 = po7  & n14829;
  assign n14831 = ~n14307 & ~n14830;
  assign n14832 = n14307 & n14830;
  assign n14833 = ~n14831 & ~n14832;
  assign n14834 = ~n14828 & ~n14833;
  assign n14835 = ~n14827 & ~n14834;
  assign n14836 = po15  & ~n14835;
  assign n14837 = ~po15  & n14835;
  assign n14838 = ~n14310 & ~n14311;
  assign n14839 = po7  & n14838;
  assign n14840 = ~n14316 & ~n14839;
  assign n14841 = n14316 & n14839;
  assign n14842 = ~n14840 & ~n14841;
  assign n14843 = ~n14837 & ~n14842;
  assign n14844 = ~n14836 & ~n14843;
  assign n14845 = po16  & ~n14844;
  assign n14846 = ~po16  & n14844;
  assign n14847 = ~n14319 & ~n14320;
  assign n14848 = po7  & n14847;
  assign n14849 = ~n14325 & ~n14848;
  assign n14850 = n14325 & n14848;
  assign n14851 = ~n14849 & ~n14850;
  assign n14852 = ~n14846 & ~n14851;
  assign n14853 = ~n14845 & ~n14852;
  assign n14854 = po17  & ~n14853;
  assign n14855 = ~po17  & n14853;
  assign n14856 = ~n14328 & ~n14329;
  assign n14857 = po7  & n14856;
  assign n14858 = ~n14334 & ~n14857;
  assign n14859 = n14334 & n14857;
  assign n14860 = ~n14858 & ~n14859;
  assign n14861 = ~n14855 & ~n14860;
  assign n14862 = ~n14854 & ~n14861;
  assign n14863 = po18  & ~n14862;
  assign n14864 = ~po18  & n14862;
  assign n14865 = ~n14337 & ~n14338;
  assign n14866 = po7  & n14865;
  assign n14867 = ~n14343 & ~n14866;
  assign n14868 = n14343 & n14866;
  assign n14869 = ~n14867 & ~n14868;
  assign n14870 = ~n14864 & ~n14869;
  assign n14871 = ~n14863 & ~n14870;
  assign n14872 = po19  & ~n14871;
  assign n14873 = ~po19  & n14871;
  assign n14874 = ~n14346 & ~n14347;
  assign n14875 = po7  & n14874;
  assign n14876 = ~n14352 & ~n14875;
  assign n14877 = n14352 & n14875;
  assign n14878 = ~n14876 & ~n14877;
  assign n14879 = ~n14873 & ~n14878;
  assign n14880 = ~n14872 & ~n14879;
  assign n14881 = po20  & ~n14880;
  assign n14882 = ~po20  & n14880;
  assign n14883 = ~n14355 & ~n14356;
  assign n14884 = po7  & n14883;
  assign n14885 = ~n14361 & ~n14884;
  assign n14886 = n14361 & n14884;
  assign n14887 = ~n14885 & ~n14886;
  assign n14888 = ~n14882 & ~n14887;
  assign n14889 = ~n14881 & ~n14888;
  assign n14890 = po21  & ~n14889;
  assign n14891 = ~po21  & n14889;
  assign n14892 = ~n14364 & ~n14365;
  assign n14893 = po7  & n14892;
  assign n14894 = ~n14370 & ~n14893;
  assign n14895 = n14370 & n14893;
  assign n14896 = ~n14894 & ~n14895;
  assign n14897 = ~n14891 & ~n14896;
  assign n14898 = ~n14890 & ~n14897;
  assign n14899 = po22  & ~n14898;
  assign n14900 = ~po22  & n14898;
  assign n14901 = ~n14373 & ~n14374;
  assign n14902 = po7  & n14901;
  assign n14903 = ~n14379 & ~n14902;
  assign n14904 = n14379 & n14902;
  assign n14905 = ~n14903 & ~n14904;
  assign n14906 = ~n14900 & ~n14905;
  assign n14907 = ~n14899 & ~n14906;
  assign n14908 = po23  & ~n14907;
  assign n14909 = ~po23  & n14907;
  assign n14910 = ~n14382 & ~n14383;
  assign n14911 = po7  & n14910;
  assign n14912 = ~n14388 & ~n14911;
  assign n14913 = n14388 & n14911;
  assign n14914 = ~n14912 & ~n14913;
  assign n14915 = ~n14909 & ~n14914;
  assign n14916 = ~n14908 & ~n14915;
  assign n14917 = po24  & ~n14916;
  assign n14918 = ~po24  & n14916;
  assign n14919 = ~n14391 & ~n14392;
  assign n14920 = po7  & n14919;
  assign n14921 = ~n14397 & ~n14920;
  assign n14922 = n14397 & n14920;
  assign n14923 = ~n14921 & ~n14922;
  assign n14924 = ~n14918 & ~n14923;
  assign n14925 = ~n14917 & ~n14924;
  assign n14926 = po25  & ~n14925;
  assign n14927 = ~po25  & n14925;
  assign n14928 = ~n14400 & ~n14401;
  assign n14929 = po7  & n14928;
  assign n14930 = ~n14406 & ~n14929;
  assign n14931 = n14406 & n14929;
  assign n14932 = ~n14930 & ~n14931;
  assign n14933 = ~n14927 & ~n14932;
  assign n14934 = ~n14926 & ~n14933;
  assign n14935 = po26  & ~n14934;
  assign n14936 = ~po26  & n14934;
  assign n14937 = ~n14409 & ~n14410;
  assign n14938 = po7  & n14937;
  assign n14939 = ~n14415 & ~n14938;
  assign n14940 = n14415 & n14938;
  assign n14941 = ~n14939 & ~n14940;
  assign n14942 = ~n14936 & ~n14941;
  assign n14943 = ~n14935 & ~n14942;
  assign n14944 = po27  & ~n14943;
  assign n14945 = ~po27  & n14943;
  assign n14946 = ~n14418 & ~n14419;
  assign n14947 = po7  & n14946;
  assign n14948 = ~n14424 & ~n14947;
  assign n14949 = n14424 & n14947;
  assign n14950 = ~n14948 & ~n14949;
  assign n14951 = ~n14945 & ~n14950;
  assign n14952 = ~n14944 & ~n14951;
  assign n14953 = po28  & ~n14952;
  assign n14954 = ~po28  & n14952;
  assign n14955 = ~n14427 & ~n14428;
  assign n14956 = po7  & n14955;
  assign n14957 = ~n14433 & ~n14956;
  assign n14958 = n14433 & n14956;
  assign n14959 = ~n14957 & ~n14958;
  assign n14960 = ~n14954 & ~n14959;
  assign n14961 = ~n14953 & ~n14960;
  assign n14962 = po29  & ~n14961;
  assign n14963 = ~po29  & n14961;
  assign n14964 = ~n14436 & ~n14437;
  assign n14965 = po7  & n14964;
  assign n14966 = ~n14442 & ~n14965;
  assign n14967 = n14442 & n14965;
  assign n14968 = ~n14966 & ~n14967;
  assign n14969 = ~n14963 & ~n14968;
  assign n14970 = ~n14962 & ~n14969;
  assign n14971 = po30  & ~n14970;
  assign n14972 = ~po30  & n14970;
  assign n14973 = ~n14445 & ~n14446;
  assign n14974 = po7  & n14973;
  assign n14975 = ~n14451 & ~n14974;
  assign n14976 = n14451 & n14974;
  assign n14977 = ~n14975 & ~n14976;
  assign n14978 = ~n14972 & ~n14977;
  assign n14979 = ~n14971 & ~n14978;
  assign n14980 = po31  & ~n14979;
  assign n14981 = ~po31  & n14979;
  assign n14982 = ~n14454 & ~n14455;
  assign n14983 = po7  & n14982;
  assign n14984 = ~n14460 & ~n14983;
  assign n14985 = n14460 & n14983;
  assign n14986 = ~n14984 & ~n14985;
  assign n14987 = ~n14981 & ~n14986;
  assign n14988 = ~n14980 & ~n14987;
  assign n14989 = po32  & ~n14988;
  assign n14990 = ~po32  & n14988;
  assign n14991 = ~n14463 & ~n14464;
  assign n14992 = po7  & n14991;
  assign n14993 = ~n14469 & ~n14992;
  assign n14994 = n14469 & n14992;
  assign n14995 = ~n14993 & ~n14994;
  assign n14996 = ~n14990 & ~n14995;
  assign n14997 = ~n14989 & ~n14996;
  assign n14998 = po33  & ~n14997;
  assign n14999 = ~po33  & n14997;
  assign n15000 = ~n14472 & ~n14473;
  assign n15001 = po7  & n15000;
  assign n15002 = ~n14478 & ~n15001;
  assign n15003 = n14478 & n15001;
  assign n15004 = ~n15002 & ~n15003;
  assign n15005 = ~n14999 & ~n15004;
  assign n15006 = ~n14998 & ~n15005;
  assign n15007 = po34  & ~n15006;
  assign n15008 = ~po34  & n15006;
  assign n15009 = ~n14481 & ~n14482;
  assign n15010 = po7  & n15009;
  assign n15011 = ~n14487 & ~n15010;
  assign n15012 = n14487 & n15010;
  assign n15013 = ~n15011 & ~n15012;
  assign n15014 = ~n15008 & ~n15013;
  assign n15015 = ~n15007 & ~n15014;
  assign n15016 = po35  & ~n15015;
  assign n15017 = ~po35  & n15015;
  assign n15018 = ~n14490 & ~n14491;
  assign n15019 = po7  & n15018;
  assign n15020 = ~n14496 & ~n15019;
  assign n15021 = n14496 & n15019;
  assign n15022 = ~n15020 & ~n15021;
  assign n15023 = ~n15017 & ~n15022;
  assign n15024 = ~n15016 & ~n15023;
  assign n15025 = po36  & ~n15024;
  assign n15026 = ~po36  & n15024;
  assign n15027 = ~n14499 & ~n14500;
  assign n15028 = po7  & n15027;
  assign n15029 = ~n14505 & ~n15028;
  assign n15030 = n14505 & n15028;
  assign n15031 = ~n15029 & ~n15030;
  assign n15032 = ~n15026 & ~n15031;
  assign n15033 = ~n15025 & ~n15032;
  assign n15034 = po37  & ~n15033;
  assign n15035 = ~po37  & n15033;
  assign n15036 = ~n14508 & ~n14509;
  assign n15037 = po7  & n15036;
  assign n15038 = ~n14514 & ~n15037;
  assign n15039 = n14514 & n15037;
  assign n15040 = ~n15038 & ~n15039;
  assign n15041 = ~n15035 & ~n15040;
  assign n15042 = ~n15034 & ~n15041;
  assign n15043 = po38  & ~n15042;
  assign n15044 = ~po38  & n15042;
  assign n15045 = ~n14517 & ~n14518;
  assign n15046 = po7  & n15045;
  assign n15047 = ~n14523 & ~n15046;
  assign n15048 = n14523 & n15046;
  assign n15049 = ~n15047 & ~n15048;
  assign n15050 = ~n15044 & ~n15049;
  assign n15051 = ~n15043 & ~n15050;
  assign n15052 = po39  & ~n15051;
  assign n15053 = ~po39  & n15051;
  assign n15054 = ~n14526 & ~n14527;
  assign n15055 = po7  & n15054;
  assign n15056 = ~n14532 & ~n15055;
  assign n15057 = n14532 & n15055;
  assign n15058 = ~n15056 & ~n15057;
  assign n15059 = ~n15053 & ~n15058;
  assign n15060 = ~n15052 & ~n15059;
  assign n15061 = po40  & ~n15060;
  assign n15062 = ~po40  & n15060;
  assign n15063 = ~n14535 & ~n14536;
  assign n15064 = po7  & n15063;
  assign n15065 = ~n14541 & ~n15064;
  assign n15066 = n14541 & n15064;
  assign n15067 = ~n15065 & ~n15066;
  assign n15068 = ~n15062 & ~n15067;
  assign n15069 = ~n15061 & ~n15068;
  assign n15070 = po41  & ~n15069;
  assign n15071 = ~po41  & n15069;
  assign n15072 = ~n14544 & ~n14545;
  assign n15073 = po7  & n15072;
  assign n15074 = ~n14550 & ~n15073;
  assign n15075 = n14550 & n15073;
  assign n15076 = ~n15074 & ~n15075;
  assign n15077 = ~n15071 & ~n15076;
  assign n15078 = ~n15070 & ~n15077;
  assign n15079 = po42  & ~n15078;
  assign n15080 = ~po42  & n15078;
  assign n15081 = ~n14553 & ~n14554;
  assign n15082 = po7  & n15081;
  assign n15083 = ~n14559 & ~n15082;
  assign n15084 = n14559 & n15082;
  assign n15085 = ~n15083 & ~n15084;
  assign n15086 = ~n15080 & ~n15085;
  assign n15087 = ~n15079 & ~n15086;
  assign n15088 = po43  & ~n15087;
  assign n15089 = ~po43  & n15087;
  assign n15090 = ~n14562 & ~n14563;
  assign n15091 = po7  & n15090;
  assign n15092 = ~n14568 & ~n15091;
  assign n15093 = n14568 & n15091;
  assign n15094 = ~n15092 & ~n15093;
  assign n15095 = ~n15089 & ~n15094;
  assign n15096 = ~n15088 & ~n15095;
  assign n15097 = po44  & ~n15096;
  assign n15098 = ~po44  & n15096;
  assign n15099 = ~n14571 & ~n14572;
  assign n15100 = po7  & n15099;
  assign n15101 = ~n14577 & ~n15100;
  assign n15102 = n14577 & n15100;
  assign n15103 = ~n15101 & ~n15102;
  assign n15104 = ~n15098 & ~n15103;
  assign n15105 = ~n15097 & ~n15104;
  assign n15106 = po45  & ~n15105;
  assign n15107 = ~po45  & n15105;
  assign n15108 = ~n14580 & ~n14581;
  assign n15109 = po7  & n15108;
  assign n15110 = ~n14586 & ~n15109;
  assign n15111 = n14586 & n15109;
  assign n15112 = ~n15110 & ~n15111;
  assign n15113 = ~n15107 & ~n15112;
  assign n15114 = ~n15106 & ~n15113;
  assign n15115 = po46  & ~n15114;
  assign n15116 = ~po46  & n15114;
  assign n15117 = ~n14589 & ~n14590;
  assign n15118 = po7  & n15117;
  assign n15119 = ~n14595 & ~n15118;
  assign n15120 = n14595 & n15118;
  assign n15121 = ~n15119 & ~n15120;
  assign n15122 = ~n15116 & ~n15121;
  assign n15123 = ~n15115 & ~n15122;
  assign n15124 = po47  & ~n15123;
  assign n15125 = ~po47  & n15123;
  assign n15126 = ~n14598 & ~n14599;
  assign n15127 = po7  & n15126;
  assign n15128 = ~n14604 & ~n15127;
  assign n15129 = n14604 & n15127;
  assign n15130 = ~n15128 & ~n15129;
  assign n15131 = ~n15125 & ~n15130;
  assign n15132 = ~n15124 & ~n15131;
  assign n15133 = po48  & ~n15132;
  assign n15134 = ~po48  & n15132;
  assign n15135 = ~n14607 & ~n14608;
  assign n15136 = po7  & n15135;
  assign n15137 = ~n14613 & ~n15136;
  assign n15138 = n14613 & n15136;
  assign n15139 = ~n15137 & ~n15138;
  assign n15140 = ~n15134 & ~n15139;
  assign n15141 = ~n15133 & ~n15140;
  assign n15142 = po49  & ~n15141;
  assign n15143 = ~po49  & n15141;
  assign n15144 = ~n14616 & ~n14617;
  assign n15145 = po7  & n15144;
  assign n15146 = ~n14622 & ~n15145;
  assign n15147 = n14622 & n15145;
  assign n15148 = ~n15146 & ~n15147;
  assign n15149 = ~n15143 & ~n15148;
  assign n15150 = ~n15142 & ~n15149;
  assign n15151 = po50  & ~n15150;
  assign n15152 = ~po50  & n15150;
  assign n15153 = ~n14625 & ~n14626;
  assign n15154 = po7  & n15153;
  assign n15155 = ~n14631 & ~n15154;
  assign n15156 = n14631 & n15154;
  assign n15157 = ~n15155 & ~n15156;
  assign n15158 = ~n15152 & ~n15157;
  assign n15159 = ~n15151 & ~n15158;
  assign n15160 = po51  & ~n15159;
  assign n15161 = ~po51  & n15159;
  assign n15162 = ~n14634 & ~n14635;
  assign n15163 = po7  & n15162;
  assign n15164 = ~n14640 & ~n15163;
  assign n15165 = n14640 & n15163;
  assign n15166 = ~n15164 & ~n15165;
  assign n15167 = ~n15161 & ~n15166;
  assign n15168 = ~n15160 & ~n15167;
  assign n15169 = po52  & ~n15168;
  assign n15170 = ~po52  & n15168;
  assign n15171 = ~n14643 & ~n14644;
  assign n15172 = po7  & n15171;
  assign n15173 = ~n14649 & ~n15172;
  assign n15174 = n14649 & n15172;
  assign n15175 = ~n15173 & ~n15174;
  assign n15176 = ~n15170 & ~n15175;
  assign n15177 = ~n15169 & ~n15176;
  assign n15178 = po53  & ~n15177;
  assign n15179 = ~po53  & n15177;
  assign n15180 = ~n14652 & ~n14653;
  assign n15181 = po7  & n15180;
  assign n15182 = ~n14658 & ~n15181;
  assign n15183 = n14658 & n15181;
  assign n15184 = ~n15182 & ~n15183;
  assign n15185 = ~n15179 & ~n15184;
  assign n15186 = ~n15178 & ~n15185;
  assign n15187 = po54  & ~n15186;
  assign n15188 = ~po54  & n15186;
  assign n15189 = ~n14661 & ~n14662;
  assign n15190 = po7  & n15189;
  assign n15191 = ~n14667 & ~n15190;
  assign n15192 = n14667 & n15190;
  assign n15193 = ~n15191 & ~n15192;
  assign n15194 = ~n15188 & ~n15193;
  assign n15195 = ~n15187 & ~n15194;
  assign n15196 = po55  & ~n15195;
  assign n15197 = ~po55  & n15195;
  assign n15198 = ~n14670 & ~n14671;
  assign n15199 = po7  & n15198;
  assign n15200 = ~n14676 & ~n15199;
  assign n15201 = n14676 & n15199;
  assign n15202 = ~n15200 & ~n15201;
  assign n15203 = ~n15197 & ~n15202;
  assign n15204 = ~n15196 & ~n15203;
  assign n15205 = po56  & ~n15204;
  assign n15206 = ~n14679 & ~n14685;
  assign n15207 = po7  & n15206;
  assign n15208 = ~n14684 & ~n15207;
  assign n15209 = n14684 & n15207;
  assign n15210 = ~n15208 & ~n15209;
  assign n15211 = ~po56  & n15204;
  assign n15212 = ~n15210 & ~n15211;
  assign n15213 = ~n15205 & ~n15212;
  assign n15214 = po57  & ~n15213;
  assign n15215 = ~po57  & n15213;
  assign n15216 = n14695 & ~po7 ;
  assign n15217 = ~n14743 & ~n14744;
  assign n15218 = po7  & n15217;
  assign n15219 = ~n14749 & ~n15218;
  assign n15220 = n14749 & n15218;
  assign n15221 = ~n15219 & ~n15220;
  assign n15222 = ~n14769 & ~n15215;
  assign n15223 = ~n15214 & ~n15222;
  assign n15224 = po58  & ~n15223;
  assign n15225 = ~po58  & n15223;
  assign n15226 = ~n14698 & ~n14699;
  assign n15227 = po7  & n15226;
  assign n15228 = ~n14704 & ~n15227;
  assign n15229 = n14704 & n15227;
  assign n15230 = ~n15228 & ~n15229;
  assign n15231 = ~n15225 & ~n15230;
  assign n15232 = ~n15224 & ~n15231;
  assign n15233 = po59  & ~n15232;
  assign n15234 = ~po59  & n15232;
  assign n15235 = ~n14707 & ~n14708;
  assign n15236 = po7  & n15235;
  assign n15237 = ~n14713 & ~n15236;
  assign n15238 = n14713 & n15236;
  assign n15239 = ~n15237 & ~n15238;
  assign n15240 = ~n15234 & ~n15239;
  assign n15241 = ~n15233 & ~n15240;
  assign n15242 = po60  & ~n15241;
  assign n15243 = ~po60  & n15241;
  assign n15244 = ~n14716 & ~n14717;
  assign n15245 = po7  & n15244;
  assign n15246 = ~n14722 & ~n15245;
  assign n15247 = n14722 & n15245;
  assign n15248 = ~n15246 & ~n15247;
  assign n15249 = ~n15243 & ~n15248;
  assign n15250 = ~n15242 & ~n15249;
  assign n15251 = po61  & ~n15250;
  assign n15252 = ~po61  & n15250;
  assign n15253 = ~n14725 & ~n14726;
  assign n15254 = po7  & n15253;
  assign n15255 = ~n14731 & ~n15254;
  assign n15256 = n14731 & n15254;
  assign n15257 = ~n15255 & ~n15256;
  assign n15258 = ~n15252 & ~n15257;
  assign n15259 = ~n15251 & ~n15258;
  assign n15260 = po62  & ~n15259;
  assign n15261 = ~po62  & n15259;
  assign n15262 = ~n14734 & ~n14735;
  assign n15263 = po7  & n15262;
  assign n15264 = ~n14740 & ~n15263;
  assign n15265 = n14740 & n15263;
  assign n15266 = ~n15264 & ~n15265;
  assign n15267 = ~n15261 & ~n15266;
  assign n15268 = ~n15260 & ~n15267;
  assign n15269 = n15221 & n15268;
  assign n15270 = ~n15221 & ~n15268;
  assign n15271 = n14753 & po7 ;
  assign n15272 = ~n14752 & ~n15271;
  assign n15273 = n15270 & n15272;
  assign n15274 = ~po63  & ~n15273;
  assign n15275 = ~n14695 & po7 ;
  assign n15276 = n14751 & ~n15275;
  assign n15277 = po63  & ~n14753;
  assign n15278 = ~n15276 & n15277;
  assign n15279 = ~n15269 & ~n15278;
  assign n15280 = ~n15274 & n15279;
  assign po6  = n15216 | ~n15280;
  assign n15282 = ~n15214 & ~n15215;
  assign n15283 = po6  & n15282;
  assign n15284 = ~n14769 & ~n15283;
  assign n15285 = n14769 & n15283;
  assign n15286 = ~n15284 & ~n15285;
  assign n15287 = pi12  & po6 ;
  assign n15288 = ~pi10  & ~pi11 ;
  assign n15289 = ~pi12  & n15288;
  assign n15290 = ~n15287 & ~n15289;
  assign n15291 = po7  & ~n15290;
  assign n15292 = ~po7  & n15290;
  assign n15293 = ~pi12  & po6 ;
  assign n15294 = pi13  & ~n15293;
  assign n15295 = ~pi13  & n15293;
  assign n15296 = ~n15294 & ~n15295;
  assign n15297 = ~n15292 & n15296;
  assign n15298 = ~n15291 & ~n15297;
  assign n15299 = po8  & ~n15298;
  assign n15300 = ~po8  & n15298;
  assign n15301 = po7  & n15280;
  assign n15302 = ~n15295 & ~n15301;
  assign n15303 = pi14  & ~n15302;
  assign n15304 = ~pi14  & n15302;
  assign n15305 = ~n15303 & ~n15304;
  assign n15306 = ~n15300 & ~n15305;
  assign n15307 = ~n15299 & ~n15306;
  assign n15308 = po9  & ~n15307;
  assign n15309 = ~po9  & n15307;
  assign n15310 = ~n14774 & ~n14775;
  assign n15311 = po6  & n15310;
  assign n15312 = n14779 & ~n15311;
  assign n15313 = ~n14779 & n15311;
  assign n15314 = ~n15312 & ~n15313;
  assign n15315 = ~n15309 & ~n15314;
  assign n15316 = ~n15308 & ~n15315;
  assign n15317 = po10  & ~n15316;
  assign n15318 = ~po10  & n15316;
  assign n15319 = ~n14782 & ~n14783;
  assign n15320 = po6  & n15319;
  assign n15321 = ~n14788 & ~n15320;
  assign n15322 = n14788 & n15320;
  assign n15323 = ~n15321 & ~n15322;
  assign n15324 = ~n15318 & ~n15323;
  assign n15325 = ~n15317 & ~n15324;
  assign n15326 = po11  & ~n15325;
  assign n15327 = ~po11  & n15325;
  assign n15328 = ~n14791 & ~n14792;
  assign n15329 = po6  & n15328;
  assign n15330 = n14797 & n15329;
  assign n15331 = ~n14797 & ~n15329;
  assign n15332 = ~n15330 & ~n15331;
  assign n15333 = ~n15327 & ~n15332;
  assign n15334 = ~n15326 & ~n15333;
  assign n15335 = po12  & ~n15334;
  assign n15336 = ~po12  & n15334;
  assign n15337 = ~n14800 & ~n14801;
  assign n15338 = po6  & n15337;
  assign n15339 = ~n14806 & ~n15338;
  assign n15340 = n14806 & n15338;
  assign n15341 = ~n15339 & ~n15340;
  assign n15342 = ~n15336 & ~n15341;
  assign n15343 = ~n15335 & ~n15342;
  assign n15344 = po13  & ~n15343;
  assign n15345 = ~po13  & n15343;
  assign n15346 = ~n14809 & ~n14810;
  assign n15347 = po6  & n15346;
  assign n15348 = ~n14815 & ~n15347;
  assign n15349 = n14815 & n15347;
  assign n15350 = ~n15348 & ~n15349;
  assign n15351 = ~n15345 & ~n15350;
  assign n15352 = ~n15344 & ~n15351;
  assign n15353 = po14  & ~n15352;
  assign n15354 = ~po14  & n15352;
  assign n15355 = ~n14818 & ~n14819;
  assign n15356 = po6  & n15355;
  assign n15357 = ~n14824 & ~n15356;
  assign n15358 = n14824 & n15356;
  assign n15359 = ~n15357 & ~n15358;
  assign n15360 = ~n15354 & ~n15359;
  assign n15361 = ~n15353 & ~n15360;
  assign n15362 = po15  & ~n15361;
  assign n15363 = ~po15  & n15361;
  assign n15364 = ~n14827 & ~n14828;
  assign n15365 = po6  & n15364;
  assign n15366 = ~n14833 & ~n15365;
  assign n15367 = n14833 & n15365;
  assign n15368 = ~n15366 & ~n15367;
  assign n15369 = ~n15363 & ~n15368;
  assign n15370 = ~n15362 & ~n15369;
  assign n15371 = po16  & ~n15370;
  assign n15372 = ~po16  & n15370;
  assign n15373 = ~n14836 & ~n14837;
  assign n15374 = po6  & n15373;
  assign n15375 = ~n14842 & ~n15374;
  assign n15376 = n14842 & n15374;
  assign n15377 = ~n15375 & ~n15376;
  assign n15378 = ~n15372 & ~n15377;
  assign n15379 = ~n15371 & ~n15378;
  assign n15380 = po17  & ~n15379;
  assign n15381 = ~po17  & n15379;
  assign n15382 = ~n14845 & ~n14846;
  assign n15383 = po6  & n15382;
  assign n15384 = ~n14851 & ~n15383;
  assign n15385 = n14851 & n15383;
  assign n15386 = ~n15384 & ~n15385;
  assign n15387 = ~n15381 & ~n15386;
  assign n15388 = ~n15380 & ~n15387;
  assign n15389 = po18  & ~n15388;
  assign n15390 = ~po18  & n15388;
  assign n15391 = ~n14854 & ~n14855;
  assign n15392 = po6  & n15391;
  assign n15393 = ~n14860 & ~n15392;
  assign n15394 = n14860 & n15392;
  assign n15395 = ~n15393 & ~n15394;
  assign n15396 = ~n15390 & ~n15395;
  assign n15397 = ~n15389 & ~n15396;
  assign n15398 = po19  & ~n15397;
  assign n15399 = ~po19  & n15397;
  assign n15400 = ~n14863 & ~n14864;
  assign n15401 = po6  & n15400;
  assign n15402 = ~n14869 & ~n15401;
  assign n15403 = n14869 & n15401;
  assign n15404 = ~n15402 & ~n15403;
  assign n15405 = ~n15399 & ~n15404;
  assign n15406 = ~n15398 & ~n15405;
  assign n15407 = po20  & ~n15406;
  assign n15408 = ~po20  & n15406;
  assign n15409 = ~n14872 & ~n14873;
  assign n15410 = po6  & n15409;
  assign n15411 = ~n14878 & ~n15410;
  assign n15412 = n14878 & n15410;
  assign n15413 = ~n15411 & ~n15412;
  assign n15414 = ~n15408 & ~n15413;
  assign n15415 = ~n15407 & ~n15414;
  assign n15416 = po21  & ~n15415;
  assign n15417 = ~po21  & n15415;
  assign n15418 = ~n14881 & ~n14882;
  assign n15419 = po6  & n15418;
  assign n15420 = ~n14887 & ~n15419;
  assign n15421 = n14887 & n15419;
  assign n15422 = ~n15420 & ~n15421;
  assign n15423 = ~n15417 & ~n15422;
  assign n15424 = ~n15416 & ~n15423;
  assign n15425 = po22  & ~n15424;
  assign n15426 = ~po22  & n15424;
  assign n15427 = ~n14890 & ~n14891;
  assign n15428 = po6  & n15427;
  assign n15429 = ~n14896 & ~n15428;
  assign n15430 = n14896 & n15428;
  assign n15431 = ~n15429 & ~n15430;
  assign n15432 = ~n15426 & ~n15431;
  assign n15433 = ~n15425 & ~n15432;
  assign n15434 = po23  & ~n15433;
  assign n15435 = ~po23  & n15433;
  assign n15436 = ~n14899 & ~n14900;
  assign n15437 = po6  & n15436;
  assign n15438 = ~n14905 & ~n15437;
  assign n15439 = n14905 & n15437;
  assign n15440 = ~n15438 & ~n15439;
  assign n15441 = ~n15435 & ~n15440;
  assign n15442 = ~n15434 & ~n15441;
  assign n15443 = po24  & ~n15442;
  assign n15444 = ~po24  & n15442;
  assign n15445 = ~n14908 & ~n14909;
  assign n15446 = po6  & n15445;
  assign n15447 = ~n14914 & ~n15446;
  assign n15448 = n14914 & n15446;
  assign n15449 = ~n15447 & ~n15448;
  assign n15450 = ~n15444 & ~n15449;
  assign n15451 = ~n15443 & ~n15450;
  assign n15452 = po25  & ~n15451;
  assign n15453 = ~po25  & n15451;
  assign n15454 = ~n14917 & ~n14918;
  assign n15455 = po6  & n15454;
  assign n15456 = ~n14923 & ~n15455;
  assign n15457 = n14923 & n15455;
  assign n15458 = ~n15456 & ~n15457;
  assign n15459 = ~n15453 & ~n15458;
  assign n15460 = ~n15452 & ~n15459;
  assign n15461 = po26  & ~n15460;
  assign n15462 = ~po26  & n15460;
  assign n15463 = ~n14926 & ~n14927;
  assign n15464 = po6  & n15463;
  assign n15465 = ~n14932 & ~n15464;
  assign n15466 = n14932 & n15464;
  assign n15467 = ~n15465 & ~n15466;
  assign n15468 = ~n15462 & ~n15467;
  assign n15469 = ~n15461 & ~n15468;
  assign n15470 = po27  & ~n15469;
  assign n15471 = ~po27  & n15469;
  assign n15472 = ~n14935 & ~n14936;
  assign n15473 = po6  & n15472;
  assign n15474 = ~n14941 & ~n15473;
  assign n15475 = n14941 & n15473;
  assign n15476 = ~n15474 & ~n15475;
  assign n15477 = ~n15471 & ~n15476;
  assign n15478 = ~n15470 & ~n15477;
  assign n15479 = po28  & ~n15478;
  assign n15480 = ~po28  & n15478;
  assign n15481 = ~n14944 & ~n14945;
  assign n15482 = po6  & n15481;
  assign n15483 = ~n14950 & ~n15482;
  assign n15484 = n14950 & n15482;
  assign n15485 = ~n15483 & ~n15484;
  assign n15486 = ~n15480 & ~n15485;
  assign n15487 = ~n15479 & ~n15486;
  assign n15488 = po29  & ~n15487;
  assign n15489 = ~po29  & n15487;
  assign n15490 = ~n14953 & ~n14954;
  assign n15491 = po6  & n15490;
  assign n15492 = ~n14959 & ~n15491;
  assign n15493 = n14959 & n15491;
  assign n15494 = ~n15492 & ~n15493;
  assign n15495 = ~n15489 & ~n15494;
  assign n15496 = ~n15488 & ~n15495;
  assign n15497 = po30  & ~n15496;
  assign n15498 = ~po30  & n15496;
  assign n15499 = ~n14962 & ~n14963;
  assign n15500 = po6  & n15499;
  assign n15501 = ~n14968 & ~n15500;
  assign n15502 = n14968 & n15500;
  assign n15503 = ~n15501 & ~n15502;
  assign n15504 = ~n15498 & ~n15503;
  assign n15505 = ~n15497 & ~n15504;
  assign n15506 = po31  & ~n15505;
  assign n15507 = ~po31  & n15505;
  assign n15508 = ~n14971 & ~n14972;
  assign n15509 = po6  & n15508;
  assign n15510 = ~n14977 & ~n15509;
  assign n15511 = n14977 & n15509;
  assign n15512 = ~n15510 & ~n15511;
  assign n15513 = ~n15507 & ~n15512;
  assign n15514 = ~n15506 & ~n15513;
  assign n15515 = po32  & ~n15514;
  assign n15516 = ~po32  & n15514;
  assign n15517 = ~n14980 & ~n14981;
  assign n15518 = po6  & n15517;
  assign n15519 = ~n14986 & ~n15518;
  assign n15520 = n14986 & n15518;
  assign n15521 = ~n15519 & ~n15520;
  assign n15522 = ~n15516 & ~n15521;
  assign n15523 = ~n15515 & ~n15522;
  assign n15524 = po33  & ~n15523;
  assign n15525 = ~po33  & n15523;
  assign n15526 = ~n14989 & ~n14990;
  assign n15527 = po6  & n15526;
  assign n15528 = ~n14995 & ~n15527;
  assign n15529 = n14995 & n15527;
  assign n15530 = ~n15528 & ~n15529;
  assign n15531 = ~n15525 & ~n15530;
  assign n15532 = ~n15524 & ~n15531;
  assign n15533 = po34  & ~n15532;
  assign n15534 = ~po34  & n15532;
  assign n15535 = ~n14998 & ~n14999;
  assign n15536 = po6  & n15535;
  assign n15537 = ~n15004 & ~n15536;
  assign n15538 = n15004 & n15536;
  assign n15539 = ~n15537 & ~n15538;
  assign n15540 = ~n15534 & ~n15539;
  assign n15541 = ~n15533 & ~n15540;
  assign n15542 = po35  & ~n15541;
  assign n15543 = ~po35  & n15541;
  assign n15544 = ~n15007 & ~n15008;
  assign n15545 = po6  & n15544;
  assign n15546 = ~n15013 & ~n15545;
  assign n15547 = n15013 & n15545;
  assign n15548 = ~n15546 & ~n15547;
  assign n15549 = ~n15543 & ~n15548;
  assign n15550 = ~n15542 & ~n15549;
  assign n15551 = po36  & ~n15550;
  assign n15552 = ~po36  & n15550;
  assign n15553 = ~n15016 & ~n15017;
  assign n15554 = po6  & n15553;
  assign n15555 = ~n15022 & ~n15554;
  assign n15556 = n15022 & n15554;
  assign n15557 = ~n15555 & ~n15556;
  assign n15558 = ~n15552 & ~n15557;
  assign n15559 = ~n15551 & ~n15558;
  assign n15560 = po37  & ~n15559;
  assign n15561 = ~po37  & n15559;
  assign n15562 = ~n15025 & ~n15026;
  assign n15563 = po6  & n15562;
  assign n15564 = ~n15031 & ~n15563;
  assign n15565 = n15031 & n15563;
  assign n15566 = ~n15564 & ~n15565;
  assign n15567 = ~n15561 & ~n15566;
  assign n15568 = ~n15560 & ~n15567;
  assign n15569 = po38  & ~n15568;
  assign n15570 = ~po38  & n15568;
  assign n15571 = ~n15034 & ~n15035;
  assign n15572 = po6  & n15571;
  assign n15573 = ~n15040 & ~n15572;
  assign n15574 = n15040 & n15572;
  assign n15575 = ~n15573 & ~n15574;
  assign n15576 = ~n15570 & ~n15575;
  assign n15577 = ~n15569 & ~n15576;
  assign n15578 = po39  & ~n15577;
  assign n15579 = ~po39  & n15577;
  assign n15580 = ~n15043 & ~n15044;
  assign n15581 = po6  & n15580;
  assign n15582 = ~n15049 & ~n15581;
  assign n15583 = n15049 & n15581;
  assign n15584 = ~n15582 & ~n15583;
  assign n15585 = ~n15579 & ~n15584;
  assign n15586 = ~n15578 & ~n15585;
  assign n15587 = po40  & ~n15586;
  assign n15588 = ~po40  & n15586;
  assign n15589 = ~n15052 & ~n15053;
  assign n15590 = po6  & n15589;
  assign n15591 = ~n15058 & ~n15590;
  assign n15592 = n15058 & n15590;
  assign n15593 = ~n15591 & ~n15592;
  assign n15594 = ~n15588 & ~n15593;
  assign n15595 = ~n15587 & ~n15594;
  assign n15596 = po41  & ~n15595;
  assign n15597 = ~po41  & n15595;
  assign n15598 = ~n15061 & ~n15062;
  assign n15599 = po6  & n15598;
  assign n15600 = ~n15067 & ~n15599;
  assign n15601 = n15067 & n15599;
  assign n15602 = ~n15600 & ~n15601;
  assign n15603 = ~n15597 & ~n15602;
  assign n15604 = ~n15596 & ~n15603;
  assign n15605 = po42  & ~n15604;
  assign n15606 = ~po42  & n15604;
  assign n15607 = ~n15070 & ~n15071;
  assign n15608 = po6  & n15607;
  assign n15609 = ~n15076 & ~n15608;
  assign n15610 = n15076 & n15608;
  assign n15611 = ~n15609 & ~n15610;
  assign n15612 = ~n15606 & ~n15611;
  assign n15613 = ~n15605 & ~n15612;
  assign n15614 = po43  & ~n15613;
  assign n15615 = ~po43  & n15613;
  assign n15616 = ~n15079 & ~n15080;
  assign n15617 = po6  & n15616;
  assign n15618 = ~n15085 & ~n15617;
  assign n15619 = n15085 & n15617;
  assign n15620 = ~n15618 & ~n15619;
  assign n15621 = ~n15615 & ~n15620;
  assign n15622 = ~n15614 & ~n15621;
  assign n15623 = po44  & ~n15622;
  assign n15624 = ~po44  & n15622;
  assign n15625 = ~n15088 & ~n15089;
  assign n15626 = po6  & n15625;
  assign n15627 = ~n15094 & ~n15626;
  assign n15628 = n15094 & n15626;
  assign n15629 = ~n15627 & ~n15628;
  assign n15630 = ~n15624 & ~n15629;
  assign n15631 = ~n15623 & ~n15630;
  assign n15632 = po45  & ~n15631;
  assign n15633 = ~po45  & n15631;
  assign n15634 = ~n15097 & ~n15098;
  assign n15635 = po6  & n15634;
  assign n15636 = ~n15103 & ~n15635;
  assign n15637 = n15103 & n15635;
  assign n15638 = ~n15636 & ~n15637;
  assign n15639 = ~n15633 & ~n15638;
  assign n15640 = ~n15632 & ~n15639;
  assign n15641 = po46  & ~n15640;
  assign n15642 = ~po46  & n15640;
  assign n15643 = ~n15106 & ~n15107;
  assign n15644 = po6  & n15643;
  assign n15645 = ~n15112 & ~n15644;
  assign n15646 = n15112 & n15644;
  assign n15647 = ~n15645 & ~n15646;
  assign n15648 = ~n15642 & ~n15647;
  assign n15649 = ~n15641 & ~n15648;
  assign n15650 = po47  & ~n15649;
  assign n15651 = ~po47  & n15649;
  assign n15652 = ~n15115 & ~n15116;
  assign n15653 = po6  & n15652;
  assign n15654 = ~n15121 & ~n15653;
  assign n15655 = n15121 & n15653;
  assign n15656 = ~n15654 & ~n15655;
  assign n15657 = ~n15651 & ~n15656;
  assign n15658 = ~n15650 & ~n15657;
  assign n15659 = po48  & ~n15658;
  assign n15660 = ~po48  & n15658;
  assign n15661 = ~n15124 & ~n15125;
  assign n15662 = po6  & n15661;
  assign n15663 = ~n15130 & ~n15662;
  assign n15664 = n15130 & n15662;
  assign n15665 = ~n15663 & ~n15664;
  assign n15666 = ~n15660 & ~n15665;
  assign n15667 = ~n15659 & ~n15666;
  assign n15668 = po49  & ~n15667;
  assign n15669 = ~po49  & n15667;
  assign n15670 = ~n15133 & ~n15134;
  assign n15671 = po6  & n15670;
  assign n15672 = ~n15139 & ~n15671;
  assign n15673 = n15139 & n15671;
  assign n15674 = ~n15672 & ~n15673;
  assign n15675 = ~n15669 & ~n15674;
  assign n15676 = ~n15668 & ~n15675;
  assign n15677 = po50  & ~n15676;
  assign n15678 = ~po50  & n15676;
  assign n15679 = ~n15142 & ~n15143;
  assign n15680 = po6  & n15679;
  assign n15681 = ~n15148 & ~n15680;
  assign n15682 = n15148 & n15680;
  assign n15683 = ~n15681 & ~n15682;
  assign n15684 = ~n15678 & ~n15683;
  assign n15685 = ~n15677 & ~n15684;
  assign n15686 = po51  & ~n15685;
  assign n15687 = ~po51  & n15685;
  assign n15688 = ~n15151 & ~n15152;
  assign n15689 = po6  & n15688;
  assign n15690 = ~n15157 & ~n15689;
  assign n15691 = n15157 & n15689;
  assign n15692 = ~n15690 & ~n15691;
  assign n15693 = ~n15687 & ~n15692;
  assign n15694 = ~n15686 & ~n15693;
  assign n15695 = po52  & ~n15694;
  assign n15696 = ~po52  & n15694;
  assign n15697 = ~n15160 & ~n15161;
  assign n15698 = po6  & n15697;
  assign n15699 = ~n15166 & ~n15698;
  assign n15700 = n15166 & n15698;
  assign n15701 = ~n15699 & ~n15700;
  assign n15702 = ~n15696 & ~n15701;
  assign n15703 = ~n15695 & ~n15702;
  assign n15704 = po53  & ~n15703;
  assign n15705 = ~po53  & n15703;
  assign n15706 = ~n15169 & ~n15170;
  assign n15707 = po6  & n15706;
  assign n15708 = ~n15175 & ~n15707;
  assign n15709 = n15175 & n15707;
  assign n15710 = ~n15708 & ~n15709;
  assign n15711 = ~n15705 & ~n15710;
  assign n15712 = ~n15704 & ~n15711;
  assign n15713 = po54  & ~n15712;
  assign n15714 = ~po54  & n15712;
  assign n15715 = ~n15178 & ~n15179;
  assign n15716 = po6  & n15715;
  assign n15717 = ~n15184 & ~n15716;
  assign n15718 = n15184 & n15716;
  assign n15719 = ~n15717 & ~n15718;
  assign n15720 = ~n15714 & ~n15719;
  assign n15721 = ~n15713 & ~n15720;
  assign n15722 = po55  & ~n15721;
  assign n15723 = ~po55  & n15721;
  assign n15724 = ~n15187 & ~n15188;
  assign n15725 = po6  & n15724;
  assign n15726 = ~n15193 & ~n15725;
  assign n15727 = n15193 & n15725;
  assign n15728 = ~n15726 & ~n15727;
  assign n15729 = ~n15723 & ~n15728;
  assign n15730 = ~n15722 & ~n15729;
  assign n15731 = po56  & ~n15730;
  assign n15732 = ~po56  & n15730;
  assign n15733 = ~n15196 & ~n15197;
  assign n15734 = po6  & n15733;
  assign n15735 = ~n15202 & ~n15734;
  assign n15736 = n15202 & n15734;
  assign n15737 = ~n15735 & ~n15736;
  assign n15738 = ~n15732 & ~n15737;
  assign n15739 = ~n15731 & ~n15738;
  assign n15740 = po57  & ~n15739;
  assign n15741 = ~n15205 & ~n15211;
  assign n15742 = po6  & n15741;
  assign n15743 = ~n15210 & ~n15742;
  assign n15744 = n15210 & n15742;
  assign n15745 = ~n15743 & ~n15744;
  assign n15746 = ~po57  & n15739;
  assign n15747 = ~n15745 & ~n15746;
  assign n15748 = ~n15740 & ~n15747;
  assign n15749 = po58  & ~n15748;
  assign n15750 = ~po58  & n15748;
  assign n15751 = ~n15260 & ~n15261;
  assign n15752 = po6  & n15751;
  assign n15753 = ~n15266 & ~n15752;
  assign n15754 = n15266 & n15752;
  assign n15755 = ~n15753 & ~n15754;
  assign n15756 = ~n15286 & ~n15750;
  assign n15757 = ~n15749 & ~n15756;
  assign n15758 = po59  & ~n15757;
  assign n15759 = ~po59  & n15757;
  assign n15760 = ~n15224 & ~n15225;
  assign n15761 = po6  & n15760;
  assign n15762 = ~n15230 & ~n15761;
  assign n15763 = n15230 & n15761;
  assign n15764 = ~n15762 & ~n15763;
  assign n15765 = ~n15759 & ~n15764;
  assign n15766 = ~n15758 & ~n15765;
  assign n15767 = po60  & ~n15766;
  assign n15768 = ~po60  & n15766;
  assign n15769 = ~n15233 & ~n15234;
  assign n15770 = po6  & n15769;
  assign n15771 = ~n15239 & ~n15770;
  assign n15772 = n15239 & n15770;
  assign n15773 = ~n15771 & ~n15772;
  assign n15774 = ~n15768 & ~n15773;
  assign n15775 = ~n15767 & ~n15774;
  assign n15776 = po61  & ~n15775;
  assign n15777 = ~po61  & n15775;
  assign n15778 = ~n15242 & ~n15243;
  assign n15779 = po6  & n15778;
  assign n15780 = ~n15248 & ~n15779;
  assign n15781 = n15248 & n15779;
  assign n15782 = ~n15780 & ~n15781;
  assign n15783 = ~n15777 & ~n15782;
  assign n15784 = ~n15776 & ~n15783;
  assign n15785 = po62  & ~n15784;
  assign n15786 = ~po62  & n15784;
  assign n15787 = ~n15251 & ~n15252;
  assign n15788 = po6  & n15787;
  assign n15789 = ~n15257 & ~n15788;
  assign n15790 = n15257 & n15788;
  assign n15791 = ~n15789 & ~n15790;
  assign n15792 = ~n15786 & ~n15791;
  assign n15793 = ~n15785 & ~n15792;
  assign n15794 = n15755 & n15793;
  assign n15795 = ~n15755 & ~n15793;
  assign n15796 = n15270 & po6 ;
  assign n15797 = ~n15269 & ~n15796;
  assign n15798 = n15795 & n15797;
  assign n15799 = ~po63  & ~n15798;
  assign n15800 = ~n15221 & po6 ;
  assign n15801 = n15268 & ~n15800;
  assign n15802 = po63  & ~n15270;
  assign n15803 = ~n15801 & n15802;
  assign n15804 = ~n15799 & ~n15803;
  assign po5  = n15794 | ~n15804;
  assign n15806 = ~n15749 & ~n15750;
  assign n15807 = po5  & n15806;
  assign n15808 = ~n15286 & ~n15807;
  assign n15809 = n15286 & n15807;
  assign n15810 = ~n15808 & ~n15809;
  assign n15811 = pi10  & po5 ;
  assign n15812 = ~pi8  & ~pi9 ;
  assign n15813 = ~pi10  & n15812;
  assign n15814 = ~n15811 & ~n15813;
  assign n15815 = po6  & ~n15814;
  assign n15816 = ~po6  & n15814;
  assign n15817 = ~pi10  & po5 ;
  assign n15818 = pi11  & ~n15817;
  assign n15819 = ~pi11  & n15817;
  assign n15820 = ~n15818 & ~n15819;
  assign n15821 = ~n15816 & n15820;
  assign n15822 = ~n15815 & ~n15821;
  assign n15823 = po7  & ~n15822;
  assign n15824 = ~po7  & n15822;
  assign n15825 = po6  & ~po5 ;
  assign n15826 = ~n15819 & ~n15825;
  assign n15827 = pi12  & ~n15826;
  assign n15828 = ~pi12  & n15826;
  assign n15829 = ~n15827 & ~n15828;
  assign n15830 = ~n15824 & ~n15829;
  assign n15831 = ~n15823 & ~n15830;
  assign n15832 = po8  & ~n15831;
  assign n15833 = ~po8  & n15831;
  assign n15834 = ~n15291 & ~n15292;
  assign n15835 = po5  & n15834;
  assign n15836 = n15296 & ~n15835;
  assign n15837 = ~n15296 & n15835;
  assign n15838 = ~n15836 & ~n15837;
  assign n15839 = ~n15833 & ~n15838;
  assign n15840 = ~n15832 & ~n15839;
  assign n15841 = po9  & ~n15840;
  assign n15842 = ~po9  & n15840;
  assign n15843 = ~n15299 & ~n15300;
  assign n15844 = po5  & n15843;
  assign n15845 = ~n15305 & ~n15844;
  assign n15846 = n15305 & n15844;
  assign n15847 = ~n15845 & ~n15846;
  assign n15848 = ~n15842 & ~n15847;
  assign n15849 = ~n15841 & ~n15848;
  assign n15850 = po10  & ~n15849;
  assign n15851 = ~po10  & n15849;
  assign n15852 = ~n15308 & ~n15309;
  assign n15853 = po5  & n15852;
  assign n15854 = n15314 & n15853;
  assign n15855 = ~n15314 & ~n15853;
  assign n15856 = ~n15854 & ~n15855;
  assign n15857 = ~n15851 & ~n15856;
  assign n15858 = ~n15850 & ~n15857;
  assign n15859 = po11  & ~n15858;
  assign n15860 = ~po11  & n15858;
  assign n15861 = ~n15317 & ~n15318;
  assign n15862 = po5  & n15861;
  assign n15863 = ~n15323 & ~n15862;
  assign n15864 = n15323 & n15862;
  assign n15865 = ~n15863 & ~n15864;
  assign n15866 = ~n15860 & ~n15865;
  assign n15867 = ~n15859 & ~n15866;
  assign n15868 = po12  & ~n15867;
  assign n15869 = ~po12  & n15867;
  assign n15870 = ~n15326 & ~n15327;
  assign n15871 = po5  & n15870;
  assign n15872 = ~n15332 & ~n15871;
  assign n15873 = n15332 & n15871;
  assign n15874 = ~n15872 & ~n15873;
  assign n15875 = ~n15869 & ~n15874;
  assign n15876 = ~n15868 & ~n15875;
  assign n15877 = po13  & ~n15876;
  assign n15878 = ~po13  & n15876;
  assign n15879 = ~n15335 & ~n15336;
  assign n15880 = po5  & n15879;
  assign n15881 = ~n15341 & ~n15880;
  assign n15882 = n15341 & n15880;
  assign n15883 = ~n15881 & ~n15882;
  assign n15884 = ~n15878 & ~n15883;
  assign n15885 = ~n15877 & ~n15884;
  assign n15886 = po14  & ~n15885;
  assign n15887 = ~po14  & n15885;
  assign n15888 = ~n15344 & ~n15345;
  assign n15889 = po5  & n15888;
  assign n15890 = ~n15350 & ~n15889;
  assign n15891 = n15350 & n15889;
  assign n15892 = ~n15890 & ~n15891;
  assign n15893 = ~n15887 & ~n15892;
  assign n15894 = ~n15886 & ~n15893;
  assign n15895 = po15  & ~n15894;
  assign n15896 = ~po15  & n15894;
  assign n15897 = ~n15353 & ~n15354;
  assign n15898 = po5  & n15897;
  assign n15899 = ~n15359 & ~n15898;
  assign n15900 = n15359 & n15898;
  assign n15901 = ~n15899 & ~n15900;
  assign n15902 = ~n15896 & ~n15901;
  assign n15903 = ~n15895 & ~n15902;
  assign n15904 = po16  & ~n15903;
  assign n15905 = ~po16  & n15903;
  assign n15906 = ~n15362 & ~n15363;
  assign n15907 = po5  & n15906;
  assign n15908 = ~n15368 & ~n15907;
  assign n15909 = n15368 & n15907;
  assign n15910 = ~n15908 & ~n15909;
  assign n15911 = ~n15905 & ~n15910;
  assign n15912 = ~n15904 & ~n15911;
  assign n15913 = po17  & ~n15912;
  assign n15914 = ~po17  & n15912;
  assign n15915 = ~n15371 & ~n15372;
  assign n15916 = po5  & n15915;
  assign n15917 = ~n15377 & ~n15916;
  assign n15918 = n15377 & n15916;
  assign n15919 = ~n15917 & ~n15918;
  assign n15920 = ~n15914 & ~n15919;
  assign n15921 = ~n15913 & ~n15920;
  assign n15922 = po18  & ~n15921;
  assign n15923 = ~po18  & n15921;
  assign n15924 = ~n15380 & ~n15381;
  assign n15925 = po5  & n15924;
  assign n15926 = ~n15386 & ~n15925;
  assign n15927 = n15386 & n15925;
  assign n15928 = ~n15926 & ~n15927;
  assign n15929 = ~n15923 & ~n15928;
  assign n15930 = ~n15922 & ~n15929;
  assign n15931 = po19  & ~n15930;
  assign n15932 = ~po19  & n15930;
  assign n15933 = ~n15389 & ~n15390;
  assign n15934 = po5  & n15933;
  assign n15935 = ~n15395 & ~n15934;
  assign n15936 = n15395 & n15934;
  assign n15937 = ~n15935 & ~n15936;
  assign n15938 = ~n15932 & ~n15937;
  assign n15939 = ~n15931 & ~n15938;
  assign n15940 = po20  & ~n15939;
  assign n15941 = ~po20  & n15939;
  assign n15942 = ~n15398 & ~n15399;
  assign n15943 = po5  & n15942;
  assign n15944 = ~n15404 & ~n15943;
  assign n15945 = n15404 & n15943;
  assign n15946 = ~n15944 & ~n15945;
  assign n15947 = ~n15941 & ~n15946;
  assign n15948 = ~n15940 & ~n15947;
  assign n15949 = po21  & ~n15948;
  assign n15950 = ~po21  & n15948;
  assign n15951 = ~n15407 & ~n15408;
  assign n15952 = po5  & n15951;
  assign n15953 = ~n15413 & ~n15952;
  assign n15954 = n15413 & n15952;
  assign n15955 = ~n15953 & ~n15954;
  assign n15956 = ~n15950 & ~n15955;
  assign n15957 = ~n15949 & ~n15956;
  assign n15958 = po22  & ~n15957;
  assign n15959 = ~po22  & n15957;
  assign n15960 = ~n15416 & ~n15417;
  assign n15961 = po5  & n15960;
  assign n15962 = ~n15422 & ~n15961;
  assign n15963 = n15422 & n15961;
  assign n15964 = ~n15962 & ~n15963;
  assign n15965 = ~n15959 & ~n15964;
  assign n15966 = ~n15958 & ~n15965;
  assign n15967 = po23  & ~n15966;
  assign n15968 = ~po23  & n15966;
  assign n15969 = ~n15425 & ~n15426;
  assign n15970 = po5  & n15969;
  assign n15971 = ~n15431 & ~n15970;
  assign n15972 = n15431 & n15970;
  assign n15973 = ~n15971 & ~n15972;
  assign n15974 = ~n15968 & ~n15973;
  assign n15975 = ~n15967 & ~n15974;
  assign n15976 = po24  & ~n15975;
  assign n15977 = ~po24  & n15975;
  assign n15978 = ~n15434 & ~n15435;
  assign n15979 = po5  & n15978;
  assign n15980 = ~n15440 & ~n15979;
  assign n15981 = n15440 & n15979;
  assign n15982 = ~n15980 & ~n15981;
  assign n15983 = ~n15977 & ~n15982;
  assign n15984 = ~n15976 & ~n15983;
  assign n15985 = po25  & ~n15984;
  assign n15986 = ~po25  & n15984;
  assign n15987 = ~n15443 & ~n15444;
  assign n15988 = po5  & n15987;
  assign n15989 = ~n15449 & ~n15988;
  assign n15990 = n15449 & n15988;
  assign n15991 = ~n15989 & ~n15990;
  assign n15992 = ~n15986 & ~n15991;
  assign n15993 = ~n15985 & ~n15992;
  assign n15994 = po26  & ~n15993;
  assign n15995 = ~po26  & n15993;
  assign n15996 = ~n15452 & ~n15453;
  assign n15997 = po5  & n15996;
  assign n15998 = ~n15458 & ~n15997;
  assign n15999 = n15458 & n15997;
  assign n16000 = ~n15998 & ~n15999;
  assign n16001 = ~n15995 & ~n16000;
  assign n16002 = ~n15994 & ~n16001;
  assign n16003 = po27  & ~n16002;
  assign n16004 = ~po27  & n16002;
  assign n16005 = ~n15461 & ~n15462;
  assign n16006 = po5  & n16005;
  assign n16007 = ~n15467 & ~n16006;
  assign n16008 = n15467 & n16006;
  assign n16009 = ~n16007 & ~n16008;
  assign n16010 = ~n16004 & ~n16009;
  assign n16011 = ~n16003 & ~n16010;
  assign n16012 = po28  & ~n16011;
  assign n16013 = ~po28  & n16011;
  assign n16014 = ~n15470 & ~n15471;
  assign n16015 = po5  & n16014;
  assign n16016 = ~n15476 & ~n16015;
  assign n16017 = n15476 & n16015;
  assign n16018 = ~n16016 & ~n16017;
  assign n16019 = ~n16013 & ~n16018;
  assign n16020 = ~n16012 & ~n16019;
  assign n16021 = po29  & ~n16020;
  assign n16022 = ~po29  & n16020;
  assign n16023 = ~n15479 & ~n15480;
  assign n16024 = po5  & n16023;
  assign n16025 = ~n15485 & ~n16024;
  assign n16026 = n15485 & n16024;
  assign n16027 = ~n16025 & ~n16026;
  assign n16028 = ~n16022 & ~n16027;
  assign n16029 = ~n16021 & ~n16028;
  assign n16030 = po30  & ~n16029;
  assign n16031 = ~po30  & n16029;
  assign n16032 = ~n15488 & ~n15489;
  assign n16033 = po5  & n16032;
  assign n16034 = ~n15494 & ~n16033;
  assign n16035 = n15494 & n16033;
  assign n16036 = ~n16034 & ~n16035;
  assign n16037 = ~n16031 & ~n16036;
  assign n16038 = ~n16030 & ~n16037;
  assign n16039 = po31  & ~n16038;
  assign n16040 = ~po31  & n16038;
  assign n16041 = ~n15497 & ~n15498;
  assign n16042 = po5  & n16041;
  assign n16043 = ~n15503 & ~n16042;
  assign n16044 = n15503 & n16042;
  assign n16045 = ~n16043 & ~n16044;
  assign n16046 = ~n16040 & ~n16045;
  assign n16047 = ~n16039 & ~n16046;
  assign n16048 = po32  & ~n16047;
  assign n16049 = ~po32  & n16047;
  assign n16050 = ~n15506 & ~n15507;
  assign n16051 = po5  & n16050;
  assign n16052 = ~n15512 & ~n16051;
  assign n16053 = n15512 & n16051;
  assign n16054 = ~n16052 & ~n16053;
  assign n16055 = ~n16049 & ~n16054;
  assign n16056 = ~n16048 & ~n16055;
  assign n16057 = po33  & ~n16056;
  assign n16058 = ~po33  & n16056;
  assign n16059 = ~n15515 & ~n15516;
  assign n16060 = po5  & n16059;
  assign n16061 = ~n15521 & ~n16060;
  assign n16062 = n15521 & n16060;
  assign n16063 = ~n16061 & ~n16062;
  assign n16064 = ~n16058 & ~n16063;
  assign n16065 = ~n16057 & ~n16064;
  assign n16066 = po34  & ~n16065;
  assign n16067 = ~po34  & n16065;
  assign n16068 = ~n15524 & ~n15525;
  assign n16069 = po5  & n16068;
  assign n16070 = ~n15530 & ~n16069;
  assign n16071 = n15530 & n16069;
  assign n16072 = ~n16070 & ~n16071;
  assign n16073 = ~n16067 & ~n16072;
  assign n16074 = ~n16066 & ~n16073;
  assign n16075 = po35  & ~n16074;
  assign n16076 = ~po35  & n16074;
  assign n16077 = ~n15533 & ~n15534;
  assign n16078 = po5  & n16077;
  assign n16079 = ~n15539 & ~n16078;
  assign n16080 = n15539 & n16078;
  assign n16081 = ~n16079 & ~n16080;
  assign n16082 = ~n16076 & ~n16081;
  assign n16083 = ~n16075 & ~n16082;
  assign n16084 = po36  & ~n16083;
  assign n16085 = ~po36  & n16083;
  assign n16086 = ~n15542 & ~n15543;
  assign n16087 = po5  & n16086;
  assign n16088 = ~n15548 & ~n16087;
  assign n16089 = n15548 & n16087;
  assign n16090 = ~n16088 & ~n16089;
  assign n16091 = ~n16085 & ~n16090;
  assign n16092 = ~n16084 & ~n16091;
  assign n16093 = po37  & ~n16092;
  assign n16094 = ~po37  & n16092;
  assign n16095 = ~n15551 & ~n15552;
  assign n16096 = po5  & n16095;
  assign n16097 = ~n15557 & ~n16096;
  assign n16098 = n15557 & n16096;
  assign n16099 = ~n16097 & ~n16098;
  assign n16100 = ~n16094 & ~n16099;
  assign n16101 = ~n16093 & ~n16100;
  assign n16102 = po38  & ~n16101;
  assign n16103 = ~po38  & n16101;
  assign n16104 = ~n15560 & ~n15561;
  assign n16105 = po5  & n16104;
  assign n16106 = ~n15566 & ~n16105;
  assign n16107 = n15566 & n16105;
  assign n16108 = ~n16106 & ~n16107;
  assign n16109 = ~n16103 & ~n16108;
  assign n16110 = ~n16102 & ~n16109;
  assign n16111 = po39  & ~n16110;
  assign n16112 = ~po39  & n16110;
  assign n16113 = ~n15569 & ~n15570;
  assign n16114 = po5  & n16113;
  assign n16115 = ~n15575 & ~n16114;
  assign n16116 = n15575 & n16114;
  assign n16117 = ~n16115 & ~n16116;
  assign n16118 = ~n16112 & ~n16117;
  assign n16119 = ~n16111 & ~n16118;
  assign n16120 = po40  & ~n16119;
  assign n16121 = ~po40  & n16119;
  assign n16122 = ~n15578 & ~n15579;
  assign n16123 = po5  & n16122;
  assign n16124 = ~n15584 & ~n16123;
  assign n16125 = n15584 & n16123;
  assign n16126 = ~n16124 & ~n16125;
  assign n16127 = ~n16121 & ~n16126;
  assign n16128 = ~n16120 & ~n16127;
  assign n16129 = po41  & ~n16128;
  assign n16130 = ~po41  & n16128;
  assign n16131 = ~n15587 & ~n15588;
  assign n16132 = po5  & n16131;
  assign n16133 = ~n15593 & ~n16132;
  assign n16134 = n15593 & n16132;
  assign n16135 = ~n16133 & ~n16134;
  assign n16136 = ~n16130 & ~n16135;
  assign n16137 = ~n16129 & ~n16136;
  assign n16138 = po42  & ~n16137;
  assign n16139 = ~po42  & n16137;
  assign n16140 = ~n15596 & ~n15597;
  assign n16141 = po5  & n16140;
  assign n16142 = ~n15602 & ~n16141;
  assign n16143 = n15602 & n16141;
  assign n16144 = ~n16142 & ~n16143;
  assign n16145 = ~n16139 & ~n16144;
  assign n16146 = ~n16138 & ~n16145;
  assign n16147 = po43  & ~n16146;
  assign n16148 = ~po43  & n16146;
  assign n16149 = ~n15605 & ~n15606;
  assign n16150 = po5  & n16149;
  assign n16151 = ~n15611 & ~n16150;
  assign n16152 = n15611 & n16150;
  assign n16153 = ~n16151 & ~n16152;
  assign n16154 = ~n16148 & ~n16153;
  assign n16155 = ~n16147 & ~n16154;
  assign n16156 = po44  & ~n16155;
  assign n16157 = ~po44  & n16155;
  assign n16158 = ~n15614 & ~n15615;
  assign n16159 = po5  & n16158;
  assign n16160 = ~n15620 & ~n16159;
  assign n16161 = n15620 & n16159;
  assign n16162 = ~n16160 & ~n16161;
  assign n16163 = ~n16157 & ~n16162;
  assign n16164 = ~n16156 & ~n16163;
  assign n16165 = po45  & ~n16164;
  assign n16166 = ~po45  & n16164;
  assign n16167 = ~n15623 & ~n15624;
  assign n16168 = po5  & n16167;
  assign n16169 = ~n15629 & ~n16168;
  assign n16170 = n15629 & n16168;
  assign n16171 = ~n16169 & ~n16170;
  assign n16172 = ~n16166 & ~n16171;
  assign n16173 = ~n16165 & ~n16172;
  assign n16174 = po46  & ~n16173;
  assign n16175 = ~po46  & n16173;
  assign n16176 = ~n15632 & ~n15633;
  assign n16177 = po5  & n16176;
  assign n16178 = ~n15638 & ~n16177;
  assign n16179 = n15638 & n16177;
  assign n16180 = ~n16178 & ~n16179;
  assign n16181 = ~n16175 & ~n16180;
  assign n16182 = ~n16174 & ~n16181;
  assign n16183 = po47  & ~n16182;
  assign n16184 = ~po47  & n16182;
  assign n16185 = ~n15641 & ~n15642;
  assign n16186 = po5  & n16185;
  assign n16187 = ~n15647 & ~n16186;
  assign n16188 = n15647 & n16186;
  assign n16189 = ~n16187 & ~n16188;
  assign n16190 = ~n16184 & ~n16189;
  assign n16191 = ~n16183 & ~n16190;
  assign n16192 = po48  & ~n16191;
  assign n16193 = ~po48  & n16191;
  assign n16194 = ~n15650 & ~n15651;
  assign n16195 = po5  & n16194;
  assign n16196 = ~n15656 & ~n16195;
  assign n16197 = n15656 & n16195;
  assign n16198 = ~n16196 & ~n16197;
  assign n16199 = ~n16193 & ~n16198;
  assign n16200 = ~n16192 & ~n16199;
  assign n16201 = po49  & ~n16200;
  assign n16202 = ~po49  & n16200;
  assign n16203 = ~n15659 & ~n15660;
  assign n16204 = po5  & n16203;
  assign n16205 = ~n15665 & ~n16204;
  assign n16206 = n15665 & n16204;
  assign n16207 = ~n16205 & ~n16206;
  assign n16208 = ~n16202 & ~n16207;
  assign n16209 = ~n16201 & ~n16208;
  assign n16210 = po50  & ~n16209;
  assign n16211 = ~po50  & n16209;
  assign n16212 = ~n15668 & ~n15669;
  assign n16213 = po5  & n16212;
  assign n16214 = ~n15674 & ~n16213;
  assign n16215 = n15674 & n16213;
  assign n16216 = ~n16214 & ~n16215;
  assign n16217 = ~n16211 & ~n16216;
  assign n16218 = ~n16210 & ~n16217;
  assign n16219 = po51  & ~n16218;
  assign n16220 = ~po51  & n16218;
  assign n16221 = ~n15677 & ~n15678;
  assign n16222 = po5  & n16221;
  assign n16223 = ~n15683 & ~n16222;
  assign n16224 = n15683 & n16222;
  assign n16225 = ~n16223 & ~n16224;
  assign n16226 = ~n16220 & ~n16225;
  assign n16227 = ~n16219 & ~n16226;
  assign n16228 = po52  & ~n16227;
  assign n16229 = ~po52  & n16227;
  assign n16230 = ~n15686 & ~n15687;
  assign n16231 = po5  & n16230;
  assign n16232 = ~n15692 & ~n16231;
  assign n16233 = n15692 & n16231;
  assign n16234 = ~n16232 & ~n16233;
  assign n16235 = ~n16229 & ~n16234;
  assign n16236 = ~n16228 & ~n16235;
  assign n16237 = po53  & ~n16236;
  assign n16238 = ~po53  & n16236;
  assign n16239 = ~n15695 & ~n15696;
  assign n16240 = po5  & n16239;
  assign n16241 = ~n15701 & ~n16240;
  assign n16242 = n15701 & n16240;
  assign n16243 = ~n16241 & ~n16242;
  assign n16244 = ~n16238 & ~n16243;
  assign n16245 = ~n16237 & ~n16244;
  assign n16246 = po54  & ~n16245;
  assign n16247 = ~po54  & n16245;
  assign n16248 = ~n15704 & ~n15705;
  assign n16249 = po5  & n16248;
  assign n16250 = ~n15710 & ~n16249;
  assign n16251 = n15710 & n16249;
  assign n16252 = ~n16250 & ~n16251;
  assign n16253 = ~n16247 & ~n16252;
  assign n16254 = ~n16246 & ~n16253;
  assign n16255 = po55  & ~n16254;
  assign n16256 = ~po55  & n16254;
  assign n16257 = ~n15713 & ~n15714;
  assign n16258 = po5  & n16257;
  assign n16259 = ~n15719 & ~n16258;
  assign n16260 = n15719 & n16258;
  assign n16261 = ~n16259 & ~n16260;
  assign n16262 = ~n16256 & ~n16261;
  assign n16263 = ~n16255 & ~n16262;
  assign n16264 = po56  & ~n16263;
  assign n16265 = ~po56  & n16263;
  assign n16266 = ~n15722 & ~n15723;
  assign n16267 = po5  & n16266;
  assign n16268 = ~n15728 & ~n16267;
  assign n16269 = n15728 & n16267;
  assign n16270 = ~n16268 & ~n16269;
  assign n16271 = ~n16265 & ~n16270;
  assign n16272 = ~n16264 & ~n16271;
  assign n16273 = po57  & ~n16272;
  assign n16274 = ~po57  & n16272;
  assign n16275 = ~n15731 & ~n15732;
  assign n16276 = po5  & n16275;
  assign n16277 = ~n15737 & ~n16276;
  assign n16278 = n15737 & n16276;
  assign n16279 = ~n16277 & ~n16278;
  assign n16280 = ~n16274 & ~n16279;
  assign n16281 = ~n16273 & ~n16280;
  assign n16282 = po58  & ~n16281;
  assign n16283 = ~n15740 & ~n15746;
  assign n16284 = po5  & n16283;
  assign n16285 = ~n15745 & ~n16284;
  assign n16286 = n15745 & n16284;
  assign n16287 = ~n16285 & ~n16286;
  assign n16288 = ~po58  & n16281;
  assign n16289 = ~n16287 & ~n16288;
  assign n16290 = ~n16282 & ~n16289;
  assign n16291 = po59  & ~n16290;
  assign n16292 = ~po59  & n16290;
  assign n16293 = ~n15785 & ~n15786;
  assign n16294 = po5  & n16293;
  assign n16295 = ~n15791 & ~n16294;
  assign n16296 = n15791 & n16294;
  assign n16297 = ~n16295 & ~n16296;
  assign n16298 = ~n15810 & ~n16292;
  assign n16299 = ~n16291 & ~n16298;
  assign n16300 = po60  & ~n16299;
  assign n16301 = ~po60  & n16299;
  assign n16302 = ~n15758 & ~n15759;
  assign n16303 = po5  & n16302;
  assign n16304 = ~n15764 & ~n16303;
  assign n16305 = n15764 & n16303;
  assign n16306 = ~n16304 & ~n16305;
  assign n16307 = ~n16301 & ~n16306;
  assign n16308 = ~n16300 & ~n16307;
  assign n16309 = po61  & ~n16308;
  assign n16310 = ~po61  & n16308;
  assign n16311 = ~n15767 & ~n15768;
  assign n16312 = po5  & n16311;
  assign n16313 = ~n15773 & ~n16312;
  assign n16314 = n15773 & n16312;
  assign n16315 = ~n16313 & ~n16314;
  assign n16316 = ~n16310 & ~n16315;
  assign n16317 = ~n16309 & ~n16316;
  assign n16318 = po62  & ~n16317;
  assign n16319 = ~po62  & n16317;
  assign n16320 = ~n15776 & ~n15777;
  assign n16321 = po5  & n16320;
  assign n16322 = ~n15782 & ~n16321;
  assign n16323 = n15782 & n16321;
  assign n16324 = ~n16322 & ~n16323;
  assign n16325 = ~n16319 & ~n16324;
  assign n16326 = ~n16318 & ~n16325;
  assign n16327 = n16297 & n16326;
  assign n16328 = ~n16297 & ~n16326;
  assign n16329 = n15795 & ~n15804;
  assign n16330 = ~n15794 & ~n16329;
  assign n16331 = n16328 & n16330;
  assign n16332 = ~po63  & ~n16331;
  assign n16333 = ~n15755 & ~n15804;
  assign n16334 = n15793 & ~n16333;
  assign n16335 = po63  & ~n15795;
  assign n16336 = ~n16334 & n16335;
  assign n16337 = ~n16332 & ~n16336;
  assign po4  = n16327 | ~n16337;
  assign n16339 = ~n16291 & ~n16292;
  assign n16340 = po4  & n16339;
  assign n16341 = ~n15810 & ~n16340;
  assign n16342 = n15810 & n16340;
  assign n16343 = ~n16341 & ~n16342;
  assign n16344 = pi8  & po4 ;
  assign n16345 = ~pi6  & ~pi7 ;
  assign n16346 = ~pi8  & n16345;
  assign n16347 = ~n16344 & ~n16346;
  assign n16348 = po5  & ~n16347;
  assign n16349 = ~po5  & n16347;
  assign n16350 = ~pi8  & po4 ;
  assign n16351 = pi9  & ~n16350;
  assign n16352 = ~pi9  & n16350;
  assign n16353 = ~n16351 & ~n16352;
  assign n16354 = ~n16349 & n16353;
  assign n16355 = ~n16348 & ~n16354;
  assign n16356 = po6  & ~n16355;
  assign n16357 = ~po6  & n16355;
  assign n16358 = po5  & ~po4 ;
  assign n16359 = ~n16352 & ~n16358;
  assign n16360 = pi10  & ~n16359;
  assign n16361 = ~pi10  & n16359;
  assign n16362 = ~n16360 & ~n16361;
  assign n16363 = ~n16357 & ~n16362;
  assign n16364 = ~n16356 & ~n16363;
  assign n16365 = po7  & ~n16364;
  assign n16366 = ~po7  & n16364;
  assign n16367 = ~n15815 & ~n15816;
  assign n16368 = po4  & n16367;
  assign n16369 = n15820 & ~n16368;
  assign n16370 = ~n15820 & n16368;
  assign n16371 = ~n16369 & ~n16370;
  assign n16372 = ~n16366 & ~n16371;
  assign n16373 = ~n16365 & ~n16372;
  assign n16374 = po8  & ~n16373;
  assign n16375 = ~po8  & n16373;
  assign n16376 = ~n15823 & ~n15824;
  assign n16377 = po4  & n16376;
  assign n16378 = ~n15829 & ~n16377;
  assign n16379 = n15829 & n16377;
  assign n16380 = ~n16378 & ~n16379;
  assign n16381 = ~n16375 & ~n16380;
  assign n16382 = ~n16374 & ~n16381;
  assign n16383 = po9  & ~n16382;
  assign n16384 = ~po9  & n16382;
  assign n16385 = ~n15832 & ~n15833;
  assign n16386 = po4  & n16385;
  assign n16387 = n15838 & n16386;
  assign n16388 = ~n15838 & ~n16386;
  assign n16389 = ~n16387 & ~n16388;
  assign n16390 = ~n16384 & ~n16389;
  assign n16391 = ~n16383 & ~n16390;
  assign n16392 = po10  & ~n16391;
  assign n16393 = ~po10  & n16391;
  assign n16394 = ~n15841 & ~n15842;
  assign n16395 = po4  & n16394;
  assign n16396 = ~n15847 & ~n16395;
  assign n16397 = n15847 & n16395;
  assign n16398 = ~n16396 & ~n16397;
  assign n16399 = ~n16393 & ~n16398;
  assign n16400 = ~n16392 & ~n16399;
  assign n16401 = po11  & ~n16400;
  assign n16402 = ~po11  & n16400;
  assign n16403 = ~n15850 & ~n15851;
  assign n16404 = po4  & n16403;
  assign n16405 = ~n15856 & ~n16404;
  assign n16406 = n15856 & n16404;
  assign n16407 = ~n16405 & ~n16406;
  assign n16408 = ~n16402 & ~n16407;
  assign n16409 = ~n16401 & ~n16408;
  assign n16410 = po12  & ~n16409;
  assign n16411 = ~po12  & n16409;
  assign n16412 = ~n15859 & ~n15860;
  assign n16413 = po4  & n16412;
  assign n16414 = ~n15865 & ~n16413;
  assign n16415 = n15865 & n16413;
  assign n16416 = ~n16414 & ~n16415;
  assign n16417 = ~n16411 & ~n16416;
  assign n16418 = ~n16410 & ~n16417;
  assign n16419 = po13  & ~n16418;
  assign n16420 = ~po13  & n16418;
  assign n16421 = ~n15868 & ~n15869;
  assign n16422 = po4  & n16421;
  assign n16423 = ~n15874 & ~n16422;
  assign n16424 = n15874 & n16422;
  assign n16425 = ~n16423 & ~n16424;
  assign n16426 = ~n16420 & ~n16425;
  assign n16427 = ~n16419 & ~n16426;
  assign n16428 = po14  & ~n16427;
  assign n16429 = ~po14  & n16427;
  assign n16430 = ~n15877 & ~n15878;
  assign n16431 = po4  & n16430;
  assign n16432 = ~n15883 & ~n16431;
  assign n16433 = n15883 & n16431;
  assign n16434 = ~n16432 & ~n16433;
  assign n16435 = ~n16429 & ~n16434;
  assign n16436 = ~n16428 & ~n16435;
  assign n16437 = po15  & ~n16436;
  assign n16438 = ~po15  & n16436;
  assign n16439 = ~n15886 & ~n15887;
  assign n16440 = po4  & n16439;
  assign n16441 = ~n15892 & ~n16440;
  assign n16442 = n15892 & n16440;
  assign n16443 = ~n16441 & ~n16442;
  assign n16444 = ~n16438 & ~n16443;
  assign n16445 = ~n16437 & ~n16444;
  assign n16446 = po16  & ~n16445;
  assign n16447 = ~po16  & n16445;
  assign n16448 = ~n15895 & ~n15896;
  assign n16449 = po4  & n16448;
  assign n16450 = ~n15901 & ~n16449;
  assign n16451 = n15901 & n16449;
  assign n16452 = ~n16450 & ~n16451;
  assign n16453 = ~n16447 & ~n16452;
  assign n16454 = ~n16446 & ~n16453;
  assign n16455 = po17  & ~n16454;
  assign n16456 = ~po17  & n16454;
  assign n16457 = ~n15904 & ~n15905;
  assign n16458 = po4  & n16457;
  assign n16459 = ~n15910 & ~n16458;
  assign n16460 = n15910 & n16458;
  assign n16461 = ~n16459 & ~n16460;
  assign n16462 = ~n16456 & ~n16461;
  assign n16463 = ~n16455 & ~n16462;
  assign n16464 = po18  & ~n16463;
  assign n16465 = ~po18  & n16463;
  assign n16466 = ~n15913 & ~n15914;
  assign n16467 = po4  & n16466;
  assign n16468 = ~n15919 & ~n16467;
  assign n16469 = n15919 & n16467;
  assign n16470 = ~n16468 & ~n16469;
  assign n16471 = ~n16465 & ~n16470;
  assign n16472 = ~n16464 & ~n16471;
  assign n16473 = po19  & ~n16472;
  assign n16474 = ~po19  & n16472;
  assign n16475 = ~n15922 & ~n15923;
  assign n16476 = po4  & n16475;
  assign n16477 = ~n15928 & ~n16476;
  assign n16478 = n15928 & n16476;
  assign n16479 = ~n16477 & ~n16478;
  assign n16480 = ~n16474 & ~n16479;
  assign n16481 = ~n16473 & ~n16480;
  assign n16482 = po20  & ~n16481;
  assign n16483 = ~po20  & n16481;
  assign n16484 = ~n15931 & ~n15932;
  assign n16485 = po4  & n16484;
  assign n16486 = ~n15937 & ~n16485;
  assign n16487 = n15937 & n16485;
  assign n16488 = ~n16486 & ~n16487;
  assign n16489 = ~n16483 & ~n16488;
  assign n16490 = ~n16482 & ~n16489;
  assign n16491 = po21  & ~n16490;
  assign n16492 = ~po21  & n16490;
  assign n16493 = ~n15940 & ~n15941;
  assign n16494 = po4  & n16493;
  assign n16495 = ~n15946 & ~n16494;
  assign n16496 = n15946 & n16494;
  assign n16497 = ~n16495 & ~n16496;
  assign n16498 = ~n16492 & ~n16497;
  assign n16499 = ~n16491 & ~n16498;
  assign n16500 = po22  & ~n16499;
  assign n16501 = ~po22  & n16499;
  assign n16502 = ~n15949 & ~n15950;
  assign n16503 = po4  & n16502;
  assign n16504 = ~n15955 & ~n16503;
  assign n16505 = n15955 & n16503;
  assign n16506 = ~n16504 & ~n16505;
  assign n16507 = ~n16501 & ~n16506;
  assign n16508 = ~n16500 & ~n16507;
  assign n16509 = po23  & ~n16508;
  assign n16510 = ~po23  & n16508;
  assign n16511 = ~n15958 & ~n15959;
  assign n16512 = po4  & n16511;
  assign n16513 = ~n15964 & ~n16512;
  assign n16514 = n15964 & n16512;
  assign n16515 = ~n16513 & ~n16514;
  assign n16516 = ~n16510 & ~n16515;
  assign n16517 = ~n16509 & ~n16516;
  assign n16518 = po24  & ~n16517;
  assign n16519 = ~po24  & n16517;
  assign n16520 = ~n15967 & ~n15968;
  assign n16521 = po4  & n16520;
  assign n16522 = ~n15973 & ~n16521;
  assign n16523 = n15973 & n16521;
  assign n16524 = ~n16522 & ~n16523;
  assign n16525 = ~n16519 & ~n16524;
  assign n16526 = ~n16518 & ~n16525;
  assign n16527 = po25  & ~n16526;
  assign n16528 = ~po25  & n16526;
  assign n16529 = ~n15976 & ~n15977;
  assign n16530 = po4  & n16529;
  assign n16531 = ~n15982 & ~n16530;
  assign n16532 = n15982 & n16530;
  assign n16533 = ~n16531 & ~n16532;
  assign n16534 = ~n16528 & ~n16533;
  assign n16535 = ~n16527 & ~n16534;
  assign n16536 = po26  & ~n16535;
  assign n16537 = ~po26  & n16535;
  assign n16538 = ~n15985 & ~n15986;
  assign n16539 = po4  & n16538;
  assign n16540 = ~n15991 & ~n16539;
  assign n16541 = n15991 & n16539;
  assign n16542 = ~n16540 & ~n16541;
  assign n16543 = ~n16537 & ~n16542;
  assign n16544 = ~n16536 & ~n16543;
  assign n16545 = po27  & ~n16544;
  assign n16546 = ~po27  & n16544;
  assign n16547 = ~n15994 & ~n15995;
  assign n16548 = po4  & n16547;
  assign n16549 = ~n16000 & ~n16548;
  assign n16550 = n16000 & n16548;
  assign n16551 = ~n16549 & ~n16550;
  assign n16552 = ~n16546 & ~n16551;
  assign n16553 = ~n16545 & ~n16552;
  assign n16554 = po28  & ~n16553;
  assign n16555 = ~po28  & n16553;
  assign n16556 = ~n16003 & ~n16004;
  assign n16557 = po4  & n16556;
  assign n16558 = ~n16009 & ~n16557;
  assign n16559 = n16009 & n16557;
  assign n16560 = ~n16558 & ~n16559;
  assign n16561 = ~n16555 & ~n16560;
  assign n16562 = ~n16554 & ~n16561;
  assign n16563 = po29  & ~n16562;
  assign n16564 = ~po29  & n16562;
  assign n16565 = ~n16012 & ~n16013;
  assign n16566 = po4  & n16565;
  assign n16567 = ~n16018 & ~n16566;
  assign n16568 = n16018 & n16566;
  assign n16569 = ~n16567 & ~n16568;
  assign n16570 = ~n16564 & ~n16569;
  assign n16571 = ~n16563 & ~n16570;
  assign n16572 = po30  & ~n16571;
  assign n16573 = ~po30  & n16571;
  assign n16574 = ~n16021 & ~n16022;
  assign n16575 = po4  & n16574;
  assign n16576 = ~n16027 & ~n16575;
  assign n16577 = n16027 & n16575;
  assign n16578 = ~n16576 & ~n16577;
  assign n16579 = ~n16573 & ~n16578;
  assign n16580 = ~n16572 & ~n16579;
  assign n16581 = po31  & ~n16580;
  assign n16582 = ~po31  & n16580;
  assign n16583 = ~n16030 & ~n16031;
  assign n16584 = po4  & n16583;
  assign n16585 = ~n16036 & ~n16584;
  assign n16586 = n16036 & n16584;
  assign n16587 = ~n16585 & ~n16586;
  assign n16588 = ~n16582 & ~n16587;
  assign n16589 = ~n16581 & ~n16588;
  assign n16590 = po32  & ~n16589;
  assign n16591 = ~po32  & n16589;
  assign n16592 = ~n16039 & ~n16040;
  assign n16593 = po4  & n16592;
  assign n16594 = ~n16045 & ~n16593;
  assign n16595 = n16045 & n16593;
  assign n16596 = ~n16594 & ~n16595;
  assign n16597 = ~n16591 & ~n16596;
  assign n16598 = ~n16590 & ~n16597;
  assign n16599 = po33  & ~n16598;
  assign n16600 = ~po33  & n16598;
  assign n16601 = ~n16048 & ~n16049;
  assign n16602 = po4  & n16601;
  assign n16603 = ~n16054 & ~n16602;
  assign n16604 = n16054 & n16602;
  assign n16605 = ~n16603 & ~n16604;
  assign n16606 = ~n16600 & ~n16605;
  assign n16607 = ~n16599 & ~n16606;
  assign n16608 = po34  & ~n16607;
  assign n16609 = ~po34  & n16607;
  assign n16610 = ~n16057 & ~n16058;
  assign n16611 = po4  & n16610;
  assign n16612 = ~n16063 & ~n16611;
  assign n16613 = n16063 & n16611;
  assign n16614 = ~n16612 & ~n16613;
  assign n16615 = ~n16609 & ~n16614;
  assign n16616 = ~n16608 & ~n16615;
  assign n16617 = po35  & ~n16616;
  assign n16618 = ~po35  & n16616;
  assign n16619 = ~n16066 & ~n16067;
  assign n16620 = po4  & n16619;
  assign n16621 = ~n16072 & ~n16620;
  assign n16622 = n16072 & n16620;
  assign n16623 = ~n16621 & ~n16622;
  assign n16624 = ~n16618 & ~n16623;
  assign n16625 = ~n16617 & ~n16624;
  assign n16626 = po36  & ~n16625;
  assign n16627 = ~po36  & n16625;
  assign n16628 = ~n16075 & ~n16076;
  assign n16629 = po4  & n16628;
  assign n16630 = ~n16081 & ~n16629;
  assign n16631 = n16081 & n16629;
  assign n16632 = ~n16630 & ~n16631;
  assign n16633 = ~n16627 & ~n16632;
  assign n16634 = ~n16626 & ~n16633;
  assign n16635 = po37  & ~n16634;
  assign n16636 = ~po37  & n16634;
  assign n16637 = ~n16084 & ~n16085;
  assign n16638 = po4  & n16637;
  assign n16639 = ~n16090 & ~n16638;
  assign n16640 = n16090 & n16638;
  assign n16641 = ~n16639 & ~n16640;
  assign n16642 = ~n16636 & ~n16641;
  assign n16643 = ~n16635 & ~n16642;
  assign n16644 = po38  & ~n16643;
  assign n16645 = ~po38  & n16643;
  assign n16646 = ~n16093 & ~n16094;
  assign n16647 = po4  & n16646;
  assign n16648 = ~n16099 & ~n16647;
  assign n16649 = n16099 & n16647;
  assign n16650 = ~n16648 & ~n16649;
  assign n16651 = ~n16645 & ~n16650;
  assign n16652 = ~n16644 & ~n16651;
  assign n16653 = po39  & ~n16652;
  assign n16654 = ~po39  & n16652;
  assign n16655 = ~n16102 & ~n16103;
  assign n16656 = po4  & n16655;
  assign n16657 = ~n16108 & ~n16656;
  assign n16658 = n16108 & n16656;
  assign n16659 = ~n16657 & ~n16658;
  assign n16660 = ~n16654 & ~n16659;
  assign n16661 = ~n16653 & ~n16660;
  assign n16662 = po40  & ~n16661;
  assign n16663 = ~po40  & n16661;
  assign n16664 = ~n16111 & ~n16112;
  assign n16665 = po4  & n16664;
  assign n16666 = ~n16117 & ~n16665;
  assign n16667 = n16117 & n16665;
  assign n16668 = ~n16666 & ~n16667;
  assign n16669 = ~n16663 & ~n16668;
  assign n16670 = ~n16662 & ~n16669;
  assign n16671 = po41  & ~n16670;
  assign n16672 = ~po41  & n16670;
  assign n16673 = ~n16120 & ~n16121;
  assign n16674 = po4  & n16673;
  assign n16675 = ~n16126 & ~n16674;
  assign n16676 = n16126 & n16674;
  assign n16677 = ~n16675 & ~n16676;
  assign n16678 = ~n16672 & ~n16677;
  assign n16679 = ~n16671 & ~n16678;
  assign n16680 = po42  & ~n16679;
  assign n16681 = ~po42  & n16679;
  assign n16682 = ~n16129 & ~n16130;
  assign n16683 = po4  & n16682;
  assign n16684 = ~n16135 & ~n16683;
  assign n16685 = n16135 & n16683;
  assign n16686 = ~n16684 & ~n16685;
  assign n16687 = ~n16681 & ~n16686;
  assign n16688 = ~n16680 & ~n16687;
  assign n16689 = po43  & ~n16688;
  assign n16690 = ~po43  & n16688;
  assign n16691 = ~n16138 & ~n16139;
  assign n16692 = po4  & n16691;
  assign n16693 = ~n16144 & ~n16692;
  assign n16694 = n16144 & n16692;
  assign n16695 = ~n16693 & ~n16694;
  assign n16696 = ~n16690 & ~n16695;
  assign n16697 = ~n16689 & ~n16696;
  assign n16698 = po44  & ~n16697;
  assign n16699 = ~po44  & n16697;
  assign n16700 = ~n16147 & ~n16148;
  assign n16701 = po4  & n16700;
  assign n16702 = ~n16153 & ~n16701;
  assign n16703 = n16153 & n16701;
  assign n16704 = ~n16702 & ~n16703;
  assign n16705 = ~n16699 & ~n16704;
  assign n16706 = ~n16698 & ~n16705;
  assign n16707 = po45  & ~n16706;
  assign n16708 = ~po45  & n16706;
  assign n16709 = ~n16156 & ~n16157;
  assign n16710 = po4  & n16709;
  assign n16711 = ~n16162 & ~n16710;
  assign n16712 = n16162 & n16710;
  assign n16713 = ~n16711 & ~n16712;
  assign n16714 = ~n16708 & ~n16713;
  assign n16715 = ~n16707 & ~n16714;
  assign n16716 = po46  & ~n16715;
  assign n16717 = ~po46  & n16715;
  assign n16718 = ~n16165 & ~n16166;
  assign n16719 = po4  & n16718;
  assign n16720 = ~n16171 & ~n16719;
  assign n16721 = n16171 & n16719;
  assign n16722 = ~n16720 & ~n16721;
  assign n16723 = ~n16717 & ~n16722;
  assign n16724 = ~n16716 & ~n16723;
  assign n16725 = po47  & ~n16724;
  assign n16726 = ~po47  & n16724;
  assign n16727 = ~n16174 & ~n16175;
  assign n16728 = po4  & n16727;
  assign n16729 = ~n16180 & ~n16728;
  assign n16730 = n16180 & n16728;
  assign n16731 = ~n16729 & ~n16730;
  assign n16732 = ~n16726 & ~n16731;
  assign n16733 = ~n16725 & ~n16732;
  assign n16734 = po48  & ~n16733;
  assign n16735 = ~po48  & n16733;
  assign n16736 = ~n16183 & ~n16184;
  assign n16737 = po4  & n16736;
  assign n16738 = ~n16189 & ~n16737;
  assign n16739 = n16189 & n16737;
  assign n16740 = ~n16738 & ~n16739;
  assign n16741 = ~n16735 & ~n16740;
  assign n16742 = ~n16734 & ~n16741;
  assign n16743 = po49  & ~n16742;
  assign n16744 = ~po49  & n16742;
  assign n16745 = ~n16192 & ~n16193;
  assign n16746 = po4  & n16745;
  assign n16747 = ~n16198 & ~n16746;
  assign n16748 = n16198 & n16746;
  assign n16749 = ~n16747 & ~n16748;
  assign n16750 = ~n16744 & ~n16749;
  assign n16751 = ~n16743 & ~n16750;
  assign n16752 = po50  & ~n16751;
  assign n16753 = ~po50  & n16751;
  assign n16754 = ~n16201 & ~n16202;
  assign n16755 = po4  & n16754;
  assign n16756 = ~n16207 & ~n16755;
  assign n16757 = n16207 & n16755;
  assign n16758 = ~n16756 & ~n16757;
  assign n16759 = ~n16753 & ~n16758;
  assign n16760 = ~n16752 & ~n16759;
  assign n16761 = po51  & ~n16760;
  assign n16762 = ~po51  & n16760;
  assign n16763 = ~n16210 & ~n16211;
  assign n16764 = po4  & n16763;
  assign n16765 = ~n16216 & ~n16764;
  assign n16766 = n16216 & n16764;
  assign n16767 = ~n16765 & ~n16766;
  assign n16768 = ~n16762 & ~n16767;
  assign n16769 = ~n16761 & ~n16768;
  assign n16770 = po52  & ~n16769;
  assign n16771 = ~po52  & n16769;
  assign n16772 = ~n16219 & ~n16220;
  assign n16773 = po4  & n16772;
  assign n16774 = ~n16225 & ~n16773;
  assign n16775 = n16225 & n16773;
  assign n16776 = ~n16774 & ~n16775;
  assign n16777 = ~n16771 & ~n16776;
  assign n16778 = ~n16770 & ~n16777;
  assign n16779 = po53  & ~n16778;
  assign n16780 = ~po53  & n16778;
  assign n16781 = ~n16228 & ~n16229;
  assign n16782 = po4  & n16781;
  assign n16783 = ~n16234 & ~n16782;
  assign n16784 = n16234 & n16782;
  assign n16785 = ~n16783 & ~n16784;
  assign n16786 = ~n16780 & ~n16785;
  assign n16787 = ~n16779 & ~n16786;
  assign n16788 = po54  & ~n16787;
  assign n16789 = ~po54  & n16787;
  assign n16790 = ~n16237 & ~n16238;
  assign n16791 = po4  & n16790;
  assign n16792 = ~n16243 & ~n16791;
  assign n16793 = n16243 & n16791;
  assign n16794 = ~n16792 & ~n16793;
  assign n16795 = ~n16789 & ~n16794;
  assign n16796 = ~n16788 & ~n16795;
  assign n16797 = po55  & ~n16796;
  assign n16798 = ~po55  & n16796;
  assign n16799 = ~n16246 & ~n16247;
  assign n16800 = po4  & n16799;
  assign n16801 = ~n16252 & ~n16800;
  assign n16802 = n16252 & n16800;
  assign n16803 = ~n16801 & ~n16802;
  assign n16804 = ~n16798 & ~n16803;
  assign n16805 = ~n16797 & ~n16804;
  assign n16806 = po56  & ~n16805;
  assign n16807 = ~po56  & n16805;
  assign n16808 = ~n16255 & ~n16256;
  assign n16809 = po4  & n16808;
  assign n16810 = ~n16261 & ~n16809;
  assign n16811 = n16261 & n16809;
  assign n16812 = ~n16810 & ~n16811;
  assign n16813 = ~n16807 & ~n16812;
  assign n16814 = ~n16806 & ~n16813;
  assign n16815 = po57  & ~n16814;
  assign n16816 = ~po57  & n16814;
  assign n16817 = ~n16264 & ~n16265;
  assign n16818 = po4  & n16817;
  assign n16819 = ~n16270 & ~n16818;
  assign n16820 = n16270 & n16818;
  assign n16821 = ~n16819 & ~n16820;
  assign n16822 = ~n16816 & ~n16821;
  assign n16823 = ~n16815 & ~n16822;
  assign n16824 = po58  & ~n16823;
  assign n16825 = ~po58  & n16823;
  assign n16826 = ~n16273 & ~n16274;
  assign n16827 = po4  & n16826;
  assign n16828 = ~n16279 & ~n16827;
  assign n16829 = n16279 & n16827;
  assign n16830 = ~n16828 & ~n16829;
  assign n16831 = ~n16825 & ~n16830;
  assign n16832 = ~n16824 & ~n16831;
  assign n16833 = po59  & ~n16832;
  assign n16834 = ~n16282 & ~n16288;
  assign n16835 = po4  & n16834;
  assign n16836 = ~n16287 & ~n16835;
  assign n16837 = n16287 & n16835;
  assign n16838 = ~n16836 & ~n16837;
  assign n16839 = ~po59  & n16832;
  assign n16840 = ~n16838 & ~n16839;
  assign n16841 = ~n16833 & ~n16840;
  assign n16842 = po60  & ~n16841;
  assign n16843 = ~po60  & n16841;
  assign n16844 = ~n16318 & ~n16319;
  assign n16845 = po4  & n16844;
  assign n16846 = ~n16324 & ~n16845;
  assign n16847 = n16324 & n16845;
  assign n16848 = ~n16846 & ~n16847;
  assign n16849 = ~n16343 & ~n16843;
  assign n16850 = ~n16842 & ~n16849;
  assign n16851 = po61  & ~n16850;
  assign n16852 = ~po61  & n16850;
  assign n16853 = ~n16300 & ~n16301;
  assign n16854 = po4  & n16853;
  assign n16855 = ~n16306 & ~n16854;
  assign n16856 = n16306 & n16854;
  assign n16857 = ~n16855 & ~n16856;
  assign n16858 = ~n16852 & ~n16857;
  assign n16859 = ~n16851 & ~n16858;
  assign n16860 = po62  & ~n16859;
  assign n16861 = ~po62  & n16859;
  assign n16862 = ~n16309 & ~n16310;
  assign n16863 = po4  & n16862;
  assign n16864 = ~n16315 & ~n16863;
  assign n16865 = n16315 & n16863;
  assign n16866 = ~n16864 & ~n16865;
  assign n16867 = ~n16861 & ~n16866;
  assign n16868 = ~n16860 & ~n16867;
  assign n16869 = n16848 & n16868;
  assign n16870 = ~n16848 & ~n16868;
  assign n16871 = n16328 & ~n16337;
  assign n16872 = ~n16327 & ~n16871;
  assign n16873 = n16870 & n16872;
  assign n16874 = ~po63  & ~n16873;
  assign n16875 = ~n16297 & ~n16337;
  assign n16876 = n16326 & ~n16875;
  assign n16877 = po63  & ~n16328;
  assign n16878 = ~n16876 & n16877;
  assign n16879 = ~n16874 & ~n16878;
  assign po3  = n16869 | ~n16879;
  assign n16881 = ~n16842 & ~n16843;
  assign n16882 = po3  & n16881;
  assign n16883 = ~n16343 & ~n16882;
  assign n16884 = n16343 & n16882;
  assign n16885 = ~n16883 & ~n16884;
  assign n16886 = pi6  & po3 ;
  assign n16887 = ~pi4  & ~pi5 ;
  assign n16888 = ~pi6  & n16887;
  assign n16889 = ~n16886 & ~n16888;
  assign n16890 = po4  & ~n16889;
  assign n16891 = ~po4  & n16889;
  assign n16892 = ~pi6  & po3 ;
  assign n16893 = pi7  & ~n16892;
  assign n16894 = ~pi7  & n16892;
  assign n16895 = ~n16893 & ~n16894;
  assign n16896 = ~n16891 & n16895;
  assign n16897 = ~n16890 & ~n16896;
  assign n16898 = po5  & ~n16897;
  assign n16899 = ~po5  & n16897;
  assign n16900 = po4  & ~po3 ;
  assign n16901 = ~n16894 & ~n16900;
  assign n16902 = pi8  & ~n16901;
  assign n16903 = ~pi8  & n16901;
  assign n16904 = ~n16902 & ~n16903;
  assign n16905 = ~n16899 & ~n16904;
  assign n16906 = ~n16898 & ~n16905;
  assign n16907 = po6  & ~n16906;
  assign n16908 = ~po6  & n16906;
  assign n16909 = ~n16348 & ~n16349;
  assign n16910 = po3  & n16909;
  assign n16911 = n16353 & ~n16910;
  assign n16912 = ~n16353 & n16910;
  assign n16913 = ~n16911 & ~n16912;
  assign n16914 = ~n16908 & ~n16913;
  assign n16915 = ~n16907 & ~n16914;
  assign n16916 = po7  & ~n16915;
  assign n16917 = ~po7  & n16915;
  assign n16918 = ~n16356 & ~n16357;
  assign n16919 = po3  & n16918;
  assign n16920 = ~n16362 & ~n16919;
  assign n16921 = n16362 & n16919;
  assign n16922 = ~n16920 & ~n16921;
  assign n16923 = ~n16917 & ~n16922;
  assign n16924 = ~n16916 & ~n16923;
  assign n16925 = po8  & ~n16924;
  assign n16926 = ~po8  & n16924;
  assign n16927 = ~n16365 & ~n16366;
  assign n16928 = po3  & n16927;
  assign n16929 = n16371 & n16928;
  assign n16930 = ~n16371 & ~n16928;
  assign n16931 = ~n16929 & ~n16930;
  assign n16932 = ~n16926 & ~n16931;
  assign n16933 = ~n16925 & ~n16932;
  assign n16934 = po9  & ~n16933;
  assign n16935 = ~po9  & n16933;
  assign n16936 = ~n16374 & ~n16375;
  assign n16937 = po3  & n16936;
  assign n16938 = ~n16380 & ~n16937;
  assign n16939 = n16380 & n16937;
  assign n16940 = ~n16938 & ~n16939;
  assign n16941 = ~n16935 & ~n16940;
  assign n16942 = ~n16934 & ~n16941;
  assign n16943 = po10  & ~n16942;
  assign n16944 = ~po10  & n16942;
  assign n16945 = ~n16383 & ~n16384;
  assign n16946 = po3  & n16945;
  assign n16947 = ~n16389 & ~n16946;
  assign n16948 = n16389 & n16946;
  assign n16949 = ~n16947 & ~n16948;
  assign n16950 = ~n16944 & ~n16949;
  assign n16951 = ~n16943 & ~n16950;
  assign n16952 = po11  & ~n16951;
  assign n16953 = ~po11  & n16951;
  assign n16954 = ~n16392 & ~n16393;
  assign n16955 = po3  & n16954;
  assign n16956 = ~n16398 & ~n16955;
  assign n16957 = n16398 & n16955;
  assign n16958 = ~n16956 & ~n16957;
  assign n16959 = ~n16953 & ~n16958;
  assign n16960 = ~n16952 & ~n16959;
  assign n16961 = po12  & ~n16960;
  assign n16962 = ~po12  & n16960;
  assign n16963 = ~n16401 & ~n16402;
  assign n16964 = po3  & n16963;
  assign n16965 = ~n16407 & ~n16964;
  assign n16966 = n16407 & n16964;
  assign n16967 = ~n16965 & ~n16966;
  assign n16968 = ~n16962 & ~n16967;
  assign n16969 = ~n16961 & ~n16968;
  assign n16970 = po13  & ~n16969;
  assign n16971 = ~po13  & n16969;
  assign n16972 = ~n16410 & ~n16411;
  assign n16973 = po3  & n16972;
  assign n16974 = ~n16416 & ~n16973;
  assign n16975 = n16416 & n16973;
  assign n16976 = ~n16974 & ~n16975;
  assign n16977 = ~n16971 & ~n16976;
  assign n16978 = ~n16970 & ~n16977;
  assign n16979 = po14  & ~n16978;
  assign n16980 = ~po14  & n16978;
  assign n16981 = ~n16419 & ~n16420;
  assign n16982 = po3  & n16981;
  assign n16983 = ~n16425 & ~n16982;
  assign n16984 = n16425 & n16982;
  assign n16985 = ~n16983 & ~n16984;
  assign n16986 = ~n16980 & ~n16985;
  assign n16987 = ~n16979 & ~n16986;
  assign n16988 = po15  & ~n16987;
  assign n16989 = ~po15  & n16987;
  assign n16990 = ~n16428 & ~n16429;
  assign n16991 = po3  & n16990;
  assign n16992 = ~n16434 & ~n16991;
  assign n16993 = n16434 & n16991;
  assign n16994 = ~n16992 & ~n16993;
  assign n16995 = ~n16989 & ~n16994;
  assign n16996 = ~n16988 & ~n16995;
  assign n16997 = po16  & ~n16996;
  assign n16998 = ~po16  & n16996;
  assign n16999 = ~n16437 & ~n16438;
  assign n17000 = po3  & n16999;
  assign n17001 = ~n16443 & ~n17000;
  assign n17002 = n16443 & n17000;
  assign n17003 = ~n17001 & ~n17002;
  assign n17004 = ~n16998 & ~n17003;
  assign n17005 = ~n16997 & ~n17004;
  assign n17006 = po17  & ~n17005;
  assign n17007 = ~po17  & n17005;
  assign n17008 = ~n16446 & ~n16447;
  assign n17009 = po3  & n17008;
  assign n17010 = ~n16452 & ~n17009;
  assign n17011 = n16452 & n17009;
  assign n17012 = ~n17010 & ~n17011;
  assign n17013 = ~n17007 & ~n17012;
  assign n17014 = ~n17006 & ~n17013;
  assign n17015 = po18  & ~n17014;
  assign n17016 = ~po18  & n17014;
  assign n17017 = ~n16455 & ~n16456;
  assign n17018 = po3  & n17017;
  assign n17019 = ~n16461 & ~n17018;
  assign n17020 = n16461 & n17018;
  assign n17021 = ~n17019 & ~n17020;
  assign n17022 = ~n17016 & ~n17021;
  assign n17023 = ~n17015 & ~n17022;
  assign n17024 = po19  & ~n17023;
  assign n17025 = ~po19  & n17023;
  assign n17026 = ~n16464 & ~n16465;
  assign n17027 = po3  & n17026;
  assign n17028 = ~n16470 & ~n17027;
  assign n17029 = n16470 & n17027;
  assign n17030 = ~n17028 & ~n17029;
  assign n17031 = ~n17025 & ~n17030;
  assign n17032 = ~n17024 & ~n17031;
  assign n17033 = po20  & ~n17032;
  assign n17034 = ~po20  & n17032;
  assign n17035 = ~n16473 & ~n16474;
  assign n17036 = po3  & n17035;
  assign n17037 = ~n16479 & ~n17036;
  assign n17038 = n16479 & n17036;
  assign n17039 = ~n17037 & ~n17038;
  assign n17040 = ~n17034 & ~n17039;
  assign n17041 = ~n17033 & ~n17040;
  assign n17042 = po21  & ~n17041;
  assign n17043 = ~po21  & n17041;
  assign n17044 = ~n16482 & ~n16483;
  assign n17045 = po3  & n17044;
  assign n17046 = ~n16488 & ~n17045;
  assign n17047 = n16488 & n17045;
  assign n17048 = ~n17046 & ~n17047;
  assign n17049 = ~n17043 & ~n17048;
  assign n17050 = ~n17042 & ~n17049;
  assign n17051 = po22  & ~n17050;
  assign n17052 = ~po22  & n17050;
  assign n17053 = ~n16491 & ~n16492;
  assign n17054 = po3  & n17053;
  assign n17055 = ~n16497 & ~n17054;
  assign n17056 = n16497 & n17054;
  assign n17057 = ~n17055 & ~n17056;
  assign n17058 = ~n17052 & ~n17057;
  assign n17059 = ~n17051 & ~n17058;
  assign n17060 = po23  & ~n17059;
  assign n17061 = ~po23  & n17059;
  assign n17062 = ~n16500 & ~n16501;
  assign n17063 = po3  & n17062;
  assign n17064 = ~n16506 & ~n17063;
  assign n17065 = n16506 & n17063;
  assign n17066 = ~n17064 & ~n17065;
  assign n17067 = ~n17061 & ~n17066;
  assign n17068 = ~n17060 & ~n17067;
  assign n17069 = po24  & ~n17068;
  assign n17070 = ~po24  & n17068;
  assign n17071 = ~n16509 & ~n16510;
  assign n17072 = po3  & n17071;
  assign n17073 = ~n16515 & ~n17072;
  assign n17074 = n16515 & n17072;
  assign n17075 = ~n17073 & ~n17074;
  assign n17076 = ~n17070 & ~n17075;
  assign n17077 = ~n17069 & ~n17076;
  assign n17078 = po25  & ~n17077;
  assign n17079 = ~po25  & n17077;
  assign n17080 = ~n16518 & ~n16519;
  assign n17081 = po3  & n17080;
  assign n17082 = ~n16524 & ~n17081;
  assign n17083 = n16524 & n17081;
  assign n17084 = ~n17082 & ~n17083;
  assign n17085 = ~n17079 & ~n17084;
  assign n17086 = ~n17078 & ~n17085;
  assign n17087 = po26  & ~n17086;
  assign n17088 = ~po26  & n17086;
  assign n17089 = ~n16527 & ~n16528;
  assign n17090 = po3  & n17089;
  assign n17091 = ~n16533 & ~n17090;
  assign n17092 = n16533 & n17090;
  assign n17093 = ~n17091 & ~n17092;
  assign n17094 = ~n17088 & ~n17093;
  assign n17095 = ~n17087 & ~n17094;
  assign n17096 = po27  & ~n17095;
  assign n17097 = ~po27  & n17095;
  assign n17098 = ~n16536 & ~n16537;
  assign n17099 = po3  & n17098;
  assign n17100 = ~n16542 & ~n17099;
  assign n17101 = n16542 & n17099;
  assign n17102 = ~n17100 & ~n17101;
  assign n17103 = ~n17097 & ~n17102;
  assign n17104 = ~n17096 & ~n17103;
  assign n17105 = po28  & ~n17104;
  assign n17106 = ~po28  & n17104;
  assign n17107 = ~n16545 & ~n16546;
  assign n17108 = po3  & n17107;
  assign n17109 = ~n16551 & ~n17108;
  assign n17110 = n16551 & n17108;
  assign n17111 = ~n17109 & ~n17110;
  assign n17112 = ~n17106 & ~n17111;
  assign n17113 = ~n17105 & ~n17112;
  assign n17114 = po29  & ~n17113;
  assign n17115 = ~po29  & n17113;
  assign n17116 = ~n16554 & ~n16555;
  assign n17117 = po3  & n17116;
  assign n17118 = ~n16560 & ~n17117;
  assign n17119 = n16560 & n17117;
  assign n17120 = ~n17118 & ~n17119;
  assign n17121 = ~n17115 & ~n17120;
  assign n17122 = ~n17114 & ~n17121;
  assign n17123 = po30  & ~n17122;
  assign n17124 = ~po30  & n17122;
  assign n17125 = ~n16563 & ~n16564;
  assign n17126 = po3  & n17125;
  assign n17127 = ~n16569 & ~n17126;
  assign n17128 = n16569 & n17126;
  assign n17129 = ~n17127 & ~n17128;
  assign n17130 = ~n17124 & ~n17129;
  assign n17131 = ~n17123 & ~n17130;
  assign n17132 = po31  & ~n17131;
  assign n17133 = ~po31  & n17131;
  assign n17134 = ~n16572 & ~n16573;
  assign n17135 = po3  & n17134;
  assign n17136 = ~n16578 & ~n17135;
  assign n17137 = n16578 & n17135;
  assign n17138 = ~n17136 & ~n17137;
  assign n17139 = ~n17133 & ~n17138;
  assign n17140 = ~n17132 & ~n17139;
  assign n17141 = po32  & ~n17140;
  assign n17142 = ~po32  & n17140;
  assign n17143 = ~n16581 & ~n16582;
  assign n17144 = po3  & n17143;
  assign n17145 = ~n16587 & ~n17144;
  assign n17146 = n16587 & n17144;
  assign n17147 = ~n17145 & ~n17146;
  assign n17148 = ~n17142 & ~n17147;
  assign n17149 = ~n17141 & ~n17148;
  assign n17150 = po33  & ~n17149;
  assign n17151 = ~po33  & n17149;
  assign n17152 = ~n16590 & ~n16591;
  assign n17153 = po3  & n17152;
  assign n17154 = ~n16596 & ~n17153;
  assign n17155 = n16596 & n17153;
  assign n17156 = ~n17154 & ~n17155;
  assign n17157 = ~n17151 & ~n17156;
  assign n17158 = ~n17150 & ~n17157;
  assign n17159 = po34  & ~n17158;
  assign n17160 = ~po34  & n17158;
  assign n17161 = ~n16599 & ~n16600;
  assign n17162 = po3  & n17161;
  assign n17163 = ~n16605 & ~n17162;
  assign n17164 = n16605 & n17162;
  assign n17165 = ~n17163 & ~n17164;
  assign n17166 = ~n17160 & ~n17165;
  assign n17167 = ~n17159 & ~n17166;
  assign n17168 = po35  & ~n17167;
  assign n17169 = ~po35  & n17167;
  assign n17170 = ~n16608 & ~n16609;
  assign n17171 = po3  & n17170;
  assign n17172 = ~n16614 & ~n17171;
  assign n17173 = n16614 & n17171;
  assign n17174 = ~n17172 & ~n17173;
  assign n17175 = ~n17169 & ~n17174;
  assign n17176 = ~n17168 & ~n17175;
  assign n17177 = po36  & ~n17176;
  assign n17178 = ~po36  & n17176;
  assign n17179 = ~n16617 & ~n16618;
  assign n17180 = po3  & n17179;
  assign n17181 = ~n16623 & ~n17180;
  assign n17182 = n16623 & n17180;
  assign n17183 = ~n17181 & ~n17182;
  assign n17184 = ~n17178 & ~n17183;
  assign n17185 = ~n17177 & ~n17184;
  assign n17186 = po37  & ~n17185;
  assign n17187 = ~po37  & n17185;
  assign n17188 = ~n16626 & ~n16627;
  assign n17189 = po3  & n17188;
  assign n17190 = ~n16632 & ~n17189;
  assign n17191 = n16632 & n17189;
  assign n17192 = ~n17190 & ~n17191;
  assign n17193 = ~n17187 & ~n17192;
  assign n17194 = ~n17186 & ~n17193;
  assign n17195 = po38  & ~n17194;
  assign n17196 = ~po38  & n17194;
  assign n17197 = ~n16635 & ~n16636;
  assign n17198 = po3  & n17197;
  assign n17199 = ~n16641 & ~n17198;
  assign n17200 = n16641 & n17198;
  assign n17201 = ~n17199 & ~n17200;
  assign n17202 = ~n17196 & ~n17201;
  assign n17203 = ~n17195 & ~n17202;
  assign n17204 = po39  & ~n17203;
  assign n17205 = ~po39  & n17203;
  assign n17206 = ~n16644 & ~n16645;
  assign n17207 = po3  & n17206;
  assign n17208 = ~n16650 & ~n17207;
  assign n17209 = n16650 & n17207;
  assign n17210 = ~n17208 & ~n17209;
  assign n17211 = ~n17205 & ~n17210;
  assign n17212 = ~n17204 & ~n17211;
  assign n17213 = po40  & ~n17212;
  assign n17214 = ~po40  & n17212;
  assign n17215 = ~n16653 & ~n16654;
  assign n17216 = po3  & n17215;
  assign n17217 = ~n16659 & ~n17216;
  assign n17218 = n16659 & n17216;
  assign n17219 = ~n17217 & ~n17218;
  assign n17220 = ~n17214 & ~n17219;
  assign n17221 = ~n17213 & ~n17220;
  assign n17222 = po41  & ~n17221;
  assign n17223 = ~po41  & n17221;
  assign n17224 = ~n16662 & ~n16663;
  assign n17225 = po3  & n17224;
  assign n17226 = ~n16668 & ~n17225;
  assign n17227 = n16668 & n17225;
  assign n17228 = ~n17226 & ~n17227;
  assign n17229 = ~n17223 & ~n17228;
  assign n17230 = ~n17222 & ~n17229;
  assign n17231 = po42  & ~n17230;
  assign n17232 = ~po42  & n17230;
  assign n17233 = ~n16671 & ~n16672;
  assign n17234 = po3  & n17233;
  assign n17235 = ~n16677 & ~n17234;
  assign n17236 = n16677 & n17234;
  assign n17237 = ~n17235 & ~n17236;
  assign n17238 = ~n17232 & ~n17237;
  assign n17239 = ~n17231 & ~n17238;
  assign n17240 = po43  & ~n17239;
  assign n17241 = ~po43  & n17239;
  assign n17242 = ~n16680 & ~n16681;
  assign n17243 = po3  & n17242;
  assign n17244 = ~n16686 & ~n17243;
  assign n17245 = n16686 & n17243;
  assign n17246 = ~n17244 & ~n17245;
  assign n17247 = ~n17241 & ~n17246;
  assign n17248 = ~n17240 & ~n17247;
  assign n17249 = po44  & ~n17248;
  assign n17250 = ~po44  & n17248;
  assign n17251 = ~n16689 & ~n16690;
  assign n17252 = po3  & n17251;
  assign n17253 = ~n16695 & ~n17252;
  assign n17254 = n16695 & n17252;
  assign n17255 = ~n17253 & ~n17254;
  assign n17256 = ~n17250 & ~n17255;
  assign n17257 = ~n17249 & ~n17256;
  assign n17258 = po45  & ~n17257;
  assign n17259 = ~po45  & n17257;
  assign n17260 = ~n16698 & ~n16699;
  assign n17261 = po3  & n17260;
  assign n17262 = ~n16704 & ~n17261;
  assign n17263 = n16704 & n17261;
  assign n17264 = ~n17262 & ~n17263;
  assign n17265 = ~n17259 & ~n17264;
  assign n17266 = ~n17258 & ~n17265;
  assign n17267 = po46  & ~n17266;
  assign n17268 = ~po46  & n17266;
  assign n17269 = ~n16707 & ~n16708;
  assign n17270 = po3  & n17269;
  assign n17271 = ~n16713 & ~n17270;
  assign n17272 = n16713 & n17270;
  assign n17273 = ~n17271 & ~n17272;
  assign n17274 = ~n17268 & ~n17273;
  assign n17275 = ~n17267 & ~n17274;
  assign n17276 = po47  & ~n17275;
  assign n17277 = ~po47  & n17275;
  assign n17278 = ~n16716 & ~n16717;
  assign n17279 = po3  & n17278;
  assign n17280 = ~n16722 & ~n17279;
  assign n17281 = n16722 & n17279;
  assign n17282 = ~n17280 & ~n17281;
  assign n17283 = ~n17277 & ~n17282;
  assign n17284 = ~n17276 & ~n17283;
  assign n17285 = po48  & ~n17284;
  assign n17286 = ~po48  & n17284;
  assign n17287 = ~n16725 & ~n16726;
  assign n17288 = po3  & n17287;
  assign n17289 = ~n16731 & ~n17288;
  assign n17290 = n16731 & n17288;
  assign n17291 = ~n17289 & ~n17290;
  assign n17292 = ~n17286 & ~n17291;
  assign n17293 = ~n17285 & ~n17292;
  assign n17294 = po49  & ~n17293;
  assign n17295 = ~po49  & n17293;
  assign n17296 = ~n16734 & ~n16735;
  assign n17297 = po3  & n17296;
  assign n17298 = ~n16740 & ~n17297;
  assign n17299 = n16740 & n17297;
  assign n17300 = ~n17298 & ~n17299;
  assign n17301 = ~n17295 & ~n17300;
  assign n17302 = ~n17294 & ~n17301;
  assign n17303 = po50  & ~n17302;
  assign n17304 = ~po50  & n17302;
  assign n17305 = ~n16743 & ~n16744;
  assign n17306 = po3  & n17305;
  assign n17307 = ~n16749 & ~n17306;
  assign n17308 = n16749 & n17306;
  assign n17309 = ~n17307 & ~n17308;
  assign n17310 = ~n17304 & ~n17309;
  assign n17311 = ~n17303 & ~n17310;
  assign n17312 = po51  & ~n17311;
  assign n17313 = ~po51  & n17311;
  assign n17314 = ~n16752 & ~n16753;
  assign n17315 = po3  & n17314;
  assign n17316 = ~n16758 & ~n17315;
  assign n17317 = n16758 & n17315;
  assign n17318 = ~n17316 & ~n17317;
  assign n17319 = ~n17313 & ~n17318;
  assign n17320 = ~n17312 & ~n17319;
  assign n17321 = po52  & ~n17320;
  assign n17322 = ~po52  & n17320;
  assign n17323 = ~n16761 & ~n16762;
  assign n17324 = po3  & n17323;
  assign n17325 = ~n16767 & ~n17324;
  assign n17326 = n16767 & n17324;
  assign n17327 = ~n17325 & ~n17326;
  assign n17328 = ~n17322 & ~n17327;
  assign n17329 = ~n17321 & ~n17328;
  assign n17330 = po53  & ~n17329;
  assign n17331 = ~po53  & n17329;
  assign n17332 = ~n16770 & ~n16771;
  assign n17333 = po3  & n17332;
  assign n17334 = ~n16776 & ~n17333;
  assign n17335 = n16776 & n17333;
  assign n17336 = ~n17334 & ~n17335;
  assign n17337 = ~n17331 & ~n17336;
  assign n17338 = ~n17330 & ~n17337;
  assign n17339 = po54  & ~n17338;
  assign n17340 = ~po54  & n17338;
  assign n17341 = ~n16779 & ~n16780;
  assign n17342 = po3  & n17341;
  assign n17343 = ~n16785 & ~n17342;
  assign n17344 = n16785 & n17342;
  assign n17345 = ~n17343 & ~n17344;
  assign n17346 = ~n17340 & ~n17345;
  assign n17347 = ~n17339 & ~n17346;
  assign n17348 = po55  & ~n17347;
  assign n17349 = ~po55  & n17347;
  assign n17350 = ~n16788 & ~n16789;
  assign n17351 = po3  & n17350;
  assign n17352 = ~n16794 & ~n17351;
  assign n17353 = n16794 & n17351;
  assign n17354 = ~n17352 & ~n17353;
  assign n17355 = ~n17349 & ~n17354;
  assign n17356 = ~n17348 & ~n17355;
  assign n17357 = po56  & ~n17356;
  assign n17358 = ~po56  & n17356;
  assign n17359 = ~n16797 & ~n16798;
  assign n17360 = po3  & n17359;
  assign n17361 = ~n16803 & ~n17360;
  assign n17362 = n16803 & n17360;
  assign n17363 = ~n17361 & ~n17362;
  assign n17364 = ~n17358 & ~n17363;
  assign n17365 = ~n17357 & ~n17364;
  assign n17366 = po57  & ~n17365;
  assign n17367 = ~po57  & n17365;
  assign n17368 = ~n16806 & ~n16807;
  assign n17369 = po3  & n17368;
  assign n17370 = ~n16812 & ~n17369;
  assign n17371 = n16812 & n17369;
  assign n17372 = ~n17370 & ~n17371;
  assign n17373 = ~n17367 & ~n17372;
  assign n17374 = ~n17366 & ~n17373;
  assign n17375 = po58  & ~n17374;
  assign n17376 = ~po58  & n17374;
  assign n17377 = ~n16815 & ~n16816;
  assign n17378 = po3  & n17377;
  assign n17379 = ~n16821 & ~n17378;
  assign n17380 = n16821 & n17378;
  assign n17381 = ~n17379 & ~n17380;
  assign n17382 = ~n17376 & ~n17381;
  assign n17383 = ~n17375 & ~n17382;
  assign n17384 = po59  & ~n17383;
  assign n17385 = ~po59  & n17383;
  assign n17386 = ~n16824 & ~n16825;
  assign n17387 = po3  & n17386;
  assign n17388 = ~n16830 & ~n17387;
  assign n17389 = n16830 & n17387;
  assign n17390 = ~n17388 & ~n17389;
  assign n17391 = ~n17385 & ~n17390;
  assign n17392 = ~n17384 & ~n17391;
  assign n17393 = po60  & ~n17392;
  assign n17394 = ~n16833 & ~n16839;
  assign n17395 = po3  & n17394;
  assign n17396 = ~n16838 & ~n17395;
  assign n17397 = n16838 & n17395;
  assign n17398 = ~n17396 & ~n17397;
  assign n17399 = ~po60  & n17392;
  assign n17400 = ~n17398 & ~n17399;
  assign n17401 = ~n17393 & ~n17400;
  assign n17402 = po61  & ~n17401;
  assign n17403 = ~po61  & n17401;
  assign n17404 = ~n16860 & ~n16861;
  assign n17405 = po3  & n17404;
  assign n17406 = ~n16866 & ~n17405;
  assign n17407 = n16866 & n17405;
  assign n17408 = ~n17406 & ~n17407;
  assign n17409 = ~n16885 & ~n17403;
  assign n17410 = ~n17402 & ~n17409;
  assign n17411 = po62  & ~n17410;
  assign n17412 = ~po62  & n17410;
  assign n17413 = ~n16851 & ~n16852;
  assign n17414 = po3  & n17413;
  assign n17415 = ~n16857 & ~n17414;
  assign n17416 = n16857 & n17414;
  assign n17417 = ~n17415 & ~n17416;
  assign n17418 = ~n17412 & ~n17417;
  assign n17419 = ~n17411 & ~n17418;
  assign n17420 = n17408 & n17419;
  assign n17421 = ~n17408 & ~n17419;
  assign n17422 = n16870 & ~n16879;
  assign n17423 = ~n16869 & ~n17422;
  assign n17424 = n17421 & n17423;
  assign n17425 = ~po63  & ~n17424;
  assign n17426 = ~n16848 & ~n16879;
  assign n17427 = n16868 & ~n17426;
  assign n17428 = po63  & ~n16870;
  assign n17429 = ~n17427 & n17428;
  assign n17430 = ~n17425 & ~n17429;
  assign po2  = n17420 | ~n17430;
  assign n17432 = ~n17402 & ~n17403;
  assign n17433 = po2  & n17432;
  assign n17434 = ~n16885 & ~n17433;
  assign n17435 = n16885 & n17433;
  assign n17436 = ~n17434 & ~n17435;
  assign n17437 = pi4  & po2 ;
  assign n17438 = ~pi2  & ~pi3 ;
  assign n17439 = ~pi4  & n17438;
  assign n17440 = ~n17437 & ~n17439;
  assign n17441 = po3  & ~n17440;
  assign n17442 = ~po3  & n17440;
  assign n17443 = ~pi4  & po2 ;
  assign n17444 = pi5  & ~n17443;
  assign n17445 = ~pi5  & n17443;
  assign n17446 = ~n17444 & ~n17445;
  assign n17447 = ~n17442 & n17446;
  assign n17448 = ~n17441 & ~n17447;
  assign n17449 = po4  & ~n17448;
  assign n17450 = ~po4  & n17448;
  assign n17451 = po3  & ~po2 ;
  assign n17452 = ~n17445 & ~n17451;
  assign n17453 = pi6  & ~n17452;
  assign n17454 = ~pi6  & n17452;
  assign n17455 = ~n17453 & ~n17454;
  assign n17456 = ~n17450 & ~n17455;
  assign n17457 = ~n17449 & ~n17456;
  assign n17458 = po5  & ~n17457;
  assign n17459 = ~po5  & n17457;
  assign n17460 = ~n16890 & ~n16891;
  assign n17461 = po2  & n17460;
  assign n17462 = n16895 & ~n17461;
  assign n17463 = ~n16895 & n17461;
  assign n17464 = ~n17462 & ~n17463;
  assign n17465 = ~n17459 & ~n17464;
  assign n17466 = ~n17458 & ~n17465;
  assign n17467 = po6  & ~n17466;
  assign n17468 = ~po6  & n17466;
  assign n17469 = ~n16898 & ~n16899;
  assign n17470 = po2  & n17469;
  assign n17471 = ~n16904 & ~n17470;
  assign n17472 = n16904 & n17470;
  assign n17473 = ~n17471 & ~n17472;
  assign n17474 = ~n17468 & ~n17473;
  assign n17475 = ~n17467 & ~n17474;
  assign n17476 = po7  & ~n17475;
  assign n17477 = ~po7  & n17475;
  assign n17478 = ~n16907 & ~n16908;
  assign n17479 = po2  & n17478;
  assign n17480 = n16913 & n17479;
  assign n17481 = ~n16913 & ~n17479;
  assign n17482 = ~n17480 & ~n17481;
  assign n17483 = ~n17477 & ~n17482;
  assign n17484 = ~n17476 & ~n17483;
  assign n17485 = po8  & ~n17484;
  assign n17486 = ~po8  & n17484;
  assign n17487 = ~n16916 & ~n16917;
  assign n17488 = po2  & n17487;
  assign n17489 = ~n16922 & ~n17488;
  assign n17490 = n16922 & n17488;
  assign n17491 = ~n17489 & ~n17490;
  assign n17492 = ~n17486 & ~n17491;
  assign n17493 = ~n17485 & ~n17492;
  assign n17494 = po9  & ~n17493;
  assign n17495 = ~po9  & n17493;
  assign n17496 = ~n16925 & ~n16926;
  assign n17497 = po2  & n17496;
  assign n17498 = ~n16931 & ~n17497;
  assign n17499 = n16931 & n17497;
  assign n17500 = ~n17498 & ~n17499;
  assign n17501 = ~n17495 & ~n17500;
  assign n17502 = ~n17494 & ~n17501;
  assign n17503 = po10  & ~n17502;
  assign n17504 = ~po10  & n17502;
  assign n17505 = ~n16934 & ~n16935;
  assign n17506 = po2  & n17505;
  assign n17507 = ~n16940 & ~n17506;
  assign n17508 = n16940 & n17506;
  assign n17509 = ~n17507 & ~n17508;
  assign n17510 = ~n17504 & ~n17509;
  assign n17511 = ~n17503 & ~n17510;
  assign n17512 = po11  & ~n17511;
  assign n17513 = ~po11  & n17511;
  assign n17514 = ~n16943 & ~n16944;
  assign n17515 = po2  & n17514;
  assign n17516 = ~n16949 & ~n17515;
  assign n17517 = n16949 & n17515;
  assign n17518 = ~n17516 & ~n17517;
  assign n17519 = ~n17513 & ~n17518;
  assign n17520 = ~n17512 & ~n17519;
  assign n17521 = po12  & ~n17520;
  assign n17522 = ~po12  & n17520;
  assign n17523 = ~n16952 & ~n16953;
  assign n17524 = po2  & n17523;
  assign n17525 = ~n16958 & ~n17524;
  assign n17526 = n16958 & n17524;
  assign n17527 = ~n17525 & ~n17526;
  assign n17528 = ~n17522 & ~n17527;
  assign n17529 = ~n17521 & ~n17528;
  assign n17530 = po13  & ~n17529;
  assign n17531 = ~po13  & n17529;
  assign n17532 = ~n16961 & ~n16962;
  assign n17533 = po2  & n17532;
  assign n17534 = ~n16967 & ~n17533;
  assign n17535 = n16967 & n17533;
  assign n17536 = ~n17534 & ~n17535;
  assign n17537 = ~n17531 & ~n17536;
  assign n17538 = ~n17530 & ~n17537;
  assign n17539 = po14  & ~n17538;
  assign n17540 = ~po14  & n17538;
  assign n17541 = ~n16970 & ~n16971;
  assign n17542 = po2  & n17541;
  assign n17543 = ~n16976 & ~n17542;
  assign n17544 = n16976 & n17542;
  assign n17545 = ~n17543 & ~n17544;
  assign n17546 = ~n17540 & ~n17545;
  assign n17547 = ~n17539 & ~n17546;
  assign n17548 = po15  & ~n17547;
  assign n17549 = ~po15  & n17547;
  assign n17550 = ~n16979 & ~n16980;
  assign n17551 = po2  & n17550;
  assign n17552 = ~n16985 & ~n17551;
  assign n17553 = n16985 & n17551;
  assign n17554 = ~n17552 & ~n17553;
  assign n17555 = ~n17549 & ~n17554;
  assign n17556 = ~n17548 & ~n17555;
  assign n17557 = po16  & ~n17556;
  assign n17558 = ~po16  & n17556;
  assign n17559 = ~n16988 & ~n16989;
  assign n17560 = po2  & n17559;
  assign n17561 = ~n16994 & ~n17560;
  assign n17562 = n16994 & n17560;
  assign n17563 = ~n17561 & ~n17562;
  assign n17564 = ~n17558 & ~n17563;
  assign n17565 = ~n17557 & ~n17564;
  assign n17566 = po17  & ~n17565;
  assign n17567 = ~po17  & n17565;
  assign n17568 = ~n16997 & ~n16998;
  assign n17569 = po2  & n17568;
  assign n17570 = ~n17003 & ~n17569;
  assign n17571 = n17003 & n17569;
  assign n17572 = ~n17570 & ~n17571;
  assign n17573 = ~n17567 & ~n17572;
  assign n17574 = ~n17566 & ~n17573;
  assign n17575 = po18  & ~n17574;
  assign n17576 = ~po18  & n17574;
  assign n17577 = ~n17006 & ~n17007;
  assign n17578 = po2  & n17577;
  assign n17579 = ~n17012 & ~n17578;
  assign n17580 = n17012 & n17578;
  assign n17581 = ~n17579 & ~n17580;
  assign n17582 = ~n17576 & ~n17581;
  assign n17583 = ~n17575 & ~n17582;
  assign n17584 = po19  & ~n17583;
  assign n17585 = ~po19  & n17583;
  assign n17586 = ~n17015 & ~n17016;
  assign n17587 = po2  & n17586;
  assign n17588 = ~n17021 & ~n17587;
  assign n17589 = n17021 & n17587;
  assign n17590 = ~n17588 & ~n17589;
  assign n17591 = ~n17585 & ~n17590;
  assign n17592 = ~n17584 & ~n17591;
  assign n17593 = po20  & ~n17592;
  assign n17594 = ~po20  & n17592;
  assign n17595 = ~n17024 & ~n17025;
  assign n17596 = po2  & n17595;
  assign n17597 = ~n17030 & ~n17596;
  assign n17598 = n17030 & n17596;
  assign n17599 = ~n17597 & ~n17598;
  assign n17600 = ~n17594 & ~n17599;
  assign n17601 = ~n17593 & ~n17600;
  assign n17602 = po21  & ~n17601;
  assign n17603 = ~po21  & n17601;
  assign n17604 = ~n17033 & ~n17034;
  assign n17605 = po2  & n17604;
  assign n17606 = ~n17039 & ~n17605;
  assign n17607 = n17039 & n17605;
  assign n17608 = ~n17606 & ~n17607;
  assign n17609 = ~n17603 & ~n17608;
  assign n17610 = ~n17602 & ~n17609;
  assign n17611 = po22  & ~n17610;
  assign n17612 = ~po22  & n17610;
  assign n17613 = ~n17042 & ~n17043;
  assign n17614 = po2  & n17613;
  assign n17615 = ~n17048 & ~n17614;
  assign n17616 = n17048 & n17614;
  assign n17617 = ~n17615 & ~n17616;
  assign n17618 = ~n17612 & ~n17617;
  assign n17619 = ~n17611 & ~n17618;
  assign n17620 = po23  & ~n17619;
  assign n17621 = ~po23  & n17619;
  assign n17622 = ~n17051 & ~n17052;
  assign n17623 = po2  & n17622;
  assign n17624 = ~n17057 & ~n17623;
  assign n17625 = n17057 & n17623;
  assign n17626 = ~n17624 & ~n17625;
  assign n17627 = ~n17621 & ~n17626;
  assign n17628 = ~n17620 & ~n17627;
  assign n17629 = po24  & ~n17628;
  assign n17630 = ~po24  & n17628;
  assign n17631 = ~n17060 & ~n17061;
  assign n17632 = po2  & n17631;
  assign n17633 = ~n17066 & ~n17632;
  assign n17634 = n17066 & n17632;
  assign n17635 = ~n17633 & ~n17634;
  assign n17636 = ~n17630 & ~n17635;
  assign n17637 = ~n17629 & ~n17636;
  assign n17638 = po25  & ~n17637;
  assign n17639 = ~po25  & n17637;
  assign n17640 = ~n17069 & ~n17070;
  assign n17641 = po2  & n17640;
  assign n17642 = ~n17075 & ~n17641;
  assign n17643 = n17075 & n17641;
  assign n17644 = ~n17642 & ~n17643;
  assign n17645 = ~n17639 & ~n17644;
  assign n17646 = ~n17638 & ~n17645;
  assign n17647 = po26  & ~n17646;
  assign n17648 = ~po26  & n17646;
  assign n17649 = ~n17078 & ~n17079;
  assign n17650 = po2  & n17649;
  assign n17651 = ~n17084 & ~n17650;
  assign n17652 = n17084 & n17650;
  assign n17653 = ~n17651 & ~n17652;
  assign n17654 = ~n17648 & ~n17653;
  assign n17655 = ~n17647 & ~n17654;
  assign n17656 = po27  & ~n17655;
  assign n17657 = ~po27  & n17655;
  assign n17658 = ~n17087 & ~n17088;
  assign n17659 = po2  & n17658;
  assign n17660 = ~n17093 & ~n17659;
  assign n17661 = n17093 & n17659;
  assign n17662 = ~n17660 & ~n17661;
  assign n17663 = ~n17657 & ~n17662;
  assign n17664 = ~n17656 & ~n17663;
  assign n17665 = po28  & ~n17664;
  assign n17666 = ~po28  & n17664;
  assign n17667 = ~n17096 & ~n17097;
  assign n17668 = po2  & n17667;
  assign n17669 = ~n17102 & ~n17668;
  assign n17670 = n17102 & n17668;
  assign n17671 = ~n17669 & ~n17670;
  assign n17672 = ~n17666 & ~n17671;
  assign n17673 = ~n17665 & ~n17672;
  assign n17674 = po29  & ~n17673;
  assign n17675 = ~po29  & n17673;
  assign n17676 = ~n17105 & ~n17106;
  assign n17677 = po2  & n17676;
  assign n17678 = ~n17111 & ~n17677;
  assign n17679 = n17111 & n17677;
  assign n17680 = ~n17678 & ~n17679;
  assign n17681 = ~n17675 & ~n17680;
  assign n17682 = ~n17674 & ~n17681;
  assign n17683 = po30  & ~n17682;
  assign n17684 = ~po30  & n17682;
  assign n17685 = ~n17114 & ~n17115;
  assign n17686 = po2  & n17685;
  assign n17687 = ~n17120 & ~n17686;
  assign n17688 = n17120 & n17686;
  assign n17689 = ~n17687 & ~n17688;
  assign n17690 = ~n17684 & ~n17689;
  assign n17691 = ~n17683 & ~n17690;
  assign n17692 = po31  & ~n17691;
  assign n17693 = ~po31  & n17691;
  assign n17694 = ~n17123 & ~n17124;
  assign n17695 = po2  & n17694;
  assign n17696 = ~n17129 & ~n17695;
  assign n17697 = n17129 & n17695;
  assign n17698 = ~n17696 & ~n17697;
  assign n17699 = ~n17693 & ~n17698;
  assign n17700 = ~n17692 & ~n17699;
  assign n17701 = po32  & ~n17700;
  assign n17702 = ~po32  & n17700;
  assign n17703 = ~n17132 & ~n17133;
  assign n17704 = po2  & n17703;
  assign n17705 = ~n17138 & ~n17704;
  assign n17706 = n17138 & n17704;
  assign n17707 = ~n17705 & ~n17706;
  assign n17708 = ~n17702 & ~n17707;
  assign n17709 = ~n17701 & ~n17708;
  assign n17710 = po33  & ~n17709;
  assign n17711 = ~po33  & n17709;
  assign n17712 = ~n17141 & ~n17142;
  assign n17713 = po2  & n17712;
  assign n17714 = ~n17147 & ~n17713;
  assign n17715 = n17147 & n17713;
  assign n17716 = ~n17714 & ~n17715;
  assign n17717 = ~n17711 & ~n17716;
  assign n17718 = ~n17710 & ~n17717;
  assign n17719 = po34  & ~n17718;
  assign n17720 = ~po34  & n17718;
  assign n17721 = ~n17150 & ~n17151;
  assign n17722 = po2  & n17721;
  assign n17723 = ~n17156 & ~n17722;
  assign n17724 = n17156 & n17722;
  assign n17725 = ~n17723 & ~n17724;
  assign n17726 = ~n17720 & ~n17725;
  assign n17727 = ~n17719 & ~n17726;
  assign n17728 = po35  & ~n17727;
  assign n17729 = ~po35  & n17727;
  assign n17730 = ~n17159 & ~n17160;
  assign n17731 = po2  & n17730;
  assign n17732 = ~n17165 & ~n17731;
  assign n17733 = n17165 & n17731;
  assign n17734 = ~n17732 & ~n17733;
  assign n17735 = ~n17729 & ~n17734;
  assign n17736 = ~n17728 & ~n17735;
  assign n17737 = po36  & ~n17736;
  assign n17738 = ~po36  & n17736;
  assign n17739 = ~n17168 & ~n17169;
  assign n17740 = po2  & n17739;
  assign n17741 = ~n17174 & ~n17740;
  assign n17742 = n17174 & n17740;
  assign n17743 = ~n17741 & ~n17742;
  assign n17744 = ~n17738 & ~n17743;
  assign n17745 = ~n17737 & ~n17744;
  assign n17746 = po37  & ~n17745;
  assign n17747 = ~po37  & n17745;
  assign n17748 = ~n17177 & ~n17178;
  assign n17749 = po2  & n17748;
  assign n17750 = ~n17183 & ~n17749;
  assign n17751 = n17183 & n17749;
  assign n17752 = ~n17750 & ~n17751;
  assign n17753 = ~n17747 & ~n17752;
  assign n17754 = ~n17746 & ~n17753;
  assign n17755 = po38  & ~n17754;
  assign n17756 = ~po38  & n17754;
  assign n17757 = ~n17186 & ~n17187;
  assign n17758 = po2  & n17757;
  assign n17759 = ~n17192 & ~n17758;
  assign n17760 = n17192 & n17758;
  assign n17761 = ~n17759 & ~n17760;
  assign n17762 = ~n17756 & ~n17761;
  assign n17763 = ~n17755 & ~n17762;
  assign n17764 = po39  & ~n17763;
  assign n17765 = ~po39  & n17763;
  assign n17766 = ~n17195 & ~n17196;
  assign n17767 = po2  & n17766;
  assign n17768 = ~n17201 & ~n17767;
  assign n17769 = n17201 & n17767;
  assign n17770 = ~n17768 & ~n17769;
  assign n17771 = ~n17765 & ~n17770;
  assign n17772 = ~n17764 & ~n17771;
  assign n17773 = po40  & ~n17772;
  assign n17774 = ~po40  & n17772;
  assign n17775 = ~n17204 & ~n17205;
  assign n17776 = po2  & n17775;
  assign n17777 = ~n17210 & ~n17776;
  assign n17778 = n17210 & n17776;
  assign n17779 = ~n17777 & ~n17778;
  assign n17780 = ~n17774 & ~n17779;
  assign n17781 = ~n17773 & ~n17780;
  assign n17782 = po41  & ~n17781;
  assign n17783 = ~po41  & n17781;
  assign n17784 = ~n17213 & ~n17214;
  assign n17785 = po2  & n17784;
  assign n17786 = ~n17219 & ~n17785;
  assign n17787 = n17219 & n17785;
  assign n17788 = ~n17786 & ~n17787;
  assign n17789 = ~n17783 & ~n17788;
  assign n17790 = ~n17782 & ~n17789;
  assign n17791 = po42  & ~n17790;
  assign n17792 = ~po42  & n17790;
  assign n17793 = ~n17222 & ~n17223;
  assign n17794 = po2  & n17793;
  assign n17795 = ~n17228 & ~n17794;
  assign n17796 = n17228 & n17794;
  assign n17797 = ~n17795 & ~n17796;
  assign n17798 = ~n17792 & ~n17797;
  assign n17799 = ~n17791 & ~n17798;
  assign n17800 = po43  & ~n17799;
  assign n17801 = ~po43  & n17799;
  assign n17802 = ~n17231 & ~n17232;
  assign n17803 = po2  & n17802;
  assign n17804 = ~n17237 & ~n17803;
  assign n17805 = n17237 & n17803;
  assign n17806 = ~n17804 & ~n17805;
  assign n17807 = ~n17801 & ~n17806;
  assign n17808 = ~n17800 & ~n17807;
  assign n17809 = po44  & ~n17808;
  assign n17810 = ~po44  & n17808;
  assign n17811 = ~n17240 & ~n17241;
  assign n17812 = po2  & n17811;
  assign n17813 = ~n17246 & ~n17812;
  assign n17814 = n17246 & n17812;
  assign n17815 = ~n17813 & ~n17814;
  assign n17816 = ~n17810 & ~n17815;
  assign n17817 = ~n17809 & ~n17816;
  assign n17818 = po45  & ~n17817;
  assign n17819 = ~po45  & n17817;
  assign n17820 = ~n17249 & ~n17250;
  assign n17821 = po2  & n17820;
  assign n17822 = ~n17255 & ~n17821;
  assign n17823 = n17255 & n17821;
  assign n17824 = ~n17822 & ~n17823;
  assign n17825 = ~n17819 & ~n17824;
  assign n17826 = ~n17818 & ~n17825;
  assign n17827 = po46  & ~n17826;
  assign n17828 = ~po46  & n17826;
  assign n17829 = ~n17258 & ~n17259;
  assign n17830 = po2  & n17829;
  assign n17831 = ~n17264 & ~n17830;
  assign n17832 = n17264 & n17830;
  assign n17833 = ~n17831 & ~n17832;
  assign n17834 = ~n17828 & ~n17833;
  assign n17835 = ~n17827 & ~n17834;
  assign n17836 = po47  & ~n17835;
  assign n17837 = ~po47  & n17835;
  assign n17838 = ~n17267 & ~n17268;
  assign n17839 = po2  & n17838;
  assign n17840 = ~n17273 & ~n17839;
  assign n17841 = n17273 & n17839;
  assign n17842 = ~n17840 & ~n17841;
  assign n17843 = ~n17837 & ~n17842;
  assign n17844 = ~n17836 & ~n17843;
  assign n17845 = po48  & ~n17844;
  assign n17846 = ~po48  & n17844;
  assign n17847 = ~n17276 & ~n17277;
  assign n17848 = po2  & n17847;
  assign n17849 = ~n17282 & ~n17848;
  assign n17850 = n17282 & n17848;
  assign n17851 = ~n17849 & ~n17850;
  assign n17852 = ~n17846 & ~n17851;
  assign n17853 = ~n17845 & ~n17852;
  assign n17854 = po49  & ~n17853;
  assign n17855 = ~po49  & n17853;
  assign n17856 = ~n17285 & ~n17286;
  assign n17857 = po2  & n17856;
  assign n17858 = ~n17291 & ~n17857;
  assign n17859 = n17291 & n17857;
  assign n17860 = ~n17858 & ~n17859;
  assign n17861 = ~n17855 & ~n17860;
  assign n17862 = ~n17854 & ~n17861;
  assign n17863 = po50  & ~n17862;
  assign n17864 = ~po50  & n17862;
  assign n17865 = ~n17294 & ~n17295;
  assign n17866 = po2  & n17865;
  assign n17867 = ~n17300 & ~n17866;
  assign n17868 = n17300 & n17866;
  assign n17869 = ~n17867 & ~n17868;
  assign n17870 = ~n17864 & ~n17869;
  assign n17871 = ~n17863 & ~n17870;
  assign n17872 = po51  & ~n17871;
  assign n17873 = ~po51  & n17871;
  assign n17874 = ~n17303 & ~n17304;
  assign n17875 = po2  & n17874;
  assign n17876 = ~n17309 & ~n17875;
  assign n17877 = n17309 & n17875;
  assign n17878 = ~n17876 & ~n17877;
  assign n17879 = ~n17873 & ~n17878;
  assign n17880 = ~n17872 & ~n17879;
  assign n17881 = po52  & ~n17880;
  assign n17882 = ~po52  & n17880;
  assign n17883 = ~n17312 & ~n17313;
  assign n17884 = po2  & n17883;
  assign n17885 = ~n17318 & ~n17884;
  assign n17886 = n17318 & n17884;
  assign n17887 = ~n17885 & ~n17886;
  assign n17888 = ~n17882 & ~n17887;
  assign n17889 = ~n17881 & ~n17888;
  assign n17890 = po53  & ~n17889;
  assign n17891 = ~po53  & n17889;
  assign n17892 = ~n17321 & ~n17322;
  assign n17893 = po2  & n17892;
  assign n17894 = ~n17327 & ~n17893;
  assign n17895 = n17327 & n17893;
  assign n17896 = ~n17894 & ~n17895;
  assign n17897 = ~n17891 & ~n17896;
  assign n17898 = ~n17890 & ~n17897;
  assign n17899 = po54  & ~n17898;
  assign n17900 = ~po54  & n17898;
  assign n17901 = ~n17330 & ~n17331;
  assign n17902 = po2  & n17901;
  assign n17903 = ~n17336 & ~n17902;
  assign n17904 = n17336 & n17902;
  assign n17905 = ~n17903 & ~n17904;
  assign n17906 = ~n17900 & ~n17905;
  assign n17907 = ~n17899 & ~n17906;
  assign n17908 = po55  & ~n17907;
  assign n17909 = ~po55  & n17907;
  assign n17910 = ~n17339 & ~n17340;
  assign n17911 = po2  & n17910;
  assign n17912 = ~n17345 & ~n17911;
  assign n17913 = n17345 & n17911;
  assign n17914 = ~n17912 & ~n17913;
  assign n17915 = ~n17909 & ~n17914;
  assign n17916 = ~n17908 & ~n17915;
  assign n17917 = po56  & ~n17916;
  assign n17918 = ~po56  & n17916;
  assign n17919 = ~n17348 & ~n17349;
  assign n17920 = po2  & n17919;
  assign n17921 = ~n17354 & ~n17920;
  assign n17922 = n17354 & n17920;
  assign n17923 = ~n17921 & ~n17922;
  assign n17924 = ~n17918 & ~n17923;
  assign n17925 = ~n17917 & ~n17924;
  assign n17926 = po57  & ~n17925;
  assign n17927 = ~po57  & n17925;
  assign n17928 = ~n17357 & ~n17358;
  assign n17929 = po2  & n17928;
  assign n17930 = ~n17363 & ~n17929;
  assign n17931 = n17363 & n17929;
  assign n17932 = ~n17930 & ~n17931;
  assign n17933 = ~n17927 & ~n17932;
  assign n17934 = ~n17926 & ~n17933;
  assign n17935 = po58  & ~n17934;
  assign n17936 = ~po58  & n17934;
  assign n17937 = ~n17366 & ~n17367;
  assign n17938 = po2  & n17937;
  assign n17939 = ~n17372 & ~n17938;
  assign n17940 = n17372 & n17938;
  assign n17941 = ~n17939 & ~n17940;
  assign n17942 = ~n17936 & ~n17941;
  assign n17943 = ~n17935 & ~n17942;
  assign n17944 = po59  & ~n17943;
  assign n17945 = ~po59  & n17943;
  assign n17946 = ~n17375 & ~n17376;
  assign n17947 = po2  & n17946;
  assign n17948 = ~n17381 & ~n17947;
  assign n17949 = n17381 & n17947;
  assign n17950 = ~n17948 & ~n17949;
  assign n17951 = ~n17945 & ~n17950;
  assign n17952 = ~n17944 & ~n17951;
  assign n17953 = po60  & ~n17952;
  assign n17954 = ~po60  & n17952;
  assign n17955 = ~n17384 & ~n17385;
  assign n17956 = po2  & n17955;
  assign n17957 = ~n17390 & ~n17956;
  assign n17958 = n17390 & n17956;
  assign n17959 = ~n17957 & ~n17958;
  assign n17960 = ~n17954 & ~n17959;
  assign n17961 = ~n17953 & ~n17960;
  assign n17962 = po61  & ~n17961;
  assign n17963 = ~n17393 & ~n17399;
  assign n17964 = po2  & n17963;
  assign n17965 = ~n17398 & ~n17964;
  assign n17966 = n17398 & n17964;
  assign n17967 = ~n17965 & ~n17966;
  assign n17968 = ~po61  & n17961;
  assign n17969 = ~n17967 & ~n17968;
  assign n17970 = ~n17962 & ~n17969;
  assign n17971 = po62  & ~n17970;
  assign n17972 = ~po62  & n17970;
  assign n17973 = ~n17411 & ~n17412;
  assign n17974 = po2  & n17973;
  assign n17975 = ~n17417 & ~n17974;
  assign n17976 = n17417 & n17974;
  assign n17977 = ~n17975 & ~n17976;
  assign n17978 = ~n17436 & ~n17972;
  assign n17979 = ~n17971 & ~n17978;
  assign n17980 = n17977 & n17979;
  assign n17981 = ~n17977 & ~n17979;
  assign n17982 = n17421 & ~n17430;
  assign n17983 = ~n17420 & ~n17982;
  assign n17984 = n17981 & n17983;
  assign n17985 = ~po63  & ~n17984;
  assign n17986 = ~n17408 & ~n17430;
  assign n17987 = n17419 & ~n17986;
  assign n17988 = po63  & ~n17421;
  assign n17989 = ~n17987 & n17988;
  assign n17990 = ~n17985 & ~n17989;
  assign po1  = n17980 | ~n17990;
  assign n17992 = ~n17971 & ~n17972;
  assign n17993 = po1  & n17992;
  assign n17994 = ~n17436 & ~n17993;
  assign n17995 = n17436 & n17993;
  assign n17996 = ~n17994 & ~n17995;
  assign n17997 = ~n17935 & ~n17936;
  assign n17998 = po1  & n17997;
  assign n17999 = ~n17941 & ~n17998;
  assign n18000 = n17941 & n17998;
  assign n18001 = ~n17999 & ~n18000;
  assign n18002 = ~pi0  & ~pi1 ;
  assign n18003 = ~pi2  & ~n18002;
  assign n18004 = pi2  & ~po1 ;
  assign n18005 = ~pi2  & po1 ;
  assign n18006 = ~pi3  & n18005;
  assign n18007 = pi3  & ~n18005;
  assign n18008 = ~n18006 & ~n18007;
  assign n18009 = ~po2  & ~n18008;
  assign n18010 = ~n18003 & ~n18004;
  assign n18011 = ~n18009 & n18010;
  assign n18012 = po2  & n18008;
  assign n18013 = ~n18011 & ~n18012;
  assign n18014 = po2  & ~po1 ;
  assign n18015 = ~n18006 & ~n18014;
  assign n18016 = pi4  & ~n18015;
  assign n18017 = ~pi4  & n18015;
  assign n18018 = ~n18016 & ~n18017;
  assign n18019 = ~po3  & n18018;
  assign n18020 = ~n18013 & ~n18019;
  assign n18021 = po3  & ~n18018;
  assign n18022 = ~n18020 & ~n18021;
  assign n18023 = ~n17441 & ~n17442;
  assign n18024 = po1  & n18023;
  assign n18025 = n17446 & ~n18024;
  assign n18026 = ~n17446 & n18024;
  assign n18027 = ~n18025 & ~n18026;
  assign n18028 = ~po4  & n18027;
  assign n18029 = ~n18022 & ~n18028;
  assign n18030 = po4  & ~n18027;
  assign n18031 = ~n18029 & ~n18030;
  assign n18032 = ~n17449 & ~n17450;
  assign n18033 = po1  & n18032;
  assign n18034 = ~n17455 & ~n18033;
  assign n18035 = n17455 & n18033;
  assign n18036 = ~n18034 & ~n18035;
  assign n18037 = ~po5  & n18036;
  assign n18038 = ~n18031 & ~n18037;
  assign n18039 = po5  & ~n18036;
  assign n18040 = ~n18038 & ~n18039;
  assign n18041 = ~n17458 & ~n17459;
  assign n18042 = po1  & n18041;
  assign n18043 = n17464 & n18042;
  assign n18044 = ~n17464 & ~n18042;
  assign n18045 = ~n18043 & ~n18044;
  assign n18046 = ~po6  & n18045;
  assign n18047 = ~n18040 & ~n18046;
  assign n18048 = po6  & ~n18045;
  assign n18049 = ~n18047 & ~n18048;
  assign n18050 = ~n17467 & ~n17468;
  assign n18051 = po1  & n18050;
  assign n18052 = ~n17473 & ~n18051;
  assign n18053 = n17473 & n18051;
  assign n18054 = ~n18052 & ~n18053;
  assign n18055 = ~po7  & n18054;
  assign n18056 = ~n18049 & ~n18055;
  assign n18057 = po7  & ~n18054;
  assign n18058 = ~n18056 & ~n18057;
  assign n18059 = ~n17476 & ~n17477;
  assign n18060 = po1  & n18059;
  assign n18061 = ~n17482 & ~n18060;
  assign n18062 = n17482 & n18060;
  assign n18063 = ~n18061 & ~n18062;
  assign n18064 = ~po8  & n18063;
  assign n18065 = ~n18058 & ~n18064;
  assign n18066 = po8  & ~n18063;
  assign n18067 = ~n18065 & ~n18066;
  assign n18068 = ~n17485 & ~n17486;
  assign n18069 = po1  & n18068;
  assign n18070 = ~n17491 & ~n18069;
  assign n18071 = n17491 & n18069;
  assign n18072 = ~n18070 & ~n18071;
  assign n18073 = ~po9  & n18072;
  assign n18074 = ~n18067 & ~n18073;
  assign n18075 = po9  & ~n18072;
  assign n18076 = ~n18074 & ~n18075;
  assign n18077 = ~n17494 & ~n17495;
  assign n18078 = po1  & n18077;
  assign n18079 = ~n17500 & ~n18078;
  assign n18080 = n17500 & n18078;
  assign n18081 = ~n18079 & ~n18080;
  assign n18082 = ~po10  & n18081;
  assign n18083 = ~n18076 & ~n18082;
  assign n18084 = po10  & ~n18081;
  assign n18085 = ~n18083 & ~n18084;
  assign n18086 = ~n17503 & ~n17504;
  assign n18087 = po1  & n18086;
  assign n18088 = ~n17509 & ~n18087;
  assign n18089 = n17509 & n18087;
  assign n18090 = ~n18088 & ~n18089;
  assign n18091 = ~po11  & n18090;
  assign n18092 = ~n18085 & ~n18091;
  assign n18093 = po11  & ~n18090;
  assign n18094 = ~n18092 & ~n18093;
  assign n18095 = ~n17512 & ~n17513;
  assign n18096 = po1  & n18095;
  assign n18097 = ~n17518 & ~n18096;
  assign n18098 = n17518 & n18096;
  assign n18099 = ~n18097 & ~n18098;
  assign n18100 = ~po12  & n18099;
  assign n18101 = ~n18094 & ~n18100;
  assign n18102 = po12  & ~n18099;
  assign n18103 = ~n18101 & ~n18102;
  assign n18104 = ~n17521 & ~n17522;
  assign n18105 = po1  & n18104;
  assign n18106 = ~n17527 & ~n18105;
  assign n18107 = n17527 & n18105;
  assign n18108 = ~n18106 & ~n18107;
  assign n18109 = ~po13  & n18108;
  assign n18110 = ~n18103 & ~n18109;
  assign n18111 = po13  & ~n18108;
  assign n18112 = ~n18110 & ~n18111;
  assign n18113 = ~n17530 & ~n17531;
  assign n18114 = po1  & n18113;
  assign n18115 = ~n17536 & ~n18114;
  assign n18116 = n17536 & n18114;
  assign n18117 = ~n18115 & ~n18116;
  assign n18118 = ~po14  & n18117;
  assign n18119 = ~n18112 & ~n18118;
  assign n18120 = po14  & ~n18117;
  assign n18121 = ~n18119 & ~n18120;
  assign n18122 = ~n17539 & ~n17540;
  assign n18123 = po1  & n18122;
  assign n18124 = ~n17545 & ~n18123;
  assign n18125 = n17545 & n18123;
  assign n18126 = ~n18124 & ~n18125;
  assign n18127 = ~po15  & n18126;
  assign n18128 = ~n18121 & ~n18127;
  assign n18129 = po15  & ~n18126;
  assign n18130 = ~n18128 & ~n18129;
  assign n18131 = ~n17548 & ~n17549;
  assign n18132 = po1  & n18131;
  assign n18133 = ~n17554 & ~n18132;
  assign n18134 = n17554 & n18132;
  assign n18135 = ~n18133 & ~n18134;
  assign n18136 = ~po16  & n18135;
  assign n18137 = ~n18130 & ~n18136;
  assign n18138 = po16  & ~n18135;
  assign n18139 = ~n18137 & ~n18138;
  assign n18140 = ~n17557 & ~n17558;
  assign n18141 = po1  & n18140;
  assign n18142 = ~n17563 & ~n18141;
  assign n18143 = n17563 & n18141;
  assign n18144 = ~n18142 & ~n18143;
  assign n18145 = ~po17  & n18144;
  assign n18146 = ~n18139 & ~n18145;
  assign n18147 = po17  & ~n18144;
  assign n18148 = ~n18146 & ~n18147;
  assign n18149 = ~n17566 & ~n17567;
  assign n18150 = po1  & n18149;
  assign n18151 = ~n17572 & ~n18150;
  assign n18152 = n17572 & n18150;
  assign n18153 = ~n18151 & ~n18152;
  assign n18154 = ~po18  & n18153;
  assign n18155 = ~n18148 & ~n18154;
  assign n18156 = po18  & ~n18153;
  assign n18157 = ~n18155 & ~n18156;
  assign n18158 = ~n17575 & ~n17576;
  assign n18159 = po1  & n18158;
  assign n18160 = ~n17581 & ~n18159;
  assign n18161 = n17581 & n18159;
  assign n18162 = ~n18160 & ~n18161;
  assign n18163 = ~po19  & n18162;
  assign n18164 = ~n18157 & ~n18163;
  assign n18165 = po19  & ~n18162;
  assign n18166 = ~n18164 & ~n18165;
  assign n18167 = ~n17584 & ~n17585;
  assign n18168 = po1  & n18167;
  assign n18169 = ~n17590 & ~n18168;
  assign n18170 = n17590 & n18168;
  assign n18171 = ~n18169 & ~n18170;
  assign n18172 = ~po20  & n18171;
  assign n18173 = ~n18166 & ~n18172;
  assign n18174 = po20  & ~n18171;
  assign n18175 = ~n18173 & ~n18174;
  assign n18176 = ~n17593 & ~n17594;
  assign n18177 = po1  & n18176;
  assign n18178 = ~n17599 & ~n18177;
  assign n18179 = n17599 & n18177;
  assign n18180 = ~n18178 & ~n18179;
  assign n18181 = ~po21  & n18180;
  assign n18182 = ~n18175 & ~n18181;
  assign n18183 = po21  & ~n18180;
  assign n18184 = ~n18182 & ~n18183;
  assign n18185 = ~n17602 & ~n17603;
  assign n18186 = po1  & n18185;
  assign n18187 = ~n17608 & ~n18186;
  assign n18188 = n17608 & n18186;
  assign n18189 = ~n18187 & ~n18188;
  assign n18190 = ~po22  & n18189;
  assign n18191 = ~n18184 & ~n18190;
  assign n18192 = po22  & ~n18189;
  assign n18193 = ~n18191 & ~n18192;
  assign n18194 = ~n17611 & ~n17612;
  assign n18195 = po1  & n18194;
  assign n18196 = ~n17617 & ~n18195;
  assign n18197 = n17617 & n18195;
  assign n18198 = ~n18196 & ~n18197;
  assign n18199 = ~po23  & n18198;
  assign n18200 = ~n18193 & ~n18199;
  assign n18201 = po23  & ~n18198;
  assign n18202 = ~n18200 & ~n18201;
  assign n18203 = ~n17620 & ~n17621;
  assign n18204 = po1  & n18203;
  assign n18205 = ~n17626 & ~n18204;
  assign n18206 = n17626 & n18204;
  assign n18207 = ~n18205 & ~n18206;
  assign n18208 = ~po24  & n18207;
  assign n18209 = ~n18202 & ~n18208;
  assign n18210 = po24  & ~n18207;
  assign n18211 = ~n18209 & ~n18210;
  assign n18212 = ~n17629 & ~n17630;
  assign n18213 = po1  & n18212;
  assign n18214 = ~n17635 & ~n18213;
  assign n18215 = n17635 & n18213;
  assign n18216 = ~n18214 & ~n18215;
  assign n18217 = ~po25  & n18216;
  assign n18218 = ~n18211 & ~n18217;
  assign n18219 = po25  & ~n18216;
  assign n18220 = ~n18218 & ~n18219;
  assign n18221 = ~n17638 & ~n17639;
  assign n18222 = po1  & n18221;
  assign n18223 = ~n17644 & ~n18222;
  assign n18224 = n17644 & n18222;
  assign n18225 = ~n18223 & ~n18224;
  assign n18226 = ~po26  & n18225;
  assign n18227 = ~n18220 & ~n18226;
  assign n18228 = po26  & ~n18225;
  assign n18229 = ~n18227 & ~n18228;
  assign n18230 = ~n17647 & ~n17648;
  assign n18231 = po1  & n18230;
  assign n18232 = ~n17653 & ~n18231;
  assign n18233 = n17653 & n18231;
  assign n18234 = ~n18232 & ~n18233;
  assign n18235 = ~po27  & n18234;
  assign n18236 = ~n18229 & ~n18235;
  assign n18237 = po27  & ~n18234;
  assign n18238 = ~n18236 & ~n18237;
  assign n18239 = ~n17656 & ~n17657;
  assign n18240 = po1  & n18239;
  assign n18241 = ~n17662 & ~n18240;
  assign n18242 = n17662 & n18240;
  assign n18243 = ~n18241 & ~n18242;
  assign n18244 = ~po28  & n18243;
  assign n18245 = ~n18238 & ~n18244;
  assign n18246 = po28  & ~n18243;
  assign n18247 = ~n18245 & ~n18246;
  assign n18248 = ~n17665 & ~n17666;
  assign n18249 = po1  & n18248;
  assign n18250 = ~n17671 & ~n18249;
  assign n18251 = n17671 & n18249;
  assign n18252 = ~n18250 & ~n18251;
  assign n18253 = ~po29  & n18252;
  assign n18254 = ~n18247 & ~n18253;
  assign n18255 = po29  & ~n18252;
  assign n18256 = ~n18254 & ~n18255;
  assign n18257 = ~n17674 & ~n17675;
  assign n18258 = po1  & n18257;
  assign n18259 = ~n17680 & ~n18258;
  assign n18260 = n17680 & n18258;
  assign n18261 = ~n18259 & ~n18260;
  assign n18262 = ~po30  & n18261;
  assign n18263 = ~n18256 & ~n18262;
  assign n18264 = po30  & ~n18261;
  assign n18265 = ~n18263 & ~n18264;
  assign n18266 = ~n17683 & ~n17684;
  assign n18267 = po1  & n18266;
  assign n18268 = ~n17689 & ~n18267;
  assign n18269 = n17689 & n18267;
  assign n18270 = ~n18268 & ~n18269;
  assign n18271 = ~po31  & n18270;
  assign n18272 = ~n18265 & ~n18271;
  assign n18273 = po31  & ~n18270;
  assign n18274 = ~n18272 & ~n18273;
  assign n18275 = ~n17692 & ~n17693;
  assign n18276 = po1  & n18275;
  assign n18277 = ~n17698 & ~n18276;
  assign n18278 = n17698 & n18276;
  assign n18279 = ~n18277 & ~n18278;
  assign n18280 = ~po32  & n18279;
  assign n18281 = ~n18274 & ~n18280;
  assign n18282 = po32  & ~n18279;
  assign n18283 = ~n18281 & ~n18282;
  assign n18284 = ~n17701 & ~n17702;
  assign n18285 = po1  & n18284;
  assign n18286 = ~n17707 & ~n18285;
  assign n18287 = n17707 & n18285;
  assign n18288 = ~n18286 & ~n18287;
  assign n18289 = ~po33  & n18288;
  assign n18290 = ~n18283 & ~n18289;
  assign n18291 = po33  & ~n18288;
  assign n18292 = ~n18290 & ~n18291;
  assign n18293 = ~n17710 & ~n17711;
  assign n18294 = po1  & n18293;
  assign n18295 = ~n17716 & ~n18294;
  assign n18296 = n17716 & n18294;
  assign n18297 = ~n18295 & ~n18296;
  assign n18298 = ~po34  & n18297;
  assign n18299 = ~n18292 & ~n18298;
  assign n18300 = po34  & ~n18297;
  assign n18301 = ~n18299 & ~n18300;
  assign n18302 = ~n17719 & ~n17720;
  assign n18303 = po1  & n18302;
  assign n18304 = ~n17725 & ~n18303;
  assign n18305 = n17725 & n18303;
  assign n18306 = ~n18304 & ~n18305;
  assign n18307 = ~po35  & n18306;
  assign n18308 = ~n18301 & ~n18307;
  assign n18309 = po35  & ~n18306;
  assign n18310 = ~n18308 & ~n18309;
  assign n18311 = ~n17728 & ~n17729;
  assign n18312 = po1  & n18311;
  assign n18313 = ~n17734 & ~n18312;
  assign n18314 = n17734 & n18312;
  assign n18315 = ~n18313 & ~n18314;
  assign n18316 = ~po36  & n18315;
  assign n18317 = ~n18310 & ~n18316;
  assign n18318 = po36  & ~n18315;
  assign n18319 = ~n18317 & ~n18318;
  assign n18320 = ~n17737 & ~n17738;
  assign n18321 = po1  & n18320;
  assign n18322 = ~n17743 & ~n18321;
  assign n18323 = n17743 & n18321;
  assign n18324 = ~n18322 & ~n18323;
  assign n18325 = ~po37  & n18324;
  assign n18326 = ~n18319 & ~n18325;
  assign n18327 = po37  & ~n18324;
  assign n18328 = ~n18326 & ~n18327;
  assign n18329 = ~n17746 & ~n17747;
  assign n18330 = po1  & n18329;
  assign n18331 = ~n17752 & ~n18330;
  assign n18332 = n17752 & n18330;
  assign n18333 = ~n18331 & ~n18332;
  assign n18334 = ~po38  & n18333;
  assign n18335 = ~n18328 & ~n18334;
  assign n18336 = po38  & ~n18333;
  assign n18337 = ~n18335 & ~n18336;
  assign n18338 = ~n17755 & ~n17756;
  assign n18339 = po1  & n18338;
  assign n18340 = ~n17761 & ~n18339;
  assign n18341 = n17761 & n18339;
  assign n18342 = ~n18340 & ~n18341;
  assign n18343 = ~po39  & n18342;
  assign n18344 = ~n18337 & ~n18343;
  assign n18345 = po39  & ~n18342;
  assign n18346 = ~n18344 & ~n18345;
  assign n18347 = ~n17764 & ~n17765;
  assign n18348 = po1  & n18347;
  assign n18349 = ~n17770 & ~n18348;
  assign n18350 = n17770 & n18348;
  assign n18351 = ~n18349 & ~n18350;
  assign n18352 = ~po40  & n18351;
  assign n18353 = ~n18346 & ~n18352;
  assign n18354 = po40  & ~n18351;
  assign n18355 = ~n18353 & ~n18354;
  assign n18356 = ~n17773 & ~n17774;
  assign n18357 = po1  & n18356;
  assign n18358 = ~n17779 & ~n18357;
  assign n18359 = n17779 & n18357;
  assign n18360 = ~n18358 & ~n18359;
  assign n18361 = ~po41  & n18360;
  assign n18362 = ~n18355 & ~n18361;
  assign n18363 = po41  & ~n18360;
  assign n18364 = ~n18362 & ~n18363;
  assign n18365 = ~n17782 & ~n17783;
  assign n18366 = po1  & n18365;
  assign n18367 = ~n17788 & ~n18366;
  assign n18368 = n17788 & n18366;
  assign n18369 = ~n18367 & ~n18368;
  assign n18370 = ~po42  & n18369;
  assign n18371 = ~n18364 & ~n18370;
  assign n18372 = po42  & ~n18369;
  assign n18373 = ~n18371 & ~n18372;
  assign n18374 = ~n17791 & ~n17792;
  assign n18375 = po1  & n18374;
  assign n18376 = ~n17797 & ~n18375;
  assign n18377 = n17797 & n18375;
  assign n18378 = ~n18376 & ~n18377;
  assign n18379 = ~po43  & n18378;
  assign n18380 = ~n18373 & ~n18379;
  assign n18381 = po43  & ~n18378;
  assign n18382 = ~n18380 & ~n18381;
  assign n18383 = ~n17800 & ~n17801;
  assign n18384 = po1  & n18383;
  assign n18385 = ~n17806 & ~n18384;
  assign n18386 = n17806 & n18384;
  assign n18387 = ~n18385 & ~n18386;
  assign n18388 = ~po44  & n18387;
  assign n18389 = ~n18382 & ~n18388;
  assign n18390 = po44  & ~n18387;
  assign n18391 = ~n18389 & ~n18390;
  assign n18392 = ~n17809 & ~n17810;
  assign n18393 = po1  & n18392;
  assign n18394 = ~n17815 & ~n18393;
  assign n18395 = n17815 & n18393;
  assign n18396 = ~n18394 & ~n18395;
  assign n18397 = ~po45  & n18396;
  assign n18398 = ~n18391 & ~n18397;
  assign n18399 = po45  & ~n18396;
  assign n18400 = ~n18398 & ~n18399;
  assign n18401 = ~n17818 & ~n17819;
  assign n18402 = po1  & n18401;
  assign n18403 = ~n17824 & ~n18402;
  assign n18404 = n17824 & n18402;
  assign n18405 = ~n18403 & ~n18404;
  assign n18406 = ~po46  & n18405;
  assign n18407 = ~n18400 & ~n18406;
  assign n18408 = po46  & ~n18405;
  assign n18409 = ~n18407 & ~n18408;
  assign n18410 = ~n17827 & ~n17828;
  assign n18411 = po1  & n18410;
  assign n18412 = ~n17833 & ~n18411;
  assign n18413 = n17833 & n18411;
  assign n18414 = ~n18412 & ~n18413;
  assign n18415 = ~po47  & n18414;
  assign n18416 = ~n18409 & ~n18415;
  assign n18417 = po47  & ~n18414;
  assign n18418 = ~n18416 & ~n18417;
  assign n18419 = ~n17836 & ~n17837;
  assign n18420 = po1  & n18419;
  assign n18421 = ~n17842 & ~n18420;
  assign n18422 = n17842 & n18420;
  assign n18423 = ~n18421 & ~n18422;
  assign n18424 = ~po48  & n18423;
  assign n18425 = ~n18418 & ~n18424;
  assign n18426 = po48  & ~n18423;
  assign n18427 = ~n18425 & ~n18426;
  assign n18428 = ~n17845 & ~n17846;
  assign n18429 = po1  & n18428;
  assign n18430 = ~n17851 & ~n18429;
  assign n18431 = n17851 & n18429;
  assign n18432 = ~n18430 & ~n18431;
  assign n18433 = ~po49  & n18432;
  assign n18434 = ~n18427 & ~n18433;
  assign n18435 = po49  & ~n18432;
  assign n18436 = ~n18434 & ~n18435;
  assign n18437 = ~n17854 & ~n17855;
  assign n18438 = po1  & n18437;
  assign n18439 = ~n17860 & ~n18438;
  assign n18440 = n17860 & n18438;
  assign n18441 = ~n18439 & ~n18440;
  assign n18442 = ~po50  & n18441;
  assign n18443 = ~n18436 & ~n18442;
  assign n18444 = po50  & ~n18441;
  assign n18445 = ~n18443 & ~n18444;
  assign n18446 = ~n17863 & ~n17864;
  assign n18447 = po1  & n18446;
  assign n18448 = ~n17869 & ~n18447;
  assign n18449 = n17869 & n18447;
  assign n18450 = ~n18448 & ~n18449;
  assign n18451 = ~po51  & n18450;
  assign n18452 = ~n18445 & ~n18451;
  assign n18453 = po51  & ~n18450;
  assign n18454 = ~n18452 & ~n18453;
  assign n18455 = ~n17872 & ~n17873;
  assign n18456 = po1  & n18455;
  assign n18457 = ~n17878 & ~n18456;
  assign n18458 = n17878 & n18456;
  assign n18459 = ~n18457 & ~n18458;
  assign n18460 = ~po52  & n18459;
  assign n18461 = ~n18454 & ~n18460;
  assign n18462 = po52  & ~n18459;
  assign n18463 = ~n18461 & ~n18462;
  assign n18464 = ~n17881 & ~n17882;
  assign n18465 = po1  & n18464;
  assign n18466 = ~n17887 & ~n18465;
  assign n18467 = n17887 & n18465;
  assign n18468 = ~n18466 & ~n18467;
  assign n18469 = ~po53  & n18468;
  assign n18470 = ~n18463 & ~n18469;
  assign n18471 = po53  & ~n18468;
  assign n18472 = ~n18470 & ~n18471;
  assign n18473 = ~n17890 & ~n17891;
  assign n18474 = po1  & n18473;
  assign n18475 = ~n17896 & ~n18474;
  assign n18476 = n17896 & n18474;
  assign n18477 = ~n18475 & ~n18476;
  assign n18478 = ~po54  & n18477;
  assign n18479 = ~n18472 & ~n18478;
  assign n18480 = po54  & ~n18477;
  assign n18481 = ~n18479 & ~n18480;
  assign n18482 = ~n17899 & ~n17900;
  assign n18483 = po1  & n18482;
  assign n18484 = ~n17905 & ~n18483;
  assign n18485 = n17905 & n18483;
  assign n18486 = ~n18484 & ~n18485;
  assign n18487 = ~po55  & n18486;
  assign n18488 = ~n18481 & ~n18487;
  assign n18489 = po55  & ~n18486;
  assign n18490 = ~n18488 & ~n18489;
  assign n18491 = ~n17908 & ~n17909;
  assign n18492 = po1  & n18491;
  assign n18493 = ~n17914 & ~n18492;
  assign n18494 = n17914 & n18492;
  assign n18495 = ~n18493 & ~n18494;
  assign n18496 = ~po56  & n18495;
  assign n18497 = ~n18490 & ~n18496;
  assign n18498 = po56  & ~n18495;
  assign n18499 = ~n18497 & ~n18498;
  assign n18500 = ~n17917 & ~n17918;
  assign n18501 = po1  & n18500;
  assign n18502 = ~n17923 & ~n18501;
  assign n18503 = n17923 & n18501;
  assign n18504 = ~n18502 & ~n18503;
  assign n18505 = ~po57  & n18504;
  assign n18506 = ~n18499 & ~n18505;
  assign n18507 = po57  & ~n18504;
  assign n18508 = ~n18506 & ~n18507;
  assign n18509 = ~n17926 & ~n17927;
  assign n18510 = po1  & n18509;
  assign n18511 = ~n17932 & ~n18510;
  assign n18512 = n17932 & n18510;
  assign n18513 = ~n18511 & ~n18512;
  assign n18514 = ~po58  & n18513;
  assign n18515 = ~n18508 & ~n18514;
  assign n18516 = po58  & ~n18513;
  assign n18517 = ~n18515 & ~n18516;
  assign n18518 = n18001 & n18517;
  assign n18519 = ~n18001 & ~n18517;
  assign n18520 = ~po59  & ~n18519;
  assign n18521 = ~n17944 & ~n17945;
  assign n18522 = po1  & n18521;
  assign n18523 = ~n17950 & ~n18522;
  assign n18524 = n17950 & n18522;
  assign n18525 = ~n18523 & ~n18524;
  assign n18526 = ~po60  & n18525;
  assign n18527 = ~n18518 & ~n18526;
  assign n18528 = ~n18520 & n18527;
  assign n18529 = po60  & ~n18525;
  assign n18530 = ~n18528 & ~n18529;
  assign n18531 = ~n17953 & ~n17954;
  assign n18532 = po1  & n18531;
  assign n18533 = ~n17959 & ~n18532;
  assign n18534 = n17959 & n18532;
  assign n18535 = ~n18533 & ~n18534;
  assign n18536 = ~po61  & n18535;
  assign n18537 = ~n18530 & ~n18536;
  assign n18538 = po61  & ~n18535;
  assign n18539 = ~n18537 & ~n18538;
  assign n18540 = ~n17962 & ~n17968;
  assign n18541 = po1  & n18540;
  assign n18542 = ~n17967 & ~n18541;
  assign n18543 = n17967 & n18541;
  assign n18544 = ~n18542 & ~n18543;
  assign n18545 = ~po62  & n18544;
  assign n18546 = ~n18539 & ~n18545;
  assign n18547 = po62  & ~n18544;
  assign n18548 = ~n18546 & ~n18547;
  assign n18549 = n17996 & n18548;
  assign n18550 = n17981 & ~n17990;
  assign n18551 = ~n17980 & ~n18550;
  assign n18552 = ~n17996 & n18551;
  assign n18553 = ~n18548 & n18552;
  assign n18554 = ~po63  & ~n18553;
  assign n18555 = ~n17977 & ~n17990;
  assign n18556 = n17979 & ~n18555;
  assign n18557 = po63  & ~n17981;
  assign n18558 = ~n18556 & n18557;
  assign n18559 = ~n18549 & ~n18558;
  assign po0  = n18554 | ~n18559;
endmodule
