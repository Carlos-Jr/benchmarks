module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 ,
    pi5 , pi6 , pi7 , pi8 , pi9 ,
    pi10 , pi11 , pi12 , pi13 , pi14 ,
    pi15 , pi16 , pi17 , pi18 , pi19 ,
    pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 ,
    pi30 , pi31 , pi32 , pi33 , pi34 ,
    pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 ,
    pi45 , pi46 , pi47 , pi48 , pi49 ,
    pi50 , pi51 , pi52 , pi53 , pi54 ,
    pi55 , pi56 , pi57 , pi58 , pi59 ,
    po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 ,
    po14 , po15 , po16 , po17 ,
    po18 , po19 , po20 , po21 ,
    po22 , po23 , po24 , po25 ,
    po26 , po27 , po28 , po29   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 ,
    pi5 , pi6 , pi7 , pi8 , pi9 ,
    pi10 , pi11 , pi12 , pi13 , pi14 ,
    pi15 , pi16 , pi17 , pi18 , pi19 ,
    pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 ,
    pi30 , pi31 , pi32 , pi33 , pi34 ,
    pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 ,
    pi45 , pi46 , pi47 , pi48 , pi49 ,
    pi50 , pi51 , pi52 , pi53 , pi54 ,
    pi55 , pi56 , pi57 , pi58 , pi59 ;
  output po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 ,
    po14 , po15 , po16 , po17 ,
    po18 , po19 , po20 , po21 ,
    po22 , po23 , po24 , po25 ,
    po26 , po27 , po28 , po29 ;
  wire n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105,
    n106, n107, n108, n109, n110, n111, n112,
    n113, n114, n115, n116, n117, n118, n119,
    n120, n121, n122, n123, n124, n125, n126,
    n127, n128, n129, n130, n131, n132, n133,
    n134, n135, n136, n137, n138, n139, n140,
    n141, n142, n143, n144, n145, n146, n147,
    n148, n149, n150, n151, n152, n153, n154,
    n155, n156, n157, n158, n159, n160, n161,
    n162, n163, n164, n165, n166, n167, n168,
    n169, n170, n171, n172, n173, n174, n175,
    n176, n177, n178, n179, n180, n181, n182,
    n183, n184, n185, n186, n187, n188, n189,
    n190, n191, n192, n193, n194, n195, n196,
    n197, n198, n199, n200, n201, n202, n203,
    n204, n205, n207, n208, n209, n210, n211,
    n212, n213, n214, n215, n216, n217, n218,
    n219, n220, n221, n222, n223, n224, n225,
    n226, n227, n228, n229, n230, n231, n232,
    n233, n234, n235, n236, n237, n238, n239,
    n240, n241, n242, n243, n244, n245, n246,
    n247, n248, n249, n250, n251, n252, n253,
    n254, n255, n256, n257, n258, n259, n260,
    n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274,
    n275, n276, n277, n278, n279, n280, n281,
    n282, n283, n284, n285, n286, n287, n288,
    n289, n290, n291, n292, n293, n294, n295,
    n296, n297, n298, n299, n300, n301, n302,
    n303, n304, n305, n306, n307, n308, n309,
    n310, n311, n312, n313, n314, n315, n316,
    n317, n318, n319, n320, n321, n322, n323,
    n324, n325, n326, n328, n329, n330;
  assign n92 = ~pi9  & ~pi10 ;
  assign n93 = pi11  & ~n92;
  assign n94 = ~pi12  & ~n93;
  assign n95 = ~pi13  & n94;
  assign n96 = pi14  & ~n95;
  assign n97 = pi15  & n96;
  assign n98 = ~pi16  & ~n97;
  assign n99 = pi17  & ~n98;
  assign n100 = ~pi18  & ~n99;
  assign n101 = pi19  & ~n100;
  assign n102 = pi20  & n101;
  assign n103 = ~pi21  & ~n102;
  assign n104 = ~pi22  & n103;
  assign n105 = pi23  & ~n104;
  assign n106 = pi24  & n105;
  assign n107 = pi25  & n106;
  assign n108 = ~pi26  & ~n107;
  assign n109 = pi27  & ~n108;
  assign n110 = pi28  & n109;
  assign n111 = pi29  & n110;
  assign n112 = ~pi11  & n92;
  assign n113 = ~n93 & ~n112;
  assign n114 = pi13  & ~n94;
  assign n115 = ~n95 & ~n114;
  assign n116 = ~pi17  & n98;
  assign n117 = ~n99 & ~n116;
  assign n118 = ~pi15  & ~n96;
  assign n119 = n117 & ~n118;
  assign n120 = ~n115 & n119;
  assign n121 = n113 & n120;
  assign n122 = pi4  & n121;
  assign n123 = pi12  & n93;
  assign n124 = ~n94 & ~n123;
  assign n125 = ~pi14  & n95;
  assign n126 = ~n96 & ~n125;
  assign n127 = pi18  & n99;
  assign n128 = ~n100 & ~n127;
  assign n129 = ~pi25  & ~n106;
  assign n130 = ~n107 & ~n129;
  assign n131 = ~pi19  & n100;
  assign n132 = ~n101 & ~n131;
  assign n133 = pi21  & n102;
  assign n134 = ~n103 & ~n133;
  assign n135 = n132 & ~n134;
  assign n136 = ~pi28  & ~n109;
  assign n137 = ~n110 & ~n136;
  assign n138 = pi22  & ~n103;
  assign n139 = ~n104 & ~n138;
  assign n140 = ~pi24  & ~n105;
  assign n141 = ~n106 & ~n140;
  assign n142 = ~n139 & n141;
  assign n143 = ~pi9  & n142;
  assign n144 = n137 & n143;
  assign n145 = n135 & n144;
  assign n146 = n130 & n145;
  assign n147 = ~n128 & n146;
  assign n148 = pi16  & n97;
  assign n149 = ~n98 & ~n148;
  assign n150 = ~pi27  & n108;
  assign n151 = ~n109 & ~n150;
  assign n152 = ~pi20  & ~n101;
  assign n153 = ~n102 & ~n152;
  assign n154 = ~pi23  & n104;
  assign n155 = ~n105 & ~n154;
  assign n156 = pi26  & n107;
  assign n157 = ~n108 & ~n156;
  assign n158 = pi29  & ~n157;
  assign n159 = n155 & n158;
  assign n160 = n153 & n159;
  assign n161 = n151 & n160;
  assign n162 = ~n149 & n161;
  assign n163 = n147 & n162;
  assign n164 = n126 & n163;
  assign n165 = ~n124 & n164;
  assign n166 = ~n97 & n165;
  assign n167 = pi6  & n166;
  assign n168 = pi2  & n167;
  assign n169 = n122 & n168;
  assign n170 = pi9  & pi10 ;
  assign n171 = ~n92 & ~n170;
  assign n172 = pi3  & ~n171;
  assign n173 = pi1  & n172;
  assign n174 = pi7  & pi8 ;
  assign n175 = pi5  & n174;
  assign n176 = pi0  & n175;
  assign n177 = n173 & n176;
  assign n178 = n169 & n177;
  assign n179 = ~n111 & ~n178;
  assign n180 = n102 & ~n127;
  assign n181 = ~n130 & n180;
  assign n182 = n139 & n181;
  assign n183 = ~n137 & n182;
  assign n184 = n97 & ~n114;
  assign n185 = pi17  & n149;
  assign n186 = ~pi1  & ~pi8 ;
  assign n187 = ~pi6  & n186;
  assign n188 = n124 & n187;
  assign n189 = ~n113 & n188;
  assign n190 = ~pi2  & ~pi3 ;
  assign n191 = ~pi7  & n190;
  assign n192 = ~pi5  & n191;
  assign n193 = ~pi4  & n192;
  assign n194 = n171 & n193;
  assign n195 = n189 & n194;
  assign n196 = n185 & n195;
  assign n197 = n184 & n196;
  assign n198 = n134 & n197;
  assign n199 = ~n155 & n198;
  assign n200 = ~n141 & n199;
  assign n201 = n157 & n200;
  assign n202 = n183 & n201;
  assign n203 = ~n151 & n202;
  assign n204 = pi9  & n203;
  assign n205 = n111 & ~n204;
  assign po0  = n179 | n205;
  assign n207 = ~pi39  & ~pi40 ;
  assign n208 = pi39  & pi40 ;
  assign n209 = ~n207 & ~n208;
  assign n210 = pi37  & pi38 ;
  assign n211 = pi35  & n210;
  assign n212 = pi41  & ~n207;
  assign n213 = ~pi41  & n207;
  assign n214 = ~n212 & ~n213;
  assign n215 = ~pi42  & ~n212;
  assign n216 = ~pi43  & n215;
  assign n217 = pi44  & ~n216;
  assign n218 = ~pi44  & n216;
  assign n219 = ~n217 & ~n218;
  assign n220 = pi45  & n217;
  assign n221 = ~pi46  & ~n220;
  assign n222 = pi47  & ~n221;
  assign n223 = ~pi48  & ~n222;
  assign n224 = pi49  & ~n223;
  assign n225 = pi50  & n224;
  assign n226 = ~pi51  & ~n225;
  assign n227 = pi51  & n225;
  assign n228 = ~n226 & ~n227;
  assign n229 = ~pi52  & n226;
  assign n230 = pi53  & ~n229;
  assign n231 = ~pi53  & n229;
  assign n232 = ~n230 & ~n231;
  assign n233 = pi54  & n230;
  assign n234 = pi55  & n233;
  assign n235 = ~pi56  & ~n234;
  assign n236 = pi57  & ~n235;
  assign n237 = ~pi57  & n235;
  assign n238 = ~n236 & ~n237;
  assign n239 = pi56  & n234;
  assign n240 = ~n235 & ~n239;
  assign n241 = pi30  & ~n240;
  assign n242 = ~pi39  & n241;
  assign n243 = n238 & n242;
  assign n244 = n232 & n243;
  assign n245 = ~pi55  & ~n233;
  assign n246 = ~n234 & ~n245;
  assign n247 = ~pi50  & ~n224;
  assign n248 = ~n225 & ~n247;
  assign n249 = n246 & n248;
  assign n250 = n244 & n249;
  assign n251 = ~pi49  & n223;
  assign n252 = ~n224 & ~n251;
  assign n253 = pi58  & n236;
  assign n254 = ~pi58  & ~n236;
  assign n255 = ~n253 & ~n254;
  assign n256 = pi52  & ~n226;
  assign n257 = ~n229 & ~n256;
  assign n258 = pi59  & ~n257;
  assign n259 = n255 & n258;
  assign n260 = n252 & n259;
  assign n261 = n250 & n260;
  assign n262 = ~n228 & n261;
  assign n263 = pi46  & n220;
  assign n264 = ~n221 & ~n263;
  assign n265 = ~pi54  & ~n230;
  assign n266 = ~n233 & ~n265;
  assign n267 = pi48  & n222;
  assign n268 = ~n223 & ~n267;
  assign n269 = n266 & ~n268;
  assign n270 = ~n264 & n269;
  assign n271 = n262 & n270;
  assign n272 = n219 & n271;
  assign n273 = ~pi47  & n221;
  assign n274 = ~n220 & ~n273;
  assign n275 = pi43  & ~n215;
  assign n276 = ~n216 & ~n275;
  assign n277 = ~pi45  & ~n217;
  assign n278 = ~n222 & ~n277;
  assign n279 = ~n276 & n278;
  assign n280 = n274 & n279;
  assign n281 = n272 & n280;
  assign n282 = n214 & n281;
  assign n283 = pi32  & n282;
  assign n284 = pi42  & n212;
  assign n285 = ~n215 & ~n284;
  assign n286 = pi36  & ~n285;
  assign n287 = pi34  & n286;
  assign n288 = pi31  & n287;
  assign n289 = n283 & n288;
  assign n290 = n211 & n289;
  assign n291 = ~n209 & n290;
  assign n292 = pi33  & n291;
  assign n293 = pi59  & n253;
  assign n294 = ~pi0  & ~pi30 ;
  assign n295 = n293 & ~n294;
  assign n296 = n225 & ~n267;
  assign n297 = ~n246 & n296;
  assign n298 = n257 & n297;
  assign n299 = ~n255 & n298;
  assign n300 = n220 & ~n275;
  assign n301 = pi47  & n264;
  assign n302 = ~pi31  & ~pi38 ;
  assign n303 = ~pi36  & n302;
  assign n304 = n285 & n303;
  assign n305 = ~n214 & n304;
  assign n306 = ~pi32  & ~pi33 ;
  assign n307 = ~pi37  & n306;
  assign n308 = ~pi35  & n307;
  assign n309 = ~pi34  & n308;
  assign n310 = n209 & n309;
  assign n311 = n305 & n310;
  assign n312 = n301 & n311;
  assign n313 = n300 & n312;
  assign n314 = n228 & n313;
  assign n315 = ~n232 & n314;
  assign n316 = ~n266 & n315;
  assign n317 = n240 & n316;
  assign n318 = n299 & n317;
  assign n319 = ~n238 & n318;
  assign n320 = pi39  & n319;
  assign n321 = n293 & ~n320;
  assign n322 = ~n295 & ~n321;
  assign n323 = ~n292 & n322;
  assign n324 = pi0  & ~n293;
  assign n325 = ~n179 & ~n324;
  assign n326 = ~n323 & n325;
  assign po1  = ~n205 & ~n326;
  assign n328 = pi0  & n293;
  assign n329 = pi30  & n328;
  assign n330 = ~n321 & ~n329;
  assign po2  = ~po0  & ~n330;
  assign po3  = 1'b0;
  assign po4  = 1'b0;
  assign po5  = 1'b0;
  assign po6  = 1'b0;
  assign po7  = 1'b0;
  assign po8  = 1'b0;
  assign po9  = 1'b0;
  assign po10  = 1'b0;
  assign po11  = 1'b0;
  assign po12  = 1'b0;
  assign po13  = 1'b0;
  assign po14  = 1'b0;
  assign po15  = 1'b0;
  assign po16  = 1'b0;
  assign po17  = 1'b0;
  assign po18  = 1'b0;
  assign po19  = 1'b0;
  assign po20  = 1'b0;
  assign po21  = 1'b0;
  assign po22  = 1'b0;
  assign po23  = 1'b0;
  assign po24  = 1'b0;
  assign po25  = 1'b0;
  assign po26  = 1'b0;
  assign po27  = 1'b0;
  assign po28  = 1'b0;
  assign po29  = 1'b0;
endmodule
