module i2c ( 
    pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8, pi9,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19,
    pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29,
    pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38, pi39,
    pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48, pi49,
    pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59,
    pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69,
    pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79,
    pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88, pi89,
    pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97, pi98, pi99,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146,
    po0, po1, po2, po3, po4, po5, po6, po7, po8, po9,
    po10, po11, po12, po13, po14, po15, po16, po17, po18, po19,
    po20, po21, po22, po23, po24, po25, po26, po27, po28, po29,
    po30, po31, po32, po33, po34, po35, po36, po37, po38, po39,
    po40, po41, po42, po43, po44, po45, po46, po47, po48, po49,
    po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66, po67, po68, po69,
    po70, po71, po72, po73, po74, po75, po76, po77, po78, po79,
    po80, po81, po82, po83, po84, po85, po86, po87, po88, po89,
    po90, po91, po92, po93, po94, po95, po96, po97, po98, po99,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141  );
  input  pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8,
    pi9, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18,
    pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28,
    pi29, pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38,
    pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48,
    pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58,
    pi59, pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68,
    pi69, pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78,
    pi79, pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88,
    pi89, pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97, pi98,
    pi99, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146;
  output po0, po1, po2, po3, po4, po5, po6, po7, po8, po9,
    po10, po11, po12, po13, po14, po15, po16, po17, po18, po19,
    po20, po21, po22, po23, po24, po25, po26, po27, po28, po29,
    po30, po31, po32, po33, po34, po35, po36, po37, po38, po39,
    po40, po41, po42, po43, po44, po45, po46, po47, po48, po49,
    po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66, po67, po68, po69,
    po70, po71, po72, po73, po74, po75, po76, po77, po78, po79,
    po80, po81, po82, po83, po84, po85, po86, po87, po88, po89,
    po90, po91, po92, po93, po94, po95, po96, po97, po98, po99,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141;
  wire n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332,
    n333, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n370, n371, n372, n373, n374, n375, n376,
    n377, n378, n379, n380, n381, n382, n383,
    n384, n385, n386, n387, n388, n389, n390,
    n391, n392, n393, n394, n395, n396, n397,
    n398, n399, n400, n401, n402, n403, n405,
    n406, n407, n408, n409, n410, n411, n412,
    n413, n414, n416, n417, n418, n419, n420,
    n421, n422, n423, n425, n426, n427, n428,
    n429, n430, n431, n432, n433, n434, n435,
    n436, n437, n439, n440, n441, n442, n443,
    n444, n445, n447, n448, n449, n450, n451,
    n452, n453, n454, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466,
    n468, n469, n470, n471, n472, n473, n475,
    n476, n477, n478, n479, n480, n482, n483,
    n484, n485, n486, n487, n488, n489, n491,
    n492, n493, n494, n495, n496, n497, n499,
    n500, n501, n502, n503, n504, n505, n506,
    n508, n509, n510, n511, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n527, n528, n529, n531,
    n532, n533, n534, n535, n536, n537, n538,
    n540, n541, n542, n543, n544, n545, n547,
    n548, n549, n550, n551, n553, n554, n555,
    n556, n557, n558, n559, n560, n561, n562,
    n563, n565, n566, n567, n568, n569, n570,
    n572, n573, n574, n575, n576, n577, n579,
    n580, n582, n583, n584, n585, n586, n587,
    n588, n589, n590, n591, n592, n593, n594,
    n595, n596, n597, n598, n599, n600, n601,
    n602, n603, n605, n606, n607, n608, n609,
    n610, n611, n612, n613, n614, n615, n616,
    n617, n618, n619, n620, n621, n622, n623,
    n624, n625, n626, n627, n628, n629, n630,
    n631, n632, n633, n634, n635, n636, n637,
    n638, n639, n640, n641, n642, n644, n645,
    n646, n647, n648, n649, n650, n652, n653,
    n654, n655, n656, n657, n658, n659, n660,
    n662, n663, n664, n665, n666, n667, n668,
    n669, n670, n671, n672, n673, n674, n675,
    n676, n677, n678, n679, n680, n681, n682,
    n683, n684, n685, n686, n687, n688, n689,
    n690, n691, n692, n693, n695, n696, n697,
    n698, n699, n700, n701, n702, n703, n704,
    n705, n706, n707, n708, n709, n710, n711,
    n712, n713, n714, n715, n716, n717, n718,
    n719, n720, n721, n723, n724, n725, n726,
    n727, n728, n730, n731, n732, n733, n734,
    n735, n737, n738, n739, n740, n741, n742,
    n744, n745, n746, n747, n748, n749, n751,
    n752, n753, n754, n755, n756, n758, n759,
    n760, n761, n762, n763, n765, n766, n767,
    n768, n769, n770, n772, n773, n774, n775,
    n776, n777, n779, n780, n781, n782, n783,
    n784, n785, n786, n787, n788, n789, n790,
    n791, n792, n793, n794, n796, n797, n798,
    n799, n800, n801, n802, n804, n805, n806,
    n807, n808, n809, n810, n811, n812, n813,
    n814, n815, n816, n817, n818, n819, n820,
    n821, n823, n824, n825, n826, n827, n828,
    n829, n830, n831, n832, n833, n834, n836,
    n837, n838, n839, n840, n841, n842, n843,
    n845, n846, n847, n848, n849, n850, n852,
    n853, n854, n855, n856, n857, n858, n860,
    n861, n862, n863, n864, n865, n866, n867,
    n868, n869, n871, n872, n873, n874, n875,
    n876, n877, n878, n880, n881, n882, n883,
    n884, n885, n886, n887, n889, n890, n891,
    n892, n893, n894, n895, n896, n897, n899,
    n900, n901, n902, n903, n904, n905, n906,
    n907, n908, n910, n911, n912, n913, n914,
    n915, n916, n917, n918, n919, n921, n922,
    n923, n925, n926, n927, n929, n930, n931,
    n935, n937, n938, n939, n940, n941, n942,
    n943, n944, n945, n946, n947, n948, n949,
    n950, n951, n952, n953, n954, n955, n957,
    n958, n959, n960, n961, n962, n963, n964,
    n965, n966, n967, n968, n969, n970, n972,
    n973, n974, n975, n976, n977, n978, n980,
    n981, n982, n983, n984, n985, n986, n987,
    n988, n989, n990, n991, n992, n993, n994,
    n995, n997, n998, n999, n1001, n1002,
    n1004, n1005, n1006, n1007, n1008, n1009,
    n1010, n1011, n1013, n1014, n1015, n1017,
    n1018, n1019, n1021, n1022, n1023, n1025,
    n1026, n1027, n1028, n1029, n1031, n1032,
    n1033, n1035, n1036, n1037, n1039, n1040,
    n1041, n1043, n1044, n1045, n1047, n1048,
    n1049, n1051, n1052, n1053, n1055, n1056,
    n1057, n1059, n1060, n1061, n1063, n1064,
    n1065, n1067, n1068, n1069, n1071, n1072,
    n1073, n1075, n1076, n1077, n1078, n1079,
    n1081, n1082, n1083, n1085, n1086, n1087,
    n1089, n1090, n1091, n1093, n1094, n1095,
    n1097, n1098, n1099, n1100, n1101, n1102,
    n1103, n1104, n1105, n1106, n1107, n1108,
    n1109, n1110, n1111, n1112, n1113, n1114,
    n1116, n1117, n1118, n1120, n1121, n1122,
    n1124, n1125, n1126, n1128, n1129, n1130,
    n1132, n1133, n1134, n1135, n1136, n1138,
    n1139, n1140, n1142, n1143, n1144, n1146,
    n1147, n1148, n1150, n1151, n1152, n1154,
    n1155, n1156, n1158, n1159, n1160, n1161,
    n1162, n1163, n1165, n1166, n1167, n1168,
    n1169, n1170, n1172, n1173, n1174, n1176,
    n1177, n1178, n1180, n1181, n1182, n1184,
    n1185, n1186, n1188, n1189, n1190, n1192,
    n1193, n1194, n1195, n1196, n1197, n1198,
    n1199, n1200, n1201, n1202, n1203, n1204,
    n1205, n1206, n1207, n1208, n1210, n1211,
    n1212, n1213, n1214, n1215, n1216, n1217,
    n1218, n1219, n1220, n1221, n1222, n1223,
    n1225, n1226, n1227, n1228, n1229, n1230,
    n1231, n1232, n1233, n1234, n1235, n1236,
    n1237, n1238, n1240, n1241, n1242, n1243,
    n1244, n1245, n1246, n1247, n1248, n1249,
    n1250, n1251, n1252, n1253, n1255, n1256,
    n1257, n1258, n1259, n1260, n1261, n1262,
    n1263, n1264, n1265, n1266, n1267, n1268,
    n1269, n1270, n1271, n1273, n1274, n1275,
    n1277, n1278, n1279, n1280, n1281, n1282,
    n1283, n1284, n1285, n1286, n1287, n1288,
    n1289, n1290, n1291, n1292, n1293, n1295,
    n1296, n1297, n1298, n1299, n1300, n1301,
    n1302, n1303, n1304, n1305, n1306, n1307,
    n1308, n1309, n1310, n1311, n1313, n1314,
    n1315, n1317, n1318, n1320, n1321, n1322,
    n1323, n1325, n1326, n1327, n1329, n1330,
    n1331, n1332, n1334, n1335, n1336, n1338,
    n1339, n1340, n1343, n1344, n1347, n1348,
    n1350, n1355, n1356, n1358;
  assign n291 = ~pi13 & ~pi14;
  assign n292 = ~pi6 & ~pi12;
  assign n293 = ~pi4 & ~pi19;
  assign n294 = ~pi18 & n293;
  assign n295 = ~pi16 & n294;
  assign n296 = ~pi5 & ~pi22;
  assign n297 = n295 & n296;
  assign n298 = ~pi9 & ~pi11;
  assign n299 = ~pi8 & ~pi21;
  assign n300 = ~pi7 & n299;
  assign n301 = ~pi17 & n298;
  assign n302 = n300 & n301;
  assign n303 = n291 & n292;
  assign n304 = n302 & n303;
  assign n305 = n297 & n304;
  assign n306 = pi54 & ~n305;
  assign n307 = ~pi0 & ~n306;
  assign n308 = ~pi56 & ~n296;
  assign n309 = ~pi7 & ~pi13;
  assign n310 = n299 & n309;
  assign n311 = ~pi14 & n310;
  assign n312 = ~pi10 & n311;
  assign n313 = pi8 & pi21;
  assign n314 = pi7 & ~n299;
  assign n315 = ~pi13 & ~n313;
  assign n316 = ~n314 & n315;
  assign n317 = ~n300 & ~n316;
  assign n318 = ~pi14 & ~n317;
  assign n319 = ~n310 & ~n318;
  assign n320 = ~pi10 & ~n319;
  assign n321 = ~n311 & ~n320;
  assign n322 = ~pi17 & n292;
  assign n323 = n297 & n322;
  assign n324 = ~n312 & n323;
  assign n325 = ~n321 & n324;
  assign n326 = ~n308 & ~n325;
  assign n327 = n298 & ~n326;
  assign n328 = ~pi56 & n296;
  assign n329 = ~n298 & n328;
  assign n330 = ~n327 & ~n329;
  assign n331 = pi54 & ~n330;
  assign n332 = ~n307 & ~n331;
  assign n333 = ~pi3 & ~pi129;
  assign po15 = n332 | ~n333;
  assign n335 = ~pi17 & pi54;
  assign n336 = ~pi5 & ~pi6;
  assign n337 = ~pi10 & ~pi22;
  assign n338 = ~pi14 & n337;
  assign n339 = n309 & n336;
  assign n340 = n338 & n339;
  assign n341 = ~pi11 & n299;
  assign n342 = ~pi12 & n341;
  assign n343 = n295 & n340;
  assign n344 = n342 & n343;
  assign n345 = n335 & ~n344;
  assign n346 = ~pi1 & ~n345;
  assign n347 = ~pi17 & n341;
  assign n348 = ~pi5 & n292;
  assign n349 = n309 & n348;
  assign n350 = pi9 & ~n349;
  assign n351 = ~pi16 & pi54;
  assign n352 = n294 & n351;
  assign n353 = n338 & n352;
  assign n354 = ~pi7 & n348;
  assign n355 = pi13 & n354;
  assign n356 = pi5 & pi6;
  assign n357 = pi12 & ~n336;
  assign n358 = ~pi7 & ~n356;
  assign n359 = ~n357 & n358;
  assign n360 = ~n348 & ~n359;
  assign n361 = ~pi13 & ~n354;
  assign n362 = ~n360 & n361;
  assign n363 = ~pi9 & ~n355;
  assign n364 = ~n362 & n363;
  assign n365 = n347 & ~n350;
  assign n366 = n353 & n365;
  assign n367 = ~n364 & n366;
  assign n368 = ~n346 & ~n367;
  assign po16 = ~n333 | n368;
  assign n370 = ~pi47 & ~pi48;
  assign n371 = ~pi40 & ~pi42;
  assign n372 = ~pi44 & n371;
  assign n373 = ~pi38 & ~pi41;
  assign n374 = ~pi46 & ~pi50;
  assign n375 = n373 & n374;
  assign n376 = n372 & n375;
  assign n377 = ~pi43 & n376;
  assign n378 = n370 & n377;
  assign n379 = pi82 & ~n378;
  assign n380 = ~pi24 & ~pi49;
  assign n381 = ~pi45 & n380;
  assign n382 = ~pi15 & n381;
  assign n383 = n370 & n382;
  assign n384 = ~pi20 & n383;
  assign n385 = pi82 & ~n384;
  assign n386 = ~pi2 & ~pi15;
  assign n387 = ~pi20 & n386;
  assign n388 = ~pi49 & n387;
  assign n389 = pi82 & ~n388;
  assign n390 = ~n385 & ~n389;
  assign n391 = pi82 & ~n376;
  assign n392 = pi122 & pi127;
  assign n393 = n390 & n392;
  assign n394 = ~n391 & ~n393;
  assign n395 = n390 & n394;
  assign n396 = ~n379 & n395;
  assign n397 = ~pi65 & n396;
  assign n398 = pi82 & ~n377;
  assign n399 = ~pi82 & n392;
  assign n400 = ~n398 & ~n399;
  assign n401 = ~n385 & n400;
  assign n402 = pi2 & ~n401;
  assign n403 = ~n397 & ~n402;
  assign po17 = ~pi129 & ~n403;
  assign n405 = pi0 & ~pi113;
  assign n406 = ~pi123 & n405;
  assign n407 = ~pi17 & ~pi18;
  assign n408 = n299 & n407;
  assign n409 = ~pi9 & n337;
  assign n410 = n408 & n409;
  assign n411 = n344 & n410;
  assign n412 = ~pi61 & ~pi118;
  assign n413 = ~n411 & n412;
  assign n414 = ~n406 & ~n413;
  assign po18 = ~pi129 & ~n414;
  assign n416 = pi4 & ~pi54;
  assign n417 = ~pi9 & ~pi14;
  assign n418 = n347 & n352;
  assign n419 = pi10 & ~pi22;
  assign n420 = n417 & n419;
  assign n421 = n349 & n420;
  assign n422 = n418 & n421;
  assign n423 = ~n416 & ~n422;
  assign po19 = n333 & ~n423;
  assign n425 = pi5 & ~pi54;
  assign n426 = ~pi13 & n337;
  assign n427 = n417 & n426;
  assign n428 = ~pi59 & n347;
  assign n429 = n427 & n428;
  assign n430 = n351 & n354;
  assign n431 = ~pi7 & ~pi25;
  assign n432 = ~pi29 & n431;
  assign n433 = n295 & n432;
  assign n434 = pi28 & n430;
  assign n435 = n433 & n434;
  assign n436 = n429 & n435;
  assign n437 = ~n425 & ~n436;
  assign po20 = n333 & ~n437;
  assign n439 = pi6 & ~pi54;
  assign n440 = pi25 & ~pi28;
  assign n441 = ~pi29 & n440;
  assign n442 = n294 & n441;
  assign n443 = n430 & n442;
  assign n444 = n429 & n443;
  assign n445 = ~n439 & ~n444;
  assign po21 = n333 & ~n445;
  assign n447 = pi7 & ~pi54;
  assign n448 = ~pi11 & n354;
  assign n449 = pi8 & ~pi17;
  assign n450 = ~pi21 & n449;
  assign n451 = n352 & n450;
  assign n452 = n427 & n451;
  assign n453 = n448 & n452;
  assign n454 = ~n447 & ~n453;
  assign po22 = n333 & ~n454;
  assign n456 = pi8 & ~pi54;
  assign n457 = n354 & n427;
  assign n458 = n293 & n351;
  assign n459 = ~pi4 & ~pi8;
  assign n460 = ~pi11 & ~pi16;
  assign n461 = n459 & n460;
  assign n462 = n407 & n461;
  assign n463 = pi21 & n458;
  assign n464 = n462 & n463;
  assign n465 = n457 & n464;
  assign n466 = ~n456 & ~n465;
  assign po23 = n333 & ~n466;
  assign n468 = pi9 & ~pi54;
  assign n469 = pi11 & n293;
  assign n470 = n408 & n469;
  assign n471 = n427 & n470;
  assign n472 = n430 & n471;
  assign n473 = ~n468 & ~n472;
  assign po24 = n333 & ~n473;
  assign n475 = pi10 & ~pi54;
  assign n476 = n410 & n458;
  assign n477 = ~pi13 & pi14;
  assign n478 = n448 & n477;
  assign n479 = n476 & n478;
  assign n480 = ~n475 & ~n479;
  assign po25 = n333 & ~n480;
  assign n482 = pi11 & ~pi54;
  assign n483 = ~pi10 & ~pi14;
  assign n484 = pi22 & n483;
  assign n485 = n298 & n484;
  assign n486 = n408 & n458;
  assign n487 = n485 & n486;
  assign n488 = n349 & n487;
  assign n489 = ~n482 & ~n488;
  assign po26 = n333 & ~n489;
  assign n491 = pi12 & ~pi54;
  assign n492 = ~pi9 & ~pi12;
  assign n493 = pi18 & n492;
  assign n494 = n458 & n493;
  assign n495 = n340 & n494;
  assign n496 = n347 & n495;
  assign n497 = ~n491 & ~n496;
  assign po27 = n333 & ~n497;
  assign n499 = pi13 & ~pi54;
  assign n500 = ~pi25 & ~pi28;
  assign n501 = pi29 & pi54;
  assign n502 = ~pi59 & n501;
  assign n503 = n500 & n502;
  assign n504 = n418 & n503;
  assign n505 = n457 & n504;
  assign n506 = ~n499 & ~n505;
  assign po28 = n333 & ~n506;
  assign n508 = pi14 & ~pi54;
  assign n509 = n302 & n353;
  assign n510 = n355 & n509;
  assign n511 = ~n508 & ~n510;
  assign po29 = n333 & ~n511;
  assign n513 = pi15 & n399;
  assign n514 = n378 & n381;
  assign n515 = pi15 & ~n514;
  assign n516 = n377 & ~n387;
  assign n517 = n383 & n516;
  assign n518 = ~n515 & ~n517;
  assign n519 = pi82 & ~n518;
  assign n520 = n378 & n382;
  assign n521 = pi82 & ~n520;
  assign n522 = ~pi70 & ~n392;
  assign n523 = ~n521 & n522;
  assign n524 = ~n513 & ~n523;
  assign n525 = ~n519 & n524;
  assign po30 = ~pi129 & ~n525;
  assign n527 = pi16 & ~pi54;
  assign n528 = pi6 & n367;
  assign n529 = ~n527 & ~n528;
  assign po31 = n333 & ~n529;
  assign n531 = pi17 & ~pi54;
  assign n532 = ~pi28 & pi59;
  assign n533 = n335 & n532;
  assign n534 = n336 & n533;
  assign n535 = n342 & n534;
  assign n536 = n427 & n535;
  assign n537 = n433 & n536;
  assign n538 = ~n531 & ~n537;
  assign po32 = n333 & ~n538;
  assign n540 = pi18 & ~pi54;
  assign n541 = n294 & n457;
  assign n542 = pi16 & n335;
  assign n543 = n341 & n542;
  assign n544 = n541 & n543;
  assign n545 = ~n540 & ~n544;
  assign po33 = n333 & ~n545;
  assign n547 = pi19 & ~pi54;
  assign n548 = pi17 & n351;
  assign n549 = n341 & n548;
  assign n550 = n541 & n549;
  assign n551 = ~n547 & ~n550;
  assign po34 = n333 & ~n551;
  assign n553 = pi20 & n399;
  assign n554 = pi20 & ~n520;
  assign n555 = ~pi20 & n520;
  assign n556 = pi2 & n555;
  assign n557 = ~n554 & ~n556;
  assign n558 = pi82 & ~n557;
  assign n559 = pi82 & ~n555;
  assign n560 = ~pi71 & ~n392;
  assign n561 = ~n559 & n560;
  assign n562 = ~n553 & ~n561;
  assign n563 = ~n558 & n562;
  assign po35 = ~pi129 & ~n563;
  assign n565 = pi21 & ~pi54;
  assign n566 = pi19 & ~pi21;
  assign n567 = pi54 & n566;
  assign n568 = n462 & n567;
  assign n569 = n457 & n568;
  assign n570 = ~n565 & ~n569;
  assign po36 = n333 & ~n570;
  assign n572 = pi22 & ~pi54;
  assign n573 = pi5 & ~pi7;
  assign n574 = ~pi11 & n573;
  assign n575 = n303 & n574;
  assign n576 = n476 & n575;
  assign n577 = ~n572 & ~n576;
  assign po37 = n333 & ~n577;
  assign n579 = ~pi23 & pi55;
  assign n580 = pi61 & ~pi129;
  assign po38 = ~n579 & n580;
  assign n582 = ~pi38 & n372;
  assign n583 = ~pi50 & n582;
  assign n584 = ~pi46 & n583;
  assign n585 = ~pi43 & ~pi47;
  assign n586 = ~pi41 & ~pi45;
  assign n587 = ~pi48 & n586;
  assign n588 = n585 & n587;
  assign n589 = n584 & n588;
  assign n590 = pi24 & pi82;
  assign n591 = n589 & n590;
  assign n592 = ~n389 & n392;
  assign n593 = pi82 & ~n589;
  assign n594 = ~n592 & ~n593;
  assign n595 = ~pi24 & ~n594;
  assign n596 = pi45 & pi82;
  assign n597 = n378 & n596;
  assign n598 = pi63 & ~n392;
  assign n599 = ~n389 & n598;
  assign n600 = ~n379 & n599;
  assign n601 = ~n597 & n600;
  assign n602 = ~pi129 & ~n591;
  assign n603 = ~n601 & n602;
  assign po39 = ~n595 & n603;
  assign n605 = pi25 & ~pi116;
  assign n606 = ~pi39 & ~pi52;
  assign n607 = ~pi51 & n606;
  assign n608 = pi116 & n607;
  assign n609 = ~n605 & ~n608;
  assign n610 = ~pi26 & ~n609;
  assign n611 = pi27 & ~n610;
  assign n612 = ~pi26 & ~pi27;
  assign n613 = pi85 & ~n612;
  assign n614 = pi116 & ~n607;
  assign n615 = pi26 & ~n605;
  assign n616 = ~n614 & n615;
  assign n617 = pi85 & pi116;
  assign n618 = ~pi85 & ~pi110;
  assign n619 = ~pi96 & n618;
  assign n620 = ~n617 & ~n619;
  assign n621 = pi100 & ~n620;
  assign n622 = pi85 & ~n605;
  assign n623 = ~pi27 & ~pi85;
  assign n624 = ~pi95 & ~pi100;
  assign n625 = ~pi97 & n624;
  assign n626 = ~pi110 & ~n625;
  assign n627 = pi25 & ~n626;
  assign n628 = ~pi26 & n623;
  assign n629 = ~n627 & n628;
  assign n630 = ~n622 & ~n629;
  assign n631 = ~n621 & ~n630;
  assign n632 = ~pi53 & ~pi58;
  assign n633 = ~n613 & n632;
  assign n634 = ~n616 & n633;
  assign n635 = ~n611 & n634;
  assign n636 = ~n631 & n635;
  assign n637 = ~pi53 & pi58;
  assign n638 = pi53 & ~pi58;
  assign n639 = ~n637 & ~n638;
  assign n640 = n605 & n628;
  assign n641 = ~n639 & n640;
  assign n642 = ~n636 & ~n641;
  assign po40 = n333 & ~n642;
  assign n644 = ~pi27 & n632;
  assign n645 = ~pi85 & ~n608;
  assign n646 = pi26 & n645;
  assign n647 = pi26 & pi116;
  assign n648 = n621 & ~n647;
  assign n649 = ~n646 & ~n648;
  assign n650 = n333 & n644;
  assign po41 = ~n649 & n650;
  assign n652 = ~pi26 & n333;
  assign n653 = pi27 & n645;
  assign n654 = pi95 & ~pi96;
  assign n655 = n618 & n654;
  assign n656 = ~n617 & ~n655;
  assign n657 = ~pi27 & ~pi100;
  assign n658 = ~n656 & n657;
  assign n659 = ~n653 & ~n658;
  assign n660 = n632 & n652;
  assign po42 = ~n659 & n660;
  assign n662 = ~pi27 & pi28;
  assign n663 = ~pi116 & n662;
  assign n664 = ~pi26 & pi53;
  assign n665 = ~pi85 & n664;
  assign n666 = n663 & n665;
  assign n667 = pi28 & ~pi116;
  assign n668 = ~pi100 & pi116;
  assign n669 = ~n667 & ~n668;
  assign n670 = n612 & ~n669;
  assign n671 = pi85 & ~n670;
  assign n672 = ~n608 & ~n667;
  assign n673 = ~pi27 & ~n672;
  assign n674 = pi26 & ~n673;
  assign n675 = ~pi100 & ~pi110;
  assign n676 = n654 & n675;
  assign n677 = pi28 & ~n626;
  assign n678 = n612 & ~n676;
  assign n679 = ~n677 & n678;
  assign n680 = pi27 & ~n667;
  assign n681 = ~n614 & n680;
  assign n682 = ~n679 & ~n681;
  assign n683 = ~n674 & n682;
  assign n684 = ~pi85 & ~n683;
  assign n685 = ~pi53 & ~n671;
  assign n686 = ~n684 & n685;
  assign n687 = ~n666 & ~n686;
  assign n688 = ~pi58 & ~n687;
  assign n689 = ~pi26 & ~pi53;
  assign n690 = ~pi85 & n689;
  assign n691 = pi58 & n663;
  assign n692 = n690 & n691;
  assign n693 = ~n688 & ~n692;
  assign po43 = n333 & ~n693;
  assign n695 = ~pi116 & ~n639;
  assign n696 = ~n626 & n632;
  assign n697 = ~n695 & ~n696;
  assign n698 = pi29 & ~n697;
  assign n699 = pi58 & pi116;
  assign n700 = ~pi58 & ~pi96;
  assign n701 = ~pi110 & n700;
  assign n702 = n624 & n701;
  assign n703 = ~n699 & ~n702;
  assign n704 = ~pi53 & pi97;
  assign n705 = ~n703 & n704;
  assign n706 = ~n698 & ~n705;
  assign n707 = ~pi27 & ~n706;
  assign n708 = pi29 & ~pi116;
  assign n709 = pi27 & n632;
  assign n710 = n708 & n709;
  assign n711 = ~n707 & ~n710;
  assign n712 = ~pi85 & ~n711;
  assign n713 = pi85 & n708;
  assign n714 = n644 & n713;
  assign n715 = ~n712 & ~n714;
  assign n716 = ~pi26 & ~n715;
  assign n717 = pi26 & ~pi27;
  assign n718 = ~pi85 & n632;
  assign n719 = n717 & n718;
  assign n720 = n708 & n719;
  assign n721 = ~n716 & ~n720;
  assign po44 = n333 & ~n721;
  assign n723 = ~pi88 & pi106;
  assign n724 = ~pi30 & ~pi109;
  assign n725 = ~pi60 & pi109;
  assign n726 = ~n724 & ~n725;
  assign n727 = ~pi106 & ~n726;
  assign n728 = ~pi129 & ~n723;
  assign po45 = ~n727 & n728;
  assign n730 = ~pi89 & pi106;
  assign n731 = ~pi31 & ~pi109;
  assign n732 = ~pi30 & pi109;
  assign n733 = ~n731 & ~n732;
  assign n734 = ~pi106 & ~n733;
  assign n735 = ~pi129 & ~n730;
  assign po46 = ~n734 & n735;
  assign n737 = ~pi99 & pi106;
  assign n738 = ~pi32 & ~pi109;
  assign n739 = ~pi31 & pi109;
  assign n740 = ~n738 & ~n739;
  assign n741 = ~pi106 & ~n740;
  assign n742 = ~pi129 & ~n737;
  assign po47 = ~n741 & n742;
  assign n744 = ~pi90 & pi106;
  assign n745 = ~pi33 & ~pi109;
  assign n746 = ~pi32 & pi109;
  assign n747 = ~n745 & ~n746;
  assign n748 = ~pi106 & ~n747;
  assign n749 = ~pi129 & ~n744;
  assign po48 = ~n748 & n749;
  assign n751 = ~pi91 & pi106;
  assign n752 = ~pi34 & ~pi109;
  assign n753 = ~pi33 & pi109;
  assign n754 = ~n752 & ~n753;
  assign n755 = ~pi106 & ~n754;
  assign n756 = ~pi129 & ~n751;
  assign po49 = ~n755 & n756;
  assign n758 = ~pi92 & pi106;
  assign n759 = ~pi35 & ~pi109;
  assign n760 = ~pi34 & pi109;
  assign n761 = ~n759 & ~n760;
  assign n762 = ~pi106 & ~n761;
  assign n763 = ~pi129 & ~n758;
  assign po50 = ~n762 & n763;
  assign n765 = ~pi98 & pi106;
  assign n766 = ~pi36 & ~pi109;
  assign n767 = ~pi35 & pi109;
  assign n768 = ~n766 & ~n767;
  assign n769 = ~pi106 & ~n768;
  assign n770 = ~pi129 & ~n765;
  assign po51 = ~n769 & n770;
  assign n772 = ~pi93 & pi106;
  assign n773 = ~pi37 & ~pi109;
  assign n774 = ~pi36 & pi109;
  assign n775 = ~n773 & ~n774;
  assign n776 = ~pi106 & ~n775;
  assign n777 = ~pi129 & ~n772;
  assign po52 = ~n776 & n777;
  assign n779 = ~pi44 & pi82;
  assign n780 = n371 & n779;
  assign n781 = pi38 & n780;
  assign n782 = n380 & n387;
  assign n783 = n588 & n782;
  assign n784 = ~pi46 & n783;
  assign n785 = ~pi50 & n784;
  assign n786 = pi82 & ~n785;
  assign n787 = n392 & ~n786;
  assign n788 = pi82 & ~n372;
  assign n789 = ~n787 & ~n788;
  assign n790 = pi74 & ~n786;
  assign n791 = n789 & n790;
  assign n792 = ~pi38 & ~n789;
  assign n793 = ~pi129 & ~n781;
  assign n794 = ~n791 & n793;
  assign po53 = ~n792 & n794;
  assign n796 = ~pi51 & ~pi52;
  assign n797 = pi109 & n796;
  assign n798 = pi39 & ~n797;
  assign n799 = ~pi51 & pi109;
  assign n800 = n606 & n799;
  assign n801 = ~pi106 & ~n800;
  assign n802 = ~n798 & n801;
  assign po54 = ~pi129 & ~n802;
  assign n804 = ~pi42 & ~pi44;
  assign n805 = pi82 & ~n804;
  assign n806 = n381 & n387;
  assign n807 = ~pi48 & n806;
  assign n808 = n585 & n807;
  assign n809 = n375 & n808;
  assign n810 = ~pi40 & n809;
  assign n811 = pi82 & ~n810;
  assign n812 = n392 & ~n811;
  assign n813 = ~n805 & ~n812;
  assign n814 = ~pi40 & ~n813;
  assign n815 = n788 & n804;
  assign n816 = n804 & n809;
  assign n817 = pi82 & ~n816;
  assign n818 = pi73 & ~n392;
  assign n819 = ~n817 & n818;
  assign n820 = ~pi129 & ~n815;
  assign n821 = ~n819 & n820;
  assign po55 = ~n814 & n821;
  assign n823 = n391 & n584;
  assign n824 = n584 & n808;
  assign n825 = pi82 & ~n824;
  assign n826 = pi76 & ~n392;
  assign n827 = ~n825 & n826;
  assign n828 = pi82 & ~n584;
  assign n829 = pi82 & ~n783;
  assign n830 = n392 & ~n829;
  assign n831 = ~n828 & ~n830;
  assign n832 = ~pi41 & ~n831;
  assign n833 = ~pi129 & ~n823;
  assign n834 = ~n827 & n833;
  assign po56 = ~n832 & n834;
  assign n836 = pi42 & n779;
  assign n837 = pi44 & pi82;
  assign n838 = ~n812 & ~n837;
  assign n839 = ~pi42 & ~n838;
  assign n840 = pi72 & ~n811;
  assign n841 = n838 & n840;
  assign n842 = ~pi129 & ~n836;
  assign n843 = ~n839 & n842;
  assign po57 = ~n841 & n843;
  assign n845 = pi43 & n375;
  assign n846 = n780 & n845;
  assign n847 = pi77 & n395;
  assign n848 = ~pi43 & ~n394;
  assign n849 = ~pi129 & ~n846;
  assign n850 = ~n848 & n849;
  assign po58 = ~n847 & n850;
  assign n852 = ~pi42 & n810;
  assign n853 = pi82 & ~n852;
  assign n854 = ~pi67 & ~n392;
  assign n855 = pi44 & n392;
  assign n856 = ~n854 & ~n855;
  assign n857 = ~n853 & n856;
  assign n858 = ~pi129 & ~n837;
  assign po59 = ~n857 & n858;
  assign n860 = n378 & n782;
  assign n861 = pi82 & ~n860;
  assign n862 = pi68 & ~n392;
  assign n863 = ~n861 & n862;
  assign n864 = pi82 & ~n807;
  assign n865 = n392 & ~n864;
  assign n866 = ~n379 & ~n865;
  assign n867 = ~pi45 & ~n866;
  assign n868 = ~pi129 & ~n597;
  assign n869 = ~n863 & n868;
  assign po60 = ~n867 & n869;
  assign n871 = n583 & n828;
  assign n872 = pi82 & ~n583;
  assign n873 = ~n830 & ~n872;
  assign n874 = pi75 & ~n829;
  assign n875 = n873 & n874;
  assign n876 = ~pi46 & ~n873;
  assign n877 = ~pi129 & ~n871;
  assign n878 = ~n875 & n877;
  assign po61 = ~n876 & n878;
  assign n880 = pi47 & pi82;
  assign n881 = n377 & n880;
  assign n882 = ~n398 & ~n865;
  assign n883 = ~pi47 & ~n882;
  assign n884 = pi64 & ~n864;
  assign n885 = n882 & n884;
  assign n886 = ~pi129 & ~n881;
  assign n887 = ~n883 & n886;
  assign po62 = ~n885 & n887;
  assign n889 = n376 & n585;
  assign n890 = n806 & n889;
  assign n891 = pi82 & ~n890;
  assign n892 = pi62 & ~n392;
  assign n893 = ~n891 & n892;
  assign n894 = ~pi48 & ~n866;
  assign n895 = n379 & n889;
  assign n896 = ~pi129 & ~n893;
  assign n897 = ~n895 & n896;
  assign po63 = ~n894 & n897;
  assign n899 = pi49 & n399;
  assign n900 = ~pi24 & n589;
  assign n901 = pi49 & ~n900;
  assign n902 = ~n514 & ~n901;
  assign n903 = n389 & ~n902;
  assign n904 = pi82 & ~n514;
  assign n905 = ~pi69 & ~n392;
  assign n906 = ~n904 & n905;
  assign n907 = ~n899 & ~n906;
  assign n908 = ~n903 & n907;
  assign po64 = ~pi129 & ~n908;
  assign n910 = pi82 & ~n582;
  assign n911 = ~n787 & ~n910;
  assign n912 = ~pi50 & ~n911;
  assign n913 = n582 & n872;
  assign n914 = pi82 & ~n784;
  assign n915 = pi66 & ~n392;
  assign n916 = ~n910 & n915;
  assign n917 = ~n914 & n916;
  assign n918 = ~pi129 & ~n913;
  assign n919 = ~n917 & n918;
  assign po65 = ~n912 & n919;
  assign n921 = pi51 & ~pi109;
  assign n922 = ~pi106 & ~n799;
  assign n923 = ~n921 & n922;
  assign po66 = ~pi129 & ~n923;
  assign n925 = pi52 & ~n799;
  assign n926 = ~pi106 & ~n797;
  assign n927 = ~n925 & n926;
  assign po67 = ~pi129 & ~n927;
  assign n929 = ~pi116 & n638;
  assign n930 = ~n705 & ~n929;
  assign n931 = n623 & n652;
  assign po68 = ~n930 & n931;
  assign po69 = pi129 | n396;
  assign po129 = pi123 | pi129;
  assign n935 = pi114 & ~pi122;
  assign po70 = ~po129 & n935;
  assign n937 = ~pi26 & pi58;
  assign n938 = ~pi58 & n647;
  assign n939 = ~n937 & ~n938;
  assign n940 = pi94 & ~n939;
  assign n941 = pi58 & ~pi116;
  assign n942 = pi37 & ~pi116;
  assign n943 = ~n937 & ~n942;
  assign n944 = ~n941 & ~n943;
  assign n945 = ~n940 & ~n944;
  assign n946 = ~pi53 & ~n945;
  assign n947 = ~pi26 & pi37;
  assign n948 = ~pi58 & n947;
  assign n949 = ~n946 & ~n948;
  assign n950 = ~pi85 & ~n949;
  assign n951 = n632 & n947;
  assign n952 = ~n950 & ~n951;
  assign n953 = ~pi27 & ~n952;
  assign n954 = n718 & n947;
  assign n955 = ~n953 & ~n954;
  assign po71 = n333 & ~n955;
  assign n957 = ~pi116 & n690;
  assign n958 = ~pi53 & ~pi85;
  assign n959 = ~n689 & ~n958;
  assign n960 = ~n665 & n959;
  assign n961 = ~pi58 & ~n960;
  assign n962 = ~n957 & ~n961;
  assign n963 = pi57 & ~n962;
  assign n964 = pi60 & n699;
  assign n965 = n690 & n964;
  assign n966 = ~n963 & ~n965;
  assign n967 = ~pi27 & ~n966;
  assign n968 = pi57 & ~pi58;
  assign n969 = n690 & n968;
  assign n970 = ~n967 & ~n969;
  assign po72 = n333 & ~n970;
  assign n972 = n612 & n941;
  assign n973 = ~pi26 & pi27;
  assign n974 = ~n717 & ~n973;
  assign n975 = ~pi58 & ~n974;
  assign n976 = n608 & n975;
  assign n977 = ~n972 & ~n976;
  assign n978 = n333 & n958;
  assign po73 = ~n977 & n978;
  assign n980 = pi59 & ~n697;
  assign n981 = pi96 & n632;
  assign n982 = n626 & n981;
  assign n983 = ~n980 & ~n982;
  assign n984 = ~pi85 & ~n983;
  assign n985 = pi59 & ~pi116;
  assign n986 = pi85 & n632;
  assign n987 = n985 & n986;
  assign n988 = ~n984 & ~n987;
  assign n989 = ~pi27 & ~n988;
  assign n990 = pi27 & n985;
  assign n991 = n718 & n990;
  assign n992 = ~n989 & ~n991;
  assign n993 = ~pi26 & ~n992;
  assign n994 = n719 & n985;
  assign n995 = ~n993 & ~n994;
  assign po74 = n333 & ~n995;
  assign n997 = ~pi117 & ~pi122;
  assign n998 = pi60 & ~n997;
  assign n999 = pi123 & n997;
  assign po75 = n998 | n999;
  assign n1001 = ~pi114 & ~pi122;
  assign n1002 = pi123 & ~pi129;
  assign po76 = n1001 & n1002;
  assign n1004 = pi136 & ~pi137;
  assign n1005 = pi131 & pi132;
  assign n1006 = pi133 & n1005;
  assign n1007 = ~pi138 & n1006;
  assign n1008 = n1004 & n1007;
  assign n1009 = ~pi62 & ~n1008;
  assign n1010 = pi140 & n1008;
  assign n1011 = ~pi129 & ~n1009;
  assign po77 = n1010 | ~n1011;
  assign n1013 = ~pi63 & ~n1008;
  assign n1014 = pi142 & n1008;
  assign n1015 = ~pi129 & ~n1013;
  assign po78 = n1014 | ~n1015;
  assign n1017 = ~pi64 & ~n1008;
  assign n1018 = pi139 & n1008;
  assign n1019 = ~pi129 & ~n1017;
  assign po79 = n1018 | ~n1019;
  assign n1021 = ~pi65 & ~n1008;
  assign n1022 = pi146 & n1008;
  assign n1023 = ~pi129 & ~n1021;
  assign po80 = n1022 | ~n1023;
  assign n1025 = ~pi136 & ~pi137;
  assign n1026 = n1007 & n1025;
  assign n1027 = ~pi66 & ~n1026;
  assign n1028 = pi143 & n1026;
  assign n1029 = ~pi129 & ~n1027;
  assign po81 = n1028 | ~n1029;
  assign n1031 = ~pi67 & ~n1026;
  assign n1032 = pi139 & n1026;
  assign n1033 = ~pi129 & ~n1031;
  assign po82 = n1032 | ~n1033;
  assign n1035 = ~pi68 & ~n1008;
  assign n1036 = pi141 & n1008;
  assign n1037 = ~pi129 & ~n1035;
  assign po83 = n1036 | ~n1037;
  assign n1039 = ~pi69 & ~n1008;
  assign n1040 = pi143 & n1008;
  assign n1041 = ~pi129 & ~n1039;
  assign po84 = n1040 | ~n1041;
  assign n1043 = ~pi70 & ~n1008;
  assign n1044 = pi144 & n1008;
  assign n1045 = ~pi129 & ~n1043;
  assign po85 = n1044 | ~n1045;
  assign n1047 = ~pi71 & ~n1008;
  assign n1048 = pi145 & n1008;
  assign n1049 = ~pi129 & ~n1047;
  assign po86 = n1048 | ~n1049;
  assign n1051 = ~pi72 & ~n1026;
  assign n1052 = pi140 & n1026;
  assign n1053 = ~pi129 & ~n1051;
  assign po87 = n1052 | ~n1053;
  assign n1055 = ~pi73 & ~n1026;
  assign n1056 = pi141 & n1026;
  assign n1057 = ~pi129 & ~n1055;
  assign po88 = n1056 | ~n1057;
  assign n1059 = ~pi74 & ~n1026;
  assign n1060 = pi142 & n1026;
  assign n1061 = ~pi129 & ~n1059;
  assign po89 = n1060 | ~n1061;
  assign n1063 = ~pi75 & ~n1026;
  assign n1064 = pi144 & n1026;
  assign n1065 = ~pi129 & ~n1063;
  assign po90 = n1064 | ~n1065;
  assign n1067 = ~pi76 & ~n1026;
  assign n1068 = pi145 & n1026;
  assign n1069 = ~pi129 & ~n1067;
  assign po91 = n1068 | ~n1069;
  assign n1071 = ~pi77 & ~n1026;
  assign n1072 = pi146 & n1026;
  assign n1073 = ~pi129 & ~n1071;
  assign po92 = n1072 | ~n1073;
  assign n1075 = ~pi136 & pi137;
  assign n1076 = n1007 & n1075;
  assign n1077 = ~pi78 & ~n1076;
  assign n1078 = ~pi142 & n1076;
  assign n1079 = ~pi129 & ~n1077;
  assign po93 = ~n1078 & n1079;
  assign n1081 = ~pi79 & ~n1076;
  assign n1082 = ~pi143 & n1076;
  assign n1083 = ~pi129 & ~n1081;
  assign po94 = ~n1082 & n1083;
  assign n1085 = ~pi80 & ~n1076;
  assign n1086 = ~pi144 & n1076;
  assign n1087 = ~pi129 & ~n1085;
  assign po95 = ~n1086 & n1087;
  assign n1089 = ~pi81 & ~n1076;
  assign n1090 = ~pi145 & n1076;
  assign n1091 = ~pi129 & ~n1089;
  assign po96 = ~n1090 & n1091;
  assign n1093 = ~pi82 & ~n1076;
  assign n1094 = ~pi146 & n1076;
  assign n1095 = ~pi129 & ~n1093;
  assign po97 = ~n1094 & n1095;
  assign n1097 = pi136 & ~pi138;
  assign n1098 = pi31 & n1097;
  assign n1099 = ~pi87 & ~pi138;
  assign n1100 = pi115 & pi138;
  assign n1101 = ~pi136 & ~n1099;
  assign n1102 = ~n1100 & n1101;
  assign n1103 = ~n1098 & ~n1102;
  assign n1104 = pi137 & ~n1103;
  assign n1105 = ~pi89 & pi138;
  assign n1106 = pi62 & ~pi138;
  assign n1107 = pi136 & ~n1105;
  assign n1108 = ~n1106 & n1107;
  assign n1109 = ~pi119 & pi138;
  assign n1110 = pi72 & ~pi138;
  assign n1111 = ~pi136 & ~n1109;
  assign n1112 = ~n1110 & n1111;
  assign n1113 = ~n1108 & ~n1112;
  assign n1114 = ~pi137 & ~n1113;
  assign po98 = n1104 | n1114;
  assign n1116 = ~pi84 & ~n1076;
  assign n1117 = ~pi141 & n1076;
  assign n1118 = ~pi129 & ~n1116;
  assign po99 = ~n1117 & n1118;
  assign n1120 = ~pi85 & ~n626;
  assign n1121 = n644 & n652;
  assign n1122 = n620 & n1121;
  assign po100 = ~n1120 & n1122;
  assign n1124 = ~pi86 & ~n1076;
  assign n1125 = ~pi139 & n1076;
  assign n1126 = ~pi129 & ~n1124;
  assign po101 = ~n1125 & n1126;
  assign n1128 = ~pi87 & ~n1076;
  assign n1129 = ~pi140 & n1076;
  assign n1130 = ~pi129 & ~n1128;
  assign po102 = ~n1129 & n1130;
  assign n1132 = pi137 & n1097;
  assign n1133 = n1006 & n1132;
  assign n1134 = ~pi88 & ~n1133;
  assign n1135 = ~pi139 & n1133;
  assign n1136 = ~pi129 & ~n1134;
  assign po103 = ~n1135 & n1136;
  assign n1138 = ~pi89 & ~n1133;
  assign n1139 = ~pi140 & n1133;
  assign n1140 = ~pi129 & ~n1138;
  assign po104 = ~n1139 & n1140;
  assign n1142 = ~pi90 & ~n1133;
  assign n1143 = ~pi142 & n1133;
  assign n1144 = ~pi129 & ~n1142;
  assign po105 = ~n1143 & n1144;
  assign n1146 = ~pi91 & ~n1133;
  assign n1147 = ~pi143 & n1133;
  assign n1148 = ~pi129 & ~n1146;
  assign po106 = ~n1147 & n1148;
  assign n1150 = ~pi92 & ~n1133;
  assign n1151 = ~pi144 & n1133;
  assign n1152 = ~pi129 & ~n1150;
  assign po107 = ~n1151 & n1152;
  assign n1154 = ~pi93 & ~n1133;
  assign n1155 = ~pi146 & n1133;
  assign n1156 = ~pi129 & ~n1154;
  assign po108 = ~n1155 & n1156;
  assign n1158 = pi82 & pi138;
  assign n1159 = n1025 & n1158;
  assign n1160 = n1006 & n1159;
  assign n1161 = ~pi94 & ~n1160;
  assign n1162 = ~pi142 & n1160;
  assign n1163 = ~pi129 & ~n1161;
  assign po109 = ~n1162 & n1163;
  assign n1165 = ~pi3 & ~pi110;
  assign n1166 = ~n1006 & ~n1165;
  assign n1167 = ~n1160 & ~n1166;
  assign n1168 = pi95 & n1167;
  assign n1169 = pi143 & n1160;
  assign n1170 = ~n1168 & ~n1169;
  assign po110 = ~pi129 & ~n1170;
  assign n1172 = pi96 & n1167;
  assign n1173 = pi146 & n1160;
  assign n1174 = ~n1172 & ~n1173;
  assign po111 = ~pi129 & ~n1174;
  assign n1176 = pi97 & n1167;
  assign n1177 = pi145 & n1160;
  assign n1178 = ~n1176 & ~n1177;
  assign po112 = ~pi129 & ~n1178;
  assign n1180 = ~pi98 & ~n1133;
  assign n1181 = ~pi145 & n1133;
  assign n1182 = ~pi129 & ~n1180;
  assign po113 = ~n1181 & n1182;
  assign n1184 = ~pi99 & ~n1133;
  assign n1185 = ~pi141 & n1133;
  assign n1186 = ~pi129 & ~n1184;
  assign po114 = ~n1185 & n1186;
  assign n1188 = pi100 & n1167;
  assign n1189 = pi144 & n1160;
  assign n1190 = ~n1188 & ~n1189;
  assign po115 = ~pi129 & ~n1190;
  assign n1192 = pi37 & n1097;
  assign n1193 = ~pi82 & ~pi138;
  assign n1194 = ~pi96 & pi138;
  assign n1195 = ~pi136 & ~n1193;
  assign n1196 = ~n1194 & n1195;
  assign n1197 = ~n1192 & ~n1196;
  assign n1198 = pi137 & ~n1197;
  assign n1199 = ~pi93 & pi138;
  assign n1200 = pi65 & ~pi138;
  assign n1201 = pi136 & ~n1199;
  assign n1202 = ~n1200 & n1201;
  assign n1203 = ~pi124 & pi138;
  assign n1204 = pi77 & ~pi138;
  assign n1205 = ~pi136 & ~n1203;
  assign n1206 = ~n1204 & n1205;
  assign n1207 = ~n1202 & ~n1206;
  assign n1208 = ~pi137 & ~n1207;
  assign po116 = n1198 | n1208;
  assign n1210 = pi91 & n1004;
  assign n1211 = pi95 & n1075;
  assign n1212 = ~n1210 & ~n1211;
  assign n1213 = pi138 & ~n1212;
  assign n1214 = ~pi79 & ~pi136;
  assign n1215 = ~pi34 & pi136;
  assign n1216 = pi137 & ~n1214;
  assign n1217 = ~n1215 & n1216;
  assign n1218 = pi66 & ~pi136;
  assign n1219 = pi69 & pi136;
  assign n1220 = ~pi137 & ~n1218;
  assign n1221 = ~n1219 & n1220;
  assign n1222 = ~n1217 & ~n1221;
  assign n1223 = ~pi138 & ~n1222;
  assign po117 = n1213 | n1223;
  assign n1225 = pi90 & n1004;
  assign n1226 = pi94 & n1075;
  assign n1227 = ~n1225 & ~n1226;
  assign n1228 = pi138 & ~n1227;
  assign n1229 = ~pi78 & ~pi136;
  assign n1230 = ~pi33 & pi136;
  assign n1231 = pi137 & ~n1229;
  assign n1232 = ~n1230 & n1231;
  assign n1233 = pi74 & ~pi136;
  assign n1234 = pi63 & pi136;
  assign n1235 = ~pi137 & ~n1233;
  assign n1236 = ~n1234 & n1235;
  assign n1237 = ~n1232 & ~n1236;
  assign n1238 = ~pi138 & ~n1237;
  assign po118 = n1228 | n1238;
  assign n1240 = pi99 & n1004;
  assign n1241 = ~pi112 & n1075;
  assign n1242 = ~n1240 & ~n1241;
  assign n1243 = pi138 & ~n1242;
  assign n1244 = ~pi84 & ~pi136;
  assign n1245 = ~pi32 & pi136;
  assign n1246 = pi137 & ~n1244;
  assign n1247 = ~n1245 & n1246;
  assign n1248 = pi73 & ~pi136;
  assign n1249 = pi68 & pi136;
  assign n1250 = ~pi137 & ~n1248;
  assign n1251 = ~n1249 & n1250;
  assign n1252 = ~n1247 & ~n1251;
  assign n1253 = ~pi138 & ~n1252;
  assign po119 = n1243 | n1253;
  assign n1255 = pi35 & n1097;
  assign n1256 = ~pi80 & ~pi138;
  assign n1257 = ~pi100 & pi138;
  assign n1258 = ~pi136 & ~n1256;
  assign n1259 = ~n1257 & n1258;
  assign n1260 = ~n1255 & ~n1259;
  assign n1261 = pi137 & ~n1260;
  assign n1262 = ~pi92 & pi138;
  assign n1263 = pi70 & ~pi138;
  assign n1264 = pi136 & ~n1262;
  assign n1265 = ~n1263 & n1264;
  assign n1266 = ~pi125 & pi138;
  assign n1267 = pi75 & ~pi138;
  assign n1268 = ~pi136 & ~n1266;
  assign n1269 = ~n1267 & n1268;
  assign n1270 = ~n1265 & ~n1269;
  assign n1271 = ~pi137 & ~n1270;
  assign po120 = n1261 | n1271;
  assign n1273 = n612 & n718;
  assign n1274 = n626 & n1273;
  assign n1275 = ~n617 & ~n1274;
  assign po121 = n333 & ~n1275;
  assign n1277 = pi36 & n1097;
  assign n1278 = ~pi81 & ~pi138;
  assign n1279 = ~pi97 & pi138;
  assign n1280 = ~pi136 & ~n1278;
  assign n1281 = ~n1279 & n1280;
  assign n1282 = ~n1277 & ~n1281;
  assign n1283 = pi137 & ~n1282;
  assign n1284 = ~pi98 & pi138;
  assign n1285 = pi71 & ~pi138;
  assign n1286 = pi136 & ~n1284;
  assign n1287 = ~n1285 & n1286;
  assign n1288 = ~pi23 & pi138;
  assign n1289 = pi76 & ~pi138;
  assign n1290 = ~pi136 & ~n1288;
  assign n1291 = ~n1289 & n1290;
  assign n1292 = ~n1287 & ~n1291;
  assign n1293 = ~pi137 & ~n1292;
  assign po122 = n1283 | n1293;
  assign n1295 = pi30 & n1097;
  assign n1296 = ~pi86 & ~pi138;
  assign n1297 = ~pi111 & pi138;
  assign n1298 = ~pi136 & ~n1296;
  assign n1299 = ~n1297 & n1298;
  assign n1300 = ~n1295 & ~n1299;
  assign n1301 = pi137 & ~n1300;
  assign n1302 = ~pi88 & pi138;
  assign n1303 = pi64 & ~pi138;
  assign n1304 = pi136 & ~n1302;
  assign n1305 = ~n1303 & n1304;
  assign n1306 = ~pi120 & pi138;
  assign n1307 = pi67 & ~pi138;
  assign n1308 = ~pi136 & ~n1306;
  assign n1309 = ~n1307 & n1308;
  assign n1310 = ~n1305 & ~n1309;
  assign n1311 = ~pi137 & ~n1310;
  assign po123 = n1301 | n1311;
  assign n1313 = pi116 & n333;
  assign n1314 = pi27 & n607;
  assign n1315 = ~n974 & n1313;
  assign po124 = ~n1314 & n1315;
  assign n1317 = ~pi97 & n637;
  assign n1318 = ~n638 & ~n1317;
  assign po125 = n1313 & ~n1318;
  assign n1320 = ~pi129 & n1006;
  assign n1321 = ~pi111 & ~n1159;
  assign n1322 = ~pi139 & n1159;
  assign n1323 = n1320 & ~n1321;
  assign po126 = ~n1322 & n1323;
  assign n1325 = ~pi141 & n1159;
  assign n1326 = pi112 & ~n1159;
  assign n1327 = n1320 & ~n1325;
  assign po127 = ~n1326 & n1327;
  assign n1329 = ~pi54 & pi113;
  assign n1330 = ~pi11 & ~pi22;
  assign n1331 = pi54 & n1330;
  assign n1332 = n333 & ~n1329;
  assign po128 = ~n1331 & n1332;
  assign n1334 = ~pi140 & n1159;
  assign n1335 = pi115 & ~n1159;
  assign n1336 = n1320 & ~n1334;
  assign po130 = ~n1335 & n1336;
  assign n1338 = ~pi4 & ~pi7;
  assign n1339 = n492 & n1338;
  assign n1340 = pi54 & n333;
  assign po131 = ~n1339 & n1340;
  assign po132 = ~pi122 | pi129;
  assign n1343 = ~pi54 & pi118;
  assign n1344 = ~n503 & ~n1343;
  assign po133 = ~pi129 & ~n1344;
  assign po134 = ~pi129 & ~n624;
  assign n1347 = ~pi120 & n1165;
  assign n1348 = ~pi111 & ~pi129;
  assign po135 = ~n1347 & n1348;
  assign n1350 = pi81 & pi120;
  assign po136 = ~pi129 & n1350;
  assign po137 = pi129 | pi134;
  assign po138 = pi129 | pi135;
  assign po139 = pi57 & ~pi129;
  assign n1355 = ~pi96 & pi125;
  assign n1356 = ~pi3 & ~n1355;
  assign po140 = ~pi129 & ~n1356;
  assign n1358 = ~pi126 & pi132;
  assign po141 = pi133 & n1358;
  assign po12 = 1'b1;
  assign po0 = pi108;
  assign po1 = pi83;
  assign po2 = pi104;
  assign po3 = pi103;
  assign po4 = pi102;
  assign po5 = pi105;
  assign po6 = pi107;
  assign po7 = pi101;
  assign po8 = pi126;
  assign po9 = pi121;
  assign po10 = pi1;
  assign po11 = pi0;
  assign po13 = pi130;
  assign po14 = pi128;
endmodule
