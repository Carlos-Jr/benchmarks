module i2c ( 
    pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8, pi9,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19,
    pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29,
    pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38, pi39,
    pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48, pi49,
    pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59,
    pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69,
    pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79,
    pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88, pi89,
    pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97, pi98, pi99,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146,
    po0, po1, po2, po3, po4, po5, po6, po7, po8, po9,
    po10, po11, po12, po13, po14, po15, po16, po17, po18, po19,
    po20, po21, po22, po23, po24, po25, po26, po27, po28, po29,
    po30, po31, po32, po33, po34, po35, po36, po37, po38, po39,
    po40, po41, po42, po43, po44, po45, po46, po47, po48, po49,
    po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66, po67, po68, po69,
    po70, po71, po72, po73, po74, po75, po76, po77, po78, po79,
    po80, po81, po82, po83, po84, po85, po86, po87, po88, po89,
    po90, po91, po92, po93, po94, po95, po96, po97, po98, po99,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141  );
  input  pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8,
    pi9, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18,
    pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28,
    pi29, pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38,
    pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48,
    pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58,
    pi59, pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68,
    pi69, pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78,
    pi79, pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88,
    pi89, pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97, pi98,
    pi99, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146;
  output po0, po1, po2, po3, po4, po5, po6, po7, po8, po9,
    po10, po11, po12, po13, po14, po15, po16, po17, po18, po19,
    po20, po21, po22, po23, po24, po25, po26, po27, po28, po29,
    po30, po31, po32, po33, po34, po35, po36, po37, po38, po39,
    po40, po41, po42, po43, po44, po45, po46, po47, po48, po49,
    po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66, po67, po68, po69,
    po70, po71, po72, po73, po74, po75, po76, po77, po78, po79,
    po80, po81, po82, po83, po84, po85, po86, po87, po88, po89,
    po90, po91, po92, po93, po94, po95, po96, po97, po98, po99,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141;
  wire n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339,
    n340, n341, n342, n343, n344, n345, n346,
    n347, n348, n349, n350, n351, n352, n353,
    n354, n355, n356, n357, n358, n359, n360,
    n361, n362, n363, n364, n365, n366, n367,
    n368, n369, n370, n371, n372, n373, n374,
    n375, n376, n377, n378, n379, n380, n381,
    n382, n383, n384, n385, n386, n387, n388,
    n389, n390, n391, n392, n393, n394, n395,
    n396, n397, n398, n399, n400, n401, n402,
    n403, n404, n405, n406, n407, n408, n409,
    n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423,
    n424, n425, n426, n427, n428, n429, n430,
    n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444,
    n445, n446, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487,
    n488, n489, n490, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501,
    n502, n503, n504, n505, n506, n507, n508,
    n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n541, n542, n543,
    n544, n545, n546, n547, n548, n549, n550,
    n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564,
    n565, n566, n567, n568, n569, n570, n571,
    n572, n573, n574, n575, n576, n577, n578,
    n580, n581, n582, n583, n584, n585, n586,
    n587, n588, n589, n590, n591, n592, n593,
    n594, n595, n596, n597, n598, n599, n600,
    n601, n602, n603, n604, n605, n606, n607,
    n608, n609, n610, n611, n612, n613, n614,
    n615, n616, n617, n618, n619, n620, n621,
    n622, n623, n625, n626, n627, n628, n629,
    n630, n631, n632, n633, n634, n635, n636,
    n637, n638, n639, n640, n641, n642, n643,
    n644, n645, n646, n647, n648, n649, n650,
    n651, n652, n653, n654, n655, n656, n657,
    n658, n659, n660, n661, n662, n663, n664,
    n665, n666, n667, n668, n669, n670, n671,
    n672, n673, n674, n675, n676, n677, n678,
    n679, n680, n681, n682, n683, n684, n685,
    n686, n687, n688, n689, n690, n691, n692,
    n693, n694, n695, n696, n697, n698, n699,
    n700, n701, n702, n703, n704, n705, n706,
    n707, n708, n709, n710, n711, n712, n713,
    n714, n715, n716, n717, n718, n719, n720,
    n721, n722, n723, n724, n725, n726, n727,
    n728, n729, n730, n731, n732, n733, n734,
    n735, n736, n737, n738, n739, n740, n741,
    n742, n743, n744, n745, n746, n747, n748,
    n749, n750, n751, n752, n753, n754, n755,
    n756, n757, n758, n759, n760, n761, n762,
    n763, n764, n765, n766, n767, n768, n769,
    n770, n771, n772, n773, n774, n775, n776,
    n777, n778, n779, n780, n781, n782, n783,
    n784, n785, n786, n787, n788, n789, n790,
    n791, n792, n793, n794, n795, n796, n797,
    n798, n799, n800, n801, n802, n803, n804,
    n805, n806, n807, n808, n809, n810, n811,
    n812, n813, n814, n815, n816, n817, n818,
    n819, n820, n821, n822, n823, n824, n825,
    n826, n827, n828, n829, n830, n831, n832,
    n833, n834, n835, n836, n837, n838, n839,
    n840, n841, n842, n843, n844, n845, n846,
    n847, n848, n849, n850, n851, n852, n853,
    n854, n855, n856, n857, n858, n859, n860,
    n861, n862, n863, n864, n865, n866, n867,
    n868, n869, n870, n871, n872, n873, n874,
    n875, n876, n877, n878, n879, n880, n881,
    n882, n883, n884, n885, n886, n887, n888,
    n889, n890, n891, n892, n893, n894, n895,
    n896, n897, n898, n899, n900, n901, n902,
    n903, n904, n905, n906, n907, n908, n909,
    n910, n911, n912, n913, n914, n915, n916,
    n917, n918, n919, n920, n921, n922, n923,
    n924, n925, n926, n927, n928, n929, n930,
    n931, n932, n933, n934, n935, n936, n937,
    n938, n939, n940, n941, n942, n943, n944,
    n945, n946, n947, n948, n949, n950, n951,
    n952, n953, n954, n955, n956, n957, n959,
    n960, n961, n962, n963, n964, n965, n966,
    n967, n968, n969, n970, n971, n972, n973,
    n974, n975, n976, n977, n978, n979, n980,
    n981, n982, n983, n984, n985, n986, n987,
    n988, n989, n990, n991, n992, n993, n994,
    n995, n996, n997, n998, n999, n1000, n1001,
    n1002, n1003, n1004, n1005, n1006, n1007,
    n1008, n1009, n1010, n1011, n1012, n1013,
    n1014, n1015, n1016, n1017, n1018, n1019,
    n1020, n1021, n1022, n1023, n1024, n1025,
    n1026, n1027, n1028, n1029, n1030, n1031,
    n1032, n1033, n1034, n1035, n1036, n1037,
    n1038, n1039, n1040, n1041, n1042, n1043,
    n1044, n1045, n1046, n1047, n1048, n1049,
    n1050, n1051, n1052, n1053, n1054, n1055,
    n1056, n1057, n1058, n1059, n1060, n1061,
    n1062, n1063, n1064, n1065, n1066, n1067,
    n1068, n1069, n1070, n1071, n1072, n1073,
    n1074, n1075, n1076, n1077, n1078, n1079,
    n1080, n1081, n1082, n1083, n1084, n1085,
    n1086, n1087, n1088, n1089, n1090, n1091,
    n1092, n1093, n1094, n1095, n1096, n1097,
    n1098, n1099, n1100, n1101, n1102, n1103,
    n1104, n1105, n1106, n1107, n1108, n1109,
    n1110, n1111, n1112, n1113, n1114, n1115,
    n1116, n1117, n1118, n1119, n1120, n1121,
    n1122, n1123, n1124, n1125, n1126, n1127,
    n1128, n1129, n1130, n1131, n1132, n1133,
    n1134, n1135, n1136, n1137, n1138, n1139,
    n1140, n1141, n1142, n1143, n1144, n1145,
    n1146, n1147, n1148, n1149, n1150, n1151,
    n1152, n1153, n1154, n1155, n1156, n1157,
    n1158, n1159, n1160, n1161, n1162, n1163,
    n1164, n1165, n1166, n1167, n1168, n1169,
    n1170, n1171, n1172, n1173, n1174, n1175,
    n1176, n1177, n1178, n1179, n1180, n1181,
    n1182, n1183, n1184, n1185, n1186, n1187,
    n1188, n1189, n1190, n1191, n1192, n1193,
    n1194, n1195, n1196, n1197, n1198, n1199,
    n1200, n1201, n1202, n1203, n1204, n1205,
    n1206, n1207, n1208, n1209, n1210, n1211,
    n1212, n1213, n1214, n1215, n1216, n1217,
    n1218, n1219, n1220, n1221, n1222, n1223,
    n1224, n1225, n1226, n1227, n1228, n1229,
    n1230, n1231, n1232, n1233, n1234, n1235,
    n1236, n1237, n1238, n1239, n1240, n1241,
    n1242, n1243, n1244, n1245, n1246, n1247,
    n1248, n1249, n1250, n1251, n1252, n1253,
    n1254, n1255, n1256, n1257, n1258, n1259,
    n1260, n1261, n1262, n1263, n1264, n1265,
    n1266, n1267, n1268, n1269, n1270, n1271,
    n1272, n1273, n1274, n1275, n1276, n1277,
    n1278, n1279, n1280, n1281, n1282, n1283,
    n1284, n1285, n1286, n1287, n1288, n1289,
    n1290, n1291, n1292, n1293, n1294, n1295,
    n1296, n1297, n1299, n1300, n1301, n1302,
    n1303, n1304, n1305, n1306, n1307, n1308,
    n1309, n1310, n1311, n1312, n1313, n1314,
    n1315, n1316, n1317, n1318, n1319, n1320,
    n1322, n1323, n1324, n1325, n1326, n1327,
    n1328, n1329, n1330, n1331, n1332, n1333,
    n1334, n1335, n1336, n1337, n1338, n1339,
    n1340, n1341, n1342, n1343, n1344, n1345,
    n1346, n1347, n1348, n1349, n1350, n1351,
    n1352, n1353, n1354, n1355, n1356, n1357,
    n1358, n1359, n1360, n1361, n1362, n1363,
    n1364, n1365, n1366, n1367, n1368, n1369,
    n1370, n1371, n1372, n1373, n1374, n1375,
    n1376, n1377, n1378, n1379, n1380, n1381,
    n1382, n1383, n1384, n1385, n1386, n1387,
    n1388, n1389, n1390, n1391, n1392, n1393,
    n1395, n1396, n1397, n1398, n1399, n1400,
    n1401, n1402, n1403, n1404, n1405, n1406,
    n1408, n1409, n1410, n1411, n1412, n1413,
    n1414, n1415, n1416, n1417, n1418, n1419,
    n1420, n1421, n1422, n1423, n1424, n1425,
    n1426, n1427, n1428, n1429, n1430, n1431,
    n1432, n1433, n1434, n1435, n1436, n1437,
    n1438, n1439, n1440, n1441, n1442, n1443,
    n1444, n1445, n1446, n1447, n1448, n1450,
    n1451, n1452, n1453, n1454, n1455, n1456,
    n1457, n1458, n1459, n1460, n1461, n1462,
    n1463, n1464, n1465, n1466, n1467, n1468,
    n1469, n1470, n1471, n1472, n1473, n1474,
    n1475, n1476, n1477, n1478, n1479, n1480,
    n1481, n1482, n1483, n1484, n1485, n1486,
    n1487, n1488, n1489, n1490, n1491, n1492,
    n1493, n1494, n1495, n1496, n1497, n1498,
    n1499, n1500, n1501, n1502, n1503, n1504,
    n1505, n1506, n1507, n1508, n1509, n1510,
    n1511, n1512, n1513, n1514, n1515, n1516,
    n1517, n1518, n1519, n1520, n1521, n1522,
    n1523, n1525, n1526, n1527, n1528, n1529,
    n1530, n1531, n1532, n1533, n1534, n1535,
    n1536, n1537, n1538, n1539, n1540, n1541,
    n1542, n1543, n1544, n1545, n1546, n1547,
    n1548, n1549, n1550, n1551, n1552, n1553,
    n1554, n1555, n1556, n1557, n1558, n1559,
    n1560, n1561, n1562, n1563, n1564, n1565,
    n1566, n1567, n1568, n1569, n1570, n1571,
    n1572, n1573, n1574, n1575, n1576, n1577,
    n1578, n1579, n1580, n1581, n1582, n1583,
    n1584, n1585, n1586, n1587, n1588, n1589,
    n1590, n1591, n1592, n1593, n1594, n1595,
    n1596, n1597, n1598, n1599, n1600, n1601,
    n1602, n1603, n1604, n1605, n1606, n1607,
    n1608, n1609, n1610, n1611, n1612, n1613,
    n1614, n1615, n1616, n1617, n1618, n1619,
    n1620, n1621, n1622, n1623, n1624, n1625,
    n1626, n1627, n1628, n1629, n1630, n1631,
    n1632, n1633, n1634, n1635, n1637, n1638,
    n1639, n1641, n1642, n1643, n1645, n1646,
    n1647, n1649, n1650, n1651, n1652, n1653,
    n1654, n1655, n1656, n1657, n1658, n1659,
    n1660, n1661, n1662, n1663, n1664, n1665,
    n1666, n1667, n1668, n1669, n1670, n1671,
    n1672, n1673, n1674, n1675, n1676, n1677,
    n1678, n1679, n1680, n1681, n1682, n1683,
    n1684, n1685, n1686, n1687, n1688, n1689,
    n1690, n1691, n1692, n1693, n1694, n1695,
    n1696, n1697, n1698, n1699, n1700, n1701,
    n1702, n1703, n1704, n1705, n1706, n1707,
    n1708, n1709, n1710, n1711, n1712, n1713,
    n1714, n1715, n1716, n1717, n1718, n1719,
    n1720, n1721, n1722, n1723, n1724, n1725,
    n1726, n1727, n1728, n1729, n1730, n1731,
    n1732, n1733, n1734, n1735, n1736, n1737,
    n1738, n1739, n1740, n1741, n1742, n1743,
    n1744, n1745, n1746, n1747, n1748, n1749,
    n1750, n1751, n1752, n1753, n1754, n1755,
    n1756, n1757, n1758, n1759, n1760, n1761,
    n1762, n1763, n1764, n1765, n1766, n1767,
    n1768, n1769, n1770, n1771, n1772, n1773,
    n1774, n1775, n1776, n1777, n1778, n1779,
    n1780, n1781, n1782, n1783, n1784, n1785,
    n1786, n1787, n1788, n1789, n1790, n1791,
    n1792, n1793, n1794, n1795, n1796, n1797,
    n1798, n1799, n1800, n1801, n1802, n1803,
    n1804, n1805, n1806, n1807, n1809, n1810,
    n1811, n1813, n1814, n1815, n1816, n1817,
    n1818, n1819, n1820, n1821, n1822, n1824,
    n1825, n1827, n1828, n1829, n1830, n1831,
    n1832, n1833, n1834, n1835, n1836, n1837,
    n1838, n1839, n1840, n1841, n1842, n1843,
    n1844, n1845, n1846, n1847, n1848, n1849,
    n1850, n1851, n1852, n1853, n1854, n1855,
    n1856, n1857, n1858, n1859, n1860, n1861,
    n1862, n1863, n1864, n1865, n1866, n1867,
    n1868, n1869, n1870, n1871, n1872, n1873,
    n1874, n1875, n1876, n1877, n1878, n1879,
    n1880, n1881, n1882, n1883, n1884, n1885,
    n1886, n1887, n1888, n1889, n1890, n1891,
    n1892, n1893, n1894, n1895, n1896, n1897,
    n1898, n1899, n1900, n1901, n1902, n1903,
    n1904, n1905, n1906, n1907, n1908, n1909,
    n1910, n1911, n1912, n1913, n1914, n1915,
    n1916, n1917, n1918, n1919, n1920, n1921,
    n1922, n1923, n1924, n1925, n1926, n1927,
    n1928, n1929, n1930, n1931, n1932, n1933,
    n1934, n1935, n1936, n1937, n1938, n1939,
    n1940, n1941, n1942, n1943, n1944, n1945,
    n1946, n1947, n1948, n1949, n1950, n1951,
    n1952, n1953, n1954, n1955, n1956, n1957,
    n1958, n1959, n1960, n1961, n1962, n1963,
    n1964, n1965, n1966, n1967, n1968, n1969,
    n1970, n1971, n1972, n1973, n1974, n1975,
    n1976, n1977, n1978, n1979, n1980, n1981,
    n1982, n1983, n1984, n1985, n1986, n1987,
    n1988, n1989, n1990, n1991, n1992, n1993,
    n1994, n1995, n1996, n1997, n1998, n1999,
    n2000, n2001, n2002, n2003, n2004, n2005,
    n2006, n2007, n2008, n2009, n2010, n2011,
    n2012, n2013, n2014, n2015, n2016, n2017,
    n2018, n2019, n2020, n2021, n2022, n2023,
    n2024, n2025, n2026, n2027, n2028, n2029,
    n2030, n2031, n2032, n2033, n2034, n2035,
    n2036, n2037, n2038, n2039, n2040, n2041,
    n2042, n2043, n2044, n2045, n2046, n2047,
    n2048, n2049, n2050, n2051, n2052, n2053,
    n2054, n2055, n2056, n2057, n2058, n2059,
    n2060, n2061, n2062, n2063, n2064, n2065,
    n2066, n2067, n2068, n2069, n2070, n2071,
    n2072, n2073, n2074, n2075, n2076, n2077,
    n2078, n2079, n2080, n2081, n2082, n2083,
    n2084, n2085, n2086, n2087, n2088, n2089,
    n2090, n2091, n2092, n2093, n2094, n2095,
    n2096, n2097, n2098, n2099, n2100, n2101,
    n2102, n2103, n2104, n2105, n2106, n2107,
    n2108, n2109, n2110, n2111, n2112, n2113,
    n2114, n2115, n2116, n2117, n2118, n2119,
    n2120, n2121, n2122, n2123, n2124, n2125,
    n2126, n2127, n2128, n2129, n2130, n2131,
    n2132, n2133, n2134, n2135, n2136, n2137,
    n2138, n2139, n2140, n2141, n2142, n2143,
    n2144, n2145, n2146, n2147, n2148, n2149,
    n2150, n2151, n2152, n2153, n2154, n2155,
    n2156, n2157, n2158, n2159, n2160, n2161,
    n2162, n2163, n2164, n2165, n2166, n2167,
    n2168, n2169, n2170, n2171, n2172, n2173,
    n2174, n2175, n2176, n2177, n2178, n2179,
    n2180, n2181, n2182, n2183, n2184, n2185,
    n2186, n2187, n2188, n2189, n2190, n2191,
    n2192, n2193, n2194, n2195, n2196, n2197,
    n2198, n2199, n2200, n2201, n2202, n2203,
    n2204, n2205, n2206, n2207, n2208, n2209,
    n2210, n2211, n2212, n2213, n2214, n2215,
    n2216, n2217, n2218, n2219, n2220, n2221,
    n2222, n2223, n2224, n2225, n2226, n2227,
    n2228, n2229, n2230, n2231, n2232, n2233,
    n2234, n2235, n2236, n2237, n2238, n2239,
    n2240, n2241, n2242, n2243, n2244, n2245,
    n2246, n2247, n2248, n2249, n2250, n2251,
    n2252, n2253, n2254, n2255, n2256, n2257,
    n2258, n2259, n2260, n2261, n2262, n2263,
    n2264, n2265, n2266, n2267, n2268, n2269,
    n2270, n2271, n2272, n2273, n2274, n2275,
    n2276, n2277, n2278, n2279, n2280, n2281,
    n2282, n2283, n2284, n2285, n2286, n2287,
    n2288, n2289, n2290, n2291, n2292, n2293,
    n2294, n2295, n2296, n2297, n2298, n2299,
    n2300, n2301, n2302, n2303, n2304, n2305,
    n2306, n2307, n2308, n2309, n2310, n2311,
    n2312, n2313, n2314, n2315, n2316, n2317,
    n2318, n2319, n2320, n2321, n2322, n2323,
    n2324, n2325, n2326, n2327, n2328, n2329,
    n2330, n2331, n2332, n2333, n2334, n2335,
    n2336, n2337, n2338, n2339, n2340, n2341,
    n2342, n2343, n2344, n2345, n2346, n2347,
    n2348, n2349, n2350, n2351, n2352, n2353,
    n2354, n2355, n2356, n2357, n2358, n2359,
    n2360, n2361, n2362, n2363, n2364, n2365,
    n2366, n2367, n2368, n2369, n2370, n2371,
    n2372, n2373, n2374, n2375, n2376, n2377,
    n2378, n2379, n2380, n2381, n2382, n2383,
    n2384, n2385, n2386, n2387, n2388, n2389,
    n2390, n2391, n2392, n2393, n2394, n2395,
    n2396, n2397, n2398, n2399, n2400, n2401,
    n2402, n2403, n2404, n2405, n2406, n2407,
    n2408, n2409, n2410, n2411, n2412, n2413,
    n2414, n2415, n2416, n2417, n2418, n2419,
    n2420, n2421, n2422, n2423, n2424, n2425,
    n2426, n2427, n2428, n2429, n2430, n2431,
    n2432, n2433, n2434, n2435, n2436, n2437,
    n2438, n2440, n2441, n2442, n2443, n2444,
    n2445, n2446, n2447, n2448, n2449, n2450,
    n2451, n2452, n2453, n2454, n2455, n2456,
    n2457, n2458, n2459, n2460, n2461, n2462,
    n2463, n2464, n2465, n2466, n2469, n2471,
    n2474, n2475, n2476, n2477, n2478, n2479,
    n2480, n2481, n2482, n2483, n2484, n2485,
    n2486, n2487, n2488, n2489, n2490, n2491,
    n2492, n2493, n2494, n2495, n2496, n2497,
    n2498, n2499, n2500, n2501, n2502, n2503,
    n2504, n2505, n2506, n2507, n2508, n2509,
    n2510, n2512, n2513, n2515, n2516, n2517,
    n2518, n2519, n2520, n2522, n2523, n2524,
    n2525, n2527, n2528, n2529, n2530, n2531,
    n2532, n2533, n2534, n2535, n2536, n2537,
    n2538, n2539, n2540, n2541, n2542, n2543,
    n2544, n2545, n2547, n2548, n2550, n2551,
    n2553, n2555, n2556, n2558, n2559, n2561,
    n2563, n2565, n2566, n2568, n2569, n2571,
    n2573, n2574, n2575, n2577, n2578, n2580,
    n2581, n2582, n2584, n2585, n2586, n2587,
    n2588, n2590, n2591, n2592, n2593, n2594,
    n2595, n2597, n2598, n2600, n2602, n2603,
    n2604, n2605, n2606, n2607, n2608, n2609,
    n2611, n2612, n2613, n2614, n2615, n2616,
    n2617, n2618, n2619, n2620, n2621, n2622,
    n2623, n2624, n2625, n2627, n2628, n2629,
    n2631, n2632, n2633, n2634, n2635, n2636,
    n2637, n2638, n2639, n2640, n2642, n2643,
    n2644, n2645, n2647, n2648, n2649, n2651,
    n2652, n2653, n2654, n2655, n2656, n2657,
    n2659, n2660, n2661, n2663, n2664, n2666,
    n2668, n2669, n2670, n2671, n2672, n2673,
    n2674, n2675, n2677, n2678, n2680, n2681,
    n2683, n2684, n2686, n2687, n2689, n2690,
    n2692, n2693, n2695, n2696, n2699, n2701,
    n2703, n2705, n2707, n2709, n2710, n2711,
    n2713, n2714, n2715, n2716, n2717, n2718,
    n2719, n2720, n2721, n2722, n2723, n2724,
    n2728, n2729, n2730, n2731, n2732, n2733,
    n2734, n2735, n2736, n2737, n2738, n2739,
    n2740, n2741, n2742, n2743, n2744, n2753,
    n2762, n2763, n2764, n2765, n2767, n2771;
  assign po12 = 1'b1;
  assign n291 = pi122 & pi127;
  assign n292 = ~pi82 & ~n291;
  assign n293 = ~pi42 & ~pi44;
  assign n294 = ~pi38 & ~pi40;
  assign n295 = ~pi46 & ~pi50;
  assign n296 = ~pi38 & ~pi46;
  assign n297 = ~pi38 & ~pi50;
  assign n298 = ~pi46 & n297;
  assign n299 = ~pi50 & n296;
  assign n300 = ~pi40 & n2474;
  assign n301 = n294 & n295;
  assign n302 = ~pi40 & n293;
  assign n303 = n2474 & n302;
  assign n304 = n295 & n302;
  assign n305 = ~pi38 & n304;
  assign n306 = n293 & n2475;
  assign n307 = ~pi45 & ~pi48;
  assign n308 = ~pi41 & ~pi43;
  assign n309 = ~pi47 & n308;
  assign n310 = n307 & n309;
  assign n311 = n293 & n294;
  assign n312 = ~pi41 & ~pi46;
  assign n313 = ~pi41 & n295;
  assign n314 = ~pi50 & n312;
  assign n315 = ~pi42 & ~pi50;
  assign n316 = ~pi40 & ~pi42;
  assign n317 = n297 & n316;
  assign n318 = ~pi38 & n316;
  assign n319 = ~pi42 & n294;
  assign n320 = ~pi50 & n2479;
  assign n321 = n294 & n315;
  assign n322 = ~pi50 & n311;
  assign n323 = n297 & n302;
  assign n324 = ~pi50 & n293;
  assign n325 = n294 & n324;
  assign n326 = ~pi44 & n2478;
  assign n327 = n312 & n2480;
  assign n328 = n311 & n2477;
  assign n329 = ~pi43 & n2481;
  assign n330 = n2476 & n308;
  assign n331 = ~pi47 & n2482;
  assign n332 = ~pi43 & ~pi47;
  assign n333 = n312 & n332;
  assign n334 = n2480 & n333;
  assign n335 = n2476 & n309;
  assign n336 = n307 & n2483;
  assign n337 = ~pi47 & ~pi48;
  assign n338 = ~pi45 & n337;
  assign n339 = ~pi43 & n312;
  assign n340 = n338 & n339;
  assign n341 = n307 & n333;
  assign n342 = n2480 & n2485;
  assign n343 = n2482 & n338;
  assign n344 = n2476 & n310;
  assign n345 = ~pi2 & ~pi20;
  assign n346 = ~pi15 & ~pi49;
  assign n347 = ~pi15 & ~pi20;
  assign n348 = ~pi2 & n347;
  assign n349 = ~pi49 & n348;
  assign n350 = n345 & n346;
  assign n351 = ~pi24 & ~pi49;
  assign n352 = n348 & n351;
  assign n353 = ~pi24 & n2486;
  assign n354 = ~n291 & n2487;
  assign n355 = n2484 & n354;
  assign n356 = ~pi15 & n351;
  assign n357 = ~pi20 & n356;
  assign n358 = n347 & n351;
  assign n359 = n307 & n332;
  assign n360 = n2488 & n359;
  assign n361 = ~pi41 & n2474;
  assign n362 = ~pi38 & n2477;
  assign n363 = n297 & n312;
  assign n364 = ~pi2 & n302;
  assign n365 = n2489 & n364;
  assign n366 = n360 & n365;
  assign n367 = ~pi2 & ~pi45;
  assign n368 = n337 & n367;
  assign n369 = ~pi49 & n347;
  assign n370 = ~pi24 & ~pi45;
  assign n371 = ~pi2 & ~pi48;
  assign n372 = n370 & n371;
  assign n373 = n307 & n2487;
  assign n374 = n369 & n372;
  assign n375 = ~pi47 & n2491;
  assign n376 = ~pi2 & n337;
  assign n377 = n2488 & n376;
  assign n378 = ~pi45 & n377;
  assign n379 = n2488 & n368;
  assign n380 = n2482 & n2492;
  assign n381 = n2484 & n2487;
  assign n382 = pi82 & ~n2490;
  assign n383 = ~n291 & ~n382;
  assign n384 = ~n292 & ~n355;
  assign n385 = ~pi65 & ~n291;
  assign n386 = ~n382 & n385;
  assign n387 = ~pi65 & n2493;
  assign n388 = pi82 & ~n2484;
  assign n389 = ~pi82 & n291;
  assign n390 = pi82 & ~n2488;
  assign n391 = ~n389 & ~n390;
  assign n392 = ~pi24 & n307;
  assign n393 = n333 & n392;
  assign n394 = ~pi50 & n294;
  assign n395 = n293 & n346;
  assign n396 = n394 & n395;
  assign n397 = n2484 & n356;
  assign n398 = n308 & n337;
  assign n399 = ~pi45 & n351;
  assign n400 = n398 & n399;
  assign n401 = ~pi15 & n2476;
  assign n402 = n400 & n401;
  assign n403 = n307 & n351;
  assign n404 = ~pi48 & n332;
  assign n405 = ~pi43 & n337;
  assign n406 = n399 & n2496;
  assign n407 = n332 & n403;
  assign n408 = n2480 & n351;
  assign n409 = n2485 & n408;
  assign n410 = n2484 & n351;
  assign n411 = n337 & n339;
  assign n412 = n312 & n2496;
  assign n413 = ~pi48 & n2478;
  assign n414 = n333 & n413;
  assign n415 = ~pi44 & n414;
  assign n416 = ~pi50 & n2499;
  assign n417 = n2477 & n2496;
  assign n418 = n311 & n2501;
  assign n419 = n2480 & n2499;
  assign n420 = ~pi44 & n394;
  assign n421 = ~pi24 & ~pi42;
  assign n422 = n420 & n421;
  assign n423 = n2485 & n422;
  assign n424 = ~pi24 & n2484;
  assign n425 = n370 & n2500;
  assign n426 = ~pi49 & n2502;
  assign n427 = n2481 & n2497;
  assign n428 = ~pi15 & n2498;
  assign n429 = ~pi15 & n403;
  assign n430 = n2483 & n429;
  assign n431 = n346 & n2502;
  assign n432 = n393 & n396;
  assign n433 = ~pi44 & n369;
  assign n434 = n2478 & n433;
  assign n435 = n393 & n434;
  assign n436 = n337 & n370;
  assign n437 = n369 & n436;
  assign n438 = n2482 & n437;
  assign n439 = n347 & n2498;
  assign n440 = n2484 & n2488;
  assign n441 = ~pi20 & n2495;
  assign n442 = pi82 & ~n2503;
  assign n443 = ~n389 & ~n442;
  assign n444 = ~n388 & n391;
  assign n445 = pi2 & ~n2504;
  assign n446 = ~n2494 & ~n445;
  assign po17 = ~pi129 & ~n446;
  assign n448 = ~pi3 & ~pi129;
  assign n449 = pi5 & ~pi54;
  assign n450 = ~pi10 & ~pi22;
  assign n451 = ~pi9 & ~pi14;
  assign n452 = n450 & n451;
  assign n453 = ~pi13 & n452;
  assign n454 = ~pi8 & ~pi11;
  assign n455 = ~pi17 & ~pi21;
  assign n456 = ~pi8 & ~pi21;
  assign n457 = ~pi11 & n456;
  assign n458 = ~pi17 & n457;
  assign n459 = ~pi8 & n455;
  assign n460 = ~pi17 & n456;
  assign n461 = ~pi11 & n2506;
  assign n462 = n454 & n455;
  assign n463 = ~pi59 & n2505;
  assign n464 = n453 & n463;
  assign n465 = ~pi5 & ~pi6;
  assign n466 = ~pi7 & ~pi12;
  assign n467 = ~pi6 & ~pi12;
  assign n468 = ~pi5 & ~pi7;
  assign n469 = n467 & n468;
  assign n470 = n465 & n466;
  assign n471 = ~pi16 & pi54;
  assign n472 = n2507 & n471;
  assign n473 = ~pi4 & ~pi19;
  assign n474 = ~pi4 & ~pi18;
  assign n475 = ~pi19 & n474;
  assign n476 = ~pi18 & n473;
  assign n477 = ~pi25 & pi28;
  assign n478 = ~pi25 & ~pi29;
  assign n479 = pi28 & n478;
  assign n480 = ~pi29 & n477;
  assign n481 = n2508 & n2509;
  assign n482 = n472 & n481;
  assign n483 = ~pi7 & n467;
  assign n484 = n2509 & n483;
  assign n485 = n453 & n484;
  assign n486 = ~pi5 & n2508;
  assign n487 = n471 & n486;
  assign n488 = n463 & n487;
  assign n489 = n485 & n488;
  assign n490 = n464 & n482;
  assign n491 = ~n449 & ~n2510;
  assign n492 = ~pi129 & ~n491;
  assign n493 = ~pi3 & n492;
  assign n494 = n448 & ~n491;
  assign n495 = pi6 & ~pi54;
  assign n496 = pi25 & ~pi28;
  assign n497 = pi25 & ~pi29;
  assign n498 = ~pi28 & n497;
  assign n499 = ~pi28 & ~pi29;
  assign n500 = pi25 & n499;
  assign n501 = ~pi29 & n496;
  assign n502 = n2508 & n2512;
  assign n503 = n472 & n502;
  assign n504 = ~pi12 & n2512;
  assign n505 = n468 & n504;
  assign n506 = n453 & n505;
  assign n507 = ~pi6 & n2508;
  assign n508 = n471 & n507;
  assign n509 = n463 & n508;
  assign n510 = n506 & n509;
  assign n511 = n464 & n503;
  assign n512 = ~n495 & ~n2513;
  assign n513 = ~pi129 & ~n512;
  assign n514 = ~pi3 & n513;
  assign n515 = n448 & ~n512;
  assign n516 = pi13 & ~pi54;
  assign n517 = ~pi13 & n2508;
  assign n518 = n471 & n517;
  assign n519 = n463 & n518;
  assign n520 = ~pi5 & n467;
  assign n521 = ~pi25 & ~pi28;
  assign n522 = ~pi25 & pi29;
  assign n523 = ~pi28 & n522;
  assign n524 = pi29 & n521;
  assign n525 = n520 & n2515;
  assign n526 = ~pi7 & n452;
  assign n527 = n525 & n526;
  assign n528 = ~pi7 & ~pi13;
  assign n529 = n465 & n528;
  assign n530 = ~pi12 & n452;
  assign n531 = n520 & n528;
  assign n532 = ~pi13 & n2507;
  assign n533 = ~pi12 & n529;
  assign n534 = n452 & n2516;
  assign n535 = n452 & n529;
  assign n536 = ~pi12 & n535;
  assign n537 = n529 & n530;
  assign n538 = n2508 & n2517;
  assign n539 = n471 & n538;
  assign n540 = n463 & n2515;
  assign n541 = n539 & n540;
  assign n542 = n471 & n473;
  assign n543 = n471 & n2508;
  assign n544 = ~pi4 & ~pi16;
  assign n545 = ~pi18 & ~pi19;
  assign n546 = ~pi16 & n2508;
  assign n547 = n544 & n545;
  assign n548 = pi54 & n2520;
  assign n549 = ~pi18 & n542;
  assign n550 = n452 & n2515;
  assign n551 = n2516 & n550;
  assign n552 = n2519 & n551;
  assign n553 = n463 & n552;
  assign n554 = n519 & n527;
  assign n555 = ~n516 & ~n2518;
  assign n556 = ~pi129 & ~n555;
  assign n557 = ~pi3 & n556;
  assign n558 = n448 & ~n555;
  assign n559 = ~pi15 & ~n345;
  assign n560 = n2482 & n559;
  assign n561 = n351 & n560;
  assign n562 = n338 & n561;
  assign n563 = ~n345 & n356;
  assign n564 = n2484 & n563;
  assign n565 = ~n345 & n2495;
  assign n566 = pi15 & ~n2498;
  assign n567 = ~n2522 & ~n566;
  assign n568 = pi82 & ~n567;
  assign n569 = pi15 & n389;
  assign n570 = pi82 & ~n2495;
  assign n571 = ~pi70 & ~n291;
  assign n572 = ~n291 & ~n570;
  assign n573 = ~pi70 & n572;
  assign n574 = ~n570 & n571;
  assign n575 = ~n569 & ~n2523;
  assign n576 = ~n568 & ~n569;
  assign n577 = ~n2523 & n576;
  assign n578 = ~n568 & n575;
  assign po30 = ~pi129 & ~n2524;
  assign n580 = pi17 & ~pi54;
  assign n581 = ~pi29 & pi59;
  assign n582 = n521 & n581;
  assign n583 = n2507 & n582;
  assign n584 = n2520 & n583;
  assign n585 = ~pi17 & pi54;
  assign n586 = n457 & n585;
  assign n587 = n453 & n586;
  assign n588 = ~pi7 & n465;
  assign n589 = ~pi12 & n521;
  assign n590 = n588 & n589;
  assign n591 = n453 & n590;
  assign n592 = ~pi16 & n585;
  assign n593 = n2508 & n592;
  assign n594 = n457 & n581;
  assign n595 = n593 & n594;
  assign n596 = n591 & n595;
  assign n597 = n2507 & n499;
  assign n598 = ~pi25 & pi59;
  assign n599 = n585 & n598;
  assign n600 = n457 & n599;
  assign n601 = n597 & n600;
  assign n602 = n453 & n2520;
  assign n603 = n601 & n602;
  assign n604 = n584 & n587;
  assign n605 = ~n580 & ~n2525;
  assign n606 = ~pi129 & ~n605;
  assign n607 = ~pi3 & n606;
  assign n608 = n448 & ~n605;
  assign n609 = pi0 & ~pi113;
  assign n610 = pi0 & ~pi123;
  assign n611 = ~pi113 & n610;
  assign n612 = ~pi123 & n609;
  assign n613 = n2505 & n2520;
  assign n614 = ~pi11 & ~pi12;
  assign n615 = ~pi8 & ~pi17;
  assign n616 = n614 & n615;
  assign n617 = ~pi21 & n2520;
  assign n618 = n616 & n617;
  assign n619 = n535 & n618;
  assign n620 = n2517 & n613;
  assign n621 = ~pi61 & ~pi118;
  assign n622 = ~n2528 & n621;
  assign n623 = ~n2527 & ~n622;
  assign po18 = ~pi129 & ~n623;
  assign n625 = ~pi5 & ~pi22;
  assign n626 = ~pi17 & n625;
  assign n627 = n467 & n625;
  assign n628 = ~pi17 & n627;
  assign n629 = n467 & n626;
  assign n630 = n2520 & n2529;
  assign n631 = ~pi14 & n528;
  assign n632 = ~pi9 & ~pi11;
  assign n633 = n456 & n632;
  assign n634 = n631 & n633;
  assign n635 = ~pi13 & ~pi14;
  assign n636 = ~pi6 & ~pi7;
  assign n637 = n635 & n636;
  assign n638 = ~pi12 & n2506;
  assign n639 = n637 & n638;
  assign n640 = n625 & n632;
  assign n641 = n2520 & n640;
  assign n642 = n639 & n641;
  assign n643 = n456 & n528;
  assign n644 = ~pi14 & ~pi17;
  assign n645 = n632 & n644;
  assign n646 = n627 & n645;
  assign n647 = n643 & n646;
  assign n648 = n2520 & n647;
  assign n649 = n630 & n634;
  assign n650 = pi54 & ~n2530;
  assign n651 = ~pi0 & ~n650;
  assign n652 = pi7 & ~n456;
  assign n653 = ~n643 & ~n652;
  assign n654 = ~pi14 & ~n653;
  assign n655 = pi14 & ~n643;
  assign n656 = ~pi7 & n456;
  assign n657 = pi8 & pi21;
  assign n658 = ~pi13 & ~n657;
  assign n659 = ~n656 & ~n658;
  assign n660 = ~pi10 & ~n659;
  assign n661 = ~n655 & n660;
  assign n662 = ~pi7 & pi13;
  assign n663 = n456 & n662;
  assign n664 = ~n652 & ~n656;
  assign n665 = n658 & n664;
  assign n666 = ~n663 & ~n665;
  assign n667 = ~pi14 & ~n666;
  assign n668 = ~pi13 & pi14;
  assign n669 = n656 & n668;
  assign n670 = ~n667 & ~n669;
  assign n671 = ~pi10 & ~n670;
  assign n672 = ~pi14 & ~n659;
  assign n673 = ~n643 & ~n672;
  assign n674 = ~pi10 & ~n654;
  assign n675 = ~n673 & n674;
  assign n676 = ~n654 & n661;
  assign n677 = ~pi14 & n456;
  assign n678 = pi10 & n528;
  assign n679 = pi10 & n635;
  assign n680 = n656 & n679;
  assign n681 = n677 & n678;
  assign n682 = ~n2531 & ~n2532;
  assign n683 = n625 & ~n682;
  assign n684 = n2520 & n683;
  assign n685 = ~pi17 & n684;
  assign n686 = n467 & n685;
  assign n687 = n630 & ~n682;
  assign n688 = ~pi56 & ~n625;
  assign n689 = n632 & ~n688;
  assign n690 = ~n2533 & n689;
  assign n691 = ~pi56 & n625;
  assign n692 = ~n632 & ~n691;
  assign n693 = pi54 & ~n692;
  assign n694 = n625 & ~n632;
  assign n695 = ~pi56 & n694;
  assign n696 = ~n2533 & ~n688;
  assign n697 = n632 & ~n696;
  assign n698 = ~n695 & ~n697;
  assign n699 = pi54 & ~n698;
  assign n700 = ~n690 & n693;
  assign n701 = ~n651 & ~n2534;
  assign n702 = ~pi129 & ~n701;
  assign n703 = ~pi3 & n702;
  assign n704 = n448 & ~n701;
  assign n705 = n450 & n614;
  assign n706 = n677 & n705;
  assign n707 = n529 & n706;
  assign n708 = n456 & n614;
  assign n709 = n2520 & n708;
  assign n710 = ~pi14 & n529;
  assign n711 = n450 & n710;
  assign n712 = n709 & n711;
  assign n713 = n2520 & n707;
  assign n714 = n585 & ~n2536;
  assign n715 = ~pi1 & ~n714;
  assign n716 = ~n467 & n468;
  assign n717 = n467 & ~n468;
  assign n718 = ~n716 & ~n717;
  assign n719 = ~n465 & ~n466;
  assign n720 = ~pi13 & ~n719;
  assign n721 = pi5 & ~n467;
  assign n722 = ~n520 & ~n721;
  assign n723 = pi6 & pi12;
  assign n724 = ~pi7 & ~n723;
  assign n725 = n722 & n724;
  assign n726 = pi7 & n520;
  assign n727 = ~n725 & ~n726;
  assign n728 = ~pi13 & ~n727;
  assign n729 = ~n718 & n720;
  assign n730 = n520 & n662;
  assign n731 = pi13 & n2507;
  assign n732 = ~pi9 & ~n2538;
  assign n733 = ~n467 & ~n468;
  assign n734 = ~pi13 & ~n733;
  assign n735 = ~n2507 & ~n734;
  assign n736 = ~n2516 & ~n719;
  assign n737 = ~n2537 & ~n2538;
  assign n738 = ~n735 & n736;
  assign n739 = ~pi9 & n2539;
  assign n740 = ~n2537 & n732;
  assign n741 = pi9 & ~n2516;
  assign n742 = ~pi14 & pi54;
  assign n743 = n450 & n742;
  assign n744 = n2520 & n743;
  assign n745 = n2505 & n744;
  assign n746 = ~n741 & n743;
  assign n747 = n613 & n746;
  assign n748 = ~n741 & n745;
  assign n749 = ~pi9 & ~n2539;
  assign n750 = pi9 & n2516;
  assign n751 = ~n749 & ~n750;
  assign n752 = n2520 & ~n751;
  assign n753 = n2505 & n752;
  assign n754 = n742 & n753;
  assign n755 = n450 & n754;
  assign n756 = ~n2540 & n2541;
  assign n757 = ~n715 & ~n2542;
  assign n758 = ~pi129 & ~n757;
  assign n759 = ~pi3 & n758;
  assign n760 = n448 & ~n757;
  assign n761 = pi4 & ~pi54;
  assign n762 = ~pi17 & ~pi18;
  assign n763 = ~pi18 & ~pi21;
  assign n764 = n615 & n763;
  assign n765 = ~pi18 & n2506;
  assign n766 = n456 & n762;
  assign n767 = ~pi11 & n473;
  assign n768 = n471 & n767;
  assign n769 = n2544 & n768;
  assign n770 = n2505 & n2519;
  assign n771 = pi10 & ~pi22;
  assign n772 = n451 & n771;
  assign n773 = n2516 & n772;
  assign n774 = n2545 & n773;
  assign n775 = ~n761 & ~n774;
  assign n776 = ~pi129 & ~n775;
  assign n777 = ~pi3 & n776;
  assign n778 = n448 & ~n775;
  assign n779 = pi7 & ~pi54;
  assign n780 = pi8 & ~pi17;
  assign n781 = ~pi21 & n780;
  assign n782 = n2519 & n781;
  assign n783 = ~pi6 & n614;
  assign n784 = n468 & n783;
  assign n785 = ~pi11 & n2507;
  assign n786 = n453 & n2547;
  assign n787 = n763 & n780;
  assign n788 = ~pi7 & n473;
  assign n789 = n471 & n788;
  assign n790 = n787 & n789;
  assign n791 = ~pi5 & n783;
  assign n792 = n453 & n791;
  assign n793 = n790 & n792;
  assign n794 = n782 & n786;
  assign n795 = ~n779 & ~n2548;
  assign n796 = ~pi129 & ~n795;
  assign n797 = ~pi3 & n796;
  assign n798 = n448 & ~n795;
  assign n799 = pi8 & ~pi54;
  assign n800 = ~pi17 & pi21;
  assign n801 = n454 & n800;
  assign n802 = ~pi11 & pi21;
  assign n803 = n762 & n802;
  assign n804 = ~pi8 & n473;
  assign n805 = n471 & n804;
  assign n806 = n803 & n805;
  assign n807 = n2519 & n801;
  assign n808 = n539 & n801;
  assign n809 = n2517 & n2550;
  assign n810 = ~n799 & ~n2551;
  assign n811 = ~pi129 & ~n810;
  assign n812 = ~pi3 & n811;
  assign n813 = n448 & ~n810;
  assign n814 = pi9 & ~pi54;
  assign n815 = n2516 & n2544;
  assign n816 = n450 & n542;
  assign n817 = pi11 & n451;
  assign n818 = n816 & n817;
  assign n819 = n450 & n635;
  assign n820 = pi11 & n468;
  assign n821 = n467 & n820;
  assign n822 = n819 & n821;
  assign n823 = ~pi9 & n473;
  assign n824 = n471 & n823;
  assign n825 = n2544 & n824;
  assign n826 = n822 & n825;
  assign n827 = n2516 & n817;
  assign n828 = n2544 & n816;
  assign n829 = n827 & n828;
  assign n830 = n815 & n818;
  assign n831 = ~n814 & ~n2553;
  assign n832 = ~pi129 & ~n831;
  assign n833 = ~pi3 & n832;
  assign n834 = n448 & ~n831;
  assign n835 = pi10 & ~pi54;
  assign n836 = ~pi11 & pi14;
  assign n837 = n2516 & n836;
  assign n838 = n668 & n2547;
  assign n839 = ~pi9 & n2544;
  assign n840 = n816 & n839;
  assign n841 = ~pi10 & n473;
  assign n842 = n471 & n841;
  assign n843 = n2544 & n842;
  assign n844 = ~pi9 & ~pi22;
  assign n845 = n668 & n844;
  assign n846 = n2547 & n845;
  assign n847 = n843 & n846;
  assign n848 = n816 & n2555;
  assign n849 = n839 & n848;
  assign n850 = n2555 & n840;
  assign n851 = ~n835 & ~n2556;
  assign n852 = ~pi129 & ~n851;
  assign n853 = ~pi3 & n852;
  assign n854 = n448 & ~n851;
  assign n855 = pi11 & ~pi54;
  assign n856 = ~pi10 & ~pi14;
  assign n857 = pi22 & n856;
  assign n858 = ~pi10 & ~pi11;
  assign n859 = pi22 & n858;
  assign n860 = n451 & n859;
  assign n861 = n632 & n857;
  assign n862 = n542 & n2558;
  assign n863 = ~pi10 & pi22;
  assign n864 = n451 & n863;
  assign n865 = n2516 & n864;
  assign n866 = n2545 & n865;
  assign n867 = n815 & n862;
  assign n868 = ~n855 & ~n2559;
  assign n869 = ~pi129 & ~n868;
  assign n870 = ~pi3 & n869;
  assign n871 = n448 & ~n868;
  assign n872 = pi12 & ~pi54;
  assign n873 = pi18 & n542;
  assign n874 = n2505 & n873;
  assign n875 = ~pi12 & n473;
  assign n876 = n471 & n875;
  assign n877 = pi18 & n2506;
  assign n878 = n876 & n877;
  assign n879 = ~pi11 & n535;
  assign n880 = n878 & n879;
  assign n881 = ~pi12 & pi18;
  assign n882 = n542 & n881;
  assign n883 = n2505 & n882;
  assign n884 = n535 & n883;
  assign n885 = n2517 & n874;
  assign n886 = ~n872 & ~n2561;
  assign n887 = ~pi129 & ~n886;
  assign n888 = ~pi3 & n887;
  assign n889 = n448 & ~n886;
  assign n890 = pi14 & ~pi54;
  assign n891 = pi13 & ~pi19;
  assign n892 = n544 & n891;
  assign n893 = n743 & n892;
  assign n894 = n2547 & n893;
  assign n895 = ~pi16 & n742;
  assign n896 = n473 & n895;
  assign n897 = n2544 & n896;
  assign n898 = ~pi9 & pi13;
  assign n899 = n450 & n898;
  assign n900 = n2547 & n899;
  assign n901 = n897 & n900;
  assign n902 = n839 & n894;
  assign n903 = ~n890 & ~n2563;
  assign n904 = ~pi129 & ~n903;
  assign n905 = ~pi3 & n904;
  assign n906 = n448 & ~n903;
  assign n907 = pi16 & ~pi54;
  assign n908 = pi6 & ~pi13;
  assign n909 = n468 & n908;
  assign n910 = ~pi5 & pi6;
  assign n911 = pi6 & ~pi12;
  assign n912 = ~pi5 & n911;
  assign n913 = ~pi12 & n910;
  assign n914 = n528 & n2565;
  assign n915 = n452 & n914;
  assign n916 = n530 & n909;
  assign n917 = n2545 & n2566;
  assign n918 = ~n907 & ~n917;
  assign n919 = ~pi129 & ~n918;
  assign n920 = ~pi3 & n919;
  assign n921 = n448 & ~n918;
  assign n922 = pi18 & ~pi54;
  assign n923 = pi16 & n585;
  assign n924 = n2508 & n923;
  assign n925 = pi16 & pi54;
  assign n926 = n2508 & n925;
  assign n927 = n2505 & n926;
  assign n928 = n457 & n924;
  assign n929 = pi16 & n586;
  assign n930 = n538 & n929;
  assign n931 = n2517 & n2568;
  assign n932 = ~n922 & ~n2569;
  assign n933 = ~pi129 & ~n932;
  assign n934 = ~pi3 & n933;
  assign n935 = n448 & ~n932;
  assign n936 = pi19 & ~pi54;
  assign n937 = pi17 & n457;
  assign n938 = n2519 & n937;
  assign n939 = n539 & n937;
  assign n940 = n2517 & n938;
  assign n941 = ~n936 & ~n2571;
  assign n942 = ~pi129 & ~n941;
  assign n943 = ~pi3 & n942;
  assign n944 = n448 & ~n941;
  assign n945 = pi2 & n2503;
  assign n946 = pi20 & ~n2495;
  assign n947 = ~n945 & ~n946;
  assign n948 = pi82 & ~n947;
  assign n949 = pi20 & n389;
  assign n950 = ~pi71 & ~n291;
  assign n951 = ~n291 & ~n442;
  assign n952 = ~pi71 & n951;
  assign n953 = ~n442 & n950;
  assign n954 = ~n949 & ~n2573;
  assign n955 = ~n948 & ~n949;
  assign n956 = ~n2573 & n955;
  assign n957 = ~n948 & n954;
  assign po35 = ~pi129 & ~n2574;
  assign n959 = pi21 & ~pi54;
  assign n960 = ~pi18 & pi19;
  assign n961 = n544 & n960;
  assign n962 = n454 & n762;
  assign n963 = ~pi21 & pi54;
  assign n964 = pi19 & n963;
  assign n965 = n544 & n964;
  assign n966 = n962 & n965;
  assign n967 = pi19 & ~pi21;
  assign n968 = ~pi18 & n967;
  assign n969 = n454 & n585;
  assign n970 = n544 & n969;
  assign n971 = n968 & n970;
  assign n972 = n586 & n961;
  assign n973 = n2517 & n2575;
  assign n974 = ~n959 & ~n973;
  assign n975 = ~pi129 & ~n974;
  assign n976 = ~pi3 & n975;
  assign n977 = n448 & ~n974;
  assign n978 = pi22 & ~pi54;
  assign n979 = pi5 & ~pi6;
  assign n980 = n614 & n979;
  assign n981 = n631 & n980;
  assign n982 = n450 & n528;
  assign n983 = n614 & n982;
  assign n984 = ~pi14 & n979;
  assign n985 = n542 & n984;
  assign n986 = n983 & n985;
  assign n987 = n816 & n981;
  assign n988 = ~pi22 & n473;
  assign n989 = n471 & n988;
  assign n990 = n2544 & n989;
  assign n991 = ~pi9 & ~pi10;
  assign n992 = n635 & n991;
  assign n993 = pi5 & ~pi7;
  assign n994 = n783 & n993;
  assign n995 = n992 & n994;
  assign n996 = n990 & n995;
  assign n997 = n839 & n2577;
  assign n998 = ~n978 & ~n2578;
  assign n999 = ~pi129 & ~n998;
  assign n1000 = ~pi3 & n999;
  assign n1001 = n448 & ~n998;
  assign n1002 = n368 & n369;
  assign n1003 = n2482 & n1002;
  assign n1004 = n2484 & n2486;
  assign n1005 = pi82 & ~n2580;
  assign n1006 = pi63 & ~n291;
  assign n1007 = ~n291 & ~n1005;
  assign n1008 = pi63 & n1007;
  assign n1009 = ~n1005 & n1006;
  assign n1010 = pi82 & ~n2486;
  assign n1011 = n291 & ~n1010;
  assign n1012 = ~n388 & ~n1011;
  assign n1013 = ~pi24 & ~n1012;
  assign n1014 = pi24 & pi82;
  assign n1015 = n293 & n1014;
  assign n1016 = n394 & n1015;
  assign n1017 = ~pi44 & pi82;
  assign n1018 = pi24 & ~pi45;
  assign n1019 = n1017 & n1018;
  assign n1020 = n414 & n1019;
  assign n1021 = pi24 & n1017;
  assign n1022 = n2485 & n1021;
  assign n1023 = n2478 & n1022;
  assign n1024 = n2485 & n1016;
  assign n1025 = ~pi129 & ~n2582;
  assign n1026 = ~n1013 & n1025;
  assign n1027 = ~n2581 & n1025;
  assign n1028 = ~n1013 & n1027;
  assign n1029 = ~n2581 & n1026;
  assign n1030 = ~pi53 & pi58;
  assign n1031 = pi53 & ~pi58;
  assign n1032 = ~n1030 & ~n1031;
  assign n1033 = ~pi96 & ~pi110;
  assign n1034 = ~pi85 & ~n1033;
  assign n1035 = pi85 & ~pi116;
  assign n1036 = pi100 & ~n1035;
  assign n1037 = pi85 & pi116;
  assign n1038 = ~pi85 & ~pi110;
  assign n1039 = ~pi96 & n1038;
  assign n1040 = ~n1037 & ~n1039;
  assign n1041 = pi100 & ~n1040;
  assign n1042 = ~n1034 & n1036;
  assign n1043 = pi25 & ~pi116;
  assign n1044 = pi85 & n1043;
  assign n1045 = pi25 & n1035;
  assign n1046 = ~n2584 & ~n2585;
  assign n1047 = ~pi26 & ~n1046;
  assign n1048 = ~pi39 & ~pi52;
  assign n1049 = ~pi51 & ~pi52;
  assign n1050 = ~pi39 & n1049;
  assign n1051 = ~pi51 & n1048;
  assign n1052 = pi116 & n2586;
  assign n1053 = ~pi85 & ~n1052;
  assign n1054 = pi26 & n1053;
  assign n1055 = ~pi25 & ~pi116;
  assign n1056 = n1054 & ~n1055;
  assign n1057 = ~n1047 & ~n1056;
  assign n1058 = ~pi27 & ~n1057;
  assign n1059 = ~n1043 & ~n1052;
  assign n1060 = pi27 & ~n1059;
  assign n1061 = pi27 & ~n2586;
  assign n1062 = ~pi95 & ~pi100;
  assign n1063 = ~pi97 & n1062;
  assign n1064 = ~pi110 & ~n1063;
  assign n1065 = pi25 & ~n1064;
  assign n1066 = ~n1061 & n1065;
  assign n1067 = ~n1060 & ~n1066;
  assign n1068 = ~pi26 & ~pi85;
  assign n1069 = ~n1067 & n1068;
  assign n1070 = pi26 & n1043;
  assign n1071 = pi26 & pi116;
  assign n1072 = ~n1065 & ~n1071;
  assign n1073 = ~n2586 & ~n1072;
  assign n1074 = ~n1070 & ~n1073;
  assign n1075 = ~pi85 & ~n1074;
  assign n1076 = ~n1047 & ~n1075;
  assign n1077 = ~pi27 & ~n1076;
  assign n1078 = n2586 & n1065;
  assign n1079 = ~n1060 & ~n1078;
  assign n1080 = n1068 & ~n1079;
  assign n1081 = ~n1077 & ~n1080;
  assign n1082 = ~n1058 & ~n1069;
  assign n1083 = ~pi53 & ~n2587;
  assign n1084 = n1032 & ~n1083;
  assign n1085 = ~pi53 & ~pi58;
  assign n1086 = ~pi27 & ~pi85;
  assign n1087 = pi25 & ~pi26;
  assign n1088 = ~pi116 & n1087;
  assign n1089 = ~pi26 & n1043;
  assign n1090 = n1086 & n2588;
  assign n1091 = ~n1085 & ~n1090;
  assign n1092 = n448 & ~n1091;
  assign n1093 = pi53 & ~pi85;
  assign n1094 = ~pi27 & n1093;
  assign n1095 = n2588 & n1094;
  assign n1096 = ~n1083 & ~n1095;
  assign n1097 = ~pi58 & ~n1096;
  assign n1098 = n1030 & n1086;
  assign n1099 = n2588 & n1098;
  assign n1100 = ~n1097 & ~n1099;
  assign n1101 = ~pi129 & ~n1100;
  assign n1102 = ~pi3 & n1101;
  assign n1103 = n448 & ~n1100;
  assign n1104 = ~n1084 & n1092;
  assign n1105 = ~pi26 & ~n2586;
  assign n1106 = ~pi27 & n2586;
  assign n1107 = ~n1105 & ~n1106;
  assign n1108 = ~n1064 & ~n1107;
  assign n1109 = ~pi26 & ~pi27;
  assign n1110 = pi26 & pi27;
  assign n1111 = pi26 & ~pi27;
  assign n1112 = ~pi26 & pi27;
  assign n1113 = ~n1111 & ~n1112;
  assign n1114 = ~n1109 & ~n1110;
  assign n1115 = ~pi116 & ~n2590;
  assign n1116 = ~n1108 & ~n1115;
  assign n1117 = pi28 & ~n1116;
  assign n1118 = ~pi26 & pi95;
  assign n1119 = ~pi100 & n1118;
  assign n1120 = pi95 & ~pi96;
  assign n1121 = ~pi26 & ~pi100;
  assign n1122 = ~pi110 & n1121;
  assign n1123 = n1120 & n1122;
  assign n1124 = n1033 & n1119;
  assign n1125 = pi26 & n1052;
  assign n1126 = n2586 & n1071;
  assign n1127 = ~n2591 & ~n2592;
  assign n1128 = ~pi27 & ~n1127;
  assign n1129 = pi27 & pi116;
  assign n1130 = n1105 & n1129;
  assign n1131 = ~pi85 & ~n1130;
  assign n1132 = ~n1128 & n1131;
  assign n1133 = ~n1117 & n1132;
  assign n1134 = pi100 & pi116;
  assign n1135 = ~pi28 & ~pi116;
  assign n1136 = n1109 & ~n1135;
  assign n1137 = ~n1134 & n1136;
  assign n1138 = pi85 & ~n1137;
  assign n1139 = ~pi53 & ~n1138;
  assign n1140 = ~n1128 & ~n1130;
  assign n1141 = ~n1117 & n1140;
  assign n1142 = ~pi85 & ~n1141;
  assign n1143 = pi28 & ~pi116;
  assign n1144 = ~pi100 & pi116;
  assign n1145 = ~n1143 & ~n1144;
  assign n1146 = pi85 & ~n1145;
  assign n1147 = n1109 & n1146;
  assign n1148 = ~n1142 & ~n1147;
  assign n1149 = ~pi53 & ~n1148;
  assign n1150 = ~n1133 & n1139;
  assign n1151 = ~pi27 & pi28;
  assign n1152 = ~pi116 & n1151;
  assign n1153 = ~pi26 & n1093;
  assign n1154 = pi53 & n1068;
  assign n1155 = n1152 & n2594;
  assign n1156 = ~n2593 & ~n1155;
  assign n1157 = ~pi58 & ~n1156;
  assign n1158 = n1030 & n1068;
  assign n1159 = ~pi26 & ~pi53;
  assign n1160 = ~pi85 & n1159;
  assign n1161 = pi58 & n1152;
  assign n1162 = n1160 & n1161;
  assign n1163 = n1152 & n1158;
  assign n1164 = ~n1157 & ~n2595;
  assign n1165 = ~pi129 & ~n1164;
  assign n1166 = ~pi3 & n1165;
  assign n1167 = n448 & ~n1164;
  assign n1168 = pi27 & n1053;
  assign n1169 = ~pi85 & pi95;
  assign n1170 = n1033 & n1169;
  assign n1171 = pi95 & ~n1035;
  assign n1172 = n1033 & n1171;
  assign n1173 = ~n1037 & ~n1172;
  assign n1174 = ~n1037 & ~n1170;
  assign n1175 = ~pi100 & ~n1129;
  assign n1176 = ~pi110 & ~n1035;
  assign n1177 = ~n1129 & n1176;
  assign n1178 = n1120 & n1177;
  assign n1179 = ~pi27 & n1037;
  assign n1180 = ~n1178 & ~n1179;
  assign n1181 = ~pi100 & ~n1180;
  assign n1182 = ~n2597 & n1175;
  assign n1183 = ~n1168 & ~n2598;
  assign n1184 = ~pi26 & n448;
  assign n1185 = n1085 & n1184;
  assign n1186 = ~pi129 & ~n1183;
  assign n1187 = ~pi3 & n1186;
  assign n1188 = ~pi26 & n1085;
  assign n1189 = n1187 & n1188;
  assign n1190 = ~n1183 & n1185;
  assign n1191 = ~n1071 & n1176;
  assign n1192 = ~pi96 & n1191;
  assign n1193 = ~pi26 & n1037;
  assign n1194 = ~n1192 & ~n1193;
  assign n1195 = pi100 & ~n1194;
  assign n1196 = n2584 & ~n1071;
  assign n1197 = ~n1054 & ~n2600;
  assign n1198 = ~pi27 & ~pi53;
  assign n1199 = ~pi58 & n1198;
  assign n1200 = n448 & n1199;
  assign n1201 = ~pi129 & ~n1197;
  assign n1202 = ~pi3 & n1201;
  assign n1203 = n1199 & n1202;
  assign n1204 = ~n1197 & n1200;
  assign n1205 = pi97 & ~n1033;
  assign n1206 = ~pi29 & ~pi97;
  assign n1207 = n1062 & ~n1206;
  assign n1208 = pi97 & ~pi110;
  assign n1209 = ~pi96 & n1208;
  assign n1210 = pi97 & n1033;
  assign n1211 = pi29 & ~pi97;
  assign n1212 = ~n2602 & ~n1211;
  assign n1213 = n1062 & ~n1212;
  assign n1214 = ~n1205 & n1207;
  assign n1215 = pi29 & pi110;
  assign n1216 = ~pi58 & ~n1215;
  assign n1217 = pi29 & ~n1064;
  assign n1218 = n1062 & n2602;
  assign n1219 = ~pi58 & ~n1218;
  assign n1220 = ~n1217 & n1219;
  assign n1221 = ~n2603 & n1216;
  assign n1222 = pi97 & pi116;
  assign n1223 = pi29 & ~pi116;
  assign n1224 = pi58 & ~n1223;
  assign n1225 = pi58 & ~n1222;
  assign n1226 = ~n1223 & n1225;
  assign n1227 = ~n1222 & n1224;
  assign n1228 = ~pi53 & ~n2605;
  assign n1229 = ~n2603 & ~n1215;
  assign n1230 = ~pi58 & ~n1229;
  assign n1231 = ~n1222 & ~n1223;
  assign n1232 = pi58 & ~n1231;
  assign n1233 = ~n1230 & ~n1232;
  assign n1234 = ~pi53 & ~n1233;
  assign n1235 = ~n2604 & n1228;
  assign n1236 = n1031 & n1223;
  assign n1237 = ~n2606 & ~n1236;
  assign n1238 = ~pi27 & ~n1237;
  assign n1239 = pi27 & n1085;
  assign n1240 = pi27 & n1223;
  assign n1241 = n1085 & n1240;
  assign n1242 = n1223 & n1239;
  assign n1243 = ~n1238 & ~n2607;
  assign n1244 = ~pi85 & ~n1243;
  assign n1245 = pi85 & n1223;
  assign n1246 = pi85 & n1199;
  assign n1247 = n1223 & n1246;
  assign n1248 = n1199 & n1245;
  assign n1249 = ~n1244 & ~n2608;
  assign n1250 = ~pi26 & ~n1249;
  assign n1251 = pi26 & n1085;
  assign n1252 = n1085 & n1086;
  assign n1253 = pi26 & n1252;
  assign n1254 = ~pi85 & n1085;
  assign n1255 = n1111 & n1254;
  assign n1256 = n1086 & n1251;
  assign n1257 = n1223 & n2609;
  assign n1258 = ~n1250 & ~n1257;
  assign n1259 = ~pi129 & ~n1258;
  assign n1260 = ~pi3 & n1259;
  assign n1261 = n448 & ~n1258;
  assign n1262 = pi82 & ~n302;
  assign n1263 = ~pi45 & n2487;
  assign n1264 = n2488 & n367;
  assign n1265 = n369 & n370;
  assign n1266 = n339 & n376;
  assign n1267 = n1265 & n1266;
  assign n1268 = n2499 & n2611;
  assign n1269 = n333 & n2491;
  assign n1270 = ~pi50 & n2612;
  assign n1271 = n2501 & n2611;
  assign n1272 = pi82 & ~n2613;
  assign n1273 = n291 & ~n1272;
  assign n1274 = ~n1262 & ~n1273;
  assign n1275 = ~pi38 & ~n1274;
  assign n1276 = n2496 & n2611;
  assign n1277 = ~pi43 & n2492;
  assign n1278 = n302 & n2477;
  assign n1279 = ~pi50 & n302;
  assign n1280 = n333 & n1279;
  assign n1281 = n2491 & n1280;
  assign n1282 = n309 & n2491;
  assign n1283 = n308 & n2492;
  assign n1284 = n304 & n2616;
  assign n1285 = n2614 & n1278;
  assign n1286 = pi82 & ~n2615;
  assign n1287 = pi74 & ~n291;
  assign n1288 = ~n291 & ~n1286;
  assign n1289 = pi74 & n1288;
  assign n1290 = ~n1286 & n1287;
  assign n1291 = pi38 & n316;
  assign n1292 = ~pi42 & n1017;
  assign n1293 = ~pi40 & n1292;
  assign n1294 = pi38 & n1293;
  assign n1295 = n1017 & n1291;
  assign n1296 = ~pi129 & ~n2618;
  assign n1297 = ~n2617 & n1296;
  assign po53 = ~n1275 & n1297;
  assign n1299 = pi82 & ~n293;
  assign n1300 = n2489 & n2614;
  assign n1301 = pi82 & ~n1300;
  assign n1302 = n291 & ~n1301;
  assign n1303 = ~n1299 & ~n1302;
  assign n1304 = ~pi40 & ~n1303;
  assign n1305 = n293 & n297;
  assign n1306 = n333 & n1305;
  assign n1307 = n293 & n1300;
  assign n1308 = n293 & n2474;
  assign n1309 = n2616 & n1308;
  assign n1310 = n2491 & n1306;
  assign n1311 = pi82 & ~n2619;
  assign n1312 = pi73 & ~n291;
  assign n1313 = ~n291 & ~n1311;
  assign n1314 = pi73 & n1313;
  assign n1315 = ~n1311 & n1312;
  assign n1316 = pi40 & pi82;
  assign n1317 = pi40 & n1292;
  assign n1318 = n293 & n1316;
  assign n1319 = ~pi129 & ~n2621;
  assign n1320 = ~n2620 & n1319;
  assign po55 = ~n1304 & n1320;
  assign n1322 = pi82 & ~n2476;
  assign n1323 = pi82 & ~n2614;
  assign n1324 = n291 & ~n1323;
  assign n1325 = ~n1322 & ~n1324;
  assign n1326 = ~pi41 & ~n1325;
  assign n1327 = n295 & n332;
  assign n1328 = n2476 & n332;
  assign n1329 = n311 & n1327;
  assign n1330 = n2476 & n2614;
  assign n1331 = n2491 & n2622;
  assign n1332 = pi82 & ~n2623;
  assign n1333 = pi76 & ~n291;
  assign n1334 = ~n291 & ~n1332;
  assign n1335 = pi76 & n1334;
  assign n1336 = ~n1332 & n1333;
  assign n1337 = pi41 & pi82;
  assign n1338 = pi41 & n1292;
  assign n1339 = n293 & n1337;
  assign n1340 = n2475 & n2625;
  assign n1341 = ~pi129 & ~n1340;
  assign n1342 = ~n2624 & n1341;
  assign n1343 = ~n1326 & n1341;
  assign n1344 = ~n2624 & n1343;
  assign n1345 = ~n1326 & n1342;
  assign n1346 = n2475 & n309;
  assign n1347 = n2475 & n2616;
  assign n1348 = n2491 & n1346;
  assign n1349 = pi82 & ~n2627;
  assign n1350 = ~pi72 & ~n291;
  assign n1351 = ~n1349 & ~n1350;
  assign n1352 = ~n1299 & ~n1351;
  assign n1353 = pi42 & ~n1017;
  assign n1354 = ~n292 & n1353;
  assign n1355 = ~n1352 & ~n1354;
  assign n1356 = pi44 & pi82;
  assign n1357 = n291 & ~n1349;
  assign n1358 = ~n1356 & ~n1357;
  assign n1359 = ~pi42 & ~n1358;
  assign n1360 = n333 & n420;
  assign n1361 = n2491 & n1360;
  assign n1362 = ~pi44 & n2627;
  assign n1363 = pi82 & ~n2628;
  assign n1364 = pi72 & ~n291;
  assign n1365 = ~n291 & ~n1363;
  assign n1366 = pi72 & n1365;
  assign n1367 = ~n1363 & n1364;
  assign n1368 = pi42 & n1017;
  assign n1369 = ~pi129 & ~n1368;
  assign n1370 = ~n2629 & n1369;
  assign n1371 = ~n1359 & n1370;
  assign n1372 = ~pi129 & ~n1355;
  assign n1373 = pi82 & ~n2481;
  assign n1374 = pi82 & ~n2492;
  assign n1375 = n291 & ~n1374;
  assign n1376 = ~n1373 & ~n1375;
  assign n1377 = ~pi43 & ~n1376;
  assign n1378 = ~pi47 & n2481;
  assign n1379 = n2491 & n1378;
  assign n1380 = n2481 & n2492;
  assign n1381 = pi82 & ~n2631;
  assign n1382 = pi77 & ~n291;
  assign n1383 = ~n291 & ~n1381;
  assign n1384 = pi77 & n1383;
  assign n1385 = ~n1381 & n1382;
  assign n1386 = pi43 & n316;
  assign n1387 = pi43 & n1293;
  assign n1388 = n1017 & n1386;
  assign n1389 = n2489 & n1293;
  assign n1390 = pi43 & n1389;
  assign n1391 = n2489 & n2633;
  assign n1392 = ~pi129 & ~n2634;
  assign n1393 = ~n2632 & n1392;
  assign po58 = ~n1377 & n1393;
  assign n1395 = n2478 & n333;
  assign n1396 = ~pi42 & n2627;
  assign n1397 = n2491 & n1395;
  assign n1398 = pi82 & ~n2635;
  assign n1399 = ~pi67 & ~n291;
  assign n1400 = pi44 & n291;
  assign n1401 = pi67 & ~n291;
  assign n1402 = ~pi44 & n291;
  assign n1403 = ~n1401 & ~n1402;
  assign n1404 = ~n1399 & ~n1400;
  assign n1405 = ~n1398 & ~n2636;
  assign n1406 = ~pi129 & ~n1356;
  assign po59 = ~n1405 & n1406;
  assign n1408 = ~pi48 & n2487;
  assign n1409 = n2482 & n377;
  assign n1410 = n2483 & n1408;
  assign n1411 = pi82 & ~n2637;
  assign n1412 = pi68 & ~n291;
  assign n1413 = ~n291 & ~n1411;
  assign n1414 = pi68 & n1413;
  assign n1415 = ~n1411 & n1412;
  assign n1416 = pi82 & ~n2487;
  assign n1417 = n291 & ~n1416;
  assign n1418 = pi82 & ~n2500;
  assign n1419 = ~n1417 & ~n1418;
  assign n1420 = ~pi45 & ~n1419;
  assign n1421 = pi45 & pi82;
  assign n1422 = pi45 & n2479;
  assign n1423 = n1017 & n1422;
  assign n1424 = n311 & n1421;
  assign n1425 = n2500 & n1421;
  assign n1426 = n2501 & n2639;
  assign n1427 = ~pi129 & ~n2640;
  assign n1428 = ~n1420 & n1427;
  assign n1429 = ~n2638 & n1427;
  assign n1430 = ~n1420 & n1429;
  assign n1431 = ~n2638 & n1428;
  assign n1432 = pi82 & ~n2480;
  assign n1433 = pi82 & ~n2616;
  assign n1434 = n291 & ~n1433;
  assign n1435 = ~n1432 & ~n1434;
  assign n1436 = ~pi46 & ~n1435;
  assign n1437 = n2480 & n2616;
  assign n1438 = pi82 & ~n1437;
  assign n1439 = pi75 & ~n291;
  assign n1440 = ~n291 & ~n1438;
  assign n1441 = pi75 & n1440;
  assign n1442 = ~n1438 & n1439;
  assign n1443 = pi46 & n1017;
  assign n1444 = pi46 & pi82;
  assign n1445 = n2480 & n1444;
  assign n1446 = n2478 & n1443;
  assign n1447 = ~pi129 & ~n2643;
  assign n1448 = ~n2642 & n1447;
  assign po61 = ~n1436 & n1448;
  assign n1450 = n2482 & n2491;
  assign n1451 = pi82 & ~n1450;
  assign n1452 = pi64 & ~n291;
  assign n1453 = ~n291 & ~n1451;
  assign n1454 = pi64 & n1453;
  assign n1455 = ~n1451 & n1452;
  assign n1456 = pi82 & ~n2482;
  assign n1457 = pi82 & ~n2491;
  assign n1458 = n291 & ~n1457;
  assign n1459 = ~n1456 & ~n1458;
  assign n1460 = ~pi47 & ~n1459;
  assign n1461 = n2474 & n308;
  assign n1462 = pi47 & n316;
  assign n1463 = n1017 & n1462;
  assign n1464 = ~pi43 & pi47;
  assign n1465 = n1389 & n1464;
  assign n1466 = pi47 & n308;
  assign n1467 = n2474 & n1466;
  assign n1468 = n1293 & n1467;
  assign n1469 = n1461 & n1463;
  assign n1470 = ~pi129 & ~n2645;
  assign n1471 = ~n1460 & n1470;
  assign n1472 = ~n2644 & n1470;
  assign n1473 = ~n1460 & n1472;
  assign n1474 = ~n2644 & n1471;
  assign n1475 = ~pi2 & ~pi47;
  assign n1476 = n1265 & n1475;
  assign n1477 = n2482 & n1476;
  assign n1478 = n2483 & n2611;
  assign n1479 = pi82 & ~n2647;
  assign n1480 = pi62 & ~n291;
  assign n1481 = ~n291 & ~n1479;
  assign n1482 = pi62 & n1481;
  assign n1483 = ~n1479 & n1480;
  assign n1484 = pi82 & ~n2611;
  assign n1485 = n291 & ~n1484;
  assign n1486 = pi82 & ~n2483;
  assign n1487 = ~n1485 & ~n1486;
  assign n1488 = ~pi48 & ~n1487;
  assign n1489 = pi48 & n1017;
  assign n1490 = n2478 & n1489;
  assign n1491 = n2477 & n332;
  assign n1492 = pi48 & n2479;
  assign n1493 = n1017 & n1492;
  assign n1494 = n1491 & n1493;
  assign n1495 = pi48 & n332;
  assign n1496 = n1017 & n1495;
  assign n1497 = n2477 & n2479;
  assign n1498 = n1496 & n1497;
  assign n1499 = n333 & n1490;
  assign n1500 = ~pi129 & ~n2649;
  assign n1501 = ~n1488 & n1500;
  assign n1502 = ~n2648 & n1500;
  assign n1503 = ~n1488 & n1502;
  assign n1504 = ~n2648 & n1501;
  assign n1505 = pi49 & ~n2502;
  assign n1506 = ~n2498 & ~n1505;
  assign n1507 = ~n348 & n408;
  assign n1508 = n333 & n1507;
  assign n1509 = n307 & n1508;
  assign n1510 = ~n348 & n2498;
  assign n1511 = ~n1505 & ~n2651;
  assign n1512 = pi82 & ~n1511;
  assign n1513 = n1010 & ~n1506;
  assign n1514 = pi82 & ~n2498;
  assign n1515 = ~pi69 & ~n291;
  assign n1516 = ~n291 & ~n1514;
  assign n1517 = ~pi69 & n1516;
  assign n1518 = ~n1514 & n1515;
  assign n1519 = pi49 & n389;
  assign n1520 = ~n2653 & ~n1519;
  assign n1521 = ~n2652 & ~n1519;
  assign n1522 = ~n2653 & n1521;
  assign n1523 = ~n2652 & n1520;
  assign po64 = ~pi129 & ~n2654;
  assign n1525 = pi82 & ~n311;
  assign n1526 = pi82 & ~n2612;
  assign n1527 = n291 & ~n1526;
  assign n1528 = ~n1525 & ~n1527;
  assign n1529 = ~pi50 & ~n1528;
  assign n1530 = n311 & n333;
  assign n1531 = n296 & n302;
  assign n1532 = n2616 & n1531;
  assign n1533 = n2491 & n1530;
  assign n1534 = pi82 & ~n2655;
  assign n1535 = pi66 & ~n291;
  assign n1536 = ~n291 & ~n1534;
  assign n1537 = pi66 & n1536;
  assign n1538 = ~n1534 & n1535;
  assign n1539 = pi50 & pi82;
  assign n1540 = pi50 & n2479;
  assign n1541 = n1017 & n1540;
  assign n1542 = n311 & n1539;
  assign n1543 = ~pi129 & ~n2657;
  assign n1544 = ~n2656 & n1543;
  assign n1545 = ~n1529 & n1543;
  assign n1546 = ~n2656 & n1545;
  assign n1547 = ~n1529 & n1544;
  assign n1548 = ~pi129 & ~n2493;
  assign n1549 = ~pi96 & n1064;
  assign n1550 = ~pi59 & ~n1064;
  assign n1551 = n1085 & ~n1550;
  assign n1552 = ~n1549 & n1551;
  assign n1553 = pi59 & ~pi116;
  assign n1554 = ~n1032 & n1553;
  assign n1555 = ~pi116 & ~n1032;
  assign n1556 = ~n1064 & n1085;
  assign n1557 = ~n1555 & ~n1556;
  assign n1558 = pi59 & ~n1557;
  assign n1559 = pi96 & n1085;
  assign n1560 = n1064 & n1085;
  assign n1561 = pi96 & n1560;
  assign n1562 = n1064 & n1559;
  assign n1563 = ~n1558 & ~n2659;
  assign n1564 = ~n1552 & ~n1554;
  assign n1565 = ~pi85 & ~n2660;
  assign n1566 = pi85 & n1085;
  assign n1567 = n1553 & n1566;
  assign n1568 = ~n1565 & ~n1567;
  assign n1569 = ~pi27 & ~n1568;
  assign n1570 = pi27 & n1553;
  assign n1571 = pi27 & n1254;
  assign n1572 = n1553 & n1571;
  assign n1573 = n1254 & n1570;
  assign n1574 = ~n1569 & ~n2661;
  assign n1575 = ~pi26 & ~n1574;
  assign n1576 = n2609 & n1553;
  assign n1577 = ~n1575 & ~n1576;
  assign n1578 = ~pi129 & ~n1577;
  assign n1579 = ~pi3 & n1578;
  assign n1580 = n448 & ~n1577;
  assign n1581 = ~pi116 & n1031;
  assign n1582 = pi58 & pi116;
  assign n1583 = ~pi58 & ~pi110;
  assign n1584 = ~pi96 & n1583;
  assign n1585 = ~pi58 & n1033;
  assign n1586 = n1062 & n2663;
  assign n1587 = ~n1582 & ~n1586;
  assign n1588 = ~pi53 & pi97;
  assign n1589 = ~pi53 & ~n1587;
  assign n1590 = pi97 & n1589;
  assign n1591 = ~n1587 & n1588;
  assign n1592 = ~n1581 & ~n2664;
  assign n1593 = n1086 & n1184;
  assign n1594 = ~pi129 & ~n1592;
  assign n1595 = ~pi3 & n1594;
  assign n1596 = n1086 & n1595;
  assign n1597 = ~pi26 & n1596;
  assign n1598 = ~n1592 & n1593;
  assign n1599 = ~pi85 & ~n1063;
  assign n1600 = ~pi110 & n1599;
  assign n1601 = ~pi85 & n1064;
  assign n1602 = pi96 & n2666;
  assign n1603 = ~n1035 & ~n1602;
  assign n1604 = n1184 & n1199;
  assign n1605 = ~pi129 & ~n1603;
  assign n1606 = ~pi3 & n1605;
  assign n1607 = n1199 & n1606;
  assign n1608 = ~pi26 & n1607;
  assign n1609 = ~n1603 & n1604;
  assign n1610 = pi131 & pi132;
  assign n1611 = pi132 & pi133;
  assign n1612 = pi131 & n1611;
  assign n1613 = pi133 & n1610;
  assign n1614 = ~pi136 & ~pi137;
  assign n1615 = pi82 & pi138;
  assign n1616 = pi82 & ~pi137;
  assign n1617 = ~pi136 & n1616;
  assign n1618 = pi138 & n1617;
  assign n1619 = pi82 & ~pi136;
  assign n1620 = ~pi137 & pi138;
  assign n1621 = n1619 & n1620;
  assign n1622 = n1614 & n1615;
  assign n1623 = pi138 & n2668;
  assign n1624 = n1617 & n1623;
  assign n1625 = n2668 & n2669;
  assign n1626 = ~pi3 & ~pi110;
  assign n1627 = ~n2668 & ~n1626;
  assign n1628 = ~pi3 & ~n2668;
  assign n1629 = ~pi110 & n1628;
  assign n1630 = n2668 & ~n2669;
  assign n1631 = ~n1629 & ~n1630;
  assign n1632 = ~n2670 & ~n1627;
  assign n1633 = pi95 & ~n2671;
  assign n1634 = pi143 & n2670;
  assign n1635 = ~n1633 & ~n1634;
  assign po110 = ~pi129 & ~n1635;
  assign n1637 = pi96 & ~n2671;
  assign n1638 = pi146 & n2670;
  assign n1639 = ~n1637 & ~n1638;
  assign po111 = ~pi129 & ~n1639;
  assign n1641 = pi97 & ~n2671;
  assign n1642 = pi145 & n2670;
  assign n1643 = ~n1641 & ~n1642;
  assign po112 = ~pi129 & ~n1643;
  assign n1645 = pi100 & ~n2671;
  assign n1646 = pi144 & n2670;
  assign n1647 = ~n1645 & ~n1646;
  assign po115 = ~pi129 & ~n1647;
  assign n1649 = pi136 & ~pi137;
  assign n1650 = pi99 & n1649;
  assign n1651 = ~pi136 & pi137;
  assign n1652 = ~pi112 & n1651;
  assign n1653 = ~n1650 & ~n1652;
  assign n1654 = pi138 & ~n1653;
  assign n1655 = ~pi32 & pi136;
  assign n1656 = ~pi84 & ~pi136;
  assign n1657 = pi137 & ~n1656;
  assign n1658 = pi84 & ~pi136;
  assign n1659 = pi32 & pi136;
  assign n1660 = ~n1658 & ~n1659;
  assign n1661 = pi137 & ~n1660;
  assign n1662 = ~n1655 & n1657;
  assign n1663 = pi68 & pi136;
  assign n1664 = pi73 & ~pi136;
  assign n1665 = ~pi137 & ~n1664;
  assign n1666 = ~pi68 & pi136;
  assign n1667 = ~pi73 & ~pi136;
  assign n1668 = ~n1666 & ~n1667;
  assign n1669 = ~pi137 & ~n1668;
  assign n1670 = ~n1663 & n1665;
  assign n1671 = ~n2672 & ~n2673;
  assign n1672 = ~pi138 & ~n1671;
  assign n1673 = ~n1654 & ~n1672;
  assign n1674 = ~pi30 & ~pi109;
  assign n1675 = ~pi60 & pi109;
  assign n1676 = pi60 & pi109;
  assign n1677 = pi30 & ~pi109;
  assign n1678 = ~n1676 & ~n1677;
  assign n1679 = ~n1674 & ~n1675;
  assign n1680 = ~pi106 & ~n1677;
  assign n1681 = ~n1676 & n1680;
  assign n1682 = ~pi106 & n2674;
  assign n1683 = ~pi88 & pi106;
  assign n1684 = ~pi129 & ~n1683;
  assign n1685 = ~pi106 & ~n2674;
  assign n1686 = pi88 & pi106;
  assign n1687 = ~n1685 & ~n1686;
  assign n1688 = ~pi129 & ~n1687;
  assign n1689 = ~n2675 & n1684;
  assign n1690 = ~pi31 & ~pi109;
  assign n1691 = ~pi30 & pi109;
  assign n1692 = pi30 & pi109;
  assign n1693 = pi31 & ~pi109;
  assign n1694 = ~n1692 & ~n1693;
  assign n1695 = ~n1690 & ~n1691;
  assign n1696 = ~pi106 & ~n1693;
  assign n1697 = ~n1692 & n1696;
  assign n1698 = ~pi106 & n2677;
  assign n1699 = ~pi89 & pi106;
  assign n1700 = ~pi129 & ~n1699;
  assign n1701 = pi89 & pi106;
  assign n1702 = ~pi106 & ~n2677;
  assign n1703 = ~n1701 & ~n1702;
  assign n1704 = ~pi129 & ~n1703;
  assign n1705 = ~n2678 & n1700;
  assign n1706 = ~pi32 & ~pi109;
  assign n1707 = ~pi31 & pi109;
  assign n1708 = pi31 & pi109;
  assign n1709 = pi32 & ~pi109;
  assign n1710 = ~n1708 & ~n1709;
  assign n1711 = ~n1706 & ~n1707;
  assign n1712 = ~pi106 & ~n1709;
  assign n1713 = ~n1708 & n1712;
  assign n1714 = ~pi106 & n2680;
  assign n1715 = ~pi99 & pi106;
  assign n1716 = ~pi129 & ~n1715;
  assign n1717 = pi99 & pi106;
  assign n1718 = ~pi106 & ~n2680;
  assign n1719 = ~n1717 & ~n1718;
  assign n1720 = ~pi129 & ~n1719;
  assign n1721 = ~n2681 & n1716;
  assign n1722 = ~pi33 & ~pi109;
  assign n1723 = ~pi32 & pi109;
  assign n1724 = pi32 & pi109;
  assign n1725 = pi33 & ~pi109;
  assign n1726 = ~n1724 & ~n1725;
  assign n1727 = ~n1722 & ~n1723;
  assign n1728 = ~pi106 & ~n1725;
  assign n1729 = ~n1724 & n1728;
  assign n1730 = ~pi106 & n2683;
  assign n1731 = ~pi90 & pi106;
  assign n1732 = ~pi129 & ~n1731;
  assign n1733 = pi90 & pi106;
  assign n1734 = ~pi106 & ~n2683;
  assign n1735 = ~n1733 & ~n1734;
  assign n1736 = ~pi129 & ~n1735;
  assign n1737 = ~n2684 & n1732;
  assign n1738 = ~pi34 & ~pi109;
  assign n1739 = ~pi33 & pi109;
  assign n1740 = pi33 & pi109;
  assign n1741 = pi34 & ~pi109;
  assign n1742 = ~n1740 & ~n1741;
  assign n1743 = ~n1738 & ~n1739;
  assign n1744 = ~pi106 & ~n1741;
  assign n1745 = ~n1740 & n1744;
  assign n1746 = ~pi106 & n2686;
  assign n1747 = ~pi91 & pi106;
  assign n1748 = ~pi129 & ~n1747;
  assign n1749 = pi91 & pi106;
  assign n1750 = ~pi106 & ~n2686;
  assign n1751 = ~n1749 & ~n1750;
  assign n1752 = ~pi129 & ~n1751;
  assign n1753 = ~n2687 & n1748;
  assign n1754 = ~pi35 & ~pi109;
  assign n1755 = ~pi34 & pi109;
  assign n1756 = pi34 & pi109;
  assign n1757 = pi35 & ~pi109;
  assign n1758 = ~n1756 & ~n1757;
  assign n1759 = ~n1754 & ~n1755;
  assign n1760 = ~pi106 & ~n1757;
  assign n1761 = ~n1756 & n1760;
  assign n1762 = ~pi106 & n2689;
  assign n1763 = ~pi92 & pi106;
  assign n1764 = ~pi129 & ~n1763;
  assign n1765 = pi92 & pi106;
  assign n1766 = ~pi106 & ~n2689;
  assign n1767 = ~n1765 & ~n1766;
  assign n1768 = ~pi129 & ~n1767;
  assign n1769 = ~n2690 & n1764;
  assign n1770 = ~pi36 & ~pi109;
  assign n1771 = ~pi35 & pi109;
  assign n1772 = pi35 & pi109;
  assign n1773 = pi36 & ~pi109;
  assign n1774 = ~n1772 & ~n1773;
  assign n1775 = ~n1770 & ~n1771;
  assign n1776 = ~pi106 & ~n1773;
  assign n1777 = ~n1772 & n1776;
  assign n1778 = ~pi106 & n2692;
  assign n1779 = ~pi98 & pi106;
  assign n1780 = ~pi129 & ~n1779;
  assign n1781 = pi98 & pi106;
  assign n1782 = ~pi106 & ~n2692;
  assign n1783 = ~n1781 & ~n1782;
  assign n1784 = ~pi129 & ~n1783;
  assign n1785 = ~n2693 & n1780;
  assign n1786 = ~pi37 & ~pi109;
  assign n1787 = ~pi36 & pi109;
  assign n1788 = pi36 & pi109;
  assign n1789 = pi37 & ~pi109;
  assign n1790 = ~n1788 & ~n1789;
  assign n1791 = ~n1786 & ~n1787;
  assign n1792 = ~pi106 & ~n1789;
  assign n1793 = ~n1788 & n1792;
  assign n1794 = ~pi106 & n2695;
  assign n1795 = ~pi93 & pi106;
  assign n1796 = ~pi129 & ~n1795;
  assign n1797 = pi93 & pi106;
  assign n1798 = ~pi106 & ~n2695;
  assign n1799 = ~n1797 & ~n1798;
  assign n1800 = ~pi129 & ~n1799;
  assign n1801 = ~n2696 & n1796;
  assign n1802 = pi109 & n1049;
  assign n1803 = pi39 & ~n1802;
  assign n1804 = ~pi51 & pi109;
  assign n1805 = n1048 & n1804;
  assign n1806 = ~pi106 & ~n1805;
  assign n1807 = ~n1803 & n1806;
  assign po54 = ~pi129 & ~n1807;
  assign n1809 = pi52 & ~n1804;
  assign n1810 = ~pi106 & ~n1802;
  assign n1811 = ~n1809 & n1810;
  assign po67 = ~pi129 & ~n1811;
  assign n1813 = ~pi23 & pi55;
  assign n1814 = pi61 & ~pi129;
  assign n1815 = ~pi129 & ~n1813;
  assign n1816 = pi61 & n1815;
  assign n1817 = ~n1813 & n1814;
  assign n1818 = pi51 & ~pi109;
  assign n1819 = ~pi106 & ~n1804;
  assign n1820 = ~n1804 & ~n1818;
  assign n1821 = ~pi106 & n1820;
  assign n1822 = ~n1818 & n1819;
  assign po66 = ~pi129 & ~n2699;
  assign n1824 = ~pi123 & ~pi129;
  assign n1825 = pi114 & ~pi122;
  assign po70 = n1824 & n1825;
  assign n1827 = ~pi117 & ~pi122;
  assign n1828 = pi60 & ~n1827;
  assign n1829 = pi123 & n1827;
  assign n1830 = ~n1828 & ~n1829;
  assign n1831 = ~pi114 & ~pi122;
  assign n1832 = pi123 & ~pi129;
  assign n1833 = ~pi114 & pi123;
  assign n1834 = ~pi122 & n1833;
  assign n1835 = ~pi129 & n1834;
  assign n1836 = n1831 & n1832;
  assign n1837 = ~pi26 & n1199;
  assign n1838 = n1188 & n2666;
  assign n1839 = ~pi27 & n1838;
  assign n1840 = n2666 & n1837;
  assign n1841 = ~n1037 & ~n2701;
  assign n1842 = ~pi129 & ~n1841;
  assign n1843 = ~pi3 & n1842;
  assign n1844 = n448 & ~n1841;
  assign n1845 = pi58 & ~pi116;
  assign n1846 = n1109 & n1845;
  assign n1847 = ~pi58 & ~n2590;
  assign n1848 = pi116 & ~n2590;
  assign n1849 = ~pi58 & n1848;
  assign n1850 = n2586 & n1849;
  assign n1851 = n1052 & n1847;
  assign n1852 = ~n1846 & ~n2703;
  assign n1853 = ~pi53 & ~pi85;
  assign n1854 = n448 & n1853;
  assign n1855 = ~pi129 & ~n1852;
  assign n1856 = ~pi3 & n1855;
  assign n1857 = ~pi53 & n1856;
  assign n1858 = ~pi85 & n1857;
  assign n1859 = ~n1852 & n1854;
  assign n1860 = ~pi26 & pi58;
  assign n1861 = pi26 & ~pi58;
  assign n1862 = pi116 & n1861;
  assign n1863 = ~pi58 & n1071;
  assign n1864 = ~n1860 & ~n2705;
  assign n1865 = pi94 & ~n1864;
  assign n1866 = pi37 & ~pi116;
  assign n1867 = ~n1860 & ~n1866;
  assign n1868 = ~n1845 & ~n1867;
  assign n1869 = ~n1865 & ~n1868;
  assign n1870 = ~pi53 & ~n1869;
  assign n1871 = ~pi26 & pi37;
  assign n1872 = ~pi58 & n1871;
  assign n1873 = ~n1870 & ~n1872;
  assign n1874 = ~pi85 & ~n1873;
  assign n1875 = n1085 & n1871;
  assign n1876 = ~n1874 & ~n1875;
  assign n1877 = ~pi27 & ~n1876;
  assign n1878 = n1254 & n1871;
  assign n1879 = ~n1877 & ~n1878;
  assign n1880 = ~pi129 & ~n1879;
  assign n1881 = ~pi3 & n1880;
  assign n1882 = n448 & ~n1879;
  assign n1883 = ~pi116 & n1160;
  assign n1884 = pi85 & ~n1159;
  assign n1885 = pi26 & pi53;
  assign n1886 = ~pi58 & ~n1885;
  assign n1887 = ~pi85 & ~n1885;
  assign n1888 = ~n1159 & ~n1887;
  assign n1889 = ~pi58 & ~n1888;
  assign n1890 = ~n1884 & n1886;
  assign n1891 = ~n1883 & ~n2707;
  assign n1892 = pi57 & ~n1891;
  assign n1893 = pi60 & n1582;
  assign n1894 = n1160 & n1893;
  assign n1895 = ~n1892 & ~n1894;
  assign n1896 = ~pi27 & ~n1895;
  assign n1897 = pi57 & ~pi58;
  assign n1898 = n1160 & n1897;
  assign n1899 = ~n1896 & ~n1898;
  assign n1900 = ~pi129 & ~n1899;
  assign n1901 = ~pi3 & n1900;
  assign n1902 = n448 & ~n1899;
  assign n1903 = pi136 & ~pi138;
  assign n1904 = pi31 & n1903;
  assign n1905 = pi115 & pi138;
  assign n1906 = ~pi87 & ~pi138;
  assign n1907 = ~pi136 & ~n1906;
  assign n1908 = ~pi115 & pi138;
  assign n1909 = pi87 & ~pi138;
  assign n1910 = ~n1908 & ~n1909;
  assign n1911 = ~pi136 & ~n1910;
  assign n1912 = ~n1905 & n1907;
  assign n1913 = ~n1904 & ~n2709;
  assign n1914 = pi137 & ~n1913;
  assign n1915 = pi62 & ~pi138;
  assign n1916 = ~pi89 & pi138;
  assign n1917 = pi136 & ~n1916;
  assign n1918 = pi89 & pi138;
  assign n1919 = ~pi62 & ~pi138;
  assign n1920 = ~n1918 & ~n1919;
  assign n1921 = pi136 & ~n1920;
  assign n1922 = ~n1915 & n1917;
  assign n1923 = pi72 & ~pi138;
  assign n1924 = ~pi119 & pi138;
  assign n1925 = ~pi136 & ~n1924;
  assign n1926 = pi119 & pi138;
  assign n1927 = ~pi72 & ~pi138;
  assign n1928 = ~n1926 & ~n1927;
  assign n1929 = ~pi136 & ~n1928;
  assign n1930 = ~n1923 & n1925;
  assign n1931 = ~n2710 & ~n2711;
  assign n1932 = ~pi137 & ~n1931;
  assign n1933 = ~n1914 & ~n1932;
  assign n1934 = ~pi142 & n2670;
  assign n1935 = ~pi94 & ~n2670;
  assign n1936 = ~pi129 & ~n1935;
  assign n1937 = pi94 & ~n2670;
  assign n1938 = pi142 & n2670;
  assign n1939 = ~n1937 & ~n1938;
  assign n1940 = ~pi129 & ~n1939;
  assign n1941 = ~n1934 & n1936;
  assign n1942 = pi37 & n1903;
  assign n1943 = ~pi96 & pi138;
  assign n1944 = ~pi82 & ~pi138;
  assign n1945 = ~pi136 & ~n1944;
  assign n1946 = pi96 & pi138;
  assign n1947 = pi82 & ~pi138;
  assign n1948 = ~n1946 & ~n1947;
  assign n1949 = ~pi136 & ~n1948;
  assign n1950 = ~n1943 & n1945;
  assign n1951 = ~n1942 & ~n2713;
  assign n1952 = pi137 & ~n1951;
  assign n1953 = pi65 & ~pi138;
  assign n1954 = ~pi93 & pi138;
  assign n1955 = pi136 & ~n1954;
  assign n1956 = ~pi65 & ~pi138;
  assign n1957 = pi93 & pi138;
  assign n1958 = ~n1956 & ~n1957;
  assign n1959 = pi136 & ~n1958;
  assign n1960 = ~n1953 & n1955;
  assign n1961 = pi77 & ~pi138;
  assign n1962 = ~pi124 & pi138;
  assign n1963 = ~pi136 & ~n1962;
  assign n1964 = pi124 & pi138;
  assign n1965 = ~pi77 & ~pi138;
  assign n1966 = ~n1964 & ~n1965;
  assign n1967 = ~pi136 & ~n1966;
  assign n1968 = ~n1961 & n1963;
  assign n1969 = ~n2714 & ~n2715;
  assign n1970 = ~pi137 & ~n1969;
  assign n1971 = ~n1952 & ~n1970;
  assign n1972 = pi35 & n1903;
  assign n1973 = ~pi100 & pi138;
  assign n1974 = ~pi80 & ~pi138;
  assign n1975 = ~pi136 & ~n1974;
  assign n1976 = pi80 & ~pi138;
  assign n1977 = pi100 & pi138;
  assign n1978 = ~n1976 & ~n1977;
  assign n1979 = ~pi136 & ~n1978;
  assign n1980 = ~n1973 & n1975;
  assign n1981 = ~n1972 & ~n2716;
  assign n1982 = pi137 & ~n1981;
  assign n1983 = pi70 & ~pi138;
  assign n1984 = ~pi92 & pi138;
  assign n1985 = pi136 & ~n1984;
  assign n1986 = pi92 & pi138;
  assign n1987 = ~pi70 & ~pi138;
  assign n1988 = ~n1986 & ~n1987;
  assign n1989 = pi136 & ~n1988;
  assign n1990 = ~n1983 & n1985;
  assign n1991 = pi75 & ~pi138;
  assign n1992 = ~pi125 & pi138;
  assign n1993 = ~pi136 & ~n1992;
  assign n1994 = pi125 & pi138;
  assign n1995 = ~pi75 & ~pi138;
  assign n1996 = ~n1994 & ~n1995;
  assign n1997 = ~pi136 & ~n1996;
  assign n1998 = ~n1991 & n1993;
  assign n1999 = ~n2717 & ~n2718;
  assign n2000 = ~pi137 & ~n1999;
  assign n2001 = ~n1982 & ~n2000;
  assign n2002 = pi36 & n1903;
  assign n2003 = ~pi97 & pi138;
  assign n2004 = ~pi81 & ~pi138;
  assign n2005 = ~pi136 & ~n2004;
  assign n2006 = pi81 & ~pi138;
  assign n2007 = pi97 & pi138;
  assign n2008 = ~n2006 & ~n2007;
  assign n2009 = ~pi136 & ~n2008;
  assign n2010 = ~n2003 & n2005;
  assign n2011 = ~n2002 & ~n2719;
  assign n2012 = pi137 & ~n2011;
  assign n2013 = pi71 & ~pi138;
  assign n2014 = ~pi98 & pi138;
  assign n2015 = pi136 & ~n2014;
  assign n2016 = pi98 & pi138;
  assign n2017 = ~pi71 & ~pi138;
  assign n2018 = ~n2016 & ~n2017;
  assign n2019 = pi136 & ~n2018;
  assign n2020 = ~n2013 & n2015;
  assign n2021 = pi76 & ~pi138;
  assign n2022 = ~pi23 & pi138;
  assign n2023 = ~pi136 & ~n2022;
  assign n2024 = ~pi76 & ~pi138;
  assign n2025 = pi23 & pi138;
  assign n2026 = ~n2024 & ~n2025;
  assign n2027 = ~pi136 & ~n2026;
  assign n2028 = ~n2021 & n2023;
  assign n2029 = ~n2720 & ~n2721;
  assign n2030 = ~pi137 & ~n2029;
  assign n2031 = ~n2012 & ~n2030;
  assign n2032 = pi30 & n1903;
  assign n2033 = ~pi111 & pi138;
  assign n2034 = ~pi86 & ~pi138;
  assign n2035 = ~pi136 & ~n2034;
  assign n2036 = pi86 & ~pi138;
  assign n2037 = pi111 & pi138;
  assign n2038 = ~n2036 & ~n2037;
  assign n2039 = ~pi136 & ~n2038;
  assign n2040 = ~n2033 & n2035;
  assign n2041 = ~n2032 & ~n2722;
  assign n2042 = pi137 & ~n2041;
  assign n2043 = pi64 & ~pi138;
  assign n2044 = ~pi88 & pi138;
  assign n2045 = pi136 & ~n2044;
  assign n2046 = pi88 & pi138;
  assign n2047 = ~pi64 & ~pi138;
  assign n2048 = ~n2046 & ~n2047;
  assign n2049 = pi136 & ~n2048;
  assign n2050 = ~n2043 & n2045;
  assign n2051 = pi67 & ~pi138;
  assign n2052 = ~pi120 & pi138;
  assign n2053 = ~pi136 & ~n2052;
  assign n2054 = pi120 & pi138;
  assign n2055 = ~pi67 & ~pi138;
  assign n2056 = ~n2054 & ~n2055;
  assign n2057 = ~pi136 & ~n2056;
  assign n2058 = ~n2051 & n2053;
  assign n2059 = ~n2723 & ~n2724;
  assign n2060 = ~pi137 & ~n2059;
  assign n2061 = ~n2042 & ~n2060;
  assign n2062 = ~pi139 & n2669;
  assign n2063 = ~pi129 & n2668;
  assign n2064 = ~pi111 & ~n2669;
  assign n2065 = n2063 & ~n2064;
  assign n2066 = pi111 & ~n2669;
  assign n2067 = ~pi136 & pi139;
  assign n2068 = pi82 & n1620;
  assign n2069 = n2067 & n2068;
  assign n2070 = ~n2066 & ~n2069;
  assign n2071 = n2668 & ~n2070;
  assign n2072 = ~pi129 & n2071;
  assign n2073 = ~n2062 & n2065;
  assign n2074 = pi112 & ~n2669;
  assign n2075 = ~pi141 & n2669;
  assign n2076 = n2063 & ~n2075;
  assign n2077 = ~pi136 & pi141;
  assign n2078 = n2068 & n2077;
  assign n2079 = ~pi112 & ~n2669;
  assign n2080 = ~n2078 & ~n2079;
  assign n2081 = n2668 & ~n2080;
  assign n2082 = ~pi129 & n2081;
  assign n2083 = ~n2074 & n2076;
  assign n2084 = pi115 & ~n2669;
  assign n2085 = ~pi140 & n2669;
  assign n2086 = n2063 & ~n2085;
  assign n2087 = ~pi136 & pi140;
  assign n2088 = n2068 & n2087;
  assign n2089 = ~pi115 & ~n2669;
  assign n2090 = ~n2088 & ~n2089;
  assign n2091 = n2668 & ~n2090;
  assign n2092 = ~pi129 & n2091;
  assign n2093 = ~n2084 & n2086;
  assign n2094 = ~pi137 & ~pi138;
  assign n2095 = pi136 & n2094;
  assign n2096 = ~pi138 & n2668;
  assign n2097 = n1649 & n2096;
  assign n2098 = n2668 & n2095;
  assign n2099 = pi140 & n2728;
  assign n2100 = ~pi62 & ~n2728;
  assign n2101 = ~pi129 & ~n2100;
  assign n2102 = pi62 & ~n2728;
  assign n2103 = ~pi140 & n1649;
  assign n2104 = n2096 & n2103;
  assign n2105 = ~n2102 & ~n2104;
  assign n2106 = ~pi129 & ~n2105;
  assign n2107 = ~n2099 & n2101;
  assign n2108 = pi142 & n2728;
  assign n2109 = ~pi63 & ~n2728;
  assign n2110 = ~pi129 & ~n2109;
  assign n2111 = pi63 & ~n2728;
  assign n2112 = ~pi142 & n1649;
  assign n2113 = n2096 & n2112;
  assign n2114 = ~n2111 & ~n2113;
  assign n2115 = ~pi129 & ~n2114;
  assign n2116 = ~n2108 & n2110;
  assign n2117 = pi139 & n2728;
  assign n2118 = ~pi64 & ~n2728;
  assign n2119 = ~pi129 & ~n2118;
  assign n2120 = pi64 & ~n2728;
  assign n2121 = ~pi139 & n1649;
  assign n2122 = n2096 & n2121;
  assign n2123 = ~n2120 & ~n2122;
  assign n2124 = ~pi129 & ~n2123;
  assign n2125 = ~n2117 & n2119;
  assign n2126 = pi146 & n2728;
  assign n2127 = ~pi65 & ~n2728;
  assign n2128 = ~pi129 & ~n2127;
  assign n2129 = pi65 & ~n2728;
  assign n2130 = ~pi146 & n1649;
  assign n2131 = n2096 & n2130;
  assign n2132 = ~n2129 & ~n2131;
  assign n2133 = ~pi129 & ~n2132;
  assign n2134 = ~n2126 & n2128;
  assign n2135 = n1614 & n2096;
  assign n2136 = pi143 & n2135;
  assign n2137 = ~pi66 & ~n2135;
  assign n2138 = ~pi129 & ~n2137;
  assign n2139 = pi66 & ~n2135;
  assign n2140 = ~pi143 & n2135;
  assign n2141 = ~n2139 & ~n2140;
  assign n2142 = ~pi129 & ~n2141;
  assign n2143 = ~n2136 & n2138;
  assign n2144 = pi139 & n2135;
  assign n2145 = ~pi67 & ~n2135;
  assign n2146 = ~pi129 & ~n2145;
  assign n2147 = pi67 & ~n2135;
  assign n2148 = ~pi139 & n2135;
  assign n2149 = ~n2147 & ~n2148;
  assign n2150 = ~pi129 & ~n2149;
  assign n2151 = ~n2144 & n2146;
  assign n2152 = pi141 & n2728;
  assign n2153 = ~pi68 & ~n2728;
  assign n2154 = ~pi129 & ~n2153;
  assign n2155 = pi68 & ~n2728;
  assign n2156 = ~pi141 & n1649;
  assign n2157 = n2096 & n2156;
  assign n2158 = ~n2155 & ~n2157;
  assign n2159 = ~pi129 & ~n2158;
  assign n2160 = ~n2152 & n2154;
  assign n2161 = pi143 & n2728;
  assign n2162 = ~pi69 & ~n2728;
  assign n2163 = ~pi129 & ~n2162;
  assign n2164 = pi69 & ~n2728;
  assign n2165 = ~pi143 & n1649;
  assign n2166 = n2096 & n2165;
  assign n2167 = ~n2164 & ~n2166;
  assign n2168 = ~pi129 & ~n2167;
  assign n2169 = ~n2161 & n2163;
  assign n2170 = pi144 & n2728;
  assign n2171 = ~pi70 & ~n2728;
  assign n2172 = ~pi129 & ~n2171;
  assign n2173 = pi70 & ~n2728;
  assign n2174 = ~pi144 & n1649;
  assign n2175 = n2096 & n2174;
  assign n2176 = ~n2173 & ~n2175;
  assign n2177 = ~pi129 & ~n2176;
  assign n2178 = ~n2170 & n2172;
  assign n2179 = pi145 & n2728;
  assign n2180 = ~pi71 & ~n2728;
  assign n2181 = ~pi129 & ~n2180;
  assign n2182 = pi71 & ~n2728;
  assign n2183 = ~pi145 & n1649;
  assign n2184 = n2096 & n2183;
  assign n2185 = ~n2182 & ~n2184;
  assign n2186 = ~pi129 & ~n2185;
  assign n2187 = ~n2179 & n2181;
  assign n2188 = pi140 & n2135;
  assign n2189 = ~pi72 & ~n2135;
  assign n2190 = ~pi129 & ~n2189;
  assign n2191 = pi72 & ~n2135;
  assign n2192 = ~pi140 & n2135;
  assign n2193 = ~n2191 & ~n2192;
  assign n2194 = ~pi129 & ~n2193;
  assign n2195 = ~n2188 & n2190;
  assign n2196 = pi141 & n2135;
  assign n2197 = ~pi73 & ~n2135;
  assign n2198 = ~pi129 & ~n2197;
  assign n2199 = pi73 & ~n2135;
  assign n2200 = ~pi141 & n2135;
  assign n2201 = ~n2199 & ~n2200;
  assign n2202 = ~pi129 & ~n2201;
  assign n2203 = ~n2196 & n2198;
  assign n2204 = pi142 & n2135;
  assign n2205 = ~pi74 & ~n2135;
  assign n2206 = ~pi129 & ~n2205;
  assign n2207 = pi74 & ~n2135;
  assign n2208 = ~pi142 & n2135;
  assign n2209 = ~n2207 & ~n2208;
  assign n2210 = ~pi129 & ~n2209;
  assign n2211 = ~n2204 & n2206;
  assign n2212 = pi144 & n2135;
  assign n2213 = ~pi75 & ~n2135;
  assign n2214 = ~pi129 & ~n2213;
  assign n2215 = pi75 & ~n2135;
  assign n2216 = ~pi144 & n2135;
  assign n2217 = ~n2215 & ~n2216;
  assign n2218 = ~pi129 & ~n2217;
  assign n2219 = ~n2212 & n2214;
  assign n2220 = pi145 & n2135;
  assign n2221 = ~pi76 & ~n2135;
  assign n2222 = ~pi129 & ~n2221;
  assign n2223 = pi76 & ~n2135;
  assign n2224 = ~pi145 & n2135;
  assign n2225 = ~n2223 & ~n2224;
  assign n2226 = ~pi129 & ~n2225;
  assign n2227 = ~n2220 & n2222;
  assign n2228 = pi146 & n2135;
  assign n2229 = ~pi77 & ~n2135;
  assign n2230 = ~pi129 & ~n2229;
  assign n2231 = pi77 & ~n2135;
  assign n2232 = ~pi146 & n2135;
  assign n2233 = ~n2231 & ~n2232;
  assign n2234 = ~pi129 & ~n2233;
  assign n2235 = ~n2228 & n2230;
  assign n2236 = n1651 & n2096;
  assign n2237 = ~pi142 & n2236;
  assign n2238 = ~pi78 & ~n2236;
  assign n2239 = ~pi129 & ~n2238;
  assign n2240 = pi78 & ~n2236;
  assign n2241 = pi142 & n2236;
  assign n2242 = ~n2240 & ~n2241;
  assign n2243 = ~pi129 & ~n2242;
  assign n2244 = ~n2237 & n2239;
  assign n2245 = ~pi143 & n2236;
  assign n2246 = ~pi79 & ~n2236;
  assign n2247 = ~pi129 & ~n2246;
  assign n2248 = pi79 & ~n2236;
  assign n2249 = pi143 & n2236;
  assign n2250 = ~n2248 & ~n2249;
  assign n2251 = ~pi129 & ~n2250;
  assign n2252 = ~n2245 & n2247;
  assign n2253 = ~pi144 & n2236;
  assign n2254 = ~pi80 & ~n2236;
  assign n2255 = ~pi129 & ~n2254;
  assign n2256 = pi80 & ~n2236;
  assign n2257 = pi144 & n2236;
  assign n2258 = ~n2256 & ~n2257;
  assign n2259 = ~pi129 & ~n2258;
  assign n2260 = ~n2253 & n2255;
  assign n2261 = ~pi145 & n2236;
  assign n2262 = ~pi81 & ~n2236;
  assign n2263 = ~pi129 & ~n2262;
  assign n2264 = pi81 & ~n2236;
  assign n2265 = pi145 & n2236;
  assign n2266 = ~n2264 & ~n2265;
  assign n2267 = ~pi129 & ~n2266;
  assign n2268 = ~n2261 & n2263;
  assign n2269 = ~pi146 & n2236;
  assign n2270 = ~pi82 & ~n2236;
  assign n2271 = ~pi129 & ~n2270;
  assign n2272 = pi82 & ~n2236;
  assign n2273 = pi146 & n2236;
  assign n2274 = ~n2272 & ~n2273;
  assign n2275 = ~pi129 & ~n2274;
  assign n2276 = ~n2269 & n2271;
  assign n2277 = ~pi141 & n2236;
  assign n2278 = ~pi84 & ~n2236;
  assign n2279 = ~pi129 & ~n2278;
  assign n2280 = pi84 & ~n2236;
  assign n2281 = pi141 & n2236;
  assign n2282 = ~n2280 & ~n2281;
  assign n2283 = ~pi129 & ~n2282;
  assign n2284 = ~n2277 & n2279;
  assign n2285 = ~pi139 & n2236;
  assign n2286 = ~pi86 & ~n2236;
  assign n2287 = ~pi129 & ~n2286;
  assign n2288 = pi86 & ~n2236;
  assign n2289 = pi139 & n2236;
  assign n2290 = ~n2288 & ~n2289;
  assign n2291 = ~pi129 & ~n2290;
  assign n2292 = ~n2285 & n2287;
  assign n2293 = ~pi140 & n2236;
  assign n2294 = ~pi87 & ~n2236;
  assign n2295 = ~pi129 & ~n2294;
  assign n2296 = pi87 & ~n2236;
  assign n2297 = pi140 & n2236;
  assign n2298 = ~n2296 & ~n2297;
  assign n2299 = ~pi129 & ~n2298;
  assign n2300 = ~n2293 & n2295;
  assign n2301 = pi137 & n1903;
  assign n2302 = pi136 & pi137;
  assign n2303 = n2096 & n2302;
  assign n2304 = n2668 & n2301;
  assign n2305 = ~pi139 & n2753;
  assign n2306 = ~pi88 & ~n2753;
  assign n2307 = ~pi129 & ~n2306;
  assign n2308 = pi88 & ~n2753;
  assign n2309 = pi139 & n2753;
  assign n2310 = ~n2308 & ~n2309;
  assign n2311 = ~pi129 & ~n2310;
  assign n2312 = ~n2305 & n2307;
  assign n2313 = ~pi140 & n2753;
  assign n2314 = ~pi89 & ~n2753;
  assign n2315 = ~pi129 & ~n2314;
  assign n2316 = pi89 & ~n2753;
  assign n2317 = pi140 & n2753;
  assign n2318 = ~n2316 & ~n2317;
  assign n2319 = ~pi129 & ~n2318;
  assign n2320 = ~n2313 & n2315;
  assign n2321 = ~pi142 & n2753;
  assign n2322 = ~pi90 & ~n2753;
  assign n2323 = ~pi129 & ~n2322;
  assign n2324 = pi90 & ~n2753;
  assign n2325 = pi142 & n2753;
  assign n2326 = ~n2324 & ~n2325;
  assign n2327 = ~pi129 & ~n2326;
  assign n2328 = ~n2321 & n2323;
  assign n2329 = ~pi143 & n2753;
  assign n2330 = ~pi91 & ~n2753;
  assign n2331 = ~pi129 & ~n2330;
  assign n2332 = pi91 & ~n2753;
  assign n2333 = pi143 & n2753;
  assign n2334 = ~n2332 & ~n2333;
  assign n2335 = ~pi129 & ~n2334;
  assign n2336 = ~n2329 & n2331;
  assign n2337 = ~pi144 & n2753;
  assign n2338 = ~pi92 & ~n2753;
  assign n2339 = ~pi129 & ~n2338;
  assign n2340 = pi92 & ~n2753;
  assign n2341 = pi144 & n2753;
  assign n2342 = ~n2340 & ~n2341;
  assign n2343 = ~pi129 & ~n2342;
  assign n2344 = ~n2337 & n2339;
  assign n2345 = ~pi146 & n2753;
  assign n2346 = ~pi93 & ~n2753;
  assign n2347 = ~pi129 & ~n2346;
  assign n2348 = pi93 & ~n2753;
  assign n2349 = pi146 & n2753;
  assign n2350 = ~n2348 & ~n2349;
  assign n2351 = ~pi129 & ~n2350;
  assign n2352 = ~n2345 & n2347;
  assign n2353 = ~pi145 & n2753;
  assign n2354 = ~pi98 & ~n2753;
  assign n2355 = ~pi129 & ~n2354;
  assign n2356 = pi98 & ~n2753;
  assign n2357 = pi145 & n2753;
  assign n2358 = ~n2356 & ~n2357;
  assign n2359 = ~pi129 & ~n2358;
  assign n2360 = ~n2353 & n2355;
  assign n2361 = ~pi141 & n2753;
  assign n2362 = ~pi99 & ~n2753;
  assign n2363 = ~pi129 & ~n2362;
  assign n2364 = pi99 & ~n2753;
  assign n2365 = pi141 & n2753;
  assign n2366 = ~n2364 & ~n2365;
  assign n2367 = ~pi129 & ~n2366;
  assign n2368 = ~n2361 & n2363;
  assign n2369 = pi91 & n1649;
  assign n2370 = pi95 & n1651;
  assign n2371 = ~n2369 & ~n2370;
  assign n2372 = pi138 & ~n2371;
  assign n2373 = ~pi34 & pi136;
  assign n2374 = ~pi79 & ~pi136;
  assign n2375 = pi137 & ~n2374;
  assign n2376 = pi79 & ~pi136;
  assign n2377 = pi34 & pi136;
  assign n2378 = ~n2376 & ~n2377;
  assign n2379 = pi137 & ~n2378;
  assign n2380 = ~n2373 & n2375;
  assign n2381 = pi69 & pi136;
  assign n2382 = pi66 & ~pi136;
  assign n2383 = ~pi137 & ~n2382;
  assign n2384 = ~pi69 & pi136;
  assign n2385 = ~pi66 & ~pi136;
  assign n2386 = ~n2384 & ~n2385;
  assign n2387 = ~pi137 & ~n2386;
  assign n2388 = ~n2381 & n2383;
  assign n2389 = ~n2762 & ~n2763;
  assign n2390 = ~pi138 & ~n2389;
  assign n2391 = ~n2372 & ~n2390;
  assign n2392 = pi90 & n1649;
  assign n2393 = pi94 & n1651;
  assign n2394 = ~n2392 & ~n2393;
  assign n2395 = pi138 & ~n2394;
  assign n2396 = ~pi33 & pi136;
  assign n2397 = ~pi78 & ~pi136;
  assign n2398 = pi137 & ~n2397;
  assign n2399 = pi78 & ~pi136;
  assign n2400 = pi33 & pi136;
  assign n2401 = ~n2399 & ~n2400;
  assign n2402 = pi137 & ~n2401;
  assign n2403 = ~n2396 & n2398;
  assign n2404 = pi63 & pi136;
  assign n2405 = pi74 & ~pi136;
  assign n2406 = ~pi137 & ~n2405;
  assign n2407 = ~pi63 & pi136;
  assign n2408 = ~pi74 & ~pi136;
  assign n2409 = ~n2407 & ~n2408;
  assign n2410 = ~pi137 & ~n2409;
  assign n2411 = ~n2404 & n2406;
  assign n2412 = ~n2764 & ~n2765;
  assign n2413 = ~pi138 & ~n2412;
  assign n2414 = ~n2395 & ~n2413;
  assign n2415 = ~pi26 & n2586;
  assign n2416 = pi116 & n448;
  assign n2417 = ~n2590 & n2416;
  assign n2418 = ~n2586 & n1112;
  assign n2419 = ~n1111 & ~n2418;
  assign n2420 = ~pi129 & ~n2419;
  assign n2421 = ~pi3 & n2420;
  assign n2422 = pi116 & n2421;
  assign n2423 = ~n2415 & n2417;
  assign n2424 = ~pi4 & ~pi9;
  assign n2425 = ~pi4 & ~pi12;
  assign n2426 = ~pi7 & ~pi9;
  assign n2427 = n2425 & n2426;
  assign n2428 = n466 & n2424;
  assign n2429 = pi54 & n448;
  assign n2430 = ~pi129 & ~n2767;
  assign n2431 = ~pi3 & n2430;
  assign n2432 = pi54 & n2431;
  assign n2433 = ~n2767 & n2429;
  assign n2434 = pi122 & ~pi129;
  assign n2435 = ~pi54 & pi118;
  assign n2436 = pi54 & ~pi59;
  assign n2437 = n2515 & n2436;
  assign n2438 = ~n2435 & ~n2437;
  assign po133 = ~pi129 & ~n2438;
  assign n2440 = ~pi97 & n1030;
  assign n2441 = ~n1031 & ~n2440;
  assign n2442 = ~pi129 & ~n2441;
  assign n2443 = ~pi3 & n2442;
  assign n2444 = pi116 & n2443;
  assign n2445 = n2416 & ~n2441;
  assign n2446 = ~pi11 & ~pi22;
  assign n2447 = pi54 & n2446;
  assign n2448 = ~pi54 & pi113;
  assign n2449 = n448 & ~n2448;
  assign n2450 = ~pi54 & ~pi113;
  assign n2451 = pi54 & ~n2446;
  assign n2452 = ~n2450 & ~n2451;
  assign n2453 = ~pi129 & ~n2452;
  assign n2454 = ~pi3 & n2453;
  assign n2455 = ~n2447 & n2449;
  assign n2456 = ~pi110 & ~pi120;
  assign n2457 = ~pi3 & n2456;
  assign n2458 = ~pi120 & n1626;
  assign n2459 = ~pi111 & ~pi129;
  assign n2460 = ~pi129 & ~n2771;
  assign n2461 = ~pi111 & n2460;
  assign n2462 = ~n2771 & n2459;
  assign n2463 = ~pi129 & ~pi134;
  assign n2464 = ~pi129 & ~pi135;
  assign n2465 = ~pi96 & pi125;
  assign n2466 = ~pi3 & ~n2465;
  assign po140 = ~pi129 & ~n2466;
  assign po134 = ~pi129 & ~n1062;
  assign n2469 = pi81 & pi120;
  assign po136 = ~pi129 & n2469;
  assign n2471 = ~pi126 & pi132;
  assign po141 = pi133 & n2471;
  assign po139 = pi57 & ~pi129;
  assign n2474 = n298 | n299;
  assign n2475 = n300 | n301;
  assign n2476 = n306 | n303 | n305;
  assign n2477 = n313 | n314;
  assign n2478 = n321 | n317 | n320;
  assign n2479 = n318 | n319;
  assign n2480 = n322 | n323 | n325 | n326;
  assign n2481 = n327 | n328;
  assign n2482 = n329 | n330;
  assign n2483 = n335 | n331 | n334;
  assign n2484 = n336 | n342 | n343 | n344;
  assign n2485 = n340 | n341;
  assign n2486 = n349 | n350;
  assign n2487 = n352 | n353;
  assign n2488 = n357 | n358;
  assign n2489 = n363 | n361 | n362;
  assign n2490 = n381 | n366 | n380;
  assign n2491 = n373 | n374;
  assign n2492 = n379 | n375 | n378;
  assign n2493 = n383 | ~n384;
  assign n2494 = n386 | n387;
  assign n2495 = n428 | n397 | n402 | n432 | n430 | n431;
  assign n2496 = n404 | n405;
  assign n2497 = n406 | n407;
  assign n2498 = n409 | n410 | n426 | n427;
  assign n2499 = n411 | n412;
  assign n2500 = n419 | n415 | n418;
  assign n2501 = n416 | n417;
  assign n2502 = n425 | n423 | n424;
  assign n2503 = n439 | n435 | n438 | n440 | n441;
  assign n2504 = n443 | n444;
  assign n2505 = n462 | n458 | n461;
  assign n2506 = n459 | n460;
  assign n2507 = n469 | n470;
  assign n2508 = n475 | n476;
  assign n2509 = n479 | n480;
  assign n2510 = n489 | n490;
  assign po20 = n493 | n494;
  assign n2512 = n501 | n498 | n500;
  assign n2513 = n510 | n511;
  assign po21 = n514 | n515;
  assign n2515 = n523 | n524;
  assign n2516 = n533 | n531 | n532;
  assign n2517 = n537 | n534 | n536;
  assign n2518 = n554 | n541 | n553;
  assign n2519 = n549 | n543 | n548;
  assign n2520 = n546 | n547;
  assign po28 = n557 | n558;
  assign n2522 = n565 | n562 | n564;
  assign n2523 = n573 | n574;
  assign n2524 = n577 | n578;
  assign n2525 = n604 | n596 | n603;
  assign po32 = n607 | n608;
  assign n2527 = n611 | n612;
  assign n2528 = n619 | n620;
  assign n2529 = n628 | n629;
  assign n2530 = n649 | n642 | n648;
  assign n2531 = n676 | n671 | n675;
  assign n2532 = n680 | n681;
  assign n2533 = n686 | n687;
  assign n2534 = n699 | n700;
  assign n2535 = n703 | n704;
  assign n2536 = n712 | n713;
  assign n2537 = n728 | n729;
  assign n2538 = n730 | n731;
  assign n2539 = n737 | ~n738;
  assign n2540 = n739 | n740;
  assign n2541 = n747 | n748;
  assign n2542 = n755 | n756;
  assign n2543 = n759 | n760;
  assign n2544 = n766 | n764 | n765;
  assign n2545 = n769 | n770;
  assign po19 = n777 | n778;
  assign n2547 = n784 | n785;
  assign n2548 = n793 | n794;
  assign po22 = n797 | n798;
  assign n2550 = n806 | n807;
  assign n2551 = n808 | n809;
  assign po23 = n812 | n813;
  assign n2553 = n830 | n826 | n829;
  assign po24 = n833 | n834;
  assign n2555 = n837 | n838;
  assign n2556 = n850 | n847 | n849;
  assign po25 = n853 | n854;
  assign n2558 = n860 | n861;
  assign n2559 = n866 | n867;
  assign po26 = n870 | n871;
  assign n2561 = n885 | n880 | n884;
  assign po27 = n888 | n889;
  assign n2563 = n901 | n902;
  assign po29 = n905 | n906;
  assign n2565 = n912 | n913;
  assign n2566 = n915 | n916;
  assign po31 = n920 | n921;
  assign n2568 = n927 | n928;
  assign n2569 = n930 | n931;
  assign po33 = n934 | n935;
  assign n2571 = n939 | n940;
  assign po34 = n943 | n944;
  assign n2573 = n952 | n953;
  assign n2574 = n956 | n957;
  assign n2575 = n972 | n966 | n971;
  assign po36 = n976 | n977;
  assign n2577 = n986 | n987;
  assign n2578 = n996 | n997;
  assign po37 = n1000 | n1001;
  assign n2580 = n1003 | n1004;
  assign n2581 = n1008 | n1009;
  assign n2582 = n1024 | n1020 | n1023;
  assign po39 = n1028 | n1029;
  assign n2584 = n1041 | n1042;
  assign n2585 = n1044 | n1045;
  assign n2586 = n1050 | n1051;
  assign n2587 = n1081 | n1082;
  assign n2588 = n1088 | n1089;
  assign po40 = n1104 | n1102 | n1103;
  assign n2590 = n1113 | ~n1114;
  assign n2591 = n1123 | n1124;
  assign n2592 = n1125 | n1126;
  assign n2593 = n1149 | n1150;
  assign n2594 = n1153 | n1154;
  assign n2595 = n1162 | n1163;
  assign po43 = n1166 | n1167;
  assign n2597 = n1173 | n1174;
  assign n2598 = n1181 | n1182;
  assign po42 = n1189 | n1190;
  assign n2600 = n1195 | n1196;
  assign po41 = n1203 | n1204;
  assign n2602 = n1209 | n1210;
  assign n2603 = n1213 | n1214;
  assign n2604 = n1220 | n1221;
  assign n2605 = n1226 | n1227;
  assign n2606 = n1234 | n1235;
  assign n2607 = n1241 | n1242;
  assign n2608 = n1247 | n1248;
  assign n2609 = n1256 | n1253 | n1255;
  assign po44 = n1260 | n1261;
  assign n2611 = n1263 | n1264;
  assign n2612 = n1269 | n1267 | n1268;
  assign n2613 = n1270 | n1271;
  assign n2614 = n1276 | n1277;
  assign n2615 = n1285 | n1281 | n1284;
  assign n2616 = n1282 | n1283;
  assign n2617 = n1289 | n1290;
  assign n2618 = n1294 | n1295;
  assign n2619 = n1310 | n1307 | n1309;
  assign n2620 = n1314 | n1315;
  assign n2621 = n1317 | n1318;
  assign n2622 = n1328 | n1329;
  assign n2623 = n1330 | n1331;
  assign n2624 = n1335 | n1336;
  assign n2625 = n1338 | n1339;
  assign po56 = n1344 | n1345;
  assign n2627 = n1347 | n1348;
  assign n2628 = n1361 | n1362;
  assign n2629 = n1366 | n1367;
  assign po57 = n1371 | n1372;
  assign n2631 = n1379 | n1380;
  assign n2632 = n1384 | n1385;
  assign n2633 = n1387 | n1388;
  assign n2634 = n1390 | n1391;
  assign n2635 = n1396 | n1397;
  assign n2636 = n1403 | ~n1404;
  assign n2637 = n1409 | n1410;
  assign n2638 = n1414 | n1415;
  assign n2639 = n1423 | n1424;
  assign n2640 = n1425 | n1426;
  assign po60 = n1430 | n1431;
  assign n2642 = n1441 | n1442;
  assign n2643 = n1445 | n1446;
  assign n2644 = n1454 | n1455;
  assign n2645 = n1469 | n1465 | n1468;
  assign po62 = n1473 | n1474;
  assign n2647 = n1477 | n1478;
  assign n2648 = n1482 | n1483;
  assign n2649 = n1499 | n1494 | n1498;
  assign po63 = n1503 | n1504;
  assign n2651 = n1509 | n1510;
  assign n2652 = n1512 | n1513;
  assign n2653 = n1517 | n1518;
  assign n2654 = n1522 | n1523;
  assign n2655 = n1532 | n1533;
  assign n2656 = n1537 | n1538;
  assign n2657 = n1541 | n1542;
  assign po65 = n1546 | n1547;
  assign n2659 = n1561 | n1562;
  assign n2660 = n1563 | n1564;
  assign n2661 = n1572 | n1573;
  assign po74 = n1579 | n1580;
  assign n2663 = n1584 | n1585;
  assign n2664 = n1590 | n1591;
  assign po68 = n1597 | n1598;
  assign n2666 = n1600 | n1601;
  assign po100 = n1608 | n1609;
  assign n2668 = n1612 | n1613;
  assign n2669 = n1622 | n1618 | n1621;
  assign n2670 = n1624 | n1625;
  assign n2671 = n1631 | ~n1632;
  assign n2672 = n1661 | n1662;
  assign n2673 = n1669 | n1670;
  assign n2674 = n1678 | ~n1679;
  assign n2675 = n1681 | n1682;
  assign po45 = n1688 | n1689;
  assign n2677 = n1694 | ~n1695;
  assign n2678 = n1697 | n1698;
  assign po46 = n1704 | n1705;
  assign n2680 = n1710 | ~n1711;
  assign n2681 = n1713 | n1714;
  assign po47 = n1720 | n1721;
  assign n2683 = n1726 | ~n1727;
  assign n2684 = n1729 | n1730;
  assign po48 = n1736 | n1737;
  assign n2686 = n1742 | ~n1743;
  assign n2687 = n1745 | n1746;
  assign po49 = n1752 | n1753;
  assign n2689 = n1758 | ~n1759;
  assign n2690 = n1761 | n1762;
  assign po50 = n1768 | n1769;
  assign n2692 = n1774 | ~n1775;
  assign n2693 = n1777 | n1778;
  assign po51 = n1784 | n1785;
  assign n2695 = n1790 | ~n1791;
  assign n2696 = n1793 | n1794;
  assign po52 = n1800 | n1801;
  assign po38 = n1816 | n1817;
  assign n2699 = n1821 | n1822;
  assign po76 = n1835 | n1836;
  assign n2701 = n1839 | n1840;
  assign po121 = n1843 | n1844;
  assign n2703 = n1850 | n1851;
  assign po73 = n1858 | n1859;
  assign n2705 = n1862 | n1863;
  assign po71 = n1881 | n1882;
  assign n2707 = n1889 | n1890;
  assign po72 = n1901 | n1902;
  assign n2709 = n1911 | n1912;
  assign n2710 = n1921 | n1922;
  assign n2711 = n1929 | n1930;
  assign po109 = n1940 | n1941;
  assign n2713 = n1949 | n1950;
  assign n2714 = n1959 | n1960;
  assign n2715 = n1967 | n1968;
  assign n2716 = n1979 | n1980;
  assign n2717 = n1989 | n1990;
  assign n2718 = n1997 | n1998;
  assign n2719 = n2009 | n2010;
  assign n2720 = n2019 | n2020;
  assign n2721 = n2027 | n2028;
  assign n2722 = n2039 | n2040;
  assign n2723 = n2049 | n2050;
  assign n2724 = n2057 | n2058;
  assign po126 = n2072 | n2073;
  assign po127 = n2082 | n2083;
  assign po130 = n2092 | n2093;
  assign n2728 = n2097 | n2098;
  assign n2729 = n2106 | n2107;
  assign n2730 = n2115 | n2116;
  assign n2731 = n2124 | n2125;
  assign n2732 = n2133 | n2134;
  assign n2733 = n2142 | n2143;
  assign n2734 = n2150 | n2151;
  assign n2735 = n2159 | n2160;
  assign n2736 = n2168 | n2169;
  assign n2737 = n2177 | n2178;
  assign n2738 = n2186 | n2187;
  assign n2739 = n2194 | n2195;
  assign n2740 = n2202 | n2203;
  assign n2741 = n2210 | n2211;
  assign n2742 = n2218 | n2219;
  assign n2743 = n2226 | n2227;
  assign n2744 = n2234 | n2235;
  assign po93 = n2243 | n2244;
  assign po94 = n2251 | n2252;
  assign po95 = n2259 | n2260;
  assign po96 = n2267 | n2268;
  assign po97 = n2275 | n2276;
  assign po99 = n2283 | n2284;
  assign po101 = n2291 | n2292;
  assign po102 = n2299 | n2300;
  assign n2753 = n2303 | n2304;
  assign po103 = n2311 | n2312;
  assign po104 = n2319 | n2320;
  assign po105 = n2327 | n2328;
  assign po106 = n2335 | n2336;
  assign po107 = n2343 | n2344;
  assign po108 = n2351 | n2352;
  assign po113 = n2359 | n2360;
  assign po114 = n2367 | n2368;
  assign n2762 = n2379 | n2380;
  assign n2763 = n2387 | n2388;
  assign n2764 = n2402 | n2403;
  assign n2765 = n2410 | n2411;
  assign po124 = n2422 | n2423;
  assign n2767 = n2427 | n2428;
  assign po131 = n2432 | n2433;
  assign po125 = n2444 | n2445;
  assign po128 = n2454 | n2455;
  assign n2771 = n2457 | n2458;
  assign po135 = n2461 | n2462;
  assign po0 = pi108;
  assign po1 = pi83;
  assign po2 = pi104;
  assign po3 = pi103;
  assign po4 = pi102;
  assign po5 = pi105;
  assign po6 = pi107;
  assign po7 = pi101;
  assign po8 = pi126;
  assign po9 = pi121;
  assign po10 = pi1;
  assign po11 = pi0;
  assign po13 = pi130;
  assign po14 = pi128;
  assign po15 = ~n2535;
  assign po16 = ~n2543;
  assign po69 = ~n1548;
  assign po75 = ~n1830;
  assign po77 = ~n2729;
  assign po78 = ~n2730;
  assign po79 = ~n2731;
  assign po80 = ~n2732;
  assign po81 = ~n2733;
  assign po82 = ~n2734;
  assign po83 = ~n2735;
  assign po84 = ~n2736;
  assign po85 = ~n2737;
  assign po86 = ~n2738;
  assign po87 = ~n2739;
  assign po88 = ~n2740;
  assign po89 = ~n2741;
  assign po90 = ~n2742;
  assign po91 = ~n2743;
  assign po92 = ~n2744;
  assign po98 = ~n1933;
  assign po116 = ~n1971;
  assign po117 = ~n2391;
  assign po118 = ~n2414;
  assign po119 = ~n1673;
  assign po120 = ~n2001;
  assign po122 = ~n2031;
  assign po123 = ~n2061;
  assign po129 = ~n1824;
  assign po132 = ~n2434;
  assign po137 = ~n2463;
  assign po138 = ~n2464;
endmodule
