module alu4_cl ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13,
    po0, po1, po2, po3, po4, po5, po6, po7  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13;
  output po0, po1, po2, po3, po4, po5, po6, po7;
  wire n23, n24, n25, n26, n27, n28, n29,
    n30, n31, n32, n33, n34, n35, n36, n37,
    n38, n39, n40, n41, n42, n43, n44, n45,
    n46, n47, n48, n49, n50, n51, n52, n53,
    n54, n55, n56, n57, n58, n59, n60, n61,
    n62, n63, n64, n65, n66, n67, n68, n69,
    n70, n71, n72, n73, n74, n75, n76, n77,
    n78, n79, n80, n81, n82, n83, n84, n85,
    n86, n87, n88, n89, n90, n91, n92, n93,
    n94, n95, n96, n97, n98, n99, n100,
    n101, n102, n103, n104, n105, n106, n107,
    n108, n109, n110, n111, n112, n113, n114,
    n115, n116, n117, n118, n119, n120, n121,
    n122, n123, n124, n125, n126, n127, n128,
    n129, n130, n131, n132, n133, n134, n135,
    n136, n137, n138, n139, n140, n141, n142,
    n143, n144, n145, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156,
    n157, n158, n159, n160, n161, n162, n163,
    n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177,
    n178, n180, n181, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192,
    n193, n194, n195, n196, n197, n198, n199,
    n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213,
    n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227,
    n228, n229, n230, n231, n232, n233, n234,
    n235, n236, n237, n238, n239, n240, n241,
    n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n327, n328, n329, n330, n331, n332, n333,
    n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403,
    n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416, n417,
    n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438,
    n439, n440, n441, n442, n443, n444, n445,
    n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n470, n472, n473, n474,
    n475, n476, n477, n478, n479, n480, n481,
    n482, n483, n484, n485, n486, n488, n489,
    n490, n491, n492, n493, n494, n495, n496,
    n497, n498, n499, n500, n501, n502, n503,
    n504, n505, n506, n507, n508, n509, n510,
    n511, n512, n513, n514, n515, n516, n517,
    n518, n519, n520, n521, n522, n523, n524,
    n525, n526, n527, n528, n529, n530, n531,
    n532, n533, n534, n535, n536, n537, n538,
    n539, n540, n541, n542, n543, n544, n545,
    n546, n547, n548, n549, n550, n551, n552,
    n553, n554, n555, n556, n557, n558, n559,
    n560, n561, n562, n563, n564, n565, n566,
    n567, n568, n569, n570, n571, n572, n573,
    n574, n575, n576, n577, n578, n579, n580,
    n581, n582, n583, n584, n585, n586, n587,
    n588, n589, n590, n591, n592, n593, n594,
    n595, n596, n597, n598, n599, n600, n601,
    n602, n603, n604, n605, n606, n608, n609,
    n610, n611, n612, n613, n614, n615, n616,
    n617, n618, n619, n620, n621, n622, n624,
    n625, n626, n627, n628, n629, n630, n631,
    n632, n633, n634, n635, n636, n637, n638,
    n639, n640, n641, n642, n643, n644, n645,
    n646, n647, n649, n650;
  assign n23 = pi00 & pi11;
  assign n24 = ~pi08 & ~pi09;
  assign n25 = ~pi10 & ~n24;
  assign n26 = n23 & ~n25;
  assign n27 = pi09 & pi11;
  assign n28 = ~pi10 & ~pi13;
  assign n29 = ~n27 & n28;
  assign n30 = ~pi08 & n29;
  assign n31 = ~pi00 & n30;
  assign n32 = ~pi00 & ~pi04;
  assign n33 = pi08 & ~pi09;
  assign n34 = ~pi10 & pi13;
  assign n35 = ~pi10 & ~pi11;
  assign n36 = ~pi13 & ~n35;
  assign n37 = n33 & ~n34;
  assign n38 = ~n36 & n37;
  assign n39 = ~n32 & n38;
  assign n40 = pi10 & ~pi11;
  assign n41 = pi08 & pi09;
  assign n42 = n40 & n41;
  assign n43 = pi08 & pi10;
  assign n44 = ~pi09 & pi11;
  assign n45 = ~pi13 & n44;
  assign n46 = n43 & n45;
  assign n47 = ~pi08 & pi09;
  assign n48 = pi13 & n47;
  assign n49 = ~n40 & n48;
  assign n50 = ~n42 & ~n46;
  assign n51 = ~n49 & n50;
  assign n52 = ~pi04 & ~n51;
  assign n53 = ~n24 & ~n41;
  assign n54 = pi11 & n34;
  assign n55 = ~n53 & n54;
  assign n56 = ~pi09 & ~pi11;
  assign n57 = ~pi08 & pi10;
  assign n58 = n56 & n57;
  assign n59 = ~n55 & ~n58;
  assign n60 = pi00 & pi04;
  assign n61 = ~n59 & n60;
  assign n62 = ~n32 & ~n60;
  assign n63 = ~pi00 & ~n40;
  assign n64 = n48 & ~n63;
  assign n65 = n62 & n64;
  assign n66 = ~n39 & ~n65;
  assign n67 = ~n61 & n66;
  assign n68 = ~n52 & n67;
  assign n69 = ~n31 & n68;
  assign n70 = ~pi08 & ~pi10;
  assign n71 = pi04 & n70;
  assign n72 = ~n25 & ~n41;
  assign n73 = ~n40 & n72;
  assign n74 = ~pi09 & n73;
  assign n75 = ~n71 & ~n74;
  assign n76 = ~n69 & ~n75;
  assign n77 = ~pi11 & ~n57;
  assign n78 = ~pi08 & pi11;
  assign n79 = ~pi00 & ~n78;
  assign n80 = pi04 & ~n77;
  assign n81 = ~n79 & n80;
  assign n82 = pi00 & ~n68;
  assign n83 = n43 & n82;
  assign n84 = ~pi08 & n40;
  assign n85 = n32 & n84;
  assign n86 = pi09 & ~n85;
  assign n87 = ~n81 & n86;
  assign n88 = ~n83 & n87;
  assign n89 = ~pi00 & pi04;
  assign n90 = pi08 & ~pi10;
  assign n91 = pi11 & n90;
  assign n92 = n89 & n91;
  assign n93 = pi08 & n35;
  assign n94 = ~n57 & ~n93;
  assign n95 = n69 & ~n94;
  assign n96 = pi08 & n40;
  assign n97 = ~n23 & ~n96;
  assign n98 = ~pi04 & ~n97;
  assign n99 = ~pi09 & ~n92;
  assign n100 = ~n98 & n99;
  assign n101 = ~n95 & n100;
  assign n102 = ~n88 & ~n101;
  assign n103 = ~n26 & ~n76;
  assign n104 = ~n102 & n103;
  assign n105 = ~pi13 & ~n104;
  assign n106 = ~pi09 & n90;
  assign n107 = n62 & n106;
  assign n108 = pi04 & n90;
  assign n109 = ~pi00 & n69;
  assign n110 = pi09 & pi13;
  assign n111 = n78 & n110;
  assign n112 = ~n109 & n111;
  assign n113 = pi13 & n40;
  assign n114 = n41 & n82;
  assign n115 = n33 & n60;
  assign n116 = n24 & n69;
  assign n117 = ~n114 & ~n115;
  assign n118 = ~n116 & n117;
  assign n119 = n113 & ~n118;
  assign n120 = ~n112 & ~n119;
  assign n121 = pi00 & ~pi08;
  assign n122 = n120 & n121;
  assign n123 = ~n108 & ~n122;
  assign n124 = n56 & ~n123;
  assign n125 = ~pi00 & n58;
  assign n126 = pi09 & n78;
  assign n127 = n34 & n126;
  assign n128 = n60 & n127;
  assign n129 = n43 & n56;
  assign n130 = pi13 & n129;
  assign n131 = n120 & n130;
  assign n132 = ~n128 & ~n131;
  assign n133 = ~pi10 & n126;
  assign n134 = n132 & n133;
  assign n135 = ~n120 & ~n125;
  assign n136 = ~n134 & n135;
  assign n137 = ~n132 & n133;
  assign n138 = ~n42 & n120;
  assign n139 = ~n137 & n138;
  assign n140 = ~n136 & ~n139;
  assign n141 = ~pi00 & pi11;
  assign n142 = ~n25 & n141;
  assign n143 = n129 & n132;
  assign n144 = ~n69 & ~n142;
  assign n145 = ~n143 & n144;
  assign n146 = n23 & ~n41;
  assign n147 = pi08 & n56;
  assign n148 = ~n132 & n147;
  assign n149 = ~n146 & ~n148;
  assign n150 = pi10 & ~n149;
  assign n151 = ~n84 & ~n90;
  assign n152 = pi09 & ~n151;
  assign n153 = ~n35 & n152;
  assign n154 = n69 & ~n153;
  assign n155 = ~n150 & n154;
  assign n156 = ~n145 & ~n155;
  assign n157 = pi09 & n43;
  assign n158 = n141 & n157;
  assign n159 = pi09 & ~n69;
  assign n160 = ~pi00 & ~n159;
  assign n161 = ~pi09 & n69;
  assign n162 = pi11 & ~n161;
  assign n163 = n70 & ~n160;
  assign n164 = ~n162 & n163;
  assign n165 = ~n107 & ~n158;
  assign n166 = ~n164 & n165;
  assign n167 = ~n124 & n166;
  assign n168 = ~n140 & n167;
  assign n169 = ~n156 & n168;
  assign n170 = pi13 & ~n169;
  assign n171 = pi12 & ~n170;
  assign n172 = ~pi12 & n170;
  assign n173 = pi13 & ~n172;
  assign n174 = ~n171 & n173;
  assign n175 = n45 & n57;
  assign n176 = n93 & n110;
  assign n177 = ~n175 & ~n176;
  assign n178 = ~n105 & n177;
  assign po0 = n174 | ~n178;
  assign n180 = ~pi08 & pi13;
  assign n181 = ~pi09 & pi10;
  assign n182 = n23 & n181;
  assign n183 = ~pi01 & ~pi05;
  assign n184 = n89 & n183;
  assign n185 = ~pi01 & ~n40;
  assign n186 = pi01 & pi05;
  assign n187 = ~n183 & ~n186;
  assign n188 = ~n89 & ~n185;
  assign n189 = n187 & n188;
  assign n190 = ~n184 & ~n189;
  assign n191 = pi09 & ~n190;
  assign n192 = ~n182 & ~n191;
  assign n193 = n180 & ~n192;
  assign n194 = ~pi09 & n40;
  assign n195 = pi13 & n194;
  assign n196 = n59 & ~n195;
  assign n197 = n64 & n89;
  assign n198 = n196 & ~n197;
  assign n199 = n186 & ~n198;
  assign n200 = ~pi05 & ~n51;
  assign n201 = n38 & ~n183;
  assign n202 = ~pi01 & n30;
  assign n203 = ~n201 & ~n202;
  assign n204 = ~n200 & n203;
  assign n205 = ~n199 & n204;
  assign n206 = ~n193 & n205;
  assign n207 = n82 & ~n206;
  assign n208 = ~n82 & n206;
  assign n209 = ~n207 & ~n208;
  assign n210 = pi11 & n72;
  assign n211 = n209 & n210;
  assign n212 = ~pi01 & n206;
  assign n213 = n111 & ~n212;
  assign n214 = pi09 & n206;
  assign n215 = ~pi05 & ~pi09;
  assign n216 = pi01 & pi08;
  assign n217 = ~n215 & n216;
  assign n218 = ~pi08 & n206;
  assign n219 = ~n217 & ~n218;
  assign n220 = n113 & ~n214;
  assign n221 = ~n219 & n220;
  assign n222 = ~n213 & ~n221;
  assign n223 = pi00 & ~n120;
  assign n224 = n222 & ~n223;
  assign n225 = ~n120 & ~n222;
  assign n226 = pi00 & n225;
  assign n227 = ~n224 & ~n226;
  assign n228 = n58 & n227;
  assign n229 = ~n211 & ~n228;
  assign n230 = ~pi01 & ~n229;
  assign n231 = n120 & n222;
  assign n232 = ~n225 & ~n231;
  assign n233 = n157 & ~n232;
  assign n234 = pi09 & n70;
  assign n235 = ~n206 & n234;
  assign n236 = ~n233 & ~n235;
  assign n237 = ~pi11 & ~n236;
  assign n238 = ~pi05 & ~n60;
  assign n239 = n106 & n238;
  assign n240 = n73 & ~n209;
  assign n241 = n23 & n157;
  assign n242 = n35 & ~n41;
  assign n243 = ~n239 & ~n242;
  assign n244 = ~n241 & n243;
  assign n245 = ~n240 & n244;
  assign n246 = pi01 & ~n245;
  assign n247 = n69 & n206;
  assign n248 = n153 & ~n247;
  assign n249 = ~pi11 & n234;
  assign n250 = ~n248 & ~n249;
  assign n251 = ~n69 & ~n206;
  assign n252 = ~n250 & n251;
  assign n253 = n153 & n247;
  assign n254 = ~pi00 & ~pi01;
  assign n255 = n157 & n254;
  assign n256 = n60 & n183;
  assign n257 = n106 & n256;
  assign n258 = ~n255 & ~n257;
  assign n259 = pi11 & ~n258;
  assign n260 = ~pi01 & pi05;
  assign n261 = ~n60 & ~n260;
  assign n262 = n60 & ~n186;
  assign n263 = n106 & ~n261;
  assign n264 = ~n262 & n263;
  assign n265 = pi01 & ~pi08;
  assign n266 = ~n227 & n265;
  assign n267 = pi05 & n90;
  assign n268 = n127 & n186;
  assign n269 = n130 & n222;
  assign n270 = ~n268 & ~n269;
  assign n271 = ~n69 & ~n132;
  assign n272 = ~n270 & n271;
  assign n273 = n270 & ~n271;
  assign n274 = ~n272 & ~n273;
  assign n275 = ~n206 & ~n274;
  assign n276 = n206 & n274;
  assign n277 = ~n275 & ~n276;
  assign n278 = n43 & ~n277;
  assign n279 = ~n266 & ~n267;
  assign n280 = ~n278 & n279;
  assign n281 = n56 & ~n280;
  assign n282 = ~n120 & n128;
  assign n283 = ~n270 & n282;
  assign n284 = n270 & ~n282;
  assign n285 = ~n283 & ~n284;
  assign n286 = n222 & ~n285;
  assign n287 = ~n222 & n285;
  assign n288 = n133 & ~n286;
  assign n289 = ~n287 & n288;
  assign n290 = ~n259 & ~n264;
  assign n291 = ~n253 & n290;
  assign n292 = ~n252 & n291;
  assign n293 = ~n246 & n292;
  assign n294 = ~n237 & n293;
  assign n295 = ~n230 & n294;
  assign n296 = ~n289 & n295;
  assign n297 = ~n281 & n296;
  assign n298 = n173 & ~n297;
  assign n299 = n172 & n297;
  assign n300 = pi01 & pi11;
  assign n301 = ~n96 & ~n300;
  assign n302 = ~pi05 & ~n301;
  assign n303 = ~n94 & n206;
  assign n304 = n91 & n260;
  assign n305 = ~pi09 & ~n304;
  assign n306 = ~n302 & n305;
  assign n307 = ~n303 & n306;
  assign n308 = ~n84 & ~n300;
  assign n309 = ~n187 & ~n308;
  assign n310 = pi05 & n78;
  assign n311 = pi09 & ~n310;
  assign n312 = ~n309 & n311;
  assign n313 = ~n307 & ~n312;
  assign n314 = pi11 & ~n25;
  assign n315 = n157 & ~n206;
  assign n316 = ~n314 & ~n315;
  assign n317 = pi01 & ~n316;
  assign n318 = pi05 & n70;
  assign n319 = ~n74 & ~n318;
  assign n320 = ~n206 & ~n319;
  assign n321 = ~n313 & ~n320;
  assign n322 = ~n317 & n321;
  assign n323 = ~pi13 & ~n322;
  assign n324 = n177 & ~n323;
  assign n325 = ~n298 & n324;
  assign po1 = n299 | ~n325;
  assign n327 = n181 & n300;
  assign n328 = pi01 & ~pi05;
  assign n329 = ~n89 & ~n260;
  assign n330 = ~n328 & ~n329;
  assign n331 = ~pi06 & ~n330;
  assign n332 = pi09 & n331;
  assign n333 = pi06 & n40;
  assign n334 = n330 & n333;
  assign n335 = ~n332 & ~n334;
  assign n336 = pi02 & ~n335;
  assign n337 = pi06 & n330;
  assign n338 = ~n330 & ~n333;
  assign n339 = ~pi02 & pi09;
  assign n340 = ~n337 & n339;
  assign n341 = ~n338 & n340;
  assign n342 = ~n327 & ~n341;
  assign n343 = ~n336 & n342;
  assign n344 = n180 & ~n343;
  assign n345 = ~pi02 & n30;
  assign n346 = pi02 & pi06;
  assign n347 = ~n196 & n346;
  assign n348 = ~pi02 & ~pi06;
  assign n349 = n38 & ~n348;
  assign n350 = ~pi06 & ~n51;
  assign n351 = ~n345 & ~n349;
  assign n352 = ~n347 & n351;
  assign n353 = ~n350 & n352;
  assign n354 = ~n344 & n353;
  assign n355 = ~n94 & n354;
  assign n356 = ~pi06 & n96;
  assign n357 = ~n355 & ~n356;
  assign n358 = ~pi09 & ~n357;
  assign n359 = ~pi02 & n44;
  assign n360 = n90 & n359;
  assign n361 = n70 & ~n354;
  assign n362 = ~n126 & ~n360;
  assign n363 = ~n361 & n362;
  assign n364 = pi06 & ~n363;
  assign n365 = pi02 & pi11;
  assign n366 = ~pi06 & ~pi09;
  assign n367 = n25 & ~n366;
  assign n368 = n365 & ~n367;
  assign n369 = pi02 & n157;
  assign n370 = ~n74 & ~n369;
  assign n371 = ~n354 & ~n370;
  assign n372 = ~n346 & ~n348;
  assign n373 = ~n84 & ~n365;
  assign n374 = pi09 & ~n372;
  assign n375 = ~n373 & n374;
  assign n376 = ~n368 & ~n375;
  assign n377 = ~n371 & n376;
  assign n378 = ~n358 & n377;
  assign n379 = ~n364 & n378;
  assign n380 = ~pi13 & ~n379;
  assign n381 = ~n250 & ~n354;
  assign n382 = pi06 & n90;
  assign n383 = n127 & n346;
  assign n384 = ~pi02 & n354;
  assign n385 = n111 & ~n384;
  assign n386 = pi09 & n354;
  assign n387 = ~pi08 & ~n354;
  assign n388 = pi02 & ~n366;
  assign n389 = pi08 & ~n388;
  assign n390 = n113 & ~n389;
  assign n391 = ~n386 & n390;
  assign n392 = ~n387 & n391;
  assign n393 = ~n385 & ~n392;
  assign n394 = n130 & n393;
  assign n395 = ~n383 & ~n394;
  assign n396 = n354 & n395;
  assign n397 = ~n354 & ~n395;
  assign n398 = ~n396 & ~n397;
  assign n399 = ~n273 & ~n276;
  assign n400 = ~n398 & n399;
  assign n401 = n398 & ~n399;
  assign n402 = ~n400 & ~n401;
  assign n403 = n43 & ~n402;
  assign n404 = pi01 & ~n224;
  assign n405 = ~n226 & ~n404;
  assign n406 = n393 & n405;
  assign n407 = ~n393 & ~n405;
  assign n408 = ~n406 & ~n407;
  assign n409 = pi02 & ~pi08;
  assign n410 = ~n408 & n409;
  assign n411 = ~n382 & ~n410;
  assign n412 = ~n403 & n411;
  assign n413 = n56 & ~n412;
  assign n414 = n58 & n408;
  assign n415 = ~pi01 & ~n207;
  assign n416 = ~n208 & ~n415;
  assign n417 = n210 & ~n354;
  assign n418 = ~n416 & n417;
  assign n419 = ~n414 & ~n418;
  assign n420 = ~pi02 & ~n419;
  assign n421 = ~n222 & ~n284;
  assign n422 = ~n283 & ~n421;
  assign n423 = n395 & n422;
  assign n424 = ~n395 & ~n422;
  assign n425 = ~n423 & ~n424;
  assign n426 = ~n393 & n425;
  assign n427 = n393 & ~n425;
  assign n428 = n133 & ~n426;
  assign n429 = ~n427 & n428;
  assign n430 = n231 & n393;
  assign n431 = ~n231 & ~n393;
  assign n432 = ~pi11 & ~n430;
  assign n433 = ~n431 & n432;
  assign n434 = ~pi02 & n254;
  assign n435 = pi02 & ~n254;
  assign n436 = pi11 & ~n434;
  assign n437 = ~n435 & n436;
  assign n438 = n157 & ~n437;
  assign n439 = ~n433 & n438;
  assign n440 = ~n354 & n416;
  assign n441 = n354 & ~n416;
  assign n442 = ~n440 & ~n441;
  assign n443 = n73 & ~n442;
  assign n444 = ~n242 & ~n443;
  assign n445 = pi02 & ~n444;
  assign n446 = ~pi02 & n210;
  assign n447 = n416 & n446;
  assign n448 = ~n253 & ~n447;
  assign n449 = n354 & ~n448;
  assign n450 = pi11 & n348;
  assign n451 = ~n346 & ~n450;
  assign n452 = ~n60 & ~n186;
  assign n453 = ~n183 & ~n452;
  assign n454 = ~n451 & n453;
  assign n455 = n372 & ~n453;
  assign n456 = ~n454 & ~n455;
  assign n457 = n106 & ~n456;
  assign n458 = ~n381 & ~n457;
  assign n459 = ~n449 & n458;
  assign n460 = ~n445 & n459;
  assign n461 = ~n439 & n460;
  assign n462 = ~n420 & n461;
  assign n463 = ~n429 & n462;
  assign n464 = ~n413 & n463;
  assign n465 = pi13 & ~n464;
  assign n466 = n172 & ~n297;
  assign n467 = n465 & n466;
  assign n468 = ~n465 & ~n466;
  assign n469 = ~n467 & ~n468;
  assign n470 = n177 & ~n380;
  assign po2 = n469 | ~n470;
  assign n472 = ~n396 & ~n401;
  assign n473 = pi02 & ~n337;
  assign n474 = ~n331 & ~n473;
  assign n475 = n113 & n474;
  assign n476 = ~n194 & ~n475;
  assign n477 = pi07 & n113;
  assign n478 = n476 & n477;
  assign n479 = ~n29 & ~n478;
  assign n480 = ~pi03 & ~n479;
  assign n481 = n181 & n365;
  assign n482 = ~pi03 & ~pi07;
  assign n483 = pi09 & n482;
  assign n484 = n474 & n483;
  assign n485 = ~n481 & ~n484;
  assign n486 = pi13 & ~n485;
  assign po5 = pi03 & pi07;
  assign n488 = ~n476 & po5;
  assign n489 = ~n486 & ~n488;
  assign n490 = ~n480 & n489;
  assign n491 = ~pi08 & ~n490;
  assign n492 = pi03 & n48;
  assign n493 = ~n474 & n492;
  assign n494 = n51 & ~n493;
  assign n495 = ~pi07 & ~n494;
  assign n496 = n38 & ~n482;
  assign n497 = ~n495 & ~n496;
  assign n498 = ~n491 & n497;
  assign n499 = ~n55 & ~n195;
  assign n500 = po5 & ~n499;
  assign n501 = n498 & ~n500;
  assign n502 = n127 & po5;
  assign n503 = ~pi03 & n498;
  assign n504 = n111 & ~n503;
  assign n505 = pi03 & ~n501;
  assign n506 = n41 & n505;
  assign n507 = n24 & n501;
  assign n508 = n33 & po5;
  assign n509 = ~n507 & ~n508;
  assign n510 = ~n506 & n509;
  assign n511 = n113 & ~n510;
  assign n512 = ~n504 & ~n511;
  assign n513 = n130 & n512;
  assign n514 = ~n502 & ~n513;
  assign n515 = n501 & n514;
  assign n516 = ~n501 & ~n514;
  assign n517 = ~n515 & ~n516;
  assign n518 = n472 & ~n517;
  assign n519 = ~n472 & n517;
  assign n520 = ~n518 & ~n519;
  assign n521 = pi08 & ~n520;
  assign n522 = pi02 & ~n406;
  assign n523 = ~n407 & ~n522;
  assign n524 = n512 & n523;
  assign n525 = ~pi08 & ~n524;
  assign n526 = ~n512 & ~n523;
  assign n527 = ~pi03 & ~n526;
  assign n528 = n525 & n527;
  assign n529 = ~n521 & ~n528;
  assign n530 = n194 & ~n529;
  assign n531 = ~n393 & ~n423;
  assign n532 = ~n424 & ~n531;
  assign n533 = n512 & n532;
  assign n534 = ~n512 & ~n532;
  assign n535 = ~n533 & ~n534;
  assign n536 = ~n514 & ~n535;
  assign n537 = n514 & n535;
  assign n538 = ~n536 & ~n537;
  assign n539 = n234 & ~n538;
  assign n540 = ~pi03 & n157;
  assign n541 = n434 & n540;
  assign n542 = ~n348 & ~n455;
  assign n543 = n106 & n482;
  assign n544 = n542 & n543;
  assign n545 = ~n541 & ~n544;
  assign n546 = ~n539 & n545;
  assign n547 = pi11 & ~n546;
  assign n548 = n430 & n512;
  assign n549 = ~n430 & ~n512;
  assign n550 = ~n548 & ~n549;
  assign n551 = n157 & ~n550;
  assign n552 = pi07 & n106;
  assign n553 = ~n524 & ~n526;
  assign n554 = pi03 & n24;
  assign n555 = ~n553 & n554;
  assign n556 = ~n551 & ~n552;
  assign n557 = ~n555 & n556;
  assign n558 = ~pi11 & ~n557;
  assign n559 = po5 & n542;
  assign n560 = ~po5 & ~n542;
  assign n561 = pi03 & n560;
  assign n562 = ~n559 & ~n561;
  assign n563 = n106 & ~n562;
  assign n564 = ~n542 & n552;
  assign n565 = ~pi02 & ~n440;
  assign n566 = ~n441 & ~n565;
  assign n567 = ~n501 & n566;
  assign n568 = n501 & ~n566;
  assign n569 = ~n567 & ~n568;
  assign n570 = n210 & n569;
  assign n571 = ~pi03 & ~n564;
  assign n572 = ~n570 & n571;
  assign n573 = n73 & ~n569;
  assign n574 = pi03 & ~n242;
  assign n575 = ~n573 & n574;
  assign n576 = ~n572 & ~n575;
  assign n577 = n249 & ~n501;
  assign n578 = n247 & n354;
  assign n579 = n501 & n578;
  assign n580 = ~n501 & ~n578;
  assign n581 = ~n579 & ~n580;
  assign n582 = n153 & ~n581;
  assign n583 = pi03 & pi11;
  assign n584 = n157 & n583;
  assign n585 = ~n434 & n584;
  assign n586 = ~n563 & ~n585;
  assign n587 = ~n577 & n586;
  assign n588 = ~n582 & n587;
  assign n589 = ~n576 & n588;
  assign n590 = ~n558 & n589;
  assign n591 = ~n547 & n590;
  assign n592 = ~n530 & n591;
  assign n593 = pi13 & ~n592;
  assign n594 = ~n467 & ~n593;
  assign n595 = n467 & ~n592;
  assign n596 = ~n594 & ~n595;
  assign n597 = pi07 & n70;
  assign n598 = ~n74 & ~n597;
  assign n599 = ~n501 & ~n598;
  assign n600 = ~pi07 & ~pi09;
  assign n601 = n25 & ~n600;
  assign n602 = n583 & ~n601;
  assign n603 = ~pi03 & n44;
  assign n604 = n90 & n603;
  assign n605 = ~n126 & ~n604;
  assign n606 = pi07 & ~n605;
  assign po4 = n482 | po5;
  assign n608 = ~n84 & ~n583;
  assign n609 = po4 & ~n608;
  assign n610 = n43 & n505;
  assign n611 = pi09 & ~n609;
  assign n612 = ~n610 & n611;
  assign n613 = ~pi07 & n96;
  assign n614 = ~n94 & n501;
  assign n615 = ~pi09 & ~n613;
  assign n616 = ~n614 & n615;
  assign n617 = ~n612 & ~n616;
  assign n618 = ~n602 & ~n606;
  assign n619 = ~n599 & n618;
  assign n620 = ~n617 & n619;
  assign n621 = ~pi13 & ~n620;
  assign n622 = n177 & ~n621;
  assign po3 = n596 | ~n622;
  assign n624 = n152 & n579;
  assign n625 = n234 & ~n533;
  assign n626 = ~n537 & n625;
  assign n627 = n106 & ~n482;
  assign n628 = ~n560 & n627;
  assign n629 = ~n503 & n566;
  assign n630 = ~n505 & ~n629;
  assign n631 = n72 & ~n630;
  assign n632 = pi11 & ~n541;
  assign n633 = ~n628 & n632;
  assign n634 = ~n631 & n633;
  assign n635 = ~n626 & n634;
  assign n636 = pi10 & ~n548;
  assign n637 = n41 & ~n636;
  assign n638 = n525 & ~n527;
  assign n639 = pi08 & ~n515;
  assign n640 = ~n519 & n639;
  assign n641 = ~n638 & ~n640;
  assign n642 = n181 & ~n641;
  assign n643 = ~pi11 & ~n637;
  assign n644 = ~n642 & n643;
  assign n645 = ~n635 & ~n644;
  assign n646 = ~n624 & ~n645;
  assign n647 = ~n595 & n646;
  assign po6 = pi13 & ~n647;
  assign n649 = ~n62 & ~n187;
  assign n650 = ~n372 & po4;
  assign po7 = n649 & n650;
endmodule
