module i2c ( 
    pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8, pi9,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19,
    pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29,
    pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38, pi39,
    pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48, pi49,
    pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59,
    pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69,
    pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79,
    pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88, pi89,
    pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97, pi98, pi99,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146,
    po0, po1, po2, po3, po4, po5, po6, po7, po8, po9,
    po10, po11, po12, po13, po14, po15, po16, po17, po18, po19,
    po20, po21, po22, po23, po24, po25, po26, po27, po28, po29,
    po30, po31, po32, po33, po34, po35, po36, po37, po38, po39,
    po40, po41, po42, po43, po44, po45, po46, po47, po48, po49,
    po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66, po67, po68, po69,
    po70, po71, po72, po73, po74, po75, po76, po77, po78, po79,
    po80, po81, po82, po83, po84, po85, po86, po87, po88, po89,
    po90, po91, po92, po93, po94, po95, po96, po97, po98, po99,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141  );
  input  pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8,
    pi9, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18,
    pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28,
    pi29, pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38,
    pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48,
    pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58,
    pi59, pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68,
    pi69, pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78,
    pi79, pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88,
    pi89, pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97, pi98,
    pi99, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146;
  output po0, po1, po2, po3, po4, po5, po6, po7, po8, po9,
    po10, po11, po12, po13, po14, po15, po16, po17, po18, po19,
    po20, po21, po22, po23, po24, po25, po26, po27, po28, po29,
    po30, po31, po32, po33, po34, po35, po36, po37, po38, po39,
    po40, po41, po42, po43, po44, po45, po46, po47, po48, po49,
    po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66, po67, po68, po69,
    po70, po71, po72, po73, po74, po75, po76, po77, po78, po79,
    po80, po81, po82, po83, po84, po85, po86, po87, po88, po89,
    po90, po91, po92, po93, po94, po95, po96, po97, po98, po99,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141;
  wire n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n339, n340,
    n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n376,
    n377, n378, n379, n380, n381, n382, n383,
    n384, n385, n386, n387, n388, n389, n390,
    n391, n392, n393, n394, n395, n396, n397,
    n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n409, n410, n411, n412,
    n413, n414, n415, n416, n417, n418, n419,
    n420, n421, n422, n424, n425, n426, n427,
    n428, n429, n430, n431, n432, n433, n434,
    n436, n437, n438, n439, n440, n441, n442,
    n443, n444, n445, n446, n447, n449, n450,
    n451, n452, n453, n454, n455, n456, n457,
    n459, n460, n461, n462, n463, n464, n465,
    n466, n467, n468, n469, n470, n472, n473,
    n474, n475, n476, n477, n478, n479, n481,
    n482, n483, n484, n485, n486, n487, n488,
    n490, n491, n492, n493, n494, n495, n496,
    n497, n499, n500, n501, n502, n503, n504,
    n505, n506, n508, n509, n510, n511, n512,
    n513, n515, n516, n517, n518, n519, n520,
    n521, n522, n523, n524, n526, n527, n528,
    n529, n530, n531, n532, n533, n535, n536,
    n537, n538, n539, n540, n541, n542, n543,
    n544, n545, n546, n547, n548, n549, n550,
    n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n564, n565,
    n566, n567, n568, n569, n570, n572, n573,
    n574, n575, n576, n577, n578, n579, n580,
    n582, n583, n584, n585, n586, n587, n589,
    n590, n591, n592, n593, n595, n596, n597,
    n598, n599, n600, n601, n602, n603, n604,
    n605, n606, n607, n608, n609, n610, n611,
    n613, n614, n615, n616, n617, n618, n620,
    n621, n622, n623, n624, n625, n627, n628,
    n630, n631, n632, n633, n634, n635, n636,
    n637, n638, n639, n640, n641, n642, n643,
    n644, n645, n646, n648, n649, n650, n651,
    n652, n653, n654, n655, n656, n657, n658,
    n659, n660, n661, n662, n663, n664, n665,
    n666, n667, n668, n669, n670, n671, n672,
    n673, n674, n675, n676, n677, n678, n679,
    n680, n681, n682, n683, n684, n685, n686,
    n687, n688, n689, n690, n691, n692, n693,
    n695, n696, n697, n698, n699, n700, n701,
    n702, n703, n704, n705, n706, n707, n709,
    n710, n711, n712, n713, n714, n715, n716,
    n717, n718, n719, n721, n722, n723, n724,
    n725, n726, n727, n728, n729, n730, n731,
    n732, n733, n734, n735, n736, n737, n738,
    n739, n740, n741, n742, n743, n744, n745,
    n746, n747, n748, n749, n750, n751, n752,
    n753, n754, n755, n756, n757, n759, n760,
    n761, n762, n763, n764, n765, n766, n767,
    n768, n769, n770, n771, n772, n773, n774,
    n775, n776, n777, n778, n779, n780, n781,
    n782, n783, n784, n785, n786, n787, n789,
    n790, n791, n792, n793, n794, n796, n797,
    n798, n799, n800, n801, n803, n804, n805,
    n806, n807, n808, n810, n811, n812, n813,
    n814, n815, n817, n818, n819, n820, n821,
    n822, n824, n825, n826, n827, n828, n829,
    n831, n832, n833, n834, n835, n836, n838,
    n839, n840, n841, n842, n843, n845, n846,
    n847, n848, n849, n850, n851, n852, n853,
    n854, n855, n856, n857, n858, n859, n860,
    n861, n862, n863, n864, n866, n867, n868,
    n869, n870, n871, n873, n874, n875, n876,
    n877, n878, n879, n880, n881, n882, n883,
    n884, n885, n886, n887, n889, n890, n891,
    n892, n893, n894, n895, n896, n897, n898,
    n899, n900, n901, n902, n903, n904, n906,
    n907, n908, n909, n910, n911, n912, n913,
    n914, n915, n916, n917, n918, n919, n920,
    n922, n923, n924, n925, n926, n927, n928,
    n929, n930, n931, n932, n933, n934, n935,
    n937, n938, n939, n940, n941, n942, n943,
    n944, n946, n947, n948, n949, n950, n951,
    n952, n953, n954, n955, n956, n957, n958,
    n959, n960, n961, n962, n963, n964, n965,
    n967, n968, n969, n970, n971, n972, n973,
    n974, n975, n976, n977, n978, n980, n981,
    n982, n983, n984, n985, n986, n987, n988,
    n989, n990, n991, n992, n993, n995, n996,
    n997, n998, n999, n1000, n1001, n1002,
    n1003, n1004, n1005, n1006, n1007, n1008,
    n1010, n1011, n1012, n1013, n1014, n1015,
    n1016, n1017, n1018, n1019, n1020, n1021,
    n1022, n1023, n1025, n1026, n1027, n1028,
    n1029, n1030, n1031, n1032, n1033, n1034,
    n1035, n1036, n1037, n1038, n1040, n1041,
    n1042, n1044, n1045, n1046, n1048, n1049,
    n1050, n1051, n1052, n1053, n1054, n1055,
    n1056, n1057, n1059, n1060, n1061, n1064,
    n1066, n1067, n1068, n1069, n1070, n1071,
    n1072, n1073, n1074, n1075, n1076, n1077,
    n1078, n1079, n1080, n1081, n1082, n1083,
    n1084, n1086, n1087, n1088, n1089, n1090,
    n1091, n1092, n1093, n1094, n1095, n1096,
    n1097, n1098, n1099, n1100, n1101, n1103,
    n1104, n1105, n1106, n1107, n1108, n1110,
    n1111, n1112, n1113, n1114, n1115, n1116,
    n1117, n1118, n1119, n1120, n1121, n1122,
    n1123, n1124, n1125, n1126, n1127, n1128,
    n1129, n1131, n1132, n1133, n1135, n1136,
    n1138, n1139, n1140, n1141, n1142, n1143,
    n1144, n1145, n1147, n1148, n1149, n1151,
    n1152, n1153, n1155, n1156, n1157, n1159,
    n1160, n1161, n1162, n1163, n1165, n1166,
    n1167, n1169, n1170, n1171, n1173, n1174,
    n1175, n1177, n1178, n1179, n1181, n1182,
    n1183, n1185, n1186, n1187, n1189, n1190,
    n1191, n1193, n1194, n1195, n1197, n1198,
    n1199, n1201, n1202, n1203, n1205, n1206,
    n1207, n1209, n1210, n1211, n1212, n1213,
    n1215, n1216, n1217, n1219, n1220, n1221,
    n1223, n1224, n1225, n1227, n1228, n1229,
    n1231, n1232, n1233, n1234, n1235, n1236,
    n1237, n1238, n1239, n1240, n1241, n1242,
    n1243, n1244, n1245, n1246, n1247, n1248,
    n1250, n1251, n1252, n1254, n1255, n1256,
    n1257, n1258, n1260, n1261, n1262, n1264,
    n1265, n1266, n1268, n1269, n1270, n1271,
    n1272, n1274, n1275, n1276, n1278, n1279,
    n1280, n1282, n1283, n1284, n1286, n1287,
    n1288, n1290, n1291, n1292, n1294, n1295,
    n1296, n1297, n1298, n1299, n1300, n1302,
    n1303, n1304, n1305, n1306, n1307, n1309,
    n1310, n1311, n1313, n1314, n1315, n1317,
    n1318, n1319, n1321, n1322, n1323, n1325,
    n1326, n1327, n1329, n1330, n1331, n1332,
    n1333, n1334, n1335, n1336, n1337, n1338,
    n1339, n1340, n1341, n1342, n1343, n1344,
    n1345, n1347, n1348, n1349, n1350, n1351,
    n1352, n1353, n1354, n1355, n1356, n1357,
    n1358, n1359, n1360, n1362, n1363, n1364,
    n1365, n1366, n1367, n1368, n1369, n1370,
    n1371, n1372, n1373, n1374, n1375, n1377,
    n1378, n1379, n1380, n1381, n1382, n1383,
    n1384, n1385, n1386, n1387, n1388, n1389,
    n1390, n1392, n1393, n1394, n1395, n1396,
    n1397, n1398, n1399, n1400, n1401, n1402,
    n1403, n1404, n1405, n1406, n1407, n1408,
    n1410, n1411, n1412, n1414, n1415, n1416,
    n1417, n1418, n1419, n1420, n1421, n1422,
    n1423, n1424, n1425, n1426, n1427, n1428,
    n1429, n1430, n1432, n1433, n1434, n1435,
    n1436, n1437, n1438, n1439, n1440, n1441,
    n1442, n1443, n1444, n1445, n1446, n1447,
    n1448, n1450, n1451, n1452, n1454, n1455,
    n1456, n1458, n1459, n1460, n1461, n1463,
    n1464, n1465, n1466, n1468, n1469, n1470,
    n1471, n1473, n1474, n1475, n1476, n1478,
    n1479, n1480, n1483, n1484, n1485, n1486,
    n1489, n1490, n1492, n1497, n1498, n1500;
  assign n291 = ~pi7 & ~pi13;
  assign n292 = ~pi8 & ~pi21;
  assign n293 = ~pi12 & ~pi17;
  assign n294 = n292 & n293;
  assign n295 = ~pi14 & n294;
  assign n296 = ~pi9 & ~pi11;
  assign n297 = ~pi5 & ~pi22;
  assign n298 = ~pi4 & ~pi19;
  assign n299 = ~pi18 & n298;
  assign n300 = ~pi16 & n299;
  assign n301 = n297 & n300;
  assign n302 = n296 & n301;
  assign n303 = ~pi6 & n302;
  assign n304 = n295 & n303;
  assign n305 = n291 & n304;
  assign n306 = pi54 & ~n305;
  assign n307 = ~pi0 & ~n306;
  assign n308 = ~pi56 & ~n297;
  assign n309 = ~pi6 & ~pi12;
  assign n310 = ~pi7 & n292;
  assign n311 = ~pi13 & ~pi14;
  assign n312 = ~n310 & ~n311;
  assign n313 = ~pi13 & pi14;
  assign n314 = pi7 & ~n292;
  assign n315 = pi8 & pi21;
  assign n316 = ~n314 & ~n315;
  assign n317 = ~n310 & n316;
  assign n318 = ~pi13 & ~n317;
  assign n319 = ~pi14 & ~n318;
  assign n320 = ~n313 & ~n319;
  assign n321 = ~pi10 & ~n320;
  assign n322 = ~n312 & n321;
  assign n323 = pi10 & ~pi14;
  assign n324 = ~pi13 & n323;
  assign n325 = n310 & n324;
  assign n326 = ~n322 & ~n325;
  assign n327 = n309 & ~n326;
  assign n328 = ~pi17 & n327;
  assign n329 = n301 & n328;
  assign n330 = ~n308 & ~n329;
  assign n331 = n296 & ~n330;
  assign n332 = ~pi56 & ~n296;
  assign n333 = n297 & n332;
  assign n334 = ~n331 & ~n333;
  assign n335 = pi54 & ~n334;
  assign n336 = ~n307 & ~n335;
  assign n337 = ~pi3 & ~pi129;
  assign po15 = n336 | ~n337;
  assign n339 = ~pi17 & pi54;
  assign n340 = ~pi5 & ~pi6;
  assign n341 = ~pi7 & n340;
  assign n342 = ~pi10 & ~pi22;
  assign n343 = n311 & n342;
  assign n344 = ~pi11 & n292;
  assign n345 = ~pi12 & n344;
  assign n346 = n300 & n345;
  assign n347 = n343 & n346;
  assign n348 = n341 & n347;
  assign n349 = n339 & ~n348;
  assign n350 = ~pi1 & ~n349;
  assign n351 = ~pi5 & n309;
  assign n352 = n291 & n351;
  assign n353 = pi9 & ~n352;
  assign n354 = n342 & ~n353;
  assign n355 = ~pi14 & n354;
  assign n356 = pi7 & ~n351;
  assign n357 = pi5 & ~n309;
  assign n358 = pi6 & pi12;
  assign n359 = ~n357 & ~n358;
  assign n360 = ~n351 & n359;
  assign n361 = ~pi7 & ~n360;
  assign n362 = ~n356 & ~n361;
  assign n363 = ~pi13 & n362;
  assign n364 = ~pi5 & ~pi7;
  assign n365 = n309 & n364;
  assign n366 = pi13 & n365;
  assign n367 = ~pi9 & ~n366;
  assign n368 = ~n363 & n367;
  assign n369 = ~pi17 & n344;
  assign n370 = n300 & n369;
  assign n371 = ~n368 & n370;
  assign n372 = pi54 & n371;
  assign n373 = n355 & n372;
  assign n374 = ~n350 & ~n373;
  assign po16 = ~n337 | n374;
  assign n376 = pi122 & pi127;
  assign n377 = ~pi82 & n376;
  assign n378 = ~pi42 & ~pi44;
  assign n379 = ~pi38 & ~pi40;
  assign n380 = ~pi50 & n379;
  assign n381 = n378 & n380;
  assign n382 = ~pi43 & ~pi47;
  assign n383 = ~pi41 & ~pi46;
  assign n384 = n382 & n383;
  assign n385 = ~pi48 & n384;
  assign n386 = n381 & n385;
  assign n387 = pi82 & ~n386;
  assign n388 = ~pi15 & ~pi20;
  assign n389 = ~pi24 & ~pi49;
  assign n390 = n388 & n389;
  assign n391 = ~pi45 & n390;
  assign n392 = pi82 & ~n391;
  assign n393 = ~n387 & ~n392;
  assign n394 = ~n377 & n393;
  assign n395 = pi2 & ~n394;
  assign n396 = ~pi40 & n378;
  assign n397 = ~pi48 & n382;
  assign n398 = n391 & n397;
  assign n399 = ~pi38 & ~pi50;
  assign n400 = n383 & n399;
  assign n401 = ~pi2 & n400;
  assign n402 = n398 & n401;
  assign n403 = n396 & n402;
  assign n404 = pi82 & ~n403;
  assign n405 = ~pi65 & ~n404;
  assign n406 = ~n376 & n405;
  assign n407 = ~n395 & ~n406;
  assign po17 = ~pi129 & ~n407;
  assign n409 = pi0 & ~pi123;
  assign n410 = ~pi113 & n409;
  assign n411 = ~pi9 & ~pi10;
  assign n412 = n311 & n411;
  assign n413 = ~pi22 & n412;
  assign n414 = n341 & n413;
  assign n415 = ~pi8 & ~pi11;
  assign n416 = n300 & n415;
  assign n417 = ~pi21 & n416;
  assign n418 = n414 & n417;
  assign n419 = n293 & n418;
  assign n420 = ~pi61 & ~n419;
  assign n421 = ~pi118 & n420;
  assign n422 = ~n410 & ~n421;
  assign po18 = ~pi129 & ~n422;
  assign n424 = pi4 & ~pi54;
  assign n425 = ~pi4 & ~pi16;
  assign n426 = pi54 & n425;
  assign n427 = ~pi19 & n426;
  assign n428 = ~pi18 & n427;
  assign n429 = n369 & n428;
  assign n430 = ~pi9 & ~pi22;
  assign n431 = n352 & n430;
  assign n432 = n429 & n431;
  assign n433 = n323 & n432;
  assign n434 = ~n424 & ~n433;
  assign po19 = n337 & ~n434;
  assign n436 = pi5 & ~pi54;
  assign n437 = ~pi59 & n369;
  assign n438 = ~pi7 & ~pi12;
  assign n439 = ~pi6 & ~pi29;
  assign n440 = n438 & n439;
  assign n441 = ~pi25 & n440;
  assign n442 = ~pi5 & n441;
  assign n443 = n437 & n442;
  assign n444 = pi28 & n413;
  assign n445 = n428 & n444;
  assign n446 = n443 & n445;
  assign n447 = ~n436 & ~n446;
  assign po20 = n337 & ~n447;
  assign n449 = pi6 & ~pi54;
  assign n450 = ~pi5 & ~pi28;
  assign n451 = n438 & n450;
  assign n452 = n413 & n451;
  assign n453 = pi25 & n452;
  assign n454 = n437 & n453;
  assign n455 = n428 & n454;
  assign n456 = n439 & n455;
  assign n457 = ~n449 & ~n456;
  assign po21 = n337 & ~n457;
  assign n459 = pi7 & ~pi54;
  assign n460 = ~pi11 & ~pi12;
  assign n461 = ~pi6 & n460;
  assign n462 = ~pi17 & ~pi18;
  assign n463 = ~pi21 & n462;
  assign n464 = ~pi7 & pi8;
  assign n465 = n463 & n464;
  assign n466 = ~pi5 & n465;
  assign n467 = n461 & n466;
  assign n468 = n413 & n467;
  assign n469 = n427 & n468;
  assign n470 = ~n459 & ~n469;
  assign po22 = n337 & ~n470;
  assign n472 = pi8 & ~pi54;
  assign n473 = n415 & n462;
  assign n474 = ~pi10 & ~pi14;
  assign n475 = n431 & n474;
  assign n476 = pi21 & n475;
  assign n477 = n473 & n476;
  assign n478 = n427 & n477;
  assign n479 = ~n472 & ~n478;
  assign po23 = n337 & ~n479;
  assign n481 = pi9 & pi54;
  assign n482 = n343 & n365;
  assign n483 = ~pi8 & n463;
  assign n484 = pi11 & n427;
  assign n485 = n483 & n484;
  assign n486 = n482 & n485;
  assign n487 = ~pi9 & ~n486;
  assign n488 = n337 & ~n487;
  assign po24 = ~n481 & n488;
  assign n490 = pi10 & ~pi54;
  assign n491 = n427 & n430;
  assign n492 = n313 & n491;
  assign n493 = n364 & n461;
  assign n494 = ~pi10 & n483;
  assign n495 = n493 & n494;
  assign n496 = n492 & n495;
  assign n497 = ~n490 & ~n496;
  assign po25 = n337 & ~n497;
  assign n499 = pi11 & ~pi54;
  assign n500 = ~pi21 & n427;
  assign n501 = n411 & n500;
  assign n502 = ~pi14 & pi22;
  assign n503 = n352 & n502;
  assign n504 = n473 & n503;
  assign n505 = n501 & n504;
  assign n506 = ~n499 & ~n505;
  assign po26 = n337 & ~n506;
  assign n508 = pi12 & ~pi54;
  assign n509 = pi18 & n293;
  assign n510 = n344 & n509;
  assign n511 = n414 & n510;
  assign n512 = n427 & n511;
  assign n513 = ~n508 & ~n512;
  assign po27 = n337 & ~n513;
  assign n515 = pi13 & ~pi54;
  assign n516 = n430 & n474;
  assign n517 = ~pi25 & pi29;
  assign n518 = ~pi28 & n517;
  assign n519 = n428 & n437;
  assign n520 = n291 & n519;
  assign n521 = n351 & n520;
  assign n522 = n518 & n521;
  assign n523 = n516 & n522;
  assign n524 = ~n515 & ~n523;
  assign po28 = n337 & ~n524;
  assign n526 = pi14 & pi54;
  assign n527 = n427 & n483;
  assign n528 = ~pi10 & pi13;
  assign n529 = n430 & n528;
  assign n530 = n493 & n529;
  assign n531 = n527 & n530;
  assign n532 = ~pi14 & ~n531;
  assign n533 = n337 & ~n532;
  assign po29 = ~n526 & n533;
  assign n535 = ~pi45 & ~pi48;
  assign n536 = n384 & n535;
  assign n537 = n389 & n536;
  assign n538 = n381 & n537;
  assign n539 = pi15 & ~n538;
  assign n540 = ~pi47 & ~pi48;
  assign n541 = ~pi45 & n540;
  assign n542 = ~pi2 & ~pi20;
  assign n543 = n381 & n383;
  assign n544 = ~pi43 & n543;
  assign n545 = ~n542 & n544;
  assign n546 = ~pi15 & n545;
  assign n547 = n389 & n546;
  assign n548 = n541 & n547;
  assign n549 = ~n539 & ~n548;
  assign n550 = pi82 & ~n549;
  assign n551 = pi15 & n377;
  assign n552 = ~n550 & ~n551;
  assign n553 = n396 & n541;
  assign n554 = ~pi43 & n383;
  assign n555 = n399 & n554;
  assign n556 = n553 & n555;
  assign n557 = ~pi15 & n556;
  assign n558 = n389 & n557;
  assign n559 = pi82 & ~n558;
  assign n560 = ~pi70 & ~n559;
  assign n561 = ~n376 & n560;
  assign n562 = n552 & ~n561;
  assign po30 = ~pi129 & ~n562;
  assign n564 = pi16 & ~pi54;
  assign n565 = ~pi13 & n438;
  assign n566 = ~pi5 & n565;
  assign n567 = pi6 & n566;
  assign n568 = n429 & n567;
  assign n569 = n516 & n568;
  assign n570 = ~n564 & ~n569;
  assign po31 = n337 & ~n570;
  assign n572 = pi17 & ~pi54;
  assign n573 = ~pi28 & n414;
  assign n574 = ~pi25 & n573;
  assign n575 = ~pi29 & n339;
  assign n576 = pi59 & n300;
  assign n577 = n575 & n576;
  assign n578 = n345 & n577;
  assign n579 = n574 & n578;
  assign n580 = ~n572 & ~n579;
  assign po32 = n337 & ~n580;
  assign n582 = pi18 & ~pi54;
  assign n583 = pi16 & n369;
  assign n584 = pi54 & n583;
  assign n585 = n299 & n584;
  assign n586 = n475 & n585;
  assign n587 = ~n582 & ~n586;
  assign po33 = n337 & ~n587;
  assign n589 = pi19 & ~pi54;
  assign n590 = pi17 & n475;
  assign n591 = n344 & n590;
  assign n592 = n428 & n591;
  assign n593 = ~n589 & ~n592;
  assign po34 = n337 & ~n593;
  assign n595 = ~pi49 & n388;
  assign n596 = ~pi24 & n535;
  assign n597 = n382 & n543;
  assign n598 = n596 & n597;
  assign n599 = n595 & n598;
  assign n600 = pi2 & n599;
  assign n601 = ~pi15 & ~pi49;
  assign n602 = n598 & n601;
  assign n603 = pi20 & ~n602;
  assign n604 = ~n600 & ~n603;
  assign n605 = pi82 & ~n604;
  assign n606 = pi20 & n377;
  assign n607 = ~n605 & ~n606;
  assign n608 = pi82 & ~n599;
  assign n609 = ~pi71 & ~n608;
  assign n610 = ~n376 & n609;
  assign n611 = n607 & ~n610;
  assign po35 = ~pi129 & ~n611;
  assign n613 = pi21 & ~pi54;
  assign n614 = ~pi21 & n475;
  assign n615 = pi19 & n614;
  assign n616 = n473 & n615;
  assign n617 = n426 & n616;
  assign n618 = ~n613 & ~n617;
  assign po36 = n337 & ~n618;
  assign n620 = pi22 & ~pi54;
  assign n621 = ~pi7 & n527;
  assign n622 = pi5 & n621;
  assign n623 = n461 & n622;
  assign n624 = n413 & n623;
  assign n625 = ~n620 & ~n624;
  assign po37 = n337 & ~n625;
  assign n627 = ~pi23 & pi55;
  assign n628 = pi61 & ~n627;
  assign po38 = ~pi129 & n628;
  assign n630 = pi82 & ~n556;
  assign n631 = n542 & n601;
  assign n632 = pi82 & ~n631;
  assign n633 = n376 & ~n632;
  assign n634 = ~n630 & ~n633;
  assign n635 = ~pi24 & ~n634;
  assign n636 = ~pi2 & n544;
  assign n637 = n541 & n636;
  assign n638 = n595 & n637;
  assign n639 = pi82 & ~n638;
  assign n640 = ~n376 & ~n639;
  assign n641 = pi63 & n640;
  assign n642 = pi24 & n536;
  assign n643 = pi82 & n381;
  assign n644 = n642 & n643;
  assign n645 = ~pi129 & ~n644;
  assign n646 = ~n641 & n645;
  assign po39 = ~n635 & n646;
  assign n648 = pi85 & ~pi116;
  assign n649 = pi25 & n648;
  assign n650 = ~pi96 & ~pi110;
  assign n651 = ~pi85 & ~n650;
  assign n652 = ~n648 & ~n651;
  assign n653 = pi100 & n652;
  assign n654 = ~n649 & ~n653;
  assign n655 = ~pi26 & ~n654;
  assign n656 = pi25 & ~pi116;
  assign n657 = pi26 & n656;
  assign n658 = ~pi95 & ~pi100;
  assign n659 = ~pi97 & n658;
  assign n660 = ~pi110 & ~n659;
  assign n661 = pi25 & ~n660;
  assign n662 = pi26 & pi116;
  assign n663 = ~n661 & ~n662;
  assign n664 = ~pi51 & ~pi52;
  assign n665 = ~pi39 & n664;
  assign n666 = ~n663 & ~n665;
  assign n667 = ~n657 & ~n666;
  assign n668 = ~pi85 & ~n667;
  assign n669 = ~n655 & ~n668;
  assign n670 = ~pi27 & ~n669;
  assign n671 = ~pi39 & ~pi52;
  assign n672 = ~pi51 & n671;
  assign n673 = pi116 & n672;
  assign n674 = ~n656 & ~n673;
  assign n675 = pi27 & ~n674;
  assign n676 = n661 & n665;
  assign n677 = ~n675 & ~n676;
  assign n678 = ~pi26 & ~pi85;
  assign n679 = ~n677 & n678;
  assign n680 = ~n670 & ~n679;
  assign n681 = ~pi53 & ~n680;
  assign n682 = pi25 & ~pi26;
  assign n683 = ~pi116 & n682;
  assign n684 = pi53 & ~pi85;
  assign n685 = ~pi27 & n684;
  assign n686 = n683 & n685;
  assign n687 = ~n681 & ~n686;
  assign n688 = ~pi58 & ~n687;
  assign n689 = ~pi27 & ~pi85;
  assign n690 = ~pi53 & pi58;
  assign n691 = n683 & n690;
  assign n692 = n689 & n691;
  assign n693 = ~n688 & ~n692;
  assign po40 = n337 & ~n693;
  assign n695 = ~pi27 & ~pi53;
  assign n696 = ~pi58 & n695;
  assign n697 = pi85 & pi116;
  assign n698 = ~pi26 & n697;
  assign n699 = ~pi110 & ~n648;
  assign n700 = ~pi96 & n699;
  assign n701 = ~n662 & n700;
  assign n702 = ~n698 & ~n701;
  assign n703 = pi100 & ~n702;
  assign n704 = ~pi85 & ~n673;
  assign n705 = pi26 & n704;
  assign n706 = ~n703 & ~n705;
  assign n707 = n337 & ~n706;
  assign po41 = n696 & n707;
  assign n709 = ~pi53 & ~pi58;
  assign n710 = ~pi26 & n709;
  assign n711 = pi27 & n704;
  assign n712 = pi95 & ~pi96;
  assign n713 = n699 & n712;
  assign n714 = ~n697 & ~n713;
  assign n715 = pi27 & pi116;
  assign n716 = ~pi100 & ~n715;
  assign n717 = ~n714 & n716;
  assign n718 = ~n711 & ~n717;
  assign n719 = n337 & ~n718;
  assign po42 = n710 & n719;
  assign n721 = ~pi26 & ~pi100;
  assign n722 = ~pi110 & n721;
  assign n723 = n712 & n722;
  assign n724 = pi26 & n673;
  assign n725 = ~n723 & ~n724;
  assign n726 = ~pi27 & ~n725;
  assign n727 = ~pi26 & ~n665;
  assign n728 = ~pi27 & n672;
  assign n729 = ~n727 & ~n728;
  assign n730 = ~n660 & ~n729;
  assign n731 = pi26 & ~pi27;
  assign n732 = ~pi26 & pi27;
  assign n733 = ~n731 & ~n732;
  assign n734 = ~pi116 & ~n733;
  assign n735 = ~n730 & ~n734;
  assign n736 = pi28 & ~n735;
  assign n737 = n715 & n727;
  assign n738 = ~n736 & ~n737;
  assign n739 = ~n726 & n738;
  assign n740 = ~pi85 & ~n739;
  assign n741 = ~pi28 & ~pi116;
  assign n742 = pi85 & ~n741;
  assign n743 = pi100 & pi116;
  assign n744 = ~pi26 & ~pi27;
  assign n745 = ~n743 & n744;
  assign n746 = n742 & n745;
  assign n747 = ~n740 & ~n746;
  assign n748 = ~pi53 & ~n747;
  assign n749 = ~pi27 & pi28;
  assign n750 = ~pi116 & n749;
  assign n751 = ~pi26 & n684;
  assign n752 = n750 & n751;
  assign n753 = ~n748 & ~n752;
  assign n754 = ~pi58 & ~n753;
  assign n755 = n678 & n690;
  assign n756 = n750 & n755;
  assign n757 = ~n754 & ~n756;
  assign po43 = n337 & ~n757;
  assign n759 = pi97 & ~n650;
  assign n760 = n658 & ~n759;
  assign n761 = ~pi110 & ~n760;
  assign n762 = pi29 & ~n761;
  assign n763 = pi97 & n760;
  assign n764 = ~pi58 & ~n763;
  assign n765 = ~n762 & n764;
  assign n766 = ~pi53 & ~n765;
  assign n767 = pi97 & pi116;
  assign n768 = pi29 & ~pi116;
  assign n769 = ~n767 & ~n768;
  assign n770 = pi58 & n769;
  assign n771 = n766 & ~n770;
  assign n772 = pi53 & ~pi58;
  assign n773 = n768 & n772;
  assign n774 = ~n771 & ~n773;
  assign n775 = ~pi27 & ~n774;
  assign n776 = pi27 & n768;
  assign n777 = n709 & n776;
  assign n778 = ~n775 & ~n777;
  assign n779 = ~pi85 & ~n778;
  assign n780 = pi85 & n696;
  assign n781 = n768 & n780;
  assign n782 = ~n779 & ~n781;
  assign n783 = ~pi26 & ~n782;
  assign n784 = ~pi85 & n709;
  assign n785 = n731 & n784;
  assign n786 = n768 & n785;
  assign n787 = ~n783 & ~n786;
  assign po44 = n337 & ~n787;
  assign n789 = pi30 & ~pi109;
  assign n790 = pi60 & pi109;
  assign n791 = ~pi106 & ~n790;
  assign n792 = ~n789 & n791;
  assign n793 = ~pi88 & pi106;
  assign n794 = ~pi129 & ~n793;
  assign po45 = ~n792 & n794;
  assign n796 = pi31 & ~pi109;
  assign n797 = pi30 & pi109;
  assign n798 = ~pi106 & ~n797;
  assign n799 = ~n796 & n798;
  assign n800 = ~pi89 & pi106;
  assign n801 = ~pi129 & ~n800;
  assign po46 = ~n799 & n801;
  assign n803 = pi32 & ~pi109;
  assign n804 = pi31 & pi109;
  assign n805 = ~pi106 & ~n804;
  assign n806 = ~n803 & n805;
  assign n807 = ~pi99 & pi106;
  assign n808 = ~pi129 & ~n807;
  assign po47 = ~n806 & n808;
  assign n810 = pi33 & ~pi109;
  assign n811 = pi32 & pi109;
  assign n812 = ~pi106 & ~n811;
  assign n813 = ~n810 & n812;
  assign n814 = ~pi90 & pi106;
  assign n815 = ~pi129 & ~n814;
  assign po48 = ~n813 & n815;
  assign n817 = pi34 & ~pi109;
  assign n818 = pi33 & pi109;
  assign n819 = ~pi106 & ~n818;
  assign n820 = ~n817 & n819;
  assign n821 = ~pi91 & pi106;
  assign n822 = ~pi129 & ~n821;
  assign po49 = ~n820 & n822;
  assign n824 = pi35 & ~pi109;
  assign n825 = pi34 & pi109;
  assign n826 = ~pi106 & ~n825;
  assign n827 = ~n824 & n826;
  assign n828 = ~pi92 & pi106;
  assign n829 = ~pi129 & ~n828;
  assign po50 = ~n827 & n829;
  assign n831 = pi36 & ~pi109;
  assign n832 = pi35 & pi109;
  assign n833 = ~pi106 & ~n832;
  assign n834 = ~n831 & n833;
  assign n835 = ~pi98 & pi106;
  assign n836 = ~pi129 & ~n835;
  assign po51 = ~n834 & n836;
  assign n838 = pi37 & ~pi109;
  assign n839 = pi36 & pi109;
  assign n840 = ~pi106 & ~n839;
  assign n841 = ~n838 & n840;
  assign n842 = ~pi93 & pi106;
  assign n843 = ~pi129 & ~n842;
  assign po52 = ~n841 & n843;
  assign n845 = pi82 & ~n396;
  assign n846 = ~pi46 & ~pi50;
  assign n847 = ~pi2 & n391;
  assign n848 = n397 & n847;
  assign n849 = ~pi41 & n848;
  assign n850 = n846 & n849;
  assign n851 = pi82 & ~n850;
  assign n852 = n376 & ~n851;
  assign n853 = ~n845 & ~n852;
  assign n854 = ~pi38 & ~n853;
  assign n855 = n396 & n850;
  assign n856 = pi82 & ~n855;
  assign n857 = ~n376 & ~n856;
  assign n858 = pi74 & n857;
  assign n859 = ~pi40 & ~pi42;
  assign n860 = ~pi44 & pi82;
  assign n861 = n859 & n860;
  assign n862 = pi38 & n861;
  assign n863 = ~pi129 & ~n862;
  assign n864 = ~n858 & n863;
  assign po53 = ~n854 & n864;
  assign n866 = pi109 & n664;
  assign n867 = pi39 & ~n866;
  assign n868 = ~pi51 & pi109;
  assign n869 = n671 & n868;
  assign n870 = ~pi106 & ~n869;
  assign n871 = ~n867 & n870;
  assign po54 = ~pi129 & ~n871;
  assign n873 = pi82 & ~n378;
  assign n874 = ~pi46 & n399;
  assign n875 = n849 & n874;
  assign n876 = pi82 & ~n875;
  assign n877 = n376 & ~n876;
  assign n878 = ~n873 & ~n877;
  assign n879 = ~pi40 & ~n878;
  assign n880 = n378 & n875;
  assign n881 = pi82 & ~n880;
  assign n882 = ~n376 & ~n881;
  assign n883 = pi73 & n882;
  assign n884 = ~pi42 & n860;
  assign n885 = pi40 & n884;
  assign n886 = ~pi129 & ~n885;
  assign n887 = ~n883 & n886;
  assign po55 = ~n879 & n887;
  assign n889 = n396 & n874;
  assign n890 = pi82 & ~n889;
  assign n891 = pi82 & ~n848;
  assign n892 = n376 & ~n891;
  assign n893 = ~n890 & ~n892;
  assign n894 = ~pi41 & ~n893;
  assign n895 = n379 & n846;
  assign n896 = n378 & n895;
  assign n897 = n848 & n896;
  assign n898 = pi82 & ~n897;
  assign n899 = ~n376 & ~n898;
  assign n900 = pi76 & n899;
  assign n901 = pi41 & n895;
  assign n902 = n884 & n901;
  assign n903 = ~pi129 & ~n902;
  assign n904 = ~n900 & n903;
  assign po56 = ~n894 & n904;
  assign n906 = pi44 & pi82;
  assign n907 = n849 & n895;
  assign n908 = pi82 & ~n907;
  assign n909 = n376 & ~n908;
  assign n910 = ~n906 & ~n909;
  assign n911 = ~pi42 & ~n910;
  assign n912 = pi42 & n860;
  assign n913 = ~pi129 & ~n912;
  assign n914 = n385 & n847;
  assign n915 = ~pi44 & n914;
  assign n916 = n380 & n915;
  assign n917 = pi82 & ~n916;
  assign n918 = ~n376 & ~n917;
  assign n919 = pi72 & n918;
  assign n920 = n913 & ~n919;
  assign po57 = ~n911 & n920;
  assign n922 = pi82 & ~n543;
  assign n923 = n540 & n847;
  assign n924 = pi82 & ~n923;
  assign n925 = n376 & ~n924;
  assign n926 = ~n922 & ~n925;
  assign n927 = ~pi43 & ~n926;
  assign n928 = n543 & n923;
  assign n929 = pi82 & ~n928;
  assign n930 = ~n376 & ~n929;
  assign n931 = pi77 & n930;
  assign n932 = pi43 & n400;
  assign n933 = n861 & n932;
  assign n934 = ~pi129 & ~n933;
  assign n935 = ~n931 & n934;
  assign po58 = ~n927 & n935;
  assign n937 = ~pi42 & n914;
  assign n938 = n380 & n937;
  assign n939 = pi82 & ~n938;
  assign n940 = ~pi67 & ~n376;
  assign n941 = pi44 & n376;
  assign n942 = ~n940 & ~n941;
  assign n943 = ~n939 & n942;
  assign n944 = ~pi129 & ~n906;
  assign po59 = ~n943 & n944;
  assign n946 = ~pi2 & n388;
  assign n947 = n389 & n946;
  assign n948 = pi82 & ~n947;
  assign n949 = n376 & ~n948;
  assign n950 = ~n387 & ~n949;
  assign n951 = ~pi45 & ~n950;
  assign n952 = ~pi2 & n540;
  assign n953 = n390 & n952;
  assign n954 = n544 & n953;
  assign n955 = pi82 & ~n954;
  assign n956 = ~n376 & ~n955;
  assign n957 = pi68 & n956;
  assign n958 = ~pi41 & n846;
  assign n959 = pi45 & n958;
  assign n960 = n397 & n959;
  assign n961 = ~pi38 & n859;
  assign n962 = n860 & n961;
  assign n963 = n960 & n962;
  assign n964 = ~pi129 & ~n963;
  assign n965 = ~n957 & n964;
  assign po60 = ~n951 & n965;
  assign n967 = pi82 & ~n381;
  assign n968 = pi82 & ~n849;
  assign n969 = n376 & ~n968;
  assign n970 = ~n967 & ~n969;
  assign n971 = ~pi46 & ~n970;
  assign n972 = n381 & n849;
  assign n973 = pi82 & ~n972;
  assign n974 = ~n376 & ~n973;
  assign n975 = pi75 & n974;
  assign n976 = pi46 & n643;
  assign n977 = ~pi129 & ~n976;
  assign n978 = ~n975 & n977;
  assign po61 = ~n971 & n978;
  assign n980 = pi82 & ~n544;
  assign n981 = ~pi48 & n847;
  assign n982 = pi82 & ~n981;
  assign n983 = n376 & ~n982;
  assign n984 = ~n980 & ~n983;
  assign n985 = ~pi47 & ~n984;
  assign n986 = pi47 & n861;
  assign n987 = n555 & n986;
  assign n988 = ~pi129 & ~n987;
  assign n989 = n544 & n981;
  assign n990 = pi82 & ~n989;
  assign n991 = ~n376 & ~n990;
  assign n992 = pi64 & n991;
  assign n993 = n988 & ~n992;
  assign po62 = ~n985 & n993;
  assign n995 = pi82 & ~n847;
  assign n996 = n376 & ~n995;
  assign n997 = pi82 & ~n597;
  assign n998 = ~n996 & ~n997;
  assign n999 = ~pi48 & ~n998;
  assign n1000 = n597 & n847;
  assign n1001 = pi82 & ~n1000;
  assign n1002 = ~n376 & ~n1001;
  assign n1003 = pi62 & n1002;
  assign n1004 = pi48 & n958;
  assign n1005 = n382 & n1004;
  assign n1006 = n962 & n1005;
  assign n1007 = ~pi129 & ~n1006;
  assign n1008 = ~n1003 & n1007;
  assign po63 = ~n999 & n1008;
  assign n1010 = n381 & n596;
  assign n1011 = n384 & n1010;
  assign n1012 = pi49 & ~n1011;
  assign n1013 = n389 & ~n946;
  assign n1014 = n535 & n1013;
  assign n1015 = n597 & n1014;
  assign n1016 = ~n1012 & ~n1015;
  assign n1017 = pi82 & ~n1016;
  assign n1018 = pi49 & n377;
  assign n1019 = ~n1017 & ~n1018;
  assign n1020 = pi82 & ~n538;
  assign n1021 = ~pi69 & ~n1020;
  assign n1022 = ~n376 & n1021;
  assign n1023 = n1019 & ~n1022;
  assign po64 = ~pi129 & ~n1023;
  assign n1025 = n378 & n379;
  assign n1026 = pi82 & ~n1025;
  assign n1027 = n554 & n923;
  assign n1028 = pi82 & ~n1027;
  assign n1029 = n376 & ~n1028;
  assign n1030 = ~n1026 & ~n1029;
  assign n1031 = ~pi50 & ~n1030;
  assign n1032 = n914 & n1025;
  assign n1033 = pi82 & ~n1032;
  assign n1034 = ~n376 & ~n1033;
  assign n1035 = pi66 & n1034;
  assign n1036 = pi50 & n962;
  assign n1037 = ~pi129 & ~n1036;
  assign n1038 = ~n1035 & n1037;
  assign po65 = ~n1031 & n1038;
  assign n1040 = pi51 & ~pi109;
  assign n1041 = ~pi106 & ~n868;
  assign n1042 = ~n1040 & n1041;
  assign po66 = ~pi129 & ~n1042;
  assign n1044 = pi52 & ~n868;
  assign n1045 = ~pi106 & ~n866;
  assign n1046 = ~n1044 & n1045;
  assign po67 = ~pi129 & ~n1046;
  assign n1048 = ~pi116 & n772;
  assign n1049 = pi58 & ~pi116;
  assign n1050 = n650 & n658;
  assign n1051 = ~pi58 & ~n1050;
  assign n1052 = pi97 & ~n1051;
  assign n1053 = ~pi53 & n1052;
  assign n1054 = ~n1049 & n1053;
  assign n1055 = ~n1048 & ~n1054;
  assign n1056 = n337 & ~n1055;
  assign n1057 = ~pi85 & n1056;
  assign po68 = n744 & n1057;
  assign n1059 = ~pi47 & n989;
  assign n1060 = pi82 & ~n1059;
  assign n1061 = ~n376 & ~n1060;
  assign po69 = pi129 | n1061;
  assign po129 = pi123 | pi129;
  assign n1064 = pi114 & ~pi122;
  assign po70 = ~po129 & n1064;
  assign n1066 = pi26 & pi58;
  assign n1067 = ~pi58 & ~n662;
  assign n1068 = pi94 & ~n1067;
  assign n1069 = ~n1066 & n1068;
  assign n1070 = pi37 & ~pi116;
  assign n1071 = ~pi58 & ~n1070;
  assign n1072 = ~n662 & ~n1071;
  assign n1073 = ~n1049 & n1072;
  assign n1074 = ~n1069 & ~n1073;
  assign n1075 = ~pi53 & ~n1074;
  assign n1076 = ~pi26 & pi37;
  assign n1077 = ~pi58 & n1076;
  assign n1078 = ~n1075 & ~n1077;
  assign n1079 = ~pi85 & ~n1078;
  assign n1080 = n709 & n1076;
  assign n1081 = ~n1079 & ~n1080;
  assign n1082 = ~pi27 & ~n1081;
  assign n1083 = n784 & n1076;
  assign n1084 = ~n1082 & ~n1083;
  assign po71 = n337 & ~n1084;
  assign n1086 = ~pi26 & ~pi53;
  assign n1087 = ~pi85 & n1086;
  assign n1088 = ~pi116 & n1087;
  assign n1089 = pi26 & pi53;
  assign n1090 = pi85 & ~n1086;
  assign n1091 = ~pi58 & ~n1090;
  assign n1092 = ~n1089 & n1091;
  assign n1093 = ~n1088 & ~n1092;
  assign n1094 = pi57 & ~n1093;
  assign n1095 = pi60 & n755;
  assign n1096 = pi116 & n1095;
  assign n1097 = ~n1094 & ~n1096;
  assign n1098 = ~pi27 & ~n1097;
  assign n1099 = pi57 & ~pi58;
  assign n1100 = n1087 & n1099;
  assign n1101 = ~n1098 & ~n1100;
  assign po72 = n337 & ~n1101;
  assign n1103 = n744 & n1049;
  assign n1104 = ~pi58 & ~n733;
  assign n1105 = n673 & n1104;
  assign n1106 = ~n1103 & ~n1105;
  assign n1107 = ~pi53 & ~n1106;
  assign n1108 = ~pi85 & n337;
  assign po73 = n1107 & n1108;
  assign n1110 = ~n690 & ~n772;
  assign n1111 = ~pi116 & ~n1110;
  assign n1112 = ~n660 & n709;
  assign n1113 = ~n1111 & ~n1112;
  assign n1114 = pi59 & ~n1113;
  assign n1115 = pi96 & n709;
  assign n1116 = n660 & n1115;
  assign n1117 = ~n1114 & ~n1116;
  assign n1118 = ~pi85 & ~n1117;
  assign n1119 = pi59 & n648;
  assign n1120 = n709 & n1119;
  assign n1121 = ~n1118 & ~n1120;
  assign n1122 = ~pi27 & ~n1121;
  assign n1123 = pi59 & ~pi116;
  assign n1124 = pi27 & n784;
  assign n1125 = n1123 & n1124;
  assign n1126 = ~n1122 & ~n1125;
  assign n1127 = ~pi26 & ~n1126;
  assign n1128 = n785 & n1123;
  assign n1129 = ~n1127 & ~n1128;
  assign po74 = n337 & ~n1129;
  assign n1131 = ~pi117 & ~pi122;
  assign n1132 = pi60 & ~n1131;
  assign n1133 = pi123 & n1131;
  assign po75 = n1132 | n1133;
  assign n1135 = ~pi114 & ~pi129;
  assign n1136 = ~pi122 & pi123;
  assign po76 = n1135 & n1136;
  assign n1138 = pi136 & ~pi137;
  assign n1139 = pi132 & pi133;
  assign n1140 = pi131 & n1139;
  assign n1141 = ~pi138 & n1140;
  assign n1142 = n1138 & n1141;
  assign n1143 = ~pi62 & ~n1142;
  assign n1144 = pi140 & n1142;
  assign n1145 = ~pi129 & ~n1144;
  assign po77 = n1143 | ~n1145;
  assign n1147 = ~pi63 & ~n1142;
  assign n1148 = pi142 & n1142;
  assign n1149 = ~pi129 & ~n1148;
  assign po78 = n1147 | ~n1149;
  assign n1151 = ~pi64 & ~n1142;
  assign n1152 = pi139 & n1142;
  assign n1153 = ~pi129 & ~n1152;
  assign po79 = n1151 | ~n1153;
  assign n1155 = ~pi65 & ~n1142;
  assign n1156 = pi146 & n1142;
  assign n1157 = ~pi129 & ~n1156;
  assign po80 = n1155 | ~n1157;
  assign n1159 = ~pi136 & n1141;
  assign n1160 = ~pi137 & n1159;
  assign n1161 = ~pi66 & ~n1160;
  assign n1162 = pi143 & n1160;
  assign n1163 = ~pi129 & ~n1162;
  assign po81 = n1161 | ~n1163;
  assign n1165 = ~pi67 & ~n1160;
  assign n1166 = pi139 & n1160;
  assign n1167 = ~pi129 & ~n1166;
  assign po82 = n1165 | ~n1167;
  assign n1169 = ~pi68 & ~n1142;
  assign n1170 = pi141 & n1142;
  assign n1171 = ~pi129 & ~n1170;
  assign po83 = n1169 | ~n1171;
  assign n1173 = ~pi69 & ~n1142;
  assign n1174 = pi143 & n1142;
  assign n1175 = ~pi129 & ~n1174;
  assign po84 = n1173 | ~n1175;
  assign n1177 = ~pi70 & ~n1142;
  assign n1178 = pi144 & n1142;
  assign n1179 = ~pi129 & ~n1178;
  assign po85 = n1177 | ~n1179;
  assign n1181 = ~pi71 & ~n1142;
  assign n1182 = pi145 & n1142;
  assign n1183 = ~pi129 & ~n1182;
  assign po86 = n1181 | ~n1183;
  assign n1185 = ~pi72 & ~n1160;
  assign n1186 = pi140 & n1160;
  assign n1187 = ~pi129 & ~n1186;
  assign po87 = n1185 | ~n1187;
  assign n1189 = ~pi73 & ~n1160;
  assign n1190 = pi141 & n1160;
  assign n1191 = ~pi129 & ~n1190;
  assign po88 = n1189 | ~n1191;
  assign n1193 = ~pi74 & ~n1160;
  assign n1194 = pi142 & n1160;
  assign n1195 = ~pi129 & ~n1194;
  assign po89 = n1193 | ~n1195;
  assign n1197 = ~pi75 & ~n1160;
  assign n1198 = pi144 & n1160;
  assign n1199 = ~pi129 & ~n1198;
  assign po90 = n1197 | ~n1199;
  assign n1201 = ~pi76 & ~n1160;
  assign n1202 = pi145 & n1160;
  assign n1203 = ~pi129 & ~n1202;
  assign po91 = n1201 | ~n1203;
  assign n1205 = ~pi77 & ~n1160;
  assign n1206 = pi146 & n1160;
  assign n1207 = ~pi129 & ~n1206;
  assign po92 = n1205 | ~n1207;
  assign n1209 = ~pi136 & pi137;
  assign n1210 = n1141 & n1209;
  assign n1211 = ~pi78 & ~n1210;
  assign n1212 = ~pi142 & n1210;
  assign n1213 = ~pi129 & ~n1212;
  assign po93 = ~n1211 & n1213;
  assign n1215 = ~pi79 & ~n1210;
  assign n1216 = ~pi143 & n1210;
  assign n1217 = ~pi129 & ~n1216;
  assign po94 = ~n1215 & n1217;
  assign n1219 = ~pi80 & ~n1210;
  assign n1220 = ~pi144 & n1210;
  assign n1221 = ~pi129 & ~n1220;
  assign po95 = ~n1219 & n1221;
  assign n1223 = ~pi81 & ~n1210;
  assign n1224 = ~pi145 & n1210;
  assign n1225 = ~pi129 & ~n1224;
  assign po96 = ~n1223 & n1225;
  assign n1227 = ~pi82 & ~n1210;
  assign n1228 = ~pi146 & n1210;
  assign n1229 = ~pi129 & ~n1228;
  assign po97 = ~n1227 & n1229;
  assign n1231 = ~pi89 & pi138;
  assign n1232 = pi62 & ~pi138;
  assign n1233 = pi136 & ~n1232;
  assign n1234 = ~n1231 & n1233;
  assign n1235 = ~pi119 & pi138;
  assign n1236 = pi72 & ~pi138;
  assign n1237 = ~pi136 & ~n1236;
  assign n1238 = ~n1235 & n1237;
  assign n1239 = ~n1234 & ~n1238;
  assign n1240 = ~pi137 & ~n1239;
  assign n1241 = pi136 & ~pi138;
  assign n1242 = pi31 & n1241;
  assign n1243 = ~pi87 & ~pi138;
  assign n1244 = pi115 & pi138;
  assign n1245 = ~pi136 & ~n1244;
  assign n1246 = ~n1243 & n1245;
  assign n1247 = ~n1242 & ~n1246;
  assign n1248 = pi137 & ~n1247;
  assign po98 = n1240 | n1248;
  assign n1250 = ~pi84 & ~n1210;
  assign n1251 = ~pi141 & n1210;
  assign n1252 = ~pi129 & ~n1251;
  assign po99 = ~n1250 & n1252;
  assign n1254 = ~pi85 & n660;
  assign n1255 = pi96 & n1254;
  assign n1256 = ~n648 & ~n1255;
  assign n1257 = n337 & ~n1256;
  assign n1258 = ~pi27 & n1257;
  assign po100 = n710 & n1258;
  assign n1260 = ~pi86 & ~n1210;
  assign n1261 = ~pi139 & n1210;
  assign n1262 = ~pi129 & ~n1261;
  assign po101 = ~n1260 & n1262;
  assign n1264 = ~pi87 & ~n1210;
  assign n1265 = ~pi140 & n1210;
  assign n1266 = ~pi129 & ~n1265;
  assign po102 = ~n1264 & n1266;
  assign n1268 = pi137 & n1241;
  assign n1269 = n1140 & n1268;
  assign n1270 = ~pi88 & ~n1269;
  assign n1271 = ~pi139 & n1269;
  assign n1272 = ~pi129 & ~n1271;
  assign po103 = ~n1270 & n1272;
  assign n1274 = ~pi89 & ~n1269;
  assign n1275 = ~pi140 & n1269;
  assign n1276 = ~pi129 & ~n1275;
  assign po104 = ~n1274 & n1276;
  assign n1278 = ~pi90 & ~n1269;
  assign n1279 = ~pi142 & n1269;
  assign n1280 = ~pi129 & ~n1279;
  assign po105 = ~n1278 & n1280;
  assign n1282 = ~pi91 & ~n1269;
  assign n1283 = ~pi143 & n1269;
  assign n1284 = ~pi129 & ~n1283;
  assign po106 = ~n1282 & n1284;
  assign n1286 = ~pi92 & ~n1269;
  assign n1287 = ~pi144 & n1269;
  assign n1288 = ~pi129 & ~n1287;
  assign po107 = ~n1286 & n1288;
  assign n1290 = ~pi93 & ~n1269;
  assign n1291 = ~pi146 & n1269;
  assign n1292 = ~pi129 & ~n1291;
  assign po108 = ~n1290 & n1292;
  assign n1294 = ~pi137 & pi138;
  assign n1295 = pi82 & ~pi136;
  assign n1296 = n1294 & n1295;
  assign n1297 = n1140 & n1296;
  assign n1298 = ~pi94 & ~n1297;
  assign n1299 = ~pi142 & n1297;
  assign n1300 = ~pi129 & ~n1299;
  assign po109 = ~n1298 & n1300;
  assign n1302 = ~pi3 & ~pi110;
  assign n1303 = ~n1140 & ~n1302;
  assign n1304 = ~n1297 & ~n1303;
  assign n1305 = pi95 & n1304;
  assign n1306 = pi143 & n1297;
  assign n1307 = ~n1305 & ~n1306;
  assign po110 = ~pi129 & ~n1307;
  assign n1309 = pi96 & n1304;
  assign n1310 = pi146 & n1297;
  assign n1311 = ~n1309 & ~n1310;
  assign po111 = ~pi129 & ~n1311;
  assign n1313 = pi97 & n1304;
  assign n1314 = pi145 & n1297;
  assign n1315 = ~n1313 & ~n1314;
  assign po112 = ~pi129 & ~n1315;
  assign n1317 = ~pi98 & ~n1269;
  assign n1318 = ~pi145 & n1269;
  assign n1319 = ~pi129 & ~n1318;
  assign po113 = ~n1317 & n1319;
  assign n1321 = ~pi99 & ~n1269;
  assign n1322 = ~pi141 & n1269;
  assign n1323 = ~pi129 & ~n1322;
  assign po114 = ~n1321 & n1323;
  assign n1325 = pi100 & n1304;
  assign n1326 = pi144 & n1297;
  assign n1327 = ~n1325 & ~n1326;
  assign po115 = ~pi129 & ~n1327;
  assign n1329 = ~pi124 & pi138;
  assign n1330 = pi77 & ~pi138;
  assign n1331 = ~pi136 & ~n1330;
  assign n1332 = ~n1329 & n1331;
  assign n1333 = ~pi93 & pi138;
  assign n1334 = pi65 & ~pi138;
  assign n1335 = pi136 & ~n1334;
  assign n1336 = ~n1333 & n1335;
  assign n1337 = ~n1332 & ~n1336;
  assign n1338 = ~pi137 & ~n1337;
  assign n1339 = pi37 & n1241;
  assign n1340 = ~pi82 & ~pi138;
  assign n1341 = ~pi96 & pi138;
  assign n1342 = ~pi136 & ~n1341;
  assign n1343 = ~n1340 & n1342;
  assign n1344 = ~n1339 & ~n1343;
  assign n1345 = pi137 & ~n1344;
  assign po116 = n1338 | n1345;
  assign n1347 = pi91 & n1138;
  assign n1348 = pi95 & n1209;
  assign n1349 = ~n1347 & ~n1348;
  assign n1350 = pi138 & ~n1349;
  assign n1351 = ~pi79 & ~pi136;
  assign n1352 = ~pi34 & pi136;
  assign n1353 = pi137 & ~n1352;
  assign n1354 = ~n1351 & n1353;
  assign n1355 = pi66 & ~pi136;
  assign n1356 = pi69 & pi136;
  assign n1357 = ~pi137 & ~n1356;
  assign n1358 = ~n1355 & n1357;
  assign n1359 = ~n1354 & ~n1358;
  assign n1360 = ~pi138 & ~n1359;
  assign po117 = n1350 | n1360;
  assign n1362 = pi90 & n1138;
  assign n1363 = pi94 & n1209;
  assign n1364 = ~n1362 & ~n1363;
  assign n1365 = pi138 & ~n1364;
  assign n1366 = ~pi78 & ~pi136;
  assign n1367 = ~pi33 & pi136;
  assign n1368 = pi137 & ~n1367;
  assign n1369 = ~n1366 & n1368;
  assign n1370 = pi74 & ~pi136;
  assign n1371 = pi63 & pi136;
  assign n1372 = ~pi137 & ~n1371;
  assign n1373 = ~n1370 & n1372;
  assign n1374 = ~n1369 & ~n1373;
  assign n1375 = ~pi138 & ~n1374;
  assign po118 = n1365 | n1375;
  assign n1377 = pi99 & n1138;
  assign n1378 = ~pi112 & n1209;
  assign n1379 = ~n1377 & ~n1378;
  assign n1380 = pi138 & ~n1379;
  assign n1381 = pi73 & ~pi136;
  assign n1382 = pi68 & pi136;
  assign n1383 = ~pi137 & ~n1382;
  assign n1384 = ~n1381 & n1383;
  assign n1385 = ~pi84 & ~pi136;
  assign n1386 = ~pi32 & pi136;
  assign n1387 = pi137 & ~n1386;
  assign n1388 = ~n1385 & n1387;
  assign n1389 = ~n1384 & ~n1388;
  assign n1390 = ~pi138 & ~n1389;
  assign po119 = n1380 | n1390;
  assign n1392 = ~pi92 & pi138;
  assign n1393 = pi70 & ~pi138;
  assign n1394 = pi136 & ~n1393;
  assign n1395 = ~n1392 & n1394;
  assign n1396 = ~pi125 & pi138;
  assign n1397 = pi75 & ~pi138;
  assign n1398 = ~pi136 & ~n1397;
  assign n1399 = ~n1396 & n1398;
  assign n1400 = ~n1395 & ~n1399;
  assign n1401 = ~pi137 & ~n1400;
  assign n1402 = pi35 & n1241;
  assign n1403 = ~pi80 & ~pi138;
  assign n1404 = ~pi100 & pi138;
  assign n1405 = ~pi136 & ~n1404;
  assign n1406 = ~n1403 & n1405;
  assign n1407 = ~n1402 & ~n1406;
  assign n1408 = pi137 & ~n1407;
  assign po120 = n1401 | n1408;
  assign n1410 = ~pi27 & n1254;
  assign n1411 = n710 & n1410;
  assign n1412 = ~n697 & ~n1411;
  assign po121 = n337 & ~n1412;
  assign n1414 = ~pi98 & pi138;
  assign n1415 = pi71 & ~pi138;
  assign n1416 = pi136 & ~n1415;
  assign n1417 = ~n1414 & n1416;
  assign n1418 = ~pi23 & pi138;
  assign n1419 = pi76 & ~pi138;
  assign n1420 = ~pi136 & ~n1419;
  assign n1421 = ~n1418 & n1420;
  assign n1422 = ~n1417 & ~n1421;
  assign n1423 = ~pi137 & ~n1422;
  assign n1424 = pi36 & n1241;
  assign n1425 = ~pi81 & ~pi138;
  assign n1426 = ~pi97 & pi138;
  assign n1427 = ~pi136 & ~n1426;
  assign n1428 = ~n1425 & n1427;
  assign n1429 = ~n1424 & ~n1428;
  assign n1430 = pi137 & ~n1429;
  assign po122 = n1423 | n1430;
  assign n1432 = ~pi88 & pi138;
  assign n1433 = pi64 & ~pi138;
  assign n1434 = pi136 & ~n1433;
  assign n1435 = ~n1432 & n1434;
  assign n1436 = ~pi120 & pi138;
  assign n1437 = pi67 & ~pi138;
  assign n1438 = ~pi136 & ~n1437;
  assign n1439 = ~n1436 & n1438;
  assign n1440 = ~n1435 & ~n1439;
  assign n1441 = ~pi137 & ~n1440;
  assign n1442 = pi30 & n1241;
  assign n1443 = ~pi86 & ~pi138;
  assign n1444 = ~pi111 & pi138;
  assign n1445 = ~pi136 & ~n1444;
  assign n1446 = ~n1443 & n1445;
  assign n1447 = ~n1442 & ~n1446;
  assign n1448 = pi137 & ~n1447;
  assign po123 = n1441 | n1448;
  assign n1450 = ~pi26 & n665;
  assign n1451 = pi116 & ~n1450;
  assign n1452 = n337 & ~n733;
  assign po124 = n1451 & n1452;
  assign n1454 = ~pi97 & n690;
  assign n1455 = ~n772 & ~n1454;
  assign n1456 = pi116 & n337;
  assign po125 = ~n1455 & n1456;
  assign n1458 = ~pi111 & ~n1296;
  assign n1459 = n1140 & ~n1458;
  assign n1460 = ~pi139 & n1296;
  assign n1461 = ~pi129 & ~n1460;
  assign po126 = n1459 & n1461;
  assign n1463 = pi112 & ~n1296;
  assign n1464 = ~pi141 & n1296;
  assign n1465 = n1140 & ~n1464;
  assign n1466 = ~pi129 & n1465;
  assign po127 = ~n1463 & n1466;
  assign n1468 = ~pi11 & pi54;
  assign n1469 = ~pi22 & n1468;
  assign n1470 = ~pi54 & pi113;
  assign n1471 = n337 & ~n1470;
  assign po128 = ~n1469 & n1471;
  assign n1473 = pi115 & ~n1296;
  assign n1474 = ~pi140 & n1296;
  assign n1475 = n1140 & ~n1474;
  assign n1476 = ~pi129 & n1475;
  assign po130 = ~n1473 & n1476;
  assign n1478 = pi54 & n337;
  assign n1479 = ~pi4 & n438;
  assign n1480 = ~pi9 & n1479;
  assign po131 = n1478 & ~n1480;
  assign po132 = ~pi122 | pi129;
  assign n1483 = ~pi54 & pi118;
  assign n1484 = pi54 & ~pi59;
  assign n1485 = n518 & n1484;
  assign n1486 = ~n1483 & ~n1485;
  assign po133 = ~pi129 & ~n1486;
  assign po134 = ~pi129 & ~n658;
  assign n1489 = ~pi120 & n1302;
  assign n1490 = ~pi111 & ~n1489;
  assign po135 = ~pi129 & n1490;
  assign n1492 = pi81 & pi120;
  assign po136 = ~pi129 & n1492;
  assign po137 = pi129 | pi134;
  assign po138 = pi129 | pi135;
  assign po139 = pi57 & ~pi129;
  assign n1497 = ~pi96 & pi125;
  assign n1498 = ~pi3 & ~n1497;
  assign po140 = ~pi129 & ~n1498;
  assign n1500 = ~pi126 & pi132;
  assign po141 = pi133 & n1500;
  assign po12 = 1'b1;
  assign po0 = pi108;
  assign po1 = pi83;
  assign po2 = pi104;
  assign po3 = pi103;
  assign po4 = pi102;
  assign po5 = pi105;
  assign po6 = pi107;
  assign po7 = pi101;
  assign po8 = pi126;
  assign po9 = pi121;
  assign po10 = pi1;
  assign po11 = pi0;
  assign po13 = pi130;
  assign po14 = pi128;
endmodule
