module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 ,
    pi5 , pi6 , pi7 , pi8 , pi9 ,
    pi10 , pi11 , pi12 , pi13 , pi14 ,
    pi15 , pi16 , pi17 , pi18 , pi19 ,
    pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 ,
    pi30 , pi31 , pi32 , pi33 , pi34 ,
    pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 ,
    pi45 , pi46 , pi47 , pi48 , pi49 ,
    pi50 , pi51 , pi52 , pi53 , pi54 ,
    pi55 , pi56 , pi57 , pi58 , pi59 ,
    po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 ,
    po14 , po15 , po16 , po17 ,
    po18 , po19 , po20 , po21 ,
    po22 , po23 , po24 , po25 ,
    po26 , po27 , po28 , po29   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 ,
    pi5 , pi6 , pi7 , pi8 , pi9 ,
    pi10 , pi11 , pi12 , pi13 , pi14 ,
    pi15 , pi16 , pi17 , pi18 , pi19 ,
    pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 ,
    pi30 , pi31 , pi32 , pi33 , pi34 ,
    pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 ,
    pi45 , pi46 , pi47 , pi48 , pi49 ,
    pi50 , pi51 , pi52 , pi53 , pi54 ,
    pi55 , pi56 , pi57 , pi58 , pi59 ;
  output po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 ,
    po14 , po15 , po16 , po17 ,
    po18 , po19 , po20 , po21 ,
    po22 , po23 , po24 , po25 ,
    po26 , po27 , po28 , po29 ;
  wire n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105,
    n106, n107, n108, n109, n110, n111, n112,
    n113, n114, n115, n116, n117, n118, n119,
    n120, n121, n122, n123, n124, n125, n126,
    n127, n128, n129, n130, n131, n132, n133,
    n134, n135, n136, n137, n138, n139, n140,
    n141, n142, n143, n144, n145, n146, n147,
    n148, n149, n150, n151, n152, n153, n154,
    n155, n156, n157, n158, n159, n160, n161,
    n162, n163, n164, n165, n166, n167, n168,
    n169, n170, n171, n172, n173, n174, n175,
    n176, n177, n178, n179, n180, n181, n182,
    n183, n184, n185, n186, n187, n188, n189,
    n190, n191, n192, n193, n194, n195, n196,
    n197, n198, n199, n200, n201, n202, n203,
    n204, n205, n206, n207, n209, n210, n211,
    n212, n213, n214, n215, n216, n217, n218,
    n219, n220, n221, n222, n223, n224, n225,
    n226, n227, n228, n229, n230, n231, n232,
    n233, n234, n235, n236, n237, n238, n239,
    n240, n241, n242, n243, n244, n245, n246,
    n247, n248, n249, n250, n251, n252, n253,
    n254, n255, n256, n257, n258, n259, n260,
    n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274,
    n275, n276, n277, n278, n279, n280, n281,
    n282, n283, n284, n285, n286, n287, n288,
    n289, n290, n291, n292, n293, n294, n295,
    n296, n297, n298, n299, n300, n301, n302,
    n303, n304, n305, n306, n307, n308, n309,
    n310, n311, n312, n313, n314, n315, n316,
    n317, n318, n319, n320, n321, n322, n323,
    n324, n325, n326, n327, n328, n329, n330,
    n331, n332, n334, n335, n336;
  assign n92 = ~pi9  & ~pi10 ;
  assign n93 = pi11  & ~n92;
  assign n94 = ~pi12  & ~n93;
  assign n95 = pi12  & n93;
  assign n96 = ~n94 & ~n95;
  assign n97 = pi6  & ~n96;
  assign n98 = pi4  & n97;
  assign n99 = ~pi11  & n92;
  assign n100 = ~n93 & ~n99;
  assign n101 = ~pi13  & n94;
  assign n102 = pi13  & ~n94;
  assign n103 = ~n101 & ~n102;
  assign n104 = pi14  & ~n101;
  assign n105 = pi15  & n104;
  assign n106 = ~pi16  & ~n105;
  assign n107 = pi16  & n105;
  assign n108 = ~n106 & ~n107;
  assign n109 = pi17  & ~n106;
  assign n110 = ~pi17  & n106;
  assign n111 = ~n109 & ~n110;
  assign n112 = ~n108 & n111;
  assign n113 = ~pi18  & n112;
  assign n114 = ~n103 & n113;
  assign n115 = ~pi14  & n101;
  assign n116 = ~n104 & ~n115;
  assign n117 = pi15  & ~n104;
  assign n118 = ~pi15  & n104;
  assign n119 = ~n117 & ~n118;
  assign n120 = ~pi18  & ~n109;
  assign n121 = pi19  & ~n120;
  assign n122 = ~pi19  & n120;
  assign n123 = ~n121 & ~n122;
  assign n124 = pi20  & ~n121;
  assign n125 = ~pi20  & n121;
  assign n126 = ~n124 & ~n125;
  assign n127 = n123 & ~n126;
  assign n128 = pi20  & n121;
  assign n129 = ~pi21  & ~n128;
  assign n130 = ~pi22  & n129;
  assign n131 = pi22  & ~n129;
  assign n132 = ~n130 & ~n131;
  assign n133 = pi21  & n128;
  assign n134 = ~n129 & ~n133;
  assign n135 = ~pi9  & pi29 ;
  assign n136 = ~n134 & n135;
  assign n137 = ~n132 & n136;
  assign n138 = pi23  & ~n130;
  assign n139 = ~pi23  & n130;
  assign n140 = ~n138 & ~n139;
  assign n141 = pi24  & ~n138;
  assign n142 = ~pi24  & n138;
  assign n143 = ~n141 & ~n142;
  assign n144 = pi24  & n138;
  assign n145 = pi25  & ~n144;
  assign n146 = ~pi25  & n144;
  assign n147 = ~n145 & ~n146;
  assign n148 = pi25  & n144;
  assign n149 = ~pi26  & ~n148;
  assign n150 = pi27  & ~n149;
  assign n151 = ~pi27  & n149;
  assign n152 = ~n150 & ~n151;
  assign n153 = pi26  & n148;
  assign n154 = ~n149 & ~n153;
  assign n155 = pi28  & ~n154;
  assign n156 = n152 & n155;
  assign n157 = ~n147 & n156;
  assign n158 = ~n143 & n157;
  assign n159 = n140 & n158;
  assign n160 = n137 & n159;
  assign n161 = n127 & n160;
  assign n162 = ~n119 & n161;
  assign n163 = n116 & n162;
  assign n164 = n114 & n163;
  assign n165 = n100 & n164;
  assign n166 = pi2  & n165;
  assign n167 = n98 & n166;
  assign n168 = pi9  & pi10 ;
  assign n169 = ~n92 & ~n168;
  assign n170 = pi3  & ~n169;
  assign n171 = pi1  & n170;
  assign n172 = pi7  & pi8 ;
  assign n173 = pi5  & n172;
  assign n174 = pi0  & n173;
  assign n175 = n171 & n174;
  assign n176 = n167 & n175;
  assign n177 = pi28  & n150;
  assign n178 = pi29  & n177;
  assign n179 = ~n176 & ~n178;
  assign n180 = pi27  & n154;
  assign n181 = pi18  & n109;
  assign n182 = n121 & ~n181;
  assign n183 = n143 & n182;
  assign n184 = n132 & n183;
  assign n185 = ~pi1  & ~pi8 ;
  assign n186 = ~pi6  & n185;
  assign n187 = n96 & n186;
  assign n188 = ~n100 & n187;
  assign n189 = n119 & n188;
  assign n190 = pi14  & n189;
  assign n191 = n108 & n190;
  assign n192 = n126 & n191;
  assign n193 = ~pi2  & ~pi3 ;
  assign n194 = ~pi7  & n193;
  assign n195 = ~pi5  & n194;
  assign n196 = ~pi4  & n195;
  assign n197 = n169 & n196;
  assign n198 = n103 & n197;
  assign n199 = pi17  & n198;
  assign n200 = n134 & n199;
  assign n201 = n192 & n200;
  assign n202 = n147 & n201;
  assign n203 = pi23  & n202;
  assign n204 = pi9  & n203;
  assign n205 = n184 & n204;
  assign n206 = n180 & n205;
  assign n207 = n178 & ~n206;
  assign po0  = n179 | n207;
  assign n209 = ~pi39  & ~pi40 ;
  assign n210 = pi39  & pi40 ;
  assign n211 = ~n209 & ~n210;
  assign n212 = pi37  & pi38 ;
  assign n213 = pi35  & n212;
  assign n214 = pi41  & ~n209;
  assign n215 = ~pi41  & n209;
  assign n216 = ~n214 & ~n215;
  assign n217 = ~pi42  & ~n214;
  assign n218 = ~pi43  & n217;
  assign n219 = pi44  & ~n218;
  assign n220 = pi43  & ~n217;
  assign n221 = ~n218 & ~n220;
  assign n222 = ~n219 & ~n221;
  assign n223 = ~pi44  & n218;
  assign n224 = pi45  & n219;
  assign n225 = ~pi46  & ~n224;
  assign n226 = pi47  & ~n225;
  assign n227 = ~pi48  & ~n226;
  assign n228 = pi46  & n224;
  assign n229 = ~pi47  & ~n228;
  assign n230 = n227 & ~n229;
  assign n231 = pi45  & ~n219;
  assign n232 = ~pi45  & n219;
  assign n233 = ~n231 & ~n232;
  assign n234 = pi49  & ~n227;
  assign n235 = pi50  & n234;
  assign n236 = ~pi51  & ~n235;
  assign n237 = ~pi52  & n236;
  assign n238 = pi52  & ~n236;
  assign n239 = ~n237 & ~n238;
  assign n240 = ~pi49  & n227;
  assign n241 = ~n234 & ~n240;
  assign n242 = ~n239 & n241;
  assign n243 = pi53  & ~n237;
  assign n244 = pi50  & ~n234;
  assign n245 = ~pi50  & n234;
  assign n246 = ~n244 & ~n245;
  assign n247 = ~pi53  & n237;
  assign n248 = pi51  & n235;
  assign n249 = ~n236 & ~n248;
  assign n250 = pi54  & n243;
  assign n251 = pi55  & ~n250;
  assign n252 = ~pi55  & n250;
  assign n253 = ~n251 & ~n252;
  assign n254 = pi59  & ~n253;
  assign n255 = ~n249 & n254;
  assign n256 = pi55  & n250;
  assign n257 = ~pi56  & ~n256;
  assign n258 = pi56  & n256;
  assign n259 = ~n257 & ~n258;
  assign n260 = pi54  & ~n243;
  assign n261 = ~pi54  & n243;
  assign n262 = ~n260 & ~n261;
  assign n263 = pi57  & ~n257;
  assign n264 = pi58  & ~n263;
  assign n265 = ~pi57  & n257;
  assign n266 = pi30  & ~pi39 ;
  assign n267 = ~n265 & n266;
  assign n268 = n264 & n267;
  assign n269 = ~n262 & n268;
  assign n270 = ~n259 & n269;
  assign n271 = n255 & n270;
  assign n272 = ~n247 & n271;
  assign n273 = ~n246 & n272;
  assign n274 = ~n243 & n273;
  assign n275 = n242 & n274;
  assign n276 = ~n233 & n275;
  assign n277 = n230 & n276;
  assign n278 = ~n223 & n277;
  assign n279 = n222 & n278;
  assign n280 = n216 & n279;
  assign n281 = pi32  & n280;
  assign n282 = pi42  & n214;
  assign n283 = ~n217 & ~n282;
  assign n284 = pi36  & ~n283;
  assign n285 = pi34  & n284;
  assign n286 = pi31  & n285;
  assign n287 = n281 & n286;
  assign n288 = n213 & n287;
  assign n289 = ~n211 & n288;
  assign n290 = pi33  & n289;
  assign n291 = ~pi0  & ~pi30 ;
  assign n292 = pi58  & n263;
  assign n293 = pi59  & n292;
  assign n294 = ~n291 & n293;
  assign n295 = ~n225 & ~n228;
  assign n296 = ~pi31  & ~pi38 ;
  assign n297 = ~pi36  & n296;
  assign n298 = n283 & n297;
  assign n299 = ~n216 & n298;
  assign n300 = n233 & n299;
  assign n301 = pi44  & n300;
  assign n302 = n295 & n301;
  assign n303 = n249 & n302;
  assign n304 = pi49  & n303;
  assign n305 = n262 & n304;
  assign n306 = n239 & n305;
  assign n307 = pi39  & n306;
  assign n308 = ~pi58  & n263;
  assign n309 = ~n264 & ~n308;
  assign n310 = pi48  & n226;
  assign n311 = ~n227 & ~n310;
  assign n312 = ~pi32  & ~pi33 ;
  assign n313 = ~pi37  & n312;
  assign n314 = ~pi35  & n313;
  assign n315 = ~pi34  & n314;
  assign n316 = n211 & n315;
  assign n317 = n221 & n316;
  assign n318 = pi47  & n317;
  assign n319 = n246 & n318;
  assign n320 = n311 & n319;
  assign n321 = n253 & n320;
  assign n322 = pi53  & n321;
  assign n323 = n309 & n322;
  assign n324 = pi57  & n323;
  assign n325 = n259 & n324;
  assign n326 = n307 & n325;
  assign n327 = n293 & ~n326;
  assign n328 = ~n294 & ~n327;
  assign n329 = ~n290 & n328;
  assign n330 = pi0  & ~n293;
  assign n331 = ~n179 & ~n330;
  assign n332 = ~n329 & n331;
  assign po1  = ~n207 & ~n332;
  assign n334 = pi0  & n293;
  assign n335 = pi30  & n334;
  assign n336 = ~n327 & ~n335;
  assign po2  = ~po0  & ~n336;
  assign po3  = 1'b0;
  assign po4  = 1'b0;
  assign po5  = 1'b0;
  assign po6  = 1'b0;
  assign po7  = 1'b0;
  assign po8  = 1'b0;
  assign po9  = 1'b0;
  assign po10  = 1'b0;
  assign po11  = 1'b0;
  assign po12  = 1'b0;
  assign po13  = 1'b0;
  assign po14  = 1'b0;
  assign po15  = 1'b0;
  assign po16  = 1'b0;
  assign po17  = 1'b0;
  assign po18  = 1'b0;
  assign po19  = 1'b0;
  assign po20  = 1'b0;
  assign po21  = 1'b0;
  assign po22  = 1'b0;
  assign po23  = 1'b0;
  assign po24  = 1'b0;
  assign po25  = 1'b0;
  assign po26  = 1'b0;
  assign po27  = 1'b0;
  assign po28  = 1'b0;
  assign po29  = 1'b0;
endmodule
