module alu4_cl ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13,
    po0, po1, po2, po3, po4, po5, po6, po7  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13;
  output po0, po1, po2, po3, po4, po5, po6, po7;
  wire n23, n24, n25, n26, n27, n28, n29,
    n30, n31, n32, n33, n34, n35, n36, n37,
    n38, n39, n40, n41, n42, n43, n44, n45,
    n46, n47, n48, n49, n50, n51, n52, n53,
    n54, n55, n56, n57, n58, n59, n60, n61,
    n62, n63, n64, n65, n66, n67, n68, n69,
    n70, n71, n72, n73, n74, n75, n76, n77,
    n78, n79, n80, n81, n82, n83, n84, n85,
    n86, n87, n88, n89, n90, n91, n92, n93,
    n94, n95, n96, n97, n98, n99, n100,
    n101, n102, n103, n104, n105, n106, n107,
    n108, n109, n110, n111, n112, n113, n114,
    n115, n116, n117, n118, n119, n120, n121,
    n122, n123, n124, n125, n126, n127, n128,
    n129, n130, n131, n132, n133, n134, n135,
    n136, n137, n138, n139, n140, n141, n142,
    n143, n144, n145, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156,
    n157, n158, n159, n160, n161, n162, n163,
    n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177,
    n178, n179, n180, n181, n182, n183, n184,
    n185, n186, n187, n188, n189, n190, n191,
    n192, n193, n194, n195, n196, n197, n198,
    n199, n200, n201, n202, n203, n204, n205,
    n206, n207, n208, n209, n210, n211, n212,
    n213, n214, n215, n216, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226,
    n227, n228, n229, n230, n231, n232, n233,
    n234, n235, n236, n237, n238, n239, n240,
    n241, n242, n243, n244, n245, n246, n247,
    n248, n249, n250, n251, n252, n253, n254,
    n255, n256, n257, n258, n259, n260, n261,
    n262, n263, n264, n265, n266, n267, n268,
    n269, n270, n271, n272, n273, n274, n275,
    n276, n277, n278, n279, n280, n281, n282,
    n283, n284, n285, n286, n287, n288, n289,
    n290, n291, n292, n293, n294, n295, n296,
    n297, n298, n299, n300, n301, n302, n303,
    n304, n305, n306, n307, n308, n309, n310,
    n311, n312, n313, n314, n315, n316, n317,
    n318, n319, n320, n321, n322, n323, n324,
    n325, n326, n327, n328, n329, n330, n331,
    n332, n333, n334, n335, n336, n337, n338,
    n339, n340, n341, n342, n343, n344, n345,
    n346, n347, n348, n349, n350, n351, n352,
    n353, n354, n355, n356, n357, n358, n359,
    n360, n361, n362, n363, n364, n365, n366,
    n367, n368, n369, n370, n371, n372, n373,
    n374, n375, n376, n377, n378, n379, n380,
    n381, n382, n383, n384, n385, n386, n387,
    n388, n389, n390, n391, n392, n393, n394,
    n395, n396, n397, n398, n399, n400, n401,
    n402, n403, n404, n405, n406, n407, n408,
    n409, n410, n411, n412, n413, n414, n415,
    n416, n417, n418, n419, n420, n421, n422,
    n423, n424, n425, n426, n427, n428, n429,
    n430, n431, n432, n433, n434, n435, n436,
    n437, n438, n439, n440, n441, n442, n443,
    n444, n445, n446, n447, n448, n449, n450,
    n451, n452, n453, n454, n455, n456, n457,
    n458, n459, n460, n461, n462, n463, n464,
    n465, n466, n467, n468, n469, n470, n471,
    n472, n473, n474, n475, n476, n477, n478,
    n479, n480, n481, n482, n483, n484, n485,
    n486, n487, n488, n489, n490, n491, n492,
    n493, n494, n495, n496, n497, n498, n499,
    n500, n501, n502, n503, n504, n505, n506,
    n507, n508, n509, n510, n511, n512, n513,
    n514, n515, n516, n517, n518, n519, n520,
    n521, n522, n523, n524, n525, n526, n527,
    n528, n529, n530, n531, n532, n533, n534,
    n535, n536, n537, n538, n539, n540, n541,
    n542, n543, n544, n545, n546, n547, n548,
    n549, n550, n551, n552, n553, n554, n555,
    n556, n557, n558, n559, n560, n561, n562,
    n563, n564, n565, n566, n567, n568, n569,
    n570, n571, n572, n573, n574, n575, n576,
    n577, n578, n579, n580, n581, n582, n583,
    n584, n585, n586, n587, n588, n589, n590,
    n591, n592, n593, n594, n595, n596, n597,
    n598, n599, n600, n601, n602, n603, n604,
    n605, n606, n607, n608, n609, n610, n611,
    n612, n613, n614, n615, n616, n617, n618,
    n619, n620, n621, n622, n623, n624, n625,
    n626, n627, n628, n629, n630, n631, n632,
    n633, n634, n635, n636, n637, n638, n639,
    n640, n641, n642, n643, n644, n645, n646,
    n647, n648, n649, n650, n651, n652, n653,
    n654, n655, n656, n657, n658, n659, n660,
    n661, n662, n663, n664, n665, n666, n667,
    n668, n669, n670, n671, n672, n673, n674,
    n675, n676, n677, n678, n680, n681, n682,
    n683, n684, n685, n686, n687, n688, n689,
    n690, n691, n692, n693, n694, n695, n696,
    n697, n698, n699, n700, n701, n702, n703,
    n704, n705, n706, n707, n708, n709, n710,
    n711, n712, n713, n714, n715, n716, n717,
    n718, n719, n720, n721, n722, n723, n724,
    n725, n726, n727, n728, n729, n730, n731,
    n732, n733, n734, n735, n736, n737, n738,
    n739, n740, n741, n742, n743, n744, n745,
    n746, n747, n748, n749, n750, n751, n752,
    n753, n754, n755, n756, n757, n758, n759,
    n760, n761, n762, n763, n764, n765, n766,
    n767, n768, n769, n770, n771, n772, n773,
    n774, n775, n776, n777, n778, n779, n780,
    n781, n782, n783, n784, n785, n786, n787,
    n788, n789, n790, n791, n792, n793, n794,
    n795, n796, n797, n798, n799, n800, n801,
    n802, n803, n804, n805, n806, n807, n808,
    n809, n810, n811, n812, n813, n814, n815,
    n816, n817, n818, n819, n820, n821, n822,
    n823, n824, n825, n826, n827, n828, n829,
    n830, n831, n832, n833, n834, n835, n836,
    n837, n838, n839, n840, n841, n842, n843,
    n844, n845, n846, n847, n848, n849, n850,
    n851, n852, n853, n854, n855, n856, n857,
    n858, n859, n860, n861, n862, n863, n864,
    n865, n866, n867, n868, n869, n870, n871,
    n872, n873, n874, n875, n876, n877, n878,
    n879, n880, n881, n882, n883, n884, n885,
    n886, n887, n888, n889, n890, n891, n892,
    n893, n894, n895, n896, n897, n898, n899,
    n900, n901, n902, n903, n904, n905, n906,
    n907, n908, n909, n910, n911, n912, n913,
    n914, n915, n916, n917, n918, n919, n920,
    n921, n922, n923, n924, n925, n926, n927,
    n928, n929, n930, n931, n932, n933, n934,
    n935, n936, n937, n938, n939, n940, n941,
    n942, n943, n944, n945, n946, n947, n948,
    n949, n950, n951, n952, n953, n954, n955,
    n956, n957, n958, n959, n960, n961, n962,
    n963, n964, n965, n966, n967, n968, n969,
    n970, n971, n972, n973, n974, n975, n976,
    n977, n978, n979, n980, n981, n982, n983,
    n984, n985, n986, n987, n988, n989, n990,
    n991, n992, n993, n994, n995, n996, n997,
    n998, n999, n1000, n1001, n1002, n1003,
    n1004, n1005, n1006, n1007, n1008, n1009,
    n1010, n1011, n1012, n1013, n1014, n1015,
    n1016, n1017, n1018, n1019, n1020, n1021,
    n1022, n1023, n1024, n1025, n1026, n1027,
    n1028, n1029, n1030, n1031, n1032, n1033,
    n1034, n1035, n1036, n1037, n1038, n1039,
    n1040, n1041, n1042, n1043, n1044, n1045,
    n1046, n1047, n1048, n1049, n1050, n1052,
    n1053, n1054, n1055, n1056, n1057, n1058,
    n1059, n1060, n1061, n1062, n1063, n1064,
    n1065, n1066, n1067, n1068, n1069, n1070,
    n1071, n1072, n1073, n1074, n1075, n1076,
    n1077, n1078, n1079, n1080, n1081, n1082,
    n1083, n1084, n1085, n1086, n1087, n1088,
    n1089, n1090, n1091, n1092, n1093, n1094,
    n1095, n1096, n1097, n1098, n1099, n1100,
    n1101, n1102, n1103, n1104, n1105, n1106,
    n1107, n1108, n1109, n1110, n1111, n1112,
    n1113, n1114, n1115, n1116, n1117, n1118,
    n1119, n1120, n1121, n1122, n1123, n1124,
    n1125, n1126, n1127, n1128, n1129, n1130,
    n1131, n1132, n1133, n1134, n1135, n1136,
    n1137, n1138, n1139, n1140, n1141, n1142,
    n1143, n1144, n1145, n1146, n1147, n1148,
    n1149, n1150, n1151, n1152, n1153, n1154,
    n1155, n1156, n1157, n1158, n1159, n1160,
    n1161, n1162, n1163, n1164, n1165, n1166,
    n1167, n1168, n1169, n1170, n1171, n1172,
    n1173, n1174, n1175, n1176, n1177, n1178,
    n1179, n1180, n1181, n1182, n1183, n1184,
    n1185, n1186, n1187, n1188, n1189, n1190,
    n1191, n1192, n1193, n1194, n1195, n1196,
    n1197, n1198, n1199, n1200, n1201, n1202,
    n1203, n1204, n1205, n1206, n1207, n1208,
    n1209, n1210, n1211, n1212, n1213, n1214,
    n1215, n1216, n1217, n1218, n1219, n1220,
    n1221, n1222, n1223, n1224, n1225, n1226,
    n1227, n1228, n1229, n1230, n1231, n1232,
    n1233, n1234, n1235, n1236, n1237, n1238,
    n1239, n1240, n1241, n1242, n1243, n1244,
    n1245, n1246, n1247, n1248, n1249, n1250,
    n1251, n1252, n1253, n1254, n1255, n1256,
    n1257, n1258, n1259, n1260, n1261, n1262,
    n1263, n1264, n1265, n1266, n1267, n1268,
    n1269, n1270, n1271, n1272, n1273, n1274,
    n1275, n1276, n1277, n1278, n1279, n1280,
    n1281, n1282, n1283, n1284, n1285, n1286,
    n1287, n1288, n1289, n1290, n1291, n1292,
    n1293, n1294, n1295, n1296, n1297, n1298,
    n1299, n1300, n1301, n1302, n1303, n1304,
    n1305, n1306, n1307, n1308, n1309, n1310,
    n1311, n1312, n1313, n1314, n1315, n1316,
    n1317, n1318, n1319, n1320, n1321, n1322,
    n1323, n1324, n1325, n1326, n1327, n1328,
    n1329, n1330, n1331, n1332, n1333, n1334,
    n1335, n1336, n1337, n1338, n1339, n1340,
    n1341, n1342, n1343, n1344, n1345, n1346,
    n1347, n1348, n1349, n1350, n1351, n1352,
    n1353, n1354, n1355, n1356, n1357, n1358,
    n1359, n1360, n1361, n1362, n1363, n1364,
    n1365, n1366, n1367, n1368, n1369, n1370,
    n1371, n1372, n1373, n1374, n1375, n1376,
    n1377, n1378, n1379, n1380, n1381, n1382,
    n1383, n1384, n1385, n1386, n1387, n1388,
    n1389, n1390, n1391, n1392, n1393, n1394,
    n1395, n1396, n1397, n1398, n1399, n1400,
    n1401, n1402, n1403, n1404, n1405, n1406,
    n1407, n1408, n1409, n1410, n1411;
  assign n23 = pi00 & pi04;
  assign n24 = ~pi10 & pi13;
  assign n25 = ~pi08 & pi11;
  assign n26 = pi09 & n25;
  assign n27 = pi09 & pi11;
  assign n28 = ~pi08 & pi13;
  assign n29 = pi09 & pi13;
  assign n30 = n25 & n29;
  assign n31 = n27 & n28;
  assign n32 = ~pi10 & n1239;
  assign n33 = n24 & n26;
  assign n34 = n23 & n1240;
  assign n35 = pi10 & ~pi11;
  assign n36 = ~pi08 & pi09;
  assign n37 = pi13 & n36;
  assign n38 = ~n35 & n36;
  assign n39 = pi13 & n38;
  assign n40 = ~n35 & n37;
  assign n41 = pi08 & pi10;
  assign n42 = ~pi09 & pi11;
  assign n43 = ~pi13 & n42;
  assign n44 = ~pi13 & n41;
  assign n45 = n42 & n44;
  assign n46 = n41 & n43;
  assign n47 = pi08 & pi09;
  assign n48 = n35 & n47;
  assign n49 = ~n1242 & ~n48;
  assign n50 = ~n1241 & ~n1242;
  assign n51 = ~n48 & n50;
  assign n52 = ~n1241 & ~n48;
  assign n53 = ~n1242 & n52;
  assign n54 = ~n1241 & n49;
  assign n55 = ~pi04 & ~n1243;
  assign n56 = ~pi08 & ~pi09;
  assign n57 = ~n47 & ~n56;
  assign n58 = ~pi10 & pi11;
  assign n59 = pi11 & ~n57;
  assign n60 = ~pi10 & n59;
  assign n61 = ~n57 & n58;
  assign n62 = pi13 & n1244;
  assign n63 = ~pi09 & ~pi11;
  assign n64 = ~pi08 & pi10;
  assign n65 = ~pi08 & n35;
  assign n66 = ~pi09 & n65;
  assign n67 = n63 & n64;
  assign n68 = ~n62 & ~n1245;
  assign n69 = n23 & ~n68;
  assign n70 = ~pi00 & ~pi04;
  assign n71 = ~pi10 & ~pi11;
  assign n72 = ~pi13 & ~n71;
  assign n73 = pi08 & ~pi09;
  assign n74 = ~n24 & n73;
  assign n75 = pi10 & pi13;
  assign n76 = ~pi13 & n71;
  assign n77 = ~n75 & ~n76;
  assign n78 = n73 & ~n77;
  assign n79 = ~n72 & n74;
  assign n80 = ~n70 & n1246;
  assign n81 = ~pi10 & ~pi13;
  assign n82 = ~pi10 & ~n27;
  assign n83 = ~pi13 & n82;
  assign n84 = ~n27 & n81;
  assign n85 = ~pi08 & ~pi10;
  assign n86 = ~pi13 & ~n27;
  assign n87 = n85 & n86;
  assign n88 = ~pi13 & n85;
  assign n89 = ~n27 & n88;
  assign n90 = ~pi08 & n1247;
  assign n91 = ~pi00 & n1248;
  assign n92 = ~pi00 & ~n35;
  assign n93 = ~pi00 & pi04;
  assign n94 = pi00 & ~pi04;
  assign n95 = ~n93 & ~n94;
  assign n96 = ~n23 & ~n70;
  assign n97 = n37 & ~n1249;
  assign n98 = n35 & n93;
  assign n99 = ~n94 & ~n98;
  assign n100 = pi13 & ~n99;
  assign n101 = n36 & n100;
  assign n102 = n37 & ~n99;
  assign n103 = ~n92 & n97;
  assign n104 = ~n91 & ~n1250;
  assign n105 = ~n80 & n104;
  assign n106 = ~n69 & n105;
  assign n107 = ~n80 & ~n1250;
  assign n108 = ~n69 & n107;
  assign n109 = ~n55 & n108;
  assign n110 = ~n91 & n109;
  assign n111 = ~n69 & ~n80;
  assign n112 = ~n55 & ~n91;
  assign n113 = n111 & n112;
  assign n114 = ~n1250 & n113;
  assign n115 = ~n55 & n106;
  assign n116 = ~pi00 & n1251;
  assign n117 = n1239 & ~n116;
  assign n118 = pi13 & n35;
  assign n119 = pi00 & ~n1251;
  assign n120 = pi00 & ~n109;
  assign n121 = n47 & n1252;
  assign n122 = n56 & n1251;
  assign n123 = n23 & n73;
  assign n124 = ~n122 & ~n123;
  assign n125 = ~n121 & ~n123;
  assign n126 = ~n122 & n125;
  assign n127 = ~n121 & n124;
  assign n128 = n118 & ~n1253;
  assign n129 = ~n117 & ~n128;
  assign n130 = pi08 & n35;
  assign n131 = ~pi09 & pi13;
  assign n132 = n130 & n131;
  assign n133 = n73 & n118;
  assign n134 = n129 & n1254;
  assign n135 = ~n34 & ~n134;
  assign n136 = pi10 & n63;
  assign n137 = ~pi09 & n35;
  assign n138 = pi08 & n1255;
  assign n139 = n35 & n73;
  assign n140 = pi08 & n135;
  assign n141 = n1255 & n140;
  assign n142 = n135 & n1256;
  assign n143 = ~pi10 & ~n56;
  assign n144 = ~pi00 & pi11;
  assign n145 = pi11 & ~n143;
  assign n146 = ~pi00 & n145;
  assign n147 = ~pi00 & ~n143;
  assign n148 = pi11 & n147;
  assign n149 = ~n143 & n144;
  assign n150 = ~n1251 & ~n1258;
  assign n151 = ~n1257 & n150;
  assign n152 = pi00 & pi11;
  assign n153 = ~n47 & n152;
  assign n154 = ~n134 & ~n153;
  assign n155 = pi10 & ~n154;
  assign n156 = ~pi10 & n47;
  assign n157 = pi11 & n156;
  assign n158 = n47 & n58;
  assign n159 = pi10 & n36;
  assign n160 = ~pi11 & n159;
  assign n161 = pi09 & n65;
  assign n162 = n35 & n36;
  assign n163 = ~n1259 & ~n1260;
  assign n164 = n1251 & n163;
  assign n165 = ~n155 & n164;
  assign n166 = ~n151 & ~n165;
  assign n167 = pi09 & ~pi10;
  assign n168 = n25 & n167;
  assign n169 = pi09 & n85;
  assign n170 = pi11 & n169;
  assign n171 = n36 & n58;
  assign n172 = n135 & n169;
  assign n173 = pi11 & n172;
  assign n174 = n135 & n1261;
  assign n175 = ~pi00 & ~pi08;
  assign n176 = n1255 & n175;
  assign n177 = ~pi00 & n1245;
  assign n178 = ~n129 & ~n1263;
  assign n179 = ~n1262 & n178;
  assign n180 = ~n48 & n129;
  assign n181 = ~n179 & ~n180;
  assign n182 = pi08 & ~pi10;
  assign n183 = pi04 & n182;
  assign n184 = pi00 & ~pi08;
  assign n185 = n129 & n184;
  assign n186 = ~n183 & ~n185;
  assign n187 = n63 & ~n186;
  assign n188 = pi09 & ~n1251;
  assign n189 = ~pi00 & ~n188;
  assign n190 = ~pi09 & n1251;
  assign n191 = pi11 & ~n190;
  assign n192 = n85 & ~n191;
  assign n193 = n85 & ~n189;
  assign n194 = ~n191 & n193;
  assign n195 = ~pi11 & ~n189;
  assign n196 = pi00 & ~pi09;
  assign n197 = n1251 & n196;
  assign n198 = ~n195 & ~n197;
  assign n199 = n85 & ~n198;
  assign n200 = ~n189 & n192;
  assign n201 = pi09 & n41;
  assign n202 = pi10 & n47;
  assign n203 = ~pi00 & n1265;
  assign n204 = pi11 & n203;
  assign n205 = n144 & n1265;
  assign n206 = ~pi10 & n73;
  assign n207 = ~pi09 & n182;
  assign n208 = ~pi10 & ~n1249;
  assign n209 = n73 & n208;
  assign n210 = ~n1249 & n1267;
  assign n211 = ~n1266 & ~n1268;
  assign n212 = ~n1264 & n211;
  assign n213 = ~n187 & n212;
  assign n214 = ~n181 & n213;
  assign n215 = ~n1262 & ~n1263;
  assign n216 = ~n129 & ~n215;
  assign n217 = ~n1257 & ~n1258;
  assign n218 = ~n1251 & ~n217;
  assign n219 = ~n155 & n163;
  assign n220 = n1251 & ~n219;
  assign n221 = ~n34 & ~n48;
  assign n222 = n129 & ~n221;
  assign n223 = ~n1266 & ~n222;
  assign n224 = ~n187 & n223;
  assign n225 = ~n220 & n224;
  assign n226 = ~n218 & n225;
  assign n227 = ~n1264 & n226;
  assign n228 = ~n216 & n227;
  assign n229 = ~n1268 & n228;
  assign n230 = n213 & ~n216;
  assign n231 = ~n218 & ~n222;
  assign n232 = n213 & ~n222;
  assign n233 = ~n216 & ~n218;
  assign n234 = n232 & n233;
  assign n235 = n230 & n231;
  assign n236 = ~n220 & n1270;
  assign n237 = ~n166 & n214;
  assign n238 = ~pi12 & pi13;
  assign n239 = pi13 & ~n1269;
  assign n240 = ~pi12 & n239;
  assign n241 = ~n1269 & n238;
  assign n242 = pi01 & pi05;
  assign n243 = pi13 & n1255;
  assign n244 = n68 & ~n243;
  assign n245 = ~pi08 & n93;
  assign n246 = n28 & n98;
  assign n247 = n118 & n245;
  assign n248 = n244 & ~n1272;
  assign n249 = n242 & ~n248;
  assign n250 = ~pi05 & ~n1243;
  assign n251 = ~pi09 & pi10;
  assign n252 = n152 & n251;
  assign n253 = ~pi01 & pi05;
  assign n254 = n35 & n253;
  assign n255 = pi01 & ~pi05;
  assign n256 = ~n93 & ~n255;
  assign n257 = ~n254 & n256;
  assign n258 = ~pi01 & ~pi05;
  assign n259 = n93 & ~n258;
  assign n260 = pi09 & ~n259;
  assign n261 = ~n254 & ~n255;
  assign n262 = ~n93 & ~n261;
  assign n263 = n93 & n258;
  assign n264 = ~n262 & ~n263;
  assign n265 = pi09 & ~n264;
  assign n266 = ~n257 & n260;
  assign n267 = ~n252 & ~n1273;
  assign n268 = ~pi08 & ~n267;
  assign n269 = pi13 & n268;
  assign n270 = n28 & ~n267;
  assign n271 = ~pi01 & n1248;
  assign n272 = n1246 & ~n258;
  assign n273 = ~n271 & ~n272;
  assign n274 = ~n1274 & n273;
  assign n275 = ~n250 & ~n271;
  assign n276 = ~n272 & n275;
  assign n277 = ~n250 & n273;
  assign n278 = ~n1274 & n1275;
  assign n279 = ~n250 & n274;
  assign n280 = ~n249 & n1275;
  assign n281 = ~n1274 & n280;
  assign n282 = ~n249 & n1276;
  assign n283 = n1240 & n242;
  assign n284 = ~pi01 & n1277;
  assign n285 = ~pi01 & n1276;
  assign n286 = n1239 & ~n1278;
  assign n287 = ~pi05 & ~pi09;
  assign n288 = pi01 & pi08;
  assign n289 = ~n287 & n288;
  assign n290 = ~pi08 & n1277;
  assign n291 = ~n289 & ~n290;
  assign n292 = pi09 & n1277;
  assign n293 = n118 & ~n292;
  assign n294 = n56 & n1277;
  assign n295 = pi09 & ~n1277;
  assign n296 = pi05 & ~pi09;
  assign n297 = ~n295 & ~n296;
  assign n298 = pi08 & ~n297;
  assign n299 = pi01 & n298;
  assign n300 = n288 & ~n297;
  assign n301 = ~n294 & ~n1279;
  assign n302 = n118 & ~n301;
  assign n303 = ~n291 & n293;
  assign n304 = ~n286 & ~n1280;
  assign n305 = n1254 & n304;
  assign n306 = ~n283 & ~n305;
  assign n307 = ~n1251 & ~n135;
  assign n308 = ~n306 & n307;
  assign n309 = n306 & ~n307;
  assign n310 = ~n306 & ~n307;
  assign n311 = n306 & n307;
  assign n312 = ~n310 & ~n311;
  assign n313 = ~n308 & ~n309;
  assign n314 = ~n1277 & ~n1281;
  assign n315 = n1277 & n1281;
  assign n316 = n41 & ~n315;
  assign n317 = ~n1277 & n1281;
  assign n318 = n1277 & ~n1281;
  assign n319 = ~n317 & ~n318;
  assign n320 = n41 & ~n319;
  assign n321 = ~n314 & n316;
  assign n322 = pi05 & n182;
  assign n323 = pi00 & ~n129;
  assign n324 = n304 & ~n323;
  assign n325 = ~n129 & ~n304;
  assign n326 = pi00 & n325;
  assign n327 = n304 & n323;
  assign n328 = ~n304 & ~n323;
  assign n329 = ~n327 & ~n328;
  assign n330 = ~n324 & ~n326;
  assign n331 = pi01 & ~pi08;
  assign n332 = ~pi08 & n1283;
  assign n333 = pi01 & n332;
  assign n334 = n1283 & n331;
  assign n335 = ~n322 & ~n1284;
  assign n336 = ~n1282 & n335;
  assign n337 = n63 & ~n336;
  assign n338 = n34 & ~n306;
  assign n339 = ~n34 & n306;
  assign n340 = n34 & n306;
  assign n341 = ~n34 & ~n306;
  assign n342 = ~n340 & ~n341;
  assign n343 = ~n338 & ~n339;
  assign n344 = ~n304 & ~n1285;
  assign n345 = n304 & n1285;
  assign n346 = n1261 & ~n345;
  assign n347 = n1261 & ~n344;
  assign n348 = ~n345 & n347;
  assign n349 = ~n304 & n1285;
  assign n350 = n304 & ~n1285;
  assign n351 = ~n349 & ~n350;
  assign n352 = n1261 & ~n351;
  assign n353 = ~n344 & n346;
  assign n354 = pi10 & ~n47;
  assign n355 = ~n56 & ~n354;
  assign n356 = pi11 & ~n355;
  assign n357 = n1252 & ~n1277;
  assign n358 = ~n1252 & n1277;
  assign n359 = n1252 & n1277;
  assign n360 = ~n1252 & ~n1277;
  assign n361 = ~n359 & ~n360;
  assign n362 = ~n357 & ~n358;
  assign n363 = n356 & ~n1287;
  assign n364 = n64 & ~n1283;
  assign n365 = n63 & n364;
  assign n366 = n1245 & ~n1283;
  assign n367 = ~n363 & ~n1288;
  assign n368 = ~pi01 & ~n367;
  assign n369 = n129 & n304;
  assign n370 = ~n325 & ~n369;
  assign n371 = n1265 & ~n370;
  assign n372 = n169 & ~n1277;
  assign n373 = ~n371 & ~n372;
  assign n374 = ~pi11 & ~n373;
  assign n375 = ~pi10 & n56;
  assign n376 = ~n356 & ~n375;
  assign n377 = ~n35 & ~n355;
  assign n378 = n1287 & ~n1289;
  assign n379 = n152 & n1265;
  assign n380 = ~pi05 & ~n23;
  assign n381 = n1267 & n380;
  assign n382 = ~n47 & n71;
  assign n383 = ~n381 & ~n382;
  assign n384 = ~n379 & ~n381;
  assign n385 = ~n382 & n384;
  assign n386 = ~n379 & ~n382;
  assign n387 = ~n381 & n386;
  assign n388 = ~n379 & n383;
  assign n389 = ~n378 & n1290;
  assign n390 = pi01 & ~n389;
  assign n391 = n1251 & n1277;
  assign n392 = ~n163 & n391;
  assign n393 = ~pi11 & n36;
  assign n394 = ~n1259 & ~n393;
  assign n395 = ~n1251 & ~n394;
  assign n396 = ~n1277 & n395;
  assign n397 = ~pi00 & ~pi01;
  assign n398 = n1265 & n397;
  assign n399 = n23 & n258;
  assign n400 = n1267 & n399;
  assign n401 = ~n398 & ~n400;
  assign n402 = pi11 & ~n401;
  assign n403 = n23 & ~n242;
  assign n404 = ~n23 & ~n253;
  assign n405 = n1267 & ~n404;
  assign n406 = ~n23 & n253;
  assign n407 = n23 & n242;
  assign n408 = ~n406 & ~n407;
  assign n409 = n1267 & ~n408;
  assign n410 = ~n403 & n405;
  assign n411 = ~n402 & ~n1291;
  assign n412 = ~n396 & n411;
  assign n413 = ~n392 & n412;
  assign n414 = ~n390 & n413;
  assign n415 = ~n374 & n414;
  assign n416 = ~n368 & n414;
  assign n417 = ~n374 & n416;
  assign n418 = ~n368 & n415;
  assign n419 = ~n1286 & n1292;
  assign n420 = ~n392 & ~n396;
  assign n421 = ~n1291 & n420;
  assign n422 = ~n374 & n421;
  assign n423 = ~n390 & n422;
  assign n424 = ~n1286 & n423;
  assign n425 = ~n402 & n424;
  assign n426 = ~n337 & n425;
  assign n427 = ~n368 & n426;
  assign n428 = ~n337 & n419;
  assign n429 = pi13 & ~n1293;
  assign n430 = n1271 & n429;
  assign n431 = n1271 & ~n1293;
  assign n432 = ~n93 & ~n253;
  assign n433 = n93 & ~n255;
  assign n434 = ~n253 & ~n433;
  assign n435 = ~n255 & ~n432;
  assign n436 = ~pi06 & pi09;
  assign n437 = ~pi06 & n1295;
  assign n438 = pi09 & n437;
  assign n439 = pi09 & n1295;
  assign n440 = ~pi06 & n439;
  assign n441 = n1295 & n436;
  assign n442 = pi06 & n35;
  assign n443 = n35 & ~n1295;
  assign n444 = pi06 & n443;
  assign n445 = ~n1295 & n442;
  assign n446 = ~n1296 & ~n1297;
  assign n447 = pi02 & ~n446;
  assign n448 = pi01 & pi11;
  assign n449 = n251 & n448;
  assign n450 = n1295 & ~n442;
  assign n451 = pi06 & ~n1295;
  assign n452 = ~pi02 & pi09;
  assign n453 = ~n451 & n452;
  assign n454 = ~pi06 & ~n1295;
  assign n455 = n35 & n1295;
  assign n456 = pi06 & n455;
  assign n457 = n1295 & n442;
  assign n458 = ~n454 & ~n1298;
  assign n459 = pi09 & ~n458;
  assign n460 = ~pi02 & n459;
  assign n461 = n452 & ~n458;
  assign n462 = ~n450 & n453;
  assign n463 = ~n449 & ~n1299;
  assign n464 = ~n447 & ~n449;
  assign n465 = ~n1299 & n464;
  assign n466 = ~n447 & n463;
  assign n467 = ~pi08 & ~n1300;
  assign n468 = pi13 & n467;
  assign n469 = n28 & ~n1300;
  assign n470 = pi02 & pi06;
  assign n471 = ~n244 & n470;
  assign n472 = ~pi06 & ~n1243;
  assign n473 = ~pi02 & n1248;
  assign n474 = ~pi02 & ~pi06;
  assign n475 = n1246 & ~n474;
  assign n476 = ~n473 & ~n475;
  assign n477 = ~n472 & n476;
  assign n478 = ~n471 & ~n472;
  assign n479 = n476 & n478;
  assign n480 = ~n471 & n477;
  assign n481 = ~n1301 & n1302;
  assign n482 = n1240 & n470;
  assign n483 = ~pi02 & n481;
  assign n484 = n1239 & ~n483;
  assign n485 = ~pi06 & ~pi09;
  assign n486 = pi02 & pi08;
  assign n487 = ~n485 & n486;
  assign n488 = ~pi08 & n481;
  assign n489 = ~n487 & ~n488;
  assign n490 = pi09 & n481;
  assign n491 = n118 & ~n490;
  assign n492 = n56 & n481;
  assign n493 = pi09 & ~n481;
  assign n494 = pi06 & ~pi09;
  assign n495 = ~n493 & ~n494;
  assign n496 = pi08 & ~n495;
  assign n497 = pi02 & n496;
  assign n498 = n486 & ~n495;
  assign n499 = ~n492 & ~n1303;
  assign n500 = n118 & ~n499;
  assign n501 = ~n489 & n491;
  assign n502 = ~n484 & ~n1304;
  assign n503 = n1254 & n502;
  assign n504 = ~n482 & ~n503;
  assign n505 = n481 & n504;
  assign n506 = ~n481 & ~n504;
  assign n507 = ~n505 & ~n506;
  assign n508 = ~n1277 & ~n309;
  assign n509 = ~n308 & ~n508;
  assign n510 = ~n507 & n509;
  assign n511 = n507 & ~n509;
  assign n512 = n41 & ~n511;
  assign n513 = n41 & ~n510;
  assign n514 = ~n511 & n513;
  assign n515 = ~n507 & ~n509;
  assign n516 = n507 & n509;
  assign n517 = ~n515 & ~n516;
  assign n518 = n41 & ~n517;
  assign n519 = ~n510 & n512;
  assign n520 = pi06 & n182;
  assign n521 = pi01 & ~n324;
  assign n522 = ~pi01 & ~n323;
  assign n523 = ~n304 & ~n522;
  assign n524 = pi01 & n323;
  assign n525 = ~n523 & ~n524;
  assign n526 = ~n326 & ~n521;
  assign n527 = ~n502 & ~n1306;
  assign n528 = n502 & n1306;
  assign n529 = ~n502 & n1306;
  assign n530 = n502 & ~n1306;
  assign n531 = ~n529 & ~n530;
  assign n532 = ~n527 & ~n528;
  assign n533 = pi02 & ~pi08;
  assign n534 = ~pi08 & n1307;
  assign n535 = pi02 & n534;
  assign n536 = n1307 & n533;
  assign n537 = ~n520 & ~n1308;
  assign n538 = ~n1305 & n537;
  assign n539 = n63 & ~n538;
  assign n540 = ~n304 & ~n339;
  assign n541 = n504 & ~n540;
  assign n542 = ~n504 & n540;
  assign n543 = ~n541 & ~n542;
  assign n544 = n502 & ~n543;
  assign n545 = ~n502 & n543;
  assign n546 = n1261 & ~n545;
  assign n547 = n1261 & ~n544;
  assign n548 = ~n545 & n547;
  assign n549 = ~n502 & n540;
  assign n550 = n502 & ~n540;
  assign n551 = ~n502 & ~n540;
  assign n552 = n502 & n540;
  assign n553 = ~n551 & ~n552;
  assign n554 = ~n549 & ~n550;
  assign n555 = ~n504 & n1310;
  assign n556 = n504 & ~n1310;
  assign n557 = ~n555 & ~n556;
  assign n558 = n1261 & ~n557;
  assign n559 = ~n544 & n546;
  assign n560 = n64 & ~n1307;
  assign n561 = n63 & n560;
  assign n562 = n1245 & ~n1307;
  assign n563 = pi01 & ~n358;
  assign n564 = ~pi01 & ~n357;
  assign n565 = ~n358 & ~n564;
  assign n566 = ~pi01 & ~n1252;
  assign n567 = ~n1277 & ~n566;
  assign n568 = pi01 & n1252;
  assign n569 = ~n567 & ~n568;
  assign n570 = ~n357 & ~n563;
  assign n571 = n356 & ~n481;
  assign n572 = n356 & ~n1312;
  assign n573 = ~n481 & n572;
  assign n574 = ~n1312 & n571;
  assign n575 = ~n1311 & ~n1313;
  assign n576 = ~pi02 & ~n575;
  assign n577 = n369 & n502;
  assign n578 = ~n369 & ~n502;
  assign n579 = ~pi11 & ~n578;
  assign n580 = ~pi11 & ~n577;
  assign n581 = ~n578 & n580;
  assign n582 = ~n577 & n579;
  assign n583 = pi02 & ~n397;
  assign n584 = ~pi02 & n397;
  assign n585 = pi11 & ~n584;
  assign n586 = pi11 & ~n583;
  assign n587 = ~n584 & n586;
  assign n588 = ~n583 & n585;
  assign n589 = n1265 & ~n1315;
  assign n590 = ~n577 & ~n578;
  assign n591 = ~pi11 & ~n590;
  assign n592 = pi11 & n584;
  assign n593 = pi02 & pi11;
  assign n594 = ~n397 & n593;
  assign n595 = ~n592 & ~n594;
  assign n596 = ~n591 & n595;
  assign n597 = n1265 & ~n596;
  assign n598 = ~n1314 & n589;
  assign n599 = ~n1289 & ~n481;
  assign n600 = ~n1289 & n1312;
  assign n601 = n356 & n1312;
  assign n602 = ~n481 & n1317;
  assign n603 = ~n481 & n1312;
  assign n604 = ~n1289 & n603;
  assign n605 = n1312 & n599;
  assign n606 = ~n382 & ~n1318;
  assign n607 = pi02 & ~n606;
  assign n608 = ~pi02 & n356;
  assign n609 = ~pi02 & n1317;
  assign n610 = n1312 & n608;
  assign n611 = pi02 & ~n1289;
  assign n612 = ~n1289 & ~n1312;
  assign n613 = pi02 & n612;
  assign n614 = ~n1312 & n611;
  assign n615 = ~n1319 & ~n1320;
  assign n616 = ~n608 & ~n612;
  assign n617 = ~pi02 & ~n1312;
  assign n618 = n481 & ~n617;
  assign n619 = ~n616 & n618;
  assign n620 = n481 & ~n615;
  assign n621 = ~pi11 & n169;
  assign n622 = ~pi10 & n393;
  assign n623 = n391 & ~n1322;
  assign n624 = ~n394 & ~n481;
  assign n625 = ~n391 & ~n394;
  assign n626 = ~n1322 & ~n625;
  assign n627 = ~n481 & ~n626;
  assign n628 = ~n623 & n624;
  assign n629 = ~n23 & ~n242;
  assign n630 = n23 & ~n258;
  assign n631 = ~n242 & ~n630;
  assign n632 = ~n258 & ~n629;
  assign n633 = pi11 & n474;
  assign n634 = ~n470 & ~n633;
  assign n635 = ~n1324 & n634;
  assign n636 = ~pi02 & pi06;
  assign n637 = pi02 & ~pi06;
  assign n638 = ~n636 & ~n637;
  assign n639 = ~n470 & ~n474;
  assign n640 = n1324 & n1325;
  assign n641 = n1267 & ~n640;
  assign n642 = ~n1324 & ~n634;
  assign n643 = n1324 & ~n1325;
  assign n644 = ~n642 & ~n643;
  assign n645 = n1267 & ~n644;
  assign n646 = ~n635 & n641;
  assign n647 = n391 & n481;
  assign n648 = ~n163 & n647;
  assign n649 = n392 & n481;
  assign n650 = ~n1326 & ~n1327;
  assign n651 = ~n1323 & n650;
  assign n652 = ~n1321 & n651;
  assign n653 = n481 & ~n1312;
  assign n654 = ~n603 & ~n653;
  assign n655 = ~n1289 & ~n654;
  assign n656 = ~n382 & ~n655;
  assign n657 = pi02 & ~n656;
  assign n658 = ~n392 & ~n1319;
  assign n659 = n481 & ~n658;
  assign n660 = ~n1323 & ~n1326;
  assign n661 = ~n659 & n660;
  assign n662 = ~n657 & n661;
  assign n663 = ~n607 & n652;
  assign n664 = ~n1316 & n1328;
  assign n665 = ~n576 & n664;
  assign n666 = ~n1309 & n665;
  assign n667 = ~n1316 & ~n1327;
  assign n668 = ~n1323 & n667;
  assign n669 = ~n607 & n668;
  assign n670 = ~n539 & n669;
  assign n671 = ~n1309 & n670;
  assign n672 = ~n576 & n671;
  assign n673 = ~n1326 & n672;
  assign n674 = ~n1321 & n673;
  assign n675 = ~n539 & n666;
  assign n676 = pi13 & ~n1329;
  assign n677 = n1294 & n676;
  assign n678 = n1294 & ~n1329;
  assign po5 = pi03 & pi07;
  assign n680 = n1295 & ~n636;
  assign n681 = pi02 & ~n451;
  assign n682 = ~n437 & ~n681;
  assign n683 = ~n637 & ~n680;
  assign n684 = n35 & n1331;
  assign n685 = pi13 & n684;
  assign n686 = n118 & n1331;
  assign n687 = ~n1255 & ~n1332;
  assign n688 = po5 & ~n687;
  assign n689 = pi07 & n35;
  assign n690 = pi07 & pi09;
  assign n691 = n118 & n690;
  assign n692 = n29 & n689;
  assign n693 = pi07 & pi13;
  assign n694 = pi09 & n35;
  assign n695 = ~n1331 & n694;
  assign n696 = n693 & n695;
  assign n697 = ~n1331 & n1333;
  assign n698 = ~n1247 & ~n1334;
  assign n699 = ~pi03 & ~n698;
  assign n700 = n251 & n593;
  assign n701 = ~pi03 & ~pi07;
  assign n702 = pi09 & n701;
  assign n703 = pi09 & n1331;
  assign n704 = n701 & n703;
  assign n705 = n1331 & n702;
  assign n706 = ~n700 & ~n1335;
  assign n707 = pi13 & ~n706;
  assign n708 = ~n699 & ~n707;
  assign n709 = ~n688 & ~n707;
  assign n710 = ~n699 & n709;
  assign n711 = ~n688 & ~n699;
  assign n712 = ~n707 & n711;
  assign n713 = ~n688 & n708;
  assign n714 = ~pi08 & ~n1336;
  assign n715 = pi03 & pi09;
  assign n716 = pi03 & n37;
  assign n717 = n28 & n715;
  assign n718 = pi09 & ~n1331;
  assign n719 = pi03 & n718;
  assign n720 = n28 & n719;
  assign n721 = ~n1331 & n1337;
  assign n722 = n1243 & ~n1338;
  assign n723 = ~pi07 & ~n722;
  assign n724 = n1246 & ~n701;
  assign n725 = ~n1244 & ~n1255;
  assign n726 = pi13 & po5;
  assign n727 = pi13 & ~n725;
  assign n728 = po5 & n727;
  assign n729 = ~n725 & n726;
  assign n730 = ~n724 & ~n1339;
  assign n731 = ~n723 & n730;
  assign n732 = ~n714 & n730;
  assign n733 = ~n723 & n732;
  assign n734 = ~n714 & n731;
  assign n735 = ~pi03 & n1340;
  assign n736 = n1239 & ~n735;
  assign n737 = pi03 & ~n1340;
  assign n738 = n47 & n737;
  assign n739 = n73 & po5;
  assign n740 = n56 & n1340;
  assign n741 = ~n739 & ~n740;
  assign n742 = ~n738 & ~n739;
  assign n743 = ~n740 & n742;
  assign n744 = ~n738 & n741;
  assign n745 = n118 & ~n1341;
  assign n746 = ~n736 & ~n745;
  assign n747 = n1240 & po5;
  assign n748 = n1254 & n746;
  assign n749 = ~n747 & ~n748;
  assign n750 = ~n502 & ~n541;
  assign n751 = n749 & ~n750;
  assign n752 = ~n749 & n750;
  assign n753 = ~n751 & ~n752;
  assign n754 = ~n746 & n753;
  assign n755 = n746 & ~n753;
  assign n756 = n169 & ~n755;
  assign n757 = ~n746 & n750;
  assign n758 = n746 & ~n750;
  assign n759 = ~n746 & ~n750;
  assign n760 = n746 & n750;
  assign n761 = ~n759 & ~n760;
  assign n762 = ~n757 & ~n758;
  assign n763 = ~n749 & n1342;
  assign n764 = n749 & ~n1342;
  assign n765 = ~n763 & ~n764;
  assign n766 = n169 & ~n765;
  assign n767 = ~n754 & n756;
  assign n768 = ~pi03 & n1265;
  assign n769 = ~pi03 & n584;
  assign n770 = n1265 & n769;
  assign n771 = n584 & n768;
  assign n772 = ~n470 & n1324;
  assign n773 = ~n474 & ~n1324;
  assign n774 = ~n470 & ~n773;
  assign n775 = ~n474 & ~n772;
  assign n776 = ~pi03 & n1267;
  assign n777 = ~pi07 & n776;
  assign n778 = n1267 & n701;
  assign n779 = n701 & ~n1345;
  assign n780 = n1267 & n779;
  assign n781 = ~pi07 & ~n1345;
  assign n782 = n776 & n781;
  assign n783 = ~n1345 & n1346;
  assign n784 = ~n1344 & ~n1347;
  assign n785 = ~n1343 & n784;
  assign n786 = pi11 & ~n785;
  assign n787 = ~pi02 & n502;
  assign n788 = ~n1306 & ~n787;
  assign n789 = pi02 & ~n502;
  assign n790 = pi02 & ~n528;
  assign n791 = ~n527 & ~n790;
  assign n792 = ~pi02 & n1306;
  assign n793 = ~n502 & ~n792;
  assign n794 = pi02 & ~n1306;
  assign n795 = ~n793 & ~n794;
  assign n796 = ~n788 & ~n789;
  assign n797 = ~n746 & ~n1348;
  assign n798 = ~pi03 & ~n797;
  assign n799 = n746 & n1348;
  assign n800 = ~pi08 & ~n799;
  assign n801 = n746 & ~n1348;
  assign n802 = ~n746 & n1348;
  assign n803 = ~n801 & ~n802;
  assign n804 = ~n797 & ~n799;
  assign n805 = ~pi08 & ~n1349;
  assign n806 = ~pi03 & n805;
  assign n807 = ~pi03 & ~pi08;
  assign n808 = ~n1349 & n807;
  assign n809 = n798 & n800;
  assign n810 = ~n1340 & ~n749;
  assign n811 = n1340 & n749;
  assign n812 = ~n1340 & n749;
  assign n813 = n1340 & ~n749;
  assign n814 = ~n812 & ~n813;
  assign n815 = ~n810 & ~n811;
  assign n816 = n504 & n509;
  assign n817 = ~n481 & ~n816;
  assign n818 = ~n504 & ~n509;
  assign n819 = ~n817 & ~n818;
  assign n820 = ~n506 & n509;
  assign n821 = ~n1351 & ~n1352;
  assign n822 = n1351 & n1352;
  assign n823 = pi08 & ~n822;
  assign n824 = n1351 & ~n1352;
  assign n825 = ~n1351 & n1352;
  assign n826 = ~n824 & ~n825;
  assign n827 = pi08 & ~n826;
  assign n828 = ~n821 & n823;
  assign n829 = ~n1350 & ~n1353;
  assign n830 = n1255 & ~n829;
  assign n831 = pi03 & n56;
  assign n832 = n56 & n1349;
  assign n833 = pi03 & n832;
  assign n834 = n1349 & n831;
  assign n835 = pi07 & n1267;
  assign n836 = n577 & n746;
  assign n837 = ~n577 & ~n746;
  assign n838 = ~n836 & ~n837;
  assign n839 = n1265 & ~n838;
  assign n840 = ~n835 & ~n839;
  assign n841 = ~n1354 & ~n835;
  assign n842 = ~n839 & n841;
  assign n843 = ~n1354 & n840;
  assign n844 = ~pi11 & ~n1355;
  assign n845 = pi02 & ~n653;
  assign n846 = ~pi02 & ~n603;
  assign n847 = ~n653 & ~n846;
  assign n848 = ~n481 & ~n617;
  assign n849 = pi02 & n1312;
  assign n850 = ~n848 & ~n849;
  assign n851 = ~n603 & ~n845;
  assign n852 = ~n1340 & ~n1356;
  assign n853 = n1340 & n1356;
  assign n854 = ~n1340 & n1356;
  assign n855 = n1340 & ~n1356;
  assign n856 = ~n854 & ~n855;
  assign n857 = ~n852 & ~n853;
  assign n858 = ~n1289 & ~n1357;
  assign n859 = ~n382 & ~n858;
  assign n860 = pi03 & ~n859;
  assign n861 = n356 & n1357;
  assign n862 = pi07 & n1345;
  assign n863 = n1267 & n862;
  assign n864 = n1345 & n835;
  assign n865 = ~n861 & ~n1358;
  assign n866 = ~pi03 & ~n865;
  assign n867 = ~n1322 & n647;
  assign n868 = ~n394 & ~n647;
  assign n869 = ~n1322 & ~n868;
  assign n870 = ~n394 & ~n867;
  assign n871 = ~n1340 & ~n1359;
  assign n872 = pi03 & ~pi07;
  assign n873 = ~pi07 & n1345;
  assign n874 = pi03 & n873;
  assign n875 = n1345 & n872;
  assign n876 = po5 & ~n1345;
  assign n877 = ~n1360 & ~n876;
  assign n878 = pi03 & n1267;
  assign n879 = ~n781 & n878;
  assign n880 = ~n862 & n879;
  assign n881 = n1267 & ~n877;
  assign n882 = pi03 & pi11;
  assign n883 = n1265 & n882;
  assign n884 = ~n584 & n882;
  assign n885 = n1265 & n884;
  assign n886 = ~n584 & n883;
  assign n887 = pi07 & ~n1345;
  assign n888 = ~n873 & ~n887;
  assign n889 = n1267 & ~n888;
  assign n890 = n1265 & n585;
  assign n891 = ~n889 & ~n890;
  assign n892 = pi03 & ~n891;
  assign n893 = ~n1361 & ~n1362;
  assign n894 = n647 & n1340;
  assign n895 = ~n163 & n894;
  assign n896 = n1327 & n1340;
  assign n897 = ~n1363 & ~n1364;
  assign n898 = ~n871 & ~n1363;
  assign n899 = ~n1364 & n898;
  assign n900 = ~n871 & n897;
  assign n901 = ~n866 & n1365;
  assign n902 = ~n860 & n1365;
  assign n903 = ~n866 & n902;
  assign n904 = ~n860 & n901;
  assign n905 = ~n844 & n1366;
  assign n906 = ~n830 & n905;
  assign n907 = ~n1362 & ~n1364;
  assign n908 = ~n860 & n907;
  assign n909 = ~n1361 & n908;
  assign n910 = ~n844 & n909;
  assign n911 = ~n866 & n910;
  assign n912 = ~n786 & n911;
  assign n913 = ~n830 & n912;
  assign n914 = ~n871 & n913;
  assign n915 = ~n786 & n906;
  assign n916 = pi13 & ~n1367;
  assign n917 = n1330 & n916;
  assign n918 = n1330 & ~n1367;
  assign n919 = ~n1330 & n1367;
  assign n920 = pi13 & ~n919;
  assign n921 = ~n1330 & n916;
  assign n922 = n1330 & ~n916;
  assign n923 = ~n921 & ~n922;
  assign n924 = ~n1368 & n920;
  assign n925 = pi08 & n71;
  assign n926 = n47 & n71;
  assign n927 = pi13 & n926;
  assign n928 = pi13 & n71;
  assign n929 = n47 & n928;
  assign n930 = n29 & n925;
  assign n931 = ~pi13 & n25;
  assign n932 = n25 & n251;
  assign n933 = ~pi13 & n932;
  assign n934 = n251 & n931;
  assign n935 = ~n1370 & ~n1371;
  assign n936 = n41 & n737;
  assign n937 = ~pi11 & ~n64;
  assign n938 = po5 & ~n937;
  assign n939 = n65 & n701;
  assign n940 = pi09 & ~n939;
  assign n941 = pi09 & ~n938;
  assign n942 = ~n939 & n941;
  assign n943 = ~n938 & n940;
  assign n944 = ~n936 & n1372;
  assign n945 = ~n64 & ~n925;
  assign n946 = n1340 & ~n945;
  assign n947 = ~pi07 & n130;
  assign n948 = ~pi09 & ~n947;
  assign n949 = ~n946 & n948;
  assign n950 = ~n938 & ~n939;
  assign n951 = ~n936 & n950;
  assign n952 = pi09 & ~n951;
  assign n953 = ~n946 & ~n947;
  assign n954 = ~pi09 & ~n953;
  assign n955 = ~n952 & ~n954;
  assign n956 = ~n944 & ~n949;
  assign n957 = ~pi09 & ~n35;
  assign n958 = pi10 & pi11;
  assign n959 = ~n85 & ~n958;
  assign n960 = ~pi09 & ~n959;
  assign n961 = ~n182 & n957;
  assign n962 = pi07 & n85;
  assign n963 = ~n1374 & ~n962;
  assign n964 = ~n1340 & ~n963;
  assign n965 = ~pi07 & ~pi09;
  assign n966 = n143 & ~n965;
  assign n967 = n882 & ~n966;
  assign n968 = pi11 & n182;
  assign n969 = ~pi03 & ~pi09;
  assign n970 = ~pi03 & n968;
  assign n971 = ~pi09 & n970;
  assign n972 = ~pi03 & n42;
  assign n973 = n182 & n972;
  assign n974 = n968 & n969;
  assign n975 = ~n26 & ~n1375;
  assign n976 = ~n36 & ~n776;
  assign n977 = pi07 & pi11;
  assign n978 = ~n976 & n977;
  assign n979 = pi07 & ~n975;
  assign n980 = pi03 & ~n966;
  assign n981 = pi07 & ~n976;
  assign n982 = ~n980 & ~n981;
  assign n983 = pi11 & ~n982;
  assign n984 = ~n967 & ~n1376;
  assign n985 = ~n964 & ~n1377;
  assign n986 = n1373 & ~n1376;
  assign n987 = ~n964 & n986;
  assign n988 = ~n967 & n987;
  assign n989 = ~n954 & n985;
  assign n990 = ~n952 & n989;
  assign n991 = n1373 & n985;
  assign n992 = ~pi13 & ~n1378;
  assign n993 = n935 & ~n992;
  assign n994 = n1369 & n993;
  assign n995 = ~pi03 & n1348;
  assign n996 = ~n746 & ~n995;
  assign n997 = pi03 & ~n1348;
  assign n998 = ~n996 & ~n997;
  assign n999 = ~pi08 & ~n998;
  assign n1000 = ~n798 & n800;
  assign n1001 = ~n749 & ~n1352;
  assign n1002 = n1340 & ~n1001;
  assign n1003 = n1340 & n1352;
  assign n1004 = n749 & n1352;
  assign n1005 = pi08 & ~n1004;
  assign n1006 = ~n1380 & n1005;
  assign n1007 = ~n749 & ~n1380;
  assign n1008 = ~n1340 & ~n1352;
  assign n1009 = ~n1007 & ~n1008;
  assign n1010 = ~n810 & n1352;
  assign n1011 = ~n1379 & ~n1381;
  assign n1012 = n251 & ~n1011;
  assign n1013 = pi10 & ~n836;
  assign n1014 = n47 & ~n1013;
  assign n1015 = n47 & n836;
  assign n1016 = ~n1012 & ~n1382;
  assign n1017 = ~pi11 & ~n1016;
  assign n1018 = n169 & ~n751;
  assign n1019 = ~n746 & n1018;
  assign n1020 = ~n746 & ~n751;
  assign n1021 = ~n737 & ~n1356;
  assign n1022 = ~n355 & ~n735;
  assign n1023 = ~n735 & n1356;
  assign n1024 = ~n737 & ~n1023;
  assign n1025 = ~n355 & ~n1024;
  assign n1026 = ~n1021 & n1022;
  assign n1027 = ~po5 & n1345;
  assign n1028 = n1267 & ~n701;
  assign n1029 = ~n701 & ~n1345;
  assign n1030 = ~po5 & ~n1029;
  assign n1031 = n1267 & ~n1030;
  assign n1032 = ~n1027 & n1028;
  assign n1033 = ~n1344 & ~n1385;
  assign n1034 = ~n1344 & ~n1384;
  assign n1035 = ~n1385 & n1034;
  assign n1036 = ~n1384 & n1033;
  assign n1037 = ~n1383 & n1386;
  assign n1038 = pi11 & ~n1037;
  assign n1039 = ~n65 & ~n182;
  assign n1040 = pi09 & ~n1039;
  assign n1041 = ~n156 & ~n1260;
  assign n1042 = n647 & n1387;
  assign n1043 = n894 & n1387;
  assign n1044 = n1340 & n1042;
  assign n1045 = ~n1038 & ~n1388;
  assign n1046 = ~n1017 & n1045;
  assign n1047 = ~n1368 & ~n1017;
  assign n1048 = ~n1038 & n1047;
  assign n1049 = ~n1388 & n1048;
  assign n1050 = ~n1368 & n1046;
  assign po6 = pi13 & ~n1389;
  assign n1052 = ~n1294 & n1329;
  assign n1053 = pi13 & ~n1330;
  assign n1054 = pi13 & ~n1052;
  assign n1055 = ~n1330 & n1054;
  assign n1056 = ~n1294 & n676;
  assign n1057 = n1294 & ~n676;
  assign n1058 = ~n1056 & ~n1057;
  assign n1059 = ~n1052 & n1053;
  assign n1060 = n481 & ~n945;
  assign n1061 = ~pi06 & n130;
  assign n1062 = ~n1060 & ~n1061;
  assign n1063 = ~pi09 & ~n1062;
  assign n1064 = pi02 & pi09;
  assign n1065 = pi02 & n1265;
  assign n1066 = pi02 & n41;
  assign n1067 = pi09 & n1066;
  assign n1068 = n41 & n1064;
  assign n1069 = pi06 & n85;
  assign n1070 = ~n1391 & ~n1069;
  assign n1071 = ~n1374 & ~n1391;
  assign n1072 = ~n1069 & n1071;
  assign n1073 = ~n1374 & ~n1069;
  assign n1074 = ~n1391 & n1073;
  assign n1075 = ~n1374 & n1070;
  assign n1076 = ~n481 & ~n1392;
  assign n1077 = n470 & ~n937;
  assign n1078 = n65 & n474;
  assign n1079 = ~n1077 & ~n1078;
  assign n1080 = pi09 & ~n1079;
  assign n1081 = n143 & ~n485;
  assign n1082 = n593 & ~n1081;
  assign n1083 = ~pi02 & n42;
  assign n1084 = ~pi02 & n968;
  assign n1085 = ~pi09 & n1084;
  assign n1086 = ~pi02 & ~pi09;
  assign n1087 = n968 & n1086;
  assign n1088 = n182 & n1083;
  assign n1089 = ~n26 & ~n1393;
  assign n1090 = pi06 & ~n1089;
  assign n1091 = ~n1082 & ~n1090;
  assign n1092 = ~n1080 & ~n1082;
  assign n1093 = ~n1090 & n1092;
  assign n1094 = ~n1080 & n1091;
  assign n1095 = ~n1076 & n1394;
  assign n1096 = n85 & ~n481;
  assign n1097 = n1089 & ~n1096;
  assign n1098 = pi06 & ~n1097;
  assign n1099 = ~n481 & ~n1071;
  assign n1100 = n1092 & ~n1099;
  assign n1101 = ~n1063 & n1100;
  assign n1102 = ~n1098 & n1101;
  assign n1103 = ~n1063 & ~n1080;
  assign n1104 = ~n1090 & n1103;
  assign n1105 = ~n1076 & n1104;
  assign n1106 = ~n1082 & n1105;
  assign n1107 = ~n1063 & n1095;
  assign n1108 = ~pi13 & ~n1395;
  assign n1109 = n935 & ~n1108;
  assign n1110 = ~n1390 & n1109;
  assign n1111 = ~n1271 & n1293;
  assign n1112 = pi13 & ~n1111;
  assign n1113 = ~n1271 & n429;
  assign n1114 = n1271 & ~n429;
  assign n1115 = ~n1113 & ~n1114;
  assign n1116 = ~n1294 & n1112;
  assign n1117 = n1277 & ~n945;
  assign n1118 = ~n130 & ~n448;
  assign n1119 = ~pi05 & ~n1118;
  assign n1120 = n253 & n968;
  assign n1121 = ~pi09 & ~n1120;
  assign n1122 = ~n1119 & n1121;
  assign n1123 = ~n1117 & n1122;
  assign n1124 = pi05 & n25;
  assign n1125 = n242 & ~n937;
  assign n1126 = pi01 & ~n937;
  assign n1127 = ~n25 & ~n1126;
  assign n1128 = pi05 & ~n1127;
  assign n1129 = ~n1124 & ~n1125;
  assign n1130 = n65 & n258;
  assign n1131 = pi09 & ~n1130;
  assign n1132 = ~n1397 & n1131;
  assign n1133 = ~pi05 & n130;
  assign n1134 = pi11 & n255;
  assign n1135 = ~n1120 & ~n1134;
  assign n1136 = ~n1119 & ~n1120;
  assign n1137 = ~n1133 & n1135;
  assign n1138 = ~n1117 & ~n1133;
  assign n1139 = n1135 & n1138;
  assign n1140 = ~n1117 & n1398;
  assign n1141 = ~pi09 & ~n1399;
  assign n1142 = ~n1125 & ~n1130;
  assign n1143 = ~n1124 & n1142;
  assign n1144 = ~n1397 & ~n1130;
  assign n1145 = pi09 & ~n1400;
  assign n1146 = ~n1141 & ~n1145;
  assign n1147 = ~n1123 & ~n1132;
  assign n1148 = pi05 & n85;
  assign n1149 = ~n1374 & ~n1148;
  assign n1150 = ~n1277 & ~n1149;
  assign n1151 = n1265 & ~n1277;
  assign n1152 = ~n145 & ~n1151;
  assign n1153 = pi01 & ~n1152;
  assign n1154 = ~n1150 & ~n1153;
  assign n1155 = ~n1145 & ~n1150;
  assign n1156 = n1401 & ~n1150;
  assign n1157 = ~n1141 & n1155;
  assign n1158 = ~n1153 & n1402;
  assign n1159 = ~n1153 & n1155;
  assign n1160 = ~n1141 & n1159;
  assign n1161 = n1401 & n1154;
  assign n1162 = ~pi13 & ~n1403;
  assign n1163 = n935 & ~n1162;
  assign n1164 = n1396 & n1163;
  assign n1165 = pi12 & n1269;
  assign n1166 = pi13 & ~n1271;
  assign n1167 = pi12 & n239;
  assign n1168 = ~pi12 & ~n239;
  assign n1169 = ~n1167 & ~n1168;
  assign n1170 = pi13 & ~n1169;
  assign n1171 = ~n1165 & n1166;
  assign n1172 = n1251 & ~n945;
  assign n1173 = ~pi00 & ~n182;
  assign n1174 = pi11 & ~n1249;
  assign n1175 = n93 & n968;
  assign n1176 = pi11 & n94;
  assign n1177 = ~n1175 & ~n1176;
  assign n1178 = ~n1173 & n1174;
  assign n1179 = ~pi04 & n130;
  assign n1180 = ~pi09 & ~n1179;
  assign n1181 = n1405 & n1180;
  assign n1182 = ~n1172 & n1181;
  assign n1183 = n41 & n1252;
  assign n1184 = ~pi00 & ~n25;
  assign n1185 = pi04 & ~n937;
  assign n1186 = ~n1184 & n1185;
  assign n1187 = n65 & n70;
  assign n1188 = pi09 & ~n1187;
  assign n1189 = ~n1186 & n1188;
  assign n1190 = ~n1183 & n1189;
  assign n1191 = ~n1182 & ~n1190;
  assign n1192 = pi04 & n85;
  assign n1193 = ~n1374 & ~n1192;
  assign n1194 = ~n1251 & ~n1193;
  assign n1195 = ~n143 & n152;
  assign n1196 = ~n1194 & ~n1195;
  assign n1197 = n23 & ~n937;
  assign n1198 = pi04 & n25;
  assign n1199 = ~n1187 & ~n1198;
  assign n1200 = ~n1186 & ~n1187;
  assign n1201 = ~n1197 & n1199;
  assign n1202 = ~n1183 & ~n1197;
  assign n1203 = n1199 & n1202;
  assign n1204 = ~n1183 & n1406;
  assign n1205 = pi09 & ~n1407;
  assign n1206 = ~n1176 & ~n1179;
  assign n1207 = n1405 & ~n1179;
  assign n1208 = ~n1175 & n1206;
  assign n1209 = ~n1172 & ~n1179;
  assign n1210 = n1405 & n1209;
  assign n1211 = ~n1172 & n1408;
  assign n1212 = ~pi09 & ~n1409;
  assign n1213 = ~n1195 & ~n1212;
  assign n1214 = ~n1205 & n1213;
  assign n1215 = ~n1194 & n1214;
  assign n1216 = n1196 & ~n1212;
  assign n1217 = ~n1205 & n1216;
  assign n1218 = ~n1191 & n1196;
  assign n1219 = ~pi13 & ~n1410;
  assign n1220 = n935 & ~n1219;
  assign n1221 = ~n1404 & n1220;
  assign n1222 = n1249 & n1325;
  assign n1223 = ~po5 & ~n701;
  assign n1224 = ~n242 & ~n258;
  assign n1225 = ~n1223 & ~n1224;
  assign n1226 = n397 & n470;
  assign n1227 = ~pi06 & n584;
  assign n1228 = ~n1226 & ~n1227;
  assign n1229 = ~pi04 & ~pi05;
  assign n1230 = ~pi05 & ~n1228;
  assign n1231 = ~pi04 & n1230;
  assign n1232 = ~n1228 & n1229;
  assign n1233 = n1249 & n242;
  assign n1234 = ~n399 & ~n1233;
  assign n1235 = n1325 & ~n1234;
  assign n1236 = ~n1411 & ~n1235;
  assign n1237 = ~n1223 & ~n1236;
  assign n1238 = n1222 & n1225;
  assign n1239 = n30 | n31;
  assign n1240 = n32 | n33;
  assign n1241 = n39 | n40;
  assign n1242 = n45 | n46;
  assign n1243 = n54 | n51 | n53;
  assign n1244 = n60 | n61;
  assign n1245 = n66 | n67;
  assign n1246 = n78 | n79;
  assign n1247 = n83 | n84;
  assign n1248 = n90 | n87 | n89;
  assign n1249 = n95 | ~n96;
  assign n1250 = n103 | n101 | n102;
  assign n1251 = n115 | n110 | n114;
  assign n1252 = n119 | n120;
  assign n1253 = n126 | n127;
  assign n1254 = n132 | n133;
  assign n1255 = n136 | n137;
  assign n1256 = n138 | n139;
  assign n1257 = n141 | n142;
  assign n1258 = n149 | n146 | n148;
  assign n1259 = n157 | n158;
  assign n1260 = n162 | n160 | n161;
  assign n1261 = n171 | n168 | n170;
  assign n1262 = n173 | n174;
  assign n1263 = n176 | n177;
  assign n1264 = n200 | n194 | n199;
  assign n1265 = n201 | n202;
  assign n1266 = n204 | n205;
  assign n1267 = n206 | n207;
  assign n1268 = n209 | n210;
  assign n1269 = n237 | n229 | n236;
  assign n1270 = n234 | n235;
  assign n1271 = n240 | n241;
  assign n1272 = n246 | n247;
  assign n1273 = n265 | n266;
  assign n1274 = n269 | n270;
  assign n1275 = n276 | n277;
  assign n1276 = n278 | n279;
  assign n1277 = n281 | n282;
  assign n1278 = n284 | n285;
  assign n1279 = n299 | n300;
  assign n1280 = n302 | n303;
  assign n1281 = n312 | ~n313;
  assign n1282 = n320 | n321;
  assign n1283 = n329 | ~n330;
  assign n1284 = n333 | n334;
  assign n1285 = n342 | ~n343;
  assign n1286 = n353 | n348 | n352;
  assign n1287 = n361 | ~n362;
  assign n1288 = n365 | n366;
  assign n1289 = n376 | ~n377;
  assign n1290 = n388 | n385 | n387;
  assign n1291 = n409 | n410;
  assign n1292 = n417 | n418;
  assign n1293 = n427 | n428;
  assign n1294 = n430 | n431;
  assign n1295 = n434 | ~n435;
  assign n1296 = n441 | n438 | n440;
  assign n1297 = n444 | n445;
  assign n1298 = n456 | n457;
  assign n1299 = n462 | n460 | n461;
  assign n1300 = n465 | n466;
  assign n1301 = n468 | n469;
  assign n1302 = n479 | n480;
  assign n1303 = n497 | n498;
  assign n1304 = n500 | n501;
  assign n1305 = n519 | n514 | n518;
  assign n1306 = n525 | n526;
  assign n1307 = n531 | ~n532;
  assign n1308 = n535 | n536;
  assign n1309 = n559 | n548 | n558;
  assign n1310 = n553 | ~n554;
  assign n1311 = n561 | n562;
  assign n1312 = ~n570 | n565 | ~n569;
  assign n1313 = n573 | n574;
  assign n1314 = n581 | n582;
  assign n1315 = n587 | n588;
  assign n1316 = n597 | n598;
  assign n1317 = n600 | n601;
  assign n1318 = n605 | n602 | n604;
  assign n1319 = n609 | n610;
  assign n1320 = n613 | n614;
  assign n1321 = n619 | n620;
  assign n1322 = n621 | n622;
  assign n1323 = n627 | n628;
  assign n1324 = n631 | ~n632;
  assign n1325 = n638 | ~n639;
  assign n1326 = n645 | n646;
  assign n1327 = n648 | n649;
  assign n1328 = n662 | n663;
  assign n1329 = n674 | n675;
  assign n1330 = n677 | n678;
  assign n1331 = n682 | n683;
  assign n1332 = n685 | n686;
  assign n1333 = n691 | n692;
  assign n1334 = n696 | n697;
  assign n1335 = n704 | n705;
  assign n1336 = n713 | n710 | n712;
  assign n1337 = n716 | n717;
  assign n1338 = n720 | n721;
  assign n1339 = n728 | n729;
  assign n1340 = n733 | n734;
  assign n1341 = n743 | n744;
  assign n1342 = n761 | ~n762;
  assign n1343 = n766 | n767;
  assign n1344 = n770 | n771;
  assign n1345 = n774 | ~n775;
  assign n1346 = n777 | n778;
  assign n1347 = n783 | n780 | n782;
  assign n1348 = n796 | n791 | n795;
  assign n1349 = n803 | ~n804;
  assign n1350 = n809 | n806 | n808;
  assign n1351 = n814 | ~n815;
  assign n1352 = n819 | n820;
  assign n1353 = n827 | n828;
  assign n1354 = n833 | n834;
  assign n1355 = n842 | n843;
  assign n1356 = ~n851 | n847 | ~n850;
  assign n1357 = n856 | ~n857;
  assign n1358 = n863 | n864;
  assign n1359 = n869 | ~n870;
  assign n1360 = n874 | n875;
  assign n1361 = n880 | n881;
  assign n1362 = n885 | n886;
  assign n1363 = n892 | ~n893;
  assign n1364 = n895 | n896;
  assign n1365 = n899 | n900;
  assign n1366 = n903 | n904;
  assign n1367 = n914 | n915;
  assign n1368 = n917 | n918;
  assign n1369 = n923 | ~n924;
  assign n1370 = n930 | n927 | n929;
  assign n1371 = n933 | n934;
  assign n1372 = n942 | n943;
  assign n1373 = n955 | ~n956;
  assign n1374 = n960 | n961;
  assign n1375 = n974 | n971 | n973;
  assign n1376 = n978 | n979;
  assign n1377 = n983 | ~n984;
  assign n1378 = n991 | n988 | n990;
  assign n1379 = n999 | n1000;
  assign n1380 = n1002 | n1003;
  assign n1381 = ~n1010 | n1006 | ~n1009;
  assign n1382 = n1014 | n1015;
  assign n1383 = n1019 | n1020;
  assign n1384 = n1025 | n1026;
  assign n1385 = n1031 | n1032;
  assign n1386 = n1035 | n1036;
  assign n1387 = n1040 | ~n1041;
  assign n1388 = n1043 | n1044;
  assign n1389 = n1049 | n1050;
  assign n1390 = n1059 | n1055 | ~n1058;
  assign n1391 = n1068 | n1065 | n1067;
  assign n1392 = n1075 | n1072 | n1074;
  assign n1393 = n1088 | n1085 | n1087;
  assign n1394 = n1093 | n1094;
  assign n1395 = n1107 | n1102 | n1106;
  assign n1396 = n1115 | ~n1116;
  assign n1397 = n1128 | ~n1129;
  assign n1398 = n1136 | n1137;
  assign n1399 = n1139 | n1140;
  assign n1400 = n1143 | n1144;
  assign n1401 = n1146 | ~n1147;
  assign n1402 = n1156 | n1157;
  assign n1403 = n1161 | n1158 | n1160;
  assign n1404 = n1170 | n1171;
  assign n1405 = n1177 | ~n1178;
  assign n1406 = n1200 | n1201;
  assign n1407 = n1203 | n1204;
  assign n1408 = n1207 | n1208;
  assign n1409 = n1210 | n1211;
  assign n1410 = n1218 | n1215 | n1217;
  assign n1411 = n1231 | n1232;
  assign po7 = n1237 | n1238;
  assign po0 = ~n1221;
  assign po1 = ~n1164;
  assign po2 = ~n1110;
  assign po3 = ~n994;
  assign po4 = ~n1223;
endmodule
