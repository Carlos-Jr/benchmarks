module alu4_cl ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13,
    po0, po1, po2, po3, po4, po5, po6, po7  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13;
  output po0, po1, po2, po3, po4, po5, po6, po7;
  wire n23, n24, n25, n26, n27, n28, n29,
    n30, n31, n32, n33, n34, n35, n36, n37,
    n38, n39, n40, n41, n42, n43, n44, n45,
    n46, n47, n48, n49, n50, n51, n52, n53,
    n54, n55, n56, n57, n58, n59, n60, n61,
    n62, n63, n64, n65, n66, n67, n68, n69,
    n70, n71, n72, n73, n74, n75, n76, n77,
    n78, n79, n80, n81, n82, n83, n84, n85,
    n86, n87, n88, n89, n90, n91, n92, n93,
    n94, n95, n96, n97, n98, n99, n100,
    n101, n102, n103, n104, n105, n106, n107,
    n108, n109, n110, n111, n112, n113, n114,
    n115, n116, n117, n118, n119, n120, n121,
    n122, n123, n124, n125, n126, n127, n128,
    n129, n130, n131, n132, n133, n134, n135,
    n136, n137, n138, n139, n140, n141, n142,
    n143, n144, n145, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156,
    n157, n158, n159, n160, n161, n162, n163,
    n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177,
    n178, n179, n180, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192,
    n193, n194, n195, n196, n197, n198, n199,
    n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213,
    n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227,
    n228, n229, n230, n231, n232, n233, n234,
    n235, n236, n237, n238, n239, n240, n241,
    n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n332, n333,
    n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403,
    n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416, n417,
    n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438,
    n439, n440, n441, n442, n443, n444, n445,
    n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n484, n485, n486, n487, n488,
    n489, n490, n491, n492, n493, n494, n495,
    n496, n497, n498, n499, n501, n502, n503,
    n504, n505, n506, n507, n508, n509, n510,
    n511, n512, n513, n514, n515, n516, n517,
    n518, n519, n520, n521, n522, n523, n524,
    n525, n526, n527, n528, n529, n530, n531,
    n532, n533, n534, n535, n536, n537, n538,
    n539, n540, n541, n542, n543, n544, n545,
    n546, n547, n548, n549, n550, n551, n552,
    n553, n554, n555, n556, n557, n558, n559,
    n560, n561, n562, n563, n564, n565, n566,
    n567, n568, n569, n570, n571, n572, n573,
    n574, n575, n576, n577, n578, n579, n580,
    n581, n582, n583, n584, n585, n586, n587,
    n588, n589, n590, n591, n592, n593, n594,
    n595, n596, n597, n598, n599, n600, n601,
    n602, n603, n604, n605, n606, n607, n608,
    n609, n610, n611, n612, n613, n614, n615,
    n616, n617, n618, n619, n620, n621, n622,
    n623, n624, n625, n626, n627, n628, n629,
    n630, n631, n632, n633, n634, n635, n636,
    n637, n638, n641, n642, n643, n644, n645,
    n646, n647, n648, n649, n650, n651, n652,
    n653, n654, n655, n656, n657, n658, n659,
    n660, n661, n662, n663, n664, n665, n666,
    n667, n668, n669, n670, n671, n673, n674;
  assign n23 = pi00 & pi11;
  assign n24 = ~pi08 & ~pi09;
  assign n25 = ~pi10 & ~n24;
  assign n26 = n23 & ~n25;
  assign n27 = pi09 & pi11;
  assign n28 = ~pi10 & ~pi13;
  assign n29 = ~n27 & n28;
  assign n30 = ~pi08 & n29;
  assign n31 = ~pi00 & n30;
  assign n32 = ~pi00 & ~pi04;
  assign n33 = pi08 & ~pi09;
  assign n34 = ~pi10 & ~pi11;
  assign n35 = ~pi13 & ~n34;
  assign n36 = ~pi10 & pi13;
  assign n37 = n33 & ~n36;
  assign n38 = ~n35 & n37;
  assign n39 = ~n32 & n38;
  assign n40 = ~pi09 & pi11;
  assign n41 = pi08 & pi10;
  assign n42 = ~pi13 & n40;
  assign n43 = n41 & n42;
  assign n44 = pi10 & ~pi11;
  assign n45 = ~pi08 & pi09;
  assign n46 = pi13 & n45;
  assign n47 = ~n44 & n46;
  assign n48 = pi08 & pi09;
  assign n49 = n44 & n48;
  assign n50 = ~n43 & ~n49;
  assign n51 = ~n47 & n50;
  assign n52 = ~pi04 & ~n51;
  assign n53 = ~n24 & ~n48;
  assign n54 = ~pi10 & pi11;
  assign n55 = ~n53 & n54;
  assign n56 = pi13 & n55;
  assign n57 = ~pi09 & ~pi11;
  assign n58 = ~pi08 & pi10;
  assign n59 = n57 & n58;
  assign n60 = ~n56 & ~n59;
  assign n61 = pi00 & pi04;
  assign n62 = ~n60 & n61;
  assign n63 = ~n32 & ~n61;
  assign n64 = ~pi00 & ~n44;
  assign n65 = n46 & n63;
  assign n66 = ~n64 & n65;
  assign n67 = ~n39 & ~n66;
  assign n68 = ~n52 & n67;
  assign n69 = ~n62 & n68;
  assign n70 = ~n31 & n69;
  assign n71 = ~pi08 & ~pi10;
  assign n72 = pi04 & n71;
  assign n73 = pi08 & ~pi10;
  assign n74 = ~pi09 & ~n44;
  assign n75 = ~n73 & n74;
  assign n76 = ~n72 & ~n75;
  assign n77 = ~n70 & ~n76;
  assign n78 = ~pi11 & ~n58;
  assign n79 = ~pi08 & pi11;
  assign n80 = ~pi00 & ~n79;
  assign n81 = pi04 & ~n78;
  assign n82 = ~n80 & n81;
  assign n83 = ~pi08 & n44;
  assign n84 = n32 & n83;
  assign n85 = pi00 & ~n69;
  assign n86 = n41 & n85;
  assign n87 = pi09 & ~n84;
  assign n88 = ~n82 & n87;
  assign n89 = ~n86 & n88;
  assign n90 = ~pi00 & pi04;
  assign n91 = pi11 & n73;
  assign n92 = n90 & n91;
  assign n93 = pi08 & n34;
  assign n94 = ~n58 & ~n93;
  assign n95 = n70 & ~n94;
  assign n96 = pi08 & n44;
  assign n97 = ~n23 & ~n96;
  assign n98 = ~pi04 & ~n97;
  assign n99 = ~pi09 & ~n92;
  assign n100 = ~n98 & n99;
  assign n101 = ~n95 & n100;
  assign n102 = ~n89 & ~n101;
  assign n103 = ~n26 & ~n77;
  assign n104 = ~n102 & n103;
  assign n105 = ~pi13 & ~n104;
  assign n106 = pi09 & pi13;
  assign n107 = n93 & n106;
  assign n108 = ~pi09 & pi10;
  assign n109 = ~pi13 & n79;
  assign n110 = n108 & n109;
  assign n111 = ~n107 & ~n110;
  assign n112 = pi10 & n48;
  assign n113 = ~pi00 & pi11;
  assign n114 = n112 & n113;
  assign n115 = pi04 & n73;
  assign n116 = ~pi00 & n70;
  assign n117 = ~pi08 & pi13;
  assign n118 = n27 & n117;
  assign n119 = ~n116 & n118;
  assign n120 = pi13 & n44;
  assign n121 = n24 & n70;
  assign n122 = n33 & n61;
  assign n123 = n48 & n85;
  assign n124 = ~n121 & ~n122;
  assign n125 = ~n123 & n124;
  assign n126 = n120 & ~n125;
  assign n127 = ~n119 & ~n126;
  assign n128 = pi00 & ~pi08;
  assign n129 = n127 & n128;
  assign n130 = ~n115 & ~n129;
  assign n131 = n57 & ~n130;
  assign n132 = ~pi00 & n59;
  assign n133 = n46 & n54;
  assign n134 = n61 & n133;
  assign n135 = n33 & n120;
  assign n136 = n127 & n135;
  assign n137 = ~n134 & ~n136;
  assign n138 = n45 & n54;
  assign n139 = n137 & n138;
  assign n140 = ~n127 & ~n132;
  assign n141 = ~n139 & n140;
  assign n142 = ~n137 & n138;
  assign n143 = ~n49 & n127;
  assign n144 = ~n142 & n143;
  assign n145 = ~n141 & ~n144;
  assign n146 = ~n25 & n113;
  assign n147 = n33 & n44;
  assign n148 = n137 & n147;
  assign n149 = ~n70 & ~n146;
  assign n150 = ~n148 & n149;
  assign n151 = n48 & n54;
  assign n152 = n44 & n45;
  assign n153 = ~n151 & ~n152;
  assign n154 = n23 & ~n48;
  assign n155 = pi08 & n57;
  assign n156 = ~n137 & n155;
  assign n157 = ~n154 & ~n156;
  assign n158 = pi10 & ~n157;
  assign n159 = n70 & n153;
  assign n160 = ~n158 & n159;
  assign n161 = ~n150 & ~n160;
  assign n162 = ~pi09 & n73;
  assign n163 = n63 & n162;
  assign n164 = pi09 & ~n70;
  assign n165 = ~pi00 & ~n164;
  assign n166 = ~pi09 & n70;
  assign n167 = pi11 & ~n166;
  assign n168 = n71 & ~n165;
  assign n169 = ~n167 & n168;
  assign n170 = ~n114 & ~n163;
  assign n171 = ~n169 & n170;
  assign n172 = ~n131 & n171;
  assign n173 = ~n145 & n172;
  assign n174 = ~n161 & n173;
  assign n175 = pi12 & n174;
  assign n176 = ~pi12 & pi13;
  assign n177 = ~n174 & n176;
  assign n178 = pi13 & ~n175;
  assign n179 = ~n177 & n178;
  assign n180 = ~n105 & n111;
  assign po0 = n179 | ~n180;
  assign n182 = ~pi01 & pi05;
  assign n183 = n91 & n182;
  assign n184 = n23 & n108;
  assign n185 = ~pi01 & ~pi05;
  assign n186 = n90 & n185;
  assign n187 = ~pi01 & ~n44;
  assign n188 = pi01 & pi05;
  assign n189 = ~n185 & ~n188;
  assign n190 = ~n90 & ~n187;
  assign n191 = n189 & n190;
  assign n192 = ~n186 & ~n191;
  assign n193 = pi09 & ~n192;
  assign n194 = ~n184 & ~n193;
  assign n195 = n117 & ~n194;
  assign n196 = n38 & ~n185;
  assign n197 = ~pi01 & n30;
  assign n198 = ~pi05 & ~n51;
  assign n199 = ~pi09 & n44;
  assign n200 = pi13 & n199;
  assign n201 = n60 & ~n200;
  assign n202 = ~pi08 & n90;
  assign n203 = n120 & n202;
  assign n204 = n201 & ~n203;
  assign n205 = n188 & ~n204;
  assign n206 = ~n196 & ~n197;
  assign n207 = ~n198 & n206;
  assign n208 = ~n195 & n207;
  assign n209 = ~n205 & n208;
  assign n210 = ~n94 & n209;
  assign n211 = pi01 & pi11;
  assign n212 = ~n96 & ~n211;
  assign n213 = ~pi05 & ~n212;
  assign n214 = ~n183 & ~n213;
  assign n215 = ~n210 & n214;
  assign n216 = ~pi09 & ~n215;
  assign n217 = n83 & n185;
  assign n218 = ~pi01 & ~n79;
  assign n219 = pi05 & ~n78;
  assign n220 = ~n218 & n219;
  assign n221 = ~n217 & ~n220;
  assign n222 = pi09 & ~n221;
  assign n223 = pi11 & ~n25;
  assign n224 = n112 & ~n209;
  assign n225 = ~n223 & ~n224;
  assign n226 = pi01 & ~n225;
  assign n227 = pi05 & n71;
  assign n228 = ~n75 & ~n227;
  assign n229 = ~n209 & ~n228;
  assign n230 = ~n222 & ~n229;
  assign n231 = ~n216 & n230;
  assign n232 = ~n226 & n231;
  assign n233 = ~pi13 & ~n232;
  assign n234 = pi05 & n73;
  assign n235 = ~n70 & ~n137;
  assign n236 = n133 & n188;
  assign n237 = ~pi01 & n209;
  assign n238 = n118 & ~n237;
  assign n239 = pi09 & n209;
  assign n240 = ~pi05 & ~pi09;
  assign n241 = pi01 & pi08;
  assign n242 = ~n240 & n241;
  assign n243 = ~pi08 & n209;
  assign n244 = ~n242 & ~n243;
  assign n245 = n120 & ~n239;
  assign n246 = ~n244 & n245;
  assign n247 = ~n238 & ~n246;
  assign n248 = n135 & n247;
  assign n249 = ~n236 & ~n248;
  assign n250 = n235 & ~n249;
  assign n251 = ~n235 & n249;
  assign n252 = ~n250 & ~n251;
  assign n253 = n209 & ~n252;
  assign n254 = ~n209 & n252;
  assign n255 = n41 & ~n253;
  assign n256 = ~n254 & n255;
  assign n257 = pi00 & ~n127;
  assign n258 = n247 & ~n257;
  assign n259 = ~n127 & ~n247;
  assign n260 = pi00 & n259;
  assign n261 = ~n258 & ~n260;
  assign n262 = pi01 & ~pi08;
  assign n263 = ~n261 & n262;
  assign n264 = ~n234 & ~n263;
  assign n265 = ~n256 & n264;
  assign n266 = n57 & ~n265;
  assign n267 = n127 & n247;
  assign n268 = ~n259 & ~n267;
  assign n269 = n112 & ~n268;
  assign n270 = pi09 & n71;
  assign n271 = ~n209 & n270;
  assign n272 = ~n269 & ~n271;
  assign n273 = ~pi11 & ~n272;
  assign n274 = ~pi05 & ~n61;
  assign n275 = n162 & n274;
  assign n276 = n85 & ~n209;
  assign n277 = ~n85 & n209;
  assign n278 = ~n276 & ~n277;
  assign n279 = pi10 & ~n48;
  assign n280 = ~n24 & ~n279;
  assign n281 = ~n44 & ~n280;
  assign n282 = ~n278 & n281;
  assign n283 = n23 & n112;
  assign n284 = n34 & ~n48;
  assign n285 = ~n275 & ~n284;
  assign n286 = ~n283 & n285;
  assign n287 = ~n282 & n286;
  assign n288 = pi01 & ~n287;
  assign n289 = ~pi00 & ~pi01;
  assign n290 = n112 & n289;
  assign n291 = n61 & n185;
  assign n292 = n162 & n291;
  assign n293 = ~n290 & ~n292;
  assign n294 = pi11 & ~n293;
  assign n295 = n70 & n209;
  assign n296 = ~n153 & n295;
  assign n297 = ~n61 & ~n182;
  assign n298 = n61 & ~n188;
  assign n299 = n162 & ~n297;
  assign n300 = ~n298 & n299;
  assign n301 = ~pi11 & n45;
  assign n302 = ~n151 & ~n301;
  assign n303 = ~n70 & ~n302;
  assign n304 = ~n209 & n303;
  assign n305 = pi11 & ~n280;
  assign n306 = n278 & n305;
  assign n307 = n59 & n261;
  assign n308 = ~n306 & ~n307;
  assign n309 = ~pi01 & ~n308;
  assign n310 = ~n127 & n134;
  assign n311 = ~n249 & n310;
  assign n312 = n249 & ~n310;
  assign n313 = ~n311 & ~n312;
  assign n314 = ~n247 & n313;
  assign n315 = n247 & ~n313;
  assign n316 = n138 & ~n314;
  assign n317 = ~n315 & n316;
  assign n318 = ~n294 & ~n300;
  assign n319 = ~n304 & n318;
  assign n320 = ~n296 & n319;
  assign n321 = ~n288 & n320;
  assign n322 = ~n273 & n321;
  assign n323 = ~n309 & n322;
  assign n324 = ~n317 & n323;
  assign n325 = ~n266 & n324;
  assign n326 = n177 & ~n325;
  assign n327 = ~n177 & n325;
  assign n328 = pi13 & ~n326;
  assign n329 = ~n327 & n328;
  assign n330 = n111 & ~n233;
  assign po1 = n329 | ~n330;
  assign n332 = ~pi02 & n30;
  assign n333 = n108 & n211;
  assign n334 = pi01 & ~pi05;
  assign n335 = ~n90 & ~n182;
  assign n336 = ~n334 & ~n335;
  assign n337 = ~pi06 & ~n336;
  assign n338 = pi09 & n337;
  assign n339 = pi06 & n44;
  assign n340 = n336 & n339;
  assign n341 = ~n338 & ~n340;
  assign n342 = pi02 & ~n341;
  assign n343 = pi06 & n336;
  assign n344 = ~n336 & ~n339;
  assign n345 = ~pi02 & pi09;
  assign n346 = ~n343 & n345;
  assign n347 = ~n344 & n346;
  assign n348 = ~n333 & ~n347;
  assign n349 = ~n342 & n348;
  assign n350 = n117 & ~n349;
  assign n351 = pi02 & pi06;
  assign n352 = ~n201 & n351;
  assign n353 = ~pi02 & ~pi06;
  assign n354 = n38 & ~n353;
  assign n355 = ~pi06 & ~n51;
  assign n356 = ~n354 & ~n355;
  assign n357 = ~n352 & n356;
  assign n358 = ~n350 & n357;
  assign n359 = ~n332 & n358;
  assign n360 = ~n94 & n359;
  assign n361 = ~pi06 & n96;
  assign n362 = ~n360 & ~n361;
  assign n363 = ~pi09 & ~n362;
  assign n364 = ~n78 & n351;
  assign n365 = n83 & n353;
  assign n366 = ~n364 & ~n365;
  assign n367 = pi09 & ~n366;
  assign n368 = pi02 & pi11;
  assign n369 = ~pi06 & ~pi09;
  assign n370 = n25 & ~n369;
  assign n371 = n368 & ~n370;
  assign n372 = pi02 & n112;
  assign n373 = ~n75 & ~n372;
  assign n374 = ~n359 & ~n373;
  assign n375 = n71 & ~n359;
  assign n376 = pi09 & n79;
  assign n377 = ~pi02 & n40;
  assign n378 = n73 & n377;
  assign n379 = ~n376 & ~n378;
  assign n380 = ~n375 & n379;
  assign n381 = pi06 & ~n380;
  assign n382 = ~n367 & ~n371;
  assign n383 = ~n374 & n382;
  assign n384 = ~n363 & n383;
  assign n385 = ~n381 & n384;
  assign n386 = ~pi13 & ~n385;
  assign n387 = pi06 & n73;
  assign n388 = n133 & n351;
  assign n389 = ~pi02 & n359;
  assign n390 = n118 & ~n389;
  assign n391 = n24 & n359;
  assign n392 = pi09 & n359;
  assign n393 = pi02 & pi08;
  assign n394 = ~n369 & n393;
  assign n395 = ~n392 & n394;
  assign n396 = ~n391 & ~n395;
  assign n397 = n120 & ~n396;
  assign n398 = ~n390 & ~n397;
  assign n399 = n135 & n398;
  assign n400 = ~n388 & ~n399;
  assign n401 = n359 & n400;
  assign n402 = ~n359 & ~n400;
  assign n403 = ~n401 & ~n402;
  assign n404 = ~n209 & ~n251;
  assign n405 = ~n250 & ~n404;
  assign n406 = ~n403 & n405;
  assign n407 = n403 & ~n405;
  assign n408 = n41 & ~n406;
  assign n409 = ~n407 & n408;
  assign n410 = pi01 & ~n258;
  assign n411 = ~n260 & ~n410;
  assign n412 = n398 & n411;
  assign n413 = ~n398 & ~n411;
  assign n414 = ~n412 & ~n413;
  assign n415 = pi02 & ~pi08;
  assign n416 = ~n414 & n415;
  assign n417 = ~n387 & ~n416;
  assign n418 = ~n409 & n417;
  assign n419 = n57 & ~n418;
  assign n420 = n59 & n414;
  assign n421 = pi01 & ~n277;
  assign n422 = ~n276 & ~n421;
  assign n423 = n305 & ~n359;
  assign n424 = n422 & n423;
  assign n425 = ~n420 & ~n424;
  assign n426 = ~pi02 & ~n425;
  assign n427 = ~pi02 & n305;
  assign n428 = ~n422 & n427;
  assign n429 = n281 & n422;
  assign n430 = ~n284 & ~n429;
  assign n431 = pi02 & ~n430;
  assign n432 = ~n296 & n359;
  assign n433 = ~n428 & n432;
  assign n434 = ~n431 & n433;
  assign n435 = ~n295 & ~n302;
  assign n436 = ~pi10 & n301;
  assign n437 = n281 & ~n422;
  assign n438 = ~n284 & ~n437;
  assign n439 = pi02 & ~n438;
  assign n440 = ~n359 & ~n436;
  assign n441 = ~n435 & n440;
  assign n442 = ~n439 & n441;
  assign n443 = ~n434 & ~n442;
  assign n444 = ~n61 & ~n188;
  assign n445 = ~n185 & ~n444;
  assign n446 = ~n351 & ~n353;
  assign n447 = ~n445 & ~n446;
  assign n448 = pi11 & n353;
  assign n449 = ~n351 & ~n448;
  assign n450 = n445 & n449;
  assign n451 = n162 & ~n447;
  assign n452 = ~n450 & n451;
  assign n453 = n267 & n398;
  assign n454 = ~n267 & ~n398;
  assign n455 = ~pi11 & ~n453;
  assign n456 = ~n454 & n455;
  assign n457 = pi02 & ~n289;
  assign n458 = ~pi02 & n289;
  assign n459 = pi11 & ~n458;
  assign n460 = ~n457 & n459;
  assign n461 = n112 & ~n460;
  assign n462 = ~n456 & n461;
  assign n463 = ~n247 & ~n312;
  assign n464 = ~n311 & ~n463;
  assign n465 = n400 & n464;
  assign n466 = ~n400 & ~n464;
  assign n467 = ~n465 & ~n466;
  assign n468 = n398 & ~n467;
  assign n469 = ~n398 & n467;
  assign n470 = n138 & ~n468;
  assign n471 = ~n469 & n470;
  assign n472 = ~n443 & ~n452;
  assign n473 = ~n462 & n472;
  assign n474 = ~n426 & n473;
  assign n475 = ~n471 & n474;
  assign n476 = ~n419 & n475;
  assign n477 = pi13 & n326;
  assign n478 = ~n476 & n477;
  assign n479 = ~n326 & n476;
  assign n480 = pi13 & ~n479;
  assign n481 = ~n478 & n480;
  assign n482 = n111 & ~n386;
  assign po2 = n481 | ~n482;
  assign n484 = pi07 & n71;
  assign n485 = ~n75 & ~n484;
  assign n486 = ~pi03 & ~pi07;
  assign n487 = n38 & ~n486;
  assign n488 = pi02 & ~n343;
  assign n489 = ~n337 & ~n488;
  assign n490 = pi07 & pi09;
  assign n491 = n120 & n490;
  assign n492 = ~n489 & n491;
  assign n493 = ~n29 & ~n492;
  assign n494 = ~pi03 & ~n493;
  assign n495 = n108 & n368;
  assign n496 = pi09 & n486;
  assign n497 = n489 & n496;
  assign n498 = ~n495 & ~n497;
  assign n499 = pi13 & ~n498;
  assign po5 = pi03 & pi07;
  assign n501 = n120 & n489;
  assign n502 = ~n199 & ~n501;
  assign n503 = po5 & ~n502;
  assign n504 = ~n494 & ~n499;
  assign n505 = ~n503 & n504;
  assign n506 = ~pi08 & ~n505;
  assign n507 = pi03 & n46;
  assign n508 = ~n489 & n507;
  assign n509 = n51 & ~n508;
  assign n510 = ~pi07 & ~n509;
  assign n511 = ~n55 & ~n199;
  assign n512 = pi13 & po5;
  assign n513 = ~n511 & n512;
  assign n514 = ~n487 & ~n513;
  assign n515 = ~n510 & n514;
  assign n516 = ~n506 & n515;
  assign n517 = ~n485 & ~n516;
  assign n518 = ~pi07 & n96;
  assign n519 = ~n94 & n516;
  assign n520 = ~pi09 & ~n518;
  assign n521 = ~n519 & n520;
  assign n522 = ~n78 & po5;
  assign n523 = pi03 & ~n516;
  assign n524 = n41 & n523;
  assign n525 = n83 & n486;
  assign n526 = pi09 & ~n522;
  assign n527 = ~n525 & n526;
  assign n528 = ~n524 & n527;
  assign n529 = ~n521 & ~n528;
  assign n530 = ~pi03 & n40;
  assign n531 = n73 & n530;
  assign n532 = ~n376 & ~n531;
  assign n533 = pi07 & ~n532;
  assign n534 = ~pi07 & ~pi09;
  assign n535 = n25 & ~n534;
  assign n536 = pi03 & pi11;
  assign n537 = ~n535 & n536;
  assign n538 = ~n533 & ~n537;
  assign n539 = ~n517 & n538;
  assign n540 = ~n529 & n539;
  assign n541 = ~pi13 & ~n540;
  assign n542 = n133 & po5;
  assign n543 = ~pi03 & n516;
  assign n544 = n118 & ~n543;
  assign n545 = n24 & n516;
  assign n546 = n48 & n523;
  assign n547 = n33 & po5;
  assign n548 = ~n545 & ~n547;
  assign n549 = ~n546 & n548;
  assign n550 = n120 & ~n549;
  assign n551 = ~n544 & ~n550;
  assign n552 = n135 & n551;
  assign n553 = ~n542 & ~n552;
  assign n554 = ~n401 & ~n405;
  assign n555 = ~n402 & ~n554;
  assign n556 = n516 & n555;
  assign n557 = ~n516 & ~n555;
  assign n558 = ~n556 & ~n557;
  assign n559 = n553 & ~n558;
  assign n560 = ~n553 & n558;
  assign n561 = pi08 & ~n559;
  assign n562 = ~n560 & n561;
  assign n563 = pi02 & ~n412;
  assign n564 = ~n413 & ~n563;
  assign n565 = n551 & n564;
  assign n566 = ~n551 & ~n564;
  assign n567 = ~pi03 & ~n566;
  assign n568 = ~pi08 & ~n565;
  assign n569 = n567 & n568;
  assign n570 = ~n562 & ~n569;
  assign n571 = n199 & ~n570;
  assign n572 = pi02 & ~n358;
  assign n573 = ~n389 & ~n422;
  assign n574 = ~n572 & ~n573;
  assign n575 = n516 & n574;
  assign n576 = ~n516 & ~n574;
  assign n577 = ~n575 & ~n576;
  assign n578 = n281 & ~n577;
  assign n579 = ~n284 & ~n578;
  assign n580 = pi03 & ~n579;
  assign n581 = n305 & n577;
  assign n582 = ~n351 & ~n445;
  assign n583 = ~n353 & ~n582;
  assign n584 = pi07 & n162;
  assign n585 = ~n583 & n584;
  assign n586 = ~n581 & ~n585;
  assign n587 = ~pi03 & ~n586;
  assign n588 = n112 & n459;
  assign n589 = pi07 & ~n583;
  assign n590 = ~pi07 & n583;
  assign n591 = n162 & ~n589;
  assign n592 = ~n590 & n591;
  assign n593 = ~n588 & ~n592;
  assign n594 = pi03 & ~n593;
  assign n595 = n296 & n359;
  assign n596 = n516 & n595;
  assign n597 = n295 & n359;
  assign n598 = ~n436 & n597;
  assign n599 = ~n302 & ~n516;
  assign n600 = ~n598 & n599;
  assign n601 = n453 & n551;
  assign n602 = ~n453 & ~n551;
  assign n603 = ~n601 & ~n602;
  assign n604 = n112 & ~n603;
  assign n605 = ~n565 & ~n566;
  assign n606 = pi03 & n24;
  assign n607 = ~n605 & n606;
  assign n608 = ~n584 & ~n604;
  assign n609 = ~n607 & n608;
  assign n610 = ~pi11 & ~n609;
  assign n611 = ~pi03 & n112;
  assign n612 = n458 & n611;
  assign n613 = ~n398 & ~n465;
  assign n614 = ~n466 & ~n613;
  assign n615 = n553 & n614;
  assign n616 = ~n553 & ~n614;
  assign n617 = ~n615 & ~n616;
  assign n618 = ~n551 & n617;
  assign n619 = n551 & ~n617;
  assign n620 = n270 & ~n618;
  assign n621 = ~n619 & n620;
  assign n622 = n162 & n486;
  assign n623 = n583 & n622;
  assign n624 = ~n612 & ~n623;
  assign n625 = ~n621 & n624;
  assign n626 = pi11 & ~n625;
  assign n627 = ~n594 & ~n596;
  assign n628 = ~n600 & n627;
  assign n629 = ~n580 & n628;
  assign n630 = ~n587 & n629;
  assign n631 = ~n610 & n630;
  assign n632 = ~n571 & n631;
  assign n633 = ~n626 & n632;
  assign n634 = n478 & ~n633;
  assign n635 = ~n478 & n633;
  assign n636 = pi13 & ~n634;
  assign n637 = ~n635 & n636;
  assign n638 = n111 & ~n541;
  assign po3 = n637 | ~n638;
  assign po4 = n486 | po5;
  assign n641 = n551 & ~n616;
  assign n642 = n270 & ~n615;
  assign n643 = ~n641 & n642;
  assign n644 = ~po5 & ~n583;
  assign n645 = n162 & ~n486;
  assign n646 = ~n644 & n645;
  assign n647 = ~n523 & n574;
  assign n648 = ~n280 & ~n543;
  assign n649 = ~n647 & n648;
  assign n650 = pi11 & ~n612;
  assign n651 = ~n646 & n650;
  assign n652 = ~n649 & n651;
  assign n653 = ~n643 & n652;
  assign n654 = pi10 & ~n601;
  assign n655 = n48 & ~n654;
  assign n656 = ~n553 & ~n556;
  assign n657 = pi08 & ~n557;
  assign n658 = ~n656 & n657;
  assign n659 = ~n565 & ~n567;
  assign n660 = ~pi08 & ~n659;
  assign n661 = n108 & ~n658;
  assign n662 = ~n660 & n661;
  assign n663 = ~pi11 & ~n655;
  assign n664 = ~n662 & n663;
  assign n665 = ~n653 & ~n664;
  assign n666 = ~n73 & ~n83;
  assign n667 = pi09 & ~n666;
  assign n668 = n597 & n667;
  assign n669 = n516 & n668;
  assign n670 = ~n665 & ~n669;
  assign n671 = ~n634 & n670;
  assign po6 = pi13 & ~n671;
  assign n673 = ~n63 & ~n189;
  assign n674 = ~n446 & po4;
  assign po7 = n673 & n674;
endmodule
