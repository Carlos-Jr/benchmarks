module alu4_cl ( 
    pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8, pi9,
    po0, po1, po2, po3, po4, po5  );
  input  pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8, pi9;
  output po0, po1, po2, po3, po4, po5;
  wire n17, n18, n19, n20, n21, n22, n23,
    n24, n25, n26, n27, n28, n29, n30, n31,
    n32, n33, n34, n35, n36, n37, n38, n39,
    n40, n41, n42, n43, n44, n45, n46, n47,
    n48, n49, n50, n51, n52, n53, n54, n55,
    n56, n57, n58, n59, n60, n61, n62, n63,
    n64, n65, n66, n67, n68, n69, n70, n71,
    n72, n73, n74, n75, n76, n77, n78, n79,
    n80, n81, n82, n83, n84, n85, n86, n87,
    n88, n89, n90, n91, n92, n93, n94, n95,
    n96, n97, n98, n99, n100, n101, n102,
    n103, n104, n105, n106, n107, n108, n109,
    n110, n111, n112, n113, n114, n115, n116,
    n117, n118, n119, n120, n121, n122, n123,
    n124, n125, n126, n127, n128, n129, n130,
    n131, n132, n133, n134, n135, n136, n137,
    n138, n139, n140, n141, n142, n143, n144,
    n145, n146, n147, n148, n149, n150, n151,
    n152, n153, n154, n155, n156, n157, n158,
    n159, n160, n161, n162, n163, n164, n165,
    n166, n167, n168, n169, n170, n171, n172,
    n173, n174, n175, n176, n177, n178, n179,
    n180, n181, n182, n183, n184, n185, n186,
    n187, n188, n189, n190, n191, n192, n193,
    n194, n195, n196, n197, n198, n199, n200,
    n201, n202, n203, n204, n205, n206, n207,
    n208, n209, n210, n211, n212, n213, n214,
    n215, n216, n217, n218, n219, n220, n221,
    n222, n223, n224, n225, n226, n227, n228,
    n229, n230, n231, n232, n233, n234, n235,
    n237, n238, n239, n240, n241, n242, n243,
    n244, n245, n246, n247, n248, n249, n250,
    n251, n252, n253, n254, n255, n256, n257,
    n258, n259, n260, n261, n262, n263, n264,
    n265, n266, n267, n268, n269, n270, n271,
    n272, n273, n274, n275, n276, n277, n278,
    n279, n280, n281, n282, n283, n284, n285,
    n286, n287, n288, n289, n290, n291, n292,
    n293, n294, n295, n296, n297, n298, n299,
    n300, n301, n302, n303, n304, n305, n306,
    n307, n308, n309, n310, n311, n312, n313,
    n314, n315, n316, n317, n318, n319, n320,
    n321, n322, n323, n324, n325, n326, n327,
    n328, n329, n330, n331, n332, n333, n334,
    n335, n336, n337, n338, n339, n340, n341,
    n342, n343, n344, n345, n346, n347, n348,
    n349, n350, n351, n352, n353, n354, n355,
    n356, n357, n358, n359, n360, n361, n362,
    n363, n364, n365, n366, n367, n368, n369,
    n370, n371, n372, n373, n374, n375, n376,
    n377, n378, n379, n380, n381, n382, n383,
    n384, n385, n386, n387, n388, n389, n390,
    n391, n392, n393, n394, n395, n396, n397,
    n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n408, n409, n410, n411,
    n412, n413, n414, n415, n416, n417, n418,
    n419, n420, n421, n422, n423, n424, n425,
    n426, n427, n428, n429, n430, n431, n432,
    n433, n434, n435, n436, n437, n438, n439,
    n440, n441, n442, n443, n444, n445, n446,
    n447, n448, n449, n450, n451, n452, n453,
    n454, n455, n456, n457, n458, n459, n460,
    n461, n462, n463, n464, n465, n466, n467,
    n468, n469, n470, n471, n472, n473, n474,
    n475, n476, n477, n478, n479, n480, n481,
    n482, n483, n484, n485, n486, n487, n488,
    n489, n490, n491, n492, n493, n494, n495,
    n496, n497, n498, n499, n500, n501, n502,
    n503, n504, n505, n506, n507, n508, n509,
    n510, n511, n512, n513, n514, n515, n516,
    n517, n518, n519, n520, n521, n522, n523,
    n524, n525, n526, n527, n528, n529, n530,
    n531, n532, n533, n534, n535, n536, n537,
    n538, n539, n540, n541, n542, n543, n544,
    n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n557, n558,
    n559, n560, n561, n562, n563, n564, n565,
    n566, n567, n568, n569, n570, n571, n572,
    n573, n574, n575, n576, n577, n578, n579,
    n580, n581, n582, n583, n584, n585, n586,
    n587, n588, n589, n590, n591, n592, n593,
    n594, n595, n596, n597, n598, n599, n600,
    n601, n602, n603, n604, n605, n606, n607,
    n608, n609, n610, n611, n612, n613, n614,
    n615, n616, n617, n618, n619, n620, n621,
    n622, n623, n624, n625, n626, n627, n628,
    n629, n630, n631, n633, n634, n635, n636,
    n637, n638, n639, n640, n641, n642, n643,
    n644, n645, n646, n647, n648, n649, n650,
    n651, n652, n653, n654, n655, n656, n657,
    n658, n659, n660, n661, n662, n663, n664,
    n665, n666, n667, n668, n669, n670, n671,
    n672, n673, n674, n675, n676, n677, n678,
    n679, n680, n681, n682, n683, n684, n685,
    n686, n687, n688, n689, n690, n691, n692,
    n693, n694, n695, n696, n697, n698, n699,
    n700, n701, n702, n703, n704, n705, n706,
    n707, n708, n710, n711, n712, n713, n714,
    n715, n716, n717, n718, n719, n720, n721,
    n722, n723, n724, n725, n726, n727, n728,
    n729, n730, n731, n732, n733, n734, n735,
    n736, n737, n738, n739, n740, n741, n742,
    n743, n744, n745, n746, n747, n748, n749,
    n750, n751, n752, n753, n754, n755, n756,
    n757, n758, n759, n760, n761, n762, n763,
    n764, n765, n766, n767, n768, n769, n770,
    n771, n772, n774, n775, n776, n777, n778,
    n779, n780, n781, n782, n783, n784, n785,
    n786, n787, n788, n789, n790, n791, n792,
    n793, n794, n795, n796, n797, n798, n799,
    n800, n801, n802, n803, n804, n805, n806,
    n807, n808, n809, n810, n811, n812, n813,
    n814, n815, n816, n817;
  assign n17 = pi4 & pi5;
  assign n18 = ~pi6 & n17;
  assign n19 = ~pi7 & n18;
  assign n20 = pi6 & ~pi7;
  assign n21 = pi5 & pi9;
  assign n22 = ~pi4 & n21;
  assign n23 = ~n20 & n21;
  assign n24 = ~pi4 & n23;
  assign n25 = ~pi4 & ~n20;
  assign n26 = n21 & n25;
  assign n27 = ~n20 & n22;
  assign n28 = n17 & n20;
  assign n29 = pi4 & ~pi9;
  assign n30 = ~pi5 & pi6;
  assign n31 = pi7 & n30;
  assign n32 = pi7 & n29;
  assign n33 = n30 & n32;
  assign n34 = n29 & n31;
  assign n35 = ~n28 & ~n711;
  assign n36 = ~n710 & ~n711;
  assign n37 = ~n28 & n36;
  assign n38 = ~n710 & ~n28;
  assign n39 = ~n711 & n38;
  assign n40 = ~n710 & n35;
  assign n41 = ~pi2 & ~n712;
  assign n42 = ~pi6 & pi7;
  assign n43 = pi9 & n42;
  assign n44 = ~pi4 & n20;
  assign n45 = ~n43 & ~n44;
  assign n46 = ~pi4 & ~pi5;
  assign n47 = ~n17 & ~n46;
  assign n48 = pi0 & pi2;
  assign n49 = ~n47 & n48;
  assign n50 = pi7 & ~n47;
  assign n51 = ~pi6 & n50;
  assign n52 = pi9 & n51;
  assign n53 = n43 & ~n47;
  assign n54 = ~pi7 & n30;
  assign n55 = ~pi5 & n20;
  assign n56 = ~pi4 & n714;
  assign n57 = n20 & n46;
  assign n58 = ~n713 & ~n715;
  assign n59 = n48 & ~n58;
  assign n60 = ~n45 & n49;
  assign n61 = pi6 & pi9;
  assign n62 = ~pi6 & ~pi9;
  assign n63 = ~pi7 & ~pi9;
  assign n64 = ~pi6 & n63;
  assign n65 = ~pi7 & n62;
  assign n66 = ~n61 & ~n717;
  assign n67 = pi4 & ~pi5;
  assign n68 = ~pi0 & ~pi2;
  assign n69 = n67 & ~n68;
  assign n70 = ~n66 & n67;
  assign n71 = ~n68 & n70;
  assign n72 = ~n66 & n69;
  assign n73 = ~n716 & ~n718;
  assign n74 = ~n41 & n73;
  assign n75 = pi5 & pi7;
  assign n76 = ~pi6 & ~n75;
  assign n77 = ~pi9 & n76;
  assign n78 = n62 & ~n75;
  assign n79 = ~pi0 & n719;
  assign n80 = ~pi0 & pi2;
  assign n81 = pi0 & ~pi2;
  assign n82 = ~n80 & ~n81;
  assign n83 = ~n48 & ~n68;
  assign n84 = ~pi0 & ~n20;
  assign n85 = n21 & ~n84;
  assign n86 = n21 & ~n720;
  assign n87 = ~n84 & n86;
  assign n88 = n20 & n80;
  assign n89 = ~n81 & ~n88;
  assign n90 = n21 & ~n89;
  assign n91 = ~n720 & n85;
  assign n92 = ~n79 & ~n721;
  assign n93 = ~pi4 & ~n92;
  assign n94 = ~n41 & ~n718;
  assign n95 = ~n93 & n94;
  assign n96 = ~n716 & n95;
  assign n97 = n73 & ~n93;
  assign n98 = ~n41 & n97;
  assign n99 = n74 & ~n93;
  assign n100 = n17 & n722;
  assign n101 = n17 & n74;
  assign n102 = ~pi6 & n723;
  assign n103 = ~pi6 & ~n46;
  assign n104 = ~pi0 & ~n103;
  assign n105 = ~n722 & n104;
  assign n106 = ~n102 & ~n105;
  assign n107 = pi7 & ~n106;
  assign n108 = ~pi4 & pi5;
  assign n109 = ~pi6 & ~n722;
  assign n110 = pi6 & n722;
  assign n111 = pi6 & ~n722;
  assign n112 = ~pi6 & n722;
  assign n113 = ~n111 & ~n112;
  assign n114 = ~n109 & ~n110;
  assign n115 = n108 & n724;
  assign n116 = ~pi0 & n722;
  assign n117 = ~pi4 & pi7;
  assign n118 = pi7 & n22;
  assign n119 = pi7 & n108;
  assign n120 = pi5 & n117;
  assign n121 = pi9 & n726;
  assign n122 = n21 & n117;
  assign n123 = ~n116 & n725;
  assign n124 = pi9 & n20;
  assign n125 = pi0 & ~n722;
  assign n126 = n17 & n125;
  assign n127 = n48 & n67;
  assign n128 = n46 & n722;
  assign n129 = ~n127 & ~n128;
  assign n130 = ~n126 & n129;
  assign n131 = n124 & ~n130;
  assign n132 = ~n123 & ~n131;
  assign n133 = pi4 & ~pi7;
  assign n134 = pi4 & n714;
  assign n135 = n30 & n133;
  assign n136 = pi9 & n727;
  assign n137 = n67 & n124;
  assign n138 = n132 & n728;
  assign n139 = n42 & n48;
  assign n140 = ~pi6 & n725;
  assign n141 = n48 & n140;
  assign n142 = ~pi6 & n48;
  assign n143 = n725 & n142;
  assign n144 = n22 & n139;
  assign n145 = ~n138 & ~n729;
  assign n146 = pi4 & n30;
  assign n147 = n67 & n111;
  assign n148 = ~n722 & n146;
  assign n149 = n30 & ~n722;
  assign n150 = pi4 & n145;
  assign n151 = n149 & n150;
  assign n152 = n145 & n730;
  assign n153 = ~n115 & ~n731;
  assign n154 = ~pi7 & ~n153;
  assign n155 = pi0 & ~pi4;
  assign n156 = ~pi7 & n132;
  assign n157 = ~pi7 & ~n131;
  assign n158 = n132 & n155;
  assign n159 = ~pi7 & n158;
  assign n160 = ~pi7 & n155;
  assign n161 = n132 & n160;
  assign n162 = n155 & n732;
  assign n163 = pi4 & ~pi6;
  assign n164 = pi4 & ~n720;
  assign n165 = ~pi6 & n164;
  assign n166 = ~n720 & n163;
  assign n167 = ~n733 & ~n734;
  assign n168 = ~pi5 & ~n167;
  assign n169 = pi6 & n17;
  assign n170 = ~pi0 & pi7;
  assign n171 = ~n732 & ~n170;
  assign n172 = n169 & ~n171;
  assign n173 = pi0 & ~n17;
  assign n174 = ~n20 & ~n42;
  assign n175 = pi0 & ~n20;
  assign n176 = ~n17 & ~n42;
  assign n177 = n175 & n176;
  assign n178 = n173 & n174;
  assign n179 = pi0 & pi6;
  assign n180 = pi7 & n179;
  assign n181 = n722 & n179;
  assign n182 = pi7 & n181;
  assign n183 = n722 & n180;
  assign n184 = pi0 & ~pi6;
  assign n185 = pi0 & ~pi7;
  assign n186 = ~pi6 & n185;
  assign n187 = ~pi7 & n184;
  assign n188 = ~n736 & ~n737;
  assign n189 = ~n17 & ~n188;
  assign n190 = ~n111 & n735;
  assign n191 = ~n172 & ~n738;
  assign n192 = ~n168 & n191;
  assign n193 = ~n154 & n192;
  assign n194 = ~pi5 & ~pi6;
  assign n195 = ~pi6 & n155;
  assign n196 = ~pi5 & n195;
  assign n197 = pi0 & n46;
  assign n198 = ~pi6 & n197;
  assign n199 = n155 & n194;
  assign n200 = ~n138 & ~n739;
  assign n201 = n722 & ~n200;
  assign n202 = ~pi0 & n714;
  assign n203 = ~pi6 & n75;
  assign n204 = n145 & n203;
  assign n205 = ~n202 & ~n204;
  assign n206 = ~pi4 & ~n132;
  assign n207 = ~pi0 & ~pi4;
  assign n208 = ~pi7 & n207;
  assign n209 = ~pi0 & ~pi7;
  assign n210 = ~pi4 & n30;
  assign n211 = n209 & n210;
  assign n212 = n714 & n207;
  assign n213 = n30 & n208;
  assign n214 = ~pi6 & n726;
  assign n215 = n42 & n108;
  assign n216 = n108 & n145;
  assign n217 = n42 & n216;
  assign n218 = n145 & n741;
  assign n219 = ~n740 & ~n742;
  assign n220 = ~n132 & ~n219;
  assign n221 = ~n205 & n206;
  assign n222 = ~n201 & ~n743;
  assign n223 = n192 & ~n743;
  assign n224 = ~n154 & ~n201;
  assign n225 = n223 & n224;
  assign n226 = n193 & n222;
  assign n227 = ~n154 & ~n168;
  assign n228 = ~n201 & n227;
  assign n229 = ~n107 & n228;
  assign n230 = ~n743 & n229;
  assign n231 = ~n172 & n230;
  assign n232 = ~n738 & n231;
  assign n233 = ~n107 & n744;
  assign n234 = pi9 & ~n745;
  assign n235 = ~pi8 & n234;
  assign po3 = pi1 & pi3;
  assign n237 = n80 & po3;
  assign n238 = ~pi1 & pi3;
  assign n239 = pi5 & ~n80;
  assign n240 = pi5 & n238;
  assign n241 = ~n80 & n240;
  assign n242 = n238 & n239;
  assign n243 = ~n237 & ~n746;
  assign n244 = n20 & ~n243;
  assign n245 = ~pi1 & ~pi3;
  assign n246 = n80 & ~n245;
  assign n247 = pi1 & ~pi3;
  assign n248 = ~n80 & ~n247;
  assign n249 = pi5 & ~n248;
  assign n250 = n80 & n245;
  assign n251 = ~n80 & n247;
  assign n252 = ~n250 & ~n251;
  assign n253 = pi5 & ~n252;
  assign n254 = ~n246 & n249;
  assign n255 = ~n244 & ~n747;
  assign n256 = pi9 & ~n255;
  assign n257 = ~pi1 & n719;
  assign n258 = ~n256 & ~n257;
  assign n259 = ~pi4 & ~n258;
  assign n260 = ~pi5 & n61;
  assign n261 = ~pi4 & pi9;
  assign n262 = ~pi5 & n179;
  assign n263 = n261 & n262;
  assign n264 = n61 & n197;
  assign n265 = pi0 & n61;
  assign n266 = n46 & n265;
  assign n267 = pi9 & n46;
  assign n268 = n179 & n267;
  assign n269 = n155 & n260;
  assign n270 = ~pi6 & po3;
  assign n271 = pi4 & n21;
  assign n272 = ~n267 & ~n271;
  assign n273 = pi9 & ~n47;
  assign n274 = n270 & ~n749;
  assign n275 = ~n748 & ~n274;
  assign n276 = pi7 & ~n275;
  assign n277 = ~pi3 & ~n712;
  assign n278 = ~n29 & po3;
  assign n279 = ~pi5 & po3;
  assign n280 = n20 & n279;
  assign n281 = ~n29 & n280;
  assign n282 = n714 & n278;
  assign n283 = n67 & ~n245;
  assign n284 = ~n66 & n283;
  assign n285 = ~n750 & ~n284;
  assign n286 = ~n277 & n285;
  assign n287 = ~n276 & n285;
  assign n288 = ~n277 & n287;
  assign n289 = ~n276 & n286;
  assign n290 = ~n277 & ~n284;
  assign n291 = ~n259 & n290;
  assign n292 = ~n276 & n291;
  assign n293 = ~n750 & n292;
  assign n294 = ~n259 & n751;
  assign n295 = n722 & n752;
  assign n296 = n17 & n295;
  assign n297 = ~pi1 & n752;
  assign n298 = n725 & ~n297;
  assign n299 = pi1 & ~n752;
  assign n300 = n17 & n299;
  assign n301 = n46 & n752;
  assign n302 = n67 & po3;
  assign n303 = ~n301 & ~n302;
  assign n304 = ~n300 & n303;
  assign n305 = n124 & ~n304;
  assign n306 = ~n298 & ~n305;
  assign n307 = n728 & n306;
  assign n308 = n140 & po3;
  assign n309 = n725 & n270;
  assign n310 = ~n307 & ~n753;
  assign n311 = n729 & ~n310;
  assign n312 = ~n729 & n310;
  assign n313 = n729 & n310;
  assign n314 = ~n729 & ~n310;
  assign n315 = ~n313 & ~n314;
  assign n316 = ~n311 & ~n312;
  assign n317 = ~n306 & ~n754;
  assign n318 = n306 & n754;
  assign n319 = n108 & ~n318;
  assign n320 = ~n306 & n754;
  assign n321 = n306 & ~n754;
  assign n322 = ~n320 & ~n321;
  assign n323 = n108 & ~n322;
  assign n324 = ~n317 & n319;
  assign n325 = ~n296 & ~n755;
  assign n326 = ~pi6 & ~n325;
  assign n327 = ~pi4 & pi6;
  assign n328 = ~n30 & ~n46;
  assign n329 = ~n30 & ~n327;
  assign n330 = ~n46 & n329;
  assign n331 = ~n327 & n328;
  assign n332 = n125 & ~n752;
  assign n333 = ~n125 & n752;
  assign n334 = ~n332 & ~n333;
  assign n335 = ~n756 & n334;
  assign n336 = ~pi0 & pi6;
  assign n337 = ~pi0 & n169;
  assign n338 = ~pi0 & n17;
  assign n339 = pi6 & n338;
  assign n340 = n17 & n336;
  assign n341 = ~n335 & ~n757;
  assign n342 = ~pi1 & ~n341;
  assign n343 = pi1 & n179;
  assign n344 = n109 & ~n752;
  assign n345 = ~n343 & ~n344;
  assign n346 = n17 & ~n345;
  assign n347 = ~n342 & ~n346;
  assign n348 = ~n326 & ~n346;
  assign n349 = ~n342 & n348;
  assign n350 = ~n326 & n347;
  assign n351 = pi7 & ~n758;
  assign n352 = ~n722 & ~n145;
  assign n353 = n752 & ~n352;
  assign n354 = ~n752 & n352;
  assign n355 = ~n353 & ~n354;
  assign n356 = ~n310 & n355;
  assign n357 = n310 & ~n355;
  assign n358 = n67 & ~n357;
  assign n359 = ~n310 & n352;
  assign n360 = n310 & ~n354;
  assign n361 = n310 & ~n352;
  assign n362 = n310 & n352;
  assign n363 = ~n310 & ~n352;
  assign n364 = ~n362 & ~n363;
  assign n365 = ~n359 & ~n759;
  assign n366 = ~n752 & n760;
  assign n367 = n752 & ~n760;
  assign n368 = ~n366 & ~n367;
  assign n369 = n67 & ~n368;
  assign n370 = ~n356 & n358;
  assign n371 = pi0 & ~n132;
  assign n372 = n306 & ~n371;
  assign n373 = ~n306 & n371;
  assign n374 = ~n306 & ~n371;
  assign n375 = n306 & n371;
  assign n376 = ~n374 & ~n375;
  assign n377 = ~n372 & ~n373;
  assign n378 = ~pi1 & n46;
  assign n379 = ~n762 & n378;
  assign n380 = n17 & n132;
  assign n381 = n132 & n306;
  assign n382 = n17 & n381;
  assign n383 = n306 & n380;
  assign n384 = n17 & ~n132;
  assign n385 = ~n132 & ~n306;
  assign n386 = n17 & n385;
  assign n387 = ~n306 & n384;
  assign n388 = ~n763 & ~n764;
  assign n389 = ~n379 & n388;
  assign n390 = ~n761 & n389;
  assign n391 = pi6 & ~n390;
  assign n392 = pi1 & ~pi4;
  assign n393 = pi1 & n46;
  assign n394 = ~pi5 & n392;
  assign n395 = ~pi5 & n762;
  assign n396 = n392 & n395;
  assign n397 = n762 & n765;
  assign n398 = n108 & ~n752;
  assign n399 = pi1 & ~n17;
  assign n400 = ~n398 & ~n399;
  assign n401 = ~pi6 & ~n17;
  assign n402 = pi5 & ~n752;
  assign n403 = ~pi1 & ~n402;
  assign n404 = n401 & ~n403;
  assign n405 = ~pi6 & ~n400;
  assign n406 = pi6 & n295;
  assign n407 = ~n722 & ~n752;
  assign n408 = ~n406 & ~n407;
  assign n409 = n108 & ~n408;
  assign n410 = ~n767 & ~n409;
  assign n411 = n46 & n762;
  assign n412 = ~n401 & ~n411;
  assign n413 = pi1 & ~n412;
  assign n414 = ~n110 & n752;
  assign n415 = n110 & ~n752;
  assign n416 = n108 & ~n415;
  assign n417 = ~pi6 & ~n752;
  assign n418 = ~n407 & ~n417;
  assign n419 = ~n406 & n418;
  assign n420 = n108 & ~n419;
  assign n421 = ~n414 & n416;
  assign n422 = ~n413 & ~n768;
  assign n423 = ~n766 & n410;
  assign n424 = ~n391 & ~n766;
  assign n425 = ~n409 & n424;
  assign n426 = ~n767 & n425;
  assign n427 = ~n391 & n769;
  assign n428 = ~pi7 & ~n770;
  assign n429 = pi1 & pi7;
  assign n430 = pi1 & ~n756;
  assign n431 = pi7 & n430;
  assign n432 = ~n756 & n429;
  assign n433 = pi1 & ~pi6;
  assign n434 = n46 & n433;
  assign n435 = n194 & n392;
  assign n436 = ~n771 & ~n772;
  assign n437 = ~n334 & ~n436;
  assign n438 = ~pi5 & n163;
  assign n439 = pi7 & n245;
  assign n440 = ~po3 & ~n439;
  assign n441 = n48 & ~n440;
  assign n442 = pi3 & ~pi7;
  assign n443 = ~n238 & ~n247;
  assign n444 = ~po3 & ~n245;
  assign n445 = ~n48 & ~po2;
  assign n446 = ~n442 & ~n445;
  assign n447 = ~n441 & n446;
  assign n448 = n48 & n438;
  assign n449 = ~n440 & n448;
  assign n450 = n438 & ~n446;
  assign n451 = ~n449 & ~n450;
  assign n452 = n438 & ~n447;
  assign n453 = ~n437 & n774;
  assign n454 = ~n428 & n453;
  assign n455 = ~n351 & ~n428;
  assign n456 = ~n450 & n455;
  assign n457 = ~n437 & n456;
  assign n458 = ~n449 & n457;
  assign n459 = ~n351 & n454;
  assign n460 = pi9 & ~n775;
  assign n461 = n235 & n460;
  assign n462 = n235 & ~n775;
  assign n463 = ~n235 & n775;
  assign n464 = ~n776 & ~n463;
  assign n465 = ~n19 & ~n464;
  assign n466 = n235 & ~n460;
  assign n467 = ~n235 & n460;
  assign n468 = ~n19 & ~n467;
  assign n469 = ~n19 & ~n466;
  assign n470 = ~n467 & n469;
  assign n471 = ~n466 & n468;
  assign n472 = pi9 & ~n777;
  assign n473 = pi9 & ~n465;
  assign n474 = pi4 & pi6;
  assign n475 = pi4 & n299;
  assign n476 = pi6 & n475;
  assign n477 = n299 & n474;
  assign n478 = n20 & n245;
  assign n479 = ~pi4 & n478;
  assign n480 = n44 & n245;
  assign n481 = po3 & n327;
  assign n482 = pi5 & ~n481;
  assign n483 = ~n780 & n482;
  assign n484 = ~n779 & n483;
  assign n485 = pi6 & ~n752;
  assign n486 = n163 & n238;
  assign n487 = ~n247 & ~n327;
  assign n488 = ~n392 & n487;
  assign n489 = ~n486 & n488;
  assign n490 = ~n485 & n489;
  assign n491 = pi7 & ~n490;
  assign n492 = ~pi4 & ~pi6;
  assign n493 = ~pi4 & n417;
  assign n494 = ~n752 & n492;
  assign n495 = pi3 & pi6;
  assign n496 = n133 & ~n495;
  assign n497 = ~pi3 & pi6;
  assign n498 = ~pi6 & n752;
  assign n499 = ~n497 & ~n498;
  assign n500 = pi4 & ~n499;
  assign n501 = ~pi7 & n500;
  assign n502 = n133 & ~n499;
  assign n503 = ~n417 & n496;
  assign n504 = n752 & n327;
  assign n505 = ~pi5 & ~n504;
  assign n506 = ~n782 & n505;
  assign n507 = ~n781 & n506;
  assign n508 = ~n247 & ~n392;
  assign n509 = ~n486 & n508;
  assign n510 = ~n247 & ~n485;
  assign n511 = ~n392 & ~n486;
  assign n512 = n510 & n511;
  assign n513 = ~n485 & n509;
  assign n514 = pi7 & ~n783;
  assign n515 = ~pi5 & ~n781;
  assign n516 = ~pi7 & ~n752;
  assign n517 = n327 & ~n516;
  assign n518 = ~n782 & ~n517;
  assign n519 = n515 & n518;
  assign n520 = ~n514 & n519;
  assign n521 = ~n491 & n507;
  assign n522 = ~n484 & ~n784;
  assign n523 = pi3 & pi5;
  assign n524 = ~pi6 & ~n523;
  assign n525 = pi1 & pi6;
  assign n526 = pi5 & po3;
  assign n527 = ~n525 & ~n526;
  assign n528 = pi7 & ~n527;
  assign n529 = n429 & ~n524;
  assign n530 = ~n75 & ~n417;
  assign n531 = ~pi4 & ~n530;
  assign n532 = ~n726 & ~n781;
  assign n533 = pi3 & n786;
  assign n534 = pi6 & n429;
  assign n535 = pi1 & n75;
  assign n536 = ~n786 & ~n535;
  assign n537 = pi3 & ~n536;
  assign n538 = ~n534 & ~n537;
  assign n539 = ~n785 & ~n533;
  assign n540 = ~n781 & ~n517;
  assign n541 = ~n782 & n540;
  assign n542 = ~n781 & ~n514;
  assign n543 = ~n517 & n542;
  assign n544 = ~n782 & n543;
  assign n545 = ~n514 & n541;
  assign n546 = ~pi5 & ~n788;
  assign n547 = ~n780 & ~n481;
  assign n548 = ~n779 & n547;
  assign n549 = pi5 & ~n548;
  assign n550 = ~n533 & ~n549;
  assign n551 = ~n785 & n550;
  assign n552 = n787 & ~n549;
  assign n553 = ~n546 & n789;
  assign n554 = ~n522 & n787;
  assign n555 = ~pi9 & ~n790;
  assign n556 = ~n778 & ~n555;
  assign n557 = pi5 & n327;
  assign n558 = ~pi7 & n557;
  assign n559 = pi5 & ~pi7;
  assign n560 = n327 & n559;
  assign n561 = n20 & n108;
  assign n562 = ~n18 & ~n791;
  assign n563 = n295 & ~n562;
  assign n564 = ~pi6 & n108;
  assign n565 = ~n312 & n564;
  assign n566 = ~n306 & n565;
  assign n567 = ~n306 & ~n312;
  assign n568 = ~n125 & ~n299;
  assign n569 = ~n297 & ~n756;
  assign n570 = n125 & ~n297;
  assign n571 = ~n299 & ~n570;
  assign n572 = ~n756 & ~n571;
  assign n573 = ~n568 & n569;
  assign n574 = ~pi0 & ~pi1;
  assign n575 = n169 & n574;
  assign n576 = ~pi1 & n757;
  assign n577 = n48 & ~n245;
  assign n578 = ~n245 & n448;
  assign n579 = n438 & n577;
  assign n580 = po3 & n438;
  assign n581 = n67 & n270;
  assign n582 = pi7 & ~n796;
  assign n583 = ~n795 & n582;
  assign n584 = ~n794 & n583;
  assign n585 = ~n793 & n584;
  assign n586 = ~n792 & n585;
  assign n587 = ~n310 & ~n353;
  assign n588 = pi4 & ~n354;
  assign n589 = ~n587 & n588;
  assign n590 = pi1 & ~n372;
  assign n591 = ~pi4 & ~n373;
  assign n592 = ~n590 & n591;
  assign n593 = n30 & ~n592;
  assign n594 = pi4 & ~n353;
  assign n595 = ~n759 & n594;
  assign n596 = ~n354 & ~n587;
  assign n597 = ~pi1 & ~n371;
  assign n598 = ~pi4 & ~n306;
  assign n599 = ~pi4 & ~n597;
  assign n600 = ~n306 & n599;
  assign n601 = ~n597 & n598;
  assign n602 = n371 & n392;
  assign n603 = ~pi1 & ~n373;
  assign n604 = ~pi4 & ~n372;
  assign n605 = ~n603 & n604;
  assign n606 = ~n798 & ~n602;
  assign n607 = ~n797 & ~n602;
  assign n608 = ~n798 & n607;
  assign n609 = ~n797 & ~n799;
  assign n610 = n30 & ~n800;
  assign n611 = ~n589 & n593;
  assign n612 = ~pi7 & ~n18;
  assign n613 = ~n763 & n612;
  assign n614 = ~n801 & n613;
  assign n615 = ~n586 & ~n614;
  assign n616 = ~n763 & ~n801;
  assign n617 = ~pi7 & ~n616;
  assign n618 = ~n794 & ~n796;
  assign n619 = ~n795 & ~n796;
  assign n620 = ~n794 & n619;
  assign n621 = ~n795 & n618;
  assign n622 = ~n793 & n802;
  assign n623 = ~n792 & n622;
  assign n624 = pi7 & ~n623;
  assign n625 = ~n563 & ~n624;
  assign n626 = ~n617 & n625;
  assign n627 = ~n563 & ~n615;
  assign n628 = ~n776 & ~n624;
  assign n629 = ~n617 & n628;
  assign n630 = ~n563 & n629;
  assign n631 = ~n776 & n803;
  assign po4 = pi9 & ~n804;
  assign n633 = pi8 & ~n234;
  assign n634 = ~n235 & ~n633;
  assign n635 = pi8 & n234;
  assign n636 = ~pi8 & ~n234;
  assign n637 = ~n19 & ~n636;
  assign n638 = ~n635 & n637;
  assign n639 = ~n19 & ~n635;
  assign n640 = ~n636 & n639;
  assign n641 = ~n19 & ~n634;
  assign n642 = pi9 & ~n805;
  assign n643 = ~pi0 & ~n163;
  assign n644 = pi2 & ~n163;
  assign n645 = ~n720 & ~n644;
  assign n646 = ~n720 & ~n643;
  assign n647 = ~n155 & ~n327;
  assign n648 = n80 & n163;
  assign n649 = ~n81 & ~n155;
  assign n650 = ~n81 & n647;
  assign n651 = ~n327 & n649;
  assign n652 = ~n648 & n807;
  assign n653 = ~n806 & n647;
  assign n654 = ~n111 & ~n648;
  assign n655 = n807 & n654;
  assign n656 = ~n111 & n808;
  assign n657 = ~pi5 & ~n809;
  assign n658 = pi5 & n48;
  assign n659 = ~n179 & ~n658;
  assign n660 = ~n657 & n659;
  assign n661 = pi7 & ~n660;
  assign n662 = ~pi4 & n724;
  assign n663 = pi2 & pi6;
  assign n664 = n133 & ~n663;
  assign n665 = ~pi2 & pi6;
  assign n666 = ~n112 & ~n665;
  assign n667 = pi4 & ~n666;
  assign n668 = ~pi7 & n667;
  assign n669 = n133 & ~n666;
  assign n670 = ~n109 & n664;
  assign n671 = ~n662 & ~n810;
  assign n672 = ~pi5 & ~n671;
  assign n673 = pi6 & n125;
  assign n674 = pi4 & n673;
  assign n675 = n125 & n474;
  assign n676 = n48 & n327;
  assign n677 = n20 & n68;
  assign n678 = ~pi4 & n677;
  assign n679 = n44 & n68;
  assign n680 = ~n676 & ~n812;
  assign n681 = ~n811 & ~n676;
  assign n682 = ~n812 & n681;
  assign n683 = ~n811 & n680;
  assign n684 = pi5 & ~n813;
  assign n685 = ~n75 & ~n109;
  assign n686 = pi2 & ~pi4;
  assign n687 = ~pi4 & n109;
  assign n688 = ~n726 & ~n687;
  assign n689 = pi2 & ~n688;
  assign n690 = ~n685 & n686;
  assign n691 = ~n684 & ~n814;
  assign n692 = ~n672 & n691;
  assign n693 = pi7 & ~n809;
  assign n694 = ~n810 & ~n693;
  assign n695 = ~n662 & ~n693;
  assign n696 = ~n810 & n695;
  assign n697 = ~n662 & n694;
  assign n698 = ~pi5 & ~n815;
  assign n699 = pi7 & ~n659;
  assign n700 = ~n814 & ~n699;
  assign n701 = n691 & ~n699;
  assign n702 = ~n684 & ~n699;
  assign n703 = ~n814 & n702;
  assign n704 = ~n684 & n700;
  assign n705 = ~n698 & n816;
  assign n706 = ~n661 & n692;
  assign n707 = ~pi9 & ~n817;
  assign n708 = ~n642 & ~n707;
  assign po5 = n720 & po2;
  assign n710 = n27 | n24 | n26;
  assign n711 = n33 | n34;
  assign n712 = n40 | n37 | n39;
  assign n713 = n52 | n53;
  assign n714 = n54 | n55;
  assign n715 = n56 | n57;
  assign n716 = n59 | n60;
  assign n717 = n64 | n65;
  assign n718 = n71 | n72;
  assign n719 = n77 | n78;
  assign n720 = n82 | ~n83;
  assign n721 = n91 | n87 | n90;
  assign n722 = n99 | n96 | n98;
  assign n723 = n100 | n101;
  assign n724 = n113 | ~n114;
  assign n725 = n122 | n118 | n121;
  assign n726 = n119 | n120;
  assign n727 = n134 | n135;
  assign n728 = n136 | n137;
  assign n729 = n144 | n141 | n143;
  assign n730 = n147 | n148;
  assign n731 = n151 | n152;
  assign n732 = n156 | n157;
  assign n733 = n162 | n159 | n161;
  assign n734 = n165 | n166;
  assign n735 = n177 | n178;
  assign n736 = n182 | n183;
  assign n737 = n186 | n187;
  assign n738 = n189 | n190;
  assign n739 = n199 | n196 | n198;
  assign n740 = n213 | n211 | n212;
  assign n741 = n214 | n215;
  assign n742 = n217 | n218;
  assign n743 = n220 | n221;
  assign n744 = n225 | n226;
  assign n745 = n232 | n233;
  assign n746 = n241 | n242;
  assign n747 = n253 | n254;
  assign n748 = n266 | n263 | n264 | n268 | n269;
  assign n749 = n272 | ~n273;
  assign n750 = n281 | n282;
  assign n751 = n288 | n289;
  assign n752 = n293 | n294;
  assign n753 = n308 | n309;
  assign n754 = n315 | ~n316;
  assign n755 = n323 | n324;
  assign n756 = n330 | n331;
  assign n757 = n340 | n337 | n339;
  assign n758 = n349 | n350;
  assign n759 = n360 | n361;
  assign n760 = n364 | ~n365;
  assign n761 = n369 | n370;
  assign n762 = n376 | ~n377;
  assign n763 = n382 | n383;
  assign n764 = n386 | n387;
  assign n765 = n393 | n394;
  assign n766 = n396 | n397;
  assign n767 = n404 | n405;
  assign n768 = n420 | n421;
  assign n769 = n422 | n423;
  assign n770 = n426 | n427;
  assign n771 = n431 | n432;
  assign n772 = n434 | n435;
  assign po2 = n443 | ~n444;
  assign n774 = n451 | ~n452;
  assign n775 = n458 | n459;
  assign n776 = n461 | n462;
  assign n777 = n470 | n471;
  assign n778 = n472 | n473;
  assign n779 = n476 | n477;
  assign n780 = n479 | n480;
  assign n781 = n493 | n494;
  assign n782 = n503 | n501 | n502;
  assign n783 = n512 | n513;
  assign n784 = n520 | n521;
  assign n785 = n528 | n529;
  assign n786 = n531 | ~n532;
  assign n787 = n538 | n539;
  assign n788 = n544 | n545;
  assign n789 = n551 | n552;
  assign n790 = n553 | n554;
  assign n791 = n561 | n558 | n560;
  assign n792 = n566 | n567;
  assign n793 = n572 | n573;
  assign n794 = n575 | n576;
  assign n795 = n578 | n579;
  assign n796 = n580 | n581;
  assign n797 = n595 | ~n596;
  assign n798 = n600 | n601;
  assign n799 = n605 | ~n606;
  assign n800 = n608 | n609;
  assign n801 = n610 | n611;
  assign n802 = n620 | n621;
  assign n803 = n626 | n627;
  assign n804 = n630 | n631;
  assign n805 = n641 | n638 | n640;
  assign n806 = n645 | n646;
  assign n807 = n650 | n651;
  assign n808 = n652 | n653;
  assign n809 = n655 | n656;
  assign n810 = n670 | n668 | n669;
  assign n811 = n674 | n675;
  assign n812 = n678 | n679;
  assign n813 = n682 | n683;
  assign n814 = n689 | n690;
  assign n815 = n696 | n697;
  assign n816 = n704 | n701 | n703;
  assign n817 = n705 | n706;
  assign po0 = ~n708;
  assign po1 = ~n556;
endmodule
